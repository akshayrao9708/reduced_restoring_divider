module divider(R_0, D, Q, R_n1);
input [13:0] R_0;
input [6:0] D;
output [7:0] Q;
output [6:0] R_n1;
wire _0_;
wire _1_;
wire _2_;
wire _3_;
wire _4_;
wire _5_;
wire _6_;
wire _7_;
wire _8_;
wire _9_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire _30_;
wire _31_;
wire _32_;
wire _33_;
wire _34_;
wire _35_;
wire _36_;
wire _37_;
wire _38_;
wire _39_;
wire _40_;
wire _41_;
wire _42_;
wire _43_;
wire _44_;
wire _45_;
wire _46_;
wire _47_;
wire _48_;
wire _49_;
wire _50_;
wire _51_;
wire _52_;
wire _53_;
wire _54_;
wire _55_;
wire _56_;
wire _57_;
wire _58_;
wire _59_;
wire _60_;
wire _61_;
wire _62_;
wire _63_;
wire _64_;
wire _65_;
wire _66_;
wire _67_;
wire _68_;
wire _69_;
wire _70_;
wire _71_;
wire _72_;
wire _73_;
wire _74_;
wire _75_;
wire _76_;
wire _77_;
wire _78_;
wire _79_;
wire _80_;
wire _81_;
wire _82_;
wire _83_;
wire _84_;
wire _85_;
wire _86_;
wire _87_;
wire _88_;
wire _89_;
wire _90_;
wire _91_;
wire _92_;
wire _93_;
wire _94_;
wire _95_;
wire _96_;
wire _97_;
wire _98_;
wire _99_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
wire _255_;
wire _256_;
wire _257_;
wire _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire _267_;
wire _268_;
wire _269_;
wire _270_;
wire _271_;
wire _272_;
wire _273_;
wire _274_;
wire _275_;
wire _276_;
wire _277_;
wire _278_;
wire _279_;
wire _280_;
wire _281_;
wire _282_;
wire _283_;
wire _284_;
wire _285_;
wire _286_;
wire _287_;
wire _288_;
wire _289_;
wire _290_;
wire _291_;
wire _292_;
wire _293_;
wire _294_;
wire _295_;
wire _296_;
wire _297_;
wire _298_;
wire _299_;
wire _300_;
wire _301_;
wire _302_;
wire _303_;
wire _304_;
wire _305_;
wire _306_;
wire _307_;
wire _308_;
wire _309_;
wire _310_;
wire _311_;
wire _312_;
wire _313_;
wire _314_;
wire _315_;
wire _316_;
wire _317_;
wire _318_;
wire _319_;
wire _320_;
wire _321_;
wire _322_;
wire _323_;
wire _324_;
wire _325_;
wire _326_;
wire _327_;
wire _328_;
wire _329_;
wire _330_;
wire _331_;
wire _332_;
wire _333_;
wire _334_;
wire _335_;
wire _336_;
wire _337_;
wire _338_;
wire _339_;
wire _340_;
wire _341_;
wire _342_;
wire _343_;
wire _344_;
wire _345_;
wire _346_;
wire _347_;
wire _348_;
wire _349_;
wire _350_;
wire _351_;
wire _352_;
wire _353_;
wire _354_;
wire _355_;
wire _356_;
wire _357_;
wire _358_;
wire _359_;
wire _360_;
wire _361_;
wire _362_;
wire _363_;
wire _364_;
wire _365_;
wire _366_;
wire _367_;
wire _368_;
wire _369_;
wire _370_;
wire _371_;
wire _372_;
wire _373_;
wire _374_;
wire _375_;
wire _376_;
wire _377_;
wire _378_;
wire _379_;
wire _380_;
wire _381_;
wire _382_;
wire _383_;
wire _384_;
wire _385_;
wire _386_;
wire _387_;
wire _388_;
wire _389_;
wire _390_;
wire _391_;
wire _392_;
wire _393_;
wire _394_;
wire _395_;
wire _396_;
wire _397_;
wire _398_;
wire _399_;
wire _400_;
wire _401_;
wire _402_;
wire _403_;
wire _404_;
wire _405_;
wire _406_;
wire _407_;
wire _408_;
wire _409_;
wire _410_;
wire _411_;
wire _412_;
wire _413_;
wire _414_;
wire _415_;
wire _416_;
wire _417_;
wire _418_;
wire _419_;
wire _420_;
wire _421_;
wire _422_;
wire _423_;
wire _424_;
wire _425_;
wire _426_;
wire _427_;
wire _428_;
wire _429_;
wire _430_;
wire _431_;
wire _432_;
wire _433_;
wire _434_;
wire _435_;
wire _436_;
wire _437_;
wire _438_;
wire _439_;
wire _440_;
wire _441_;
wire _442_;
wire _443_;
wire _444_;
wire _445_;
wire _446_;
wire _447_;
wire _448_;
wire _449_;
wire _450_;
wire _451_;
wire _452_;
wire _453_;
wire _454_;
wire _455_;
wire _456_;
wire _457_;
wire _458_;
wire _459_;
wire _460_;
wire _461_;
wire _462_;
wire _463_;
wire _464_;
wire _465_;
wire _466_;
wire _467_;
wire _468_;
wire _469_;
wire _470_;
wire _471_;
wire _472_;
wire _473_;
wire _474_;
wire _475_;
wire _476_;
wire _477_;
wire _478_;
wire _479_;
wire _480_;
wire _481_;
wire _482_;
wire _483_;
wire _484_;
wire _485_;
wire _486_;
wire _487_;
wire _488_;
wire _489_;
wire _490_;
wire _491_;
wire _492_;
wire _493_;
wire _494_;
wire _495_;
wire _496_;
wire _497_;
wire _498_;
wire _499_;
wire _500_;
wire _501_;
wire _502_;
wire _503_;
wire _504_;
wire _505_;
wire _506_;
wire _507_;
wire _508_;
wire _509_;
wire _510_;
wire _511_;
wire _512_;
wire _513_;
wire _514_;
wire _515_;
wire _516_;
wire _517_;
wire _518_;
wire _519_;
wire _520_;
wire _521_;
wire _522_;
wire _523_;
wire _524_;
wire _525_;
wire _526_;
wire _527_;
wire _528_;
wire _529_;
wire _530_;
wire _531_;
wire _532_;
wire _533_;
wire _534_;
wire _535_;
wire _536_;
wire _537_;
wire _538_;
wire _539_;
wire _540_;
wire _541_;
wire _542_;
wire _543_;
wire _544_;
wire _545_;
wire _546_;
wire _547_;
wire _548_;
wire _549_;
wire _550_;
wire _551_;
wire _552_;
wire _553_;
wire _554_;
wire _555_;
wire _556_;
wire _557_;
wire _558_;
wire _559_;
wire _560_;
wire _561_;
wire _562_;
wire _563_;
wire _564_;
wire _565_;
wire _566_;
wire _567_;
wire _568_;
wire _569_;
wire _570_;
wire _571_;
wire _572_;
wire _573_;
wire _574_;
wire _575_;
wire _576_;
wire _577_;
wire _578_;
wire _579_;
wire _580_;
wire _581_;
wire _582_;
wire _583_;
wire _584_;
wire _585_;
wire _586_;
wire _587_;
wire _588_;
wire _589_;
wire _590_;
wire _591_;
wire _592_;
wire _593_;
wire _594_;
wire _595_;
wire _596_;
wire _597_;
wire _598_;
wire _599_;
wire _600_;
wire _601_;
wire _602_;
wire _603_;
wire _604_;
wire _605_;
wire _606_;
wire _607_;
wire _608_;
wire _609_;
wire _610_;
wire _611_;
wire _612_;
wire _613_;
wire _614_;
wire _615_;
wire _616_;
wire _617_;
wire _618_;
wire _619_;
wire _620_;
wire _621_;
wire _622_;
wire _623_;
wire _624_;
wire _625_;
wire _626_;
wire _627_;
wire _628_;
wire _629_;
wire _630_;
wire _631_;
wire _632_;
wire _633_;
wire _634_;
wire _635_;
wire _636_;
wire _637_;
wire _638_;
wire _639_;
wire _640_;
wire _641_;
wire _642_;
wire _643_;
wire _644_;
wire _645_;
wire _646_;
wire _647_;
wire _648_;
wire _649_;
wire _650_;
wire _651_;
wire _652_;
wire _653_;
wire _654_;
wire _655_;
wire _656_;
wire _657_;
wire _658_;
wire _659_;
wire _660_;
wire _661_;
wire _662_;
wire _663_;
wire _664_;
wire _665_;
wire _666_;
wire _667_;
wire _668_;
wire _669_;
wire _670_;
wire _671_;
wire _672_;
wire _673_;
wire _674_;
wire _675_;
wire _676_;
wire _677_;
wire _678_;
wire _679_;
wire _680_;
wire _681_;
wire _682_;
wire _683_;
wire _684_;
wire _685_;
wire _686_;
wire _687_;
wire _688_;
wire _689_;
wire _690_;
wire _691_;
wire _692_;
wire _693_;
wire _694_;
wire _695_;
wire _696_;
wire _697_;
wire _698_;
wire _699_;
wire _700_;
wire _701_;
wire _702_;
wire _703_;
wire _704_;
wire _705_;
wire _706_;
wire _707_;
wire _708_;
wire _709_;
wire _710_;
wire _711_;
wire _712_;
wire _713_;
wire _714_;
wire _715_;
wire _716_;
wire _717_;
wire _718_;
wire _719_;
wire _720_;
wire _721_;
wire _722_;
wire _723_;
wire _724_;
wire _725_;
wire _726_;
wire _727_;
wire _728_;
wire _729_;
wire _730_;
wire _731_;
wire _732_;
wire _733_;
wire _734_;
wire _735_;
wire _736_;
wire _737_;
wire _738_;
wire _739_;
wire _740_;
wire _741_;
wire _742_;
wire _743_;
wire _744_;
wire _745_;
wire _746_;
wire _747_;
wire _748_;
wire _749_;
wire _750_;
wire _751_;
wire _752_;
wire _753_;
wire _754_;
wire _755_;
wire _756_;
wire _757_;
wire _758_;
wire _759_;
wire _760_;
wire _761_;
wire _762_;
wire _763_;
wire _764_;
wire _765_;
wire _766_;
wire _767_;
wire _768_;
wire _769_;
wire _770_;
wire _771_;
wire _772_;
wire _773_;
wire _774_;
wire _775_;
wire _776_;
wire _777_;
wire _778_;
wire _779_;
wire _780_;
wire _781_;
wire _782_;
wire _783_;
wire _784_;
wire _785_;
wire _786_;
wire _787_;
wire _788_;
wire _789_;
wire _790_;
wire _791_;
wire _792_;
wire _793_;
wire _794_;
wire _795_;
wire _796_;
wire _797_;
wire _798_;
wire _799_;
wire _800_;
wire _801_;
wire _802_;
wire _803_;
wire _804_;
wire _805_;
wire _806_;
wire _807_;
wire _808_;
wire _809_;
wire _810_;
wire _811_;
wire _812_;
wire _813_;
wire _814_;
wire _815_;
wire _816_;
wire _817_;
wire _818_;
wire _819_;
wire _820_;
wire _821_;
wire _822_;
wire _823_;
wire _824_;
wire _825_;
wire _826_;
wire _827_;
wire _828_;
wire _829_;
wire _830_;
wire _831_;
wire _832_;
wire _833_;
wire _834_;
wire _835_;
wire _836_;
wire _837_;
wire _838_;
wire _839_;
wire _840_;
wire _841_;
wire _842_;
wire _843_;
wire _844_;
wire _845_;
wire _846_;
wire _847_;
wire _848_;
wire _849_;
wire _850_;
wire _851_;
wire _852_;
wire _853_;
wire _854_;
wire _855_;
wire _856_;
wire _857_;
wire _858_;
wire _859_;
wire _860_;
wire _861_;
wire _862_;
wire _863_;
wire _864_;
wire _865_;
wire _866_;
wire _867_;
wire _868_;
wire _869_;
wire _870_;
wire _871_;
wire _872_;
wire _873_;
wire _874_;
wire _875_;
wire _876_;
wire _877_;
wire _878_;
wire _879_;
wire _880_;
wire _881_;
wire _882_;
wire _883_;
wire _884_;
wire _885_;
wire _886_;
wire _887_;
wire _888_;
wire _889_;
wire _890_;
wire _891_;
wire _892_;
wire _893_;
wire _894_;
wire _895_;
wire _896_;
wire _897_;
wire _898_;
wire _899_;
wire _900_;
wire _901_;
wire _902_;
wire _903_;
wire _904_;
wire _905_;
wire _906_;
wire _907_;
wire _908_;
wire _909_;
wire _910_;
wire _911_;
wire _912_;
wire _913_;
wire _914_;
wire _915_;
wire _916_;
wire _917_;
wire _918_;
wire _919_;
wire _920_;
wire _921_;
wire _922_;
wire _923_;
wire _924_;
wire _925_;
wire _926_;
wire _927_;
wire _928_;
wire _929_;
wire _930_;
wire _931_;
wire _932_;
wire _933_;
wire _934_;
wire _935_;
wire _936_;
wire _937_;
wire _938_;
wire _939_;
wire _940_;
wire _941_;
wire _942_;
wire _943_;
wire _944_;
wire _945_;
wire _946_;
wire _947_;
wire _948_;
wire _949_;
wire _950_;
wire _951_;
wire _952_;
wire _953_;
wire _954_;
wire _955_;
wire _956_;
wire _957_;
wire _958_;
wire _959_;
wire _960_;
wire _961_;
wire _962_;
wire _963_;
wire _964_;
wire _965_;
wire _966_;
wire _967_;
wire _968_;
wire _969_;
wire _970_;
wire _971_;
wire _972_;
wire _973_;
wire _974_;
wire _975_;
wire _976_;
wire _977_;
wire _978_;
wire _979_;
wire _980_;
wire _981_;
wire _982_;
wire _983_;
wire _984_;
wire _985_;
wire _986_;
wire _987_;
wire _988_;
wire _989_;
wire _990_;
wire _991_;
wire _992_;
wire _993_;
wire _994_;
wire _995_;
wire _996_;
wire _997_;
wire _998_;
wire _999_;
wire _1000_;
wire _1001_;
wire _1002_;
wire _1003_;
wire _1004_;
wire _1005_;
wire _1006_;
wire _1007_;
wire _1008_;
wire _1009_;
wire _1010_;
wire _1011_;
wire _1012_;
wire _1013_;
wire _1014_;
wire _1015_;
wire _1016_;
wire _1017_;
wire _1018_;
wire _1019_;
wire _1020_;
wire _1021_;
wire _1022_;
wire _1023_;
wire _1024_;
wire _1025_;
wire _1026_;
wire _1027_;
wire _1028_;
wire _1029_;
wire _1030_;
wire _1031_;
wire _1032_;
wire _1033_;
wire _1034_;
wire _1035_;
wire _1036_;
wire _1037_;
wire _1038_;
wire _1039_;
wire _1040_;
wire _1041_;
wire _1042_;
wire _1043_;
wire _1044_;
wire _1045_;
wire _1046_;
wire _1047_;
wire _1048_;
wire _1049_;
wire _1050_;
wire _1051_;
wire _1052_;
wire _1053_;
wire _1054_;
wire _1055_;
wire _1056_;
wire _1057_;
wire _1058_;
wire _1059_;
wire _1060_;
wire _1061_;
wire _1062_;
wire _1063_;
wire _1064_;
wire _1065_;
wire _1066_;
wire _1067_;
wire _1068_;
wire _1069_;
wire _1070_;
wire _1071_;
wire _1072_;
wire _1073_;
wire _1074_;
wire _1075_;
wire _1076_;
wire _1077_;
wire _1078_;
wire _1079_;
wire _1080_;
wire _1081_;
wire _1082_;
wire _1083_;
wire _1084_;
wire _1085_;
wire _1086_;
wire _1087_;
wire _1088_;
wire _1089_;
wire _1090_;
wire _1091_;
wire _1092_;
wire _1093_;
wire _1094_;
wire _1095_;
wire _1096_;
wire _1097_;
wire _1098_;
wire _1099_;
wire _1100_;
wire _1101_;
wire _1102_;
wire _1103_;
wire _1104_;
wire _1105_;
wire _1106_;
wire _1107_;
wire _1108_;
wire _1109_;
wire _1110_;
wire _1111_;
wire _1112_;
wire _1113_;
wire _1114_;
wire _1115_;
wire _1116_;
wire _1117_;
wire _1118_;
wire _1119_;
wire _1120_;
wire _1121_;
wire _1122_;
wire _1123_;
wire _1124_;
wire _1125_;
wire _1126_;
wire _1127_;
wire _1128_;
wire _1129_;
wire _1130_;
wire _1131_;
wire _1132_;
wire _1133_;
wire _1134_;
wire _1135_;
wire _1136_;
wire _1137_;
wire _1138_;
wire _1139_;
wire _1140_;
wire _1141_;
wire _1142_;
wire _1143_;
wire _1144_;
wire _1145_;
wire _1146_;
wire _1147_;
wire _1148_;
wire _1149_;
wire _1150_;
wire _1151_;
wire _1152_;
wire _1153_;
wire _1154_;
wire _1155_;
wire _1156_;
wire _1157_;
wire _1158_;
wire _1159_;
wire _1160_;
wire _1161_;
wire _1162_;
wire _1163_;
wire _1164_;
wire _1165_;
wire _1166_;
wire _1167_;
wire _1168_;
wire _1169_;
wire _1170_;
wire _1171_;
wire _1172_;
wire _1173_;
wire _1174_;
wire _1175_;
wire _1176_;
wire _1177_;
wire _1178_;
wire _1179_;
wire _1180_;
wire _1181_;
wire _1182_;
wire _1183_;
wire _1184_;
wire _1185_;
wire _1186_;
wire _1187_;
wire _1188_;
wire _1189_;
wire _1190_;
wire _1191_;
wire _1192_;
wire _1193_;
wire _1194_;
wire _1195_;
wire _1196_;
wire _1197_;
wire _1198_;
wire _1199_;
wire _1200_;
wire _1201_;
wire _1202_;
wire _1203_;
wire _1204_;
wire _1205_;
wire _1206_;
wire _1207_;
wire _1208_;
wire _1209_;
wire _1210_;
wire _1211_;
wire _1212_;
wire _1213_;
wire _1214_;
wire _1215_;
wire _1216_;
wire _1217_;
wire _1218_;
wire _1219_;
wire _1220_;
wire _1221_;
wire _1222_;
wire _1223_;
wire _1224_;
wire _1225_;
wire _1226_;
wire _1227_;
wire _1228_;
wire _1229_;
wire _1230_;
wire _1231_;
wire _1232_;
wire _1233_;
wire _1234_;
wire _1235_;
wire _1236_;
wire _1237_;
wire _1238_;
wire _1239_;
wire _1240_;
wire _1241_;
wire _1242_;
wire _1243_;
wire _1244_;
wire _1245_;
wire _1246_;
wire _1247_;
wire _1248_;
wire _1249_;
wire _1250_;
wire _1251_;
wire _1252_;
wire _1253_;
wire _1254_;
wire _1255_;
wire _1256_;
wire _1257_;
wire _1258_;
wire _1259_;
wire _1260_;
wire _1261_;
wire _1262_;
wire _1263_;
wire _1264_;
wire _1265_;
wire _1266_;
wire _1267_;
wire _1268_;
wire _1269_;
wire _1270_;
wire _1271_;
wire _1272_;
wire _1273_;
wire _1274_;
wire _1275_;
wire _1276_;
wire _1277_;
wire _1278_;
wire _1279_;
wire _1280_;
wire _1281_;
wire _1282_;
wire _1283_;
wire _1284_;
wire _1285_;
wire _1286_;
wire _1287_;
wire _1288_;
wire _1289_;
wire _1290_;
wire _1291_;
wire _1292_;
wire _1293_;
wire _1294_;
wire _1295_;
wire _1296_;
wire _1297_;
wire _1298_;
wire _1299_;
wire _1300_;
wire _1301_;
wire _1302_;
wire _1303_;
wire _1304_;
wire _1305_;
wire _1306_;
wire _1307_;
wire _1308_;
wire _1309_;
wire _1310_;
wire _1311_;
wire _1312_;
wire _1313_;
wire _1314_;
wire _1315_;
wire _1316_;
wire _1317_;
wire _1318_;
wire _1319_;
wire _1320_;
wire _1321_;
wire _1322_;
wire _1323_;
wire _1324_;
wire _1325_;
wire _1326_;
wire _1327_;
wire _1328_;
wire _1329_;
wire _1330_;
wire _1331_;
wire _1332_;
wire _1333_;
wire _1334_;
wire _1335_;
wire _1336_;
wire _1337_;
wire _1338_;
wire _1339_;
wire _1340_;
wire _1341_;
wire _1342_;
wire _1343_;
wire _1344_;
wire _1345_;
wire _1346_;
wire _1347_;
wire _1348_;
wire _1349_;
wire _1350_;
wire _1351_;
wire _1352_;
wire _1353_;
wire _1354_;
wire _1355_;
wire _1356_;
wire _1357_;
wire _1358_;
wire _1359_;
wire _1360_;
wire _1361_;
wire _1362_;
wire _1363_;
wire _1364_;
wire _1365_;
wire _1366_;
wire _1367_;
wire _1368_;
wire _1369_;
wire _1370_;
wire _1371_;
wire _1372_;
wire _1373_;
wire _1374_;
wire _1375_;
wire _1376_;
wire _1377_;
wire _1378_;
wire _1379_;
wire _1380_;
wire _1381_;
wire _1382_;
wire _1383_;
wire _1384_;
wire _1385_;
wire _1386_;
wire _1387_;
wire _1388_;
wire _1389_;
wire _1390_;
wire _1391_;
wire _1392_;
wire _1393_;
wire _1394_;
wire _1395_;
wire _1396_;
wire _1397_;
wire _1398_;
wire _1399_;
wire _1400_;
wire _1401_;
wire _1402_;
wire _1403_;
wire _1404_;
wire _1405_;
wire _1406_;
wire _1407_;
wire _1408_;
wire _1409_;
wire _1410_;
wire _1411_;
wire _1412_;
wire _1413_;
wire _1414_;
wire _1415_;
wire _1416_;
wire _1417_;
wire _1418_;
wire _1419_;
wire _1420_;
wire _1421_;
wire _1422_;
wire _1423_;
wire _1424_;
wire _1425_;
wire _1426_;
wire _1427_;
wire _1428_;
wire _1429_;
wire _1430_;
wire _1431_;
wire _1432_;
wire _1433_;
wire _1434_;
wire _1435_;
wire _1436_;
wire _1437_;
wire _1438_;
wire _1439_;
wire _1440_;
wire _1441_;
wire _1442_;
wire _1443_;
wire _1444_;
wire _1445_;
wire _1446_;
wire _1447_;
wire _1448_;
wire _1449_;
wire _1450_;
wire _1451_;
wire _1452_;
wire _1453_;
wire _1454_;
wire _1455_;
wire _1456_;
wire _1457_;
wire _1458_;
wire _1459_;
wire _1460_;
wire _1461_;
wire _1462_;
wire _1463_;
wire _1464_;
wire _1465_;
wire _1466_;
wire _1467_;
wire _1468_;
wire _1469_;
wire _1470_;
wire _1471_;
wire _1472_;
wire _1473_;
wire zeroWire;
wire oneWire;
assign zeroWire = 1'b0 /*1730*/;
assign oneWire = 1'b1 /*1730*/;
assign _13_ = ~D[0] /*1680*/;
assign _10_ = R_0[7] & _13_ /*1676*/;
assign _11_ = R_0[7] ^ _13_ /*1679*/;
assign _12_ = oneWire & _11_ /*1677*/;
assign _0_ = oneWire ^ _11_ /*1678*/;
assign _9_ = _10_ | _12_ /*1675*/;
assign _18_ = ~D[1] /*1674*/;
assign _15_ = R_0[8] & _18_ /*1670*/;
assign _16_ = R_0[8] ^ _18_ /*1673*/;
assign _17_ = _9_ & _16_ /*1671*/;
assign _1_ = _9_ ^ _16_ /*1672*/;
assign _14_ = _15_ | _17_ /*1669*/;
assign _23_ = ~D[2] /*1668*/;
assign _20_ = R_0[9] & _23_ /*1664*/;
assign _21_ = R_0[9] ^ _23_ /*1667*/;
assign _22_ = _14_ & _21_ /*1665*/;
assign _2_ = _14_ ^ _21_ /*1666*/;
assign _19_ = _20_ | _22_ /*1663*/;
assign _28_ = ~D[3] /*1662*/;
assign _25_ = R_0[10] & _28_ /*1658*/;
assign _26_ = R_0[10] ^ _28_ /*1661*/;
assign _27_ = _19_ & _26_ /*1659*/;
assign _3_ = _19_ ^ _26_ /*1660*/;
assign _24_ = _25_ | _27_ /*1657*/;
assign _33_ = ~D[4] /*1656*/;
assign _30_ = R_0[11] & _33_ /*1652*/;
assign _31_ = R_0[11] ^ _33_ /*1655*/;
assign _32_ = _24_ & _31_ /*1653*/;
assign _4_ = _24_ ^ _31_ /*1654*/;
assign _29_ = _30_ | _32_ /*1651*/;
assign _38_ = ~D[5] /*1650*/;
assign _35_ = R_0[12] & _38_ /*1646*/;
assign _36_ = R_0[12] ^ _38_ /*1649*/;
assign _37_ = _29_ & _36_ /*1647*/;
assign _5_ = _29_ ^ _36_ /*1648*/;
assign _34_ = _35_ | _37_ /*1645*/;
assign _43_ = ~D[6] /*1644*/;
assign _40_ = R_0[13] & _43_ /*1640*/;
assign _41_ = R_0[13] ^ _43_ /*1643*/;
assign _42_ = _34_ & _41_ /*1641*/;
assign _6_ = _34_ ^ _41_ /*1642*/;
assign _39_ = _40_ | _42_ /*1639*/;
assign _44_ = zeroWire & oneWire /*1634*/;
assign _45_ = zeroWire ^ oneWire /*1637*/;
assign _46_ = _39_ & _45_ /*1635*/;
assign _7_ = _39_ ^ _45_ /*1636*/;
assign Q[7] = _44_ | _46_ /*1633*/;
assign _59_ = ~Q[7] /*1585*/;
assign _58_ = _59_ & D[0] /*1584*/;
assign _61_ = _0_ & _58_ /*1579*/;
assign _62_ = _0_ ^ _58_ /*1582*/;
assign _63_ = zeroWire & _62_ /*1580*/;
assign _49_ = zeroWire ^ _62_ /*1581*/;
assign _60_ = _61_ | _63_ /*1578*/;
assign _65_ = ~Q[7] /*1577*/;
assign _64_ = _65_ & D[1] /*1576*/;
assign _67_ = _1_ & _64_ /*1571*/;
assign _68_ = _1_ ^ _64_ /*1574*/;
assign _69_ = _60_ & _68_ /*1572*/;
assign _50_ = _60_ ^ _68_ /*1573*/;
assign _66_ = _67_ | _69_ /*1570*/;
assign _71_ = ~Q[7] /*1569*/;
assign _70_ = _71_ & D[2] /*1568*/;
assign _73_ = _2_ & _70_ /*1563*/;
assign _74_ = _2_ ^ _70_ /*1566*/;
assign _75_ = _66_ & _74_ /*1564*/;
assign _51_ = _66_ ^ _74_ /*1565*/;
assign _72_ = _73_ | _75_ /*1562*/;
assign _77_ = ~Q[7] /*1561*/;
assign _76_ = _77_ & D[3] /*1560*/;
assign _79_ = _3_ & _76_ /*1555*/;
assign _80_ = _3_ ^ _76_ /*1558*/;
assign _81_ = _72_ & _80_ /*1556*/;
assign _52_ = _72_ ^ _80_ /*1557*/;
assign _78_ = _79_ | _81_ /*1554*/;
assign _83_ = ~Q[7] /*1553*/;
assign _82_ = _83_ & D[4] /*1552*/;
assign _85_ = _4_ & _82_ /*1547*/;
assign _86_ = _4_ ^ _82_ /*1550*/;
assign _87_ = _78_ & _86_ /*1548*/;
assign _53_ = _78_ ^ _86_ /*1549*/;
assign _84_ = _85_ | _87_ /*1546*/;
assign _89_ = ~Q[7] /*1545*/;
assign _88_ = _89_ & D[5] /*1544*/;
assign _91_ = _5_ & _88_ /*1539*/;
assign _92_ = _5_ ^ _88_ /*1542*/;
assign _93_ = _84_ & _92_ /*1540*/;
assign _54_ = _84_ ^ _92_ /*1541*/;
assign _90_ = _91_ | _93_ /*1538*/;
assign _95_ = ~Q[7] /*1537*/;
assign _94_ = _95_ & D[6] /*1536*/;
assign _97_ = _6_ & _94_ /*1531*/;
assign _98_ = _6_ ^ _94_ /*1534*/;
assign _99_ = _90_ & _98_ /*1532*/;
assign _55_ = _90_ ^ _98_ /*1533*/;
assign _96_ = _97_ | _99_ /*1530*/;
assign _101_ = ~Q[7] /*1529*/;
assign _100_ = _101_ & zeroWire /*1528*/;
assign _102_ = _7_ ^ _100_ /*1526*/;
assign _56_ = _102_ ^ _96_ /*1525*/;
assign _117_ = ~D[0] /*1495*/;
assign _114_ = R_0[6] & _117_ /*1491*/;
assign _115_ = R_0[6] ^ _117_ /*1494*/;
assign _116_ = oneWire & _115_ /*1492*/;
assign _105_ = oneWire ^ _115_ /*1493*/;
assign _113_ = _114_ | _116_ /*1490*/;
assign _122_ = ~D[1] /*1489*/;
assign _119_ = _49_ & _122_ /*1485*/;
assign _120_ = _49_ ^ _122_ /*1488*/;
assign _121_ = _113_ & _120_ /*1486*/;
assign _106_ = _113_ ^ _120_ /*1487*/;
assign _118_ = _119_ | _121_ /*1484*/;
assign _127_ = ~D[2] /*1483*/;
assign _124_ = _50_ & _127_ /*1479*/;
assign _125_ = _50_ ^ _127_ /*1482*/;
assign _126_ = _118_ & _125_ /*1480*/;
assign _107_ = _118_ ^ _125_ /*1481*/;
assign _123_ = _124_ | _126_ /*1478*/;
assign _132_ = ~D[3] /*1477*/;
assign _129_ = _51_ & _132_ /*1473*/;
assign _130_ = _51_ ^ _132_ /*1476*/;
assign _131_ = _123_ & _130_ /*1474*/;
assign _108_ = _123_ ^ _130_ /*1475*/;
assign _128_ = _129_ | _131_ /*1472*/;
assign _137_ = ~D[4] /*1471*/;
assign _134_ = _52_ & _137_ /*1467*/;
assign _135_ = _52_ ^ _137_ /*1470*/;
assign _136_ = _128_ & _135_ /*1468*/;
assign _109_ = _128_ ^ _135_ /*1469*/;
assign _133_ = _134_ | _136_ /*1466*/;
assign _142_ = ~D[5] /*1465*/;
assign _139_ = _53_ & _142_ /*1461*/;
assign _140_ = _53_ ^ _142_ /*1464*/;
assign _141_ = _133_ & _140_ /*1462*/;
assign _110_ = _133_ ^ _140_ /*1463*/;
assign _138_ = _139_ | _141_ /*1460*/;
assign _147_ = ~D[6] /*1459*/;
assign _144_ = _54_ & _147_ /*1455*/;
assign _145_ = _54_ ^ _147_ /*1458*/;
assign _146_ = _138_ & _145_ /*1456*/;
assign _111_ = _138_ ^ _145_ /*1457*/;
assign _143_ = _144_ | _146_ /*1454*/;
assign _148_ = _55_ & oneWire /*1449*/;
assign _149_ = _55_ ^ oneWire /*1452*/;
assign _150_ = _143_ & _149_ /*1450*/;
assign _112_ = _143_ ^ _149_ /*1451*/;
assign Q[6] = _148_ | _150_ /*1448*/;
assign _171_ = ~Q[6] /*1399*/;
assign _170_ = _171_ & D[0] /*1398*/;
assign _173_ = _105_ & _170_ /*1393*/;
assign _174_ = _105_ ^ _170_ /*1396*/;
assign _175_ = zeroWire & _174_ /*1394*/;
assign _161_ = zeroWire ^ _174_ /*1395*/;
assign _172_ = _173_ | _175_ /*1392*/;
assign _177_ = ~Q[6] /*1391*/;
assign _176_ = _177_ & D[1] /*1390*/;
assign _179_ = _106_ & _176_ /*1385*/;
assign _180_ = _106_ ^ _176_ /*1388*/;
assign _181_ = _172_ & _180_ /*1386*/;
assign _162_ = _172_ ^ _180_ /*1387*/;
assign _178_ = _179_ | _181_ /*1384*/;
assign _183_ = ~Q[6] /*1383*/;
assign _182_ = _183_ & D[2] /*1382*/;
assign _185_ = _107_ & _182_ /*1377*/;
assign _186_ = _107_ ^ _182_ /*1380*/;
assign _187_ = _178_ & _186_ /*1378*/;
assign _163_ = _178_ ^ _186_ /*1379*/;
assign _184_ = _185_ | _187_ /*1376*/;
assign _189_ = ~Q[6] /*1375*/;
assign _188_ = _189_ & D[3] /*1374*/;
assign _191_ = _108_ & _188_ /*1369*/;
assign _192_ = _108_ ^ _188_ /*1372*/;
assign _193_ = _184_ & _192_ /*1370*/;
assign _164_ = _184_ ^ _192_ /*1371*/;
assign _190_ = _191_ | _193_ /*1368*/;
assign _195_ = ~Q[6] /*1367*/;
assign _194_ = _195_ & D[4] /*1366*/;
assign _197_ = _109_ & _194_ /*1361*/;
assign _198_ = _109_ ^ _194_ /*1364*/;
assign _199_ = _190_ & _198_ /*1362*/;
assign _165_ = _190_ ^ _198_ /*1363*/;
assign _196_ = _197_ | _199_ /*1360*/;
assign _201_ = ~Q[6] /*1359*/;
assign _200_ = _201_ & D[5] /*1358*/;
assign _203_ = _110_ & _200_ /*1353*/;
assign _204_ = _110_ ^ _200_ /*1356*/;
assign _205_ = _196_ & _204_ /*1354*/;
assign _166_ = _196_ ^ _204_ /*1355*/;
assign _202_ = _203_ | _205_ /*1352*/;
assign _207_ = ~Q[6] /*1351*/;
assign _206_ = _207_ & D[6] /*1350*/;
assign _209_ = _111_ & _206_ /*1345*/;
assign _210_ = _111_ ^ _206_ /*1348*/;
assign _211_ = _202_ & _210_ /*1346*/;
assign _167_ = _202_ ^ _210_ /*1347*/;
assign _208_ = _209_ | _211_ /*1344*/;
assign _213_ = ~Q[6] /*1343*/;
assign _212_ = _213_ & zeroWire /*1342*/;
assign _214_ = _112_ ^ _212_ /*1340*/;
assign _168_ = _214_ ^ _208_ /*1339*/;
assign _229_ = ~D[0] /*1309*/;
assign _226_ = R_0[5] & _229_ /*1305*/;
assign _227_ = R_0[5] ^ _229_ /*1308*/;
assign _228_ = oneWire & _227_ /*1306*/;
assign _217_ = oneWire ^ _227_ /*1307*/;
assign _225_ = _226_ | _228_ /*1304*/;
assign _234_ = ~D[1] /*1303*/;
assign _231_ = _161_ & _234_ /*1299*/;
assign _232_ = _161_ ^ _234_ /*1302*/;
assign _233_ = _225_ & _232_ /*1300*/;
assign _218_ = _225_ ^ _232_ /*1301*/;
assign _230_ = _231_ | _233_ /*1298*/;
assign _239_ = ~D[2] /*1297*/;
assign _236_ = _162_ & _239_ /*1293*/;
assign _237_ = _162_ ^ _239_ /*1296*/;
assign _238_ = _230_ & _237_ /*1294*/;
assign _219_ = _230_ ^ _237_ /*1295*/;
assign _235_ = _236_ | _238_ /*1292*/;
assign _244_ = ~D[3] /*1291*/;
assign _241_ = _163_ & _244_ /*1287*/;
assign _242_ = _163_ ^ _244_ /*1290*/;
assign _243_ = _235_ & _242_ /*1288*/;
assign _220_ = _235_ ^ _242_ /*1289*/;
assign _240_ = _241_ | _243_ /*1286*/;
assign _249_ = ~D[4] /*1285*/;
assign _246_ = _164_ & _249_ /*1281*/;
assign _247_ = _164_ ^ _249_ /*1284*/;
assign _248_ = _240_ & _247_ /*1282*/;
assign _221_ = _240_ ^ _247_ /*1283*/;
assign _245_ = _246_ | _248_ /*1280*/;
assign _254_ = ~D[5] /*1279*/;
assign _251_ = _165_ & _254_ /*1275*/;
assign _252_ = _165_ ^ _254_ /*1278*/;
assign _253_ = _245_ & _252_ /*1276*/;
assign _222_ = _245_ ^ _252_ /*1277*/;
assign _250_ = _251_ | _253_ /*1274*/;
assign _259_ = ~D[6] /*1273*/;
assign _256_ = _166_ & _259_ /*1269*/;
assign _257_ = _166_ ^ _259_ /*1272*/;
assign _258_ = _250_ & _257_ /*1270*/;
assign _223_ = _250_ ^ _257_ /*1271*/;
assign _255_ = _256_ | _258_ /*1268*/;
assign _260_ = _167_ & oneWire /*1263*/;
assign _261_ = _167_ ^ oneWire /*1266*/;
assign _262_ = _255_ & _261_ /*1264*/;
assign _224_ = _255_ ^ _261_ /*1265*/;
assign Q[5] = _260_ | _262_ /*1262*/;
assign _283_ = ~Q[5] /*1213*/;
assign _282_ = _283_ & D[0] /*1212*/;
assign _285_ = _217_ & _282_ /*1207*/;
assign _286_ = _217_ ^ _282_ /*1210*/;
assign _287_ = zeroWire & _286_ /*1208*/;
assign _273_ = zeroWire ^ _286_ /*1209*/;
assign _284_ = _285_ | _287_ /*1206*/;
assign _289_ = ~Q[5] /*1205*/;
assign _288_ = _289_ & D[1] /*1204*/;
assign _291_ = _218_ & _288_ /*1199*/;
assign _292_ = _218_ ^ _288_ /*1202*/;
assign _293_ = _284_ & _292_ /*1200*/;
assign _274_ = _284_ ^ _292_ /*1201*/;
assign _290_ = _291_ | _293_ /*1198*/;
assign _295_ = ~Q[5] /*1197*/;
assign _294_ = _295_ & D[2] /*1196*/;
assign _297_ = _219_ & _294_ /*1191*/;
assign _298_ = _219_ ^ _294_ /*1194*/;
assign _299_ = _290_ & _298_ /*1192*/;
assign _275_ = _290_ ^ _298_ /*1193*/;
assign _296_ = _297_ | _299_ /*1190*/;
assign _301_ = ~Q[5] /*1189*/;
assign _300_ = _301_ & D[3] /*1188*/;
assign _303_ = _220_ & _300_ /*1183*/;
assign _304_ = _220_ ^ _300_ /*1186*/;
assign _305_ = _296_ & _304_ /*1184*/;
assign _276_ = _296_ ^ _304_ /*1185*/;
assign _302_ = _303_ | _305_ /*1182*/;
assign _307_ = ~Q[5] /*1181*/;
assign _306_ = _307_ & D[4] /*1180*/;
assign _309_ = _221_ & _306_ /*1175*/;
assign _310_ = _221_ ^ _306_ /*1178*/;
assign _311_ = _302_ & _310_ /*1176*/;
assign _277_ = _302_ ^ _310_ /*1177*/;
assign _308_ = _309_ | _311_ /*1174*/;
assign _313_ = ~Q[5] /*1173*/;
assign _312_ = _313_ & D[5] /*1172*/;
assign _315_ = _222_ & _312_ /*1167*/;
assign _316_ = _222_ ^ _312_ /*1170*/;
assign _317_ = _308_ & _316_ /*1168*/;
assign _278_ = _308_ ^ _316_ /*1169*/;
assign _314_ = _315_ | _317_ /*1166*/;
assign _319_ = ~Q[5] /*1165*/;
assign _318_ = _319_ & D[6] /*1164*/;
assign _321_ = _223_ & _318_ /*1159*/;
assign _322_ = _223_ ^ _318_ /*1162*/;
assign _323_ = _314_ & _322_ /*1160*/;
assign _279_ = _314_ ^ _322_ /*1161*/;
assign _320_ = _321_ | _323_ /*1158*/;
assign _325_ = ~Q[5] /*1157*/;
assign _324_ = _325_ & zeroWire /*1156*/;
assign _326_ = _224_ ^ _324_ /*1154*/;
assign _280_ = _326_ ^ _320_ /*1153*/;
assign _341_ = ~D[0] /*1123*/;
assign _338_ = R_0[4] & _341_ /*1119*/;
assign _339_ = R_0[4] ^ _341_ /*1122*/;
assign _340_ = oneWire & _339_ /*1120*/;
assign _329_ = oneWire ^ _339_ /*1121*/;
assign _337_ = _338_ | _340_ /*1118*/;
assign _346_ = ~D[1] /*1117*/;
assign _343_ = _273_ & _346_ /*1113*/;
assign _344_ = _273_ ^ _346_ /*1116*/;
assign _345_ = _337_ & _344_ /*1114*/;
assign _330_ = _337_ ^ _344_ /*1115*/;
assign _342_ = _343_ | _345_ /*1112*/;
assign _351_ = ~D[2] /*1111*/;
assign _348_ = _274_ & _351_ /*1107*/;
assign _349_ = _274_ ^ _351_ /*1110*/;
assign _350_ = _342_ & _349_ /*1108*/;
assign _331_ = _342_ ^ _349_ /*1109*/;
assign _347_ = _348_ | _350_ /*1106*/;
assign _356_ = ~D[3] /*1105*/;
assign _353_ = _275_ & _356_ /*1101*/;
assign _354_ = _275_ ^ _356_ /*1104*/;
assign _355_ = _347_ & _354_ /*1102*/;
assign _332_ = _347_ ^ _354_ /*1103*/;
assign _352_ = _353_ | _355_ /*1100*/;
assign _361_ = ~D[4] /*1099*/;
assign _358_ = _276_ & _361_ /*1095*/;
assign _359_ = _276_ ^ _361_ /*1098*/;
assign _360_ = _352_ & _359_ /*1096*/;
assign _333_ = _352_ ^ _359_ /*1097*/;
assign _357_ = _358_ | _360_ /*1094*/;
assign _366_ = ~D[5] /*1093*/;
assign _363_ = _277_ & _366_ /*1089*/;
assign _364_ = _277_ ^ _366_ /*1092*/;
assign _365_ = _357_ & _364_ /*1090*/;
assign _334_ = _357_ ^ _364_ /*1091*/;
assign _362_ = _363_ | _365_ /*1088*/;
assign _371_ = ~D[6] /*1087*/;
assign _368_ = _278_ & _371_ /*1083*/;
assign _369_ = _278_ ^ _371_ /*1086*/;
assign _370_ = _362_ & _369_ /*1084*/;
assign _335_ = _362_ ^ _369_ /*1085*/;
assign _367_ = _368_ | _370_ /*1082*/;
assign _372_ = _279_ & oneWire /*1077*/;
assign _373_ = _279_ ^ oneWire /*1080*/;
assign _374_ = _367_ & _373_ /*1078*/;
assign _336_ = _367_ ^ _373_ /*1079*/;
assign Q[4] = _372_ | _374_ /*1076*/;
assign _395_ = ~Q[4] /*1027*/;
assign _394_ = _395_ & D[0] /*1026*/;
assign _397_ = _329_ & _394_ /*1021*/;
assign _398_ = _329_ ^ _394_ /*1024*/;
assign _399_ = zeroWire & _398_ /*1022*/;
assign _385_ = zeroWire ^ _398_ /*1023*/;
assign _396_ = _397_ | _399_ /*1020*/;
assign _401_ = ~Q[4] /*1019*/;
assign _400_ = _401_ & D[1] /*1018*/;
assign _403_ = _330_ & _400_ /*1013*/;
assign _404_ = _330_ ^ _400_ /*1016*/;
assign _405_ = _396_ & _404_ /*1014*/;
assign _386_ = _396_ ^ _404_ /*1015*/;
assign _402_ = _403_ | _405_ /*1012*/;
assign _407_ = ~Q[4] /*1011*/;
assign _406_ = _407_ & D[2] /*1010*/;
assign _409_ = _331_ & _406_ /*1005*/;
assign _410_ = _331_ ^ _406_ /*1008*/;
assign _411_ = _402_ & _410_ /*1006*/;
assign _387_ = _402_ ^ _410_ /*1007*/;
assign _408_ = _409_ | _411_ /*1004*/;
assign _413_ = ~Q[4] /*1003*/;
assign _412_ = _413_ & D[3] /*1002*/;
assign _415_ = _332_ & _412_ /*997*/;
assign _416_ = _332_ ^ _412_ /*1000*/;
assign _417_ = _408_ & _416_ /*998*/;
assign _388_ = _408_ ^ _416_ /*999*/;
assign _414_ = _415_ | _417_ /*996*/;
assign _419_ = ~Q[4] /*995*/;
assign _418_ = _419_ & D[4] /*994*/;
assign _421_ = _333_ & _418_ /*989*/;
assign _422_ = _333_ ^ _418_ /*992*/;
assign _423_ = _414_ & _422_ /*990*/;
assign _389_ = _414_ ^ _422_ /*991*/;
assign _420_ = _421_ | _423_ /*988*/;
assign _425_ = ~Q[4] /*987*/;
assign _424_ = _425_ & D[5] /*986*/;
assign _427_ = _334_ & _424_ /*981*/;
assign _428_ = _334_ ^ _424_ /*984*/;
assign _429_ = _420_ & _428_ /*982*/;
assign _390_ = _420_ ^ _428_ /*983*/;
assign _426_ = _427_ | _429_ /*980*/;
assign _431_ = ~Q[4] /*979*/;
assign _430_ = _431_ & D[6] /*978*/;
assign _433_ = _335_ & _430_ /*973*/;
assign _434_ = _335_ ^ _430_ /*976*/;
assign _435_ = _426_ & _434_ /*974*/;
assign _391_ = _426_ ^ _434_ /*975*/;
assign _432_ = _433_ | _435_ /*972*/;
assign _437_ = ~Q[4] /*971*/;
assign _436_ = _437_ & zeroWire /*970*/;
assign _438_ = _336_ ^ _436_ /*968*/;
assign _392_ = _438_ ^ _432_ /*967*/;
assign _453_ = ~D[0] /*937*/;
assign _450_ = R_0[3] & _453_ /*933*/;
assign _451_ = R_0[3] ^ _453_ /*936*/;
assign _452_ = oneWire & _451_ /*934*/;
assign _441_ = oneWire ^ _451_ /*935*/;
assign _449_ = _450_ | _452_ /*932*/;
assign _458_ = ~D[1] /*931*/;
assign _455_ = _385_ & _458_ /*927*/;
assign _456_ = _385_ ^ _458_ /*930*/;
assign _457_ = _449_ & _456_ /*928*/;
assign _442_ = _449_ ^ _456_ /*929*/;
assign _454_ = _455_ | _457_ /*926*/;
assign _463_ = ~D[2] /*925*/;
assign _460_ = _386_ & _463_ /*921*/;
assign _461_ = _386_ ^ _463_ /*924*/;
assign _462_ = _454_ & _461_ /*922*/;
assign _443_ = _454_ ^ _461_ /*923*/;
assign _459_ = _460_ | _462_ /*920*/;
assign _468_ = ~D[3] /*919*/;
assign _465_ = _387_ & _468_ /*915*/;
assign _466_ = _387_ ^ _468_ /*918*/;
assign _467_ = _459_ & _466_ /*916*/;
assign _444_ = _459_ ^ _466_ /*917*/;
assign _464_ = _465_ | _467_ /*914*/;
assign _473_ = ~D[4] /*913*/;
assign _470_ = _388_ & _473_ /*909*/;
assign _471_ = _388_ ^ _473_ /*912*/;
assign _472_ = _464_ & _471_ /*910*/;
assign _445_ = _464_ ^ _471_ /*911*/;
assign _469_ = _470_ | _472_ /*908*/;
assign _478_ = ~D[5] /*907*/;
assign _475_ = _389_ & _478_ /*903*/;
assign _476_ = _389_ ^ _478_ /*906*/;
assign _477_ = _469_ & _476_ /*904*/;
assign _446_ = _469_ ^ _476_ /*905*/;
assign _474_ = _475_ | _477_ /*902*/;
assign _483_ = ~D[6] /*901*/;
assign _480_ = _390_ & _483_ /*897*/;
assign _481_ = _390_ ^ _483_ /*900*/;
assign _482_ = _474_ & _481_ /*898*/;
assign _447_ = _474_ ^ _481_ /*899*/;
assign _479_ = _480_ | _482_ /*896*/;
assign _484_ = _391_ & oneWire /*891*/;
assign _485_ = _391_ ^ oneWire /*894*/;
assign _486_ = _479_ & _485_ /*892*/;
assign _448_ = _479_ ^ _485_ /*893*/;
assign Q[3] = _484_ | _486_ /*890*/;
assign _507_ = ~Q[3] /*841*/;
assign _506_ = _507_ & D[0] /*840*/;
assign _509_ = _441_ & _506_ /*835*/;
assign _510_ = _441_ ^ _506_ /*838*/;
assign _511_ = zeroWire & _510_ /*836*/;
assign _497_ = zeroWire ^ _510_ /*837*/;
assign _508_ = _509_ | _511_ /*834*/;
assign _513_ = ~Q[3] /*833*/;
assign _512_ = _513_ & D[1] /*832*/;
assign _515_ = _442_ & _512_ /*827*/;
assign _516_ = _442_ ^ _512_ /*830*/;
assign _517_ = _508_ & _516_ /*828*/;
assign _498_ = _508_ ^ _516_ /*829*/;
assign _514_ = _515_ | _517_ /*826*/;
assign _519_ = ~Q[3] /*825*/;
assign _518_ = _519_ & D[2] /*824*/;
assign _521_ = _443_ & _518_ /*819*/;
assign _522_ = _443_ ^ _518_ /*822*/;
assign _523_ = _514_ & _522_ /*820*/;
assign _499_ = _514_ ^ _522_ /*821*/;
assign _520_ = _521_ | _523_ /*818*/;
assign _525_ = ~Q[3] /*817*/;
assign _524_ = _525_ & D[3] /*816*/;
assign _527_ = _444_ & _524_ /*811*/;
assign _528_ = _444_ ^ _524_ /*814*/;
assign _529_ = _520_ & _528_ /*812*/;
assign _500_ = _520_ ^ _528_ /*813*/;
assign _526_ = _527_ | _529_ /*810*/;
assign _531_ = ~Q[3] /*809*/;
assign _530_ = _531_ & D[4] /*808*/;
assign _533_ = _445_ & _530_ /*803*/;
assign _534_ = _445_ ^ _530_ /*806*/;
assign _535_ = _526_ & _534_ /*804*/;
assign _501_ = _526_ ^ _534_ /*805*/;
assign _532_ = _533_ | _535_ /*802*/;
assign _537_ = ~Q[3] /*801*/;
assign _536_ = _537_ & D[5] /*800*/;
assign _539_ = _446_ & _536_ /*795*/;
assign _540_ = _446_ ^ _536_ /*798*/;
assign _541_ = _532_ & _540_ /*796*/;
assign _502_ = _532_ ^ _540_ /*797*/;
assign _538_ = _539_ | _541_ /*794*/;
assign _543_ = ~Q[3] /*793*/;
assign _542_ = _543_ & D[6] /*792*/;
assign _545_ = _447_ & _542_ /*787*/;
assign _546_ = _447_ ^ _542_ /*790*/;
assign _547_ = _538_ & _546_ /*788*/;
assign _503_ = _538_ ^ _546_ /*789*/;
assign _544_ = _545_ | _547_ /*786*/;
assign _549_ = ~Q[3] /*785*/;
assign _548_ = _549_ & zeroWire /*784*/;
assign _550_ = _448_ ^ _548_ /*782*/;
assign _504_ = _550_ ^ _544_ /*781*/;
assign _565_ = ~D[0] /*751*/;
assign _562_ = R_0[2] & _565_ /*747*/;
assign _563_ = R_0[2] ^ _565_ /*750*/;
assign _564_ = oneWire & _563_ /*748*/;
assign _553_ = oneWire ^ _563_ /*749*/;
assign _561_ = _562_ | _564_ /*746*/;
assign _570_ = ~D[1] /*745*/;
assign _567_ = _497_ & _570_ /*741*/;
assign _568_ = _497_ ^ _570_ /*744*/;
assign _569_ = _561_ & _568_ /*742*/;
assign _554_ = _561_ ^ _568_ /*743*/;
assign _566_ = _567_ | _569_ /*740*/;
assign _575_ = ~D[2] /*739*/;
assign _572_ = _498_ & _575_ /*735*/;
assign _573_ = _498_ ^ _575_ /*738*/;
assign _574_ = _566_ & _573_ /*736*/;
assign _555_ = _566_ ^ _573_ /*737*/;
assign _571_ = _572_ | _574_ /*734*/;
assign _580_ = ~D[3] /*733*/;
assign _577_ = _499_ & _580_ /*729*/;
assign _578_ = _499_ ^ _580_ /*732*/;
assign _579_ = _571_ & _578_ /*730*/;
assign _556_ = _571_ ^ _578_ /*731*/;
assign _576_ = _577_ | _579_ /*728*/;
assign _585_ = ~D[4] /*727*/;
assign _582_ = _500_ & _585_ /*723*/;
assign _583_ = _500_ ^ _585_ /*726*/;
assign _584_ = _576_ & _583_ /*724*/;
assign _557_ = _576_ ^ _583_ /*725*/;
assign _581_ = _582_ | _584_ /*722*/;
assign _590_ = ~D[5] /*721*/;
assign _587_ = _501_ & _590_ /*717*/;
assign _588_ = _501_ ^ _590_ /*720*/;
assign _589_ = _581_ & _588_ /*718*/;
assign _558_ = _581_ ^ _588_ /*719*/;
assign _586_ = _587_ | _589_ /*716*/;
assign _595_ = ~D[6] /*715*/;
assign _592_ = _502_ & _595_ /*711*/;
assign _593_ = _502_ ^ _595_ /*714*/;
assign _594_ = _586_ & _593_ /*712*/;
assign _559_ = _586_ ^ _593_ /*713*/;
assign _591_ = _592_ | _594_ /*710*/;
assign _596_ = _503_ & oneWire /*705*/;
assign _597_ = _503_ ^ oneWire /*708*/;
assign _598_ = _591_ & _597_ /*706*/;
assign _560_ = _591_ ^ _597_ /*707*/;
assign Q[2] = _596_ | _598_ /*704*/;
assign _619_ = ~Q[2] /*655*/;
assign _618_ = _619_ & D[0] /*654*/;
assign _621_ = _553_ & _618_ /*649*/;
assign _622_ = _553_ ^ _618_ /*652*/;
assign _623_ = zeroWire & _622_ /*650*/;
assign _609_ = zeroWire ^ _622_ /*651*/;
assign _620_ = _621_ | _623_ /*648*/;
assign _625_ = ~Q[2] /*647*/;
assign _624_ = _625_ & D[1] /*646*/;
assign _627_ = _554_ & _624_ /*641*/;
assign _628_ = _554_ ^ _624_ /*644*/;
assign _629_ = _620_ & _628_ /*642*/;
assign _610_ = _620_ ^ _628_ /*643*/;
assign _626_ = _627_ | _629_ /*640*/;
assign _631_ = ~Q[2] /*639*/;
assign _630_ = _631_ & D[2] /*638*/;
assign _633_ = _555_ & _630_ /*633*/;
assign _634_ = _555_ ^ _630_ /*636*/;
assign _635_ = _626_ & _634_ /*634*/;
assign _611_ = _626_ ^ _634_ /*635*/;
assign _632_ = _633_ | _635_ /*632*/;
assign _637_ = ~Q[2] /*631*/;
assign _636_ = _637_ & D[3] /*630*/;
assign _639_ = _556_ & _636_ /*625*/;
assign _640_ = _556_ ^ _636_ /*628*/;
assign _641_ = _632_ & _640_ /*626*/;
assign _612_ = _632_ ^ _640_ /*627*/;
assign _638_ = _639_ | _641_ /*624*/;
assign _643_ = ~Q[2] /*623*/;
assign _642_ = _643_ & D[4] /*622*/;
assign _645_ = _557_ & _642_ /*617*/;
assign _646_ = _557_ ^ _642_ /*620*/;
assign _647_ = _638_ & _646_ /*618*/;
assign _613_ = _638_ ^ _646_ /*619*/;
assign _644_ = _645_ | _647_ /*616*/;
assign _649_ = ~Q[2] /*615*/;
assign _648_ = _649_ & D[5] /*614*/;
assign _651_ = _558_ & _648_ /*609*/;
assign _652_ = _558_ ^ _648_ /*612*/;
assign _653_ = _644_ & _652_ /*610*/;
assign _614_ = _644_ ^ _652_ /*611*/;
assign _650_ = _651_ | _653_ /*608*/;
assign _655_ = ~Q[2] /*607*/;
assign _654_ = _655_ & D[6] /*606*/;
assign _657_ = _559_ & _654_ /*601*/;
assign _658_ = _559_ ^ _654_ /*604*/;
assign _659_ = _650_ & _658_ /*602*/;
assign _615_ = _650_ ^ _658_ /*603*/;
assign _656_ = _657_ | _659_ /*600*/;
assign _661_ = ~Q[2] /*599*/;
assign _660_ = _661_ & zeroWire /*598*/;
assign _662_ = _560_ ^ _660_ /*596*/;
assign _616_ = _662_ ^ _656_ /*595*/;
assign _677_ = ~D[0] /*565*/;
assign _674_ = R_0[1] & _677_ /*561*/;
assign _675_ = R_0[1] ^ _677_ /*564*/;
assign _676_ = oneWire & _675_ /*562*/;
assign _665_ = oneWire ^ _675_ /*563*/;
assign _673_ = _674_ | _676_ /*560*/;
assign _682_ = ~D[1] /*559*/;
assign _679_ = _609_ & _682_ /*555*/;
assign _680_ = _609_ ^ _682_ /*558*/;
assign _681_ = _673_ & _680_ /*556*/;
assign _666_ = _673_ ^ _680_ /*557*/;
assign _678_ = _679_ | _681_ /*554*/;
assign _687_ = ~D[2] /*553*/;
assign _684_ = _610_ & _687_ /*549*/;
assign _685_ = _610_ ^ _687_ /*552*/;
assign _686_ = _678_ & _685_ /*550*/;
assign _667_ = _678_ ^ _685_ /*551*/;
assign _683_ = _684_ | _686_ /*548*/;
assign _692_ = ~D[3] /*547*/;
assign _689_ = _611_ & _692_ /*543*/;
assign _690_ = _611_ ^ _692_ /*546*/;
assign _691_ = _683_ & _690_ /*544*/;
assign _668_ = _683_ ^ _690_ /*545*/;
assign _688_ = _689_ | _691_ /*542*/;
assign _697_ = ~D[4] /*541*/;
assign _694_ = _612_ & _697_ /*537*/;
assign _695_ = _612_ ^ _697_ /*540*/;
assign _696_ = _688_ & _695_ /*538*/;
assign _669_ = _688_ ^ _695_ /*539*/;
assign _693_ = _694_ | _696_ /*536*/;
assign _702_ = ~D[5] /*535*/;
assign _699_ = _613_ & _702_ /*531*/;
assign _700_ = _613_ ^ _702_ /*534*/;
assign _701_ = _693_ & _700_ /*532*/;
assign _670_ = _693_ ^ _700_ /*533*/;
assign _698_ = _699_ | _701_ /*530*/;
assign _707_ = ~D[6] /*529*/;
assign _704_ = _614_ & _707_ /*525*/;
assign _705_ = _614_ ^ _707_ /*528*/;
assign _706_ = _698_ & _705_ /*526*/;
assign _671_ = _698_ ^ _705_ /*527*/;
assign _703_ = _704_ | _706_ /*524*/;
assign _708_ = _615_ & oneWire /*519*/;
assign _709_ = _615_ ^ oneWire /*522*/;
assign _710_ = _703_ & _709_ /*520*/;
assign _672_ = _703_ ^ _709_ /*521*/;
assign Q[1] = _708_ | _710_ /*518*/;
assign _731_ = ~Q[1] /*469*/;
assign _730_ = _731_ & D[0] /*468*/;
assign _733_ = _665_ & _730_ /*463*/;
assign _734_ = _665_ ^ _730_ /*466*/;
assign _735_ = zeroWire & _734_ /*464*/;
assign _721_ = zeroWire ^ _734_ /*465*/;
assign _732_ = _733_ | _735_ /*462*/;
assign _737_ = ~Q[1] /*461*/;
assign _736_ = _737_ & D[1] /*460*/;
assign _739_ = _666_ & _736_ /*455*/;
assign _740_ = _666_ ^ _736_ /*458*/;
assign _741_ = _732_ & _740_ /*456*/;
assign _722_ = _732_ ^ _740_ /*457*/;
assign _738_ = _739_ | _741_ /*454*/;
assign _743_ = ~Q[1] /*453*/;
assign _742_ = _743_ & D[2] /*452*/;
assign _745_ = _667_ & _742_ /*447*/;
assign _746_ = _667_ ^ _742_ /*450*/;
assign _747_ = _738_ & _746_ /*448*/;
assign _723_ = _738_ ^ _746_ /*449*/;
assign _744_ = _745_ | _747_ /*446*/;
assign _749_ = ~Q[1] /*445*/;
assign _748_ = _749_ & D[3] /*444*/;
assign _751_ = _668_ & _748_ /*439*/;
assign _752_ = _668_ ^ _748_ /*442*/;
assign _753_ = _744_ & _752_ /*440*/;
assign _724_ = _744_ ^ _752_ /*441*/;
assign _750_ = _751_ | _753_ /*438*/;
assign _755_ = ~Q[1] /*437*/;
assign _754_ = _755_ & D[4] /*436*/;
assign _757_ = _669_ & _754_ /*431*/;
assign _758_ = _669_ ^ _754_ /*434*/;
assign _759_ = _750_ & _758_ /*432*/;
assign _725_ = _750_ ^ _758_ /*433*/;
assign _756_ = _757_ | _759_ /*430*/;
assign _761_ = ~Q[1] /*429*/;
assign _760_ = _761_ & D[5] /*428*/;
assign _763_ = _670_ & _760_ /*423*/;
assign _764_ = _670_ ^ _760_ /*426*/;
assign _765_ = _756_ & _764_ /*424*/;
assign _726_ = _756_ ^ _764_ /*425*/;
assign _762_ = _763_ | _765_ /*422*/;
assign _767_ = ~Q[1] /*421*/;
assign _766_ = _767_ & D[6] /*420*/;
assign _769_ = _671_ & _766_ /*415*/;
assign _770_ = _671_ ^ _766_ /*418*/;
assign _771_ = _762_ & _770_ /*416*/;
assign _727_ = _762_ ^ _770_ /*417*/;
assign _768_ = _769_ | _771_ /*414*/;
assign _773_ = ~Q[1] /*413*/;
assign _772_ = _773_ & zeroWire /*412*/;
assign _774_ = _672_ ^ _772_ /*410*/;
assign _728_ = _774_ ^ _768_ /*409*/;
assign _789_ = ~D[0] /*379*/;
assign _786_ = R_0[0] & _789_ /*375*/;
assign _787_ = R_0[0] ^ _789_ /*378*/;
assign _788_ = oneWire & _787_ /*376*/;
assign _777_ = oneWire ^ _787_ /*377*/;
assign _785_ = _786_ | _788_ /*374*/;
assign _794_ = ~D[1] /*373*/;
assign _791_ = _721_ & _794_ /*369*/;
assign _792_ = _721_ ^ _794_ /*372*/;
assign _793_ = _785_ & _792_ /*370*/;
assign _778_ = _785_ ^ _792_ /*371*/;
assign _790_ = _791_ | _793_ /*368*/;
assign _799_ = ~D[2] /*367*/;
assign _796_ = _722_ & _799_ /*363*/;
assign _797_ = _722_ ^ _799_ /*366*/;
assign _798_ = _790_ & _797_ /*364*/;
assign _779_ = _790_ ^ _797_ /*365*/;
assign _795_ = _796_ | _798_ /*362*/;
assign _804_ = ~D[3] /*361*/;
assign _801_ = _723_ & _804_ /*357*/;
assign _802_ = _723_ ^ _804_ /*360*/;
assign _803_ = _795_ & _802_ /*358*/;
assign _780_ = _795_ ^ _802_ /*359*/;
assign _800_ = _801_ | _803_ /*356*/;
assign _809_ = ~D[4] /*355*/;
assign _806_ = _724_ & _809_ /*351*/;
assign _807_ = _724_ ^ _809_ /*354*/;
assign _808_ = _800_ & _807_ /*352*/;
assign _781_ = _800_ ^ _807_ /*353*/;
assign _805_ = _806_ | _808_ /*350*/;
assign _814_ = ~D[5] /*349*/;
assign _811_ = _725_ & _814_ /*345*/;
assign _812_ = _725_ ^ _814_ /*348*/;
assign _813_ = _805_ & _812_ /*346*/;
assign _782_ = _805_ ^ _812_ /*347*/;
assign _810_ = _811_ | _813_ /*344*/;
assign _819_ = ~D[6] /*343*/;
assign _816_ = _726_ & _819_ /*339*/;
assign _817_ = _726_ ^ _819_ /*342*/;
assign _818_ = _810_ & _817_ /*340*/;
assign _783_ = _810_ ^ _817_ /*341*/;
assign _815_ = _816_ | _818_ /*338*/;
assign _820_ = _727_ & oneWire /*333*/;
assign _821_ = _727_ ^ oneWire /*336*/;
assign _822_ = _815_ & _821_ /*334*/;
assign _784_ = _815_ ^ _821_ /*335*/;
assign Q[0] = _820_ | _822_ /*332*/;
assign _843_ = ~Q[0] /*283*/;
assign _842_ = _843_ & D[0] /*282*/;
assign _845_ = _777_ & _842_ /*277*/;
assign _846_ = _777_ ^ _842_ /*280*/;
assign _847_ = zeroWire & _846_ /*278*/;
assign R_n1[0] = zeroWire ^ _846_ /*279*/;
assign _844_ = _845_ | _847_ /*276*/;
assign _849_ = ~Q[0] /*275*/;
assign _848_ = _849_ & D[1] /*274*/;
assign _851_ = _778_ & _848_ /*269*/;
assign _852_ = _778_ ^ _848_ /*272*/;
assign _853_ = _844_ & _852_ /*270*/;
assign R_n1[1] = _844_ ^ _852_ /*271*/;
assign _850_ = _851_ | _853_ /*268*/;
assign _855_ = ~Q[0] /*267*/;
assign _854_ = _855_ & D[2] /*266*/;
assign _857_ = _779_ & _854_ /*261*/;
assign _858_ = _779_ ^ _854_ /*264*/;
assign _859_ = _850_ & _858_ /*262*/;
assign R_n1[2] = _850_ ^ _858_ /*263*/;
assign _856_ = _857_ | _859_ /*260*/;
assign _861_ = ~Q[0] /*259*/;
assign _860_ = _861_ & D[3] /*258*/;
assign _863_ = _780_ & _860_ /*253*/;
assign _864_ = _780_ ^ _860_ /*256*/;
assign _865_ = _856_ & _864_ /*254*/;
assign R_n1[3] = _856_ ^ _864_ /*255*/;
assign _862_ = _863_ | _865_ /*252*/;
assign _867_ = ~Q[0] /*251*/;
assign _866_ = _867_ & D[4] /*250*/;
assign _869_ = _781_ & _866_ /*245*/;
assign _870_ = _781_ ^ _866_ /*248*/;
assign _871_ = _862_ & _870_ /*246*/;
assign R_n1[4] = _862_ ^ _870_ /*247*/;
assign _868_ = _869_ | _871_ /*244*/;
assign _873_ = ~Q[0] /*243*/;
assign _872_ = _873_ & D[5] /*242*/;
assign _875_ = _782_ & _872_ /*237*/;
assign _876_ = _782_ ^ _872_ /*240*/;
assign _877_ = _868_ & _876_ /*238*/;
assign R_n1[5] = _868_ ^ _876_ /*239*/;
assign _874_ = _875_ | _877_ /*236*/;
assign _879_ = ~Q[0] /*235*/;
assign _878_ = _879_ & D[6] /*234*/;
assign _881_ = _783_ & _878_ /*229*/;
assign _882_ = _783_ ^ _878_ /*232*/;
assign _883_ = _874_ & _882_ /*230*/;
assign R_n1[6] = _874_ ^ _882_ /*231*/;
assign _880_ = _881_ | _883_ /*228*/;
endmodule
