module divider(q, rout, rin, div);
  wire _0_;
  wire _1_;
  wire _2_;
  wire _3_;
  wire _4_;
  wire _5_;
  wire _6_;
  wire _7_;
  wire _8_;
  wire _9_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire [2:0] r_0;
  wire [2:0] r_1;
  wire [1:0] m_1;
  wire [1:0] sum_1;
  wire [1:0] inv_1;
  wire [1:0] r_2;
  wire [1:0] m_2;
  wire [1:0] sum_2;
  wire [1:0] inv_2;
  wire zeroWire;
  wire oneWire;
  input [1:0] rin;
  input [0:0] div;
  output [1:0] q;
  output [1:0] rout;
  assign zeroWire = 1'b0 /*0*/;
  assign oneWire = 1'b1 /*0*/;
  assign r_0[0] = rin[0] /*65*/;
  assign r_0[1] = rin[1] /*64*/;
  assign r_0[2] = zeroWire /*63*/;
  assign inv_1[0] = ~div[0] /*62*/;
assign inv_1[1] = oneWire /*61*/;
  assign _0_ = inv_1[0] ^ r_0[1] /*59*/;
  assign sum_1[0] = _0_ ^ oneWire /*58*/;
  assign _1_ = _0_ & oneWire /*57*/;
  assign _2_ = inv_1[0] & r_0[1] /*56*/;
  assign _3_ = _1_ | _2_ /*55*/;
  assign _4_ = inv_1[1] ^ r_0[2] /*54*/;
  assign sum_1[1] = _4_ ^ _3_ /*53*/;
  assign _5_ = _4_ & _3_ /*52*/;
  assign _6_ = inv_1[1] & r_0[2] /*51*/;
  assign _7_ = _5_ | _6_ /*50*/;
  assign q[1] = ~sum_1[1] /*47*/;
  assign m_1[0] = r_0[1] /*46*/;
  assign m_1[1] = r_0[2] /*45*/;
  assign _8_ = ~q[1] /*43*/;
  assign _9_ = sum_1[0] & q[1] /*42*/;
  assign _10_ = m_1[0] & _8_ /*41*/;
  assign r_1[1] = _10_ | _9_ /*40*/;
  assign _11_ = ~q[1] /*39*/;
  assign _12_ = sum_1[1] & q[1] /*38*/;
  assign _13_ = m_1[1] & _11_ /*37*/;
  assign r_1[2] = _13_ | _12_ /*36*/;
assign r_1[0]= r_0[0] /*35*/;
  assign inv_2[0] = ~div[0] /*32*/;
assign inv_2[1] = oneWire /*31*/;
  assign _14_ = inv_2[0] ^ r_1[0] /*29*/;
  assign sum_2[0] = _14_ ^ oneWire /*28*/;
  assign _15_ = _14_ & oneWire /*27*/;
  assign _16_ = inv_2[0] & r_1[0] /*26*/;
  assign _17_ = _15_ | _16_ /*25*/;
  assign _18_ = inv_2[1] ^ r_1[1] /*24*/;
  assign sum_2[1] = _18_ ^ _17_ /*23*/;
  assign _19_ = _18_ & _17_ /*22*/;
  assign _20_ = inv_2[1] & r_1[1] /*21*/;
  assign _21_ = _19_ | _20_ /*20*/;
  assign q[0] = ~sum_2[1] /*17*/;
  assign m_2[0] = r_1[0] /*16*/;
  assign m_2[1] = r_1[1] /*15*/;
  assign _22_ = ~q[0] /*13*/;
  assign _23_ = sum_2[0] & q[0] /*12*/;
  assign _24_ = m_2[0] & _22_ /*11*/;
  assign r_2[0] = _24_ | _23_ /*10*/;
  assign _25_ = ~q[0] /*9*/;
  assign _26_ = sum_2[1] & q[0] /*8*/;
  assign _27_ = m_2[1] & _25_ /*7*/;
  assign r_2[1] = _27_ | _26_ /*6*/;
  assign rout[0] = r_2[0] /*0*/;
  assign rout[1] = r_2[1] /*1*/;
endmodule