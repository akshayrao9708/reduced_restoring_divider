module divider(q, rout, rin, div);
  wire _0_;
  wire _1_;
  wire _2_;
  wire _3_;
  wire _4_;
  wire _5_;
  wire _6_;
  wire _7_;
  wire _8_;
  wire _9_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  wire _38_;
  wire _39_;
  wire _40_;
  wire _41_;
  wire _42_;
  wire _43_;
  wire _44_;
  wire _45_;
  wire _46_;
  wire _47_;
  wire _48_;
  wire _49_;
  wire _50_;
  wire _51_;
  wire _52_;
  wire _53_;
  wire _54_;
  wire _55_;
  wire _56_;
  wire _57_;
  wire _58_;
  wire _59_;
  wire _60_;
  wire _61_;
  wire _62_;
  wire [4:0] r_0;
  wire [4:0] r_1;
  wire [2:0] m_1;
  wire [2:0] sum_1;
  wire [2:0] inv_1;
  wire [3:0] r_2;
  wire [2:0] m_2;
  wire [2:0] sum_2;
  wire [2:0] inv_2;
  wire [2:0] r_3;
  wire [2:0] m_3;
  wire [2:0] sum_3;
  wire [2:0] inv_3;
  wire zeroWire;
  wire oneWire;
  input [3:0] rin;
  input [1:0] div;
  output [2:0] q;
  output [2:0] rout;
  assign zeroWire = 1'b0 /*0*/;
  assign oneWire = 1'b1 /*0*/;
  assign r_0[0] = rin[0] /*149*/;
  assign r_0[1] = rin[1] /*148*/;
  assign r_0[2] = rin[2] /*147*/;
  assign r_0[3] = rin[3] /*146*/;
  assign r_0[4] = zeroWire /*145*/;
  assign inv_1[0] = ~div[0] /*144*/;
  assign inv_1[1] = ~div[1] /*143*/;
assign inv_1[2] = oneWire /*142*/;
  assign _0_ = inv_1[0] ^ r_0[2] /*140*/;
  assign sum_1[0] = _0_ ^ oneWire /*139*/;
  assign _1_ = _0_ & oneWire /*138*/;
  assign _2_ = inv_1[0] & r_0[2] /*137*/;
  assign _3_ = _1_ | _2_ /*136*/;
  assign _4_ = inv_1[1] ^ r_0[3] /*135*/;
  assign sum_1[1] = _4_ ^ _3_ /*134*/;
  assign _5_ = _4_ & _3_ /*133*/;
  assign _6_ = inv_1[1] & r_0[3] /*132*/;
  assign _7_ = _5_ | _6_ /*131*/;
  assign _8_ = inv_1[2] ^ r_0[4] /*129*/;
  assign sum_1[2] = _8_ ^ _7_ /*128*/;
  assign _9_ = _8_ & _7_ /*127*/;
  assign _10_ = inv_1[2] & r_0[4] /*126*/;
  assign _11_ = _9_ | _10_ /*125*/;
  assign q[2] = ~sum_1[2] /*123*/;
  assign m_1[0] = r_0[2] /*122*/;
  assign m_1[1] = r_0[3] /*121*/;
  assign m_1[2] = r_0[4] /*120*/;
  assign _12_ = ~q[2] /*118*/;
  assign _13_ = sum_1[0] & q[2] /*117*/;
  assign _14_ = m_1[0] & _12_ /*116*/;
  assign r_1[2] = _14_ | _13_ /*115*/;
  assign _15_ = ~q[2] /*114*/;
  assign _16_ = sum_1[1] & q[2] /*113*/;
  assign _17_ = m_1[1] & _15_ /*112*/;
  assign r_1[3] = _17_ | _16_ /*111*/;
  assign _18_ = ~q[2] /*110*/;
  assign _19_ = sum_1[2] & q[2] /*109*/;
  assign _20_ = m_1[2] & _18_ /*108*/;
  assign r_1[4] = _20_ | _19_ /*107*/;
assign r_1[0]= r_0[0] /*106*/;
assign r_1[1]= r_0[1] /*105*/;
  assign inv_2[0] = ~div[0] /*102*/;
  assign inv_2[1] = ~div[1] /*101*/;
assign inv_2[2] = oneWire /*100*/;
  assign _21_ = inv_2[0] ^ r_1[1] /*98*/;
  assign sum_2[0] = _21_ ^ oneWire /*97*/;
  assign _22_ = _21_ & oneWire /*96*/;
  assign _23_ = inv_2[0] & r_1[1] /*95*/;
  assign _24_ = _22_ | _23_ /*94*/;
  assign _25_ = inv_2[1] ^ r_1[2] /*93*/;
  assign sum_2[1] = _25_ ^ _24_ /*92*/;
  assign _26_ = _25_ & _24_ /*91*/;
  assign _27_ = inv_2[1] & r_1[2] /*90*/;
  assign _28_ = _26_ | _27_ /*89*/;
  assign _29_ = inv_2[2] ^ r_1[3] /*87*/;
  assign sum_2[2] = _29_ ^ _28_ /*86*/;
  assign _30_ = _29_ & _28_ /*85*/;
  assign _31_ = inv_2[2] & r_1[3] /*84*/;
  assign _32_ = _30_ | _31_ /*83*/;
  assign q[1] = ~sum_2[2] /*81*/;
  assign m_2[0] = r_1[1] /*80*/;
  assign m_2[1] = r_1[2] /*79*/;
  assign m_2[2] = r_1[3] /*78*/;
  assign _33_ = ~q[1] /*76*/;
  assign _34_ = sum_2[0] & q[1] /*75*/;
  assign _35_ = m_2[0] & _33_ /*74*/;
  assign r_2[1] = _35_ | _34_ /*73*/;
  assign _36_ = ~q[1] /*72*/;
  assign _37_ = sum_2[1] & q[1] /*71*/;
  assign _38_ = m_2[1] & _36_ /*70*/;
  assign r_2[2] = _38_ | _37_ /*69*/;
  assign _39_ = ~q[1] /*68*/;
  assign _40_ = sum_2[2] & q[1] /*67*/;
  assign _41_ = m_2[2] & _39_ /*66*/;
  assign r_2[3] = _41_ | _40_ /*65*/;
  assign r_2[0]= r_1[0] /*64*/;
  assign inv_3[0] = ~div[0] /*60*/;
  assign inv_3[1] = ~div[1] /*59*/;
  assign inv_3[2] = oneWire /*58*/;
  assign _42_ = inv_3[0] ^ r_2[0] /*56*/;
  assign sum_3[0] = _42_ ^ oneWire /*55*/;
  assign _43_ = _42_ & oneWire /*54*/;
  assign _44_ = inv_3[0] & r_2[0] /*53*/;
  assign _45_ = _43_ | _44_ /*52*/;
  assign _46_ = inv_3[1] ^ r_2[1] /*51*/;
  assign sum_3[1] = _46_ ^ _45_ /*50*/;
  assign _47_ = _46_ & _45_ /*49*/;
  assign _48_ = inv_3[1] & r_2[1] /*48*/;
  assign _49_ = _47_ | _48_ /*47*/;
  assign _50_ = inv_3[2] ^ r_2[2] /*45*/;
  assign sum_3[2] = _50_ ^ _49_ /*44*/;
  assign _51_ = _50_ & _49_ /*43*/;
  assign _52_ = inv_3[2] & r_2[2] /*42*/;
  assign _53_ = _51_ | _52_ /*41*/;
  assign q[0] = ~sum_3[2] /*39*/;
  assign m_3[0] = r_2[0] /*38*/;
  assign m_3[1] = r_2[1] /*37*/;
  assign m_3[2] = r_2[2] /*36*/;
  assign _54_ = ~q[0] /*34*/;
  assign _55_ = sum_3[0] & q[0] /*33*/;
  assign _56_ = m_3[0] & _54_ /*32*/;
  assign r_3[0] = _56_ | _55_ /*31*/;
  assign _57_ = ~q[0] /*30*/;
  assign _58_ = sum_3[1] & q[0] /*29*/;
  assign _59_ = m_3[1] & _57_ /*28*/;
  assign r_3[1] = _59_ | _58_ /*27*/;
  assign _60_ = ~q[0] /*26*/;
  assign _61_ = sum_3[2] & q[0] /*25*/;
  assign _62_ = m_3[2] & _60_ /*24*/;
  assign r_3[2] = _62_ | _61_ /*23*/;
  assign rout[0] = r_3[0] /*0*/;
  assign rout[1] = r_3[1] /*1*/;
  assign rout[2] = r_3[2] /*2*/;
endmodule