module nonresdivReduced(R_0, D, Q, R_n1);
input [13:0] R_0;
input [6:0] D;
output [7:0] Q;
output [6:0] R_n1;
wire _0_;
wire _1_;
wire _2_;
wire _3_;
wire _4_;
wire _5_;
wire _6_;
wire _7_;
wire _8_;
wire _9_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire _30_;
wire _31_;
wire _32_;
wire _33_;
wire _34_;
wire _35_;
wire _36_;
wire _37_;
wire _38_;
wire _39_;
wire _40_;
wire _41_;
wire _42_;
wire _43_;
wire _44_;
wire _45_;
wire _46_;
wire _47_;
wire _48_;
wire _49_;
wire _50_;
wire _51_;
wire _52_;
wire _53_;
wire _54_;
wire _55_;
wire _56_;
wire _57_;
wire _58_;
wire _59_;
wire _60_;
wire _61_;
wire _62_;
wire _63_;
wire _64_;
wire _65_;
wire _66_;
wire _67_;
wire _68_;
wire _69_;
wire _70_;
wire _71_;
wire _72_;
wire _73_;
wire _74_;
wire _75_;
wire _76_;
wire _77_;
wire _78_;
wire _79_;
wire _80_;
wire _81_;
wire _82_;
wire _83_;
wire _84_;
wire _85_;
wire _86_;
wire _87_;
wire _88_;
wire _89_;
wire _90_;
wire _91_;
wire _92_;
wire _93_;
wire _94_;
wire _95_;
wire _96_;
wire _97_;
wire _98_;
wire _99_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
wire _255_;
wire _256_;
wire _257_;
wire _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire _267_;
wire _268_;
wire _269_;
wire _270_;
wire _271_;
wire _272_;
wire _273_;
wire _274_;
wire _275_;
wire _276_;
wire _277_;
wire _278_;
wire _279_;
wire _280_;
wire _281_;
wire _282_;
wire _283_;
wire _284_;
wire _285_;
wire _286_;
wire _287_;
wire _288_;
wire _289_;
wire _290_;
wire _291_;
wire _292_;
wire _293_;
wire _294_;
wire _295_;
wire _296_;
wire _297_;
wire _298_;
wire _299_;
wire _300_;
wire _301_;
wire _302_;
wire _303_;
wire _304_;
wire _305_;
wire _306_;
wire _307_;
wire _308_;
wire _309_;
wire _310_;
wire _311_;
wire _312_;
wire _313_;
wire _314_;
wire _315_;
wire _316_;
wire _317_;
wire _318_;
wire _319_;
wire _320_;
wire _321_;
wire _322_;
wire _323_;
wire _324_;
wire _325_;
wire _326_;
wire _327_;
wire _328_;
wire _329_;
wire _330_;
wire _331_;
wire _332_;
wire _333_;
wire _334_;
wire _335_;
wire _336_;
wire _337_;
wire _338_;
wire _339_;
wire _340_;
wire _341_;
wire _342_;
wire _343_;
wire _344_;
wire _345_;
wire _346_;
wire _347_;
wire _348_;
wire _349_;
wire _350_;
wire _351_;
wire _352_;
wire _353_;
wire _354_;
wire _355_;
wire _356_;
wire _357_;
wire _358_;
wire _359_;
wire _360_;
wire _361_;
wire _362_;
wire _363_;
wire _364_;
wire _365_;
wire _366_;
wire _367_;
wire _368_;
wire _369_;
wire _370_;
wire _371_;
wire _372_;
wire _373_;
wire _374_;
wire _375_;
wire _376_;
wire _377_;
wire _378_;
wire _379_;
wire _380_;
wire _381_;
wire _382_;
wire _383_;
wire _384_;
wire _385_;
wire _386_;
wire _387_;
wire _388_;
wire _389_;
wire _390_;
wire _391_;
wire _392_;
wire _393_;
wire _394_;
wire _395_;
wire _396_;
wire _397_;
wire _398_;
wire _399_;
wire _400_;
wire _401_;
wire _402_;
wire _403_;
wire _404_;
wire _405_;
wire _406_;
wire _407_;
wire _408_;
wire _409_;
wire _410_;
wire _411_;
wire _412_;
wire _413_;
wire _414_;
wire _415_;
wire _416_;
wire _417_;
wire _418_;
wire _419_;
wire _420_;
wire _421_;
wire _422_;
wire _423_;
wire _424_;
wire _425_;
wire _426_;
wire _427_;
wire _428_;
wire _429_;
wire _430_;
wire _431_;
wire _432_;
wire _433_;
wire _434_;
wire _435_;
wire _436_;
wire _437_;
wire _438_;
wire _439_;
wire _440_;
wire _441_;
wire _442_;
wire _443_;
wire _444_;
wire _445_;
wire _446_;
wire _447_;
wire _448_;
wire _449_;
wire _450_;
wire _451_;
wire _452_;
wire _453_;
wire _454_;
wire _455_;
wire _456_;
wire _457_;
wire _458_;
wire _459_;
wire _460_;
wire _461_;
wire _462_;
wire _463_;
wire _464_;
wire _465_;
wire _466_;
wire _467_;
wire _468_;
wire _469_;
wire _470_;
wire _471_;
wire _472_;
wire _473_;
wire _474_;
wire _475_;
wire _476_;
wire _477_;
wire _478_;
wire _479_;
wire _480_;
wire _481_;
wire _482_;
wire _483_;
wire _484_;
wire _485_;
wire _486_;
wire zeroWire;
wire oneWire;
assign zeroWire = 1'b0 /*899*/;
assign oneWire = 1'b1 /*899*/;
assign _13_ = ~D[0] /*849*/;
assign _10_ = R_0[7] & _13_ /*845*/;
assign _11_ = R_0[7] ^ _13_ /*848*/;
assign _12_ = oneWire & _11_ /*846*/;
assign _0_ = oneWire ^ _11_ /*847*/;
assign _9_ = _10_ | _12_ /*844*/;
assign _18_ = ~D[1] /*843*/;
assign _15_ = R_0[8] & _18_ /*839*/;
assign _16_ = R_0[8] ^ _18_ /*842*/;
assign _17_ = _9_ & _16_ /*840*/;
assign _1_ = _9_ ^ _16_ /*841*/;
assign _14_ = _15_ | _17_ /*838*/;
assign _23_ = ~D[2] /*837*/;
assign _20_ = R_0[9] & _23_ /*833*/;
assign _21_ = R_0[9] ^ _23_ /*836*/;
assign _22_ = _14_ & _21_ /*834*/;
assign _2_ = _14_ ^ _21_ /*835*/;
assign _19_ = _20_ | _22_ /*832*/;
assign _28_ = ~D[3] /*831*/;
assign _25_ = R_0[10] & _28_ /*827*/;
assign _26_ = R_0[10] ^ _28_ /*830*/;
assign _27_ = _19_ & _26_ /*828*/;
assign _3_ = _19_ ^ _26_ /*829*/;
assign _24_ = _25_ | _27_ /*826*/;
assign _33_ = ~D[4] /*825*/;
assign _30_ = R_0[11] & _33_ /*821*/;
assign _31_ = R_0[11] ^ _33_ /*824*/;
assign _32_ = _24_ & _31_ /*822*/;
assign _4_ = _24_ ^ _31_ /*823*/;
assign _29_ = _30_ | _32_ /*820*/;
assign _38_ = ~D[5] /*819*/;
assign _35_ = R_0[12] & _38_ /*815*/;
assign _36_ = R_0[12] ^ _38_ /*818*/;
assign _37_ = _29_ & _36_ /*816*/;
assign _5_ = _29_ ^ _36_ /*817*/;
assign _34_ = _35_ | _37_ /*814*/;
assign _43_ = ~D[6] /*813*/;
assign _40_ = R_0[13] & _43_ /*809*/;
assign _41_ = R_0[13] ^ _43_ /*812*/;
assign _42_ = _34_ & _41_ /*810*/;
assign _6_ = _34_ ^ _41_ /*811*/;
assign _39_ = _40_ | _42_ /*808*/;
assign _44_ = zeroWire & oneWire /*803*/;
assign _45_ = zeroWire ^ oneWire /*806*/;
assign _46_ = _39_ & _45_ /*804*/;
assign _7_ = _39_ ^ _45_ /*805*/;
assign Q[7] = _44_ | _46_ /*802*/;
assign _62_ = D[0] ^ Q[7] /*754*/;
assign _59_ = R_0[6] & _62_ /*750*/;
assign _60_ = R_0[6] ^ _62_ /*753*/;
assign _61_ = Q[7] & _60_ /*751*/;
assign _49_ = Q[7] ^ _60_ /*752*/;
assign _58_ = _59_ | _61_ /*749*/;
assign _67_ = D[1] ^ Q[7] /*748*/;
assign _64_ = _0_ & _67_ /*744*/;
assign _65_ = _0_ ^ _67_ /*747*/;
assign _66_ = _58_ & _65_ /*745*/;
assign _50_ = _58_ ^ _65_ /*746*/;
assign _63_ = _64_ | _66_ /*743*/;
assign _72_ = D[2] ^ Q[7] /*742*/;
assign _69_ = _1_ & _72_ /*738*/;
assign _70_ = _1_ ^ _72_ /*741*/;
assign _71_ = _63_ & _70_ /*739*/;
assign _51_ = _63_ ^ _70_ /*740*/;
assign _68_ = _69_ | _71_ /*737*/;
assign _77_ = D[3] ^ Q[7] /*736*/;
assign _74_ = _2_ & _77_ /*732*/;
assign _75_ = _2_ ^ _77_ /*735*/;
assign _76_ = _68_ & _75_ /*733*/;
assign _52_ = _68_ ^ _75_ /*734*/;
assign _73_ = _74_ | _76_ /*731*/;
assign _82_ = D[4] ^ Q[7] /*730*/;
assign _79_ = _3_ & _82_ /*726*/;
assign _80_ = _3_ ^ _82_ /*729*/;
assign _81_ = _73_ & _80_ /*727*/;
assign _53_ = _73_ ^ _80_ /*728*/;
assign _78_ = _79_ | _81_ /*725*/;
assign _87_ = D[5] ^ Q[7] /*724*/;
assign _84_ = _4_ & _87_ /*720*/;
assign _85_ = _4_ ^ _87_ /*723*/;
assign _86_ = _78_ & _85_ /*721*/;
assign _54_ = _78_ ^ _85_ /*722*/;
assign _83_ = _84_ | _86_ /*719*/;
assign _92_ = D[6] ^ Q[7] /*718*/;
assign _89_ = _5_ & _92_ /*714*/;
assign _90_ = _5_ ^ _92_ /*717*/;
assign _91_ = _83_ & _90_ /*715*/;
assign _55_ = _83_ ^ _90_ /*716*/;
assign _88_ = _89_ | _91_ /*713*/;
assign _96_ = zeroWire ^ Q[7] /*712*/;
assign _93_ = _6_ & _96_ /*708*/;
assign _94_ = _6_ ^ _96_ /*711*/;
assign _95_ = _88_ & _94_ /*709*/;
assign _56_ = _88_ ^ _94_ /*710*/;
assign Q[6] = _93_ | _95_ /*707*/;
assign _111_ = D[0] ^ Q[6] /*657*/;
assign _108_ = R_0[5] & _111_ /*653*/;
assign _109_ = R_0[5] ^ _111_ /*656*/;
assign _110_ = Q[6] & _109_ /*654*/;
assign _98_ = Q[6] ^ _109_ /*655*/;
assign _107_ = _108_ | _110_ /*652*/;
assign _116_ = D[1] ^ Q[6] /*651*/;
assign _113_ = _49_ & _116_ /*647*/;
assign _114_ = _49_ ^ _116_ /*650*/;
assign _115_ = _107_ & _114_ /*648*/;
assign _99_ = _107_ ^ _114_ /*649*/;
assign _112_ = _113_ | _115_ /*646*/;
assign _121_ = D[2] ^ Q[6] /*645*/;
assign _118_ = _50_ & _121_ /*641*/;
assign _119_ = _50_ ^ _121_ /*644*/;
assign _120_ = _112_ & _119_ /*642*/;
assign _100_ = _112_ ^ _119_ /*643*/;
assign _117_ = _118_ | _120_ /*640*/;
assign _126_ = D[3] ^ Q[6] /*639*/;
assign _123_ = _51_ & _126_ /*635*/;
assign _124_ = _51_ ^ _126_ /*638*/;
assign _125_ = _117_ & _124_ /*636*/;
assign _101_ = _117_ ^ _124_ /*637*/;
assign _122_ = _123_ | _125_ /*634*/;
assign _131_ = D[4] ^ Q[6] /*633*/;
assign _128_ = _52_ & _131_ /*629*/;
assign _129_ = _52_ ^ _131_ /*632*/;
assign _130_ = _122_ & _129_ /*630*/;
assign _102_ = _122_ ^ _129_ /*631*/;
assign _127_ = _128_ | _130_ /*628*/;
assign _136_ = D[5] ^ Q[6] /*627*/;
assign _133_ = _53_ & _136_ /*623*/;
assign _134_ = _53_ ^ _136_ /*626*/;
assign _135_ = _127_ & _134_ /*624*/;
assign _103_ = _127_ ^ _134_ /*625*/;
assign _132_ = _133_ | _135_ /*622*/;
assign _141_ = D[6] ^ Q[6] /*621*/;
assign _138_ = _54_ & _141_ /*617*/;
assign _139_ = _54_ ^ _141_ /*620*/;
assign _140_ = _132_ & _139_ /*618*/;
assign _104_ = _132_ ^ _139_ /*619*/;
assign _137_ = _138_ | _140_ /*616*/;
assign _145_ = zeroWire ^ Q[6] /*615*/;
assign _142_ = _55_ & _145_ /*611*/;
assign _143_ = _55_ ^ _145_ /*614*/;
assign _144_ = _137_ & _143_ /*612*/;
assign _105_ = _137_ ^ _143_ /*613*/;
assign Q[5] = _142_ | _144_ /*610*/;
assign _160_ = D[0] ^ Q[5] /*560*/;
assign _157_ = R_0[4] & _160_ /*556*/;
assign _158_ = R_0[4] ^ _160_ /*559*/;
assign _159_ = Q[5] & _158_ /*557*/;
assign _147_ = Q[5] ^ _158_ /*558*/;
assign _156_ = _157_ | _159_ /*555*/;
assign _165_ = D[1] ^ Q[5] /*554*/;
assign _162_ = _98_ & _165_ /*550*/;
assign _163_ = _98_ ^ _165_ /*553*/;
assign _164_ = _156_ & _163_ /*551*/;
assign _148_ = _156_ ^ _163_ /*552*/;
assign _161_ = _162_ | _164_ /*549*/;
assign _170_ = D[2] ^ Q[5] /*548*/;
assign _167_ = _99_ & _170_ /*544*/;
assign _168_ = _99_ ^ _170_ /*547*/;
assign _169_ = _161_ & _168_ /*545*/;
assign _149_ = _161_ ^ _168_ /*546*/;
assign _166_ = _167_ | _169_ /*543*/;
assign _175_ = D[3] ^ Q[5] /*542*/;
assign _172_ = _100_ & _175_ /*538*/;
assign _173_ = _100_ ^ _175_ /*541*/;
assign _174_ = _166_ & _173_ /*539*/;
assign _150_ = _166_ ^ _173_ /*540*/;
assign _171_ = _172_ | _174_ /*537*/;
assign _180_ = D[4] ^ Q[5] /*536*/;
assign _177_ = _101_ & _180_ /*532*/;
assign _178_ = _101_ ^ _180_ /*535*/;
assign _179_ = _171_ & _178_ /*533*/;
assign _151_ = _171_ ^ _178_ /*534*/;
assign _176_ = _177_ | _179_ /*531*/;
assign _185_ = D[5] ^ Q[5] /*530*/;
assign _182_ = _102_ & _185_ /*526*/;
assign _183_ = _102_ ^ _185_ /*529*/;
assign _184_ = _176_ & _183_ /*527*/;
assign _152_ = _176_ ^ _183_ /*528*/;
assign _181_ = _182_ | _184_ /*525*/;
assign _190_ = D[6] ^ Q[5] /*524*/;
assign _187_ = _103_ & _190_ /*520*/;
assign _188_ = _103_ ^ _190_ /*523*/;
assign _189_ = _181_ & _188_ /*521*/;
assign _153_ = _181_ ^ _188_ /*522*/;
assign _186_ = _187_ | _189_ /*519*/;
assign _194_ = zeroWire ^ Q[5] /*518*/;
assign _191_ = _104_ & _194_ /*514*/;
assign _192_ = _104_ ^ _194_ /*517*/;
assign _193_ = _186_ & _192_ /*515*/;
assign _154_ = _186_ ^ _192_ /*516*/;
assign Q[4] = _191_ | _193_ /*513*/;
assign _209_ = D[0] ^ Q[4] /*463*/;
assign _206_ = R_0[3] & _209_ /*459*/;
assign _207_ = R_0[3] ^ _209_ /*462*/;
assign _208_ = Q[4] & _207_ /*460*/;
assign _196_ = Q[4] ^ _207_ /*461*/;
assign _205_ = _206_ | _208_ /*458*/;
assign _214_ = D[1] ^ Q[4] /*457*/;
assign _211_ = _147_ & _214_ /*453*/;
assign _212_ = _147_ ^ _214_ /*456*/;
assign _213_ = _205_ & _212_ /*454*/;
assign _197_ = _205_ ^ _212_ /*455*/;
assign _210_ = _211_ | _213_ /*452*/;
assign _219_ = D[2] ^ Q[4] /*451*/;
assign _216_ = _148_ & _219_ /*447*/;
assign _217_ = _148_ ^ _219_ /*450*/;
assign _218_ = _210_ & _217_ /*448*/;
assign _198_ = _210_ ^ _217_ /*449*/;
assign _215_ = _216_ | _218_ /*446*/;
assign _224_ = D[3] ^ Q[4] /*445*/;
assign _221_ = _149_ & _224_ /*441*/;
assign _222_ = _149_ ^ _224_ /*444*/;
assign _223_ = _215_ & _222_ /*442*/;
assign _199_ = _215_ ^ _222_ /*443*/;
assign _220_ = _221_ | _223_ /*440*/;
assign _229_ = D[4] ^ Q[4] /*439*/;
assign _226_ = _150_ & _229_ /*435*/;
assign _227_ = _150_ ^ _229_ /*438*/;
assign _228_ = _220_ & _227_ /*436*/;
assign _200_ = _220_ ^ _227_ /*437*/;
assign _225_ = _226_ | _228_ /*434*/;
assign _234_ = D[5] ^ Q[4] /*433*/;
assign _231_ = _151_ & _234_ /*429*/;
assign _232_ = _151_ ^ _234_ /*432*/;
assign _233_ = _225_ & _232_ /*430*/;
assign _201_ = _225_ ^ _232_ /*431*/;
assign _230_ = _231_ | _233_ /*428*/;
assign _239_ = D[6] ^ Q[4] /*427*/;
assign _236_ = _152_ & _239_ /*423*/;
assign _237_ = _152_ ^ _239_ /*426*/;
assign _238_ = _230_ & _237_ /*424*/;
assign _202_ = _230_ ^ _237_ /*425*/;
assign _235_ = _236_ | _238_ /*422*/;
assign _243_ = zeroWire ^ Q[4] /*421*/;
assign _240_ = _153_ & _243_ /*417*/;
assign _241_ = _153_ ^ _243_ /*420*/;
assign _242_ = _235_ & _241_ /*418*/;
assign _203_ = _235_ ^ _241_ /*419*/;
assign Q[3] = _240_ | _242_ /*416*/;
assign _258_ = D[0] ^ Q[3] /*366*/;
assign _255_ = R_0[2] & _258_ /*362*/;
assign _256_ = R_0[2] ^ _258_ /*365*/;
assign _257_ = Q[3] & _256_ /*363*/;
assign _245_ = Q[3] ^ _256_ /*364*/;
assign _254_ = _255_ | _257_ /*361*/;
assign _263_ = D[1] ^ Q[3] /*360*/;
assign _260_ = _196_ & _263_ /*356*/;
assign _261_ = _196_ ^ _263_ /*359*/;
assign _262_ = _254_ & _261_ /*357*/;
assign _246_ = _254_ ^ _261_ /*358*/;
assign _259_ = _260_ | _262_ /*355*/;
assign _268_ = D[2] ^ Q[3] /*354*/;
assign _265_ = _197_ & _268_ /*350*/;
assign _266_ = _197_ ^ _268_ /*353*/;
assign _267_ = _259_ & _266_ /*351*/;
assign _247_ = _259_ ^ _266_ /*352*/;
assign _264_ = _265_ | _267_ /*349*/;
assign _273_ = D[3] ^ Q[3] /*348*/;
assign _270_ = _198_ & _273_ /*344*/;
assign _271_ = _198_ ^ _273_ /*347*/;
assign _272_ = _264_ & _271_ /*345*/;
assign _248_ = _264_ ^ _271_ /*346*/;
assign _269_ = _270_ | _272_ /*343*/;
assign _278_ = D[4] ^ Q[3] /*342*/;
assign _275_ = _199_ & _278_ /*338*/;
assign _276_ = _199_ ^ _278_ /*341*/;
assign _277_ = _269_ & _276_ /*339*/;
assign _249_ = _269_ ^ _276_ /*340*/;
assign _274_ = _275_ | _277_ /*337*/;
assign _283_ = D[5] ^ Q[3] /*336*/;
assign _280_ = _200_ & _283_ /*332*/;
assign _281_ = _200_ ^ _283_ /*335*/;
assign _282_ = _274_ & _281_ /*333*/;
assign _250_ = _274_ ^ _281_ /*334*/;
assign _279_ = _280_ | _282_ /*331*/;
assign _288_ = D[6] ^ Q[3] /*330*/;
assign _285_ = _201_ & _288_ /*326*/;
assign _286_ = _201_ ^ _288_ /*329*/;
assign _287_ = _279_ & _286_ /*327*/;
assign _251_ = _279_ ^ _286_ /*328*/;
assign _284_ = _285_ | _287_ /*325*/;
assign _292_ = zeroWire ^ Q[3] /*324*/;
assign _289_ = _202_ & _292_ /*320*/;
assign _290_ = _202_ ^ _292_ /*323*/;
assign _291_ = _284_ & _290_ /*321*/;
assign _252_ = _284_ ^ _290_ /*322*/;
assign Q[2] = _289_ | _291_ /*319*/;
assign _307_ = D[0] ^ Q[2] /*269*/;
assign _304_ = R_0[1] & _307_ /*265*/;
assign _305_ = R_0[1] ^ _307_ /*268*/;
assign _306_ = Q[2] & _305_ /*266*/;
assign _294_ = Q[2] ^ _305_ /*267*/;
assign _303_ = _304_ | _306_ /*264*/;
assign _312_ = D[1] ^ Q[2] /*263*/;
assign _309_ = _245_ & _312_ /*259*/;
assign _310_ = _245_ ^ _312_ /*262*/;
assign _311_ = _303_ & _310_ /*260*/;
assign _295_ = _303_ ^ _310_ /*261*/;
assign _308_ = _309_ | _311_ /*258*/;
assign _317_ = D[2] ^ Q[2] /*257*/;
assign _314_ = _246_ & _317_ /*253*/;
assign _315_ = _246_ ^ _317_ /*256*/;
assign _316_ = _308_ & _315_ /*254*/;
assign _296_ = _308_ ^ _315_ /*255*/;
assign _313_ = _314_ | _316_ /*252*/;
assign _322_ = D[3] ^ Q[2] /*251*/;
assign _319_ = _247_ & _322_ /*247*/;
assign _320_ = _247_ ^ _322_ /*250*/;
assign _321_ = _313_ & _320_ /*248*/;
assign _297_ = _313_ ^ _320_ /*249*/;
assign _318_ = _319_ | _321_ /*246*/;
assign _327_ = D[4] ^ Q[2] /*245*/;
assign _324_ = _248_ & _327_ /*241*/;
assign _325_ = _248_ ^ _327_ /*244*/;
assign _326_ = _318_ & _325_ /*242*/;
assign _298_ = _318_ ^ _325_ /*243*/;
assign _323_ = _324_ | _326_ /*240*/;
assign _332_ = D[5] ^ Q[2] /*239*/;
assign _329_ = _249_ & _332_ /*235*/;
assign _330_ = _249_ ^ _332_ /*238*/;
assign _331_ = _323_ & _330_ /*236*/;
assign _299_ = _323_ ^ _330_ /*237*/;
assign _328_ = _329_ | _331_ /*234*/;
assign _337_ = D[6] ^ Q[2] /*233*/;
assign _334_ = _250_ & _337_ /*229*/;
assign _335_ = _250_ ^ _337_ /*232*/;
assign _336_ = _328_ & _335_ /*230*/;
assign _300_ = _328_ ^ _335_ /*231*/;
assign _333_ = _334_ | _336_ /*228*/;
assign _341_ = zeroWire ^ Q[2] /*227*/;
assign _338_ = _251_ & _341_ /*223*/;
assign _339_ = _251_ ^ _341_ /*226*/;
assign _340_ = _333_ & _339_ /*224*/;
assign _301_ = _333_ ^ _339_ /*225*/;
assign Q[1] = _338_ | _340_ /*222*/;
assign _356_ = D[0] ^ Q[1] /*172*/;
assign _353_ = R_0[0] & _356_ /*168*/;
assign _354_ = R_0[0] ^ _356_ /*171*/;
assign _355_ = Q[1] & _354_ /*169*/;
assign _343_ = Q[1] ^ _354_ /*170*/;
assign _352_ = _353_ | _355_ /*167*/;
assign _361_ = D[1] ^ Q[1] /*166*/;
assign _358_ = _294_ & _361_ /*162*/;
assign _359_ = _294_ ^ _361_ /*165*/;
assign _360_ = _352_ & _359_ /*163*/;
assign _344_ = _352_ ^ _359_ /*164*/;
assign _357_ = _358_ | _360_ /*161*/;
assign _366_ = D[2] ^ Q[1] /*160*/;
assign _363_ = _295_ & _366_ /*156*/;
assign _364_ = _295_ ^ _366_ /*159*/;
assign _365_ = _357_ & _364_ /*157*/;
assign _345_ = _357_ ^ _364_ /*158*/;
assign _362_ = _363_ | _365_ /*155*/;
assign _371_ = D[3] ^ Q[1] /*154*/;
assign _368_ = _296_ & _371_ /*150*/;
assign _369_ = _296_ ^ _371_ /*153*/;
assign _370_ = _362_ & _369_ /*151*/;
assign _346_ = _362_ ^ _369_ /*152*/;
assign _367_ = _368_ | _370_ /*149*/;
assign _376_ = D[4] ^ Q[1] /*148*/;
assign _373_ = _297_ & _376_ /*144*/;
assign _374_ = _297_ ^ _376_ /*147*/;
assign _375_ = _367_ & _374_ /*145*/;
assign _347_ = _367_ ^ _374_ /*146*/;
assign _372_ = _373_ | _375_ /*143*/;
assign _381_ = D[5] ^ Q[1] /*142*/;
assign _378_ = _298_ & _381_ /*138*/;
assign _379_ = _298_ ^ _381_ /*141*/;
assign _380_ = _372_ & _379_ /*139*/;
assign _348_ = _372_ ^ _379_ /*140*/;
assign _377_ = _378_ | _380_ /*137*/;
assign _386_ = D[6] ^ Q[1] /*136*/;
assign _383_ = _299_ & _386_ /*132*/;
assign _384_ = _299_ ^ _386_ /*135*/;
assign _385_ = _377_ & _384_ /*133*/;
assign _349_ = _377_ ^ _384_ /*134*/;
assign _382_ = _383_ | _385_ /*131*/;
assign _390_ = zeroWire ^ Q[1] /*130*/;
assign _387_ = _300_ & _390_ /*126*/;
assign _388_ = _300_ ^ _390_ /*129*/;
assign _389_ = _382_ & _388_ /*127*/;
assign _350_ = _382_ ^ _388_ /*128*/;
assign Q[0] = _387_ | _389_ /*125*/;
assign _394_ = ~Q[0] /*74*/;
assign _393_ = _394_ & D[0] /*73*/;
assign _396_ = _343_ & _393_ /*68*/;
assign _397_ = _343_ ^ _393_ /*71*/;
assign _398_ = zeroWire & _397_ /*69*/;
assign R_n1[0] = zeroWire ^ _397_ /*70*/;
assign _395_ = _396_ | _398_ /*67*/;
assign _400_ = ~Q[0] /*66*/;
assign _399_ = _400_ & D[1] /*65*/;
assign _402_ = _344_ & _399_ /*60*/;
assign _403_ = _344_ ^ _399_ /*63*/;
assign _404_ = _395_ & _403_ /*61*/;
assign R_n1[1] = _395_ ^ _403_ /*62*/;
assign _401_ = _402_ | _404_ /*59*/;
assign _406_ = ~Q[0] /*58*/;
assign _405_ = _406_ & D[2] /*57*/;
assign _408_ = _345_ & _405_ /*52*/;
assign _409_ = _345_ ^ _405_ /*55*/;
assign _410_ = _401_ & _409_ /*53*/;
assign R_n1[2] = _401_ ^ _409_ /*54*/;
assign _407_ = _408_ | _410_ /*51*/;
assign _412_ = ~Q[0] /*50*/;
assign _411_ = _412_ & D[3] /*49*/;
assign _414_ = _346_ & _411_ /*44*/;
assign _415_ = _346_ ^ _411_ /*47*/;
assign _416_ = _407_ & _415_ /*45*/;
assign R_n1[3] = _407_ ^ _415_ /*46*/;
assign _413_ = _414_ | _416_ /*43*/;
assign _418_ = ~Q[0] /*42*/;
assign _417_ = _418_ & D[4] /*41*/;
assign _420_ = _347_ & _417_ /*36*/;
assign _421_ = _347_ ^ _417_ /*39*/;
assign _422_ = _413_ & _421_ /*37*/;
assign R_n1[4] = _413_ ^ _421_ /*38*/;
assign _419_ = _420_ | _422_ /*35*/;
assign _424_ = ~Q[0] /*34*/;
assign _423_ = _424_ & D[5] /*33*/;
assign _426_ = _348_ & _423_ /*28*/;
assign _427_ = _348_ ^ _423_ /*31*/;
assign _428_ = _419_ & _427_ /*29*/;
assign R_n1[5] = _419_ ^ _427_ /*30*/;
assign _425_ = _426_ | _428_ /*27*/;
assign _430_ = ~Q[0] /*26*/;
assign _429_ = _430_ & D[6] /*25*/;
assign _432_ = _349_ & _429_ /*20*/;
assign _433_ = _349_ ^ _429_ /*23*/;
assign _434_ = _425_ & _433_ /*21*/;
assign R_n1[6] = _425_ ^ _433_ /*22*/;
assign _431_ = _432_ | _434_ /*19*/;
endmodule
