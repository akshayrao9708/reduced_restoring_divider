module divider(Q, R_n1, R_0, D);
  wire _0_;
  wire _1_;
  wire _2_;
  wire _3_;
  wire _4_;
  wire _5_;
  wire _6_;
  wire _7_;
  wire _8_;
  wire _9_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  wire _38_;
  wire _39_;
  wire _40_;
  wire _41_;
  wire _42_;
  wire _43_;
  wire _44_;
  wire _45_;
  wire _46_;
  wire _47_;
  wire _48_;
  wire _49_;
  wire _50_;
  wire _51_;
  wire _52_;
  wire _53_;
  wire _54_;
  wire _55_;
  wire _56_;
  wire _57_;
  wire _58_;
  wire _59_;
  wire _60_;
  wire _61_;
  wire _62_;
  wire _63_;
  wire _64_;
  wire _65_;
  wire _66_;
  wire _67_;
  wire _68_;
  wire _69_;
  wire _70_;
  wire _71_;
  wire _72_;
  wire _73_;
  wire _74_;
  wire _75_;
  wire _76_;
  wire _77_;
  wire _78_;
  wire _79_;
  wire _80_;
  wire _81_;
  wire _82_;
  wire _83_;
  wire _84_;
  wire _85_;
  wire _86_;
  wire _87_;
  wire _88_;
  wire _89_;
  wire _90_;
  wire _91_;
  wire _92_;
  wire _93_;
  wire _94_;
  wire _95_;
  wire _96_;
  wire _97_;
  wire _98_;
  wire _99_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire _304_;
  wire _305_;
  wire _306_;
  wire _307_;
  wire _308_;
  wire _309_;
  wire _310_;
  wire _311_;
  wire _312_;
  wire _313_;
  wire _314_;
  wire _315_;
  wire _316_;
  wire _317_;
  wire _318_;
  wire _319_;
  wire _320_;
  wire _321_;
  wire _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire _326_;
  wire _327_;
  wire _328_;
  wire _329_;
  wire _330_;
  wire _331_;
  wire _332_;
  wire _333_;
  wire _334_;
  wire _335_;
  wire _336_;
  wire _337_;
  wire _338_;
  wire _339_;
  wire _340_;
  wire _341_;
  wire _342_;
  wire _343_;
  wire _344_;
  wire _345_;
  wire _346_;
  wire _347_;
  wire _348_;
  wire _349_;
  wire _350_;
  wire _351_;
  wire _352_;
  wire _353_;
  wire _354_;
  wire _355_;
  wire _356_;
  wire _357_;
  wire _358_;
  wire _359_;
  wire _360_;
  wire _361_;
  wire _362_;
  wire _363_;
  wire _364_;
  wire _365_;
  wire _366_;
  wire _367_;
  wire _368_;
  wire _369_;
  wire _370_;
  wire _371_;
  wire _372_;
  wire _373_;
  wire _374_;
  wire _375_;
  wire _376_;
  wire _377_;
  wire _378_;
  wire _379_;
  wire _380_;
  wire _381_;
  wire _382_;
  wire _383_;
  wire _384_;
  wire _385_;
  wire _386_;
  wire _387_;
  wire _388_;
  wire _389_;
  wire _390_;
  wire _391_;
  wire _392_;
  wire _393_;
  wire _394_;
  wire _395_;
  wire _396_;
  wire _397_;
  wire _398_;
  wire _399_;
  wire _400_;
  wire _401_;
  wire _402_;
  wire _403_;
  wire _404_;
  wire _405_;
  wire _406_;
  wire _407_;
  wire _408_;
  wire _409_;
  wire _410_;
  wire _411_;
  wire _412_;
  wire _413_;
  wire _414_;
  wire _415_;
  wire _416_;
  wire _417_;
  wire _418_;
  wire _419_;
  wire _420_;
  wire _421_;
  wire _422_;
  wire _423_;
  wire _424_;
  wire _425_;
  wire _426_;
  wire _427_;
  wire _428_;
  wire _429_;
  wire _430_;
  wire _431_;
  wire _432_;
  wire _433_;
  wire _434_;
  wire _435_;
  wire _436_;
  wire _437_;
  wire _438_;
  wire _439_;
  wire _440_;
  wire _441_;
  wire _442_;
  wire _443_;
  wire _444_;
  wire _445_;
  wire _446_;
  wire _447_;
  wire [14:0] r_0;
  wire [14:0] r_1;
  wire [7:0] m_1;
  wire [7:0] sum_1;
  wire [7:0] inv_1;
  wire [13:0] r_2;
  wire [7:0] m_2;
  wire [7:0] sum_2;
  wire [7:0] inv_2;
  wire [12:0] r_3;
  wire [7:0] m_3;
  wire [7:0] sum_3;
  wire [7:0] inv_3;
  wire [11:0] r_4;
  wire [7:0] m_4;
  wire [7:0] sum_4;
  wire [7:0] inv_4;
  wire [10:0] r_5;
  wire [7:0] m_5;
  wire [7:0] sum_5;
  wire [7:0] inv_5;
  wire [9:0] r_6;
  wire [7:0] m_6;
  wire [7:0] sum_6;
  wire [7:0] inv_6;
  wire [8:0] r_7;
  wire [7:0] m_7;
  wire [7:0] sum_7;
  wire [7:0] inv_7;
  wire [7:0] r_8;
  wire [7:0] m_8;
  wire [7:0] sum_8;
  wire [7:0] inv_8;
  wire zeroWire;
  wire oneWire;
  input [13:0] R_0;
  input [6:0] D;
  output [7:0] Q;
  output [7:0] R_n1;
  assign zeroWire = 1'b0 /*0*/;
  assign oneWire = 1'b1 /*0*/;
  assign r_0[0] = R_0[0] /*1199*/;
  assign r_0[1] = R_0[1] /*1198*/;
  assign r_0[2] = R_0[2] /*1197*/;
  assign r_0[3] = R_0[3] /*1196*/;
  assign r_0[4] = R_0[4] /*1195*/;
  assign r_0[5] = R_0[5] /*1194*/;
  assign r_0[6] = R_0[6] /*1193*/;
  assign r_0[7] = R_0[7] /*1192*/;
  assign r_0[8] = R_0[8] /*1191*/;
  assign r_0[9] = R_0[9] /*1190*/;
  assign r_0[10] = R_0[10] /*1189*/;
  assign r_0[11] = R_0[11] /*1188*/;
  assign r_0[12] = R_0[12] /*1187*/;
  assign r_0[13] = R_0[13] /*1186*/;
  assign r_0[14] = zeroWire /*1185*/;
  assign inv_1[0] = ~D[0] /*1184*/;
  assign inv_1[1] = ~D[1] /*1183*/;
  assign inv_1[2] = ~D[2] /*1182*/;
  assign inv_1[3] = ~D[3] /*1181*/;
  assign inv_1[4] = ~D[4] /*1180*/;
  assign inv_1[5] = ~D[5] /*1179*/;
  assign inv_1[6] = ~D[6] /*1178*/;
assign inv_1[7] = oneWire /*1177*/;
  assign _0_ = inv_1[0] ^ r_0[7] /*1175*/;
  assign sum_1[0] = _0_ ^ oneWire /*1174*/;
  assign _1_ = _0_ & oneWire /*1173*/;
  assign _2_ = inv_1[0] & r_0[7] /*1172*/;
  assign _3_ = _1_ | _2_ /*1171*/;
  assign _4_ = inv_1[1] ^ r_0[8] /*1169*/;
  assign sum_1[1] = _4_ ^ _3_ /*1168*/;
  assign _5_ = _4_ & _3_ /*1167*/;
  assign _6_ = inv_1[1] & r_0[8] /*1166*/;
  assign _7_ = _5_ | _6_ /*1165*/;
  assign _8_ = inv_1[2] ^ r_0[9] /*1164*/;
  assign sum_1[2] = _8_ ^ _7_ /*1163*/;
  assign _9_ = _8_ & _7_ /*1162*/;
  assign _10_ = inv_1[2] & r_0[9] /*1161*/;
  assign _11_ = _9_ | _10_ /*1160*/;
  assign _12_ = inv_1[3] ^ r_0[10] /*1159*/;
  assign sum_1[3] = _12_ ^ _11_ /*1158*/;
  assign _13_ = _12_ & _11_ /*1157*/;
  assign _14_ = inv_1[3] & r_0[10] /*1156*/;
  assign _15_ = _13_ | _14_ /*1155*/;
  assign _16_ = inv_1[4] ^ r_0[11] /*1154*/;
  assign sum_1[4] = _16_ ^ _15_ /*1153*/;
  assign _17_ = _16_ & _15_ /*1152*/;
  assign _18_ = inv_1[4] & r_0[11] /*1151*/;
  assign _19_ = _17_ | _18_ /*1150*/;
  assign _20_ = inv_1[5] ^ r_0[12] /*1149*/;
  assign sum_1[5] = _20_ ^ _19_ /*1148*/;
  assign _21_ = _20_ & _19_ /*1147*/;
  assign _22_ = inv_1[5] & r_0[12] /*1146*/;
  assign _23_ = _21_ | _22_ /*1145*/;
  assign _24_ = inv_1[6] ^ r_0[13] /*1144*/;
  assign sum_1[6] = _24_ ^ _23_ /*1143*/;
  assign _25_ = _24_ & _23_ /*1142*/;
  assign _26_ = inv_1[6] & r_0[13] /*1141*/;
  assign _27_ = _25_ | _26_ /*1140*/;
  assign _28_ = inv_1[7] ^ r_0[14] /*1139*/;
  assign sum_1[7] = _28_ ^ _27_ /*1138*/;
  assign _29_ = _28_ & _27_ /*1137*/;
  assign _30_ = inv_1[7] & r_0[14] /*1136*/;
  assign _31_ = _29_ | _30_ /*1135*/;
  assign Q[7] = ~sum_1[7] /*1133*/;
  assign m_1[0] = r_0[7] /*1132*/;
  assign m_1[1] = r_0[8] /*1131*/;
  assign m_1[2] = r_0[9] /*1130*/;
  assign m_1[3] = r_0[10] /*1129*/;
  assign m_1[4] = r_0[11] /*1128*/;
  assign m_1[5] = r_0[12] /*1127*/;
  assign m_1[6] = r_0[13] /*1126*/;
  assign m_1[7] = r_0[14] /*1125*/;
  assign _32_ = ~Q[7] /*1123*/;
  assign _33_ = sum_1[0] & Q[7] /*1122*/;
  assign _34_ = m_1[0] & _32_ /*1121*/;
  assign r_1[7] = _34_ | _33_ /*1120*/;
  assign _35_ = ~Q[7] /*1119*/;
  assign _36_ = sum_1[1] & Q[7] /*1118*/;
  assign _37_ = m_1[1] & _35_ /*1117*/;
  assign r_1[8] = _37_ | _36_ /*1116*/;
  assign _38_ = ~Q[7] /*1115*/;
  assign _39_ = sum_1[2] & Q[7] /*1114*/;
  assign _40_ = m_1[2] & _38_ /*1113*/;
  assign r_1[9] = _40_ | _39_ /*1112*/;
  assign _41_ = ~Q[7] /*1111*/;
  assign _42_ = sum_1[3] & Q[7] /*1110*/;
  assign _43_ = m_1[3] & _41_ /*1109*/;
  assign r_1[10] = _43_ | _42_ /*1108*/;
  assign _44_ = ~Q[7] /*1107*/;
  assign _45_ = sum_1[4] & Q[7] /*1106*/;
  assign _46_ = m_1[4] & _44_ /*1105*/;
  assign r_1[11] = _46_ | _45_ /*1104*/;
  assign _47_ = ~Q[7] /*1103*/;
  assign _48_ = sum_1[5] & Q[7] /*1102*/;
  assign _49_ = m_1[5] & _47_ /*1101*/;
  assign r_1[12] = _49_ | _48_ /*1100*/;
  assign _50_ = ~Q[7] /*1099*/;
  assign _51_ = sum_1[6] & Q[7] /*1098*/;
  assign _52_ = m_1[6] & _50_ /*1097*/;
  assign r_1[13] = _52_ | _51_ /*1096*/;
  assign _53_ = ~Q[7] /*1095*/;
  assign _54_ = sum_1[7] & Q[7] /*1094*/;
  assign _55_ = m_1[7] & _53_ /*1093*/;
  assign r_1[14] = _55_ | _54_ /*1092*/;
assign r_1[0]= r_0[0] /*1091*/;
assign r_1[1]= r_0[1] /*1090*/;
assign r_1[2]= r_0[2] /*1089*/;
assign r_1[3]= r_0[3] /*1088*/;
assign r_1[4]= r_0[4] /*1087*/;
assign r_1[5]= r_0[5] /*1086*/;
assign r_1[6]= r_0[6] /*1085*/;
  assign inv_2[0] = ~D[0] /*1072*/;
  assign inv_2[1] = ~D[1] /*1071*/;
  assign inv_2[2] = ~D[2] /*1070*/;
  assign inv_2[3] = ~D[3] /*1069*/;
  assign inv_2[4] = ~D[4] /*1068*/;
  assign inv_2[5] = ~D[5] /*1067*/;
  assign inv_2[6] = ~D[6] /*1066*/;
assign inv_2[7] = oneWire /*1065*/;
  assign _56_ = inv_2[0] ^ r_1[6] /*1063*/;
  assign sum_2[0] = _56_ ^ oneWire /*1062*/;
  assign _57_ = _56_ & oneWire /*1061*/;
  assign _58_ = inv_2[0] & r_1[6] /*1060*/;
  assign _59_ = _57_ | _58_ /*1059*/;
  assign _60_ = inv_2[1] ^ r_1[7] /*1057*/;
  assign sum_2[1] = _60_ ^ _59_ /*1056*/;
  assign _61_ = _60_ & _59_ /*1055*/;
  assign _62_ = inv_2[1] & r_1[7] /*1054*/;
  assign _63_ = _61_ | _62_ /*1053*/;
  assign _64_ = inv_2[2] ^ r_1[8] /*1052*/;
  assign sum_2[2] = _64_ ^ _63_ /*1051*/;
  assign _65_ = _64_ & _63_ /*1050*/;
  assign _66_ = inv_2[2] & r_1[8] /*1049*/;
  assign _67_ = _65_ | _66_ /*1048*/;
  assign _68_ = inv_2[3] ^ r_1[9] /*1047*/;
  assign sum_2[3] = _68_ ^ _67_ /*1046*/;
  assign _69_ = _68_ & _67_ /*1045*/;
  assign _70_ = inv_2[3] & r_1[9] /*1044*/;
  assign _71_ = _69_ | _70_ /*1043*/;
  assign _72_ = inv_2[4] ^ r_1[10] /*1042*/;
  assign sum_2[4] = _72_ ^ _71_ /*1041*/;
  assign _73_ = _72_ & _71_ /*1040*/;
  assign _74_ = inv_2[4] & r_1[10] /*1039*/;
  assign _75_ = _73_ | _74_ /*1038*/;
  assign _76_ = inv_2[5] ^ r_1[11] /*1037*/;
  assign sum_2[5] = _76_ ^ _75_ /*1036*/;
  assign _77_ = _76_ & _75_ /*1035*/;
  assign _78_ = inv_2[5] & r_1[11] /*1034*/;
  assign _79_ = _77_ | _78_ /*1033*/;
  assign _80_ = inv_2[6] ^ r_1[12] /*1032*/;
  assign sum_2[6] = _80_ ^ _79_ /*1031*/;
  assign _81_ = _80_ & _79_ /*1030*/;
  assign _82_ = inv_2[6] & r_1[12] /*1029*/;
  assign _83_ = _81_ | _82_ /*1028*/;
  assign _84_ = inv_2[7] ^ r_1[13] /*1027*/;
  assign sum_2[7] = _84_ ^ _83_ /*1026*/;
  assign _85_ = _84_ & _83_ /*1025*/;
  assign _86_ = inv_2[7] & r_1[13] /*1024*/;
  assign _87_ = _85_ | _86_ /*1023*/;
  assign Q[6] = ~sum_2[7] /*1021*/;
  assign m_2[0] = r_1[6] /*1020*/;
  assign m_2[1] = r_1[7] /*1019*/;
  assign m_2[2] = r_1[8] /*1018*/;
  assign m_2[3] = r_1[9] /*1017*/;
  assign m_2[4] = r_1[10] /*1016*/;
  assign m_2[5] = r_1[11] /*1015*/;
  assign m_2[6] = r_1[12] /*1014*/;
  assign m_2[7] = r_1[13] /*1013*/;
  assign _88_ = ~Q[6] /*1011*/;
  assign _89_ = sum_2[0] & Q[6] /*1010*/;
  assign _90_ = m_2[0] & _88_ /*1009*/;
  assign r_2[6] = _90_ | _89_ /*1008*/;
  assign _91_ = ~Q[6] /*1007*/;
  assign _92_ = sum_2[1] & Q[6] /*1006*/;
  assign _93_ = m_2[1] & _91_ /*1005*/;
  assign r_2[7] = _93_ | _92_ /*1004*/;
  assign _94_ = ~Q[6] /*1003*/;
  assign _95_ = sum_2[2] & Q[6] /*1002*/;
  assign _96_ = m_2[2] & _94_ /*1001*/;
  assign r_2[8] = _96_ | _95_ /*1000*/;
  assign _97_ = ~Q[6] /*999*/;
  assign _98_ = sum_2[3] & Q[6] /*998*/;
  assign _99_ = m_2[3] & _97_ /*997*/;
  assign r_2[9] = _99_ | _98_ /*996*/;
  assign _100_ = ~Q[6] /*995*/;
  assign _101_ = sum_2[4] & Q[6] /*994*/;
  assign _102_ = m_2[4] & _100_ /*993*/;
  assign r_2[10] = _102_ | _101_ /*992*/;
  assign _103_ = ~Q[6] /*991*/;
  assign _104_ = sum_2[5] & Q[6] /*990*/;
  assign _105_ = m_2[5] & _103_ /*989*/;
  assign r_2[11] = _105_ | _104_ /*988*/;
  assign _106_ = ~Q[6] /*987*/;
  assign _107_ = sum_2[6] & Q[6] /*986*/;
  assign _108_ = m_2[6] & _106_ /*985*/;
  assign r_2[12] = _108_ | _107_ /*984*/;
  assign _109_ = ~Q[6] /*983*/;
  assign _110_ = sum_2[7] & Q[6] /*982*/;
  assign _111_ = m_2[7] & _109_ /*981*/;
  assign r_2[13] = _111_ | _110_ /*980*/;
assign r_2[0]= r_1[0] /*979*/;
assign r_2[1]= r_1[1] /*978*/;
assign r_2[2]= r_1[2] /*977*/;
assign r_2[3]= r_1[3] /*976*/;
assign r_2[4]= r_1[4] /*975*/;
assign r_2[5]= r_1[5] /*974*/;
  assign inv_3[0] = ~D[0] /*960*/;
  assign inv_3[1] = ~D[1] /*959*/;
  assign inv_3[2] = ~D[2] /*958*/;
  assign inv_3[3] = ~D[3] /*957*/;
  assign inv_3[4] = ~D[4] /*956*/;
  assign inv_3[5] = ~D[5] /*955*/;
  assign inv_3[6] = ~D[6] /*954*/;
assign inv_3[7] = oneWire /*953*/;
  assign _112_ = inv_3[0] ^ r_2[5] /*951*/;
  assign sum_3[0] = _112_ ^ oneWire /*950*/;
  assign _113_ = _112_ & oneWire /*949*/;
  assign _114_ = inv_3[0] & r_2[5] /*948*/;
  assign _115_ = _113_ | _114_ /*947*/;
  assign _116_ = inv_3[1] ^ r_2[6] /*945*/;
  assign sum_3[1] = _116_ ^ _115_ /*944*/;
  assign _117_ = _116_ & _115_ /*943*/;
  assign _118_ = inv_3[1] & r_2[6] /*942*/;
  assign _119_ = _117_ | _118_ /*941*/;
  assign _120_ = inv_3[2] ^ r_2[7] /*940*/;
  assign sum_3[2] = _120_ ^ _119_ /*939*/;
  assign _121_ = _120_ & _119_ /*938*/;
  assign _122_ = inv_3[2] & r_2[7] /*937*/;
  assign _123_ = _121_ | _122_ /*936*/;
  assign _124_ = inv_3[3] ^ r_2[8] /*935*/;
  assign sum_3[3] = _124_ ^ _123_ /*934*/;
  assign _125_ = _124_ & _123_ /*933*/;
  assign _126_ = inv_3[3] & r_2[8] /*932*/;
  assign _127_ = _125_ | _126_ /*931*/;
  assign _128_ = inv_3[4] ^ r_2[9] /*930*/;
  assign sum_3[4] = _128_ ^ _127_ /*929*/;
  assign _129_ = _128_ & _127_ /*928*/;
  assign _130_ = inv_3[4] & r_2[9] /*927*/;
  assign _131_ = _129_ | _130_ /*926*/;
  assign _132_ = inv_3[5] ^ r_2[10] /*925*/;
  assign sum_3[5] = _132_ ^ _131_ /*924*/;
  assign _133_ = _132_ & _131_ /*923*/;
  assign _134_ = inv_3[5] & r_2[10] /*922*/;
  assign _135_ = _133_ | _134_ /*921*/;
  assign _136_ = inv_3[6] ^ r_2[11] /*920*/;
  assign sum_3[6] = _136_ ^ _135_ /*919*/;
  assign _137_ = _136_ & _135_ /*918*/;
  assign _138_ = inv_3[6] & r_2[11] /*917*/;
  assign _139_ = _137_ | _138_ /*916*/;
  assign _140_ = inv_3[7] ^ r_2[12] /*915*/;
  assign sum_3[7] = _140_ ^ _139_ /*914*/;
  assign _141_ = _140_ & _139_ /*913*/;
  assign _142_ = inv_3[7] & r_2[12] /*912*/;
  assign _143_ = _141_ | _142_ /*911*/;
  assign Q[5] = ~sum_3[7] /*909*/;
  assign m_3[0] = r_2[5] /*908*/;
  assign m_3[1] = r_2[6] /*907*/;
  assign m_3[2] = r_2[7] /*906*/;
  assign m_3[3] = r_2[8] /*905*/;
  assign m_3[4] = r_2[9] /*904*/;
  assign m_3[5] = r_2[10] /*903*/;
  assign m_3[6] = r_2[11] /*902*/;
  assign m_3[7] = r_2[12] /*901*/;
  assign _144_ = ~Q[5] /*899*/;
  assign _145_ = sum_3[0] & Q[5] /*898*/;
  assign _146_ = m_3[0] & _144_ /*897*/;
  assign r_3[5] = _146_ | _145_ /*896*/;
  assign _147_ = ~Q[5] /*895*/;
  assign _148_ = sum_3[1] & Q[5] /*894*/;
  assign _149_ = m_3[1] & _147_ /*893*/;
  assign r_3[6] = _149_ | _148_ /*892*/;
  assign _150_ = ~Q[5] /*891*/;
  assign _151_ = sum_3[2] & Q[5] /*890*/;
  assign _152_ = m_3[2] & _150_ /*889*/;
  assign r_3[7] = _152_ | _151_ /*888*/;
  assign _153_ = ~Q[5] /*887*/;
  assign _154_ = sum_3[3] & Q[5] /*886*/;
  assign _155_ = m_3[3] & _153_ /*885*/;
  assign r_3[8] = _155_ | _154_ /*884*/;
  assign _156_ = ~Q[5] /*883*/;
  assign _157_ = sum_3[4] & Q[5] /*882*/;
  assign _158_ = m_3[4] & _156_ /*881*/;
  assign r_3[9] = _158_ | _157_ /*880*/;
  assign _159_ = ~Q[5] /*879*/;
  assign _160_ = sum_3[5] & Q[5] /*878*/;
  assign _161_ = m_3[5] & _159_ /*877*/;
  assign r_3[10] = _161_ | _160_ /*876*/;
  assign _162_ = ~Q[5] /*875*/;
  assign _163_ = sum_3[6] & Q[5] /*874*/;
  assign _164_ = m_3[6] & _162_ /*873*/;
  assign r_3[11] = _164_ | _163_ /*872*/;
  assign _165_ = ~Q[5] /*871*/;
  assign _166_ = sum_3[7] & Q[5] /*870*/;
  assign _167_ = m_3[7] & _165_ /*869*/;
  assign r_3[12] = _167_ | _166_ /*868*/;
assign r_3[0]= r_2[0] /*867*/;
assign r_3[1]= r_2[1] /*866*/;
assign r_3[2]= r_2[2] /*865*/;
assign r_3[3]= r_2[3] /*864*/;
assign r_3[4]= r_2[4] /*863*/;
  assign inv_4[0] = ~D[0] /*848*/;
  assign inv_4[1] = ~D[1] /*847*/;
  assign inv_4[2] = ~D[2] /*846*/;
  assign inv_4[3] = ~D[3] /*845*/;
  assign inv_4[4] = ~D[4] /*844*/;
  assign inv_4[5] = ~D[5] /*843*/;
  assign inv_4[6] = ~D[6] /*842*/;
assign inv_4[7] = oneWire /*841*/;
  assign _168_ = inv_4[0] ^ r_3[4] /*839*/;
  assign sum_4[0] = _168_ ^ oneWire /*838*/;
  assign _169_ = _168_ & oneWire /*837*/;
  assign _170_ = inv_4[0] & r_3[4] /*836*/;
  assign _171_ = _169_ | _170_ /*835*/;
  assign _172_ = inv_4[1] ^ r_3[5] /*833*/;
  assign sum_4[1] = _172_ ^ _171_ /*832*/;
  assign _173_ = _172_ & _171_ /*831*/;
  assign _174_ = inv_4[1] & r_3[5] /*830*/;
  assign _175_ = _173_ | _174_ /*829*/;
  assign _176_ = inv_4[2] ^ r_3[6] /*828*/;
  assign sum_4[2] = _176_ ^ _175_ /*827*/;
  assign _177_ = _176_ & _175_ /*826*/;
  assign _178_ = inv_4[2] & r_3[6] /*825*/;
  assign _179_ = _177_ | _178_ /*824*/;
  assign _180_ = inv_4[3] ^ r_3[7] /*823*/;
  assign sum_4[3] = _180_ ^ _179_ /*822*/;
  assign _181_ = _180_ & _179_ /*821*/;
  assign _182_ = inv_4[3] & r_3[7] /*820*/;
  assign _183_ = _181_ | _182_ /*819*/;
  assign _184_ = inv_4[4] ^ r_3[8] /*818*/;
  assign sum_4[4] = _184_ ^ _183_ /*817*/;
  assign _185_ = _184_ & _183_ /*816*/;
  assign _186_ = inv_4[4] & r_3[8] /*815*/;
  assign _187_ = _185_ | _186_ /*814*/;
  assign _188_ = inv_4[5] ^ r_3[9] /*813*/;
  assign sum_4[5] = _188_ ^ _187_ /*812*/;
  assign _189_ = _188_ & _187_ /*811*/;
  assign _190_ = inv_4[5] & r_3[9] /*810*/;
  assign _191_ = _189_ | _190_ /*809*/;
  assign _192_ = inv_4[6] ^ r_3[10] /*808*/;
  assign sum_4[6] = _192_ ^ _191_ /*807*/;
  assign _193_ = _192_ & _191_ /*806*/;
  assign _194_ = inv_4[6] & r_3[10] /*805*/;
  assign _195_ = _193_ | _194_ /*804*/;
  assign _196_ = inv_4[7] ^ r_3[11] /*803*/;
  assign sum_4[7] = _196_ ^ _195_ /*802*/;
  assign _197_ = _196_ & _195_ /*801*/;
  assign _198_ = inv_4[7] & r_3[11] /*800*/;
  assign _199_ = _197_ | _198_ /*799*/;
  assign Q[4] = ~sum_4[7] /*797*/;
  assign m_4[0] = r_3[4] /*796*/;
  assign m_4[1] = r_3[5] /*795*/;
  assign m_4[2] = r_3[6] /*794*/;
  assign m_4[3] = r_3[7] /*793*/;
  assign m_4[4] = r_3[8] /*792*/;
  assign m_4[5] = r_3[9] /*791*/;
  assign m_4[6] = r_3[10] /*790*/;
  assign m_4[7] = r_3[11] /*789*/;
  assign _200_ = ~Q[4] /*787*/;
  assign _201_ = sum_4[0] & Q[4] /*786*/;
  assign _202_ = m_4[0] & _200_ /*785*/;
  assign r_4[4] = _202_ | _201_ /*784*/;
  assign _203_ = ~Q[4] /*783*/;
  assign _204_ = sum_4[1] & Q[4] /*782*/;
  assign _205_ = m_4[1] & _203_ /*781*/;
  assign r_4[5] = _205_ | _204_ /*780*/;
  assign _206_ = ~Q[4] /*779*/;
  assign _207_ = sum_4[2] & Q[4] /*778*/;
  assign _208_ = m_4[2] & _206_ /*777*/;
  assign r_4[6] = _208_ | _207_ /*776*/;
  assign _209_ = ~Q[4] /*775*/;
  assign _210_ = sum_4[3] & Q[4] /*774*/;
  assign _211_ = m_4[3] & _209_ /*773*/;
  assign r_4[7] = _211_ | _210_ /*772*/;
  assign _212_ = ~Q[4] /*771*/;
  assign _213_ = sum_4[4] & Q[4] /*770*/;
  assign _214_ = m_4[4] & _212_ /*769*/;
  assign r_4[8] = _214_ | _213_ /*768*/;
  assign _215_ = ~Q[4] /*767*/;
  assign _216_ = sum_4[5] & Q[4] /*766*/;
  assign _217_ = m_4[5] & _215_ /*765*/;
  assign r_4[9] = _217_ | _216_ /*764*/;
  assign _218_ = ~Q[4] /*763*/;
  assign _219_ = sum_4[6] & Q[4] /*762*/;
  assign _220_ = m_4[6] & _218_ /*761*/;
  assign r_4[10] = _220_ | _219_ /*760*/;
  assign _221_ = ~Q[4] /*759*/;
  assign _222_ = sum_4[7] & Q[4] /*758*/;
  assign _223_ = m_4[7] & _221_ /*757*/;
  assign r_4[11] = _223_ | _222_ /*756*/;
assign r_4[0]= r_3[0] /*755*/;
assign r_4[1]= r_3[1] /*754*/;
assign r_4[2]= r_3[2] /*753*/;
assign r_4[3]= r_3[3] /*752*/;
  assign inv_5[0] = ~D[0] /*736*/;
  assign inv_5[1] = ~D[1] /*735*/;
  assign inv_5[2] = ~D[2] /*734*/;
  assign inv_5[3] = ~D[3] /*733*/;
  assign inv_5[4] = ~D[4] /*732*/;
  assign inv_5[5] = ~D[5] /*731*/;
  assign inv_5[6] = ~D[6] /*730*/;
assign inv_5[7] = oneWire /*729*/;
  assign _224_ = inv_5[0] ^ r_4[3] /*727*/;
  assign sum_5[0] = _224_ ^ oneWire /*726*/;
  assign _225_ = _224_ & oneWire /*725*/;
  assign _226_ = inv_5[0] & r_4[3] /*724*/;
  assign _227_ = _225_ | _226_ /*723*/;
  assign _228_ = inv_5[1] ^ r_4[4] /*721*/;
  assign sum_5[1] = _228_ ^ _227_ /*720*/;
  assign _229_ = _228_ & _227_ /*719*/;
  assign _230_ = inv_5[1] & r_4[4] /*718*/;
  assign _231_ = _229_ | _230_ /*717*/;
  assign _232_ = inv_5[2] ^ r_4[5] /*716*/;
  assign sum_5[2] = _232_ ^ _231_ /*715*/;
  assign _233_ = _232_ & _231_ /*714*/;
  assign _234_ = inv_5[2] & r_4[5] /*713*/;
  assign _235_ = _233_ | _234_ /*712*/;
  assign _236_ = inv_5[3] ^ r_4[6] /*711*/;
  assign sum_5[3] = _236_ ^ _235_ /*710*/;
  assign _237_ = _236_ & _235_ /*709*/;
  assign _238_ = inv_5[3] & r_4[6] /*708*/;
  assign _239_ = _237_ | _238_ /*707*/;
  assign _240_ = inv_5[4] ^ r_4[7] /*706*/;
  assign sum_5[4] = _240_ ^ _239_ /*705*/;
  assign _241_ = _240_ & _239_ /*704*/;
  assign _242_ = inv_5[4] & r_4[7] /*703*/;
  assign _243_ = _241_ | _242_ /*702*/;
  assign _244_ = inv_5[5] ^ r_4[8] /*701*/;
  assign sum_5[5] = _244_ ^ _243_ /*700*/;
  assign _245_ = _244_ & _243_ /*699*/;
  assign _246_ = inv_5[5] & r_4[8] /*698*/;
  assign _247_ = _245_ | _246_ /*697*/;
  assign _248_ = inv_5[6] ^ r_4[9] /*696*/;
  assign sum_5[6] = _248_ ^ _247_ /*695*/;
  assign _249_ = _248_ & _247_ /*694*/;
  assign _250_ = inv_5[6] & r_4[9] /*693*/;
  assign _251_ = _249_ | _250_ /*692*/;
  assign _252_ = inv_5[7] ^ r_4[10] /*691*/;
  assign sum_5[7] = _252_ ^ _251_ /*690*/;
  assign _253_ = _252_ & _251_ /*689*/;
  assign _254_ = inv_5[7] & r_4[10] /*688*/;
  assign _255_ = _253_ | _254_ /*687*/;
  assign Q[3] = ~sum_5[7] /*685*/;
  assign m_5[0] = r_4[3] /*684*/;
  assign m_5[1] = r_4[4] /*683*/;
  assign m_5[2] = r_4[5] /*682*/;
  assign m_5[3] = r_4[6] /*681*/;
  assign m_5[4] = r_4[7] /*680*/;
  assign m_5[5] = r_4[8] /*679*/;
  assign m_5[6] = r_4[9] /*678*/;
  assign m_5[7] = r_4[10] /*677*/;
  assign _256_ = ~Q[3] /*675*/;
  assign _257_ = sum_5[0] & Q[3] /*674*/;
  assign _258_ = m_5[0] & _256_ /*673*/;
  assign r_5[3] = _258_ | _257_ /*672*/;
  assign _259_ = ~Q[3] /*671*/;
  assign _260_ = sum_5[1] & Q[3] /*670*/;
  assign _261_ = m_5[1] & _259_ /*669*/;
  assign r_5[4] = _261_ | _260_ /*668*/;
  assign _262_ = ~Q[3] /*667*/;
  assign _263_ = sum_5[2] & Q[3] /*666*/;
  assign _264_ = m_5[2] & _262_ /*665*/;
  assign r_5[5] = _264_ | _263_ /*664*/;
  assign _265_ = ~Q[3] /*663*/;
  assign _266_ = sum_5[3] & Q[3] /*662*/;
  assign _267_ = m_5[3] & _265_ /*661*/;
  assign r_5[6] = _267_ | _266_ /*660*/;
  assign _268_ = ~Q[3] /*659*/;
  assign _269_ = sum_5[4] & Q[3] /*658*/;
  assign _270_ = m_5[4] & _268_ /*657*/;
  assign r_5[7] = _270_ | _269_ /*656*/;
  assign _271_ = ~Q[3] /*655*/;
  assign _272_ = sum_5[5] & Q[3] /*654*/;
  assign _273_ = m_5[5] & _271_ /*653*/;
  assign r_5[8] = _273_ | _272_ /*652*/;
  assign _274_ = ~Q[3] /*651*/;
  assign _275_ = sum_5[6] & Q[3] /*650*/;
  assign _276_ = m_5[6] & _274_ /*649*/;
  assign r_5[9] = _276_ | _275_ /*648*/;
  assign _277_ = ~Q[3] /*647*/;
  assign _278_ = sum_5[7] & Q[3] /*646*/;
  assign _279_ = m_5[7] & _277_ /*645*/;
  assign r_5[10] = _279_ | _278_ /*644*/;
assign r_5[0]= r_4[0] /*643*/;
assign r_5[1]= r_4[1] /*642*/;
assign r_5[2]= r_4[2] /*641*/;
  assign inv_6[0] = ~D[0] /*624*/;
  assign inv_6[1] = ~D[1] /*623*/;
  assign inv_6[2] = ~D[2] /*622*/;
  assign inv_6[3] = ~D[3] /*621*/;
  assign inv_6[4] = ~D[4] /*620*/;
  assign inv_6[5] = ~D[5] /*619*/;
  assign inv_6[6] = ~D[6] /*618*/;
assign inv_6[7] = oneWire /*617*/;
  assign _280_ = inv_6[0] ^ r_5[2] /*615*/;
  assign sum_6[0] = _280_ ^ oneWire /*614*/;
  assign _281_ = _280_ & oneWire /*613*/;
  assign _282_ = inv_6[0] & r_5[2] /*612*/;
  assign _283_ = _281_ | _282_ /*611*/;
  assign _284_ = inv_6[1] ^ r_5[3] /*609*/;
  assign sum_6[1] = _284_ ^ _283_ /*608*/;
  assign _285_ = _284_ & _283_ /*607*/;
  assign _286_ = inv_6[1] & r_5[3] /*606*/;
  assign _287_ = _285_ | _286_ /*605*/;
  assign _288_ = inv_6[2] ^ r_5[4] /*604*/;
  assign sum_6[2] = _288_ ^ _287_ /*603*/;
  assign _289_ = _288_ & _287_ /*602*/;
  assign _290_ = inv_6[2] & r_5[4] /*601*/;
  assign _291_ = _289_ | _290_ /*600*/;
  assign _292_ = inv_6[3] ^ r_5[5] /*599*/;
  assign sum_6[3] = _292_ ^ _291_ /*598*/;
  assign _293_ = _292_ & _291_ /*597*/;
  assign _294_ = inv_6[3] & r_5[5] /*596*/;
  assign _295_ = _293_ | _294_ /*595*/;
  assign _296_ = inv_6[4] ^ r_5[6] /*594*/;
  assign sum_6[4] = _296_ ^ _295_ /*593*/;
  assign _297_ = _296_ & _295_ /*592*/;
  assign _298_ = inv_6[4] & r_5[6] /*591*/;
  assign _299_ = _297_ | _298_ /*590*/;
  assign _300_ = inv_6[5] ^ r_5[7] /*589*/;
  assign sum_6[5] = _300_ ^ _299_ /*588*/;
  assign _301_ = _300_ & _299_ /*587*/;
  assign _302_ = inv_6[5] & r_5[7] /*586*/;
  assign _303_ = _301_ | _302_ /*585*/;
  assign _304_ = inv_6[6] ^ r_5[8] /*584*/;
  assign sum_6[6] = _304_ ^ _303_ /*583*/;
  assign _305_ = _304_ & _303_ /*582*/;
  assign _306_ = inv_6[6] & r_5[8] /*581*/;
  assign _307_ = _305_ | _306_ /*580*/;
  assign _308_ = inv_6[7] ^ r_5[9] /*579*/;
  assign sum_6[7] = _308_ ^ _307_ /*578*/;
  assign _309_ = _308_ & _307_ /*577*/;
  assign _310_ = inv_6[7] & r_5[9] /*576*/;
  assign _311_ = _309_ | _310_ /*575*/;
  assign Q[2] = ~sum_6[7] /*573*/;
  assign m_6[0] = r_5[2] /*572*/;
  assign m_6[1] = r_5[3] /*571*/;
  assign m_6[2] = r_5[4] /*570*/;
  assign m_6[3] = r_5[5] /*569*/;
  assign m_6[4] = r_5[6] /*568*/;
  assign m_6[5] = r_5[7] /*567*/;
  assign m_6[6] = r_5[8] /*566*/;
  assign m_6[7] = r_5[9] /*565*/;
  assign _312_ = ~Q[2] /*563*/;
  assign _313_ = sum_6[0] & Q[2] /*562*/;
  assign _314_ = m_6[0] & _312_ /*561*/;
  assign r_6[2] = _314_ | _313_ /*560*/;
  assign _315_ = ~Q[2] /*559*/;
  assign _316_ = sum_6[1] & Q[2] /*558*/;
  assign _317_ = m_6[1] & _315_ /*557*/;
  assign r_6[3] = _317_ | _316_ /*556*/;
  assign _318_ = ~Q[2] /*555*/;
  assign _319_ = sum_6[2] & Q[2] /*554*/;
  assign _320_ = m_6[2] & _318_ /*553*/;
  assign r_6[4] = _320_ | _319_ /*552*/;
  assign _321_ = ~Q[2] /*551*/;
  assign _322_ = sum_6[3] & Q[2] /*550*/;
  assign _323_ = m_6[3] & _321_ /*549*/;
  assign r_6[5] = _323_ | _322_ /*548*/;
  assign _324_ = ~Q[2] /*547*/;
  assign _325_ = sum_6[4] & Q[2] /*546*/;
  assign _326_ = m_6[4] & _324_ /*545*/;
  assign r_6[6] = _326_ | _325_ /*544*/;
  assign _327_ = ~Q[2] /*543*/;
  assign _328_ = sum_6[5] & Q[2] /*542*/;
  assign _329_ = m_6[5] & _327_ /*541*/;
  assign r_6[7] = _329_ | _328_ /*540*/;
  assign _330_ = ~Q[2] /*539*/;
  assign _331_ = sum_6[6] & Q[2] /*538*/;
  assign _332_ = m_6[6] & _330_ /*537*/;
  assign r_6[8] = _332_ | _331_ /*536*/;
  assign _333_ = ~Q[2] /*535*/;
  assign _334_ = sum_6[7] & Q[2] /*534*/;
  assign _335_ = m_6[7] & _333_ /*533*/;
  assign r_6[9] = _335_ | _334_ /*532*/;
assign r_6[0]= r_5[0] /*531*/;
assign r_6[1]= r_5[1] /*530*/;
  assign inv_7[0] = ~D[0] /*512*/;
  assign inv_7[1] = ~D[1] /*511*/;
  assign inv_7[2] = ~D[2] /*510*/;
  assign inv_7[3] = ~D[3] /*509*/;
  assign inv_7[4] = ~D[4] /*508*/;
  assign inv_7[5] = ~D[5] /*507*/;
  assign inv_7[6] = ~D[6] /*506*/;
assign inv_7[7] = oneWire /*505*/;
  assign _336_ = inv_7[0] ^ r_6[1] /*503*/;
  assign sum_7[0] = _336_ ^ oneWire /*502*/;
  assign _337_ = _336_ & oneWire /*501*/;
  assign _338_ = inv_7[0] & r_6[1] /*500*/;
  assign _339_ = _337_ | _338_ /*499*/;
  assign _340_ = inv_7[1] ^ r_6[2] /*497*/;
  assign sum_7[1] = _340_ ^ _339_ /*496*/;
  assign _341_ = _340_ & _339_ /*495*/;
  assign _342_ = inv_7[1] & r_6[2] /*494*/;
  assign _343_ = _341_ | _342_ /*493*/;
  assign _344_ = inv_7[2] ^ r_6[3] /*492*/;
  assign sum_7[2] = _344_ ^ _343_ /*491*/;
  assign _345_ = _344_ & _343_ /*490*/;
  assign _346_ = inv_7[2] & r_6[3] /*489*/;
  assign _347_ = _345_ | _346_ /*488*/;
  assign _348_ = inv_7[3] ^ r_6[4] /*487*/;
  assign sum_7[3] = _348_ ^ _347_ /*486*/;
  assign _349_ = _348_ & _347_ /*485*/;
  assign _350_ = inv_7[3] & r_6[4] /*484*/;
  assign _351_ = _349_ | _350_ /*483*/;
  assign _352_ = inv_7[4] ^ r_6[5] /*482*/;
  assign sum_7[4] = _352_ ^ _351_ /*481*/;
  assign _353_ = _352_ & _351_ /*480*/;
  assign _354_ = inv_7[4] & r_6[5] /*479*/;
  assign _355_ = _353_ | _354_ /*478*/;
  assign _356_ = inv_7[5] ^ r_6[6] /*477*/;
  assign sum_7[5] = _356_ ^ _355_ /*476*/;
  assign _357_ = _356_ & _355_ /*475*/;
  assign _358_ = inv_7[5] & r_6[6] /*474*/;
  assign _359_ = _357_ | _358_ /*473*/;
  assign _360_ = inv_7[6] ^ r_6[7] /*472*/;
  assign sum_7[6] = _360_ ^ _359_ /*471*/;
  assign _361_ = _360_ & _359_ /*470*/;
  assign _362_ = inv_7[6] & r_6[7] /*469*/;
  assign _363_ = _361_ | _362_ /*468*/;
  assign _364_ = inv_7[7] ^ r_6[8] /*467*/;
  assign sum_7[7] = _364_ ^ _363_ /*466*/;
  assign _365_ = _364_ & _363_ /*465*/;
  assign _366_ = inv_7[7] & r_6[8] /*464*/;
  assign _367_ = _365_ | _366_ /*463*/;
  assign Q[1] = ~sum_7[7] /*461*/;
  assign m_7[0] = r_6[1] /*460*/;
  assign m_7[1] = r_6[2] /*459*/;
  assign m_7[2] = r_6[3] /*458*/;
  assign m_7[3] = r_6[4] /*457*/;
  assign m_7[4] = r_6[5] /*456*/;
  assign m_7[5] = r_6[6] /*455*/;
  assign m_7[6] = r_6[7] /*454*/;
  assign m_7[7] = r_6[8] /*453*/;
  assign _368_ = ~Q[1] /*451*/;
  assign _369_ = sum_7[0] & Q[1] /*450*/;
  assign _370_ = m_7[0] & _368_ /*449*/;
  assign r_7[1] = _370_ | _369_ /*448*/;
  assign _371_ = ~Q[1] /*447*/;
  assign _372_ = sum_7[1] & Q[1] /*446*/;
  assign _373_ = m_7[1] & _371_ /*445*/;
  assign r_7[2] = _373_ | _372_ /*444*/;
  assign _374_ = ~Q[1] /*443*/;
  assign _375_ = sum_7[2] & Q[1] /*442*/;
  assign _376_ = m_7[2] & _374_ /*441*/;
  assign r_7[3] = _376_ | _375_ /*440*/;
  assign _377_ = ~Q[1] /*439*/;
  assign _378_ = sum_7[3] & Q[1] /*438*/;
  assign _379_ = m_7[3] & _377_ /*437*/;
  assign r_7[4] = _379_ | _378_ /*436*/;
  assign _380_ = ~Q[1] /*435*/;
  assign _381_ = sum_7[4] & Q[1] /*434*/;
  assign _382_ = m_7[4] & _380_ /*433*/;
  assign r_7[5] = _382_ | _381_ /*432*/;
  assign _383_ = ~Q[1] /*431*/;
  assign _384_ = sum_7[5] & Q[1] /*430*/;
  assign _385_ = m_7[5] & _383_ /*429*/;
  assign r_7[6] = _385_ | _384_ /*428*/;
  assign _386_ = ~Q[1] /*427*/;
  assign _387_ = sum_7[6] & Q[1] /*426*/;
  assign _388_ = m_7[6] & _386_ /*425*/;
  assign r_7[7] = _388_ | _387_ /*424*/;
  assign _389_ = ~Q[1] /*423*/;
  assign _390_ = sum_7[7] & Q[1] /*422*/;
  assign _391_ = m_7[7] & _389_ /*421*/;
  assign r_7[8] = _391_ | _390_ /*420*/;
assign r_7[0]= r_6[0] /*419*/;
  assign inv_8[0] = ~D[0] /*400*/;
  assign inv_8[1] = ~D[1] /*399*/;
  assign inv_8[2] = ~D[2] /*398*/;
  assign inv_8[3] = ~D[3] /*397*/;
  assign inv_8[4] = ~D[4] /*396*/;
  assign inv_8[5] = ~D[5] /*395*/;
  assign inv_8[6] = ~D[6] /*394*/;
assign inv_8[7] = oneWire /*393*/;
  assign _392_ = inv_8[0] ^ r_7[0] /*391*/;
  assign sum_8[0] = _392_ ^ oneWire /*390*/;
  assign _393_ = _392_ & oneWire /*389*/;
  assign _394_ = inv_8[0] & r_7[0] /*388*/;
  assign _395_ = _393_ | _394_ /*387*/;
  assign _396_ = inv_8[1] ^ r_7[1] /*385*/;
  assign sum_8[1] = _396_ ^ _395_ /*384*/;
  assign _397_ = _396_ & _395_ /*383*/;
  assign _398_ = inv_8[1] & r_7[1] /*382*/;
  assign _399_ = _397_ | _398_ /*381*/;
  assign _400_ = inv_8[2] ^ r_7[2] /*380*/;
  assign sum_8[2] = _400_ ^ _399_ /*379*/;
  assign _401_ = _400_ & _399_ /*378*/;
  assign _402_ = inv_8[2] & r_7[2] /*377*/;
  assign _403_ = _401_ | _402_ /*376*/;
  assign _404_ = inv_8[3] ^ r_7[3] /*375*/;
  assign sum_8[3] = _404_ ^ _403_ /*374*/;
  assign _405_ = _404_ & _403_ /*373*/;
  assign _406_ = inv_8[3] & r_7[3] /*372*/;
  assign _407_ = _405_ | _406_ /*371*/;
  assign _408_ = inv_8[4] ^ r_7[4] /*370*/;
  assign sum_8[4] = _408_ ^ _407_ /*369*/;
  assign _409_ = _408_ & _407_ /*368*/;
  assign _410_ = inv_8[4] & r_7[4] /*367*/;
  assign _411_ = _409_ | _410_ /*366*/;
  assign _412_ = inv_8[5] ^ r_7[5] /*365*/;
  assign sum_8[5] = _412_ ^ _411_ /*364*/;
  assign _413_ = _412_ & _411_ /*363*/;
  assign _414_ = inv_8[5] & r_7[5] /*362*/;
  assign _415_ = _413_ | _414_ /*361*/;
  assign _416_ = inv_8[6] ^ r_7[6] /*360*/;
  assign sum_8[6] = _416_ ^ _415_ /*359*/;
  assign _417_ = _416_ & _415_ /*358*/;
  assign _418_ = inv_8[6] & r_7[6] /*357*/;
  assign _419_ = _417_ | _418_ /*356*/;
  assign _420_ = inv_8[7] ^ r_7[7] /*355*/;
  assign sum_8[7] = _420_ ^ _419_ /*354*/;
  assign _421_ = _420_ & _419_ /*353*/;
  assign _422_ = inv_8[7] & r_7[7] /*352*/;
  assign _423_ = _421_ | _422_ /*351*/;
  assign Q[0] = ~sum_8[7] /*349*/;
  assign m_8[0] = r_7[0] /*348*/;
  assign m_8[1] = r_7[1] /*347*/;
  assign m_8[2] = r_7[2] /*346*/;
  assign m_8[3] = r_7[3] /*345*/;
  assign m_8[4] = r_7[4] /*344*/;
  assign m_8[5] = r_7[5] /*343*/;
  assign m_8[6] = r_7[6] /*342*/;
  assign m_8[7] = r_7[7] /*341*/;
  assign _424_ = ~Q[0] /*339*/;
  assign _425_ = sum_8[0] & Q[0] /*338*/;
  assign _426_ = m_8[0] & _424_ /*337*/;
  assign r_8[0] = _426_ | _425_ /*336*/;
  assign _427_ = ~Q[0] /*335*/;
  assign _428_ = sum_8[1] & Q[0] /*334*/;
  assign _429_ = m_8[1] & _427_ /*333*/;
  assign r_8[1] = _429_ | _428_ /*332*/;
  assign _430_ = ~Q[0] /*331*/;
  assign _431_ = sum_8[2] & Q[0] /*330*/;
  assign _432_ = m_8[2] & _430_ /*329*/;
  assign r_8[2] = _432_ | _431_ /*328*/;
  assign _433_ = ~Q[0] /*327*/;
  assign _434_ = sum_8[3] & Q[0] /*326*/;
  assign _435_ = m_8[3] & _433_ /*325*/;
  assign r_8[3] = _435_ | _434_ /*324*/;
  assign _436_ = ~Q[0] /*323*/;
  assign _437_ = sum_8[4] & Q[0] /*322*/;
  assign _438_ = m_8[4] & _436_ /*321*/;
  assign r_8[4] = _438_ | _437_ /*320*/;
  assign _439_ = ~Q[0] /*319*/;
  assign _440_ = sum_8[5] & Q[0] /*318*/;
  assign _441_ = m_8[5] & _439_ /*317*/;
  assign r_8[5] = _441_ | _440_ /*316*/;
  assign _442_ = ~Q[0] /*315*/;
  assign _443_ = sum_8[6] & Q[0] /*314*/;
  assign _444_ = m_8[6] & _442_ /*313*/;
  assign r_8[6] = _444_ | _443_ /*312*/;
  assign _445_ = ~Q[0] /*311*/;
  assign _446_ = sum_8[7] & Q[0] /*310*/;
  assign _447_ = m_8[7] & _445_ /*309*/;
  assign r_8[7] = _447_ | _446_ /*308*/;
  assign R_n1[0] = r_8[0] /*0*/;
  assign R_n1[1] = r_8[1] /*1*/;
  assign R_n1[2] = r_8[2] /*2*/;
  assign R_n1[3] = r_8[3] /*3*/;
  assign R_n1[4] = r_8[4] /*4*/;
  assign R_n1[5] = r_8[5] /*5*/;
  assign R_n1[6] = r_8[6] /*6*/;
  assign R_n1[7] = r_8[7] /*7*/;
endmodule