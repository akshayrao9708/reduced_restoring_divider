module nonresdivReduced(R_0, D, Q, R_n1);
input [13:0] R_0;
input [6:0] D;
output [7:0] Q;
output [7:0] R_n1;
wire _0_;
wire _1_;
wire _2_;
wire _3_;
wire _4_;
wire _5_;
wire _6_;
wire _7_;
wire _8_;
wire _9_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire _30_;
wire _31_;
wire _32_;
wire _33_;
wire _34_;
wire _35_;
wire _36_;
wire _37_;
wire _38_;
wire _39_;
wire _40_;
wire _41_;
wire _42_;
wire _43_;
wire _44_;
wire _45_;
wire _46_;
wire _47_;
wire _48_;
wire _49_;
wire _50_;
wire _51_;
wire _52_;
wire _53_;
wire _54_;
wire _55_;
wire _56_;
wire _57_;
wire _58_;
wire _59_;
wire _60_;
wire _61_;
wire _62_;
wire _63_;
wire _64_;
wire _65_;
wire _66_;
wire _67_;
wire _68_;
wire _69_;
wire _70_;
wire _71_;
wire _72_;
wire _73_;
wire _74_;
wire _75_;
wire _76_;
wire _77_;
wire _78_;
wire _79_;
wire _80_;
wire _81_;
wire _82_;
wire _83_;
wire _84_;
wire _85_;
wire _86_;
wire _87_;
wire _88_;
wire _89_;
wire _90_;
wire _91_;
wire _92_;
wire _93_;
wire _94_;
wire _95_;
wire _96_;
wire _97_;
wire _98_;
wire _99_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
wire _255_;
wire _256_;
wire _257_;
wire _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire _267_;
wire _268_;
wire _269_;
wire _270_;
wire _271_;
wire _272_;
wire _273_;
wire _274_;
wire _275_;
wire _276_;
wire _277_;
wire _278_;
wire _279_;
wire _280_;
wire _281_;
wire _282_;
wire _283_;
wire _284_;
wire _285_;
wire _286_;
wire _287_;
wire _288_;
wire _289_;
wire _290_;
wire _291_;
wire _292_;
wire _293_;
wire _294_;
wire _295_;
wire _296_;
wire _297_;
wire _298_;
wire _299_;
wire _300_;
wire _301_;
wire _302_;
wire _303_;
wire _304_;
wire _305_;
wire _306_;
wire _307_;
wire _308_;
wire _309_;
wire _310_;
wire _311_;
wire _312_;
wire _313_;
wire _314_;
wire _315_;
wire _316_;
wire _317_;
wire _318_;
wire _319_;
wire _320_;
wire _321_;
wire _322_;
wire _323_;
wire _324_;
wire _325_;
wire _326_;
wire _327_;
wire _328_;
wire _329_;
wire _330_;
wire _331_;
wire _332_;
wire _333_;
wire _334_;
wire _335_;
wire _336_;
wire _337_;
wire _338_;
wire _339_;
wire _340_;
wire _341_;
wire _342_;
wire _343_;
wire _344_;
wire _345_;
wire _346_;
wire _347_;
wire _348_;
wire _349_;
wire _350_;
wire _351_;
wire _352_;
wire _353_;
wire _354_;
wire _355_;
wire _356_;
wire _357_;
wire _358_;
wire _359_;
wire _360_;
wire _361_;
wire _362_;
wire _363_;
wire _364_;
wire _365_;
wire _366_;
wire _367_;
wire _368_;
wire _369_;
wire _370_;
wire _371_;
wire _372_;
wire _373_;
wire _374_;
wire _375_;
wire _376_;
wire _377_;
wire _378_;
wire _379_;
wire _380_;
wire _381_;
wire _382_;
wire _383_;
wire _384_;
wire _385_;
wire _386_;
wire _387_;
wire _388_;
wire _389_;
wire _390_;
wire _391_;
wire _392_;
wire _393_;
wire _394_;
wire _395_;
wire _396_;
wire _397_;
wire _398_;
wire _399_;
wire _400_;
wire _401_;
wire _402_;
wire _403_;
wire _404_;
wire _405_;
wire _406_;
wire _407_;
wire _408_;
wire _409_;
wire _410_;
wire _411_;
wire _412_;
wire _413_;
wire _414_;
wire _415_;
wire _416_;
wire _417_;
wire _418_;
wire _419_;
wire _420_;
wire _421_;
wire _422_;
wire _423_;
wire _424_;
wire _425_;
wire _426_;
wire _427_;
wire _428_;
wire _429_;
wire zeroWire;
wire oneWire;
assign zeroWire = 1'b0 /*867*/;
assign oneWire = 1'b1 /*867*/;
assign _11_ = ~D[0] /*817*/;
assign _9_ = R_0[7] | _11_ /*814*/;
assign _10_ = R_0[7] ^ _11_ /*816*/;
assign _0_ = ~_10_ /*815*/;
assign _18_ = ~D[1] /*813*/;
assign _15_ = R_0[8] & _18_ /*809*/;
assign _16_ = R_0[8] ^ _18_ /*812*/;
assign _17_ = _9_ & _16_ /*810*/;
assign _14_ = _15_ | _17_ /*808*/;
assign _1_ = _9_ ^ _16_ /*811*/;
assign _23_ = ~D[2] /*807*/;
assign _20_ = R_0[9] & _23_ /*803*/;
assign _21_ = R_0[9] ^ _23_ /*806*/;
assign _22_ = _14_ & _21_ /*804*/;
assign _19_ = _20_ | _22_ /*802*/;
assign _2_ = _14_ ^ _21_ /*805*/;
assign _28_ = ~D[3] /*801*/;
assign _25_ = R_0[10] & _28_ /*797*/;
assign _26_ = R_0[10] ^ _28_ /*800*/;
assign _27_ = _19_ & _26_ /*798*/;
assign _24_ = _25_ | _27_ /*796*/;
assign _3_ = _19_ ^ _26_ /*799*/;
assign _33_ = ~D[4] /*795*/;
assign _30_ = R_0[11] & _33_ /*791*/;
assign _31_ = R_0[11] ^ _33_ /*794*/;
assign _32_ = _24_ & _31_ /*792*/;
assign _29_ = _30_ | _32_ /*790*/;
assign _4_ = _24_ ^ _31_ /*793*/;
assign _38_ = ~D[5] /*789*/;
assign _35_ = R_0[12] & _38_ /*785*/;
assign _36_ = R_0[12] ^ _38_ /*788*/;
assign _37_ = _29_ & _36_ /*786*/;
assign _34_ = _35_ | _37_ /*784*/;
assign _5_ = _29_ ^ _36_ /*787*/;
assign _43_ = ~D[6] /*783*/;
assign _40_ = R_0[13] & _43_ /*779*/;
assign _41_ = R_0[13] ^ _43_ /*782*/;
assign _42_ = _34_ & _41_ /*780*/;
assign _39_ = _40_ | _42_ /*778*/;
assign _6_ = _34_ ^ _41_ /*781*/;
assign _44_ = zeroWire & oneWire /*773*/;
assign _45_ = zeroWire ^ oneWire /*776*/;
assign _46_ = _39_ & _45_ /*774*/;
assign Q[7] = _44_ | _46_ /*772*/;
assign _7_ = _39_ ^ _45_ /*775*/;
assign _62_ = D[0] ^ Q[7] /*722*/;
assign _59_ = R_0[6] & _62_ /*718*/;
assign _60_ = R_0[6] ^ _62_ /*721*/;
assign _61_ = Q[7] & _60_ /*719*/;
assign _58_ = _59_ | _61_ /*717*/;
assign _49_ = Q[7] ^ _60_ /*720*/;
assign _67_ = D[1] ^ Q[7] /*716*/;
assign _64_ = _0_ & _67_ /*712*/;
assign _65_ = _0_ ^ _67_ /*715*/;
assign _66_ = _58_ & _65_ /*713*/;
assign _63_ = _64_ | _66_ /*711*/;
assign _50_ = _58_ ^ _65_ /*714*/;
assign _72_ = D[2] ^ Q[7] /*710*/;
assign _69_ = _1_ & _72_ /*706*/;
assign _70_ = _1_ ^ _72_ /*709*/;
assign _71_ = _63_ & _70_ /*707*/;
assign _68_ = _69_ | _71_ /*705*/;
assign _51_ = _63_ ^ _70_ /*708*/;
assign _77_ = D[3] ^ Q[7] /*704*/;
assign _74_ = _2_ & _77_ /*700*/;
assign _75_ = _2_ ^ _77_ /*703*/;
assign _76_ = _68_ & _75_ /*701*/;
assign _73_ = _74_ | _76_ /*699*/;
assign _52_ = _68_ ^ _75_ /*702*/;
assign _82_ = D[4] ^ Q[7] /*698*/;
assign _79_ = _3_ & _82_ /*694*/;
assign _80_ = _3_ ^ _82_ /*697*/;
assign _81_ = _73_ & _80_ /*695*/;
assign _78_ = _79_ | _81_ /*693*/;
assign _53_ = _73_ ^ _80_ /*696*/;
assign _87_ = D[5] ^ Q[7] /*692*/;
assign _84_ = _4_ & _87_ /*688*/;
assign _85_ = _4_ ^ _87_ /*691*/;
assign _86_ = _78_ & _85_ /*689*/;
assign _83_ = _84_ | _86_ /*687*/;
assign _54_ = _78_ ^ _85_ /*690*/;
assign _92_ = D[6] ^ Q[7] /*686*/;
assign _89_ = _5_ & _92_ /*682*/;
assign _90_ = _5_ ^ _92_ /*685*/;
assign _91_ = _83_ & _90_ /*683*/;
assign _88_ = _89_ | _91_ /*681*/;
assign _55_ = _83_ ^ _90_ /*684*/;
assign _96_ = zeroWire ^ Q[7] /*680*/;
assign _93_ = _6_ & _96_ /*676*/;
assign _94_ = _6_ ^ _96_ /*679*/;
assign _95_ = _88_ & _94_ /*677*/;
assign Q[6] = _93_ | _95_ /*675*/;
assign _56_ = _88_ ^ _94_ /*678*/;
assign _111_ = D[0] ^ Q[6] /*625*/;
assign _108_ = R_0[5] & _111_ /*621*/;
assign _109_ = R_0[5] ^ _111_ /*624*/;
assign _110_ = Q[6] & _109_ /*622*/;
assign _107_ = _108_ | _110_ /*620*/;
assign _98_ = Q[6] ^ _109_ /*623*/;
assign _116_ = D[1] ^ Q[6] /*619*/;
assign _113_ = _49_ & _116_ /*615*/;
assign _114_ = _49_ ^ _116_ /*618*/;
assign _115_ = _107_ & _114_ /*616*/;
assign _112_ = _113_ | _115_ /*614*/;
assign _99_ = _107_ ^ _114_ /*617*/;
assign _121_ = D[2] ^ Q[6] /*613*/;
assign _118_ = _50_ & _121_ /*609*/;
assign _119_ = _50_ ^ _121_ /*612*/;
assign _120_ = _112_ & _119_ /*610*/;
assign _117_ = _118_ | _120_ /*608*/;
assign _100_ = _112_ ^ _119_ /*611*/;
assign _126_ = D[3] ^ Q[6] /*607*/;
assign _123_ = _51_ & _126_ /*603*/;
assign _124_ = _51_ ^ _126_ /*606*/;
assign _125_ = _117_ & _124_ /*604*/;
assign _122_ = _123_ | _125_ /*602*/;
assign _101_ = _117_ ^ _124_ /*605*/;
assign _131_ = D[4] ^ Q[6] /*601*/;
assign _128_ = _52_ & _131_ /*597*/;
assign _129_ = _52_ ^ _131_ /*600*/;
assign _130_ = _122_ & _129_ /*598*/;
assign _127_ = _128_ | _130_ /*596*/;
assign _102_ = _122_ ^ _129_ /*599*/;
assign _136_ = D[5] ^ Q[6] /*595*/;
assign _133_ = _53_ & _136_ /*591*/;
assign _134_ = _53_ ^ _136_ /*594*/;
assign _135_ = _127_ & _134_ /*592*/;
assign _132_ = _133_ | _135_ /*590*/;
assign _103_ = _127_ ^ _134_ /*593*/;
assign _141_ = D[6] ^ Q[6] /*589*/;
assign _138_ = _54_ & _141_ /*585*/;
assign _139_ = _54_ ^ _141_ /*588*/;
assign _140_ = _132_ & _139_ /*586*/;
assign _137_ = _138_ | _140_ /*584*/;
assign _104_ = _132_ ^ _139_ /*587*/;
assign _145_ = zeroWire ^ Q[6] /*583*/;
assign _142_ = _55_ & _145_ /*579*/;
assign _143_ = _55_ ^ _145_ /*582*/;
assign _144_ = _137_ & _143_ /*580*/;
assign Q[5] = _142_ | _144_ /*578*/;
assign _105_ = _137_ ^ _143_ /*581*/;
assign _160_ = D[0] ^ Q[5] /*528*/;
assign _157_ = R_0[4] & _160_ /*524*/;
assign _158_ = R_0[4] ^ _160_ /*527*/;
assign _159_ = Q[5] & _158_ /*525*/;
assign _156_ = _157_ | _159_ /*523*/;
assign _147_ = Q[5] ^ _158_ /*526*/;
assign _165_ = D[1] ^ Q[5] /*522*/;
assign _162_ = _98_ & _165_ /*518*/;
assign _163_ = _98_ ^ _165_ /*521*/;
assign _164_ = _156_ & _163_ /*519*/;
assign _161_ = _162_ | _164_ /*517*/;
assign _148_ = _156_ ^ _163_ /*520*/;
assign _170_ = D[2] ^ Q[5] /*516*/;
assign _167_ = _99_ & _170_ /*512*/;
assign _168_ = _99_ ^ _170_ /*515*/;
assign _169_ = _161_ & _168_ /*513*/;
assign _166_ = _167_ | _169_ /*511*/;
assign _149_ = _161_ ^ _168_ /*514*/;
assign _175_ = D[3] ^ Q[5] /*510*/;
assign _172_ = _100_ & _175_ /*506*/;
assign _173_ = _100_ ^ _175_ /*509*/;
assign _174_ = _166_ & _173_ /*507*/;
assign _171_ = _172_ | _174_ /*505*/;
assign _150_ = _166_ ^ _173_ /*508*/;
assign _180_ = D[4] ^ Q[5] /*504*/;
assign _177_ = _101_ & _180_ /*500*/;
assign _178_ = _101_ ^ _180_ /*503*/;
assign _179_ = _171_ & _178_ /*501*/;
assign _176_ = _177_ | _179_ /*499*/;
assign _151_ = _171_ ^ _178_ /*502*/;
assign _185_ = D[5] ^ Q[5] /*498*/;
assign _182_ = _102_ & _185_ /*494*/;
assign _183_ = _102_ ^ _185_ /*497*/;
assign _184_ = _176_ & _183_ /*495*/;
assign _181_ = _182_ | _184_ /*493*/;
assign _152_ = _176_ ^ _183_ /*496*/;
assign _190_ = D[6] ^ Q[5] /*492*/;
assign _187_ = _103_ & _190_ /*488*/;
assign _188_ = _103_ ^ _190_ /*491*/;
assign _189_ = _181_ & _188_ /*489*/;
assign _186_ = _187_ | _189_ /*487*/;
assign _153_ = _181_ ^ _188_ /*490*/;
assign _194_ = zeroWire ^ Q[5] /*486*/;
assign _191_ = _104_ & _194_ /*482*/;
assign _192_ = _104_ ^ _194_ /*485*/;
assign _193_ = _186_ & _192_ /*483*/;
assign Q[4] = _191_ | _193_ /*481*/;
assign _154_ = _186_ ^ _192_ /*484*/;
assign _209_ = D[0] ^ Q[4] /*431*/;
assign _206_ = R_0[3] & _209_ /*427*/;
assign _207_ = R_0[3] ^ _209_ /*430*/;
assign _208_ = Q[4] & _207_ /*428*/;
assign _205_ = _206_ | _208_ /*426*/;
assign _196_ = Q[4] ^ _207_ /*429*/;
assign _214_ = D[1] ^ Q[4] /*425*/;
assign _211_ = _147_ & _214_ /*421*/;
assign _212_ = _147_ ^ _214_ /*424*/;
assign _213_ = _205_ & _212_ /*422*/;
assign _210_ = _211_ | _213_ /*420*/;
assign _197_ = _205_ ^ _212_ /*423*/;
assign _219_ = D[2] ^ Q[4] /*419*/;
assign _216_ = _148_ & _219_ /*415*/;
assign _217_ = _148_ ^ _219_ /*418*/;
assign _218_ = _210_ & _217_ /*416*/;
assign _215_ = _216_ | _218_ /*414*/;
assign _198_ = _210_ ^ _217_ /*417*/;
assign _224_ = D[3] ^ Q[4] /*413*/;
assign _221_ = _149_ & _224_ /*409*/;
assign _222_ = _149_ ^ _224_ /*412*/;
assign _223_ = _215_ & _222_ /*410*/;
assign _220_ = _221_ | _223_ /*408*/;
assign _199_ = _215_ ^ _222_ /*411*/;
assign _229_ = D[4] ^ Q[4] /*407*/;
assign _226_ = _150_ & _229_ /*403*/;
assign _227_ = _150_ ^ _229_ /*406*/;
assign _228_ = _220_ & _227_ /*404*/;
assign _225_ = _226_ | _228_ /*402*/;
assign _200_ = _220_ ^ _227_ /*405*/;
assign _234_ = D[5] ^ Q[4] /*401*/;
assign _231_ = _151_ & _234_ /*397*/;
assign _232_ = _151_ ^ _234_ /*400*/;
assign _233_ = _225_ & _232_ /*398*/;
assign _230_ = _231_ | _233_ /*396*/;
assign _201_ = _225_ ^ _232_ /*399*/;
assign _239_ = D[6] ^ Q[4] /*395*/;
assign _236_ = _152_ & _239_ /*391*/;
assign _237_ = _152_ ^ _239_ /*394*/;
assign _238_ = _230_ & _237_ /*392*/;
assign _235_ = _236_ | _238_ /*390*/;
assign _202_ = _230_ ^ _237_ /*393*/;
assign _243_ = zeroWire ^ Q[4] /*389*/;
assign _240_ = _153_ & _243_ /*385*/;
assign _241_ = _153_ ^ _243_ /*388*/;
assign _242_ = _235_ & _241_ /*386*/;
assign Q[3] = _240_ | _242_ /*384*/;
assign _203_ = _235_ ^ _241_ /*387*/;
assign _258_ = D[0] ^ Q[3] /*334*/;
assign _255_ = R_0[2] & _258_ /*330*/;
assign _256_ = R_0[2] ^ _258_ /*333*/;
assign _257_ = Q[3] & _256_ /*331*/;
assign _254_ = _255_ | _257_ /*329*/;
assign _245_ = Q[3] ^ _256_ /*332*/;
assign _263_ = D[1] ^ Q[3] /*328*/;
assign _260_ = _196_ & _263_ /*324*/;
assign _261_ = _196_ ^ _263_ /*327*/;
assign _262_ = _254_ & _261_ /*325*/;
assign _259_ = _260_ | _262_ /*323*/;
assign _246_ = _254_ ^ _261_ /*326*/;
assign _268_ = D[2] ^ Q[3] /*322*/;
assign _265_ = _197_ & _268_ /*318*/;
assign _266_ = _197_ ^ _268_ /*321*/;
assign _267_ = _259_ & _266_ /*319*/;
assign _264_ = _265_ | _267_ /*317*/;
assign _247_ = _259_ ^ _266_ /*320*/;
assign _273_ = D[3] ^ Q[3] /*316*/;
assign _270_ = _198_ & _273_ /*312*/;
assign _271_ = _198_ ^ _273_ /*315*/;
assign _272_ = _264_ & _271_ /*313*/;
assign _269_ = _270_ | _272_ /*311*/;
assign _248_ = _264_ ^ _271_ /*314*/;
assign _278_ = D[4] ^ Q[3] /*310*/;
assign _275_ = _199_ & _278_ /*306*/;
assign _276_ = _199_ ^ _278_ /*309*/;
assign _277_ = _269_ & _276_ /*307*/;
assign _274_ = _275_ | _277_ /*305*/;
assign _249_ = _269_ ^ _276_ /*308*/;
assign _283_ = D[5] ^ Q[3] /*304*/;
assign _280_ = _200_ & _283_ /*300*/;
assign _281_ = _200_ ^ _283_ /*303*/;
assign _282_ = _274_ & _281_ /*301*/;
assign _279_ = _280_ | _282_ /*299*/;
assign _250_ = _274_ ^ _281_ /*302*/;
assign _288_ = D[6] ^ Q[3] /*298*/;
assign _285_ = _201_ & _288_ /*294*/;
assign _286_ = _201_ ^ _288_ /*297*/;
assign _287_ = _279_ & _286_ /*295*/;
assign _284_ = _285_ | _287_ /*293*/;
assign _251_ = _279_ ^ _286_ /*296*/;
assign _292_ = zeroWire ^ Q[3] /*292*/;
assign _289_ = _202_ & _292_ /*288*/;
assign _290_ = _202_ ^ _292_ /*291*/;
assign _291_ = _284_ & _290_ /*289*/;
assign Q[2] = _289_ | _291_ /*287*/;
assign _252_ = _284_ ^ _290_ /*290*/;
assign _307_ = D[0] ^ Q[2] /*237*/;
assign _304_ = R_0[1] & _307_ /*233*/;
assign _305_ = R_0[1] ^ _307_ /*236*/;
assign _306_ = Q[2] & _305_ /*234*/;
assign _303_ = _304_ | _306_ /*232*/;
assign _294_ = Q[2] ^ _305_ /*235*/;
assign _312_ = D[1] ^ Q[2] /*231*/;
assign _309_ = _245_ & _312_ /*227*/;
assign _310_ = _245_ ^ _312_ /*230*/;
assign _311_ = _303_ & _310_ /*228*/;
assign _308_ = _309_ | _311_ /*226*/;
assign _295_ = _303_ ^ _310_ /*229*/;
assign _317_ = D[2] ^ Q[2] /*225*/;
assign _314_ = _246_ & _317_ /*221*/;
assign _315_ = _246_ ^ _317_ /*224*/;
assign _316_ = _308_ & _315_ /*222*/;
assign _313_ = _314_ | _316_ /*220*/;
assign _296_ = _308_ ^ _315_ /*223*/;
assign _322_ = D[3] ^ Q[2] /*219*/;
assign _319_ = _247_ & _322_ /*215*/;
assign _320_ = _247_ ^ _322_ /*218*/;
assign _321_ = _313_ & _320_ /*216*/;
assign _318_ = _319_ | _321_ /*214*/;
assign _297_ = _313_ ^ _320_ /*217*/;
assign _327_ = D[4] ^ Q[2] /*213*/;
assign _324_ = _248_ & _327_ /*209*/;
assign _325_ = _248_ ^ _327_ /*212*/;
assign _326_ = _318_ & _325_ /*210*/;
assign _323_ = _324_ | _326_ /*208*/;
assign _298_ = _318_ ^ _325_ /*211*/;
assign _332_ = D[5] ^ Q[2] /*207*/;
assign _329_ = _249_ & _332_ /*203*/;
assign _330_ = _249_ ^ _332_ /*206*/;
assign _331_ = _323_ & _330_ /*204*/;
assign _328_ = _329_ | _331_ /*202*/;
assign _299_ = _323_ ^ _330_ /*205*/;
assign _337_ = D[6] ^ Q[2] /*201*/;
assign _334_ = _250_ & _337_ /*197*/;
assign _335_ = _250_ ^ _337_ /*200*/;
assign _336_ = _328_ & _335_ /*198*/;
assign _333_ = _334_ | _336_ /*196*/;
assign _300_ = _328_ ^ _335_ /*199*/;
assign _341_ = zeroWire ^ Q[2] /*195*/;
assign _338_ = _251_ & _341_ /*191*/;
assign _339_ = _251_ ^ _341_ /*194*/;
assign _340_ = _333_ & _339_ /*192*/;
assign Q[1] = _338_ | _340_ /*190*/;
assign _301_ = _333_ ^ _339_ /*193*/;
assign _356_ = D[0] ^ Q[1] /*140*/;
assign _353_ = R_0[0] & _356_ /*136*/;
assign _354_ = R_0[0] ^ _356_ /*139*/;
assign _355_ = Q[1] & _354_ /*137*/;
assign _352_ = _353_ | _355_ /*135*/;
assign _343_ = Q[1] ^ _354_ /*138*/;
assign _361_ = D[1] ^ Q[1] /*134*/;
assign _358_ = _294_ & _361_ /*130*/;
assign _359_ = _294_ ^ _361_ /*133*/;
assign _360_ = _352_ & _359_ /*131*/;
assign _357_ = _358_ | _360_ /*129*/;
assign _344_ = _352_ ^ _359_ /*132*/;
assign _366_ = D[2] ^ Q[1] /*128*/;
assign _363_ = _295_ & _366_ /*124*/;
assign _364_ = _295_ ^ _366_ /*127*/;
assign _365_ = _357_ & _364_ /*125*/;
assign _362_ = _363_ | _365_ /*123*/;
assign _345_ = _357_ ^ _364_ /*126*/;
assign _371_ = D[3] ^ Q[1] /*122*/;
assign _368_ = _296_ & _371_ /*118*/;
assign _369_ = _296_ ^ _371_ /*121*/;
assign _370_ = _362_ & _369_ /*119*/;
assign _367_ = _368_ | _370_ /*117*/;
assign _346_ = _362_ ^ _369_ /*120*/;
assign _376_ = D[4] ^ Q[1] /*116*/;
assign _373_ = _297_ & _376_ /*112*/;
assign _374_ = _297_ ^ _376_ /*115*/;
assign _375_ = _367_ & _374_ /*113*/;
assign _372_ = _373_ | _375_ /*111*/;
assign _347_ = _367_ ^ _374_ /*114*/;
assign _381_ = D[5] ^ Q[1] /*110*/;
assign _378_ = _298_ & _381_ /*106*/;
assign _379_ = _298_ ^ _381_ /*109*/;
assign _380_ = _372_ & _379_ /*107*/;
assign _377_ = _378_ | _380_ /*105*/;
assign _348_ = _372_ ^ _379_ /*108*/;
assign _386_ = D[6] ^ Q[1] /*104*/;
assign _383_ = _299_ & _386_ /*100*/;
assign _384_ = _299_ ^ _386_ /*103*/;
assign _385_ = _377_ & _384_ /*101*/;
assign _382_ = _383_ | _385_ /*99*/;
assign _349_ = _377_ ^ _384_ /*102*/;
assign _390_ = zeroWire ^ Q[1] /*98*/;
assign _387_ = _300_ & _390_ /*94*/;
assign _388_ = _300_ ^ _390_ /*97*/;
assign _389_ = _382_ & _388_ /*95*/;
assign Q[0] = _387_ | _389_ /*93*/;
assign _350_ = _382_ ^ _388_ /*92*/;
assign _392_ = ~Q[0] /*43*/;
assign _393_ = _392_ & D[0] /*42*/;
assign _394_ = _343_ & _393_ /*40*/;
assign R_n1[0] = _343_ ^ _393_ /*41*/;
assign _398_ = _392_ & D[1] /*39*/;
assign _400_ = _344_ & _398_ /*35*/;
assign _401_ = _344_ ^ _398_ /*38*/;
assign _402_ = _394_ & _401_ /*36*/;
assign _399_ = _400_ | _402_ /*34*/;
assign R_n1[1] = _394_ ^ _401_ /*37*/;
assign _403_ = _392_ & D[2] /*33*/;
assign _405_ = _345_ & _403_ /*29*/;
assign _406_ = _345_ ^ _403_ /*32*/;
assign _407_ = _399_ & _406_ /*30*/;
assign _404_ = _405_ | _407_ /*28*/;
assign R_n1[2] = _399_ ^ _406_ /*31*/;
assign _408_ = _392_ & D[3] /*27*/;
assign _410_ = _346_ & _408_ /*23*/;
assign _411_ = _346_ ^ _408_ /*26*/;
assign _412_ = _404_ & _411_ /*24*/;
assign _409_ = _410_ | _412_ /*22*/;
assign R_n1[3] = _404_ ^ _411_ /*25*/;
assign _413_ = _392_ & D[4] /*21*/;
assign _415_ = _347_ & _413_ /*17*/;
assign _416_ = _347_ ^ _413_ /*20*/;
assign _417_ = _409_ & _416_ /*18*/;
assign _414_ = _415_ | _417_ /*16*/;
assign R_n1[4] = _409_ ^ _416_ /*19*/;
assign _418_ = _392_ & D[5] /*15*/;
assign _420_ = _348_ & _418_ /*11*/;
assign _421_ = _348_ ^ _418_ /*14*/;
assign _422_ = _414_ & _421_ /*12*/;
assign _419_ = _420_ | _422_ /*10*/;
assign R_n1[5] = _414_ ^ _421_ /*13*/;
assign _423_ = _392_ & D[6] /*9*/;
assign _425_ = _349_ & _423_ /*5*/;
assign _426_ = _349_ ^ _423_ /*8*/;
assign _427_ = _419_ & _426_ /*6*/;
assign _424_ = _425_ | _427_ /*4*/;
assign R_n1[6] = _419_ ^ _426_ /*7*/;
assign _428_ = _392_ & zeroWire /*3*/;
assign _429_ = _350_ ^ _428_ /*2*/;
assign R_n1[7] = _429_ ^ _424_ /*1*/;
endmodule
