module divider(R_0, D, Q, R_n1);
input [29:0] R_0;
input [14:0] D;
output [15:0] Q;
output [14:0] R_n1;
wire _0_;
wire _1_;
wire _2_;
wire _3_;
wire _4_;
wire _5_;
wire _6_;
wire _7_;
wire _8_;
wire _9_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire _30_;
wire _31_;
wire _32_;
wire _33_;
wire _34_;
wire _35_;
wire _36_;
wire _37_;
wire _38_;
wire _39_;
wire _40_;
wire _41_;
wire _42_;
wire _43_;
wire _44_;
wire _45_;
wire _46_;
wire _47_;
wire _48_;
wire _49_;
wire _50_;
wire _51_;
wire _52_;
wire _53_;
wire _54_;
wire _55_;
wire _56_;
wire _57_;
wire _58_;
wire _59_;
wire _60_;
wire _61_;
wire _62_;
wire _63_;
wire _64_;
wire _65_;
wire _66_;
wire _67_;
wire _68_;
wire _69_;
wire _70_;
wire _71_;
wire _72_;
wire _73_;
wire _74_;
wire _75_;
wire _76_;
wire _77_;
wire _78_;
wire _79_;
wire _80_;
wire _81_;
wire _82_;
wire _83_;
wire _84_;
wire _85_;
wire _86_;
wire _87_;
wire _88_;
wire _89_;
wire _90_;
wire _91_;
wire _92_;
wire _93_;
wire _94_;
wire _95_;
wire _96_;
wire _97_;
wire _98_;
wire _99_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
wire _255_;
wire _256_;
wire _257_;
wire _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire _267_;
wire _268_;
wire _269_;
wire _270_;
wire _271_;
wire _272_;
wire _273_;
wire _274_;
wire _275_;
wire _276_;
wire _277_;
wire _278_;
wire _279_;
wire _280_;
wire _281_;
wire _282_;
wire _283_;
wire _284_;
wire _285_;
wire _286_;
wire _287_;
wire _288_;
wire _289_;
wire _290_;
wire _291_;
wire _292_;
wire _293_;
wire _294_;
wire _295_;
wire _296_;
wire _297_;
wire _298_;
wire _299_;
wire _300_;
wire _301_;
wire _302_;
wire _303_;
wire _304_;
wire _305_;
wire _306_;
wire _307_;
wire _308_;
wire _309_;
wire _310_;
wire _311_;
wire _312_;
wire _313_;
wire _314_;
wire _315_;
wire _316_;
wire _317_;
wire _318_;
wire _319_;
wire _320_;
wire _321_;
wire _322_;
wire _323_;
wire _324_;
wire _325_;
wire _326_;
wire _327_;
wire _328_;
wire _329_;
wire _330_;
wire _331_;
wire _332_;
wire _333_;
wire _334_;
wire _335_;
wire _336_;
wire _337_;
wire _338_;
wire _339_;
wire _340_;
wire _341_;
wire _342_;
wire _343_;
wire _344_;
wire _345_;
wire _346_;
wire _347_;
wire _348_;
wire _349_;
wire _350_;
wire _351_;
wire _352_;
wire _353_;
wire _354_;
wire _355_;
wire _356_;
wire _357_;
wire _358_;
wire _359_;
wire _360_;
wire _361_;
wire _362_;
wire _363_;
wire _364_;
wire _365_;
wire _366_;
wire _367_;
wire _368_;
wire _369_;
wire _370_;
wire _371_;
wire _372_;
wire _373_;
wire _374_;
wire _375_;
wire _376_;
wire _377_;
wire _378_;
wire _379_;
wire _380_;
wire _381_;
wire _382_;
wire _383_;
wire _384_;
wire _385_;
wire _386_;
wire _387_;
wire _388_;
wire _389_;
wire _390_;
wire _391_;
wire _392_;
wire _393_;
wire _394_;
wire _395_;
wire _396_;
wire _397_;
wire _398_;
wire _399_;
wire _400_;
wire _401_;
wire _402_;
wire _403_;
wire _404_;
wire _405_;
wire _406_;
wire _407_;
wire _408_;
wire _409_;
wire _410_;
wire _411_;
wire _412_;
wire _413_;
wire _414_;
wire _415_;
wire _416_;
wire _417_;
wire _418_;
wire _419_;
wire _420_;
wire _421_;
wire _422_;
wire _423_;
wire _424_;
wire _425_;
wire _426_;
wire _427_;
wire _428_;
wire _429_;
wire _430_;
wire _431_;
wire _432_;
wire _433_;
wire _434_;
wire _435_;
wire _436_;
wire _437_;
wire _438_;
wire _439_;
wire _440_;
wire _441_;
wire _442_;
wire _443_;
wire _444_;
wire _445_;
wire _446_;
wire _447_;
wire _448_;
wire _449_;
wire _450_;
wire _451_;
wire _452_;
wire _453_;
wire _454_;
wire _455_;
wire _456_;
wire _457_;
wire _458_;
wire _459_;
wire _460_;
wire _461_;
wire _462_;
wire _463_;
wire _464_;
wire _465_;
wire _466_;
wire _467_;
wire _468_;
wire _469_;
wire _470_;
wire _471_;
wire _472_;
wire _473_;
wire _474_;
wire _475_;
wire _476_;
wire _477_;
wire _478_;
wire _479_;
wire _480_;
wire _481_;
wire _482_;
wire _483_;
wire _484_;
wire _485_;
wire _486_;
wire _487_;
wire _488_;
wire _489_;
wire _490_;
wire _491_;
wire _492_;
wire _493_;
wire _494_;
wire _495_;
wire _496_;
wire _497_;
wire _498_;
wire _499_;
wire _500_;
wire _501_;
wire _502_;
wire _503_;
wire _504_;
wire _505_;
wire _506_;
wire _507_;
wire _508_;
wire _509_;
wire _510_;
wire _511_;
wire _512_;
wire _513_;
wire _514_;
wire _515_;
wire _516_;
wire _517_;
wire _518_;
wire _519_;
wire _520_;
wire _521_;
wire _522_;
wire _523_;
wire _524_;
wire _525_;
wire _526_;
wire _527_;
wire _528_;
wire _529_;
wire _530_;
wire _531_;
wire _532_;
wire _533_;
wire _534_;
wire _535_;
wire _536_;
wire _537_;
wire _538_;
wire _539_;
wire _540_;
wire _541_;
wire _542_;
wire _543_;
wire _544_;
wire _545_;
wire _546_;
wire _547_;
wire _548_;
wire _549_;
wire _550_;
wire _551_;
wire _552_;
wire _553_;
wire _554_;
wire _555_;
wire _556_;
wire _557_;
wire _558_;
wire _559_;
wire _560_;
wire _561_;
wire _562_;
wire _563_;
wire _564_;
wire _565_;
wire _566_;
wire _567_;
wire _568_;
wire _569_;
wire _570_;
wire _571_;
wire _572_;
wire _573_;
wire _574_;
wire _575_;
wire _576_;
wire _577_;
wire _578_;
wire _579_;
wire _580_;
wire _581_;
wire _582_;
wire _583_;
wire _584_;
wire _585_;
wire _586_;
wire _587_;
wire _588_;
wire _589_;
wire _590_;
wire _591_;
wire _592_;
wire _593_;
wire _594_;
wire _595_;
wire _596_;
wire _597_;
wire _598_;
wire _599_;
wire _600_;
wire _601_;
wire _602_;
wire _603_;
wire _604_;
wire _605_;
wire _606_;
wire _607_;
wire _608_;
wire _609_;
wire _610_;
wire _611_;
wire _612_;
wire _613_;
wire _614_;
wire _615_;
wire _616_;
wire _617_;
wire _618_;
wire _619_;
wire _620_;
wire _621_;
wire _622_;
wire _623_;
wire _624_;
wire _625_;
wire _626_;
wire _627_;
wire _628_;
wire _629_;
wire _630_;
wire _631_;
wire _632_;
wire _633_;
wire _634_;
wire _635_;
wire _636_;
wire _637_;
wire _638_;
wire _639_;
wire _640_;
wire _641_;
wire _642_;
wire _643_;
wire _644_;
wire _645_;
wire _646_;
wire _647_;
wire _648_;
wire _649_;
wire _650_;
wire _651_;
wire _652_;
wire _653_;
wire _654_;
wire _655_;
wire _656_;
wire _657_;
wire _658_;
wire _659_;
wire _660_;
wire _661_;
wire _662_;
wire _663_;
wire _664_;
wire _665_;
wire _666_;
wire _667_;
wire _668_;
wire _669_;
wire _670_;
wire _671_;
wire _672_;
wire _673_;
wire _674_;
wire _675_;
wire _676_;
wire _677_;
wire _678_;
wire _679_;
wire _680_;
wire _681_;
wire _682_;
wire _683_;
wire _684_;
wire _685_;
wire _686_;
wire _687_;
wire _688_;
wire _689_;
wire _690_;
wire _691_;
wire _692_;
wire _693_;
wire _694_;
wire _695_;
wire _696_;
wire _697_;
wire _698_;
wire _699_;
wire _700_;
wire _701_;
wire _702_;
wire _703_;
wire _704_;
wire _705_;
wire _706_;
wire _707_;
wire _708_;
wire _709_;
wire _710_;
wire _711_;
wire _712_;
wire _713_;
wire _714_;
wire _715_;
wire _716_;
wire _717_;
wire _718_;
wire _719_;
wire _720_;
wire _721_;
wire _722_;
wire _723_;
wire _724_;
wire _725_;
wire _726_;
wire _727_;
wire _728_;
wire _729_;
wire _730_;
wire _731_;
wire _732_;
wire _733_;
wire _734_;
wire _735_;
wire _736_;
wire _737_;
wire _738_;
wire _739_;
wire _740_;
wire _741_;
wire _742_;
wire _743_;
wire _744_;
wire _745_;
wire _746_;
wire _747_;
wire _748_;
wire _749_;
wire _750_;
wire _751_;
wire _752_;
wire _753_;
wire _754_;
wire _755_;
wire _756_;
wire _757_;
wire _758_;
wire _759_;
wire _760_;
wire _761_;
wire _762_;
wire _763_;
wire _764_;
wire _765_;
wire _766_;
wire _767_;
wire _768_;
wire _769_;
wire _770_;
wire _771_;
wire _772_;
wire _773_;
wire _774_;
wire _775_;
wire _776_;
wire _777_;
wire _778_;
wire _779_;
wire _780_;
wire _781_;
wire _782_;
wire _783_;
wire _784_;
wire _785_;
wire _786_;
wire _787_;
wire _788_;
wire _789_;
wire _790_;
wire _791_;
wire _792_;
wire _793_;
wire _794_;
wire _795_;
wire _796_;
wire _797_;
wire _798_;
wire _799_;
wire _800_;
wire _801_;
wire _802_;
wire _803_;
wire _804_;
wire _805_;
wire _806_;
wire _807_;
wire _808_;
wire _809_;
wire _810_;
wire _811_;
wire _812_;
wire _813_;
wire _814_;
wire _815_;
wire _816_;
wire _817_;
wire _818_;
wire _819_;
wire _820_;
wire _821_;
wire _822_;
wire _823_;
wire _824_;
wire _825_;
wire _826_;
wire _827_;
wire _828_;
wire _829_;
wire _830_;
wire _831_;
wire _832_;
wire _833_;
wire _834_;
wire _835_;
wire _836_;
wire _837_;
wire _838_;
wire _839_;
wire _840_;
wire _841_;
wire _842_;
wire _843_;
wire _844_;
wire _845_;
wire _846_;
wire _847_;
wire _848_;
wire _849_;
wire _850_;
wire _851_;
wire _852_;
wire _853_;
wire _854_;
wire _855_;
wire _856_;
wire _857_;
wire _858_;
wire _859_;
wire _860_;
wire _861_;
wire _862_;
wire _863_;
wire _864_;
wire _865_;
wire _866_;
wire _867_;
wire _868_;
wire _869_;
wire _870_;
wire _871_;
wire _872_;
wire _873_;
wire _874_;
wire _875_;
wire _876_;
wire _877_;
wire _878_;
wire _879_;
wire _880_;
wire _881_;
wire _882_;
wire _883_;
wire _884_;
wire _885_;
wire _886_;
wire _887_;
wire _888_;
wire _889_;
wire _890_;
wire _891_;
wire _892_;
wire _893_;
wire _894_;
wire _895_;
wire _896_;
wire _897_;
wire _898_;
wire _899_;
wire _900_;
wire _901_;
wire _902_;
wire _903_;
wire _904_;
wire _905_;
wire _906_;
wire _907_;
wire _908_;
wire _909_;
wire _910_;
wire _911_;
wire _912_;
wire _913_;
wire _914_;
wire _915_;
wire _916_;
wire _917_;
wire _918_;
wire _919_;
wire _920_;
wire _921_;
wire _922_;
wire _923_;
wire _924_;
wire _925_;
wire _926_;
wire _927_;
wire _928_;
wire _929_;
wire _930_;
wire _931_;
wire _932_;
wire _933_;
wire _934_;
wire _935_;
wire _936_;
wire _937_;
wire _938_;
wire _939_;
wire _940_;
wire _941_;
wire _942_;
wire _943_;
wire _944_;
wire _945_;
wire _946_;
wire _947_;
wire _948_;
wire _949_;
wire _950_;
wire _951_;
wire _952_;
wire _953_;
wire _954_;
wire _955_;
wire _956_;
wire _957_;
wire _958_;
wire _959_;
wire _960_;
wire _961_;
wire _962_;
wire _963_;
wire _964_;
wire _965_;
wire _966_;
wire _967_;
wire _968_;
wire _969_;
wire _970_;
wire _971_;
wire _972_;
wire _973_;
wire _974_;
wire _975_;
wire _976_;
wire _977_;
wire _978_;
wire _979_;
wire _980_;
wire _981_;
wire _982_;
wire _983_;
wire _984_;
wire _985_;
wire _986_;
wire _987_;
wire _988_;
wire _989_;
wire _990_;
wire _991_;
wire _992_;
wire _993_;
wire _994_;
wire _995_;
wire _996_;
wire _997_;
wire _998_;
wire _999_;
wire _1000_;
wire _1001_;
wire _1002_;
wire _1003_;
wire _1004_;
wire _1005_;
wire _1006_;
wire _1007_;
wire _1008_;
wire _1009_;
wire _1010_;
wire _1011_;
wire _1012_;
wire _1013_;
wire _1014_;
wire _1015_;
wire _1016_;
wire _1017_;
wire _1018_;
wire _1019_;
wire _1020_;
wire _1021_;
wire _1022_;
wire _1023_;
wire _1024_;
wire _1025_;
wire _1026_;
wire _1027_;
wire _1028_;
wire _1029_;
wire _1030_;
wire _1031_;
wire _1032_;
wire _1033_;
wire _1034_;
wire _1035_;
wire _1036_;
wire _1037_;
wire _1038_;
wire _1039_;
wire _1040_;
wire _1041_;
wire _1042_;
wire _1043_;
wire _1044_;
wire _1045_;
wire _1046_;
wire _1047_;
wire _1048_;
wire _1049_;
wire _1050_;
wire _1051_;
wire _1052_;
wire _1053_;
wire _1054_;
wire _1055_;
wire _1056_;
wire _1057_;
wire _1058_;
wire _1059_;
wire _1060_;
wire _1061_;
wire _1062_;
wire _1063_;
wire _1064_;
wire _1065_;
wire _1066_;
wire _1067_;
wire _1068_;
wire _1069_;
wire _1070_;
wire _1071_;
wire _1072_;
wire _1073_;
wire _1074_;
wire _1075_;
wire _1076_;
wire _1077_;
wire _1078_;
wire _1079_;
wire _1080_;
wire _1081_;
wire _1082_;
wire _1083_;
wire _1084_;
wire _1085_;
wire _1086_;
wire _1087_;
wire _1088_;
wire _1089_;
wire _1090_;
wire _1091_;
wire _1092_;
wire _1093_;
wire _1094_;
wire _1095_;
wire _1096_;
wire _1097_;
wire _1098_;
wire _1099_;
wire _1100_;
wire _1101_;
wire _1102_;
wire _1103_;
wire _1104_;
wire _1105_;
wire _1106_;
wire _1107_;
wire _1108_;
wire _1109_;
wire _1110_;
wire _1111_;
wire _1112_;
wire _1113_;
wire _1114_;
wire _1115_;
wire _1116_;
wire _1117_;
wire _1118_;
wire _1119_;
wire _1120_;
wire _1121_;
wire _1122_;
wire _1123_;
wire _1124_;
wire _1125_;
wire _1126_;
wire _1127_;
wire _1128_;
wire _1129_;
wire _1130_;
wire _1131_;
wire _1132_;
wire _1133_;
wire _1134_;
wire _1135_;
wire _1136_;
wire _1137_;
wire _1138_;
wire _1139_;
wire _1140_;
wire _1141_;
wire _1142_;
wire _1143_;
wire _1144_;
wire _1145_;
wire _1146_;
wire _1147_;
wire _1148_;
wire _1149_;
wire _1150_;
wire _1151_;
wire _1152_;
wire _1153_;
wire _1154_;
wire _1155_;
wire _1156_;
wire _1157_;
wire _1158_;
wire _1159_;
wire _1160_;
wire _1161_;
wire _1162_;
wire _1163_;
wire _1164_;
wire _1165_;
wire _1166_;
wire _1167_;
wire _1168_;
wire _1169_;
wire _1170_;
wire _1171_;
wire _1172_;
wire _1173_;
wire _1174_;
wire _1175_;
wire _1176_;
wire _1177_;
wire _1178_;
wire _1179_;
wire _1180_;
wire _1181_;
wire _1182_;
wire _1183_;
wire _1184_;
wire _1185_;
wire _1186_;
wire _1187_;
wire _1188_;
wire _1189_;
wire _1190_;
wire _1191_;
wire _1192_;
wire _1193_;
wire _1194_;
wire _1195_;
wire _1196_;
wire _1197_;
wire _1198_;
wire _1199_;
wire _1200_;
wire _1201_;
wire _1202_;
wire _1203_;
wire _1204_;
wire _1205_;
wire _1206_;
wire _1207_;
wire _1208_;
wire _1209_;
wire _1210_;
wire _1211_;
wire _1212_;
wire _1213_;
wire _1214_;
wire _1215_;
wire _1216_;
wire _1217_;
wire _1218_;
wire _1219_;
wire _1220_;
wire _1221_;
wire _1222_;
wire _1223_;
wire _1224_;
wire _1225_;
wire _1226_;
wire _1227_;
wire _1228_;
wire _1229_;
wire _1230_;
wire _1231_;
wire _1232_;
wire _1233_;
wire _1234_;
wire _1235_;
wire _1236_;
wire _1237_;
wire _1238_;
wire _1239_;
wire _1240_;
wire _1241_;
wire _1242_;
wire _1243_;
wire _1244_;
wire _1245_;
wire _1246_;
wire _1247_;
wire _1248_;
wire _1249_;
wire _1250_;
wire _1251_;
wire _1252_;
wire _1253_;
wire _1254_;
wire _1255_;
wire _1256_;
wire _1257_;
wire _1258_;
wire _1259_;
wire _1260_;
wire _1261_;
wire _1262_;
wire _1263_;
wire _1264_;
wire _1265_;
wire _1266_;
wire _1267_;
wire _1268_;
wire _1269_;
wire _1270_;
wire _1271_;
wire _1272_;
wire _1273_;
wire _1274_;
wire _1275_;
wire _1276_;
wire _1277_;
wire _1278_;
wire _1279_;
wire _1280_;
wire _1281_;
wire _1282_;
wire _1283_;
wire _1284_;
wire _1285_;
wire _1286_;
wire _1287_;
wire _1288_;
wire _1289_;
wire _1290_;
wire _1291_;
wire _1292_;
wire _1293_;
wire _1294_;
wire _1295_;
wire _1296_;
wire _1297_;
wire _1298_;
wire _1299_;
wire _1300_;
wire _1301_;
wire _1302_;
wire _1303_;
wire _1304_;
wire _1305_;
wire _1306_;
wire _1307_;
wire _1308_;
wire _1309_;
wire _1310_;
wire _1311_;
wire _1312_;
wire _1313_;
wire _1314_;
wire _1315_;
wire _1316_;
wire _1317_;
wire _1318_;
wire _1319_;
wire _1320_;
wire _1321_;
wire _1322_;
wire _1323_;
wire _1324_;
wire _1325_;
wire _1326_;
wire _1327_;
wire _1328_;
wire _1329_;
wire _1330_;
wire _1331_;
wire _1332_;
wire _1333_;
wire _1334_;
wire _1335_;
wire _1336_;
wire _1337_;
wire _1338_;
wire _1339_;
wire _1340_;
wire _1341_;
wire _1342_;
wire _1343_;
wire _1344_;
wire _1345_;
wire _1346_;
wire _1347_;
wire _1348_;
wire _1349_;
wire _1350_;
wire _1351_;
wire _1352_;
wire _1353_;
wire _1354_;
wire _1355_;
wire _1356_;
wire _1357_;
wire _1358_;
wire _1359_;
wire _1360_;
wire _1361_;
wire _1362_;
wire _1363_;
wire _1364_;
wire _1365_;
wire _1366_;
wire _1367_;
wire _1368_;
wire _1369_;
wire _1370_;
wire _1371_;
wire _1372_;
wire _1373_;
wire _1374_;
wire _1375_;
wire _1376_;
wire _1377_;
wire _1378_;
wire _1379_;
wire _1380_;
wire _1381_;
wire _1382_;
wire _1383_;
wire _1384_;
wire _1385_;
wire _1386_;
wire _1387_;
wire _1388_;
wire _1389_;
wire _1390_;
wire _1391_;
wire _1392_;
wire _1393_;
wire _1394_;
wire _1395_;
wire _1396_;
wire _1397_;
wire _1398_;
wire _1399_;
wire _1400_;
wire _1401_;
wire _1402_;
wire _1403_;
wire _1404_;
wire _1405_;
wire _1406_;
wire _1407_;
wire _1408_;
wire _1409_;
wire _1410_;
wire _1411_;
wire _1412_;
wire _1413_;
wire _1414_;
wire _1415_;
wire _1416_;
wire _1417_;
wire _1418_;
wire _1419_;
wire _1420_;
wire _1421_;
wire _1422_;
wire _1423_;
wire _1424_;
wire _1425_;
wire _1426_;
wire _1427_;
wire _1428_;
wire _1429_;
wire _1430_;
wire _1431_;
wire _1432_;
wire _1433_;
wire _1434_;
wire _1435_;
wire _1436_;
wire _1437_;
wire _1438_;
wire _1439_;
wire _1440_;
wire _1441_;
wire _1442_;
wire _1443_;
wire _1444_;
wire _1445_;
wire _1446_;
wire _1447_;
wire _1448_;
wire _1449_;
wire _1450_;
wire _1451_;
wire _1452_;
wire _1453_;
wire _1454_;
wire _1455_;
wire _1456_;
wire _1457_;
wire _1458_;
wire _1459_;
wire _1460_;
wire _1461_;
wire _1462_;
wire _1463_;
wire _1464_;
wire _1465_;
wire _1466_;
wire _1467_;
wire _1468_;
wire _1469_;
wire _1470_;
wire _1471_;
wire _1472_;
wire _1473_;
wire _1474_;
wire _1475_;
wire _1476_;
wire _1477_;
wire _1478_;
wire _1479_;
wire _1480_;
wire _1481_;
wire _1482_;
wire _1483_;
wire _1484_;
wire _1485_;
wire _1486_;
wire _1487_;
wire _1488_;
wire _1489_;
wire _1490_;
wire _1491_;
wire _1492_;
wire _1493_;
wire _1494_;
wire _1495_;
wire _1496_;
wire _1497_;
wire _1498_;
wire _1499_;
wire _1500_;
wire _1501_;
wire _1502_;
wire _1503_;
wire _1504_;
wire _1505_;
wire _1506_;
wire _1507_;
wire _1508_;
wire _1509_;
wire _1510_;
wire _1511_;
wire _1512_;
wire _1513_;
wire _1514_;
wire _1515_;
wire _1516_;
wire _1517_;
wire _1518_;
wire _1519_;
wire _1520_;
wire _1521_;
wire _1522_;
wire _1523_;
wire _1524_;
wire _1525_;
wire _1526_;
wire _1527_;
wire _1528_;
wire _1529_;
wire _1530_;
wire _1531_;
wire _1532_;
wire _1533_;
wire _1534_;
wire _1535_;
wire _1536_;
wire _1537_;
wire _1538_;
wire _1539_;
wire _1540_;
wire _1541_;
wire _1542_;
wire _1543_;
wire _1544_;
wire _1545_;
wire _1546_;
wire _1547_;
wire _1548_;
wire _1549_;
wire _1550_;
wire _1551_;
wire _1552_;
wire _1553_;
wire _1554_;
wire _1555_;
wire _1556_;
wire _1557_;
wire _1558_;
wire _1559_;
wire _1560_;
wire _1561_;
wire _1562_;
wire _1563_;
wire _1564_;
wire _1565_;
wire _1566_;
wire _1567_;
wire _1568_;
wire _1569_;
wire _1570_;
wire _1571_;
wire _1572_;
wire _1573_;
wire _1574_;
wire _1575_;
wire _1576_;
wire _1577_;
wire _1578_;
wire _1579_;
wire _1580_;
wire _1581_;
wire _1582_;
wire _1583_;
wire _1584_;
wire _1585_;
wire _1586_;
wire _1587_;
wire _1588_;
wire _1589_;
wire _1590_;
wire _1591_;
wire _1592_;
wire _1593_;
wire _1594_;
wire _1595_;
wire _1596_;
wire _1597_;
wire _1598_;
wire _1599_;
wire _1600_;
wire _1601_;
wire _1602_;
wire _1603_;
wire _1604_;
wire _1605_;
wire _1606_;
wire _1607_;
wire _1608_;
wire _1609_;
wire _1610_;
wire _1611_;
wire _1612_;
wire _1613_;
wire _1614_;
wire _1615_;
wire _1616_;
wire _1617_;
wire _1618_;
wire _1619_;
wire _1620_;
wire _1621_;
wire _1622_;
wire _1623_;
wire _1624_;
wire _1625_;
wire _1626_;
wire _1627_;
wire _1628_;
wire _1629_;
wire _1630_;
wire _1631_;
wire _1632_;
wire _1633_;
wire _1634_;
wire _1635_;
wire _1636_;
wire _1637_;
wire _1638_;
wire _1639_;
wire _1640_;
wire _1641_;
wire _1642_;
wire _1643_;
wire _1644_;
wire _1645_;
wire _1646_;
wire _1647_;
wire _1648_;
wire _1649_;
wire _1650_;
wire _1651_;
wire _1652_;
wire _1653_;
wire _1654_;
wire _1655_;
wire _1656_;
wire _1657_;
wire _1658_;
wire _1659_;
wire _1660_;
wire _1661_;
wire _1662_;
wire _1663_;
wire _1664_;
wire _1665_;
wire _1666_;
wire _1667_;
wire _1668_;
wire _1669_;
wire _1670_;
wire _1671_;
wire _1672_;
wire _1673_;
wire _1674_;
wire _1675_;
wire _1676_;
wire _1677_;
wire _1678_;
wire _1679_;
wire _1680_;
wire _1681_;
wire _1682_;
wire _1683_;
wire _1684_;
wire _1685_;
wire _1686_;
wire _1687_;
wire _1688_;
wire _1689_;
wire _1690_;
wire _1691_;
wire _1692_;
wire _1693_;
wire _1694_;
wire _1695_;
wire _1696_;
wire _1697_;
wire _1698_;
wire _1699_;
wire _1700_;
wire _1701_;
wire _1702_;
wire _1703_;
wire _1704_;
wire _1705_;
wire _1706_;
wire _1707_;
wire _1708_;
wire _1709_;
wire _1710_;
wire _1711_;
wire _1712_;
wire _1713_;
wire _1714_;
wire _1715_;
wire _1716_;
wire _1717_;
wire _1718_;
wire _1719_;
wire _1720_;
wire _1721_;
wire _1722_;
wire _1723_;
wire _1724_;
wire _1725_;
wire _1726_;
wire _1727_;
wire _1728_;
wire _1729_;
wire _1730_;
wire _1731_;
wire _1732_;
wire _1733_;
wire _1734_;
wire _1735_;
wire _1736_;
wire _1737_;
wire _1738_;
wire _1739_;
wire _1740_;
wire _1741_;
wire _1742_;
wire _1743_;
wire _1744_;
wire _1745_;
wire _1746_;
wire _1747_;
wire _1748_;
wire _1749_;
wire _1750_;
wire _1751_;
wire _1752_;
wire _1753_;
wire _1754_;
wire _1755_;
wire _1756_;
wire _1757_;
wire _1758_;
wire _1759_;
wire _1760_;
wire _1761_;
wire _1762_;
wire _1763_;
wire _1764_;
wire _1765_;
wire _1766_;
wire _1767_;
wire _1768_;
wire _1769_;
wire _1770_;
wire _1771_;
wire _1772_;
wire _1773_;
wire _1774_;
wire _1775_;
wire _1776_;
wire _1777_;
wire _1778_;
wire _1779_;
wire _1780_;
wire _1781_;
wire _1782_;
wire _1783_;
wire _1784_;
wire _1785_;
wire _1786_;
wire _1787_;
wire _1788_;
wire _1789_;
wire _1790_;
wire _1791_;
wire _1792_;
wire _1793_;
wire _1794_;
wire _1795_;
wire _1796_;
wire _1797_;
wire _1798_;
wire _1799_;
wire _1800_;
wire _1801_;
wire _1802_;
wire _1803_;
wire _1804_;
wire _1805_;
wire _1806_;
wire _1807_;
wire _1808_;
wire _1809_;
wire _1810_;
wire _1811_;
wire _1812_;
wire _1813_;
wire _1814_;
wire _1815_;
wire _1816_;
wire _1817_;
wire _1818_;
wire _1819_;
wire _1820_;
wire _1821_;
wire _1822_;
wire _1823_;
wire _1824_;
wire _1825_;
wire _1826_;
wire _1827_;
wire _1828_;
wire _1829_;
wire _1830_;
wire _1831_;
wire _1832_;
wire _1833_;
wire _1834_;
wire _1835_;
wire _1836_;
wire _1837_;
wire _1838_;
wire _1839_;
wire _1840_;
wire _1841_;
wire _1842_;
wire _1843_;
wire _1844_;
wire _1845_;
wire _1846_;
wire _1847_;
wire _1848_;
wire _1849_;
wire _1850_;
wire _1851_;
wire _1852_;
wire _1853_;
wire _1854_;
wire _1855_;
wire _1856_;
wire _1857_;
wire _1858_;
wire _1859_;
wire _1860_;
wire _1861_;
wire _1862_;
wire _1863_;
wire _1864_;
wire _1865_;
wire _1866_;
wire _1867_;
wire _1868_;
wire _1869_;
wire _1870_;
wire _1871_;
wire _1872_;
wire _1873_;
wire _1874_;
wire _1875_;
wire _1876_;
wire _1877_;
wire _1878_;
wire _1879_;
wire _1880_;
wire _1881_;
wire _1882_;
wire _1883_;
wire _1884_;
wire _1885_;
wire _1886_;
wire _1887_;
wire _1888_;
wire _1889_;
wire _1890_;
wire _1891_;
wire _1892_;
wire _1893_;
wire _1894_;
wire _1895_;
wire _1896_;
wire _1897_;
wire _1898_;
wire _1899_;
wire _1900_;
wire _1901_;
wire _1902_;
wire _1903_;
wire _1904_;
wire _1905_;
wire _1906_;
wire _1907_;
wire _1908_;
wire _1909_;
wire _1910_;
wire _1911_;
wire _1912_;
wire _1913_;
wire _1914_;
wire _1915_;
wire _1916_;
wire _1917_;
wire _1918_;
wire _1919_;
wire _1920_;
wire _1921_;
wire _1922_;
wire _1923_;
wire _1924_;
wire _1925_;
wire _1926_;
wire _1927_;
wire _1928_;
wire _1929_;
wire _1930_;
wire _1931_;
wire _1932_;
wire _1933_;
wire _1934_;
wire _1935_;
wire _1936_;
wire _1937_;
wire _1938_;
wire _1939_;
wire _1940_;
wire _1941_;
wire _1942_;
wire _1943_;
wire _1944_;
wire _1945_;
wire _1946_;
wire _1947_;
wire _1948_;
wire _1949_;
wire _1950_;
wire _1951_;
wire _1952_;
wire _1953_;
wire _1954_;
wire _1955_;
wire _1956_;
wire _1957_;
wire _1958_;
wire _1959_;
wire _1960_;
wire _1961_;
wire _1962_;
wire _1963_;
wire _1964_;
wire _1965_;
wire _1966_;
wire _1967_;
wire _1968_;
wire _1969_;
wire _1970_;
wire _1971_;
wire _1972_;
wire _1973_;
wire _1974_;
wire _1975_;
wire _1976_;
wire _1977_;
wire _1978_;
wire _1979_;
wire _1980_;
wire _1981_;
wire _1982_;
wire _1983_;
wire _1984_;
wire _1985_;
wire _1986_;
wire _1987_;
wire _1988_;
wire _1989_;
wire _1990_;
wire _1991_;
wire _1992_;
wire _1993_;
wire _1994_;
wire _1995_;
wire _1996_;
wire _1997_;
wire _1998_;
wire _1999_;
wire _2000_;
wire _2001_;
wire _2002_;
wire _2003_;
wire _2004_;
wire _2005_;
wire _2006_;
wire _2007_;
wire _2008_;
wire _2009_;
wire _2010_;
wire _2011_;
wire _2012_;
wire _2013_;
wire _2014_;
wire _2015_;
wire _2016_;
wire _2017_;
wire _2018_;
wire _2019_;
wire _2020_;
wire _2021_;
wire _2022_;
wire _2023_;
wire _2024_;
wire _2025_;
wire _2026_;
wire _2027_;
wire _2028_;
wire _2029_;
wire _2030_;
wire _2031_;
wire _2032_;
wire _2033_;
wire _2034_;
wire _2035_;
wire _2036_;
wire _2037_;
wire _2038_;
wire _2039_;
wire _2040_;
wire _2041_;
wire _2042_;
wire _2043_;
wire _2044_;
wire _2045_;
wire _2046_;
wire _2047_;
wire _2048_;
wire _2049_;
wire _2050_;
wire _2051_;
wire _2052_;
wire _2053_;
wire _2054_;
wire _2055_;
wire _2056_;
wire _2057_;
wire _2058_;
wire _2059_;
wire _2060_;
wire _2061_;
wire _2062_;
wire _2063_;
wire _2064_;
wire _2065_;
wire _2066_;
wire _2067_;
wire _2068_;
wire _2069_;
wire _2070_;
wire _2071_;
wire _2072_;
wire _2073_;
wire _2074_;
wire _2075_;
wire _2076_;
wire _2077_;
wire _2078_;
wire _2079_;
wire _2080_;
wire _2081_;
wire _2082_;
wire _2083_;
wire _2084_;
wire _2085_;
wire _2086_;
wire _2087_;
wire _2088_;
wire _2089_;
wire _2090_;
wire _2091_;
wire _2092_;
wire _2093_;
wire _2094_;
wire _2095_;
wire _2096_;
wire _2097_;
wire _2098_;
wire _2099_;
wire _2100_;
wire _2101_;
wire _2102_;
wire _2103_;
wire _2104_;
wire _2105_;
wire _2106_;
wire _2107_;
wire _2108_;
wire _2109_;
wire _2110_;
wire _2111_;
wire _2112_;
wire _2113_;
wire _2114_;
wire _2115_;
wire _2116_;
wire _2117_;
wire _2118_;
wire _2119_;
wire _2120_;
wire _2121_;
wire _2122_;
wire _2123_;
wire _2124_;
wire _2125_;
wire _2126_;
wire _2127_;
wire _2128_;
wire _2129_;
wire _2130_;
wire _2131_;
wire _2132_;
wire _2133_;
wire _2134_;
wire _2135_;
wire _2136_;
wire _2137_;
wire _2138_;
wire _2139_;
wire _2140_;
wire _2141_;
wire _2142_;
wire _2143_;
wire _2144_;
wire _2145_;
wire _2146_;
wire _2147_;
wire _2148_;
wire _2149_;
wire _2150_;
wire _2151_;
wire _2152_;
wire _2153_;
wire _2154_;
wire _2155_;
wire _2156_;
wire _2157_;
wire _2158_;
wire _2159_;
wire _2160_;
wire _2161_;
wire _2162_;
wire _2163_;
wire _2164_;
wire _2165_;
wire _2166_;
wire _2167_;
wire _2168_;
wire _2169_;
wire _2170_;
wire _2171_;
wire _2172_;
wire _2173_;
wire _2174_;
wire _2175_;
wire _2176_;
wire _2177_;
wire _2178_;
wire _2179_;
wire _2180_;
wire _2181_;
wire _2182_;
wire _2183_;
wire _2184_;
wire _2185_;
wire _2186_;
wire _2187_;
wire _2188_;
wire _2189_;
wire _2190_;
wire _2191_;
wire _2192_;
wire _2193_;
wire _2194_;
wire _2195_;
wire _2196_;
wire _2197_;
wire _2198_;
wire _2199_;
wire _2200_;
wire _2201_;
wire _2202_;
wire _2203_;
wire _2204_;
wire _2205_;
wire _2206_;
wire _2207_;
wire _2208_;
wire _2209_;
wire _2210_;
wire _2211_;
wire _2212_;
wire _2213_;
wire _2214_;
wire _2215_;
wire _2216_;
wire _2217_;
wire _2218_;
wire _2219_;
wire _2220_;
wire _2221_;
wire _2222_;
wire _2223_;
wire _2224_;
wire _2225_;
wire _2226_;
wire _2227_;
wire _2228_;
wire _2229_;
wire _2230_;
wire _2231_;
wire _2232_;
wire _2233_;
wire _2234_;
wire _2235_;
wire _2236_;
wire _2237_;
wire _2238_;
wire _2239_;
wire _2240_;
wire _2241_;
wire _2242_;
wire _2243_;
wire _2244_;
wire _2245_;
wire _2246_;
wire _2247_;
wire _2248_;
wire _2249_;
wire _2250_;
wire _2251_;
wire _2252_;
wire _2253_;
wire _2254_;
wire _2255_;
wire _2256_;
wire _2257_;
wire _2258_;
wire _2259_;
wire _2260_;
wire _2261_;
wire _2262_;
wire _2263_;
wire _2264_;
wire _2265_;
wire _2266_;
wire _2267_;
wire _2268_;
wire _2269_;
wire _2270_;
wire _2271_;
wire _2272_;
wire _2273_;
wire _2274_;
wire _2275_;
wire _2276_;
wire _2277_;
wire _2278_;
wire _2279_;
wire _2280_;
wire _2281_;
wire _2282_;
wire _2283_;
wire _2284_;
wire _2285_;
wire _2286_;
wire _2287_;
wire _2288_;
wire _2289_;
wire _2290_;
wire _2291_;
wire _2292_;
wire _2293_;
wire _2294_;
wire _2295_;
wire _2296_;
wire _2297_;
wire _2298_;
wire _2299_;
wire _2300_;
wire _2301_;
wire _2302_;
wire _2303_;
wire _2304_;
wire _2305_;
wire _2306_;
wire _2307_;
wire _2308_;
wire _2309_;
wire _2310_;
wire _2311_;
wire _2312_;
wire _2313_;
wire _2314_;
wire _2315_;
wire _2316_;
wire _2317_;
wire _2318_;
wire _2319_;
wire _2320_;
wire _2321_;
wire _2322_;
wire _2323_;
wire _2324_;
wire _2325_;
wire _2326_;
wire _2327_;
wire _2328_;
wire _2329_;
wire _2330_;
wire _2331_;
wire _2332_;
wire _2333_;
wire _2334_;
wire _2335_;
wire _2336_;
wire _2337_;
wire _2338_;
wire _2339_;
wire _2340_;
wire _2341_;
wire _2342_;
wire _2343_;
wire _2344_;
wire _2345_;
wire _2346_;
wire _2347_;
wire _2348_;
wire _2349_;
wire _2350_;
wire _2351_;
wire _2352_;
wire _2353_;
wire _2354_;
wire _2355_;
wire _2356_;
wire _2357_;
wire _2358_;
wire _2359_;
wire _2360_;
wire _2361_;
wire _2362_;
wire _2363_;
wire _2364_;
wire _2365_;
wire _2366_;
wire _2367_;
wire _2368_;
wire _2369_;
wire _2370_;
wire _2371_;
wire _2372_;
wire _2373_;
wire _2374_;
wire _2375_;
wire _2376_;
wire _2377_;
wire _2378_;
wire _2379_;
wire _2380_;
wire _2381_;
wire _2382_;
wire _2383_;
wire _2384_;
wire _2385_;
wire _2386_;
wire _2387_;
wire _2388_;
wire _2389_;
wire _2390_;
wire _2391_;
wire _2392_;
wire _2393_;
wire _2394_;
wire _2395_;
wire _2396_;
wire _2397_;
wire _2398_;
wire _2399_;
wire _2400_;
wire _2401_;
wire _2402_;
wire _2403_;
wire _2404_;
wire _2405_;
wire _2406_;
wire _2407_;
wire _2408_;
wire _2409_;
wire _2410_;
wire _2411_;
wire _2412_;
wire _2413_;
wire _2414_;
wire _2415_;
wire _2416_;
wire _2417_;
wire _2418_;
wire _2419_;
wire _2420_;
wire _2421_;
wire _2422_;
wire _2423_;
wire _2424_;
wire _2425_;
wire _2426_;
wire _2427_;
wire _2428_;
wire _2429_;
wire _2430_;
wire _2431_;
wire _2432_;
wire _2433_;
wire _2434_;
wire _2435_;
wire _2436_;
wire _2437_;
wire _2438_;
wire _2439_;
wire _2440_;
wire _2441_;
wire _2442_;
wire _2443_;
wire _2444_;
wire _2445_;
wire _2446_;
wire _2447_;
wire _2448_;
wire _2449_;
wire _2450_;
wire _2451_;
wire _2452_;
wire _2453_;
wire _2454_;
wire _2455_;
wire _2456_;
wire _2457_;
wire _2458_;
wire _2459_;
wire _2460_;
wire _2461_;
wire _2462_;
wire _2463_;
wire _2464_;
wire _2465_;
wire _2466_;
wire _2467_;
wire _2468_;
wire _2469_;
wire _2470_;
wire _2471_;
wire _2472_;
wire _2473_;
wire _2474_;
wire _2475_;
wire _2476_;
wire _2477_;
wire _2478_;
wire _2479_;
wire _2480_;
wire _2481_;
wire _2482_;
wire _2483_;
wire _2484_;
wire _2485_;
wire _2486_;
wire _2487_;
wire _2488_;
wire _2489_;
wire _2490_;
wire _2491_;
wire _2492_;
wire _2493_;
wire _2494_;
wire _2495_;
wire _2496_;
wire _2497_;
wire _2498_;
wire _2499_;
wire _2500_;
wire _2501_;
wire _2502_;
wire _2503_;
wire _2504_;
wire _2505_;
wire _2506_;
wire _2507_;
wire _2508_;
wire _2509_;
wire _2510_;
wire _2511_;
wire _2512_;
wire _2513_;
wire _2514_;
wire _2515_;
wire _2516_;
wire _2517_;
wire _2518_;
wire _2519_;
wire _2520_;
wire _2521_;
wire _2522_;
wire _2523_;
wire _2524_;
wire _2525_;
wire _2526_;
wire _2527_;
wire _2528_;
wire _2529_;
wire _2530_;
wire _2531_;
wire _2532_;
wire _2533_;
wire _2534_;
wire _2535_;
wire _2536_;
wire _2537_;
wire _2538_;
wire _2539_;
wire _2540_;
wire _2541_;
wire _2542_;
wire _2543_;
wire _2544_;
wire _2545_;
wire _2546_;
wire _2547_;
wire _2548_;
wire _2549_;
wire _2550_;
wire _2551_;
wire _2552_;
wire _2553_;
wire _2554_;
wire _2555_;
wire _2556_;
wire _2557_;
wire _2558_;
wire _2559_;
wire _2560_;
wire _2561_;
wire _2562_;
wire _2563_;
wire _2564_;
wire _2565_;
wire _2566_;
wire _2567_;
wire _2568_;
wire _2569_;
wire _2570_;
wire _2571_;
wire _2572_;
wire _2573_;
wire _2574_;
wire _2575_;
wire _2576_;
wire _2577_;
wire _2578_;
wire _2579_;
wire _2580_;
wire _2581_;
wire _2582_;
wire _2583_;
wire _2584_;
wire _2585_;
wire _2586_;
wire _2587_;
wire _2588_;
wire _2589_;
wire _2590_;
wire _2591_;
wire _2592_;
wire _2593_;
wire _2594_;
wire _2595_;
wire _2596_;
wire _2597_;
wire _2598_;
wire _2599_;
wire _2600_;
wire _2601_;
wire _2602_;
wire _2603_;
wire _2604_;
wire _2605_;
wire _2606_;
wire _2607_;
wire _2608_;
wire _2609_;
wire _2610_;
wire _2611_;
wire _2612_;
wire _2613_;
wire _2614_;
wire _2615_;
wire _2616_;
wire _2617_;
wire _2618_;
wire _2619_;
wire _2620_;
wire _2621_;
wire _2622_;
wire _2623_;
wire _2624_;
wire _2625_;
wire _2626_;
wire _2627_;
wire _2628_;
wire _2629_;
wire _2630_;
wire _2631_;
wire _2632_;
wire _2633_;
wire _2634_;
wire _2635_;
wire _2636_;
wire _2637_;
wire _2638_;
wire _2639_;
wire _2640_;
wire _2641_;
wire _2642_;
wire _2643_;
wire _2644_;
wire _2645_;
wire _2646_;
wire _2647_;
wire _2648_;
wire _2649_;
wire _2650_;
wire _2651_;
wire _2652_;
wire _2653_;
wire _2654_;
wire _2655_;
wire _2656_;
wire _2657_;
wire _2658_;
wire _2659_;
wire _2660_;
wire _2661_;
wire _2662_;
wire _2663_;
wire _2664_;
wire _2665_;
wire _2666_;
wire _2667_;
wire _2668_;
wire _2669_;
wire _2670_;
wire _2671_;
wire _2672_;
wire _2673_;
wire _2674_;
wire _2675_;
wire _2676_;
wire _2677_;
wire _2678_;
wire _2679_;
wire _2680_;
wire _2681_;
wire _2682_;
wire _2683_;
wire _2684_;
wire _2685_;
wire _2686_;
wire _2687_;
wire _2688_;
wire _2689_;
wire _2690_;
wire _2691_;
wire _2692_;
wire _2693_;
wire _2694_;
wire _2695_;
wire _2696_;
wire _2697_;
wire _2698_;
wire _2699_;
wire _2700_;
wire _2701_;
wire _2702_;
wire _2703_;
wire _2704_;
wire _2705_;
wire _2706_;
wire _2707_;
wire _2708_;
wire _2709_;
wire _2710_;
wire _2711_;
wire _2712_;
wire _2713_;
wire _2714_;
wire _2715_;
wire _2716_;
wire _2717_;
wire _2718_;
wire _2719_;
wire _2720_;
wire _2721_;
wire _2722_;
wire _2723_;
wire _2724_;
wire _2725_;
wire _2726_;
wire _2727_;
wire _2728_;
wire _2729_;
wire _2730_;
wire _2731_;
wire _2732_;
wire _2733_;
wire _2734_;
wire _2735_;
wire _2736_;
wire _2737_;
wire _2738_;
wire _2739_;
wire _2740_;
wire _2741_;
wire _2742_;
wire _2743_;
wire _2744_;
wire _2745_;
wire _2746_;
wire _2747_;
wire _2748_;
wire _2749_;
wire _2750_;
wire _2751_;
wire _2752_;
wire _2753_;
wire _2754_;
wire _2755_;
wire _2756_;
wire _2757_;
wire _2758_;
wire _2759_;
wire _2760_;
wire _2761_;
wire _2762_;
wire _2763_;
wire _2764_;
wire _2765_;
wire _2766_;
wire _2767_;
wire _2768_;
wire _2769_;
wire _2770_;
wire _2771_;
wire _2772_;
wire _2773_;
wire _2774_;
wire _2775_;
wire _2776_;
wire _2777_;
wire _2778_;
wire _2779_;
wire _2780_;
wire _2781_;
wire _2782_;
wire _2783_;
wire _2784_;
wire _2785_;
wire _2786_;
wire _2787_;
wire _2788_;
wire _2789_;
wire _2790_;
wire _2791_;
wire _2792_;
wire _2793_;
wire _2794_;
wire _2795_;
wire _2796_;
wire _2797_;
wire _2798_;
wire _2799_;
wire _2800_;
wire _2801_;
wire _2802_;
wire _2803_;
wire _2804_;
wire _2805_;
wire _2806_;
wire _2807_;
wire _2808_;
wire _2809_;
wire _2810_;
wire _2811_;
wire _2812_;
wire _2813_;
wire _2814_;
wire _2815_;
wire _2816_;
wire _2817_;
wire _2818_;
wire _2819_;
wire _2820_;
wire _2821_;
wire _2822_;
wire _2823_;
wire _2824_;
wire _2825_;
wire _2826_;
wire _2827_;
wire _2828_;
wire _2829_;
wire _2830_;
wire _2831_;
wire _2832_;
wire _2833_;
wire _2834_;
wire _2835_;
wire _2836_;
wire _2837_;
wire _2838_;
wire _2839_;
wire _2840_;
wire _2841_;
wire _2842_;
wire _2843_;
wire _2844_;
wire _2845_;
wire _2846_;
wire _2847_;
wire _2848_;
wire _2849_;
wire _2850_;
wire _2851_;
wire _2852_;
wire _2853_;
wire _2854_;
wire _2855_;
wire _2856_;
wire _2857_;
wire _2858_;
wire _2859_;
wire _2860_;
wire _2861_;
wire _2862_;
wire _2863_;
wire _2864_;
wire _2865_;
wire _2866_;
wire _2867_;
wire _2868_;
wire _2869_;
wire _2870_;
wire _2871_;
wire _2872_;
wire _2873_;
wire _2874_;
wire _2875_;
wire _2876_;
wire _2877_;
wire _2878_;
wire _2879_;
wire _2880_;
wire _2881_;
wire _2882_;
wire _2883_;
wire _2884_;
wire _2885_;
wire _2886_;
wire _2887_;
wire _2888_;
wire _2889_;
wire _2890_;
wire _2891_;
wire _2892_;
wire _2893_;
wire _2894_;
wire _2895_;
wire _2896_;
wire _2897_;
wire _2898_;
wire _2899_;
wire _2900_;
wire _2901_;
wire _2902_;
wire _2903_;
wire _2904_;
wire _2905_;
wire _2906_;
wire _2907_;
wire _2908_;
wire _2909_;
wire _2910_;
wire _2911_;
wire _2912_;
wire _2913_;
wire _2914_;
wire _2915_;
wire _2916_;
wire _2917_;
wire _2918_;
wire _2919_;
wire _2920_;
wire _2921_;
wire _2922_;
wire _2923_;
wire _2924_;
wire _2925_;
wire _2926_;
wire _2927_;
wire _2928_;
wire _2929_;
wire _2930_;
wire _2931_;
wire _2932_;
wire _2933_;
wire _2934_;
wire _2935_;
wire _2936_;
wire _2937_;
wire _2938_;
wire _2939_;
wire _2940_;
wire _2941_;
wire _2942_;
wire _2943_;
wire _2944_;
wire _2945_;
wire _2946_;
wire _2947_;
wire _2948_;
wire _2949_;
wire _2950_;
wire _2951_;
wire _2952_;
wire _2953_;
wire _2954_;
wire _2955_;
wire _2956_;
wire _2957_;
wire _2958_;
wire _2959_;
wire _2960_;
wire _2961_;
wire _2962_;
wire _2963_;
wire _2964_;
wire _2965_;
wire _2966_;
wire _2967_;
wire _2968_;
wire _2969_;
wire _2970_;
wire _2971_;
wire _2972_;
wire _2973_;
wire _2974_;
wire _2975_;
wire _2976_;
wire _2977_;
wire _2978_;
wire _2979_;
wire _2980_;
wire _2981_;
wire _2982_;
wire _2983_;
wire _2984_;
wire _2985_;
wire _2986_;
wire _2987_;
wire _2988_;
wire _2989_;
wire _2990_;
wire _2991_;
wire _2992_;
wire _2993_;
wire _2994_;
wire _2995_;
wire _2996_;
wire _2997_;
wire _2998_;
wire _2999_;
wire _3000_;
wire _3001_;
wire _3002_;
wire _3003_;
wire _3004_;
wire _3005_;
wire _3006_;
wire _3007_;
wire _3008_;
wire _3009_;
wire _3010_;
wire _3011_;
wire _3012_;
wire _3013_;
wire _3014_;
wire _3015_;
wire _3016_;
wire _3017_;
wire _3018_;
wire _3019_;
wire _3020_;
wire _3021_;
wire _3022_;
wire _3023_;
wire _3024_;
wire _3025_;
wire _3026_;
wire _3027_;
wire _3028_;
wire _3029_;
wire _3030_;
wire _3031_;
wire _3032_;
wire _3033_;
wire _3034_;
wire _3035_;
wire _3036_;
wire _3037_;
wire _3038_;
wire _3039_;
wire _3040_;
wire _3041_;
wire _3042_;
wire _3043_;
wire _3044_;
wire _3045_;
wire _3046_;
wire _3047_;
wire _3048_;
wire _3049_;
wire _3050_;
wire _3051_;
wire _3052_;
wire _3053_;
wire _3054_;
wire _3055_;
wire _3056_;
wire _3057_;
wire _3058_;
wire _3059_;
wire _3060_;
wire _3061_;
wire _3062_;
wire _3063_;
wire _3064_;
wire _3065_;
wire _3066_;
wire _3067_;
wire _3068_;
wire _3069_;
wire _3070_;
wire _3071_;
wire _3072_;
wire _3073_;
wire _3074_;
wire _3075_;
wire _3076_;
wire _3077_;
wire _3078_;
wire _3079_;
wire _3080_;
wire _3081_;
wire _3082_;
wire _3083_;
wire _3084_;
wire _3085_;
wire _3086_;
wire _3087_;
wire _3088_;
wire _3089_;
wire _3090_;
wire _3091_;
wire _3092_;
wire _3093_;
wire _3094_;
wire _3095_;
wire _3096_;
wire _3097_;
wire _3098_;
wire _3099_;
wire _3100_;
wire _3101_;
wire _3102_;
wire _3103_;
wire _3104_;
wire _3105_;
wire _3106_;
wire _3107_;
wire _3108_;
wire _3109_;
wire _3110_;
wire _3111_;
wire _3112_;
wire _3113_;
wire _3114_;
wire _3115_;
wire _3116_;
wire _3117_;
wire _3118_;
wire _3119_;
wire _3120_;
wire _3121_;
wire _3122_;
wire _3123_;
wire _3124_;
wire _3125_;
wire _3126_;
wire _3127_;
wire _3128_;
wire _3129_;
wire _3130_;
wire _3131_;
wire _3132_;
wire _3133_;
wire _3134_;
wire _3135_;
wire _3136_;
wire _3137_;
wire _3138_;
wire _3139_;
wire _3140_;
wire _3141_;
wire _3142_;
wire _3143_;
wire _3144_;
wire _3145_;
wire _3146_;
wire _3147_;
wire _3148_;
wire _3149_;
wire _3150_;
wire _3151_;
wire _3152_;
wire _3153_;
wire _3154_;
wire _3155_;
wire _3156_;
wire _3157_;
wire _3158_;
wire _3159_;
wire _3160_;
wire _3161_;
wire _3162_;
wire _3163_;
wire _3164_;
wire _3165_;
wire _3166_;
wire _3167_;
wire _3168_;
wire _3169_;
wire _3170_;
wire _3171_;
wire _3172_;
wire _3173_;
wire _3174_;
wire _3175_;
wire _3176_;
wire _3177_;
wire _3178_;
wire _3179_;
wire _3180_;
wire _3181_;
wire _3182_;
wire _3183_;
wire _3184_;
wire _3185_;
wire _3186_;
wire _3187_;
wire _3188_;
wire _3189_;
wire _3190_;
wire _3191_;
wire _3192_;
wire _3193_;
wire _3194_;
wire _3195_;
wire _3196_;
wire _3197_;
wire _3198_;
wire _3199_;
wire _3200_;
wire _3201_;
wire _3202_;
wire _3203_;
wire _3204_;
wire _3205_;
wire _3206_;
wire _3207_;
wire _3208_;
wire _3209_;
wire _3210_;
wire _3211_;
wire _3212_;
wire _3213_;
wire _3214_;
wire _3215_;
wire _3216_;
wire _3217_;
wire _3218_;
wire _3219_;
wire _3220_;
wire _3221_;
wire _3222_;
wire _3223_;
wire _3224_;
wire _3225_;
wire _3226_;
wire _3227_;
wire _3228_;
wire _3229_;
wire _3230_;
wire _3231_;
wire _3232_;
wire _3233_;
wire _3234_;
wire _3235_;
wire _3236_;
wire _3237_;
wire _3238_;
wire _3239_;
wire _3240_;
wire _3241_;
wire _3242_;
wire _3243_;
wire _3244_;
wire _3245_;
wire _3246_;
wire _3247_;
wire _3248_;
wire _3249_;
wire _3250_;
wire _3251_;
wire _3252_;
wire _3253_;
wire _3254_;
wire _3255_;
wire _3256_;
wire _3257_;
wire _3258_;
wire _3259_;
wire _3260_;
wire _3261_;
wire _3262_;
wire _3263_;
wire _3264_;
wire _3265_;
wire _3266_;
wire _3267_;
wire _3268_;
wire _3269_;
wire _3270_;
wire _3271_;
wire _3272_;
wire _3273_;
wire _3274_;
wire _3275_;
wire _3276_;
wire _3277_;
wire _3278_;
wire _3279_;
wire _3280_;
wire _3281_;
wire _3282_;
wire _3283_;
wire _3284_;
wire _3285_;
wire _3286_;
wire _3287_;
wire _3288_;
wire _3289_;
wire _3290_;
wire _3291_;
wire _3292_;
wire _3293_;
wire _3294_;
wire _3295_;
wire _3296_;
wire _3297_;
wire _3298_;
wire _3299_;
wire _3300_;
wire _3301_;
wire _3302_;
wire _3303_;
wire _3304_;
wire _3305_;
wire _3306_;
wire _3307_;
wire _3308_;
wire _3309_;
wire _3310_;
wire _3311_;
wire _3312_;
wire _3313_;
wire _3314_;
wire _3315_;
wire _3316_;
wire _3317_;
wire _3318_;
wire _3319_;
wire _3320_;
wire _3321_;
wire _3322_;
wire _3323_;
wire _3324_;
wire _3325_;
wire _3326_;
wire _3327_;
wire _3328_;
wire _3329_;
wire _3330_;
wire _3331_;
wire _3332_;
wire _3333_;
wire _3334_;
wire _3335_;
wire _3336_;
wire _3337_;
wire _3338_;
wire _3339_;
wire _3340_;
wire _3341_;
wire _3342_;
wire _3343_;
wire _3344_;
wire _3345_;
wire _3346_;
wire _3347_;
wire _3348_;
wire _3349_;
wire _3350_;
wire _3351_;
wire _3352_;
wire _3353_;
wire _3354_;
wire _3355_;
wire _3356_;
wire _3357_;
wire _3358_;
wire _3359_;
wire _3360_;
wire _3361_;
wire _3362_;
wire _3363_;
wire _3364_;
wire _3365_;
wire _3366_;
wire _3367_;
wire _3368_;
wire _3369_;
wire _3370_;
wire _3371_;
wire _3372_;
wire _3373_;
wire _3374_;
wire _3375_;
wire _3376_;
wire _3377_;
wire _3378_;
wire _3379_;
wire _3380_;
wire _3381_;
wire _3382_;
wire _3383_;
wire _3384_;
wire _3385_;
wire _3386_;
wire _3387_;
wire _3388_;
wire _3389_;
wire _3390_;
wire _3391_;
wire _3392_;
wire _3393_;
wire _3394_;
wire _3395_;
wire _3396_;
wire _3397_;
wire _3398_;
wire _3399_;
wire _3400_;
wire _3401_;
wire _3402_;
wire _3403_;
wire _3404_;
wire _3405_;
wire _3406_;
wire _3407_;
wire _3408_;
wire _3409_;
wire _3410_;
wire _3411_;
wire _3412_;
wire _3413_;
wire _3414_;
wire _3415_;
wire _3416_;
wire _3417_;
wire _3418_;
wire _3419_;
wire _3420_;
wire _3421_;
wire _3422_;
wire _3423_;
wire _3424_;
wire _3425_;
wire _3426_;
wire _3427_;
wire _3428_;
wire _3429_;
wire _3430_;
wire _3431_;
wire _3432_;
wire _3433_;
wire _3434_;
wire _3435_;
wire _3436_;
wire _3437_;
wire _3438_;
wire _3439_;
wire _3440_;
wire _3441_;
wire _3442_;
wire _3443_;
wire _3444_;
wire _3445_;
wire _3446_;
wire _3447_;
wire _3448_;
wire _3449_;
wire _3450_;
wire _3451_;
wire _3452_;
wire _3453_;
wire _3454_;
wire _3455_;
wire _3456_;
wire _3457_;
wire _3458_;
wire _3459_;
wire _3460_;
wire _3461_;
wire _3462_;
wire _3463_;
wire _3464_;
wire _3465_;
wire _3466_;
wire _3467_;
wire _3468_;
wire _3469_;
wire _3470_;
wire _3471_;
wire _3472_;
wire _3473_;
wire _3474_;
wire _3475_;
wire _3476_;
wire _3477_;
wire _3478_;
wire _3479_;
wire _3480_;
wire _3481_;
wire _3482_;
wire _3483_;
wire _3484_;
wire _3485_;
wire _3486_;
wire _3487_;
wire _3488_;
wire _3489_;
wire _3490_;
wire _3491_;
wire _3492_;
wire _3493_;
wire _3494_;
wire _3495_;
wire _3496_;
wire _3497_;
wire _3498_;
wire _3499_;
wire _3500_;
wire _3501_;
wire _3502_;
wire _3503_;
wire _3504_;
wire _3505_;
wire _3506_;
wire _3507_;
wire _3508_;
wire _3509_;
wire _3510_;
wire _3511_;
wire _3512_;
wire _3513_;
wire _3514_;
wire _3515_;
wire _3516_;
wire _3517_;
wire _3518_;
wire _3519_;
wire _3520_;
wire _3521_;
wire _3522_;
wire _3523_;
wire _3524_;
wire _3525_;
wire _3526_;
wire _3527_;
wire _3528_;
wire _3529_;
wire _3530_;
wire _3531_;
wire _3532_;
wire _3533_;
wire _3534_;
wire _3535_;
wire _3536_;
wire _3537_;
wire _3538_;
wire _3539_;
wire _3540_;
wire _3541_;
wire _3542_;
wire _3543_;
wire _3544_;
wire _3545_;
wire _3546_;
wire _3547_;
wire _3548_;
wire _3549_;
wire _3550_;
wire _3551_;
wire _3552_;
wire _3553_;
wire _3554_;
wire _3555_;
wire _3556_;
wire _3557_;
wire _3558_;
wire _3559_;
wire _3560_;
wire _3561_;
wire _3562_;
wire _3563_;
wire _3564_;
wire _3565_;
wire _3566_;
wire _3567_;
wire _3568_;
wire _3569_;
wire _3570_;
wire _3571_;
wire _3572_;
wire _3573_;
wire _3574_;
wire _3575_;
wire _3576_;
wire _3577_;
wire _3578_;
wire _3579_;
wire _3580_;
wire _3581_;
wire _3582_;
wire _3583_;
wire _3584_;
wire _3585_;
wire _3586_;
wire _3587_;
wire _3588_;
wire _3589_;
wire _3590_;
wire _3591_;
wire _3592_;
wire _3593_;
wire _3594_;
wire _3595_;
wire _3596_;
wire _3597_;
wire _3598_;
wire _3599_;
wire _3600_;
wire _3601_;
wire _3602_;
wire _3603_;
wire _3604_;
wire _3605_;
wire _3606_;
wire _3607_;
wire _3608_;
wire _3609_;
wire _3610_;
wire _3611_;
wire _3612_;
wire _3613_;
wire _3614_;
wire _3615_;
wire _3616_;
wire _3617_;
wire _3618_;
wire _3619_;
wire _3620_;
wire _3621_;
wire _3622_;
wire _3623_;
wire _3624_;
wire _3625_;
wire _3626_;
wire _3627_;
wire _3628_;
wire _3629_;
wire _3630_;
wire _3631_;
wire _3632_;
wire _3633_;
wire _3634_;
wire _3635_;
wire _3636_;
wire _3637_;
wire _3638_;
wire _3639_;
wire _3640_;
wire _3641_;
wire _3642_;
wire _3643_;
wire _3644_;
wire _3645_;
wire _3646_;
wire _3647_;
wire _3648_;
wire _3649_;
wire _3650_;
wire _3651_;
wire _3652_;
wire _3653_;
wire _3654_;
wire _3655_;
wire _3656_;
wire _3657_;
wire _3658_;
wire _3659_;
wire _3660_;
wire _3661_;
wire _3662_;
wire _3663_;
wire _3664_;
wire _3665_;
wire _3666_;
wire _3667_;
wire _3668_;
wire _3669_;
wire _3670_;
wire _3671_;
wire _3672_;
wire _3673_;
wire _3674_;
wire _3675_;
wire _3676_;
wire _3677_;
wire _3678_;
wire _3679_;
wire _3680_;
wire _3681_;
wire _3682_;
wire _3683_;
wire _3684_;
wire _3685_;
wire _3686_;
wire _3687_;
wire _3688_;
wire _3689_;
wire _3690_;
wire _3691_;
wire _3692_;
wire _3693_;
wire _3694_;
wire _3695_;
wire _3696_;
wire _3697_;
wire _3698_;
wire _3699_;
wire _3700_;
wire _3701_;
wire _3702_;
wire _3703_;
wire _3704_;
wire _3705_;
wire _3706_;
wire _3707_;
wire _3708_;
wire _3709_;
wire _3710_;
wire _3711_;
wire _3712_;
wire _3713_;
wire _3714_;
wire _3715_;
wire _3716_;
wire _3717_;
wire _3718_;
wire _3719_;
wire _3720_;
wire _3721_;
wire _3722_;
wire _3723_;
wire _3724_;
wire _3725_;
wire _3726_;
wire _3727_;
wire _3728_;
wire _3729_;
wire _3730_;
wire _3731_;
wire _3732_;
wire _3733_;
wire _3734_;
wire _3735_;
wire _3736_;
wire _3737_;
wire _3738_;
wire _3739_;
wire _3740_;
wire _3741_;
wire _3742_;
wire _3743_;
wire _3744_;
wire _3745_;
wire _3746_;
wire _3747_;
wire _3748_;
wire _3749_;
wire _3750_;
wire _3751_;
wire _3752_;
wire _3753_;
wire _3754_;
wire _3755_;
wire _3756_;
wire _3757_;
wire _3758_;
wire _3759_;
wire _3760_;
wire _3761_;
wire _3762_;
wire _3763_;
wire _3764_;
wire _3765_;
wire _3766_;
wire _3767_;
wire _3768_;
wire _3769_;
wire _3770_;
wire _3771_;
wire _3772_;
wire _3773_;
wire _3774_;
wire _3775_;
wire _3776_;
wire _3777_;
wire _3778_;
wire _3779_;
wire _3780_;
wire _3781_;
wire _3782_;
wire _3783_;
wire _3784_;
wire _3785_;
wire _3786_;
wire _3787_;
wire _3788_;
wire _3789_;
wire _3790_;
wire _3791_;
wire _3792_;
wire _3793_;
wire _3794_;
wire _3795_;
wire _3796_;
wire _3797_;
wire _3798_;
wire _3799_;
wire _3800_;
wire _3801_;
wire _3802_;
wire _3803_;
wire _3804_;
wire _3805_;
wire _3806_;
wire _3807_;
wire _3808_;
wire _3809_;
wire _3810_;
wire _3811_;
wire _3812_;
wire _3813_;
wire _3814_;
wire _3815_;
wire _3816_;
wire _3817_;
wire _3818_;
wire _3819_;
wire _3820_;
wire _3821_;
wire _3822_;
wire _3823_;
wire _3824_;
wire _3825_;
wire _3826_;
wire _3827_;
wire _3828_;
wire _3829_;
wire _3830_;
wire _3831_;
wire _3832_;
wire _3833_;
wire _3834_;
wire _3835_;
wire _3836_;
wire _3837_;
wire _3838_;
wire _3839_;
wire _3840_;
wire _3841_;
wire _3842_;
wire _3843_;
wire _3844_;
wire _3845_;
wire _3846_;
wire _3847_;
wire _3848_;
wire _3849_;
wire _3850_;
wire _3851_;
wire _3852_;
wire _3853_;
wire _3854_;
wire _3855_;
wire _3856_;
wire _3857_;
wire _3858_;
wire _3859_;
wire _3860_;
wire _3861_;
wire _3862_;
wire _3863_;
wire _3864_;
wire _3865_;
wire _3866_;
wire _3867_;
wire _3868_;
wire _3869_;
wire _3870_;
wire _3871_;
wire _3872_;
wire _3873_;
wire _3874_;
wire _3875_;
wire _3876_;
wire _3877_;
wire _3878_;
wire _3879_;
wire _3880_;
wire _3881_;
wire _3882_;
wire _3883_;
wire _3884_;
wire _3885_;
wire _3886_;
wire _3887_;
wire _3888_;
wire _3889_;
wire _3890_;
wire _3891_;
wire _3892_;
wire _3893_;
wire _3894_;
wire _3895_;
wire _3896_;
wire _3897_;
wire _3898_;
wire _3899_;
wire _3900_;
wire _3901_;
wire _3902_;
wire _3903_;
wire _3904_;
wire _3905_;
wire _3906_;
wire _3907_;
wire _3908_;
wire _3909_;
wire _3910_;
wire _3911_;
wire _3912_;
wire _3913_;
wire _3914_;
wire _3915_;
wire _3916_;
wire _3917_;
wire _3918_;
wire _3919_;
wire _3920_;
wire _3921_;
wire _3922_;
wire _3923_;
wire _3924_;
wire _3925_;
wire _3926_;
wire _3927_;
wire _3928_;
wire _3929_;
wire _3930_;
wire _3931_;
wire _3932_;
wire _3933_;
wire _3934_;
wire _3935_;
wire _3936_;
wire _3937_;
wire _3938_;
wire _3939_;
wire _3940_;
wire _3941_;
wire _3942_;
wire _3943_;
wire _3944_;
wire _3945_;
wire _3946_;
wire _3947_;
wire _3948_;
wire _3949_;
wire _3950_;
wire _3951_;
wire _3952_;
wire _3953_;
wire _3954_;
wire _3955_;
wire _3956_;
wire _3957_;
wire _3958_;
wire _3959_;
wire _3960_;
wire _3961_;
wire _3962_;
wire _3963_;
wire _3964_;
wire _3965_;
wire _3966_;
wire _3967_;
wire _3968_;
wire _3969_;
wire _3970_;
wire _3971_;
wire _3972_;
wire _3973_;
wire _3974_;
wire _3975_;
wire _3976_;
wire _3977_;
wire _3978_;
wire _3979_;
wire _3980_;
wire _3981_;
wire _3982_;
wire _3983_;
wire _3984_;
wire _3985_;
wire _3986_;
wire _3987_;
wire _3988_;
wire _3989_;
wire _3990_;
wire _3991_;
wire _3992_;
wire _3993_;
wire _3994_;
wire _3995_;
wire _3996_;
wire _3997_;
wire _3998_;
wire _3999_;
wire _4000_;
wire _4001_;
wire _4002_;
wire _4003_;
wire _4004_;
wire _4005_;
wire _4006_;
wire _4007_;
wire _4008_;
wire _4009_;
wire _4010_;
wire _4011_;
wire _4012_;
wire _4013_;
wire _4014_;
wire _4015_;
wire _4016_;
wire _4017_;
wire _4018_;
wire _4019_;
wire _4020_;
wire _4021_;
wire _4022_;
wire _4023_;
wire _4024_;
wire _4025_;
wire _4026_;
wire _4027_;
wire _4028_;
wire _4029_;
wire _4030_;
wire _4031_;
wire _4032_;
wire _4033_;
wire _4034_;
wire _4035_;
wire _4036_;
wire _4037_;
wire _4038_;
wire _4039_;
wire _4040_;
wire _4041_;
wire _4042_;
wire _4043_;
wire _4044_;
wire _4045_;
wire _4046_;
wire _4047_;
wire _4048_;
wire _4049_;
wire _4050_;
wire _4051_;
wire _4052_;
wire _4053_;
wire _4054_;
wire _4055_;
wire _4056_;
wire _4057_;
wire _4058_;
wire _4059_;
wire _4060_;
wire _4061_;
wire _4062_;
wire _4063_;
wire _4064_;
wire _4065_;
wire _4066_;
wire _4067_;
wire _4068_;
wire _4069_;
wire _4070_;
wire _4071_;
wire _4072_;
wire _4073_;
wire _4074_;
wire _4075_;
wire _4076_;
wire _4077_;
wire _4078_;
wire _4079_;
wire _4080_;
wire _4081_;
wire _4082_;
wire _4083_;
wire _4084_;
wire _4085_;
wire _4086_;
wire _4087_;
wire _4088_;
wire _4089_;
wire _4090_;
wire _4091_;
wire _4092_;
wire _4093_;
wire _4094_;
wire _4095_;
wire _4096_;
wire _4097_;
wire _4098_;
wire _4099_;
wire _4100_;
wire _4101_;
wire _4102_;
wire _4103_;
wire _4104_;
wire _4105_;
wire _4106_;
wire _4107_;
wire _4108_;
wire _4109_;
wire _4110_;
wire _4111_;
wire _4112_;
wire _4113_;
wire _4114_;
wire _4115_;
wire _4116_;
wire _4117_;
wire _4118_;
wire _4119_;
wire _4120_;
wire _4121_;
wire _4122_;
wire _4123_;
wire _4124_;
wire _4125_;
wire _4126_;
wire _4127_;
wire _4128_;
wire _4129_;
wire _4130_;
wire _4131_;
wire _4132_;
wire _4133_;
wire _4134_;
wire _4135_;
wire _4136_;
wire _4137_;
wire _4138_;
wire _4139_;
wire _4140_;
wire _4141_;
wire _4142_;
wire _4143_;
wire _4144_;
wire _4145_;
wire _4146_;
wire _4147_;
wire _4148_;
wire _4149_;
wire _4150_;
wire _4151_;
wire _4152_;
wire _4153_;
wire _4154_;
wire _4155_;
wire _4156_;
wire _4157_;
wire _4158_;
wire _4159_;
wire _4160_;
wire _4161_;
wire _4162_;
wire _4163_;
wire _4164_;
wire _4165_;
wire _4166_;
wire _4167_;
wire _4168_;
wire _4169_;
wire _4170_;
wire _4171_;
wire _4172_;
wire _4173_;
wire _4174_;
wire _4175_;
wire _4176_;
wire _4177_;
wire _4178_;
wire _4179_;
wire _4180_;
wire _4181_;
wire _4182_;
wire _4183_;
wire _4184_;
wire _4185_;
wire _4186_;
wire _4187_;
wire _4188_;
wire _4189_;
wire _4190_;
wire _4191_;
wire _4192_;
wire _4193_;
wire _4194_;
wire _4195_;
wire _4196_;
wire _4197_;
wire _4198_;
wire _4199_;
wire _4200_;
wire _4201_;
wire _4202_;
wire _4203_;
wire _4204_;
wire _4205_;
wire _4206_;
wire _4207_;
wire _4208_;
wire _4209_;
wire _4210_;
wire _4211_;
wire _4212_;
wire _4213_;
wire _4214_;
wire _4215_;
wire _4216_;
wire _4217_;
wire _4218_;
wire _4219_;
wire _4220_;
wire _4221_;
wire _4222_;
wire _4223_;
wire _4224_;
wire _4225_;
wire _4226_;
wire _4227_;
wire _4228_;
wire _4229_;
wire _4230_;
wire _4231_;
wire _4232_;
wire _4233_;
wire _4234_;
wire _4235_;
wire _4236_;
wire _4237_;
wire _4238_;
wire _4239_;
wire _4240_;
wire _4241_;
wire _4242_;
wire _4243_;
wire _4244_;
wire _4245_;
wire _4246_;
wire _4247_;
wire _4248_;
wire _4249_;
wire _4250_;
wire _4251_;
wire _4252_;
wire _4253_;
wire _4254_;
wire _4255_;
wire _4256_;
wire _4257_;
wire _4258_;
wire _4259_;
wire _4260_;
wire _4261_;
wire _4262_;
wire _4263_;
wire _4264_;
wire _4265_;
wire _4266_;
wire _4267_;
wire _4268_;
wire _4269_;
wire _4270_;
wire _4271_;
wire _4272_;
wire _4273_;
wire _4274_;
wire _4275_;
wire _4276_;
wire _4277_;
wire _4278_;
wire _4279_;
wire _4280_;
wire _4281_;
wire _4282_;
wire _4283_;
wire _4284_;
wire _4285_;
wire _4286_;
wire _4287_;
wire _4288_;
wire _4289_;
wire _4290_;
wire _4291_;
wire _4292_;
wire _4293_;
wire _4294_;
wire _4295_;
wire _4296_;
wire _4297_;
wire _4298_;
wire _4299_;
wire _4300_;
wire _4301_;
wire _4302_;
wire _4303_;
wire _4304_;
wire _4305_;
wire _4306_;
wire _4307_;
wire _4308_;
wire _4309_;
wire _4310_;
wire _4311_;
wire _4312_;
wire _4313_;
wire _4314_;
wire _4315_;
wire _4316_;
wire _4317_;
wire _4318_;
wire _4319_;
wire _4320_;
wire _4321_;
wire _4322_;
wire _4323_;
wire _4324_;
wire _4325_;
wire _4326_;
wire _4327_;
wire _4328_;
wire _4329_;
wire _4330_;
wire _4331_;
wire _4332_;
wire _4333_;
wire _4334_;
wire _4335_;
wire _4336_;
wire _4337_;
wire _4338_;
wire _4339_;
wire _4340_;
wire _4341_;
wire _4342_;
wire _4343_;
wire _4344_;
wire _4345_;
wire _4346_;
wire _4347_;
wire _4348_;
wire _4349_;
wire _4350_;
wire _4351_;
wire _4352_;
wire _4353_;
wire _4354_;
wire _4355_;
wire _4356_;
wire _4357_;
wire _4358_;
wire _4359_;
wire _4360_;
wire _4361_;
wire _4362_;
wire _4363_;
wire _4364_;
wire _4365_;
wire _4366_;
wire _4367_;
wire _4368_;
wire _4369_;
wire _4370_;
wire _4371_;
wire _4372_;
wire _4373_;
wire _4374_;
wire _4375_;
wire _4376_;
wire _4377_;
wire _4378_;
wire _4379_;
wire _4380_;
wire _4381_;
wire _4382_;
wire _4383_;
wire _4384_;
wire _4385_;
wire _4386_;
wire _4387_;
wire _4388_;
wire _4389_;
wire _4390_;
wire _4391_;
wire _4392_;
wire _4393_;
wire _4394_;
wire _4395_;
wire _4396_;
wire _4397_;
wire _4398_;
wire _4399_;
wire _4400_;
wire _4401_;
wire _4402_;
wire _4403_;
wire _4404_;
wire _4405_;
wire _4406_;
wire _4407_;
wire _4408_;
wire _4409_;
wire _4410_;
wire _4411_;
wire _4412_;
wire _4413_;
wire _4414_;
wire _4415_;
wire _4416_;
wire _4417_;
wire _4418_;
wire _4419_;
wire _4420_;
wire _4421_;
wire _4422_;
wire _4423_;
wire _4424_;
wire _4425_;
wire _4426_;
wire _4427_;
wire _4428_;
wire _4429_;
wire _4430_;
wire _4431_;
wire _4432_;
wire _4433_;
wire _4434_;
wire _4435_;
wire _4436_;
wire _4437_;
wire _4438_;
wire _4439_;
wire _4440_;
wire _4441_;
wire _4442_;
wire _4443_;
wire _4444_;
wire _4445_;
wire _4446_;
wire _4447_;
wire _4448_;
wire _4449_;
wire _4450_;
wire _4451_;
wire _4452_;
wire _4453_;
wire _4454_;
wire _4455_;
wire _4456_;
wire _4457_;
wire _4458_;
wire _4459_;
wire _4460_;
wire _4461_;
wire _4462_;
wire _4463_;
wire _4464_;
wire _4465_;
wire _4466_;
wire _4467_;
wire _4468_;
wire _4469_;
wire _4470_;
wire _4471_;
wire _4472_;
wire _4473_;
wire _4474_;
wire _4475_;
wire _4476_;
wire _4477_;
wire _4478_;
wire _4479_;
wire _4480_;
wire _4481_;
wire _4482_;
wire _4483_;
wire _4484_;
wire _4485_;
wire _4486_;
wire _4487_;
wire _4488_;
wire _4489_;
wire _4490_;
wire _4491_;
wire _4492_;
wire _4493_;
wire _4494_;
wire _4495_;
wire _4496_;
wire _4497_;
wire _4498_;
wire _4499_;
wire _4500_;
wire _4501_;
wire _4502_;
wire _4503_;
wire _4504_;
wire _4505_;
wire _4506_;
wire _4507_;
wire _4508_;
wire _4509_;
wire _4510_;
wire _4511_;
wire _4512_;
wire _4513_;
wire _4514_;
wire _4515_;
wire _4516_;
wire _4517_;
wire _4518_;
wire _4519_;
wire _4520_;
wire _4521_;
wire _4522_;
wire _4523_;
wire _4524_;
wire _4525_;
wire _4526_;
wire _4527_;
wire _4528_;
wire _4529_;
wire _4530_;
wire _4531_;
wire _4532_;
wire _4533_;
wire _4534_;
wire _4535_;
wire _4536_;
wire _4537_;
wire _4538_;
wire _4539_;
wire _4540_;
wire _4541_;
wire _4542_;
wire _4543_;
wire _4544_;
wire _4545_;
wire _4546_;
wire _4547_;
wire _4548_;
wire _4549_;
wire _4550_;
wire _4551_;
wire _4552_;
wire _4553_;
wire _4554_;
wire _4555_;
wire _4556_;
wire _4557_;
wire _4558_;
wire _4559_;
wire _4560_;
wire _4561_;
wire _4562_;
wire _4563_;
wire _4564_;
wire _4565_;
wire _4566_;
wire _4567_;
wire _4568_;
wire _4569_;
wire _4570_;
wire _4571_;
wire _4572_;
wire _4573_;
wire _4574_;
wire _4575_;
wire _4576_;
wire _4577_;
wire _4578_;
wire _4579_;
wire _4580_;
wire _4581_;
wire _4582_;
wire _4583_;
wire _4584_;
wire _4585_;
wire _4586_;
wire _4587_;
wire _4588_;
wire _4589_;
wire _4590_;
wire _4591_;
wire _4592_;
wire _4593_;
wire _4594_;
wire _4595_;
wire _4596_;
wire _4597_;
wire _4598_;
wire _4599_;
wire _4600_;
wire _4601_;
wire _4602_;
wire _4603_;
wire _4604_;
wire _4605_;
wire _4606_;
wire _4607_;
wire _4608_;
wire _4609_;
wire _4610_;
wire _4611_;
wire _4612_;
wire _4613_;
wire _4614_;
wire _4615_;
wire _4616_;
wire _4617_;
wire _4618_;
wire _4619_;
wire _4620_;
wire _4621_;
wire _4622_;
wire _4623_;
wire _4624_;
wire _4625_;
wire _4626_;
wire _4627_;
wire _4628_;
wire _4629_;
wire _4630_;
wire _4631_;
wire _4632_;
wire _4633_;
wire _4634_;
wire _4635_;
wire _4636_;
wire _4637_;
wire _4638_;
wire _4639_;
wire _4640_;
wire _4641_;
wire _4642_;
wire _4643_;
wire _4644_;
wire _4645_;
wire _4646_;
wire _4647_;
wire _4648_;
wire _4649_;
wire _4650_;
wire _4651_;
wire _4652_;
wire _4653_;
wire _4654_;
wire _4655_;
wire _4656_;
wire _4657_;
wire _4658_;
wire _4659_;
wire _4660_;
wire _4661_;
wire _4662_;
wire _4663_;
wire _4664_;
wire _4665_;
wire _4666_;
wire _4667_;
wire _4668_;
wire _4669_;
wire _4670_;
wire _4671_;
wire _4672_;
wire _4673_;
wire _4674_;
wire _4675_;
wire _4676_;
wire _4677_;
wire _4678_;
wire _4679_;
wire _4680_;
wire _4681_;
wire _4682_;
wire _4683_;
wire _4684_;
wire _4685_;
wire _4686_;
wire _4687_;
wire _4688_;
wire _4689_;
wire _4690_;
wire _4691_;
wire _4692_;
wire _4693_;
wire _4694_;
wire _4695_;
wire _4696_;
wire _4697_;
wire _4698_;
wire _4699_;
wire _4700_;
wire _4701_;
wire _4702_;
wire _4703_;
wire _4704_;
wire _4705_;
wire _4706_;
wire _4707_;
wire _4708_;
wire _4709_;
wire _4710_;
wire _4711_;
wire _4712_;
wire _4713_;
wire _4714_;
wire _4715_;
wire _4716_;
wire _4717_;
wire _4718_;
wire _4719_;
wire _4720_;
wire _4721_;
wire _4722_;
wire _4723_;
wire _4724_;
wire _4725_;
wire _4726_;
wire _4727_;
wire _4728_;
wire _4729_;
wire _4730_;
wire _4731_;
wire _4732_;
wire _4733_;
wire _4734_;
wire _4735_;
wire _4736_;
wire _4737_;
wire _4738_;
wire _4739_;
wire _4740_;
wire _4741_;
wire _4742_;
wire _4743_;
wire _4744_;
wire _4745_;
wire _4746_;
wire _4747_;
wire _4748_;
wire _4749_;
wire _4750_;
wire _4751_;
wire _4752_;
wire _4753_;
wire _4754_;
wire _4755_;
wire _4756_;
wire _4757_;
wire _4758_;
wire _4759_;
wire _4760_;
wire _4761_;
wire _4762_;
wire _4763_;
wire _4764_;
wire _4765_;
wire _4766_;
wire _4767_;
wire _4768_;
wire _4769_;
wire _4770_;
wire _4771_;
wire _4772_;
wire _4773_;
wire _4774_;
wire _4775_;
wire _4776_;
wire _4777_;
wire _4778_;
wire _4779_;
wire _4780_;
wire _4781_;
wire _4782_;
wire _4783_;
wire _4784_;
wire _4785_;
wire _4786_;
wire _4787_;
wire _4788_;
wire _4789_;
wire _4790_;
wire _4791_;
wire _4792_;
wire _4793_;
wire _4794_;
wire _4795_;
wire _4796_;
wire _4797_;
wire _4798_;
wire _4799_;
wire _4800_;
wire _4801_;
wire _4802_;
wire _4803_;
wire _4804_;
wire _4805_;
wire _4806_;
wire _4807_;
wire _4808_;
wire _4809_;
wire _4810_;
wire _4811_;
wire _4812_;
wire _4813_;
wire _4814_;
wire _4815_;
wire _4816_;
wire _4817_;
wire _4818_;
wire _4819_;
wire _4820_;
wire _4821_;
wire _4822_;
wire _4823_;
wire _4824_;
wire _4825_;
wire _4826_;
wire _4827_;
wire _4828_;
wire _4829_;
wire _4830_;
wire _4831_;
wire _4832_;
wire _4833_;
wire _4834_;
wire _4835_;
wire _4836_;
wire _4837_;
wire _4838_;
wire _4839_;
wire _4840_;
wire _4841_;
wire _4842_;
wire _4843_;
wire _4844_;
wire _4845_;
wire _4846_;
wire _4847_;
wire _4848_;
wire _4849_;
wire _4850_;
wire _4851_;
wire _4852_;
wire _4853_;
wire _4854_;
wire _4855_;
wire _4856_;
wire _4857_;
wire _4858_;
wire _4859_;
wire _4860_;
wire _4861_;
wire _4862_;
wire _4863_;
wire _4864_;
wire _4865_;
wire _4866_;
wire _4867_;
wire _4868_;
wire _4869_;
wire _4870_;
wire _4871_;
wire _4872_;
wire _4873_;
wire _4874_;
wire _4875_;
wire _4876_;
wire _4877_;
wire _4878_;
wire _4879_;
wire _4880_;
wire _4881_;
wire _4882_;
wire _4883_;
wire _4884_;
wire _4885_;
wire _4886_;
wire _4887_;
wire _4888_;
wire _4889_;
wire _4890_;
wire _4891_;
wire _4892_;
wire _4893_;
wire _4894_;
wire _4895_;
wire _4896_;
wire _4897_;
wire _4898_;
wire _4899_;
wire _4900_;
wire _4901_;
wire _4902_;
wire _4903_;
wire _4904_;
wire _4905_;
wire _4906_;
wire _4907_;
wire _4908_;
wire _4909_;
wire _4910_;
wire _4911_;
wire _4912_;
wire _4913_;
wire _4914_;
wire _4915_;
wire _4916_;
wire _4917_;
wire _4918_;
wire _4919_;
wire _4920_;
wire _4921_;
wire _4922_;
wire _4923_;
wire _4924_;
wire _4925_;
wire _4926_;
wire _4927_;
wire _4928_;
wire _4929_;
wire _4930_;
wire _4931_;
wire _4932_;
wire _4933_;
wire _4934_;
wire _4935_;
wire _4936_;
wire _4937_;
wire _4938_;
wire _4939_;
wire _4940_;
wire _4941_;
wire _4942_;
wire _4943_;
wire _4944_;
wire _4945_;
wire _4946_;
wire _4947_;
wire _4948_;
wire _4949_;
wire _4950_;
wire _4951_;
wire _4952_;
wire _4953_;
wire _4954_;
wire _4955_;
wire _4956_;
wire _4957_;
wire _4958_;
wire _4959_;
wire _4960_;
wire _4961_;
wire _4962_;
wire _4963_;
wire _4964_;
wire _4965_;
wire _4966_;
wire _4967_;
wire _4968_;
wire _4969_;
wire _4970_;
wire _4971_;
wire _4972_;
wire _4973_;
wire _4974_;
wire _4975_;
wire _4976_;
wire _4977_;
wire _4978_;
wire _4979_;
wire _4980_;
wire _4981_;
wire _4982_;
wire _4983_;
wire _4984_;
wire _4985_;
wire _4986_;
wire _4987_;
wire _4988_;
wire _4989_;
wire _4990_;
wire _4991_;
wire _4992_;
wire _4993_;
wire _4994_;
wire _4995_;
wire _4996_;
wire _4997_;
wire _4998_;
wire _4999_;
wire _5000_;
wire _5001_;
wire _5002_;
wire _5003_;
wire _5004_;
wire _5005_;
wire _5006_;
wire _5007_;
wire _5008_;
wire _5009_;
wire _5010_;
wire _5011_;
wire _5012_;
wire _5013_;
wire _5014_;
wire _5015_;
wire _5016_;
wire _5017_;
wire _5018_;
wire _5019_;
wire _5020_;
wire _5021_;
wire _5022_;
wire _5023_;
wire _5024_;
wire _5025_;
wire _5026_;
wire _5027_;
wire _5028_;
wire _5029_;
wire _5030_;
wire _5031_;
wire _5032_;
wire _5033_;
wire _5034_;
wire _5035_;
wire _5036_;
wire _5037_;
wire _5038_;
wire _5039_;
wire _5040_;
wire _5041_;
wire _5042_;
wire _5043_;
wire _5044_;
wire _5045_;
wire _5046_;
wire _5047_;
wire _5048_;
wire _5049_;
wire _5050_;
wire _5051_;
wire _5052_;
wire _5053_;
wire _5054_;
wire _5055_;
wire _5056_;
wire _5057_;
wire _5058_;
wire _5059_;
wire _5060_;
wire _5061_;
wire _5062_;
wire _5063_;
wire _5064_;
wire _5065_;
wire _5066_;
wire _5067_;
wire _5068_;
wire _5069_;
wire _5070_;
wire _5071_;
wire _5072_;
wire _5073_;
wire _5074_;
wire _5075_;
wire _5076_;
wire _5077_;
wire _5078_;
wire _5079_;
wire _5080_;
wire _5081_;
wire _5082_;
wire _5083_;
wire _5084_;
wire _5085_;
wire _5086_;
wire _5087_;
wire _5088_;
wire _5089_;
wire _5090_;
wire _5091_;
wire _5092_;
wire _5093_;
wire _5094_;
wire _5095_;
wire _5096_;
wire _5097_;
wire _5098_;
wire _5099_;
wire _5100_;
wire _5101_;
wire _5102_;
wire _5103_;
wire _5104_;
wire _5105_;
wire _5106_;
wire _5107_;
wire _5108_;
wire _5109_;
wire _5110_;
wire _5111_;
wire _5112_;
wire _5113_;
wire _5114_;
wire _5115_;
wire _5116_;
wire _5117_;
wire _5118_;
wire _5119_;
wire _5120_;
wire _5121_;
wire _5122_;
wire _5123_;
wire _5124_;
wire _5125_;
wire _5126_;
wire _5127_;
wire _5128_;
wire _5129_;
wire _5130_;
wire _5131_;
wire _5132_;
wire _5133_;
wire _5134_;
wire _5135_;
wire _5136_;
wire _5137_;
wire _5138_;
wire _5139_;
wire _5140_;
wire _5141_;
wire _5142_;
wire _5143_;
wire _5144_;
wire _5145_;
wire _5146_;
wire _5147_;
wire _5148_;
wire _5149_;
wire _5150_;
wire _5151_;
wire _5152_;
wire _5153_;
wire _5154_;
wire _5155_;
wire _5156_;
wire _5157_;
wire _5158_;
wire _5159_;
wire _5160_;
wire _5161_;
wire _5162_;
wire _5163_;
wire _5164_;
wire _5165_;
wire _5166_;
wire _5167_;
wire _5168_;
wire _5169_;
wire _5170_;
wire _5171_;
wire _5172_;
wire _5173_;
wire _5174_;
wire _5175_;
wire _5176_;
wire _5177_;
wire _5178_;
wire _5179_;
wire _5180_;
wire _5181_;
wire _5182_;
wire _5183_;
wire _5184_;
wire _5185_;
wire _5186_;
wire _5187_;
wire _5188_;
wire _5189_;
wire _5190_;
wire _5191_;
wire _5192_;
wire _5193_;
wire _5194_;
wire _5195_;
wire _5196_;
wire _5197_;
wire _5198_;
wire _5199_;
wire _5200_;
wire _5201_;
wire _5202_;
wire _5203_;
wire _5204_;
wire _5205_;
wire _5206_;
wire _5207_;
wire _5208_;
wire _5209_;
wire _5210_;
wire _5211_;
wire _5212_;
wire _5213_;
wire _5214_;
wire _5215_;
wire _5216_;
wire _5217_;
wire _5218_;
wire _5219_;
wire _5220_;
wire _5221_;
wire _5222_;
wire _5223_;
wire _5224_;
wire _5225_;
wire _5226_;
wire _5227_;
wire _5228_;
wire _5229_;
wire _5230_;
wire _5231_;
wire _5232_;
wire _5233_;
wire _5234_;
wire _5235_;
wire _5236_;
wire _5237_;
wire _5238_;
wire _5239_;
wire _5240_;
wire _5241_;
wire _5242_;
wire _5243_;
wire _5244_;
wire _5245_;
wire _5246_;
wire _5247_;
wire _5248_;
wire _5249_;
wire _5250_;
wire _5251_;
wire _5252_;
wire _5253_;
wire _5254_;
wire _5255_;
wire _5256_;
wire _5257_;
wire _5258_;
wire _5259_;
wire _5260_;
wire _5261_;
wire _5262_;
wire _5263_;
wire _5264_;
wire _5265_;
wire _5266_;
wire _5267_;
wire _5268_;
wire _5269_;
wire _5270_;
wire _5271_;
wire _5272_;
wire _5273_;
wire _5274_;
wire _5275_;
wire _5276_;
wire _5277_;
wire _5278_;
wire _5279_;
wire _5280_;
wire _5281_;
wire _5282_;
wire _5283_;
wire _5284_;
wire _5285_;
wire _5286_;
wire _5287_;
wire _5288_;
wire _5289_;
wire _5290_;
wire _5291_;
wire _5292_;
wire _5293_;
wire _5294_;
wire _5295_;
wire _5296_;
wire _5297_;
wire _5298_;
wire _5299_;
wire _5300_;
wire _5301_;
wire _5302_;
wire _5303_;
wire _5304_;
wire _5305_;
wire _5306_;
wire _5307_;
wire _5308_;
wire _5309_;
wire _5310_;
wire _5311_;
wire _5312_;
wire _5313_;
wire _5314_;
wire _5315_;
wire _5316_;
wire _5317_;
wire _5318_;
wire _5319_;
wire _5320_;
wire _5321_;
wire _5322_;
wire _5323_;
wire _5324_;
wire _5325_;
wire _5326_;
wire _5327_;
wire _5328_;
wire _5329_;
wire _5330_;
wire _5331_;
wire _5332_;
wire _5333_;
wire _5334_;
wire _5335_;
wire _5336_;
wire _5337_;
wire _5338_;
wire _5339_;
wire _5340_;
wire _5341_;
wire _5342_;
wire _5343_;
wire _5344_;
wire _5345_;
wire _5346_;
wire _5347_;
wire _5348_;
wire _5349_;
wire _5350_;
wire _5351_;
wire _5352_;
wire _5353_;
wire _5354_;
wire _5355_;
wire _5356_;
wire _5357_;
wire _5358_;
wire _5359_;
wire _5360_;
wire _5361_;
wire _5362_;
wire _5363_;
wire _5364_;
wire _5365_;
wire _5366_;
wire _5367_;
wire _5368_;
wire _5369_;
wire _5370_;
wire _5371_;
wire _5372_;
wire _5373_;
wire _5374_;
wire _5375_;
wire _5376_;
wire _5377_;
wire _5378_;
wire _5379_;
wire _5380_;
wire _5381_;
wire _5382_;
wire _5383_;
wire _5384_;
wire _5385_;
wire _5386_;
wire _5387_;
wire _5388_;
wire _5389_;
wire _5390_;
wire _5391_;
wire _5392_;
wire _5393_;
wire _5394_;
wire _5395_;
wire _5396_;
wire _5397_;
wire _5398_;
wire _5399_;
wire _5400_;
wire _5401_;
wire _5402_;
wire _5403_;
wire _5404_;
wire _5405_;
wire _5406_;
wire _5407_;
wire _5408_;
wire _5409_;
wire _5410_;
wire _5411_;
wire _5412_;
wire _5413_;
wire _5414_;
wire _5415_;
wire _5416_;
wire _5417_;
wire _5418_;
wire _5419_;
wire _5420_;
wire _5421_;
wire _5422_;
wire _5423_;
wire _5424_;
wire _5425_;
wire _5426_;
wire _5427_;
wire _5428_;
wire _5429_;
wire _5430_;
wire _5431_;
wire _5432_;
wire _5433_;
wire _5434_;
wire _5435_;
wire _5436_;
wire _5437_;
wire _5438_;
wire _5439_;
wire _5440_;
wire _5441_;
wire _5442_;
wire _5443_;
wire _5444_;
wire _5445_;
wire _5446_;
wire _5447_;
wire _5448_;
wire _5449_;
wire _5450_;
wire _5451_;
wire _5452_;
wire _5453_;
wire _5454_;
wire _5455_;
wire _5456_;
wire _5457_;
wire zeroWire;
wire oneWire;
assign zeroWire = 1'b0 /*6482*/;
assign oneWire = 1'b1 /*6482*/;
assign _21_ = ~D[0] /*6384*/;
assign _18_ = R_0[15] & _21_ /*6380*/;
assign _19_ = R_0[15] ^ _21_ /*6383*/;
assign _20_ = oneWire & _19_ /*6381*/;
assign _0_ = oneWire ^ _19_ /*6382*/;
assign _17_ = _18_ | _20_ /*6379*/;
assign _26_ = ~D[1] /*6378*/;
assign _23_ = R_0[16] & _26_ /*6374*/;
assign _24_ = R_0[16] ^ _26_ /*6377*/;
assign _25_ = _17_ & _24_ /*6375*/;
assign _1_ = _17_ ^ _24_ /*6376*/;
assign _22_ = _23_ | _25_ /*6373*/;
assign _31_ = ~D[2] /*6372*/;
assign _28_ = R_0[17] & _31_ /*6368*/;
assign _29_ = R_0[17] ^ _31_ /*6371*/;
assign _30_ = _22_ & _29_ /*6369*/;
assign _2_ = _22_ ^ _29_ /*6370*/;
assign _27_ = _28_ | _30_ /*6367*/;
assign _36_ = ~D[3] /*6366*/;
assign _33_ = R_0[18] & _36_ /*6362*/;
assign _34_ = R_0[18] ^ _36_ /*6365*/;
assign _35_ = _27_ & _34_ /*6363*/;
assign _3_ = _27_ ^ _34_ /*6364*/;
assign _32_ = _33_ | _35_ /*6361*/;
assign _41_ = ~D[4] /*6360*/;
assign _38_ = R_0[19] & _41_ /*6356*/;
assign _39_ = R_0[19] ^ _41_ /*6359*/;
assign _40_ = _32_ & _39_ /*6357*/;
assign _4_ = _32_ ^ _39_ /*6358*/;
assign _37_ = _38_ | _40_ /*6355*/;
assign _46_ = ~D[5] /*6354*/;
assign _43_ = R_0[20] & _46_ /*6350*/;
assign _44_ = R_0[20] ^ _46_ /*6353*/;
assign _45_ = _37_ & _44_ /*6351*/;
assign _5_ = _37_ ^ _44_ /*6352*/;
assign _42_ = _43_ | _45_ /*6349*/;
assign _51_ = ~D[6] /*6348*/;
assign _48_ = R_0[21] & _51_ /*6344*/;
assign _49_ = R_0[21] ^ _51_ /*6347*/;
assign _50_ = _42_ & _49_ /*6345*/;
assign _6_ = _42_ ^ _49_ /*6346*/;
assign _47_ = _48_ | _50_ /*6343*/;
assign _56_ = ~D[7] /*6342*/;
assign _53_ = R_0[22] & _56_ /*6338*/;
assign _54_ = R_0[22] ^ _56_ /*6341*/;
assign _55_ = _47_ & _54_ /*6339*/;
assign _7_ = _47_ ^ _54_ /*6340*/;
assign _52_ = _53_ | _55_ /*6337*/;
assign _61_ = ~D[8] /*6336*/;
assign _58_ = R_0[23] & _61_ /*6332*/;
assign _59_ = R_0[23] ^ _61_ /*6335*/;
assign _60_ = _52_ & _59_ /*6333*/;
assign _8_ = _52_ ^ _59_ /*6334*/;
assign _57_ = _58_ | _60_ /*6331*/;
assign _66_ = ~D[9] /*6330*/;
assign _63_ = R_0[24] & _66_ /*6326*/;
assign _64_ = R_0[24] ^ _66_ /*6329*/;
assign _65_ = _57_ & _64_ /*6327*/;
assign _9_ = _57_ ^ _64_ /*6328*/;
assign _62_ = _63_ | _65_ /*6325*/;
assign _71_ = ~D[10] /*6324*/;
assign _68_ = R_0[25] & _71_ /*6320*/;
assign _69_ = R_0[25] ^ _71_ /*6323*/;
assign _70_ = _62_ & _69_ /*6321*/;
assign _10_ = _62_ ^ _69_ /*6322*/;
assign _67_ = _68_ | _70_ /*6319*/;
assign _76_ = ~D[11] /*6318*/;
assign _73_ = R_0[26] & _76_ /*6314*/;
assign _74_ = R_0[26] ^ _76_ /*6317*/;
assign _75_ = _67_ & _74_ /*6315*/;
assign _11_ = _67_ ^ _74_ /*6316*/;
assign _72_ = _73_ | _75_ /*6313*/;
assign _81_ = ~D[12] /*6312*/;
assign _78_ = R_0[27] & _81_ /*6308*/;
assign _79_ = R_0[27] ^ _81_ /*6311*/;
assign _80_ = _72_ & _79_ /*6309*/;
assign _12_ = _72_ ^ _79_ /*6310*/;
assign _77_ = _78_ | _80_ /*6307*/;
assign _86_ = ~D[13] /*6306*/;
assign _83_ = R_0[28] & _86_ /*6302*/;
assign _84_ = R_0[28] ^ _86_ /*6305*/;
assign _85_ = _77_ & _84_ /*6303*/;
assign _13_ = _77_ ^ _84_ /*6304*/;
assign _82_ = _83_ | _85_ /*6301*/;
assign _91_ = ~D[14] /*6300*/;
assign _88_ = R_0[29] & _91_ /*6296*/;
assign _89_ = R_0[29] ^ _91_ /*6299*/;
assign _90_ = _82_ & _89_ /*6297*/;
assign _14_ = _82_ ^ _89_ /*6298*/;
assign _87_ = _88_ | _90_ /*6295*/;
assign _92_ = zeroWire & oneWire /*6290*/;
assign _93_ = zeroWire ^ oneWire /*6293*/;
assign _94_ = _87_ & _93_ /*6291*/;
assign _15_ = _87_ ^ _93_ /*6292*/;
assign Q[15] = _92_ | _94_ /*6289*/;
assign _115_ = ~Q[15] /*6193*/;
assign _114_ = _115_ & D[0] /*6192*/;
assign _117_ = _0_ & _114_ /*6187*/;
assign _118_ = _0_ ^ _114_ /*6190*/;
assign _119_ = zeroWire & _118_ /*6188*/;
assign _97_ = zeroWire ^ _118_ /*6189*/;
assign _116_ = _117_ | _119_ /*6186*/;
assign _121_ = ~Q[15] /*6185*/;
assign _120_ = _121_ & D[1] /*6184*/;
assign _123_ = _1_ & _120_ /*6179*/;
assign _124_ = _1_ ^ _120_ /*6182*/;
assign _125_ = _116_ & _124_ /*6180*/;
assign _98_ = _116_ ^ _124_ /*6181*/;
assign _122_ = _123_ | _125_ /*6178*/;
assign _127_ = ~Q[15] /*6177*/;
assign _126_ = _127_ & D[2] /*6176*/;
assign _129_ = _2_ & _126_ /*6171*/;
assign _130_ = _2_ ^ _126_ /*6174*/;
assign _131_ = _122_ & _130_ /*6172*/;
assign _99_ = _122_ ^ _130_ /*6173*/;
assign _128_ = _129_ | _131_ /*6170*/;
assign _133_ = ~Q[15] /*6169*/;
assign _132_ = _133_ & D[3] /*6168*/;
assign _135_ = _3_ & _132_ /*6163*/;
assign _136_ = _3_ ^ _132_ /*6166*/;
assign _137_ = _128_ & _136_ /*6164*/;
assign _100_ = _128_ ^ _136_ /*6165*/;
assign _134_ = _135_ | _137_ /*6162*/;
assign _139_ = ~Q[15] /*6161*/;
assign _138_ = _139_ & D[4] /*6160*/;
assign _141_ = _4_ & _138_ /*6155*/;
assign _142_ = _4_ ^ _138_ /*6158*/;
assign _143_ = _134_ & _142_ /*6156*/;
assign _101_ = _134_ ^ _142_ /*6157*/;
assign _140_ = _141_ | _143_ /*6154*/;
assign _145_ = ~Q[15] /*6153*/;
assign _144_ = _145_ & D[5] /*6152*/;
assign _147_ = _5_ & _144_ /*6147*/;
assign _148_ = _5_ ^ _144_ /*6150*/;
assign _149_ = _140_ & _148_ /*6148*/;
assign _102_ = _140_ ^ _148_ /*6149*/;
assign _146_ = _147_ | _149_ /*6146*/;
assign _151_ = ~Q[15] /*6145*/;
assign _150_ = _151_ & D[6] /*6144*/;
assign _153_ = _6_ & _150_ /*6139*/;
assign _154_ = _6_ ^ _150_ /*6142*/;
assign _155_ = _146_ & _154_ /*6140*/;
assign _103_ = _146_ ^ _154_ /*6141*/;
assign _152_ = _153_ | _155_ /*6138*/;
assign _157_ = ~Q[15] /*6137*/;
assign _156_ = _157_ & D[7] /*6136*/;
assign _159_ = _7_ & _156_ /*6131*/;
assign _160_ = _7_ ^ _156_ /*6134*/;
assign _161_ = _152_ & _160_ /*6132*/;
assign _104_ = _152_ ^ _160_ /*6133*/;
assign _158_ = _159_ | _161_ /*6130*/;
assign _163_ = ~Q[15] /*6129*/;
assign _162_ = _163_ & D[8] /*6128*/;
assign _165_ = _8_ & _162_ /*6123*/;
assign _166_ = _8_ ^ _162_ /*6126*/;
assign _167_ = _158_ & _166_ /*6124*/;
assign _105_ = _158_ ^ _166_ /*6125*/;
assign _164_ = _165_ | _167_ /*6122*/;
assign _169_ = ~Q[15] /*6121*/;
assign _168_ = _169_ & D[9] /*6120*/;
assign _171_ = _9_ & _168_ /*6115*/;
assign _172_ = _9_ ^ _168_ /*6118*/;
assign _173_ = _164_ & _172_ /*6116*/;
assign _106_ = _164_ ^ _172_ /*6117*/;
assign _170_ = _171_ | _173_ /*6114*/;
assign _175_ = ~Q[15] /*6113*/;
assign _174_ = _175_ & D[10] /*6112*/;
assign _177_ = _10_ & _174_ /*6107*/;
assign _178_ = _10_ ^ _174_ /*6110*/;
assign _179_ = _170_ & _178_ /*6108*/;
assign _107_ = _170_ ^ _178_ /*6109*/;
assign _176_ = _177_ | _179_ /*6106*/;
assign _181_ = ~Q[15] /*6105*/;
assign _180_ = _181_ & D[11] /*6104*/;
assign _183_ = _11_ & _180_ /*6099*/;
assign _184_ = _11_ ^ _180_ /*6102*/;
assign _185_ = _176_ & _184_ /*6100*/;
assign _108_ = _176_ ^ _184_ /*6101*/;
assign _182_ = _183_ | _185_ /*6098*/;
assign _187_ = ~Q[15] /*6097*/;
assign _186_ = _187_ & D[12] /*6096*/;
assign _189_ = _12_ & _186_ /*6091*/;
assign _190_ = _12_ ^ _186_ /*6094*/;
assign _191_ = _182_ & _190_ /*6092*/;
assign _109_ = _182_ ^ _190_ /*6093*/;
assign _188_ = _189_ | _191_ /*6090*/;
assign _193_ = ~Q[15] /*6089*/;
assign _192_ = _193_ & D[13] /*6088*/;
assign _195_ = _13_ & _192_ /*6083*/;
assign _196_ = _13_ ^ _192_ /*6086*/;
assign _197_ = _188_ & _196_ /*6084*/;
assign _110_ = _188_ ^ _196_ /*6085*/;
assign _194_ = _195_ | _197_ /*6082*/;
assign _199_ = ~Q[15] /*6081*/;
assign _198_ = _199_ & D[14] /*6080*/;
assign _201_ = _14_ & _198_ /*6075*/;
assign _202_ = _14_ ^ _198_ /*6078*/;
assign _203_ = _194_ & _202_ /*6076*/;
assign _111_ = _194_ ^ _202_ /*6077*/;
assign _200_ = _201_ | _203_ /*6074*/;
assign _205_ = ~Q[15] /*6073*/;
assign _204_ = _205_ & zeroWire /*6072*/;
assign _206_ = _15_ ^ _204_ /*6070*/;
assign _112_ = _206_ ^ _200_ /*6069*/;
assign _229_ = ~D[0] /*6007*/;
assign _226_ = R_0[14] & _229_ /*6003*/;
assign _227_ = R_0[14] ^ _229_ /*6006*/;
assign _228_ = oneWire & _227_ /*6004*/;
assign _209_ = oneWire ^ _227_ /*6005*/;
assign _225_ = _226_ | _228_ /*6002*/;
assign _234_ = ~D[1] /*6001*/;
assign _231_ = _97_ & _234_ /*5997*/;
assign _232_ = _97_ ^ _234_ /*6000*/;
assign _233_ = _225_ & _232_ /*5998*/;
assign _210_ = _225_ ^ _232_ /*5999*/;
assign _230_ = _231_ | _233_ /*5996*/;
assign _239_ = ~D[2] /*5995*/;
assign _236_ = _98_ & _239_ /*5991*/;
assign _237_ = _98_ ^ _239_ /*5994*/;
assign _238_ = _230_ & _237_ /*5992*/;
assign _211_ = _230_ ^ _237_ /*5993*/;
assign _235_ = _236_ | _238_ /*5990*/;
assign _244_ = ~D[3] /*5989*/;
assign _241_ = _99_ & _244_ /*5985*/;
assign _242_ = _99_ ^ _244_ /*5988*/;
assign _243_ = _235_ & _242_ /*5986*/;
assign _212_ = _235_ ^ _242_ /*5987*/;
assign _240_ = _241_ | _243_ /*5984*/;
assign _249_ = ~D[4] /*5983*/;
assign _246_ = _100_ & _249_ /*5979*/;
assign _247_ = _100_ ^ _249_ /*5982*/;
assign _248_ = _240_ & _247_ /*5980*/;
assign _213_ = _240_ ^ _247_ /*5981*/;
assign _245_ = _246_ | _248_ /*5978*/;
assign _254_ = ~D[5] /*5977*/;
assign _251_ = _101_ & _254_ /*5973*/;
assign _252_ = _101_ ^ _254_ /*5976*/;
assign _253_ = _245_ & _252_ /*5974*/;
assign _214_ = _245_ ^ _252_ /*5975*/;
assign _250_ = _251_ | _253_ /*5972*/;
assign _259_ = ~D[6] /*5971*/;
assign _256_ = _102_ & _259_ /*5967*/;
assign _257_ = _102_ ^ _259_ /*5970*/;
assign _258_ = _250_ & _257_ /*5968*/;
assign _215_ = _250_ ^ _257_ /*5969*/;
assign _255_ = _256_ | _258_ /*5966*/;
assign _264_ = ~D[7] /*5965*/;
assign _261_ = _103_ & _264_ /*5961*/;
assign _262_ = _103_ ^ _264_ /*5964*/;
assign _263_ = _255_ & _262_ /*5962*/;
assign _216_ = _255_ ^ _262_ /*5963*/;
assign _260_ = _261_ | _263_ /*5960*/;
assign _269_ = ~D[8] /*5959*/;
assign _266_ = _104_ & _269_ /*5955*/;
assign _267_ = _104_ ^ _269_ /*5958*/;
assign _268_ = _260_ & _267_ /*5956*/;
assign _217_ = _260_ ^ _267_ /*5957*/;
assign _265_ = _266_ | _268_ /*5954*/;
assign _274_ = ~D[9] /*5953*/;
assign _271_ = _105_ & _274_ /*5949*/;
assign _272_ = _105_ ^ _274_ /*5952*/;
assign _273_ = _265_ & _272_ /*5950*/;
assign _218_ = _265_ ^ _272_ /*5951*/;
assign _270_ = _271_ | _273_ /*5948*/;
assign _279_ = ~D[10] /*5947*/;
assign _276_ = _106_ & _279_ /*5943*/;
assign _277_ = _106_ ^ _279_ /*5946*/;
assign _278_ = _270_ & _277_ /*5944*/;
assign _219_ = _270_ ^ _277_ /*5945*/;
assign _275_ = _276_ | _278_ /*5942*/;
assign _284_ = ~D[11] /*5941*/;
assign _281_ = _107_ & _284_ /*5937*/;
assign _282_ = _107_ ^ _284_ /*5940*/;
assign _283_ = _275_ & _282_ /*5938*/;
assign _220_ = _275_ ^ _282_ /*5939*/;
assign _280_ = _281_ | _283_ /*5936*/;
assign _289_ = ~D[12] /*5935*/;
assign _286_ = _108_ & _289_ /*5931*/;
assign _287_ = _108_ ^ _289_ /*5934*/;
assign _288_ = _280_ & _287_ /*5932*/;
assign _221_ = _280_ ^ _287_ /*5933*/;
assign _285_ = _286_ | _288_ /*5930*/;
assign _294_ = ~D[13] /*5929*/;
assign _291_ = _109_ & _294_ /*5925*/;
assign _292_ = _109_ ^ _294_ /*5928*/;
assign _293_ = _285_ & _292_ /*5926*/;
assign _222_ = _285_ ^ _292_ /*5927*/;
assign _290_ = _291_ | _293_ /*5924*/;
assign _299_ = ~D[14] /*5923*/;
assign _296_ = _110_ & _299_ /*5919*/;
assign _297_ = _110_ ^ _299_ /*5922*/;
assign _298_ = _290_ & _297_ /*5920*/;
assign _223_ = _290_ ^ _297_ /*5921*/;
assign _295_ = _296_ | _298_ /*5918*/;
assign _300_ = _111_ & oneWire /*5913*/;
assign _301_ = _111_ ^ oneWire /*5916*/;
assign _302_ = _295_ & _301_ /*5914*/;
assign _224_ = _295_ ^ _301_ /*5915*/;
assign Q[14] = _300_ | _302_ /*5912*/;
assign _339_ = ~Q[14] /*5815*/;
assign _338_ = _339_ & D[0] /*5814*/;
assign _341_ = _209_ & _338_ /*5809*/;
assign _342_ = _209_ ^ _338_ /*5812*/;
assign _343_ = zeroWire & _342_ /*5810*/;
assign _321_ = zeroWire ^ _342_ /*5811*/;
assign _340_ = _341_ | _343_ /*5808*/;
assign _345_ = ~Q[14] /*5807*/;
assign _344_ = _345_ & D[1] /*5806*/;
assign _347_ = _210_ & _344_ /*5801*/;
assign _348_ = _210_ ^ _344_ /*5804*/;
assign _349_ = _340_ & _348_ /*5802*/;
assign _322_ = _340_ ^ _348_ /*5803*/;
assign _346_ = _347_ | _349_ /*5800*/;
assign _351_ = ~Q[14] /*5799*/;
assign _350_ = _351_ & D[2] /*5798*/;
assign _353_ = _211_ & _350_ /*5793*/;
assign _354_ = _211_ ^ _350_ /*5796*/;
assign _355_ = _346_ & _354_ /*5794*/;
assign _323_ = _346_ ^ _354_ /*5795*/;
assign _352_ = _353_ | _355_ /*5792*/;
assign _357_ = ~Q[14] /*5791*/;
assign _356_ = _357_ & D[3] /*5790*/;
assign _359_ = _212_ & _356_ /*5785*/;
assign _360_ = _212_ ^ _356_ /*5788*/;
assign _361_ = _352_ & _360_ /*5786*/;
assign _324_ = _352_ ^ _360_ /*5787*/;
assign _358_ = _359_ | _361_ /*5784*/;
assign _363_ = ~Q[14] /*5783*/;
assign _362_ = _363_ & D[4] /*5782*/;
assign _365_ = _213_ & _362_ /*5777*/;
assign _366_ = _213_ ^ _362_ /*5780*/;
assign _367_ = _358_ & _366_ /*5778*/;
assign _325_ = _358_ ^ _366_ /*5779*/;
assign _364_ = _365_ | _367_ /*5776*/;
assign _369_ = ~Q[14] /*5775*/;
assign _368_ = _369_ & D[5] /*5774*/;
assign _371_ = _214_ & _368_ /*5769*/;
assign _372_ = _214_ ^ _368_ /*5772*/;
assign _373_ = _364_ & _372_ /*5770*/;
assign _326_ = _364_ ^ _372_ /*5771*/;
assign _370_ = _371_ | _373_ /*5768*/;
assign _375_ = ~Q[14] /*5767*/;
assign _374_ = _375_ & D[6] /*5766*/;
assign _377_ = _215_ & _374_ /*5761*/;
assign _378_ = _215_ ^ _374_ /*5764*/;
assign _379_ = _370_ & _378_ /*5762*/;
assign _327_ = _370_ ^ _378_ /*5763*/;
assign _376_ = _377_ | _379_ /*5760*/;
assign _381_ = ~Q[14] /*5759*/;
assign _380_ = _381_ & D[7] /*5758*/;
assign _383_ = _216_ & _380_ /*5753*/;
assign _384_ = _216_ ^ _380_ /*5756*/;
assign _385_ = _376_ & _384_ /*5754*/;
assign _328_ = _376_ ^ _384_ /*5755*/;
assign _382_ = _383_ | _385_ /*5752*/;
assign _387_ = ~Q[14] /*5751*/;
assign _386_ = _387_ & D[8] /*5750*/;
assign _389_ = _217_ & _386_ /*5745*/;
assign _390_ = _217_ ^ _386_ /*5748*/;
assign _391_ = _382_ & _390_ /*5746*/;
assign _329_ = _382_ ^ _390_ /*5747*/;
assign _388_ = _389_ | _391_ /*5744*/;
assign _393_ = ~Q[14] /*5743*/;
assign _392_ = _393_ & D[9] /*5742*/;
assign _395_ = _218_ & _392_ /*5737*/;
assign _396_ = _218_ ^ _392_ /*5740*/;
assign _397_ = _388_ & _396_ /*5738*/;
assign _330_ = _388_ ^ _396_ /*5739*/;
assign _394_ = _395_ | _397_ /*5736*/;
assign _399_ = ~Q[14] /*5735*/;
assign _398_ = _399_ & D[10] /*5734*/;
assign _401_ = _219_ & _398_ /*5729*/;
assign _402_ = _219_ ^ _398_ /*5732*/;
assign _403_ = _394_ & _402_ /*5730*/;
assign _331_ = _394_ ^ _402_ /*5731*/;
assign _400_ = _401_ | _403_ /*5728*/;
assign _405_ = ~Q[14] /*5727*/;
assign _404_ = _405_ & D[11] /*5726*/;
assign _407_ = _220_ & _404_ /*5721*/;
assign _408_ = _220_ ^ _404_ /*5724*/;
assign _409_ = _400_ & _408_ /*5722*/;
assign _332_ = _400_ ^ _408_ /*5723*/;
assign _406_ = _407_ | _409_ /*5720*/;
assign _411_ = ~Q[14] /*5719*/;
assign _410_ = _411_ & D[12] /*5718*/;
assign _413_ = _221_ & _410_ /*5713*/;
assign _414_ = _221_ ^ _410_ /*5716*/;
assign _415_ = _406_ & _414_ /*5714*/;
assign _333_ = _406_ ^ _414_ /*5715*/;
assign _412_ = _413_ | _415_ /*5712*/;
assign _417_ = ~Q[14] /*5711*/;
assign _416_ = _417_ & D[13] /*5710*/;
assign _419_ = _222_ & _416_ /*5705*/;
assign _420_ = _222_ ^ _416_ /*5708*/;
assign _421_ = _412_ & _420_ /*5706*/;
assign _334_ = _412_ ^ _420_ /*5707*/;
assign _418_ = _419_ | _421_ /*5704*/;
assign _423_ = ~Q[14] /*5703*/;
assign _422_ = _423_ & D[14] /*5702*/;
assign _425_ = _223_ & _422_ /*5697*/;
assign _426_ = _223_ ^ _422_ /*5700*/;
assign _427_ = _418_ & _426_ /*5698*/;
assign _335_ = _418_ ^ _426_ /*5699*/;
assign _424_ = _425_ | _427_ /*5696*/;
assign _429_ = ~Q[14] /*5695*/;
assign _428_ = _429_ & zeroWire /*5694*/;
assign _430_ = _224_ ^ _428_ /*5692*/;
assign _336_ = _430_ ^ _424_ /*5691*/;
assign _453_ = ~D[0] /*5629*/;
assign _450_ = R_0[13] & _453_ /*5625*/;
assign _451_ = R_0[13] ^ _453_ /*5628*/;
assign _452_ = oneWire & _451_ /*5626*/;
assign _433_ = oneWire ^ _451_ /*5627*/;
assign _449_ = _450_ | _452_ /*5624*/;
assign _458_ = ~D[1] /*5623*/;
assign _455_ = _321_ & _458_ /*5619*/;
assign _456_ = _321_ ^ _458_ /*5622*/;
assign _457_ = _449_ & _456_ /*5620*/;
assign _434_ = _449_ ^ _456_ /*5621*/;
assign _454_ = _455_ | _457_ /*5618*/;
assign _463_ = ~D[2] /*5617*/;
assign _460_ = _322_ & _463_ /*5613*/;
assign _461_ = _322_ ^ _463_ /*5616*/;
assign _462_ = _454_ & _461_ /*5614*/;
assign _435_ = _454_ ^ _461_ /*5615*/;
assign _459_ = _460_ | _462_ /*5612*/;
assign _468_ = ~D[3] /*5611*/;
assign _465_ = _323_ & _468_ /*5607*/;
assign _466_ = _323_ ^ _468_ /*5610*/;
assign _467_ = _459_ & _466_ /*5608*/;
assign _436_ = _459_ ^ _466_ /*5609*/;
assign _464_ = _465_ | _467_ /*5606*/;
assign _473_ = ~D[4] /*5605*/;
assign _470_ = _324_ & _473_ /*5601*/;
assign _471_ = _324_ ^ _473_ /*5604*/;
assign _472_ = _464_ & _471_ /*5602*/;
assign _437_ = _464_ ^ _471_ /*5603*/;
assign _469_ = _470_ | _472_ /*5600*/;
assign _478_ = ~D[5] /*5599*/;
assign _475_ = _325_ & _478_ /*5595*/;
assign _476_ = _325_ ^ _478_ /*5598*/;
assign _477_ = _469_ & _476_ /*5596*/;
assign _438_ = _469_ ^ _476_ /*5597*/;
assign _474_ = _475_ | _477_ /*5594*/;
assign _483_ = ~D[6] /*5593*/;
assign _480_ = _326_ & _483_ /*5589*/;
assign _481_ = _326_ ^ _483_ /*5592*/;
assign _482_ = _474_ & _481_ /*5590*/;
assign _439_ = _474_ ^ _481_ /*5591*/;
assign _479_ = _480_ | _482_ /*5588*/;
assign _488_ = ~D[7] /*5587*/;
assign _485_ = _327_ & _488_ /*5583*/;
assign _486_ = _327_ ^ _488_ /*5586*/;
assign _487_ = _479_ & _486_ /*5584*/;
assign _440_ = _479_ ^ _486_ /*5585*/;
assign _484_ = _485_ | _487_ /*5582*/;
assign _493_ = ~D[8] /*5581*/;
assign _490_ = _328_ & _493_ /*5577*/;
assign _491_ = _328_ ^ _493_ /*5580*/;
assign _492_ = _484_ & _491_ /*5578*/;
assign _441_ = _484_ ^ _491_ /*5579*/;
assign _489_ = _490_ | _492_ /*5576*/;
assign _498_ = ~D[9] /*5575*/;
assign _495_ = _329_ & _498_ /*5571*/;
assign _496_ = _329_ ^ _498_ /*5574*/;
assign _497_ = _489_ & _496_ /*5572*/;
assign _442_ = _489_ ^ _496_ /*5573*/;
assign _494_ = _495_ | _497_ /*5570*/;
assign _503_ = ~D[10] /*5569*/;
assign _500_ = _330_ & _503_ /*5565*/;
assign _501_ = _330_ ^ _503_ /*5568*/;
assign _502_ = _494_ & _501_ /*5566*/;
assign _443_ = _494_ ^ _501_ /*5567*/;
assign _499_ = _500_ | _502_ /*5564*/;
assign _508_ = ~D[11] /*5563*/;
assign _505_ = _331_ & _508_ /*5559*/;
assign _506_ = _331_ ^ _508_ /*5562*/;
assign _507_ = _499_ & _506_ /*5560*/;
assign _444_ = _499_ ^ _506_ /*5561*/;
assign _504_ = _505_ | _507_ /*5558*/;
assign _513_ = ~D[12] /*5557*/;
assign _510_ = _332_ & _513_ /*5553*/;
assign _511_ = _332_ ^ _513_ /*5556*/;
assign _512_ = _504_ & _511_ /*5554*/;
assign _445_ = _504_ ^ _511_ /*5555*/;
assign _509_ = _510_ | _512_ /*5552*/;
assign _518_ = ~D[13] /*5551*/;
assign _515_ = _333_ & _518_ /*5547*/;
assign _516_ = _333_ ^ _518_ /*5550*/;
assign _517_ = _509_ & _516_ /*5548*/;
assign _446_ = _509_ ^ _516_ /*5549*/;
assign _514_ = _515_ | _517_ /*5546*/;
assign _523_ = ~D[14] /*5545*/;
assign _520_ = _334_ & _523_ /*5541*/;
assign _521_ = _334_ ^ _523_ /*5544*/;
assign _522_ = _514_ & _521_ /*5542*/;
assign _447_ = _514_ ^ _521_ /*5543*/;
assign _519_ = _520_ | _522_ /*5540*/;
assign _524_ = _335_ & oneWire /*5535*/;
assign _525_ = _335_ ^ oneWire /*5538*/;
assign _526_ = _519_ & _525_ /*5536*/;
assign _448_ = _519_ ^ _525_ /*5537*/;
assign Q[13] = _524_ | _526_ /*5534*/;
assign _563_ = ~Q[13] /*5437*/;
assign _562_ = _563_ & D[0] /*5436*/;
assign _565_ = _433_ & _562_ /*5431*/;
assign _566_ = _433_ ^ _562_ /*5434*/;
assign _567_ = zeroWire & _566_ /*5432*/;
assign _545_ = zeroWire ^ _566_ /*5433*/;
assign _564_ = _565_ | _567_ /*5430*/;
assign _569_ = ~Q[13] /*5429*/;
assign _568_ = _569_ & D[1] /*5428*/;
assign _571_ = _434_ & _568_ /*5423*/;
assign _572_ = _434_ ^ _568_ /*5426*/;
assign _573_ = _564_ & _572_ /*5424*/;
assign _546_ = _564_ ^ _572_ /*5425*/;
assign _570_ = _571_ | _573_ /*5422*/;
assign _575_ = ~Q[13] /*5421*/;
assign _574_ = _575_ & D[2] /*5420*/;
assign _577_ = _435_ & _574_ /*5415*/;
assign _578_ = _435_ ^ _574_ /*5418*/;
assign _579_ = _570_ & _578_ /*5416*/;
assign _547_ = _570_ ^ _578_ /*5417*/;
assign _576_ = _577_ | _579_ /*5414*/;
assign _581_ = ~Q[13] /*5413*/;
assign _580_ = _581_ & D[3] /*5412*/;
assign _583_ = _436_ & _580_ /*5407*/;
assign _584_ = _436_ ^ _580_ /*5410*/;
assign _585_ = _576_ & _584_ /*5408*/;
assign _548_ = _576_ ^ _584_ /*5409*/;
assign _582_ = _583_ | _585_ /*5406*/;
assign _587_ = ~Q[13] /*5405*/;
assign _586_ = _587_ & D[4] /*5404*/;
assign _589_ = _437_ & _586_ /*5399*/;
assign _590_ = _437_ ^ _586_ /*5402*/;
assign _591_ = _582_ & _590_ /*5400*/;
assign _549_ = _582_ ^ _590_ /*5401*/;
assign _588_ = _589_ | _591_ /*5398*/;
assign _593_ = ~Q[13] /*5397*/;
assign _592_ = _593_ & D[5] /*5396*/;
assign _595_ = _438_ & _592_ /*5391*/;
assign _596_ = _438_ ^ _592_ /*5394*/;
assign _597_ = _588_ & _596_ /*5392*/;
assign _550_ = _588_ ^ _596_ /*5393*/;
assign _594_ = _595_ | _597_ /*5390*/;
assign _599_ = ~Q[13] /*5389*/;
assign _598_ = _599_ & D[6] /*5388*/;
assign _601_ = _439_ & _598_ /*5383*/;
assign _602_ = _439_ ^ _598_ /*5386*/;
assign _603_ = _594_ & _602_ /*5384*/;
assign _551_ = _594_ ^ _602_ /*5385*/;
assign _600_ = _601_ | _603_ /*5382*/;
assign _605_ = ~Q[13] /*5381*/;
assign _604_ = _605_ & D[7] /*5380*/;
assign _607_ = _440_ & _604_ /*5375*/;
assign _608_ = _440_ ^ _604_ /*5378*/;
assign _609_ = _600_ & _608_ /*5376*/;
assign _552_ = _600_ ^ _608_ /*5377*/;
assign _606_ = _607_ | _609_ /*5374*/;
assign _611_ = ~Q[13] /*5373*/;
assign _610_ = _611_ & D[8] /*5372*/;
assign _613_ = _441_ & _610_ /*5367*/;
assign _614_ = _441_ ^ _610_ /*5370*/;
assign _615_ = _606_ & _614_ /*5368*/;
assign _553_ = _606_ ^ _614_ /*5369*/;
assign _612_ = _613_ | _615_ /*5366*/;
assign _617_ = ~Q[13] /*5365*/;
assign _616_ = _617_ & D[9] /*5364*/;
assign _619_ = _442_ & _616_ /*5359*/;
assign _620_ = _442_ ^ _616_ /*5362*/;
assign _621_ = _612_ & _620_ /*5360*/;
assign _554_ = _612_ ^ _620_ /*5361*/;
assign _618_ = _619_ | _621_ /*5358*/;
assign _623_ = ~Q[13] /*5357*/;
assign _622_ = _623_ & D[10] /*5356*/;
assign _625_ = _443_ & _622_ /*5351*/;
assign _626_ = _443_ ^ _622_ /*5354*/;
assign _627_ = _618_ & _626_ /*5352*/;
assign _555_ = _618_ ^ _626_ /*5353*/;
assign _624_ = _625_ | _627_ /*5350*/;
assign _629_ = ~Q[13] /*5349*/;
assign _628_ = _629_ & D[11] /*5348*/;
assign _631_ = _444_ & _628_ /*5343*/;
assign _632_ = _444_ ^ _628_ /*5346*/;
assign _633_ = _624_ & _632_ /*5344*/;
assign _556_ = _624_ ^ _632_ /*5345*/;
assign _630_ = _631_ | _633_ /*5342*/;
assign _635_ = ~Q[13] /*5341*/;
assign _634_ = _635_ & D[12] /*5340*/;
assign _637_ = _445_ & _634_ /*5335*/;
assign _638_ = _445_ ^ _634_ /*5338*/;
assign _639_ = _630_ & _638_ /*5336*/;
assign _557_ = _630_ ^ _638_ /*5337*/;
assign _636_ = _637_ | _639_ /*5334*/;
assign _641_ = ~Q[13] /*5333*/;
assign _640_ = _641_ & D[13] /*5332*/;
assign _643_ = _446_ & _640_ /*5327*/;
assign _644_ = _446_ ^ _640_ /*5330*/;
assign _645_ = _636_ & _644_ /*5328*/;
assign _558_ = _636_ ^ _644_ /*5329*/;
assign _642_ = _643_ | _645_ /*5326*/;
assign _647_ = ~Q[13] /*5325*/;
assign _646_ = _647_ & D[14] /*5324*/;
assign _649_ = _447_ & _646_ /*5319*/;
assign _650_ = _447_ ^ _646_ /*5322*/;
assign _651_ = _642_ & _650_ /*5320*/;
assign _559_ = _642_ ^ _650_ /*5321*/;
assign _648_ = _649_ | _651_ /*5318*/;
assign _653_ = ~Q[13] /*5317*/;
assign _652_ = _653_ & zeroWire /*5316*/;
assign _654_ = _448_ ^ _652_ /*5314*/;
assign _560_ = _654_ ^ _648_ /*5313*/;
assign _677_ = ~D[0] /*5251*/;
assign _674_ = R_0[12] & _677_ /*5247*/;
assign _675_ = R_0[12] ^ _677_ /*5250*/;
assign _676_ = oneWire & _675_ /*5248*/;
assign _657_ = oneWire ^ _675_ /*5249*/;
assign _673_ = _674_ | _676_ /*5246*/;
assign _682_ = ~D[1] /*5245*/;
assign _679_ = _545_ & _682_ /*5241*/;
assign _680_ = _545_ ^ _682_ /*5244*/;
assign _681_ = _673_ & _680_ /*5242*/;
assign _658_ = _673_ ^ _680_ /*5243*/;
assign _678_ = _679_ | _681_ /*5240*/;
assign _687_ = ~D[2] /*5239*/;
assign _684_ = _546_ & _687_ /*5235*/;
assign _685_ = _546_ ^ _687_ /*5238*/;
assign _686_ = _678_ & _685_ /*5236*/;
assign _659_ = _678_ ^ _685_ /*5237*/;
assign _683_ = _684_ | _686_ /*5234*/;
assign _692_ = ~D[3] /*5233*/;
assign _689_ = _547_ & _692_ /*5229*/;
assign _690_ = _547_ ^ _692_ /*5232*/;
assign _691_ = _683_ & _690_ /*5230*/;
assign _660_ = _683_ ^ _690_ /*5231*/;
assign _688_ = _689_ | _691_ /*5228*/;
assign _697_ = ~D[4] /*5227*/;
assign _694_ = _548_ & _697_ /*5223*/;
assign _695_ = _548_ ^ _697_ /*5226*/;
assign _696_ = _688_ & _695_ /*5224*/;
assign _661_ = _688_ ^ _695_ /*5225*/;
assign _693_ = _694_ | _696_ /*5222*/;
assign _702_ = ~D[5] /*5221*/;
assign _699_ = _549_ & _702_ /*5217*/;
assign _700_ = _549_ ^ _702_ /*5220*/;
assign _701_ = _693_ & _700_ /*5218*/;
assign _662_ = _693_ ^ _700_ /*5219*/;
assign _698_ = _699_ | _701_ /*5216*/;
assign _707_ = ~D[6] /*5215*/;
assign _704_ = _550_ & _707_ /*5211*/;
assign _705_ = _550_ ^ _707_ /*5214*/;
assign _706_ = _698_ & _705_ /*5212*/;
assign _663_ = _698_ ^ _705_ /*5213*/;
assign _703_ = _704_ | _706_ /*5210*/;
assign _712_ = ~D[7] /*5209*/;
assign _709_ = _551_ & _712_ /*5205*/;
assign _710_ = _551_ ^ _712_ /*5208*/;
assign _711_ = _703_ & _710_ /*5206*/;
assign _664_ = _703_ ^ _710_ /*5207*/;
assign _708_ = _709_ | _711_ /*5204*/;
assign _717_ = ~D[8] /*5203*/;
assign _714_ = _552_ & _717_ /*5199*/;
assign _715_ = _552_ ^ _717_ /*5202*/;
assign _716_ = _708_ & _715_ /*5200*/;
assign _665_ = _708_ ^ _715_ /*5201*/;
assign _713_ = _714_ | _716_ /*5198*/;
assign _722_ = ~D[9] /*5197*/;
assign _719_ = _553_ & _722_ /*5193*/;
assign _720_ = _553_ ^ _722_ /*5196*/;
assign _721_ = _713_ & _720_ /*5194*/;
assign _666_ = _713_ ^ _720_ /*5195*/;
assign _718_ = _719_ | _721_ /*5192*/;
assign _727_ = ~D[10] /*5191*/;
assign _724_ = _554_ & _727_ /*5187*/;
assign _725_ = _554_ ^ _727_ /*5190*/;
assign _726_ = _718_ & _725_ /*5188*/;
assign _667_ = _718_ ^ _725_ /*5189*/;
assign _723_ = _724_ | _726_ /*5186*/;
assign _732_ = ~D[11] /*5185*/;
assign _729_ = _555_ & _732_ /*5181*/;
assign _730_ = _555_ ^ _732_ /*5184*/;
assign _731_ = _723_ & _730_ /*5182*/;
assign _668_ = _723_ ^ _730_ /*5183*/;
assign _728_ = _729_ | _731_ /*5180*/;
assign _737_ = ~D[12] /*5179*/;
assign _734_ = _556_ & _737_ /*5175*/;
assign _735_ = _556_ ^ _737_ /*5178*/;
assign _736_ = _728_ & _735_ /*5176*/;
assign _669_ = _728_ ^ _735_ /*5177*/;
assign _733_ = _734_ | _736_ /*5174*/;
assign _742_ = ~D[13] /*5173*/;
assign _739_ = _557_ & _742_ /*5169*/;
assign _740_ = _557_ ^ _742_ /*5172*/;
assign _741_ = _733_ & _740_ /*5170*/;
assign _670_ = _733_ ^ _740_ /*5171*/;
assign _738_ = _739_ | _741_ /*5168*/;
assign _747_ = ~D[14] /*5167*/;
assign _744_ = _558_ & _747_ /*5163*/;
assign _745_ = _558_ ^ _747_ /*5166*/;
assign _746_ = _738_ & _745_ /*5164*/;
assign _671_ = _738_ ^ _745_ /*5165*/;
assign _743_ = _744_ | _746_ /*5162*/;
assign _748_ = _559_ & oneWire /*5157*/;
assign _749_ = _559_ ^ oneWire /*5160*/;
assign _750_ = _743_ & _749_ /*5158*/;
assign _672_ = _743_ ^ _749_ /*5159*/;
assign Q[12] = _748_ | _750_ /*5156*/;
assign _787_ = ~Q[12] /*5059*/;
assign _786_ = _787_ & D[0] /*5058*/;
assign _789_ = _657_ & _786_ /*5053*/;
assign _790_ = _657_ ^ _786_ /*5056*/;
assign _791_ = zeroWire & _790_ /*5054*/;
assign _769_ = zeroWire ^ _790_ /*5055*/;
assign _788_ = _789_ | _791_ /*5052*/;
assign _793_ = ~Q[12] /*5051*/;
assign _792_ = _793_ & D[1] /*5050*/;
assign _795_ = _658_ & _792_ /*5045*/;
assign _796_ = _658_ ^ _792_ /*5048*/;
assign _797_ = _788_ & _796_ /*5046*/;
assign _770_ = _788_ ^ _796_ /*5047*/;
assign _794_ = _795_ | _797_ /*5044*/;
assign _799_ = ~Q[12] /*5043*/;
assign _798_ = _799_ & D[2] /*5042*/;
assign _801_ = _659_ & _798_ /*5037*/;
assign _802_ = _659_ ^ _798_ /*5040*/;
assign _803_ = _794_ & _802_ /*5038*/;
assign _771_ = _794_ ^ _802_ /*5039*/;
assign _800_ = _801_ | _803_ /*5036*/;
assign _805_ = ~Q[12] /*5035*/;
assign _804_ = _805_ & D[3] /*5034*/;
assign _807_ = _660_ & _804_ /*5029*/;
assign _808_ = _660_ ^ _804_ /*5032*/;
assign _809_ = _800_ & _808_ /*5030*/;
assign _772_ = _800_ ^ _808_ /*5031*/;
assign _806_ = _807_ | _809_ /*5028*/;
assign _811_ = ~Q[12] /*5027*/;
assign _810_ = _811_ & D[4] /*5026*/;
assign _813_ = _661_ & _810_ /*5021*/;
assign _814_ = _661_ ^ _810_ /*5024*/;
assign _815_ = _806_ & _814_ /*5022*/;
assign _773_ = _806_ ^ _814_ /*5023*/;
assign _812_ = _813_ | _815_ /*5020*/;
assign _817_ = ~Q[12] /*5019*/;
assign _816_ = _817_ & D[5] /*5018*/;
assign _819_ = _662_ & _816_ /*5013*/;
assign _820_ = _662_ ^ _816_ /*5016*/;
assign _821_ = _812_ & _820_ /*5014*/;
assign _774_ = _812_ ^ _820_ /*5015*/;
assign _818_ = _819_ | _821_ /*5012*/;
assign _823_ = ~Q[12] /*5011*/;
assign _822_ = _823_ & D[6] /*5010*/;
assign _825_ = _663_ & _822_ /*5005*/;
assign _826_ = _663_ ^ _822_ /*5008*/;
assign _827_ = _818_ & _826_ /*5006*/;
assign _775_ = _818_ ^ _826_ /*5007*/;
assign _824_ = _825_ | _827_ /*5004*/;
assign _829_ = ~Q[12] /*5003*/;
assign _828_ = _829_ & D[7] /*5002*/;
assign _831_ = _664_ & _828_ /*4997*/;
assign _832_ = _664_ ^ _828_ /*5000*/;
assign _833_ = _824_ & _832_ /*4998*/;
assign _776_ = _824_ ^ _832_ /*4999*/;
assign _830_ = _831_ | _833_ /*4996*/;
assign _835_ = ~Q[12] /*4995*/;
assign _834_ = _835_ & D[8] /*4994*/;
assign _837_ = _665_ & _834_ /*4989*/;
assign _838_ = _665_ ^ _834_ /*4992*/;
assign _839_ = _830_ & _838_ /*4990*/;
assign _777_ = _830_ ^ _838_ /*4991*/;
assign _836_ = _837_ | _839_ /*4988*/;
assign _841_ = ~Q[12] /*4987*/;
assign _840_ = _841_ & D[9] /*4986*/;
assign _843_ = _666_ & _840_ /*4981*/;
assign _844_ = _666_ ^ _840_ /*4984*/;
assign _845_ = _836_ & _844_ /*4982*/;
assign _778_ = _836_ ^ _844_ /*4983*/;
assign _842_ = _843_ | _845_ /*4980*/;
assign _847_ = ~Q[12] /*4979*/;
assign _846_ = _847_ & D[10] /*4978*/;
assign _849_ = _667_ & _846_ /*4973*/;
assign _850_ = _667_ ^ _846_ /*4976*/;
assign _851_ = _842_ & _850_ /*4974*/;
assign _779_ = _842_ ^ _850_ /*4975*/;
assign _848_ = _849_ | _851_ /*4972*/;
assign _853_ = ~Q[12] /*4971*/;
assign _852_ = _853_ & D[11] /*4970*/;
assign _855_ = _668_ & _852_ /*4965*/;
assign _856_ = _668_ ^ _852_ /*4968*/;
assign _857_ = _848_ & _856_ /*4966*/;
assign _780_ = _848_ ^ _856_ /*4967*/;
assign _854_ = _855_ | _857_ /*4964*/;
assign _859_ = ~Q[12] /*4963*/;
assign _858_ = _859_ & D[12] /*4962*/;
assign _861_ = _669_ & _858_ /*4957*/;
assign _862_ = _669_ ^ _858_ /*4960*/;
assign _863_ = _854_ & _862_ /*4958*/;
assign _781_ = _854_ ^ _862_ /*4959*/;
assign _860_ = _861_ | _863_ /*4956*/;
assign _865_ = ~Q[12] /*4955*/;
assign _864_ = _865_ & D[13] /*4954*/;
assign _867_ = _670_ & _864_ /*4949*/;
assign _868_ = _670_ ^ _864_ /*4952*/;
assign _869_ = _860_ & _868_ /*4950*/;
assign _782_ = _860_ ^ _868_ /*4951*/;
assign _866_ = _867_ | _869_ /*4948*/;
assign _871_ = ~Q[12] /*4947*/;
assign _870_ = _871_ & D[14] /*4946*/;
assign _873_ = _671_ & _870_ /*4941*/;
assign _874_ = _671_ ^ _870_ /*4944*/;
assign _875_ = _866_ & _874_ /*4942*/;
assign _783_ = _866_ ^ _874_ /*4943*/;
assign _872_ = _873_ | _875_ /*4940*/;
assign _877_ = ~Q[12] /*4939*/;
assign _876_ = _877_ & zeroWire /*4938*/;
assign _878_ = _672_ ^ _876_ /*4936*/;
assign _784_ = _878_ ^ _872_ /*4935*/;
assign _901_ = ~D[0] /*4873*/;
assign _898_ = R_0[11] & _901_ /*4869*/;
assign _899_ = R_0[11] ^ _901_ /*4872*/;
assign _900_ = oneWire & _899_ /*4870*/;
assign _881_ = oneWire ^ _899_ /*4871*/;
assign _897_ = _898_ | _900_ /*4868*/;
assign _906_ = ~D[1] /*4867*/;
assign _903_ = _769_ & _906_ /*4863*/;
assign _904_ = _769_ ^ _906_ /*4866*/;
assign _905_ = _897_ & _904_ /*4864*/;
assign _882_ = _897_ ^ _904_ /*4865*/;
assign _902_ = _903_ | _905_ /*4862*/;
assign _911_ = ~D[2] /*4861*/;
assign _908_ = _770_ & _911_ /*4857*/;
assign _909_ = _770_ ^ _911_ /*4860*/;
assign _910_ = _902_ & _909_ /*4858*/;
assign _883_ = _902_ ^ _909_ /*4859*/;
assign _907_ = _908_ | _910_ /*4856*/;
assign _916_ = ~D[3] /*4855*/;
assign _913_ = _771_ & _916_ /*4851*/;
assign _914_ = _771_ ^ _916_ /*4854*/;
assign _915_ = _907_ & _914_ /*4852*/;
assign _884_ = _907_ ^ _914_ /*4853*/;
assign _912_ = _913_ | _915_ /*4850*/;
assign _921_ = ~D[4] /*4849*/;
assign _918_ = _772_ & _921_ /*4845*/;
assign _919_ = _772_ ^ _921_ /*4848*/;
assign _920_ = _912_ & _919_ /*4846*/;
assign _885_ = _912_ ^ _919_ /*4847*/;
assign _917_ = _918_ | _920_ /*4844*/;
assign _926_ = ~D[5] /*4843*/;
assign _923_ = _773_ & _926_ /*4839*/;
assign _924_ = _773_ ^ _926_ /*4842*/;
assign _925_ = _917_ & _924_ /*4840*/;
assign _886_ = _917_ ^ _924_ /*4841*/;
assign _922_ = _923_ | _925_ /*4838*/;
assign _931_ = ~D[6] /*4837*/;
assign _928_ = _774_ & _931_ /*4833*/;
assign _929_ = _774_ ^ _931_ /*4836*/;
assign _930_ = _922_ & _929_ /*4834*/;
assign _887_ = _922_ ^ _929_ /*4835*/;
assign _927_ = _928_ | _930_ /*4832*/;
assign _936_ = ~D[7] /*4831*/;
assign _933_ = _775_ & _936_ /*4827*/;
assign _934_ = _775_ ^ _936_ /*4830*/;
assign _935_ = _927_ & _934_ /*4828*/;
assign _888_ = _927_ ^ _934_ /*4829*/;
assign _932_ = _933_ | _935_ /*4826*/;
assign _941_ = ~D[8] /*4825*/;
assign _938_ = _776_ & _941_ /*4821*/;
assign _939_ = _776_ ^ _941_ /*4824*/;
assign _940_ = _932_ & _939_ /*4822*/;
assign _889_ = _932_ ^ _939_ /*4823*/;
assign _937_ = _938_ | _940_ /*4820*/;
assign _946_ = ~D[9] /*4819*/;
assign _943_ = _777_ & _946_ /*4815*/;
assign _944_ = _777_ ^ _946_ /*4818*/;
assign _945_ = _937_ & _944_ /*4816*/;
assign _890_ = _937_ ^ _944_ /*4817*/;
assign _942_ = _943_ | _945_ /*4814*/;
assign _951_ = ~D[10] /*4813*/;
assign _948_ = _778_ & _951_ /*4809*/;
assign _949_ = _778_ ^ _951_ /*4812*/;
assign _950_ = _942_ & _949_ /*4810*/;
assign _891_ = _942_ ^ _949_ /*4811*/;
assign _947_ = _948_ | _950_ /*4808*/;
assign _956_ = ~D[11] /*4807*/;
assign _953_ = _779_ & _956_ /*4803*/;
assign _954_ = _779_ ^ _956_ /*4806*/;
assign _955_ = _947_ & _954_ /*4804*/;
assign _892_ = _947_ ^ _954_ /*4805*/;
assign _952_ = _953_ | _955_ /*4802*/;
assign _961_ = ~D[12] /*4801*/;
assign _958_ = _780_ & _961_ /*4797*/;
assign _959_ = _780_ ^ _961_ /*4800*/;
assign _960_ = _952_ & _959_ /*4798*/;
assign _893_ = _952_ ^ _959_ /*4799*/;
assign _957_ = _958_ | _960_ /*4796*/;
assign _966_ = ~D[13] /*4795*/;
assign _963_ = _781_ & _966_ /*4791*/;
assign _964_ = _781_ ^ _966_ /*4794*/;
assign _965_ = _957_ & _964_ /*4792*/;
assign _894_ = _957_ ^ _964_ /*4793*/;
assign _962_ = _963_ | _965_ /*4790*/;
assign _971_ = ~D[14] /*4789*/;
assign _968_ = _782_ & _971_ /*4785*/;
assign _969_ = _782_ ^ _971_ /*4788*/;
assign _970_ = _962_ & _969_ /*4786*/;
assign _895_ = _962_ ^ _969_ /*4787*/;
assign _967_ = _968_ | _970_ /*4784*/;
assign _972_ = _783_ & oneWire /*4779*/;
assign _973_ = _783_ ^ oneWire /*4782*/;
assign _974_ = _967_ & _973_ /*4780*/;
assign _896_ = _967_ ^ _973_ /*4781*/;
assign Q[11] = _972_ | _974_ /*4778*/;
assign _1011_ = ~Q[11] /*4681*/;
assign _1010_ = _1011_ & D[0] /*4680*/;
assign _1013_ = _881_ & _1010_ /*4675*/;
assign _1014_ = _881_ ^ _1010_ /*4678*/;
assign _1015_ = zeroWire & _1014_ /*4676*/;
assign _993_ = zeroWire ^ _1014_ /*4677*/;
assign _1012_ = _1013_ | _1015_ /*4674*/;
assign _1017_ = ~Q[11] /*4673*/;
assign _1016_ = _1017_ & D[1] /*4672*/;
assign _1019_ = _882_ & _1016_ /*4667*/;
assign _1020_ = _882_ ^ _1016_ /*4670*/;
assign _1021_ = _1012_ & _1020_ /*4668*/;
assign _994_ = _1012_ ^ _1020_ /*4669*/;
assign _1018_ = _1019_ | _1021_ /*4666*/;
assign _1023_ = ~Q[11] /*4665*/;
assign _1022_ = _1023_ & D[2] /*4664*/;
assign _1025_ = _883_ & _1022_ /*4659*/;
assign _1026_ = _883_ ^ _1022_ /*4662*/;
assign _1027_ = _1018_ & _1026_ /*4660*/;
assign _995_ = _1018_ ^ _1026_ /*4661*/;
assign _1024_ = _1025_ | _1027_ /*4658*/;
assign _1029_ = ~Q[11] /*4657*/;
assign _1028_ = _1029_ & D[3] /*4656*/;
assign _1031_ = _884_ & _1028_ /*4651*/;
assign _1032_ = _884_ ^ _1028_ /*4654*/;
assign _1033_ = _1024_ & _1032_ /*4652*/;
assign _996_ = _1024_ ^ _1032_ /*4653*/;
assign _1030_ = _1031_ | _1033_ /*4650*/;
assign _1035_ = ~Q[11] /*4649*/;
assign _1034_ = _1035_ & D[4] /*4648*/;
assign _1037_ = _885_ & _1034_ /*4643*/;
assign _1038_ = _885_ ^ _1034_ /*4646*/;
assign _1039_ = _1030_ & _1038_ /*4644*/;
assign _997_ = _1030_ ^ _1038_ /*4645*/;
assign _1036_ = _1037_ | _1039_ /*4642*/;
assign _1041_ = ~Q[11] /*4641*/;
assign _1040_ = _1041_ & D[5] /*4640*/;
assign _1043_ = _886_ & _1040_ /*4635*/;
assign _1044_ = _886_ ^ _1040_ /*4638*/;
assign _1045_ = _1036_ & _1044_ /*4636*/;
assign _998_ = _1036_ ^ _1044_ /*4637*/;
assign _1042_ = _1043_ | _1045_ /*4634*/;
assign _1047_ = ~Q[11] /*4633*/;
assign _1046_ = _1047_ & D[6] /*4632*/;
assign _1049_ = _887_ & _1046_ /*4627*/;
assign _1050_ = _887_ ^ _1046_ /*4630*/;
assign _1051_ = _1042_ & _1050_ /*4628*/;
assign _999_ = _1042_ ^ _1050_ /*4629*/;
assign _1048_ = _1049_ | _1051_ /*4626*/;
assign _1053_ = ~Q[11] /*4625*/;
assign _1052_ = _1053_ & D[7] /*4624*/;
assign _1055_ = _888_ & _1052_ /*4619*/;
assign _1056_ = _888_ ^ _1052_ /*4622*/;
assign _1057_ = _1048_ & _1056_ /*4620*/;
assign _1000_ = _1048_ ^ _1056_ /*4621*/;
assign _1054_ = _1055_ | _1057_ /*4618*/;
assign _1059_ = ~Q[11] /*4617*/;
assign _1058_ = _1059_ & D[8] /*4616*/;
assign _1061_ = _889_ & _1058_ /*4611*/;
assign _1062_ = _889_ ^ _1058_ /*4614*/;
assign _1063_ = _1054_ & _1062_ /*4612*/;
assign _1001_ = _1054_ ^ _1062_ /*4613*/;
assign _1060_ = _1061_ | _1063_ /*4610*/;
assign _1065_ = ~Q[11] /*4609*/;
assign _1064_ = _1065_ & D[9] /*4608*/;
assign _1067_ = _890_ & _1064_ /*4603*/;
assign _1068_ = _890_ ^ _1064_ /*4606*/;
assign _1069_ = _1060_ & _1068_ /*4604*/;
assign _1002_ = _1060_ ^ _1068_ /*4605*/;
assign _1066_ = _1067_ | _1069_ /*4602*/;
assign _1071_ = ~Q[11] /*4601*/;
assign _1070_ = _1071_ & D[10] /*4600*/;
assign _1073_ = _891_ & _1070_ /*4595*/;
assign _1074_ = _891_ ^ _1070_ /*4598*/;
assign _1075_ = _1066_ & _1074_ /*4596*/;
assign _1003_ = _1066_ ^ _1074_ /*4597*/;
assign _1072_ = _1073_ | _1075_ /*4594*/;
assign _1077_ = ~Q[11] /*4593*/;
assign _1076_ = _1077_ & D[11] /*4592*/;
assign _1079_ = _892_ & _1076_ /*4587*/;
assign _1080_ = _892_ ^ _1076_ /*4590*/;
assign _1081_ = _1072_ & _1080_ /*4588*/;
assign _1004_ = _1072_ ^ _1080_ /*4589*/;
assign _1078_ = _1079_ | _1081_ /*4586*/;
assign _1083_ = ~Q[11] /*4585*/;
assign _1082_ = _1083_ & D[12] /*4584*/;
assign _1085_ = _893_ & _1082_ /*4579*/;
assign _1086_ = _893_ ^ _1082_ /*4582*/;
assign _1087_ = _1078_ & _1086_ /*4580*/;
assign _1005_ = _1078_ ^ _1086_ /*4581*/;
assign _1084_ = _1085_ | _1087_ /*4578*/;
assign _1089_ = ~Q[11] /*4577*/;
assign _1088_ = _1089_ & D[13] /*4576*/;
assign _1091_ = _894_ & _1088_ /*4571*/;
assign _1092_ = _894_ ^ _1088_ /*4574*/;
assign _1093_ = _1084_ & _1092_ /*4572*/;
assign _1006_ = _1084_ ^ _1092_ /*4573*/;
assign _1090_ = _1091_ | _1093_ /*4570*/;
assign _1095_ = ~Q[11] /*4569*/;
assign _1094_ = _1095_ & D[14] /*4568*/;
assign _1097_ = _895_ & _1094_ /*4563*/;
assign _1098_ = _895_ ^ _1094_ /*4566*/;
assign _1099_ = _1090_ & _1098_ /*4564*/;
assign _1007_ = _1090_ ^ _1098_ /*4565*/;
assign _1096_ = _1097_ | _1099_ /*4562*/;
assign _1101_ = ~Q[11] /*4561*/;
assign _1100_ = _1101_ & zeroWire /*4560*/;
assign _1102_ = _896_ ^ _1100_ /*4558*/;
assign _1008_ = _1102_ ^ _1096_ /*4557*/;
assign _1125_ = ~D[0] /*4495*/;
assign _1122_ = R_0[10] & _1125_ /*4491*/;
assign _1123_ = R_0[10] ^ _1125_ /*4494*/;
assign _1124_ = oneWire & _1123_ /*4492*/;
assign _1105_ = oneWire ^ _1123_ /*4493*/;
assign _1121_ = _1122_ | _1124_ /*4490*/;
assign _1130_ = ~D[1] /*4489*/;
assign _1127_ = _993_ & _1130_ /*4485*/;
assign _1128_ = _993_ ^ _1130_ /*4488*/;
assign _1129_ = _1121_ & _1128_ /*4486*/;
assign _1106_ = _1121_ ^ _1128_ /*4487*/;
assign _1126_ = _1127_ | _1129_ /*4484*/;
assign _1135_ = ~D[2] /*4483*/;
assign _1132_ = _994_ & _1135_ /*4479*/;
assign _1133_ = _994_ ^ _1135_ /*4482*/;
assign _1134_ = _1126_ & _1133_ /*4480*/;
assign _1107_ = _1126_ ^ _1133_ /*4481*/;
assign _1131_ = _1132_ | _1134_ /*4478*/;
assign _1140_ = ~D[3] /*4477*/;
assign _1137_ = _995_ & _1140_ /*4473*/;
assign _1138_ = _995_ ^ _1140_ /*4476*/;
assign _1139_ = _1131_ & _1138_ /*4474*/;
assign _1108_ = _1131_ ^ _1138_ /*4475*/;
assign _1136_ = _1137_ | _1139_ /*4472*/;
assign _1145_ = ~D[4] /*4471*/;
assign _1142_ = _996_ & _1145_ /*4467*/;
assign _1143_ = _996_ ^ _1145_ /*4470*/;
assign _1144_ = _1136_ & _1143_ /*4468*/;
assign _1109_ = _1136_ ^ _1143_ /*4469*/;
assign _1141_ = _1142_ | _1144_ /*4466*/;
assign _1150_ = ~D[5] /*4465*/;
assign _1147_ = _997_ & _1150_ /*4461*/;
assign _1148_ = _997_ ^ _1150_ /*4464*/;
assign _1149_ = _1141_ & _1148_ /*4462*/;
assign _1110_ = _1141_ ^ _1148_ /*4463*/;
assign _1146_ = _1147_ | _1149_ /*4460*/;
assign _1155_ = ~D[6] /*4459*/;
assign _1152_ = _998_ & _1155_ /*4455*/;
assign _1153_ = _998_ ^ _1155_ /*4458*/;
assign _1154_ = _1146_ & _1153_ /*4456*/;
assign _1111_ = _1146_ ^ _1153_ /*4457*/;
assign _1151_ = _1152_ | _1154_ /*4454*/;
assign _1160_ = ~D[7] /*4453*/;
assign _1157_ = _999_ & _1160_ /*4449*/;
assign _1158_ = _999_ ^ _1160_ /*4452*/;
assign _1159_ = _1151_ & _1158_ /*4450*/;
assign _1112_ = _1151_ ^ _1158_ /*4451*/;
assign _1156_ = _1157_ | _1159_ /*4448*/;
assign _1165_ = ~D[8] /*4447*/;
assign _1162_ = _1000_ & _1165_ /*4443*/;
assign _1163_ = _1000_ ^ _1165_ /*4446*/;
assign _1164_ = _1156_ & _1163_ /*4444*/;
assign _1113_ = _1156_ ^ _1163_ /*4445*/;
assign _1161_ = _1162_ | _1164_ /*4442*/;
assign _1170_ = ~D[9] /*4441*/;
assign _1167_ = _1001_ & _1170_ /*4437*/;
assign _1168_ = _1001_ ^ _1170_ /*4440*/;
assign _1169_ = _1161_ & _1168_ /*4438*/;
assign _1114_ = _1161_ ^ _1168_ /*4439*/;
assign _1166_ = _1167_ | _1169_ /*4436*/;
assign _1175_ = ~D[10] /*4435*/;
assign _1172_ = _1002_ & _1175_ /*4431*/;
assign _1173_ = _1002_ ^ _1175_ /*4434*/;
assign _1174_ = _1166_ & _1173_ /*4432*/;
assign _1115_ = _1166_ ^ _1173_ /*4433*/;
assign _1171_ = _1172_ | _1174_ /*4430*/;
assign _1180_ = ~D[11] /*4429*/;
assign _1177_ = _1003_ & _1180_ /*4425*/;
assign _1178_ = _1003_ ^ _1180_ /*4428*/;
assign _1179_ = _1171_ & _1178_ /*4426*/;
assign _1116_ = _1171_ ^ _1178_ /*4427*/;
assign _1176_ = _1177_ | _1179_ /*4424*/;
assign _1185_ = ~D[12] /*4423*/;
assign _1182_ = _1004_ & _1185_ /*4419*/;
assign _1183_ = _1004_ ^ _1185_ /*4422*/;
assign _1184_ = _1176_ & _1183_ /*4420*/;
assign _1117_ = _1176_ ^ _1183_ /*4421*/;
assign _1181_ = _1182_ | _1184_ /*4418*/;
assign _1190_ = ~D[13] /*4417*/;
assign _1187_ = _1005_ & _1190_ /*4413*/;
assign _1188_ = _1005_ ^ _1190_ /*4416*/;
assign _1189_ = _1181_ & _1188_ /*4414*/;
assign _1118_ = _1181_ ^ _1188_ /*4415*/;
assign _1186_ = _1187_ | _1189_ /*4412*/;
assign _1195_ = ~D[14] /*4411*/;
assign _1192_ = _1006_ & _1195_ /*4407*/;
assign _1193_ = _1006_ ^ _1195_ /*4410*/;
assign _1194_ = _1186_ & _1193_ /*4408*/;
assign _1119_ = _1186_ ^ _1193_ /*4409*/;
assign _1191_ = _1192_ | _1194_ /*4406*/;
assign _1196_ = _1007_ & oneWire /*4401*/;
assign _1197_ = _1007_ ^ oneWire /*4404*/;
assign _1198_ = _1191_ & _1197_ /*4402*/;
assign _1120_ = _1191_ ^ _1197_ /*4403*/;
assign Q[10] = _1196_ | _1198_ /*4400*/;
assign _1235_ = ~Q[10] /*4303*/;
assign _1234_ = _1235_ & D[0] /*4302*/;
assign _1237_ = _1105_ & _1234_ /*4297*/;
assign _1238_ = _1105_ ^ _1234_ /*4300*/;
assign _1239_ = zeroWire & _1238_ /*4298*/;
assign _1217_ = zeroWire ^ _1238_ /*4299*/;
assign _1236_ = _1237_ | _1239_ /*4296*/;
assign _1241_ = ~Q[10] /*4295*/;
assign _1240_ = _1241_ & D[1] /*4294*/;
assign _1243_ = _1106_ & _1240_ /*4289*/;
assign _1244_ = _1106_ ^ _1240_ /*4292*/;
assign _1245_ = _1236_ & _1244_ /*4290*/;
assign _1218_ = _1236_ ^ _1244_ /*4291*/;
assign _1242_ = _1243_ | _1245_ /*4288*/;
assign _1247_ = ~Q[10] /*4287*/;
assign _1246_ = _1247_ & D[2] /*4286*/;
assign _1249_ = _1107_ & _1246_ /*4281*/;
assign _1250_ = _1107_ ^ _1246_ /*4284*/;
assign _1251_ = _1242_ & _1250_ /*4282*/;
assign _1219_ = _1242_ ^ _1250_ /*4283*/;
assign _1248_ = _1249_ | _1251_ /*4280*/;
assign _1253_ = ~Q[10] /*4279*/;
assign _1252_ = _1253_ & D[3] /*4278*/;
assign _1255_ = _1108_ & _1252_ /*4273*/;
assign _1256_ = _1108_ ^ _1252_ /*4276*/;
assign _1257_ = _1248_ & _1256_ /*4274*/;
assign _1220_ = _1248_ ^ _1256_ /*4275*/;
assign _1254_ = _1255_ | _1257_ /*4272*/;
assign _1259_ = ~Q[10] /*4271*/;
assign _1258_ = _1259_ & D[4] /*4270*/;
assign _1261_ = _1109_ & _1258_ /*4265*/;
assign _1262_ = _1109_ ^ _1258_ /*4268*/;
assign _1263_ = _1254_ & _1262_ /*4266*/;
assign _1221_ = _1254_ ^ _1262_ /*4267*/;
assign _1260_ = _1261_ | _1263_ /*4264*/;
assign _1265_ = ~Q[10] /*4263*/;
assign _1264_ = _1265_ & D[5] /*4262*/;
assign _1267_ = _1110_ & _1264_ /*4257*/;
assign _1268_ = _1110_ ^ _1264_ /*4260*/;
assign _1269_ = _1260_ & _1268_ /*4258*/;
assign _1222_ = _1260_ ^ _1268_ /*4259*/;
assign _1266_ = _1267_ | _1269_ /*4256*/;
assign _1271_ = ~Q[10] /*4255*/;
assign _1270_ = _1271_ & D[6] /*4254*/;
assign _1273_ = _1111_ & _1270_ /*4249*/;
assign _1274_ = _1111_ ^ _1270_ /*4252*/;
assign _1275_ = _1266_ & _1274_ /*4250*/;
assign _1223_ = _1266_ ^ _1274_ /*4251*/;
assign _1272_ = _1273_ | _1275_ /*4248*/;
assign _1277_ = ~Q[10] /*4247*/;
assign _1276_ = _1277_ & D[7] /*4246*/;
assign _1279_ = _1112_ & _1276_ /*4241*/;
assign _1280_ = _1112_ ^ _1276_ /*4244*/;
assign _1281_ = _1272_ & _1280_ /*4242*/;
assign _1224_ = _1272_ ^ _1280_ /*4243*/;
assign _1278_ = _1279_ | _1281_ /*4240*/;
assign _1283_ = ~Q[10] /*4239*/;
assign _1282_ = _1283_ & D[8] /*4238*/;
assign _1285_ = _1113_ & _1282_ /*4233*/;
assign _1286_ = _1113_ ^ _1282_ /*4236*/;
assign _1287_ = _1278_ & _1286_ /*4234*/;
assign _1225_ = _1278_ ^ _1286_ /*4235*/;
assign _1284_ = _1285_ | _1287_ /*4232*/;
assign _1289_ = ~Q[10] /*4231*/;
assign _1288_ = _1289_ & D[9] /*4230*/;
assign _1291_ = _1114_ & _1288_ /*4225*/;
assign _1292_ = _1114_ ^ _1288_ /*4228*/;
assign _1293_ = _1284_ & _1292_ /*4226*/;
assign _1226_ = _1284_ ^ _1292_ /*4227*/;
assign _1290_ = _1291_ | _1293_ /*4224*/;
assign _1295_ = ~Q[10] /*4223*/;
assign _1294_ = _1295_ & D[10] /*4222*/;
assign _1297_ = _1115_ & _1294_ /*4217*/;
assign _1298_ = _1115_ ^ _1294_ /*4220*/;
assign _1299_ = _1290_ & _1298_ /*4218*/;
assign _1227_ = _1290_ ^ _1298_ /*4219*/;
assign _1296_ = _1297_ | _1299_ /*4216*/;
assign _1301_ = ~Q[10] /*4215*/;
assign _1300_ = _1301_ & D[11] /*4214*/;
assign _1303_ = _1116_ & _1300_ /*4209*/;
assign _1304_ = _1116_ ^ _1300_ /*4212*/;
assign _1305_ = _1296_ & _1304_ /*4210*/;
assign _1228_ = _1296_ ^ _1304_ /*4211*/;
assign _1302_ = _1303_ | _1305_ /*4208*/;
assign _1307_ = ~Q[10] /*4207*/;
assign _1306_ = _1307_ & D[12] /*4206*/;
assign _1309_ = _1117_ & _1306_ /*4201*/;
assign _1310_ = _1117_ ^ _1306_ /*4204*/;
assign _1311_ = _1302_ & _1310_ /*4202*/;
assign _1229_ = _1302_ ^ _1310_ /*4203*/;
assign _1308_ = _1309_ | _1311_ /*4200*/;
assign _1313_ = ~Q[10] /*4199*/;
assign _1312_ = _1313_ & D[13] /*4198*/;
assign _1315_ = _1118_ & _1312_ /*4193*/;
assign _1316_ = _1118_ ^ _1312_ /*4196*/;
assign _1317_ = _1308_ & _1316_ /*4194*/;
assign _1230_ = _1308_ ^ _1316_ /*4195*/;
assign _1314_ = _1315_ | _1317_ /*4192*/;
assign _1319_ = ~Q[10] /*4191*/;
assign _1318_ = _1319_ & D[14] /*4190*/;
assign _1321_ = _1119_ & _1318_ /*4185*/;
assign _1322_ = _1119_ ^ _1318_ /*4188*/;
assign _1323_ = _1314_ & _1322_ /*4186*/;
assign _1231_ = _1314_ ^ _1322_ /*4187*/;
assign _1320_ = _1321_ | _1323_ /*4184*/;
assign _1325_ = ~Q[10] /*4183*/;
assign _1324_ = _1325_ & zeroWire /*4182*/;
assign _1326_ = _1120_ ^ _1324_ /*4180*/;
assign _1232_ = _1326_ ^ _1320_ /*4179*/;
assign _1349_ = ~D[0] /*4117*/;
assign _1346_ = R_0[9] & _1349_ /*4113*/;
assign _1347_ = R_0[9] ^ _1349_ /*4116*/;
assign _1348_ = oneWire & _1347_ /*4114*/;
assign _1329_ = oneWire ^ _1347_ /*4115*/;
assign _1345_ = _1346_ | _1348_ /*4112*/;
assign _1354_ = ~D[1] /*4111*/;
assign _1351_ = _1217_ & _1354_ /*4107*/;
assign _1352_ = _1217_ ^ _1354_ /*4110*/;
assign _1353_ = _1345_ & _1352_ /*4108*/;
assign _1330_ = _1345_ ^ _1352_ /*4109*/;
assign _1350_ = _1351_ | _1353_ /*4106*/;
assign _1359_ = ~D[2] /*4105*/;
assign _1356_ = _1218_ & _1359_ /*4101*/;
assign _1357_ = _1218_ ^ _1359_ /*4104*/;
assign _1358_ = _1350_ & _1357_ /*4102*/;
assign _1331_ = _1350_ ^ _1357_ /*4103*/;
assign _1355_ = _1356_ | _1358_ /*4100*/;
assign _1364_ = ~D[3] /*4099*/;
assign _1361_ = _1219_ & _1364_ /*4095*/;
assign _1362_ = _1219_ ^ _1364_ /*4098*/;
assign _1363_ = _1355_ & _1362_ /*4096*/;
assign _1332_ = _1355_ ^ _1362_ /*4097*/;
assign _1360_ = _1361_ | _1363_ /*4094*/;
assign _1369_ = ~D[4] /*4093*/;
assign _1366_ = _1220_ & _1369_ /*4089*/;
assign _1367_ = _1220_ ^ _1369_ /*4092*/;
assign _1368_ = _1360_ & _1367_ /*4090*/;
assign _1333_ = _1360_ ^ _1367_ /*4091*/;
assign _1365_ = _1366_ | _1368_ /*4088*/;
assign _1374_ = ~D[5] /*4087*/;
assign _1371_ = _1221_ & _1374_ /*4083*/;
assign _1372_ = _1221_ ^ _1374_ /*4086*/;
assign _1373_ = _1365_ & _1372_ /*4084*/;
assign _1334_ = _1365_ ^ _1372_ /*4085*/;
assign _1370_ = _1371_ | _1373_ /*4082*/;
assign _1379_ = ~D[6] /*4081*/;
assign _1376_ = _1222_ & _1379_ /*4077*/;
assign _1377_ = _1222_ ^ _1379_ /*4080*/;
assign _1378_ = _1370_ & _1377_ /*4078*/;
assign _1335_ = _1370_ ^ _1377_ /*4079*/;
assign _1375_ = _1376_ | _1378_ /*4076*/;
assign _1384_ = ~D[7] /*4075*/;
assign _1381_ = _1223_ & _1384_ /*4071*/;
assign _1382_ = _1223_ ^ _1384_ /*4074*/;
assign _1383_ = _1375_ & _1382_ /*4072*/;
assign _1336_ = _1375_ ^ _1382_ /*4073*/;
assign _1380_ = _1381_ | _1383_ /*4070*/;
assign _1389_ = ~D[8] /*4069*/;
assign _1386_ = _1224_ & _1389_ /*4065*/;
assign _1387_ = _1224_ ^ _1389_ /*4068*/;
assign _1388_ = _1380_ & _1387_ /*4066*/;
assign _1337_ = _1380_ ^ _1387_ /*4067*/;
assign _1385_ = _1386_ | _1388_ /*4064*/;
assign _1394_ = ~D[9] /*4063*/;
assign _1391_ = _1225_ & _1394_ /*4059*/;
assign _1392_ = _1225_ ^ _1394_ /*4062*/;
assign _1393_ = _1385_ & _1392_ /*4060*/;
assign _1338_ = _1385_ ^ _1392_ /*4061*/;
assign _1390_ = _1391_ | _1393_ /*4058*/;
assign _1399_ = ~D[10] /*4057*/;
assign _1396_ = _1226_ & _1399_ /*4053*/;
assign _1397_ = _1226_ ^ _1399_ /*4056*/;
assign _1398_ = _1390_ & _1397_ /*4054*/;
assign _1339_ = _1390_ ^ _1397_ /*4055*/;
assign _1395_ = _1396_ | _1398_ /*4052*/;
assign _1404_ = ~D[11] /*4051*/;
assign _1401_ = _1227_ & _1404_ /*4047*/;
assign _1402_ = _1227_ ^ _1404_ /*4050*/;
assign _1403_ = _1395_ & _1402_ /*4048*/;
assign _1340_ = _1395_ ^ _1402_ /*4049*/;
assign _1400_ = _1401_ | _1403_ /*4046*/;
assign _1409_ = ~D[12] /*4045*/;
assign _1406_ = _1228_ & _1409_ /*4041*/;
assign _1407_ = _1228_ ^ _1409_ /*4044*/;
assign _1408_ = _1400_ & _1407_ /*4042*/;
assign _1341_ = _1400_ ^ _1407_ /*4043*/;
assign _1405_ = _1406_ | _1408_ /*4040*/;
assign _1414_ = ~D[13] /*4039*/;
assign _1411_ = _1229_ & _1414_ /*4035*/;
assign _1412_ = _1229_ ^ _1414_ /*4038*/;
assign _1413_ = _1405_ & _1412_ /*4036*/;
assign _1342_ = _1405_ ^ _1412_ /*4037*/;
assign _1410_ = _1411_ | _1413_ /*4034*/;
assign _1419_ = ~D[14] /*4033*/;
assign _1416_ = _1230_ & _1419_ /*4029*/;
assign _1417_ = _1230_ ^ _1419_ /*4032*/;
assign _1418_ = _1410_ & _1417_ /*4030*/;
assign _1343_ = _1410_ ^ _1417_ /*4031*/;
assign _1415_ = _1416_ | _1418_ /*4028*/;
assign _1420_ = _1231_ & oneWire /*4023*/;
assign _1421_ = _1231_ ^ oneWire /*4026*/;
assign _1422_ = _1415_ & _1421_ /*4024*/;
assign _1344_ = _1415_ ^ _1421_ /*4025*/;
assign Q[9] = _1420_ | _1422_ /*4022*/;
assign _1459_ = ~Q[9] /*3925*/;
assign _1458_ = _1459_ & D[0] /*3924*/;
assign _1461_ = _1329_ & _1458_ /*3919*/;
assign _1462_ = _1329_ ^ _1458_ /*3922*/;
assign _1463_ = zeroWire & _1462_ /*3920*/;
assign _1441_ = zeroWire ^ _1462_ /*3921*/;
assign _1460_ = _1461_ | _1463_ /*3918*/;
assign _1465_ = ~Q[9] /*3917*/;
assign _1464_ = _1465_ & D[1] /*3916*/;
assign _1467_ = _1330_ & _1464_ /*3911*/;
assign _1468_ = _1330_ ^ _1464_ /*3914*/;
assign _1469_ = _1460_ & _1468_ /*3912*/;
assign _1442_ = _1460_ ^ _1468_ /*3913*/;
assign _1466_ = _1467_ | _1469_ /*3910*/;
assign _1471_ = ~Q[9] /*3909*/;
assign _1470_ = _1471_ & D[2] /*3908*/;
assign _1473_ = _1331_ & _1470_ /*3903*/;
assign _1474_ = _1331_ ^ _1470_ /*3906*/;
assign _1475_ = _1466_ & _1474_ /*3904*/;
assign _1443_ = _1466_ ^ _1474_ /*3905*/;
assign _1472_ = _1473_ | _1475_ /*3902*/;
assign _1477_ = ~Q[9] /*3901*/;
assign _1476_ = _1477_ & D[3] /*3900*/;
assign _1479_ = _1332_ & _1476_ /*3895*/;
assign _1480_ = _1332_ ^ _1476_ /*3898*/;
assign _1481_ = _1472_ & _1480_ /*3896*/;
assign _1444_ = _1472_ ^ _1480_ /*3897*/;
assign _1478_ = _1479_ | _1481_ /*3894*/;
assign _1483_ = ~Q[9] /*3893*/;
assign _1482_ = _1483_ & D[4] /*3892*/;
assign _1485_ = _1333_ & _1482_ /*3887*/;
assign _1486_ = _1333_ ^ _1482_ /*3890*/;
assign _1487_ = _1478_ & _1486_ /*3888*/;
assign _1445_ = _1478_ ^ _1486_ /*3889*/;
assign _1484_ = _1485_ | _1487_ /*3886*/;
assign _1489_ = ~Q[9] /*3885*/;
assign _1488_ = _1489_ & D[5] /*3884*/;
assign _1491_ = _1334_ & _1488_ /*3879*/;
assign _1492_ = _1334_ ^ _1488_ /*3882*/;
assign _1493_ = _1484_ & _1492_ /*3880*/;
assign _1446_ = _1484_ ^ _1492_ /*3881*/;
assign _1490_ = _1491_ | _1493_ /*3878*/;
assign _1495_ = ~Q[9] /*3877*/;
assign _1494_ = _1495_ & D[6] /*3876*/;
assign _1497_ = _1335_ & _1494_ /*3871*/;
assign _1498_ = _1335_ ^ _1494_ /*3874*/;
assign _1499_ = _1490_ & _1498_ /*3872*/;
assign _1447_ = _1490_ ^ _1498_ /*3873*/;
assign _1496_ = _1497_ | _1499_ /*3870*/;
assign _1501_ = ~Q[9] /*3869*/;
assign _1500_ = _1501_ & D[7] /*3868*/;
assign _1503_ = _1336_ & _1500_ /*3863*/;
assign _1504_ = _1336_ ^ _1500_ /*3866*/;
assign _1505_ = _1496_ & _1504_ /*3864*/;
assign _1448_ = _1496_ ^ _1504_ /*3865*/;
assign _1502_ = _1503_ | _1505_ /*3862*/;
assign _1507_ = ~Q[9] /*3861*/;
assign _1506_ = _1507_ & D[8] /*3860*/;
assign _1509_ = _1337_ & _1506_ /*3855*/;
assign _1510_ = _1337_ ^ _1506_ /*3858*/;
assign _1511_ = _1502_ & _1510_ /*3856*/;
assign _1449_ = _1502_ ^ _1510_ /*3857*/;
assign _1508_ = _1509_ | _1511_ /*3854*/;
assign _1513_ = ~Q[9] /*3853*/;
assign _1512_ = _1513_ & D[9] /*3852*/;
assign _1515_ = _1338_ & _1512_ /*3847*/;
assign _1516_ = _1338_ ^ _1512_ /*3850*/;
assign _1517_ = _1508_ & _1516_ /*3848*/;
assign _1450_ = _1508_ ^ _1516_ /*3849*/;
assign _1514_ = _1515_ | _1517_ /*3846*/;
assign _1519_ = ~Q[9] /*3845*/;
assign _1518_ = _1519_ & D[10] /*3844*/;
assign _1521_ = _1339_ & _1518_ /*3839*/;
assign _1522_ = _1339_ ^ _1518_ /*3842*/;
assign _1523_ = _1514_ & _1522_ /*3840*/;
assign _1451_ = _1514_ ^ _1522_ /*3841*/;
assign _1520_ = _1521_ | _1523_ /*3838*/;
assign _1525_ = ~Q[9] /*3837*/;
assign _1524_ = _1525_ & D[11] /*3836*/;
assign _1527_ = _1340_ & _1524_ /*3831*/;
assign _1528_ = _1340_ ^ _1524_ /*3834*/;
assign _1529_ = _1520_ & _1528_ /*3832*/;
assign _1452_ = _1520_ ^ _1528_ /*3833*/;
assign _1526_ = _1527_ | _1529_ /*3830*/;
assign _1531_ = ~Q[9] /*3829*/;
assign _1530_ = _1531_ & D[12] /*3828*/;
assign _1533_ = _1341_ & _1530_ /*3823*/;
assign _1534_ = _1341_ ^ _1530_ /*3826*/;
assign _1535_ = _1526_ & _1534_ /*3824*/;
assign _1453_ = _1526_ ^ _1534_ /*3825*/;
assign _1532_ = _1533_ | _1535_ /*3822*/;
assign _1537_ = ~Q[9] /*3821*/;
assign _1536_ = _1537_ & D[13] /*3820*/;
assign _1539_ = _1342_ & _1536_ /*3815*/;
assign _1540_ = _1342_ ^ _1536_ /*3818*/;
assign _1541_ = _1532_ & _1540_ /*3816*/;
assign _1454_ = _1532_ ^ _1540_ /*3817*/;
assign _1538_ = _1539_ | _1541_ /*3814*/;
assign _1543_ = ~Q[9] /*3813*/;
assign _1542_ = _1543_ & D[14] /*3812*/;
assign _1545_ = _1343_ & _1542_ /*3807*/;
assign _1546_ = _1343_ ^ _1542_ /*3810*/;
assign _1547_ = _1538_ & _1546_ /*3808*/;
assign _1455_ = _1538_ ^ _1546_ /*3809*/;
assign _1544_ = _1545_ | _1547_ /*3806*/;
assign _1549_ = ~Q[9] /*3805*/;
assign _1548_ = _1549_ & zeroWire /*3804*/;
assign _1550_ = _1344_ ^ _1548_ /*3802*/;
assign _1456_ = _1550_ ^ _1544_ /*3801*/;
assign _1573_ = ~D[0] /*3739*/;
assign _1570_ = R_0[8] & _1573_ /*3735*/;
assign _1571_ = R_0[8] ^ _1573_ /*3738*/;
assign _1572_ = oneWire & _1571_ /*3736*/;
assign _1553_ = oneWire ^ _1571_ /*3737*/;
assign _1569_ = _1570_ | _1572_ /*3734*/;
assign _1578_ = ~D[1] /*3733*/;
assign _1575_ = _1441_ & _1578_ /*3729*/;
assign _1576_ = _1441_ ^ _1578_ /*3732*/;
assign _1577_ = _1569_ & _1576_ /*3730*/;
assign _1554_ = _1569_ ^ _1576_ /*3731*/;
assign _1574_ = _1575_ | _1577_ /*3728*/;
assign _1583_ = ~D[2] /*3727*/;
assign _1580_ = _1442_ & _1583_ /*3723*/;
assign _1581_ = _1442_ ^ _1583_ /*3726*/;
assign _1582_ = _1574_ & _1581_ /*3724*/;
assign _1555_ = _1574_ ^ _1581_ /*3725*/;
assign _1579_ = _1580_ | _1582_ /*3722*/;
assign _1588_ = ~D[3] /*3721*/;
assign _1585_ = _1443_ & _1588_ /*3717*/;
assign _1586_ = _1443_ ^ _1588_ /*3720*/;
assign _1587_ = _1579_ & _1586_ /*3718*/;
assign _1556_ = _1579_ ^ _1586_ /*3719*/;
assign _1584_ = _1585_ | _1587_ /*3716*/;
assign _1593_ = ~D[4] /*3715*/;
assign _1590_ = _1444_ & _1593_ /*3711*/;
assign _1591_ = _1444_ ^ _1593_ /*3714*/;
assign _1592_ = _1584_ & _1591_ /*3712*/;
assign _1557_ = _1584_ ^ _1591_ /*3713*/;
assign _1589_ = _1590_ | _1592_ /*3710*/;
assign _1598_ = ~D[5] /*3709*/;
assign _1595_ = _1445_ & _1598_ /*3705*/;
assign _1596_ = _1445_ ^ _1598_ /*3708*/;
assign _1597_ = _1589_ & _1596_ /*3706*/;
assign _1558_ = _1589_ ^ _1596_ /*3707*/;
assign _1594_ = _1595_ | _1597_ /*3704*/;
assign _1603_ = ~D[6] /*3703*/;
assign _1600_ = _1446_ & _1603_ /*3699*/;
assign _1601_ = _1446_ ^ _1603_ /*3702*/;
assign _1602_ = _1594_ & _1601_ /*3700*/;
assign _1559_ = _1594_ ^ _1601_ /*3701*/;
assign _1599_ = _1600_ | _1602_ /*3698*/;
assign _1608_ = ~D[7] /*3697*/;
assign _1605_ = _1447_ & _1608_ /*3693*/;
assign _1606_ = _1447_ ^ _1608_ /*3696*/;
assign _1607_ = _1599_ & _1606_ /*3694*/;
assign _1560_ = _1599_ ^ _1606_ /*3695*/;
assign _1604_ = _1605_ | _1607_ /*3692*/;
assign _1613_ = ~D[8] /*3691*/;
assign _1610_ = _1448_ & _1613_ /*3687*/;
assign _1611_ = _1448_ ^ _1613_ /*3690*/;
assign _1612_ = _1604_ & _1611_ /*3688*/;
assign _1561_ = _1604_ ^ _1611_ /*3689*/;
assign _1609_ = _1610_ | _1612_ /*3686*/;
assign _1618_ = ~D[9] /*3685*/;
assign _1615_ = _1449_ & _1618_ /*3681*/;
assign _1616_ = _1449_ ^ _1618_ /*3684*/;
assign _1617_ = _1609_ & _1616_ /*3682*/;
assign _1562_ = _1609_ ^ _1616_ /*3683*/;
assign _1614_ = _1615_ | _1617_ /*3680*/;
assign _1623_ = ~D[10] /*3679*/;
assign _1620_ = _1450_ & _1623_ /*3675*/;
assign _1621_ = _1450_ ^ _1623_ /*3678*/;
assign _1622_ = _1614_ & _1621_ /*3676*/;
assign _1563_ = _1614_ ^ _1621_ /*3677*/;
assign _1619_ = _1620_ | _1622_ /*3674*/;
assign _1628_ = ~D[11] /*3673*/;
assign _1625_ = _1451_ & _1628_ /*3669*/;
assign _1626_ = _1451_ ^ _1628_ /*3672*/;
assign _1627_ = _1619_ & _1626_ /*3670*/;
assign _1564_ = _1619_ ^ _1626_ /*3671*/;
assign _1624_ = _1625_ | _1627_ /*3668*/;
assign _1633_ = ~D[12] /*3667*/;
assign _1630_ = _1452_ & _1633_ /*3663*/;
assign _1631_ = _1452_ ^ _1633_ /*3666*/;
assign _1632_ = _1624_ & _1631_ /*3664*/;
assign _1565_ = _1624_ ^ _1631_ /*3665*/;
assign _1629_ = _1630_ | _1632_ /*3662*/;
assign _1638_ = ~D[13] /*3661*/;
assign _1635_ = _1453_ & _1638_ /*3657*/;
assign _1636_ = _1453_ ^ _1638_ /*3660*/;
assign _1637_ = _1629_ & _1636_ /*3658*/;
assign _1566_ = _1629_ ^ _1636_ /*3659*/;
assign _1634_ = _1635_ | _1637_ /*3656*/;
assign _1643_ = ~D[14] /*3655*/;
assign _1640_ = _1454_ & _1643_ /*3651*/;
assign _1641_ = _1454_ ^ _1643_ /*3654*/;
assign _1642_ = _1634_ & _1641_ /*3652*/;
assign _1567_ = _1634_ ^ _1641_ /*3653*/;
assign _1639_ = _1640_ | _1642_ /*3650*/;
assign _1644_ = _1455_ & oneWire /*3645*/;
assign _1645_ = _1455_ ^ oneWire /*3648*/;
assign _1646_ = _1639_ & _1645_ /*3646*/;
assign _1568_ = _1639_ ^ _1645_ /*3647*/;
assign Q[8] = _1644_ | _1646_ /*3644*/;
assign _1683_ = ~Q[8] /*3547*/;
assign _1682_ = _1683_ & D[0] /*3546*/;
assign _1685_ = _1553_ & _1682_ /*3541*/;
assign _1686_ = _1553_ ^ _1682_ /*3544*/;
assign _1687_ = zeroWire & _1686_ /*3542*/;
assign _1665_ = zeroWire ^ _1686_ /*3543*/;
assign _1684_ = _1685_ | _1687_ /*3540*/;
assign _1689_ = ~Q[8] /*3539*/;
assign _1688_ = _1689_ & D[1] /*3538*/;
assign _1691_ = _1554_ & _1688_ /*3533*/;
assign _1692_ = _1554_ ^ _1688_ /*3536*/;
assign _1693_ = _1684_ & _1692_ /*3534*/;
assign _1666_ = _1684_ ^ _1692_ /*3535*/;
assign _1690_ = _1691_ | _1693_ /*3532*/;
assign _1695_ = ~Q[8] /*3531*/;
assign _1694_ = _1695_ & D[2] /*3530*/;
assign _1697_ = _1555_ & _1694_ /*3525*/;
assign _1698_ = _1555_ ^ _1694_ /*3528*/;
assign _1699_ = _1690_ & _1698_ /*3526*/;
assign _1667_ = _1690_ ^ _1698_ /*3527*/;
assign _1696_ = _1697_ | _1699_ /*3524*/;
assign _1701_ = ~Q[8] /*3523*/;
assign _1700_ = _1701_ & D[3] /*3522*/;
assign _1703_ = _1556_ & _1700_ /*3517*/;
assign _1704_ = _1556_ ^ _1700_ /*3520*/;
assign _1705_ = _1696_ & _1704_ /*3518*/;
assign _1668_ = _1696_ ^ _1704_ /*3519*/;
assign _1702_ = _1703_ | _1705_ /*3516*/;
assign _1707_ = ~Q[8] /*3515*/;
assign _1706_ = _1707_ & D[4] /*3514*/;
assign _1709_ = _1557_ & _1706_ /*3509*/;
assign _1710_ = _1557_ ^ _1706_ /*3512*/;
assign _1711_ = _1702_ & _1710_ /*3510*/;
assign _1669_ = _1702_ ^ _1710_ /*3511*/;
assign _1708_ = _1709_ | _1711_ /*3508*/;
assign _1713_ = ~Q[8] /*3507*/;
assign _1712_ = _1713_ & D[5] /*3506*/;
assign _1715_ = _1558_ & _1712_ /*3501*/;
assign _1716_ = _1558_ ^ _1712_ /*3504*/;
assign _1717_ = _1708_ & _1716_ /*3502*/;
assign _1670_ = _1708_ ^ _1716_ /*3503*/;
assign _1714_ = _1715_ | _1717_ /*3500*/;
assign _1719_ = ~Q[8] /*3499*/;
assign _1718_ = _1719_ & D[6] /*3498*/;
assign _1721_ = _1559_ & _1718_ /*3493*/;
assign _1722_ = _1559_ ^ _1718_ /*3496*/;
assign _1723_ = _1714_ & _1722_ /*3494*/;
assign _1671_ = _1714_ ^ _1722_ /*3495*/;
assign _1720_ = _1721_ | _1723_ /*3492*/;
assign _1725_ = ~Q[8] /*3491*/;
assign _1724_ = _1725_ & D[7] /*3490*/;
assign _1727_ = _1560_ & _1724_ /*3485*/;
assign _1728_ = _1560_ ^ _1724_ /*3488*/;
assign _1729_ = _1720_ & _1728_ /*3486*/;
assign _1672_ = _1720_ ^ _1728_ /*3487*/;
assign _1726_ = _1727_ | _1729_ /*3484*/;
assign _1731_ = ~Q[8] /*3483*/;
assign _1730_ = _1731_ & D[8] /*3482*/;
assign _1733_ = _1561_ & _1730_ /*3477*/;
assign _1734_ = _1561_ ^ _1730_ /*3480*/;
assign _1735_ = _1726_ & _1734_ /*3478*/;
assign _1673_ = _1726_ ^ _1734_ /*3479*/;
assign _1732_ = _1733_ | _1735_ /*3476*/;
assign _1737_ = ~Q[8] /*3475*/;
assign _1736_ = _1737_ & D[9] /*3474*/;
assign _1739_ = _1562_ & _1736_ /*3469*/;
assign _1740_ = _1562_ ^ _1736_ /*3472*/;
assign _1741_ = _1732_ & _1740_ /*3470*/;
assign _1674_ = _1732_ ^ _1740_ /*3471*/;
assign _1738_ = _1739_ | _1741_ /*3468*/;
assign _1743_ = ~Q[8] /*3467*/;
assign _1742_ = _1743_ & D[10] /*3466*/;
assign _1745_ = _1563_ & _1742_ /*3461*/;
assign _1746_ = _1563_ ^ _1742_ /*3464*/;
assign _1747_ = _1738_ & _1746_ /*3462*/;
assign _1675_ = _1738_ ^ _1746_ /*3463*/;
assign _1744_ = _1745_ | _1747_ /*3460*/;
assign _1749_ = ~Q[8] /*3459*/;
assign _1748_ = _1749_ & D[11] /*3458*/;
assign _1751_ = _1564_ & _1748_ /*3453*/;
assign _1752_ = _1564_ ^ _1748_ /*3456*/;
assign _1753_ = _1744_ & _1752_ /*3454*/;
assign _1676_ = _1744_ ^ _1752_ /*3455*/;
assign _1750_ = _1751_ | _1753_ /*3452*/;
assign _1755_ = ~Q[8] /*3451*/;
assign _1754_ = _1755_ & D[12] /*3450*/;
assign _1757_ = _1565_ & _1754_ /*3445*/;
assign _1758_ = _1565_ ^ _1754_ /*3448*/;
assign _1759_ = _1750_ & _1758_ /*3446*/;
assign _1677_ = _1750_ ^ _1758_ /*3447*/;
assign _1756_ = _1757_ | _1759_ /*3444*/;
assign _1761_ = ~Q[8] /*3443*/;
assign _1760_ = _1761_ & D[13] /*3442*/;
assign _1763_ = _1566_ & _1760_ /*3437*/;
assign _1764_ = _1566_ ^ _1760_ /*3440*/;
assign _1765_ = _1756_ & _1764_ /*3438*/;
assign _1678_ = _1756_ ^ _1764_ /*3439*/;
assign _1762_ = _1763_ | _1765_ /*3436*/;
assign _1767_ = ~Q[8] /*3435*/;
assign _1766_ = _1767_ & D[14] /*3434*/;
assign _1769_ = _1567_ & _1766_ /*3429*/;
assign _1770_ = _1567_ ^ _1766_ /*3432*/;
assign _1771_ = _1762_ & _1770_ /*3430*/;
assign _1679_ = _1762_ ^ _1770_ /*3431*/;
assign _1768_ = _1769_ | _1771_ /*3428*/;
assign _1773_ = ~Q[8] /*3427*/;
assign _1772_ = _1773_ & zeroWire /*3426*/;
assign _1774_ = _1568_ ^ _1772_ /*3424*/;
assign _1680_ = _1774_ ^ _1768_ /*3423*/;
assign _1797_ = ~D[0] /*3361*/;
assign _1794_ = R_0[7] & _1797_ /*3357*/;
assign _1795_ = R_0[7] ^ _1797_ /*3360*/;
assign _1796_ = oneWire & _1795_ /*3358*/;
assign _1777_ = oneWire ^ _1795_ /*3359*/;
assign _1793_ = _1794_ | _1796_ /*3356*/;
assign _1802_ = ~D[1] /*3355*/;
assign _1799_ = _1665_ & _1802_ /*3351*/;
assign _1800_ = _1665_ ^ _1802_ /*3354*/;
assign _1801_ = _1793_ & _1800_ /*3352*/;
assign _1778_ = _1793_ ^ _1800_ /*3353*/;
assign _1798_ = _1799_ | _1801_ /*3350*/;
assign _1807_ = ~D[2] /*3349*/;
assign _1804_ = _1666_ & _1807_ /*3345*/;
assign _1805_ = _1666_ ^ _1807_ /*3348*/;
assign _1806_ = _1798_ & _1805_ /*3346*/;
assign _1779_ = _1798_ ^ _1805_ /*3347*/;
assign _1803_ = _1804_ | _1806_ /*3344*/;
assign _1812_ = ~D[3] /*3343*/;
assign _1809_ = _1667_ & _1812_ /*3339*/;
assign _1810_ = _1667_ ^ _1812_ /*3342*/;
assign _1811_ = _1803_ & _1810_ /*3340*/;
assign _1780_ = _1803_ ^ _1810_ /*3341*/;
assign _1808_ = _1809_ | _1811_ /*3338*/;
assign _1817_ = ~D[4] /*3337*/;
assign _1814_ = _1668_ & _1817_ /*3333*/;
assign _1815_ = _1668_ ^ _1817_ /*3336*/;
assign _1816_ = _1808_ & _1815_ /*3334*/;
assign _1781_ = _1808_ ^ _1815_ /*3335*/;
assign _1813_ = _1814_ | _1816_ /*3332*/;
assign _1822_ = ~D[5] /*3331*/;
assign _1819_ = _1669_ & _1822_ /*3327*/;
assign _1820_ = _1669_ ^ _1822_ /*3330*/;
assign _1821_ = _1813_ & _1820_ /*3328*/;
assign _1782_ = _1813_ ^ _1820_ /*3329*/;
assign _1818_ = _1819_ | _1821_ /*3326*/;
assign _1827_ = ~D[6] /*3325*/;
assign _1824_ = _1670_ & _1827_ /*3321*/;
assign _1825_ = _1670_ ^ _1827_ /*3324*/;
assign _1826_ = _1818_ & _1825_ /*3322*/;
assign _1783_ = _1818_ ^ _1825_ /*3323*/;
assign _1823_ = _1824_ | _1826_ /*3320*/;
assign _1832_ = ~D[7] /*3319*/;
assign _1829_ = _1671_ & _1832_ /*3315*/;
assign _1830_ = _1671_ ^ _1832_ /*3318*/;
assign _1831_ = _1823_ & _1830_ /*3316*/;
assign _1784_ = _1823_ ^ _1830_ /*3317*/;
assign _1828_ = _1829_ | _1831_ /*3314*/;
assign _1837_ = ~D[8] /*3313*/;
assign _1834_ = _1672_ & _1837_ /*3309*/;
assign _1835_ = _1672_ ^ _1837_ /*3312*/;
assign _1836_ = _1828_ & _1835_ /*3310*/;
assign _1785_ = _1828_ ^ _1835_ /*3311*/;
assign _1833_ = _1834_ | _1836_ /*3308*/;
assign _1842_ = ~D[9] /*3307*/;
assign _1839_ = _1673_ & _1842_ /*3303*/;
assign _1840_ = _1673_ ^ _1842_ /*3306*/;
assign _1841_ = _1833_ & _1840_ /*3304*/;
assign _1786_ = _1833_ ^ _1840_ /*3305*/;
assign _1838_ = _1839_ | _1841_ /*3302*/;
assign _1847_ = ~D[10] /*3301*/;
assign _1844_ = _1674_ & _1847_ /*3297*/;
assign _1845_ = _1674_ ^ _1847_ /*3300*/;
assign _1846_ = _1838_ & _1845_ /*3298*/;
assign _1787_ = _1838_ ^ _1845_ /*3299*/;
assign _1843_ = _1844_ | _1846_ /*3296*/;
assign _1852_ = ~D[11] /*3295*/;
assign _1849_ = _1675_ & _1852_ /*3291*/;
assign _1850_ = _1675_ ^ _1852_ /*3294*/;
assign _1851_ = _1843_ & _1850_ /*3292*/;
assign _1788_ = _1843_ ^ _1850_ /*3293*/;
assign _1848_ = _1849_ | _1851_ /*3290*/;
assign _1857_ = ~D[12] /*3289*/;
assign _1854_ = _1676_ & _1857_ /*3285*/;
assign _1855_ = _1676_ ^ _1857_ /*3288*/;
assign _1856_ = _1848_ & _1855_ /*3286*/;
assign _1789_ = _1848_ ^ _1855_ /*3287*/;
assign _1853_ = _1854_ | _1856_ /*3284*/;
assign _1862_ = ~D[13] /*3283*/;
assign _1859_ = _1677_ & _1862_ /*3279*/;
assign _1860_ = _1677_ ^ _1862_ /*3282*/;
assign _1861_ = _1853_ & _1860_ /*3280*/;
assign _1790_ = _1853_ ^ _1860_ /*3281*/;
assign _1858_ = _1859_ | _1861_ /*3278*/;
assign _1867_ = ~D[14] /*3277*/;
assign _1864_ = _1678_ & _1867_ /*3273*/;
assign _1865_ = _1678_ ^ _1867_ /*3276*/;
assign _1866_ = _1858_ & _1865_ /*3274*/;
assign _1791_ = _1858_ ^ _1865_ /*3275*/;
assign _1863_ = _1864_ | _1866_ /*3272*/;
assign _1868_ = _1679_ & oneWire /*3267*/;
assign _1869_ = _1679_ ^ oneWire /*3270*/;
assign _1870_ = _1863_ & _1869_ /*3268*/;
assign _1792_ = _1863_ ^ _1869_ /*3269*/;
assign Q[7] = _1868_ | _1870_ /*3266*/;
assign _1907_ = ~Q[7] /*3169*/;
assign _1906_ = _1907_ & D[0] /*3168*/;
assign _1909_ = _1777_ & _1906_ /*3163*/;
assign _1910_ = _1777_ ^ _1906_ /*3166*/;
assign _1911_ = zeroWire & _1910_ /*3164*/;
assign _1889_ = zeroWire ^ _1910_ /*3165*/;
assign _1908_ = _1909_ | _1911_ /*3162*/;
assign _1913_ = ~Q[7] /*3161*/;
assign _1912_ = _1913_ & D[1] /*3160*/;
assign _1915_ = _1778_ & _1912_ /*3155*/;
assign _1916_ = _1778_ ^ _1912_ /*3158*/;
assign _1917_ = _1908_ & _1916_ /*3156*/;
assign _1890_ = _1908_ ^ _1916_ /*3157*/;
assign _1914_ = _1915_ | _1917_ /*3154*/;
assign _1919_ = ~Q[7] /*3153*/;
assign _1918_ = _1919_ & D[2] /*3152*/;
assign _1921_ = _1779_ & _1918_ /*3147*/;
assign _1922_ = _1779_ ^ _1918_ /*3150*/;
assign _1923_ = _1914_ & _1922_ /*3148*/;
assign _1891_ = _1914_ ^ _1922_ /*3149*/;
assign _1920_ = _1921_ | _1923_ /*3146*/;
assign _1925_ = ~Q[7] /*3145*/;
assign _1924_ = _1925_ & D[3] /*3144*/;
assign _1927_ = _1780_ & _1924_ /*3139*/;
assign _1928_ = _1780_ ^ _1924_ /*3142*/;
assign _1929_ = _1920_ & _1928_ /*3140*/;
assign _1892_ = _1920_ ^ _1928_ /*3141*/;
assign _1926_ = _1927_ | _1929_ /*3138*/;
assign _1931_ = ~Q[7] /*3137*/;
assign _1930_ = _1931_ & D[4] /*3136*/;
assign _1933_ = _1781_ & _1930_ /*3131*/;
assign _1934_ = _1781_ ^ _1930_ /*3134*/;
assign _1935_ = _1926_ & _1934_ /*3132*/;
assign _1893_ = _1926_ ^ _1934_ /*3133*/;
assign _1932_ = _1933_ | _1935_ /*3130*/;
assign _1937_ = ~Q[7] /*3129*/;
assign _1936_ = _1937_ & D[5] /*3128*/;
assign _1939_ = _1782_ & _1936_ /*3123*/;
assign _1940_ = _1782_ ^ _1936_ /*3126*/;
assign _1941_ = _1932_ & _1940_ /*3124*/;
assign _1894_ = _1932_ ^ _1940_ /*3125*/;
assign _1938_ = _1939_ | _1941_ /*3122*/;
assign _1943_ = ~Q[7] /*3121*/;
assign _1942_ = _1943_ & D[6] /*3120*/;
assign _1945_ = _1783_ & _1942_ /*3115*/;
assign _1946_ = _1783_ ^ _1942_ /*3118*/;
assign _1947_ = _1938_ & _1946_ /*3116*/;
assign _1895_ = _1938_ ^ _1946_ /*3117*/;
assign _1944_ = _1945_ | _1947_ /*3114*/;
assign _1949_ = ~Q[7] /*3113*/;
assign _1948_ = _1949_ & D[7] /*3112*/;
assign _1951_ = _1784_ & _1948_ /*3107*/;
assign _1952_ = _1784_ ^ _1948_ /*3110*/;
assign _1953_ = _1944_ & _1952_ /*3108*/;
assign _1896_ = _1944_ ^ _1952_ /*3109*/;
assign _1950_ = _1951_ | _1953_ /*3106*/;
assign _1955_ = ~Q[7] /*3105*/;
assign _1954_ = _1955_ & D[8] /*3104*/;
assign _1957_ = _1785_ & _1954_ /*3099*/;
assign _1958_ = _1785_ ^ _1954_ /*3102*/;
assign _1959_ = _1950_ & _1958_ /*3100*/;
assign _1897_ = _1950_ ^ _1958_ /*3101*/;
assign _1956_ = _1957_ | _1959_ /*3098*/;
assign _1961_ = ~Q[7] /*3097*/;
assign _1960_ = _1961_ & D[9] /*3096*/;
assign _1963_ = _1786_ & _1960_ /*3091*/;
assign _1964_ = _1786_ ^ _1960_ /*3094*/;
assign _1965_ = _1956_ & _1964_ /*3092*/;
assign _1898_ = _1956_ ^ _1964_ /*3093*/;
assign _1962_ = _1963_ | _1965_ /*3090*/;
assign _1967_ = ~Q[7] /*3089*/;
assign _1966_ = _1967_ & D[10] /*3088*/;
assign _1969_ = _1787_ & _1966_ /*3083*/;
assign _1970_ = _1787_ ^ _1966_ /*3086*/;
assign _1971_ = _1962_ & _1970_ /*3084*/;
assign _1899_ = _1962_ ^ _1970_ /*3085*/;
assign _1968_ = _1969_ | _1971_ /*3082*/;
assign _1973_ = ~Q[7] /*3081*/;
assign _1972_ = _1973_ & D[11] /*3080*/;
assign _1975_ = _1788_ & _1972_ /*3075*/;
assign _1976_ = _1788_ ^ _1972_ /*3078*/;
assign _1977_ = _1968_ & _1976_ /*3076*/;
assign _1900_ = _1968_ ^ _1976_ /*3077*/;
assign _1974_ = _1975_ | _1977_ /*3074*/;
assign _1979_ = ~Q[7] /*3073*/;
assign _1978_ = _1979_ & D[12] /*3072*/;
assign _1981_ = _1789_ & _1978_ /*3067*/;
assign _1982_ = _1789_ ^ _1978_ /*3070*/;
assign _1983_ = _1974_ & _1982_ /*3068*/;
assign _1901_ = _1974_ ^ _1982_ /*3069*/;
assign _1980_ = _1981_ | _1983_ /*3066*/;
assign _1985_ = ~Q[7] /*3065*/;
assign _1984_ = _1985_ & D[13] /*3064*/;
assign _1987_ = _1790_ & _1984_ /*3059*/;
assign _1988_ = _1790_ ^ _1984_ /*3062*/;
assign _1989_ = _1980_ & _1988_ /*3060*/;
assign _1902_ = _1980_ ^ _1988_ /*3061*/;
assign _1986_ = _1987_ | _1989_ /*3058*/;
assign _1991_ = ~Q[7] /*3057*/;
assign _1990_ = _1991_ & D[14] /*3056*/;
assign _1993_ = _1791_ & _1990_ /*3051*/;
assign _1994_ = _1791_ ^ _1990_ /*3054*/;
assign _1995_ = _1986_ & _1994_ /*3052*/;
assign _1903_ = _1986_ ^ _1994_ /*3053*/;
assign _1992_ = _1993_ | _1995_ /*3050*/;
assign _1997_ = ~Q[7] /*3049*/;
assign _1996_ = _1997_ & zeroWire /*3048*/;
assign _1998_ = _1792_ ^ _1996_ /*3046*/;
assign _1904_ = _1998_ ^ _1992_ /*3045*/;
assign _2021_ = ~D[0] /*2983*/;
assign _2018_ = R_0[6] & _2021_ /*2979*/;
assign _2019_ = R_0[6] ^ _2021_ /*2982*/;
assign _2020_ = oneWire & _2019_ /*2980*/;
assign _2001_ = oneWire ^ _2019_ /*2981*/;
assign _2017_ = _2018_ | _2020_ /*2978*/;
assign _2026_ = ~D[1] /*2977*/;
assign _2023_ = _1889_ & _2026_ /*2973*/;
assign _2024_ = _1889_ ^ _2026_ /*2976*/;
assign _2025_ = _2017_ & _2024_ /*2974*/;
assign _2002_ = _2017_ ^ _2024_ /*2975*/;
assign _2022_ = _2023_ | _2025_ /*2972*/;
assign _2031_ = ~D[2] /*2971*/;
assign _2028_ = _1890_ & _2031_ /*2967*/;
assign _2029_ = _1890_ ^ _2031_ /*2970*/;
assign _2030_ = _2022_ & _2029_ /*2968*/;
assign _2003_ = _2022_ ^ _2029_ /*2969*/;
assign _2027_ = _2028_ | _2030_ /*2966*/;
assign _2036_ = ~D[3] /*2965*/;
assign _2033_ = _1891_ & _2036_ /*2961*/;
assign _2034_ = _1891_ ^ _2036_ /*2964*/;
assign _2035_ = _2027_ & _2034_ /*2962*/;
assign _2004_ = _2027_ ^ _2034_ /*2963*/;
assign _2032_ = _2033_ | _2035_ /*2960*/;
assign _2041_ = ~D[4] /*2959*/;
assign _2038_ = _1892_ & _2041_ /*2955*/;
assign _2039_ = _1892_ ^ _2041_ /*2958*/;
assign _2040_ = _2032_ & _2039_ /*2956*/;
assign _2005_ = _2032_ ^ _2039_ /*2957*/;
assign _2037_ = _2038_ | _2040_ /*2954*/;
assign _2046_ = ~D[5] /*2953*/;
assign _2043_ = _1893_ & _2046_ /*2949*/;
assign _2044_ = _1893_ ^ _2046_ /*2952*/;
assign _2045_ = _2037_ & _2044_ /*2950*/;
assign _2006_ = _2037_ ^ _2044_ /*2951*/;
assign _2042_ = _2043_ | _2045_ /*2948*/;
assign _2051_ = ~D[6] /*2947*/;
assign _2048_ = _1894_ & _2051_ /*2943*/;
assign _2049_ = _1894_ ^ _2051_ /*2946*/;
assign _2050_ = _2042_ & _2049_ /*2944*/;
assign _2007_ = _2042_ ^ _2049_ /*2945*/;
assign _2047_ = _2048_ | _2050_ /*2942*/;
assign _2056_ = ~D[7] /*2941*/;
assign _2053_ = _1895_ & _2056_ /*2937*/;
assign _2054_ = _1895_ ^ _2056_ /*2940*/;
assign _2055_ = _2047_ & _2054_ /*2938*/;
assign _2008_ = _2047_ ^ _2054_ /*2939*/;
assign _2052_ = _2053_ | _2055_ /*2936*/;
assign _2061_ = ~D[8] /*2935*/;
assign _2058_ = _1896_ & _2061_ /*2931*/;
assign _2059_ = _1896_ ^ _2061_ /*2934*/;
assign _2060_ = _2052_ & _2059_ /*2932*/;
assign _2009_ = _2052_ ^ _2059_ /*2933*/;
assign _2057_ = _2058_ | _2060_ /*2930*/;
assign _2066_ = ~D[9] /*2929*/;
assign _2063_ = _1897_ & _2066_ /*2925*/;
assign _2064_ = _1897_ ^ _2066_ /*2928*/;
assign _2065_ = _2057_ & _2064_ /*2926*/;
assign _2010_ = _2057_ ^ _2064_ /*2927*/;
assign _2062_ = _2063_ | _2065_ /*2924*/;
assign _2071_ = ~D[10] /*2923*/;
assign _2068_ = _1898_ & _2071_ /*2919*/;
assign _2069_ = _1898_ ^ _2071_ /*2922*/;
assign _2070_ = _2062_ & _2069_ /*2920*/;
assign _2011_ = _2062_ ^ _2069_ /*2921*/;
assign _2067_ = _2068_ | _2070_ /*2918*/;
assign _2076_ = ~D[11] /*2917*/;
assign _2073_ = _1899_ & _2076_ /*2913*/;
assign _2074_ = _1899_ ^ _2076_ /*2916*/;
assign _2075_ = _2067_ & _2074_ /*2914*/;
assign _2012_ = _2067_ ^ _2074_ /*2915*/;
assign _2072_ = _2073_ | _2075_ /*2912*/;
assign _2081_ = ~D[12] /*2911*/;
assign _2078_ = _1900_ & _2081_ /*2907*/;
assign _2079_ = _1900_ ^ _2081_ /*2910*/;
assign _2080_ = _2072_ & _2079_ /*2908*/;
assign _2013_ = _2072_ ^ _2079_ /*2909*/;
assign _2077_ = _2078_ | _2080_ /*2906*/;
assign _2086_ = ~D[13] /*2905*/;
assign _2083_ = _1901_ & _2086_ /*2901*/;
assign _2084_ = _1901_ ^ _2086_ /*2904*/;
assign _2085_ = _2077_ & _2084_ /*2902*/;
assign _2014_ = _2077_ ^ _2084_ /*2903*/;
assign _2082_ = _2083_ | _2085_ /*2900*/;
assign _2091_ = ~D[14] /*2899*/;
assign _2088_ = _1902_ & _2091_ /*2895*/;
assign _2089_ = _1902_ ^ _2091_ /*2898*/;
assign _2090_ = _2082_ & _2089_ /*2896*/;
assign _2015_ = _2082_ ^ _2089_ /*2897*/;
assign _2087_ = _2088_ | _2090_ /*2894*/;
assign _2092_ = _1903_ & oneWire /*2889*/;
assign _2093_ = _1903_ ^ oneWire /*2892*/;
assign _2094_ = _2087_ & _2093_ /*2890*/;
assign _2016_ = _2087_ ^ _2093_ /*2891*/;
assign Q[6] = _2092_ | _2094_ /*2888*/;
assign _2131_ = ~Q[6] /*2791*/;
assign _2130_ = _2131_ & D[0] /*2790*/;
assign _2133_ = _2001_ & _2130_ /*2785*/;
assign _2134_ = _2001_ ^ _2130_ /*2788*/;
assign _2135_ = zeroWire & _2134_ /*2786*/;
assign _2113_ = zeroWire ^ _2134_ /*2787*/;
assign _2132_ = _2133_ | _2135_ /*2784*/;
assign _2137_ = ~Q[6] /*2783*/;
assign _2136_ = _2137_ & D[1] /*2782*/;
assign _2139_ = _2002_ & _2136_ /*2777*/;
assign _2140_ = _2002_ ^ _2136_ /*2780*/;
assign _2141_ = _2132_ & _2140_ /*2778*/;
assign _2114_ = _2132_ ^ _2140_ /*2779*/;
assign _2138_ = _2139_ | _2141_ /*2776*/;
assign _2143_ = ~Q[6] /*2775*/;
assign _2142_ = _2143_ & D[2] /*2774*/;
assign _2145_ = _2003_ & _2142_ /*2769*/;
assign _2146_ = _2003_ ^ _2142_ /*2772*/;
assign _2147_ = _2138_ & _2146_ /*2770*/;
assign _2115_ = _2138_ ^ _2146_ /*2771*/;
assign _2144_ = _2145_ | _2147_ /*2768*/;
assign _2149_ = ~Q[6] /*2767*/;
assign _2148_ = _2149_ & D[3] /*2766*/;
assign _2151_ = _2004_ & _2148_ /*2761*/;
assign _2152_ = _2004_ ^ _2148_ /*2764*/;
assign _2153_ = _2144_ & _2152_ /*2762*/;
assign _2116_ = _2144_ ^ _2152_ /*2763*/;
assign _2150_ = _2151_ | _2153_ /*2760*/;
assign _2155_ = ~Q[6] /*2759*/;
assign _2154_ = _2155_ & D[4] /*2758*/;
assign _2157_ = _2005_ & _2154_ /*2753*/;
assign _2158_ = _2005_ ^ _2154_ /*2756*/;
assign _2159_ = _2150_ & _2158_ /*2754*/;
assign _2117_ = _2150_ ^ _2158_ /*2755*/;
assign _2156_ = _2157_ | _2159_ /*2752*/;
assign _2161_ = ~Q[6] /*2751*/;
assign _2160_ = _2161_ & D[5] /*2750*/;
assign _2163_ = _2006_ & _2160_ /*2745*/;
assign _2164_ = _2006_ ^ _2160_ /*2748*/;
assign _2165_ = _2156_ & _2164_ /*2746*/;
assign _2118_ = _2156_ ^ _2164_ /*2747*/;
assign _2162_ = _2163_ | _2165_ /*2744*/;
assign _2167_ = ~Q[6] /*2743*/;
assign _2166_ = _2167_ & D[6] /*2742*/;
assign _2169_ = _2007_ & _2166_ /*2737*/;
assign _2170_ = _2007_ ^ _2166_ /*2740*/;
assign _2171_ = _2162_ & _2170_ /*2738*/;
assign _2119_ = _2162_ ^ _2170_ /*2739*/;
assign _2168_ = _2169_ | _2171_ /*2736*/;
assign _2173_ = ~Q[6] /*2735*/;
assign _2172_ = _2173_ & D[7] /*2734*/;
assign _2175_ = _2008_ & _2172_ /*2729*/;
assign _2176_ = _2008_ ^ _2172_ /*2732*/;
assign _2177_ = _2168_ & _2176_ /*2730*/;
assign _2120_ = _2168_ ^ _2176_ /*2731*/;
assign _2174_ = _2175_ | _2177_ /*2728*/;
assign _2179_ = ~Q[6] /*2727*/;
assign _2178_ = _2179_ & D[8] /*2726*/;
assign _2181_ = _2009_ & _2178_ /*2721*/;
assign _2182_ = _2009_ ^ _2178_ /*2724*/;
assign _2183_ = _2174_ & _2182_ /*2722*/;
assign _2121_ = _2174_ ^ _2182_ /*2723*/;
assign _2180_ = _2181_ | _2183_ /*2720*/;
assign _2185_ = ~Q[6] /*2719*/;
assign _2184_ = _2185_ & D[9] /*2718*/;
assign _2187_ = _2010_ & _2184_ /*2713*/;
assign _2188_ = _2010_ ^ _2184_ /*2716*/;
assign _2189_ = _2180_ & _2188_ /*2714*/;
assign _2122_ = _2180_ ^ _2188_ /*2715*/;
assign _2186_ = _2187_ | _2189_ /*2712*/;
assign _2191_ = ~Q[6] /*2711*/;
assign _2190_ = _2191_ & D[10] /*2710*/;
assign _2193_ = _2011_ & _2190_ /*2705*/;
assign _2194_ = _2011_ ^ _2190_ /*2708*/;
assign _2195_ = _2186_ & _2194_ /*2706*/;
assign _2123_ = _2186_ ^ _2194_ /*2707*/;
assign _2192_ = _2193_ | _2195_ /*2704*/;
assign _2197_ = ~Q[6] /*2703*/;
assign _2196_ = _2197_ & D[11] /*2702*/;
assign _2199_ = _2012_ & _2196_ /*2697*/;
assign _2200_ = _2012_ ^ _2196_ /*2700*/;
assign _2201_ = _2192_ & _2200_ /*2698*/;
assign _2124_ = _2192_ ^ _2200_ /*2699*/;
assign _2198_ = _2199_ | _2201_ /*2696*/;
assign _2203_ = ~Q[6] /*2695*/;
assign _2202_ = _2203_ & D[12] /*2694*/;
assign _2205_ = _2013_ & _2202_ /*2689*/;
assign _2206_ = _2013_ ^ _2202_ /*2692*/;
assign _2207_ = _2198_ & _2206_ /*2690*/;
assign _2125_ = _2198_ ^ _2206_ /*2691*/;
assign _2204_ = _2205_ | _2207_ /*2688*/;
assign _2209_ = ~Q[6] /*2687*/;
assign _2208_ = _2209_ & D[13] /*2686*/;
assign _2211_ = _2014_ & _2208_ /*2681*/;
assign _2212_ = _2014_ ^ _2208_ /*2684*/;
assign _2213_ = _2204_ & _2212_ /*2682*/;
assign _2126_ = _2204_ ^ _2212_ /*2683*/;
assign _2210_ = _2211_ | _2213_ /*2680*/;
assign _2215_ = ~Q[6] /*2679*/;
assign _2214_ = _2215_ & D[14] /*2678*/;
assign _2217_ = _2015_ & _2214_ /*2673*/;
assign _2218_ = _2015_ ^ _2214_ /*2676*/;
assign _2219_ = _2210_ & _2218_ /*2674*/;
assign _2127_ = _2210_ ^ _2218_ /*2675*/;
assign _2216_ = _2217_ | _2219_ /*2672*/;
assign _2221_ = ~Q[6] /*2671*/;
assign _2220_ = _2221_ & zeroWire /*2670*/;
assign _2222_ = _2016_ ^ _2220_ /*2668*/;
assign _2128_ = _2222_ ^ _2216_ /*2667*/;
assign _2245_ = ~D[0] /*2605*/;
assign _2242_ = R_0[5] & _2245_ /*2601*/;
assign _2243_ = R_0[5] ^ _2245_ /*2604*/;
assign _2244_ = oneWire & _2243_ /*2602*/;
assign _2225_ = oneWire ^ _2243_ /*2603*/;
assign _2241_ = _2242_ | _2244_ /*2600*/;
assign _2250_ = ~D[1] /*2599*/;
assign _2247_ = _2113_ & _2250_ /*2595*/;
assign _2248_ = _2113_ ^ _2250_ /*2598*/;
assign _2249_ = _2241_ & _2248_ /*2596*/;
assign _2226_ = _2241_ ^ _2248_ /*2597*/;
assign _2246_ = _2247_ | _2249_ /*2594*/;
assign _2255_ = ~D[2] /*2593*/;
assign _2252_ = _2114_ & _2255_ /*2589*/;
assign _2253_ = _2114_ ^ _2255_ /*2592*/;
assign _2254_ = _2246_ & _2253_ /*2590*/;
assign _2227_ = _2246_ ^ _2253_ /*2591*/;
assign _2251_ = _2252_ | _2254_ /*2588*/;
assign _2260_ = ~D[3] /*2587*/;
assign _2257_ = _2115_ & _2260_ /*2583*/;
assign _2258_ = _2115_ ^ _2260_ /*2586*/;
assign _2259_ = _2251_ & _2258_ /*2584*/;
assign _2228_ = _2251_ ^ _2258_ /*2585*/;
assign _2256_ = _2257_ | _2259_ /*2582*/;
assign _2265_ = ~D[4] /*2581*/;
assign _2262_ = _2116_ & _2265_ /*2577*/;
assign _2263_ = _2116_ ^ _2265_ /*2580*/;
assign _2264_ = _2256_ & _2263_ /*2578*/;
assign _2229_ = _2256_ ^ _2263_ /*2579*/;
assign _2261_ = _2262_ | _2264_ /*2576*/;
assign _2270_ = ~D[5] /*2575*/;
assign _2267_ = _2117_ & _2270_ /*2571*/;
assign _2268_ = _2117_ ^ _2270_ /*2574*/;
assign _2269_ = _2261_ & _2268_ /*2572*/;
assign _2230_ = _2261_ ^ _2268_ /*2573*/;
assign _2266_ = _2267_ | _2269_ /*2570*/;
assign _2275_ = ~D[6] /*2569*/;
assign _2272_ = _2118_ & _2275_ /*2565*/;
assign _2273_ = _2118_ ^ _2275_ /*2568*/;
assign _2274_ = _2266_ & _2273_ /*2566*/;
assign _2231_ = _2266_ ^ _2273_ /*2567*/;
assign _2271_ = _2272_ | _2274_ /*2564*/;
assign _2280_ = ~D[7] /*2563*/;
assign _2277_ = _2119_ & _2280_ /*2559*/;
assign _2278_ = _2119_ ^ _2280_ /*2562*/;
assign _2279_ = _2271_ & _2278_ /*2560*/;
assign _2232_ = _2271_ ^ _2278_ /*2561*/;
assign _2276_ = _2277_ | _2279_ /*2558*/;
assign _2285_ = ~D[8] /*2557*/;
assign _2282_ = _2120_ & _2285_ /*2553*/;
assign _2283_ = _2120_ ^ _2285_ /*2556*/;
assign _2284_ = _2276_ & _2283_ /*2554*/;
assign _2233_ = _2276_ ^ _2283_ /*2555*/;
assign _2281_ = _2282_ | _2284_ /*2552*/;
assign _2290_ = ~D[9] /*2551*/;
assign _2287_ = _2121_ & _2290_ /*2547*/;
assign _2288_ = _2121_ ^ _2290_ /*2550*/;
assign _2289_ = _2281_ & _2288_ /*2548*/;
assign _2234_ = _2281_ ^ _2288_ /*2549*/;
assign _2286_ = _2287_ | _2289_ /*2546*/;
assign _2295_ = ~D[10] /*2545*/;
assign _2292_ = _2122_ & _2295_ /*2541*/;
assign _2293_ = _2122_ ^ _2295_ /*2544*/;
assign _2294_ = _2286_ & _2293_ /*2542*/;
assign _2235_ = _2286_ ^ _2293_ /*2543*/;
assign _2291_ = _2292_ | _2294_ /*2540*/;
assign _2300_ = ~D[11] /*2539*/;
assign _2297_ = _2123_ & _2300_ /*2535*/;
assign _2298_ = _2123_ ^ _2300_ /*2538*/;
assign _2299_ = _2291_ & _2298_ /*2536*/;
assign _2236_ = _2291_ ^ _2298_ /*2537*/;
assign _2296_ = _2297_ | _2299_ /*2534*/;
assign _2305_ = ~D[12] /*2533*/;
assign _2302_ = _2124_ & _2305_ /*2529*/;
assign _2303_ = _2124_ ^ _2305_ /*2532*/;
assign _2304_ = _2296_ & _2303_ /*2530*/;
assign _2237_ = _2296_ ^ _2303_ /*2531*/;
assign _2301_ = _2302_ | _2304_ /*2528*/;
assign _2310_ = ~D[13] /*2527*/;
assign _2307_ = _2125_ & _2310_ /*2523*/;
assign _2308_ = _2125_ ^ _2310_ /*2526*/;
assign _2309_ = _2301_ & _2308_ /*2524*/;
assign _2238_ = _2301_ ^ _2308_ /*2525*/;
assign _2306_ = _2307_ | _2309_ /*2522*/;
assign _2315_ = ~D[14] /*2521*/;
assign _2312_ = _2126_ & _2315_ /*2517*/;
assign _2313_ = _2126_ ^ _2315_ /*2520*/;
assign _2314_ = _2306_ & _2313_ /*2518*/;
assign _2239_ = _2306_ ^ _2313_ /*2519*/;
assign _2311_ = _2312_ | _2314_ /*2516*/;
assign _2316_ = _2127_ & oneWire /*2511*/;
assign _2317_ = _2127_ ^ oneWire /*2514*/;
assign _2318_ = _2311_ & _2317_ /*2512*/;
assign _2240_ = _2311_ ^ _2317_ /*2513*/;
assign Q[5] = _2316_ | _2318_ /*2510*/;
assign _2355_ = ~Q[5] /*2413*/;
assign _2354_ = _2355_ & D[0] /*2412*/;
assign _2357_ = _2225_ & _2354_ /*2407*/;
assign _2358_ = _2225_ ^ _2354_ /*2410*/;
assign _2359_ = zeroWire & _2358_ /*2408*/;
assign _2337_ = zeroWire ^ _2358_ /*2409*/;
assign _2356_ = _2357_ | _2359_ /*2406*/;
assign _2361_ = ~Q[5] /*2405*/;
assign _2360_ = _2361_ & D[1] /*2404*/;
assign _2363_ = _2226_ & _2360_ /*2399*/;
assign _2364_ = _2226_ ^ _2360_ /*2402*/;
assign _2365_ = _2356_ & _2364_ /*2400*/;
assign _2338_ = _2356_ ^ _2364_ /*2401*/;
assign _2362_ = _2363_ | _2365_ /*2398*/;
assign _2367_ = ~Q[5] /*2397*/;
assign _2366_ = _2367_ & D[2] /*2396*/;
assign _2369_ = _2227_ & _2366_ /*2391*/;
assign _2370_ = _2227_ ^ _2366_ /*2394*/;
assign _2371_ = _2362_ & _2370_ /*2392*/;
assign _2339_ = _2362_ ^ _2370_ /*2393*/;
assign _2368_ = _2369_ | _2371_ /*2390*/;
assign _2373_ = ~Q[5] /*2389*/;
assign _2372_ = _2373_ & D[3] /*2388*/;
assign _2375_ = _2228_ & _2372_ /*2383*/;
assign _2376_ = _2228_ ^ _2372_ /*2386*/;
assign _2377_ = _2368_ & _2376_ /*2384*/;
assign _2340_ = _2368_ ^ _2376_ /*2385*/;
assign _2374_ = _2375_ | _2377_ /*2382*/;
assign _2379_ = ~Q[5] /*2381*/;
assign _2378_ = _2379_ & D[4] /*2380*/;
assign _2381_ = _2229_ & _2378_ /*2375*/;
assign _2382_ = _2229_ ^ _2378_ /*2378*/;
assign _2383_ = _2374_ & _2382_ /*2376*/;
assign _2341_ = _2374_ ^ _2382_ /*2377*/;
assign _2380_ = _2381_ | _2383_ /*2374*/;
assign _2385_ = ~Q[5] /*2373*/;
assign _2384_ = _2385_ & D[5] /*2372*/;
assign _2387_ = _2230_ & _2384_ /*2367*/;
assign _2388_ = _2230_ ^ _2384_ /*2370*/;
assign _2389_ = _2380_ & _2388_ /*2368*/;
assign _2342_ = _2380_ ^ _2388_ /*2369*/;
assign _2386_ = _2387_ | _2389_ /*2366*/;
assign _2391_ = ~Q[5] /*2365*/;
assign _2390_ = _2391_ & D[6] /*2364*/;
assign _2393_ = _2231_ & _2390_ /*2359*/;
assign _2394_ = _2231_ ^ _2390_ /*2362*/;
assign _2395_ = _2386_ & _2394_ /*2360*/;
assign _2343_ = _2386_ ^ _2394_ /*2361*/;
assign _2392_ = _2393_ | _2395_ /*2358*/;
assign _2397_ = ~Q[5] /*2357*/;
assign _2396_ = _2397_ & D[7] /*2356*/;
assign _2399_ = _2232_ & _2396_ /*2351*/;
assign _2400_ = _2232_ ^ _2396_ /*2354*/;
assign _2401_ = _2392_ & _2400_ /*2352*/;
assign _2344_ = _2392_ ^ _2400_ /*2353*/;
assign _2398_ = _2399_ | _2401_ /*2350*/;
assign _2403_ = ~Q[5] /*2349*/;
assign _2402_ = _2403_ & D[8] /*2348*/;
assign _2405_ = _2233_ & _2402_ /*2343*/;
assign _2406_ = _2233_ ^ _2402_ /*2346*/;
assign _2407_ = _2398_ & _2406_ /*2344*/;
assign _2345_ = _2398_ ^ _2406_ /*2345*/;
assign _2404_ = _2405_ | _2407_ /*2342*/;
assign _2409_ = ~Q[5] /*2341*/;
assign _2408_ = _2409_ & D[9] /*2340*/;
assign _2411_ = _2234_ & _2408_ /*2335*/;
assign _2412_ = _2234_ ^ _2408_ /*2338*/;
assign _2413_ = _2404_ & _2412_ /*2336*/;
assign _2346_ = _2404_ ^ _2412_ /*2337*/;
assign _2410_ = _2411_ | _2413_ /*2334*/;
assign _2415_ = ~Q[5] /*2333*/;
assign _2414_ = _2415_ & D[10] /*2332*/;
assign _2417_ = _2235_ & _2414_ /*2327*/;
assign _2418_ = _2235_ ^ _2414_ /*2330*/;
assign _2419_ = _2410_ & _2418_ /*2328*/;
assign _2347_ = _2410_ ^ _2418_ /*2329*/;
assign _2416_ = _2417_ | _2419_ /*2326*/;
assign _2421_ = ~Q[5] /*2325*/;
assign _2420_ = _2421_ & D[11] /*2324*/;
assign _2423_ = _2236_ & _2420_ /*2319*/;
assign _2424_ = _2236_ ^ _2420_ /*2322*/;
assign _2425_ = _2416_ & _2424_ /*2320*/;
assign _2348_ = _2416_ ^ _2424_ /*2321*/;
assign _2422_ = _2423_ | _2425_ /*2318*/;
assign _2427_ = ~Q[5] /*2317*/;
assign _2426_ = _2427_ & D[12] /*2316*/;
assign _2429_ = _2237_ & _2426_ /*2311*/;
assign _2430_ = _2237_ ^ _2426_ /*2314*/;
assign _2431_ = _2422_ & _2430_ /*2312*/;
assign _2349_ = _2422_ ^ _2430_ /*2313*/;
assign _2428_ = _2429_ | _2431_ /*2310*/;
assign _2433_ = ~Q[5] /*2309*/;
assign _2432_ = _2433_ & D[13] /*2308*/;
assign _2435_ = _2238_ & _2432_ /*2303*/;
assign _2436_ = _2238_ ^ _2432_ /*2306*/;
assign _2437_ = _2428_ & _2436_ /*2304*/;
assign _2350_ = _2428_ ^ _2436_ /*2305*/;
assign _2434_ = _2435_ | _2437_ /*2302*/;
assign _2439_ = ~Q[5] /*2301*/;
assign _2438_ = _2439_ & D[14] /*2300*/;
assign _2441_ = _2239_ & _2438_ /*2295*/;
assign _2442_ = _2239_ ^ _2438_ /*2298*/;
assign _2443_ = _2434_ & _2442_ /*2296*/;
assign _2351_ = _2434_ ^ _2442_ /*2297*/;
assign _2440_ = _2441_ | _2443_ /*2294*/;
assign _2445_ = ~Q[5] /*2293*/;
assign _2444_ = _2445_ & zeroWire /*2292*/;
assign _2446_ = _2240_ ^ _2444_ /*2290*/;
assign _2352_ = _2446_ ^ _2440_ /*2289*/;
assign _2469_ = ~D[0] /*2227*/;
assign _2466_ = R_0[4] & _2469_ /*2223*/;
assign _2467_ = R_0[4] ^ _2469_ /*2226*/;
assign _2468_ = oneWire & _2467_ /*2224*/;
assign _2449_ = oneWire ^ _2467_ /*2225*/;
assign _2465_ = _2466_ | _2468_ /*2222*/;
assign _2474_ = ~D[1] /*2221*/;
assign _2471_ = _2337_ & _2474_ /*2217*/;
assign _2472_ = _2337_ ^ _2474_ /*2220*/;
assign _2473_ = _2465_ & _2472_ /*2218*/;
assign _2450_ = _2465_ ^ _2472_ /*2219*/;
assign _2470_ = _2471_ | _2473_ /*2216*/;
assign _2479_ = ~D[2] /*2215*/;
assign _2476_ = _2338_ & _2479_ /*2211*/;
assign _2477_ = _2338_ ^ _2479_ /*2214*/;
assign _2478_ = _2470_ & _2477_ /*2212*/;
assign _2451_ = _2470_ ^ _2477_ /*2213*/;
assign _2475_ = _2476_ | _2478_ /*2210*/;
assign _2484_ = ~D[3] /*2209*/;
assign _2481_ = _2339_ & _2484_ /*2205*/;
assign _2482_ = _2339_ ^ _2484_ /*2208*/;
assign _2483_ = _2475_ & _2482_ /*2206*/;
assign _2452_ = _2475_ ^ _2482_ /*2207*/;
assign _2480_ = _2481_ | _2483_ /*2204*/;
assign _2489_ = ~D[4] /*2203*/;
assign _2486_ = _2340_ & _2489_ /*2199*/;
assign _2487_ = _2340_ ^ _2489_ /*2202*/;
assign _2488_ = _2480_ & _2487_ /*2200*/;
assign _2453_ = _2480_ ^ _2487_ /*2201*/;
assign _2485_ = _2486_ | _2488_ /*2198*/;
assign _2494_ = ~D[5] /*2197*/;
assign _2491_ = _2341_ & _2494_ /*2193*/;
assign _2492_ = _2341_ ^ _2494_ /*2196*/;
assign _2493_ = _2485_ & _2492_ /*2194*/;
assign _2454_ = _2485_ ^ _2492_ /*2195*/;
assign _2490_ = _2491_ | _2493_ /*2192*/;
assign _2499_ = ~D[6] /*2191*/;
assign _2496_ = _2342_ & _2499_ /*2187*/;
assign _2497_ = _2342_ ^ _2499_ /*2190*/;
assign _2498_ = _2490_ & _2497_ /*2188*/;
assign _2455_ = _2490_ ^ _2497_ /*2189*/;
assign _2495_ = _2496_ | _2498_ /*2186*/;
assign _2504_ = ~D[7] /*2185*/;
assign _2501_ = _2343_ & _2504_ /*2181*/;
assign _2502_ = _2343_ ^ _2504_ /*2184*/;
assign _2503_ = _2495_ & _2502_ /*2182*/;
assign _2456_ = _2495_ ^ _2502_ /*2183*/;
assign _2500_ = _2501_ | _2503_ /*2180*/;
assign _2509_ = ~D[8] /*2179*/;
assign _2506_ = _2344_ & _2509_ /*2175*/;
assign _2507_ = _2344_ ^ _2509_ /*2178*/;
assign _2508_ = _2500_ & _2507_ /*2176*/;
assign _2457_ = _2500_ ^ _2507_ /*2177*/;
assign _2505_ = _2506_ | _2508_ /*2174*/;
assign _2514_ = ~D[9] /*2173*/;
assign _2511_ = _2345_ & _2514_ /*2169*/;
assign _2512_ = _2345_ ^ _2514_ /*2172*/;
assign _2513_ = _2505_ & _2512_ /*2170*/;
assign _2458_ = _2505_ ^ _2512_ /*2171*/;
assign _2510_ = _2511_ | _2513_ /*2168*/;
assign _2519_ = ~D[10] /*2167*/;
assign _2516_ = _2346_ & _2519_ /*2163*/;
assign _2517_ = _2346_ ^ _2519_ /*2166*/;
assign _2518_ = _2510_ & _2517_ /*2164*/;
assign _2459_ = _2510_ ^ _2517_ /*2165*/;
assign _2515_ = _2516_ | _2518_ /*2162*/;
assign _2524_ = ~D[11] /*2161*/;
assign _2521_ = _2347_ & _2524_ /*2157*/;
assign _2522_ = _2347_ ^ _2524_ /*2160*/;
assign _2523_ = _2515_ & _2522_ /*2158*/;
assign _2460_ = _2515_ ^ _2522_ /*2159*/;
assign _2520_ = _2521_ | _2523_ /*2156*/;
assign _2529_ = ~D[12] /*2155*/;
assign _2526_ = _2348_ & _2529_ /*2151*/;
assign _2527_ = _2348_ ^ _2529_ /*2154*/;
assign _2528_ = _2520_ & _2527_ /*2152*/;
assign _2461_ = _2520_ ^ _2527_ /*2153*/;
assign _2525_ = _2526_ | _2528_ /*2150*/;
assign _2534_ = ~D[13] /*2149*/;
assign _2531_ = _2349_ & _2534_ /*2145*/;
assign _2532_ = _2349_ ^ _2534_ /*2148*/;
assign _2533_ = _2525_ & _2532_ /*2146*/;
assign _2462_ = _2525_ ^ _2532_ /*2147*/;
assign _2530_ = _2531_ | _2533_ /*2144*/;
assign _2539_ = ~D[14] /*2143*/;
assign _2536_ = _2350_ & _2539_ /*2139*/;
assign _2537_ = _2350_ ^ _2539_ /*2142*/;
assign _2538_ = _2530_ & _2537_ /*2140*/;
assign _2463_ = _2530_ ^ _2537_ /*2141*/;
assign _2535_ = _2536_ | _2538_ /*2138*/;
assign _2540_ = _2351_ & oneWire /*2133*/;
assign _2541_ = _2351_ ^ oneWire /*2136*/;
assign _2542_ = _2535_ & _2541_ /*2134*/;
assign _2464_ = _2535_ ^ _2541_ /*2135*/;
assign Q[4] = _2540_ | _2542_ /*2132*/;
assign _2579_ = ~Q[4] /*2035*/;
assign _2578_ = _2579_ & D[0] /*2034*/;
assign _2581_ = _2449_ & _2578_ /*2029*/;
assign _2582_ = _2449_ ^ _2578_ /*2032*/;
assign _2583_ = zeroWire & _2582_ /*2030*/;
assign _2561_ = zeroWire ^ _2582_ /*2031*/;
assign _2580_ = _2581_ | _2583_ /*2028*/;
assign _2585_ = ~Q[4] /*2027*/;
assign _2584_ = _2585_ & D[1] /*2026*/;
assign _2587_ = _2450_ & _2584_ /*2021*/;
assign _2588_ = _2450_ ^ _2584_ /*2024*/;
assign _2589_ = _2580_ & _2588_ /*2022*/;
assign _2562_ = _2580_ ^ _2588_ /*2023*/;
assign _2586_ = _2587_ | _2589_ /*2020*/;
assign _2591_ = ~Q[4] /*2019*/;
assign _2590_ = _2591_ & D[2] /*2018*/;
assign _2593_ = _2451_ & _2590_ /*2013*/;
assign _2594_ = _2451_ ^ _2590_ /*2016*/;
assign _2595_ = _2586_ & _2594_ /*2014*/;
assign _2563_ = _2586_ ^ _2594_ /*2015*/;
assign _2592_ = _2593_ | _2595_ /*2012*/;
assign _2597_ = ~Q[4] /*2011*/;
assign _2596_ = _2597_ & D[3] /*2010*/;
assign _2599_ = _2452_ & _2596_ /*2005*/;
assign _2600_ = _2452_ ^ _2596_ /*2008*/;
assign _2601_ = _2592_ & _2600_ /*2006*/;
assign _2564_ = _2592_ ^ _2600_ /*2007*/;
assign _2598_ = _2599_ | _2601_ /*2004*/;
assign _2603_ = ~Q[4] /*2003*/;
assign _2602_ = _2603_ & D[4] /*2002*/;
assign _2605_ = _2453_ & _2602_ /*1997*/;
assign _2606_ = _2453_ ^ _2602_ /*2000*/;
assign _2607_ = _2598_ & _2606_ /*1998*/;
assign _2565_ = _2598_ ^ _2606_ /*1999*/;
assign _2604_ = _2605_ | _2607_ /*1996*/;
assign _2609_ = ~Q[4] /*1995*/;
assign _2608_ = _2609_ & D[5] /*1994*/;
assign _2611_ = _2454_ & _2608_ /*1989*/;
assign _2612_ = _2454_ ^ _2608_ /*1992*/;
assign _2613_ = _2604_ & _2612_ /*1990*/;
assign _2566_ = _2604_ ^ _2612_ /*1991*/;
assign _2610_ = _2611_ | _2613_ /*1988*/;
assign _2615_ = ~Q[4] /*1987*/;
assign _2614_ = _2615_ & D[6] /*1986*/;
assign _2617_ = _2455_ & _2614_ /*1981*/;
assign _2618_ = _2455_ ^ _2614_ /*1984*/;
assign _2619_ = _2610_ & _2618_ /*1982*/;
assign _2567_ = _2610_ ^ _2618_ /*1983*/;
assign _2616_ = _2617_ | _2619_ /*1980*/;
assign _2621_ = ~Q[4] /*1979*/;
assign _2620_ = _2621_ & D[7] /*1978*/;
assign _2623_ = _2456_ & _2620_ /*1973*/;
assign _2624_ = _2456_ ^ _2620_ /*1976*/;
assign _2625_ = _2616_ & _2624_ /*1974*/;
assign _2568_ = _2616_ ^ _2624_ /*1975*/;
assign _2622_ = _2623_ | _2625_ /*1972*/;
assign _2627_ = ~Q[4] /*1971*/;
assign _2626_ = _2627_ & D[8] /*1970*/;
assign _2629_ = _2457_ & _2626_ /*1965*/;
assign _2630_ = _2457_ ^ _2626_ /*1968*/;
assign _2631_ = _2622_ & _2630_ /*1966*/;
assign _2569_ = _2622_ ^ _2630_ /*1967*/;
assign _2628_ = _2629_ | _2631_ /*1964*/;
assign _2633_ = ~Q[4] /*1963*/;
assign _2632_ = _2633_ & D[9] /*1962*/;
assign _2635_ = _2458_ & _2632_ /*1957*/;
assign _2636_ = _2458_ ^ _2632_ /*1960*/;
assign _2637_ = _2628_ & _2636_ /*1958*/;
assign _2570_ = _2628_ ^ _2636_ /*1959*/;
assign _2634_ = _2635_ | _2637_ /*1956*/;
assign _2639_ = ~Q[4] /*1955*/;
assign _2638_ = _2639_ & D[10] /*1954*/;
assign _2641_ = _2459_ & _2638_ /*1949*/;
assign _2642_ = _2459_ ^ _2638_ /*1952*/;
assign _2643_ = _2634_ & _2642_ /*1950*/;
assign _2571_ = _2634_ ^ _2642_ /*1951*/;
assign _2640_ = _2641_ | _2643_ /*1948*/;
assign _2645_ = ~Q[4] /*1947*/;
assign _2644_ = _2645_ & D[11] /*1946*/;
assign _2647_ = _2460_ & _2644_ /*1941*/;
assign _2648_ = _2460_ ^ _2644_ /*1944*/;
assign _2649_ = _2640_ & _2648_ /*1942*/;
assign _2572_ = _2640_ ^ _2648_ /*1943*/;
assign _2646_ = _2647_ | _2649_ /*1940*/;
assign _2651_ = ~Q[4] /*1939*/;
assign _2650_ = _2651_ & D[12] /*1938*/;
assign _2653_ = _2461_ & _2650_ /*1933*/;
assign _2654_ = _2461_ ^ _2650_ /*1936*/;
assign _2655_ = _2646_ & _2654_ /*1934*/;
assign _2573_ = _2646_ ^ _2654_ /*1935*/;
assign _2652_ = _2653_ | _2655_ /*1932*/;
assign _2657_ = ~Q[4] /*1931*/;
assign _2656_ = _2657_ & D[13] /*1930*/;
assign _2659_ = _2462_ & _2656_ /*1925*/;
assign _2660_ = _2462_ ^ _2656_ /*1928*/;
assign _2661_ = _2652_ & _2660_ /*1926*/;
assign _2574_ = _2652_ ^ _2660_ /*1927*/;
assign _2658_ = _2659_ | _2661_ /*1924*/;
assign _2663_ = ~Q[4] /*1923*/;
assign _2662_ = _2663_ & D[14] /*1922*/;
assign _2665_ = _2463_ & _2662_ /*1917*/;
assign _2666_ = _2463_ ^ _2662_ /*1920*/;
assign _2667_ = _2658_ & _2666_ /*1918*/;
assign _2575_ = _2658_ ^ _2666_ /*1919*/;
assign _2664_ = _2665_ | _2667_ /*1916*/;
assign _2669_ = ~Q[4] /*1915*/;
assign _2668_ = _2669_ & zeroWire /*1914*/;
assign _2670_ = _2464_ ^ _2668_ /*1912*/;
assign _2576_ = _2670_ ^ _2664_ /*1911*/;
assign _2693_ = ~D[0] /*1849*/;
assign _2690_ = R_0[3] & _2693_ /*1845*/;
assign _2691_ = R_0[3] ^ _2693_ /*1848*/;
assign _2692_ = oneWire & _2691_ /*1846*/;
assign _2673_ = oneWire ^ _2691_ /*1847*/;
assign _2689_ = _2690_ | _2692_ /*1844*/;
assign _2698_ = ~D[1] /*1843*/;
assign _2695_ = _2561_ & _2698_ /*1839*/;
assign _2696_ = _2561_ ^ _2698_ /*1842*/;
assign _2697_ = _2689_ & _2696_ /*1840*/;
assign _2674_ = _2689_ ^ _2696_ /*1841*/;
assign _2694_ = _2695_ | _2697_ /*1838*/;
assign _2703_ = ~D[2] /*1837*/;
assign _2700_ = _2562_ & _2703_ /*1833*/;
assign _2701_ = _2562_ ^ _2703_ /*1836*/;
assign _2702_ = _2694_ & _2701_ /*1834*/;
assign _2675_ = _2694_ ^ _2701_ /*1835*/;
assign _2699_ = _2700_ | _2702_ /*1832*/;
assign _2708_ = ~D[3] /*1831*/;
assign _2705_ = _2563_ & _2708_ /*1827*/;
assign _2706_ = _2563_ ^ _2708_ /*1830*/;
assign _2707_ = _2699_ & _2706_ /*1828*/;
assign _2676_ = _2699_ ^ _2706_ /*1829*/;
assign _2704_ = _2705_ | _2707_ /*1826*/;
assign _2713_ = ~D[4] /*1825*/;
assign _2710_ = _2564_ & _2713_ /*1821*/;
assign _2711_ = _2564_ ^ _2713_ /*1824*/;
assign _2712_ = _2704_ & _2711_ /*1822*/;
assign _2677_ = _2704_ ^ _2711_ /*1823*/;
assign _2709_ = _2710_ | _2712_ /*1820*/;
assign _2718_ = ~D[5] /*1819*/;
assign _2715_ = _2565_ & _2718_ /*1815*/;
assign _2716_ = _2565_ ^ _2718_ /*1818*/;
assign _2717_ = _2709_ & _2716_ /*1816*/;
assign _2678_ = _2709_ ^ _2716_ /*1817*/;
assign _2714_ = _2715_ | _2717_ /*1814*/;
assign _2723_ = ~D[6] /*1813*/;
assign _2720_ = _2566_ & _2723_ /*1809*/;
assign _2721_ = _2566_ ^ _2723_ /*1812*/;
assign _2722_ = _2714_ & _2721_ /*1810*/;
assign _2679_ = _2714_ ^ _2721_ /*1811*/;
assign _2719_ = _2720_ | _2722_ /*1808*/;
assign _2728_ = ~D[7] /*1807*/;
assign _2725_ = _2567_ & _2728_ /*1803*/;
assign _2726_ = _2567_ ^ _2728_ /*1806*/;
assign _2727_ = _2719_ & _2726_ /*1804*/;
assign _2680_ = _2719_ ^ _2726_ /*1805*/;
assign _2724_ = _2725_ | _2727_ /*1802*/;
assign _2733_ = ~D[8] /*1801*/;
assign _2730_ = _2568_ & _2733_ /*1797*/;
assign _2731_ = _2568_ ^ _2733_ /*1800*/;
assign _2732_ = _2724_ & _2731_ /*1798*/;
assign _2681_ = _2724_ ^ _2731_ /*1799*/;
assign _2729_ = _2730_ | _2732_ /*1796*/;
assign _2738_ = ~D[9] /*1795*/;
assign _2735_ = _2569_ & _2738_ /*1791*/;
assign _2736_ = _2569_ ^ _2738_ /*1794*/;
assign _2737_ = _2729_ & _2736_ /*1792*/;
assign _2682_ = _2729_ ^ _2736_ /*1793*/;
assign _2734_ = _2735_ | _2737_ /*1790*/;
assign _2743_ = ~D[10] /*1789*/;
assign _2740_ = _2570_ & _2743_ /*1785*/;
assign _2741_ = _2570_ ^ _2743_ /*1788*/;
assign _2742_ = _2734_ & _2741_ /*1786*/;
assign _2683_ = _2734_ ^ _2741_ /*1787*/;
assign _2739_ = _2740_ | _2742_ /*1784*/;
assign _2748_ = ~D[11] /*1783*/;
assign _2745_ = _2571_ & _2748_ /*1779*/;
assign _2746_ = _2571_ ^ _2748_ /*1782*/;
assign _2747_ = _2739_ & _2746_ /*1780*/;
assign _2684_ = _2739_ ^ _2746_ /*1781*/;
assign _2744_ = _2745_ | _2747_ /*1778*/;
assign _2753_ = ~D[12] /*1777*/;
assign _2750_ = _2572_ & _2753_ /*1773*/;
assign _2751_ = _2572_ ^ _2753_ /*1776*/;
assign _2752_ = _2744_ & _2751_ /*1774*/;
assign _2685_ = _2744_ ^ _2751_ /*1775*/;
assign _2749_ = _2750_ | _2752_ /*1772*/;
assign _2758_ = ~D[13] /*1771*/;
assign _2755_ = _2573_ & _2758_ /*1767*/;
assign _2756_ = _2573_ ^ _2758_ /*1770*/;
assign _2757_ = _2749_ & _2756_ /*1768*/;
assign _2686_ = _2749_ ^ _2756_ /*1769*/;
assign _2754_ = _2755_ | _2757_ /*1766*/;
assign _2763_ = ~D[14] /*1765*/;
assign _2760_ = _2574_ & _2763_ /*1761*/;
assign _2761_ = _2574_ ^ _2763_ /*1764*/;
assign _2762_ = _2754_ & _2761_ /*1762*/;
assign _2687_ = _2754_ ^ _2761_ /*1763*/;
assign _2759_ = _2760_ | _2762_ /*1760*/;
assign _2764_ = _2575_ & oneWire /*1755*/;
assign _2765_ = _2575_ ^ oneWire /*1758*/;
assign _2766_ = _2759_ & _2765_ /*1756*/;
assign _2688_ = _2759_ ^ _2765_ /*1757*/;
assign Q[3] = _2764_ | _2766_ /*1754*/;
assign _2803_ = ~Q[3] /*1657*/;
assign _2802_ = _2803_ & D[0] /*1656*/;
assign _2805_ = _2673_ & _2802_ /*1651*/;
assign _2806_ = _2673_ ^ _2802_ /*1654*/;
assign _2807_ = zeroWire & _2806_ /*1652*/;
assign _2785_ = zeroWire ^ _2806_ /*1653*/;
assign _2804_ = _2805_ | _2807_ /*1650*/;
assign _2809_ = ~Q[3] /*1649*/;
assign _2808_ = _2809_ & D[1] /*1648*/;
assign _2811_ = _2674_ & _2808_ /*1643*/;
assign _2812_ = _2674_ ^ _2808_ /*1646*/;
assign _2813_ = _2804_ & _2812_ /*1644*/;
assign _2786_ = _2804_ ^ _2812_ /*1645*/;
assign _2810_ = _2811_ | _2813_ /*1642*/;
assign _2815_ = ~Q[3] /*1641*/;
assign _2814_ = _2815_ & D[2] /*1640*/;
assign _2817_ = _2675_ & _2814_ /*1635*/;
assign _2818_ = _2675_ ^ _2814_ /*1638*/;
assign _2819_ = _2810_ & _2818_ /*1636*/;
assign _2787_ = _2810_ ^ _2818_ /*1637*/;
assign _2816_ = _2817_ | _2819_ /*1634*/;
assign _2821_ = ~Q[3] /*1633*/;
assign _2820_ = _2821_ & D[3] /*1632*/;
assign _2823_ = _2676_ & _2820_ /*1627*/;
assign _2824_ = _2676_ ^ _2820_ /*1630*/;
assign _2825_ = _2816_ & _2824_ /*1628*/;
assign _2788_ = _2816_ ^ _2824_ /*1629*/;
assign _2822_ = _2823_ | _2825_ /*1626*/;
assign _2827_ = ~Q[3] /*1625*/;
assign _2826_ = _2827_ & D[4] /*1624*/;
assign _2829_ = _2677_ & _2826_ /*1619*/;
assign _2830_ = _2677_ ^ _2826_ /*1622*/;
assign _2831_ = _2822_ & _2830_ /*1620*/;
assign _2789_ = _2822_ ^ _2830_ /*1621*/;
assign _2828_ = _2829_ | _2831_ /*1618*/;
assign _2833_ = ~Q[3] /*1617*/;
assign _2832_ = _2833_ & D[5] /*1616*/;
assign _2835_ = _2678_ & _2832_ /*1611*/;
assign _2836_ = _2678_ ^ _2832_ /*1614*/;
assign _2837_ = _2828_ & _2836_ /*1612*/;
assign _2790_ = _2828_ ^ _2836_ /*1613*/;
assign _2834_ = _2835_ | _2837_ /*1610*/;
assign _2839_ = ~Q[3] /*1609*/;
assign _2838_ = _2839_ & D[6] /*1608*/;
assign _2841_ = _2679_ & _2838_ /*1603*/;
assign _2842_ = _2679_ ^ _2838_ /*1606*/;
assign _2843_ = _2834_ & _2842_ /*1604*/;
assign _2791_ = _2834_ ^ _2842_ /*1605*/;
assign _2840_ = _2841_ | _2843_ /*1602*/;
assign _2845_ = ~Q[3] /*1601*/;
assign _2844_ = _2845_ & D[7] /*1600*/;
assign _2847_ = _2680_ & _2844_ /*1595*/;
assign _2848_ = _2680_ ^ _2844_ /*1598*/;
assign _2849_ = _2840_ & _2848_ /*1596*/;
assign _2792_ = _2840_ ^ _2848_ /*1597*/;
assign _2846_ = _2847_ | _2849_ /*1594*/;
assign _2851_ = ~Q[3] /*1593*/;
assign _2850_ = _2851_ & D[8] /*1592*/;
assign _2853_ = _2681_ & _2850_ /*1587*/;
assign _2854_ = _2681_ ^ _2850_ /*1590*/;
assign _2855_ = _2846_ & _2854_ /*1588*/;
assign _2793_ = _2846_ ^ _2854_ /*1589*/;
assign _2852_ = _2853_ | _2855_ /*1586*/;
assign _2857_ = ~Q[3] /*1585*/;
assign _2856_ = _2857_ & D[9] /*1584*/;
assign _2859_ = _2682_ & _2856_ /*1579*/;
assign _2860_ = _2682_ ^ _2856_ /*1582*/;
assign _2861_ = _2852_ & _2860_ /*1580*/;
assign _2794_ = _2852_ ^ _2860_ /*1581*/;
assign _2858_ = _2859_ | _2861_ /*1578*/;
assign _2863_ = ~Q[3] /*1577*/;
assign _2862_ = _2863_ & D[10] /*1576*/;
assign _2865_ = _2683_ & _2862_ /*1571*/;
assign _2866_ = _2683_ ^ _2862_ /*1574*/;
assign _2867_ = _2858_ & _2866_ /*1572*/;
assign _2795_ = _2858_ ^ _2866_ /*1573*/;
assign _2864_ = _2865_ | _2867_ /*1570*/;
assign _2869_ = ~Q[3] /*1569*/;
assign _2868_ = _2869_ & D[11] /*1568*/;
assign _2871_ = _2684_ & _2868_ /*1563*/;
assign _2872_ = _2684_ ^ _2868_ /*1566*/;
assign _2873_ = _2864_ & _2872_ /*1564*/;
assign _2796_ = _2864_ ^ _2872_ /*1565*/;
assign _2870_ = _2871_ | _2873_ /*1562*/;
assign _2875_ = ~Q[3] /*1561*/;
assign _2874_ = _2875_ & D[12] /*1560*/;
assign _2877_ = _2685_ & _2874_ /*1555*/;
assign _2878_ = _2685_ ^ _2874_ /*1558*/;
assign _2879_ = _2870_ & _2878_ /*1556*/;
assign _2797_ = _2870_ ^ _2878_ /*1557*/;
assign _2876_ = _2877_ | _2879_ /*1554*/;
assign _2881_ = ~Q[3] /*1553*/;
assign _2880_ = _2881_ & D[13] /*1552*/;
assign _2883_ = _2686_ & _2880_ /*1547*/;
assign _2884_ = _2686_ ^ _2880_ /*1550*/;
assign _2885_ = _2876_ & _2884_ /*1548*/;
assign _2798_ = _2876_ ^ _2884_ /*1549*/;
assign _2882_ = _2883_ | _2885_ /*1546*/;
assign _2887_ = ~Q[3] /*1545*/;
assign _2886_ = _2887_ & D[14] /*1544*/;
assign _2889_ = _2687_ & _2886_ /*1539*/;
assign _2890_ = _2687_ ^ _2886_ /*1542*/;
assign _2891_ = _2882_ & _2890_ /*1540*/;
assign _2799_ = _2882_ ^ _2890_ /*1541*/;
assign _2888_ = _2889_ | _2891_ /*1538*/;
assign _2893_ = ~Q[3] /*1537*/;
assign _2892_ = _2893_ & zeroWire /*1536*/;
assign _2894_ = _2688_ ^ _2892_ /*1534*/;
assign _2800_ = _2894_ ^ _2888_ /*1533*/;
assign _2917_ = ~D[0] /*1471*/;
assign _2914_ = R_0[2] & _2917_ /*1467*/;
assign _2915_ = R_0[2] ^ _2917_ /*1470*/;
assign _2916_ = oneWire & _2915_ /*1468*/;
assign _2897_ = oneWire ^ _2915_ /*1469*/;
assign _2913_ = _2914_ | _2916_ /*1466*/;
assign _2922_ = ~D[1] /*1465*/;
assign _2919_ = _2785_ & _2922_ /*1461*/;
assign _2920_ = _2785_ ^ _2922_ /*1464*/;
assign _2921_ = _2913_ & _2920_ /*1462*/;
assign _2898_ = _2913_ ^ _2920_ /*1463*/;
assign _2918_ = _2919_ | _2921_ /*1460*/;
assign _2927_ = ~D[2] /*1459*/;
assign _2924_ = _2786_ & _2927_ /*1455*/;
assign _2925_ = _2786_ ^ _2927_ /*1458*/;
assign _2926_ = _2918_ & _2925_ /*1456*/;
assign _2899_ = _2918_ ^ _2925_ /*1457*/;
assign _2923_ = _2924_ | _2926_ /*1454*/;
assign _2932_ = ~D[3] /*1453*/;
assign _2929_ = _2787_ & _2932_ /*1449*/;
assign _2930_ = _2787_ ^ _2932_ /*1452*/;
assign _2931_ = _2923_ & _2930_ /*1450*/;
assign _2900_ = _2923_ ^ _2930_ /*1451*/;
assign _2928_ = _2929_ | _2931_ /*1448*/;
assign _2937_ = ~D[4] /*1447*/;
assign _2934_ = _2788_ & _2937_ /*1443*/;
assign _2935_ = _2788_ ^ _2937_ /*1446*/;
assign _2936_ = _2928_ & _2935_ /*1444*/;
assign _2901_ = _2928_ ^ _2935_ /*1445*/;
assign _2933_ = _2934_ | _2936_ /*1442*/;
assign _2942_ = ~D[5] /*1441*/;
assign _2939_ = _2789_ & _2942_ /*1437*/;
assign _2940_ = _2789_ ^ _2942_ /*1440*/;
assign _2941_ = _2933_ & _2940_ /*1438*/;
assign _2902_ = _2933_ ^ _2940_ /*1439*/;
assign _2938_ = _2939_ | _2941_ /*1436*/;
assign _2947_ = ~D[6] /*1435*/;
assign _2944_ = _2790_ & _2947_ /*1431*/;
assign _2945_ = _2790_ ^ _2947_ /*1434*/;
assign _2946_ = _2938_ & _2945_ /*1432*/;
assign _2903_ = _2938_ ^ _2945_ /*1433*/;
assign _2943_ = _2944_ | _2946_ /*1430*/;
assign _2952_ = ~D[7] /*1429*/;
assign _2949_ = _2791_ & _2952_ /*1425*/;
assign _2950_ = _2791_ ^ _2952_ /*1428*/;
assign _2951_ = _2943_ & _2950_ /*1426*/;
assign _2904_ = _2943_ ^ _2950_ /*1427*/;
assign _2948_ = _2949_ | _2951_ /*1424*/;
assign _2957_ = ~D[8] /*1423*/;
assign _2954_ = _2792_ & _2957_ /*1419*/;
assign _2955_ = _2792_ ^ _2957_ /*1422*/;
assign _2956_ = _2948_ & _2955_ /*1420*/;
assign _2905_ = _2948_ ^ _2955_ /*1421*/;
assign _2953_ = _2954_ | _2956_ /*1418*/;
assign _2962_ = ~D[9] /*1417*/;
assign _2959_ = _2793_ & _2962_ /*1413*/;
assign _2960_ = _2793_ ^ _2962_ /*1416*/;
assign _2961_ = _2953_ & _2960_ /*1414*/;
assign _2906_ = _2953_ ^ _2960_ /*1415*/;
assign _2958_ = _2959_ | _2961_ /*1412*/;
assign _2967_ = ~D[10] /*1411*/;
assign _2964_ = _2794_ & _2967_ /*1407*/;
assign _2965_ = _2794_ ^ _2967_ /*1410*/;
assign _2966_ = _2958_ & _2965_ /*1408*/;
assign _2907_ = _2958_ ^ _2965_ /*1409*/;
assign _2963_ = _2964_ | _2966_ /*1406*/;
assign _2972_ = ~D[11] /*1405*/;
assign _2969_ = _2795_ & _2972_ /*1401*/;
assign _2970_ = _2795_ ^ _2972_ /*1404*/;
assign _2971_ = _2963_ & _2970_ /*1402*/;
assign _2908_ = _2963_ ^ _2970_ /*1403*/;
assign _2968_ = _2969_ | _2971_ /*1400*/;
assign _2977_ = ~D[12] /*1399*/;
assign _2974_ = _2796_ & _2977_ /*1395*/;
assign _2975_ = _2796_ ^ _2977_ /*1398*/;
assign _2976_ = _2968_ & _2975_ /*1396*/;
assign _2909_ = _2968_ ^ _2975_ /*1397*/;
assign _2973_ = _2974_ | _2976_ /*1394*/;
assign _2982_ = ~D[13] /*1393*/;
assign _2979_ = _2797_ & _2982_ /*1389*/;
assign _2980_ = _2797_ ^ _2982_ /*1392*/;
assign _2981_ = _2973_ & _2980_ /*1390*/;
assign _2910_ = _2973_ ^ _2980_ /*1391*/;
assign _2978_ = _2979_ | _2981_ /*1388*/;
assign _2987_ = ~D[14] /*1387*/;
assign _2984_ = _2798_ & _2987_ /*1383*/;
assign _2985_ = _2798_ ^ _2987_ /*1386*/;
assign _2986_ = _2978_ & _2985_ /*1384*/;
assign _2911_ = _2978_ ^ _2985_ /*1385*/;
assign _2983_ = _2984_ | _2986_ /*1382*/;
assign _2988_ = _2799_ & oneWire /*1377*/;
assign _2989_ = _2799_ ^ oneWire /*1380*/;
assign _2990_ = _2983_ & _2989_ /*1378*/;
assign _2912_ = _2983_ ^ _2989_ /*1379*/;
assign Q[2] = _2988_ | _2990_ /*1376*/;
assign _3027_ = ~Q[2] /*1279*/;
assign _3026_ = _3027_ & D[0] /*1278*/;
assign _3029_ = _2897_ & _3026_ /*1273*/;
assign _3030_ = _2897_ ^ _3026_ /*1276*/;
assign _3031_ = zeroWire & _3030_ /*1274*/;
assign _3009_ = zeroWire ^ _3030_ /*1275*/;
assign _3028_ = _3029_ | _3031_ /*1272*/;
assign _3033_ = ~Q[2] /*1271*/;
assign _3032_ = _3033_ & D[1] /*1270*/;
assign _3035_ = _2898_ & _3032_ /*1265*/;
assign _3036_ = _2898_ ^ _3032_ /*1268*/;
assign _3037_ = _3028_ & _3036_ /*1266*/;
assign _3010_ = _3028_ ^ _3036_ /*1267*/;
assign _3034_ = _3035_ | _3037_ /*1264*/;
assign _3039_ = ~Q[2] /*1263*/;
assign _3038_ = _3039_ & D[2] /*1262*/;
assign _3041_ = _2899_ & _3038_ /*1257*/;
assign _3042_ = _2899_ ^ _3038_ /*1260*/;
assign _3043_ = _3034_ & _3042_ /*1258*/;
assign _3011_ = _3034_ ^ _3042_ /*1259*/;
assign _3040_ = _3041_ | _3043_ /*1256*/;
assign _3045_ = ~Q[2] /*1255*/;
assign _3044_ = _3045_ & D[3] /*1254*/;
assign _3047_ = _2900_ & _3044_ /*1249*/;
assign _3048_ = _2900_ ^ _3044_ /*1252*/;
assign _3049_ = _3040_ & _3048_ /*1250*/;
assign _3012_ = _3040_ ^ _3048_ /*1251*/;
assign _3046_ = _3047_ | _3049_ /*1248*/;
assign _3051_ = ~Q[2] /*1247*/;
assign _3050_ = _3051_ & D[4] /*1246*/;
assign _3053_ = _2901_ & _3050_ /*1241*/;
assign _3054_ = _2901_ ^ _3050_ /*1244*/;
assign _3055_ = _3046_ & _3054_ /*1242*/;
assign _3013_ = _3046_ ^ _3054_ /*1243*/;
assign _3052_ = _3053_ | _3055_ /*1240*/;
assign _3057_ = ~Q[2] /*1239*/;
assign _3056_ = _3057_ & D[5] /*1238*/;
assign _3059_ = _2902_ & _3056_ /*1233*/;
assign _3060_ = _2902_ ^ _3056_ /*1236*/;
assign _3061_ = _3052_ & _3060_ /*1234*/;
assign _3014_ = _3052_ ^ _3060_ /*1235*/;
assign _3058_ = _3059_ | _3061_ /*1232*/;
assign _3063_ = ~Q[2] /*1231*/;
assign _3062_ = _3063_ & D[6] /*1230*/;
assign _3065_ = _2903_ & _3062_ /*1225*/;
assign _3066_ = _2903_ ^ _3062_ /*1228*/;
assign _3067_ = _3058_ & _3066_ /*1226*/;
assign _3015_ = _3058_ ^ _3066_ /*1227*/;
assign _3064_ = _3065_ | _3067_ /*1224*/;
assign _3069_ = ~Q[2] /*1223*/;
assign _3068_ = _3069_ & D[7] /*1222*/;
assign _3071_ = _2904_ & _3068_ /*1217*/;
assign _3072_ = _2904_ ^ _3068_ /*1220*/;
assign _3073_ = _3064_ & _3072_ /*1218*/;
assign _3016_ = _3064_ ^ _3072_ /*1219*/;
assign _3070_ = _3071_ | _3073_ /*1216*/;
assign _3075_ = ~Q[2] /*1215*/;
assign _3074_ = _3075_ & D[8] /*1214*/;
assign _3077_ = _2905_ & _3074_ /*1209*/;
assign _3078_ = _2905_ ^ _3074_ /*1212*/;
assign _3079_ = _3070_ & _3078_ /*1210*/;
assign _3017_ = _3070_ ^ _3078_ /*1211*/;
assign _3076_ = _3077_ | _3079_ /*1208*/;
assign _3081_ = ~Q[2] /*1207*/;
assign _3080_ = _3081_ & D[9] /*1206*/;
assign _3083_ = _2906_ & _3080_ /*1201*/;
assign _3084_ = _2906_ ^ _3080_ /*1204*/;
assign _3085_ = _3076_ & _3084_ /*1202*/;
assign _3018_ = _3076_ ^ _3084_ /*1203*/;
assign _3082_ = _3083_ | _3085_ /*1200*/;
assign _3087_ = ~Q[2] /*1199*/;
assign _3086_ = _3087_ & D[10] /*1198*/;
assign _3089_ = _2907_ & _3086_ /*1193*/;
assign _3090_ = _2907_ ^ _3086_ /*1196*/;
assign _3091_ = _3082_ & _3090_ /*1194*/;
assign _3019_ = _3082_ ^ _3090_ /*1195*/;
assign _3088_ = _3089_ | _3091_ /*1192*/;
assign _3093_ = ~Q[2] /*1191*/;
assign _3092_ = _3093_ & D[11] /*1190*/;
assign _3095_ = _2908_ & _3092_ /*1185*/;
assign _3096_ = _2908_ ^ _3092_ /*1188*/;
assign _3097_ = _3088_ & _3096_ /*1186*/;
assign _3020_ = _3088_ ^ _3096_ /*1187*/;
assign _3094_ = _3095_ | _3097_ /*1184*/;
assign _3099_ = ~Q[2] /*1183*/;
assign _3098_ = _3099_ & D[12] /*1182*/;
assign _3101_ = _2909_ & _3098_ /*1177*/;
assign _3102_ = _2909_ ^ _3098_ /*1180*/;
assign _3103_ = _3094_ & _3102_ /*1178*/;
assign _3021_ = _3094_ ^ _3102_ /*1179*/;
assign _3100_ = _3101_ | _3103_ /*1176*/;
assign _3105_ = ~Q[2] /*1175*/;
assign _3104_ = _3105_ & D[13] /*1174*/;
assign _3107_ = _2910_ & _3104_ /*1169*/;
assign _3108_ = _2910_ ^ _3104_ /*1172*/;
assign _3109_ = _3100_ & _3108_ /*1170*/;
assign _3022_ = _3100_ ^ _3108_ /*1171*/;
assign _3106_ = _3107_ | _3109_ /*1168*/;
assign _3111_ = ~Q[2] /*1167*/;
assign _3110_ = _3111_ & D[14] /*1166*/;
assign _3113_ = _2911_ & _3110_ /*1161*/;
assign _3114_ = _2911_ ^ _3110_ /*1164*/;
assign _3115_ = _3106_ & _3114_ /*1162*/;
assign _3023_ = _3106_ ^ _3114_ /*1163*/;
assign _3112_ = _3113_ | _3115_ /*1160*/;
assign _3117_ = ~Q[2] /*1159*/;
assign _3116_ = _3117_ & zeroWire /*1158*/;
assign _3118_ = _2912_ ^ _3116_ /*1156*/;
assign _3024_ = _3118_ ^ _3112_ /*1155*/;
assign _3141_ = ~D[0] /*1093*/;
assign _3138_ = R_0[1] & _3141_ /*1089*/;
assign _3139_ = R_0[1] ^ _3141_ /*1092*/;
assign _3140_ = oneWire & _3139_ /*1090*/;
assign _3121_ = oneWire ^ _3139_ /*1091*/;
assign _3137_ = _3138_ | _3140_ /*1088*/;
assign _3146_ = ~D[1] /*1087*/;
assign _3143_ = _3009_ & _3146_ /*1083*/;
assign _3144_ = _3009_ ^ _3146_ /*1086*/;
assign _3145_ = _3137_ & _3144_ /*1084*/;
assign _3122_ = _3137_ ^ _3144_ /*1085*/;
assign _3142_ = _3143_ | _3145_ /*1082*/;
assign _3151_ = ~D[2] /*1081*/;
assign _3148_ = _3010_ & _3151_ /*1077*/;
assign _3149_ = _3010_ ^ _3151_ /*1080*/;
assign _3150_ = _3142_ & _3149_ /*1078*/;
assign _3123_ = _3142_ ^ _3149_ /*1079*/;
assign _3147_ = _3148_ | _3150_ /*1076*/;
assign _3156_ = ~D[3] /*1075*/;
assign _3153_ = _3011_ & _3156_ /*1071*/;
assign _3154_ = _3011_ ^ _3156_ /*1074*/;
assign _3155_ = _3147_ & _3154_ /*1072*/;
assign _3124_ = _3147_ ^ _3154_ /*1073*/;
assign _3152_ = _3153_ | _3155_ /*1070*/;
assign _3161_ = ~D[4] /*1069*/;
assign _3158_ = _3012_ & _3161_ /*1065*/;
assign _3159_ = _3012_ ^ _3161_ /*1068*/;
assign _3160_ = _3152_ & _3159_ /*1066*/;
assign _3125_ = _3152_ ^ _3159_ /*1067*/;
assign _3157_ = _3158_ | _3160_ /*1064*/;
assign _3166_ = ~D[5] /*1063*/;
assign _3163_ = _3013_ & _3166_ /*1059*/;
assign _3164_ = _3013_ ^ _3166_ /*1062*/;
assign _3165_ = _3157_ & _3164_ /*1060*/;
assign _3126_ = _3157_ ^ _3164_ /*1061*/;
assign _3162_ = _3163_ | _3165_ /*1058*/;
assign _3171_ = ~D[6] /*1057*/;
assign _3168_ = _3014_ & _3171_ /*1053*/;
assign _3169_ = _3014_ ^ _3171_ /*1056*/;
assign _3170_ = _3162_ & _3169_ /*1054*/;
assign _3127_ = _3162_ ^ _3169_ /*1055*/;
assign _3167_ = _3168_ | _3170_ /*1052*/;
assign _3176_ = ~D[7] /*1051*/;
assign _3173_ = _3015_ & _3176_ /*1047*/;
assign _3174_ = _3015_ ^ _3176_ /*1050*/;
assign _3175_ = _3167_ & _3174_ /*1048*/;
assign _3128_ = _3167_ ^ _3174_ /*1049*/;
assign _3172_ = _3173_ | _3175_ /*1046*/;
assign _3181_ = ~D[8] /*1045*/;
assign _3178_ = _3016_ & _3181_ /*1041*/;
assign _3179_ = _3016_ ^ _3181_ /*1044*/;
assign _3180_ = _3172_ & _3179_ /*1042*/;
assign _3129_ = _3172_ ^ _3179_ /*1043*/;
assign _3177_ = _3178_ | _3180_ /*1040*/;
assign _3186_ = ~D[9] /*1039*/;
assign _3183_ = _3017_ & _3186_ /*1035*/;
assign _3184_ = _3017_ ^ _3186_ /*1038*/;
assign _3185_ = _3177_ & _3184_ /*1036*/;
assign _3130_ = _3177_ ^ _3184_ /*1037*/;
assign _3182_ = _3183_ | _3185_ /*1034*/;
assign _3191_ = ~D[10] /*1033*/;
assign _3188_ = _3018_ & _3191_ /*1029*/;
assign _3189_ = _3018_ ^ _3191_ /*1032*/;
assign _3190_ = _3182_ & _3189_ /*1030*/;
assign _3131_ = _3182_ ^ _3189_ /*1031*/;
assign _3187_ = _3188_ | _3190_ /*1028*/;
assign _3196_ = ~D[11] /*1027*/;
assign _3193_ = _3019_ & _3196_ /*1023*/;
assign _3194_ = _3019_ ^ _3196_ /*1026*/;
assign _3195_ = _3187_ & _3194_ /*1024*/;
assign _3132_ = _3187_ ^ _3194_ /*1025*/;
assign _3192_ = _3193_ | _3195_ /*1022*/;
assign _3201_ = ~D[12] /*1021*/;
assign _3198_ = _3020_ & _3201_ /*1017*/;
assign _3199_ = _3020_ ^ _3201_ /*1020*/;
assign _3200_ = _3192_ & _3199_ /*1018*/;
assign _3133_ = _3192_ ^ _3199_ /*1019*/;
assign _3197_ = _3198_ | _3200_ /*1016*/;
assign _3206_ = ~D[13] /*1015*/;
assign _3203_ = _3021_ & _3206_ /*1011*/;
assign _3204_ = _3021_ ^ _3206_ /*1014*/;
assign _3205_ = _3197_ & _3204_ /*1012*/;
assign _3134_ = _3197_ ^ _3204_ /*1013*/;
assign _3202_ = _3203_ | _3205_ /*1010*/;
assign _3211_ = ~D[14] /*1009*/;
assign _3208_ = _3022_ & _3211_ /*1005*/;
assign _3209_ = _3022_ ^ _3211_ /*1008*/;
assign _3210_ = _3202_ & _3209_ /*1006*/;
assign _3135_ = _3202_ ^ _3209_ /*1007*/;
assign _3207_ = _3208_ | _3210_ /*1004*/;
assign _3212_ = _3023_ & oneWire /*999*/;
assign _3213_ = _3023_ ^ oneWire /*1002*/;
assign _3214_ = _3207_ & _3213_ /*1000*/;
assign _3136_ = _3207_ ^ _3213_ /*1001*/;
assign Q[1] = _3212_ | _3214_ /*998*/;
assign _3251_ = ~Q[1] /*901*/;
assign _3250_ = _3251_ & D[0] /*900*/;
assign _3253_ = _3121_ & _3250_ /*895*/;
assign _3254_ = _3121_ ^ _3250_ /*898*/;
assign _3255_ = zeroWire & _3254_ /*896*/;
assign _3233_ = zeroWire ^ _3254_ /*897*/;
assign _3252_ = _3253_ | _3255_ /*894*/;
assign _3257_ = ~Q[1] /*893*/;
assign _3256_ = _3257_ & D[1] /*892*/;
assign _3259_ = _3122_ & _3256_ /*887*/;
assign _3260_ = _3122_ ^ _3256_ /*890*/;
assign _3261_ = _3252_ & _3260_ /*888*/;
assign _3234_ = _3252_ ^ _3260_ /*889*/;
assign _3258_ = _3259_ | _3261_ /*886*/;
assign _3263_ = ~Q[1] /*885*/;
assign _3262_ = _3263_ & D[2] /*884*/;
assign _3265_ = _3123_ & _3262_ /*879*/;
assign _3266_ = _3123_ ^ _3262_ /*882*/;
assign _3267_ = _3258_ & _3266_ /*880*/;
assign _3235_ = _3258_ ^ _3266_ /*881*/;
assign _3264_ = _3265_ | _3267_ /*878*/;
assign _3269_ = ~Q[1] /*877*/;
assign _3268_ = _3269_ & D[3] /*876*/;
assign _3271_ = _3124_ & _3268_ /*871*/;
assign _3272_ = _3124_ ^ _3268_ /*874*/;
assign _3273_ = _3264_ & _3272_ /*872*/;
assign _3236_ = _3264_ ^ _3272_ /*873*/;
assign _3270_ = _3271_ | _3273_ /*870*/;
assign _3275_ = ~Q[1] /*869*/;
assign _3274_ = _3275_ & D[4] /*868*/;
assign _3277_ = _3125_ & _3274_ /*863*/;
assign _3278_ = _3125_ ^ _3274_ /*866*/;
assign _3279_ = _3270_ & _3278_ /*864*/;
assign _3237_ = _3270_ ^ _3278_ /*865*/;
assign _3276_ = _3277_ | _3279_ /*862*/;
assign _3281_ = ~Q[1] /*861*/;
assign _3280_ = _3281_ & D[5] /*860*/;
assign _3283_ = _3126_ & _3280_ /*855*/;
assign _3284_ = _3126_ ^ _3280_ /*858*/;
assign _3285_ = _3276_ & _3284_ /*856*/;
assign _3238_ = _3276_ ^ _3284_ /*857*/;
assign _3282_ = _3283_ | _3285_ /*854*/;
assign _3287_ = ~Q[1] /*853*/;
assign _3286_ = _3287_ & D[6] /*852*/;
assign _3289_ = _3127_ & _3286_ /*847*/;
assign _3290_ = _3127_ ^ _3286_ /*850*/;
assign _3291_ = _3282_ & _3290_ /*848*/;
assign _3239_ = _3282_ ^ _3290_ /*849*/;
assign _3288_ = _3289_ | _3291_ /*846*/;
assign _3293_ = ~Q[1] /*845*/;
assign _3292_ = _3293_ & D[7] /*844*/;
assign _3295_ = _3128_ & _3292_ /*839*/;
assign _3296_ = _3128_ ^ _3292_ /*842*/;
assign _3297_ = _3288_ & _3296_ /*840*/;
assign _3240_ = _3288_ ^ _3296_ /*841*/;
assign _3294_ = _3295_ | _3297_ /*838*/;
assign _3299_ = ~Q[1] /*837*/;
assign _3298_ = _3299_ & D[8] /*836*/;
assign _3301_ = _3129_ & _3298_ /*831*/;
assign _3302_ = _3129_ ^ _3298_ /*834*/;
assign _3303_ = _3294_ & _3302_ /*832*/;
assign _3241_ = _3294_ ^ _3302_ /*833*/;
assign _3300_ = _3301_ | _3303_ /*830*/;
assign _3305_ = ~Q[1] /*829*/;
assign _3304_ = _3305_ & D[9] /*828*/;
assign _3307_ = _3130_ & _3304_ /*823*/;
assign _3308_ = _3130_ ^ _3304_ /*826*/;
assign _3309_ = _3300_ & _3308_ /*824*/;
assign _3242_ = _3300_ ^ _3308_ /*825*/;
assign _3306_ = _3307_ | _3309_ /*822*/;
assign _3311_ = ~Q[1] /*821*/;
assign _3310_ = _3311_ & D[10] /*820*/;
assign _3313_ = _3131_ & _3310_ /*815*/;
assign _3314_ = _3131_ ^ _3310_ /*818*/;
assign _3315_ = _3306_ & _3314_ /*816*/;
assign _3243_ = _3306_ ^ _3314_ /*817*/;
assign _3312_ = _3313_ | _3315_ /*814*/;
assign _3317_ = ~Q[1] /*813*/;
assign _3316_ = _3317_ & D[11] /*812*/;
assign _3319_ = _3132_ & _3316_ /*807*/;
assign _3320_ = _3132_ ^ _3316_ /*810*/;
assign _3321_ = _3312_ & _3320_ /*808*/;
assign _3244_ = _3312_ ^ _3320_ /*809*/;
assign _3318_ = _3319_ | _3321_ /*806*/;
assign _3323_ = ~Q[1] /*805*/;
assign _3322_ = _3323_ & D[12] /*804*/;
assign _3325_ = _3133_ & _3322_ /*799*/;
assign _3326_ = _3133_ ^ _3322_ /*802*/;
assign _3327_ = _3318_ & _3326_ /*800*/;
assign _3245_ = _3318_ ^ _3326_ /*801*/;
assign _3324_ = _3325_ | _3327_ /*798*/;
assign _3329_ = ~Q[1] /*797*/;
assign _3328_ = _3329_ & D[13] /*796*/;
assign _3331_ = _3134_ & _3328_ /*791*/;
assign _3332_ = _3134_ ^ _3328_ /*794*/;
assign _3333_ = _3324_ & _3332_ /*792*/;
assign _3246_ = _3324_ ^ _3332_ /*793*/;
assign _3330_ = _3331_ | _3333_ /*790*/;
assign _3335_ = ~Q[1] /*789*/;
assign _3334_ = _3335_ & D[14] /*788*/;
assign _3337_ = _3135_ & _3334_ /*783*/;
assign _3338_ = _3135_ ^ _3334_ /*786*/;
assign _3339_ = _3330_ & _3338_ /*784*/;
assign _3247_ = _3330_ ^ _3338_ /*785*/;
assign _3336_ = _3337_ | _3339_ /*782*/;
assign _3341_ = ~Q[1] /*781*/;
assign _3340_ = _3341_ & zeroWire /*780*/;
assign _3342_ = _3136_ ^ _3340_ /*778*/;
assign _3248_ = _3342_ ^ _3336_ /*777*/;
assign _3365_ = ~D[0] /*715*/;
assign _3362_ = R_0[0] & _3365_ /*711*/;
assign _3363_ = R_0[0] ^ _3365_ /*714*/;
assign _3364_ = oneWire & _3363_ /*712*/;
assign _3345_ = oneWire ^ _3363_ /*713*/;
assign _3361_ = _3362_ | _3364_ /*710*/;
assign _3370_ = ~D[1] /*709*/;
assign _3367_ = _3233_ & _3370_ /*705*/;
assign _3368_ = _3233_ ^ _3370_ /*708*/;
assign _3369_ = _3361_ & _3368_ /*706*/;
assign _3346_ = _3361_ ^ _3368_ /*707*/;
assign _3366_ = _3367_ | _3369_ /*704*/;
assign _3375_ = ~D[2] /*703*/;
assign _3372_ = _3234_ & _3375_ /*699*/;
assign _3373_ = _3234_ ^ _3375_ /*702*/;
assign _3374_ = _3366_ & _3373_ /*700*/;
assign _3347_ = _3366_ ^ _3373_ /*701*/;
assign _3371_ = _3372_ | _3374_ /*698*/;
assign _3380_ = ~D[3] /*697*/;
assign _3377_ = _3235_ & _3380_ /*693*/;
assign _3378_ = _3235_ ^ _3380_ /*696*/;
assign _3379_ = _3371_ & _3378_ /*694*/;
assign _3348_ = _3371_ ^ _3378_ /*695*/;
assign _3376_ = _3377_ | _3379_ /*692*/;
assign _3385_ = ~D[4] /*691*/;
assign _3382_ = _3236_ & _3385_ /*687*/;
assign _3383_ = _3236_ ^ _3385_ /*690*/;
assign _3384_ = _3376_ & _3383_ /*688*/;
assign _3349_ = _3376_ ^ _3383_ /*689*/;
assign _3381_ = _3382_ | _3384_ /*686*/;
assign _3390_ = ~D[5] /*685*/;
assign _3387_ = _3237_ & _3390_ /*681*/;
assign _3388_ = _3237_ ^ _3390_ /*684*/;
assign _3389_ = _3381_ & _3388_ /*682*/;
assign _3350_ = _3381_ ^ _3388_ /*683*/;
assign _3386_ = _3387_ | _3389_ /*680*/;
assign _3395_ = ~D[6] /*679*/;
assign _3392_ = _3238_ & _3395_ /*675*/;
assign _3393_ = _3238_ ^ _3395_ /*678*/;
assign _3394_ = _3386_ & _3393_ /*676*/;
assign _3351_ = _3386_ ^ _3393_ /*677*/;
assign _3391_ = _3392_ | _3394_ /*674*/;
assign _3400_ = ~D[7] /*673*/;
assign _3397_ = _3239_ & _3400_ /*669*/;
assign _3398_ = _3239_ ^ _3400_ /*672*/;
assign _3399_ = _3391_ & _3398_ /*670*/;
assign _3352_ = _3391_ ^ _3398_ /*671*/;
assign _3396_ = _3397_ | _3399_ /*668*/;
assign _3405_ = ~D[8] /*667*/;
assign _3402_ = _3240_ & _3405_ /*663*/;
assign _3403_ = _3240_ ^ _3405_ /*666*/;
assign _3404_ = _3396_ & _3403_ /*664*/;
assign _3353_ = _3396_ ^ _3403_ /*665*/;
assign _3401_ = _3402_ | _3404_ /*662*/;
assign _3410_ = ~D[9] /*661*/;
assign _3407_ = _3241_ & _3410_ /*657*/;
assign _3408_ = _3241_ ^ _3410_ /*660*/;
assign _3409_ = _3401_ & _3408_ /*658*/;
assign _3354_ = _3401_ ^ _3408_ /*659*/;
assign _3406_ = _3407_ | _3409_ /*656*/;
assign _3415_ = ~D[10] /*655*/;
assign _3412_ = _3242_ & _3415_ /*651*/;
assign _3413_ = _3242_ ^ _3415_ /*654*/;
assign _3414_ = _3406_ & _3413_ /*652*/;
assign _3355_ = _3406_ ^ _3413_ /*653*/;
assign _3411_ = _3412_ | _3414_ /*650*/;
assign _3420_ = ~D[11] /*649*/;
assign _3417_ = _3243_ & _3420_ /*645*/;
assign _3418_ = _3243_ ^ _3420_ /*648*/;
assign _3419_ = _3411_ & _3418_ /*646*/;
assign _3356_ = _3411_ ^ _3418_ /*647*/;
assign _3416_ = _3417_ | _3419_ /*644*/;
assign _3425_ = ~D[12] /*643*/;
assign _3422_ = _3244_ & _3425_ /*639*/;
assign _3423_ = _3244_ ^ _3425_ /*642*/;
assign _3424_ = _3416_ & _3423_ /*640*/;
assign _3357_ = _3416_ ^ _3423_ /*641*/;
assign _3421_ = _3422_ | _3424_ /*638*/;
assign _3430_ = ~D[13] /*637*/;
assign _3427_ = _3245_ & _3430_ /*633*/;
assign _3428_ = _3245_ ^ _3430_ /*636*/;
assign _3429_ = _3421_ & _3428_ /*634*/;
assign _3358_ = _3421_ ^ _3428_ /*635*/;
assign _3426_ = _3427_ | _3429_ /*632*/;
assign _3435_ = ~D[14] /*631*/;
assign _3432_ = _3246_ & _3435_ /*627*/;
assign _3433_ = _3246_ ^ _3435_ /*630*/;
assign _3434_ = _3426_ & _3433_ /*628*/;
assign _3359_ = _3426_ ^ _3433_ /*629*/;
assign _3431_ = _3432_ | _3434_ /*626*/;
assign _3436_ = _3247_ & oneWire /*621*/;
assign _3437_ = _3247_ ^ oneWire /*624*/;
assign _3438_ = _3431_ & _3437_ /*622*/;
assign _3360_ = _3431_ ^ _3437_ /*623*/;
assign Q[0] = _3436_ | _3438_ /*620*/;
assign _3475_ = ~Q[0] /*523*/;
assign _3474_ = _3475_ & D[0] /*522*/;
assign _3477_ = _3345_ & _3474_ /*517*/;
assign _3478_ = _3345_ ^ _3474_ /*520*/;
assign _3479_ = zeroWire & _3478_ /*518*/;
assign R_n1[0] = zeroWire ^ _3478_ /*519*/;
assign _3476_ = _3477_ | _3479_ /*516*/;
assign _3481_ = ~Q[0] /*515*/;
assign _3480_ = _3481_ & D[1] /*514*/;
assign _3483_ = _3346_ & _3480_ /*509*/;
assign _3484_ = _3346_ ^ _3480_ /*512*/;
assign _3485_ = _3476_ & _3484_ /*510*/;
assign R_n1[1] = _3476_ ^ _3484_ /*511*/;
assign _3482_ = _3483_ | _3485_ /*508*/;
assign _3487_ = ~Q[0] /*507*/;
assign _3486_ = _3487_ & D[2] /*506*/;
assign _3489_ = _3347_ & _3486_ /*501*/;
assign _3490_ = _3347_ ^ _3486_ /*504*/;
assign _3491_ = _3482_ & _3490_ /*502*/;
assign R_n1[2] = _3482_ ^ _3490_ /*503*/;
assign _3488_ = _3489_ | _3491_ /*500*/;
assign _3493_ = ~Q[0] /*499*/;
assign _3492_ = _3493_ & D[3] /*498*/;
assign _3495_ = _3348_ & _3492_ /*493*/;
assign _3496_ = _3348_ ^ _3492_ /*496*/;
assign _3497_ = _3488_ & _3496_ /*494*/;
assign R_n1[3] = _3488_ ^ _3496_ /*495*/;
assign _3494_ = _3495_ | _3497_ /*492*/;
assign _3499_ = ~Q[0] /*491*/;
assign _3498_ = _3499_ & D[4] /*490*/;
assign _3501_ = _3349_ & _3498_ /*485*/;
assign _3502_ = _3349_ ^ _3498_ /*488*/;
assign _3503_ = _3494_ & _3502_ /*486*/;
assign R_n1[4] = _3494_ ^ _3502_ /*487*/;
assign _3500_ = _3501_ | _3503_ /*484*/;
assign _3505_ = ~Q[0] /*483*/;
assign _3504_ = _3505_ & D[5] /*482*/;
assign _3507_ = _3350_ & _3504_ /*477*/;
assign _3508_ = _3350_ ^ _3504_ /*480*/;
assign _3509_ = _3500_ & _3508_ /*478*/;
assign R_n1[5] = _3500_ ^ _3508_ /*479*/;
assign _3506_ = _3507_ | _3509_ /*476*/;
assign _3511_ = ~Q[0] /*475*/;
assign _3510_ = _3511_ & D[6] /*474*/;
assign _3513_ = _3351_ & _3510_ /*469*/;
assign _3514_ = _3351_ ^ _3510_ /*472*/;
assign _3515_ = _3506_ & _3514_ /*470*/;
assign R_n1[6] = _3506_ ^ _3514_ /*471*/;
assign _3512_ = _3513_ | _3515_ /*468*/;
assign _3517_ = ~Q[0] /*467*/;
assign _3516_ = _3517_ & D[7] /*466*/;
assign _3519_ = _3352_ & _3516_ /*461*/;
assign _3520_ = _3352_ ^ _3516_ /*464*/;
assign _3521_ = _3512_ & _3520_ /*462*/;
assign R_n1[7] = _3512_ ^ _3520_ /*463*/;
assign _3518_ = _3519_ | _3521_ /*460*/;
assign _3523_ = ~Q[0] /*459*/;
assign _3522_ = _3523_ & D[8] /*458*/;
assign _3525_ = _3353_ & _3522_ /*453*/;
assign _3526_ = _3353_ ^ _3522_ /*456*/;
assign _3527_ = _3518_ & _3526_ /*454*/;
assign R_n1[8] = _3518_ ^ _3526_ /*455*/;
assign _3524_ = _3525_ | _3527_ /*452*/;
assign _3529_ = ~Q[0] /*451*/;
assign _3528_ = _3529_ & D[9] /*450*/;
assign _3531_ = _3354_ & _3528_ /*445*/;
assign _3532_ = _3354_ ^ _3528_ /*448*/;
assign _3533_ = _3524_ & _3532_ /*446*/;
assign R_n1[9] = _3524_ ^ _3532_ /*447*/;
assign _3530_ = _3531_ | _3533_ /*444*/;
assign _3535_ = ~Q[0] /*443*/;
assign _3534_ = _3535_ & D[10] /*442*/;
assign _3537_ = _3355_ & _3534_ /*437*/;
assign _3538_ = _3355_ ^ _3534_ /*440*/;
assign _3539_ = _3530_ & _3538_ /*438*/;
assign R_n1[10] = _3530_ ^ _3538_ /*439*/;
assign _3536_ = _3537_ | _3539_ /*436*/;
assign _3541_ = ~Q[0] /*435*/;
assign _3540_ = _3541_ & D[11] /*434*/;
assign _3543_ = _3356_ & _3540_ /*429*/;
assign _3544_ = _3356_ ^ _3540_ /*432*/;
assign _3545_ = _3536_ & _3544_ /*430*/;
assign R_n1[11] = _3536_ ^ _3544_ /*431*/;
assign _3542_ = _3543_ | _3545_ /*428*/;
assign _3547_ = ~Q[0] /*427*/;
assign _3546_ = _3547_ & D[12] /*426*/;
assign _3549_ = _3357_ & _3546_ /*421*/;
assign _3550_ = _3357_ ^ _3546_ /*424*/;
assign _3551_ = _3542_ & _3550_ /*422*/;
assign R_n1[12] = _3542_ ^ _3550_ /*423*/;
assign _3548_ = _3549_ | _3551_ /*420*/;
assign _3553_ = ~Q[0] /*419*/;
assign _3552_ = _3553_ & D[13] /*418*/;
assign _3555_ = _3358_ & _3552_ /*413*/;
assign _3556_ = _3358_ ^ _3552_ /*416*/;
assign _3557_ = _3548_ & _3556_ /*414*/;
assign R_n1[13] = _3548_ ^ _3556_ /*415*/;
assign _3554_ = _3555_ | _3557_ /*412*/;
assign _3559_ = ~Q[0] /*411*/;
assign _3558_ = _3559_ & D[14] /*410*/;
assign _3561_ = _3359_ & _3558_ /*405*/;
assign _3562_ = _3359_ ^ _3558_ /*408*/;
assign _3563_ = _3554_ & _3562_ /*406*/;
assign R_n1[14] = _3554_ ^ _3562_ /*407*/;
assign _3560_ = _3561_ | _3563_ /*404*/;
endmodule
