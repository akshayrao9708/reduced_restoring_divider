module divider(R_0, D, Q, R_n1);
input [5:0] R_0;
input [2:0] D;
output [3:0] Q;
output [2:0] R_n1;
wire _0_;
wire _1_;
wire _2_;
wire _3_;
wire _4_;
wire _5_;
wire _6_;
wire _7_;
wire _8_;
wire _9_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire _30_;
wire _31_;
wire _32_;
wire _33_;
wire _34_;
wire _35_;
wire _36_;
wire _37_;
wire _38_;
wire _39_;
wire _40_;
wire _41_;
wire _42_;
wire _43_;
wire _44_;
wire _45_;
wire _46_;
wire _47_;
wire _48_;
wire _49_;
wire _50_;
wire _51_;
wire _52_;
wire _53_;
wire _54_;
wire _55_;
wire _56_;
wire _57_;
wire _58_;
wire _59_;
wire _60_;
wire _61_;
wire _62_;
wire _63_;
wire _64_;
wire _65_;
wire _66_;
wire _67_;
wire _68_;
wire _69_;
wire _70_;
wire _71_;
wire _72_;
wire _73_;
wire _74_;
wire _75_;
wire _76_;
wire _77_;
wire _78_;
wire _79_;
wire _80_;
wire _81_;
wire _82_;
wire _83_;
wire _84_;
wire _85_;
wire _86_;
wire _87_;
wire _88_;
wire _89_;
wire _90_;
wire _91_;
wire _92_;
wire _93_;
wire _94_;
wire _95_;
wire _96_;
wire _97_;
wire _98_;
wire _99_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
wire _255_;
wire _256_;
wire _257_;
wire _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire _267_;
wire _268_;
wire _269_;
wire _270_;
wire _271_;
wire _272_;
wire _273_;
wire _274_;
wire _275_;
wire _276_;
wire _277_;
wire _278_;
wire _279_;
wire _280_;
wire _281_;
wire _282_;
wire _283_;
wire _284_;
wire _285_;
wire _286_;
wire _287_;
wire _288_;
wire _289_;
wire _290_;
wire _291_;
wire _292_;
wire _293_;
wire _294_;
wire _295_;
wire _296_;
wire _297_;
wire _298_;
wire _299_;
wire _300_;
wire _301_;
wire _302_;
wire _303_;
wire _304_;
wire _305_;
wire _306_;
wire _307_;
wire _308_;
wire _309_;
wire _310_;
wire _311_;
wire _312_;
wire _313_;
wire _314_;
wire _315_;
wire _316_;
wire _317_;
wire _318_;
wire _319_;
wire _320_;
wire _321_;
wire _322_;
wire _323_;
wire _324_;
wire _325_;
wire _326_;
wire _327_;
wire _328_;
wire _329_;
wire _330_;
wire _331_;
wire _332_;
wire _333_;
wire _334_;
wire _335_;
wire _336_;
wire _337_;
wire _338_;
wire _339_;
wire _340_;
wire _341_;
wire _342_;
wire _343_;
wire _344_;
wire _345_;
wire _346_;
wire _347_;
wire _348_;
wire _349_;
wire _350_;
wire _351_;
wire _352_;
wire _353_;
wire _354_;
wire _355_;
wire _356_;
wire _357_;
wire _358_;
wire _359_;
wire _360_;
wire _361_;
wire _362_;
wire _363_;
wire _364_;
wire _365_;
wire _366_;
wire _367_;
wire _368_;
wire _369_;
wire _370_;
wire _371_;
wire _372_;
wire _373_;
wire _374_;
wire _375_;
wire _376_;
wire _377_;
wire _378_;
wire _379_;
wire _380_;
wire _381_;
wire _382_;
wire _383_;
wire _384_;
wire _385_;
wire _386_;
wire _387_;
wire _388_;
wire _389_;
wire _390_;
wire _391_;
wire _392_;
wire _393_;
wire _394_;
wire _395_;
wire _396_;
wire _397_;
wire _398_;
wire _399_;
wire _400_;
wire _401_;
wire _402_;
wire _403_;
wire _404_;
wire _405_;
wire _406_;
wire _407_;
wire _408_;
wire _409_;
wire _410_;
wire _411_;
wire _412_;
wire _413_;
wire _414_;
wire _415_;
wire _416_;
wire _417_;
wire _418_;
wire _419_;
wire _420_;
wire _421_;
wire _422_;
wire _423_;
wire _424_;
wire _425_;
wire _426_;
wire _427_;
wire _428_;
wire _429_;
wire _430_;
wire _431_;
wire _432_;
wire _433_;
wire _434_;
wire _435_;
wire _436_;
wire _437_;
wire _438_;
wire _439_;
wire _440_;
wire _441_;
wire zeroWire;
wire oneWire;
assign zeroWire = 1'b0 /*506*/;
assign oneWire = 1'b1 /*506*/;
assign _9_ = ~D[0] /*480*/;
assign _6_ = R_0[3] & _9_ /*476*/;
assign _7_ = R_0[3] ^ _9_ /*479*/;
assign _8_ = oneWire & _7_ /*477*/;
assign _0_ = oneWire ^ _7_ /*478*/;
assign _5_ = _6_ | _8_ /*475*/;
assign _14_ = ~D[1] /*474*/;
assign _11_ = R_0[4] & _14_ /*470*/;
assign _12_ = R_0[4] ^ _14_ /*473*/;
assign _13_ = _5_ & _12_ /*471*/;
assign _1_ = _5_ ^ _12_ /*472*/;
assign _10_ = _11_ | _13_ /*469*/;
assign _19_ = ~D[2] /*468*/;
assign _16_ = R_0[5] & _19_ /*464*/;
assign _17_ = R_0[5] ^ _19_ /*467*/;
assign _18_ = _10_ & _17_ /*465*/;
assign _2_ = _10_ ^ _17_ /*466*/;
assign _15_ = _16_ | _18_ /*463*/;
assign _20_ = zeroWire & oneWire /*458*/;
assign _21_ = zeroWire ^ oneWire /*461*/;
assign _22_ = _15_ & _21_ /*459*/;
assign _3_ = _15_ ^ _21_ /*460*/;
assign Q[3] = _20_ | _22_ /*457*/;
assign _31_ = ~Q[3] /*433*/;
assign _30_ = _31_ & D[0] /*432*/;
assign _33_ = _0_ & _30_ /*427*/;
assign _34_ = _0_ ^ _30_ /*430*/;
assign _35_ = zeroWire & _34_ /*428*/;
assign _25_ = zeroWire ^ _34_ /*429*/;
assign _32_ = _33_ | _35_ /*426*/;
assign _37_ = ~Q[3] /*425*/;
assign _36_ = _37_ & D[1] /*424*/;
assign _39_ = _1_ & _36_ /*419*/;
assign _40_ = _1_ ^ _36_ /*422*/;
assign _41_ = _32_ & _40_ /*420*/;
assign _26_ = _32_ ^ _40_ /*421*/;
assign _38_ = _39_ | _41_ /*418*/;
assign _43_ = ~Q[3] /*417*/;
assign _42_ = _43_ & D[2] /*416*/;
assign _45_ = _2_ & _42_ /*411*/;
assign _46_ = _2_ ^ _42_ /*414*/;
assign _47_ = _38_ & _46_ /*412*/;
assign _27_ = _38_ ^ _46_ /*413*/;
assign _44_ = _45_ | _47_ /*410*/;
assign _49_ = ~Q[3] /*409*/;
assign _48_ = _49_ & zeroWire /*408*/;
assign _50_ = _3_ ^ _48_ /*406*/;
assign _28_ = _50_ ^ _44_ /*405*/;
assign _61_ = ~D[0] /*391*/;
assign _58_ = R_0[2] & _61_ /*387*/;
assign _59_ = R_0[2] ^ _61_ /*390*/;
assign _60_ = oneWire & _59_ /*388*/;
assign _53_ = oneWire ^ _59_ /*389*/;
assign _57_ = _58_ | _60_ /*386*/;
assign _66_ = ~D[1] /*385*/;
assign _63_ = _25_ & _66_ /*381*/;
assign _64_ = _25_ ^ _66_ /*384*/;
assign _65_ = _57_ & _64_ /*382*/;
assign _54_ = _57_ ^ _64_ /*383*/;
assign _62_ = _63_ | _65_ /*380*/;
assign _71_ = ~D[2] /*379*/;
assign _68_ = _26_ & _71_ /*375*/;
assign _69_ = _26_ ^ _71_ /*378*/;
assign _70_ = _62_ & _69_ /*376*/;
assign _55_ = _62_ ^ _69_ /*377*/;
assign _67_ = _68_ | _70_ /*374*/;
assign _72_ = _27_ & oneWire /*369*/;
assign _73_ = _27_ ^ oneWire /*372*/;
assign _74_ = _67_ & _73_ /*370*/;
assign _56_ = _67_ ^ _73_ /*371*/;
assign Q[2] = _72_ | _74_ /*368*/;
assign _87_ = ~Q[2] /*343*/;
assign _86_ = _87_ & D[0] /*342*/;
assign _89_ = _53_ & _86_ /*337*/;
assign _90_ = _53_ ^ _86_ /*340*/;
assign _91_ = zeroWire & _90_ /*338*/;
assign _81_ = zeroWire ^ _90_ /*339*/;
assign _88_ = _89_ | _91_ /*336*/;
assign _93_ = ~Q[2] /*335*/;
assign _92_ = _93_ & D[1] /*334*/;
assign _95_ = _54_ & _92_ /*329*/;
assign _96_ = _54_ ^ _92_ /*332*/;
assign _97_ = _88_ & _96_ /*330*/;
assign _82_ = _88_ ^ _96_ /*331*/;
assign _94_ = _95_ | _97_ /*328*/;
assign _99_ = ~Q[2] /*327*/;
assign _98_ = _99_ & D[2] /*326*/;
assign _101_ = _55_ & _98_ /*321*/;
assign _102_ = _55_ ^ _98_ /*324*/;
assign _103_ = _94_ & _102_ /*322*/;
assign _83_ = _94_ ^ _102_ /*323*/;
assign _100_ = _101_ | _103_ /*320*/;
assign _105_ = ~Q[2] /*319*/;
assign _104_ = _105_ & zeroWire /*318*/;
assign _106_ = _56_ ^ _104_ /*316*/;
assign _84_ = _106_ ^ _100_ /*315*/;
assign _117_ = ~D[0] /*301*/;
assign _114_ = R_0[1] & _117_ /*297*/;
assign _115_ = R_0[1] ^ _117_ /*300*/;
assign _116_ = oneWire & _115_ /*298*/;
assign _109_ = oneWire ^ _115_ /*299*/;
assign _113_ = _114_ | _116_ /*296*/;
assign _122_ = ~D[1] /*295*/;
assign _119_ = _81_ & _122_ /*291*/;
assign _120_ = _81_ ^ _122_ /*294*/;
assign _121_ = _113_ & _120_ /*292*/;
assign _110_ = _113_ ^ _120_ /*293*/;
assign _118_ = _119_ | _121_ /*290*/;
assign _127_ = ~D[2] /*289*/;
assign _124_ = _82_ & _127_ /*285*/;
assign _125_ = _82_ ^ _127_ /*288*/;
assign _126_ = _118_ & _125_ /*286*/;
assign _111_ = _118_ ^ _125_ /*287*/;
assign _123_ = _124_ | _126_ /*284*/;
assign _128_ = _83_ & oneWire /*279*/;
assign _129_ = _83_ ^ oneWire /*282*/;
assign _130_ = _123_ & _129_ /*280*/;
assign _112_ = _123_ ^ _129_ /*281*/;
assign Q[1] = _128_ | _130_ /*278*/;
assign _143_ = ~Q[1] /*253*/;
assign _142_ = _143_ & D[0] /*252*/;
assign _145_ = _109_ & _142_ /*247*/;
assign _146_ = _109_ ^ _142_ /*250*/;
assign _147_ = zeroWire & _146_ /*248*/;
assign _137_ = zeroWire ^ _146_ /*249*/;
assign _144_ = _145_ | _147_ /*246*/;
assign _149_ = ~Q[1] /*245*/;
assign _148_ = _149_ & D[1] /*244*/;
assign _151_ = _110_ & _148_ /*239*/;
assign _152_ = _110_ ^ _148_ /*242*/;
assign _153_ = _144_ & _152_ /*240*/;
assign _138_ = _144_ ^ _152_ /*241*/;
assign _150_ = _151_ | _153_ /*238*/;
assign _155_ = ~Q[1] /*237*/;
assign _154_ = _155_ & D[2] /*236*/;
assign _157_ = _111_ & _154_ /*231*/;
assign _158_ = _111_ ^ _154_ /*234*/;
assign _159_ = _150_ & _158_ /*232*/;
assign _139_ = _150_ ^ _158_ /*233*/;
assign _156_ = _157_ | _159_ /*230*/;
assign _161_ = ~Q[1] /*229*/;
assign _160_ = _161_ & zeroWire /*228*/;
assign _162_ = _112_ ^ _160_ /*226*/;
assign _140_ = _162_ ^ _156_ /*225*/;
assign _173_ = ~D[0] /*211*/;
assign _170_ = R_0[0] & _173_ /*207*/;
assign _171_ = R_0[0] ^ _173_ /*210*/;
assign _172_ = oneWire & _171_ /*208*/;
assign _165_ = oneWire ^ _171_ /*209*/;
assign _169_ = _170_ | _172_ /*206*/;
assign _178_ = ~D[1] /*205*/;
assign _175_ = _137_ & _178_ /*201*/;
assign _176_ = _137_ ^ _178_ /*204*/;
assign _177_ = _169_ & _176_ /*202*/;
assign _166_ = _169_ ^ _176_ /*203*/;
assign _174_ = _175_ | _177_ /*200*/;
assign _183_ = ~D[2] /*199*/;
assign _180_ = _138_ & _183_ /*195*/;
assign _181_ = _138_ ^ _183_ /*198*/;
assign _182_ = _174_ & _181_ /*196*/;
assign _167_ = _174_ ^ _181_ /*197*/;
assign _179_ = _180_ | _182_ /*194*/;
assign _184_ = _139_ & oneWire /*189*/;
assign _185_ = _139_ ^ oneWire /*192*/;
assign _186_ = _179_ & _185_ /*190*/;
assign _168_ = _179_ ^ _185_ /*191*/;
assign Q[0] = _184_ | _186_ /*188*/;
assign _199_ = ~Q[0] /*163*/;
assign _198_ = _199_ & D[0] /*162*/;
assign _201_ = _165_ & _198_ /*157*/;
assign _202_ = _165_ ^ _198_ /*160*/;
assign _203_ = zeroWire & _202_ /*158*/;
assign R_n1[0] = zeroWire ^ _202_ /*159*/;
assign _200_ = _201_ | _203_ /*156*/;
assign _205_ = ~Q[0] /*155*/;
assign _204_ = _205_ & D[1] /*154*/;
assign _207_ = _166_ & _204_ /*149*/;
assign _208_ = _166_ ^ _204_ /*152*/;
assign _209_ = _200_ & _208_ /*150*/;
assign R_n1[1] = _200_ ^ _208_ /*151*/;
assign _206_ = _207_ | _209_ /*148*/;
assign _211_ = ~Q[0] /*147*/;
assign _210_ = _211_ & D[2] /*146*/;
assign _213_ = _167_ & _210_ /*141*/;
assign _214_ = _167_ ^ _210_ /*144*/;
assign _215_ = _206_ & _214_ /*142*/;
assign R_n1[2] = _206_ ^ _214_ /*143*/;
assign _212_ = _213_ | _215_ /*140*/;
endmodule
