module divider(q, rout, rin, div);
  wire _0_;
  wire _1_;
  wire _2_;
  wire _3_;
  wire _4_;
  wire _5_;
  wire _6_;
  wire _7_;
  wire _8_;
  wire _9_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  wire _38_;
  wire _39_;
  wire _40_;
  wire _41_;
  wire _42_;
  wire _43_;
  wire _44_;
  wire _45_;
  wire _46_;
  wire _47_;
  wire _48_;
  wire _49_;
  wire _50_;
  wire _51_;
  wire _52_;
  wire _53_;
  wire _54_;
  wire _55_;
  wire _56_;
  wire _57_;
  wire _58_;
  wire _59_;
  wire _60_;
  wire _61_;
  wire _62_;
  wire _63_;
  wire _64_;
  wire _65_;
  wire _66_;
  wire _67_;
  wire _68_;
  wire _69_;
  wire _70_;
  wire _71_;
  wire _72_;
  wire _73_;
  wire _74_;
  wire _75_;
  wire _76_;
  wire _77_;
  wire _78_;
  wire _79_;
  wire _80_;
  wire _81_;
  wire _82_;
  wire _83_;
  wire _84_;
  wire _85_;
  wire _86_;
  wire _87_;
  wire _88_;
  wire _89_;
  wire _90_;
  wire _91_;
  wire _92_;
  wire _93_;
  wire _94_;
  wire _95_;
  wire _96_;
  wire _97_;
  wire _98_;
  wire _99_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire [6:0] r_0;
  wire [7:0] r_1;
  wire [7:0] m_1;
  wire [7:0] sum_1;
  wire [6:0] inv_1;
  wire [8:0] r_2;
  wire [8:0] m_2;
  wire [8:0] sum_2;
  wire [7:0] inv_2;
  wire [9:0] r_3;
  wire [9:0] m_3;
  wire [9:0] sum_3;
  wire [8:0] inv_3;
  wire [10:0] r_4;
  wire [10:0] m_4;
  wire [10:0] sum_4;
  wire [9:0] inv_4;
  wire zeroWire;
  wire oneWire;
  input [5:0] rin;
  input [2:0] div;
  output [3:0] q;
  output [10:0] rout;
  assign zeroWire = 1'b0 /*0*/;
  assign oneWire = 1'b1 /*0*/;
  assign r_0[0] = rin[0] /*660*/;
  assign r_0[1] = rin[1] /*659*/;
  assign r_0[2] = rin[2] /*658*/;
  assign r_0[3] = rin[3] /*657*/;
  assign r_0[4] = rin[4] /*656*/;
  assign r_0[5] = rin[5] /*655*/;
  assign r_0[6] = zeroWire /*654*/;
  assign inv_1[0] = oneWire /*504*/;
  assign inv_1[1] = oneWire /*498*/;
  assign inv_1[2] = oneWire /*492*/;
  assign inv_1[3] = ~div[0] /*486*/;
  assign inv_1[4] = ~div[1] /*480*/;
  assign inv_1[5] = ~div[2] /*474*/;
  assign inv_1[6] = oneWire /*468*/;
  assign _0_ = inv_1[0] ^ r_0[0] /*503*/;
  assign sum_1[0] = _0_ ^ oneWire /*502*/;
  assign _1_ = _0_ & oneWire /*501*/;
  assign _2_ = inv_1[0] & r_0[0] /*500*/;
  assign _3_ = _1_ | _2_ /*499*/;
  assign _4_ = inv_1[1] ^ r_0[1] /*497*/;
  assign sum_1[1] = _4_ ^ _3_ /*496*/;
  assign _5_ = _4_ & _3_ /*495*/;
  assign _6_ = inv_1[1] & r_0[1] /*494*/;
  assign _7_ = _5_ | _6_ /*493*/;
  assign _8_ = inv_1[2] ^ r_0[2] /*491*/;
  assign sum_1[2] = _8_ ^ _7_ /*490*/;
  assign _9_ = _8_ & _7_ /*489*/;
  assign _10_ = inv_1[2] & r_0[2] /*488*/;
  assign _11_ = _9_ | _10_ /*487*/;
  assign _12_ = inv_1[3] ^ r_0[3] /*485*/;
  assign sum_1[3] = _12_ ^ _11_ /*484*/;
  assign _13_ = _12_ & _11_ /*483*/;
  assign _14_ = inv_1[3] & r_0[3] /*482*/;
  assign _15_ = _13_ | _14_ /*481*/;
  assign _16_ = inv_1[4] ^ r_0[4] /*479*/;
  assign sum_1[4] = _16_ ^ _15_ /*478*/;
  assign _17_ = _16_ & _15_ /*477*/;
  assign _18_ = inv_1[4] & r_0[4] /*476*/;
  assign _19_ = _17_ | _18_ /*475*/;
  assign _20_ = inv_1[5] ^ r_0[5] /*473*/;
  assign sum_1[5] = _20_ ^ _19_ /*472*/;
  assign _21_ = _20_ & _19_ /*471*/;
  assign _22_ = inv_1[5] & r_0[5] /*470*/;
  assign _23_ = _21_ | _22_ /*469*/;
  assign _24_ = inv_1[6] ^ r_0[6] /*467*/;
  assign sum_1[6] = _24_ ^ _23_ /*466*/;
  assign _25_ = _24_ & _23_ /*465*/;
  assign _26_ = inv_1[6] & r_0[6] /*464*/;
  assign _27_ = _25_ | _26_ /*463*/;
  assign _28_ = _27_ ^ _23_ /*462*/;
  assign _29_ = ~_28_ /*461*/;
  assign _30_ = sum_1[6] & _29_ /*460*/;
  assign _31_ = _28_ & _27_ /*459*/;
  assign sum_1[7] = _31_ | _30_ /*458*/;
  assign q[3] = ~sum_1[7] /*457*/;
  assign m_1[0] = r_0[0] /*456*/;
  assign m_1[1] = r_0[1] /*455*/;
  assign m_1[2] = r_0[2] /*454*/;
  assign m_1[3] = r_0[3] /*453*/;
  assign m_1[4] = r_0[4] /*452*/;
  assign m_1[5] = r_0[5] /*451*/;
  assign m_1[6] = r_0[6] /*450*/;
  assign m_1[7] = r_0[6] /*449*/;
  assign _33_ = ~q[3] /*448*/;
  assign _34_ = sum_1[0] & q[3] /*447*/;
  assign _35_ = m_1[0] & _33_ /*446*/;
  assign r_1[0] = _35_ | _34_ /*445*/;
  assign _36_ = ~q[3] /*444*/;
  assign _37_ = sum_1[1] & q[3] /*443*/;
  assign _38_ = m_1[1] & _36_ /*442*/;
  assign r_1[1] = _38_ | _37_ /*441*/;
  assign _39_ = ~q[3] /*440*/;
  assign _40_ = sum_1[2] & q[3] /*439*/;
  assign _41_ = m_1[2] & _39_ /*438*/;
  assign r_1[2] = _41_ | _40_ /*437*/;
  assign _42_ = ~q[3] /*436*/;
  assign _43_ = sum_1[3] & q[3] /*435*/;
  assign _44_ = m_1[3] & _42_ /*434*/;
  assign r_1[3] = _44_ | _43_ /*433*/;
  assign _45_ = ~q[3] /*432*/;
  assign _46_ = sum_1[4] & q[3] /*431*/;
  assign _47_ = m_1[4] & _45_ /*430*/;
  assign r_1[4] = _47_ | _46_ /*429*/;
  assign _48_ = ~q[3] /*428*/;
  assign _49_ = sum_1[5] & q[3] /*427*/;
  assign _50_ = m_1[5] & _48_ /*426*/;
  assign r_1[5] = _50_ | _49_ /*425*/;
  assign _51_ = ~q[3] /*424*/;
  assign _52_ = sum_1[6] & q[3] /*423*/;
  assign _53_ = m_1[6] & _51_ /*422*/;
  assign r_1[6] = _53_ | _52_ /*421*/;
  assign _54_ = ~q[3] /*420*/;
  assign _55_ = sum_1[7] & q[3] /*419*/;
  assign _56_ = m_1[7] & _54_ /*418*/;
  assign r_1[7] = _56_ | _55_ /*417*/;
  assign inv_2[0] = oneWire /*380*/;
  assign inv_2[1] = oneWire /*374*/;
  assign inv_2[2] = ~div[0] /*368*/;
  assign inv_2[3] = ~div[1] /*362*/;
  assign inv_2[4] = ~div[2] /*356*/;
  assign inv_2[5] = oneWire /*350*/;
  assign inv_2[6] = oneWire /*344*/;
  assign inv_2[7] = oneWire /*338*/;
  assign _57_ = inv_2[0] ^ r_1[0] /*379*/;
  assign sum_2[0] = _57_ ^ oneWire /*378*/;
  assign _58_ = _57_ & oneWire /*377*/;
  assign _59_ = inv_2[0] & r_1[0] /*376*/;
  assign _60_ = _58_ | _59_ /*375*/;
  assign _61_ = inv_2[1] ^ r_1[1] /*373*/;
  assign sum_2[1] = _61_ ^ _60_ /*372*/;
  assign _62_ = _61_ & _60_ /*371*/;
  assign _63_ = inv_2[1] & r_1[1] /*370*/;
  assign _64_ = _62_ | _63_ /*369*/;
  assign _65_ = inv_2[2] ^ r_1[2] /*367*/;
  assign sum_2[2] = _65_ ^ _64_ /*366*/;
  assign _66_ = _65_ & _64_ /*365*/;
  assign _67_ = inv_2[2] & r_1[2] /*364*/;
  assign _68_ = _66_ | _67_ /*363*/;
  assign _69_ = inv_2[3] ^ r_1[3] /*361*/;
  assign sum_2[3] = _69_ ^ _68_ /*360*/;
  assign _70_ = _69_ & _68_ /*359*/;
  assign _71_ = inv_2[3] & r_1[3] /*358*/;
  assign _72_ = _70_ | _71_ /*357*/;
  assign _73_ = inv_2[4] ^ r_1[4] /*355*/;
  assign sum_2[4] = _73_ ^ _72_ /*354*/;
  assign _74_ = _73_ & _72_ /*353*/;
  assign _75_ = inv_2[4] & r_1[4] /*352*/;
  assign _76_ = _74_ | _75_ /*351*/;
  assign _77_ = inv_2[5] ^ r_1[5] /*349*/;
  assign sum_2[5] = _77_ ^ _76_ /*348*/;
  assign _78_ = _77_ & _76_ /*347*/;
  assign _79_ = inv_2[5] & r_1[5] /*346*/;
  assign _80_ = _78_ | _79_ /*345*/;
  assign _81_ = inv_2[6] ^ r_1[6] /*343*/;
  assign sum_2[6] = _81_ ^ _80_ /*342*/;
  assign _82_ = _81_ & _80_ /*341*/;
  assign _83_ = inv_2[6] & r_1[6] /*340*/;
  assign _84_ = _82_ | _83_ /*339*/;
  assign _85_ = inv_2[7] ^ r_1[7] /*337*/;
  assign sum_2[7] = _85_ ^ _84_ /*336*/;
  assign _86_ = _85_ & _84_ /*335*/;
  assign _87_ = inv_2[7] & r_1[7] /*334*/;
  assign _88_ = _86_ | _87_ /*333*/;
  assign _89_ = _88_ ^ _84_ /*332*/;
  assign _90_ = ~_89_ /*331*/;
  assign _91_ = sum_2[7] & _90_ /*330*/;
  assign _92_ = _89_ & _88_ /*329*/;
  assign sum_2[8] = _92_ | _91_ /*328*/;
  assign q[2] = ~sum_2[8] /*327*/;
  assign m_2[0] = r_1[0] /*326*/;
  assign m_2[1] = r_1[1] /*325*/;
  assign m_2[2] = r_1[2] /*324*/;
  assign m_2[3] = r_1[3] /*323*/;
  assign m_2[4] = r_1[4] /*322*/;
  assign m_2[5] = r_1[5] /*321*/;
  assign m_2[6] = r_1[6] /*320*/;
  assign m_2[7] = r_1[7] /*319*/;
  assign m_2[8] = r_1[7] /*318*/;
  assign _94_ = ~q[2] /*317*/;
  assign _95_ = sum_2[0] & q[2] /*316*/;
  assign _96_ = m_2[0] & _94_ /*315*/;
  assign r_2[0] = _96_ | _95_ /*314*/;
  assign _97_ = ~q[2] /*313*/;
  assign _98_ = sum_2[1] & q[2] /*312*/;
  assign _99_ = m_2[1] & _97_ /*311*/;
  assign r_2[1] = _99_ | _98_ /*310*/;
  assign _100_ = ~q[2] /*309*/;
  assign _101_ = sum_2[2] & q[2] /*308*/;
  assign _102_ = m_2[2] & _100_ /*307*/;
  assign r_2[2] = _102_ | _101_ /*306*/;
  assign _103_ = ~q[2] /*305*/;
  assign _104_ = sum_2[3] & q[2] /*304*/;
  assign _105_ = m_2[3] & _103_ /*303*/;
  assign r_2[3] = _105_ | _104_ /*302*/;
  assign _106_ = ~q[2] /*301*/;
  assign _107_ = sum_2[4] & q[2] /*300*/;
  assign _108_ = m_2[4] & _106_ /*299*/;
  assign r_2[4] = _108_ | _107_ /*298*/;
  assign _109_ = ~q[2] /*297*/;
  assign _110_ = sum_2[5] & q[2] /*296*/;
  assign _111_ = m_2[5] & _109_ /*295*/;
  assign r_2[5] = _111_ | _110_ /*294*/;
  assign _112_ = ~q[2] /*293*/;
  assign _113_ = sum_2[6] & q[2] /*292*/;
  assign _114_ = m_2[6] & _112_ /*291*/;
  assign r_2[6] = _114_ | _113_ /*290*/;
  assign _115_ = ~q[2] /*289*/;
  assign _116_ = sum_2[7] & q[2] /*288*/;
  assign _117_ = m_2[7] & _115_ /*287*/;
  assign r_2[7] = _117_ | _116_ /*286*/;
  assign _118_ = ~q[2] /*285*/;
  assign _119_ = sum_2[8] & q[2] /*284*/;
  assign _120_ = m_2[8] & _118_ /*283*/;
  assign r_2[8] = _120_ | _119_ /*282*/;
  assign inv_3[0] = oneWire /*256*/;
  assign inv_3[1] = ~div[0] /*250*/;
  assign inv_3[2] = ~div[1] /*244*/;
  assign inv_3[3] = ~div[2] /*238*/;
  assign inv_3[4] = oneWire /*232*/;
  assign inv_3[5] = oneWire /*226*/;
  assign inv_3[6] = oneWire /*220*/;
  assign inv_3[7] = oneWire /*214*/;
  assign inv_3[8] = oneWire /*208*/;
  assign _121_ = inv_3[0] ^ r_2[0] /*255*/;
  assign sum_3[0] = _121_ ^ oneWire /*254*/;
  assign _122_ = _121_ & oneWire /*253*/;
  assign _123_ = inv_3[0] & r_2[0] /*252*/;
  assign _124_ = _122_ | _123_ /*251*/;
  assign _125_ = inv_3[1] ^ r_2[1] /*249*/;
  assign sum_3[1] = _125_ ^ _124_ /*248*/;
  assign _126_ = _125_ & _124_ /*247*/;
  assign _127_ = inv_3[1] & r_2[1] /*246*/;
  assign _128_ = _126_ | _127_ /*245*/;
  assign _129_ = inv_3[2] ^ r_2[2] /*243*/;
  assign sum_3[2] = _129_ ^ _128_ /*242*/;
  assign _130_ = _129_ & _128_ /*241*/;
  assign _131_ = inv_3[2] & r_2[2] /*240*/;
  assign _132_ = _130_ | _131_ /*239*/;
  assign _133_ = inv_3[3] ^ r_2[3] /*237*/;
  assign sum_3[3] = _133_ ^ _132_ /*236*/;
  assign _134_ = _133_ & _132_ /*235*/;
  assign _135_ = inv_3[3] & r_2[3] /*234*/;
  assign _136_ = _134_ | _135_ /*233*/;
  assign _137_ = inv_3[4] ^ r_2[4] /*231*/;
  assign sum_3[4] = _137_ ^ _136_ /*230*/;
  assign _138_ = _137_ & _136_ /*229*/;
  assign _139_ = inv_3[4] & r_2[4] /*228*/;
  assign _140_ = _138_ | _139_ /*227*/;
  assign _141_ = inv_3[5] ^ r_2[5] /*225*/;
  assign sum_3[5] = _141_ ^ _140_ /*224*/;
  assign _142_ = _141_ & _140_ /*223*/;
  assign _143_ = inv_3[5] & r_2[5] /*222*/;
  assign _144_ = _142_ | _143_ /*221*/;
  assign _145_ = inv_3[6] ^ r_2[6] /*219*/;
  assign sum_3[6] = _145_ ^ _144_ /*218*/;
  assign _146_ = _145_ & _144_ /*217*/;
  assign _147_ = inv_3[6] & r_2[6] /*216*/;
  assign _148_ = _146_ | _147_ /*215*/;
  assign _149_ = inv_3[7] ^ r_2[7] /*213*/;
  assign sum_3[7] = _149_ ^ _148_ /*212*/;
  assign _150_ = _149_ & _148_ /*211*/;
  assign _151_ = inv_3[7] & r_2[7] /*210*/;
  assign _152_ = _150_ | _151_ /*209*/;
  assign _153_ = inv_3[8] ^ r_2[8] /*207*/;
  assign sum_3[8] = _153_ ^ _152_ /*206*/;
  assign _154_ = _153_ & _152_ /*205*/;
  assign _155_ = inv_3[8] & r_2[8] /*204*/;
  assign _156_ = _154_ | _155_ /*203*/;
  assign _157_ = _156_ ^ _152_ /*202*/;
  assign _158_ = ~_157_ /*201*/;
  assign _159_ = sum_3[8] & _158_ /*200*/;
  assign _160_ = _157_ & _156_ /*199*/;
  assign sum_3[9] = _160_ | _159_ /*198*/;
  assign q[1] = ~sum_3[9] /*197*/;
  assign m_3[0] = r_2[0] /*196*/;
  assign m_3[1] = r_2[1] /*195*/;
  assign m_3[2] = r_2[2] /*194*/;
  assign m_3[3] = r_2[3] /*193*/;
  assign m_3[4] = r_2[4] /*192*/;
  assign m_3[5] = r_2[5] /*191*/;
  assign m_3[6] = r_2[6] /*190*/;
  assign m_3[7] = r_2[7] /*189*/;
  assign m_3[8] = r_2[8] /*188*/;
  assign m_3[9] = r_2[8] /*187*/;
  assign _162_ = ~q[1] /*186*/;
  assign _163_ = sum_3[0] & q[1] /*185*/;
  assign _164_ = m_3[0] & _162_ /*184*/;
  assign r_3[0] = _164_ | _163_ /*183*/;
  assign _165_ = ~q[1] /*182*/;
  assign _166_ = sum_3[1] & q[1] /*181*/;
  assign _167_ = m_3[1] & _165_ /*180*/;
  assign r_3[1] = _167_ | _166_ /*179*/;
  assign _168_ = ~q[1] /*178*/;
  assign _169_ = sum_3[2] & q[1] /*177*/;
  assign _170_ = m_3[2] & _168_ /*176*/;
  assign r_3[2] = _170_ | _169_ /*175*/;
  assign _171_ = ~q[1] /*174*/;
  assign _172_ = sum_3[3] & q[1] /*173*/;
  assign _173_ = m_3[3] & _171_ /*172*/;
  assign r_3[3] = _173_ | _172_ /*171*/;
  assign _174_ = ~q[1] /*170*/;
  assign _175_ = sum_3[4] & q[1] /*169*/;
  assign _176_ = m_3[4] & _174_ /*168*/;
  assign r_3[4] = _176_ | _175_ /*167*/;
  assign _177_ = ~q[1] /*166*/;
  assign _178_ = sum_3[5] & q[1] /*165*/;
  assign _179_ = m_3[5] & _177_ /*164*/;
  assign r_3[5] = _179_ | _178_ /*163*/;
  assign _180_ = ~q[1] /*162*/;
  assign _181_ = sum_3[6] & q[1] /*161*/;
  assign _182_ = m_3[6] & _180_ /*160*/;
  assign r_3[6] = _182_ | _181_ /*159*/;
  assign _183_ = ~q[1] /*158*/;
  assign _184_ = sum_3[7] & q[1] /*157*/;
  assign _185_ = m_3[7] & _183_ /*156*/;
  assign r_3[7] = _185_ | _184_ /*155*/;
  assign _186_ = ~q[1] /*154*/;
  assign _187_ = sum_3[8] & q[1] /*153*/;
  assign _188_ = m_3[8] & _186_ /*152*/;
  assign r_3[8] = _188_ | _187_ /*151*/;
  assign _189_ = ~q[1] /*150*/;
  assign _190_ = sum_3[9] & q[1] /*149*/;
  assign _191_ = m_3[9] & _189_ /*148*/;
  assign r_3[9] = _191_ | _190_ /*147*/;
  assign inv_4[0] = ~div[0] /*132*/;
  assign inv_4[1] = ~div[1] /*126*/;
  assign inv_4[2] = ~div[2] /*120*/;
  assign inv_4[3] = oneWire /*114*/;
  assign inv_4[4] = oneWire /*108*/;
  assign inv_4[5] = oneWire /*102*/;
  assign inv_4[6] = oneWire /*96*/;
  assign inv_4[7] = oneWire /*90*/;
  assign inv_4[8] = oneWire /*84*/;
  assign inv_4[9] = oneWire /*78*/;
  assign _192_ = inv_4[0] ^ r_3[0] /*131*/;
  assign sum_4[0] = _192_ ^ oneWire /*130*/;
  assign _193_ = _192_ & oneWire /*129*/;
  assign _194_ = inv_4[0] & r_3[0] /*128*/;
  assign _195_ = _193_ | _194_ /*127*/;
  assign _196_ = inv_4[1] ^ r_3[1] /*125*/;
  assign sum_4[1] = _196_ ^ _195_ /*124*/;
  assign _197_ = _196_ & _195_ /*123*/;
  assign _198_ = inv_4[1] & r_3[1] /*122*/;
  assign _199_ = _197_ | _198_ /*121*/;
  assign _200_ = inv_4[2] ^ r_3[2] /*119*/;
  assign sum_4[2] = _200_ ^ _199_ /*118*/;
  assign _201_ = _200_ & _199_ /*117*/;
  assign _202_ = inv_4[2] & r_3[2] /*116*/;
  assign _203_ = _201_ | _202_ /*115*/;
  assign _204_ = inv_4[3] ^ r_3[3] /*113*/;
  assign sum_4[3] = _204_ ^ _203_ /*112*/;
  assign _205_ = _204_ & _203_ /*111*/;
  assign _206_ = inv_4[3] & r_3[3] /*110*/;
  assign _207_ = _205_ | _206_ /*109*/;
  assign _208_ = inv_4[4] ^ r_3[4] /*107*/;
  assign sum_4[4] = _208_ ^ _207_ /*106*/;
  assign _209_ = _208_ & _207_ /*105*/;
  assign _210_ = inv_4[4] & r_3[4] /*104*/;
  assign _211_ = _209_ | _210_ /*103*/;
  assign _212_ = inv_4[5] ^ r_3[5] /*101*/;
  assign sum_4[5] = _212_ ^ _211_ /*100*/;
  assign _213_ = _212_ & _211_ /*99*/;
  assign _214_ = inv_4[5] & r_3[5] /*98*/;
  assign _215_ = _213_ | _214_ /*97*/;
  assign _216_ = inv_4[6] ^ r_3[6] /*95*/;
  assign sum_4[6] = _216_ ^ _215_ /*94*/;
  assign _217_ = _216_ & _215_ /*93*/;
  assign _218_ = inv_4[6] & r_3[6] /*92*/;
  assign _219_ = _217_ | _218_ /*91*/;
  assign _220_ = inv_4[7] ^ r_3[7] /*89*/;
  assign sum_4[7] = _220_ ^ _219_ /*88*/;
  assign _221_ = _220_ & _219_ /*87*/;
  assign _222_ = inv_4[7] & r_3[7] /*86*/;
  assign _223_ = _221_ | _222_ /*85*/;
  assign _224_ = inv_4[8] ^ r_3[8] /*83*/;
  assign sum_4[8] = _224_ ^ _223_ /*82*/;
  assign _225_ = _224_ & _223_ /*81*/;
  assign _226_ = inv_4[8] & r_3[8] /*80*/;
  assign _227_ = _225_ | _226_ /*79*/;
  assign _228_ = inv_4[9] ^ r_3[9] /*77*/;
  assign sum_4[9] = _228_ ^ _227_ /*76*/;
  assign _229_ = _228_ & _227_ /*75*/;
  assign _230_ = inv_4[9] & r_3[9] /*74*/;
  assign _231_ = _229_ | _230_ /*73*/;
  assign _232_ = _231_ ^ _227_ /*72*/;
  assign _233_ = ~_232_ /*71*/;
  assign _234_ = sum_4[9] & _233_ /*70*/;
  assign _235_ = _232_ & _231_ /*69*/;
  assign sum_4[10] = _235_ | _234_ /*68*/;
  assign q[0] = ~sum_4[10] /*67*/;
  assign m_4[0] = r_3[0] /*66*/;
  assign m_4[1] = r_3[1] /*65*/;
  assign m_4[2] = r_3[2] /*64*/;
  assign m_4[3] = r_3[3] /*63*/;
  assign m_4[4] = r_3[4] /*62*/;
  assign m_4[5] = r_3[5] /*61*/;
  assign m_4[6] = r_3[6] /*60*/;
  assign m_4[7] = r_3[7] /*59*/;
  assign m_4[8] = r_3[8] /*58*/;
  assign m_4[9] = r_3[9] /*57*/;
  assign m_4[10] = r_3[9] /*56*/;
  assign _237_ = ~q[0] /*55*/;
  assign _238_ = sum_4[0] & q[0] /*54*/;
  assign _239_ = m_4[0] & _237_ /*53*/;
  assign r_4[0] = _239_ | _238_ /*52*/;
  assign _240_ = ~q[0] /*51*/;
  assign _241_ = sum_4[1] & q[0] /*50*/;
  assign _242_ = m_4[1] & _240_ /*49*/;
  assign r_4[1] = _242_ | _241_ /*48*/;
  assign _243_ = ~q[0] /*47*/;
  assign _244_ = sum_4[2] & q[0] /*46*/;
  assign _245_ = m_4[2] & _243_ /*45*/;
  assign r_4[2] = _245_ | _244_ /*44*/;
  assign _246_ = ~q[0] /*43*/;
  assign _247_ = sum_4[3] & q[0] /*42*/;
  assign _248_ = m_4[3] & _246_ /*41*/;
  assign r_4[3] = _248_ | _247_ /*40*/;
  assign _249_ = ~q[0] /*39*/;
  assign _250_ = sum_4[4] & q[0] /*38*/;
  assign _251_ = m_4[4] & _249_ /*37*/;
  assign r_4[4] = _251_ | _250_ /*36*/;
  assign _252_ = ~q[0] /*35*/;
  assign _253_ = sum_4[5] & q[0] /*34*/;
  assign _254_ = m_4[5] & _252_ /*33*/;
  assign r_4[5] = _254_ | _253_ /*32*/;
  assign _255_ = ~q[0] /*31*/;
  assign _256_ = sum_4[6] & q[0] /*30*/;
  assign _257_ = m_4[6] & _255_ /*29*/;
  assign r_4[6] = _257_ | _256_ /*28*/;
  assign _258_ = ~q[0] /*27*/;
  assign _259_ = sum_4[7] & q[0] /*26*/;
  assign _260_ = m_4[7] & _258_ /*25*/;
  assign r_4[7] = _260_ | _259_ /*24*/;
  assign _261_ = ~q[0] /*23*/;
  assign _262_ = sum_4[8] & q[0] /*22*/;
  assign _263_ = m_4[8] & _261_ /*21*/;
  assign r_4[8] = _263_ | _262_ /*20*/;
  assign _264_ = ~q[0] /*19*/;
  assign _265_ = sum_4[9] & q[0] /*18*/;
  assign _266_ = m_4[9] & _264_ /*17*/;
  assign r_4[9] = _266_ | _265_ /*16*/;
  assign _267_ = ~q[0] /*15*/;
  assign _268_ = sum_4[10] & q[0] /*14*/;
  assign _269_ = m_4[10] & _267_ /*13*/;
  assign r_4[10] = _269_ | _268_ /*12*/;
  assign rout[0] = r_4[0] /*0*/;
  assign rout[1] = r_4[1] /*1*/;
  assign rout[2] = r_4[2] /*2*/;
  assign rout[3] = r_4[3] /*3*/;
  assign rout[4] = r_4[4] /*4*/;
  assign rout[5] = r_4[5] /*5*/;
  assign rout[6] = r_4[6] /*6*/;
  assign rout[7] = r_4[7] /*7*/;
  assign rout[8] = r_4[8] /*8*/;
  assign rout[9] = r_4[9] /*9*/;
  assign rout[10] = r_4[10] /*10*/;
endmodule