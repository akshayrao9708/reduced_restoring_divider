module divider(q, rout, rin, div);
  wire _0_;
  wire _1_;
  wire _2_;
  wire _3_;
  wire _4_;
  wire _5_;
  wire _6_;
  wire _7_;
  wire _8_;
  wire _9_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  wire _38_;
  wire _39_;
  wire _40_;
  wire _41_;
  wire _42_;
  wire _43_;
  wire _44_;
  wire _45_;
  wire _46_;
  wire _47_;
  wire _48_;
  wire _49_;
  wire _50_;
  wire _51_;
  wire _52_;
  wire _53_;
  wire _54_;
  wire _55_;
  wire _56_;
  wire _57_;
  wire _58_;
  wire _59_;
  wire _60_;
  wire _61_;
  wire _62_;
  wire _63_;
  wire _64_;
  wire _65_;
  wire _66_;
  wire _67_;
  wire _68_;
  wire _69_;
  wire _70_;
  wire _71_;
  wire _72_;
  wire _73_;
  wire _74_;
  wire _75_;
  wire _76_;
  wire _77_;
  wire _78_;
  wire _79_;
  wire _80_;
  wire _81_;
  wire _82_;
  wire _83_;
  wire _84_;
  wire _85_;
  wire _86_;
  wire _87_;
  wire _88_;
  wire _89_;
  wire _90_;
  wire _91_;
  wire _92_;
  wire _93_;
  wire _94_;
  wire _95_;
  wire _96_;
  wire _97_;
  wire _98_;
  wire _99_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire [4:0] r_0;
  wire [5:0] r_1;
  wire [5:0] m_1;
  wire [5:0] sum_1;
  wire [4:0] inv_1;
  wire [6:0] r_2;
  wire [6:0] m_2;
  wire [6:0] sum_2;
  wire [5:0] inv_2;
  wire [7:0] r_3;
  wire [7:0] m_3;
  wire [7:0] sum_3;
  wire [6:0] inv_3;
  wire zeroWire;
  wire oneWire;
  input [3:0] rin;
  input [1:0] div;
  output [2:0] q;
  output [7:0] rout;
  assign zeroWire = 1'b0 /*0*/;
  assign oneWire = 1'b1 /*0*/;
  assign r_0[0] = rin[0] /*393*/;
  assign r_0[1] = rin[1] /*392*/;
  assign r_0[2] = rin[2] /*391*/;
  assign r_0[3] = rin[3] /*390*/;
  assign r_0[4] = zeroWire /*389*/;
  assign inv_1[0] = oneWire /*276*/;
  assign inv_1[1] = oneWire /*270*/;
  assign inv_1[2] = ~div[0] /*264*/;
  assign inv_1[3] = ~div[1] /*258*/;
  assign inv_1[4] = oneWire /*252*/;
  assign _0_ = inv_1[0] ^ r_0[0] /*275*/;
  assign sum_1[0] = _0_ ^ oneWire /*274*/;
  assign _1_ = _0_ & oneWire /*273*/;
  assign _2_ = inv_1[0] & r_0[0] /*272*/;
  assign _3_ = _1_ | _2_ /*271*/;
  assign _4_ = inv_1[1] ^ r_0[1] /*269*/;
  assign sum_1[1] = _4_ ^ _3_ /*268*/;
  assign _5_ = _4_ & _3_ /*267*/;
  assign _6_ = inv_1[1] & r_0[1] /*266*/;
  assign _7_ = _5_ | _6_ /*265*/;
  assign _8_ = inv_1[2] ^ r_0[2] /*263*/;
  assign sum_1[2] = _8_ ^ _7_ /*262*/;
  assign _9_ = _8_ & _7_ /*261*/;
  assign _10_ = inv_1[2] & r_0[2] /*260*/;
  assign _11_ = _9_ | _10_ /*259*/;
  assign _12_ = inv_1[3] ^ r_0[3] /*257*/;
  assign sum_1[3] = _12_ ^ _11_ /*256*/;
  assign _13_ = _12_ & _11_ /*255*/;
  assign _14_ = inv_1[3] & r_0[3] /*254*/;
  assign _15_ = _13_ | _14_ /*253*/;
  assign _16_ = inv_1[4] ^ r_0[4] /*251*/;
  assign sum_1[4] = _16_ ^ _15_ /*250*/;
  assign _17_ = _16_ & _15_ /*249*/;
  assign _18_ = inv_1[4] & r_0[4] /*248*/;
  assign _19_ = _17_ | _18_ /*247*/;
  assign _20_ = _19_ ^ _15_ /*246*/;
  assign _21_ = ~_20_ /*245*/;
  assign _22_ = sum_1[4] & _21_ /*244*/;
  assign _23_ = _20_ & _19_ /*243*/;
  assign sum_1[5] = _23_ | _22_ /*242*/;
  assign q[2] = ~sum_1[5] /*241*/;
  assign m_1[0] = r_0[0] /*240*/;
  assign m_1[1] = r_0[1] /*239*/;
  assign m_1[2] = r_0[2] /*238*/;
  assign m_1[3] = r_0[3] /*237*/;
  assign m_1[4] = r_0[4] /*236*/;
  assign m_1[5] = r_0[4] /*235*/;
  assign _25_ = ~q[2] /*234*/;
  assign _26_ = sum_1[0] & q[2] /*233*/;
  assign _27_ = m_1[0] & _25_ /*232*/;
  assign r_1[0] = _27_ | _26_ /*231*/;
  assign _28_ = ~q[2] /*230*/;
  assign _29_ = sum_1[1] & q[2] /*229*/;
  assign _30_ = m_1[1] & _28_ /*228*/;
  assign r_1[1] = _30_ | _29_ /*227*/;
  assign _31_ = ~q[2] /*226*/;
  assign _32_ = sum_1[2] & q[2] /*225*/;
  assign _33_ = m_1[2] & _31_ /*224*/;
  assign r_1[2] = _33_ | _32_ /*223*/;
  assign _34_ = ~q[2] /*222*/;
  assign _35_ = sum_1[3] & q[2] /*221*/;
  assign _36_ = m_1[3] & _34_ /*220*/;
  assign r_1[3] = _36_ | _35_ /*219*/;
  assign _37_ = ~q[2] /*218*/;
  assign _38_ = sum_1[4] & q[2] /*217*/;
  assign _39_ = m_1[4] & _37_ /*216*/;
  assign r_1[4] = _39_ | _38_ /*215*/;
  assign _40_ = ~q[2] /*214*/;
  assign _41_ = sum_1[5] & q[2] /*213*/;
  assign _42_ = m_1[5] & _40_ /*212*/;
  assign r_1[5] = _42_ | _41_ /*211*/;
  assign inv_2[0] = oneWire /*186*/;
  assign inv_2[1] = ~div[0] /*180*/;
  assign inv_2[2] = ~div[1] /*174*/;
  assign inv_2[3] = oneWire /*168*/;
  assign inv_2[4] = oneWire /*162*/;
  assign inv_2[5] = oneWire /*156*/;
  assign _43_ = inv_2[0] ^ r_1[0] /*185*/;
  assign sum_2[0] = _43_ ^ oneWire /*184*/;
  assign _44_ = _43_ & oneWire /*183*/;
  assign _45_ = inv_2[0] & r_1[0] /*182*/;
  assign _46_ = _44_ | _45_ /*181*/;
  assign _47_ = inv_2[1] ^ r_1[1] /*179*/;
  assign sum_2[1] = _47_ ^ _46_ /*178*/;
  assign _48_ = _47_ & _46_ /*177*/;
  assign _49_ = inv_2[1] & r_1[1] /*176*/;
  assign _50_ = _48_ | _49_ /*175*/;
  assign _51_ = inv_2[2] ^ r_1[2] /*173*/;
  assign sum_2[2] = _51_ ^ _50_ /*172*/;
  assign _52_ = _51_ & _50_ /*171*/;
  assign _53_ = inv_2[2] & r_1[2] /*170*/;
  assign _54_ = _52_ | _53_ /*169*/;
  assign _55_ = inv_2[3] ^ r_1[3] /*167*/;
  assign sum_2[3] = _55_ ^ _54_ /*166*/;
  assign _56_ = _55_ & _54_ /*165*/;
  assign _57_ = inv_2[3] & r_1[3] /*164*/;
  assign _58_ = _56_ | _57_ /*163*/;
  assign _59_ = inv_2[4] ^ r_1[4] /*161*/;
  assign sum_2[4] = _59_ ^ _58_ /*160*/;
  assign _60_ = _59_ & _58_ /*159*/;
  assign _61_ = inv_2[4] & r_1[4] /*158*/;
  assign _62_ = _60_ | _61_ /*157*/;
  assign _63_ = inv_2[5] ^ r_1[5] /*155*/;
  assign sum_2[5] = _63_ ^ _62_ /*154*/;
  assign _64_ = _63_ & _62_ /*153*/;
  assign _65_ = inv_2[5] & r_1[5] /*152*/;
  assign _66_ = _64_ | _65_ /*151*/;
  assign _67_ = _66_ ^ _62_ /*150*/;
  assign _68_ = ~_67_ /*149*/;
  assign _69_ = sum_2[5] & _68_ /*148*/;
  assign _70_ = _67_ & _66_ /*147*/;
  assign sum_2[6] = _70_ | _69_ /*146*/;
  assign q[1] = ~sum_2[6] /*145*/;
  assign m_2[0] = r_1[0] /*144*/;
  assign m_2[1] = r_1[1] /*143*/;
  assign m_2[2] = r_1[2] /*142*/;
  assign m_2[3] = r_1[3] /*141*/;
  assign m_2[4] = r_1[4] /*140*/;
  assign m_2[5] = r_1[5] /*139*/;
  assign m_2[6] = r_1[5] /*138*/;
  assign _72_ = ~q[1] /*137*/;
  assign _73_ = sum_2[0] & q[1] /*136*/;
  assign _74_ = m_2[0] & _72_ /*135*/;
  assign r_2[0] = _74_ | _73_ /*134*/;
  assign _75_ = ~q[1] /*133*/;
  assign _76_ = sum_2[1] & q[1] /*132*/;
  assign _77_ = m_2[1] & _75_ /*131*/;
  assign r_2[1] = _77_ | _76_ /*130*/;
  assign _78_ = ~q[1] /*129*/;
  assign _79_ = sum_2[2] & q[1] /*128*/;
  assign _80_ = m_2[2] & _78_ /*127*/;
  assign r_2[2] = _80_ | _79_ /*126*/;
  assign _81_ = ~q[1] /*125*/;
  assign _82_ = sum_2[3] & q[1] /*124*/;
  assign _83_ = m_2[3] & _81_ /*123*/;
  assign r_2[3] = _83_ | _82_ /*122*/;
  assign _84_ = ~q[1] /*121*/;
  assign _85_ = sum_2[4] & q[1] /*120*/;
  assign _86_ = m_2[4] & _84_ /*119*/;
  assign r_2[4] = _86_ | _85_ /*118*/;
  assign _87_ = ~q[1] /*117*/;
  assign _88_ = sum_2[5] & q[1] /*116*/;
  assign _89_ = m_2[5] & _87_ /*115*/;
  assign r_2[5] = _89_ | _88_ /*114*/;
  assign _90_ = ~q[1] /*113*/;
  assign _91_ = sum_2[6] & q[1] /*112*/;
  assign _92_ = m_2[6] & _90_ /*111*/;
  assign r_2[6] = _92_ | _91_ /*110*/;
  assign inv_3[0] = ~div[0] /*96*/;
  assign inv_3[1] = ~div[1] /*90*/;
  assign inv_3[2] = oneWire /*84*/;
  assign inv_3[3] = oneWire /*78*/;
  assign inv_3[4] = oneWire /*72*/;
  assign inv_3[5] = oneWire /*66*/;
  assign inv_3[6] = oneWire /*60*/;
  assign _93_ = inv_3[0] ^ r_2[0] /*95*/;
  assign sum_3[0] = _93_ ^ oneWire /*94*/;
  assign _94_ = _93_ & oneWire /*93*/;
  assign _95_ = inv_3[0] & r_2[0] /*92*/;
  assign _96_ = _94_ | _95_ /*91*/;
  assign _97_ = inv_3[1] ^ r_2[1] /*89*/;
  assign sum_3[1] = _97_ ^ _96_ /*88*/;
  assign _98_ = _97_ & _96_ /*87*/;
  assign _99_ = inv_3[1] & r_2[1] /*86*/;
  assign _100_ = _98_ | _99_ /*85*/;
  assign _101_ = inv_3[2] ^ r_2[2] /*83*/;
  assign sum_3[2] = _101_ ^ _100_ /*82*/;
  assign _102_ = _101_ & _100_ /*81*/;
  assign _103_ = inv_3[2] & r_2[2] /*80*/;
  assign _104_ = _102_ | _103_ /*79*/;
  assign _105_ = inv_3[3] ^ r_2[3] /*77*/;
  assign sum_3[3] = _105_ ^ _104_ /*76*/;
  assign _106_ = _105_ & _104_ /*75*/;
  assign _107_ = inv_3[3] & r_2[3] /*74*/;
  assign _108_ = _106_ | _107_ /*73*/;
  assign _109_ = inv_3[4] ^ r_2[4] /*71*/;
  assign sum_3[4] = _109_ ^ _108_ /*70*/;
  assign _110_ = _109_ & _108_ /*69*/;
  assign _111_ = inv_3[4] & r_2[4] /*68*/;
  assign _112_ = _110_ | _111_ /*67*/;
  assign _113_ = inv_3[5] ^ r_2[5] /*65*/;
  assign sum_3[5] = _113_ ^ _112_ /*64*/;
  assign _114_ = _113_ & _112_ /*63*/;
  assign _115_ = inv_3[5] & r_2[5] /*62*/;
  assign _116_ = _114_ | _115_ /*61*/;
  assign _117_ = inv_3[6] ^ r_2[6] /*59*/;
  assign sum_3[6] = _117_ ^ _116_ /*58*/;
  assign _118_ = _117_ & _116_ /*57*/;
  assign _119_ = inv_3[6] & r_2[6] /*56*/;
  assign _120_ = _118_ | _119_ /*55*/;
  assign _121_ = _120_ ^ _116_ /*54*/;
  assign _122_ = ~_121_ /*53*/;
  assign _123_ = sum_3[6] & _122_ /*52*/;
  assign _124_ = _121_ & _120_ /*51*/;
  assign sum_3[7] = _124_ | _123_ /*50*/;
  assign q[0] = ~sum_3[7] /*49*/;
  assign m_3[0] = r_2[0] /*48*/;
  assign m_3[1] = r_2[1] /*47*/;
  assign m_3[2] = r_2[2] /*46*/;
  assign m_3[3] = r_2[3] /*45*/;
  assign m_3[4] = r_2[4] /*44*/;
  assign m_3[5] = r_2[5] /*43*/;
  assign m_3[6] = r_2[6] /*42*/;
  assign m_3[7] = r_2[6] /*41*/;
  assign _126_ = ~q[0] /*40*/;
  assign _127_ = sum_3[0] & q[0] /*39*/;
  assign _128_ = m_3[0] & _126_ /*38*/;
  assign r_3[0] = _128_ | _127_ /*37*/;
  assign _129_ = ~q[0] /*36*/;
  assign _130_ = sum_3[1] & q[0] /*35*/;
  assign _131_ = m_3[1] & _129_ /*34*/;
  assign r_3[1] = _131_ | _130_ /*33*/;
  assign _132_ = ~q[0] /*32*/;
  assign _133_ = sum_3[2] & q[0] /*31*/;
  assign _134_ = m_3[2] & _132_ /*30*/;
  assign r_3[2] = _134_ | _133_ /*29*/;
  assign _135_ = ~q[0] /*28*/;
  assign _136_ = sum_3[3] & q[0] /*27*/;
  assign _137_ = m_3[3] & _135_ /*26*/;
  assign r_3[3] = _137_ | _136_ /*25*/;
  assign _138_ = ~q[0] /*24*/;
  assign _139_ = sum_3[4] & q[0] /*23*/;
  assign _140_ = m_3[4] & _138_ /*22*/;
  assign r_3[4] = _140_ | _139_ /*21*/;
  assign _141_ = ~q[0] /*20*/;
  assign _142_ = sum_3[5] & q[0] /*19*/;
  assign _143_ = m_3[5] & _141_ /*18*/;
  assign r_3[5] = _143_ | _142_ /*17*/;
  assign _144_ = ~q[0] /*16*/;
  assign _145_ = sum_3[6] & q[0] /*15*/;
  assign _146_ = m_3[6] & _144_ /*14*/;
  assign r_3[6] = _146_ | _145_ /*13*/;
  assign _147_ = ~q[0] /*12*/;
  assign _148_ = sum_3[7] & q[0] /*11*/;
  assign _149_ = m_3[7] & _147_ /*10*/;
  assign r_3[7] = _149_ | _148_ /*9*/;
  assign rout[0] = r_3[0] /*0*/;
  assign rout[1] = r_3[1] /*1*/;
  assign rout[2] = r_3[2] /*2*/;
  assign rout[3] = r_3[3] /*3*/;
  assign rout[4] = r_3[4] /*4*/;
  assign rout[5] = r_3[5] /*5*/;
  assign rout[6] = r_3[6] /*6*/;
  assign rout[7] = r_3[7] /*7*/;
endmodule