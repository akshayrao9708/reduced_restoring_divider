module nonresdivReduced(R_0, D, Q, R_n1);
input [125:0] R_0;
input [62:0] D;
output [63:0] Q;
output [63:0] R_n1;
wire _0_;
wire _1_;
wire _2_;
wire _3_;
wire _4_;
wire _5_;
wire _6_;
wire _7_;
wire _8_;
wire _9_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire _30_;
wire _31_;
wire _32_;
wire _33_;
wire _34_;
wire _35_;
wire _36_;
wire _37_;
wire _38_;
wire _39_;
wire _40_;
wire _41_;
wire _42_;
wire _43_;
wire _44_;
wire _45_;
wire _46_;
wire _47_;
wire _48_;
wire _49_;
wire _50_;
wire _51_;
wire _52_;
wire _53_;
wire _54_;
wire _55_;
wire _56_;
wire _57_;
wire _58_;
wire _59_;
wire _60_;
wire _61_;
wire _62_;
wire _63_;
wire _64_;
wire _65_;
wire _66_;
wire _67_;
wire _68_;
wire _69_;
wire _70_;
wire _71_;
wire _72_;
wire _73_;
wire _74_;
wire _75_;
wire _76_;
wire _77_;
wire _78_;
wire _79_;
wire _80_;
wire _81_;
wire _82_;
wire _83_;
wire _84_;
wire _85_;
wire _86_;
wire _87_;
wire _88_;
wire _89_;
wire _90_;
wire _91_;
wire _92_;
wire _93_;
wire _94_;
wire _95_;
wire _96_;
wire _97_;
wire _98_;
wire _99_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
wire _255_;
wire _256_;
wire _257_;
wire _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire _267_;
wire _268_;
wire _269_;
wire _270_;
wire _271_;
wire _272_;
wire _273_;
wire _274_;
wire _275_;
wire _276_;
wire _277_;
wire _278_;
wire _279_;
wire _280_;
wire _281_;
wire _282_;
wire _283_;
wire _284_;
wire _285_;
wire _286_;
wire _287_;
wire _288_;
wire _289_;
wire _290_;
wire _291_;
wire _292_;
wire _293_;
wire _294_;
wire _295_;
wire _296_;
wire _297_;
wire _298_;
wire _299_;
wire _300_;
wire _301_;
wire _302_;
wire _303_;
wire _304_;
wire _305_;
wire _306_;
wire _307_;
wire _308_;
wire _309_;
wire _310_;
wire _311_;
wire _312_;
wire _313_;
wire _314_;
wire _315_;
wire _316_;
wire _317_;
wire _318_;
wire _319_;
wire _320_;
wire _321_;
wire _322_;
wire _323_;
wire _324_;
wire _325_;
wire _326_;
wire _327_;
wire _328_;
wire _329_;
wire _330_;
wire _331_;
wire _332_;
wire _333_;
wire _334_;
wire _335_;
wire _336_;
wire _337_;
wire _338_;
wire _339_;
wire _340_;
wire _341_;
wire _342_;
wire _343_;
wire _344_;
wire _345_;
wire _346_;
wire _347_;
wire _348_;
wire _349_;
wire _350_;
wire _351_;
wire _352_;
wire _353_;
wire _354_;
wire _355_;
wire _356_;
wire _357_;
wire _358_;
wire _359_;
wire _360_;
wire _361_;
wire _362_;
wire _363_;
wire _364_;
wire _365_;
wire _366_;
wire _367_;
wire _368_;
wire _369_;
wire _370_;
wire _371_;
wire _372_;
wire _373_;
wire _374_;
wire _375_;
wire _376_;
wire _377_;
wire _378_;
wire _379_;
wire _380_;
wire _381_;
wire _382_;
wire _383_;
wire _384_;
wire _385_;
wire _386_;
wire _387_;
wire _388_;
wire _389_;
wire _390_;
wire _391_;
wire _392_;
wire _393_;
wire _394_;
wire _395_;
wire _396_;
wire _397_;
wire _398_;
wire _399_;
wire _400_;
wire _401_;
wire _402_;
wire _403_;
wire _404_;
wire _405_;
wire _406_;
wire _407_;
wire _408_;
wire _409_;
wire _410_;
wire _411_;
wire _412_;
wire _413_;
wire _414_;
wire _415_;
wire _416_;
wire _417_;
wire _418_;
wire _419_;
wire _420_;
wire _421_;
wire _422_;
wire _423_;
wire _424_;
wire _425_;
wire _426_;
wire _427_;
wire _428_;
wire _429_;
wire _430_;
wire _431_;
wire _432_;
wire _433_;
wire _434_;
wire _435_;
wire _436_;
wire _437_;
wire _438_;
wire _439_;
wire _440_;
wire _441_;
wire _442_;
wire _443_;
wire _444_;
wire _445_;
wire _446_;
wire _447_;
wire _448_;
wire _449_;
wire _450_;
wire _451_;
wire _452_;
wire _453_;
wire _454_;
wire _455_;
wire _456_;
wire _457_;
wire _458_;
wire _459_;
wire _460_;
wire _461_;
wire _462_;
wire _463_;
wire _464_;
wire _465_;
wire _466_;
wire _467_;
wire _468_;
wire _469_;
wire _470_;
wire _471_;
wire _472_;
wire _473_;
wire _474_;
wire _475_;
wire _476_;
wire _477_;
wire _478_;
wire _479_;
wire _480_;
wire _481_;
wire _482_;
wire _483_;
wire _484_;
wire _485_;
wire _486_;
wire _487_;
wire _488_;
wire _489_;
wire _490_;
wire _491_;
wire _492_;
wire _493_;
wire _494_;
wire _495_;
wire _496_;
wire _497_;
wire _498_;
wire _499_;
wire _500_;
wire _501_;
wire _502_;
wire _503_;
wire _504_;
wire _505_;
wire _506_;
wire _507_;
wire _508_;
wire _509_;
wire _510_;
wire _511_;
wire _512_;
wire _513_;
wire _514_;
wire _515_;
wire _516_;
wire _517_;
wire _518_;
wire _519_;
wire _520_;
wire _521_;
wire _522_;
wire _523_;
wire _524_;
wire _525_;
wire _526_;
wire _527_;
wire _528_;
wire _529_;
wire _530_;
wire _531_;
wire _532_;
wire _533_;
wire _534_;
wire _535_;
wire _536_;
wire _537_;
wire _538_;
wire _539_;
wire _540_;
wire _541_;
wire _542_;
wire _543_;
wire _544_;
wire _545_;
wire _546_;
wire _547_;
wire _548_;
wire _549_;
wire _550_;
wire _551_;
wire _552_;
wire _553_;
wire _554_;
wire _555_;
wire _556_;
wire _557_;
wire _558_;
wire _559_;
wire _560_;
wire _561_;
wire _562_;
wire _563_;
wire _564_;
wire _565_;
wire _566_;
wire _567_;
wire _568_;
wire _569_;
wire _570_;
wire _571_;
wire _572_;
wire _573_;
wire _574_;
wire _575_;
wire _576_;
wire _577_;
wire _578_;
wire _579_;
wire _580_;
wire _581_;
wire _582_;
wire _583_;
wire _584_;
wire _585_;
wire _586_;
wire _587_;
wire _588_;
wire _589_;
wire _590_;
wire _591_;
wire _592_;
wire _593_;
wire _594_;
wire _595_;
wire _596_;
wire _597_;
wire _598_;
wire _599_;
wire _600_;
wire _601_;
wire _602_;
wire _603_;
wire _604_;
wire _605_;
wire _606_;
wire _607_;
wire _608_;
wire _609_;
wire _610_;
wire _611_;
wire _612_;
wire _613_;
wire _614_;
wire _615_;
wire _616_;
wire _617_;
wire _618_;
wire _619_;
wire _620_;
wire _621_;
wire _622_;
wire _623_;
wire _624_;
wire _625_;
wire _626_;
wire _627_;
wire _628_;
wire _629_;
wire _630_;
wire _631_;
wire _632_;
wire _633_;
wire _634_;
wire _635_;
wire _636_;
wire _637_;
wire _638_;
wire _639_;
wire _640_;
wire _641_;
wire _642_;
wire _643_;
wire _644_;
wire _645_;
wire _646_;
wire _647_;
wire _648_;
wire _649_;
wire _650_;
wire _651_;
wire _652_;
wire _653_;
wire _654_;
wire _655_;
wire _656_;
wire _657_;
wire _658_;
wire _659_;
wire _660_;
wire _661_;
wire _662_;
wire _663_;
wire _664_;
wire _665_;
wire _666_;
wire _667_;
wire _668_;
wire _669_;
wire _670_;
wire _671_;
wire _672_;
wire _673_;
wire _674_;
wire _675_;
wire _676_;
wire _677_;
wire _678_;
wire _679_;
wire _680_;
wire _681_;
wire _682_;
wire _683_;
wire _684_;
wire _685_;
wire _686_;
wire _687_;
wire _688_;
wire _689_;
wire _690_;
wire _691_;
wire _692_;
wire _693_;
wire _694_;
wire _695_;
wire _696_;
wire _697_;
wire _698_;
wire _699_;
wire _700_;
wire _701_;
wire _702_;
wire _703_;
wire _704_;
wire _705_;
wire _706_;
wire _707_;
wire _708_;
wire _709_;
wire _710_;
wire _711_;
wire _712_;
wire _713_;
wire _714_;
wire _715_;
wire _716_;
wire _717_;
wire _718_;
wire _719_;
wire _720_;
wire _721_;
wire _722_;
wire _723_;
wire _724_;
wire _725_;
wire _726_;
wire _727_;
wire _728_;
wire _729_;
wire _730_;
wire _731_;
wire _732_;
wire _733_;
wire _734_;
wire _735_;
wire _736_;
wire _737_;
wire _738_;
wire _739_;
wire _740_;
wire _741_;
wire _742_;
wire _743_;
wire _744_;
wire _745_;
wire _746_;
wire _747_;
wire _748_;
wire _749_;
wire _750_;
wire _751_;
wire _752_;
wire _753_;
wire _754_;
wire _755_;
wire _756_;
wire _757_;
wire _758_;
wire _759_;
wire _760_;
wire _761_;
wire _762_;
wire _763_;
wire _764_;
wire _765_;
wire _766_;
wire _767_;
wire _768_;
wire _769_;
wire _770_;
wire _771_;
wire _772_;
wire _773_;
wire _774_;
wire _775_;
wire _776_;
wire _777_;
wire _778_;
wire _779_;
wire _780_;
wire _781_;
wire _782_;
wire _783_;
wire _784_;
wire _785_;
wire _786_;
wire _787_;
wire _788_;
wire _789_;
wire _790_;
wire _791_;
wire _792_;
wire _793_;
wire _794_;
wire _795_;
wire _796_;
wire _797_;
wire _798_;
wire _799_;
wire _800_;
wire _801_;
wire _802_;
wire _803_;
wire _804_;
wire _805_;
wire _806_;
wire _807_;
wire _808_;
wire _809_;
wire _810_;
wire _811_;
wire _812_;
wire _813_;
wire _814_;
wire _815_;
wire _816_;
wire _817_;
wire _818_;
wire _819_;
wire _820_;
wire _821_;
wire _822_;
wire _823_;
wire _824_;
wire _825_;
wire _826_;
wire _827_;
wire _828_;
wire _829_;
wire _830_;
wire _831_;
wire _832_;
wire _833_;
wire _834_;
wire _835_;
wire _836_;
wire _837_;
wire _838_;
wire _839_;
wire _840_;
wire _841_;
wire _842_;
wire _843_;
wire _844_;
wire _845_;
wire _846_;
wire _847_;
wire _848_;
wire _849_;
wire _850_;
wire _851_;
wire _852_;
wire _853_;
wire _854_;
wire _855_;
wire _856_;
wire _857_;
wire _858_;
wire _859_;
wire _860_;
wire _861_;
wire _862_;
wire _863_;
wire _864_;
wire _865_;
wire _866_;
wire _867_;
wire _868_;
wire _869_;
wire _870_;
wire _871_;
wire _872_;
wire _873_;
wire _874_;
wire _875_;
wire _876_;
wire _877_;
wire _878_;
wire _879_;
wire _880_;
wire _881_;
wire _882_;
wire _883_;
wire _884_;
wire _885_;
wire _886_;
wire _887_;
wire _888_;
wire _889_;
wire _890_;
wire _891_;
wire _892_;
wire _893_;
wire _894_;
wire _895_;
wire _896_;
wire _897_;
wire _898_;
wire _899_;
wire _900_;
wire _901_;
wire _902_;
wire _903_;
wire _904_;
wire _905_;
wire _906_;
wire _907_;
wire _908_;
wire _909_;
wire _910_;
wire _911_;
wire _912_;
wire _913_;
wire _914_;
wire _915_;
wire _916_;
wire _917_;
wire _918_;
wire _919_;
wire _920_;
wire _921_;
wire _922_;
wire _923_;
wire _924_;
wire _925_;
wire _926_;
wire _927_;
wire _928_;
wire _929_;
wire _930_;
wire _931_;
wire _932_;
wire _933_;
wire _934_;
wire _935_;
wire _936_;
wire _937_;
wire _938_;
wire _939_;
wire _940_;
wire _941_;
wire _942_;
wire _943_;
wire _944_;
wire _945_;
wire _946_;
wire _947_;
wire _948_;
wire _949_;
wire _950_;
wire _951_;
wire _952_;
wire _953_;
wire _954_;
wire _955_;
wire _956_;
wire _957_;
wire _958_;
wire _959_;
wire _960_;
wire _961_;
wire _962_;
wire _963_;
wire _964_;
wire _965_;
wire _966_;
wire _967_;
wire _968_;
wire _969_;
wire _970_;
wire _971_;
wire _972_;
wire _973_;
wire _974_;
wire _975_;
wire _976_;
wire _977_;
wire _978_;
wire _979_;
wire _980_;
wire _981_;
wire _982_;
wire _983_;
wire _984_;
wire _985_;
wire _986_;
wire _987_;
wire _988_;
wire _989_;
wire _990_;
wire _991_;
wire _992_;
wire _993_;
wire _994_;
wire _995_;
wire _996_;
wire _997_;
wire _998_;
wire _999_;
wire _1000_;
wire _1001_;
wire _1002_;
wire _1003_;
wire _1004_;
wire _1005_;
wire _1006_;
wire _1007_;
wire _1008_;
wire _1009_;
wire _1010_;
wire _1011_;
wire _1012_;
wire _1013_;
wire _1014_;
wire _1015_;
wire _1016_;
wire _1017_;
wire _1018_;
wire _1019_;
wire _1020_;
wire _1021_;
wire _1022_;
wire _1023_;
wire _1024_;
wire _1025_;
wire _1026_;
wire _1027_;
wire _1028_;
wire _1029_;
wire _1030_;
wire _1031_;
wire _1032_;
wire _1033_;
wire _1034_;
wire _1035_;
wire _1036_;
wire _1037_;
wire _1038_;
wire _1039_;
wire _1040_;
wire _1041_;
wire _1042_;
wire _1043_;
wire _1044_;
wire _1045_;
wire _1046_;
wire _1047_;
wire _1048_;
wire _1049_;
wire _1050_;
wire _1051_;
wire _1052_;
wire _1053_;
wire _1054_;
wire _1055_;
wire _1056_;
wire _1057_;
wire _1058_;
wire _1059_;
wire _1060_;
wire _1061_;
wire _1062_;
wire _1063_;
wire _1064_;
wire _1065_;
wire _1066_;
wire _1067_;
wire _1068_;
wire _1069_;
wire _1070_;
wire _1071_;
wire _1072_;
wire _1073_;
wire _1074_;
wire _1075_;
wire _1076_;
wire _1077_;
wire _1078_;
wire _1079_;
wire _1080_;
wire _1081_;
wire _1082_;
wire _1083_;
wire _1084_;
wire _1085_;
wire _1086_;
wire _1087_;
wire _1088_;
wire _1089_;
wire _1090_;
wire _1091_;
wire _1092_;
wire _1093_;
wire _1094_;
wire _1095_;
wire _1096_;
wire _1097_;
wire _1098_;
wire _1099_;
wire _1100_;
wire _1101_;
wire _1102_;
wire _1103_;
wire _1104_;
wire _1105_;
wire _1106_;
wire _1107_;
wire _1108_;
wire _1109_;
wire _1110_;
wire _1111_;
wire _1112_;
wire _1113_;
wire _1114_;
wire _1115_;
wire _1116_;
wire _1117_;
wire _1118_;
wire _1119_;
wire _1120_;
wire _1121_;
wire _1122_;
wire _1123_;
wire _1124_;
wire _1125_;
wire _1126_;
wire _1127_;
wire _1128_;
wire _1129_;
wire _1130_;
wire _1131_;
wire _1132_;
wire _1133_;
wire _1134_;
wire _1135_;
wire _1136_;
wire _1137_;
wire _1138_;
wire _1139_;
wire _1140_;
wire _1141_;
wire _1142_;
wire _1143_;
wire _1144_;
wire _1145_;
wire _1146_;
wire _1147_;
wire _1148_;
wire _1149_;
wire _1150_;
wire _1151_;
wire _1152_;
wire _1153_;
wire _1154_;
wire _1155_;
wire _1156_;
wire _1157_;
wire _1158_;
wire _1159_;
wire _1160_;
wire _1161_;
wire _1162_;
wire _1163_;
wire _1164_;
wire _1165_;
wire _1166_;
wire _1167_;
wire _1168_;
wire _1169_;
wire _1170_;
wire _1171_;
wire _1172_;
wire _1173_;
wire _1174_;
wire _1175_;
wire _1176_;
wire _1177_;
wire _1178_;
wire _1179_;
wire _1180_;
wire _1181_;
wire _1182_;
wire _1183_;
wire _1184_;
wire _1185_;
wire _1186_;
wire _1187_;
wire _1188_;
wire _1189_;
wire _1190_;
wire _1191_;
wire _1192_;
wire _1193_;
wire _1194_;
wire _1195_;
wire _1196_;
wire _1197_;
wire _1198_;
wire _1199_;
wire _1200_;
wire _1201_;
wire _1202_;
wire _1203_;
wire _1204_;
wire _1205_;
wire _1206_;
wire _1207_;
wire _1208_;
wire _1209_;
wire _1210_;
wire _1211_;
wire _1212_;
wire _1213_;
wire _1214_;
wire _1215_;
wire _1216_;
wire _1217_;
wire _1218_;
wire _1219_;
wire _1220_;
wire _1221_;
wire _1222_;
wire _1223_;
wire _1224_;
wire _1225_;
wire _1226_;
wire _1227_;
wire _1228_;
wire _1229_;
wire _1230_;
wire _1231_;
wire _1232_;
wire _1233_;
wire _1234_;
wire _1235_;
wire _1236_;
wire _1237_;
wire _1238_;
wire _1239_;
wire _1240_;
wire _1241_;
wire _1242_;
wire _1243_;
wire _1244_;
wire _1245_;
wire _1246_;
wire _1247_;
wire _1248_;
wire _1249_;
wire _1250_;
wire _1251_;
wire _1252_;
wire _1253_;
wire _1254_;
wire _1255_;
wire _1256_;
wire _1257_;
wire _1258_;
wire _1259_;
wire _1260_;
wire _1261_;
wire _1262_;
wire _1263_;
wire _1264_;
wire _1265_;
wire _1266_;
wire _1267_;
wire _1268_;
wire _1269_;
wire _1270_;
wire _1271_;
wire _1272_;
wire _1273_;
wire _1274_;
wire _1275_;
wire _1276_;
wire _1277_;
wire _1278_;
wire _1279_;
wire _1280_;
wire _1281_;
wire _1282_;
wire _1283_;
wire _1284_;
wire _1285_;
wire _1286_;
wire _1287_;
wire _1288_;
wire _1289_;
wire _1290_;
wire _1291_;
wire _1292_;
wire _1293_;
wire _1294_;
wire _1295_;
wire _1296_;
wire _1297_;
wire _1298_;
wire _1299_;
wire _1300_;
wire _1301_;
wire _1302_;
wire _1303_;
wire _1304_;
wire _1305_;
wire _1306_;
wire _1307_;
wire _1308_;
wire _1309_;
wire _1310_;
wire _1311_;
wire _1312_;
wire _1313_;
wire _1314_;
wire _1315_;
wire _1316_;
wire _1317_;
wire _1318_;
wire _1319_;
wire _1320_;
wire _1321_;
wire _1322_;
wire _1323_;
wire _1324_;
wire _1325_;
wire _1326_;
wire _1327_;
wire _1328_;
wire _1329_;
wire _1330_;
wire _1331_;
wire _1332_;
wire _1333_;
wire _1334_;
wire _1335_;
wire _1336_;
wire _1337_;
wire _1338_;
wire _1339_;
wire _1340_;
wire _1341_;
wire _1342_;
wire _1343_;
wire _1344_;
wire _1345_;
wire _1346_;
wire _1347_;
wire _1348_;
wire _1349_;
wire _1350_;
wire _1351_;
wire _1352_;
wire _1353_;
wire _1354_;
wire _1355_;
wire _1356_;
wire _1357_;
wire _1358_;
wire _1359_;
wire _1360_;
wire _1361_;
wire _1362_;
wire _1363_;
wire _1364_;
wire _1365_;
wire _1366_;
wire _1367_;
wire _1368_;
wire _1369_;
wire _1370_;
wire _1371_;
wire _1372_;
wire _1373_;
wire _1374_;
wire _1375_;
wire _1376_;
wire _1377_;
wire _1378_;
wire _1379_;
wire _1380_;
wire _1381_;
wire _1382_;
wire _1383_;
wire _1384_;
wire _1385_;
wire _1386_;
wire _1387_;
wire _1388_;
wire _1389_;
wire _1390_;
wire _1391_;
wire _1392_;
wire _1393_;
wire _1394_;
wire _1395_;
wire _1396_;
wire _1397_;
wire _1398_;
wire _1399_;
wire _1400_;
wire _1401_;
wire _1402_;
wire _1403_;
wire _1404_;
wire _1405_;
wire _1406_;
wire _1407_;
wire _1408_;
wire _1409_;
wire _1410_;
wire _1411_;
wire _1412_;
wire _1413_;
wire _1414_;
wire _1415_;
wire _1416_;
wire _1417_;
wire _1418_;
wire _1419_;
wire _1420_;
wire _1421_;
wire _1422_;
wire _1423_;
wire _1424_;
wire _1425_;
wire _1426_;
wire _1427_;
wire _1428_;
wire _1429_;
wire _1430_;
wire _1431_;
wire _1432_;
wire _1433_;
wire _1434_;
wire _1435_;
wire _1436_;
wire _1437_;
wire _1438_;
wire _1439_;
wire _1440_;
wire _1441_;
wire _1442_;
wire _1443_;
wire _1444_;
wire _1445_;
wire _1446_;
wire _1447_;
wire _1448_;
wire _1449_;
wire _1450_;
wire _1451_;
wire _1452_;
wire _1453_;
wire _1454_;
wire _1455_;
wire _1456_;
wire _1457_;
wire _1458_;
wire _1459_;
wire _1460_;
wire _1461_;
wire _1462_;
wire _1463_;
wire _1464_;
wire _1465_;
wire _1466_;
wire _1467_;
wire _1468_;
wire _1469_;
wire _1470_;
wire _1471_;
wire _1472_;
wire _1473_;
wire _1474_;
wire _1475_;
wire _1476_;
wire _1477_;
wire _1478_;
wire _1479_;
wire _1480_;
wire _1481_;
wire _1482_;
wire _1483_;
wire _1484_;
wire _1485_;
wire _1486_;
wire _1487_;
wire _1488_;
wire _1489_;
wire _1490_;
wire _1491_;
wire _1492_;
wire _1493_;
wire _1494_;
wire _1495_;
wire _1496_;
wire _1497_;
wire _1498_;
wire _1499_;
wire _1500_;
wire _1501_;
wire _1502_;
wire _1503_;
wire _1504_;
wire _1505_;
wire _1506_;
wire _1507_;
wire _1508_;
wire _1509_;
wire _1510_;
wire _1511_;
wire _1512_;
wire _1513_;
wire _1514_;
wire _1515_;
wire _1516_;
wire _1517_;
wire _1518_;
wire _1519_;
wire _1520_;
wire _1521_;
wire _1522_;
wire _1523_;
wire _1524_;
wire _1525_;
wire _1526_;
wire _1527_;
wire _1528_;
wire _1529_;
wire _1530_;
wire _1531_;
wire _1532_;
wire _1533_;
wire _1534_;
wire _1535_;
wire _1536_;
wire _1537_;
wire _1538_;
wire _1539_;
wire _1540_;
wire _1541_;
wire _1542_;
wire _1543_;
wire _1544_;
wire _1545_;
wire _1546_;
wire _1547_;
wire _1548_;
wire _1549_;
wire _1550_;
wire _1551_;
wire _1552_;
wire _1553_;
wire _1554_;
wire _1555_;
wire _1556_;
wire _1557_;
wire _1558_;
wire _1559_;
wire _1560_;
wire _1561_;
wire _1562_;
wire _1563_;
wire _1564_;
wire _1565_;
wire _1566_;
wire _1567_;
wire _1568_;
wire _1569_;
wire _1570_;
wire _1571_;
wire _1572_;
wire _1573_;
wire _1574_;
wire _1575_;
wire _1576_;
wire _1577_;
wire _1578_;
wire _1579_;
wire _1580_;
wire _1581_;
wire _1582_;
wire _1583_;
wire _1584_;
wire _1585_;
wire _1586_;
wire _1587_;
wire _1588_;
wire _1589_;
wire _1590_;
wire _1591_;
wire _1592_;
wire _1593_;
wire _1594_;
wire _1595_;
wire _1596_;
wire _1597_;
wire _1598_;
wire _1599_;
wire _1600_;
wire _1601_;
wire _1602_;
wire _1603_;
wire _1604_;
wire _1605_;
wire _1606_;
wire _1607_;
wire _1608_;
wire _1609_;
wire _1610_;
wire _1611_;
wire _1612_;
wire _1613_;
wire _1614_;
wire _1615_;
wire _1616_;
wire _1617_;
wire _1618_;
wire _1619_;
wire _1620_;
wire _1621_;
wire _1622_;
wire _1623_;
wire _1624_;
wire _1625_;
wire _1626_;
wire _1627_;
wire _1628_;
wire _1629_;
wire _1630_;
wire _1631_;
wire _1632_;
wire _1633_;
wire _1634_;
wire _1635_;
wire _1636_;
wire _1637_;
wire _1638_;
wire _1639_;
wire _1640_;
wire _1641_;
wire _1642_;
wire _1643_;
wire _1644_;
wire _1645_;
wire _1646_;
wire _1647_;
wire _1648_;
wire _1649_;
wire _1650_;
wire _1651_;
wire _1652_;
wire _1653_;
wire _1654_;
wire _1655_;
wire _1656_;
wire _1657_;
wire _1658_;
wire _1659_;
wire _1660_;
wire _1661_;
wire _1662_;
wire _1663_;
wire _1664_;
wire _1665_;
wire _1666_;
wire _1667_;
wire _1668_;
wire _1669_;
wire _1670_;
wire _1671_;
wire _1672_;
wire _1673_;
wire _1674_;
wire _1675_;
wire _1676_;
wire _1677_;
wire _1678_;
wire _1679_;
wire _1680_;
wire _1681_;
wire _1682_;
wire _1683_;
wire _1684_;
wire _1685_;
wire _1686_;
wire _1687_;
wire _1688_;
wire _1689_;
wire _1690_;
wire _1691_;
wire _1692_;
wire _1693_;
wire _1694_;
wire _1695_;
wire _1696_;
wire _1697_;
wire _1698_;
wire _1699_;
wire _1700_;
wire _1701_;
wire _1702_;
wire _1703_;
wire _1704_;
wire _1705_;
wire _1706_;
wire _1707_;
wire _1708_;
wire _1709_;
wire _1710_;
wire _1711_;
wire _1712_;
wire _1713_;
wire _1714_;
wire _1715_;
wire _1716_;
wire _1717_;
wire _1718_;
wire _1719_;
wire _1720_;
wire _1721_;
wire _1722_;
wire _1723_;
wire _1724_;
wire _1725_;
wire _1726_;
wire _1727_;
wire _1728_;
wire _1729_;
wire _1730_;
wire _1731_;
wire _1732_;
wire _1733_;
wire _1734_;
wire _1735_;
wire _1736_;
wire _1737_;
wire _1738_;
wire _1739_;
wire _1740_;
wire _1741_;
wire _1742_;
wire _1743_;
wire _1744_;
wire _1745_;
wire _1746_;
wire _1747_;
wire _1748_;
wire _1749_;
wire _1750_;
wire _1751_;
wire _1752_;
wire _1753_;
wire _1754_;
wire _1755_;
wire _1756_;
wire _1757_;
wire _1758_;
wire _1759_;
wire _1760_;
wire _1761_;
wire _1762_;
wire _1763_;
wire _1764_;
wire _1765_;
wire _1766_;
wire _1767_;
wire _1768_;
wire _1769_;
wire _1770_;
wire _1771_;
wire _1772_;
wire _1773_;
wire _1774_;
wire _1775_;
wire _1776_;
wire _1777_;
wire _1778_;
wire _1779_;
wire _1780_;
wire _1781_;
wire _1782_;
wire _1783_;
wire _1784_;
wire _1785_;
wire _1786_;
wire _1787_;
wire _1788_;
wire _1789_;
wire _1790_;
wire _1791_;
wire _1792_;
wire _1793_;
wire _1794_;
wire _1795_;
wire _1796_;
wire _1797_;
wire _1798_;
wire _1799_;
wire _1800_;
wire _1801_;
wire _1802_;
wire _1803_;
wire _1804_;
wire _1805_;
wire _1806_;
wire _1807_;
wire _1808_;
wire _1809_;
wire _1810_;
wire _1811_;
wire _1812_;
wire _1813_;
wire _1814_;
wire _1815_;
wire _1816_;
wire _1817_;
wire _1818_;
wire _1819_;
wire _1820_;
wire _1821_;
wire _1822_;
wire _1823_;
wire _1824_;
wire _1825_;
wire _1826_;
wire _1827_;
wire _1828_;
wire _1829_;
wire _1830_;
wire _1831_;
wire _1832_;
wire _1833_;
wire _1834_;
wire _1835_;
wire _1836_;
wire _1837_;
wire _1838_;
wire _1839_;
wire _1840_;
wire _1841_;
wire _1842_;
wire _1843_;
wire _1844_;
wire _1845_;
wire _1846_;
wire _1847_;
wire _1848_;
wire _1849_;
wire _1850_;
wire _1851_;
wire _1852_;
wire _1853_;
wire _1854_;
wire _1855_;
wire _1856_;
wire _1857_;
wire _1858_;
wire _1859_;
wire _1860_;
wire _1861_;
wire _1862_;
wire _1863_;
wire _1864_;
wire _1865_;
wire _1866_;
wire _1867_;
wire _1868_;
wire _1869_;
wire _1870_;
wire _1871_;
wire _1872_;
wire _1873_;
wire _1874_;
wire _1875_;
wire _1876_;
wire _1877_;
wire _1878_;
wire _1879_;
wire _1880_;
wire _1881_;
wire _1882_;
wire _1883_;
wire _1884_;
wire _1885_;
wire _1886_;
wire _1887_;
wire _1888_;
wire _1889_;
wire _1890_;
wire _1891_;
wire _1892_;
wire _1893_;
wire _1894_;
wire _1895_;
wire _1896_;
wire _1897_;
wire _1898_;
wire _1899_;
wire _1900_;
wire _1901_;
wire _1902_;
wire _1903_;
wire _1904_;
wire _1905_;
wire _1906_;
wire _1907_;
wire _1908_;
wire _1909_;
wire _1910_;
wire _1911_;
wire _1912_;
wire _1913_;
wire _1914_;
wire _1915_;
wire _1916_;
wire _1917_;
wire _1918_;
wire _1919_;
wire _1920_;
wire _1921_;
wire _1922_;
wire _1923_;
wire _1924_;
wire _1925_;
wire _1926_;
wire _1927_;
wire _1928_;
wire _1929_;
wire _1930_;
wire _1931_;
wire _1932_;
wire _1933_;
wire _1934_;
wire _1935_;
wire _1936_;
wire _1937_;
wire _1938_;
wire _1939_;
wire _1940_;
wire _1941_;
wire _1942_;
wire _1943_;
wire _1944_;
wire _1945_;
wire _1946_;
wire _1947_;
wire _1948_;
wire _1949_;
wire _1950_;
wire _1951_;
wire _1952_;
wire _1953_;
wire _1954_;
wire _1955_;
wire _1956_;
wire _1957_;
wire _1958_;
wire _1959_;
wire _1960_;
wire _1961_;
wire _1962_;
wire _1963_;
wire _1964_;
wire _1965_;
wire _1966_;
wire _1967_;
wire _1968_;
wire _1969_;
wire _1970_;
wire _1971_;
wire _1972_;
wire _1973_;
wire _1974_;
wire _1975_;
wire _1976_;
wire _1977_;
wire _1978_;
wire _1979_;
wire _1980_;
wire _1981_;
wire _1982_;
wire _1983_;
wire _1984_;
wire _1985_;
wire _1986_;
wire _1987_;
wire _1988_;
wire _1989_;
wire _1990_;
wire _1991_;
wire _1992_;
wire _1993_;
wire _1994_;
wire _1995_;
wire _1996_;
wire _1997_;
wire _1998_;
wire _1999_;
wire _2000_;
wire _2001_;
wire _2002_;
wire _2003_;
wire _2004_;
wire _2005_;
wire _2006_;
wire _2007_;
wire _2008_;
wire _2009_;
wire _2010_;
wire _2011_;
wire _2012_;
wire _2013_;
wire _2014_;
wire _2015_;
wire _2016_;
wire _2017_;
wire _2018_;
wire _2019_;
wire _2020_;
wire _2021_;
wire _2022_;
wire _2023_;
wire _2024_;
wire _2025_;
wire _2026_;
wire _2027_;
wire _2028_;
wire _2029_;
wire _2030_;
wire _2031_;
wire _2032_;
wire _2033_;
wire _2034_;
wire _2035_;
wire _2036_;
wire _2037_;
wire _2038_;
wire _2039_;
wire _2040_;
wire _2041_;
wire _2042_;
wire _2043_;
wire _2044_;
wire _2045_;
wire _2046_;
wire _2047_;
wire _2048_;
wire _2049_;
wire _2050_;
wire _2051_;
wire _2052_;
wire _2053_;
wire _2054_;
wire _2055_;
wire _2056_;
wire _2057_;
wire _2058_;
wire _2059_;
wire _2060_;
wire _2061_;
wire _2062_;
wire _2063_;
wire _2064_;
wire _2065_;
wire _2066_;
wire _2067_;
wire _2068_;
wire _2069_;
wire _2070_;
wire _2071_;
wire _2072_;
wire _2073_;
wire _2074_;
wire _2075_;
wire _2076_;
wire _2077_;
wire _2078_;
wire _2079_;
wire _2080_;
wire _2081_;
wire _2082_;
wire _2083_;
wire _2084_;
wire _2085_;
wire _2086_;
wire _2087_;
wire _2088_;
wire _2089_;
wire _2090_;
wire _2091_;
wire _2092_;
wire _2093_;
wire _2094_;
wire _2095_;
wire _2096_;
wire _2097_;
wire _2098_;
wire _2099_;
wire _2100_;
wire _2101_;
wire _2102_;
wire _2103_;
wire _2104_;
wire _2105_;
wire _2106_;
wire _2107_;
wire _2108_;
wire _2109_;
wire _2110_;
wire _2111_;
wire _2112_;
wire _2113_;
wire _2114_;
wire _2115_;
wire _2116_;
wire _2117_;
wire _2118_;
wire _2119_;
wire _2120_;
wire _2121_;
wire _2122_;
wire _2123_;
wire _2124_;
wire _2125_;
wire _2126_;
wire _2127_;
wire _2128_;
wire _2129_;
wire _2130_;
wire _2131_;
wire _2132_;
wire _2133_;
wire _2134_;
wire _2135_;
wire _2136_;
wire _2137_;
wire _2138_;
wire _2139_;
wire _2140_;
wire _2141_;
wire _2142_;
wire _2143_;
wire _2144_;
wire _2145_;
wire _2146_;
wire _2147_;
wire _2148_;
wire _2149_;
wire _2150_;
wire _2151_;
wire _2152_;
wire _2153_;
wire _2154_;
wire _2155_;
wire _2156_;
wire _2157_;
wire _2158_;
wire _2159_;
wire _2160_;
wire _2161_;
wire _2162_;
wire _2163_;
wire _2164_;
wire _2165_;
wire _2166_;
wire _2167_;
wire _2168_;
wire _2169_;
wire _2170_;
wire _2171_;
wire _2172_;
wire _2173_;
wire _2174_;
wire _2175_;
wire _2176_;
wire _2177_;
wire _2178_;
wire _2179_;
wire _2180_;
wire _2181_;
wire _2182_;
wire _2183_;
wire _2184_;
wire _2185_;
wire _2186_;
wire _2187_;
wire _2188_;
wire _2189_;
wire _2190_;
wire _2191_;
wire _2192_;
wire _2193_;
wire _2194_;
wire _2195_;
wire _2196_;
wire _2197_;
wire _2198_;
wire _2199_;
wire _2200_;
wire _2201_;
wire _2202_;
wire _2203_;
wire _2204_;
wire _2205_;
wire _2206_;
wire _2207_;
wire _2208_;
wire _2209_;
wire _2210_;
wire _2211_;
wire _2212_;
wire _2213_;
wire _2214_;
wire _2215_;
wire _2216_;
wire _2217_;
wire _2218_;
wire _2219_;
wire _2220_;
wire _2221_;
wire _2222_;
wire _2223_;
wire _2224_;
wire _2225_;
wire _2226_;
wire _2227_;
wire _2228_;
wire _2229_;
wire _2230_;
wire _2231_;
wire _2232_;
wire _2233_;
wire _2234_;
wire _2235_;
wire _2236_;
wire _2237_;
wire _2238_;
wire _2239_;
wire _2240_;
wire _2241_;
wire _2242_;
wire _2243_;
wire _2244_;
wire _2245_;
wire _2246_;
wire _2247_;
wire _2248_;
wire _2249_;
wire _2250_;
wire _2251_;
wire _2252_;
wire _2253_;
wire _2254_;
wire _2255_;
wire _2256_;
wire _2257_;
wire _2258_;
wire _2259_;
wire _2260_;
wire _2261_;
wire _2262_;
wire _2263_;
wire _2264_;
wire _2265_;
wire _2266_;
wire _2267_;
wire _2268_;
wire _2269_;
wire _2270_;
wire _2271_;
wire _2272_;
wire _2273_;
wire _2274_;
wire _2275_;
wire _2276_;
wire _2277_;
wire _2278_;
wire _2279_;
wire _2280_;
wire _2281_;
wire _2282_;
wire _2283_;
wire _2284_;
wire _2285_;
wire _2286_;
wire _2287_;
wire _2288_;
wire _2289_;
wire _2290_;
wire _2291_;
wire _2292_;
wire _2293_;
wire _2294_;
wire _2295_;
wire _2296_;
wire _2297_;
wire _2298_;
wire _2299_;
wire _2300_;
wire _2301_;
wire _2302_;
wire _2303_;
wire _2304_;
wire _2305_;
wire _2306_;
wire _2307_;
wire _2308_;
wire _2309_;
wire _2310_;
wire _2311_;
wire _2312_;
wire _2313_;
wire _2314_;
wire _2315_;
wire _2316_;
wire _2317_;
wire _2318_;
wire _2319_;
wire _2320_;
wire _2321_;
wire _2322_;
wire _2323_;
wire _2324_;
wire _2325_;
wire _2326_;
wire _2327_;
wire _2328_;
wire _2329_;
wire _2330_;
wire _2331_;
wire _2332_;
wire _2333_;
wire _2334_;
wire _2335_;
wire _2336_;
wire _2337_;
wire _2338_;
wire _2339_;
wire _2340_;
wire _2341_;
wire _2342_;
wire _2343_;
wire _2344_;
wire _2345_;
wire _2346_;
wire _2347_;
wire _2348_;
wire _2349_;
wire _2350_;
wire _2351_;
wire _2352_;
wire _2353_;
wire _2354_;
wire _2355_;
wire _2356_;
wire _2357_;
wire _2358_;
wire _2359_;
wire _2360_;
wire _2361_;
wire _2362_;
wire _2363_;
wire _2364_;
wire _2365_;
wire _2366_;
wire _2367_;
wire _2368_;
wire _2369_;
wire _2370_;
wire _2371_;
wire _2372_;
wire _2373_;
wire _2374_;
wire _2375_;
wire _2376_;
wire _2377_;
wire _2378_;
wire _2379_;
wire _2380_;
wire _2381_;
wire _2382_;
wire _2383_;
wire _2384_;
wire _2385_;
wire _2386_;
wire _2387_;
wire _2388_;
wire _2389_;
wire _2390_;
wire _2391_;
wire _2392_;
wire _2393_;
wire _2394_;
wire _2395_;
wire _2396_;
wire _2397_;
wire _2398_;
wire _2399_;
wire _2400_;
wire _2401_;
wire _2402_;
wire _2403_;
wire _2404_;
wire _2405_;
wire _2406_;
wire _2407_;
wire _2408_;
wire _2409_;
wire _2410_;
wire _2411_;
wire _2412_;
wire _2413_;
wire _2414_;
wire _2415_;
wire _2416_;
wire _2417_;
wire _2418_;
wire _2419_;
wire _2420_;
wire _2421_;
wire _2422_;
wire _2423_;
wire _2424_;
wire _2425_;
wire _2426_;
wire _2427_;
wire _2428_;
wire _2429_;
wire _2430_;
wire _2431_;
wire _2432_;
wire _2433_;
wire _2434_;
wire _2435_;
wire _2436_;
wire _2437_;
wire _2438_;
wire _2439_;
wire _2440_;
wire _2441_;
wire _2442_;
wire _2443_;
wire _2444_;
wire _2445_;
wire _2446_;
wire _2447_;
wire _2448_;
wire _2449_;
wire _2450_;
wire _2451_;
wire _2452_;
wire _2453_;
wire _2454_;
wire _2455_;
wire _2456_;
wire _2457_;
wire _2458_;
wire _2459_;
wire _2460_;
wire _2461_;
wire _2462_;
wire _2463_;
wire _2464_;
wire _2465_;
wire _2466_;
wire _2467_;
wire _2468_;
wire _2469_;
wire _2470_;
wire _2471_;
wire _2472_;
wire _2473_;
wire _2474_;
wire _2475_;
wire _2476_;
wire _2477_;
wire _2478_;
wire _2479_;
wire _2480_;
wire _2481_;
wire _2482_;
wire _2483_;
wire _2484_;
wire _2485_;
wire _2486_;
wire _2487_;
wire _2488_;
wire _2489_;
wire _2490_;
wire _2491_;
wire _2492_;
wire _2493_;
wire _2494_;
wire _2495_;
wire _2496_;
wire _2497_;
wire _2498_;
wire _2499_;
wire _2500_;
wire _2501_;
wire _2502_;
wire _2503_;
wire _2504_;
wire _2505_;
wire _2506_;
wire _2507_;
wire _2508_;
wire _2509_;
wire _2510_;
wire _2511_;
wire _2512_;
wire _2513_;
wire _2514_;
wire _2515_;
wire _2516_;
wire _2517_;
wire _2518_;
wire _2519_;
wire _2520_;
wire _2521_;
wire _2522_;
wire _2523_;
wire _2524_;
wire _2525_;
wire _2526_;
wire _2527_;
wire _2528_;
wire _2529_;
wire _2530_;
wire _2531_;
wire _2532_;
wire _2533_;
wire _2534_;
wire _2535_;
wire _2536_;
wire _2537_;
wire _2538_;
wire _2539_;
wire _2540_;
wire _2541_;
wire _2542_;
wire _2543_;
wire _2544_;
wire _2545_;
wire _2546_;
wire _2547_;
wire _2548_;
wire _2549_;
wire _2550_;
wire _2551_;
wire _2552_;
wire _2553_;
wire _2554_;
wire _2555_;
wire _2556_;
wire _2557_;
wire _2558_;
wire _2559_;
wire _2560_;
wire _2561_;
wire _2562_;
wire _2563_;
wire _2564_;
wire _2565_;
wire _2566_;
wire _2567_;
wire _2568_;
wire _2569_;
wire _2570_;
wire _2571_;
wire _2572_;
wire _2573_;
wire _2574_;
wire _2575_;
wire _2576_;
wire _2577_;
wire _2578_;
wire _2579_;
wire _2580_;
wire _2581_;
wire _2582_;
wire _2583_;
wire _2584_;
wire _2585_;
wire _2586_;
wire _2587_;
wire _2588_;
wire _2589_;
wire _2590_;
wire _2591_;
wire _2592_;
wire _2593_;
wire _2594_;
wire _2595_;
wire _2596_;
wire _2597_;
wire _2598_;
wire _2599_;
wire _2600_;
wire _2601_;
wire _2602_;
wire _2603_;
wire _2604_;
wire _2605_;
wire _2606_;
wire _2607_;
wire _2608_;
wire _2609_;
wire _2610_;
wire _2611_;
wire _2612_;
wire _2613_;
wire _2614_;
wire _2615_;
wire _2616_;
wire _2617_;
wire _2618_;
wire _2619_;
wire _2620_;
wire _2621_;
wire _2622_;
wire _2623_;
wire _2624_;
wire _2625_;
wire _2626_;
wire _2627_;
wire _2628_;
wire _2629_;
wire _2630_;
wire _2631_;
wire _2632_;
wire _2633_;
wire _2634_;
wire _2635_;
wire _2636_;
wire _2637_;
wire _2638_;
wire _2639_;
wire _2640_;
wire _2641_;
wire _2642_;
wire _2643_;
wire _2644_;
wire _2645_;
wire _2646_;
wire _2647_;
wire _2648_;
wire _2649_;
wire _2650_;
wire _2651_;
wire _2652_;
wire _2653_;
wire _2654_;
wire _2655_;
wire _2656_;
wire _2657_;
wire _2658_;
wire _2659_;
wire _2660_;
wire _2661_;
wire _2662_;
wire _2663_;
wire _2664_;
wire _2665_;
wire _2666_;
wire _2667_;
wire _2668_;
wire _2669_;
wire _2670_;
wire _2671_;
wire _2672_;
wire _2673_;
wire _2674_;
wire _2675_;
wire _2676_;
wire _2677_;
wire _2678_;
wire _2679_;
wire _2680_;
wire _2681_;
wire _2682_;
wire _2683_;
wire _2684_;
wire _2685_;
wire _2686_;
wire _2687_;
wire _2688_;
wire _2689_;
wire _2690_;
wire _2691_;
wire _2692_;
wire _2693_;
wire _2694_;
wire _2695_;
wire _2696_;
wire _2697_;
wire _2698_;
wire _2699_;
wire _2700_;
wire _2701_;
wire _2702_;
wire _2703_;
wire _2704_;
wire _2705_;
wire _2706_;
wire _2707_;
wire _2708_;
wire _2709_;
wire _2710_;
wire _2711_;
wire _2712_;
wire _2713_;
wire _2714_;
wire _2715_;
wire _2716_;
wire _2717_;
wire _2718_;
wire _2719_;
wire _2720_;
wire _2721_;
wire _2722_;
wire _2723_;
wire _2724_;
wire _2725_;
wire _2726_;
wire _2727_;
wire _2728_;
wire _2729_;
wire _2730_;
wire _2731_;
wire _2732_;
wire _2733_;
wire _2734_;
wire _2735_;
wire _2736_;
wire _2737_;
wire _2738_;
wire _2739_;
wire _2740_;
wire _2741_;
wire _2742_;
wire _2743_;
wire _2744_;
wire _2745_;
wire _2746_;
wire _2747_;
wire _2748_;
wire _2749_;
wire _2750_;
wire _2751_;
wire _2752_;
wire _2753_;
wire _2754_;
wire _2755_;
wire _2756_;
wire _2757_;
wire _2758_;
wire _2759_;
wire _2760_;
wire _2761_;
wire _2762_;
wire _2763_;
wire _2764_;
wire _2765_;
wire _2766_;
wire _2767_;
wire _2768_;
wire _2769_;
wire _2770_;
wire _2771_;
wire _2772_;
wire _2773_;
wire _2774_;
wire _2775_;
wire _2776_;
wire _2777_;
wire _2778_;
wire _2779_;
wire _2780_;
wire _2781_;
wire _2782_;
wire _2783_;
wire _2784_;
wire _2785_;
wire _2786_;
wire _2787_;
wire _2788_;
wire _2789_;
wire _2790_;
wire _2791_;
wire _2792_;
wire _2793_;
wire _2794_;
wire _2795_;
wire _2796_;
wire _2797_;
wire _2798_;
wire _2799_;
wire _2800_;
wire _2801_;
wire _2802_;
wire _2803_;
wire _2804_;
wire _2805_;
wire _2806_;
wire _2807_;
wire _2808_;
wire _2809_;
wire _2810_;
wire _2811_;
wire _2812_;
wire _2813_;
wire _2814_;
wire _2815_;
wire _2816_;
wire _2817_;
wire _2818_;
wire _2819_;
wire _2820_;
wire _2821_;
wire _2822_;
wire _2823_;
wire _2824_;
wire _2825_;
wire _2826_;
wire _2827_;
wire _2828_;
wire _2829_;
wire _2830_;
wire _2831_;
wire _2832_;
wire _2833_;
wire _2834_;
wire _2835_;
wire _2836_;
wire _2837_;
wire _2838_;
wire _2839_;
wire _2840_;
wire _2841_;
wire _2842_;
wire _2843_;
wire _2844_;
wire _2845_;
wire _2846_;
wire _2847_;
wire _2848_;
wire _2849_;
wire _2850_;
wire _2851_;
wire _2852_;
wire _2853_;
wire _2854_;
wire _2855_;
wire _2856_;
wire _2857_;
wire _2858_;
wire _2859_;
wire _2860_;
wire _2861_;
wire _2862_;
wire _2863_;
wire _2864_;
wire _2865_;
wire _2866_;
wire _2867_;
wire _2868_;
wire _2869_;
wire _2870_;
wire _2871_;
wire _2872_;
wire _2873_;
wire _2874_;
wire _2875_;
wire _2876_;
wire _2877_;
wire _2878_;
wire _2879_;
wire _2880_;
wire _2881_;
wire _2882_;
wire _2883_;
wire _2884_;
wire _2885_;
wire _2886_;
wire _2887_;
wire _2888_;
wire _2889_;
wire _2890_;
wire _2891_;
wire _2892_;
wire _2893_;
wire _2894_;
wire _2895_;
wire _2896_;
wire _2897_;
wire _2898_;
wire _2899_;
wire _2900_;
wire _2901_;
wire _2902_;
wire _2903_;
wire _2904_;
wire _2905_;
wire _2906_;
wire _2907_;
wire _2908_;
wire _2909_;
wire _2910_;
wire _2911_;
wire _2912_;
wire _2913_;
wire _2914_;
wire _2915_;
wire _2916_;
wire _2917_;
wire _2918_;
wire _2919_;
wire _2920_;
wire _2921_;
wire _2922_;
wire _2923_;
wire _2924_;
wire _2925_;
wire _2926_;
wire _2927_;
wire _2928_;
wire _2929_;
wire _2930_;
wire _2931_;
wire _2932_;
wire _2933_;
wire _2934_;
wire _2935_;
wire _2936_;
wire _2937_;
wire _2938_;
wire _2939_;
wire _2940_;
wire _2941_;
wire _2942_;
wire _2943_;
wire _2944_;
wire _2945_;
wire _2946_;
wire _2947_;
wire _2948_;
wire _2949_;
wire _2950_;
wire _2951_;
wire _2952_;
wire _2953_;
wire _2954_;
wire _2955_;
wire _2956_;
wire _2957_;
wire _2958_;
wire _2959_;
wire _2960_;
wire _2961_;
wire _2962_;
wire _2963_;
wire _2964_;
wire _2965_;
wire _2966_;
wire _2967_;
wire _2968_;
wire _2969_;
wire _2970_;
wire _2971_;
wire _2972_;
wire _2973_;
wire _2974_;
wire _2975_;
wire _2976_;
wire _2977_;
wire _2978_;
wire _2979_;
wire _2980_;
wire _2981_;
wire _2982_;
wire _2983_;
wire _2984_;
wire _2985_;
wire _2986_;
wire _2987_;
wire _2988_;
wire _2989_;
wire _2990_;
wire _2991_;
wire _2992_;
wire _2993_;
wire _2994_;
wire _2995_;
wire _2996_;
wire _2997_;
wire _2998_;
wire _2999_;
wire _3000_;
wire _3001_;
wire _3002_;
wire _3003_;
wire _3004_;
wire _3005_;
wire _3006_;
wire _3007_;
wire _3008_;
wire _3009_;
wire _3010_;
wire _3011_;
wire _3012_;
wire _3013_;
wire _3014_;
wire _3015_;
wire _3016_;
wire _3017_;
wire _3018_;
wire _3019_;
wire _3020_;
wire _3021_;
wire _3022_;
wire _3023_;
wire _3024_;
wire _3025_;
wire _3026_;
wire _3027_;
wire _3028_;
wire _3029_;
wire _3030_;
wire _3031_;
wire _3032_;
wire _3033_;
wire _3034_;
wire _3035_;
wire _3036_;
wire _3037_;
wire _3038_;
wire _3039_;
wire _3040_;
wire _3041_;
wire _3042_;
wire _3043_;
wire _3044_;
wire _3045_;
wire _3046_;
wire _3047_;
wire _3048_;
wire _3049_;
wire _3050_;
wire _3051_;
wire _3052_;
wire _3053_;
wire _3054_;
wire _3055_;
wire _3056_;
wire _3057_;
wire _3058_;
wire _3059_;
wire _3060_;
wire _3061_;
wire _3062_;
wire _3063_;
wire _3064_;
wire _3065_;
wire _3066_;
wire _3067_;
wire _3068_;
wire _3069_;
wire _3070_;
wire _3071_;
wire _3072_;
wire _3073_;
wire _3074_;
wire _3075_;
wire _3076_;
wire _3077_;
wire _3078_;
wire _3079_;
wire _3080_;
wire _3081_;
wire _3082_;
wire _3083_;
wire _3084_;
wire _3085_;
wire _3086_;
wire _3087_;
wire _3088_;
wire _3089_;
wire _3090_;
wire _3091_;
wire _3092_;
wire _3093_;
wire _3094_;
wire _3095_;
wire _3096_;
wire _3097_;
wire _3098_;
wire _3099_;
wire _3100_;
wire _3101_;
wire _3102_;
wire _3103_;
wire _3104_;
wire _3105_;
wire _3106_;
wire _3107_;
wire _3108_;
wire _3109_;
wire _3110_;
wire _3111_;
wire _3112_;
wire _3113_;
wire _3114_;
wire _3115_;
wire _3116_;
wire _3117_;
wire _3118_;
wire _3119_;
wire _3120_;
wire _3121_;
wire _3122_;
wire _3123_;
wire _3124_;
wire _3125_;
wire _3126_;
wire _3127_;
wire _3128_;
wire _3129_;
wire _3130_;
wire _3131_;
wire _3132_;
wire _3133_;
wire _3134_;
wire _3135_;
wire _3136_;
wire _3137_;
wire _3138_;
wire _3139_;
wire _3140_;
wire _3141_;
wire _3142_;
wire _3143_;
wire _3144_;
wire _3145_;
wire _3146_;
wire _3147_;
wire _3148_;
wire _3149_;
wire _3150_;
wire _3151_;
wire _3152_;
wire _3153_;
wire _3154_;
wire _3155_;
wire _3156_;
wire _3157_;
wire _3158_;
wire _3159_;
wire _3160_;
wire _3161_;
wire _3162_;
wire _3163_;
wire _3164_;
wire _3165_;
wire _3166_;
wire _3167_;
wire _3168_;
wire _3169_;
wire _3170_;
wire _3171_;
wire _3172_;
wire _3173_;
wire _3174_;
wire _3175_;
wire _3176_;
wire _3177_;
wire _3178_;
wire _3179_;
wire _3180_;
wire _3181_;
wire _3182_;
wire _3183_;
wire _3184_;
wire _3185_;
wire _3186_;
wire _3187_;
wire _3188_;
wire _3189_;
wire _3190_;
wire _3191_;
wire _3192_;
wire _3193_;
wire _3194_;
wire _3195_;
wire _3196_;
wire _3197_;
wire _3198_;
wire _3199_;
wire _3200_;
wire _3201_;
wire _3202_;
wire _3203_;
wire _3204_;
wire _3205_;
wire _3206_;
wire _3207_;
wire _3208_;
wire _3209_;
wire _3210_;
wire _3211_;
wire _3212_;
wire _3213_;
wire _3214_;
wire _3215_;
wire _3216_;
wire _3217_;
wire _3218_;
wire _3219_;
wire _3220_;
wire _3221_;
wire _3222_;
wire _3223_;
wire _3224_;
wire _3225_;
wire _3226_;
wire _3227_;
wire _3228_;
wire _3229_;
wire _3230_;
wire _3231_;
wire _3232_;
wire _3233_;
wire _3234_;
wire _3235_;
wire _3236_;
wire _3237_;
wire _3238_;
wire _3239_;
wire _3240_;
wire _3241_;
wire _3242_;
wire _3243_;
wire _3244_;
wire _3245_;
wire _3246_;
wire _3247_;
wire _3248_;
wire _3249_;
wire _3250_;
wire _3251_;
wire _3252_;
wire _3253_;
wire _3254_;
wire _3255_;
wire _3256_;
wire _3257_;
wire _3258_;
wire _3259_;
wire _3260_;
wire _3261_;
wire _3262_;
wire _3263_;
wire _3264_;
wire _3265_;
wire _3266_;
wire _3267_;
wire _3268_;
wire _3269_;
wire _3270_;
wire _3271_;
wire _3272_;
wire _3273_;
wire _3274_;
wire _3275_;
wire _3276_;
wire _3277_;
wire _3278_;
wire _3279_;
wire _3280_;
wire _3281_;
wire _3282_;
wire _3283_;
wire _3284_;
wire _3285_;
wire _3286_;
wire _3287_;
wire _3288_;
wire _3289_;
wire _3290_;
wire _3291_;
wire _3292_;
wire _3293_;
wire _3294_;
wire _3295_;
wire _3296_;
wire _3297_;
wire _3298_;
wire _3299_;
wire _3300_;
wire _3301_;
wire _3302_;
wire _3303_;
wire _3304_;
wire _3305_;
wire _3306_;
wire _3307_;
wire _3308_;
wire _3309_;
wire _3310_;
wire _3311_;
wire _3312_;
wire _3313_;
wire _3314_;
wire _3315_;
wire _3316_;
wire _3317_;
wire _3318_;
wire _3319_;
wire _3320_;
wire _3321_;
wire _3322_;
wire _3323_;
wire _3324_;
wire _3325_;
wire _3326_;
wire _3327_;
wire _3328_;
wire _3329_;
wire _3330_;
wire _3331_;
wire _3332_;
wire _3333_;
wire _3334_;
wire _3335_;
wire _3336_;
wire _3337_;
wire _3338_;
wire _3339_;
wire _3340_;
wire _3341_;
wire _3342_;
wire _3343_;
wire _3344_;
wire _3345_;
wire _3346_;
wire _3347_;
wire _3348_;
wire _3349_;
wire _3350_;
wire _3351_;
wire _3352_;
wire _3353_;
wire _3354_;
wire _3355_;
wire _3356_;
wire _3357_;
wire _3358_;
wire _3359_;
wire _3360_;
wire _3361_;
wire _3362_;
wire _3363_;
wire _3364_;
wire _3365_;
wire _3366_;
wire _3367_;
wire _3368_;
wire _3369_;
wire _3370_;
wire _3371_;
wire _3372_;
wire _3373_;
wire _3374_;
wire _3375_;
wire _3376_;
wire _3377_;
wire _3378_;
wire _3379_;
wire _3380_;
wire _3381_;
wire _3382_;
wire _3383_;
wire _3384_;
wire _3385_;
wire _3386_;
wire _3387_;
wire _3388_;
wire _3389_;
wire _3390_;
wire _3391_;
wire _3392_;
wire _3393_;
wire _3394_;
wire _3395_;
wire _3396_;
wire _3397_;
wire _3398_;
wire _3399_;
wire _3400_;
wire _3401_;
wire _3402_;
wire _3403_;
wire _3404_;
wire _3405_;
wire _3406_;
wire _3407_;
wire _3408_;
wire _3409_;
wire _3410_;
wire _3411_;
wire _3412_;
wire _3413_;
wire _3414_;
wire _3415_;
wire _3416_;
wire _3417_;
wire _3418_;
wire _3419_;
wire _3420_;
wire _3421_;
wire _3422_;
wire _3423_;
wire _3424_;
wire _3425_;
wire _3426_;
wire _3427_;
wire _3428_;
wire _3429_;
wire _3430_;
wire _3431_;
wire _3432_;
wire _3433_;
wire _3434_;
wire _3435_;
wire _3436_;
wire _3437_;
wire _3438_;
wire _3439_;
wire _3440_;
wire _3441_;
wire _3442_;
wire _3443_;
wire _3444_;
wire _3445_;
wire _3446_;
wire _3447_;
wire _3448_;
wire _3449_;
wire _3450_;
wire _3451_;
wire _3452_;
wire _3453_;
wire _3454_;
wire _3455_;
wire _3456_;
wire _3457_;
wire _3458_;
wire _3459_;
wire _3460_;
wire _3461_;
wire _3462_;
wire _3463_;
wire _3464_;
wire _3465_;
wire _3466_;
wire _3467_;
wire _3468_;
wire _3469_;
wire _3470_;
wire _3471_;
wire _3472_;
wire _3473_;
wire _3474_;
wire _3475_;
wire _3476_;
wire _3477_;
wire _3478_;
wire _3479_;
wire _3480_;
wire _3481_;
wire _3482_;
wire _3483_;
wire _3484_;
wire _3485_;
wire _3486_;
wire _3487_;
wire _3488_;
wire _3489_;
wire _3490_;
wire _3491_;
wire _3492_;
wire _3493_;
wire _3494_;
wire _3495_;
wire _3496_;
wire _3497_;
wire _3498_;
wire _3499_;
wire _3500_;
wire _3501_;
wire _3502_;
wire _3503_;
wire _3504_;
wire _3505_;
wire _3506_;
wire _3507_;
wire _3508_;
wire _3509_;
wire _3510_;
wire _3511_;
wire _3512_;
wire _3513_;
wire _3514_;
wire _3515_;
wire _3516_;
wire _3517_;
wire _3518_;
wire _3519_;
wire _3520_;
wire _3521_;
wire _3522_;
wire _3523_;
wire _3524_;
wire _3525_;
wire _3526_;
wire _3527_;
wire _3528_;
wire _3529_;
wire _3530_;
wire _3531_;
wire _3532_;
wire _3533_;
wire _3534_;
wire _3535_;
wire _3536_;
wire _3537_;
wire _3538_;
wire _3539_;
wire _3540_;
wire _3541_;
wire _3542_;
wire _3543_;
wire _3544_;
wire _3545_;
wire _3546_;
wire _3547_;
wire _3548_;
wire _3549_;
wire _3550_;
wire _3551_;
wire _3552_;
wire _3553_;
wire _3554_;
wire _3555_;
wire _3556_;
wire _3557_;
wire _3558_;
wire _3559_;
wire _3560_;
wire _3561_;
wire _3562_;
wire _3563_;
wire _3564_;
wire _3565_;
wire _3566_;
wire _3567_;
wire _3568_;
wire _3569_;
wire _3570_;
wire _3571_;
wire _3572_;
wire _3573_;
wire _3574_;
wire _3575_;
wire _3576_;
wire _3577_;
wire _3578_;
wire _3579_;
wire _3580_;
wire _3581_;
wire _3582_;
wire _3583_;
wire _3584_;
wire _3585_;
wire _3586_;
wire _3587_;
wire _3588_;
wire _3589_;
wire _3590_;
wire _3591_;
wire _3592_;
wire _3593_;
wire _3594_;
wire _3595_;
wire _3596_;
wire _3597_;
wire _3598_;
wire _3599_;
wire _3600_;
wire _3601_;
wire _3602_;
wire _3603_;
wire _3604_;
wire _3605_;
wire _3606_;
wire _3607_;
wire _3608_;
wire _3609_;
wire _3610_;
wire _3611_;
wire _3612_;
wire _3613_;
wire _3614_;
wire _3615_;
wire _3616_;
wire _3617_;
wire _3618_;
wire _3619_;
wire _3620_;
wire _3621_;
wire _3622_;
wire _3623_;
wire _3624_;
wire _3625_;
wire _3626_;
wire _3627_;
wire _3628_;
wire _3629_;
wire _3630_;
wire _3631_;
wire _3632_;
wire _3633_;
wire _3634_;
wire _3635_;
wire _3636_;
wire _3637_;
wire _3638_;
wire _3639_;
wire _3640_;
wire _3641_;
wire _3642_;
wire _3643_;
wire _3644_;
wire _3645_;
wire _3646_;
wire _3647_;
wire _3648_;
wire _3649_;
wire _3650_;
wire _3651_;
wire _3652_;
wire _3653_;
wire _3654_;
wire _3655_;
wire _3656_;
wire _3657_;
wire _3658_;
wire _3659_;
wire _3660_;
wire _3661_;
wire _3662_;
wire _3663_;
wire _3664_;
wire _3665_;
wire _3666_;
wire _3667_;
wire _3668_;
wire _3669_;
wire _3670_;
wire _3671_;
wire _3672_;
wire _3673_;
wire _3674_;
wire _3675_;
wire _3676_;
wire _3677_;
wire _3678_;
wire _3679_;
wire _3680_;
wire _3681_;
wire _3682_;
wire _3683_;
wire _3684_;
wire _3685_;
wire _3686_;
wire _3687_;
wire _3688_;
wire _3689_;
wire _3690_;
wire _3691_;
wire _3692_;
wire _3693_;
wire _3694_;
wire _3695_;
wire _3696_;
wire _3697_;
wire _3698_;
wire _3699_;
wire _3700_;
wire _3701_;
wire _3702_;
wire _3703_;
wire _3704_;
wire _3705_;
wire _3706_;
wire _3707_;
wire _3708_;
wire _3709_;
wire _3710_;
wire _3711_;
wire _3712_;
wire _3713_;
wire _3714_;
wire _3715_;
wire _3716_;
wire _3717_;
wire _3718_;
wire _3719_;
wire _3720_;
wire _3721_;
wire _3722_;
wire _3723_;
wire _3724_;
wire _3725_;
wire _3726_;
wire _3727_;
wire _3728_;
wire _3729_;
wire _3730_;
wire _3731_;
wire _3732_;
wire _3733_;
wire _3734_;
wire _3735_;
wire _3736_;
wire _3737_;
wire _3738_;
wire _3739_;
wire _3740_;
wire _3741_;
wire _3742_;
wire _3743_;
wire _3744_;
wire _3745_;
wire _3746_;
wire _3747_;
wire _3748_;
wire _3749_;
wire _3750_;
wire _3751_;
wire _3752_;
wire _3753_;
wire _3754_;
wire _3755_;
wire _3756_;
wire _3757_;
wire _3758_;
wire _3759_;
wire _3760_;
wire _3761_;
wire _3762_;
wire _3763_;
wire _3764_;
wire _3765_;
wire _3766_;
wire _3767_;
wire _3768_;
wire _3769_;
wire _3770_;
wire _3771_;
wire _3772_;
wire _3773_;
wire _3774_;
wire _3775_;
wire _3776_;
wire _3777_;
wire _3778_;
wire _3779_;
wire _3780_;
wire _3781_;
wire _3782_;
wire _3783_;
wire _3784_;
wire _3785_;
wire _3786_;
wire _3787_;
wire _3788_;
wire _3789_;
wire _3790_;
wire _3791_;
wire _3792_;
wire _3793_;
wire _3794_;
wire _3795_;
wire _3796_;
wire _3797_;
wire _3798_;
wire _3799_;
wire _3800_;
wire _3801_;
wire _3802_;
wire _3803_;
wire _3804_;
wire _3805_;
wire _3806_;
wire _3807_;
wire _3808_;
wire _3809_;
wire _3810_;
wire _3811_;
wire _3812_;
wire _3813_;
wire _3814_;
wire _3815_;
wire _3816_;
wire _3817_;
wire _3818_;
wire _3819_;
wire _3820_;
wire _3821_;
wire _3822_;
wire _3823_;
wire _3824_;
wire _3825_;
wire _3826_;
wire _3827_;
wire _3828_;
wire _3829_;
wire _3830_;
wire _3831_;
wire _3832_;
wire _3833_;
wire _3834_;
wire _3835_;
wire _3836_;
wire _3837_;
wire _3838_;
wire _3839_;
wire _3840_;
wire _3841_;
wire _3842_;
wire _3843_;
wire _3844_;
wire _3845_;
wire _3846_;
wire _3847_;
wire _3848_;
wire _3849_;
wire _3850_;
wire _3851_;
wire _3852_;
wire _3853_;
wire _3854_;
wire _3855_;
wire _3856_;
wire _3857_;
wire _3858_;
wire _3859_;
wire _3860_;
wire _3861_;
wire _3862_;
wire _3863_;
wire _3864_;
wire _3865_;
wire _3866_;
wire _3867_;
wire _3868_;
wire _3869_;
wire _3870_;
wire _3871_;
wire _3872_;
wire _3873_;
wire _3874_;
wire _3875_;
wire _3876_;
wire _3877_;
wire _3878_;
wire _3879_;
wire _3880_;
wire _3881_;
wire _3882_;
wire _3883_;
wire _3884_;
wire _3885_;
wire _3886_;
wire _3887_;
wire _3888_;
wire _3889_;
wire _3890_;
wire _3891_;
wire _3892_;
wire _3893_;
wire _3894_;
wire _3895_;
wire _3896_;
wire _3897_;
wire _3898_;
wire _3899_;
wire _3900_;
wire _3901_;
wire _3902_;
wire _3903_;
wire _3904_;
wire _3905_;
wire _3906_;
wire _3907_;
wire _3908_;
wire _3909_;
wire _3910_;
wire _3911_;
wire _3912_;
wire _3913_;
wire _3914_;
wire _3915_;
wire _3916_;
wire _3917_;
wire _3918_;
wire _3919_;
wire _3920_;
wire _3921_;
wire _3922_;
wire _3923_;
wire _3924_;
wire _3925_;
wire _3926_;
wire _3927_;
wire _3928_;
wire _3929_;
wire _3930_;
wire _3931_;
wire _3932_;
wire _3933_;
wire _3934_;
wire _3935_;
wire _3936_;
wire _3937_;
wire _3938_;
wire _3939_;
wire _3940_;
wire _3941_;
wire _3942_;
wire _3943_;
wire _3944_;
wire _3945_;
wire _3946_;
wire _3947_;
wire _3948_;
wire _3949_;
wire _3950_;
wire _3951_;
wire _3952_;
wire _3953_;
wire _3954_;
wire _3955_;
wire _3956_;
wire _3957_;
wire _3958_;
wire _3959_;
wire _3960_;
wire _3961_;
wire _3962_;
wire _3963_;
wire _3964_;
wire _3965_;
wire _3966_;
wire _3967_;
wire _3968_;
wire _3969_;
wire _3970_;
wire _3971_;
wire _3972_;
wire _3973_;
wire _3974_;
wire _3975_;
wire _3976_;
wire _3977_;
wire _3978_;
wire _3979_;
wire _3980_;
wire _3981_;
wire _3982_;
wire _3983_;
wire _3984_;
wire _3985_;
wire _3986_;
wire _3987_;
wire _3988_;
wire _3989_;
wire _3990_;
wire _3991_;
wire _3992_;
wire _3993_;
wire _3994_;
wire _3995_;
wire _3996_;
wire _3997_;
wire _3998_;
wire _3999_;
wire _4000_;
wire _4001_;
wire _4002_;
wire _4003_;
wire _4004_;
wire _4005_;
wire _4006_;
wire _4007_;
wire _4008_;
wire _4009_;
wire _4010_;
wire _4011_;
wire _4012_;
wire _4013_;
wire _4014_;
wire _4015_;
wire _4016_;
wire _4017_;
wire _4018_;
wire _4019_;
wire _4020_;
wire _4021_;
wire _4022_;
wire _4023_;
wire _4024_;
wire _4025_;
wire _4026_;
wire _4027_;
wire _4028_;
wire _4029_;
wire _4030_;
wire _4031_;
wire _4032_;
wire _4033_;
wire _4034_;
wire _4035_;
wire _4036_;
wire _4037_;
wire _4038_;
wire _4039_;
wire _4040_;
wire _4041_;
wire _4042_;
wire _4043_;
wire _4044_;
wire _4045_;
wire _4046_;
wire _4047_;
wire _4048_;
wire _4049_;
wire _4050_;
wire _4051_;
wire _4052_;
wire _4053_;
wire _4054_;
wire _4055_;
wire _4056_;
wire _4057_;
wire _4058_;
wire _4059_;
wire _4060_;
wire _4061_;
wire _4062_;
wire _4063_;
wire _4064_;
wire _4065_;
wire _4066_;
wire _4067_;
wire _4068_;
wire _4069_;
wire _4070_;
wire _4071_;
wire _4072_;
wire _4073_;
wire _4074_;
wire _4075_;
wire _4076_;
wire _4077_;
wire _4078_;
wire _4079_;
wire _4080_;
wire _4081_;
wire _4082_;
wire _4083_;
wire _4084_;
wire _4085_;
wire _4086_;
wire _4087_;
wire _4088_;
wire _4089_;
wire _4090_;
wire _4091_;
wire _4092_;
wire _4093_;
wire _4094_;
wire _4095_;
wire _4096_;
wire _4097_;
wire _4098_;
wire _4099_;
wire _4100_;
wire _4101_;
wire _4102_;
wire _4103_;
wire _4104_;
wire _4105_;
wire _4106_;
wire _4107_;
wire _4108_;
wire _4109_;
wire _4110_;
wire _4111_;
wire _4112_;
wire _4113_;
wire _4114_;
wire _4115_;
wire _4116_;
wire _4117_;
wire _4118_;
wire _4119_;
wire _4120_;
wire _4121_;
wire _4122_;
wire _4123_;
wire _4124_;
wire _4125_;
wire _4126_;
wire _4127_;
wire _4128_;
wire _4129_;
wire _4130_;
wire _4131_;
wire _4132_;
wire _4133_;
wire _4134_;
wire _4135_;
wire _4136_;
wire _4137_;
wire _4138_;
wire _4139_;
wire _4140_;
wire _4141_;
wire _4142_;
wire _4143_;
wire _4144_;
wire _4145_;
wire _4146_;
wire _4147_;
wire _4148_;
wire _4149_;
wire _4150_;
wire _4151_;
wire _4152_;
wire _4153_;
wire _4154_;
wire _4155_;
wire _4156_;
wire _4157_;
wire _4158_;
wire _4159_;
wire _4160_;
wire _4161_;
wire _4162_;
wire _4163_;
wire _4164_;
wire _4165_;
wire _4166_;
wire _4167_;
wire _4168_;
wire _4169_;
wire _4170_;
wire _4171_;
wire _4172_;
wire _4173_;
wire _4174_;
wire _4175_;
wire _4176_;
wire _4177_;
wire _4178_;
wire _4179_;
wire _4180_;
wire _4181_;
wire _4182_;
wire _4183_;
wire _4184_;
wire _4185_;
wire _4186_;
wire _4187_;
wire _4188_;
wire _4189_;
wire _4190_;
wire _4191_;
wire _4192_;
wire _4193_;
wire _4194_;
wire _4195_;
wire _4196_;
wire _4197_;
wire _4198_;
wire _4199_;
wire _4200_;
wire _4201_;
wire _4202_;
wire _4203_;
wire _4204_;
wire _4205_;
wire _4206_;
wire _4207_;
wire _4208_;
wire _4209_;
wire _4210_;
wire _4211_;
wire _4212_;
wire _4213_;
wire _4214_;
wire _4215_;
wire _4216_;
wire _4217_;
wire _4218_;
wire _4219_;
wire _4220_;
wire _4221_;
wire _4222_;
wire _4223_;
wire _4224_;
wire _4225_;
wire _4226_;
wire _4227_;
wire _4228_;
wire _4229_;
wire _4230_;
wire _4231_;
wire _4232_;
wire _4233_;
wire _4234_;
wire _4235_;
wire _4236_;
wire _4237_;
wire _4238_;
wire _4239_;
wire _4240_;
wire _4241_;
wire _4242_;
wire _4243_;
wire _4244_;
wire _4245_;
wire _4246_;
wire _4247_;
wire _4248_;
wire _4249_;
wire _4250_;
wire _4251_;
wire _4252_;
wire _4253_;
wire _4254_;
wire _4255_;
wire _4256_;
wire _4257_;
wire _4258_;
wire _4259_;
wire _4260_;
wire _4261_;
wire _4262_;
wire _4263_;
wire _4264_;
wire _4265_;
wire _4266_;
wire _4267_;
wire _4268_;
wire _4269_;
wire _4270_;
wire _4271_;
wire _4272_;
wire _4273_;
wire _4274_;
wire _4275_;
wire _4276_;
wire _4277_;
wire _4278_;
wire _4279_;
wire _4280_;
wire _4281_;
wire _4282_;
wire _4283_;
wire _4284_;
wire _4285_;
wire _4286_;
wire _4287_;
wire _4288_;
wire _4289_;
wire _4290_;
wire _4291_;
wire _4292_;
wire _4293_;
wire _4294_;
wire _4295_;
wire _4296_;
wire _4297_;
wire _4298_;
wire _4299_;
wire _4300_;
wire _4301_;
wire _4302_;
wire _4303_;
wire _4304_;
wire _4305_;
wire _4306_;
wire _4307_;
wire _4308_;
wire _4309_;
wire _4310_;
wire _4311_;
wire _4312_;
wire _4313_;
wire _4314_;
wire _4315_;
wire _4316_;
wire _4317_;
wire _4318_;
wire _4319_;
wire _4320_;
wire _4321_;
wire _4322_;
wire _4323_;
wire _4324_;
wire _4325_;
wire _4326_;
wire _4327_;
wire _4328_;
wire _4329_;
wire _4330_;
wire _4331_;
wire _4332_;
wire _4333_;
wire _4334_;
wire _4335_;
wire _4336_;
wire _4337_;
wire _4338_;
wire _4339_;
wire _4340_;
wire _4341_;
wire _4342_;
wire _4343_;
wire _4344_;
wire _4345_;
wire _4346_;
wire _4347_;
wire _4348_;
wire _4349_;
wire _4350_;
wire _4351_;
wire _4352_;
wire _4353_;
wire _4354_;
wire _4355_;
wire _4356_;
wire _4357_;
wire _4358_;
wire _4359_;
wire _4360_;
wire _4361_;
wire _4362_;
wire _4363_;
wire _4364_;
wire _4365_;
wire _4366_;
wire _4367_;
wire _4368_;
wire _4369_;
wire _4370_;
wire _4371_;
wire _4372_;
wire _4373_;
wire _4374_;
wire _4375_;
wire _4376_;
wire _4377_;
wire _4378_;
wire _4379_;
wire _4380_;
wire _4381_;
wire _4382_;
wire _4383_;
wire _4384_;
wire _4385_;
wire _4386_;
wire _4387_;
wire _4388_;
wire _4389_;
wire _4390_;
wire _4391_;
wire _4392_;
wire _4393_;
wire _4394_;
wire _4395_;
wire _4396_;
wire _4397_;
wire _4398_;
wire _4399_;
wire _4400_;
wire _4401_;
wire _4402_;
wire _4403_;
wire _4404_;
wire _4405_;
wire _4406_;
wire _4407_;
wire _4408_;
wire _4409_;
wire _4410_;
wire _4411_;
wire _4412_;
wire _4413_;
wire _4414_;
wire _4415_;
wire _4416_;
wire _4417_;
wire _4418_;
wire _4419_;
wire _4420_;
wire _4421_;
wire _4422_;
wire _4423_;
wire _4424_;
wire _4425_;
wire _4426_;
wire _4427_;
wire _4428_;
wire _4429_;
wire _4430_;
wire _4431_;
wire _4432_;
wire _4433_;
wire _4434_;
wire _4435_;
wire _4436_;
wire _4437_;
wire _4438_;
wire _4439_;
wire _4440_;
wire _4441_;
wire _4442_;
wire _4443_;
wire _4444_;
wire _4445_;
wire _4446_;
wire _4447_;
wire _4448_;
wire _4449_;
wire _4450_;
wire _4451_;
wire _4452_;
wire _4453_;
wire _4454_;
wire _4455_;
wire _4456_;
wire _4457_;
wire _4458_;
wire _4459_;
wire _4460_;
wire _4461_;
wire _4462_;
wire _4463_;
wire _4464_;
wire _4465_;
wire _4466_;
wire _4467_;
wire _4468_;
wire _4469_;
wire _4470_;
wire _4471_;
wire _4472_;
wire _4473_;
wire _4474_;
wire _4475_;
wire _4476_;
wire _4477_;
wire _4478_;
wire _4479_;
wire _4480_;
wire _4481_;
wire _4482_;
wire _4483_;
wire _4484_;
wire _4485_;
wire _4486_;
wire _4487_;
wire _4488_;
wire _4489_;
wire _4490_;
wire _4491_;
wire _4492_;
wire _4493_;
wire _4494_;
wire _4495_;
wire _4496_;
wire _4497_;
wire _4498_;
wire _4499_;
wire _4500_;
wire _4501_;
wire _4502_;
wire _4503_;
wire _4504_;
wire _4505_;
wire _4506_;
wire _4507_;
wire _4508_;
wire _4509_;
wire _4510_;
wire _4511_;
wire _4512_;
wire _4513_;
wire _4514_;
wire _4515_;
wire _4516_;
wire _4517_;
wire _4518_;
wire _4519_;
wire _4520_;
wire _4521_;
wire _4522_;
wire _4523_;
wire _4524_;
wire _4525_;
wire _4526_;
wire _4527_;
wire _4528_;
wire _4529_;
wire _4530_;
wire _4531_;
wire _4532_;
wire _4533_;
wire _4534_;
wire _4535_;
wire _4536_;
wire _4537_;
wire _4538_;
wire _4539_;
wire _4540_;
wire _4541_;
wire _4542_;
wire _4543_;
wire _4544_;
wire _4545_;
wire _4546_;
wire _4547_;
wire _4548_;
wire _4549_;
wire _4550_;
wire _4551_;
wire _4552_;
wire _4553_;
wire _4554_;
wire _4555_;
wire _4556_;
wire _4557_;
wire _4558_;
wire _4559_;
wire _4560_;
wire _4561_;
wire _4562_;
wire _4563_;
wire _4564_;
wire _4565_;
wire _4566_;
wire _4567_;
wire _4568_;
wire _4569_;
wire _4570_;
wire _4571_;
wire _4572_;
wire _4573_;
wire _4574_;
wire _4575_;
wire _4576_;
wire _4577_;
wire _4578_;
wire _4579_;
wire _4580_;
wire _4581_;
wire _4582_;
wire _4583_;
wire _4584_;
wire _4585_;
wire _4586_;
wire _4587_;
wire _4588_;
wire _4589_;
wire _4590_;
wire _4591_;
wire _4592_;
wire _4593_;
wire _4594_;
wire _4595_;
wire _4596_;
wire _4597_;
wire _4598_;
wire _4599_;
wire _4600_;
wire _4601_;
wire _4602_;
wire _4603_;
wire _4604_;
wire _4605_;
wire _4606_;
wire _4607_;
wire _4608_;
wire _4609_;
wire _4610_;
wire _4611_;
wire _4612_;
wire _4613_;
wire _4614_;
wire _4615_;
wire _4616_;
wire _4617_;
wire _4618_;
wire _4619_;
wire _4620_;
wire _4621_;
wire _4622_;
wire _4623_;
wire _4624_;
wire _4625_;
wire _4626_;
wire _4627_;
wire _4628_;
wire _4629_;
wire _4630_;
wire _4631_;
wire _4632_;
wire _4633_;
wire _4634_;
wire _4635_;
wire _4636_;
wire _4637_;
wire _4638_;
wire _4639_;
wire _4640_;
wire _4641_;
wire _4642_;
wire _4643_;
wire _4644_;
wire _4645_;
wire _4646_;
wire _4647_;
wire _4648_;
wire _4649_;
wire _4650_;
wire _4651_;
wire _4652_;
wire _4653_;
wire _4654_;
wire _4655_;
wire _4656_;
wire _4657_;
wire _4658_;
wire _4659_;
wire _4660_;
wire _4661_;
wire _4662_;
wire _4663_;
wire _4664_;
wire _4665_;
wire _4666_;
wire _4667_;
wire _4668_;
wire _4669_;
wire _4670_;
wire _4671_;
wire _4672_;
wire _4673_;
wire _4674_;
wire _4675_;
wire _4676_;
wire _4677_;
wire _4678_;
wire _4679_;
wire _4680_;
wire _4681_;
wire _4682_;
wire _4683_;
wire _4684_;
wire _4685_;
wire _4686_;
wire _4687_;
wire _4688_;
wire _4689_;
wire _4690_;
wire _4691_;
wire _4692_;
wire _4693_;
wire _4694_;
wire _4695_;
wire _4696_;
wire _4697_;
wire _4698_;
wire _4699_;
wire _4700_;
wire _4701_;
wire _4702_;
wire _4703_;
wire _4704_;
wire _4705_;
wire _4706_;
wire _4707_;
wire _4708_;
wire _4709_;
wire _4710_;
wire _4711_;
wire _4712_;
wire _4713_;
wire _4714_;
wire _4715_;
wire _4716_;
wire _4717_;
wire _4718_;
wire _4719_;
wire _4720_;
wire _4721_;
wire _4722_;
wire _4723_;
wire _4724_;
wire _4725_;
wire _4726_;
wire _4727_;
wire _4728_;
wire _4729_;
wire _4730_;
wire _4731_;
wire _4732_;
wire _4733_;
wire _4734_;
wire _4735_;
wire _4736_;
wire _4737_;
wire _4738_;
wire _4739_;
wire _4740_;
wire _4741_;
wire _4742_;
wire _4743_;
wire _4744_;
wire _4745_;
wire _4746_;
wire _4747_;
wire _4748_;
wire _4749_;
wire _4750_;
wire _4751_;
wire _4752_;
wire _4753_;
wire _4754_;
wire _4755_;
wire _4756_;
wire _4757_;
wire _4758_;
wire _4759_;
wire _4760_;
wire _4761_;
wire _4762_;
wire _4763_;
wire _4764_;
wire _4765_;
wire _4766_;
wire _4767_;
wire _4768_;
wire _4769_;
wire _4770_;
wire _4771_;
wire _4772_;
wire _4773_;
wire _4774_;
wire _4775_;
wire _4776_;
wire _4777_;
wire _4778_;
wire _4779_;
wire _4780_;
wire _4781_;
wire _4782_;
wire _4783_;
wire _4784_;
wire _4785_;
wire _4786_;
wire _4787_;
wire _4788_;
wire _4789_;
wire _4790_;
wire _4791_;
wire _4792_;
wire _4793_;
wire _4794_;
wire _4795_;
wire _4796_;
wire _4797_;
wire _4798_;
wire _4799_;
wire _4800_;
wire _4801_;
wire _4802_;
wire _4803_;
wire _4804_;
wire _4805_;
wire _4806_;
wire _4807_;
wire _4808_;
wire _4809_;
wire _4810_;
wire _4811_;
wire _4812_;
wire _4813_;
wire _4814_;
wire _4815_;
wire _4816_;
wire _4817_;
wire _4818_;
wire _4819_;
wire _4820_;
wire _4821_;
wire _4822_;
wire _4823_;
wire _4824_;
wire _4825_;
wire _4826_;
wire _4827_;
wire _4828_;
wire _4829_;
wire _4830_;
wire _4831_;
wire _4832_;
wire _4833_;
wire _4834_;
wire _4835_;
wire _4836_;
wire _4837_;
wire _4838_;
wire _4839_;
wire _4840_;
wire _4841_;
wire _4842_;
wire _4843_;
wire _4844_;
wire _4845_;
wire _4846_;
wire _4847_;
wire _4848_;
wire _4849_;
wire _4850_;
wire _4851_;
wire _4852_;
wire _4853_;
wire _4854_;
wire _4855_;
wire _4856_;
wire _4857_;
wire _4858_;
wire _4859_;
wire _4860_;
wire _4861_;
wire _4862_;
wire _4863_;
wire _4864_;
wire _4865_;
wire _4866_;
wire _4867_;
wire _4868_;
wire _4869_;
wire _4870_;
wire _4871_;
wire _4872_;
wire _4873_;
wire _4874_;
wire _4875_;
wire _4876_;
wire _4877_;
wire _4878_;
wire _4879_;
wire _4880_;
wire _4881_;
wire _4882_;
wire _4883_;
wire _4884_;
wire _4885_;
wire _4886_;
wire _4887_;
wire _4888_;
wire _4889_;
wire _4890_;
wire _4891_;
wire _4892_;
wire _4893_;
wire _4894_;
wire _4895_;
wire _4896_;
wire _4897_;
wire _4898_;
wire _4899_;
wire _4900_;
wire _4901_;
wire _4902_;
wire _4903_;
wire _4904_;
wire _4905_;
wire _4906_;
wire _4907_;
wire _4908_;
wire _4909_;
wire _4910_;
wire _4911_;
wire _4912_;
wire _4913_;
wire _4914_;
wire _4915_;
wire _4916_;
wire _4917_;
wire _4918_;
wire _4919_;
wire _4920_;
wire _4921_;
wire _4922_;
wire _4923_;
wire _4924_;
wire _4925_;
wire _4926_;
wire _4927_;
wire _4928_;
wire _4929_;
wire _4930_;
wire _4931_;
wire _4932_;
wire _4933_;
wire _4934_;
wire _4935_;
wire _4936_;
wire _4937_;
wire _4938_;
wire _4939_;
wire _4940_;
wire _4941_;
wire _4942_;
wire _4943_;
wire _4944_;
wire _4945_;
wire _4946_;
wire _4947_;
wire _4948_;
wire _4949_;
wire _4950_;
wire _4951_;
wire _4952_;
wire _4953_;
wire _4954_;
wire _4955_;
wire _4956_;
wire _4957_;
wire _4958_;
wire _4959_;
wire _4960_;
wire _4961_;
wire _4962_;
wire _4963_;
wire _4964_;
wire _4965_;
wire _4966_;
wire _4967_;
wire _4968_;
wire _4969_;
wire _4970_;
wire _4971_;
wire _4972_;
wire _4973_;
wire _4974_;
wire _4975_;
wire _4976_;
wire _4977_;
wire _4978_;
wire _4979_;
wire _4980_;
wire _4981_;
wire _4982_;
wire _4983_;
wire _4984_;
wire _4985_;
wire _4986_;
wire _4987_;
wire _4988_;
wire _4989_;
wire _4990_;
wire _4991_;
wire _4992_;
wire _4993_;
wire _4994_;
wire _4995_;
wire _4996_;
wire _4997_;
wire _4998_;
wire _4999_;
wire _5000_;
wire _5001_;
wire _5002_;
wire _5003_;
wire _5004_;
wire _5005_;
wire _5006_;
wire _5007_;
wire _5008_;
wire _5009_;
wire _5010_;
wire _5011_;
wire _5012_;
wire _5013_;
wire _5014_;
wire _5015_;
wire _5016_;
wire _5017_;
wire _5018_;
wire _5019_;
wire _5020_;
wire _5021_;
wire _5022_;
wire _5023_;
wire _5024_;
wire _5025_;
wire _5026_;
wire _5027_;
wire _5028_;
wire _5029_;
wire _5030_;
wire _5031_;
wire _5032_;
wire _5033_;
wire _5034_;
wire _5035_;
wire _5036_;
wire _5037_;
wire _5038_;
wire _5039_;
wire _5040_;
wire _5041_;
wire _5042_;
wire _5043_;
wire _5044_;
wire _5045_;
wire _5046_;
wire _5047_;
wire _5048_;
wire _5049_;
wire _5050_;
wire _5051_;
wire _5052_;
wire _5053_;
wire _5054_;
wire _5055_;
wire _5056_;
wire _5057_;
wire _5058_;
wire _5059_;
wire _5060_;
wire _5061_;
wire _5062_;
wire _5063_;
wire _5064_;
wire _5065_;
wire _5066_;
wire _5067_;
wire _5068_;
wire _5069_;
wire _5070_;
wire _5071_;
wire _5072_;
wire _5073_;
wire _5074_;
wire _5075_;
wire _5076_;
wire _5077_;
wire _5078_;
wire _5079_;
wire _5080_;
wire _5081_;
wire _5082_;
wire _5083_;
wire _5084_;
wire _5085_;
wire _5086_;
wire _5087_;
wire _5088_;
wire _5089_;
wire _5090_;
wire _5091_;
wire _5092_;
wire _5093_;
wire _5094_;
wire _5095_;
wire _5096_;
wire _5097_;
wire _5098_;
wire _5099_;
wire _5100_;
wire _5101_;
wire _5102_;
wire _5103_;
wire _5104_;
wire _5105_;
wire _5106_;
wire _5107_;
wire _5108_;
wire _5109_;
wire _5110_;
wire _5111_;
wire _5112_;
wire _5113_;
wire _5114_;
wire _5115_;
wire _5116_;
wire _5117_;
wire _5118_;
wire _5119_;
wire _5120_;
wire _5121_;
wire _5122_;
wire _5123_;
wire _5124_;
wire _5125_;
wire _5126_;
wire _5127_;
wire _5128_;
wire _5129_;
wire _5130_;
wire _5131_;
wire _5132_;
wire _5133_;
wire _5134_;
wire _5135_;
wire _5136_;
wire _5137_;
wire _5138_;
wire _5139_;
wire _5140_;
wire _5141_;
wire _5142_;
wire _5143_;
wire _5144_;
wire _5145_;
wire _5146_;
wire _5147_;
wire _5148_;
wire _5149_;
wire _5150_;
wire _5151_;
wire _5152_;
wire _5153_;
wire _5154_;
wire _5155_;
wire _5156_;
wire _5157_;
wire _5158_;
wire _5159_;
wire _5160_;
wire _5161_;
wire _5162_;
wire _5163_;
wire _5164_;
wire _5165_;
wire _5166_;
wire _5167_;
wire _5168_;
wire _5169_;
wire _5170_;
wire _5171_;
wire _5172_;
wire _5173_;
wire _5174_;
wire _5175_;
wire _5176_;
wire _5177_;
wire _5178_;
wire _5179_;
wire _5180_;
wire _5181_;
wire _5182_;
wire _5183_;
wire _5184_;
wire _5185_;
wire _5186_;
wire _5187_;
wire _5188_;
wire _5189_;
wire _5190_;
wire _5191_;
wire _5192_;
wire _5193_;
wire _5194_;
wire _5195_;
wire _5196_;
wire _5197_;
wire _5198_;
wire _5199_;
wire _5200_;
wire _5201_;
wire _5202_;
wire _5203_;
wire _5204_;
wire _5205_;
wire _5206_;
wire _5207_;
wire _5208_;
wire _5209_;
wire _5210_;
wire _5211_;
wire _5212_;
wire _5213_;
wire _5214_;
wire _5215_;
wire _5216_;
wire _5217_;
wire _5218_;
wire _5219_;
wire _5220_;
wire _5221_;
wire _5222_;
wire _5223_;
wire _5224_;
wire _5225_;
wire _5226_;
wire _5227_;
wire _5228_;
wire _5229_;
wire _5230_;
wire _5231_;
wire _5232_;
wire _5233_;
wire _5234_;
wire _5235_;
wire _5236_;
wire _5237_;
wire _5238_;
wire _5239_;
wire _5240_;
wire _5241_;
wire _5242_;
wire _5243_;
wire _5244_;
wire _5245_;
wire _5246_;
wire _5247_;
wire _5248_;
wire _5249_;
wire _5250_;
wire _5251_;
wire _5252_;
wire _5253_;
wire _5254_;
wire _5255_;
wire _5256_;
wire _5257_;
wire _5258_;
wire _5259_;
wire _5260_;
wire _5261_;
wire _5262_;
wire _5263_;
wire _5264_;
wire _5265_;
wire _5266_;
wire _5267_;
wire _5268_;
wire _5269_;
wire _5270_;
wire _5271_;
wire _5272_;
wire _5273_;
wire _5274_;
wire _5275_;
wire _5276_;
wire _5277_;
wire _5278_;
wire _5279_;
wire _5280_;
wire _5281_;
wire _5282_;
wire _5283_;
wire _5284_;
wire _5285_;
wire _5286_;
wire _5287_;
wire _5288_;
wire _5289_;
wire _5290_;
wire _5291_;
wire _5292_;
wire _5293_;
wire _5294_;
wire _5295_;
wire _5296_;
wire _5297_;
wire _5298_;
wire _5299_;
wire _5300_;
wire _5301_;
wire _5302_;
wire _5303_;
wire _5304_;
wire _5305_;
wire _5306_;
wire _5307_;
wire _5308_;
wire _5309_;
wire _5310_;
wire _5311_;
wire _5312_;
wire _5313_;
wire _5314_;
wire _5315_;
wire _5316_;
wire _5317_;
wire _5318_;
wire _5319_;
wire _5320_;
wire _5321_;
wire _5322_;
wire _5323_;
wire _5324_;
wire _5325_;
wire _5326_;
wire _5327_;
wire _5328_;
wire _5329_;
wire _5330_;
wire _5331_;
wire _5332_;
wire _5333_;
wire _5334_;
wire _5335_;
wire _5336_;
wire _5337_;
wire _5338_;
wire _5339_;
wire _5340_;
wire _5341_;
wire _5342_;
wire _5343_;
wire _5344_;
wire _5345_;
wire _5346_;
wire _5347_;
wire _5348_;
wire _5349_;
wire _5350_;
wire _5351_;
wire _5352_;
wire _5353_;
wire _5354_;
wire _5355_;
wire _5356_;
wire _5357_;
wire _5358_;
wire _5359_;
wire _5360_;
wire _5361_;
wire _5362_;
wire _5363_;
wire _5364_;
wire _5365_;
wire _5366_;
wire _5367_;
wire _5368_;
wire _5369_;
wire _5370_;
wire _5371_;
wire _5372_;
wire _5373_;
wire _5374_;
wire _5375_;
wire _5376_;
wire _5377_;
wire _5378_;
wire _5379_;
wire _5380_;
wire _5381_;
wire _5382_;
wire _5383_;
wire _5384_;
wire _5385_;
wire _5386_;
wire _5387_;
wire _5388_;
wire _5389_;
wire _5390_;
wire _5391_;
wire _5392_;
wire _5393_;
wire _5394_;
wire _5395_;
wire _5396_;
wire _5397_;
wire _5398_;
wire _5399_;
wire _5400_;
wire _5401_;
wire _5402_;
wire _5403_;
wire _5404_;
wire _5405_;
wire _5406_;
wire _5407_;
wire _5408_;
wire _5409_;
wire _5410_;
wire _5411_;
wire _5412_;
wire _5413_;
wire _5414_;
wire _5415_;
wire _5416_;
wire _5417_;
wire _5418_;
wire _5419_;
wire _5420_;
wire _5421_;
wire _5422_;
wire _5423_;
wire _5424_;
wire _5425_;
wire _5426_;
wire _5427_;
wire _5428_;
wire _5429_;
wire _5430_;
wire _5431_;
wire _5432_;
wire _5433_;
wire _5434_;
wire _5435_;
wire _5436_;
wire _5437_;
wire _5438_;
wire _5439_;
wire _5440_;
wire _5441_;
wire _5442_;
wire _5443_;
wire _5444_;
wire _5445_;
wire _5446_;
wire _5447_;
wire _5448_;
wire _5449_;
wire _5450_;
wire _5451_;
wire _5452_;
wire _5453_;
wire _5454_;
wire _5455_;
wire _5456_;
wire _5457_;
wire _5458_;
wire _5459_;
wire _5460_;
wire _5461_;
wire _5462_;
wire _5463_;
wire _5464_;
wire _5465_;
wire _5466_;
wire _5467_;
wire _5468_;
wire _5469_;
wire _5470_;
wire _5471_;
wire _5472_;
wire _5473_;
wire _5474_;
wire _5475_;
wire _5476_;
wire _5477_;
wire _5478_;
wire _5479_;
wire _5480_;
wire _5481_;
wire _5482_;
wire _5483_;
wire _5484_;
wire _5485_;
wire _5486_;
wire _5487_;
wire _5488_;
wire _5489_;
wire _5490_;
wire _5491_;
wire _5492_;
wire _5493_;
wire _5494_;
wire _5495_;
wire _5496_;
wire _5497_;
wire _5498_;
wire _5499_;
wire _5500_;
wire _5501_;
wire _5502_;
wire _5503_;
wire _5504_;
wire _5505_;
wire _5506_;
wire _5507_;
wire _5508_;
wire _5509_;
wire _5510_;
wire _5511_;
wire _5512_;
wire _5513_;
wire _5514_;
wire _5515_;
wire _5516_;
wire _5517_;
wire _5518_;
wire _5519_;
wire _5520_;
wire _5521_;
wire _5522_;
wire _5523_;
wire _5524_;
wire _5525_;
wire _5526_;
wire _5527_;
wire _5528_;
wire _5529_;
wire _5530_;
wire _5531_;
wire _5532_;
wire _5533_;
wire _5534_;
wire _5535_;
wire _5536_;
wire _5537_;
wire _5538_;
wire _5539_;
wire _5540_;
wire _5541_;
wire _5542_;
wire _5543_;
wire _5544_;
wire _5545_;
wire _5546_;
wire _5547_;
wire _5548_;
wire _5549_;
wire _5550_;
wire _5551_;
wire _5552_;
wire _5553_;
wire _5554_;
wire _5555_;
wire _5556_;
wire _5557_;
wire _5558_;
wire _5559_;
wire _5560_;
wire _5561_;
wire _5562_;
wire _5563_;
wire _5564_;
wire _5565_;
wire _5566_;
wire _5567_;
wire _5568_;
wire _5569_;
wire _5570_;
wire _5571_;
wire _5572_;
wire _5573_;
wire _5574_;
wire _5575_;
wire _5576_;
wire _5577_;
wire _5578_;
wire _5579_;
wire _5580_;
wire _5581_;
wire _5582_;
wire _5583_;
wire _5584_;
wire _5585_;
wire _5586_;
wire _5587_;
wire _5588_;
wire _5589_;
wire _5590_;
wire _5591_;
wire _5592_;
wire _5593_;
wire _5594_;
wire _5595_;
wire _5596_;
wire _5597_;
wire _5598_;
wire _5599_;
wire _5600_;
wire _5601_;
wire _5602_;
wire _5603_;
wire _5604_;
wire _5605_;
wire _5606_;
wire _5607_;
wire _5608_;
wire _5609_;
wire _5610_;
wire _5611_;
wire _5612_;
wire _5613_;
wire _5614_;
wire _5615_;
wire _5616_;
wire _5617_;
wire _5618_;
wire _5619_;
wire _5620_;
wire _5621_;
wire _5622_;
wire _5623_;
wire _5624_;
wire _5625_;
wire _5626_;
wire _5627_;
wire _5628_;
wire _5629_;
wire _5630_;
wire _5631_;
wire _5632_;
wire _5633_;
wire _5634_;
wire _5635_;
wire _5636_;
wire _5637_;
wire _5638_;
wire _5639_;
wire _5640_;
wire _5641_;
wire _5642_;
wire _5643_;
wire _5644_;
wire _5645_;
wire _5646_;
wire _5647_;
wire _5648_;
wire _5649_;
wire _5650_;
wire _5651_;
wire _5652_;
wire _5653_;
wire _5654_;
wire _5655_;
wire _5656_;
wire _5657_;
wire _5658_;
wire _5659_;
wire _5660_;
wire _5661_;
wire _5662_;
wire _5663_;
wire _5664_;
wire _5665_;
wire _5666_;
wire _5667_;
wire _5668_;
wire _5669_;
wire _5670_;
wire _5671_;
wire _5672_;
wire _5673_;
wire _5674_;
wire _5675_;
wire _5676_;
wire _5677_;
wire _5678_;
wire _5679_;
wire _5680_;
wire _5681_;
wire _5682_;
wire _5683_;
wire _5684_;
wire _5685_;
wire _5686_;
wire _5687_;
wire _5688_;
wire _5689_;
wire _5690_;
wire _5691_;
wire _5692_;
wire _5693_;
wire _5694_;
wire _5695_;
wire _5696_;
wire _5697_;
wire _5698_;
wire _5699_;
wire _5700_;
wire _5701_;
wire _5702_;
wire _5703_;
wire _5704_;
wire _5705_;
wire _5706_;
wire _5707_;
wire _5708_;
wire _5709_;
wire _5710_;
wire _5711_;
wire _5712_;
wire _5713_;
wire _5714_;
wire _5715_;
wire _5716_;
wire _5717_;
wire _5718_;
wire _5719_;
wire _5720_;
wire _5721_;
wire _5722_;
wire _5723_;
wire _5724_;
wire _5725_;
wire _5726_;
wire _5727_;
wire _5728_;
wire _5729_;
wire _5730_;
wire _5731_;
wire _5732_;
wire _5733_;
wire _5734_;
wire _5735_;
wire _5736_;
wire _5737_;
wire _5738_;
wire _5739_;
wire _5740_;
wire _5741_;
wire _5742_;
wire _5743_;
wire _5744_;
wire _5745_;
wire _5746_;
wire _5747_;
wire _5748_;
wire _5749_;
wire _5750_;
wire _5751_;
wire _5752_;
wire _5753_;
wire _5754_;
wire _5755_;
wire _5756_;
wire _5757_;
wire _5758_;
wire _5759_;
wire _5760_;
wire _5761_;
wire _5762_;
wire _5763_;
wire _5764_;
wire _5765_;
wire _5766_;
wire _5767_;
wire _5768_;
wire _5769_;
wire _5770_;
wire _5771_;
wire _5772_;
wire _5773_;
wire _5774_;
wire _5775_;
wire _5776_;
wire _5777_;
wire _5778_;
wire _5779_;
wire _5780_;
wire _5781_;
wire _5782_;
wire _5783_;
wire _5784_;
wire _5785_;
wire _5786_;
wire _5787_;
wire _5788_;
wire _5789_;
wire _5790_;
wire _5791_;
wire _5792_;
wire _5793_;
wire _5794_;
wire _5795_;
wire _5796_;
wire _5797_;
wire _5798_;
wire _5799_;
wire _5800_;
wire _5801_;
wire _5802_;
wire _5803_;
wire _5804_;
wire _5805_;
wire _5806_;
wire _5807_;
wire _5808_;
wire _5809_;
wire _5810_;
wire _5811_;
wire _5812_;
wire _5813_;
wire _5814_;
wire _5815_;
wire _5816_;
wire _5817_;
wire _5818_;
wire _5819_;
wire _5820_;
wire _5821_;
wire _5822_;
wire _5823_;
wire _5824_;
wire _5825_;
wire _5826_;
wire _5827_;
wire _5828_;
wire _5829_;
wire _5830_;
wire _5831_;
wire _5832_;
wire _5833_;
wire _5834_;
wire _5835_;
wire _5836_;
wire _5837_;
wire _5838_;
wire _5839_;
wire _5840_;
wire _5841_;
wire _5842_;
wire _5843_;
wire _5844_;
wire _5845_;
wire _5846_;
wire _5847_;
wire _5848_;
wire _5849_;
wire _5850_;
wire _5851_;
wire _5852_;
wire _5853_;
wire _5854_;
wire _5855_;
wire _5856_;
wire _5857_;
wire _5858_;
wire _5859_;
wire _5860_;
wire _5861_;
wire _5862_;
wire _5863_;
wire _5864_;
wire _5865_;
wire _5866_;
wire _5867_;
wire _5868_;
wire _5869_;
wire _5870_;
wire _5871_;
wire _5872_;
wire _5873_;
wire _5874_;
wire _5875_;
wire _5876_;
wire _5877_;
wire _5878_;
wire _5879_;
wire _5880_;
wire _5881_;
wire _5882_;
wire _5883_;
wire _5884_;
wire _5885_;
wire _5886_;
wire _5887_;
wire _5888_;
wire _5889_;
wire _5890_;
wire _5891_;
wire _5892_;
wire _5893_;
wire _5894_;
wire _5895_;
wire _5896_;
wire _5897_;
wire _5898_;
wire _5899_;
wire _5900_;
wire _5901_;
wire _5902_;
wire _5903_;
wire _5904_;
wire _5905_;
wire _5906_;
wire _5907_;
wire _5908_;
wire _5909_;
wire _5910_;
wire _5911_;
wire _5912_;
wire _5913_;
wire _5914_;
wire _5915_;
wire _5916_;
wire _5917_;
wire _5918_;
wire _5919_;
wire _5920_;
wire _5921_;
wire _5922_;
wire _5923_;
wire _5924_;
wire _5925_;
wire _5926_;
wire _5927_;
wire _5928_;
wire _5929_;
wire _5930_;
wire _5931_;
wire _5932_;
wire _5933_;
wire _5934_;
wire _5935_;
wire _5936_;
wire _5937_;
wire _5938_;
wire _5939_;
wire _5940_;
wire _5941_;
wire _5942_;
wire _5943_;
wire _5944_;
wire _5945_;
wire _5946_;
wire _5947_;
wire _5948_;
wire _5949_;
wire _5950_;
wire _5951_;
wire _5952_;
wire _5953_;
wire _5954_;
wire _5955_;
wire _5956_;
wire _5957_;
wire _5958_;
wire _5959_;
wire _5960_;
wire _5961_;
wire _5962_;
wire _5963_;
wire _5964_;
wire _5965_;
wire _5966_;
wire _5967_;
wire _5968_;
wire _5969_;
wire _5970_;
wire _5971_;
wire _5972_;
wire _5973_;
wire _5974_;
wire _5975_;
wire _5976_;
wire _5977_;
wire _5978_;
wire _5979_;
wire _5980_;
wire _5981_;
wire _5982_;
wire _5983_;
wire _5984_;
wire _5985_;
wire _5986_;
wire _5987_;
wire _5988_;
wire _5989_;
wire _5990_;
wire _5991_;
wire _5992_;
wire _5993_;
wire _5994_;
wire _5995_;
wire _5996_;
wire _5997_;
wire _5998_;
wire _5999_;
wire _6000_;
wire _6001_;
wire _6002_;
wire _6003_;
wire _6004_;
wire _6005_;
wire _6006_;
wire _6007_;
wire _6008_;
wire _6009_;
wire _6010_;
wire _6011_;
wire _6012_;
wire _6013_;
wire _6014_;
wire _6015_;
wire _6016_;
wire _6017_;
wire _6018_;
wire _6019_;
wire _6020_;
wire _6021_;
wire _6022_;
wire _6023_;
wire _6024_;
wire _6025_;
wire _6026_;
wire _6027_;
wire _6028_;
wire _6029_;
wire _6030_;
wire _6031_;
wire _6032_;
wire _6033_;
wire _6034_;
wire _6035_;
wire _6036_;
wire _6037_;
wire _6038_;
wire _6039_;
wire _6040_;
wire _6041_;
wire _6042_;
wire _6043_;
wire _6044_;
wire _6045_;
wire _6046_;
wire _6047_;
wire _6048_;
wire _6049_;
wire _6050_;
wire _6051_;
wire _6052_;
wire _6053_;
wire _6054_;
wire _6055_;
wire _6056_;
wire _6057_;
wire _6058_;
wire _6059_;
wire _6060_;
wire _6061_;
wire _6062_;
wire _6063_;
wire _6064_;
wire _6065_;
wire _6066_;
wire _6067_;
wire _6068_;
wire _6069_;
wire _6070_;
wire _6071_;
wire _6072_;
wire _6073_;
wire _6074_;
wire _6075_;
wire _6076_;
wire _6077_;
wire _6078_;
wire _6079_;
wire _6080_;
wire _6081_;
wire _6082_;
wire _6083_;
wire _6084_;
wire _6085_;
wire _6086_;
wire _6087_;
wire _6088_;
wire _6089_;
wire _6090_;
wire _6091_;
wire _6092_;
wire _6093_;
wire _6094_;
wire _6095_;
wire _6096_;
wire _6097_;
wire _6098_;
wire _6099_;
wire _6100_;
wire _6101_;
wire _6102_;
wire _6103_;
wire _6104_;
wire _6105_;
wire _6106_;
wire _6107_;
wire _6108_;
wire _6109_;
wire _6110_;
wire _6111_;
wire _6112_;
wire _6113_;
wire _6114_;
wire _6115_;
wire _6116_;
wire _6117_;
wire _6118_;
wire _6119_;
wire _6120_;
wire _6121_;
wire _6122_;
wire _6123_;
wire _6124_;
wire _6125_;
wire _6126_;
wire _6127_;
wire _6128_;
wire _6129_;
wire _6130_;
wire _6131_;
wire _6132_;
wire _6133_;
wire _6134_;
wire _6135_;
wire _6136_;
wire _6137_;
wire _6138_;
wire _6139_;
wire _6140_;
wire _6141_;
wire _6142_;
wire _6143_;
wire _6144_;
wire _6145_;
wire _6146_;
wire _6147_;
wire _6148_;
wire _6149_;
wire _6150_;
wire _6151_;
wire _6152_;
wire _6153_;
wire _6154_;
wire _6155_;
wire _6156_;
wire _6157_;
wire _6158_;
wire _6159_;
wire _6160_;
wire _6161_;
wire _6162_;
wire _6163_;
wire _6164_;
wire _6165_;
wire _6166_;
wire _6167_;
wire _6168_;
wire _6169_;
wire _6170_;
wire _6171_;
wire _6172_;
wire _6173_;
wire _6174_;
wire _6175_;
wire _6176_;
wire _6177_;
wire _6178_;
wire _6179_;
wire _6180_;
wire _6181_;
wire _6182_;
wire _6183_;
wire _6184_;
wire _6185_;
wire _6186_;
wire _6187_;
wire _6188_;
wire _6189_;
wire _6190_;
wire _6191_;
wire _6192_;
wire _6193_;
wire _6194_;
wire _6195_;
wire _6196_;
wire _6197_;
wire _6198_;
wire _6199_;
wire _6200_;
wire _6201_;
wire _6202_;
wire _6203_;
wire _6204_;
wire _6205_;
wire _6206_;
wire _6207_;
wire _6208_;
wire _6209_;
wire _6210_;
wire _6211_;
wire _6212_;
wire _6213_;
wire _6214_;
wire _6215_;
wire _6216_;
wire _6217_;
wire _6218_;
wire _6219_;
wire _6220_;
wire _6221_;
wire _6222_;
wire _6223_;
wire _6224_;
wire _6225_;
wire _6226_;
wire _6227_;
wire _6228_;
wire _6229_;
wire _6230_;
wire _6231_;
wire _6232_;
wire _6233_;
wire _6234_;
wire _6235_;
wire _6236_;
wire _6237_;
wire _6238_;
wire _6239_;
wire _6240_;
wire _6241_;
wire _6242_;
wire _6243_;
wire _6244_;
wire _6245_;
wire _6246_;
wire _6247_;
wire _6248_;
wire _6249_;
wire _6250_;
wire _6251_;
wire _6252_;
wire _6253_;
wire _6254_;
wire _6255_;
wire _6256_;
wire _6257_;
wire _6258_;
wire _6259_;
wire _6260_;
wire _6261_;
wire _6262_;
wire _6263_;
wire _6264_;
wire _6265_;
wire _6266_;
wire _6267_;
wire _6268_;
wire _6269_;
wire _6270_;
wire _6271_;
wire _6272_;
wire _6273_;
wire _6274_;
wire _6275_;
wire _6276_;
wire _6277_;
wire _6278_;
wire _6279_;
wire _6280_;
wire _6281_;
wire _6282_;
wire _6283_;
wire _6284_;
wire _6285_;
wire _6286_;
wire _6287_;
wire _6288_;
wire _6289_;
wire _6290_;
wire _6291_;
wire _6292_;
wire _6293_;
wire _6294_;
wire _6295_;
wire _6296_;
wire _6297_;
wire _6298_;
wire _6299_;
wire _6300_;
wire _6301_;
wire _6302_;
wire _6303_;
wire _6304_;
wire _6305_;
wire _6306_;
wire _6307_;
wire _6308_;
wire _6309_;
wire _6310_;
wire _6311_;
wire _6312_;
wire _6313_;
wire _6314_;
wire _6315_;
wire _6316_;
wire _6317_;
wire _6318_;
wire _6319_;
wire _6320_;
wire _6321_;
wire _6322_;
wire _6323_;
wire _6324_;
wire _6325_;
wire _6326_;
wire _6327_;
wire _6328_;
wire _6329_;
wire _6330_;
wire _6331_;
wire _6332_;
wire _6333_;
wire _6334_;
wire _6335_;
wire _6336_;
wire _6337_;
wire _6338_;
wire _6339_;
wire _6340_;
wire _6341_;
wire _6342_;
wire _6343_;
wire _6344_;
wire _6345_;
wire _6346_;
wire _6347_;
wire _6348_;
wire _6349_;
wire _6350_;
wire _6351_;
wire _6352_;
wire _6353_;
wire _6354_;
wire _6355_;
wire _6356_;
wire _6357_;
wire _6358_;
wire _6359_;
wire _6360_;
wire _6361_;
wire _6362_;
wire _6363_;
wire _6364_;
wire _6365_;
wire _6366_;
wire _6367_;
wire _6368_;
wire _6369_;
wire _6370_;
wire _6371_;
wire _6372_;
wire _6373_;
wire _6374_;
wire _6375_;
wire _6376_;
wire _6377_;
wire _6378_;
wire _6379_;
wire _6380_;
wire _6381_;
wire _6382_;
wire _6383_;
wire _6384_;
wire _6385_;
wire _6386_;
wire _6387_;
wire _6388_;
wire _6389_;
wire _6390_;
wire _6391_;
wire _6392_;
wire _6393_;
wire _6394_;
wire _6395_;
wire _6396_;
wire _6397_;
wire _6398_;
wire _6399_;
wire _6400_;
wire _6401_;
wire _6402_;
wire _6403_;
wire _6404_;
wire _6405_;
wire _6406_;
wire _6407_;
wire _6408_;
wire _6409_;
wire _6410_;
wire _6411_;
wire _6412_;
wire _6413_;
wire _6414_;
wire _6415_;
wire _6416_;
wire _6417_;
wire _6418_;
wire _6419_;
wire _6420_;
wire _6421_;
wire _6422_;
wire _6423_;
wire _6424_;
wire _6425_;
wire _6426_;
wire _6427_;
wire _6428_;
wire _6429_;
wire _6430_;
wire _6431_;
wire _6432_;
wire _6433_;
wire _6434_;
wire _6435_;
wire _6436_;
wire _6437_;
wire _6438_;
wire _6439_;
wire _6440_;
wire _6441_;
wire _6442_;
wire _6443_;
wire _6444_;
wire _6445_;
wire _6446_;
wire _6447_;
wire _6448_;
wire _6449_;
wire _6450_;
wire _6451_;
wire _6452_;
wire _6453_;
wire _6454_;
wire _6455_;
wire _6456_;
wire _6457_;
wire _6458_;
wire _6459_;
wire _6460_;
wire _6461_;
wire _6462_;
wire _6463_;
wire _6464_;
wire _6465_;
wire _6466_;
wire _6467_;
wire _6468_;
wire _6469_;
wire _6470_;
wire _6471_;
wire _6472_;
wire _6473_;
wire _6474_;
wire _6475_;
wire _6476_;
wire _6477_;
wire _6478_;
wire _6479_;
wire _6480_;
wire _6481_;
wire _6482_;
wire _6483_;
wire _6484_;
wire _6485_;
wire _6486_;
wire _6487_;
wire _6488_;
wire _6489_;
wire _6490_;
wire _6491_;
wire _6492_;
wire _6493_;
wire _6494_;
wire _6495_;
wire _6496_;
wire _6497_;
wire _6498_;
wire _6499_;
wire _6500_;
wire _6501_;
wire _6502_;
wire _6503_;
wire _6504_;
wire _6505_;
wire _6506_;
wire _6507_;
wire _6508_;
wire _6509_;
wire _6510_;
wire _6511_;
wire _6512_;
wire _6513_;
wire _6514_;
wire _6515_;
wire _6516_;
wire _6517_;
wire _6518_;
wire _6519_;
wire _6520_;
wire _6521_;
wire _6522_;
wire _6523_;
wire _6524_;
wire _6525_;
wire _6526_;
wire _6527_;
wire _6528_;
wire _6529_;
wire _6530_;
wire _6531_;
wire _6532_;
wire _6533_;
wire _6534_;
wire _6535_;
wire _6536_;
wire _6537_;
wire _6538_;
wire _6539_;
wire _6540_;
wire _6541_;
wire _6542_;
wire _6543_;
wire _6544_;
wire _6545_;
wire _6546_;
wire _6547_;
wire _6548_;
wire _6549_;
wire _6550_;
wire _6551_;
wire _6552_;
wire _6553_;
wire _6554_;
wire _6555_;
wire _6556_;
wire _6557_;
wire _6558_;
wire _6559_;
wire _6560_;
wire _6561_;
wire _6562_;
wire _6563_;
wire _6564_;
wire _6565_;
wire _6566_;
wire _6567_;
wire _6568_;
wire _6569_;
wire _6570_;
wire _6571_;
wire _6572_;
wire _6573_;
wire _6574_;
wire _6575_;
wire _6576_;
wire _6577_;
wire _6578_;
wire _6579_;
wire _6580_;
wire _6581_;
wire _6582_;
wire _6583_;
wire _6584_;
wire _6585_;
wire _6586_;
wire _6587_;
wire _6588_;
wire _6589_;
wire _6590_;
wire _6591_;
wire _6592_;
wire _6593_;
wire _6594_;
wire _6595_;
wire _6596_;
wire _6597_;
wire _6598_;
wire _6599_;
wire _6600_;
wire _6601_;
wire _6602_;
wire _6603_;
wire _6604_;
wire _6605_;
wire _6606_;
wire _6607_;
wire _6608_;
wire _6609_;
wire _6610_;
wire _6611_;
wire _6612_;
wire _6613_;
wire _6614_;
wire _6615_;
wire _6616_;
wire _6617_;
wire _6618_;
wire _6619_;
wire _6620_;
wire _6621_;
wire _6622_;
wire _6623_;
wire _6624_;
wire _6625_;
wire _6626_;
wire _6627_;
wire _6628_;
wire _6629_;
wire _6630_;
wire _6631_;
wire _6632_;
wire _6633_;
wire _6634_;
wire _6635_;
wire _6636_;
wire _6637_;
wire _6638_;
wire _6639_;
wire _6640_;
wire _6641_;
wire _6642_;
wire _6643_;
wire _6644_;
wire _6645_;
wire _6646_;
wire _6647_;
wire _6648_;
wire _6649_;
wire _6650_;
wire _6651_;
wire _6652_;
wire _6653_;
wire _6654_;
wire _6655_;
wire _6656_;
wire _6657_;
wire _6658_;
wire _6659_;
wire _6660_;
wire _6661_;
wire _6662_;
wire _6663_;
wire _6664_;
wire _6665_;
wire _6666_;
wire _6667_;
wire _6668_;
wire _6669_;
wire _6670_;
wire _6671_;
wire _6672_;
wire _6673_;
wire _6674_;
wire _6675_;
wire _6676_;
wire _6677_;
wire _6678_;
wire _6679_;
wire _6680_;
wire _6681_;
wire _6682_;
wire _6683_;
wire _6684_;
wire _6685_;
wire _6686_;
wire _6687_;
wire _6688_;
wire _6689_;
wire _6690_;
wire _6691_;
wire _6692_;
wire _6693_;
wire _6694_;
wire _6695_;
wire _6696_;
wire _6697_;
wire _6698_;
wire _6699_;
wire _6700_;
wire _6701_;
wire _6702_;
wire _6703_;
wire _6704_;
wire _6705_;
wire _6706_;
wire _6707_;
wire _6708_;
wire _6709_;
wire _6710_;
wire _6711_;
wire _6712_;
wire _6713_;
wire _6714_;
wire _6715_;
wire _6716_;
wire _6717_;
wire _6718_;
wire _6719_;
wire _6720_;
wire _6721_;
wire _6722_;
wire _6723_;
wire _6724_;
wire _6725_;
wire _6726_;
wire _6727_;
wire _6728_;
wire _6729_;
wire _6730_;
wire _6731_;
wire _6732_;
wire _6733_;
wire _6734_;
wire _6735_;
wire _6736_;
wire _6737_;
wire _6738_;
wire _6739_;
wire _6740_;
wire _6741_;
wire _6742_;
wire _6743_;
wire _6744_;
wire _6745_;
wire _6746_;
wire _6747_;
wire _6748_;
wire _6749_;
wire _6750_;
wire _6751_;
wire _6752_;
wire _6753_;
wire _6754_;
wire _6755_;
wire _6756_;
wire _6757_;
wire _6758_;
wire _6759_;
wire _6760_;
wire _6761_;
wire _6762_;
wire _6763_;
wire _6764_;
wire _6765_;
wire _6766_;
wire _6767_;
wire _6768_;
wire _6769_;
wire _6770_;
wire _6771_;
wire _6772_;
wire _6773_;
wire _6774_;
wire _6775_;
wire _6776_;
wire _6777_;
wire _6778_;
wire _6779_;
wire _6780_;
wire _6781_;
wire _6782_;
wire _6783_;
wire _6784_;
wire _6785_;
wire _6786_;
wire _6787_;
wire _6788_;
wire _6789_;
wire _6790_;
wire _6791_;
wire _6792_;
wire _6793_;
wire _6794_;
wire _6795_;
wire _6796_;
wire _6797_;
wire _6798_;
wire _6799_;
wire _6800_;
wire _6801_;
wire _6802_;
wire _6803_;
wire _6804_;
wire _6805_;
wire _6806_;
wire _6807_;
wire _6808_;
wire _6809_;
wire _6810_;
wire _6811_;
wire _6812_;
wire _6813_;
wire _6814_;
wire _6815_;
wire _6816_;
wire _6817_;
wire _6818_;
wire _6819_;
wire _6820_;
wire _6821_;
wire _6822_;
wire _6823_;
wire _6824_;
wire _6825_;
wire _6826_;
wire _6827_;
wire _6828_;
wire _6829_;
wire _6830_;
wire _6831_;
wire _6832_;
wire _6833_;
wire _6834_;
wire _6835_;
wire _6836_;
wire _6837_;
wire _6838_;
wire _6839_;
wire _6840_;
wire _6841_;
wire _6842_;
wire _6843_;
wire _6844_;
wire _6845_;
wire _6846_;
wire _6847_;
wire _6848_;
wire _6849_;
wire _6850_;
wire _6851_;
wire _6852_;
wire _6853_;
wire _6854_;
wire _6855_;
wire _6856_;
wire _6857_;
wire _6858_;
wire _6859_;
wire _6860_;
wire _6861_;
wire _6862_;
wire _6863_;
wire _6864_;
wire _6865_;
wire _6866_;
wire _6867_;
wire _6868_;
wire _6869_;
wire _6870_;
wire _6871_;
wire _6872_;
wire _6873_;
wire _6874_;
wire _6875_;
wire _6876_;
wire _6877_;
wire _6878_;
wire _6879_;
wire _6880_;
wire _6881_;
wire _6882_;
wire _6883_;
wire _6884_;
wire _6885_;
wire _6886_;
wire _6887_;
wire _6888_;
wire _6889_;
wire _6890_;
wire _6891_;
wire _6892_;
wire _6893_;
wire _6894_;
wire _6895_;
wire _6896_;
wire _6897_;
wire _6898_;
wire _6899_;
wire _6900_;
wire _6901_;
wire _6902_;
wire _6903_;
wire _6904_;
wire _6905_;
wire _6906_;
wire _6907_;
wire _6908_;
wire _6909_;
wire _6910_;
wire _6911_;
wire _6912_;
wire _6913_;
wire _6914_;
wire _6915_;
wire _6916_;
wire _6917_;
wire _6918_;
wire _6919_;
wire _6920_;
wire _6921_;
wire _6922_;
wire _6923_;
wire _6924_;
wire _6925_;
wire _6926_;
wire _6927_;
wire _6928_;
wire _6929_;
wire _6930_;
wire _6931_;
wire _6932_;
wire _6933_;
wire _6934_;
wire _6935_;
wire _6936_;
wire _6937_;
wire _6938_;
wire _6939_;
wire _6940_;
wire _6941_;
wire _6942_;
wire _6943_;
wire _6944_;
wire _6945_;
wire _6946_;
wire _6947_;
wire _6948_;
wire _6949_;
wire _6950_;
wire _6951_;
wire _6952_;
wire _6953_;
wire _6954_;
wire _6955_;
wire _6956_;
wire _6957_;
wire _6958_;
wire _6959_;
wire _6960_;
wire _6961_;
wire _6962_;
wire _6963_;
wire _6964_;
wire _6965_;
wire _6966_;
wire _6967_;
wire _6968_;
wire _6969_;
wire _6970_;
wire _6971_;
wire _6972_;
wire _6973_;
wire _6974_;
wire _6975_;
wire _6976_;
wire _6977_;
wire _6978_;
wire _6979_;
wire _6980_;
wire _6981_;
wire _6982_;
wire _6983_;
wire _6984_;
wire _6985_;
wire _6986_;
wire _6987_;
wire _6988_;
wire _6989_;
wire _6990_;
wire _6991_;
wire _6992_;
wire _6993_;
wire _6994_;
wire _6995_;
wire _6996_;
wire _6997_;
wire _6998_;
wire _6999_;
wire _7000_;
wire _7001_;
wire _7002_;
wire _7003_;
wire _7004_;
wire _7005_;
wire _7006_;
wire _7007_;
wire _7008_;
wire _7009_;
wire _7010_;
wire _7011_;
wire _7012_;
wire _7013_;
wire _7014_;
wire _7015_;
wire _7016_;
wire _7017_;
wire _7018_;
wire _7019_;
wire _7020_;
wire _7021_;
wire _7022_;
wire _7023_;
wire _7024_;
wire _7025_;
wire _7026_;
wire _7027_;
wire _7028_;
wire _7029_;
wire _7030_;
wire _7031_;
wire _7032_;
wire _7033_;
wire _7034_;
wire _7035_;
wire _7036_;
wire _7037_;
wire _7038_;
wire _7039_;
wire _7040_;
wire _7041_;
wire _7042_;
wire _7043_;
wire _7044_;
wire _7045_;
wire _7046_;
wire _7047_;
wire _7048_;
wire _7049_;
wire _7050_;
wire _7051_;
wire _7052_;
wire _7053_;
wire _7054_;
wire _7055_;
wire _7056_;
wire _7057_;
wire _7058_;
wire _7059_;
wire _7060_;
wire _7061_;
wire _7062_;
wire _7063_;
wire _7064_;
wire _7065_;
wire _7066_;
wire _7067_;
wire _7068_;
wire _7069_;
wire _7070_;
wire _7071_;
wire _7072_;
wire _7073_;
wire _7074_;
wire _7075_;
wire _7076_;
wire _7077_;
wire _7078_;
wire _7079_;
wire _7080_;
wire _7081_;
wire _7082_;
wire _7083_;
wire _7084_;
wire _7085_;
wire _7086_;
wire _7087_;
wire _7088_;
wire _7089_;
wire _7090_;
wire _7091_;
wire _7092_;
wire _7093_;
wire _7094_;
wire _7095_;
wire _7096_;
wire _7097_;
wire _7098_;
wire _7099_;
wire _7100_;
wire _7101_;
wire _7102_;
wire _7103_;
wire _7104_;
wire _7105_;
wire _7106_;
wire _7107_;
wire _7108_;
wire _7109_;
wire _7110_;
wire _7111_;
wire _7112_;
wire _7113_;
wire _7114_;
wire _7115_;
wire _7116_;
wire _7117_;
wire _7118_;
wire _7119_;
wire _7120_;
wire _7121_;
wire _7122_;
wire _7123_;
wire _7124_;
wire _7125_;
wire _7126_;
wire _7127_;
wire _7128_;
wire _7129_;
wire _7130_;
wire _7131_;
wire _7132_;
wire _7133_;
wire _7134_;
wire _7135_;
wire _7136_;
wire _7137_;
wire _7138_;
wire _7139_;
wire _7140_;
wire _7141_;
wire _7142_;
wire _7143_;
wire _7144_;
wire _7145_;
wire _7146_;
wire _7147_;
wire _7148_;
wire _7149_;
wire _7150_;
wire _7151_;
wire _7152_;
wire _7153_;
wire _7154_;
wire _7155_;
wire _7156_;
wire _7157_;
wire _7158_;
wire _7159_;
wire _7160_;
wire _7161_;
wire _7162_;
wire _7163_;
wire _7164_;
wire _7165_;
wire _7166_;
wire _7167_;
wire _7168_;
wire _7169_;
wire _7170_;
wire _7171_;
wire _7172_;
wire _7173_;
wire _7174_;
wire _7175_;
wire _7176_;
wire _7177_;
wire _7178_;
wire _7179_;
wire _7180_;
wire _7181_;
wire _7182_;
wire _7183_;
wire _7184_;
wire _7185_;
wire _7186_;
wire _7187_;
wire _7188_;
wire _7189_;
wire _7190_;
wire _7191_;
wire _7192_;
wire _7193_;
wire _7194_;
wire _7195_;
wire _7196_;
wire _7197_;
wire _7198_;
wire _7199_;
wire _7200_;
wire _7201_;
wire _7202_;
wire _7203_;
wire _7204_;
wire _7205_;
wire _7206_;
wire _7207_;
wire _7208_;
wire _7209_;
wire _7210_;
wire _7211_;
wire _7212_;
wire _7213_;
wire _7214_;
wire _7215_;
wire _7216_;
wire _7217_;
wire _7218_;
wire _7219_;
wire _7220_;
wire _7221_;
wire _7222_;
wire _7223_;
wire _7224_;
wire _7225_;
wire _7226_;
wire _7227_;
wire _7228_;
wire _7229_;
wire _7230_;
wire _7231_;
wire _7232_;
wire _7233_;
wire _7234_;
wire _7235_;
wire _7236_;
wire _7237_;
wire _7238_;
wire _7239_;
wire _7240_;
wire _7241_;
wire _7242_;
wire _7243_;
wire _7244_;
wire _7245_;
wire _7246_;
wire _7247_;
wire _7248_;
wire _7249_;
wire _7250_;
wire _7251_;
wire _7252_;
wire _7253_;
wire _7254_;
wire _7255_;
wire _7256_;
wire _7257_;
wire _7258_;
wire _7259_;
wire _7260_;
wire _7261_;
wire _7262_;
wire _7263_;
wire _7264_;
wire _7265_;
wire _7266_;
wire _7267_;
wire _7268_;
wire _7269_;
wire _7270_;
wire _7271_;
wire _7272_;
wire _7273_;
wire _7274_;
wire _7275_;
wire _7276_;
wire _7277_;
wire _7278_;
wire _7279_;
wire _7280_;
wire _7281_;
wire _7282_;
wire _7283_;
wire _7284_;
wire _7285_;
wire _7286_;
wire _7287_;
wire _7288_;
wire _7289_;
wire _7290_;
wire _7291_;
wire _7292_;
wire _7293_;
wire _7294_;
wire _7295_;
wire _7296_;
wire _7297_;
wire _7298_;
wire _7299_;
wire _7300_;
wire _7301_;
wire _7302_;
wire _7303_;
wire _7304_;
wire _7305_;
wire _7306_;
wire _7307_;
wire _7308_;
wire _7309_;
wire _7310_;
wire _7311_;
wire _7312_;
wire _7313_;
wire _7314_;
wire _7315_;
wire _7316_;
wire _7317_;
wire _7318_;
wire _7319_;
wire _7320_;
wire _7321_;
wire _7322_;
wire _7323_;
wire _7324_;
wire _7325_;
wire _7326_;
wire _7327_;
wire _7328_;
wire _7329_;
wire _7330_;
wire _7331_;
wire _7332_;
wire _7333_;
wire _7334_;
wire _7335_;
wire _7336_;
wire _7337_;
wire _7338_;
wire _7339_;
wire _7340_;
wire _7341_;
wire _7342_;
wire _7343_;
wire _7344_;
wire _7345_;
wire _7346_;
wire _7347_;
wire _7348_;
wire _7349_;
wire _7350_;
wire _7351_;
wire _7352_;
wire _7353_;
wire _7354_;
wire _7355_;
wire _7356_;
wire _7357_;
wire _7358_;
wire _7359_;
wire _7360_;
wire _7361_;
wire _7362_;
wire _7363_;
wire _7364_;
wire _7365_;
wire _7366_;
wire _7367_;
wire _7368_;
wire _7369_;
wire _7370_;
wire _7371_;
wire _7372_;
wire _7373_;
wire _7374_;
wire _7375_;
wire _7376_;
wire _7377_;
wire _7378_;
wire _7379_;
wire _7380_;
wire _7381_;
wire _7382_;
wire _7383_;
wire _7384_;
wire _7385_;
wire _7386_;
wire _7387_;
wire _7388_;
wire _7389_;
wire _7390_;
wire _7391_;
wire _7392_;
wire _7393_;
wire _7394_;
wire _7395_;
wire _7396_;
wire _7397_;
wire _7398_;
wire _7399_;
wire _7400_;
wire _7401_;
wire _7402_;
wire _7403_;
wire _7404_;
wire _7405_;
wire _7406_;
wire _7407_;
wire _7408_;
wire _7409_;
wire _7410_;
wire _7411_;
wire _7412_;
wire _7413_;
wire _7414_;
wire _7415_;
wire _7416_;
wire _7417_;
wire _7418_;
wire _7419_;
wire _7420_;
wire _7421_;
wire _7422_;
wire _7423_;
wire _7424_;
wire _7425_;
wire _7426_;
wire _7427_;
wire _7428_;
wire _7429_;
wire _7430_;
wire _7431_;
wire _7432_;
wire _7433_;
wire _7434_;
wire _7435_;
wire _7436_;
wire _7437_;
wire _7438_;
wire _7439_;
wire _7440_;
wire _7441_;
wire _7442_;
wire _7443_;
wire _7444_;
wire _7445_;
wire _7446_;
wire _7447_;
wire _7448_;
wire _7449_;
wire _7450_;
wire _7451_;
wire _7452_;
wire _7453_;
wire _7454_;
wire _7455_;
wire _7456_;
wire _7457_;
wire _7458_;
wire _7459_;
wire _7460_;
wire _7461_;
wire _7462_;
wire _7463_;
wire _7464_;
wire _7465_;
wire _7466_;
wire _7467_;
wire _7468_;
wire _7469_;
wire _7470_;
wire _7471_;
wire _7472_;
wire _7473_;
wire _7474_;
wire _7475_;
wire _7476_;
wire _7477_;
wire _7478_;
wire _7479_;
wire _7480_;
wire _7481_;
wire _7482_;
wire _7483_;
wire _7484_;
wire _7485_;
wire _7486_;
wire _7487_;
wire _7488_;
wire _7489_;
wire _7490_;
wire _7491_;
wire _7492_;
wire _7493_;
wire _7494_;
wire _7495_;
wire _7496_;
wire _7497_;
wire _7498_;
wire _7499_;
wire _7500_;
wire _7501_;
wire _7502_;
wire _7503_;
wire _7504_;
wire _7505_;
wire _7506_;
wire _7507_;
wire _7508_;
wire _7509_;
wire _7510_;
wire _7511_;
wire _7512_;
wire _7513_;
wire _7514_;
wire _7515_;
wire _7516_;
wire _7517_;
wire _7518_;
wire _7519_;
wire _7520_;
wire _7521_;
wire _7522_;
wire _7523_;
wire _7524_;
wire _7525_;
wire _7526_;
wire _7527_;
wire _7528_;
wire _7529_;
wire _7530_;
wire _7531_;
wire _7532_;
wire _7533_;
wire _7534_;
wire _7535_;
wire _7536_;
wire _7537_;
wire _7538_;
wire _7539_;
wire _7540_;
wire _7541_;
wire _7542_;
wire _7543_;
wire _7544_;
wire _7545_;
wire _7546_;
wire _7547_;
wire _7548_;
wire _7549_;
wire _7550_;
wire _7551_;
wire _7552_;
wire _7553_;
wire _7554_;
wire _7555_;
wire _7556_;
wire _7557_;
wire _7558_;
wire _7559_;
wire _7560_;
wire _7561_;
wire _7562_;
wire _7563_;
wire _7564_;
wire _7565_;
wire _7566_;
wire _7567_;
wire _7568_;
wire _7569_;
wire _7570_;
wire _7571_;
wire _7572_;
wire _7573_;
wire _7574_;
wire _7575_;
wire _7576_;
wire _7577_;
wire _7578_;
wire _7579_;
wire _7580_;
wire _7581_;
wire _7582_;
wire _7583_;
wire _7584_;
wire _7585_;
wire _7586_;
wire _7587_;
wire _7588_;
wire _7589_;
wire _7590_;
wire _7591_;
wire _7592_;
wire _7593_;
wire _7594_;
wire _7595_;
wire _7596_;
wire _7597_;
wire _7598_;
wire _7599_;
wire _7600_;
wire _7601_;
wire _7602_;
wire _7603_;
wire _7604_;
wire _7605_;
wire _7606_;
wire _7607_;
wire _7608_;
wire _7609_;
wire _7610_;
wire _7611_;
wire _7612_;
wire _7613_;
wire _7614_;
wire _7615_;
wire _7616_;
wire _7617_;
wire _7618_;
wire _7619_;
wire _7620_;
wire _7621_;
wire _7622_;
wire _7623_;
wire _7624_;
wire _7625_;
wire _7626_;
wire _7627_;
wire _7628_;
wire _7629_;
wire _7630_;
wire _7631_;
wire _7632_;
wire _7633_;
wire _7634_;
wire _7635_;
wire _7636_;
wire _7637_;
wire _7638_;
wire _7639_;
wire _7640_;
wire _7641_;
wire _7642_;
wire _7643_;
wire _7644_;
wire _7645_;
wire _7646_;
wire _7647_;
wire _7648_;
wire _7649_;
wire _7650_;
wire _7651_;
wire _7652_;
wire _7653_;
wire _7654_;
wire _7655_;
wire _7656_;
wire _7657_;
wire _7658_;
wire _7659_;
wire _7660_;
wire _7661_;
wire _7662_;
wire _7663_;
wire _7664_;
wire _7665_;
wire _7666_;
wire _7667_;
wire _7668_;
wire _7669_;
wire _7670_;
wire _7671_;
wire _7672_;
wire _7673_;
wire _7674_;
wire _7675_;
wire _7676_;
wire _7677_;
wire _7678_;
wire _7679_;
wire _7680_;
wire _7681_;
wire _7682_;
wire _7683_;
wire _7684_;
wire _7685_;
wire _7686_;
wire _7687_;
wire _7688_;
wire _7689_;
wire _7690_;
wire _7691_;
wire _7692_;
wire _7693_;
wire _7694_;
wire _7695_;
wire _7696_;
wire _7697_;
wire _7698_;
wire _7699_;
wire _7700_;
wire _7701_;
wire _7702_;
wire _7703_;
wire _7704_;
wire _7705_;
wire _7706_;
wire _7707_;
wire _7708_;
wire _7709_;
wire _7710_;
wire _7711_;
wire _7712_;
wire _7713_;
wire _7714_;
wire _7715_;
wire _7716_;
wire _7717_;
wire _7718_;
wire _7719_;
wire _7720_;
wire _7721_;
wire _7722_;
wire _7723_;
wire _7724_;
wire _7725_;
wire _7726_;
wire _7727_;
wire _7728_;
wire _7729_;
wire _7730_;
wire _7731_;
wire _7732_;
wire _7733_;
wire _7734_;
wire _7735_;
wire _7736_;
wire _7737_;
wire _7738_;
wire _7739_;
wire _7740_;
wire _7741_;
wire _7742_;
wire _7743_;
wire _7744_;
wire _7745_;
wire _7746_;
wire _7747_;
wire _7748_;
wire _7749_;
wire _7750_;
wire _7751_;
wire _7752_;
wire _7753_;
wire _7754_;
wire _7755_;
wire _7756_;
wire _7757_;
wire _7758_;
wire _7759_;
wire _7760_;
wire _7761_;
wire _7762_;
wire _7763_;
wire _7764_;
wire _7765_;
wire _7766_;
wire _7767_;
wire _7768_;
wire _7769_;
wire _7770_;
wire _7771_;
wire _7772_;
wire _7773_;
wire _7774_;
wire _7775_;
wire _7776_;
wire _7777_;
wire _7778_;
wire _7779_;
wire _7780_;
wire _7781_;
wire _7782_;
wire _7783_;
wire _7784_;
wire _7785_;
wire _7786_;
wire _7787_;
wire _7788_;
wire _7789_;
wire _7790_;
wire _7791_;
wire _7792_;
wire _7793_;
wire _7794_;
wire _7795_;
wire _7796_;
wire _7797_;
wire _7798_;
wire _7799_;
wire _7800_;
wire _7801_;
wire _7802_;
wire _7803_;
wire _7804_;
wire _7805_;
wire _7806_;
wire _7807_;
wire _7808_;
wire _7809_;
wire _7810_;
wire _7811_;
wire _7812_;
wire _7813_;
wire _7814_;
wire _7815_;
wire _7816_;
wire _7817_;
wire _7818_;
wire _7819_;
wire _7820_;
wire _7821_;
wire _7822_;
wire _7823_;
wire _7824_;
wire _7825_;
wire _7826_;
wire _7827_;
wire _7828_;
wire _7829_;
wire _7830_;
wire _7831_;
wire _7832_;
wire _7833_;
wire _7834_;
wire _7835_;
wire _7836_;
wire _7837_;
wire _7838_;
wire _7839_;
wire _7840_;
wire _7841_;
wire _7842_;
wire _7843_;
wire _7844_;
wire _7845_;
wire _7846_;
wire _7847_;
wire _7848_;
wire _7849_;
wire _7850_;
wire _7851_;
wire _7852_;
wire _7853_;
wire _7854_;
wire _7855_;
wire _7856_;
wire _7857_;
wire _7858_;
wire _7859_;
wire _7860_;
wire _7861_;
wire _7862_;
wire _7863_;
wire _7864_;
wire _7865_;
wire _7866_;
wire _7867_;
wire _7868_;
wire _7869_;
wire _7870_;
wire _7871_;
wire _7872_;
wire _7873_;
wire _7874_;
wire _7875_;
wire _7876_;
wire _7877_;
wire _7878_;
wire _7879_;
wire _7880_;
wire _7881_;
wire _7882_;
wire _7883_;
wire _7884_;
wire _7885_;
wire _7886_;
wire _7887_;
wire _7888_;
wire _7889_;
wire _7890_;
wire _7891_;
wire _7892_;
wire _7893_;
wire _7894_;
wire _7895_;
wire _7896_;
wire _7897_;
wire _7898_;
wire _7899_;
wire _7900_;
wire _7901_;
wire _7902_;
wire _7903_;
wire _7904_;
wire _7905_;
wire _7906_;
wire _7907_;
wire _7908_;
wire _7909_;
wire _7910_;
wire _7911_;
wire _7912_;
wire _7913_;
wire _7914_;
wire _7915_;
wire _7916_;
wire _7917_;
wire _7918_;
wire _7919_;
wire _7920_;
wire _7921_;
wire _7922_;
wire _7923_;
wire _7924_;
wire _7925_;
wire _7926_;
wire _7927_;
wire _7928_;
wire _7929_;
wire _7930_;
wire _7931_;
wire _7932_;
wire _7933_;
wire _7934_;
wire _7935_;
wire _7936_;
wire _7937_;
wire _7938_;
wire _7939_;
wire _7940_;
wire _7941_;
wire _7942_;
wire _7943_;
wire _7944_;
wire _7945_;
wire _7946_;
wire _7947_;
wire _7948_;
wire _7949_;
wire _7950_;
wire _7951_;
wire _7952_;
wire _7953_;
wire _7954_;
wire _7955_;
wire _7956_;
wire _7957_;
wire _7958_;
wire _7959_;
wire _7960_;
wire _7961_;
wire _7962_;
wire _7963_;
wire _7964_;
wire _7965_;
wire _7966_;
wire _7967_;
wire _7968_;
wire _7969_;
wire _7970_;
wire _7971_;
wire _7972_;
wire _7973_;
wire _7974_;
wire _7975_;
wire _7976_;
wire _7977_;
wire _7978_;
wire _7979_;
wire _7980_;
wire _7981_;
wire _7982_;
wire _7983_;
wire _7984_;
wire _7985_;
wire _7986_;
wire _7987_;
wire _7988_;
wire _7989_;
wire _7990_;
wire _7991_;
wire _7992_;
wire _7993_;
wire _7994_;
wire _7995_;
wire _7996_;
wire _7997_;
wire _7998_;
wire _7999_;
wire _8000_;
wire _8001_;
wire _8002_;
wire _8003_;
wire _8004_;
wire _8005_;
wire _8006_;
wire _8007_;
wire _8008_;
wire _8009_;
wire _8010_;
wire _8011_;
wire _8012_;
wire _8013_;
wire _8014_;
wire _8015_;
wire _8016_;
wire _8017_;
wire _8018_;
wire _8019_;
wire _8020_;
wire _8021_;
wire _8022_;
wire _8023_;
wire _8024_;
wire _8025_;
wire _8026_;
wire _8027_;
wire _8028_;
wire _8029_;
wire _8030_;
wire _8031_;
wire _8032_;
wire _8033_;
wire _8034_;
wire _8035_;
wire _8036_;
wire _8037_;
wire _8038_;
wire _8039_;
wire _8040_;
wire _8041_;
wire _8042_;
wire _8043_;
wire _8044_;
wire _8045_;
wire _8046_;
wire _8047_;
wire _8048_;
wire _8049_;
wire _8050_;
wire _8051_;
wire _8052_;
wire _8053_;
wire _8054_;
wire _8055_;
wire _8056_;
wire _8057_;
wire _8058_;
wire _8059_;
wire _8060_;
wire _8061_;
wire _8062_;
wire _8063_;
wire _8064_;
wire _8065_;
wire _8066_;
wire _8067_;
wire _8068_;
wire _8069_;
wire _8070_;
wire _8071_;
wire _8072_;
wire _8073_;
wire _8074_;
wire _8075_;
wire _8076_;
wire _8077_;
wire _8078_;
wire _8079_;
wire _8080_;
wire _8081_;
wire _8082_;
wire _8083_;
wire _8084_;
wire _8085_;
wire _8086_;
wire _8087_;
wire _8088_;
wire _8089_;
wire _8090_;
wire _8091_;
wire _8092_;
wire _8093_;
wire _8094_;
wire _8095_;
wire _8096_;
wire _8097_;
wire _8098_;
wire _8099_;
wire _8100_;
wire _8101_;
wire _8102_;
wire _8103_;
wire _8104_;
wire _8105_;
wire _8106_;
wire _8107_;
wire _8108_;
wire _8109_;
wire _8110_;
wire _8111_;
wire _8112_;
wire _8113_;
wire _8114_;
wire _8115_;
wire _8116_;
wire _8117_;
wire _8118_;
wire _8119_;
wire _8120_;
wire _8121_;
wire _8122_;
wire _8123_;
wire _8124_;
wire _8125_;
wire _8126_;
wire _8127_;
wire _8128_;
wire _8129_;
wire _8130_;
wire _8131_;
wire _8132_;
wire _8133_;
wire _8134_;
wire _8135_;
wire _8136_;
wire _8137_;
wire _8138_;
wire _8139_;
wire _8140_;
wire _8141_;
wire _8142_;
wire _8143_;
wire _8144_;
wire _8145_;
wire _8146_;
wire _8147_;
wire _8148_;
wire _8149_;
wire _8150_;
wire _8151_;
wire _8152_;
wire _8153_;
wire _8154_;
wire _8155_;
wire _8156_;
wire _8157_;
wire _8158_;
wire _8159_;
wire _8160_;
wire _8161_;
wire _8162_;
wire _8163_;
wire _8164_;
wire _8165_;
wire _8166_;
wire _8167_;
wire _8168_;
wire _8169_;
wire _8170_;
wire _8171_;
wire _8172_;
wire _8173_;
wire _8174_;
wire _8175_;
wire _8176_;
wire _8177_;
wire _8178_;
wire _8179_;
wire _8180_;
wire _8181_;
wire _8182_;
wire _8183_;
wire _8184_;
wire _8185_;
wire _8186_;
wire _8187_;
wire _8188_;
wire _8189_;
wire _8190_;
wire _8191_;
wire _8192_;
wire _8193_;
wire _8194_;
wire _8195_;
wire _8196_;
wire _8197_;
wire _8198_;
wire _8199_;
wire _8200_;
wire _8201_;
wire _8202_;
wire _8203_;
wire _8204_;
wire _8205_;
wire _8206_;
wire _8207_;
wire _8208_;
wire _8209_;
wire _8210_;
wire _8211_;
wire _8212_;
wire _8213_;
wire _8214_;
wire _8215_;
wire _8216_;
wire _8217_;
wire _8218_;
wire _8219_;
wire _8220_;
wire _8221_;
wire _8222_;
wire _8223_;
wire _8224_;
wire _8225_;
wire _8226_;
wire _8227_;
wire _8228_;
wire _8229_;
wire _8230_;
wire _8231_;
wire _8232_;
wire _8233_;
wire _8234_;
wire _8235_;
wire _8236_;
wire _8237_;
wire _8238_;
wire _8239_;
wire _8240_;
wire _8241_;
wire _8242_;
wire _8243_;
wire _8244_;
wire _8245_;
wire _8246_;
wire _8247_;
wire _8248_;
wire _8249_;
wire _8250_;
wire _8251_;
wire _8252_;
wire _8253_;
wire _8254_;
wire _8255_;
wire _8256_;
wire _8257_;
wire _8258_;
wire _8259_;
wire _8260_;
wire _8261_;
wire _8262_;
wire _8263_;
wire _8264_;
wire _8265_;
wire _8266_;
wire _8267_;
wire _8268_;
wire _8269_;
wire _8270_;
wire _8271_;
wire _8272_;
wire _8273_;
wire _8274_;
wire _8275_;
wire _8276_;
wire _8277_;
wire _8278_;
wire _8279_;
wire _8280_;
wire _8281_;
wire _8282_;
wire _8283_;
wire _8284_;
wire _8285_;
wire _8286_;
wire _8287_;
wire _8288_;
wire _8289_;
wire _8290_;
wire _8291_;
wire _8292_;
wire _8293_;
wire _8294_;
wire _8295_;
wire _8296_;
wire _8297_;
wire _8298_;
wire _8299_;
wire _8300_;
wire _8301_;
wire _8302_;
wire _8303_;
wire _8304_;
wire _8305_;
wire _8306_;
wire _8307_;
wire _8308_;
wire _8309_;
wire _8310_;
wire _8311_;
wire _8312_;
wire _8313_;
wire _8314_;
wire _8315_;
wire _8316_;
wire _8317_;
wire _8318_;
wire _8319_;
wire _8320_;
wire _8321_;
wire _8322_;
wire _8323_;
wire _8324_;
wire _8325_;
wire _8326_;
wire _8327_;
wire _8328_;
wire _8329_;
wire _8330_;
wire _8331_;
wire _8332_;
wire _8333_;
wire _8334_;
wire _8335_;
wire _8336_;
wire _8337_;
wire _8338_;
wire _8339_;
wire _8340_;
wire _8341_;
wire _8342_;
wire _8343_;
wire _8344_;
wire _8345_;
wire _8346_;
wire _8347_;
wire _8348_;
wire _8349_;
wire _8350_;
wire _8351_;
wire _8352_;
wire _8353_;
wire _8354_;
wire _8355_;
wire _8356_;
wire _8357_;
wire _8358_;
wire _8359_;
wire _8360_;
wire _8361_;
wire _8362_;
wire _8363_;
wire _8364_;
wire _8365_;
wire _8366_;
wire _8367_;
wire _8368_;
wire _8369_;
wire _8370_;
wire _8371_;
wire _8372_;
wire _8373_;
wire _8374_;
wire _8375_;
wire _8376_;
wire _8377_;
wire _8378_;
wire _8379_;
wire _8380_;
wire _8381_;
wire _8382_;
wire _8383_;
wire _8384_;
wire _8385_;
wire _8386_;
wire _8387_;
wire _8388_;
wire _8389_;
wire _8390_;
wire _8391_;
wire _8392_;
wire _8393_;
wire _8394_;
wire _8395_;
wire _8396_;
wire _8397_;
wire _8398_;
wire _8399_;
wire _8400_;
wire _8401_;
wire _8402_;
wire _8403_;
wire _8404_;
wire _8405_;
wire _8406_;
wire _8407_;
wire _8408_;
wire _8409_;
wire _8410_;
wire _8411_;
wire _8412_;
wire _8413_;
wire _8414_;
wire _8415_;
wire _8416_;
wire _8417_;
wire _8418_;
wire _8419_;
wire _8420_;
wire _8421_;
wire _8422_;
wire _8423_;
wire _8424_;
wire _8425_;
wire _8426_;
wire _8427_;
wire _8428_;
wire _8429_;
wire _8430_;
wire _8431_;
wire _8432_;
wire _8433_;
wire _8434_;
wire _8435_;
wire _8436_;
wire _8437_;
wire _8438_;
wire _8439_;
wire _8440_;
wire _8441_;
wire _8442_;
wire _8443_;
wire _8444_;
wire _8445_;
wire _8446_;
wire _8447_;
wire _8448_;
wire _8449_;
wire _8450_;
wire _8451_;
wire _8452_;
wire _8453_;
wire _8454_;
wire _8455_;
wire _8456_;
wire _8457_;
wire _8458_;
wire _8459_;
wire _8460_;
wire _8461_;
wire _8462_;
wire _8463_;
wire _8464_;
wire _8465_;
wire _8466_;
wire _8467_;
wire _8468_;
wire _8469_;
wire _8470_;
wire _8471_;
wire _8472_;
wire _8473_;
wire _8474_;
wire _8475_;
wire _8476_;
wire _8477_;
wire _8478_;
wire _8479_;
wire _8480_;
wire _8481_;
wire _8482_;
wire _8483_;
wire _8484_;
wire _8485_;
wire _8486_;
wire _8487_;
wire _8488_;
wire _8489_;
wire _8490_;
wire _8491_;
wire _8492_;
wire _8493_;
wire _8494_;
wire _8495_;
wire _8496_;
wire _8497_;
wire _8498_;
wire _8499_;
wire _8500_;
wire _8501_;
wire _8502_;
wire _8503_;
wire _8504_;
wire _8505_;
wire _8506_;
wire _8507_;
wire _8508_;
wire _8509_;
wire _8510_;
wire _8511_;
wire _8512_;
wire _8513_;
wire _8514_;
wire _8515_;
wire _8516_;
wire _8517_;
wire _8518_;
wire _8519_;
wire _8520_;
wire _8521_;
wire _8522_;
wire _8523_;
wire _8524_;
wire _8525_;
wire _8526_;
wire _8527_;
wire _8528_;
wire _8529_;
wire _8530_;
wire _8531_;
wire _8532_;
wire _8533_;
wire _8534_;
wire _8535_;
wire _8536_;
wire _8537_;
wire _8538_;
wire _8539_;
wire _8540_;
wire _8541_;
wire _8542_;
wire _8543_;
wire _8544_;
wire _8545_;
wire _8546_;
wire _8547_;
wire _8548_;
wire _8549_;
wire _8550_;
wire _8551_;
wire _8552_;
wire _8553_;
wire _8554_;
wire _8555_;
wire _8556_;
wire _8557_;
wire _8558_;
wire _8559_;
wire _8560_;
wire _8561_;
wire _8562_;
wire _8563_;
wire _8564_;
wire _8565_;
wire _8566_;
wire _8567_;
wire _8568_;
wire _8569_;
wire _8570_;
wire _8571_;
wire _8572_;
wire _8573_;
wire _8574_;
wire _8575_;
wire _8576_;
wire _8577_;
wire _8578_;
wire _8579_;
wire _8580_;
wire _8581_;
wire _8582_;
wire _8583_;
wire _8584_;
wire _8585_;
wire _8586_;
wire _8587_;
wire _8588_;
wire _8589_;
wire _8590_;
wire _8591_;
wire _8592_;
wire _8593_;
wire _8594_;
wire _8595_;
wire _8596_;
wire _8597_;
wire _8598_;
wire _8599_;
wire _8600_;
wire _8601_;
wire _8602_;
wire _8603_;
wire _8604_;
wire _8605_;
wire _8606_;
wire _8607_;
wire _8608_;
wire _8609_;
wire _8610_;
wire _8611_;
wire _8612_;
wire _8613_;
wire _8614_;
wire _8615_;
wire _8616_;
wire _8617_;
wire _8618_;
wire _8619_;
wire _8620_;
wire _8621_;
wire _8622_;
wire _8623_;
wire _8624_;
wire _8625_;
wire _8626_;
wire _8627_;
wire _8628_;
wire _8629_;
wire _8630_;
wire _8631_;
wire _8632_;
wire _8633_;
wire _8634_;
wire _8635_;
wire _8636_;
wire _8637_;
wire _8638_;
wire _8639_;
wire _8640_;
wire _8641_;
wire _8642_;
wire _8643_;
wire _8644_;
wire _8645_;
wire _8646_;
wire _8647_;
wire _8648_;
wire _8649_;
wire _8650_;
wire _8651_;
wire _8652_;
wire _8653_;
wire _8654_;
wire _8655_;
wire _8656_;
wire _8657_;
wire _8658_;
wire _8659_;
wire _8660_;
wire _8661_;
wire _8662_;
wire _8663_;
wire _8664_;
wire _8665_;
wire _8666_;
wire _8667_;
wire _8668_;
wire _8669_;
wire _8670_;
wire _8671_;
wire _8672_;
wire _8673_;
wire _8674_;
wire _8675_;
wire _8676_;
wire _8677_;
wire _8678_;
wire _8679_;
wire _8680_;
wire _8681_;
wire _8682_;
wire _8683_;
wire _8684_;
wire _8685_;
wire _8686_;
wire _8687_;
wire _8688_;
wire _8689_;
wire _8690_;
wire _8691_;
wire _8692_;
wire _8693_;
wire _8694_;
wire _8695_;
wire _8696_;
wire _8697_;
wire _8698_;
wire _8699_;
wire _8700_;
wire _8701_;
wire _8702_;
wire _8703_;
wire _8704_;
wire _8705_;
wire _8706_;
wire _8707_;
wire _8708_;
wire _8709_;
wire _8710_;
wire _8711_;
wire _8712_;
wire _8713_;
wire _8714_;
wire _8715_;
wire _8716_;
wire _8717_;
wire _8718_;
wire _8719_;
wire _8720_;
wire _8721_;
wire _8722_;
wire _8723_;
wire _8724_;
wire _8725_;
wire _8726_;
wire _8727_;
wire _8728_;
wire _8729_;
wire _8730_;
wire _8731_;
wire _8732_;
wire _8733_;
wire _8734_;
wire _8735_;
wire _8736_;
wire _8737_;
wire _8738_;
wire _8739_;
wire _8740_;
wire _8741_;
wire _8742_;
wire _8743_;
wire _8744_;
wire _8745_;
wire _8746_;
wire _8747_;
wire _8748_;
wire _8749_;
wire _8750_;
wire _8751_;
wire _8752_;
wire _8753_;
wire _8754_;
wire _8755_;
wire _8756_;
wire _8757_;
wire _8758_;
wire _8759_;
wire _8760_;
wire _8761_;
wire _8762_;
wire _8763_;
wire _8764_;
wire _8765_;
wire _8766_;
wire _8767_;
wire _8768_;
wire _8769_;
wire _8770_;
wire _8771_;
wire _8772_;
wire _8773_;
wire _8774_;
wire _8775_;
wire _8776_;
wire _8777_;
wire _8778_;
wire _8779_;
wire _8780_;
wire _8781_;
wire _8782_;
wire _8783_;
wire _8784_;
wire _8785_;
wire _8786_;
wire _8787_;
wire _8788_;
wire _8789_;
wire _8790_;
wire _8791_;
wire _8792_;
wire _8793_;
wire _8794_;
wire _8795_;
wire _8796_;
wire _8797_;
wire _8798_;
wire _8799_;
wire _8800_;
wire _8801_;
wire _8802_;
wire _8803_;
wire _8804_;
wire _8805_;
wire _8806_;
wire _8807_;
wire _8808_;
wire _8809_;
wire _8810_;
wire _8811_;
wire _8812_;
wire _8813_;
wire _8814_;
wire _8815_;
wire _8816_;
wire _8817_;
wire _8818_;
wire _8819_;
wire _8820_;
wire _8821_;
wire _8822_;
wire _8823_;
wire _8824_;
wire _8825_;
wire _8826_;
wire _8827_;
wire _8828_;
wire _8829_;
wire _8830_;
wire _8831_;
wire _8832_;
wire _8833_;
wire _8834_;
wire _8835_;
wire _8836_;
wire _8837_;
wire _8838_;
wire _8839_;
wire _8840_;
wire _8841_;
wire _8842_;
wire _8843_;
wire _8844_;
wire _8845_;
wire _8846_;
wire _8847_;
wire _8848_;
wire _8849_;
wire _8850_;
wire _8851_;
wire _8852_;
wire _8853_;
wire _8854_;
wire _8855_;
wire _8856_;
wire _8857_;
wire _8858_;
wire _8859_;
wire _8860_;
wire _8861_;
wire _8862_;
wire _8863_;
wire _8864_;
wire _8865_;
wire _8866_;
wire _8867_;
wire _8868_;
wire _8869_;
wire _8870_;
wire _8871_;
wire _8872_;
wire _8873_;
wire _8874_;
wire _8875_;
wire _8876_;
wire _8877_;
wire _8878_;
wire _8879_;
wire _8880_;
wire _8881_;
wire _8882_;
wire _8883_;
wire _8884_;
wire _8885_;
wire _8886_;
wire _8887_;
wire _8888_;
wire _8889_;
wire _8890_;
wire _8891_;
wire _8892_;
wire _8893_;
wire _8894_;
wire _8895_;
wire _8896_;
wire _8897_;
wire _8898_;
wire _8899_;
wire _8900_;
wire _8901_;
wire _8902_;
wire _8903_;
wire _8904_;
wire _8905_;
wire _8906_;
wire _8907_;
wire _8908_;
wire _8909_;
wire _8910_;
wire _8911_;
wire _8912_;
wire _8913_;
wire _8914_;
wire _8915_;
wire _8916_;
wire _8917_;
wire _8918_;
wire _8919_;
wire _8920_;
wire _8921_;
wire _8922_;
wire _8923_;
wire _8924_;
wire _8925_;
wire _8926_;
wire _8927_;
wire _8928_;
wire _8929_;
wire _8930_;
wire _8931_;
wire _8932_;
wire _8933_;
wire _8934_;
wire _8935_;
wire _8936_;
wire _8937_;
wire _8938_;
wire _8939_;
wire _8940_;
wire _8941_;
wire _8942_;
wire _8943_;
wire _8944_;
wire _8945_;
wire _8946_;
wire _8947_;
wire _8948_;
wire _8949_;
wire _8950_;
wire _8951_;
wire _8952_;
wire _8953_;
wire _8954_;
wire _8955_;
wire _8956_;
wire _8957_;
wire _8958_;
wire _8959_;
wire _8960_;
wire _8961_;
wire _8962_;
wire _8963_;
wire _8964_;
wire _8965_;
wire _8966_;
wire _8967_;
wire _8968_;
wire _8969_;
wire _8970_;
wire _8971_;
wire _8972_;
wire _8973_;
wire _8974_;
wire _8975_;
wire _8976_;
wire _8977_;
wire _8978_;
wire _8979_;
wire _8980_;
wire _8981_;
wire _8982_;
wire _8983_;
wire _8984_;
wire _8985_;
wire _8986_;
wire _8987_;
wire _8988_;
wire _8989_;
wire _8990_;
wire _8991_;
wire _8992_;
wire _8993_;
wire _8994_;
wire _8995_;
wire _8996_;
wire _8997_;
wire _8998_;
wire _8999_;
wire _9000_;
wire _9001_;
wire _9002_;
wire _9003_;
wire _9004_;
wire _9005_;
wire _9006_;
wire _9007_;
wire _9008_;
wire _9009_;
wire _9010_;
wire _9011_;
wire _9012_;
wire _9013_;
wire _9014_;
wire _9015_;
wire _9016_;
wire _9017_;
wire _9018_;
wire _9019_;
wire _9020_;
wire _9021_;
wire _9022_;
wire _9023_;
wire _9024_;
wire _9025_;
wire _9026_;
wire _9027_;
wire _9028_;
wire _9029_;
wire _9030_;
wire _9031_;
wire _9032_;
wire _9033_;
wire _9034_;
wire _9035_;
wire _9036_;
wire _9037_;
wire _9038_;
wire _9039_;
wire _9040_;
wire _9041_;
wire _9042_;
wire _9043_;
wire _9044_;
wire _9045_;
wire _9046_;
wire _9047_;
wire _9048_;
wire _9049_;
wire _9050_;
wire _9051_;
wire _9052_;
wire _9053_;
wire _9054_;
wire _9055_;
wire _9056_;
wire _9057_;
wire _9058_;
wire _9059_;
wire _9060_;
wire _9061_;
wire _9062_;
wire _9063_;
wire _9064_;
wire _9065_;
wire _9066_;
wire _9067_;
wire _9068_;
wire _9069_;
wire _9070_;
wire _9071_;
wire _9072_;
wire _9073_;
wire _9074_;
wire _9075_;
wire _9076_;
wire _9077_;
wire _9078_;
wire _9079_;
wire _9080_;
wire _9081_;
wire _9082_;
wire _9083_;
wire _9084_;
wire _9085_;
wire _9086_;
wire _9087_;
wire _9088_;
wire _9089_;
wire _9090_;
wire _9091_;
wire _9092_;
wire _9093_;
wire _9094_;
wire _9095_;
wire _9096_;
wire _9097_;
wire _9098_;
wire _9099_;
wire _9100_;
wire _9101_;
wire _9102_;
wire _9103_;
wire _9104_;
wire _9105_;
wire _9106_;
wire _9107_;
wire _9108_;
wire _9109_;
wire _9110_;
wire _9111_;
wire _9112_;
wire _9113_;
wire _9114_;
wire _9115_;
wire _9116_;
wire _9117_;
wire _9118_;
wire _9119_;
wire _9120_;
wire _9121_;
wire _9122_;
wire _9123_;
wire _9124_;
wire _9125_;
wire _9126_;
wire _9127_;
wire _9128_;
wire _9129_;
wire _9130_;
wire _9131_;
wire _9132_;
wire _9133_;
wire _9134_;
wire _9135_;
wire _9136_;
wire _9137_;
wire _9138_;
wire _9139_;
wire _9140_;
wire _9141_;
wire _9142_;
wire _9143_;
wire _9144_;
wire _9145_;
wire _9146_;
wire _9147_;
wire _9148_;
wire _9149_;
wire _9150_;
wire _9151_;
wire _9152_;
wire _9153_;
wire _9154_;
wire _9155_;
wire _9156_;
wire _9157_;
wire _9158_;
wire _9159_;
wire _9160_;
wire _9161_;
wire _9162_;
wire _9163_;
wire _9164_;
wire _9165_;
wire _9166_;
wire _9167_;
wire _9168_;
wire _9169_;
wire _9170_;
wire _9171_;
wire _9172_;
wire _9173_;
wire _9174_;
wire _9175_;
wire _9176_;
wire _9177_;
wire _9178_;
wire _9179_;
wire _9180_;
wire _9181_;
wire _9182_;
wire _9183_;
wire _9184_;
wire _9185_;
wire _9186_;
wire _9187_;
wire _9188_;
wire _9189_;
wire _9190_;
wire _9191_;
wire _9192_;
wire _9193_;
wire _9194_;
wire _9195_;
wire _9196_;
wire _9197_;
wire _9198_;
wire _9199_;
wire _9200_;
wire _9201_;
wire _9202_;
wire _9203_;
wire _9204_;
wire _9205_;
wire _9206_;
wire _9207_;
wire _9208_;
wire _9209_;
wire _9210_;
wire _9211_;
wire _9212_;
wire _9213_;
wire _9214_;
wire _9215_;
wire _9216_;
wire _9217_;
wire _9218_;
wire _9219_;
wire _9220_;
wire _9221_;
wire _9222_;
wire _9223_;
wire _9224_;
wire _9225_;
wire _9226_;
wire _9227_;
wire _9228_;
wire _9229_;
wire _9230_;
wire _9231_;
wire _9232_;
wire _9233_;
wire _9234_;
wire _9235_;
wire _9236_;
wire _9237_;
wire _9238_;
wire _9239_;
wire _9240_;
wire _9241_;
wire _9242_;
wire _9243_;
wire _9244_;
wire _9245_;
wire _9246_;
wire _9247_;
wire _9248_;
wire _9249_;
wire _9250_;
wire _9251_;
wire _9252_;
wire _9253_;
wire _9254_;
wire _9255_;
wire _9256_;
wire _9257_;
wire _9258_;
wire _9259_;
wire _9260_;
wire _9261_;
wire _9262_;
wire _9263_;
wire _9264_;
wire _9265_;
wire _9266_;
wire _9267_;
wire _9268_;
wire _9269_;
wire _9270_;
wire _9271_;
wire _9272_;
wire _9273_;
wire _9274_;
wire _9275_;
wire _9276_;
wire _9277_;
wire _9278_;
wire _9279_;
wire _9280_;
wire _9281_;
wire _9282_;
wire _9283_;
wire _9284_;
wire _9285_;
wire _9286_;
wire _9287_;
wire _9288_;
wire _9289_;
wire _9290_;
wire _9291_;
wire _9292_;
wire _9293_;
wire _9294_;
wire _9295_;
wire _9296_;
wire _9297_;
wire _9298_;
wire _9299_;
wire _9300_;
wire _9301_;
wire _9302_;
wire _9303_;
wire _9304_;
wire _9305_;
wire _9306_;
wire _9307_;
wire _9308_;
wire _9309_;
wire _9310_;
wire _9311_;
wire _9312_;
wire _9313_;
wire _9314_;
wire _9315_;
wire _9316_;
wire _9317_;
wire _9318_;
wire _9319_;
wire _9320_;
wire _9321_;
wire _9322_;
wire _9323_;
wire _9324_;
wire _9325_;
wire _9326_;
wire _9327_;
wire _9328_;
wire _9329_;
wire _9330_;
wire _9331_;
wire _9332_;
wire _9333_;
wire _9334_;
wire _9335_;
wire _9336_;
wire _9337_;
wire _9338_;
wire _9339_;
wire _9340_;
wire _9341_;
wire _9342_;
wire _9343_;
wire _9344_;
wire _9345_;
wire _9346_;
wire _9347_;
wire _9348_;
wire _9349_;
wire _9350_;
wire _9351_;
wire _9352_;
wire _9353_;
wire _9354_;
wire _9355_;
wire _9356_;
wire _9357_;
wire _9358_;
wire _9359_;
wire _9360_;
wire _9361_;
wire _9362_;
wire _9363_;
wire _9364_;
wire _9365_;
wire _9366_;
wire _9367_;
wire _9368_;
wire _9369_;
wire _9370_;
wire _9371_;
wire _9372_;
wire _9373_;
wire _9374_;
wire _9375_;
wire _9376_;
wire _9377_;
wire _9378_;
wire _9379_;
wire _9380_;
wire _9381_;
wire _9382_;
wire _9383_;
wire _9384_;
wire _9385_;
wire _9386_;
wire _9387_;
wire _9388_;
wire _9389_;
wire _9390_;
wire _9391_;
wire _9392_;
wire _9393_;
wire _9394_;
wire _9395_;
wire _9396_;
wire _9397_;
wire _9398_;
wire _9399_;
wire _9400_;
wire _9401_;
wire _9402_;
wire _9403_;
wire _9404_;
wire _9405_;
wire _9406_;
wire _9407_;
wire _9408_;
wire _9409_;
wire _9410_;
wire _9411_;
wire _9412_;
wire _9413_;
wire _9414_;
wire _9415_;
wire _9416_;
wire _9417_;
wire _9418_;
wire _9419_;
wire _9420_;
wire _9421_;
wire _9422_;
wire _9423_;
wire _9424_;
wire _9425_;
wire _9426_;
wire _9427_;
wire _9428_;
wire _9429_;
wire _9430_;
wire _9431_;
wire _9432_;
wire _9433_;
wire _9434_;
wire _9435_;
wire _9436_;
wire _9437_;
wire _9438_;
wire _9439_;
wire _9440_;
wire _9441_;
wire _9442_;
wire _9443_;
wire _9444_;
wire _9445_;
wire _9446_;
wire _9447_;
wire _9448_;
wire _9449_;
wire _9450_;
wire _9451_;
wire _9452_;
wire _9453_;
wire _9454_;
wire _9455_;
wire _9456_;
wire _9457_;
wire _9458_;
wire _9459_;
wire _9460_;
wire _9461_;
wire _9462_;
wire _9463_;
wire _9464_;
wire _9465_;
wire _9466_;
wire _9467_;
wire _9468_;
wire _9469_;
wire _9470_;
wire _9471_;
wire _9472_;
wire _9473_;
wire _9474_;
wire _9475_;
wire _9476_;
wire _9477_;
wire _9478_;
wire _9479_;
wire _9480_;
wire _9481_;
wire _9482_;
wire _9483_;
wire _9484_;
wire _9485_;
wire _9486_;
wire _9487_;
wire _9488_;
wire _9489_;
wire _9490_;
wire _9491_;
wire _9492_;
wire _9493_;
wire _9494_;
wire _9495_;
wire _9496_;
wire _9497_;
wire _9498_;
wire _9499_;
wire _9500_;
wire _9501_;
wire _9502_;
wire _9503_;
wire _9504_;
wire _9505_;
wire _9506_;
wire _9507_;
wire _9508_;
wire _9509_;
wire _9510_;
wire _9511_;
wire _9512_;
wire _9513_;
wire _9514_;
wire _9515_;
wire _9516_;
wire _9517_;
wire _9518_;
wire _9519_;
wire _9520_;
wire _9521_;
wire _9522_;
wire _9523_;
wire _9524_;
wire _9525_;
wire _9526_;
wire _9527_;
wire _9528_;
wire _9529_;
wire _9530_;
wire _9531_;
wire _9532_;
wire _9533_;
wire _9534_;
wire _9535_;
wire _9536_;
wire _9537_;
wire _9538_;
wire _9539_;
wire _9540_;
wire _9541_;
wire _9542_;
wire _9543_;
wire _9544_;
wire _9545_;
wire _9546_;
wire _9547_;
wire _9548_;
wire _9549_;
wire _9550_;
wire _9551_;
wire _9552_;
wire _9553_;
wire _9554_;
wire _9555_;
wire _9556_;
wire _9557_;
wire _9558_;
wire _9559_;
wire _9560_;
wire _9561_;
wire _9562_;
wire _9563_;
wire _9564_;
wire _9565_;
wire _9566_;
wire _9567_;
wire _9568_;
wire _9569_;
wire _9570_;
wire _9571_;
wire _9572_;
wire _9573_;
wire _9574_;
wire _9575_;
wire _9576_;
wire _9577_;
wire _9578_;
wire _9579_;
wire _9580_;
wire _9581_;
wire _9582_;
wire _9583_;
wire _9584_;
wire _9585_;
wire _9586_;
wire _9587_;
wire _9588_;
wire _9589_;
wire _9590_;
wire _9591_;
wire _9592_;
wire _9593_;
wire _9594_;
wire _9595_;
wire _9596_;
wire _9597_;
wire _9598_;
wire _9599_;
wire _9600_;
wire _9601_;
wire _9602_;
wire _9603_;
wire _9604_;
wire _9605_;
wire _9606_;
wire _9607_;
wire _9608_;
wire _9609_;
wire _9610_;
wire _9611_;
wire _9612_;
wire _9613_;
wire _9614_;
wire _9615_;
wire _9616_;
wire _9617_;
wire _9618_;
wire _9619_;
wire _9620_;
wire _9621_;
wire _9622_;
wire _9623_;
wire _9624_;
wire _9625_;
wire _9626_;
wire _9627_;
wire _9628_;
wire _9629_;
wire _9630_;
wire _9631_;
wire _9632_;
wire _9633_;
wire _9634_;
wire _9635_;
wire _9636_;
wire _9637_;
wire _9638_;
wire _9639_;
wire _9640_;
wire _9641_;
wire _9642_;
wire _9643_;
wire _9644_;
wire _9645_;
wire _9646_;
wire _9647_;
wire _9648_;
wire _9649_;
wire _9650_;
wire _9651_;
wire _9652_;
wire _9653_;
wire _9654_;
wire _9655_;
wire _9656_;
wire _9657_;
wire _9658_;
wire _9659_;
wire _9660_;
wire _9661_;
wire _9662_;
wire _9663_;
wire _9664_;
wire _9665_;
wire _9666_;
wire _9667_;
wire _9668_;
wire _9669_;
wire _9670_;
wire _9671_;
wire _9672_;
wire _9673_;
wire _9674_;
wire _9675_;
wire _9676_;
wire _9677_;
wire _9678_;
wire _9679_;
wire _9680_;
wire _9681_;
wire _9682_;
wire _9683_;
wire _9684_;
wire _9685_;
wire _9686_;
wire _9687_;
wire _9688_;
wire _9689_;
wire _9690_;
wire _9691_;
wire _9692_;
wire _9693_;
wire _9694_;
wire _9695_;
wire _9696_;
wire _9697_;
wire _9698_;
wire _9699_;
wire _9700_;
wire _9701_;
wire _9702_;
wire _9703_;
wire _9704_;
wire _9705_;
wire _9706_;
wire _9707_;
wire _9708_;
wire _9709_;
wire _9710_;
wire _9711_;
wire _9712_;
wire _9713_;
wire _9714_;
wire _9715_;
wire _9716_;
wire _9717_;
wire _9718_;
wire _9719_;
wire _9720_;
wire _9721_;
wire _9722_;
wire _9723_;
wire _9724_;
wire _9725_;
wire _9726_;
wire _9727_;
wire _9728_;
wire _9729_;
wire _9730_;
wire _9731_;
wire _9732_;
wire _9733_;
wire _9734_;
wire _9735_;
wire _9736_;
wire _9737_;
wire _9738_;
wire _9739_;
wire _9740_;
wire _9741_;
wire _9742_;
wire _9743_;
wire _9744_;
wire _9745_;
wire _9746_;
wire _9747_;
wire _9748_;
wire _9749_;
wire _9750_;
wire _9751_;
wire _9752_;
wire _9753_;
wire _9754_;
wire _9755_;
wire _9756_;
wire _9757_;
wire _9758_;
wire _9759_;
wire _9760_;
wire _9761_;
wire _9762_;
wire _9763_;
wire _9764_;
wire _9765_;
wire _9766_;
wire _9767_;
wire _9768_;
wire _9769_;
wire _9770_;
wire _9771_;
wire _9772_;
wire _9773_;
wire _9774_;
wire _9775_;
wire _9776_;
wire _9777_;
wire _9778_;
wire _9779_;
wire _9780_;
wire _9781_;
wire _9782_;
wire _9783_;
wire _9784_;
wire _9785_;
wire _9786_;
wire _9787_;
wire _9788_;
wire _9789_;
wire _9790_;
wire _9791_;
wire _9792_;
wire _9793_;
wire _9794_;
wire _9795_;
wire _9796_;
wire _9797_;
wire _9798_;
wire _9799_;
wire _9800_;
wire _9801_;
wire _9802_;
wire _9803_;
wire _9804_;
wire _9805_;
wire _9806_;
wire _9807_;
wire _9808_;
wire _9809_;
wire _9810_;
wire _9811_;
wire _9812_;
wire _9813_;
wire _9814_;
wire _9815_;
wire _9816_;
wire _9817_;
wire _9818_;
wire _9819_;
wire _9820_;
wire _9821_;
wire _9822_;
wire _9823_;
wire _9824_;
wire _9825_;
wire _9826_;
wire _9827_;
wire _9828_;
wire _9829_;
wire _9830_;
wire _9831_;
wire _9832_;
wire _9833_;
wire _9834_;
wire _9835_;
wire _9836_;
wire _9837_;
wire _9838_;
wire _9839_;
wire _9840_;
wire _9841_;
wire _9842_;
wire _9843_;
wire _9844_;
wire _9845_;
wire _9846_;
wire _9847_;
wire _9848_;
wire _9849_;
wire _9850_;
wire _9851_;
wire _9852_;
wire _9853_;
wire _9854_;
wire _9855_;
wire _9856_;
wire _9857_;
wire _9858_;
wire _9859_;
wire _9860_;
wire _9861_;
wire _9862_;
wire _9863_;
wire _9864_;
wire _9865_;
wire _9866_;
wire _9867_;
wire _9868_;
wire _9869_;
wire _9870_;
wire _9871_;
wire _9872_;
wire _9873_;
wire _9874_;
wire _9875_;
wire _9876_;
wire _9877_;
wire _9878_;
wire _9879_;
wire _9880_;
wire _9881_;
wire _9882_;
wire _9883_;
wire _9884_;
wire _9885_;
wire _9886_;
wire _9887_;
wire _9888_;
wire _9889_;
wire _9890_;
wire _9891_;
wire _9892_;
wire _9893_;
wire _9894_;
wire _9895_;
wire _9896_;
wire _9897_;
wire _9898_;
wire _9899_;
wire _9900_;
wire _9901_;
wire _9902_;
wire _9903_;
wire _9904_;
wire _9905_;
wire _9906_;
wire _9907_;
wire _9908_;
wire _9909_;
wire _9910_;
wire _9911_;
wire _9912_;
wire _9913_;
wire _9914_;
wire _9915_;
wire _9916_;
wire _9917_;
wire _9918_;
wire _9919_;
wire _9920_;
wire _9921_;
wire _9922_;
wire _9923_;
wire _9924_;
wire _9925_;
wire _9926_;
wire _9927_;
wire _9928_;
wire _9929_;
wire _9930_;
wire _9931_;
wire _9932_;
wire _9933_;
wire _9934_;
wire _9935_;
wire _9936_;
wire _9937_;
wire _9938_;
wire _9939_;
wire _9940_;
wire _9941_;
wire _9942_;
wire _9943_;
wire _9944_;
wire _9945_;
wire _9946_;
wire _9947_;
wire _9948_;
wire _9949_;
wire _9950_;
wire _9951_;
wire _9952_;
wire _9953_;
wire _9954_;
wire _9955_;
wire _9956_;
wire _9957_;
wire _9958_;
wire _9959_;
wire _9960_;
wire _9961_;
wire _9962_;
wire _9963_;
wire _9964_;
wire _9965_;
wire _9966_;
wire _9967_;
wire _9968_;
wire _9969_;
wire _9970_;
wire _9971_;
wire _9972_;
wire _9973_;
wire _9974_;
wire _9975_;
wire _9976_;
wire _9977_;
wire _9978_;
wire _9979_;
wire _9980_;
wire _9981_;
wire _9982_;
wire _9983_;
wire _9984_;
wire _9985_;
wire _9986_;
wire _9987_;
wire _9988_;
wire _9989_;
wire _9990_;
wire _9991_;
wire _9992_;
wire _9993_;
wire _9994_;
wire _9995_;
wire _9996_;
wire _9997_;
wire _9998_;
wire _9999_;
wire _10000_;
wire _10001_;
wire _10002_;
wire _10003_;
wire _10004_;
wire _10005_;
wire _10006_;
wire _10007_;
wire _10008_;
wire _10009_;
wire _10010_;
wire _10011_;
wire _10012_;
wire _10013_;
wire _10014_;
wire _10015_;
wire _10016_;
wire _10017_;
wire _10018_;
wire _10019_;
wire _10020_;
wire _10021_;
wire _10022_;
wire _10023_;
wire _10024_;
wire _10025_;
wire _10026_;
wire _10027_;
wire _10028_;
wire _10029_;
wire _10030_;
wire _10031_;
wire _10032_;
wire _10033_;
wire _10034_;
wire _10035_;
wire _10036_;
wire _10037_;
wire _10038_;
wire _10039_;
wire _10040_;
wire _10041_;
wire _10042_;
wire _10043_;
wire _10044_;
wire _10045_;
wire _10046_;
wire _10047_;
wire _10048_;
wire _10049_;
wire _10050_;
wire _10051_;
wire _10052_;
wire _10053_;
wire _10054_;
wire _10055_;
wire _10056_;
wire _10057_;
wire _10058_;
wire _10059_;
wire _10060_;
wire _10061_;
wire _10062_;
wire _10063_;
wire _10064_;
wire _10065_;
wire _10066_;
wire _10067_;
wire _10068_;
wire _10069_;
wire _10070_;
wire _10071_;
wire _10072_;
wire _10073_;
wire _10074_;
wire _10075_;
wire _10076_;
wire _10077_;
wire _10078_;
wire _10079_;
wire _10080_;
wire _10081_;
wire _10082_;
wire _10083_;
wire _10084_;
wire _10085_;
wire _10086_;
wire _10087_;
wire _10088_;
wire _10089_;
wire _10090_;
wire _10091_;
wire _10092_;
wire _10093_;
wire _10094_;
wire _10095_;
wire _10096_;
wire _10097_;
wire _10098_;
wire _10099_;
wire _10100_;
wire _10101_;
wire _10102_;
wire _10103_;
wire _10104_;
wire _10105_;
wire _10106_;
wire _10107_;
wire _10108_;
wire _10109_;
wire _10110_;
wire _10111_;
wire _10112_;
wire _10113_;
wire _10114_;
wire _10115_;
wire _10116_;
wire _10117_;
wire _10118_;
wire _10119_;
wire _10120_;
wire _10121_;
wire _10122_;
wire _10123_;
wire _10124_;
wire _10125_;
wire _10126_;
wire _10127_;
wire _10128_;
wire _10129_;
wire _10130_;
wire _10131_;
wire _10132_;
wire _10133_;
wire _10134_;
wire _10135_;
wire _10136_;
wire _10137_;
wire _10138_;
wire _10139_;
wire _10140_;
wire _10141_;
wire _10142_;
wire _10143_;
wire _10144_;
wire _10145_;
wire _10146_;
wire _10147_;
wire _10148_;
wire _10149_;
wire _10150_;
wire _10151_;
wire _10152_;
wire _10153_;
wire _10154_;
wire _10155_;
wire _10156_;
wire _10157_;
wire _10158_;
wire _10159_;
wire _10160_;
wire _10161_;
wire _10162_;
wire _10163_;
wire _10164_;
wire _10165_;
wire _10166_;
wire _10167_;
wire _10168_;
wire _10169_;
wire _10170_;
wire _10171_;
wire _10172_;
wire _10173_;
wire _10174_;
wire _10175_;
wire _10176_;
wire _10177_;
wire _10178_;
wire _10179_;
wire _10180_;
wire _10181_;
wire _10182_;
wire _10183_;
wire _10184_;
wire _10185_;
wire _10186_;
wire _10187_;
wire _10188_;
wire _10189_;
wire _10190_;
wire _10191_;
wire _10192_;
wire _10193_;
wire _10194_;
wire _10195_;
wire _10196_;
wire _10197_;
wire _10198_;
wire _10199_;
wire _10200_;
wire _10201_;
wire _10202_;
wire _10203_;
wire _10204_;
wire _10205_;
wire _10206_;
wire _10207_;
wire _10208_;
wire _10209_;
wire _10210_;
wire _10211_;
wire _10212_;
wire _10213_;
wire _10214_;
wire _10215_;
wire _10216_;
wire _10217_;
wire _10218_;
wire _10219_;
wire _10220_;
wire _10221_;
wire _10222_;
wire _10223_;
wire _10224_;
wire _10225_;
wire _10226_;
wire _10227_;
wire _10228_;
wire _10229_;
wire _10230_;
wire _10231_;
wire _10232_;
wire _10233_;
wire _10234_;
wire _10235_;
wire _10236_;
wire _10237_;
wire _10238_;
wire _10239_;
wire _10240_;
wire _10241_;
wire _10242_;
wire _10243_;
wire _10244_;
wire _10245_;
wire _10246_;
wire _10247_;
wire _10248_;
wire _10249_;
wire _10250_;
wire _10251_;
wire _10252_;
wire _10253_;
wire _10254_;
wire _10255_;
wire _10256_;
wire _10257_;
wire _10258_;
wire _10259_;
wire _10260_;
wire _10261_;
wire _10262_;
wire _10263_;
wire _10264_;
wire _10265_;
wire _10266_;
wire _10267_;
wire _10268_;
wire _10269_;
wire _10270_;
wire _10271_;
wire _10272_;
wire _10273_;
wire _10274_;
wire _10275_;
wire _10276_;
wire _10277_;
wire _10278_;
wire _10279_;
wire _10280_;
wire _10281_;
wire _10282_;
wire _10283_;
wire _10284_;
wire _10285_;
wire _10286_;
wire _10287_;
wire _10288_;
wire _10289_;
wire _10290_;
wire _10291_;
wire _10292_;
wire _10293_;
wire _10294_;
wire _10295_;
wire _10296_;
wire _10297_;
wire _10298_;
wire _10299_;
wire _10300_;
wire _10301_;
wire _10302_;
wire _10303_;
wire _10304_;
wire _10305_;
wire _10306_;
wire _10307_;
wire _10308_;
wire _10309_;
wire _10310_;
wire _10311_;
wire _10312_;
wire _10313_;
wire _10314_;
wire _10315_;
wire _10316_;
wire _10317_;
wire _10318_;
wire _10319_;
wire _10320_;
wire _10321_;
wire _10322_;
wire _10323_;
wire _10324_;
wire _10325_;
wire _10326_;
wire _10327_;
wire _10328_;
wire _10329_;
wire _10330_;
wire _10331_;
wire _10332_;
wire _10333_;
wire _10334_;
wire _10335_;
wire _10336_;
wire _10337_;
wire _10338_;
wire _10339_;
wire _10340_;
wire _10341_;
wire _10342_;
wire _10343_;
wire _10344_;
wire _10345_;
wire _10346_;
wire _10347_;
wire _10348_;
wire _10349_;
wire _10350_;
wire _10351_;
wire _10352_;
wire _10353_;
wire _10354_;
wire _10355_;
wire _10356_;
wire _10357_;
wire _10358_;
wire _10359_;
wire _10360_;
wire _10361_;
wire _10362_;
wire _10363_;
wire _10364_;
wire _10365_;
wire _10366_;
wire _10367_;
wire _10368_;
wire _10369_;
wire _10370_;
wire _10371_;
wire _10372_;
wire _10373_;
wire _10374_;
wire _10375_;
wire _10376_;
wire _10377_;
wire _10378_;
wire _10379_;
wire _10380_;
wire _10381_;
wire _10382_;
wire _10383_;
wire _10384_;
wire _10385_;
wire _10386_;
wire _10387_;
wire _10388_;
wire _10389_;
wire _10390_;
wire _10391_;
wire _10392_;
wire _10393_;
wire _10394_;
wire _10395_;
wire _10396_;
wire _10397_;
wire _10398_;
wire _10399_;
wire _10400_;
wire _10401_;
wire _10402_;
wire _10403_;
wire _10404_;
wire _10405_;
wire _10406_;
wire _10407_;
wire _10408_;
wire _10409_;
wire _10410_;
wire _10411_;
wire _10412_;
wire _10413_;
wire _10414_;
wire _10415_;
wire _10416_;
wire _10417_;
wire _10418_;
wire _10419_;
wire _10420_;
wire _10421_;
wire _10422_;
wire _10423_;
wire _10424_;
wire _10425_;
wire _10426_;
wire _10427_;
wire _10428_;
wire _10429_;
wire _10430_;
wire _10431_;
wire _10432_;
wire _10433_;
wire _10434_;
wire _10435_;
wire _10436_;
wire _10437_;
wire _10438_;
wire _10439_;
wire _10440_;
wire _10441_;
wire _10442_;
wire _10443_;
wire _10444_;
wire _10445_;
wire _10446_;
wire _10447_;
wire _10448_;
wire _10449_;
wire _10450_;
wire _10451_;
wire _10452_;
wire _10453_;
wire _10454_;
wire _10455_;
wire _10456_;
wire _10457_;
wire _10458_;
wire _10459_;
wire _10460_;
wire _10461_;
wire _10462_;
wire _10463_;
wire _10464_;
wire _10465_;
wire _10466_;
wire _10467_;
wire _10468_;
wire _10469_;
wire _10470_;
wire _10471_;
wire _10472_;
wire _10473_;
wire _10474_;
wire _10475_;
wire _10476_;
wire _10477_;
wire _10478_;
wire _10479_;
wire _10480_;
wire _10481_;
wire _10482_;
wire _10483_;
wire _10484_;
wire _10485_;
wire _10486_;
wire _10487_;
wire _10488_;
wire _10489_;
wire _10490_;
wire _10491_;
wire _10492_;
wire _10493_;
wire _10494_;
wire _10495_;
wire _10496_;
wire _10497_;
wire _10498_;
wire _10499_;
wire _10500_;
wire _10501_;
wire _10502_;
wire _10503_;
wire _10504_;
wire _10505_;
wire _10506_;
wire _10507_;
wire _10508_;
wire _10509_;
wire _10510_;
wire _10511_;
wire _10512_;
wire _10513_;
wire _10514_;
wire _10515_;
wire _10516_;
wire _10517_;
wire _10518_;
wire _10519_;
wire _10520_;
wire _10521_;
wire _10522_;
wire _10523_;
wire _10524_;
wire _10525_;
wire _10526_;
wire _10527_;
wire _10528_;
wire _10529_;
wire _10530_;
wire _10531_;
wire _10532_;
wire _10533_;
wire _10534_;
wire _10535_;
wire _10536_;
wire _10537_;
wire _10538_;
wire _10539_;
wire _10540_;
wire _10541_;
wire _10542_;
wire _10543_;
wire _10544_;
wire _10545_;
wire _10546_;
wire _10547_;
wire _10548_;
wire _10549_;
wire _10550_;
wire _10551_;
wire _10552_;
wire _10553_;
wire _10554_;
wire _10555_;
wire _10556_;
wire _10557_;
wire _10558_;
wire _10559_;
wire _10560_;
wire _10561_;
wire _10562_;
wire _10563_;
wire _10564_;
wire _10565_;
wire _10566_;
wire _10567_;
wire _10568_;
wire _10569_;
wire _10570_;
wire _10571_;
wire _10572_;
wire _10573_;
wire _10574_;
wire _10575_;
wire _10576_;
wire _10577_;
wire _10578_;
wire _10579_;
wire _10580_;
wire _10581_;
wire _10582_;
wire _10583_;
wire _10584_;
wire _10585_;
wire _10586_;
wire _10587_;
wire _10588_;
wire _10589_;
wire _10590_;
wire _10591_;
wire _10592_;
wire _10593_;
wire _10594_;
wire _10595_;
wire _10596_;
wire _10597_;
wire _10598_;
wire _10599_;
wire _10600_;
wire _10601_;
wire _10602_;
wire _10603_;
wire _10604_;
wire _10605_;
wire _10606_;
wire _10607_;
wire _10608_;
wire _10609_;
wire _10610_;
wire _10611_;
wire _10612_;
wire _10613_;
wire _10614_;
wire _10615_;
wire _10616_;
wire _10617_;
wire _10618_;
wire _10619_;
wire _10620_;
wire _10621_;
wire _10622_;
wire _10623_;
wire _10624_;
wire _10625_;
wire _10626_;
wire _10627_;
wire _10628_;
wire _10629_;
wire _10630_;
wire _10631_;
wire _10632_;
wire _10633_;
wire _10634_;
wire _10635_;
wire _10636_;
wire _10637_;
wire _10638_;
wire _10639_;
wire _10640_;
wire _10641_;
wire _10642_;
wire _10643_;
wire _10644_;
wire _10645_;
wire _10646_;
wire _10647_;
wire _10648_;
wire _10649_;
wire _10650_;
wire _10651_;
wire _10652_;
wire _10653_;
wire _10654_;
wire _10655_;
wire _10656_;
wire _10657_;
wire _10658_;
wire _10659_;
wire _10660_;
wire _10661_;
wire _10662_;
wire _10663_;
wire _10664_;
wire _10665_;
wire _10666_;
wire _10667_;
wire _10668_;
wire _10669_;
wire _10670_;
wire _10671_;
wire _10672_;
wire _10673_;
wire _10674_;
wire _10675_;
wire _10676_;
wire _10677_;
wire _10678_;
wire _10679_;
wire _10680_;
wire _10681_;
wire _10682_;
wire _10683_;
wire _10684_;
wire _10685_;
wire _10686_;
wire _10687_;
wire _10688_;
wire _10689_;
wire _10690_;
wire _10691_;
wire _10692_;
wire _10693_;
wire _10694_;
wire _10695_;
wire _10696_;
wire _10697_;
wire _10698_;
wire _10699_;
wire _10700_;
wire _10701_;
wire _10702_;
wire _10703_;
wire _10704_;
wire _10705_;
wire _10706_;
wire _10707_;
wire _10708_;
wire _10709_;
wire _10710_;
wire _10711_;
wire _10712_;
wire _10713_;
wire _10714_;
wire _10715_;
wire _10716_;
wire _10717_;
wire _10718_;
wire _10719_;
wire _10720_;
wire _10721_;
wire _10722_;
wire _10723_;
wire _10724_;
wire _10725_;
wire _10726_;
wire _10727_;
wire _10728_;
wire _10729_;
wire _10730_;
wire _10731_;
wire _10732_;
wire _10733_;
wire _10734_;
wire _10735_;
wire _10736_;
wire _10737_;
wire _10738_;
wire _10739_;
wire _10740_;
wire _10741_;
wire _10742_;
wire _10743_;
wire _10744_;
wire _10745_;
wire _10746_;
wire _10747_;
wire _10748_;
wire _10749_;
wire _10750_;
wire _10751_;
wire _10752_;
wire _10753_;
wire _10754_;
wire _10755_;
wire _10756_;
wire _10757_;
wire _10758_;
wire _10759_;
wire _10760_;
wire _10761_;
wire _10762_;
wire _10763_;
wire _10764_;
wire _10765_;
wire _10766_;
wire _10767_;
wire _10768_;
wire _10769_;
wire _10770_;
wire _10771_;
wire _10772_;
wire _10773_;
wire _10774_;
wire _10775_;
wire _10776_;
wire _10777_;
wire _10778_;
wire _10779_;
wire _10780_;
wire _10781_;
wire _10782_;
wire _10783_;
wire _10784_;
wire _10785_;
wire _10786_;
wire _10787_;
wire _10788_;
wire _10789_;
wire _10790_;
wire _10791_;
wire _10792_;
wire _10793_;
wire _10794_;
wire _10795_;
wire _10796_;
wire _10797_;
wire _10798_;
wire _10799_;
wire _10800_;
wire _10801_;
wire _10802_;
wire _10803_;
wire _10804_;
wire _10805_;
wire _10806_;
wire _10807_;
wire _10808_;
wire _10809_;
wire _10810_;
wire _10811_;
wire _10812_;
wire _10813_;
wire _10814_;
wire _10815_;
wire _10816_;
wire _10817_;
wire _10818_;
wire _10819_;
wire _10820_;
wire _10821_;
wire _10822_;
wire _10823_;
wire _10824_;
wire _10825_;
wire _10826_;
wire _10827_;
wire _10828_;
wire _10829_;
wire _10830_;
wire _10831_;
wire _10832_;
wire _10833_;
wire _10834_;
wire _10835_;
wire _10836_;
wire _10837_;
wire _10838_;
wire _10839_;
wire _10840_;
wire _10841_;
wire _10842_;
wire _10843_;
wire _10844_;
wire _10845_;
wire _10846_;
wire _10847_;
wire _10848_;
wire _10849_;
wire _10850_;
wire _10851_;
wire _10852_;
wire _10853_;
wire _10854_;
wire _10855_;
wire _10856_;
wire _10857_;
wire _10858_;
wire _10859_;
wire _10860_;
wire _10861_;
wire _10862_;
wire _10863_;
wire _10864_;
wire _10865_;
wire _10866_;
wire _10867_;
wire _10868_;
wire _10869_;
wire _10870_;
wire _10871_;
wire _10872_;
wire _10873_;
wire _10874_;
wire _10875_;
wire _10876_;
wire _10877_;
wire _10878_;
wire _10879_;
wire _10880_;
wire _10881_;
wire _10882_;
wire _10883_;
wire _10884_;
wire _10885_;
wire _10886_;
wire _10887_;
wire _10888_;
wire _10889_;
wire _10890_;
wire _10891_;
wire _10892_;
wire _10893_;
wire _10894_;
wire _10895_;
wire _10896_;
wire _10897_;
wire _10898_;
wire _10899_;
wire _10900_;
wire _10901_;
wire _10902_;
wire _10903_;
wire _10904_;
wire _10905_;
wire _10906_;
wire _10907_;
wire _10908_;
wire _10909_;
wire _10910_;
wire _10911_;
wire _10912_;
wire _10913_;
wire _10914_;
wire _10915_;
wire _10916_;
wire _10917_;
wire _10918_;
wire _10919_;
wire _10920_;
wire _10921_;
wire _10922_;
wire _10923_;
wire _10924_;
wire _10925_;
wire _10926_;
wire _10927_;
wire _10928_;
wire _10929_;
wire _10930_;
wire _10931_;
wire _10932_;
wire _10933_;
wire _10934_;
wire _10935_;
wire _10936_;
wire _10937_;
wire _10938_;
wire _10939_;
wire _10940_;
wire _10941_;
wire _10942_;
wire _10943_;
wire _10944_;
wire _10945_;
wire _10946_;
wire _10947_;
wire _10948_;
wire _10949_;
wire _10950_;
wire _10951_;
wire _10952_;
wire _10953_;
wire _10954_;
wire _10955_;
wire _10956_;
wire _10957_;
wire _10958_;
wire _10959_;
wire _10960_;
wire _10961_;
wire _10962_;
wire _10963_;
wire _10964_;
wire _10965_;
wire _10966_;
wire _10967_;
wire _10968_;
wire _10969_;
wire _10970_;
wire _10971_;
wire _10972_;
wire _10973_;
wire _10974_;
wire _10975_;
wire _10976_;
wire _10977_;
wire _10978_;
wire _10979_;
wire _10980_;
wire _10981_;
wire _10982_;
wire _10983_;
wire _10984_;
wire _10985_;
wire _10986_;
wire _10987_;
wire _10988_;
wire _10989_;
wire _10990_;
wire _10991_;
wire _10992_;
wire _10993_;
wire _10994_;
wire _10995_;
wire _10996_;
wire _10997_;
wire _10998_;
wire _10999_;
wire _11000_;
wire _11001_;
wire _11002_;
wire _11003_;
wire _11004_;
wire _11005_;
wire _11006_;
wire _11007_;
wire _11008_;
wire _11009_;
wire _11010_;
wire _11011_;
wire _11012_;
wire _11013_;
wire _11014_;
wire _11015_;
wire _11016_;
wire _11017_;
wire _11018_;
wire _11019_;
wire _11020_;
wire _11021_;
wire _11022_;
wire _11023_;
wire _11024_;
wire _11025_;
wire _11026_;
wire _11027_;
wire _11028_;
wire _11029_;
wire _11030_;
wire _11031_;
wire _11032_;
wire _11033_;
wire _11034_;
wire _11035_;
wire _11036_;
wire _11037_;
wire _11038_;
wire _11039_;
wire _11040_;
wire _11041_;
wire _11042_;
wire _11043_;
wire _11044_;
wire _11045_;
wire _11046_;
wire _11047_;
wire _11048_;
wire _11049_;
wire _11050_;
wire _11051_;
wire _11052_;
wire _11053_;
wire _11054_;
wire _11055_;
wire _11056_;
wire _11057_;
wire _11058_;
wire _11059_;
wire _11060_;
wire _11061_;
wire _11062_;
wire _11063_;
wire _11064_;
wire _11065_;
wire _11066_;
wire _11067_;
wire _11068_;
wire _11069_;
wire _11070_;
wire _11071_;
wire _11072_;
wire _11073_;
wire _11074_;
wire _11075_;
wire _11076_;
wire _11077_;
wire _11078_;
wire _11079_;
wire _11080_;
wire _11081_;
wire _11082_;
wire _11083_;
wire _11084_;
wire _11085_;
wire _11086_;
wire _11087_;
wire _11088_;
wire _11089_;
wire _11090_;
wire _11091_;
wire _11092_;
wire _11093_;
wire _11094_;
wire _11095_;
wire _11096_;
wire _11097_;
wire _11098_;
wire _11099_;
wire _11100_;
wire _11101_;
wire _11102_;
wire _11103_;
wire _11104_;
wire _11105_;
wire _11106_;
wire _11107_;
wire _11108_;
wire _11109_;
wire _11110_;
wire _11111_;
wire _11112_;
wire _11113_;
wire _11114_;
wire _11115_;
wire _11116_;
wire _11117_;
wire _11118_;
wire _11119_;
wire _11120_;
wire _11121_;
wire _11122_;
wire _11123_;
wire _11124_;
wire _11125_;
wire _11126_;
wire _11127_;
wire _11128_;
wire _11129_;
wire _11130_;
wire _11131_;
wire _11132_;
wire _11133_;
wire _11134_;
wire _11135_;
wire _11136_;
wire _11137_;
wire _11138_;
wire _11139_;
wire _11140_;
wire _11141_;
wire _11142_;
wire _11143_;
wire _11144_;
wire _11145_;
wire _11146_;
wire _11147_;
wire _11148_;
wire _11149_;
wire _11150_;
wire _11151_;
wire _11152_;
wire _11153_;
wire _11154_;
wire _11155_;
wire _11156_;
wire _11157_;
wire _11158_;
wire _11159_;
wire _11160_;
wire _11161_;
wire _11162_;
wire _11163_;
wire _11164_;
wire _11165_;
wire _11166_;
wire _11167_;
wire _11168_;
wire _11169_;
wire _11170_;
wire _11171_;
wire _11172_;
wire _11173_;
wire _11174_;
wire _11175_;
wire _11176_;
wire _11177_;
wire _11178_;
wire _11179_;
wire _11180_;
wire _11181_;
wire _11182_;
wire _11183_;
wire _11184_;
wire _11185_;
wire _11186_;
wire _11187_;
wire _11188_;
wire _11189_;
wire _11190_;
wire _11191_;
wire _11192_;
wire _11193_;
wire _11194_;
wire _11195_;
wire _11196_;
wire _11197_;
wire _11198_;
wire _11199_;
wire _11200_;
wire _11201_;
wire _11202_;
wire _11203_;
wire _11204_;
wire _11205_;
wire _11206_;
wire _11207_;
wire _11208_;
wire _11209_;
wire _11210_;
wire _11211_;
wire _11212_;
wire _11213_;
wire _11214_;
wire _11215_;
wire _11216_;
wire _11217_;
wire _11218_;
wire _11219_;
wire _11220_;
wire _11221_;
wire _11222_;
wire _11223_;
wire _11224_;
wire _11225_;
wire _11226_;
wire _11227_;
wire _11228_;
wire _11229_;
wire _11230_;
wire _11231_;
wire _11232_;
wire _11233_;
wire _11234_;
wire _11235_;
wire _11236_;
wire _11237_;
wire _11238_;
wire _11239_;
wire _11240_;
wire _11241_;
wire _11242_;
wire _11243_;
wire _11244_;
wire _11245_;
wire _11246_;
wire _11247_;
wire _11248_;
wire _11249_;
wire _11250_;
wire _11251_;
wire _11252_;
wire _11253_;
wire _11254_;
wire _11255_;
wire _11256_;
wire _11257_;
wire _11258_;
wire _11259_;
wire _11260_;
wire _11261_;
wire _11262_;
wire _11263_;
wire _11264_;
wire _11265_;
wire _11266_;
wire _11267_;
wire _11268_;
wire _11269_;
wire _11270_;
wire _11271_;
wire _11272_;
wire _11273_;
wire _11274_;
wire _11275_;
wire _11276_;
wire _11277_;
wire _11278_;
wire _11279_;
wire _11280_;
wire _11281_;
wire _11282_;
wire _11283_;
wire _11284_;
wire _11285_;
wire _11286_;
wire _11287_;
wire _11288_;
wire _11289_;
wire _11290_;
wire _11291_;
wire _11292_;
wire _11293_;
wire _11294_;
wire _11295_;
wire _11296_;
wire _11297_;
wire _11298_;
wire _11299_;
wire _11300_;
wire _11301_;
wire _11302_;
wire _11303_;
wire _11304_;
wire _11305_;
wire _11306_;
wire _11307_;
wire _11308_;
wire _11309_;
wire _11310_;
wire _11311_;
wire _11312_;
wire _11313_;
wire _11314_;
wire _11315_;
wire _11316_;
wire _11317_;
wire _11318_;
wire _11319_;
wire _11320_;
wire _11321_;
wire _11322_;
wire _11323_;
wire _11324_;
wire _11325_;
wire _11326_;
wire _11327_;
wire _11328_;
wire _11329_;
wire _11330_;
wire _11331_;
wire _11332_;
wire _11333_;
wire _11334_;
wire _11335_;
wire _11336_;
wire _11337_;
wire _11338_;
wire _11339_;
wire _11340_;
wire _11341_;
wire _11342_;
wire _11343_;
wire _11344_;
wire _11345_;
wire _11346_;
wire _11347_;
wire _11348_;
wire _11349_;
wire _11350_;
wire _11351_;
wire _11352_;
wire _11353_;
wire _11354_;
wire _11355_;
wire _11356_;
wire _11357_;
wire _11358_;
wire _11359_;
wire _11360_;
wire _11361_;
wire _11362_;
wire _11363_;
wire _11364_;
wire _11365_;
wire _11366_;
wire _11367_;
wire _11368_;
wire _11369_;
wire _11370_;
wire _11371_;
wire _11372_;
wire _11373_;
wire _11374_;
wire _11375_;
wire _11376_;
wire _11377_;
wire _11378_;
wire _11379_;
wire _11380_;
wire _11381_;
wire _11382_;
wire _11383_;
wire _11384_;
wire _11385_;
wire _11386_;
wire _11387_;
wire _11388_;
wire _11389_;
wire _11390_;
wire _11391_;
wire _11392_;
wire _11393_;
wire _11394_;
wire _11395_;
wire _11396_;
wire _11397_;
wire _11398_;
wire _11399_;
wire _11400_;
wire _11401_;
wire _11402_;
wire _11403_;
wire _11404_;
wire _11405_;
wire _11406_;
wire _11407_;
wire _11408_;
wire _11409_;
wire _11410_;
wire _11411_;
wire _11412_;
wire _11413_;
wire _11414_;
wire _11415_;
wire _11416_;
wire _11417_;
wire _11418_;
wire _11419_;
wire _11420_;
wire _11421_;
wire _11422_;
wire _11423_;
wire _11424_;
wire _11425_;
wire _11426_;
wire _11427_;
wire _11428_;
wire _11429_;
wire _11430_;
wire _11431_;
wire _11432_;
wire _11433_;
wire _11434_;
wire _11435_;
wire _11436_;
wire _11437_;
wire _11438_;
wire _11439_;
wire _11440_;
wire _11441_;
wire _11442_;
wire _11443_;
wire _11444_;
wire _11445_;
wire _11446_;
wire _11447_;
wire _11448_;
wire _11449_;
wire _11450_;
wire _11451_;
wire _11452_;
wire _11453_;
wire _11454_;
wire _11455_;
wire _11456_;
wire _11457_;
wire _11458_;
wire _11459_;
wire _11460_;
wire _11461_;
wire _11462_;
wire _11463_;
wire _11464_;
wire _11465_;
wire _11466_;
wire _11467_;
wire _11468_;
wire _11469_;
wire _11470_;
wire _11471_;
wire _11472_;
wire _11473_;
wire _11474_;
wire _11475_;
wire _11476_;
wire _11477_;
wire _11478_;
wire _11479_;
wire _11480_;
wire _11481_;
wire _11482_;
wire _11483_;
wire _11484_;
wire _11485_;
wire _11486_;
wire _11487_;
wire _11488_;
wire _11489_;
wire _11490_;
wire _11491_;
wire _11492_;
wire _11493_;
wire _11494_;
wire _11495_;
wire _11496_;
wire _11497_;
wire _11498_;
wire _11499_;
wire _11500_;
wire _11501_;
wire _11502_;
wire _11503_;
wire _11504_;
wire _11505_;
wire _11506_;
wire _11507_;
wire _11508_;
wire _11509_;
wire _11510_;
wire _11511_;
wire _11512_;
wire _11513_;
wire _11514_;
wire _11515_;
wire _11516_;
wire _11517_;
wire _11518_;
wire _11519_;
wire _11520_;
wire _11521_;
wire _11522_;
wire _11523_;
wire _11524_;
wire _11525_;
wire _11526_;
wire _11527_;
wire _11528_;
wire _11529_;
wire _11530_;
wire _11531_;
wire _11532_;
wire _11533_;
wire _11534_;
wire _11535_;
wire _11536_;
wire _11537_;
wire _11538_;
wire _11539_;
wire _11540_;
wire _11541_;
wire _11542_;
wire _11543_;
wire _11544_;
wire _11545_;
wire _11546_;
wire _11547_;
wire _11548_;
wire _11549_;
wire _11550_;
wire _11551_;
wire _11552_;
wire _11553_;
wire _11554_;
wire _11555_;
wire _11556_;
wire _11557_;
wire _11558_;
wire _11559_;
wire _11560_;
wire _11561_;
wire _11562_;
wire _11563_;
wire _11564_;
wire _11565_;
wire _11566_;
wire _11567_;
wire _11568_;
wire _11569_;
wire _11570_;
wire _11571_;
wire _11572_;
wire _11573_;
wire _11574_;
wire _11575_;
wire _11576_;
wire _11577_;
wire _11578_;
wire _11579_;
wire _11580_;
wire _11581_;
wire _11582_;
wire _11583_;
wire _11584_;
wire _11585_;
wire _11586_;
wire _11587_;
wire _11588_;
wire _11589_;
wire _11590_;
wire _11591_;
wire _11592_;
wire _11593_;
wire _11594_;
wire _11595_;
wire _11596_;
wire _11597_;
wire _11598_;
wire _11599_;
wire _11600_;
wire _11601_;
wire _11602_;
wire _11603_;
wire _11604_;
wire _11605_;
wire _11606_;
wire _11607_;
wire _11608_;
wire _11609_;
wire _11610_;
wire _11611_;
wire _11612_;
wire _11613_;
wire _11614_;
wire _11615_;
wire _11616_;
wire _11617_;
wire _11618_;
wire _11619_;
wire _11620_;
wire _11621_;
wire _11622_;
wire _11623_;
wire _11624_;
wire _11625_;
wire _11626_;
wire _11627_;
wire _11628_;
wire _11629_;
wire _11630_;
wire _11631_;
wire _11632_;
wire _11633_;
wire _11634_;
wire _11635_;
wire _11636_;
wire _11637_;
wire _11638_;
wire _11639_;
wire _11640_;
wire _11641_;
wire _11642_;
wire _11643_;
wire _11644_;
wire _11645_;
wire _11646_;
wire _11647_;
wire _11648_;
wire _11649_;
wire _11650_;
wire _11651_;
wire _11652_;
wire _11653_;
wire _11654_;
wire _11655_;
wire _11656_;
wire _11657_;
wire _11658_;
wire _11659_;
wire _11660_;
wire _11661_;
wire _11662_;
wire _11663_;
wire _11664_;
wire _11665_;
wire _11666_;
wire _11667_;
wire _11668_;
wire _11669_;
wire _11670_;
wire _11671_;
wire _11672_;
wire _11673_;
wire _11674_;
wire _11675_;
wire _11676_;
wire _11677_;
wire _11678_;
wire _11679_;
wire _11680_;
wire _11681_;
wire _11682_;
wire _11683_;
wire _11684_;
wire _11685_;
wire _11686_;
wire _11687_;
wire _11688_;
wire _11689_;
wire _11690_;
wire _11691_;
wire _11692_;
wire _11693_;
wire _11694_;
wire _11695_;
wire _11696_;
wire _11697_;
wire _11698_;
wire _11699_;
wire _11700_;
wire _11701_;
wire _11702_;
wire _11703_;
wire _11704_;
wire _11705_;
wire _11706_;
wire _11707_;
wire _11708_;
wire _11709_;
wire _11710_;
wire _11711_;
wire _11712_;
wire _11713_;
wire _11714_;
wire _11715_;
wire _11716_;
wire _11717_;
wire _11718_;
wire _11719_;
wire _11720_;
wire _11721_;
wire _11722_;
wire _11723_;
wire _11724_;
wire _11725_;
wire _11726_;
wire _11727_;
wire _11728_;
wire _11729_;
wire _11730_;
wire _11731_;
wire _11732_;
wire _11733_;
wire _11734_;
wire _11735_;
wire _11736_;
wire _11737_;
wire _11738_;
wire _11739_;
wire _11740_;
wire _11741_;
wire _11742_;
wire _11743_;
wire _11744_;
wire _11745_;
wire _11746_;
wire _11747_;
wire _11748_;
wire _11749_;
wire _11750_;
wire _11751_;
wire _11752_;
wire _11753_;
wire _11754_;
wire _11755_;
wire _11756_;
wire _11757_;
wire _11758_;
wire _11759_;
wire _11760_;
wire _11761_;
wire _11762_;
wire _11763_;
wire _11764_;
wire _11765_;
wire _11766_;
wire _11767_;
wire _11768_;
wire _11769_;
wire _11770_;
wire _11771_;
wire _11772_;
wire _11773_;
wire _11774_;
wire _11775_;
wire _11776_;
wire _11777_;
wire _11778_;
wire _11779_;
wire _11780_;
wire _11781_;
wire _11782_;
wire _11783_;
wire _11784_;
wire _11785_;
wire _11786_;
wire _11787_;
wire _11788_;
wire _11789_;
wire _11790_;
wire _11791_;
wire _11792_;
wire _11793_;
wire _11794_;
wire _11795_;
wire _11796_;
wire _11797_;
wire _11798_;
wire _11799_;
wire _11800_;
wire _11801_;
wire _11802_;
wire _11803_;
wire _11804_;
wire _11805_;
wire _11806_;
wire _11807_;
wire _11808_;
wire _11809_;
wire _11810_;
wire _11811_;
wire _11812_;
wire _11813_;
wire _11814_;
wire _11815_;
wire _11816_;
wire _11817_;
wire _11818_;
wire _11819_;
wire _11820_;
wire _11821_;
wire _11822_;
wire _11823_;
wire _11824_;
wire _11825_;
wire _11826_;
wire _11827_;
wire _11828_;
wire _11829_;
wire _11830_;
wire _11831_;
wire _11832_;
wire _11833_;
wire _11834_;
wire _11835_;
wire _11836_;
wire _11837_;
wire _11838_;
wire _11839_;
wire _11840_;
wire _11841_;
wire _11842_;
wire _11843_;
wire _11844_;
wire _11845_;
wire _11846_;
wire _11847_;
wire _11848_;
wire _11849_;
wire _11850_;
wire _11851_;
wire _11852_;
wire _11853_;
wire _11854_;
wire _11855_;
wire _11856_;
wire _11857_;
wire _11858_;
wire _11859_;
wire _11860_;
wire _11861_;
wire _11862_;
wire _11863_;
wire _11864_;
wire _11865_;
wire _11866_;
wire _11867_;
wire _11868_;
wire _11869_;
wire _11870_;
wire _11871_;
wire _11872_;
wire _11873_;
wire _11874_;
wire _11875_;
wire _11876_;
wire _11877_;
wire _11878_;
wire _11879_;
wire _11880_;
wire _11881_;
wire _11882_;
wire _11883_;
wire _11884_;
wire _11885_;
wire _11886_;
wire _11887_;
wire _11888_;
wire _11889_;
wire _11890_;
wire _11891_;
wire _11892_;
wire _11893_;
wire _11894_;
wire _11895_;
wire _11896_;
wire _11897_;
wire _11898_;
wire _11899_;
wire _11900_;
wire _11901_;
wire _11902_;
wire _11903_;
wire _11904_;
wire _11905_;
wire _11906_;
wire _11907_;
wire _11908_;
wire _11909_;
wire _11910_;
wire _11911_;
wire _11912_;
wire _11913_;
wire _11914_;
wire _11915_;
wire _11916_;
wire _11917_;
wire _11918_;
wire _11919_;
wire _11920_;
wire _11921_;
wire _11922_;
wire _11923_;
wire _11924_;
wire _11925_;
wire _11926_;
wire _11927_;
wire _11928_;
wire _11929_;
wire _11930_;
wire _11931_;
wire _11932_;
wire _11933_;
wire _11934_;
wire _11935_;
wire _11936_;
wire _11937_;
wire _11938_;
wire _11939_;
wire _11940_;
wire _11941_;
wire _11942_;
wire _11943_;
wire _11944_;
wire _11945_;
wire _11946_;
wire _11947_;
wire _11948_;
wire _11949_;
wire _11950_;
wire _11951_;
wire _11952_;
wire _11953_;
wire _11954_;
wire _11955_;
wire _11956_;
wire _11957_;
wire _11958_;
wire _11959_;
wire _11960_;
wire _11961_;
wire _11962_;
wire _11963_;
wire _11964_;
wire _11965_;
wire _11966_;
wire _11967_;
wire _11968_;
wire _11969_;
wire _11970_;
wire _11971_;
wire _11972_;
wire _11973_;
wire _11974_;
wire _11975_;
wire _11976_;
wire _11977_;
wire _11978_;
wire _11979_;
wire _11980_;
wire _11981_;
wire _11982_;
wire _11983_;
wire _11984_;
wire _11985_;
wire _11986_;
wire _11987_;
wire _11988_;
wire _11989_;
wire _11990_;
wire _11991_;
wire _11992_;
wire _11993_;
wire _11994_;
wire _11995_;
wire _11996_;
wire _11997_;
wire _11998_;
wire _11999_;
wire _12000_;
wire _12001_;
wire _12002_;
wire _12003_;
wire _12004_;
wire _12005_;
wire _12006_;
wire _12007_;
wire _12008_;
wire _12009_;
wire _12010_;
wire _12011_;
wire _12012_;
wire _12013_;
wire _12014_;
wire _12015_;
wire _12016_;
wire _12017_;
wire _12018_;
wire _12019_;
wire _12020_;
wire _12021_;
wire _12022_;
wire _12023_;
wire _12024_;
wire _12025_;
wire _12026_;
wire _12027_;
wire _12028_;
wire _12029_;
wire _12030_;
wire _12031_;
wire _12032_;
wire _12033_;
wire _12034_;
wire _12035_;
wire _12036_;
wire _12037_;
wire _12038_;
wire _12039_;
wire _12040_;
wire _12041_;
wire _12042_;
wire _12043_;
wire _12044_;
wire _12045_;
wire _12046_;
wire _12047_;
wire _12048_;
wire _12049_;
wire _12050_;
wire _12051_;
wire _12052_;
wire _12053_;
wire _12054_;
wire _12055_;
wire _12056_;
wire _12057_;
wire _12058_;
wire _12059_;
wire _12060_;
wire _12061_;
wire _12062_;
wire _12063_;
wire _12064_;
wire _12065_;
wire _12066_;
wire _12067_;
wire _12068_;
wire _12069_;
wire _12070_;
wire _12071_;
wire _12072_;
wire _12073_;
wire _12074_;
wire _12075_;
wire _12076_;
wire _12077_;
wire _12078_;
wire _12079_;
wire _12080_;
wire _12081_;
wire _12082_;
wire _12083_;
wire _12084_;
wire _12085_;
wire _12086_;
wire _12087_;
wire _12088_;
wire _12089_;
wire _12090_;
wire _12091_;
wire _12092_;
wire _12093_;
wire _12094_;
wire _12095_;
wire _12096_;
wire _12097_;
wire _12098_;
wire _12099_;
wire _12100_;
wire _12101_;
wire _12102_;
wire _12103_;
wire _12104_;
wire _12105_;
wire _12106_;
wire _12107_;
wire _12108_;
wire _12109_;
wire _12110_;
wire _12111_;
wire _12112_;
wire _12113_;
wire _12114_;
wire _12115_;
wire _12116_;
wire _12117_;
wire _12118_;
wire _12119_;
wire _12120_;
wire _12121_;
wire _12122_;
wire _12123_;
wire _12124_;
wire _12125_;
wire _12126_;
wire _12127_;
wire _12128_;
wire _12129_;
wire _12130_;
wire _12131_;
wire _12132_;
wire _12133_;
wire _12134_;
wire _12135_;
wire _12136_;
wire _12137_;
wire _12138_;
wire _12139_;
wire _12140_;
wire _12141_;
wire _12142_;
wire _12143_;
wire _12144_;
wire _12145_;
wire _12146_;
wire _12147_;
wire _12148_;
wire _12149_;
wire _12150_;
wire _12151_;
wire _12152_;
wire _12153_;
wire _12154_;
wire _12155_;
wire _12156_;
wire _12157_;
wire _12158_;
wire _12159_;
wire _12160_;
wire _12161_;
wire _12162_;
wire _12163_;
wire _12164_;
wire _12165_;
wire _12166_;
wire _12167_;
wire _12168_;
wire _12169_;
wire _12170_;
wire _12171_;
wire _12172_;
wire _12173_;
wire _12174_;
wire _12175_;
wire _12176_;
wire _12177_;
wire _12178_;
wire _12179_;
wire _12180_;
wire _12181_;
wire _12182_;
wire _12183_;
wire _12184_;
wire _12185_;
wire _12186_;
wire _12187_;
wire _12188_;
wire _12189_;
wire _12190_;
wire _12191_;
wire _12192_;
wire _12193_;
wire _12194_;
wire _12195_;
wire _12196_;
wire _12197_;
wire _12198_;
wire _12199_;
wire _12200_;
wire _12201_;
wire _12202_;
wire _12203_;
wire _12204_;
wire _12205_;
wire _12206_;
wire _12207_;
wire _12208_;
wire _12209_;
wire _12210_;
wire _12211_;
wire _12212_;
wire _12213_;
wire _12214_;
wire _12215_;
wire _12216_;
wire _12217_;
wire _12218_;
wire _12219_;
wire _12220_;
wire _12221_;
wire _12222_;
wire _12223_;
wire _12224_;
wire _12225_;
wire _12226_;
wire _12227_;
wire _12228_;
wire _12229_;
wire _12230_;
wire _12231_;
wire _12232_;
wire _12233_;
wire _12234_;
wire _12235_;
wire _12236_;
wire _12237_;
wire _12238_;
wire _12239_;
wire _12240_;
wire _12241_;
wire _12242_;
wire _12243_;
wire _12244_;
wire _12245_;
wire _12246_;
wire _12247_;
wire _12248_;
wire _12249_;
wire _12250_;
wire _12251_;
wire _12252_;
wire _12253_;
wire _12254_;
wire _12255_;
wire _12256_;
wire _12257_;
wire _12258_;
wire _12259_;
wire _12260_;
wire _12261_;
wire _12262_;
wire _12263_;
wire _12264_;
wire _12265_;
wire _12266_;
wire _12267_;
wire _12268_;
wire _12269_;
wire _12270_;
wire _12271_;
wire _12272_;
wire _12273_;
wire _12274_;
wire _12275_;
wire _12276_;
wire _12277_;
wire _12278_;
wire _12279_;
wire _12280_;
wire _12281_;
wire _12282_;
wire _12283_;
wire _12284_;
wire _12285_;
wire _12286_;
wire _12287_;
wire _12288_;
wire _12289_;
wire _12290_;
wire _12291_;
wire _12292_;
wire _12293_;
wire _12294_;
wire _12295_;
wire _12296_;
wire _12297_;
wire _12298_;
wire _12299_;
wire _12300_;
wire _12301_;
wire _12302_;
wire _12303_;
wire _12304_;
wire _12305_;
wire _12306_;
wire _12307_;
wire _12308_;
wire _12309_;
wire _12310_;
wire _12311_;
wire _12312_;
wire _12313_;
wire _12314_;
wire _12315_;
wire _12316_;
wire _12317_;
wire _12318_;
wire _12319_;
wire _12320_;
wire _12321_;
wire _12322_;
wire _12323_;
wire _12324_;
wire _12325_;
wire _12326_;
wire _12327_;
wire _12328_;
wire _12329_;
wire _12330_;
wire _12331_;
wire _12332_;
wire _12333_;
wire _12334_;
wire _12335_;
wire _12336_;
wire _12337_;
wire _12338_;
wire _12339_;
wire _12340_;
wire _12341_;
wire _12342_;
wire _12343_;
wire _12344_;
wire _12345_;
wire _12346_;
wire _12347_;
wire _12348_;
wire _12349_;
wire _12350_;
wire _12351_;
wire _12352_;
wire _12353_;
wire _12354_;
wire _12355_;
wire _12356_;
wire _12357_;
wire _12358_;
wire _12359_;
wire _12360_;
wire _12361_;
wire _12362_;
wire _12363_;
wire _12364_;
wire _12365_;
wire _12366_;
wire _12367_;
wire _12368_;
wire _12369_;
wire _12370_;
wire _12371_;
wire _12372_;
wire _12373_;
wire _12374_;
wire _12375_;
wire _12376_;
wire _12377_;
wire _12378_;
wire _12379_;
wire _12380_;
wire _12381_;
wire _12382_;
wire _12383_;
wire _12384_;
wire _12385_;
wire _12386_;
wire _12387_;
wire _12388_;
wire _12389_;
wire _12390_;
wire _12391_;
wire _12392_;
wire _12393_;
wire _12394_;
wire _12395_;
wire _12396_;
wire _12397_;
wire _12398_;
wire _12399_;
wire _12400_;
wire _12401_;
wire _12402_;
wire _12403_;
wire _12404_;
wire _12405_;
wire _12406_;
wire _12407_;
wire _12408_;
wire _12409_;
wire _12410_;
wire _12411_;
wire _12412_;
wire _12413_;
wire _12414_;
wire _12415_;
wire _12416_;
wire _12417_;
wire _12418_;
wire _12419_;
wire _12420_;
wire _12421_;
wire _12422_;
wire _12423_;
wire _12424_;
wire _12425_;
wire _12426_;
wire _12427_;
wire _12428_;
wire _12429_;
wire _12430_;
wire _12431_;
wire _12432_;
wire _12433_;
wire _12434_;
wire _12435_;
wire _12436_;
wire _12437_;
wire _12438_;
wire _12439_;
wire _12440_;
wire _12441_;
wire _12442_;
wire _12443_;
wire _12444_;
wire _12445_;
wire _12446_;
wire _12447_;
wire _12448_;
wire _12449_;
wire _12450_;
wire _12451_;
wire _12452_;
wire _12453_;
wire _12454_;
wire _12455_;
wire _12456_;
wire _12457_;
wire _12458_;
wire _12459_;
wire _12460_;
wire _12461_;
wire _12462_;
wire _12463_;
wire _12464_;
wire _12465_;
wire _12466_;
wire _12467_;
wire _12468_;
wire _12469_;
wire _12470_;
wire _12471_;
wire _12472_;
wire _12473_;
wire _12474_;
wire _12475_;
wire _12476_;
wire _12477_;
wire _12478_;
wire _12479_;
wire _12480_;
wire _12481_;
wire _12482_;
wire _12483_;
wire _12484_;
wire _12485_;
wire _12486_;
wire _12487_;
wire _12488_;
wire _12489_;
wire _12490_;
wire _12491_;
wire _12492_;
wire _12493_;
wire _12494_;
wire _12495_;
wire _12496_;
wire _12497_;
wire _12498_;
wire _12499_;
wire _12500_;
wire _12501_;
wire _12502_;
wire _12503_;
wire _12504_;
wire _12505_;
wire _12506_;
wire _12507_;
wire _12508_;
wire _12509_;
wire _12510_;
wire _12511_;
wire _12512_;
wire _12513_;
wire _12514_;
wire _12515_;
wire _12516_;
wire _12517_;
wire _12518_;
wire _12519_;
wire _12520_;
wire _12521_;
wire _12522_;
wire _12523_;
wire _12524_;
wire _12525_;
wire _12526_;
wire _12527_;
wire _12528_;
wire _12529_;
wire _12530_;
wire _12531_;
wire _12532_;
wire _12533_;
wire _12534_;
wire _12535_;
wire _12536_;
wire _12537_;
wire _12538_;
wire _12539_;
wire _12540_;
wire _12541_;
wire _12542_;
wire _12543_;
wire _12544_;
wire _12545_;
wire _12546_;
wire _12547_;
wire _12548_;
wire _12549_;
wire _12550_;
wire _12551_;
wire _12552_;
wire _12553_;
wire _12554_;
wire _12555_;
wire _12556_;
wire _12557_;
wire _12558_;
wire _12559_;
wire _12560_;
wire _12561_;
wire _12562_;
wire _12563_;
wire _12564_;
wire _12565_;
wire _12566_;
wire _12567_;
wire _12568_;
wire _12569_;
wire _12570_;
wire _12571_;
wire _12572_;
wire _12573_;
wire _12574_;
wire _12575_;
wire _12576_;
wire _12577_;
wire _12578_;
wire _12579_;
wire _12580_;
wire _12581_;
wire _12582_;
wire _12583_;
wire _12584_;
wire _12585_;
wire _12586_;
wire _12587_;
wire _12588_;
wire _12589_;
wire _12590_;
wire _12591_;
wire _12592_;
wire _12593_;
wire _12594_;
wire _12595_;
wire _12596_;
wire _12597_;
wire _12598_;
wire _12599_;
wire _12600_;
wire _12601_;
wire _12602_;
wire _12603_;
wire _12604_;
wire _12605_;
wire _12606_;
wire _12607_;
wire _12608_;
wire _12609_;
wire _12610_;
wire _12611_;
wire _12612_;
wire _12613_;
wire _12614_;
wire _12615_;
wire _12616_;
wire _12617_;
wire _12618_;
wire _12619_;
wire _12620_;
wire _12621_;
wire _12622_;
wire _12623_;
wire _12624_;
wire _12625_;
wire _12626_;
wire _12627_;
wire _12628_;
wire _12629_;
wire _12630_;
wire _12631_;
wire _12632_;
wire _12633_;
wire _12634_;
wire _12635_;
wire _12636_;
wire _12637_;
wire _12638_;
wire _12639_;
wire _12640_;
wire _12641_;
wire _12642_;
wire _12643_;
wire _12644_;
wire _12645_;
wire _12646_;
wire _12647_;
wire _12648_;
wire _12649_;
wire _12650_;
wire _12651_;
wire _12652_;
wire _12653_;
wire _12654_;
wire _12655_;
wire _12656_;
wire _12657_;
wire _12658_;
wire _12659_;
wire _12660_;
wire _12661_;
wire _12662_;
wire _12663_;
wire _12664_;
wire _12665_;
wire _12666_;
wire _12667_;
wire _12668_;
wire _12669_;
wire _12670_;
wire _12671_;
wire _12672_;
wire _12673_;
wire _12674_;
wire _12675_;
wire _12676_;
wire _12677_;
wire _12678_;
wire _12679_;
wire _12680_;
wire _12681_;
wire _12682_;
wire _12683_;
wire _12684_;
wire _12685_;
wire _12686_;
wire _12687_;
wire _12688_;
wire _12689_;
wire _12690_;
wire _12691_;
wire _12692_;
wire _12693_;
wire _12694_;
wire _12695_;
wire _12696_;
wire _12697_;
wire _12698_;
wire _12699_;
wire _12700_;
wire _12701_;
wire _12702_;
wire _12703_;
wire _12704_;
wire _12705_;
wire _12706_;
wire _12707_;
wire _12708_;
wire _12709_;
wire _12710_;
wire _12711_;
wire _12712_;
wire _12713_;
wire _12714_;
wire _12715_;
wire _12716_;
wire _12717_;
wire _12718_;
wire _12719_;
wire _12720_;
wire _12721_;
wire _12722_;
wire _12723_;
wire _12724_;
wire _12725_;
wire _12726_;
wire _12727_;
wire _12728_;
wire _12729_;
wire _12730_;
wire _12731_;
wire _12732_;
wire _12733_;
wire _12734_;
wire _12735_;
wire _12736_;
wire _12737_;
wire _12738_;
wire _12739_;
wire _12740_;
wire _12741_;
wire _12742_;
wire _12743_;
wire _12744_;
wire _12745_;
wire _12746_;
wire _12747_;
wire _12748_;
wire _12749_;
wire _12750_;
wire _12751_;
wire _12752_;
wire _12753_;
wire _12754_;
wire _12755_;
wire _12756_;
wire _12757_;
wire _12758_;
wire _12759_;
wire _12760_;
wire _12761_;
wire _12762_;
wire _12763_;
wire _12764_;
wire _12765_;
wire _12766_;
wire _12767_;
wire _12768_;
wire _12769_;
wire _12770_;
wire _12771_;
wire _12772_;
wire _12773_;
wire _12774_;
wire _12775_;
wire _12776_;
wire _12777_;
wire _12778_;
wire _12779_;
wire _12780_;
wire _12781_;
wire _12782_;
wire _12783_;
wire _12784_;
wire _12785_;
wire _12786_;
wire _12787_;
wire _12788_;
wire _12789_;
wire _12790_;
wire _12791_;
wire _12792_;
wire _12793_;
wire _12794_;
wire _12795_;
wire _12796_;
wire _12797_;
wire _12798_;
wire _12799_;
wire _12800_;
wire _12801_;
wire _12802_;
wire _12803_;
wire _12804_;
wire _12805_;
wire _12806_;
wire _12807_;
wire _12808_;
wire _12809_;
wire _12810_;
wire _12811_;
wire _12812_;
wire _12813_;
wire _12814_;
wire _12815_;
wire _12816_;
wire _12817_;
wire _12818_;
wire _12819_;
wire _12820_;
wire _12821_;
wire _12822_;
wire _12823_;
wire _12824_;
wire _12825_;
wire _12826_;
wire _12827_;
wire _12828_;
wire _12829_;
wire _12830_;
wire _12831_;
wire _12832_;
wire _12833_;
wire _12834_;
wire _12835_;
wire _12836_;
wire _12837_;
wire _12838_;
wire _12839_;
wire _12840_;
wire _12841_;
wire _12842_;
wire _12843_;
wire _12844_;
wire _12845_;
wire _12846_;
wire _12847_;
wire _12848_;
wire _12849_;
wire _12850_;
wire _12851_;
wire _12852_;
wire _12853_;
wire _12854_;
wire _12855_;
wire _12856_;
wire _12857_;
wire _12858_;
wire _12859_;
wire _12860_;
wire _12861_;
wire _12862_;
wire _12863_;
wire _12864_;
wire _12865_;
wire _12866_;
wire _12867_;
wire _12868_;
wire _12869_;
wire _12870_;
wire _12871_;
wire _12872_;
wire _12873_;
wire _12874_;
wire _12875_;
wire _12876_;
wire _12877_;
wire _12878_;
wire _12879_;
wire _12880_;
wire _12881_;
wire _12882_;
wire _12883_;
wire _12884_;
wire _12885_;
wire _12886_;
wire _12887_;
wire _12888_;
wire _12889_;
wire _12890_;
wire _12891_;
wire _12892_;
wire _12893_;
wire _12894_;
wire _12895_;
wire _12896_;
wire _12897_;
wire _12898_;
wire _12899_;
wire _12900_;
wire _12901_;
wire _12902_;
wire _12903_;
wire _12904_;
wire _12905_;
wire _12906_;
wire _12907_;
wire _12908_;
wire _12909_;
wire _12910_;
wire _12911_;
wire _12912_;
wire _12913_;
wire _12914_;
wire _12915_;
wire _12916_;
wire _12917_;
wire _12918_;
wire _12919_;
wire _12920_;
wire _12921_;
wire _12922_;
wire _12923_;
wire _12924_;
wire _12925_;
wire _12926_;
wire _12927_;
wire _12928_;
wire _12929_;
wire _12930_;
wire _12931_;
wire _12932_;
wire _12933_;
wire _12934_;
wire _12935_;
wire _12936_;
wire _12937_;
wire _12938_;
wire _12939_;
wire _12940_;
wire _12941_;
wire _12942_;
wire _12943_;
wire _12944_;
wire _12945_;
wire _12946_;
wire _12947_;
wire _12948_;
wire _12949_;
wire _12950_;
wire _12951_;
wire _12952_;
wire _12953_;
wire _12954_;
wire _12955_;
wire _12956_;
wire _12957_;
wire _12958_;
wire _12959_;
wire _12960_;
wire _12961_;
wire _12962_;
wire _12963_;
wire _12964_;
wire _12965_;
wire _12966_;
wire _12967_;
wire _12968_;
wire _12969_;
wire _12970_;
wire _12971_;
wire _12972_;
wire _12973_;
wire _12974_;
wire _12975_;
wire _12976_;
wire _12977_;
wire _12978_;
wire _12979_;
wire _12980_;
wire _12981_;
wire _12982_;
wire _12983_;
wire _12984_;
wire _12985_;
wire _12986_;
wire _12987_;
wire _12988_;
wire _12989_;
wire _12990_;
wire _12991_;
wire _12992_;
wire _12993_;
wire _12994_;
wire _12995_;
wire _12996_;
wire _12997_;
wire _12998_;
wire _12999_;
wire _13000_;
wire _13001_;
wire _13002_;
wire _13003_;
wire _13004_;
wire _13005_;
wire _13006_;
wire _13007_;
wire _13008_;
wire _13009_;
wire _13010_;
wire _13011_;
wire _13012_;
wire _13013_;
wire _13014_;
wire _13015_;
wire _13016_;
wire _13017_;
wire _13018_;
wire _13019_;
wire _13020_;
wire _13021_;
wire _13022_;
wire _13023_;
wire _13024_;
wire _13025_;
wire _13026_;
wire _13027_;
wire _13028_;
wire _13029_;
wire _13030_;
wire _13031_;
wire _13032_;
wire _13033_;
wire _13034_;
wire _13035_;
wire _13036_;
wire _13037_;
wire _13038_;
wire _13039_;
wire _13040_;
wire _13041_;
wire _13042_;
wire _13043_;
wire _13044_;
wire _13045_;
wire _13046_;
wire _13047_;
wire _13048_;
wire _13049_;
wire _13050_;
wire _13051_;
wire _13052_;
wire _13053_;
wire _13054_;
wire _13055_;
wire _13056_;
wire _13057_;
wire _13058_;
wire _13059_;
wire _13060_;
wire _13061_;
wire _13062_;
wire _13063_;
wire _13064_;
wire _13065_;
wire _13066_;
wire _13067_;
wire _13068_;
wire _13069_;
wire _13070_;
wire _13071_;
wire _13072_;
wire _13073_;
wire _13074_;
wire _13075_;
wire _13076_;
wire _13077_;
wire _13078_;
wire _13079_;
wire _13080_;
wire _13081_;
wire _13082_;
wire _13083_;
wire _13084_;
wire _13085_;
wire _13086_;
wire _13087_;
wire _13088_;
wire _13089_;
wire _13090_;
wire _13091_;
wire _13092_;
wire _13093_;
wire _13094_;
wire _13095_;
wire _13096_;
wire _13097_;
wire _13098_;
wire _13099_;
wire _13100_;
wire _13101_;
wire _13102_;
wire _13103_;
wire _13104_;
wire _13105_;
wire _13106_;
wire _13107_;
wire _13108_;
wire _13109_;
wire _13110_;
wire _13111_;
wire _13112_;
wire _13113_;
wire _13114_;
wire _13115_;
wire _13116_;
wire _13117_;
wire _13118_;
wire _13119_;
wire _13120_;
wire _13121_;
wire _13122_;
wire _13123_;
wire _13124_;
wire _13125_;
wire _13126_;
wire _13127_;
wire _13128_;
wire _13129_;
wire _13130_;
wire _13131_;
wire _13132_;
wire _13133_;
wire _13134_;
wire _13135_;
wire _13136_;
wire _13137_;
wire _13138_;
wire _13139_;
wire _13140_;
wire _13141_;
wire _13142_;
wire _13143_;
wire _13144_;
wire _13145_;
wire _13146_;
wire _13147_;
wire _13148_;
wire _13149_;
wire _13150_;
wire _13151_;
wire _13152_;
wire _13153_;
wire _13154_;
wire _13155_;
wire _13156_;
wire _13157_;
wire _13158_;
wire _13159_;
wire _13160_;
wire _13161_;
wire _13162_;
wire _13163_;
wire _13164_;
wire _13165_;
wire _13166_;
wire _13167_;
wire _13168_;
wire _13169_;
wire _13170_;
wire _13171_;
wire _13172_;
wire _13173_;
wire _13174_;
wire _13175_;
wire _13176_;
wire _13177_;
wire _13178_;
wire _13179_;
wire _13180_;
wire _13181_;
wire _13182_;
wire _13183_;
wire _13184_;
wire _13185_;
wire _13186_;
wire _13187_;
wire _13188_;
wire _13189_;
wire _13190_;
wire _13191_;
wire _13192_;
wire _13193_;
wire _13194_;
wire _13195_;
wire _13196_;
wire _13197_;
wire _13198_;
wire _13199_;
wire _13200_;
wire _13201_;
wire _13202_;
wire _13203_;
wire _13204_;
wire _13205_;
wire _13206_;
wire _13207_;
wire _13208_;
wire _13209_;
wire _13210_;
wire _13211_;
wire _13212_;
wire _13213_;
wire _13214_;
wire _13215_;
wire _13216_;
wire _13217_;
wire _13218_;
wire _13219_;
wire _13220_;
wire _13221_;
wire _13222_;
wire _13223_;
wire _13224_;
wire _13225_;
wire _13226_;
wire _13227_;
wire _13228_;
wire _13229_;
wire _13230_;
wire _13231_;
wire _13232_;
wire _13233_;
wire _13234_;
wire _13235_;
wire _13236_;
wire _13237_;
wire _13238_;
wire _13239_;
wire _13240_;
wire _13241_;
wire _13242_;
wire _13243_;
wire _13244_;
wire _13245_;
wire _13246_;
wire _13247_;
wire _13248_;
wire _13249_;
wire _13250_;
wire _13251_;
wire _13252_;
wire _13253_;
wire _13254_;
wire _13255_;
wire _13256_;
wire _13257_;
wire _13258_;
wire _13259_;
wire _13260_;
wire _13261_;
wire _13262_;
wire _13263_;
wire _13264_;
wire _13265_;
wire _13266_;
wire _13267_;
wire _13268_;
wire _13269_;
wire _13270_;
wire _13271_;
wire _13272_;
wire _13273_;
wire _13274_;
wire _13275_;
wire _13276_;
wire _13277_;
wire _13278_;
wire _13279_;
wire _13280_;
wire _13281_;
wire _13282_;
wire _13283_;
wire _13284_;
wire _13285_;
wire _13286_;
wire _13287_;
wire _13288_;
wire _13289_;
wire _13290_;
wire _13291_;
wire _13292_;
wire _13293_;
wire _13294_;
wire _13295_;
wire _13296_;
wire _13297_;
wire _13298_;
wire _13299_;
wire _13300_;
wire _13301_;
wire _13302_;
wire _13303_;
wire _13304_;
wire _13305_;
wire _13306_;
wire _13307_;
wire _13308_;
wire _13309_;
wire _13310_;
wire _13311_;
wire _13312_;
wire _13313_;
wire _13314_;
wire _13315_;
wire _13316_;
wire _13317_;
wire _13318_;
wire _13319_;
wire _13320_;
wire _13321_;
wire _13322_;
wire _13323_;
wire _13324_;
wire _13325_;
wire _13326_;
wire _13327_;
wire _13328_;
wire _13329_;
wire _13330_;
wire _13331_;
wire _13332_;
wire _13333_;
wire _13334_;
wire _13335_;
wire _13336_;
wire _13337_;
wire _13338_;
wire _13339_;
wire _13340_;
wire _13341_;
wire _13342_;
wire _13343_;
wire _13344_;
wire _13345_;
wire _13346_;
wire _13347_;
wire _13348_;
wire _13349_;
wire _13350_;
wire _13351_;
wire _13352_;
wire _13353_;
wire _13354_;
wire _13355_;
wire _13356_;
wire _13357_;
wire _13358_;
wire _13359_;
wire _13360_;
wire _13361_;
wire _13362_;
wire _13363_;
wire _13364_;
wire _13365_;
wire _13366_;
wire _13367_;
wire _13368_;
wire _13369_;
wire _13370_;
wire _13371_;
wire _13372_;
wire _13373_;
wire _13374_;
wire _13375_;
wire _13376_;
wire _13377_;
wire _13378_;
wire _13379_;
wire _13380_;
wire _13381_;
wire _13382_;
wire _13383_;
wire _13384_;
wire _13385_;
wire _13386_;
wire _13387_;
wire _13388_;
wire _13389_;
wire _13390_;
wire _13391_;
wire _13392_;
wire _13393_;
wire _13394_;
wire _13395_;
wire _13396_;
wire _13397_;
wire _13398_;
wire _13399_;
wire _13400_;
wire _13401_;
wire _13402_;
wire _13403_;
wire _13404_;
wire _13405_;
wire _13406_;
wire _13407_;
wire _13408_;
wire _13409_;
wire _13410_;
wire _13411_;
wire _13412_;
wire _13413_;
wire _13414_;
wire _13415_;
wire _13416_;
wire _13417_;
wire _13418_;
wire _13419_;
wire _13420_;
wire _13421_;
wire _13422_;
wire _13423_;
wire _13424_;
wire _13425_;
wire _13426_;
wire _13427_;
wire _13428_;
wire _13429_;
wire _13430_;
wire _13431_;
wire _13432_;
wire _13433_;
wire _13434_;
wire _13435_;
wire _13436_;
wire _13437_;
wire _13438_;
wire _13439_;
wire _13440_;
wire _13441_;
wire _13442_;
wire _13443_;
wire _13444_;
wire _13445_;
wire _13446_;
wire _13447_;
wire _13448_;
wire _13449_;
wire _13450_;
wire _13451_;
wire _13452_;
wire _13453_;
wire _13454_;
wire _13455_;
wire _13456_;
wire _13457_;
wire _13458_;
wire _13459_;
wire _13460_;
wire _13461_;
wire _13462_;
wire _13463_;
wire _13464_;
wire _13465_;
wire _13466_;
wire _13467_;
wire _13468_;
wire _13469_;
wire _13470_;
wire _13471_;
wire _13472_;
wire _13473_;
wire _13474_;
wire _13475_;
wire _13476_;
wire _13477_;
wire _13478_;
wire _13479_;
wire _13480_;
wire _13481_;
wire _13482_;
wire _13483_;
wire _13484_;
wire _13485_;
wire _13486_;
wire _13487_;
wire _13488_;
wire _13489_;
wire _13490_;
wire _13491_;
wire _13492_;
wire _13493_;
wire _13494_;
wire _13495_;
wire _13496_;
wire _13497_;
wire _13498_;
wire _13499_;
wire _13500_;
wire _13501_;
wire _13502_;
wire _13503_;
wire _13504_;
wire _13505_;
wire _13506_;
wire _13507_;
wire _13508_;
wire _13509_;
wire _13510_;
wire _13511_;
wire _13512_;
wire _13513_;
wire _13514_;
wire _13515_;
wire _13516_;
wire _13517_;
wire _13518_;
wire _13519_;
wire _13520_;
wire _13521_;
wire _13522_;
wire _13523_;
wire _13524_;
wire _13525_;
wire _13526_;
wire _13527_;
wire _13528_;
wire _13529_;
wire _13530_;
wire _13531_;
wire _13532_;
wire _13533_;
wire _13534_;
wire _13535_;
wire _13536_;
wire _13537_;
wire _13538_;
wire _13539_;
wire _13540_;
wire _13541_;
wire _13542_;
wire _13543_;
wire _13544_;
wire _13545_;
wire _13546_;
wire _13547_;
wire _13548_;
wire _13549_;
wire _13550_;
wire _13551_;
wire _13552_;
wire _13553_;
wire _13554_;
wire _13555_;
wire _13556_;
wire _13557_;
wire _13558_;
wire _13559_;
wire _13560_;
wire _13561_;
wire _13562_;
wire _13563_;
wire _13564_;
wire _13565_;
wire _13566_;
wire _13567_;
wire _13568_;
wire _13569_;
wire _13570_;
wire _13571_;
wire _13572_;
wire _13573_;
wire _13574_;
wire _13575_;
wire _13576_;
wire _13577_;
wire _13578_;
wire _13579_;
wire _13580_;
wire _13581_;
wire _13582_;
wire _13583_;
wire _13584_;
wire _13585_;
wire _13586_;
wire _13587_;
wire _13588_;
wire _13589_;
wire _13590_;
wire _13591_;
wire _13592_;
wire _13593_;
wire _13594_;
wire _13595_;
wire _13596_;
wire _13597_;
wire _13598_;
wire _13599_;
wire _13600_;
wire _13601_;
wire _13602_;
wire _13603_;
wire _13604_;
wire _13605_;
wire _13606_;
wire _13607_;
wire _13608_;
wire _13609_;
wire _13610_;
wire _13611_;
wire _13612_;
wire _13613_;
wire _13614_;
wire _13615_;
wire _13616_;
wire _13617_;
wire _13618_;
wire _13619_;
wire _13620_;
wire _13621_;
wire _13622_;
wire _13623_;
wire _13624_;
wire _13625_;
wire _13626_;
wire _13627_;
wire _13628_;
wire _13629_;
wire _13630_;
wire _13631_;
wire _13632_;
wire _13633_;
wire _13634_;
wire _13635_;
wire _13636_;
wire _13637_;
wire _13638_;
wire _13639_;
wire _13640_;
wire _13641_;
wire _13642_;
wire _13643_;
wire _13644_;
wire _13645_;
wire _13646_;
wire _13647_;
wire _13648_;
wire _13649_;
wire _13650_;
wire _13651_;
wire _13652_;
wire _13653_;
wire _13654_;
wire _13655_;
wire _13656_;
wire _13657_;
wire _13658_;
wire _13659_;
wire _13660_;
wire _13661_;
wire _13662_;
wire _13663_;
wire _13664_;
wire _13665_;
wire _13666_;
wire _13667_;
wire _13668_;
wire _13669_;
wire _13670_;
wire _13671_;
wire _13672_;
wire _13673_;
wire _13674_;
wire _13675_;
wire _13676_;
wire _13677_;
wire _13678_;
wire _13679_;
wire _13680_;
wire _13681_;
wire _13682_;
wire _13683_;
wire _13684_;
wire _13685_;
wire _13686_;
wire _13687_;
wire _13688_;
wire _13689_;
wire _13690_;
wire _13691_;
wire _13692_;
wire _13693_;
wire _13694_;
wire _13695_;
wire _13696_;
wire _13697_;
wire _13698_;
wire _13699_;
wire _13700_;
wire _13701_;
wire _13702_;
wire _13703_;
wire _13704_;
wire _13705_;
wire _13706_;
wire _13707_;
wire _13708_;
wire _13709_;
wire _13710_;
wire _13711_;
wire _13712_;
wire _13713_;
wire _13714_;
wire _13715_;
wire _13716_;
wire _13717_;
wire _13718_;
wire _13719_;
wire _13720_;
wire _13721_;
wire _13722_;
wire _13723_;
wire _13724_;
wire _13725_;
wire _13726_;
wire _13727_;
wire _13728_;
wire _13729_;
wire _13730_;
wire _13731_;
wire _13732_;
wire _13733_;
wire _13734_;
wire _13735_;
wire _13736_;
wire _13737_;
wire _13738_;
wire _13739_;
wire _13740_;
wire _13741_;
wire _13742_;
wire _13743_;
wire _13744_;
wire _13745_;
wire _13746_;
wire _13747_;
wire _13748_;
wire _13749_;
wire _13750_;
wire _13751_;
wire _13752_;
wire _13753_;
wire _13754_;
wire _13755_;
wire _13756_;
wire _13757_;
wire _13758_;
wire _13759_;
wire _13760_;
wire _13761_;
wire _13762_;
wire _13763_;
wire _13764_;
wire _13765_;
wire _13766_;
wire _13767_;
wire _13768_;
wire _13769_;
wire _13770_;
wire _13771_;
wire _13772_;
wire _13773_;
wire _13774_;
wire _13775_;
wire _13776_;
wire _13777_;
wire _13778_;
wire _13779_;
wire _13780_;
wire _13781_;
wire _13782_;
wire _13783_;
wire _13784_;
wire _13785_;
wire _13786_;
wire _13787_;
wire _13788_;
wire _13789_;
wire _13790_;
wire _13791_;
wire _13792_;
wire _13793_;
wire _13794_;
wire _13795_;
wire _13796_;
wire _13797_;
wire _13798_;
wire _13799_;
wire _13800_;
wire _13801_;
wire _13802_;
wire _13803_;
wire _13804_;
wire _13805_;
wire _13806_;
wire _13807_;
wire _13808_;
wire _13809_;
wire _13810_;
wire _13811_;
wire _13812_;
wire _13813_;
wire _13814_;
wire _13815_;
wire _13816_;
wire _13817_;
wire _13818_;
wire _13819_;
wire _13820_;
wire _13821_;
wire _13822_;
wire _13823_;
wire _13824_;
wire _13825_;
wire _13826_;
wire _13827_;
wire _13828_;
wire _13829_;
wire _13830_;
wire _13831_;
wire _13832_;
wire _13833_;
wire _13834_;
wire _13835_;
wire _13836_;
wire _13837_;
wire _13838_;
wire _13839_;
wire _13840_;
wire _13841_;
wire _13842_;
wire _13843_;
wire _13844_;
wire _13845_;
wire _13846_;
wire _13847_;
wire _13848_;
wire _13849_;
wire _13850_;
wire _13851_;
wire _13852_;
wire _13853_;
wire _13854_;
wire _13855_;
wire _13856_;
wire _13857_;
wire _13858_;
wire _13859_;
wire _13860_;
wire _13861_;
wire _13862_;
wire _13863_;
wire _13864_;
wire _13865_;
wire _13866_;
wire _13867_;
wire _13868_;
wire _13869_;
wire _13870_;
wire _13871_;
wire _13872_;
wire _13873_;
wire _13874_;
wire _13875_;
wire _13876_;
wire _13877_;
wire _13878_;
wire _13879_;
wire _13880_;
wire _13881_;
wire _13882_;
wire _13883_;
wire _13884_;
wire _13885_;
wire _13886_;
wire _13887_;
wire _13888_;
wire _13889_;
wire _13890_;
wire _13891_;
wire _13892_;
wire _13893_;
wire _13894_;
wire _13895_;
wire _13896_;
wire _13897_;
wire _13898_;
wire _13899_;
wire _13900_;
wire _13901_;
wire _13902_;
wire _13903_;
wire _13904_;
wire _13905_;
wire _13906_;
wire _13907_;
wire _13908_;
wire _13909_;
wire _13910_;
wire _13911_;
wire _13912_;
wire _13913_;
wire _13914_;
wire _13915_;
wire _13916_;
wire _13917_;
wire _13918_;
wire _13919_;
wire _13920_;
wire _13921_;
wire _13922_;
wire _13923_;
wire _13924_;
wire _13925_;
wire _13926_;
wire _13927_;
wire _13928_;
wire _13929_;
wire _13930_;
wire _13931_;
wire _13932_;
wire _13933_;
wire _13934_;
wire _13935_;
wire _13936_;
wire _13937_;
wire _13938_;
wire _13939_;
wire _13940_;
wire _13941_;
wire _13942_;
wire _13943_;
wire _13944_;
wire _13945_;
wire _13946_;
wire _13947_;
wire _13948_;
wire _13949_;
wire _13950_;
wire _13951_;
wire _13952_;
wire _13953_;
wire _13954_;
wire _13955_;
wire _13956_;
wire _13957_;
wire _13958_;
wire _13959_;
wire _13960_;
wire _13961_;
wire _13962_;
wire _13963_;
wire _13964_;
wire _13965_;
wire _13966_;
wire _13967_;
wire _13968_;
wire _13969_;
wire _13970_;
wire _13971_;
wire _13972_;
wire _13973_;
wire _13974_;
wire _13975_;
wire _13976_;
wire _13977_;
wire _13978_;
wire _13979_;
wire _13980_;
wire _13981_;
wire _13982_;
wire _13983_;
wire _13984_;
wire _13985_;
wire _13986_;
wire _13987_;
wire _13988_;
wire _13989_;
wire _13990_;
wire _13991_;
wire _13992_;
wire _13993_;
wire _13994_;
wire _13995_;
wire _13996_;
wire _13997_;
wire _13998_;
wire _13999_;
wire _14000_;
wire _14001_;
wire _14002_;
wire _14003_;
wire _14004_;
wire _14005_;
wire _14006_;
wire _14007_;
wire _14008_;
wire _14009_;
wire _14010_;
wire _14011_;
wire _14012_;
wire _14013_;
wire _14014_;
wire _14015_;
wire _14016_;
wire _14017_;
wire _14018_;
wire _14019_;
wire _14020_;
wire _14021_;
wire _14022_;
wire _14023_;
wire _14024_;
wire _14025_;
wire _14026_;
wire _14027_;
wire _14028_;
wire _14029_;
wire _14030_;
wire _14031_;
wire _14032_;
wire _14033_;
wire _14034_;
wire _14035_;
wire _14036_;
wire _14037_;
wire _14038_;
wire _14039_;
wire _14040_;
wire _14041_;
wire _14042_;
wire _14043_;
wire _14044_;
wire _14045_;
wire _14046_;
wire _14047_;
wire _14048_;
wire _14049_;
wire _14050_;
wire _14051_;
wire _14052_;
wire _14053_;
wire _14054_;
wire _14055_;
wire _14056_;
wire _14057_;
wire _14058_;
wire _14059_;
wire _14060_;
wire _14061_;
wire _14062_;
wire _14063_;
wire _14064_;
wire _14065_;
wire _14066_;
wire _14067_;
wire _14068_;
wire _14069_;
wire _14070_;
wire _14071_;
wire _14072_;
wire _14073_;
wire _14074_;
wire _14075_;
wire _14076_;
wire _14077_;
wire _14078_;
wire _14079_;
wire _14080_;
wire _14081_;
wire _14082_;
wire _14083_;
wire _14084_;
wire _14085_;
wire _14086_;
wire _14087_;
wire _14088_;
wire _14089_;
wire _14090_;
wire _14091_;
wire _14092_;
wire _14093_;
wire _14094_;
wire _14095_;
wire _14096_;
wire _14097_;
wire _14098_;
wire _14099_;
wire _14100_;
wire _14101_;
wire _14102_;
wire _14103_;
wire _14104_;
wire _14105_;
wire _14106_;
wire _14107_;
wire _14108_;
wire _14109_;
wire _14110_;
wire _14111_;
wire _14112_;
wire _14113_;
wire _14114_;
wire _14115_;
wire _14116_;
wire _14117_;
wire _14118_;
wire _14119_;
wire _14120_;
wire _14121_;
wire _14122_;
wire _14123_;
wire _14124_;
wire _14125_;
wire _14126_;
wire _14127_;
wire _14128_;
wire _14129_;
wire _14130_;
wire _14131_;
wire _14132_;
wire _14133_;
wire _14134_;
wire _14135_;
wire _14136_;
wire _14137_;
wire _14138_;
wire _14139_;
wire _14140_;
wire _14141_;
wire _14142_;
wire _14143_;
wire _14144_;
wire _14145_;
wire _14146_;
wire _14147_;
wire _14148_;
wire _14149_;
wire _14150_;
wire _14151_;
wire _14152_;
wire _14153_;
wire _14154_;
wire _14155_;
wire _14156_;
wire _14157_;
wire _14158_;
wire _14159_;
wire _14160_;
wire _14161_;
wire _14162_;
wire _14163_;
wire _14164_;
wire _14165_;
wire _14166_;
wire _14167_;
wire _14168_;
wire _14169_;
wire _14170_;
wire _14171_;
wire _14172_;
wire _14173_;
wire _14174_;
wire _14175_;
wire _14176_;
wire _14177_;
wire _14178_;
wire _14179_;
wire _14180_;
wire _14181_;
wire _14182_;
wire _14183_;
wire _14184_;
wire _14185_;
wire _14186_;
wire _14187_;
wire _14188_;
wire _14189_;
wire _14190_;
wire _14191_;
wire _14192_;
wire _14193_;
wire _14194_;
wire _14195_;
wire _14196_;
wire _14197_;
wire _14198_;
wire _14199_;
wire _14200_;
wire _14201_;
wire _14202_;
wire _14203_;
wire _14204_;
wire _14205_;
wire _14206_;
wire _14207_;
wire _14208_;
wire _14209_;
wire _14210_;
wire _14211_;
wire _14212_;
wire _14213_;
wire _14214_;
wire _14215_;
wire _14216_;
wire _14217_;
wire _14218_;
wire _14219_;
wire _14220_;
wire _14221_;
wire _14222_;
wire _14223_;
wire _14224_;
wire _14225_;
wire _14226_;
wire _14227_;
wire _14228_;
wire _14229_;
wire _14230_;
wire _14231_;
wire _14232_;
wire _14233_;
wire _14234_;
wire _14235_;
wire _14236_;
wire _14237_;
wire _14238_;
wire _14239_;
wire _14240_;
wire _14241_;
wire _14242_;
wire _14243_;
wire _14244_;
wire _14245_;
wire _14246_;
wire _14247_;
wire _14248_;
wire _14249_;
wire _14250_;
wire _14251_;
wire _14252_;
wire _14253_;
wire _14254_;
wire _14255_;
wire _14256_;
wire _14257_;
wire _14258_;
wire _14259_;
wire _14260_;
wire _14261_;
wire _14262_;
wire _14263_;
wire _14264_;
wire _14265_;
wire _14266_;
wire _14267_;
wire _14268_;
wire _14269_;
wire _14270_;
wire _14271_;
wire _14272_;
wire _14273_;
wire _14274_;
wire _14275_;
wire _14276_;
wire _14277_;
wire _14278_;
wire _14279_;
wire _14280_;
wire _14281_;
wire _14282_;
wire _14283_;
wire _14284_;
wire _14285_;
wire _14286_;
wire _14287_;
wire _14288_;
wire _14289_;
wire _14290_;
wire _14291_;
wire _14292_;
wire _14293_;
wire _14294_;
wire _14295_;
wire _14296_;
wire _14297_;
wire _14298_;
wire _14299_;
wire _14300_;
wire _14301_;
wire _14302_;
wire _14303_;
wire _14304_;
wire _14305_;
wire _14306_;
wire _14307_;
wire _14308_;
wire _14309_;
wire _14310_;
wire _14311_;
wire _14312_;
wire _14313_;
wire _14314_;
wire _14315_;
wire _14316_;
wire _14317_;
wire _14318_;
wire _14319_;
wire _14320_;
wire _14321_;
wire _14322_;
wire _14323_;
wire _14324_;
wire _14325_;
wire _14326_;
wire _14327_;
wire _14328_;
wire _14329_;
wire _14330_;
wire _14331_;
wire _14332_;
wire _14333_;
wire _14334_;
wire _14335_;
wire _14336_;
wire _14337_;
wire _14338_;
wire _14339_;
wire _14340_;
wire _14341_;
wire _14342_;
wire _14343_;
wire _14344_;
wire _14345_;
wire _14346_;
wire _14347_;
wire _14348_;
wire _14349_;
wire _14350_;
wire _14351_;
wire _14352_;
wire _14353_;
wire _14354_;
wire _14355_;
wire _14356_;
wire _14357_;
wire _14358_;
wire _14359_;
wire _14360_;
wire _14361_;
wire _14362_;
wire _14363_;
wire _14364_;
wire _14365_;
wire _14366_;
wire _14367_;
wire _14368_;
wire _14369_;
wire _14370_;
wire _14371_;
wire _14372_;
wire _14373_;
wire _14374_;
wire _14375_;
wire _14376_;
wire _14377_;
wire _14378_;
wire _14379_;
wire _14380_;
wire _14381_;
wire _14382_;
wire _14383_;
wire _14384_;
wire _14385_;
wire _14386_;
wire _14387_;
wire _14388_;
wire _14389_;
wire _14390_;
wire _14391_;
wire _14392_;
wire _14393_;
wire _14394_;
wire _14395_;
wire _14396_;
wire _14397_;
wire _14398_;
wire _14399_;
wire _14400_;
wire _14401_;
wire _14402_;
wire _14403_;
wire _14404_;
wire _14405_;
wire _14406_;
wire _14407_;
wire _14408_;
wire _14409_;
wire _14410_;
wire _14411_;
wire _14412_;
wire _14413_;
wire _14414_;
wire _14415_;
wire _14416_;
wire _14417_;
wire _14418_;
wire _14419_;
wire _14420_;
wire _14421_;
wire _14422_;
wire _14423_;
wire _14424_;
wire _14425_;
wire _14426_;
wire _14427_;
wire _14428_;
wire _14429_;
wire _14430_;
wire _14431_;
wire _14432_;
wire _14433_;
wire _14434_;
wire _14435_;
wire _14436_;
wire _14437_;
wire _14438_;
wire _14439_;
wire _14440_;
wire _14441_;
wire _14442_;
wire _14443_;
wire _14444_;
wire _14445_;
wire _14446_;
wire _14447_;
wire _14448_;
wire _14449_;
wire _14450_;
wire _14451_;
wire _14452_;
wire _14453_;
wire _14454_;
wire _14455_;
wire _14456_;
wire _14457_;
wire _14458_;
wire _14459_;
wire _14460_;
wire _14461_;
wire _14462_;
wire _14463_;
wire _14464_;
wire _14465_;
wire _14466_;
wire _14467_;
wire _14468_;
wire _14469_;
wire _14470_;
wire _14471_;
wire _14472_;
wire _14473_;
wire _14474_;
wire _14475_;
wire _14476_;
wire _14477_;
wire _14478_;
wire _14479_;
wire _14480_;
wire _14481_;
wire _14482_;
wire _14483_;
wire _14484_;
wire _14485_;
wire _14486_;
wire _14487_;
wire _14488_;
wire _14489_;
wire _14490_;
wire _14491_;
wire _14492_;
wire _14493_;
wire _14494_;
wire _14495_;
wire _14496_;
wire _14497_;
wire _14498_;
wire _14499_;
wire _14500_;
wire _14501_;
wire _14502_;
wire _14503_;
wire _14504_;
wire _14505_;
wire _14506_;
wire _14507_;
wire _14508_;
wire _14509_;
wire _14510_;
wire _14511_;
wire _14512_;
wire _14513_;
wire _14514_;
wire _14515_;
wire _14516_;
wire _14517_;
wire _14518_;
wire _14519_;
wire _14520_;
wire _14521_;
wire _14522_;
wire _14523_;
wire _14524_;
wire _14525_;
wire _14526_;
wire _14527_;
wire _14528_;
wire _14529_;
wire _14530_;
wire _14531_;
wire _14532_;
wire _14533_;
wire _14534_;
wire _14535_;
wire _14536_;
wire _14537_;
wire _14538_;
wire _14539_;
wire _14540_;
wire _14541_;
wire _14542_;
wire _14543_;
wire _14544_;
wire _14545_;
wire _14546_;
wire _14547_;
wire _14548_;
wire _14549_;
wire _14550_;
wire _14551_;
wire _14552_;
wire _14553_;
wire _14554_;
wire _14555_;
wire _14556_;
wire _14557_;
wire _14558_;
wire _14559_;
wire _14560_;
wire _14561_;
wire _14562_;
wire _14563_;
wire _14564_;
wire _14565_;
wire _14566_;
wire _14567_;
wire _14568_;
wire _14569_;
wire _14570_;
wire _14571_;
wire _14572_;
wire _14573_;
wire _14574_;
wire _14575_;
wire _14576_;
wire _14577_;
wire _14578_;
wire _14579_;
wire _14580_;
wire _14581_;
wire _14582_;
wire _14583_;
wire _14584_;
wire _14585_;
wire _14586_;
wire _14587_;
wire _14588_;
wire _14589_;
wire _14590_;
wire _14591_;
wire _14592_;
wire _14593_;
wire _14594_;
wire _14595_;
wire _14596_;
wire _14597_;
wire _14598_;
wire _14599_;
wire _14600_;
wire _14601_;
wire _14602_;
wire _14603_;
wire _14604_;
wire _14605_;
wire _14606_;
wire _14607_;
wire _14608_;
wire _14609_;
wire _14610_;
wire _14611_;
wire _14612_;
wire _14613_;
wire _14614_;
wire _14615_;
wire _14616_;
wire _14617_;
wire _14618_;
wire _14619_;
wire _14620_;
wire _14621_;
wire _14622_;
wire _14623_;
wire _14624_;
wire _14625_;
wire _14626_;
wire _14627_;
wire _14628_;
wire _14629_;
wire _14630_;
wire _14631_;
wire _14632_;
wire _14633_;
wire _14634_;
wire _14635_;
wire _14636_;
wire _14637_;
wire _14638_;
wire _14639_;
wire _14640_;
wire _14641_;
wire _14642_;
wire _14643_;
wire _14644_;
wire _14645_;
wire _14646_;
wire _14647_;
wire _14648_;
wire _14649_;
wire _14650_;
wire _14651_;
wire _14652_;
wire _14653_;
wire _14654_;
wire _14655_;
wire _14656_;
wire _14657_;
wire _14658_;
wire _14659_;
wire _14660_;
wire _14661_;
wire _14662_;
wire _14663_;
wire _14664_;
wire _14665_;
wire _14666_;
wire _14667_;
wire _14668_;
wire _14669_;
wire _14670_;
wire _14671_;
wire _14672_;
wire _14673_;
wire _14674_;
wire _14675_;
wire _14676_;
wire _14677_;
wire _14678_;
wire _14679_;
wire _14680_;
wire _14681_;
wire _14682_;
wire _14683_;
wire _14684_;
wire _14685_;
wire _14686_;
wire _14687_;
wire _14688_;
wire _14689_;
wire _14690_;
wire _14691_;
wire _14692_;
wire _14693_;
wire _14694_;
wire _14695_;
wire _14696_;
wire _14697_;
wire _14698_;
wire _14699_;
wire _14700_;
wire _14701_;
wire _14702_;
wire _14703_;
wire _14704_;
wire _14705_;
wire _14706_;
wire _14707_;
wire _14708_;
wire _14709_;
wire _14710_;
wire _14711_;
wire _14712_;
wire _14713_;
wire _14714_;
wire _14715_;
wire _14716_;
wire _14717_;
wire _14718_;
wire _14719_;
wire _14720_;
wire _14721_;
wire _14722_;
wire _14723_;
wire _14724_;
wire _14725_;
wire _14726_;
wire _14727_;
wire _14728_;
wire _14729_;
wire _14730_;
wire _14731_;
wire _14732_;
wire _14733_;
wire _14734_;
wire _14735_;
wire _14736_;
wire _14737_;
wire _14738_;
wire _14739_;
wire _14740_;
wire _14741_;
wire _14742_;
wire _14743_;
wire _14744_;
wire _14745_;
wire _14746_;
wire _14747_;
wire _14748_;
wire _14749_;
wire _14750_;
wire _14751_;
wire _14752_;
wire _14753_;
wire _14754_;
wire _14755_;
wire _14756_;
wire _14757_;
wire _14758_;
wire _14759_;
wire _14760_;
wire _14761_;
wire _14762_;
wire _14763_;
wire _14764_;
wire _14765_;
wire _14766_;
wire _14767_;
wire _14768_;
wire _14769_;
wire _14770_;
wire _14771_;
wire _14772_;
wire _14773_;
wire _14774_;
wire _14775_;
wire _14776_;
wire _14777_;
wire _14778_;
wire _14779_;
wire _14780_;
wire _14781_;
wire _14782_;
wire _14783_;
wire _14784_;
wire _14785_;
wire _14786_;
wire _14787_;
wire _14788_;
wire _14789_;
wire _14790_;
wire _14791_;
wire _14792_;
wire _14793_;
wire _14794_;
wire _14795_;
wire _14796_;
wire _14797_;
wire _14798_;
wire _14799_;
wire _14800_;
wire _14801_;
wire _14802_;
wire _14803_;
wire _14804_;
wire _14805_;
wire _14806_;
wire _14807_;
wire _14808_;
wire _14809_;
wire _14810_;
wire _14811_;
wire _14812_;
wire _14813_;
wire _14814_;
wire _14815_;
wire _14816_;
wire _14817_;
wire _14818_;
wire _14819_;
wire _14820_;
wire _14821_;
wire _14822_;
wire _14823_;
wire _14824_;
wire _14825_;
wire _14826_;
wire _14827_;
wire _14828_;
wire _14829_;
wire _14830_;
wire _14831_;
wire _14832_;
wire _14833_;
wire _14834_;
wire _14835_;
wire _14836_;
wire _14837_;
wire _14838_;
wire _14839_;
wire _14840_;
wire _14841_;
wire _14842_;
wire _14843_;
wire _14844_;
wire _14845_;
wire _14846_;
wire _14847_;
wire _14848_;
wire _14849_;
wire _14850_;
wire _14851_;
wire _14852_;
wire _14853_;
wire _14854_;
wire _14855_;
wire _14856_;
wire _14857_;
wire _14858_;
wire _14859_;
wire _14860_;
wire _14861_;
wire _14862_;
wire _14863_;
wire _14864_;
wire _14865_;
wire _14866_;
wire _14867_;
wire _14868_;
wire _14869_;
wire _14870_;
wire _14871_;
wire _14872_;
wire _14873_;
wire _14874_;
wire _14875_;
wire _14876_;
wire _14877_;
wire _14878_;
wire _14879_;
wire _14880_;
wire _14881_;
wire _14882_;
wire _14883_;
wire _14884_;
wire _14885_;
wire _14886_;
wire _14887_;
wire _14888_;
wire _14889_;
wire _14890_;
wire _14891_;
wire _14892_;
wire _14893_;
wire _14894_;
wire _14895_;
wire _14896_;
wire _14897_;
wire _14898_;
wire _14899_;
wire _14900_;
wire _14901_;
wire _14902_;
wire _14903_;
wire _14904_;
wire _14905_;
wire _14906_;
wire _14907_;
wire _14908_;
wire _14909_;
wire _14910_;
wire _14911_;
wire _14912_;
wire _14913_;
wire _14914_;
wire _14915_;
wire _14916_;
wire _14917_;
wire _14918_;
wire _14919_;
wire _14920_;
wire _14921_;
wire _14922_;
wire _14923_;
wire _14924_;
wire _14925_;
wire _14926_;
wire _14927_;
wire _14928_;
wire _14929_;
wire _14930_;
wire _14931_;
wire _14932_;
wire _14933_;
wire _14934_;
wire _14935_;
wire _14936_;
wire _14937_;
wire _14938_;
wire _14939_;
wire _14940_;
wire _14941_;
wire _14942_;
wire _14943_;
wire _14944_;
wire _14945_;
wire _14946_;
wire _14947_;
wire _14948_;
wire _14949_;
wire _14950_;
wire _14951_;
wire _14952_;
wire _14953_;
wire _14954_;
wire _14955_;
wire _14956_;
wire _14957_;
wire _14958_;
wire _14959_;
wire _14960_;
wire _14961_;
wire _14962_;
wire _14963_;
wire _14964_;
wire _14965_;
wire _14966_;
wire _14967_;
wire _14968_;
wire _14969_;
wire _14970_;
wire _14971_;
wire _14972_;
wire _14973_;
wire _14974_;
wire _14975_;
wire _14976_;
wire _14977_;
wire _14978_;
wire _14979_;
wire _14980_;
wire _14981_;
wire _14982_;
wire _14983_;
wire _14984_;
wire _14985_;
wire _14986_;
wire _14987_;
wire _14988_;
wire _14989_;
wire _14990_;
wire _14991_;
wire _14992_;
wire _14993_;
wire _14994_;
wire _14995_;
wire _14996_;
wire _14997_;
wire _14998_;
wire _14999_;
wire _15000_;
wire _15001_;
wire _15002_;
wire _15003_;
wire _15004_;
wire _15005_;
wire _15006_;
wire _15007_;
wire _15008_;
wire _15009_;
wire _15010_;
wire _15011_;
wire _15012_;
wire _15013_;
wire _15014_;
wire _15015_;
wire _15016_;
wire _15017_;
wire _15018_;
wire _15019_;
wire _15020_;
wire _15021_;
wire _15022_;
wire _15023_;
wire _15024_;
wire _15025_;
wire _15026_;
wire _15027_;
wire _15028_;
wire _15029_;
wire _15030_;
wire _15031_;
wire _15032_;
wire _15033_;
wire _15034_;
wire _15035_;
wire _15036_;
wire _15037_;
wire _15038_;
wire _15039_;
wire _15040_;
wire _15041_;
wire _15042_;
wire _15043_;
wire _15044_;
wire _15045_;
wire _15046_;
wire _15047_;
wire _15048_;
wire _15049_;
wire _15050_;
wire _15051_;
wire _15052_;
wire _15053_;
wire _15054_;
wire _15055_;
wire _15056_;
wire _15057_;
wire _15058_;
wire _15059_;
wire _15060_;
wire _15061_;
wire _15062_;
wire _15063_;
wire _15064_;
wire _15065_;
wire _15066_;
wire _15067_;
wire _15068_;
wire _15069_;
wire _15070_;
wire _15071_;
wire _15072_;
wire _15073_;
wire _15074_;
wire _15075_;
wire _15076_;
wire _15077_;
wire _15078_;
wire _15079_;
wire _15080_;
wire _15081_;
wire _15082_;
wire _15083_;
wire _15084_;
wire _15085_;
wire _15086_;
wire _15087_;
wire _15088_;
wire _15089_;
wire _15090_;
wire _15091_;
wire _15092_;
wire _15093_;
wire _15094_;
wire _15095_;
wire _15096_;
wire _15097_;
wire _15098_;
wire _15099_;
wire _15100_;
wire _15101_;
wire _15102_;
wire _15103_;
wire _15104_;
wire _15105_;
wire _15106_;
wire _15107_;
wire _15108_;
wire _15109_;
wire _15110_;
wire _15111_;
wire _15112_;
wire _15113_;
wire _15114_;
wire _15115_;
wire _15116_;
wire _15117_;
wire _15118_;
wire _15119_;
wire _15120_;
wire _15121_;
wire _15122_;
wire _15123_;
wire _15124_;
wire _15125_;
wire _15126_;
wire _15127_;
wire _15128_;
wire _15129_;
wire _15130_;
wire _15131_;
wire _15132_;
wire _15133_;
wire _15134_;
wire _15135_;
wire _15136_;
wire _15137_;
wire _15138_;
wire _15139_;
wire _15140_;
wire _15141_;
wire _15142_;
wire _15143_;
wire _15144_;
wire _15145_;
wire _15146_;
wire _15147_;
wire _15148_;
wire _15149_;
wire _15150_;
wire _15151_;
wire _15152_;
wire _15153_;
wire _15154_;
wire _15155_;
wire _15156_;
wire _15157_;
wire _15158_;
wire _15159_;
wire _15160_;
wire _15161_;
wire _15162_;
wire _15163_;
wire _15164_;
wire _15165_;
wire _15166_;
wire _15167_;
wire _15168_;
wire _15169_;
wire _15170_;
wire _15171_;
wire _15172_;
wire _15173_;
wire _15174_;
wire _15175_;
wire _15176_;
wire _15177_;
wire _15178_;
wire _15179_;
wire _15180_;
wire _15181_;
wire _15182_;
wire _15183_;
wire _15184_;
wire _15185_;
wire _15186_;
wire _15187_;
wire _15188_;
wire _15189_;
wire _15190_;
wire _15191_;
wire _15192_;
wire _15193_;
wire _15194_;
wire _15195_;
wire _15196_;
wire _15197_;
wire _15198_;
wire _15199_;
wire _15200_;
wire _15201_;
wire _15202_;
wire _15203_;
wire _15204_;
wire _15205_;
wire _15206_;
wire _15207_;
wire _15208_;
wire _15209_;
wire _15210_;
wire _15211_;
wire _15212_;
wire _15213_;
wire _15214_;
wire _15215_;
wire _15216_;
wire _15217_;
wire _15218_;
wire _15219_;
wire _15220_;
wire _15221_;
wire _15222_;
wire _15223_;
wire _15224_;
wire _15225_;
wire _15226_;
wire _15227_;
wire _15228_;
wire _15229_;
wire _15230_;
wire _15231_;
wire _15232_;
wire _15233_;
wire _15234_;
wire _15235_;
wire _15236_;
wire _15237_;
wire _15238_;
wire _15239_;
wire _15240_;
wire _15241_;
wire _15242_;
wire _15243_;
wire _15244_;
wire _15245_;
wire _15246_;
wire _15247_;
wire _15248_;
wire _15249_;
wire _15250_;
wire _15251_;
wire _15252_;
wire _15253_;
wire _15254_;
wire _15255_;
wire _15256_;
wire _15257_;
wire _15258_;
wire _15259_;
wire _15260_;
wire _15261_;
wire _15262_;
wire _15263_;
wire _15264_;
wire _15265_;
wire _15266_;
wire _15267_;
wire _15268_;
wire _15269_;
wire _15270_;
wire _15271_;
wire _15272_;
wire _15273_;
wire _15274_;
wire _15275_;
wire _15276_;
wire _15277_;
wire _15278_;
wire _15279_;
wire _15280_;
wire _15281_;
wire _15282_;
wire _15283_;
wire _15284_;
wire _15285_;
wire _15286_;
wire _15287_;
wire _15288_;
wire _15289_;
wire _15290_;
wire _15291_;
wire _15292_;
wire _15293_;
wire _15294_;
wire _15295_;
wire _15296_;
wire _15297_;
wire _15298_;
wire _15299_;
wire _15300_;
wire _15301_;
wire _15302_;
wire _15303_;
wire _15304_;
wire _15305_;
wire _15306_;
wire _15307_;
wire _15308_;
wire _15309_;
wire _15310_;
wire _15311_;
wire _15312_;
wire _15313_;
wire _15314_;
wire _15315_;
wire _15316_;
wire _15317_;
wire _15318_;
wire _15319_;
wire _15320_;
wire _15321_;
wire _15322_;
wire _15323_;
wire _15324_;
wire _15325_;
wire _15326_;
wire _15327_;
wire _15328_;
wire _15329_;
wire _15330_;
wire _15331_;
wire _15332_;
wire _15333_;
wire _15334_;
wire _15335_;
wire _15336_;
wire _15337_;
wire _15338_;
wire _15339_;
wire _15340_;
wire _15341_;
wire _15342_;
wire _15343_;
wire _15344_;
wire _15345_;
wire _15346_;
wire _15347_;
wire _15348_;
wire _15349_;
wire _15350_;
wire _15351_;
wire _15352_;
wire _15353_;
wire _15354_;
wire _15355_;
wire _15356_;
wire _15357_;
wire _15358_;
wire _15359_;
wire _15360_;
wire _15361_;
wire _15362_;
wire _15363_;
wire _15364_;
wire _15365_;
wire _15366_;
wire _15367_;
wire _15368_;
wire _15369_;
wire _15370_;
wire _15371_;
wire _15372_;
wire _15373_;
wire _15374_;
wire _15375_;
wire _15376_;
wire _15377_;
wire _15378_;
wire _15379_;
wire _15380_;
wire _15381_;
wire _15382_;
wire _15383_;
wire _15384_;
wire _15385_;
wire _15386_;
wire _15387_;
wire _15388_;
wire _15389_;
wire _15390_;
wire _15391_;
wire _15392_;
wire _15393_;
wire _15394_;
wire _15395_;
wire _15396_;
wire _15397_;
wire _15398_;
wire _15399_;
wire _15400_;
wire _15401_;
wire _15402_;
wire _15403_;
wire _15404_;
wire _15405_;
wire _15406_;
wire _15407_;
wire _15408_;
wire _15409_;
wire _15410_;
wire _15411_;
wire _15412_;
wire _15413_;
wire _15414_;
wire _15415_;
wire _15416_;
wire _15417_;
wire _15418_;
wire _15419_;
wire _15420_;
wire _15421_;
wire _15422_;
wire _15423_;
wire _15424_;
wire _15425_;
wire _15426_;
wire _15427_;
wire _15428_;
wire _15429_;
wire _15430_;
wire _15431_;
wire _15432_;
wire _15433_;
wire _15434_;
wire _15435_;
wire _15436_;
wire _15437_;
wire _15438_;
wire _15439_;
wire _15440_;
wire _15441_;
wire _15442_;
wire _15443_;
wire _15444_;
wire _15445_;
wire _15446_;
wire _15447_;
wire _15448_;
wire _15449_;
wire _15450_;
wire _15451_;
wire _15452_;
wire _15453_;
wire _15454_;
wire _15455_;
wire _15456_;
wire _15457_;
wire _15458_;
wire _15459_;
wire _15460_;
wire _15461_;
wire _15462_;
wire _15463_;
wire _15464_;
wire _15465_;
wire _15466_;
wire _15467_;
wire _15468_;
wire _15469_;
wire _15470_;
wire _15471_;
wire _15472_;
wire _15473_;
wire _15474_;
wire _15475_;
wire _15476_;
wire _15477_;
wire _15478_;
wire _15479_;
wire _15480_;
wire _15481_;
wire _15482_;
wire _15483_;
wire _15484_;
wire _15485_;
wire _15486_;
wire _15487_;
wire _15488_;
wire _15489_;
wire _15490_;
wire _15491_;
wire _15492_;
wire _15493_;
wire _15494_;
wire _15495_;
wire _15496_;
wire _15497_;
wire _15498_;
wire _15499_;
wire _15500_;
wire _15501_;
wire _15502_;
wire _15503_;
wire _15504_;
wire _15505_;
wire _15506_;
wire _15507_;
wire _15508_;
wire _15509_;
wire _15510_;
wire _15511_;
wire _15512_;
wire _15513_;
wire _15514_;
wire _15515_;
wire _15516_;
wire _15517_;
wire _15518_;
wire _15519_;
wire _15520_;
wire _15521_;
wire _15522_;
wire _15523_;
wire _15524_;
wire _15525_;
wire _15526_;
wire _15527_;
wire _15528_;
wire _15529_;
wire _15530_;
wire _15531_;
wire _15532_;
wire _15533_;
wire _15534_;
wire _15535_;
wire _15536_;
wire _15537_;
wire _15538_;
wire _15539_;
wire _15540_;
wire _15541_;
wire _15542_;
wire _15543_;
wire _15544_;
wire _15545_;
wire _15546_;
wire _15547_;
wire _15548_;
wire _15549_;
wire _15550_;
wire _15551_;
wire _15552_;
wire _15553_;
wire _15554_;
wire _15555_;
wire _15556_;
wire _15557_;
wire _15558_;
wire _15559_;
wire _15560_;
wire _15561_;
wire _15562_;
wire _15563_;
wire _15564_;
wire _15565_;
wire _15566_;
wire _15567_;
wire _15568_;
wire _15569_;
wire _15570_;
wire _15571_;
wire _15572_;
wire _15573_;
wire _15574_;
wire _15575_;
wire _15576_;
wire _15577_;
wire _15578_;
wire _15579_;
wire _15580_;
wire _15581_;
wire _15582_;
wire _15583_;
wire _15584_;
wire _15585_;
wire _15586_;
wire _15587_;
wire _15588_;
wire _15589_;
wire _15590_;
wire _15591_;
wire _15592_;
wire _15593_;
wire _15594_;
wire _15595_;
wire _15596_;
wire _15597_;
wire _15598_;
wire _15599_;
wire _15600_;
wire _15601_;
wire _15602_;
wire _15603_;
wire _15604_;
wire _15605_;
wire _15606_;
wire _15607_;
wire _15608_;
wire _15609_;
wire _15610_;
wire _15611_;
wire _15612_;
wire _15613_;
wire _15614_;
wire _15615_;
wire _15616_;
wire _15617_;
wire _15618_;
wire _15619_;
wire _15620_;
wire _15621_;
wire _15622_;
wire _15623_;
wire _15624_;
wire _15625_;
wire _15626_;
wire _15627_;
wire _15628_;
wire _15629_;
wire _15630_;
wire _15631_;
wire _15632_;
wire _15633_;
wire _15634_;
wire _15635_;
wire _15636_;
wire _15637_;
wire _15638_;
wire _15639_;
wire _15640_;
wire _15641_;
wire _15642_;
wire _15643_;
wire _15644_;
wire _15645_;
wire _15646_;
wire _15647_;
wire _15648_;
wire _15649_;
wire _15650_;
wire _15651_;
wire _15652_;
wire _15653_;
wire _15654_;
wire _15655_;
wire _15656_;
wire _15657_;
wire _15658_;
wire _15659_;
wire _15660_;
wire _15661_;
wire _15662_;
wire _15663_;
wire _15664_;
wire _15665_;
wire _15666_;
wire _15667_;
wire _15668_;
wire _15669_;
wire _15670_;
wire _15671_;
wire _15672_;
wire _15673_;
wire _15674_;
wire _15675_;
wire _15676_;
wire _15677_;
wire _15678_;
wire _15679_;
wire _15680_;
wire _15681_;
wire _15682_;
wire _15683_;
wire _15684_;
wire _15685_;
wire _15686_;
wire _15687_;
wire _15688_;
wire _15689_;
wire _15690_;
wire _15691_;
wire _15692_;
wire _15693_;
wire _15694_;
wire _15695_;
wire _15696_;
wire _15697_;
wire _15698_;
wire _15699_;
wire _15700_;
wire _15701_;
wire _15702_;
wire _15703_;
wire _15704_;
wire _15705_;
wire _15706_;
wire _15707_;
wire _15708_;
wire _15709_;
wire _15710_;
wire _15711_;
wire _15712_;
wire _15713_;
wire _15714_;
wire _15715_;
wire _15716_;
wire _15717_;
wire _15718_;
wire _15719_;
wire _15720_;
wire _15721_;
wire _15722_;
wire _15723_;
wire _15724_;
wire _15725_;
wire _15726_;
wire _15727_;
wire _15728_;
wire _15729_;
wire _15730_;
wire _15731_;
wire _15732_;
wire _15733_;
wire _15734_;
wire _15735_;
wire _15736_;
wire _15737_;
wire _15738_;
wire _15739_;
wire _15740_;
wire _15741_;
wire _15742_;
wire _15743_;
wire _15744_;
wire _15745_;
wire _15746_;
wire _15747_;
wire _15748_;
wire _15749_;
wire _15750_;
wire _15751_;
wire _15752_;
wire _15753_;
wire _15754_;
wire _15755_;
wire _15756_;
wire _15757_;
wire _15758_;
wire _15759_;
wire _15760_;
wire _15761_;
wire _15762_;
wire _15763_;
wire _15764_;
wire _15765_;
wire _15766_;
wire _15767_;
wire _15768_;
wire _15769_;
wire _15770_;
wire _15771_;
wire _15772_;
wire _15773_;
wire _15774_;
wire _15775_;
wire _15776_;
wire _15777_;
wire _15778_;
wire _15779_;
wire _15780_;
wire _15781_;
wire _15782_;
wire _15783_;
wire _15784_;
wire _15785_;
wire _15786_;
wire _15787_;
wire _15788_;
wire _15789_;
wire _15790_;
wire _15791_;
wire _15792_;
wire _15793_;
wire _15794_;
wire _15795_;
wire _15796_;
wire _15797_;
wire _15798_;
wire _15799_;
wire _15800_;
wire _15801_;
wire _15802_;
wire _15803_;
wire _15804_;
wire _15805_;
wire _15806_;
wire _15807_;
wire _15808_;
wire _15809_;
wire _15810_;
wire _15811_;
wire _15812_;
wire _15813_;
wire _15814_;
wire _15815_;
wire _15816_;
wire _15817_;
wire _15818_;
wire _15819_;
wire _15820_;
wire _15821_;
wire _15822_;
wire _15823_;
wire _15824_;
wire _15825_;
wire _15826_;
wire _15827_;
wire _15828_;
wire _15829_;
wire _15830_;
wire _15831_;
wire _15832_;
wire _15833_;
wire _15834_;
wire _15835_;
wire _15836_;
wire _15837_;
wire _15838_;
wire _15839_;
wire _15840_;
wire _15841_;
wire _15842_;
wire _15843_;
wire _15844_;
wire _15845_;
wire _15846_;
wire _15847_;
wire _15848_;
wire _15849_;
wire _15850_;
wire _15851_;
wire _15852_;
wire _15853_;
wire _15854_;
wire _15855_;
wire _15856_;
wire _15857_;
wire _15858_;
wire _15859_;
wire _15860_;
wire _15861_;
wire _15862_;
wire _15863_;
wire _15864_;
wire _15865_;
wire _15866_;
wire _15867_;
wire _15868_;
wire _15869_;
wire _15870_;
wire _15871_;
wire _15872_;
wire _15873_;
wire _15874_;
wire _15875_;
wire _15876_;
wire _15877_;
wire _15878_;
wire _15879_;
wire _15880_;
wire _15881_;
wire _15882_;
wire _15883_;
wire _15884_;
wire _15885_;
wire _15886_;
wire _15887_;
wire _15888_;
wire _15889_;
wire _15890_;
wire _15891_;
wire _15892_;
wire _15893_;
wire _15894_;
wire _15895_;
wire _15896_;
wire _15897_;
wire _15898_;
wire _15899_;
wire _15900_;
wire _15901_;
wire _15902_;
wire _15903_;
wire _15904_;
wire _15905_;
wire _15906_;
wire _15907_;
wire _15908_;
wire _15909_;
wire _15910_;
wire _15911_;
wire _15912_;
wire _15913_;
wire _15914_;
wire _15915_;
wire _15916_;
wire _15917_;
wire _15918_;
wire _15919_;
wire _15920_;
wire _15921_;
wire _15922_;
wire _15923_;
wire _15924_;
wire _15925_;
wire _15926_;
wire _15927_;
wire _15928_;
wire _15929_;
wire _15930_;
wire _15931_;
wire _15932_;
wire _15933_;
wire _15934_;
wire _15935_;
wire _15936_;
wire _15937_;
wire _15938_;
wire _15939_;
wire _15940_;
wire _15941_;
wire _15942_;
wire _15943_;
wire _15944_;
wire _15945_;
wire _15946_;
wire _15947_;
wire _15948_;
wire _15949_;
wire _15950_;
wire _15951_;
wire _15952_;
wire _15953_;
wire _15954_;
wire _15955_;
wire _15956_;
wire _15957_;
wire _15958_;
wire _15959_;
wire _15960_;
wire _15961_;
wire _15962_;
wire _15963_;
wire _15964_;
wire _15965_;
wire _15966_;
wire _15967_;
wire _15968_;
wire _15969_;
wire _15970_;
wire _15971_;
wire _15972_;
wire _15973_;
wire _15974_;
wire _15975_;
wire _15976_;
wire _15977_;
wire _15978_;
wire _15979_;
wire _15980_;
wire _15981_;
wire _15982_;
wire _15983_;
wire _15984_;
wire _15985_;
wire _15986_;
wire _15987_;
wire _15988_;
wire _15989_;
wire _15990_;
wire _15991_;
wire _15992_;
wire _15993_;
wire _15994_;
wire _15995_;
wire _15996_;
wire _15997_;
wire _15998_;
wire _15999_;
wire _16000_;
wire _16001_;
wire _16002_;
wire _16003_;
wire _16004_;
wire _16005_;
wire _16006_;
wire _16007_;
wire _16008_;
wire _16009_;
wire _16010_;
wire _16011_;
wire _16012_;
wire _16013_;
wire _16014_;
wire _16015_;
wire _16016_;
wire _16017_;
wire _16018_;
wire _16019_;
wire _16020_;
wire _16021_;
wire _16022_;
wire _16023_;
wire _16024_;
wire _16025_;
wire _16026_;
wire _16027_;
wire _16028_;
wire _16029_;
wire _16030_;
wire _16031_;
wire _16032_;
wire _16033_;
wire _16034_;
wire _16035_;
wire _16036_;
wire _16037_;
wire _16038_;
wire _16039_;
wire _16040_;
wire _16041_;
wire _16042_;
wire _16043_;
wire _16044_;
wire _16045_;
wire _16046_;
wire _16047_;
wire _16048_;
wire _16049_;
wire _16050_;
wire _16051_;
wire _16052_;
wire _16053_;
wire _16054_;
wire _16055_;
wire _16056_;
wire _16057_;
wire _16058_;
wire _16059_;
wire _16060_;
wire _16061_;
wire _16062_;
wire _16063_;
wire _16064_;
wire _16065_;
wire _16066_;
wire _16067_;
wire _16068_;
wire _16069_;
wire _16070_;
wire _16071_;
wire _16072_;
wire _16073_;
wire _16074_;
wire _16075_;
wire _16076_;
wire _16077_;
wire _16078_;
wire _16079_;
wire _16080_;
wire _16081_;
wire _16082_;
wire _16083_;
wire _16084_;
wire _16085_;
wire _16086_;
wire _16087_;
wire _16088_;
wire _16089_;
wire _16090_;
wire _16091_;
wire _16092_;
wire _16093_;
wire _16094_;
wire _16095_;
wire _16096_;
wire _16097_;
wire _16098_;
wire _16099_;
wire _16100_;
wire _16101_;
wire _16102_;
wire _16103_;
wire _16104_;
wire _16105_;
wire _16106_;
wire _16107_;
wire _16108_;
wire _16109_;
wire _16110_;
wire _16111_;
wire _16112_;
wire _16113_;
wire _16114_;
wire _16115_;
wire _16116_;
wire _16117_;
wire _16118_;
wire _16119_;
wire _16120_;
wire _16121_;
wire _16122_;
wire _16123_;
wire _16124_;
wire _16125_;
wire _16126_;
wire _16127_;
wire _16128_;
wire _16129_;
wire _16130_;
wire _16131_;
wire _16132_;
wire _16133_;
wire _16134_;
wire _16135_;
wire _16136_;
wire _16137_;
wire _16138_;
wire _16139_;
wire _16140_;
wire _16141_;
wire _16142_;
wire _16143_;
wire _16144_;
wire _16145_;
wire _16146_;
wire _16147_;
wire _16148_;
wire _16149_;
wire _16150_;
wire _16151_;
wire _16152_;
wire _16153_;
wire _16154_;
wire _16155_;
wire _16156_;
wire _16157_;
wire _16158_;
wire _16159_;
wire _16160_;
wire _16161_;
wire _16162_;
wire _16163_;
wire _16164_;
wire _16165_;
wire _16166_;
wire _16167_;
wire _16168_;
wire _16169_;
wire _16170_;
wire _16171_;
wire _16172_;
wire _16173_;
wire _16174_;
wire _16175_;
wire _16176_;
wire _16177_;
wire _16178_;
wire _16179_;
wire _16180_;
wire _16181_;
wire _16182_;
wire _16183_;
wire _16184_;
wire _16185_;
wire _16186_;
wire _16187_;
wire _16188_;
wire _16189_;
wire _16190_;
wire _16191_;
wire _16192_;
wire _16193_;
wire _16194_;
wire _16195_;
wire _16196_;
wire _16197_;
wire _16198_;
wire _16199_;
wire _16200_;
wire _16201_;
wire _16202_;
wire _16203_;
wire _16204_;
wire _16205_;
wire _16206_;
wire _16207_;
wire _16208_;
wire _16209_;
wire _16210_;
wire _16211_;
wire _16212_;
wire _16213_;
wire _16214_;
wire _16215_;
wire _16216_;
wire _16217_;
wire _16218_;
wire _16219_;
wire _16220_;
wire _16221_;
wire _16222_;
wire _16223_;
wire _16224_;
wire _16225_;
wire _16226_;
wire _16227_;
wire _16228_;
wire _16229_;
wire _16230_;
wire _16231_;
wire _16232_;
wire _16233_;
wire _16234_;
wire _16235_;
wire _16236_;
wire _16237_;
wire _16238_;
wire _16239_;
wire _16240_;
wire _16241_;
wire _16242_;
wire _16243_;
wire _16244_;
wire _16245_;
wire _16246_;
wire _16247_;
wire _16248_;
wire _16249_;
wire _16250_;
wire _16251_;
wire _16252_;
wire _16253_;
wire _16254_;
wire _16255_;
wire _16256_;
wire _16257_;
wire _16258_;
wire _16259_;
wire _16260_;
wire _16261_;
wire _16262_;
wire _16263_;
wire _16264_;
wire _16265_;
wire _16266_;
wire _16267_;
wire _16268_;
wire _16269_;
wire _16270_;
wire _16271_;
wire _16272_;
wire _16273_;
wire _16274_;
wire _16275_;
wire _16276_;
wire _16277_;
wire _16278_;
wire _16279_;
wire _16280_;
wire _16281_;
wire _16282_;
wire _16283_;
wire _16284_;
wire _16285_;
wire _16286_;
wire _16287_;
wire _16288_;
wire _16289_;
wire _16290_;
wire _16291_;
wire _16292_;
wire _16293_;
wire _16294_;
wire _16295_;
wire _16296_;
wire _16297_;
wire _16298_;
wire _16299_;
wire _16300_;
wire _16301_;
wire _16302_;
wire _16303_;
wire _16304_;
wire _16305_;
wire _16306_;
wire _16307_;
wire _16308_;
wire _16309_;
wire _16310_;
wire _16311_;
wire _16312_;
wire _16313_;
wire _16314_;
wire _16315_;
wire _16316_;
wire _16317_;
wire _16318_;
wire _16319_;
wire _16320_;
wire _16321_;
wire _16322_;
wire _16323_;
wire _16324_;
wire _16325_;
wire _16326_;
wire _16327_;
wire _16328_;
wire _16329_;
wire _16330_;
wire _16331_;
wire _16332_;
wire _16333_;
wire _16334_;
wire _16335_;
wire _16336_;
wire _16337_;
wire _16338_;
wire _16339_;
wire _16340_;
wire _16341_;
wire _16342_;
wire _16343_;
wire _16344_;
wire _16345_;
wire _16346_;
wire _16347_;
wire _16348_;
wire _16349_;
wire _16350_;
wire _16351_;
wire _16352_;
wire _16353_;
wire _16354_;
wire _16355_;
wire _16356_;
wire _16357_;
wire _16358_;
wire _16359_;
wire _16360_;
wire _16361_;
wire _16362_;
wire _16363_;
wire _16364_;
wire _16365_;
wire _16366_;
wire _16367_;
wire _16368_;
wire _16369_;
wire _16370_;
wire _16371_;
wire _16372_;
wire _16373_;
wire _16374_;
wire _16375_;
wire _16376_;
wire _16377_;
wire _16378_;
wire _16379_;
wire _16380_;
wire _16381_;
wire _16382_;
wire _16383_;
wire _16384_;
wire _16385_;
wire _16386_;
wire _16387_;
wire _16388_;
wire _16389_;
wire _16390_;
wire _16391_;
wire _16392_;
wire _16393_;
wire _16394_;
wire _16395_;
wire _16396_;
wire _16397_;
wire _16398_;
wire _16399_;
wire _16400_;
wire _16401_;
wire _16402_;
wire _16403_;
wire _16404_;
wire _16405_;
wire _16406_;
wire _16407_;
wire _16408_;
wire _16409_;
wire _16410_;
wire _16411_;
wire _16412_;
wire _16413_;
wire _16414_;
wire _16415_;
wire _16416_;
wire _16417_;
wire _16418_;
wire _16419_;
wire _16420_;
wire _16421_;
wire _16422_;
wire _16423_;
wire _16424_;
wire _16425_;
wire _16426_;
wire _16427_;
wire _16428_;
wire _16429_;
wire _16430_;
wire _16431_;
wire _16432_;
wire _16433_;
wire _16434_;
wire _16435_;
wire _16436_;
wire _16437_;
wire _16438_;
wire _16439_;
wire _16440_;
wire _16441_;
wire _16442_;
wire _16443_;
wire _16444_;
wire _16445_;
wire _16446_;
wire _16447_;
wire _16448_;
wire _16449_;
wire _16450_;
wire _16451_;
wire _16452_;
wire _16453_;
wire _16454_;
wire _16455_;
wire _16456_;
wire _16457_;
wire _16458_;
wire _16459_;
wire _16460_;
wire _16461_;
wire _16462_;
wire _16463_;
wire _16464_;
wire _16465_;
wire _16466_;
wire _16467_;
wire _16468_;
wire _16469_;
wire _16470_;
wire _16471_;
wire _16472_;
wire _16473_;
wire _16474_;
wire _16475_;
wire _16476_;
wire _16477_;
wire _16478_;
wire _16479_;
wire _16480_;
wire _16481_;
wire _16482_;
wire _16483_;
wire _16484_;
wire _16485_;
wire _16486_;
wire _16487_;
wire _16488_;
wire _16489_;
wire _16490_;
wire _16491_;
wire _16492_;
wire _16493_;
wire _16494_;
wire _16495_;
wire _16496_;
wire _16497_;
wire _16498_;
wire _16499_;
wire _16500_;
wire _16501_;
wire _16502_;
wire _16503_;
wire _16504_;
wire _16505_;
wire _16506_;
wire _16507_;
wire _16508_;
wire _16509_;
wire _16510_;
wire _16511_;
wire _16512_;
wire _16513_;
wire _16514_;
wire _16515_;
wire _16516_;
wire _16517_;
wire _16518_;
wire _16519_;
wire _16520_;
wire _16521_;
wire _16522_;
wire _16523_;
wire _16524_;
wire _16525_;
wire _16526_;
wire _16527_;
wire _16528_;
wire _16529_;
wire _16530_;
wire _16531_;
wire _16532_;
wire _16533_;
wire _16534_;
wire _16535_;
wire _16536_;
wire _16537_;
wire _16538_;
wire _16539_;
wire _16540_;
wire _16541_;
wire _16542_;
wire _16543_;
wire _16544_;
wire _16545_;
wire _16546_;
wire _16547_;
wire _16548_;
wire _16549_;
wire _16550_;
wire _16551_;
wire _16552_;
wire _16553_;
wire _16554_;
wire _16555_;
wire _16556_;
wire _16557_;
wire _16558_;
wire _16559_;
wire _16560_;
wire _16561_;
wire _16562_;
wire _16563_;
wire _16564_;
wire _16565_;
wire _16566_;
wire _16567_;
wire _16568_;
wire _16569_;
wire _16570_;
wire _16571_;
wire _16572_;
wire _16573_;
wire _16574_;
wire _16575_;
wire _16576_;
wire _16577_;
wire _16578_;
wire _16579_;
wire _16580_;
wire _16581_;
wire _16582_;
wire _16583_;
wire _16584_;
wire _16585_;
wire _16586_;
wire _16587_;
wire _16588_;
wire _16589_;
wire _16590_;
wire _16591_;
wire _16592_;
wire _16593_;
wire _16594_;
wire _16595_;
wire _16596_;
wire _16597_;
wire _16598_;
wire _16599_;
wire _16600_;
wire _16601_;
wire _16602_;
wire _16603_;
wire _16604_;
wire _16605_;
wire _16606_;
wire _16607_;
wire _16608_;
wire _16609_;
wire _16610_;
wire _16611_;
wire _16612_;
wire _16613_;
wire _16614_;
wire _16615_;
wire _16616_;
wire _16617_;
wire _16618_;
wire _16619_;
wire _16620_;
wire _16621_;
wire _16622_;
wire _16623_;
wire _16624_;
wire _16625_;
wire _16626_;
wire _16627_;
wire _16628_;
wire _16629_;
wire _16630_;
wire _16631_;
wire _16632_;
wire _16633_;
wire _16634_;
wire _16635_;
wire _16636_;
wire _16637_;
wire _16638_;
wire _16639_;
wire _16640_;
wire _16641_;
wire _16642_;
wire _16643_;
wire _16644_;
wire _16645_;
wire _16646_;
wire _16647_;
wire _16648_;
wire _16649_;
wire _16650_;
wire _16651_;
wire _16652_;
wire _16653_;
wire _16654_;
wire _16655_;
wire _16656_;
wire _16657_;
wire _16658_;
wire _16659_;
wire _16660_;
wire _16661_;
wire _16662_;
wire _16663_;
wire _16664_;
wire _16665_;
wire _16666_;
wire _16667_;
wire _16668_;
wire _16669_;
wire _16670_;
wire _16671_;
wire _16672_;
wire _16673_;
wire _16674_;
wire _16675_;
wire _16676_;
wire _16677_;
wire _16678_;
wire _16679_;
wire _16680_;
wire _16681_;
wire _16682_;
wire _16683_;
wire _16684_;
wire _16685_;
wire _16686_;
wire _16687_;
wire _16688_;
wire _16689_;
wire _16690_;
wire _16691_;
wire _16692_;
wire _16693_;
wire _16694_;
wire _16695_;
wire _16696_;
wire _16697_;
wire _16698_;
wire _16699_;
wire _16700_;
wire _16701_;
wire _16702_;
wire _16703_;
wire _16704_;
wire _16705_;
wire _16706_;
wire _16707_;
wire _16708_;
wire _16709_;
wire _16710_;
wire _16711_;
wire _16712_;
wire _16713_;
wire _16714_;
wire _16715_;
wire _16716_;
wire _16717_;
wire _16718_;
wire _16719_;
wire _16720_;
wire _16721_;
wire _16722_;
wire _16723_;
wire _16724_;
wire _16725_;
wire _16726_;
wire _16727_;
wire _16728_;
wire _16729_;
wire _16730_;
wire _16731_;
wire _16732_;
wire _16733_;
wire _16734_;
wire _16735_;
wire _16736_;
wire _16737_;
wire _16738_;
wire _16739_;
wire _16740_;
wire _16741_;
wire _16742_;
wire _16743_;
wire _16744_;
wire _16745_;
wire _16746_;
wire _16747_;
wire _16748_;
wire _16749_;
wire _16750_;
wire _16751_;
wire _16752_;
wire _16753_;
wire _16754_;
wire _16755_;
wire _16756_;
wire _16757_;
wire _16758_;
wire _16759_;
wire _16760_;
wire _16761_;
wire _16762_;
wire _16763_;
wire _16764_;
wire _16765_;
wire _16766_;
wire _16767_;
wire _16768_;
wire _16769_;
wire _16770_;
wire _16771_;
wire _16772_;
wire _16773_;
wire _16774_;
wire _16775_;
wire _16776_;
wire _16777_;
wire _16778_;
wire _16779_;
wire _16780_;
wire _16781_;
wire _16782_;
wire _16783_;
wire _16784_;
wire _16785_;
wire _16786_;
wire _16787_;
wire _16788_;
wire _16789_;
wire _16790_;
wire _16791_;
wire _16792_;
wire _16793_;
wire _16794_;
wire _16795_;
wire _16796_;
wire _16797_;
wire _16798_;
wire _16799_;
wire _16800_;
wire _16801_;
wire _16802_;
wire _16803_;
wire _16804_;
wire _16805_;
wire _16806_;
wire _16807_;
wire _16808_;
wire _16809_;
wire _16810_;
wire _16811_;
wire _16812_;
wire _16813_;
wire _16814_;
wire _16815_;
wire _16816_;
wire _16817_;
wire _16818_;
wire _16819_;
wire _16820_;
wire _16821_;
wire _16822_;
wire _16823_;
wire _16824_;
wire _16825_;
wire _16826_;
wire _16827_;
wire _16828_;
wire _16829_;
wire _16830_;
wire _16831_;
wire _16832_;
wire _16833_;
wire _16834_;
wire _16835_;
wire _16836_;
wire _16837_;
wire _16838_;
wire _16839_;
wire _16840_;
wire _16841_;
wire _16842_;
wire _16843_;
wire _16844_;
wire _16845_;
wire _16846_;
wire _16847_;
wire _16848_;
wire _16849_;
wire _16850_;
wire _16851_;
wire _16852_;
wire _16853_;
wire _16854_;
wire _16855_;
wire _16856_;
wire _16857_;
wire _16858_;
wire _16859_;
wire _16860_;
wire _16861_;
wire _16862_;
wire _16863_;
wire _16864_;
wire _16865_;
wire _16866_;
wire _16867_;
wire _16868_;
wire _16869_;
wire _16870_;
wire _16871_;
wire _16872_;
wire _16873_;
wire _16874_;
wire _16875_;
wire _16876_;
wire _16877_;
wire _16878_;
wire _16879_;
wire _16880_;
wire _16881_;
wire _16882_;
wire _16883_;
wire _16884_;
wire _16885_;
wire _16886_;
wire _16887_;
wire _16888_;
wire _16889_;
wire _16890_;
wire _16891_;
wire _16892_;
wire _16893_;
wire _16894_;
wire _16895_;
wire _16896_;
wire _16897_;
wire _16898_;
wire _16899_;
wire _16900_;
wire _16901_;
wire _16902_;
wire _16903_;
wire _16904_;
wire _16905_;
wire _16906_;
wire _16907_;
wire _16908_;
wire _16909_;
wire _16910_;
wire _16911_;
wire _16912_;
wire _16913_;
wire _16914_;
wire _16915_;
wire _16916_;
wire _16917_;
wire _16918_;
wire _16919_;
wire _16920_;
wire _16921_;
wire _16922_;
wire _16923_;
wire _16924_;
wire _16925_;
wire _16926_;
wire _16927_;
wire _16928_;
wire _16929_;
wire _16930_;
wire _16931_;
wire _16932_;
wire _16933_;
wire _16934_;
wire _16935_;
wire _16936_;
wire _16937_;
wire _16938_;
wire _16939_;
wire _16940_;
wire _16941_;
wire _16942_;
wire _16943_;
wire _16944_;
wire _16945_;
wire _16946_;
wire _16947_;
wire _16948_;
wire _16949_;
wire _16950_;
wire _16951_;
wire _16952_;
wire _16953_;
wire _16954_;
wire _16955_;
wire _16956_;
wire _16957_;
wire _16958_;
wire _16959_;
wire _16960_;
wire _16961_;
wire _16962_;
wire _16963_;
wire _16964_;
wire _16965_;
wire _16966_;
wire _16967_;
wire _16968_;
wire _16969_;
wire _16970_;
wire _16971_;
wire _16972_;
wire _16973_;
wire _16974_;
wire _16975_;
wire _16976_;
wire _16977_;
wire _16978_;
wire _16979_;
wire _16980_;
wire _16981_;
wire _16982_;
wire _16983_;
wire _16984_;
wire _16985_;
wire _16986_;
wire _16987_;
wire _16988_;
wire _16989_;
wire _16990_;
wire _16991_;
wire _16992_;
wire _16993_;
wire _16994_;
wire _16995_;
wire _16996_;
wire _16997_;
wire _16998_;
wire _16999_;
wire _17000_;
wire _17001_;
wire _17002_;
wire _17003_;
wire _17004_;
wire _17005_;
wire _17006_;
wire _17007_;
wire _17008_;
wire _17009_;
wire _17010_;
wire _17011_;
wire _17012_;
wire _17013_;
wire _17014_;
wire _17015_;
wire _17016_;
wire _17017_;
wire _17018_;
wire _17019_;
wire _17020_;
wire _17021_;
wire _17022_;
wire _17023_;
wire _17024_;
wire _17025_;
wire _17026_;
wire _17027_;
wire _17028_;
wire _17029_;
wire _17030_;
wire _17031_;
wire _17032_;
wire _17033_;
wire _17034_;
wire _17035_;
wire _17036_;
wire _17037_;
wire _17038_;
wire _17039_;
wire _17040_;
wire _17041_;
wire _17042_;
wire _17043_;
wire _17044_;
wire _17045_;
wire _17046_;
wire _17047_;
wire _17048_;
wire _17049_;
wire _17050_;
wire _17051_;
wire _17052_;
wire _17053_;
wire _17054_;
wire _17055_;
wire _17056_;
wire _17057_;
wire _17058_;
wire _17059_;
wire _17060_;
wire _17061_;
wire _17062_;
wire _17063_;
wire _17064_;
wire _17065_;
wire _17066_;
wire _17067_;
wire _17068_;
wire _17069_;
wire _17070_;
wire _17071_;
wire _17072_;
wire _17073_;
wire _17074_;
wire _17075_;
wire _17076_;
wire _17077_;
wire _17078_;
wire _17079_;
wire _17080_;
wire _17081_;
wire _17082_;
wire _17083_;
wire _17084_;
wire _17085_;
wire _17086_;
wire _17087_;
wire _17088_;
wire _17089_;
wire _17090_;
wire _17091_;
wire _17092_;
wire _17093_;
wire _17094_;
wire _17095_;
wire _17096_;
wire _17097_;
wire _17098_;
wire _17099_;
wire _17100_;
wire _17101_;
wire _17102_;
wire _17103_;
wire _17104_;
wire _17105_;
wire _17106_;
wire _17107_;
wire _17108_;
wire _17109_;
wire _17110_;
wire _17111_;
wire _17112_;
wire _17113_;
wire _17114_;
wire _17115_;
wire _17116_;
wire _17117_;
wire _17118_;
wire _17119_;
wire _17120_;
wire _17121_;
wire _17122_;
wire _17123_;
wire _17124_;
wire _17125_;
wire _17126_;
wire _17127_;
wire _17128_;
wire _17129_;
wire _17130_;
wire _17131_;
wire _17132_;
wire _17133_;
wire _17134_;
wire _17135_;
wire _17136_;
wire _17137_;
wire _17138_;
wire _17139_;
wire _17140_;
wire _17141_;
wire _17142_;
wire _17143_;
wire _17144_;
wire _17145_;
wire _17146_;
wire _17147_;
wire _17148_;
wire _17149_;
wire _17150_;
wire _17151_;
wire _17152_;
wire _17153_;
wire _17154_;
wire _17155_;
wire _17156_;
wire _17157_;
wire _17158_;
wire _17159_;
wire _17160_;
wire _17161_;
wire _17162_;
wire _17163_;
wire _17164_;
wire _17165_;
wire _17166_;
wire _17167_;
wire _17168_;
wire _17169_;
wire _17170_;
wire _17171_;
wire _17172_;
wire _17173_;
wire _17174_;
wire _17175_;
wire _17176_;
wire _17177_;
wire _17178_;
wire _17179_;
wire _17180_;
wire _17181_;
wire _17182_;
wire _17183_;
wire _17184_;
wire _17185_;
wire _17186_;
wire _17187_;
wire _17188_;
wire _17189_;
wire _17190_;
wire _17191_;
wire _17192_;
wire _17193_;
wire _17194_;
wire _17195_;
wire _17196_;
wire _17197_;
wire _17198_;
wire _17199_;
wire _17200_;
wire _17201_;
wire _17202_;
wire _17203_;
wire _17204_;
wire _17205_;
wire _17206_;
wire _17207_;
wire _17208_;
wire _17209_;
wire _17210_;
wire _17211_;
wire _17212_;
wire _17213_;
wire _17214_;
wire _17215_;
wire _17216_;
wire _17217_;
wire _17218_;
wire _17219_;
wire _17220_;
wire _17221_;
wire _17222_;
wire _17223_;
wire _17224_;
wire _17225_;
wire _17226_;
wire _17227_;
wire _17228_;
wire _17229_;
wire _17230_;
wire _17231_;
wire _17232_;
wire _17233_;
wire _17234_;
wire _17235_;
wire _17236_;
wire _17237_;
wire _17238_;
wire _17239_;
wire _17240_;
wire _17241_;
wire _17242_;
wire _17243_;
wire _17244_;
wire _17245_;
wire _17246_;
wire _17247_;
wire _17248_;
wire _17249_;
wire _17250_;
wire _17251_;
wire _17252_;
wire _17253_;
wire _17254_;
wire _17255_;
wire _17256_;
wire _17257_;
wire _17258_;
wire _17259_;
wire _17260_;
wire _17261_;
wire _17262_;
wire _17263_;
wire _17264_;
wire _17265_;
wire _17266_;
wire _17267_;
wire _17268_;
wire _17269_;
wire _17270_;
wire _17271_;
wire _17272_;
wire _17273_;
wire _17274_;
wire _17275_;
wire _17276_;
wire _17277_;
wire _17278_;
wire _17279_;
wire _17280_;
wire _17281_;
wire _17282_;
wire _17283_;
wire _17284_;
wire _17285_;
wire _17286_;
wire _17287_;
wire _17288_;
wire _17289_;
wire _17290_;
wire _17291_;
wire _17292_;
wire _17293_;
wire _17294_;
wire _17295_;
wire _17296_;
wire _17297_;
wire _17298_;
wire _17299_;
wire _17300_;
wire _17301_;
wire _17302_;
wire _17303_;
wire _17304_;
wire _17305_;
wire _17306_;
wire _17307_;
wire _17308_;
wire _17309_;
wire _17310_;
wire _17311_;
wire _17312_;
wire _17313_;
wire _17314_;
wire _17315_;
wire _17316_;
wire _17317_;
wire _17318_;
wire _17319_;
wire _17320_;
wire _17321_;
wire _17322_;
wire _17323_;
wire _17324_;
wire _17325_;
wire _17326_;
wire _17327_;
wire _17328_;
wire _17329_;
wire _17330_;
wire _17331_;
wire _17332_;
wire _17333_;
wire _17334_;
wire _17335_;
wire _17336_;
wire _17337_;
wire _17338_;
wire _17339_;
wire _17340_;
wire _17341_;
wire _17342_;
wire _17343_;
wire _17344_;
wire _17345_;
wire _17346_;
wire _17347_;
wire _17348_;
wire _17349_;
wire _17350_;
wire _17351_;
wire _17352_;
wire _17353_;
wire _17354_;
wire _17355_;
wire _17356_;
wire _17357_;
wire _17358_;
wire _17359_;
wire _17360_;
wire _17361_;
wire _17362_;
wire _17363_;
wire _17364_;
wire _17365_;
wire _17366_;
wire _17367_;
wire _17368_;
wire _17369_;
wire _17370_;
wire _17371_;
wire _17372_;
wire _17373_;
wire _17374_;
wire _17375_;
wire _17376_;
wire _17377_;
wire _17378_;
wire _17379_;
wire _17380_;
wire _17381_;
wire _17382_;
wire _17383_;
wire _17384_;
wire _17385_;
wire _17386_;
wire _17387_;
wire _17388_;
wire _17389_;
wire _17390_;
wire _17391_;
wire _17392_;
wire _17393_;
wire _17394_;
wire _17395_;
wire _17396_;
wire _17397_;
wire _17398_;
wire _17399_;
wire _17400_;
wire _17401_;
wire _17402_;
wire _17403_;
wire _17404_;
wire _17405_;
wire _17406_;
wire _17407_;
wire _17408_;
wire _17409_;
wire _17410_;
wire _17411_;
wire _17412_;
wire _17413_;
wire _17414_;
wire _17415_;
wire _17416_;
wire _17417_;
wire _17418_;
wire _17419_;
wire _17420_;
wire _17421_;
wire _17422_;
wire _17423_;
wire _17424_;
wire _17425_;
wire _17426_;
wire _17427_;
wire _17428_;
wire _17429_;
wire _17430_;
wire _17431_;
wire _17432_;
wire _17433_;
wire _17434_;
wire _17435_;
wire _17436_;
wire _17437_;
wire _17438_;
wire _17439_;
wire _17440_;
wire _17441_;
wire _17442_;
wire _17443_;
wire _17444_;
wire _17445_;
wire _17446_;
wire _17447_;
wire _17448_;
wire _17449_;
wire _17450_;
wire _17451_;
wire _17452_;
wire _17453_;
wire _17454_;
wire _17455_;
wire _17456_;
wire _17457_;
wire _17458_;
wire _17459_;
wire _17460_;
wire _17461_;
wire _17462_;
wire _17463_;
wire _17464_;
wire _17465_;
wire _17466_;
wire _17467_;
wire _17468_;
wire _17469_;
wire _17470_;
wire _17471_;
wire _17472_;
wire _17473_;
wire _17474_;
wire _17475_;
wire _17476_;
wire _17477_;
wire _17478_;
wire _17479_;
wire _17480_;
wire _17481_;
wire _17482_;
wire _17483_;
wire _17484_;
wire _17485_;
wire _17486_;
wire _17487_;
wire _17488_;
wire _17489_;
wire _17490_;
wire _17491_;
wire _17492_;
wire _17493_;
wire _17494_;
wire _17495_;
wire _17496_;
wire _17497_;
wire _17498_;
wire _17499_;
wire _17500_;
wire _17501_;
wire _17502_;
wire _17503_;
wire _17504_;
wire _17505_;
wire _17506_;
wire _17507_;
wire _17508_;
wire _17509_;
wire _17510_;
wire _17511_;
wire _17512_;
wire _17513_;
wire _17514_;
wire _17515_;
wire _17516_;
wire _17517_;
wire _17518_;
wire _17519_;
wire _17520_;
wire _17521_;
wire _17522_;
wire _17523_;
wire _17524_;
wire _17525_;
wire _17526_;
wire _17527_;
wire _17528_;
wire _17529_;
wire _17530_;
wire _17531_;
wire _17532_;
wire _17533_;
wire _17534_;
wire _17535_;
wire _17536_;
wire _17537_;
wire _17538_;
wire _17539_;
wire _17540_;
wire _17541_;
wire _17542_;
wire _17543_;
wire _17544_;
wire _17545_;
wire _17546_;
wire _17547_;
wire _17548_;
wire _17549_;
wire _17550_;
wire _17551_;
wire _17552_;
wire _17553_;
wire _17554_;
wire _17555_;
wire _17556_;
wire _17557_;
wire _17558_;
wire _17559_;
wire _17560_;
wire _17561_;
wire _17562_;
wire _17563_;
wire _17564_;
wire _17565_;
wire _17566_;
wire _17567_;
wire _17568_;
wire _17569_;
wire _17570_;
wire _17571_;
wire _17572_;
wire _17573_;
wire _17574_;
wire _17575_;
wire _17576_;
wire _17577_;
wire _17578_;
wire _17579_;
wire _17580_;
wire _17581_;
wire _17582_;
wire _17583_;
wire _17584_;
wire _17585_;
wire _17586_;
wire _17587_;
wire _17588_;
wire _17589_;
wire _17590_;
wire _17591_;
wire _17592_;
wire _17593_;
wire _17594_;
wire _17595_;
wire _17596_;
wire _17597_;
wire _17598_;
wire _17599_;
wire _17600_;
wire _17601_;
wire _17602_;
wire _17603_;
wire _17604_;
wire _17605_;
wire _17606_;
wire _17607_;
wire _17608_;
wire _17609_;
wire _17610_;
wire _17611_;
wire _17612_;
wire _17613_;
wire _17614_;
wire _17615_;
wire _17616_;
wire _17617_;
wire _17618_;
wire _17619_;
wire _17620_;
wire _17621_;
wire _17622_;
wire _17623_;
wire _17624_;
wire _17625_;
wire _17626_;
wire _17627_;
wire _17628_;
wire _17629_;
wire _17630_;
wire _17631_;
wire _17632_;
wire _17633_;
wire _17634_;
wire _17635_;
wire _17636_;
wire _17637_;
wire _17638_;
wire _17639_;
wire _17640_;
wire _17641_;
wire _17642_;
wire _17643_;
wire _17644_;
wire _17645_;
wire _17646_;
wire _17647_;
wire _17648_;
wire _17649_;
wire _17650_;
wire _17651_;
wire _17652_;
wire _17653_;
wire _17654_;
wire _17655_;
wire _17656_;
wire _17657_;
wire _17658_;
wire _17659_;
wire _17660_;
wire _17661_;
wire _17662_;
wire _17663_;
wire _17664_;
wire _17665_;
wire _17666_;
wire _17667_;
wire _17668_;
wire _17669_;
wire _17670_;
wire _17671_;
wire _17672_;
wire _17673_;
wire _17674_;
wire _17675_;
wire _17676_;
wire _17677_;
wire _17678_;
wire _17679_;
wire _17680_;
wire _17681_;
wire _17682_;
wire _17683_;
wire _17684_;
wire _17685_;
wire _17686_;
wire _17687_;
wire _17688_;
wire _17689_;
wire _17690_;
wire _17691_;
wire _17692_;
wire _17693_;
wire _17694_;
wire _17695_;
wire _17696_;
wire _17697_;
wire _17698_;
wire _17699_;
wire _17700_;
wire _17701_;
wire _17702_;
wire _17703_;
wire _17704_;
wire _17705_;
wire _17706_;
wire _17707_;
wire _17708_;
wire _17709_;
wire _17710_;
wire _17711_;
wire _17712_;
wire _17713_;
wire _17714_;
wire _17715_;
wire _17716_;
wire _17717_;
wire _17718_;
wire _17719_;
wire _17720_;
wire _17721_;
wire _17722_;
wire _17723_;
wire _17724_;
wire _17725_;
wire _17726_;
wire _17727_;
wire _17728_;
wire _17729_;
wire _17730_;
wire _17731_;
wire _17732_;
wire _17733_;
wire _17734_;
wire _17735_;
wire _17736_;
wire _17737_;
wire _17738_;
wire _17739_;
wire _17740_;
wire _17741_;
wire _17742_;
wire _17743_;
wire _17744_;
wire _17745_;
wire _17746_;
wire _17747_;
wire _17748_;
wire _17749_;
wire _17750_;
wire _17751_;
wire _17752_;
wire _17753_;
wire _17754_;
wire _17755_;
wire _17756_;
wire _17757_;
wire _17758_;
wire _17759_;
wire _17760_;
wire _17761_;
wire _17762_;
wire _17763_;
wire _17764_;
wire _17765_;
wire _17766_;
wire _17767_;
wire _17768_;
wire _17769_;
wire _17770_;
wire _17771_;
wire _17772_;
wire _17773_;
wire _17774_;
wire _17775_;
wire _17776_;
wire _17777_;
wire _17778_;
wire _17779_;
wire _17780_;
wire _17781_;
wire _17782_;
wire _17783_;
wire _17784_;
wire _17785_;
wire _17786_;
wire _17787_;
wire _17788_;
wire _17789_;
wire _17790_;
wire _17791_;
wire _17792_;
wire _17793_;
wire _17794_;
wire _17795_;
wire _17796_;
wire _17797_;
wire _17798_;
wire _17799_;
wire _17800_;
wire _17801_;
wire _17802_;
wire _17803_;
wire _17804_;
wire _17805_;
wire _17806_;
wire _17807_;
wire _17808_;
wire _17809_;
wire _17810_;
wire _17811_;
wire _17812_;
wire _17813_;
wire _17814_;
wire _17815_;
wire _17816_;
wire _17817_;
wire _17818_;
wire _17819_;
wire _17820_;
wire _17821_;
wire _17822_;
wire _17823_;
wire _17824_;
wire _17825_;
wire _17826_;
wire _17827_;
wire _17828_;
wire _17829_;
wire _17830_;
wire _17831_;
wire _17832_;
wire _17833_;
wire _17834_;
wire _17835_;
wire _17836_;
wire _17837_;
wire _17838_;
wire _17839_;
wire _17840_;
wire _17841_;
wire _17842_;
wire _17843_;
wire _17844_;
wire _17845_;
wire _17846_;
wire _17847_;
wire _17848_;
wire _17849_;
wire _17850_;
wire _17851_;
wire _17852_;
wire _17853_;
wire _17854_;
wire _17855_;
wire _17856_;
wire _17857_;
wire _17858_;
wire _17859_;
wire _17860_;
wire _17861_;
wire _17862_;
wire _17863_;
wire _17864_;
wire _17865_;
wire _17866_;
wire _17867_;
wire _17868_;
wire _17869_;
wire _17870_;
wire _17871_;
wire _17872_;
wire _17873_;
wire _17874_;
wire _17875_;
wire _17876_;
wire _17877_;
wire _17878_;
wire _17879_;
wire _17880_;
wire _17881_;
wire _17882_;
wire _17883_;
wire _17884_;
wire _17885_;
wire _17886_;
wire _17887_;
wire _17888_;
wire _17889_;
wire _17890_;
wire _17891_;
wire _17892_;
wire _17893_;
wire _17894_;
wire _17895_;
wire _17896_;
wire _17897_;
wire _17898_;
wire _17899_;
wire _17900_;
wire _17901_;
wire _17902_;
wire _17903_;
wire _17904_;
wire _17905_;
wire _17906_;
wire _17907_;
wire _17908_;
wire _17909_;
wire _17910_;
wire _17911_;
wire _17912_;
wire _17913_;
wire _17914_;
wire _17915_;
wire _17916_;
wire _17917_;
wire _17918_;
wire _17919_;
wire _17920_;
wire _17921_;
wire _17922_;
wire _17923_;
wire _17924_;
wire _17925_;
wire _17926_;
wire _17927_;
wire _17928_;
wire _17929_;
wire _17930_;
wire _17931_;
wire _17932_;
wire _17933_;
wire _17934_;
wire _17935_;
wire _17936_;
wire _17937_;
wire _17938_;
wire _17939_;
wire _17940_;
wire _17941_;
wire _17942_;
wire _17943_;
wire _17944_;
wire _17945_;
wire _17946_;
wire _17947_;
wire _17948_;
wire _17949_;
wire _17950_;
wire _17951_;
wire _17952_;
wire _17953_;
wire _17954_;
wire _17955_;
wire _17956_;
wire _17957_;
wire _17958_;
wire _17959_;
wire _17960_;
wire _17961_;
wire _17962_;
wire _17963_;
wire _17964_;
wire _17965_;
wire _17966_;
wire _17967_;
wire _17968_;
wire _17969_;
wire _17970_;
wire _17971_;
wire _17972_;
wire _17973_;
wire _17974_;
wire _17975_;
wire _17976_;
wire _17977_;
wire _17978_;
wire _17979_;
wire _17980_;
wire _17981_;
wire _17982_;
wire _17983_;
wire _17984_;
wire _17985_;
wire _17986_;
wire _17987_;
wire _17988_;
wire _17989_;
wire _17990_;
wire _17991_;
wire _17992_;
wire _17993_;
wire _17994_;
wire _17995_;
wire _17996_;
wire _17997_;
wire _17998_;
wire _17999_;
wire _18000_;
wire _18001_;
wire _18002_;
wire _18003_;
wire _18004_;
wire _18005_;
wire _18006_;
wire _18007_;
wire _18008_;
wire _18009_;
wire _18010_;
wire _18011_;
wire _18012_;
wire _18013_;
wire _18014_;
wire _18015_;
wire _18016_;
wire _18017_;
wire _18018_;
wire _18019_;
wire _18020_;
wire _18021_;
wire _18022_;
wire _18023_;
wire _18024_;
wire _18025_;
wire _18026_;
wire _18027_;
wire _18028_;
wire _18029_;
wire _18030_;
wire _18031_;
wire _18032_;
wire _18033_;
wire _18034_;
wire _18035_;
wire _18036_;
wire _18037_;
wire _18038_;
wire _18039_;
wire _18040_;
wire _18041_;
wire _18042_;
wire _18043_;
wire _18044_;
wire _18045_;
wire _18046_;
wire _18047_;
wire _18048_;
wire _18049_;
wire _18050_;
wire _18051_;
wire _18052_;
wire _18053_;
wire _18054_;
wire _18055_;
wire _18056_;
wire _18057_;
wire _18058_;
wire _18059_;
wire _18060_;
wire _18061_;
wire _18062_;
wire _18063_;
wire _18064_;
wire _18065_;
wire _18066_;
wire _18067_;
wire _18068_;
wire _18069_;
wire _18070_;
wire _18071_;
wire _18072_;
wire _18073_;
wire _18074_;
wire _18075_;
wire _18076_;
wire _18077_;
wire _18078_;
wire _18079_;
wire _18080_;
wire _18081_;
wire _18082_;
wire _18083_;
wire _18084_;
wire _18085_;
wire _18086_;
wire _18087_;
wire _18088_;
wire _18089_;
wire _18090_;
wire _18091_;
wire _18092_;
wire _18093_;
wire _18094_;
wire _18095_;
wire _18096_;
wire _18097_;
wire _18098_;
wire _18099_;
wire _18100_;
wire _18101_;
wire _18102_;
wire _18103_;
wire _18104_;
wire _18105_;
wire _18106_;
wire _18107_;
wire _18108_;
wire _18109_;
wire _18110_;
wire _18111_;
wire _18112_;
wire _18113_;
wire _18114_;
wire _18115_;
wire _18116_;
wire _18117_;
wire _18118_;
wire _18119_;
wire _18120_;
wire _18121_;
wire _18122_;
wire _18123_;
wire _18124_;
wire _18125_;
wire _18126_;
wire _18127_;
wire _18128_;
wire _18129_;
wire _18130_;
wire _18131_;
wire _18132_;
wire _18133_;
wire _18134_;
wire _18135_;
wire _18136_;
wire _18137_;
wire _18138_;
wire _18139_;
wire _18140_;
wire _18141_;
wire _18142_;
wire _18143_;
wire _18144_;
wire _18145_;
wire _18146_;
wire _18147_;
wire _18148_;
wire _18149_;
wire _18150_;
wire _18151_;
wire _18152_;
wire _18153_;
wire _18154_;
wire _18155_;
wire _18156_;
wire _18157_;
wire _18158_;
wire _18159_;
wire _18160_;
wire _18161_;
wire _18162_;
wire _18163_;
wire _18164_;
wire _18165_;
wire _18166_;
wire _18167_;
wire _18168_;
wire _18169_;
wire _18170_;
wire _18171_;
wire _18172_;
wire _18173_;
wire _18174_;
wire _18175_;
wire _18176_;
wire _18177_;
wire _18178_;
wire _18179_;
wire _18180_;
wire _18181_;
wire _18182_;
wire _18183_;
wire _18184_;
wire _18185_;
wire _18186_;
wire _18187_;
wire _18188_;
wire _18189_;
wire _18190_;
wire _18191_;
wire _18192_;
wire _18193_;
wire _18194_;
wire _18195_;
wire _18196_;
wire _18197_;
wire _18198_;
wire _18199_;
wire _18200_;
wire _18201_;
wire _18202_;
wire _18203_;
wire _18204_;
wire _18205_;
wire _18206_;
wire _18207_;
wire _18208_;
wire _18209_;
wire _18210_;
wire _18211_;
wire _18212_;
wire _18213_;
wire _18214_;
wire _18215_;
wire _18216_;
wire _18217_;
wire _18218_;
wire _18219_;
wire _18220_;
wire _18221_;
wire _18222_;
wire _18223_;
wire _18224_;
wire _18225_;
wire _18226_;
wire _18227_;
wire _18228_;
wire _18229_;
wire _18230_;
wire _18231_;
wire _18232_;
wire _18233_;
wire _18234_;
wire _18235_;
wire _18236_;
wire _18237_;
wire _18238_;
wire _18239_;
wire _18240_;
wire _18241_;
wire _18242_;
wire _18243_;
wire _18244_;
wire _18245_;
wire _18246_;
wire _18247_;
wire _18248_;
wire _18249_;
wire _18250_;
wire _18251_;
wire _18252_;
wire _18253_;
wire _18254_;
wire _18255_;
wire _18256_;
wire _18257_;
wire _18258_;
wire _18259_;
wire _18260_;
wire _18261_;
wire _18262_;
wire _18263_;
wire _18264_;
wire _18265_;
wire _18266_;
wire _18267_;
wire _18268_;
wire _18269_;
wire _18270_;
wire _18271_;
wire _18272_;
wire _18273_;
wire _18274_;
wire _18275_;
wire _18276_;
wire _18277_;
wire _18278_;
wire _18279_;
wire _18280_;
wire _18281_;
wire _18282_;
wire _18283_;
wire _18284_;
wire _18285_;
wire _18286_;
wire _18287_;
wire _18288_;
wire _18289_;
wire _18290_;
wire _18291_;
wire _18292_;
wire _18293_;
wire _18294_;
wire _18295_;
wire _18296_;
wire _18297_;
wire _18298_;
wire _18299_;
wire _18300_;
wire _18301_;
wire _18302_;
wire _18303_;
wire _18304_;
wire _18305_;
wire _18306_;
wire _18307_;
wire _18308_;
wire _18309_;
wire _18310_;
wire _18311_;
wire _18312_;
wire _18313_;
wire _18314_;
wire _18315_;
wire _18316_;
wire _18317_;
wire _18318_;
wire _18319_;
wire _18320_;
wire _18321_;
wire _18322_;
wire _18323_;
wire _18324_;
wire _18325_;
wire _18326_;
wire _18327_;
wire _18328_;
wire _18329_;
wire _18330_;
wire _18331_;
wire _18332_;
wire _18333_;
wire _18334_;
wire _18335_;
wire _18336_;
wire _18337_;
wire _18338_;
wire _18339_;
wire _18340_;
wire _18341_;
wire _18342_;
wire _18343_;
wire _18344_;
wire _18345_;
wire _18346_;
wire _18347_;
wire _18348_;
wire _18349_;
wire _18350_;
wire _18351_;
wire _18352_;
wire _18353_;
wire _18354_;
wire _18355_;
wire _18356_;
wire _18357_;
wire _18358_;
wire _18359_;
wire _18360_;
wire _18361_;
wire _18362_;
wire _18363_;
wire _18364_;
wire _18365_;
wire _18366_;
wire _18367_;
wire _18368_;
wire _18369_;
wire _18370_;
wire _18371_;
wire _18372_;
wire _18373_;
wire _18374_;
wire _18375_;
wire _18376_;
wire _18377_;
wire _18378_;
wire _18379_;
wire _18380_;
wire _18381_;
wire _18382_;
wire _18383_;
wire _18384_;
wire _18385_;
wire _18386_;
wire _18387_;
wire _18388_;
wire _18389_;
wire _18390_;
wire _18391_;
wire _18392_;
wire _18393_;
wire _18394_;
wire _18395_;
wire _18396_;
wire _18397_;
wire _18398_;
wire _18399_;
wire _18400_;
wire _18401_;
wire _18402_;
wire _18403_;
wire _18404_;
wire _18405_;
wire _18406_;
wire _18407_;
wire _18408_;
wire _18409_;
wire _18410_;
wire _18411_;
wire _18412_;
wire _18413_;
wire _18414_;
wire _18415_;
wire _18416_;
wire _18417_;
wire _18418_;
wire _18419_;
wire _18420_;
wire _18421_;
wire _18422_;
wire _18423_;
wire _18424_;
wire _18425_;
wire _18426_;
wire _18427_;
wire _18428_;
wire _18429_;
wire _18430_;
wire _18431_;
wire _18432_;
wire _18433_;
wire _18434_;
wire _18435_;
wire _18436_;
wire _18437_;
wire _18438_;
wire _18439_;
wire _18440_;
wire _18441_;
wire _18442_;
wire _18443_;
wire _18444_;
wire _18445_;
wire _18446_;
wire _18447_;
wire _18448_;
wire _18449_;
wire _18450_;
wire _18451_;
wire _18452_;
wire _18453_;
wire _18454_;
wire _18455_;
wire _18456_;
wire _18457_;
wire _18458_;
wire _18459_;
wire _18460_;
wire _18461_;
wire _18462_;
wire _18463_;
wire _18464_;
wire _18465_;
wire _18466_;
wire _18467_;
wire _18468_;
wire _18469_;
wire _18470_;
wire _18471_;
wire _18472_;
wire _18473_;
wire _18474_;
wire _18475_;
wire _18476_;
wire _18477_;
wire _18478_;
wire _18479_;
wire _18480_;
wire _18481_;
wire _18482_;
wire _18483_;
wire _18484_;
wire _18485_;
wire _18486_;
wire _18487_;
wire _18488_;
wire _18489_;
wire _18490_;
wire _18491_;
wire _18492_;
wire _18493_;
wire _18494_;
wire _18495_;
wire _18496_;
wire _18497_;
wire _18498_;
wire _18499_;
wire _18500_;
wire _18501_;
wire _18502_;
wire _18503_;
wire _18504_;
wire _18505_;
wire _18506_;
wire _18507_;
wire _18508_;
wire _18509_;
wire _18510_;
wire _18511_;
wire _18512_;
wire _18513_;
wire _18514_;
wire _18515_;
wire _18516_;
wire _18517_;
wire _18518_;
wire _18519_;
wire _18520_;
wire _18521_;
wire _18522_;
wire _18523_;
wire _18524_;
wire _18525_;
wire _18526_;
wire _18527_;
wire _18528_;
wire _18529_;
wire _18530_;
wire _18531_;
wire _18532_;
wire _18533_;
wire _18534_;
wire _18535_;
wire _18536_;
wire _18537_;
wire _18538_;
wire _18539_;
wire _18540_;
wire _18541_;
wire _18542_;
wire _18543_;
wire _18544_;
wire _18545_;
wire _18546_;
wire _18547_;
wire _18548_;
wire _18549_;
wire _18550_;
wire _18551_;
wire _18552_;
wire _18553_;
wire _18554_;
wire _18555_;
wire _18556_;
wire _18557_;
wire _18558_;
wire _18559_;
wire _18560_;
wire _18561_;
wire _18562_;
wire _18563_;
wire _18564_;
wire _18565_;
wire _18566_;
wire _18567_;
wire _18568_;
wire _18569_;
wire _18570_;
wire _18571_;
wire _18572_;
wire _18573_;
wire _18574_;
wire _18575_;
wire _18576_;
wire _18577_;
wire _18578_;
wire _18579_;
wire _18580_;
wire _18581_;
wire _18582_;
wire _18583_;
wire _18584_;
wire _18585_;
wire _18586_;
wire _18587_;
wire _18588_;
wire _18589_;
wire _18590_;
wire _18591_;
wire _18592_;
wire _18593_;
wire _18594_;
wire _18595_;
wire _18596_;
wire _18597_;
wire _18598_;
wire _18599_;
wire _18600_;
wire _18601_;
wire _18602_;
wire _18603_;
wire _18604_;
wire _18605_;
wire _18606_;
wire _18607_;
wire _18608_;
wire _18609_;
wire _18610_;
wire _18611_;
wire _18612_;
wire _18613_;
wire _18614_;
wire _18615_;
wire _18616_;
wire _18617_;
wire _18618_;
wire _18619_;
wire _18620_;
wire _18621_;
wire _18622_;
wire _18623_;
wire _18624_;
wire _18625_;
wire _18626_;
wire _18627_;
wire _18628_;
wire _18629_;
wire _18630_;
wire _18631_;
wire _18632_;
wire _18633_;
wire _18634_;
wire _18635_;
wire _18636_;
wire _18637_;
wire _18638_;
wire _18639_;
wire _18640_;
wire _18641_;
wire _18642_;
wire _18643_;
wire _18644_;
wire _18645_;
wire _18646_;
wire _18647_;
wire _18648_;
wire _18649_;
wire _18650_;
wire _18651_;
wire _18652_;
wire _18653_;
wire _18654_;
wire _18655_;
wire _18656_;
wire _18657_;
wire _18658_;
wire _18659_;
wire _18660_;
wire _18661_;
wire _18662_;
wire _18663_;
wire _18664_;
wire _18665_;
wire _18666_;
wire _18667_;
wire _18668_;
wire _18669_;
wire _18670_;
wire _18671_;
wire _18672_;
wire _18673_;
wire _18674_;
wire _18675_;
wire _18676_;
wire _18677_;
wire _18678_;
wire _18679_;
wire _18680_;
wire _18681_;
wire _18682_;
wire _18683_;
wire _18684_;
wire _18685_;
wire _18686_;
wire _18687_;
wire _18688_;
wire _18689_;
wire _18690_;
wire _18691_;
wire _18692_;
wire _18693_;
wire _18694_;
wire _18695_;
wire _18696_;
wire _18697_;
wire _18698_;
wire _18699_;
wire _18700_;
wire _18701_;
wire _18702_;
wire _18703_;
wire _18704_;
wire _18705_;
wire _18706_;
wire _18707_;
wire _18708_;
wire _18709_;
wire _18710_;
wire _18711_;
wire _18712_;
wire _18713_;
wire _18714_;
wire _18715_;
wire _18716_;
wire _18717_;
wire _18718_;
wire _18719_;
wire _18720_;
wire _18721_;
wire _18722_;
wire _18723_;
wire _18724_;
wire _18725_;
wire _18726_;
wire _18727_;
wire _18728_;
wire _18729_;
wire _18730_;
wire _18731_;
wire _18732_;
wire _18733_;
wire _18734_;
wire _18735_;
wire _18736_;
wire _18737_;
wire _18738_;
wire _18739_;
wire _18740_;
wire _18741_;
wire _18742_;
wire _18743_;
wire _18744_;
wire _18745_;
wire _18746_;
wire _18747_;
wire _18748_;
wire _18749_;
wire _18750_;
wire _18751_;
wire _18752_;
wire _18753_;
wire _18754_;
wire _18755_;
wire _18756_;
wire _18757_;
wire _18758_;
wire _18759_;
wire _18760_;
wire _18761_;
wire _18762_;
wire _18763_;
wire _18764_;
wire _18765_;
wire _18766_;
wire _18767_;
wire _18768_;
wire _18769_;
wire _18770_;
wire _18771_;
wire _18772_;
wire _18773_;
wire _18774_;
wire _18775_;
wire _18776_;
wire _18777_;
wire _18778_;
wire _18779_;
wire _18780_;
wire _18781_;
wire _18782_;
wire _18783_;
wire _18784_;
wire _18785_;
wire _18786_;
wire _18787_;
wire _18788_;
wire _18789_;
wire _18790_;
wire _18791_;
wire _18792_;
wire _18793_;
wire _18794_;
wire _18795_;
wire _18796_;
wire _18797_;
wire _18798_;
wire _18799_;
wire _18800_;
wire _18801_;
wire _18802_;
wire _18803_;
wire _18804_;
wire _18805_;
wire _18806_;
wire _18807_;
wire _18808_;
wire _18809_;
wire _18810_;
wire _18811_;
wire _18812_;
wire _18813_;
wire _18814_;
wire _18815_;
wire _18816_;
wire _18817_;
wire _18818_;
wire _18819_;
wire _18820_;
wire _18821_;
wire _18822_;
wire _18823_;
wire _18824_;
wire _18825_;
wire _18826_;
wire _18827_;
wire _18828_;
wire _18829_;
wire _18830_;
wire _18831_;
wire _18832_;
wire _18833_;
wire _18834_;
wire _18835_;
wire _18836_;
wire _18837_;
wire _18838_;
wire _18839_;
wire _18840_;
wire _18841_;
wire _18842_;
wire _18843_;
wire _18844_;
wire _18845_;
wire _18846_;
wire _18847_;
wire _18848_;
wire _18849_;
wire _18850_;
wire _18851_;
wire _18852_;
wire _18853_;
wire _18854_;
wire _18855_;
wire _18856_;
wire _18857_;
wire _18858_;
wire _18859_;
wire _18860_;
wire _18861_;
wire _18862_;
wire _18863_;
wire _18864_;
wire _18865_;
wire _18866_;
wire _18867_;
wire _18868_;
wire _18869_;
wire _18870_;
wire _18871_;
wire _18872_;
wire _18873_;
wire _18874_;
wire _18875_;
wire _18876_;
wire _18877_;
wire _18878_;
wire _18879_;
wire _18880_;
wire _18881_;
wire _18882_;
wire _18883_;
wire _18884_;
wire _18885_;
wire _18886_;
wire _18887_;
wire _18888_;
wire _18889_;
wire _18890_;
wire _18891_;
wire _18892_;
wire _18893_;
wire _18894_;
wire _18895_;
wire _18896_;
wire _18897_;
wire _18898_;
wire _18899_;
wire _18900_;
wire _18901_;
wire _18902_;
wire _18903_;
wire _18904_;
wire _18905_;
wire _18906_;
wire _18907_;
wire _18908_;
wire _18909_;
wire _18910_;
wire _18911_;
wire _18912_;
wire _18913_;
wire _18914_;
wire _18915_;
wire _18916_;
wire _18917_;
wire _18918_;
wire _18919_;
wire _18920_;
wire _18921_;
wire _18922_;
wire _18923_;
wire _18924_;
wire _18925_;
wire _18926_;
wire _18927_;
wire _18928_;
wire _18929_;
wire _18930_;
wire _18931_;
wire _18932_;
wire _18933_;
wire _18934_;
wire _18935_;
wire _18936_;
wire _18937_;
wire _18938_;
wire _18939_;
wire _18940_;
wire _18941_;
wire _18942_;
wire _18943_;
wire _18944_;
wire _18945_;
wire _18946_;
wire _18947_;
wire _18948_;
wire _18949_;
wire _18950_;
wire _18951_;
wire _18952_;
wire _18953_;
wire _18954_;
wire _18955_;
wire _18956_;
wire _18957_;
wire _18958_;
wire _18959_;
wire _18960_;
wire _18961_;
wire _18962_;
wire _18963_;
wire _18964_;
wire _18965_;
wire _18966_;
wire _18967_;
wire _18968_;
wire _18969_;
wire _18970_;
wire _18971_;
wire _18972_;
wire _18973_;
wire _18974_;
wire _18975_;
wire _18976_;
wire _18977_;
wire _18978_;
wire _18979_;
wire _18980_;
wire _18981_;
wire _18982_;
wire _18983_;
wire _18984_;
wire _18985_;
wire _18986_;
wire _18987_;
wire _18988_;
wire _18989_;
wire _18990_;
wire _18991_;
wire _18992_;
wire _18993_;
wire _18994_;
wire _18995_;
wire _18996_;
wire _18997_;
wire _18998_;
wire _18999_;
wire _19000_;
wire _19001_;
wire _19002_;
wire _19003_;
wire _19004_;
wire _19005_;
wire _19006_;
wire _19007_;
wire _19008_;
wire _19009_;
wire _19010_;
wire _19011_;
wire _19012_;
wire _19013_;
wire _19014_;
wire _19015_;
wire _19016_;
wire _19017_;
wire _19018_;
wire _19019_;
wire _19020_;
wire _19021_;
wire _19022_;
wire _19023_;
wire _19024_;
wire _19025_;
wire _19026_;
wire _19027_;
wire _19028_;
wire _19029_;
wire _19030_;
wire _19031_;
wire _19032_;
wire _19033_;
wire _19034_;
wire _19035_;
wire _19036_;
wire _19037_;
wire _19038_;
wire _19039_;
wire _19040_;
wire _19041_;
wire _19042_;
wire _19043_;
wire _19044_;
wire _19045_;
wire _19046_;
wire _19047_;
wire _19048_;
wire _19049_;
wire _19050_;
wire _19051_;
wire _19052_;
wire _19053_;
wire _19054_;
wire _19055_;
wire _19056_;
wire _19057_;
wire _19058_;
wire _19059_;
wire _19060_;
wire _19061_;
wire _19062_;
wire _19063_;
wire _19064_;
wire _19065_;
wire _19066_;
wire _19067_;
wire _19068_;
wire _19069_;
wire _19070_;
wire _19071_;
wire _19072_;
wire _19073_;
wire _19074_;
wire _19075_;
wire _19076_;
wire _19077_;
wire _19078_;
wire _19079_;
wire _19080_;
wire _19081_;
wire _19082_;
wire _19083_;
wire _19084_;
wire _19085_;
wire _19086_;
wire _19087_;
wire _19088_;
wire _19089_;
wire _19090_;
wire _19091_;
wire _19092_;
wire _19093_;
wire _19094_;
wire _19095_;
wire _19096_;
wire _19097_;
wire _19098_;
wire _19099_;
wire _19100_;
wire _19101_;
wire _19102_;
wire _19103_;
wire _19104_;
wire _19105_;
wire _19106_;
wire _19107_;
wire _19108_;
wire _19109_;
wire _19110_;
wire _19111_;
wire _19112_;
wire _19113_;
wire _19114_;
wire _19115_;
wire _19116_;
wire _19117_;
wire _19118_;
wire _19119_;
wire _19120_;
wire _19121_;
wire _19122_;
wire _19123_;
wire _19124_;
wire _19125_;
wire _19126_;
wire _19127_;
wire _19128_;
wire _19129_;
wire _19130_;
wire _19131_;
wire _19132_;
wire _19133_;
wire _19134_;
wire _19135_;
wire _19136_;
wire _19137_;
wire _19138_;
wire _19139_;
wire _19140_;
wire _19141_;
wire _19142_;
wire _19143_;
wire _19144_;
wire _19145_;
wire _19146_;
wire _19147_;
wire _19148_;
wire _19149_;
wire _19150_;
wire _19151_;
wire _19152_;
wire _19153_;
wire _19154_;
wire _19155_;
wire _19156_;
wire _19157_;
wire _19158_;
wire _19159_;
wire _19160_;
wire _19161_;
wire _19162_;
wire _19163_;
wire _19164_;
wire _19165_;
wire _19166_;
wire _19167_;
wire _19168_;
wire _19169_;
wire _19170_;
wire _19171_;
wire _19172_;
wire _19173_;
wire _19174_;
wire _19175_;
wire _19176_;
wire _19177_;
wire _19178_;
wire _19179_;
wire _19180_;
wire _19181_;
wire _19182_;
wire _19183_;
wire _19184_;
wire _19185_;
wire _19186_;
wire _19187_;
wire _19188_;
wire _19189_;
wire _19190_;
wire _19191_;
wire _19192_;
wire _19193_;
wire _19194_;
wire _19195_;
wire _19196_;
wire _19197_;
wire _19198_;
wire _19199_;
wire _19200_;
wire _19201_;
wire _19202_;
wire _19203_;
wire _19204_;
wire _19205_;
wire _19206_;
wire _19207_;
wire _19208_;
wire _19209_;
wire _19210_;
wire _19211_;
wire _19212_;
wire _19213_;
wire _19214_;
wire _19215_;
wire _19216_;
wire _19217_;
wire _19218_;
wire _19219_;
wire _19220_;
wire _19221_;
wire _19222_;
wire _19223_;
wire _19224_;
wire _19225_;
wire _19226_;
wire _19227_;
wire _19228_;
wire _19229_;
wire _19230_;
wire _19231_;
wire _19232_;
wire _19233_;
wire _19234_;
wire _19235_;
wire _19236_;
wire _19237_;
wire _19238_;
wire _19239_;
wire _19240_;
wire _19241_;
wire _19242_;
wire _19243_;
wire _19244_;
wire _19245_;
wire _19246_;
wire _19247_;
wire _19248_;
wire _19249_;
wire _19250_;
wire _19251_;
wire _19252_;
wire _19253_;
wire _19254_;
wire _19255_;
wire _19256_;
wire _19257_;
wire _19258_;
wire _19259_;
wire _19260_;
wire _19261_;
wire _19262_;
wire _19263_;
wire _19264_;
wire _19265_;
wire _19266_;
wire _19267_;
wire _19268_;
wire _19269_;
wire _19270_;
wire _19271_;
wire _19272_;
wire _19273_;
wire _19274_;
wire _19275_;
wire _19276_;
wire _19277_;
wire _19278_;
wire _19279_;
wire _19280_;
wire _19281_;
wire _19282_;
wire _19283_;
wire _19284_;
wire _19285_;
wire _19286_;
wire _19287_;
wire _19288_;
wire _19289_;
wire _19290_;
wire _19291_;
wire _19292_;
wire _19293_;
wire _19294_;
wire _19295_;
wire _19296_;
wire _19297_;
wire _19298_;
wire _19299_;
wire _19300_;
wire _19301_;
wire _19302_;
wire _19303_;
wire _19304_;
wire _19305_;
wire _19306_;
wire _19307_;
wire _19308_;
wire _19309_;
wire _19310_;
wire _19311_;
wire _19312_;
wire _19313_;
wire _19314_;
wire _19315_;
wire _19316_;
wire _19317_;
wire _19318_;
wire _19319_;
wire _19320_;
wire _19321_;
wire _19322_;
wire _19323_;
wire _19324_;
wire _19325_;
wire _19326_;
wire _19327_;
wire _19328_;
wire _19329_;
wire _19330_;
wire _19331_;
wire _19332_;
wire _19333_;
wire _19334_;
wire _19335_;
wire _19336_;
wire _19337_;
wire _19338_;
wire _19339_;
wire _19340_;
wire _19341_;
wire _19342_;
wire _19343_;
wire _19344_;
wire _19345_;
wire _19346_;
wire _19347_;
wire _19348_;
wire _19349_;
wire _19350_;
wire _19351_;
wire _19352_;
wire _19353_;
wire _19354_;
wire _19355_;
wire _19356_;
wire _19357_;
wire _19358_;
wire _19359_;
wire _19360_;
wire _19361_;
wire _19362_;
wire _19363_;
wire _19364_;
wire _19365_;
wire _19366_;
wire _19367_;
wire _19368_;
wire _19369_;
wire _19370_;
wire _19371_;
wire _19372_;
wire _19373_;
wire _19374_;
wire _19375_;
wire _19376_;
wire _19377_;
wire _19378_;
wire _19379_;
wire _19380_;
wire _19381_;
wire _19382_;
wire _19383_;
wire _19384_;
wire _19385_;
wire _19386_;
wire _19387_;
wire _19388_;
wire _19389_;
wire _19390_;
wire _19391_;
wire _19392_;
wire _19393_;
wire _19394_;
wire _19395_;
wire _19396_;
wire _19397_;
wire _19398_;
wire _19399_;
wire _19400_;
wire _19401_;
wire _19402_;
wire _19403_;
wire _19404_;
wire _19405_;
wire _19406_;
wire _19407_;
wire _19408_;
wire _19409_;
wire _19410_;
wire _19411_;
wire _19412_;
wire _19413_;
wire _19414_;
wire _19415_;
wire _19416_;
wire _19417_;
wire _19418_;
wire _19419_;
wire _19420_;
wire _19421_;
wire _19422_;
wire _19423_;
wire _19424_;
wire _19425_;
wire _19426_;
wire _19427_;
wire _19428_;
wire _19429_;
wire _19430_;
wire _19431_;
wire _19432_;
wire _19433_;
wire _19434_;
wire _19435_;
wire _19436_;
wire _19437_;
wire _19438_;
wire _19439_;
wire _19440_;
wire _19441_;
wire _19442_;
wire _19443_;
wire _19444_;
wire _19445_;
wire _19446_;
wire _19447_;
wire _19448_;
wire _19449_;
wire _19450_;
wire _19451_;
wire _19452_;
wire _19453_;
wire _19454_;
wire _19455_;
wire _19456_;
wire _19457_;
wire _19458_;
wire _19459_;
wire _19460_;
wire _19461_;
wire _19462_;
wire _19463_;
wire _19464_;
wire _19465_;
wire _19466_;
wire _19467_;
wire _19468_;
wire _19469_;
wire _19470_;
wire _19471_;
wire _19472_;
wire _19473_;
wire _19474_;
wire _19475_;
wire _19476_;
wire _19477_;
wire _19478_;
wire _19479_;
wire _19480_;
wire _19481_;
wire _19482_;
wire _19483_;
wire _19484_;
wire _19485_;
wire _19486_;
wire _19487_;
wire _19488_;
wire _19489_;
wire _19490_;
wire _19491_;
wire _19492_;
wire _19493_;
wire _19494_;
wire _19495_;
wire _19496_;
wire _19497_;
wire _19498_;
wire _19499_;
wire _19500_;
wire _19501_;
wire _19502_;
wire _19503_;
wire _19504_;
wire _19505_;
wire _19506_;
wire _19507_;
wire _19508_;
wire _19509_;
wire _19510_;
wire _19511_;
wire _19512_;
wire _19513_;
wire _19514_;
wire _19515_;
wire _19516_;
wire _19517_;
wire _19518_;
wire _19519_;
wire _19520_;
wire _19521_;
wire _19522_;
wire _19523_;
wire _19524_;
wire _19525_;
wire _19526_;
wire _19527_;
wire _19528_;
wire _19529_;
wire _19530_;
wire _19531_;
wire _19532_;
wire _19533_;
wire _19534_;
wire _19535_;
wire _19536_;
wire _19537_;
wire _19538_;
wire _19539_;
wire _19540_;
wire _19541_;
wire _19542_;
wire _19543_;
wire _19544_;
wire _19545_;
wire _19546_;
wire _19547_;
wire _19548_;
wire _19549_;
wire _19550_;
wire _19551_;
wire _19552_;
wire _19553_;
wire _19554_;
wire _19555_;
wire _19556_;
wire _19557_;
wire _19558_;
wire _19559_;
wire _19560_;
wire _19561_;
wire _19562_;
wire _19563_;
wire _19564_;
wire _19565_;
wire _19566_;
wire _19567_;
wire _19568_;
wire _19569_;
wire _19570_;
wire _19571_;
wire _19572_;
wire _19573_;
wire _19574_;
wire _19575_;
wire _19576_;
wire _19577_;
wire _19578_;
wire _19579_;
wire _19580_;
wire _19581_;
wire _19582_;
wire _19583_;
wire _19584_;
wire _19585_;
wire _19586_;
wire _19587_;
wire _19588_;
wire _19589_;
wire _19590_;
wire _19591_;
wire _19592_;
wire _19593_;
wire _19594_;
wire _19595_;
wire _19596_;
wire _19597_;
wire _19598_;
wire _19599_;
wire _19600_;
wire _19601_;
wire _19602_;
wire _19603_;
wire _19604_;
wire _19605_;
wire _19606_;
wire _19607_;
wire _19608_;
wire _19609_;
wire _19610_;
wire _19611_;
wire _19612_;
wire _19613_;
wire _19614_;
wire _19615_;
wire _19616_;
wire _19617_;
wire _19618_;
wire _19619_;
wire _19620_;
wire _19621_;
wire _19622_;
wire _19623_;
wire _19624_;
wire _19625_;
wire _19626_;
wire _19627_;
wire _19628_;
wire _19629_;
wire _19630_;
wire _19631_;
wire _19632_;
wire _19633_;
wire _19634_;
wire _19635_;
wire _19636_;
wire _19637_;
wire _19638_;
wire _19639_;
wire _19640_;
wire _19641_;
wire _19642_;
wire _19643_;
wire _19644_;
wire _19645_;
wire _19646_;
wire _19647_;
wire _19648_;
wire _19649_;
wire _19650_;
wire _19651_;
wire _19652_;
wire _19653_;
wire _19654_;
wire _19655_;
wire _19656_;
wire _19657_;
wire _19658_;
wire _19659_;
wire _19660_;
wire _19661_;
wire _19662_;
wire _19663_;
wire _19664_;
wire _19665_;
wire _19666_;
wire _19667_;
wire _19668_;
wire _19669_;
wire _19670_;
wire _19671_;
wire _19672_;
wire _19673_;
wire _19674_;
wire _19675_;
wire _19676_;
wire _19677_;
wire _19678_;
wire _19679_;
wire _19680_;
wire _19681_;
wire _19682_;
wire _19683_;
wire _19684_;
wire _19685_;
wire _19686_;
wire _19687_;
wire _19688_;
wire _19689_;
wire _19690_;
wire _19691_;
wire _19692_;
wire _19693_;
wire _19694_;
wire _19695_;
wire _19696_;
wire _19697_;
wire _19698_;
wire _19699_;
wire _19700_;
wire _19701_;
wire _19702_;
wire _19703_;
wire _19704_;
wire _19705_;
wire _19706_;
wire _19707_;
wire _19708_;
wire _19709_;
wire _19710_;
wire _19711_;
wire _19712_;
wire _19713_;
wire _19714_;
wire _19715_;
wire _19716_;
wire _19717_;
wire _19718_;
wire _19719_;
wire _19720_;
wire _19721_;
wire _19722_;
wire _19723_;
wire _19724_;
wire _19725_;
wire _19726_;
wire _19727_;
wire _19728_;
wire _19729_;
wire _19730_;
wire _19731_;
wire _19732_;
wire _19733_;
wire _19734_;
wire _19735_;
wire _19736_;
wire _19737_;
wire _19738_;
wire _19739_;
wire _19740_;
wire _19741_;
wire _19742_;
wire _19743_;
wire _19744_;
wire _19745_;
wire _19746_;
wire _19747_;
wire _19748_;
wire _19749_;
wire _19750_;
wire _19751_;
wire _19752_;
wire _19753_;
wire _19754_;
wire _19755_;
wire _19756_;
wire _19757_;
wire _19758_;
wire _19759_;
wire _19760_;
wire _19761_;
wire _19762_;
wire _19763_;
wire _19764_;
wire _19765_;
wire _19766_;
wire _19767_;
wire _19768_;
wire _19769_;
wire _19770_;
wire _19771_;
wire _19772_;
wire _19773_;
wire _19774_;
wire _19775_;
wire _19776_;
wire _19777_;
wire _19778_;
wire _19779_;
wire _19780_;
wire _19781_;
wire _19782_;
wire _19783_;
wire _19784_;
wire _19785_;
wire _19786_;
wire _19787_;
wire _19788_;
wire _19789_;
wire _19790_;
wire _19791_;
wire _19792_;
wire _19793_;
wire _19794_;
wire _19795_;
wire _19796_;
wire _19797_;
wire _19798_;
wire _19799_;
wire _19800_;
wire _19801_;
wire _19802_;
wire _19803_;
wire _19804_;
wire _19805_;
wire _19806_;
wire _19807_;
wire _19808_;
wire _19809_;
wire _19810_;
wire _19811_;
wire _19812_;
wire _19813_;
wire _19814_;
wire _19815_;
wire _19816_;
wire _19817_;
wire _19818_;
wire _19819_;
wire _19820_;
wire _19821_;
wire _19822_;
wire _19823_;
wire _19824_;
wire _19825_;
wire _19826_;
wire _19827_;
wire _19828_;
wire _19829_;
wire _19830_;
wire _19831_;
wire _19832_;
wire _19833_;
wire _19834_;
wire _19835_;
wire _19836_;
wire _19837_;
wire _19838_;
wire _19839_;
wire _19840_;
wire _19841_;
wire _19842_;
wire _19843_;
wire _19844_;
wire _19845_;
wire _19846_;
wire _19847_;
wire _19848_;
wire _19849_;
wire _19850_;
wire _19851_;
wire _19852_;
wire _19853_;
wire _19854_;
wire _19855_;
wire _19856_;
wire _19857_;
wire _19858_;
wire _19859_;
wire _19860_;
wire _19861_;
wire _19862_;
wire _19863_;
wire _19864_;
wire _19865_;
wire _19866_;
wire _19867_;
wire _19868_;
wire _19869_;
wire _19870_;
wire _19871_;
wire _19872_;
wire _19873_;
wire _19874_;
wire _19875_;
wire _19876_;
wire _19877_;
wire _19878_;
wire _19879_;
wire _19880_;
wire _19881_;
wire _19882_;
wire _19883_;
wire _19884_;
wire _19885_;
wire _19886_;
wire _19887_;
wire _19888_;
wire _19889_;
wire _19890_;
wire _19891_;
wire _19892_;
wire _19893_;
wire _19894_;
wire _19895_;
wire _19896_;
wire _19897_;
wire _19898_;
wire _19899_;
wire _19900_;
wire _19901_;
wire _19902_;
wire _19903_;
wire _19904_;
wire _19905_;
wire _19906_;
wire _19907_;
wire _19908_;
wire _19909_;
wire _19910_;
wire _19911_;
wire _19912_;
wire _19913_;
wire _19914_;
wire _19915_;
wire _19916_;
wire _19917_;
wire _19918_;
wire _19919_;
wire _19920_;
wire _19921_;
wire _19922_;
wire _19923_;
wire _19924_;
wire _19925_;
wire _19926_;
wire _19927_;
wire _19928_;
wire _19929_;
wire _19930_;
wire _19931_;
wire _19932_;
wire _19933_;
wire _19934_;
wire _19935_;
wire _19936_;
wire _19937_;
wire _19938_;
wire _19939_;
wire _19940_;
wire _19941_;
wire _19942_;
wire _19943_;
wire _19944_;
wire _19945_;
wire _19946_;
wire _19947_;
wire _19948_;
wire _19949_;
wire _19950_;
wire _19951_;
wire _19952_;
wire _19953_;
wire _19954_;
wire _19955_;
wire _19956_;
wire _19957_;
wire _19958_;
wire _19959_;
wire _19960_;
wire _19961_;
wire _19962_;
wire _19963_;
wire _19964_;
wire _19965_;
wire _19966_;
wire _19967_;
wire _19968_;
wire _19969_;
wire _19970_;
wire _19971_;
wire _19972_;
wire _19973_;
wire _19974_;
wire _19975_;
wire _19976_;
wire _19977_;
wire _19978_;
wire _19979_;
wire _19980_;
wire _19981_;
wire _19982_;
wire _19983_;
wire _19984_;
wire _19985_;
wire _19986_;
wire _19987_;
wire _19988_;
wire _19989_;
wire _19990_;
wire _19991_;
wire _19992_;
wire _19993_;
wire _19994_;
wire _19995_;
wire _19996_;
wire _19997_;
wire _19998_;
wire _19999_;
wire _20000_;
wire _20001_;
wire _20002_;
wire _20003_;
wire _20004_;
wire _20005_;
wire _20006_;
wire _20007_;
wire _20008_;
wire _20009_;
wire _20010_;
wire _20011_;
wire _20012_;
wire _20013_;
wire _20014_;
wire _20015_;
wire _20016_;
wire _20017_;
wire _20018_;
wire _20019_;
wire _20020_;
wire _20021_;
wire _20022_;
wire _20023_;
wire _20024_;
wire _20025_;
wire _20026_;
wire _20027_;
wire _20028_;
wire _20029_;
wire _20030_;
wire _20031_;
wire _20032_;
wire _20033_;
wire _20034_;
wire _20035_;
wire _20036_;
wire _20037_;
wire _20038_;
wire _20039_;
wire _20040_;
wire _20041_;
wire _20042_;
wire _20043_;
wire _20044_;
wire _20045_;
wire _20046_;
wire _20047_;
wire _20048_;
wire _20049_;
wire _20050_;
wire _20051_;
wire _20052_;
wire _20053_;
wire _20054_;
wire _20055_;
wire _20056_;
wire _20057_;
wire _20058_;
wire _20059_;
wire _20060_;
wire _20061_;
wire _20062_;
wire _20063_;
wire _20064_;
wire _20065_;
wire _20066_;
wire _20067_;
wire _20068_;
wire _20069_;
wire _20070_;
wire _20071_;
wire _20072_;
wire _20073_;
wire _20074_;
wire _20075_;
wire _20076_;
wire _20077_;
wire _20078_;
wire _20079_;
wire _20080_;
wire _20081_;
wire _20082_;
wire _20083_;
wire _20084_;
wire _20085_;
wire _20086_;
wire _20087_;
wire _20088_;
wire _20089_;
wire _20090_;
wire _20091_;
wire _20092_;
wire _20093_;
wire _20094_;
wire _20095_;
wire _20096_;
wire _20097_;
wire _20098_;
wire _20099_;
wire _20100_;
wire _20101_;
wire _20102_;
wire _20103_;
wire _20104_;
wire _20105_;
wire _20106_;
wire _20107_;
wire _20108_;
wire _20109_;
wire _20110_;
wire _20111_;
wire _20112_;
wire _20113_;
wire _20114_;
wire _20115_;
wire _20116_;
wire _20117_;
wire _20118_;
wire _20119_;
wire _20120_;
wire _20121_;
wire _20122_;
wire _20123_;
wire _20124_;
wire _20125_;
wire _20126_;
wire _20127_;
wire _20128_;
wire _20129_;
wire _20130_;
wire _20131_;
wire _20132_;
wire _20133_;
wire _20134_;
wire _20135_;
wire _20136_;
wire _20137_;
wire _20138_;
wire _20139_;
wire _20140_;
wire _20141_;
wire _20142_;
wire _20143_;
wire _20144_;
wire _20145_;
wire _20146_;
wire _20147_;
wire _20148_;
wire _20149_;
wire _20150_;
wire _20151_;
wire _20152_;
wire _20153_;
wire _20154_;
wire _20155_;
wire _20156_;
wire _20157_;
wire _20158_;
wire _20159_;
wire _20160_;
wire _20161_;
wire _20162_;
wire _20163_;
wire _20164_;
wire _20165_;
wire _20166_;
wire _20167_;
wire _20168_;
wire _20169_;
wire _20170_;
wire _20171_;
wire _20172_;
wire _20173_;
wire _20174_;
wire _20175_;
wire _20176_;
wire _20177_;
wire _20178_;
wire _20179_;
wire _20180_;
wire _20181_;
wire _20182_;
wire _20183_;
wire _20184_;
wire _20185_;
wire _20186_;
wire _20187_;
wire _20188_;
wire _20189_;
wire _20190_;
wire _20191_;
wire _20192_;
wire _20193_;
wire _20194_;
wire _20195_;
wire _20196_;
wire _20197_;
wire _20198_;
wire _20199_;
wire _20200_;
wire _20201_;
wire _20202_;
wire _20203_;
wire _20204_;
wire _20205_;
wire _20206_;
wire _20207_;
wire _20208_;
wire _20209_;
wire _20210_;
wire _20211_;
wire _20212_;
wire _20213_;
wire _20214_;
wire _20215_;
wire _20216_;
wire _20217_;
wire _20218_;
wire _20219_;
wire _20220_;
wire _20221_;
wire _20222_;
wire _20223_;
wire _20224_;
wire _20225_;
wire _20226_;
wire _20227_;
wire _20228_;
wire _20229_;
wire _20230_;
wire _20231_;
wire _20232_;
wire _20233_;
wire _20234_;
wire _20235_;
wire _20236_;
wire _20237_;
wire _20238_;
wire _20239_;
wire _20240_;
wire _20241_;
wire _20242_;
wire _20243_;
wire _20244_;
wire _20245_;
wire _20246_;
wire _20247_;
wire _20248_;
wire _20249_;
wire _20250_;
wire _20251_;
wire _20252_;
wire _20253_;
wire _20254_;
wire _20255_;
wire _20256_;
wire _20257_;
wire _20258_;
wire _20259_;
wire _20260_;
wire _20261_;
wire _20262_;
wire _20263_;
wire _20264_;
wire _20265_;
wire _20266_;
wire _20267_;
wire _20268_;
wire _20269_;
wire _20270_;
wire _20271_;
wire _20272_;
wire _20273_;
wire _20274_;
wire _20275_;
wire _20276_;
wire _20277_;
wire _20278_;
wire _20279_;
wire _20280_;
wire _20281_;
wire _20282_;
wire _20283_;
wire _20284_;
wire _20285_;
wire _20286_;
wire _20287_;
wire _20288_;
wire _20289_;
wire _20290_;
wire _20291_;
wire _20292_;
wire _20293_;
wire _20294_;
wire _20295_;
wire _20296_;
wire _20297_;
wire _20298_;
wire _20299_;
wire _20300_;
wire _20301_;
wire _20302_;
wire _20303_;
wire _20304_;
wire _20305_;
wire _20306_;
wire _20307_;
wire _20308_;
wire _20309_;
wire _20310_;
wire _20311_;
wire _20312_;
wire _20313_;
wire _20314_;
wire _20315_;
wire _20316_;
wire _20317_;
wire _20318_;
wire _20319_;
wire _20320_;
wire _20321_;
wire _20322_;
wire _20323_;
wire _20324_;
wire _20325_;
wire _20326_;
wire _20327_;
wire _20328_;
wire _20329_;
wire _20330_;
wire _20331_;
wire _20332_;
wire _20333_;
wire _20334_;
wire _20335_;
wire _20336_;
wire _20337_;
wire _20338_;
wire _20339_;
wire _20340_;
wire _20341_;
wire _20342_;
wire _20343_;
wire _20344_;
wire _20345_;
wire _20346_;
wire _20347_;
wire _20348_;
wire _20349_;
wire _20350_;
wire _20351_;
wire _20352_;
wire _20353_;
wire _20354_;
wire _20355_;
wire _20356_;
wire _20357_;
wire _20358_;
wire _20359_;
wire _20360_;
wire _20361_;
wire _20362_;
wire _20363_;
wire _20364_;
wire _20365_;
wire _20366_;
wire _20367_;
wire _20368_;
wire _20369_;
wire _20370_;
wire _20371_;
wire _20372_;
wire _20373_;
wire _20374_;
wire _20375_;
wire _20376_;
wire _20377_;
wire _20378_;
wire _20379_;
wire _20380_;
wire _20381_;
wire _20382_;
wire _20383_;
wire _20384_;
wire _20385_;
wire _20386_;
wire _20387_;
wire _20388_;
wire _20389_;
wire _20390_;
wire _20391_;
wire _20392_;
wire _20393_;
wire _20394_;
wire _20395_;
wire _20396_;
wire _20397_;
wire _20398_;
wire _20399_;
wire _20400_;
wire _20401_;
wire _20402_;
wire _20403_;
wire _20404_;
wire _20405_;
wire _20406_;
wire _20407_;
wire _20408_;
wire _20409_;
wire _20410_;
wire _20411_;
wire _20412_;
wire _20413_;
wire _20414_;
wire _20415_;
wire _20416_;
wire _20417_;
wire _20418_;
wire _20419_;
wire _20420_;
wire _20421_;
wire _20422_;
wire _20423_;
wire _20424_;
wire _20425_;
wire _20426_;
wire _20427_;
wire _20428_;
wire _20429_;
wire _20430_;
wire _20431_;
wire _20432_;
wire _20433_;
wire _20434_;
wire _20435_;
wire _20436_;
wire _20437_;
wire _20438_;
wire _20439_;
wire _20440_;
wire _20441_;
wire _20442_;
wire _20443_;
wire _20444_;
wire _20445_;
wire _20446_;
wire _20447_;
wire _20448_;
wire _20449_;
wire _20450_;
wire _20451_;
wire _20452_;
wire _20453_;
wire _20454_;
wire _20455_;
wire _20456_;
wire _20457_;
wire _20458_;
wire _20459_;
wire _20460_;
wire _20461_;
wire _20462_;
wire _20463_;
wire _20464_;
wire _20465_;
wire _20466_;
wire _20467_;
wire _20468_;
wire _20469_;
wire _20470_;
wire _20471_;
wire _20472_;
wire _20473_;
wire _20474_;
wire _20475_;
wire _20476_;
wire _20477_;
wire _20478_;
wire _20479_;
wire _20480_;
wire _20481_;
wire _20482_;
wire _20483_;
wire _20484_;
wire _20485_;
wire _20486_;
wire _20487_;
wire _20488_;
wire _20489_;
wire _20490_;
wire _20491_;
wire _20492_;
wire _20493_;
wire _20494_;
wire _20495_;
wire _20496_;
wire _20497_;
wire _20498_;
wire _20499_;
wire _20500_;
wire _20501_;
wire _20502_;
wire _20503_;
wire _20504_;
wire _20505_;
wire _20506_;
wire _20507_;
wire _20508_;
wire _20509_;
wire _20510_;
wire _20511_;
wire _20512_;
wire _20513_;
wire _20514_;
wire _20515_;
wire _20516_;
wire _20517_;
wire _20518_;
wire _20519_;
wire _20520_;
wire _20521_;
wire _20522_;
wire _20523_;
wire _20524_;
wire _20525_;
wire _20526_;
wire _20527_;
wire _20528_;
wire _20529_;
wire _20530_;
wire _20531_;
wire _20532_;
wire _20533_;
wire _20534_;
wire _20535_;
wire _20536_;
wire _20537_;
wire _20538_;
wire _20539_;
wire _20540_;
wire _20541_;
wire _20542_;
wire _20543_;
wire _20544_;
wire _20545_;
wire _20546_;
wire _20547_;
wire _20548_;
wire _20549_;
wire _20550_;
wire _20551_;
wire _20552_;
wire _20553_;
wire _20554_;
wire _20555_;
wire _20556_;
wire _20557_;
wire _20558_;
wire _20559_;
wire _20560_;
wire _20561_;
wire _20562_;
wire _20563_;
wire _20564_;
wire _20565_;
wire _20566_;
wire _20567_;
wire _20568_;
wire _20569_;
wire _20570_;
wire _20571_;
wire _20572_;
wire _20573_;
wire _20574_;
wire _20575_;
wire _20576_;
wire _20577_;
wire _20578_;
wire _20579_;
wire _20580_;
wire _20581_;
wire _20582_;
wire _20583_;
wire _20584_;
wire _20585_;
wire _20586_;
wire _20587_;
wire _20588_;
wire _20589_;
wire _20590_;
wire _20591_;
wire _20592_;
wire _20593_;
wire _20594_;
wire _20595_;
wire _20596_;
wire _20597_;
wire _20598_;
wire _20599_;
wire _20600_;
wire _20601_;
wire _20602_;
wire _20603_;
wire _20604_;
wire _20605_;
wire _20606_;
wire _20607_;
wire _20608_;
wire _20609_;
wire _20610_;
wire _20611_;
wire _20612_;
wire _20613_;
wire _20614_;
wire _20615_;
wire _20616_;
wire _20617_;
wire _20618_;
wire _20619_;
wire _20620_;
wire _20621_;
wire _20622_;
wire _20623_;
wire _20624_;
wire _20625_;
wire _20626_;
wire _20627_;
wire _20628_;
wire _20629_;
wire _20630_;
wire _20631_;
wire _20632_;
wire _20633_;
wire _20634_;
wire _20635_;
wire _20636_;
wire _20637_;
wire _20638_;
wire _20639_;
wire _20640_;
wire _20641_;
wire _20642_;
wire _20643_;
wire _20644_;
wire _20645_;
wire _20646_;
wire _20647_;
wire _20648_;
wire _20649_;
wire _20650_;
wire _20651_;
wire _20652_;
wire _20653_;
wire _20654_;
wire _20655_;
wire _20656_;
wire _20657_;
wire _20658_;
wire _20659_;
wire _20660_;
wire _20661_;
wire _20662_;
wire _20663_;
wire _20664_;
wire _20665_;
wire _20666_;
wire _20667_;
wire _20668_;
wire _20669_;
wire _20670_;
wire _20671_;
wire _20672_;
wire _20673_;
wire _20674_;
wire _20675_;
wire _20676_;
wire _20677_;
wire _20678_;
wire _20679_;
wire _20680_;
wire _20681_;
wire _20682_;
wire _20683_;
wire _20684_;
wire _20685_;
wire _20686_;
wire _20687_;
wire _20688_;
wire _20689_;
wire _20690_;
wire _20691_;
wire _20692_;
wire _20693_;
wire _20694_;
wire _20695_;
wire _20696_;
wire _20697_;
wire _20698_;
wire _20699_;
wire _20700_;
wire _20701_;
wire _20702_;
wire _20703_;
wire _20704_;
wire _20705_;
wire _20706_;
wire _20707_;
wire _20708_;
wire _20709_;
wire _20710_;
wire _20711_;
wire _20712_;
wire _20713_;
wire _20714_;
wire _20715_;
wire _20716_;
wire _20717_;
wire _20718_;
wire _20719_;
wire _20720_;
wire _20721_;
wire _20722_;
wire _20723_;
wire _20724_;
wire _20725_;
wire _20726_;
wire _20727_;
wire _20728_;
wire _20729_;
wire _20730_;
wire _20731_;
wire _20732_;
wire _20733_;
wire _20734_;
wire _20735_;
wire _20736_;
wire _20737_;
wire _20738_;
wire _20739_;
wire _20740_;
wire _20741_;
wire _20742_;
wire _20743_;
wire _20744_;
wire _20745_;
wire _20746_;
wire _20747_;
wire _20748_;
wire _20749_;
wire _20750_;
wire _20751_;
wire _20752_;
wire _20753_;
wire _20754_;
wire _20755_;
wire _20756_;
wire _20757_;
wire _20758_;
wire _20759_;
wire _20760_;
wire _20761_;
wire _20762_;
wire _20763_;
wire _20764_;
wire _20765_;
wire _20766_;
wire _20767_;
wire _20768_;
wire _20769_;
wire _20770_;
wire _20771_;
wire _20772_;
wire _20773_;
wire _20774_;
wire _20775_;
wire _20776_;
wire _20777_;
wire _20778_;
wire _20779_;
wire _20780_;
wire _20781_;
wire _20782_;
wire _20783_;
wire _20784_;
wire _20785_;
wire _20786_;
wire _20787_;
wire _20788_;
wire _20789_;
wire _20790_;
wire _20791_;
wire _20792_;
wire _20793_;
wire _20794_;
wire _20795_;
wire _20796_;
wire _20797_;
wire _20798_;
wire _20799_;
wire _20800_;
wire _20801_;
wire _20802_;
wire _20803_;
wire _20804_;
wire _20805_;
wire _20806_;
wire _20807_;
wire _20808_;
wire _20809_;
wire _20810_;
wire _20811_;
wire _20812_;
wire _20813_;
wire _20814_;
wire _20815_;
wire _20816_;
wire _20817_;
wire _20818_;
wire _20819_;
wire _20820_;
wire _20821_;
wire _20822_;
wire _20823_;
wire _20824_;
wire _20825_;
wire _20826_;
wire _20827_;
wire _20828_;
wire _20829_;
wire _20830_;
wire _20831_;
wire _20832_;
wire _20833_;
wire _20834_;
wire _20835_;
wire _20836_;
wire _20837_;
wire _20838_;
wire _20839_;
wire _20840_;
wire _20841_;
wire _20842_;
wire _20843_;
wire _20844_;
wire _20845_;
wire _20846_;
wire _20847_;
wire _20848_;
wire _20849_;
wire _20850_;
wire _20851_;
wire _20852_;
wire _20853_;
wire _20854_;
wire _20855_;
wire _20856_;
wire _20857_;
wire _20858_;
wire _20859_;
wire _20860_;
wire _20861_;
wire _20862_;
wire _20863_;
wire _20864_;
wire _20865_;
wire _20866_;
wire _20867_;
wire _20868_;
wire _20869_;
wire _20870_;
wire _20871_;
wire _20872_;
wire _20873_;
wire _20874_;
wire _20875_;
wire _20876_;
wire _20877_;
wire _20878_;
wire _20879_;
wire _20880_;
wire _20881_;
wire _20882_;
wire _20883_;
wire _20884_;
wire _20885_;
wire _20886_;
wire _20887_;
wire _20888_;
wire _20889_;
wire _20890_;
wire _20891_;
wire _20892_;
wire _20893_;
wire _20894_;
wire _20895_;
wire _20896_;
wire _20897_;
wire _20898_;
wire _20899_;
wire _20900_;
wire _20901_;
wire _20902_;
wire _20903_;
wire _20904_;
wire _20905_;
wire _20906_;
wire _20907_;
wire _20908_;
wire _20909_;
wire _20910_;
wire _20911_;
wire _20912_;
wire _20913_;
wire _20914_;
wire _20915_;
wire _20916_;
wire _20917_;
wire _20918_;
wire _20919_;
wire _20920_;
wire _20921_;
wire _20922_;
wire _20923_;
wire _20924_;
wire _20925_;
wire _20926_;
wire _20927_;
wire _20928_;
wire _20929_;
wire _20930_;
wire _20931_;
wire _20932_;
wire _20933_;
wire _20934_;
wire _20935_;
wire _20936_;
wire _20937_;
wire _20938_;
wire _20939_;
wire _20940_;
wire _20941_;
wire _20942_;
wire _20943_;
wire _20944_;
wire _20945_;
wire _20946_;
wire _20947_;
wire _20948_;
wire _20949_;
wire _20950_;
wire _20951_;
wire _20952_;
wire _20953_;
wire _20954_;
wire _20955_;
wire _20956_;
wire _20957_;
wire _20958_;
wire _20959_;
wire _20960_;
wire _20961_;
wire _20962_;
wire _20963_;
wire _20964_;
wire _20965_;
wire _20966_;
wire _20967_;
wire _20968_;
wire _20969_;
wire _20970_;
wire _20971_;
wire _20972_;
wire _20973_;
wire _20974_;
wire _20975_;
wire _20976_;
wire _20977_;
wire _20978_;
wire _20979_;
wire _20980_;
wire _20981_;
wire _20982_;
wire _20983_;
wire _20984_;
wire _20985_;
wire _20986_;
wire _20987_;
wire _20988_;
wire _20989_;
wire _20990_;
wire _20991_;
wire _20992_;
wire _20993_;
wire _20994_;
wire _20995_;
wire _20996_;
wire _20997_;
wire _20998_;
wire _20999_;
wire _21000_;
wire _21001_;
wire _21002_;
wire _21003_;
wire _21004_;
wire _21005_;
wire _21006_;
wire _21007_;
wire _21008_;
wire _21009_;
wire _21010_;
wire _21011_;
wire _21012_;
wire _21013_;
wire _21014_;
wire _21015_;
wire _21016_;
wire _21017_;
wire _21018_;
wire _21019_;
wire _21020_;
wire _21021_;
wire _21022_;
wire _21023_;
wire _21024_;
wire _21025_;
wire _21026_;
wire _21027_;
wire _21028_;
wire _21029_;
wire _21030_;
wire _21031_;
wire _21032_;
wire _21033_;
wire _21034_;
wire _21035_;
wire _21036_;
wire _21037_;
wire _21038_;
wire _21039_;
wire _21040_;
wire _21041_;
wire _21042_;
wire _21043_;
wire _21044_;
wire _21045_;
wire _21046_;
wire _21047_;
wire _21048_;
wire _21049_;
wire _21050_;
wire _21051_;
wire _21052_;
wire _21053_;
wire _21054_;
wire _21055_;
wire _21056_;
wire _21057_;
wire _21058_;
wire _21059_;
wire _21060_;
wire _21061_;
wire _21062_;
wire _21063_;
wire _21064_;
wire _21065_;
wire _21066_;
wire _21067_;
wire _21068_;
wire _21069_;
wire _21070_;
wire _21071_;
wire _21072_;
wire _21073_;
wire _21074_;
wire _21075_;
wire _21076_;
wire _21077_;
wire _21078_;
wire _21079_;
wire _21080_;
wire _21081_;
wire _21082_;
wire _21083_;
wire _21084_;
wire _21085_;
wire _21086_;
wire _21087_;
wire _21088_;
wire _21089_;
wire _21090_;
wire _21091_;
wire _21092_;
wire _21093_;
wire _21094_;
wire _21095_;
wire _21096_;
wire _21097_;
wire _21098_;
wire _21099_;
wire _21100_;
wire _21101_;
wire _21102_;
wire _21103_;
wire _21104_;
wire _21105_;
wire _21106_;
wire _21107_;
wire _21108_;
wire _21109_;
wire _21110_;
wire _21111_;
wire _21112_;
wire _21113_;
wire _21114_;
wire _21115_;
wire _21116_;
wire _21117_;
wire _21118_;
wire _21119_;
wire _21120_;
wire _21121_;
wire _21122_;
wire _21123_;
wire _21124_;
wire _21125_;
wire _21126_;
wire _21127_;
wire _21128_;
wire _21129_;
wire _21130_;
wire _21131_;
wire _21132_;
wire _21133_;
wire _21134_;
wire _21135_;
wire _21136_;
wire _21137_;
wire _21138_;
wire _21139_;
wire _21140_;
wire _21141_;
wire _21142_;
wire _21143_;
wire _21144_;
wire _21145_;
wire _21146_;
wire _21147_;
wire _21148_;
wire _21149_;
wire _21150_;
wire _21151_;
wire _21152_;
wire _21153_;
wire _21154_;
wire _21155_;
wire _21156_;
wire _21157_;
wire _21158_;
wire _21159_;
wire _21160_;
wire _21161_;
wire _21162_;
wire _21163_;
wire _21164_;
wire _21165_;
wire _21166_;
wire _21167_;
wire _21168_;
wire _21169_;
wire _21170_;
wire _21171_;
wire _21172_;
wire _21173_;
wire _21174_;
wire _21175_;
wire _21176_;
wire _21177_;
wire _21178_;
wire _21179_;
wire _21180_;
wire _21181_;
wire _21182_;
wire _21183_;
wire _21184_;
wire _21185_;
wire _21186_;
wire _21187_;
wire _21188_;
wire _21189_;
wire _21190_;
wire _21191_;
wire _21192_;
wire _21193_;
wire _21194_;
wire _21195_;
wire _21196_;
wire _21197_;
wire _21198_;
wire _21199_;
wire _21200_;
wire _21201_;
wire _21202_;
wire _21203_;
wire _21204_;
wire _21205_;
wire _21206_;
wire _21207_;
wire _21208_;
wire _21209_;
wire _21210_;
wire _21211_;
wire _21212_;
wire _21213_;
wire _21214_;
wire _21215_;
wire _21216_;
wire _21217_;
wire _21218_;
wire _21219_;
wire _21220_;
wire _21221_;
wire _21222_;
wire _21223_;
wire _21224_;
wire _21225_;
wire _21226_;
wire _21227_;
wire _21228_;
wire _21229_;
wire _21230_;
wire _21231_;
wire _21232_;
wire _21233_;
wire _21234_;
wire _21235_;
wire _21236_;
wire _21237_;
wire _21238_;
wire _21239_;
wire _21240_;
wire _21241_;
wire _21242_;
wire _21243_;
wire _21244_;
wire _21245_;
wire _21246_;
wire _21247_;
wire _21248_;
wire _21249_;
wire _21250_;
wire _21251_;
wire _21252_;
wire _21253_;
wire _21254_;
wire _21255_;
wire _21256_;
wire _21257_;
wire _21258_;
wire _21259_;
wire _21260_;
wire _21261_;
wire _21262_;
wire _21263_;
wire _21264_;
wire _21265_;
wire _21266_;
wire _21267_;
wire _21268_;
wire _21269_;
wire _21270_;
wire _21271_;
wire _21272_;
wire _21273_;
wire _21274_;
wire _21275_;
wire _21276_;
wire _21277_;
wire _21278_;
wire _21279_;
wire _21280_;
wire _21281_;
wire _21282_;
wire _21283_;
wire _21284_;
wire _21285_;
wire _21286_;
wire _21287_;
wire _21288_;
wire _21289_;
wire _21290_;
wire _21291_;
wire _21292_;
wire _21293_;
wire _21294_;
wire _21295_;
wire _21296_;
wire _21297_;
wire _21298_;
wire _21299_;
wire _21300_;
wire _21301_;
wire _21302_;
wire _21303_;
wire _21304_;
wire _21305_;
wire _21306_;
wire _21307_;
wire _21308_;
wire _21309_;
wire _21310_;
wire _21311_;
wire _21312_;
wire _21313_;
wire _21314_;
wire _21315_;
wire _21316_;
wire _21317_;
wire _21318_;
wire _21319_;
wire _21320_;
wire _21321_;
wire _21322_;
wire _21323_;
wire _21324_;
wire _21325_;
wire _21326_;
wire _21327_;
wire _21328_;
wire _21329_;
wire _21330_;
wire _21331_;
wire _21332_;
wire _21333_;
wire _21334_;
wire _21335_;
wire _21336_;
wire _21337_;
wire _21338_;
wire _21339_;
wire _21340_;
wire _21341_;
wire _21342_;
wire _21343_;
wire _21344_;
wire _21345_;
wire _21346_;
wire _21347_;
wire _21348_;
wire _21349_;
wire _21350_;
wire _21351_;
wire _21352_;
wire _21353_;
wire _21354_;
wire _21355_;
wire _21356_;
wire _21357_;
wire _21358_;
wire _21359_;
wire _21360_;
wire _21361_;
wire _21362_;
wire _21363_;
wire _21364_;
wire _21365_;
wire _21366_;
wire _21367_;
wire _21368_;
wire _21369_;
wire _21370_;
wire _21371_;
wire _21372_;
wire _21373_;
wire _21374_;
wire _21375_;
wire _21376_;
wire _21377_;
wire _21378_;
wire _21379_;
wire _21380_;
wire _21381_;
wire _21382_;
wire _21383_;
wire _21384_;
wire _21385_;
wire _21386_;
wire _21387_;
wire _21388_;
wire _21389_;
wire _21390_;
wire _21391_;
wire _21392_;
wire _21393_;
wire _21394_;
wire _21395_;
wire _21396_;
wire _21397_;
wire _21398_;
wire _21399_;
wire _21400_;
wire _21401_;
wire _21402_;
wire _21403_;
wire _21404_;
wire _21405_;
wire _21406_;
wire _21407_;
wire _21408_;
wire _21409_;
wire _21410_;
wire _21411_;
wire _21412_;
wire _21413_;
wire _21414_;
wire _21415_;
wire _21416_;
wire _21417_;
wire _21418_;
wire _21419_;
wire _21420_;
wire _21421_;
wire _21422_;
wire _21423_;
wire _21424_;
wire _21425_;
wire _21426_;
wire _21427_;
wire _21428_;
wire _21429_;
wire _21430_;
wire _21431_;
wire _21432_;
wire _21433_;
wire _21434_;
wire _21435_;
wire _21436_;
wire _21437_;
wire _21438_;
wire _21439_;
wire _21440_;
wire _21441_;
wire _21442_;
wire _21443_;
wire _21444_;
wire _21445_;
wire _21446_;
wire _21447_;
wire _21448_;
wire _21449_;
wire _21450_;
wire _21451_;
wire _21452_;
wire _21453_;
wire _21454_;
wire _21455_;
wire _21456_;
wire _21457_;
wire _21458_;
wire _21459_;
wire _21460_;
wire _21461_;
wire _21462_;
wire _21463_;
wire _21464_;
wire _21465_;
wire _21466_;
wire _21467_;
wire _21468_;
wire _21469_;
wire _21470_;
wire _21471_;
wire _21472_;
wire _21473_;
wire _21474_;
wire _21475_;
wire _21476_;
wire _21477_;
wire _21478_;
wire _21479_;
wire _21480_;
wire _21481_;
wire _21482_;
wire _21483_;
wire _21484_;
wire _21485_;
wire _21486_;
wire _21487_;
wire _21488_;
wire _21489_;
wire _21490_;
wire _21491_;
wire _21492_;
wire _21493_;
wire _21494_;
wire _21495_;
wire _21496_;
wire _21497_;
wire _21498_;
wire _21499_;
wire _21500_;
wire _21501_;
wire _21502_;
wire _21503_;
wire _21504_;
wire _21505_;
wire _21506_;
wire _21507_;
wire _21508_;
wire _21509_;
wire _21510_;
wire _21511_;
wire _21512_;
wire _21513_;
wire _21514_;
wire _21515_;
wire _21516_;
wire _21517_;
wire _21518_;
wire _21519_;
wire _21520_;
wire _21521_;
wire _21522_;
wire _21523_;
wire _21524_;
wire _21525_;
wire _21526_;
wire _21527_;
wire _21528_;
wire _21529_;
wire _21530_;
wire _21531_;
wire _21532_;
wire _21533_;
wire _21534_;
wire _21535_;
wire _21536_;
wire _21537_;
wire _21538_;
wire _21539_;
wire _21540_;
wire _21541_;
wire _21542_;
wire _21543_;
wire _21544_;
wire _21545_;
wire _21546_;
wire _21547_;
wire _21548_;
wire _21549_;
wire _21550_;
wire _21551_;
wire _21552_;
wire _21553_;
wire _21554_;
wire _21555_;
wire _21556_;
wire _21557_;
wire _21558_;
wire _21559_;
wire _21560_;
wire _21561_;
wire _21562_;
wire _21563_;
wire _21564_;
wire _21565_;
wire _21566_;
wire _21567_;
wire _21568_;
wire _21569_;
wire _21570_;
wire _21571_;
wire _21572_;
wire _21573_;
wire _21574_;
wire _21575_;
wire _21576_;
wire _21577_;
wire _21578_;
wire _21579_;
wire _21580_;
wire _21581_;
wire _21582_;
wire _21583_;
wire _21584_;
wire _21585_;
wire _21586_;
wire _21587_;
wire _21588_;
wire _21589_;
wire _21590_;
wire _21591_;
wire _21592_;
wire _21593_;
wire _21594_;
wire _21595_;
wire _21596_;
wire _21597_;
wire _21598_;
wire _21599_;
wire _21600_;
wire _21601_;
wire _21602_;
wire _21603_;
wire _21604_;
wire _21605_;
wire _21606_;
wire _21607_;
wire _21608_;
wire _21609_;
wire _21610_;
wire _21611_;
wire _21612_;
wire _21613_;
wire _21614_;
wire _21615_;
wire _21616_;
wire _21617_;
wire _21618_;
wire _21619_;
wire _21620_;
wire _21621_;
wire _21622_;
wire _21623_;
wire _21624_;
wire _21625_;
wire _21626_;
wire _21627_;
wire _21628_;
wire _21629_;
wire _21630_;
wire _21631_;
wire _21632_;
wire _21633_;
wire _21634_;
wire _21635_;
wire _21636_;
wire _21637_;
wire _21638_;
wire _21639_;
wire _21640_;
wire _21641_;
wire _21642_;
wire _21643_;
wire _21644_;
wire _21645_;
wire _21646_;
wire _21647_;
wire _21648_;
wire _21649_;
wire _21650_;
wire _21651_;
wire _21652_;
wire _21653_;
wire _21654_;
wire _21655_;
wire _21656_;
wire _21657_;
wire _21658_;
wire _21659_;
wire _21660_;
wire _21661_;
wire _21662_;
wire _21663_;
wire _21664_;
wire _21665_;
wire _21666_;
wire _21667_;
wire _21668_;
wire _21669_;
wire _21670_;
wire _21671_;
wire _21672_;
wire _21673_;
wire _21674_;
wire _21675_;
wire _21676_;
wire _21677_;
wire _21678_;
wire _21679_;
wire _21680_;
wire _21681_;
wire _21682_;
wire _21683_;
wire _21684_;
wire _21685_;
wire _21686_;
wire _21687_;
wire _21688_;
wire _21689_;
wire _21690_;
wire _21691_;
wire _21692_;
wire _21693_;
wire _21694_;
wire _21695_;
wire _21696_;
wire _21697_;
wire _21698_;
wire _21699_;
wire _21700_;
wire _21701_;
wire _21702_;
wire _21703_;
wire _21704_;
wire _21705_;
wire _21706_;
wire _21707_;
wire _21708_;
wire _21709_;
wire _21710_;
wire _21711_;
wire _21712_;
wire _21713_;
wire _21714_;
wire _21715_;
wire _21716_;
wire _21717_;
wire _21718_;
wire _21719_;
wire _21720_;
wire _21721_;
wire _21722_;
wire _21723_;
wire _21724_;
wire _21725_;
wire _21726_;
wire _21727_;
wire _21728_;
wire _21729_;
wire _21730_;
wire _21731_;
wire _21732_;
wire _21733_;
wire _21734_;
wire _21735_;
wire _21736_;
wire _21737_;
wire _21738_;
wire _21739_;
wire _21740_;
wire _21741_;
wire _21742_;
wire _21743_;
wire _21744_;
wire _21745_;
wire _21746_;
wire _21747_;
wire _21748_;
wire _21749_;
wire _21750_;
wire _21751_;
wire _21752_;
wire _21753_;
wire _21754_;
wire _21755_;
wire _21756_;
wire _21757_;
wire _21758_;
wire _21759_;
wire _21760_;
wire _21761_;
wire _21762_;
wire _21763_;
wire _21764_;
wire _21765_;
wire _21766_;
wire _21767_;
wire _21768_;
wire _21769_;
wire _21770_;
wire _21771_;
wire _21772_;
wire _21773_;
wire _21774_;
wire _21775_;
wire _21776_;
wire _21777_;
wire _21778_;
wire _21779_;
wire _21780_;
wire _21781_;
wire _21782_;
wire _21783_;
wire _21784_;
wire _21785_;
wire _21786_;
wire _21787_;
wire _21788_;
wire _21789_;
wire _21790_;
wire _21791_;
wire _21792_;
wire _21793_;
wire _21794_;
wire _21795_;
wire _21796_;
wire _21797_;
wire _21798_;
wire _21799_;
wire _21800_;
wire _21801_;
wire _21802_;
wire _21803_;
wire _21804_;
wire _21805_;
wire _21806_;
wire _21807_;
wire _21808_;
wire _21809_;
wire _21810_;
wire _21811_;
wire _21812_;
wire _21813_;
wire _21814_;
wire _21815_;
wire _21816_;
wire _21817_;
wire _21818_;
wire _21819_;
wire _21820_;
wire _21821_;
wire _21822_;
wire _21823_;
wire _21824_;
wire _21825_;
wire _21826_;
wire _21827_;
wire _21828_;
wire _21829_;
wire _21830_;
wire _21831_;
wire _21832_;
wire _21833_;
wire _21834_;
wire _21835_;
wire _21836_;
wire _21837_;
wire _21838_;
wire _21839_;
wire _21840_;
wire _21841_;
wire _21842_;
wire _21843_;
wire _21844_;
wire _21845_;
wire _21846_;
wire _21847_;
wire _21848_;
wire _21849_;
wire _21850_;
wire _21851_;
wire _21852_;
wire _21853_;
wire _21854_;
wire _21855_;
wire _21856_;
wire _21857_;
wire _21858_;
wire _21859_;
wire _21860_;
wire _21861_;
wire _21862_;
wire _21863_;
wire _21864_;
wire _21865_;
wire _21866_;
wire _21867_;
wire _21868_;
wire _21869_;
wire _21870_;
wire _21871_;
wire _21872_;
wire _21873_;
wire _21874_;
wire _21875_;
wire _21876_;
wire _21877_;
wire _21878_;
wire _21879_;
wire _21880_;
wire _21881_;
wire _21882_;
wire _21883_;
wire _21884_;
wire _21885_;
wire _21886_;
wire _21887_;
wire _21888_;
wire _21889_;
wire _21890_;
wire _21891_;
wire _21892_;
wire _21893_;
wire _21894_;
wire _21895_;
wire _21896_;
wire _21897_;
wire _21898_;
wire _21899_;
wire _21900_;
wire _21901_;
wire _21902_;
wire _21903_;
wire _21904_;
wire _21905_;
wire _21906_;
wire _21907_;
wire _21908_;
wire _21909_;
wire _21910_;
wire _21911_;
wire _21912_;
wire _21913_;
wire _21914_;
wire _21915_;
wire _21916_;
wire _21917_;
wire _21918_;
wire _21919_;
wire _21920_;
wire _21921_;
wire _21922_;
wire _21923_;
wire _21924_;
wire _21925_;
wire _21926_;
wire _21927_;
wire _21928_;
wire _21929_;
wire _21930_;
wire _21931_;
wire _21932_;
wire _21933_;
wire _21934_;
wire _21935_;
wire _21936_;
wire _21937_;
wire _21938_;
wire _21939_;
wire _21940_;
wire _21941_;
wire _21942_;
wire _21943_;
wire _21944_;
wire _21945_;
wire _21946_;
wire _21947_;
wire _21948_;
wire _21949_;
wire _21950_;
wire _21951_;
wire _21952_;
wire _21953_;
wire _21954_;
wire _21955_;
wire _21956_;
wire _21957_;
wire _21958_;
wire _21959_;
wire _21960_;
wire _21961_;
wire _21962_;
wire _21963_;
wire _21964_;
wire _21965_;
wire _21966_;
wire _21967_;
wire _21968_;
wire _21969_;
wire _21970_;
wire _21971_;
wire _21972_;
wire _21973_;
wire _21974_;
wire _21975_;
wire _21976_;
wire _21977_;
wire _21978_;
wire _21979_;
wire _21980_;
wire _21981_;
wire _21982_;
wire _21983_;
wire _21984_;
wire _21985_;
wire _21986_;
wire _21987_;
wire _21988_;
wire _21989_;
wire _21990_;
wire _21991_;
wire _21992_;
wire _21993_;
wire _21994_;
wire _21995_;
wire _21996_;
wire _21997_;
wire _21998_;
wire _21999_;
wire _22000_;
wire _22001_;
wire _22002_;
wire _22003_;
wire _22004_;
wire _22005_;
wire _22006_;
wire _22007_;
wire _22008_;
wire _22009_;
wire _22010_;
wire _22011_;
wire _22012_;
wire _22013_;
wire _22014_;
wire _22015_;
wire _22016_;
wire _22017_;
wire _22018_;
wire _22019_;
wire _22020_;
wire _22021_;
wire _22022_;
wire _22023_;
wire _22024_;
wire _22025_;
wire _22026_;
wire _22027_;
wire _22028_;
wire _22029_;
wire _22030_;
wire _22031_;
wire _22032_;
wire _22033_;
wire _22034_;
wire _22035_;
wire _22036_;
wire _22037_;
wire _22038_;
wire _22039_;
wire _22040_;
wire _22041_;
wire _22042_;
wire _22043_;
wire _22044_;
wire _22045_;
wire _22046_;
wire _22047_;
wire _22048_;
wire _22049_;
wire _22050_;
wire _22051_;
wire _22052_;
wire _22053_;
wire _22054_;
wire _22055_;
wire _22056_;
wire _22057_;
wire _22058_;
wire _22059_;
wire _22060_;
wire _22061_;
wire _22062_;
wire _22063_;
wire _22064_;
wire _22065_;
wire _22066_;
wire _22067_;
wire _22068_;
wire _22069_;
wire _22070_;
wire _22071_;
wire _22072_;
wire _22073_;
wire _22074_;
wire _22075_;
wire _22076_;
wire _22077_;
wire _22078_;
wire _22079_;
wire _22080_;
wire _22081_;
wire _22082_;
wire _22083_;
wire _22084_;
wire _22085_;
wire _22086_;
wire _22087_;
wire _22088_;
wire _22089_;
wire _22090_;
wire _22091_;
wire _22092_;
wire _22093_;
wire _22094_;
wire _22095_;
wire _22096_;
wire _22097_;
wire _22098_;
wire _22099_;
wire _22100_;
wire _22101_;
wire _22102_;
wire _22103_;
wire _22104_;
wire _22105_;
wire _22106_;
wire _22107_;
wire _22108_;
wire _22109_;
wire _22110_;
wire _22111_;
wire _22112_;
wire _22113_;
wire _22114_;
wire _22115_;
wire _22116_;
wire _22117_;
wire _22118_;
wire _22119_;
wire _22120_;
wire _22121_;
wire _22122_;
wire _22123_;
wire _22124_;
wire _22125_;
wire _22126_;
wire _22127_;
wire _22128_;
wire _22129_;
wire _22130_;
wire _22131_;
wire _22132_;
wire _22133_;
wire _22134_;
wire _22135_;
wire _22136_;
wire _22137_;
wire _22138_;
wire _22139_;
wire _22140_;
wire _22141_;
wire _22142_;
wire _22143_;
wire _22144_;
wire _22145_;
wire _22146_;
wire _22147_;
wire _22148_;
wire _22149_;
wire _22150_;
wire _22151_;
wire _22152_;
wire _22153_;
wire _22154_;
wire _22155_;
wire _22156_;
wire _22157_;
wire _22158_;
wire _22159_;
wire _22160_;
wire _22161_;
wire _22162_;
wire _22163_;
wire _22164_;
wire _22165_;
wire _22166_;
wire _22167_;
wire _22168_;
wire _22169_;
wire _22170_;
wire _22171_;
wire _22172_;
wire _22173_;
wire _22174_;
wire _22175_;
wire _22176_;
wire _22177_;
wire _22178_;
wire _22179_;
wire _22180_;
wire _22181_;
wire _22182_;
wire _22183_;
wire _22184_;
wire _22185_;
wire _22186_;
wire _22187_;
wire _22188_;
wire _22189_;
wire _22190_;
wire _22191_;
wire _22192_;
wire _22193_;
wire _22194_;
wire _22195_;
wire _22196_;
wire _22197_;
wire _22198_;
wire _22199_;
wire _22200_;
wire _22201_;
wire _22202_;
wire _22203_;
wire _22204_;
wire _22205_;
wire _22206_;
wire _22207_;
wire _22208_;
wire _22209_;
wire _22210_;
wire _22211_;
wire _22212_;
wire _22213_;
wire _22214_;
wire _22215_;
wire _22216_;
wire _22217_;
wire _22218_;
wire _22219_;
wire _22220_;
wire _22221_;
wire _22222_;
wire _22223_;
wire _22224_;
wire _22225_;
wire _22226_;
wire _22227_;
wire _22228_;
wire _22229_;
wire _22230_;
wire _22231_;
wire _22232_;
wire _22233_;
wire _22234_;
wire _22235_;
wire _22236_;
wire _22237_;
wire _22238_;
wire _22239_;
wire _22240_;
wire _22241_;
wire _22242_;
wire _22243_;
wire _22244_;
wire _22245_;
wire _22246_;
wire _22247_;
wire _22248_;
wire _22249_;
wire _22250_;
wire _22251_;
wire _22252_;
wire _22253_;
wire _22254_;
wire _22255_;
wire _22256_;
wire _22257_;
wire _22258_;
wire _22259_;
wire _22260_;
wire _22261_;
wire _22262_;
wire _22263_;
wire _22264_;
wire _22265_;
wire _22266_;
wire _22267_;
wire _22268_;
wire _22269_;
wire _22270_;
wire _22271_;
wire _22272_;
wire _22273_;
wire _22274_;
wire _22275_;
wire _22276_;
wire _22277_;
wire _22278_;
wire _22279_;
wire _22280_;
wire _22281_;
wire _22282_;
wire _22283_;
wire _22284_;
wire _22285_;
wire _22286_;
wire _22287_;
wire _22288_;
wire _22289_;
wire _22290_;
wire _22291_;
wire _22292_;
wire _22293_;
wire _22294_;
wire _22295_;
wire _22296_;
wire _22297_;
wire _22298_;
wire _22299_;
wire _22300_;
wire _22301_;
wire _22302_;
wire _22303_;
wire _22304_;
wire _22305_;
wire _22306_;
wire _22307_;
wire _22308_;
wire _22309_;
wire _22310_;
wire _22311_;
wire _22312_;
wire _22313_;
wire _22314_;
wire _22315_;
wire _22316_;
wire _22317_;
wire _22318_;
wire _22319_;
wire _22320_;
wire _22321_;
wire _22322_;
wire _22323_;
wire _22324_;
wire _22325_;
wire _22326_;
wire _22327_;
wire _22328_;
wire _22329_;
wire _22330_;
wire _22331_;
wire _22332_;
wire _22333_;
wire _22334_;
wire _22335_;
wire _22336_;
wire _22337_;
wire _22338_;
wire _22339_;
wire _22340_;
wire _22341_;
wire _22342_;
wire _22343_;
wire _22344_;
wire _22345_;
wire _22346_;
wire _22347_;
wire _22348_;
wire _22349_;
wire _22350_;
wire _22351_;
wire _22352_;
wire _22353_;
wire _22354_;
wire _22355_;
wire _22356_;
wire _22357_;
wire _22358_;
wire _22359_;
wire _22360_;
wire _22361_;
wire _22362_;
wire _22363_;
wire _22364_;
wire _22365_;
wire _22366_;
wire _22367_;
wire _22368_;
wire _22369_;
wire _22370_;
wire _22371_;
wire _22372_;
wire _22373_;
wire _22374_;
wire _22375_;
wire _22376_;
wire _22377_;
wire _22378_;
wire _22379_;
wire _22380_;
wire _22381_;
wire _22382_;
wire _22383_;
wire _22384_;
wire _22385_;
wire _22386_;
wire _22387_;
wire _22388_;
wire _22389_;
wire _22390_;
wire _22391_;
wire _22392_;
wire _22393_;
wire _22394_;
wire _22395_;
wire _22396_;
wire _22397_;
wire _22398_;
wire _22399_;
wire _22400_;
wire _22401_;
wire _22402_;
wire _22403_;
wire _22404_;
wire _22405_;
wire _22406_;
wire _22407_;
wire _22408_;
wire _22409_;
wire _22410_;
wire _22411_;
wire _22412_;
wire _22413_;
wire _22414_;
wire _22415_;
wire _22416_;
wire _22417_;
wire _22418_;
wire _22419_;
wire _22420_;
wire _22421_;
wire _22422_;
wire _22423_;
wire _22424_;
wire _22425_;
wire _22426_;
wire _22427_;
wire _22428_;
wire _22429_;
wire _22430_;
wire _22431_;
wire _22432_;
wire _22433_;
wire _22434_;
wire _22435_;
wire _22436_;
wire _22437_;
wire _22438_;
wire _22439_;
wire _22440_;
wire _22441_;
wire _22442_;
wire _22443_;
wire _22444_;
wire _22445_;
wire _22446_;
wire _22447_;
wire _22448_;
wire _22449_;
wire _22450_;
wire _22451_;
wire _22452_;
wire _22453_;
wire _22454_;
wire _22455_;
wire _22456_;
wire _22457_;
wire _22458_;
wire _22459_;
wire _22460_;
wire _22461_;
wire _22462_;
wire _22463_;
wire _22464_;
wire _22465_;
wire _22466_;
wire _22467_;
wire _22468_;
wire _22469_;
wire _22470_;
wire _22471_;
wire _22472_;
wire _22473_;
wire _22474_;
wire _22475_;
wire _22476_;
wire _22477_;
wire _22478_;
wire _22479_;
wire _22480_;
wire _22481_;
wire _22482_;
wire _22483_;
wire _22484_;
wire _22485_;
wire _22486_;
wire _22487_;
wire _22488_;
wire _22489_;
wire _22490_;
wire _22491_;
wire _22492_;
wire _22493_;
wire _22494_;
wire _22495_;
wire _22496_;
wire _22497_;
wire _22498_;
wire _22499_;
wire _22500_;
wire _22501_;
wire _22502_;
wire _22503_;
wire _22504_;
wire _22505_;
wire _22506_;
wire _22507_;
wire _22508_;
wire _22509_;
wire _22510_;
wire _22511_;
wire _22512_;
wire _22513_;
wire _22514_;
wire _22515_;
wire _22516_;
wire _22517_;
wire _22518_;
wire _22519_;
wire _22520_;
wire _22521_;
wire _22522_;
wire _22523_;
wire _22524_;
wire _22525_;
wire _22526_;
wire _22527_;
wire _22528_;
wire _22529_;
wire _22530_;
wire _22531_;
wire _22532_;
wire _22533_;
wire _22534_;
wire _22535_;
wire _22536_;
wire _22537_;
wire _22538_;
wire _22539_;
wire _22540_;
wire _22541_;
wire _22542_;
wire _22543_;
wire _22544_;
wire _22545_;
wire _22546_;
wire _22547_;
wire _22548_;
wire _22549_;
wire _22550_;
wire _22551_;
wire _22552_;
wire _22553_;
wire _22554_;
wire _22555_;
wire _22556_;
wire _22557_;
wire _22558_;
wire _22559_;
wire _22560_;
wire _22561_;
wire _22562_;
wire _22563_;
wire _22564_;
wire _22565_;
wire _22566_;
wire _22567_;
wire _22568_;
wire _22569_;
wire _22570_;
wire _22571_;
wire _22572_;
wire _22573_;
wire _22574_;
wire _22575_;
wire _22576_;
wire _22577_;
wire _22578_;
wire _22579_;
wire _22580_;
wire _22581_;
wire _22582_;
wire _22583_;
wire _22584_;
wire _22585_;
wire _22586_;
wire _22587_;
wire _22588_;
wire _22589_;
wire _22590_;
wire _22591_;
wire _22592_;
wire _22593_;
wire _22594_;
wire _22595_;
wire _22596_;
wire _22597_;
wire _22598_;
wire _22599_;
wire _22600_;
wire _22601_;
wire _22602_;
wire _22603_;
wire _22604_;
wire _22605_;
wire _22606_;
wire _22607_;
wire _22608_;
wire _22609_;
wire _22610_;
wire _22611_;
wire _22612_;
wire _22613_;
wire _22614_;
wire _22615_;
wire _22616_;
wire _22617_;
wire _22618_;
wire _22619_;
wire _22620_;
wire _22621_;
wire _22622_;
wire _22623_;
wire _22624_;
wire _22625_;
wire _22626_;
wire _22627_;
wire _22628_;
wire _22629_;
wire _22630_;
wire _22631_;
wire _22632_;
wire _22633_;
wire _22634_;
wire _22635_;
wire _22636_;
wire _22637_;
wire _22638_;
wire _22639_;
wire _22640_;
wire _22641_;
wire _22642_;
wire _22643_;
wire _22644_;
wire _22645_;
wire _22646_;
wire _22647_;
wire _22648_;
wire _22649_;
wire _22650_;
wire _22651_;
wire _22652_;
wire _22653_;
wire _22654_;
wire _22655_;
wire _22656_;
wire _22657_;
wire _22658_;
wire _22659_;
wire _22660_;
wire _22661_;
wire _22662_;
wire _22663_;
wire _22664_;
wire _22665_;
wire _22666_;
wire _22667_;
wire _22668_;
wire _22669_;
wire _22670_;
wire _22671_;
wire _22672_;
wire _22673_;
wire _22674_;
wire _22675_;
wire _22676_;
wire _22677_;
wire _22678_;
wire _22679_;
wire _22680_;
wire _22681_;
wire _22682_;
wire _22683_;
wire _22684_;
wire _22685_;
wire _22686_;
wire _22687_;
wire _22688_;
wire _22689_;
wire _22690_;
wire _22691_;
wire _22692_;
wire _22693_;
wire _22694_;
wire _22695_;
wire _22696_;
wire _22697_;
wire _22698_;
wire _22699_;
wire _22700_;
wire _22701_;
wire _22702_;
wire _22703_;
wire _22704_;
wire _22705_;
wire _22706_;
wire _22707_;
wire _22708_;
wire _22709_;
wire _22710_;
wire _22711_;
wire _22712_;
wire _22713_;
wire _22714_;
wire _22715_;
wire _22716_;
wire _22717_;
wire _22718_;
wire _22719_;
wire _22720_;
wire _22721_;
wire _22722_;
wire _22723_;
wire _22724_;
wire _22725_;
wire _22726_;
wire _22727_;
wire _22728_;
wire _22729_;
wire _22730_;
wire _22731_;
wire _22732_;
wire _22733_;
wire _22734_;
wire _22735_;
wire _22736_;
wire _22737_;
wire _22738_;
wire _22739_;
wire _22740_;
wire _22741_;
wire _22742_;
wire _22743_;
wire _22744_;
wire _22745_;
wire _22746_;
wire _22747_;
wire _22748_;
wire _22749_;
wire _22750_;
wire _22751_;
wire _22752_;
wire _22753_;
wire _22754_;
wire _22755_;
wire _22756_;
wire _22757_;
wire _22758_;
wire _22759_;
wire _22760_;
wire _22761_;
wire _22762_;
wire _22763_;
wire _22764_;
wire _22765_;
wire _22766_;
wire _22767_;
wire _22768_;
wire _22769_;
wire _22770_;
wire _22771_;
wire _22772_;
wire _22773_;
wire _22774_;
wire _22775_;
wire _22776_;
wire _22777_;
wire _22778_;
wire _22779_;
wire _22780_;
wire _22781_;
wire _22782_;
wire _22783_;
wire _22784_;
wire _22785_;
wire _22786_;
wire _22787_;
wire _22788_;
wire _22789_;
wire _22790_;
wire _22791_;
wire _22792_;
wire _22793_;
wire _22794_;
wire _22795_;
wire _22796_;
wire _22797_;
wire _22798_;
wire _22799_;
wire _22800_;
wire _22801_;
wire _22802_;
wire _22803_;
wire _22804_;
wire _22805_;
wire _22806_;
wire _22807_;
wire _22808_;
wire _22809_;
wire _22810_;
wire _22811_;
wire _22812_;
wire _22813_;
wire _22814_;
wire _22815_;
wire _22816_;
wire _22817_;
wire _22818_;
wire _22819_;
wire _22820_;
wire _22821_;
wire _22822_;
wire _22823_;
wire _22824_;
wire _22825_;
wire _22826_;
wire _22827_;
wire _22828_;
wire _22829_;
wire _22830_;
wire _22831_;
wire _22832_;
wire _22833_;
wire _22834_;
wire _22835_;
wire _22836_;
wire _22837_;
wire _22838_;
wire _22839_;
wire _22840_;
wire _22841_;
wire _22842_;
wire _22843_;
wire _22844_;
wire _22845_;
wire _22846_;
wire _22847_;
wire _22848_;
wire _22849_;
wire _22850_;
wire _22851_;
wire _22852_;
wire _22853_;
wire _22854_;
wire _22855_;
wire _22856_;
wire _22857_;
wire _22858_;
wire _22859_;
wire _22860_;
wire _22861_;
wire _22862_;
wire _22863_;
wire _22864_;
wire _22865_;
wire _22866_;
wire _22867_;
wire _22868_;
wire _22869_;
wire _22870_;
wire _22871_;
wire _22872_;
wire _22873_;
wire _22874_;
wire _22875_;
wire _22876_;
wire _22877_;
wire _22878_;
wire _22879_;
wire _22880_;
wire _22881_;
wire _22882_;
wire _22883_;
wire _22884_;
wire _22885_;
wire _22886_;
wire _22887_;
wire _22888_;
wire _22889_;
wire _22890_;
wire _22891_;
wire _22892_;
wire _22893_;
wire _22894_;
wire _22895_;
wire _22896_;
wire _22897_;
wire _22898_;
wire _22899_;
wire _22900_;
wire _22901_;
wire _22902_;
wire _22903_;
wire _22904_;
wire _22905_;
wire _22906_;
wire _22907_;
wire _22908_;
wire _22909_;
wire _22910_;
wire _22911_;
wire _22912_;
wire _22913_;
wire _22914_;
wire _22915_;
wire _22916_;
wire _22917_;
wire _22918_;
wire _22919_;
wire _22920_;
wire _22921_;
wire _22922_;
wire _22923_;
wire _22924_;
wire _22925_;
wire _22926_;
wire _22927_;
wire _22928_;
wire _22929_;
wire _22930_;
wire _22931_;
wire _22932_;
wire _22933_;
wire _22934_;
wire _22935_;
wire _22936_;
wire _22937_;
wire _22938_;
wire _22939_;
wire _22940_;
wire _22941_;
wire _22942_;
wire _22943_;
wire _22944_;
wire _22945_;
wire _22946_;
wire _22947_;
wire _22948_;
wire _22949_;
wire _22950_;
wire _22951_;
wire _22952_;
wire _22953_;
wire _22954_;
wire _22955_;
wire _22956_;
wire _22957_;
wire _22958_;
wire _22959_;
wire _22960_;
wire _22961_;
wire _22962_;
wire _22963_;
wire _22964_;
wire _22965_;
wire _22966_;
wire _22967_;
wire _22968_;
wire _22969_;
wire _22970_;
wire _22971_;
wire _22972_;
wire _22973_;
wire _22974_;
wire _22975_;
wire _22976_;
wire _22977_;
wire _22978_;
wire _22979_;
wire _22980_;
wire _22981_;
wire _22982_;
wire _22983_;
wire _22984_;
wire _22985_;
wire _22986_;
wire _22987_;
wire _22988_;
wire _22989_;
wire _22990_;
wire _22991_;
wire _22992_;
wire _22993_;
wire _22994_;
wire _22995_;
wire _22996_;
wire _22997_;
wire _22998_;
wire _22999_;
wire _23000_;
wire _23001_;
wire _23002_;
wire _23003_;
wire _23004_;
wire _23005_;
wire _23006_;
wire _23007_;
wire _23008_;
wire _23009_;
wire _23010_;
wire _23011_;
wire _23012_;
wire _23013_;
wire _23014_;
wire _23015_;
wire _23016_;
wire _23017_;
wire _23018_;
wire _23019_;
wire _23020_;
wire _23021_;
wire _23022_;
wire _23023_;
wire _23024_;
wire _23025_;
wire _23026_;
wire _23027_;
wire _23028_;
wire _23029_;
wire _23030_;
wire _23031_;
wire _23032_;
wire _23033_;
wire _23034_;
wire _23035_;
wire _23036_;
wire _23037_;
wire _23038_;
wire _23039_;
wire _23040_;
wire _23041_;
wire _23042_;
wire _23043_;
wire _23044_;
wire _23045_;
wire _23046_;
wire _23047_;
wire _23048_;
wire _23049_;
wire _23050_;
wire _23051_;
wire _23052_;
wire _23053_;
wire _23054_;
wire _23055_;
wire _23056_;
wire _23057_;
wire _23058_;
wire _23059_;
wire _23060_;
wire _23061_;
wire _23062_;
wire _23063_;
wire _23064_;
wire _23065_;
wire _23066_;
wire _23067_;
wire _23068_;
wire _23069_;
wire _23070_;
wire _23071_;
wire _23072_;
wire _23073_;
wire _23074_;
wire _23075_;
wire _23076_;
wire _23077_;
wire _23078_;
wire _23079_;
wire _23080_;
wire _23081_;
wire _23082_;
wire _23083_;
wire _23084_;
wire _23085_;
wire _23086_;
wire _23087_;
wire _23088_;
wire _23089_;
wire _23090_;
wire _23091_;
wire _23092_;
wire _23093_;
wire _23094_;
wire _23095_;
wire _23096_;
wire _23097_;
wire _23098_;
wire _23099_;
wire _23100_;
wire _23101_;
wire _23102_;
wire _23103_;
wire _23104_;
wire _23105_;
wire _23106_;
wire _23107_;
wire _23108_;
wire _23109_;
wire _23110_;
wire _23111_;
wire _23112_;
wire _23113_;
wire _23114_;
wire _23115_;
wire _23116_;
wire _23117_;
wire _23118_;
wire _23119_;
wire _23120_;
wire _23121_;
wire _23122_;
wire _23123_;
wire _23124_;
wire _23125_;
wire _23126_;
wire _23127_;
wire _23128_;
wire _23129_;
wire _23130_;
wire _23131_;
wire _23132_;
wire _23133_;
wire _23134_;
wire _23135_;
wire _23136_;
wire _23137_;
wire _23138_;
wire _23139_;
wire _23140_;
wire _23141_;
wire _23142_;
wire _23143_;
wire _23144_;
wire _23145_;
wire _23146_;
wire _23147_;
wire _23148_;
wire _23149_;
wire _23150_;
wire _23151_;
wire _23152_;
wire _23153_;
wire _23154_;
wire _23155_;
wire _23156_;
wire _23157_;
wire _23158_;
wire _23159_;
wire _23160_;
wire _23161_;
wire _23162_;
wire _23163_;
wire _23164_;
wire _23165_;
wire _23166_;
wire _23167_;
wire _23168_;
wire _23169_;
wire _23170_;
wire _23171_;
wire _23172_;
wire _23173_;
wire _23174_;
wire _23175_;
wire _23176_;
wire _23177_;
wire _23178_;
wire _23179_;
wire _23180_;
wire _23181_;
wire _23182_;
wire _23183_;
wire _23184_;
wire _23185_;
wire _23186_;
wire _23187_;
wire _23188_;
wire _23189_;
wire _23190_;
wire _23191_;
wire _23192_;
wire _23193_;
wire _23194_;
wire _23195_;
wire _23196_;
wire _23197_;
wire _23198_;
wire _23199_;
wire _23200_;
wire _23201_;
wire _23202_;
wire _23203_;
wire _23204_;
wire _23205_;
wire _23206_;
wire _23207_;
wire _23208_;
wire _23209_;
wire _23210_;
wire _23211_;
wire _23212_;
wire _23213_;
wire _23214_;
wire _23215_;
wire _23216_;
wire _23217_;
wire _23218_;
wire _23219_;
wire _23220_;
wire _23221_;
wire _23222_;
wire _23223_;
wire _23224_;
wire _23225_;
wire _23226_;
wire _23227_;
wire _23228_;
wire _23229_;
wire _23230_;
wire _23231_;
wire _23232_;
wire _23233_;
wire _23234_;
wire _23235_;
wire _23236_;
wire _23237_;
wire _23238_;
wire _23239_;
wire _23240_;
wire _23241_;
wire _23242_;
wire _23243_;
wire _23244_;
wire _23245_;
wire _23246_;
wire _23247_;
wire _23248_;
wire _23249_;
wire _23250_;
wire _23251_;
wire _23252_;
wire _23253_;
wire _23254_;
wire _23255_;
wire _23256_;
wire _23257_;
wire _23258_;
wire _23259_;
wire _23260_;
wire _23261_;
wire _23262_;
wire _23263_;
wire _23264_;
wire _23265_;
wire _23266_;
wire _23267_;
wire _23268_;
wire _23269_;
wire _23270_;
wire _23271_;
wire _23272_;
wire _23273_;
wire _23274_;
wire _23275_;
wire _23276_;
wire _23277_;
wire _23278_;
wire _23279_;
wire _23280_;
wire _23281_;
wire _23282_;
wire _23283_;
wire _23284_;
wire _23285_;
wire _23286_;
wire _23287_;
wire _23288_;
wire _23289_;
wire _23290_;
wire _23291_;
wire _23292_;
wire _23293_;
wire _23294_;
wire _23295_;
wire _23296_;
wire _23297_;
wire _23298_;
wire _23299_;
wire _23300_;
wire _23301_;
wire _23302_;
wire _23303_;
wire _23304_;
wire _23305_;
wire _23306_;
wire _23307_;
wire _23308_;
wire _23309_;
wire _23310_;
wire _23311_;
wire _23312_;
wire _23313_;
wire _23314_;
wire _23315_;
wire _23316_;
wire _23317_;
wire _23318_;
wire _23319_;
wire _23320_;
wire _23321_;
wire _23322_;
wire _23323_;
wire _23324_;
wire _23325_;
wire _23326_;
wire _23327_;
wire _23328_;
wire _23329_;
wire _23330_;
wire _23331_;
wire _23332_;
wire _23333_;
wire _23334_;
wire _23335_;
wire _23336_;
wire _23337_;
wire _23338_;
wire _23339_;
wire _23340_;
wire _23341_;
wire _23342_;
wire _23343_;
wire _23344_;
wire _23345_;
wire _23346_;
wire _23347_;
wire _23348_;
wire _23349_;
wire _23350_;
wire _23351_;
wire _23352_;
wire _23353_;
wire _23354_;
wire _23355_;
wire _23356_;
wire _23357_;
wire _23358_;
wire _23359_;
wire _23360_;
wire _23361_;
wire _23362_;
wire _23363_;
wire _23364_;
wire _23365_;
wire _23366_;
wire _23367_;
wire _23368_;
wire _23369_;
wire _23370_;
wire _23371_;
wire _23372_;
wire _23373_;
wire _23374_;
wire _23375_;
wire _23376_;
wire _23377_;
wire _23378_;
wire _23379_;
wire _23380_;
wire _23381_;
wire _23382_;
wire _23383_;
wire _23384_;
wire _23385_;
wire _23386_;
wire _23387_;
wire _23388_;
wire _23389_;
wire _23390_;
wire _23391_;
wire _23392_;
wire _23393_;
wire _23394_;
wire _23395_;
wire _23396_;
wire _23397_;
wire _23398_;
wire _23399_;
wire _23400_;
wire _23401_;
wire _23402_;
wire _23403_;
wire _23404_;
wire _23405_;
wire _23406_;
wire _23407_;
wire _23408_;
wire _23409_;
wire _23410_;
wire _23411_;
wire _23412_;
wire _23413_;
wire _23414_;
wire _23415_;
wire _23416_;
wire _23417_;
wire _23418_;
wire _23419_;
wire _23420_;
wire _23421_;
wire _23422_;
wire _23423_;
wire _23424_;
wire _23425_;
wire _23426_;
wire _23427_;
wire _23428_;
wire _23429_;
wire _23430_;
wire _23431_;
wire _23432_;
wire _23433_;
wire _23434_;
wire _23435_;
wire _23436_;
wire _23437_;
wire _23438_;
wire _23439_;
wire _23440_;
wire _23441_;
wire _23442_;
wire _23443_;
wire _23444_;
wire _23445_;
wire _23446_;
wire _23447_;
wire _23448_;
wire _23449_;
wire _23450_;
wire _23451_;
wire _23452_;
wire _23453_;
wire _23454_;
wire _23455_;
wire _23456_;
wire _23457_;
wire _23458_;
wire _23459_;
wire _23460_;
wire _23461_;
wire _23462_;
wire _23463_;
wire _23464_;
wire _23465_;
wire _23466_;
wire _23467_;
wire _23468_;
wire _23469_;
wire _23470_;
wire _23471_;
wire _23472_;
wire _23473_;
wire _23474_;
wire _23475_;
wire _23476_;
wire _23477_;
wire _23478_;
wire _23479_;
wire _23480_;
wire _23481_;
wire _23482_;
wire _23483_;
wire _23484_;
wire _23485_;
wire _23486_;
wire _23487_;
wire _23488_;
wire _23489_;
wire _23490_;
wire _23491_;
wire _23492_;
wire _23493_;
wire _23494_;
wire _23495_;
wire _23496_;
wire _23497_;
wire _23498_;
wire _23499_;
wire _23500_;
wire _23501_;
wire _23502_;
wire _23503_;
wire _23504_;
wire _23505_;
wire _23506_;
wire _23507_;
wire _23508_;
wire _23509_;
wire _23510_;
wire _23511_;
wire _23512_;
wire _23513_;
wire _23514_;
wire _23515_;
wire _23516_;
wire _23517_;
wire _23518_;
wire _23519_;
wire _23520_;
wire _23521_;
wire _23522_;
wire _23523_;
wire _23524_;
wire _23525_;
wire _23526_;
wire _23527_;
wire _23528_;
wire _23529_;
wire _23530_;
wire _23531_;
wire _23532_;
wire _23533_;
wire _23534_;
wire _23535_;
wire _23536_;
wire _23537_;
wire _23538_;
wire _23539_;
wire _23540_;
wire _23541_;
wire _23542_;
wire _23543_;
wire _23544_;
wire _23545_;
wire _23546_;
wire _23547_;
wire _23548_;
wire _23549_;
wire _23550_;
wire _23551_;
wire _23552_;
wire _23553_;
wire _23554_;
wire _23555_;
wire _23556_;
wire _23557_;
wire _23558_;
wire _23559_;
wire _23560_;
wire _23561_;
wire _23562_;
wire _23563_;
wire _23564_;
wire _23565_;
wire _23566_;
wire _23567_;
wire _23568_;
wire _23569_;
wire _23570_;
wire _23571_;
wire _23572_;
wire _23573_;
wire _23574_;
wire _23575_;
wire _23576_;
wire _23577_;
wire _23578_;
wire _23579_;
wire _23580_;
wire _23581_;
wire _23582_;
wire _23583_;
wire _23584_;
wire _23585_;
wire _23586_;
wire _23587_;
wire _23588_;
wire _23589_;
wire _23590_;
wire _23591_;
wire _23592_;
wire _23593_;
wire _23594_;
wire _23595_;
wire _23596_;
wire _23597_;
wire _23598_;
wire _23599_;
wire _23600_;
wire _23601_;
wire _23602_;
wire _23603_;
wire _23604_;
wire _23605_;
wire _23606_;
wire _23607_;
wire _23608_;
wire _23609_;
wire _23610_;
wire _23611_;
wire _23612_;
wire _23613_;
wire _23614_;
wire _23615_;
wire _23616_;
wire _23617_;
wire _23618_;
wire _23619_;
wire _23620_;
wire _23621_;
wire _23622_;
wire _23623_;
wire _23624_;
wire _23625_;
wire _23626_;
wire _23627_;
wire _23628_;
wire _23629_;
wire _23630_;
wire _23631_;
wire _23632_;
wire _23633_;
wire _23634_;
wire _23635_;
wire _23636_;
wire _23637_;
wire _23638_;
wire _23639_;
wire _23640_;
wire _23641_;
wire _23642_;
wire _23643_;
wire _23644_;
wire _23645_;
wire _23646_;
wire _23647_;
wire _23648_;
wire _23649_;
wire _23650_;
wire _23651_;
wire _23652_;
wire _23653_;
wire _23654_;
wire _23655_;
wire _23656_;
wire _23657_;
wire _23658_;
wire _23659_;
wire _23660_;
wire _23661_;
wire _23662_;
wire _23663_;
wire _23664_;
wire _23665_;
wire _23666_;
wire _23667_;
wire _23668_;
wire _23669_;
wire _23670_;
wire _23671_;
wire _23672_;
wire _23673_;
wire _23674_;
wire _23675_;
wire _23676_;
wire _23677_;
wire _23678_;
wire _23679_;
wire _23680_;
wire _23681_;
wire _23682_;
wire _23683_;
wire _23684_;
wire _23685_;
wire _23686_;
wire _23687_;
wire _23688_;
wire _23689_;
wire _23690_;
wire _23691_;
wire _23692_;
wire _23693_;
wire _23694_;
wire _23695_;
wire _23696_;
wire _23697_;
wire _23698_;
wire _23699_;
wire _23700_;
wire _23701_;
wire _23702_;
wire _23703_;
wire _23704_;
wire _23705_;
wire _23706_;
wire _23707_;
wire _23708_;
wire _23709_;
wire _23710_;
wire _23711_;
wire _23712_;
wire _23713_;
wire _23714_;
wire _23715_;
wire _23716_;
wire _23717_;
wire _23718_;
wire _23719_;
wire _23720_;
wire _23721_;
wire _23722_;
wire _23723_;
wire _23724_;
wire _23725_;
wire _23726_;
wire _23727_;
wire _23728_;
wire _23729_;
wire _23730_;
wire _23731_;
wire _23732_;
wire _23733_;
wire _23734_;
wire _23735_;
wire _23736_;
wire _23737_;
wire _23738_;
wire _23739_;
wire _23740_;
wire _23741_;
wire _23742_;
wire _23743_;
wire _23744_;
wire _23745_;
wire _23746_;
wire _23747_;
wire _23748_;
wire _23749_;
wire _23750_;
wire _23751_;
wire _23752_;
wire _23753_;
wire _23754_;
wire _23755_;
wire _23756_;
wire _23757_;
wire _23758_;
wire _23759_;
wire _23760_;
wire _23761_;
wire _23762_;
wire _23763_;
wire _23764_;
wire _23765_;
wire _23766_;
wire _23767_;
wire _23768_;
wire _23769_;
wire _23770_;
wire _23771_;
wire _23772_;
wire _23773_;
wire _23774_;
wire _23775_;
wire _23776_;
wire _23777_;
wire _23778_;
wire _23779_;
wire _23780_;
wire _23781_;
wire _23782_;
wire _23783_;
wire _23784_;
wire _23785_;
wire _23786_;
wire _23787_;
wire _23788_;
wire _23789_;
wire _23790_;
wire _23791_;
wire _23792_;
wire _23793_;
wire _23794_;
wire _23795_;
wire _23796_;
wire _23797_;
wire _23798_;
wire _23799_;
wire _23800_;
wire _23801_;
wire _23802_;
wire _23803_;
wire _23804_;
wire _23805_;
wire _23806_;
wire _23807_;
wire _23808_;
wire _23809_;
wire _23810_;
wire _23811_;
wire _23812_;
wire _23813_;
wire _23814_;
wire _23815_;
wire _23816_;
wire _23817_;
wire _23818_;
wire _23819_;
wire _23820_;
wire _23821_;
wire _23822_;
wire _23823_;
wire _23824_;
wire _23825_;
wire _23826_;
wire _23827_;
wire _23828_;
wire _23829_;
wire _23830_;
wire _23831_;
wire _23832_;
wire _23833_;
wire _23834_;
wire _23835_;
wire _23836_;
wire _23837_;
wire _23838_;
wire _23839_;
wire _23840_;
wire _23841_;
wire _23842_;
wire _23843_;
wire _23844_;
wire _23845_;
wire _23846_;
wire _23847_;
wire _23848_;
wire _23849_;
wire _23850_;
wire _23851_;
wire _23852_;
wire _23853_;
wire _23854_;
wire _23855_;
wire _23856_;
wire _23857_;
wire _23858_;
wire _23859_;
wire _23860_;
wire _23861_;
wire _23862_;
wire _23863_;
wire _23864_;
wire _23865_;
wire _23866_;
wire _23867_;
wire _23868_;
wire _23869_;
wire _23870_;
wire _23871_;
wire _23872_;
wire _23873_;
wire _23874_;
wire _23875_;
wire _23876_;
wire _23877_;
wire _23878_;
wire _23879_;
wire _23880_;
wire _23881_;
wire _23882_;
wire _23883_;
wire _23884_;
wire _23885_;
wire _23886_;
wire _23887_;
wire _23888_;
wire _23889_;
wire _23890_;
wire _23891_;
wire _23892_;
wire _23893_;
wire _23894_;
wire _23895_;
wire _23896_;
wire _23897_;
wire _23898_;
wire _23899_;
wire _23900_;
wire _23901_;
wire _23902_;
wire _23903_;
wire _23904_;
wire _23905_;
wire _23906_;
wire _23907_;
wire _23908_;
wire _23909_;
wire _23910_;
wire _23911_;
wire _23912_;
wire _23913_;
wire _23914_;
wire _23915_;
wire _23916_;
wire _23917_;
wire _23918_;
wire _23919_;
wire _23920_;
wire _23921_;
wire _23922_;
wire _23923_;
wire _23924_;
wire _23925_;
wire _23926_;
wire _23927_;
wire _23928_;
wire _23929_;
wire _23930_;
wire _23931_;
wire _23932_;
wire _23933_;
wire _23934_;
wire _23935_;
wire _23936_;
wire _23937_;
wire _23938_;
wire _23939_;
wire _23940_;
wire _23941_;
wire _23942_;
wire _23943_;
wire _23944_;
wire _23945_;
wire _23946_;
wire _23947_;
wire _23948_;
wire _23949_;
wire _23950_;
wire _23951_;
wire _23952_;
wire _23953_;
wire _23954_;
wire _23955_;
wire _23956_;
wire _23957_;
wire _23958_;
wire _23959_;
wire _23960_;
wire _23961_;
wire _23962_;
wire _23963_;
wire _23964_;
wire _23965_;
wire _23966_;
wire _23967_;
wire _23968_;
wire _23969_;
wire _23970_;
wire _23971_;
wire _23972_;
wire _23973_;
wire _23974_;
wire _23975_;
wire _23976_;
wire _23977_;
wire _23978_;
wire _23979_;
wire _23980_;
wire _23981_;
wire _23982_;
wire _23983_;
wire _23984_;
wire _23985_;
wire _23986_;
wire _23987_;
wire _23988_;
wire _23989_;
wire _23990_;
wire _23991_;
wire _23992_;
wire _23993_;
wire _23994_;
wire _23995_;
wire _23996_;
wire _23997_;
wire _23998_;
wire _23999_;
wire _24000_;
wire _24001_;
wire _24002_;
wire _24003_;
wire _24004_;
wire _24005_;
wire _24006_;
wire _24007_;
wire _24008_;
wire _24009_;
wire _24010_;
wire _24011_;
wire _24012_;
wire _24013_;
wire _24014_;
wire _24015_;
wire _24016_;
wire _24017_;
wire _24018_;
wire _24019_;
wire _24020_;
wire _24021_;
wire _24022_;
wire _24023_;
wire _24024_;
wire _24025_;
wire _24026_;
wire _24027_;
wire _24028_;
wire _24029_;
wire _24030_;
wire _24031_;
wire _24032_;
wire _24033_;
wire _24034_;
wire _24035_;
wire _24036_;
wire _24037_;
wire _24038_;
wire _24039_;
wire _24040_;
wire _24041_;
wire _24042_;
wire _24043_;
wire _24044_;
wire _24045_;
wire _24046_;
wire _24047_;
wire _24048_;
wire _24049_;
wire _24050_;
wire _24051_;
wire _24052_;
wire _24053_;
wire _24054_;
wire _24055_;
wire _24056_;
wire _24057_;
wire _24058_;
wire _24059_;
wire _24060_;
wire _24061_;
wire _24062_;
wire _24063_;
wire _24064_;
wire _24065_;
wire _24066_;
wire _24067_;
wire _24068_;
wire _24069_;
wire _24070_;
wire _24071_;
wire _24072_;
wire _24073_;
wire _24074_;
wire _24075_;
wire _24076_;
wire _24077_;
wire _24078_;
wire _24079_;
wire _24080_;
wire _24081_;
wire _24082_;
wire _24083_;
wire _24084_;
wire _24085_;
wire _24086_;
wire _24087_;
wire _24088_;
wire _24089_;
wire _24090_;
wire _24091_;
wire _24092_;
wire _24093_;
wire _24094_;
wire _24095_;
wire _24096_;
wire _24097_;
wire _24098_;
wire _24099_;
wire _24100_;
wire _24101_;
wire _24102_;
wire _24103_;
wire _24104_;
wire _24105_;
wire _24106_;
wire _24107_;
wire _24108_;
wire _24109_;
wire _24110_;
wire _24111_;
wire _24112_;
wire _24113_;
wire _24114_;
wire _24115_;
wire _24116_;
wire _24117_;
wire _24118_;
wire _24119_;
wire _24120_;
wire _24121_;
wire _24122_;
wire _24123_;
wire _24124_;
wire _24125_;
wire _24126_;
wire _24127_;
wire _24128_;
wire _24129_;
wire _24130_;
wire _24131_;
wire _24132_;
wire _24133_;
wire _24134_;
wire _24135_;
wire _24136_;
wire _24137_;
wire _24138_;
wire _24139_;
wire _24140_;
wire _24141_;
wire _24142_;
wire _24143_;
wire _24144_;
wire _24145_;
wire _24146_;
wire _24147_;
wire _24148_;
wire _24149_;
wire _24150_;
wire _24151_;
wire _24152_;
wire _24153_;
wire _24154_;
wire _24155_;
wire _24156_;
wire _24157_;
wire _24158_;
wire _24159_;
wire _24160_;
wire _24161_;
wire _24162_;
wire _24163_;
wire _24164_;
wire _24165_;
wire _24166_;
wire _24167_;
wire _24168_;
wire _24169_;
wire _24170_;
wire _24171_;
wire _24172_;
wire _24173_;
wire _24174_;
wire _24175_;
wire _24176_;
wire _24177_;
wire _24178_;
wire _24179_;
wire _24180_;
wire _24181_;
wire _24182_;
wire _24183_;
wire _24184_;
wire _24185_;
wire _24186_;
wire _24187_;
wire _24188_;
wire _24189_;
wire _24190_;
wire _24191_;
wire _24192_;
wire _24193_;
wire _24194_;
wire _24195_;
wire _24196_;
wire _24197_;
wire _24198_;
wire _24199_;
wire _24200_;
wire _24201_;
wire _24202_;
wire _24203_;
wire _24204_;
wire _24205_;
wire _24206_;
wire _24207_;
wire _24208_;
wire _24209_;
wire _24210_;
wire _24211_;
wire _24212_;
wire _24213_;
wire _24214_;
wire _24215_;
wire _24216_;
wire _24217_;
wire _24218_;
wire _24219_;
wire _24220_;
wire _24221_;
wire _24222_;
wire _24223_;
wire _24224_;
wire _24225_;
wire _24226_;
wire _24227_;
wire _24228_;
wire _24229_;
wire _24230_;
wire _24231_;
wire _24232_;
wire _24233_;
wire _24234_;
wire _24235_;
wire _24236_;
wire _24237_;
wire _24238_;
wire _24239_;
wire _24240_;
wire _24241_;
wire _24242_;
wire _24243_;
wire _24244_;
wire _24245_;
wire _24246_;
wire _24247_;
wire _24248_;
wire _24249_;
wire _24250_;
wire _24251_;
wire _24252_;
wire _24253_;
wire _24254_;
wire _24255_;
wire _24256_;
wire _24257_;
wire _24258_;
wire _24259_;
wire _24260_;
wire _24261_;
wire _24262_;
wire _24263_;
wire _24264_;
wire _24265_;
wire _24266_;
wire _24267_;
wire _24268_;
wire _24269_;
wire _24270_;
wire _24271_;
wire _24272_;
wire _24273_;
wire _24274_;
wire _24275_;
wire _24276_;
wire _24277_;
wire _24278_;
wire _24279_;
wire _24280_;
wire _24281_;
wire _24282_;
wire _24283_;
wire _24284_;
wire _24285_;
wire _24286_;
wire _24287_;
wire _24288_;
wire _24289_;
wire _24290_;
wire _24291_;
wire _24292_;
wire _24293_;
wire _24294_;
wire _24295_;
wire _24296_;
wire _24297_;
wire _24298_;
wire _24299_;
wire _24300_;
wire _24301_;
wire _24302_;
wire _24303_;
wire _24304_;
wire _24305_;
wire _24306_;
wire _24307_;
wire _24308_;
wire _24309_;
wire _24310_;
wire _24311_;
wire _24312_;
wire _24313_;
wire _24314_;
wire _24315_;
wire _24316_;
wire _24317_;
wire _24318_;
wire _24319_;
wire _24320_;
wire _24321_;
wire _24322_;
wire _24323_;
wire _24324_;
wire _24325_;
wire _24326_;
wire _24327_;
wire _24328_;
wire _24329_;
wire _24330_;
wire _24331_;
wire _24332_;
wire _24333_;
wire _24334_;
wire _24335_;
wire _24336_;
wire _24337_;
wire _24338_;
wire _24339_;
wire _24340_;
wire _24341_;
wire _24342_;
wire _24343_;
wire _24344_;
wire _24345_;
wire _24346_;
wire _24347_;
wire _24348_;
wire _24349_;
wire _24350_;
wire _24351_;
wire _24352_;
wire _24353_;
wire _24354_;
wire _24355_;
wire _24356_;
wire _24357_;
wire _24358_;
wire _24359_;
wire _24360_;
wire _24361_;
wire _24362_;
wire _24363_;
wire _24364_;
wire _24365_;
wire _24366_;
wire _24367_;
wire _24368_;
wire _24369_;
wire _24370_;
wire _24371_;
wire _24372_;
wire _24373_;
wire _24374_;
wire _24375_;
wire _24376_;
wire _24377_;
wire _24378_;
wire _24379_;
wire _24380_;
wire _24381_;
wire _24382_;
wire _24383_;
wire _24384_;
wire _24385_;
wire _24386_;
wire _24387_;
wire _24388_;
wire _24389_;
wire _24390_;
wire _24391_;
wire _24392_;
wire _24393_;
wire _24394_;
wire _24395_;
wire _24396_;
wire _24397_;
wire _24398_;
wire _24399_;
wire _24400_;
wire _24401_;
wire _24402_;
wire _24403_;
wire _24404_;
wire _24405_;
wire _24406_;
wire _24407_;
wire _24408_;
wire _24409_;
wire _24410_;
wire _24411_;
wire _24412_;
wire _24413_;
wire _24414_;
wire _24415_;
wire _24416_;
wire _24417_;
wire _24418_;
wire _24419_;
wire _24420_;
wire _24421_;
wire _24422_;
wire _24423_;
wire _24424_;
wire _24425_;
wire _24426_;
wire _24427_;
wire _24428_;
wire _24429_;
wire _24430_;
wire _24431_;
wire _24432_;
wire _24433_;
wire _24434_;
wire _24435_;
wire _24436_;
wire _24437_;
wire _24438_;
wire _24439_;
wire _24440_;
wire _24441_;
wire _24442_;
wire _24443_;
wire _24444_;
wire _24445_;
wire _24446_;
wire _24447_;
wire _24448_;
wire _24449_;
wire _24450_;
wire _24451_;
wire _24452_;
wire _24453_;
wire _24454_;
wire _24455_;
wire _24456_;
wire _24457_;
wire _24458_;
wire _24459_;
wire _24460_;
wire _24461_;
wire _24462_;
wire _24463_;
wire _24464_;
wire _24465_;
wire _24466_;
wire _24467_;
wire _24468_;
wire _24469_;
wire _24470_;
wire _24471_;
wire _24472_;
wire _24473_;
wire _24474_;
wire _24475_;
wire _24476_;
wire _24477_;
wire _24478_;
wire _24479_;
wire _24480_;
wire _24481_;
wire _24482_;
wire _24483_;
wire _24484_;
wire _24485_;
wire _24486_;
wire _24487_;
wire _24488_;
wire _24489_;
wire _24490_;
wire _24491_;
wire _24492_;
wire _24493_;
wire _24494_;
wire _24495_;
wire _24496_;
wire _24497_;
wire _24498_;
wire _24499_;
wire _24500_;
wire _24501_;
wire _24502_;
wire _24503_;
wire _24504_;
wire _24505_;
wire _24506_;
wire _24507_;
wire _24508_;
wire _24509_;
wire _24510_;
wire _24511_;
wire _24512_;
wire _24513_;
wire _24514_;
wire _24515_;
wire _24516_;
wire _24517_;
wire _24518_;
wire _24519_;
wire _24520_;
wire _24521_;
wire _24522_;
wire _24523_;
wire _24524_;
wire _24525_;
wire _24526_;
wire _24527_;
wire _24528_;
wire _24529_;
wire _24530_;
wire _24531_;
wire _24532_;
wire _24533_;
wire _24534_;
wire _24535_;
wire _24536_;
wire _24537_;
wire _24538_;
wire _24539_;
wire _24540_;
wire _24541_;
wire _24542_;
wire _24543_;
wire _24544_;
wire _24545_;
wire _24546_;
wire _24547_;
wire _24548_;
wire _24549_;
wire _24550_;
wire _24551_;
wire _24552_;
wire _24553_;
wire _24554_;
wire _24555_;
wire _24556_;
wire _24557_;
wire _24558_;
wire _24559_;
wire _24560_;
wire _24561_;
wire _24562_;
wire _24563_;
wire _24564_;
wire _24565_;
wire _24566_;
wire _24567_;
wire _24568_;
wire _24569_;
wire _24570_;
wire _24571_;
wire _24572_;
wire _24573_;
wire _24574_;
wire _24575_;
wire _24576_;
wire _24577_;
wire _24578_;
wire _24579_;
wire _24580_;
wire _24581_;
wire _24582_;
wire _24583_;
wire _24584_;
wire _24585_;
wire _24586_;
wire _24587_;
wire _24588_;
wire _24589_;
wire _24590_;
wire _24591_;
wire _24592_;
wire _24593_;
wire _24594_;
wire _24595_;
wire _24596_;
wire _24597_;
wire _24598_;
wire _24599_;
wire _24600_;
wire _24601_;
wire _24602_;
wire _24603_;
wire _24604_;
wire _24605_;
wire _24606_;
wire _24607_;
wire _24608_;
wire _24609_;
wire _24610_;
wire _24611_;
wire _24612_;
wire _24613_;
wire _24614_;
wire _24615_;
wire _24616_;
wire _24617_;
wire _24618_;
wire _24619_;
wire _24620_;
wire _24621_;
wire _24622_;
wire _24623_;
wire _24624_;
wire _24625_;
wire _24626_;
wire _24627_;
wire _24628_;
wire _24629_;
wire _24630_;
wire _24631_;
wire _24632_;
wire _24633_;
wire _24634_;
wire _24635_;
wire _24636_;
wire _24637_;
wire _24638_;
wire _24639_;
wire _24640_;
wire _24641_;
wire _24642_;
wire _24643_;
wire _24644_;
wire _24645_;
wire _24646_;
wire _24647_;
wire _24648_;
wire _24649_;
wire _24650_;
wire _24651_;
wire _24652_;
wire _24653_;
wire _24654_;
wire _24655_;
wire _24656_;
wire _24657_;
wire _24658_;
wire _24659_;
wire _24660_;
wire _24661_;
wire _24662_;
wire _24663_;
wire _24664_;
wire _24665_;
wire _24666_;
wire _24667_;
wire _24668_;
wire _24669_;
wire _24670_;
wire _24671_;
wire _24672_;
wire _24673_;
wire _24674_;
wire _24675_;
wire _24676_;
wire _24677_;
wire _24678_;
wire _24679_;
wire _24680_;
wire _24681_;
wire _24682_;
wire _24683_;
wire _24684_;
wire _24685_;
wire _24686_;
wire _24687_;
wire _24688_;
wire _24689_;
wire _24690_;
wire _24691_;
wire _24692_;
wire _24693_;
wire _24694_;
wire _24695_;
wire _24696_;
wire _24697_;
wire _24698_;
wire _24699_;
wire _24700_;
wire _24701_;
wire _24702_;
wire _24703_;
wire _24704_;
wire _24705_;
wire _24706_;
wire _24707_;
wire _24708_;
wire _24709_;
wire _24710_;
wire _24711_;
wire _24712_;
wire _24713_;
wire _24714_;
wire _24715_;
wire _24716_;
wire _24717_;
wire _24718_;
wire _24719_;
wire _24720_;
wire _24721_;
wire _24722_;
wire _24723_;
wire _24724_;
wire _24725_;
wire _24726_;
wire _24727_;
wire _24728_;
wire _24729_;
wire _24730_;
wire _24731_;
wire _24732_;
wire _24733_;
wire _24734_;
wire _24735_;
wire _24736_;
wire _24737_;
wire _24738_;
wire _24739_;
wire _24740_;
wire _24741_;
wire _24742_;
wire _24743_;
wire _24744_;
wire _24745_;
wire _24746_;
wire _24747_;
wire _24748_;
wire _24749_;
wire _24750_;
wire _24751_;
wire _24752_;
wire _24753_;
wire _24754_;
wire _24755_;
wire _24756_;
wire _24757_;
wire _24758_;
wire _24759_;
wire _24760_;
wire _24761_;
wire _24762_;
wire _24763_;
wire _24764_;
wire _24765_;
wire _24766_;
wire _24767_;
wire _24768_;
wire _24769_;
wire _24770_;
wire _24771_;
wire _24772_;
wire _24773_;
wire _24774_;
wire _24775_;
wire _24776_;
wire _24777_;
wire _24778_;
wire _24779_;
wire _24780_;
wire _24781_;
wire _24782_;
wire _24783_;
wire _24784_;
wire _24785_;
wire _24786_;
wire _24787_;
wire _24788_;
wire _24789_;
wire _24790_;
wire _24791_;
wire _24792_;
wire _24793_;
wire _24794_;
wire _24795_;
wire _24796_;
wire _24797_;
wire _24798_;
wire _24799_;
wire _24800_;
wire _24801_;
wire _24802_;
wire _24803_;
wire _24804_;
wire _24805_;
wire _24806_;
wire _24807_;
wire _24808_;
wire _24809_;
wire _24810_;
wire _24811_;
wire _24812_;
wire _24813_;
wire _24814_;
wire _24815_;
wire _24816_;
wire _24817_;
wire _24818_;
wire _24819_;
wire _24820_;
wire _24821_;
wire _24822_;
wire _24823_;
wire _24824_;
wire _24825_;
wire _24826_;
wire _24827_;
wire _24828_;
wire _24829_;
wire _24830_;
wire _24831_;
wire _24832_;
wire _24833_;
wire _24834_;
wire _24835_;
wire _24836_;
wire _24837_;
wire _24838_;
wire _24839_;
wire _24840_;
wire _24841_;
wire _24842_;
wire _24843_;
wire _24844_;
wire _24845_;
wire _24846_;
wire _24847_;
wire _24848_;
wire _24849_;
wire _24850_;
wire _24851_;
wire _24852_;
wire _24853_;
wire _24854_;
wire _24855_;
wire _24856_;
wire _24857_;
wire _24858_;
wire _24859_;
wire _24860_;
wire _24861_;
wire _24862_;
wire _24863_;
wire _24864_;
wire _24865_;
wire _24866_;
wire _24867_;
wire _24868_;
wire _24869_;
wire _24870_;
wire _24871_;
wire _24872_;
wire _24873_;
wire _24874_;
wire _24875_;
wire _24876_;
wire _24877_;
wire _24878_;
wire _24879_;
wire _24880_;
wire _24881_;
wire _24882_;
wire _24883_;
wire _24884_;
wire _24885_;
wire _24886_;
wire _24887_;
wire _24888_;
wire _24889_;
wire _24890_;
wire _24891_;
wire _24892_;
wire _24893_;
wire _24894_;
wire _24895_;
wire _24896_;
wire _24897_;
wire _24898_;
wire _24899_;
wire _24900_;
wire _24901_;
wire _24902_;
wire _24903_;
wire _24904_;
wire _24905_;
wire _24906_;
wire _24907_;
wire _24908_;
wire _24909_;
wire _24910_;
wire _24911_;
wire _24912_;
wire _24913_;
wire _24914_;
wire _24915_;
wire _24916_;
wire _24917_;
wire _24918_;
wire _24919_;
wire _24920_;
wire _24921_;
wire _24922_;
wire _24923_;
wire _24924_;
wire _24925_;
wire _24926_;
wire _24927_;
wire _24928_;
wire _24929_;
wire _24930_;
wire _24931_;
wire _24932_;
wire _24933_;
wire _24934_;
wire _24935_;
wire _24936_;
wire _24937_;
wire _24938_;
wire _24939_;
wire _24940_;
wire _24941_;
wire _24942_;
wire _24943_;
wire _24944_;
wire _24945_;
wire _24946_;
wire _24947_;
wire _24948_;
wire _24949_;
wire _24950_;
wire _24951_;
wire _24952_;
wire _24953_;
wire _24954_;
wire _24955_;
wire _24956_;
wire _24957_;
wire _24958_;
wire _24959_;
wire _24960_;
wire _24961_;
wire _24962_;
wire _24963_;
wire _24964_;
wire _24965_;
wire _24966_;
wire _24967_;
wire _24968_;
wire _24969_;
wire _24970_;
wire _24971_;
wire _24972_;
wire _24973_;
wire _24974_;
wire _24975_;
wire _24976_;
wire _24977_;
wire _24978_;
wire _24979_;
wire _24980_;
wire _24981_;
wire _24982_;
wire _24983_;
wire _24984_;
wire _24985_;
wire _24986_;
wire _24987_;
wire _24988_;
wire _24989_;
wire _24990_;
wire _24991_;
wire _24992_;
wire _24993_;
wire _24994_;
wire _24995_;
wire _24996_;
wire _24997_;
wire _24998_;
wire _24999_;
wire _25000_;
wire _25001_;
wire _25002_;
wire _25003_;
wire _25004_;
wire _25005_;
wire _25006_;
wire _25007_;
wire _25008_;
wire _25009_;
wire _25010_;
wire _25011_;
wire _25012_;
wire _25013_;
wire _25014_;
wire _25015_;
wire _25016_;
wire _25017_;
wire _25018_;
wire _25019_;
wire _25020_;
wire _25021_;
wire _25022_;
wire _25023_;
wire _25024_;
wire _25025_;
wire _25026_;
wire _25027_;
wire _25028_;
wire _25029_;
wire _25030_;
wire _25031_;
wire _25032_;
wire _25033_;
wire _25034_;
wire _25035_;
wire _25036_;
wire _25037_;
wire _25038_;
wire _25039_;
wire _25040_;
wire _25041_;
wire _25042_;
wire _25043_;
wire _25044_;
wire _25045_;
wire _25046_;
wire _25047_;
wire _25048_;
wire _25049_;
wire _25050_;
wire _25051_;
wire _25052_;
wire _25053_;
wire _25054_;
wire _25055_;
wire _25056_;
wire _25057_;
wire _25058_;
wire _25059_;
wire _25060_;
wire _25061_;
wire _25062_;
wire _25063_;
wire _25064_;
wire _25065_;
wire _25066_;
wire _25067_;
wire _25068_;
wire _25069_;
wire _25070_;
wire _25071_;
wire _25072_;
wire _25073_;
wire _25074_;
wire _25075_;
wire _25076_;
wire _25077_;
wire _25078_;
wire _25079_;
wire _25080_;
wire _25081_;
wire _25082_;
wire _25083_;
wire _25084_;
wire _25085_;
wire _25086_;
wire _25087_;
wire _25088_;
wire _25089_;
wire _25090_;
wire _25091_;
wire _25092_;
wire _25093_;
wire _25094_;
wire _25095_;
wire _25096_;
wire _25097_;
wire _25098_;
wire _25099_;
wire _25100_;
wire _25101_;
wire _25102_;
wire _25103_;
wire _25104_;
wire _25105_;
wire _25106_;
wire _25107_;
wire _25108_;
wire _25109_;
wire _25110_;
wire _25111_;
wire _25112_;
wire _25113_;
wire _25114_;
wire _25115_;
wire _25116_;
wire _25117_;
wire _25118_;
wire _25119_;
wire _25120_;
wire _25121_;
wire _25122_;
wire _25123_;
wire _25124_;
wire _25125_;
wire _25126_;
wire _25127_;
wire _25128_;
wire _25129_;
wire _25130_;
wire _25131_;
wire _25132_;
wire _25133_;
wire _25134_;
wire _25135_;
wire _25136_;
wire _25137_;
wire _25138_;
wire _25139_;
wire _25140_;
wire _25141_;
wire _25142_;
wire _25143_;
wire _25144_;
wire _25145_;
wire _25146_;
wire _25147_;
wire _25148_;
wire _25149_;
wire _25150_;
wire _25151_;
wire _25152_;
wire _25153_;
wire _25154_;
wire _25155_;
wire _25156_;
wire _25157_;
wire _25158_;
wire _25159_;
wire _25160_;
wire _25161_;
wire _25162_;
wire _25163_;
wire _25164_;
wire _25165_;
wire _25166_;
wire _25167_;
wire _25168_;
wire _25169_;
wire _25170_;
wire _25171_;
wire _25172_;
wire _25173_;
wire _25174_;
wire _25175_;
wire _25176_;
wire _25177_;
wire _25178_;
wire _25179_;
wire _25180_;
wire _25181_;
wire _25182_;
wire _25183_;
wire _25184_;
wire _25185_;
wire _25186_;
wire _25187_;
wire _25188_;
wire _25189_;
wire _25190_;
wire _25191_;
wire _25192_;
wire _25193_;
wire _25194_;
wire _25195_;
wire _25196_;
wire _25197_;
wire _25198_;
wire _25199_;
wire _25200_;
wire _25201_;
wire _25202_;
wire _25203_;
wire _25204_;
wire _25205_;
wire _25206_;
wire _25207_;
wire _25208_;
wire _25209_;
wire _25210_;
wire _25211_;
wire _25212_;
wire _25213_;
wire _25214_;
wire _25215_;
wire _25216_;
wire _25217_;
wire _25218_;
wire _25219_;
wire _25220_;
wire _25221_;
wire _25222_;
wire _25223_;
wire _25224_;
wire _25225_;
wire _25226_;
wire _25227_;
wire _25228_;
wire _25229_;
wire _25230_;
wire _25231_;
wire _25232_;
wire _25233_;
wire _25234_;
wire _25235_;
wire _25236_;
wire _25237_;
wire _25238_;
wire _25239_;
wire _25240_;
wire _25241_;
wire _25242_;
wire _25243_;
wire _25244_;
wire _25245_;
wire _25246_;
wire _25247_;
wire _25248_;
wire _25249_;
wire _25250_;
wire _25251_;
wire _25252_;
wire _25253_;
wire _25254_;
wire _25255_;
wire _25256_;
wire _25257_;
wire _25258_;
wire _25259_;
wire _25260_;
wire _25261_;
wire _25262_;
wire _25263_;
wire _25264_;
wire _25265_;
wire _25266_;
wire _25267_;
wire _25268_;
wire _25269_;
wire _25270_;
wire _25271_;
wire _25272_;
wire _25273_;
wire _25274_;
wire _25275_;
wire _25276_;
wire _25277_;
wire _25278_;
wire _25279_;
wire _25280_;
wire _25281_;
wire _25282_;
wire _25283_;
wire _25284_;
wire _25285_;
wire _25286_;
wire _25287_;
wire _25288_;
wire _25289_;
wire _25290_;
wire _25291_;
wire _25292_;
wire _25293_;
wire _25294_;
wire _25295_;
wire _25296_;
wire _25297_;
wire _25298_;
wire _25299_;
wire _25300_;
wire _25301_;
wire _25302_;
wire _25303_;
wire _25304_;
wire _25305_;
wire _25306_;
wire _25307_;
wire _25308_;
wire _25309_;
wire _25310_;
wire _25311_;
wire _25312_;
wire _25313_;
wire _25314_;
wire _25315_;
wire _25316_;
wire _25317_;
wire _25318_;
wire _25319_;
wire _25320_;
wire _25321_;
wire _25322_;
wire _25323_;
wire _25324_;
wire _25325_;
wire _25326_;
wire _25327_;
wire _25328_;
wire _25329_;
wire _25330_;
wire _25331_;
wire _25332_;
wire _25333_;
wire _25334_;
wire _25335_;
wire _25336_;
wire _25337_;
wire _25338_;
wire _25339_;
wire _25340_;
wire _25341_;
wire _25342_;
wire _25343_;
wire _25344_;
wire _25345_;
wire _25346_;
wire _25347_;
wire _25348_;
wire _25349_;
wire _25350_;
wire _25351_;
wire _25352_;
wire _25353_;
wire _25354_;
wire _25355_;
wire _25356_;
wire _25357_;
wire _25358_;
wire _25359_;
wire _25360_;
wire _25361_;
wire _25362_;
wire _25363_;
wire _25364_;
wire _25365_;
wire _25366_;
wire _25367_;
wire _25368_;
wire _25369_;
wire _25370_;
wire _25371_;
wire _25372_;
wire _25373_;
wire _25374_;
wire _25375_;
wire _25376_;
wire _25377_;
wire _25378_;
wire _25379_;
wire _25380_;
wire _25381_;
wire _25382_;
wire _25383_;
wire _25384_;
wire _25385_;
wire _25386_;
wire _25387_;
wire _25388_;
wire _25389_;
wire _25390_;
wire _25391_;
wire _25392_;
wire _25393_;
wire _25394_;
wire _25395_;
wire _25396_;
wire _25397_;
wire _25398_;
wire _25399_;
wire _25400_;
wire _25401_;
wire _25402_;
wire _25403_;
wire _25404_;
wire _25405_;
wire _25406_;
wire _25407_;
wire _25408_;
wire _25409_;
wire _25410_;
wire _25411_;
wire _25412_;
wire _25413_;
wire _25414_;
wire _25415_;
wire _25416_;
wire _25417_;
wire _25418_;
wire _25419_;
wire _25420_;
wire _25421_;
wire _25422_;
wire _25423_;
wire _25424_;
wire _25425_;
wire _25426_;
wire _25427_;
wire _25428_;
wire _25429_;
wire _25430_;
wire _25431_;
wire _25432_;
wire _25433_;
wire _25434_;
wire _25435_;
wire _25436_;
wire _25437_;
wire _25438_;
wire _25439_;
wire _25440_;
wire _25441_;
wire _25442_;
wire _25443_;
wire _25444_;
wire _25445_;
wire _25446_;
wire _25447_;
wire _25448_;
wire _25449_;
wire _25450_;
wire _25451_;
wire _25452_;
wire _25453_;
wire _25454_;
wire _25455_;
wire _25456_;
wire _25457_;
wire _25458_;
wire _25459_;
wire _25460_;
wire _25461_;
wire _25462_;
wire _25463_;
wire _25464_;
wire _25465_;
wire _25466_;
wire _25467_;
wire _25468_;
wire _25469_;
wire _25470_;
wire _25471_;
wire _25472_;
wire _25473_;
wire _25474_;
wire _25475_;
wire _25476_;
wire _25477_;
wire _25478_;
wire _25479_;
wire _25480_;
wire _25481_;
wire _25482_;
wire _25483_;
wire _25484_;
wire _25485_;
wire _25486_;
wire _25487_;
wire _25488_;
wire _25489_;
wire _25490_;
wire _25491_;
wire _25492_;
wire _25493_;
wire _25494_;
wire _25495_;
wire _25496_;
wire _25497_;
wire _25498_;
wire _25499_;
wire _25500_;
wire _25501_;
wire _25502_;
wire _25503_;
wire _25504_;
wire _25505_;
wire _25506_;
wire _25507_;
wire _25508_;
wire _25509_;
wire _25510_;
wire _25511_;
wire _25512_;
wire _25513_;
wire _25514_;
wire _25515_;
wire _25516_;
wire _25517_;
wire _25518_;
wire _25519_;
wire _25520_;
wire _25521_;
wire _25522_;
wire _25523_;
wire _25524_;
wire _25525_;
wire _25526_;
wire _25527_;
wire _25528_;
wire _25529_;
wire _25530_;
wire _25531_;
wire _25532_;
wire _25533_;
wire _25534_;
wire _25535_;
wire _25536_;
wire _25537_;
wire _25538_;
wire _25539_;
wire _25540_;
wire _25541_;
wire _25542_;
wire _25543_;
wire _25544_;
wire _25545_;
wire _25546_;
wire _25547_;
wire _25548_;
wire _25549_;
wire _25550_;
wire _25551_;
wire _25552_;
wire _25553_;
wire _25554_;
wire _25555_;
wire _25556_;
wire _25557_;
wire _25558_;
wire _25559_;
wire _25560_;
wire _25561_;
wire _25562_;
wire _25563_;
wire _25564_;
wire _25565_;
wire _25566_;
wire _25567_;
wire _25568_;
wire _25569_;
wire _25570_;
wire _25571_;
wire _25572_;
wire _25573_;
wire _25574_;
wire _25575_;
wire _25576_;
wire _25577_;
wire _25578_;
wire _25579_;
wire _25580_;
wire _25581_;
wire _25582_;
wire _25583_;
wire _25584_;
wire _25585_;
wire _25586_;
wire _25587_;
wire _25588_;
wire _25589_;
wire _25590_;
wire _25591_;
wire _25592_;
wire _25593_;
wire _25594_;
wire _25595_;
wire _25596_;
wire _25597_;
wire _25598_;
wire _25599_;
wire _25600_;
wire _25601_;
wire _25602_;
wire _25603_;
wire _25604_;
wire _25605_;
wire _25606_;
wire _25607_;
wire _25608_;
wire _25609_;
wire _25610_;
wire _25611_;
wire _25612_;
wire _25613_;
wire _25614_;
wire _25615_;
wire _25616_;
wire _25617_;
wire _25618_;
wire _25619_;
wire _25620_;
wire _25621_;
wire _25622_;
wire _25623_;
wire _25624_;
wire _25625_;
wire _25626_;
wire _25627_;
wire _25628_;
wire _25629_;
wire _25630_;
wire _25631_;
wire _25632_;
wire _25633_;
wire _25634_;
wire _25635_;
wire _25636_;
wire _25637_;
wire _25638_;
wire _25639_;
wire _25640_;
wire _25641_;
wire _25642_;
wire _25643_;
wire _25644_;
wire _25645_;
wire _25646_;
wire _25647_;
wire _25648_;
wire _25649_;
wire _25650_;
wire _25651_;
wire _25652_;
wire _25653_;
wire _25654_;
wire _25655_;
wire _25656_;
wire _25657_;
wire _25658_;
wire _25659_;
wire _25660_;
wire _25661_;
wire _25662_;
wire _25663_;
wire _25664_;
wire _25665_;
wire _25666_;
wire _25667_;
wire _25668_;
wire _25669_;
wire _25670_;
wire _25671_;
wire _25672_;
wire _25673_;
wire _25674_;
wire _25675_;
wire _25676_;
wire _25677_;
wire _25678_;
wire _25679_;
wire _25680_;
wire _25681_;
wire _25682_;
wire _25683_;
wire _25684_;
wire _25685_;
wire _25686_;
wire _25687_;
wire _25688_;
wire _25689_;
wire _25690_;
wire _25691_;
wire _25692_;
wire _25693_;
wire _25694_;
wire _25695_;
wire _25696_;
wire _25697_;
wire _25698_;
wire _25699_;
wire _25700_;
wire _25701_;
wire _25702_;
wire _25703_;
wire _25704_;
wire _25705_;
wire _25706_;
wire _25707_;
wire _25708_;
wire _25709_;
wire _25710_;
wire _25711_;
wire _25712_;
wire _25713_;
wire _25714_;
wire _25715_;
wire _25716_;
wire _25717_;
wire _25718_;
wire _25719_;
wire _25720_;
wire _25721_;
wire _25722_;
wire _25723_;
wire _25724_;
wire _25725_;
wire _25726_;
wire _25727_;
wire _25728_;
wire _25729_;
wire _25730_;
wire _25731_;
wire _25732_;
wire _25733_;
wire _25734_;
wire _25735_;
wire _25736_;
wire _25737_;
wire _25738_;
wire _25739_;
wire _25740_;
wire _25741_;
wire _25742_;
wire _25743_;
wire _25744_;
wire _25745_;
wire _25746_;
wire _25747_;
wire _25748_;
wire _25749_;
wire _25750_;
wire _25751_;
wire _25752_;
wire _25753_;
wire _25754_;
wire _25755_;
wire _25756_;
wire _25757_;
wire _25758_;
wire _25759_;
wire _25760_;
wire _25761_;
wire _25762_;
wire _25763_;
wire _25764_;
wire _25765_;
wire _25766_;
wire _25767_;
wire _25768_;
wire _25769_;
wire _25770_;
wire _25771_;
wire _25772_;
wire _25773_;
wire _25774_;
wire _25775_;
wire _25776_;
wire _25777_;
wire _25778_;
wire _25779_;
wire _25780_;
wire _25781_;
wire _25782_;
wire _25783_;
wire _25784_;
wire _25785_;
wire _25786_;
wire _25787_;
wire _25788_;
wire _25789_;
wire _25790_;
wire _25791_;
wire _25792_;
wire _25793_;
wire _25794_;
wire _25795_;
wire _25796_;
wire _25797_;
wire _25798_;
wire _25799_;
wire _25800_;
wire _25801_;
wire _25802_;
wire _25803_;
wire _25804_;
wire _25805_;
wire _25806_;
wire _25807_;
wire _25808_;
wire _25809_;
wire _25810_;
wire _25811_;
wire _25812_;
wire _25813_;
wire _25814_;
wire _25815_;
wire _25816_;
wire _25817_;
wire _25818_;
wire _25819_;
wire _25820_;
wire _25821_;
wire _25822_;
wire _25823_;
wire _25824_;
wire _25825_;
wire _25826_;
wire _25827_;
wire _25828_;
wire _25829_;
wire _25830_;
wire _25831_;
wire _25832_;
wire _25833_;
wire _25834_;
wire _25835_;
wire _25836_;
wire _25837_;
wire _25838_;
wire _25839_;
wire _25840_;
wire _25841_;
wire _25842_;
wire _25843_;
wire _25844_;
wire _25845_;
wire _25846_;
wire _25847_;
wire _25848_;
wire _25849_;
wire _25850_;
wire _25851_;
wire _25852_;
wire _25853_;
wire _25854_;
wire _25855_;
wire _25856_;
wire _25857_;
wire _25858_;
wire _25859_;
wire _25860_;
wire _25861_;
wire _25862_;
wire _25863_;
wire _25864_;
wire _25865_;
wire _25866_;
wire _25867_;
wire _25868_;
wire _25869_;
wire _25870_;
wire _25871_;
wire _25872_;
wire _25873_;
wire _25874_;
wire _25875_;
wire _25876_;
wire _25877_;
wire _25878_;
wire _25879_;
wire _25880_;
wire _25881_;
wire _25882_;
wire _25883_;
wire _25884_;
wire _25885_;
wire _25886_;
wire _25887_;
wire _25888_;
wire _25889_;
wire _25890_;
wire _25891_;
wire _25892_;
wire _25893_;
wire _25894_;
wire _25895_;
wire _25896_;
wire _25897_;
wire _25898_;
wire _25899_;
wire _25900_;
wire _25901_;
wire _25902_;
wire _25903_;
wire _25904_;
wire _25905_;
wire _25906_;
wire _25907_;
wire _25908_;
wire _25909_;
wire _25910_;
wire _25911_;
wire _25912_;
wire _25913_;
wire _25914_;
wire _25915_;
wire _25916_;
wire _25917_;
wire _25918_;
wire _25919_;
wire _25920_;
wire _25921_;
wire _25922_;
wire _25923_;
wire _25924_;
wire _25925_;
wire _25926_;
wire _25927_;
wire _25928_;
wire _25929_;
wire _25930_;
wire _25931_;
wire _25932_;
wire _25933_;
wire _25934_;
wire _25935_;
wire _25936_;
wire _25937_;
wire _25938_;
wire _25939_;
wire _25940_;
wire _25941_;
wire _25942_;
wire _25943_;
wire _25944_;
wire _25945_;
wire _25946_;
wire _25947_;
wire _25948_;
wire _25949_;
wire _25950_;
wire _25951_;
wire _25952_;
wire _25953_;
wire _25954_;
wire _25955_;
wire _25956_;
wire _25957_;
wire _25958_;
wire _25959_;
wire _25960_;
wire _25961_;
wire _25962_;
wire _25963_;
wire _25964_;
wire _25965_;
wire _25966_;
wire _25967_;
wire _25968_;
wire _25969_;
wire _25970_;
wire _25971_;
wire _25972_;
wire _25973_;
wire _25974_;
wire _25975_;
wire _25976_;
wire _25977_;
wire _25978_;
wire _25979_;
wire _25980_;
wire _25981_;
wire _25982_;
wire _25983_;
wire _25984_;
wire _25985_;
wire _25986_;
wire _25987_;
wire _25988_;
wire _25989_;
wire _25990_;
wire _25991_;
wire _25992_;
wire _25993_;
wire _25994_;
wire _25995_;
wire _25996_;
wire _25997_;
wire _25998_;
wire _25999_;
wire _26000_;
wire _26001_;
wire _26002_;
wire _26003_;
wire _26004_;
wire _26005_;
wire _26006_;
wire _26007_;
wire _26008_;
wire _26009_;
wire _26010_;
wire _26011_;
wire _26012_;
wire _26013_;
wire _26014_;
wire _26015_;
wire _26016_;
wire _26017_;
wire _26018_;
wire _26019_;
wire _26020_;
wire _26021_;
wire _26022_;
wire _26023_;
wire _26024_;
wire _26025_;
wire _26026_;
wire _26027_;
wire _26028_;
wire _26029_;
wire _26030_;
wire _26031_;
wire _26032_;
wire _26033_;
wire _26034_;
wire _26035_;
wire _26036_;
wire _26037_;
wire _26038_;
wire _26039_;
wire _26040_;
wire _26041_;
wire _26042_;
wire _26043_;
wire _26044_;
wire _26045_;
wire _26046_;
wire _26047_;
wire _26048_;
wire _26049_;
wire _26050_;
wire _26051_;
wire _26052_;
wire _26053_;
wire _26054_;
wire _26055_;
wire _26056_;
wire _26057_;
wire _26058_;
wire _26059_;
wire _26060_;
wire _26061_;
wire _26062_;
wire _26063_;
wire _26064_;
wire _26065_;
wire _26066_;
wire _26067_;
wire _26068_;
wire _26069_;
wire _26070_;
wire _26071_;
wire _26072_;
wire _26073_;
wire _26074_;
wire _26075_;
wire _26076_;
wire _26077_;
wire _26078_;
wire _26079_;
wire _26080_;
wire _26081_;
wire _26082_;
wire _26083_;
wire _26084_;
wire _26085_;
wire _26086_;
wire _26087_;
wire _26088_;
wire _26089_;
wire _26090_;
wire _26091_;
wire _26092_;
wire _26093_;
wire _26094_;
wire _26095_;
wire _26096_;
wire _26097_;
wire _26098_;
wire _26099_;
wire _26100_;
wire _26101_;
wire _26102_;
wire _26103_;
wire _26104_;
wire _26105_;
wire _26106_;
wire _26107_;
wire _26108_;
wire _26109_;
wire _26110_;
wire _26111_;
wire _26112_;
wire _26113_;
wire _26114_;
wire _26115_;
wire _26116_;
wire _26117_;
wire _26118_;
wire _26119_;
wire _26120_;
wire _26121_;
wire _26122_;
wire _26123_;
wire _26124_;
wire _26125_;
wire _26126_;
wire _26127_;
wire _26128_;
wire _26129_;
wire _26130_;
wire _26131_;
wire _26132_;
wire _26133_;
wire _26134_;
wire _26135_;
wire _26136_;
wire _26137_;
wire _26138_;
wire _26139_;
wire _26140_;
wire _26141_;
wire _26142_;
wire _26143_;
wire _26144_;
wire _26145_;
wire _26146_;
wire _26147_;
wire _26148_;
wire _26149_;
wire _26150_;
wire _26151_;
wire _26152_;
wire _26153_;
wire _26154_;
wire _26155_;
wire _26156_;
wire _26157_;
wire _26158_;
wire _26159_;
wire _26160_;
wire _26161_;
wire _26162_;
wire _26163_;
wire _26164_;
wire _26165_;
wire _26166_;
wire _26167_;
wire _26168_;
wire _26169_;
wire _26170_;
wire _26171_;
wire _26172_;
wire _26173_;
wire _26174_;
wire _26175_;
wire _26176_;
wire _26177_;
wire _26178_;
wire _26179_;
wire _26180_;
wire _26181_;
wire _26182_;
wire _26183_;
wire _26184_;
wire _26185_;
wire _26186_;
wire _26187_;
wire _26188_;
wire _26189_;
wire _26190_;
wire _26191_;
wire _26192_;
wire _26193_;
wire _26194_;
wire _26195_;
wire _26196_;
wire _26197_;
wire _26198_;
wire _26199_;
wire _26200_;
wire _26201_;
wire _26202_;
wire _26203_;
wire _26204_;
wire _26205_;
wire _26206_;
wire _26207_;
wire _26208_;
wire _26209_;
wire _26210_;
wire _26211_;
wire _26212_;
wire _26213_;
wire _26214_;
wire _26215_;
wire _26216_;
wire _26217_;
wire _26218_;
wire _26219_;
wire _26220_;
wire _26221_;
wire _26222_;
wire _26223_;
wire _26224_;
wire _26225_;
wire _26226_;
wire _26227_;
wire _26228_;
wire _26229_;
wire _26230_;
wire _26231_;
wire _26232_;
wire _26233_;
wire _26234_;
wire _26235_;
wire _26236_;
wire _26237_;
wire _26238_;
wire _26239_;
wire _26240_;
wire _26241_;
wire _26242_;
wire _26243_;
wire _26244_;
wire _26245_;
wire _26246_;
wire _26247_;
wire _26248_;
wire _26249_;
wire _26250_;
wire _26251_;
wire _26252_;
wire _26253_;
wire _26254_;
wire _26255_;
wire _26256_;
wire _26257_;
wire _26258_;
wire _26259_;
wire _26260_;
wire _26261_;
wire _26262_;
wire _26263_;
wire _26264_;
wire _26265_;
wire _26266_;
wire _26267_;
wire _26268_;
wire _26269_;
wire _26270_;
wire _26271_;
wire _26272_;
wire _26273_;
wire _26274_;
wire _26275_;
wire _26276_;
wire _26277_;
wire _26278_;
wire _26279_;
wire _26280_;
wire _26281_;
wire _26282_;
wire _26283_;
wire _26284_;
wire _26285_;
wire _26286_;
wire _26287_;
wire _26288_;
wire _26289_;
wire _26290_;
wire _26291_;
wire _26292_;
wire _26293_;
wire _26294_;
wire _26295_;
wire _26296_;
wire _26297_;
wire _26298_;
wire _26299_;
wire _26300_;
wire _26301_;
wire _26302_;
wire _26303_;
wire _26304_;
wire _26305_;
wire _26306_;
wire _26307_;
wire _26308_;
wire _26309_;
wire _26310_;
wire _26311_;
wire _26312_;
wire _26313_;
wire _26314_;
wire _26315_;
wire _26316_;
wire _26317_;
wire _26318_;
wire _26319_;
wire _26320_;
wire _26321_;
wire _26322_;
wire _26323_;
wire _26324_;
wire _26325_;
wire _26326_;
wire _26327_;
wire _26328_;
wire _26329_;
wire _26330_;
wire _26331_;
wire _26332_;
wire _26333_;
wire _26334_;
wire _26335_;
wire _26336_;
wire _26337_;
wire _26338_;
wire _26339_;
wire _26340_;
wire _26341_;
wire _26342_;
wire _26343_;
wire _26344_;
wire _26345_;
wire _26346_;
wire _26347_;
wire _26348_;
wire _26349_;
wire _26350_;
wire _26351_;
wire _26352_;
wire _26353_;
wire _26354_;
wire _26355_;
wire _26356_;
wire _26357_;
wire _26358_;
wire _26359_;
wire _26360_;
wire _26361_;
wire _26362_;
wire _26363_;
wire _26364_;
wire _26365_;
wire _26366_;
wire _26367_;
wire _26368_;
wire _26369_;
wire _26370_;
wire _26371_;
wire _26372_;
wire _26373_;
wire _26374_;
wire _26375_;
wire _26376_;
wire _26377_;
wire _26378_;
wire _26379_;
wire _26380_;
wire _26381_;
wire _26382_;
wire _26383_;
wire _26384_;
wire _26385_;
wire _26386_;
wire _26387_;
wire _26388_;
wire _26389_;
wire _26390_;
wire _26391_;
wire _26392_;
wire _26393_;
wire _26394_;
wire _26395_;
wire _26396_;
wire _26397_;
wire _26398_;
wire _26399_;
wire _26400_;
wire _26401_;
wire _26402_;
wire _26403_;
wire _26404_;
wire _26405_;
wire _26406_;
wire _26407_;
wire _26408_;
wire _26409_;
wire _26410_;
wire _26411_;
wire _26412_;
wire _26413_;
wire _26414_;
wire _26415_;
wire _26416_;
wire _26417_;
wire _26418_;
wire _26419_;
wire _26420_;
wire _26421_;
wire _26422_;
wire _26423_;
wire _26424_;
wire _26425_;
wire _26426_;
wire _26427_;
wire _26428_;
wire _26429_;
wire _26430_;
wire _26431_;
wire _26432_;
wire _26433_;
wire _26434_;
wire _26435_;
wire _26436_;
wire _26437_;
wire _26438_;
wire _26439_;
wire _26440_;
wire _26441_;
wire _26442_;
wire _26443_;
wire _26444_;
wire _26445_;
wire _26446_;
wire _26447_;
wire _26448_;
wire _26449_;
wire _26450_;
wire _26451_;
wire _26452_;
wire _26453_;
wire _26454_;
wire _26455_;
wire _26456_;
wire _26457_;
wire _26458_;
wire _26459_;
wire _26460_;
wire _26461_;
wire _26462_;
wire _26463_;
wire _26464_;
wire _26465_;
wire _26466_;
wire _26467_;
wire _26468_;
wire _26469_;
wire _26470_;
wire _26471_;
wire _26472_;
wire _26473_;
wire _26474_;
wire _26475_;
wire _26476_;
wire _26477_;
wire _26478_;
wire _26479_;
wire _26480_;
wire _26481_;
wire _26482_;
wire _26483_;
wire _26484_;
wire _26485_;
wire _26486_;
wire _26487_;
wire _26488_;
wire _26489_;
wire _26490_;
wire _26491_;
wire _26492_;
wire _26493_;
wire _26494_;
wire _26495_;
wire _26496_;
wire _26497_;
wire _26498_;
wire _26499_;
wire _26500_;
wire _26501_;
wire _26502_;
wire _26503_;
wire _26504_;
wire _26505_;
wire _26506_;
wire _26507_;
wire _26508_;
wire _26509_;
wire _26510_;
wire _26511_;
wire _26512_;
wire _26513_;
wire _26514_;
wire _26515_;
wire _26516_;
wire _26517_;
wire _26518_;
wire _26519_;
wire _26520_;
wire _26521_;
wire _26522_;
wire _26523_;
wire _26524_;
wire _26525_;
wire _26526_;
wire _26527_;
wire _26528_;
wire _26529_;
wire _26530_;
wire _26531_;
wire _26532_;
wire _26533_;
wire _26534_;
wire _26535_;
wire _26536_;
wire _26537_;
wire _26538_;
wire _26539_;
wire _26540_;
wire _26541_;
wire _26542_;
wire _26543_;
wire _26544_;
wire _26545_;
wire _26546_;
wire _26547_;
wire _26548_;
wire _26549_;
wire _26550_;
wire _26551_;
wire _26552_;
wire _26553_;
wire _26554_;
wire _26555_;
wire _26556_;
wire _26557_;
wire _26558_;
wire _26559_;
wire _26560_;
wire _26561_;
wire _26562_;
wire _26563_;
wire _26564_;
wire _26565_;
wire _26566_;
wire _26567_;
wire _26568_;
wire _26569_;
wire _26570_;
wire _26571_;
wire _26572_;
wire _26573_;
wire _26574_;
wire _26575_;
wire _26576_;
wire _26577_;
wire _26578_;
wire _26579_;
wire _26580_;
wire _26581_;
wire _26582_;
wire _26583_;
wire _26584_;
wire _26585_;
wire _26586_;
wire _26587_;
wire _26588_;
wire _26589_;
wire _26590_;
wire _26591_;
wire _26592_;
wire _26593_;
wire _26594_;
wire _26595_;
wire _26596_;
wire _26597_;
wire _26598_;
wire _26599_;
wire _26600_;
wire _26601_;
wire _26602_;
wire _26603_;
wire _26604_;
wire _26605_;
wire _26606_;
wire _26607_;
wire _26608_;
wire _26609_;
wire _26610_;
wire _26611_;
wire _26612_;
wire _26613_;
wire _26614_;
wire _26615_;
wire _26616_;
wire _26617_;
wire _26618_;
wire _26619_;
wire _26620_;
wire _26621_;
wire _26622_;
wire _26623_;
wire _26624_;
wire _26625_;
wire _26626_;
wire _26627_;
wire _26628_;
wire _26629_;
wire _26630_;
wire _26631_;
wire _26632_;
wire _26633_;
wire _26634_;
wire _26635_;
wire _26636_;
wire _26637_;
wire _26638_;
wire _26639_;
wire _26640_;
wire _26641_;
wire _26642_;
wire _26643_;
wire _26644_;
wire _26645_;
wire _26646_;
wire _26647_;
wire _26648_;
wire _26649_;
wire _26650_;
wire _26651_;
wire _26652_;
wire _26653_;
wire _26654_;
wire _26655_;
wire _26656_;
wire _26657_;
wire _26658_;
wire _26659_;
wire _26660_;
wire _26661_;
wire _26662_;
wire _26663_;
wire _26664_;
wire _26665_;
wire _26666_;
wire _26667_;
wire _26668_;
wire _26669_;
wire _26670_;
wire _26671_;
wire _26672_;
wire _26673_;
wire _26674_;
wire _26675_;
wire _26676_;
wire _26677_;
wire _26678_;
wire _26679_;
wire _26680_;
wire _26681_;
wire _26682_;
wire _26683_;
wire _26684_;
wire _26685_;
wire _26686_;
wire _26687_;
wire _26688_;
wire _26689_;
wire _26690_;
wire _26691_;
wire _26692_;
wire _26693_;
wire _26694_;
wire _26695_;
wire _26696_;
wire _26697_;
wire _26698_;
wire _26699_;
wire _26700_;
wire _26701_;
wire _26702_;
wire _26703_;
wire _26704_;
wire _26705_;
wire _26706_;
wire _26707_;
wire _26708_;
wire _26709_;
wire _26710_;
wire _26711_;
wire _26712_;
wire _26713_;
wire _26714_;
wire _26715_;
wire _26716_;
wire _26717_;
wire _26718_;
wire _26719_;
wire _26720_;
wire _26721_;
wire _26722_;
wire _26723_;
wire _26724_;
wire _26725_;
wire _26726_;
wire _26727_;
wire _26728_;
wire _26729_;
wire _26730_;
wire _26731_;
wire _26732_;
wire _26733_;
wire _26734_;
wire _26735_;
wire _26736_;
wire _26737_;
wire _26738_;
wire _26739_;
wire _26740_;
wire _26741_;
wire _26742_;
wire _26743_;
wire _26744_;
wire _26745_;
wire _26746_;
wire _26747_;
wire _26748_;
wire _26749_;
wire _26750_;
wire _26751_;
wire _26752_;
wire _26753_;
wire _26754_;
wire _26755_;
wire _26756_;
wire _26757_;
wire _26758_;
wire _26759_;
wire _26760_;
wire _26761_;
wire _26762_;
wire _26763_;
wire _26764_;
wire _26765_;
wire _26766_;
wire _26767_;
wire _26768_;
wire _26769_;
wire _26770_;
wire _26771_;
wire _26772_;
wire _26773_;
wire _26774_;
wire _26775_;
wire _26776_;
wire _26777_;
wire _26778_;
wire _26779_;
wire _26780_;
wire _26781_;
wire _26782_;
wire _26783_;
wire _26784_;
wire _26785_;
wire _26786_;
wire _26787_;
wire _26788_;
wire _26789_;
wire _26790_;
wire _26791_;
wire _26792_;
wire _26793_;
wire _26794_;
wire _26795_;
wire _26796_;
wire _26797_;
wire _26798_;
wire _26799_;
wire _26800_;
wire _26801_;
wire _26802_;
wire _26803_;
wire _26804_;
wire _26805_;
wire _26806_;
wire _26807_;
wire _26808_;
wire _26809_;
wire _26810_;
wire _26811_;
wire _26812_;
wire _26813_;
wire _26814_;
wire _26815_;
wire _26816_;
wire _26817_;
wire _26818_;
wire _26819_;
wire _26820_;
wire _26821_;
wire _26822_;
wire _26823_;
wire _26824_;
wire _26825_;
wire _26826_;
wire _26827_;
wire _26828_;
wire _26829_;
wire _26830_;
wire _26831_;
wire _26832_;
wire _26833_;
wire _26834_;
wire _26835_;
wire _26836_;
wire _26837_;
wire _26838_;
wire _26839_;
wire _26840_;
wire _26841_;
wire _26842_;
wire _26843_;
wire _26844_;
wire _26845_;
wire _26846_;
wire _26847_;
wire _26848_;
wire _26849_;
wire _26850_;
wire _26851_;
wire _26852_;
wire _26853_;
wire _26854_;
wire _26855_;
wire _26856_;
wire _26857_;
wire _26858_;
wire _26859_;
wire _26860_;
wire _26861_;
wire _26862_;
wire _26863_;
wire _26864_;
wire _26865_;
wire _26866_;
wire _26867_;
wire _26868_;
wire _26869_;
wire _26870_;
wire _26871_;
wire _26872_;
wire _26873_;
wire _26874_;
wire _26875_;
wire _26876_;
wire _26877_;
wire _26878_;
wire _26879_;
wire _26880_;
wire _26881_;
wire _26882_;
wire _26883_;
wire _26884_;
wire _26885_;
wire _26886_;
wire _26887_;
wire _26888_;
wire _26889_;
wire _26890_;
wire _26891_;
wire _26892_;
wire _26893_;
wire _26894_;
wire _26895_;
wire _26896_;
wire _26897_;
wire _26898_;
wire _26899_;
wire _26900_;
wire _26901_;
wire _26902_;
wire _26903_;
wire _26904_;
wire _26905_;
wire _26906_;
wire _26907_;
wire _26908_;
wire _26909_;
wire _26910_;
wire _26911_;
wire _26912_;
wire _26913_;
wire _26914_;
wire _26915_;
wire _26916_;
wire _26917_;
wire _26918_;
wire _26919_;
wire _26920_;
wire _26921_;
wire _26922_;
wire _26923_;
wire _26924_;
wire _26925_;
wire _26926_;
wire _26927_;
wire _26928_;
wire _26929_;
wire _26930_;
wire _26931_;
wire _26932_;
wire _26933_;
wire _26934_;
wire _26935_;
wire _26936_;
wire _26937_;
wire _26938_;
wire _26939_;
wire _26940_;
wire _26941_;
wire _26942_;
wire _26943_;
wire _26944_;
wire _26945_;
wire _26946_;
wire _26947_;
wire _26948_;
wire _26949_;
wire _26950_;
wire _26951_;
wire _26952_;
wire _26953_;
wire _26954_;
wire _26955_;
wire _26956_;
wire _26957_;
wire _26958_;
wire _26959_;
wire _26960_;
wire _26961_;
wire _26962_;
wire _26963_;
wire _26964_;
wire _26965_;
wire _26966_;
wire _26967_;
wire _26968_;
wire _26969_;
wire _26970_;
wire _26971_;
wire _26972_;
wire _26973_;
wire _26974_;
wire _26975_;
wire _26976_;
wire _26977_;
wire _26978_;
wire _26979_;
wire _26980_;
wire _26981_;
wire _26982_;
wire _26983_;
wire _26984_;
wire _26985_;
wire _26986_;
wire _26987_;
wire _26988_;
wire _26989_;
wire _26990_;
wire _26991_;
wire _26992_;
wire _26993_;
wire _26994_;
wire _26995_;
wire _26996_;
wire _26997_;
wire _26998_;
wire _26999_;
wire _27000_;
wire _27001_;
wire _27002_;
wire _27003_;
wire _27004_;
wire _27005_;
wire _27006_;
wire _27007_;
wire _27008_;
wire _27009_;
wire _27010_;
wire _27011_;
wire _27012_;
wire _27013_;
wire _27014_;
wire _27015_;
wire _27016_;
wire _27017_;
wire _27018_;
wire _27019_;
wire _27020_;
wire _27021_;
wire _27022_;
wire _27023_;
wire _27024_;
wire _27025_;
wire _27026_;
wire _27027_;
wire _27028_;
wire _27029_;
wire _27030_;
wire _27031_;
wire _27032_;
wire _27033_;
wire _27034_;
wire _27035_;
wire _27036_;
wire _27037_;
wire _27038_;
wire _27039_;
wire _27040_;
wire _27041_;
wire _27042_;
wire _27043_;
wire _27044_;
wire _27045_;
wire _27046_;
wire _27047_;
wire _27048_;
wire _27049_;
wire _27050_;
wire _27051_;
wire _27052_;
wire _27053_;
wire _27054_;
wire _27055_;
wire _27056_;
wire _27057_;
wire _27058_;
wire _27059_;
wire _27060_;
wire _27061_;
wire _27062_;
wire _27063_;
wire _27064_;
wire _27065_;
wire _27066_;
wire _27067_;
wire _27068_;
wire _27069_;
wire _27070_;
wire _27071_;
wire _27072_;
wire _27073_;
wire _27074_;
wire _27075_;
wire _27076_;
wire _27077_;
wire _27078_;
wire _27079_;
wire _27080_;
wire _27081_;
wire _27082_;
wire _27083_;
wire _27084_;
wire _27085_;
wire _27086_;
wire _27087_;
wire _27088_;
wire _27089_;
wire _27090_;
wire _27091_;
wire _27092_;
wire _27093_;
wire _27094_;
wire _27095_;
wire _27096_;
wire _27097_;
wire _27098_;
wire _27099_;
wire _27100_;
wire _27101_;
wire _27102_;
wire _27103_;
wire _27104_;
wire _27105_;
wire _27106_;
wire _27107_;
wire _27108_;
wire _27109_;
wire _27110_;
wire _27111_;
wire _27112_;
wire _27113_;
wire _27114_;
wire _27115_;
wire _27116_;
wire _27117_;
wire _27118_;
wire _27119_;
wire _27120_;
wire _27121_;
wire _27122_;
wire _27123_;
wire _27124_;
wire _27125_;
wire _27126_;
wire _27127_;
wire _27128_;
wire _27129_;
wire _27130_;
wire _27131_;
wire _27132_;
wire _27133_;
wire _27134_;
wire _27135_;
wire _27136_;
wire _27137_;
wire _27138_;
wire _27139_;
wire _27140_;
wire _27141_;
wire _27142_;
wire _27143_;
wire _27144_;
wire _27145_;
wire _27146_;
wire _27147_;
wire _27148_;
wire _27149_;
wire _27150_;
wire _27151_;
wire _27152_;
wire _27153_;
wire _27154_;
wire _27155_;
wire _27156_;
wire _27157_;
wire _27158_;
wire _27159_;
wire _27160_;
wire _27161_;
wire _27162_;
wire _27163_;
wire _27164_;
wire _27165_;
wire _27166_;
wire _27167_;
wire _27168_;
wire _27169_;
wire _27170_;
wire _27171_;
wire _27172_;
wire _27173_;
wire _27174_;
wire _27175_;
wire _27176_;
wire _27177_;
wire _27178_;
wire _27179_;
wire _27180_;
wire _27181_;
wire _27182_;
wire _27183_;
wire _27184_;
wire _27185_;
wire _27186_;
wire _27187_;
wire _27188_;
wire _27189_;
wire _27190_;
wire _27191_;
wire _27192_;
wire _27193_;
wire _27194_;
wire _27195_;
wire _27196_;
wire _27197_;
wire _27198_;
wire _27199_;
wire _27200_;
wire _27201_;
wire _27202_;
wire _27203_;
wire _27204_;
wire _27205_;
wire _27206_;
wire _27207_;
wire _27208_;
wire _27209_;
wire _27210_;
wire _27211_;
wire _27212_;
wire _27213_;
wire _27214_;
wire _27215_;
wire _27216_;
wire _27217_;
wire _27218_;
wire _27219_;
wire _27220_;
wire _27221_;
wire _27222_;
wire _27223_;
wire _27224_;
wire _27225_;
wire _27226_;
wire _27227_;
wire _27228_;
wire _27229_;
wire _27230_;
wire _27231_;
wire _27232_;
wire _27233_;
wire _27234_;
wire _27235_;
wire _27236_;
wire _27237_;
wire _27238_;
wire _27239_;
wire _27240_;
wire _27241_;
wire _27242_;
wire _27243_;
wire _27244_;
wire _27245_;
wire _27246_;
wire _27247_;
wire _27248_;
wire _27249_;
wire _27250_;
wire _27251_;
wire _27252_;
wire _27253_;
wire _27254_;
wire _27255_;
wire _27256_;
wire _27257_;
wire _27258_;
wire _27259_;
wire _27260_;
wire _27261_;
wire _27262_;
wire _27263_;
wire _27264_;
wire _27265_;
wire _27266_;
wire _27267_;
wire _27268_;
wire _27269_;
wire _27270_;
wire _27271_;
wire _27272_;
wire _27273_;
wire _27274_;
wire _27275_;
wire _27276_;
wire _27277_;
wire _27278_;
wire _27279_;
wire _27280_;
wire _27281_;
wire _27282_;
wire _27283_;
wire _27284_;
wire _27285_;
wire _27286_;
wire _27287_;
wire _27288_;
wire _27289_;
wire _27290_;
wire _27291_;
wire _27292_;
wire _27293_;
wire _27294_;
wire _27295_;
wire _27296_;
wire _27297_;
wire _27298_;
wire _27299_;
wire _27300_;
wire _27301_;
wire _27302_;
wire _27303_;
wire _27304_;
wire _27305_;
wire _27306_;
wire _27307_;
wire _27308_;
wire _27309_;
wire _27310_;
wire _27311_;
wire _27312_;
wire _27313_;
wire _27314_;
wire _27315_;
wire _27316_;
wire _27317_;
wire _27318_;
wire _27319_;
wire _27320_;
wire _27321_;
wire _27322_;
wire _27323_;
wire _27324_;
wire _27325_;
wire _27326_;
wire _27327_;
wire _27328_;
wire _27329_;
wire _27330_;
wire _27331_;
wire _27332_;
wire _27333_;
wire _27334_;
wire _27335_;
wire _27336_;
wire _27337_;
wire _27338_;
wire _27339_;
wire _27340_;
wire _27341_;
wire _27342_;
wire _27343_;
wire _27344_;
wire _27345_;
wire _27346_;
wire _27347_;
wire _27348_;
wire _27349_;
wire _27350_;
wire _27351_;
wire _27352_;
wire _27353_;
wire _27354_;
wire _27355_;
wire _27356_;
wire _27357_;
wire _27358_;
wire _27359_;
wire _27360_;
wire _27361_;
wire _27362_;
wire _27363_;
wire _27364_;
wire _27365_;
wire _27366_;
wire _27367_;
wire _27368_;
wire _27369_;
wire _27370_;
wire _27371_;
wire _27372_;
wire _27373_;
wire _27374_;
wire _27375_;
wire _27376_;
wire _27377_;
wire _27378_;
wire _27379_;
wire _27380_;
wire _27381_;
wire _27382_;
wire _27383_;
wire _27384_;
wire _27385_;
wire _27386_;
wire _27387_;
wire _27388_;
wire _27389_;
wire _27390_;
wire _27391_;
wire _27392_;
wire _27393_;
wire _27394_;
wire _27395_;
wire _27396_;
wire _27397_;
wire _27398_;
wire _27399_;
wire _27400_;
wire _27401_;
wire _27402_;
wire _27403_;
wire _27404_;
wire _27405_;
wire _27406_;
wire _27407_;
wire _27408_;
wire _27409_;
wire _27410_;
wire _27411_;
wire _27412_;
wire _27413_;
wire _27414_;
wire _27415_;
wire _27416_;
wire _27417_;
wire _27418_;
wire _27419_;
wire _27420_;
wire _27421_;
wire _27422_;
wire _27423_;
wire _27424_;
wire _27425_;
wire _27426_;
wire _27427_;
wire _27428_;
wire _27429_;
wire _27430_;
wire _27431_;
wire _27432_;
wire _27433_;
wire _27434_;
wire _27435_;
wire _27436_;
wire _27437_;
wire _27438_;
wire _27439_;
wire _27440_;
wire _27441_;
wire _27442_;
wire _27443_;
wire _27444_;
wire _27445_;
wire _27446_;
wire _27447_;
wire _27448_;
wire _27449_;
wire _27450_;
wire _27451_;
wire _27452_;
wire _27453_;
wire _27454_;
wire _27455_;
wire _27456_;
wire _27457_;
wire _27458_;
wire _27459_;
wire _27460_;
wire _27461_;
wire _27462_;
wire _27463_;
wire _27464_;
wire _27465_;
wire _27466_;
wire _27467_;
wire _27468_;
wire _27469_;
wire _27470_;
wire _27471_;
wire _27472_;
wire _27473_;
wire _27474_;
wire _27475_;
wire _27476_;
wire _27477_;
wire _27478_;
wire _27479_;
wire _27480_;
wire _27481_;
wire _27482_;
wire _27483_;
wire _27484_;
wire _27485_;
wire _27486_;
wire _27487_;
wire _27488_;
wire _27489_;
wire _27490_;
wire _27491_;
wire _27492_;
wire _27493_;
wire _27494_;
wire _27495_;
wire _27496_;
wire _27497_;
wire _27498_;
wire _27499_;
wire _27500_;
wire _27501_;
wire _27502_;
wire _27503_;
wire _27504_;
wire _27505_;
wire _27506_;
wire _27507_;
wire _27508_;
wire _27509_;
wire _27510_;
wire _27511_;
wire _27512_;
wire _27513_;
wire _27514_;
wire _27515_;
wire _27516_;
wire _27517_;
wire _27518_;
wire _27519_;
wire _27520_;
wire _27521_;
wire _27522_;
wire _27523_;
wire _27524_;
wire _27525_;
wire _27526_;
wire _27527_;
wire _27528_;
wire _27529_;
wire _27530_;
wire _27531_;
wire _27532_;
wire _27533_;
wire _27534_;
wire _27535_;
wire _27536_;
wire _27537_;
wire _27538_;
wire _27539_;
wire _27540_;
wire _27541_;
wire _27542_;
wire _27543_;
wire _27544_;
wire _27545_;
wire _27546_;
wire _27547_;
wire _27548_;
wire _27549_;
wire _27550_;
wire _27551_;
wire _27552_;
wire _27553_;
wire _27554_;
wire _27555_;
wire _27556_;
wire _27557_;
wire _27558_;
wire _27559_;
wire _27560_;
wire _27561_;
wire _27562_;
wire _27563_;
wire _27564_;
wire _27565_;
wire _27566_;
wire _27567_;
wire _27568_;
wire _27569_;
wire _27570_;
wire _27571_;
wire _27572_;
wire _27573_;
wire _27574_;
wire _27575_;
wire _27576_;
wire _27577_;
wire _27578_;
wire _27579_;
wire _27580_;
wire _27581_;
wire _27582_;
wire _27583_;
wire _27584_;
wire _27585_;
wire _27586_;
wire _27587_;
wire _27588_;
wire _27589_;
wire _27590_;
wire _27591_;
wire _27592_;
wire _27593_;
wire _27594_;
wire _27595_;
wire _27596_;
wire _27597_;
wire _27598_;
wire _27599_;
wire _27600_;
wire _27601_;
wire _27602_;
wire _27603_;
wire _27604_;
wire _27605_;
wire _27606_;
wire _27607_;
wire _27608_;
wire _27609_;
wire _27610_;
wire _27611_;
wire _27612_;
wire _27613_;
wire _27614_;
wire _27615_;
wire _27616_;
wire _27617_;
wire _27618_;
wire _27619_;
wire _27620_;
wire _27621_;
wire _27622_;
wire _27623_;
wire _27624_;
wire _27625_;
wire _27626_;
wire _27627_;
wire _27628_;
wire _27629_;
wire _27630_;
wire _27631_;
wire _27632_;
wire _27633_;
wire _27634_;
wire _27635_;
wire _27636_;
wire _27637_;
wire _27638_;
wire _27639_;
wire _27640_;
wire _27641_;
wire _27642_;
wire _27643_;
wire _27644_;
wire _27645_;
wire _27646_;
wire _27647_;
wire _27648_;
wire _27649_;
wire _27650_;
wire _27651_;
wire _27652_;
wire _27653_;
wire _27654_;
wire _27655_;
wire _27656_;
wire _27657_;
wire _27658_;
wire _27659_;
wire _27660_;
wire _27661_;
wire _27662_;
wire _27663_;
wire _27664_;
wire _27665_;
wire _27666_;
wire _27667_;
wire _27668_;
wire _27669_;
wire _27670_;
wire _27671_;
wire _27672_;
wire _27673_;
wire _27674_;
wire _27675_;
wire _27676_;
wire _27677_;
wire _27678_;
wire _27679_;
wire _27680_;
wire _27681_;
wire _27682_;
wire _27683_;
wire _27684_;
wire _27685_;
wire _27686_;
wire _27687_;
wire _27688_;
wire _27689_;
wire _27690_;
wire _27691_;
wire _27692_;
wire _27693_;
wire _27694_;
wire _27695_;
wire _27696_;
wire _27697_;
wire _27698_;
wire _27699_;
wire _27700_;
wire _27701_;
wire _27702_;
wire _27703_;
wire _27704_;
wire _27705_;
wire _27706_;
wire _27707_;
wire _27708_;
wire _27709_;
wire _27710_;
wire _27711_;
wire _27712_;
wire _27713_;
wire _27714_;
wire _27715_;
wire _27716_;
wire _27717_;
wire _27718_;
wire _27719_;
wire _27720_;
wire _27721_;
wire _27722_;
wire _27723_;
wire _27724_;
wire _27725_;
wire _27726_;
wire _27727_;
wire _27728_;
wire _27729_;
wire _27730_;
wire _27731_;
wire _27732_;
wire _27733_;
wire _27734_;
wire _27735_;
wire _27736_;
wire _27737_;
wire _27738_;
wire _27739_;
wire _27740_;
wire _27741_;
wire _27742_;
wire _27743_;
wire _27744_;
wire _27745_;
wire _27746_;
wire _27747_;
wire _27748_;
wire _27749_;
wire _27750_;
wire _27751_;
wire _27752_;
wire _27753_;
wire _27754_;
wire _27755_;
wire _27756_;
wire _27757_;
wire _27758_;
wire _27759_;
wire _27760_;
wire _27761_;
wire _27762_;
wire _27763_;
wire _27764_;
wire _27765_;
wire _27766_;
wire _27767_;
wire _27768_;
wire _27769_;
wire _27770_;
wire _27771_;
wire _27772_;
wire _27773_;
wire _27774_;
wire _27775_;
wire _27776_;
wire _27777_;
wire _27778_;
wire _27779_;
wire _27780_;
wire _27781_;
wire _27782_;
wire _27783_;
wire _27784_;
wire _27785_;
wire _27786_;
wire _27787_;
wire _27788_;
wire _27789_;
wire _27790_;
wire _27791_;
wire _27792_;
wire _27793_;
wire _27794_;
wire _27795_;
wire _27796_;
wire _27797_;
wire _27798_;
wire _27799_;
wire _27800_;
wire _27801_;
wire _27802_;
wire _27803_;
wire _27804_;
wire _27805_;
wire _27806_;
wire _27807_;
wire _27808_;
wire _27809_;
wire _27810_;
wire _27811_;
wire _27812_;
wire _27813_;
wire _27814_;
wire _27815_;
wire _27816_;
wire _27817_;
wire _27818_;
wire _27819_;
wire _27820_;
wire _27821_;
wire _27822_;
wire _27823_;
wire _27824_;
wire _27825_;
wire _27826_;
wire _27827_;
wire _27828_;
wire _27829_;
wire _27830_;
wire _27831_;
wire _27832_;
wire _27833_;
wire _27834_;
wire _27835_;
wire _27836_;
wire _27837_;
wire _27838_;
wire _27839_;
wire _27840_;
wire _27841_;
wire _27842_;
wire _27843_;
wire _27844_;
wire _27845_;
wire _27846_;
wire _27847_;
wire _27848_;
wire _27849_;
wire _27850_;
wire _27851_;
wire _27852_;
wire _27853_;
wire _27854_;
wire _27855_;
wire _27856_;
wire _27857_;
wire _27858_;
wire _27859_;
wire _27860_;
wire _27861_;
wire _27862_;
wire _27863_;
wire _27864_;
wire _27865_;
wire _27866_;
wire _27867_;
wire _27868_;
wire _27869_;
wire _27870_;
wire _27871_;
wire _27872_;
wire _27873_;
wire _27874_;
wire _27875_;
wire _27876_;
wire _27877_;
wire _27878_;
wire _27879_;
wire _27880_;
wire _27881_;
wire _27882_;
wire _27883_;
wire _27884_;
wire _27885_;
wire _27886_;
wire _27887_;
wire _27888_;
wire _27889_;
wire _27890_;
wire _27891_;
wire _27892_;
wire _27893_;
wire _27894_;
wire _27895_;
wire _27896_;
wire _27897_;
wire _27898_;
wire _27899_;
wire _27900_;
wire _27901_;
wire _27902_;
wire _27903_;
wire _27904_;
wire _27905_;
wire _27906_;
wire _27907_;
wire _27908_;
wire _27909_;
wire _27910_;
wire _27911_;
wire _27912_;
wire _27913_;
wire _27914_;
wire _27915_;
wire _27916_;
wire _27917_;
wire _27918_;
wire _27919_;
wire _27920_;
wire _27921_;
wire _27922_;
wire _27923_;
wire _27924_;
wire _27925_;
wire _27926_;
wire _27927_;
wire _27928_;
wire _27929_;
wire _27930_;
wire _27931_;
wire _27932_;
wire _27933_;
wire _27934_;
wire _27935_;
wire _27936_;
wire _27937_;
wire _27938_;
wire _27939_;
wire _27940_;
wire _27941_;
wire _27942_;
wire _27943_;
wire _27944_;
wire _27945_;
wire _27946_;
wire _27947_;
wire _27948_;
wire _27949_;
wire _27950_;
wire _27951_;
wire _27952_;
wire _27953_;
wire _27954_;
wire _27955_;
wire _27956_;
wire _27957_;
wire _27958_;
wire _27959_;
wire _27960_;
wire _27961_;
wire _27962_;
wire _27963_;
wire _27964_;
wire _27965_;
wire _27966_;
wire _27967_;
wire _27968_;
wire _27969_;
wire _27970_;
wire _27971_;
wire _27972_;
wire _27973_;
wire _27974_;
wire _27975_;
wire _27976_;
wire _27977_;
wire _27978_;
wire _27979_;
wire _27980_;
wire _27981_;
wire _27982_;
wire _27983_;
wire _27984_;
wire _27985_;
wire _27986_;
wire _27987_;
wire _27988_;
wire _27989_;
wire _27990_;
wire _27991_;
wire _27992_;
wire _27993_;
wire _27994_;
wire _27995_;
wire _27996_;
wire _27997_;
wire _27998_;
wire _27999_;
wire _28000_;
wire _28001_;
wire _28002_;
wire _28003_;
wire _28004_;
wire _28005_;
wire _28006_;
wire _28007_;
wire _28008_;
wire _28009_;
wire _28010_;
wire _28011_;
wire _28012_;
wire _28013_;
wire _28014_;
wire _28015_;
wire _28016_;
wire _28017_;
wire _28018_;
wire _28019_;
wire _28020_;
wire _28021_;
wire _28022_;
wire _28023_;
wire _28024_;
wire _28025_;
wire _28026_;
wire _28027_;
wire _28028_;
wire _28029_;
wire _28030_;
wire _28031_;
wire _28032_;
wire _28033_;
wire _28034_;
wire _28035_;
wire _28036_;
wire _28037_;
wire _28038_;
wire _28039_;
wire _28040_;
wire _28041_;
wire _28042_;
wire _28043_;
wire _28044_;
wire _28045_;
wire _28046_;
wire _28047_;
wire _28048_;
wire _28049_;
wire _28050_;
wire _28051_;
wire _28052_;
wire _28053_;
wire _28054_;
wire _28055_;
wire _28056_;
wire _28057_;
wire _28058_;
wire _28059_;
wire _28060_;
wire _28061_;
wire _28062_;
wire _28063_;
wire _28064_;
wire _28065_;
wire _28066_;
wire _28067_;
wire _28068_;
wire _28069_;
wire _28070_;
wire _28071_;
wire _28072_;
wire _28073_;
wire _28074_;
wire _28075_;
wire _28076_;
wire _28077_;
wire _28078_;
wire _28079_;
wire _28080_;
wire _28081_;
wire _28082_;
wire _28083_;
wire _28084_;
wire _28085_;
wire _28086_;
wire _28087_;
wire _28088_;
wire _28089_;
wire _28090_;
wire _28091_;
wire _28092_;
wire _28093_;
wire _28094_;
wire _28095_;
wire _28096_;
wire _28097_;
wire _28098_;
wire _28099_;
wire _28100_;
wire _28101_;
wire _28102_;
wire _28103_;
wire _28104_;
wire _28105_;
wire _28106_;
wire _28107_;
wire _28108_;
wire _28109_;
wire _28110_;
wire _28111_;
wire _28112_;
wire _28113_;
wire _28114_;
wire _28115_;
wire _28116_;
wire _28117_;
wire _28118_;
wire _28119_;
wire _28120_;
wire _28121_;
wire _28122_;
wire _28123_;
wire _28124_;
wire _28125_;
wire _28126_;
wire _28127_;
wire _28128_;
wire _28129_;
wire _28130_;
wire _28131_;
wire _28132_;
wire _28133_;
wire _28134_;
wire _28135_;
wire _28136_;
wire _28137_;
wire _28138_;
wire _28139_;
wire _28140_;
wire _28141_;
wire _28142_;
wire _28143_;
wire _28144_;
wire _28145_;
wire _28146_;
wire _28147_;
wire _28148_;
wire _28149_;
wire _28150_;
wire _28151_;
wire _28152_;
wire _28153_;
wire _28154_;
wire _28155_;
wire _28156_;
wire _28157_;
wire _28158_;
wire _28159_;
wire _28160_;
wire _28161_;
wire _28162_;
wire _28163_;
wire _28164_;
wire _28165_;
wire _28166_;
wire _28167_;
wire _28168_;
wire _28169_;
wire _28170_;
wire _28171_;
wire _28172_;
wire _28173_;
wire _28174_;
wire _28175_;
wire _28176_;
wire _28177_;
wire _28178_;
wire _28179_;
wire _28180_;
wire _28181_;
wire _28182_;
wire _28183_;
wire _28184_;
wire _28185_;
wire _28186_;
wire _28187_;
wire _28188_;
wire _28189_;
wire _28190_;
wire _28191_;
wire _28192_;
wire _28193_;
wire _28194_;
wire _28195_;
wire _28196_;
wire _28197_;
wire _28198_;
wire _28199_;
wire _28200_;
wire _28201_;
wire _28202_;
wire _28203_;
wire _28204_;
wire _28205_;
wire _28206_;
wire _28207_;
wire _28208_;
wire _28209_;
wire _28210_;
wire _28211_;
wire _28212_;
wire _28213_;
wire _28214_;
wire _28215_;
wire _28216_;
wire _28217_;
wire _28218_;
wire _28219_;
wire _28220_;
wire _28221_;
wire _28222_;
wire _28223_;
wire _28224_;
wire _28225_;
wire _28226_;
wire _28227_;
wire _28228_;
wire _28229_;
wire _28230_;
wire _28231_;
wire _28232_;
wire _28233_;
wire _28234_;
wire _28235_;
wire _28236_;
wire _28237_;
wire _28238_;
wire _28239_;
wire _28240_;
wire _28241_;
wire _28242_;
wire _28243_;
wire _28244_;
wire _28245_;
wire _28246_;
wire _28247_;
wire _28248_;
wire _28249_;
wire _28250_;
wire _28251_;
wire _28252_;
wire _28253_;
wire _28254_;
wire _28255_;
wire _28256_;
wire _28257_;
wire _28258_;
wire _28259_;
wire _28260_;
wire _28261_;
wire _28262_;
wire _28263_;
wire _28264_;
wire _28265_;
wire _28266_;
wire _28267_;
wire _28268_;
wire _28269_;
wire _28270_;
wire _28271_;
wire _28272_;
wire _28273_;
wire _28274_;
wire _28275_;
wire _28276_;
wire _28277_;
wire _28278_;
wire _28279_;
wire _28280_;
wire _28281_;
wire _28282_;
wire _28283_;
wire _28284_;
wire _28285_;
wire _28286_;
wire _28287_;
wire _28288_;
wire _28289_;
wire _28290_;
wire _28291_;
wire _28292_;
wire _28293_;
wire _28294_;
wire _28295_;
wire _28296_;
wire _28297_;
wire _28298_;
wire _28299_;
wire _28300_;
wire _28301_;
wire _28302_;
wire _28303_;
wire _28304_;
wire _28305_;
wire _28306_;
wire _28307_;
wire _28308_;
wire _28309_;
wire _28310_;
wire _28311_;
wire _28312_;
wire _28313_;
wire _28314_;
wire _28315_;
wire _28316_;
wire _28317_;
wire _28318_;
wire _28319_;
wire _28320_;
wire _28321_;
wire _28322_;
wire _28323_;
wire _28324_;
wire _28325_;
wire _28326_;
wire _28327_;
wire _28328_;
wire _28329_;
wire _28330_;
wire _28331_;
wire _28332_;
wire _28333_;
wire _28334_;
wire _28335_;
wire _28336_;
wire _28337_;
wire _28338_;
wire _28339_;
wire _28340_;
wire _28341_;
wire _28342_;
wire _28343_;
wire _28344_;
wire _28345_;
wire _28346_;
wire _28347_;
wire _28348_;
wire _28349_;
wire _28350_;
wire _28351_;
wire _28352_;
wire _28353_;
wire _28354_;
wire _28355_;
wire _28356_;
wire _28357_;
wire _28358_;
wire _28359_;
wire _28360_;
wire _28361_;
wire _28362_;
wire _28363_;
wire _28364_;
wire _28365_;
wire _28366_;
wire _28367_;
wire _28368_;
wire _28369_;
wire _28370_;
wire _28371_;
wire _28372_;
wire _28373_;
wire _28374_;
wire _28375_;
wire _28376_;
wire _28377_;
wire _28378_;
wire _28379_;
wire _28380_;
wire _28381_;
wire _28382_;
wire _28383_;
wire _28384_;
wire _28385_;
wire _28386_;
wire _28387_;
wire _28388_;
wire _28389_;
wire _28390_;
wire _28391_;
wire _28392_;
wire _28393_;
wire _28394_;
wire _28395_;
wire _28396_;
wire _28397_;
wire _28398_;
wire _28399_;
wire _28400_;
wire _28401_;
wire _28402_;
wire _28403_;
wire _28404_;
wire _28405_;
wire _28406_;
wire _28407_;
wire _28408_;
wire _28409_;
wire _28410_;
wire _28411_;
wire _28412_;
wire _28413_;
wire _28414_;
wire _28415_;
wire _28416_;
wire _28417_;
wire _28418_;
wire _28419_;
wire _28420_;
wire _28421_;
wire _28422_;
wire _28423_;
wire _28424_;
wire _28425_;
wire _28426_;
wire _28427_;
wire _28428_;
wire _28429_;
wire _28430_;
wire _28431_;
wire _28432_;
wire _28433_;
wire _28434_;
wire _28435_;
wire _28436_;
wire _28437_;
wire _28438_;
wire _28439_;
wire _28440_;
wire _28441_;
wire _28442_;
wire _28443_;
wire _28444_;
wire _28445_;
wire _28446_;
wire _28447_;
wire _28448_;
wire _28449_;
wire _28450_;
wire _28451_;
wire _28452_;
wire _28453_;
wire _28454_;
wire _28455_;
wire _28456_;
wire _28457_;
wire _28458_;
wire _28459_;
wire _28460_;
wire _28461_;
wire _28462_;
wire _28463_;
wire _28464_;
wire _28465_;
wire _28466_;
wire _28467_;
wire _28468_;
wire _28469_;
wire _28470_;
wire _28471_;
wire _28472_;
wire _28473_;
wire _28474_;
wire _28475_;
wire _28476_;
wire _28477_;
wire _28478_;
wire _28479_;
wire _28480_;
wire _28481_;
wire _28482_;
wire _28483_;
wire _28484_;
wire _28485_;
wire _28486_;
wire _28487_;
wire _28488_;
wire _28489_;
wire _28490_;
wire _28491_;
wire _28492_;
wire _28493_;
wire _28494_;
wire _28495_;
wire _28496_;
wire _28497_;
wire _28498_;
wire _28499_;
wire _28500_;
wire _28501_;
wire _28502_;
wire _28503_;
wire _28504_;
wire _28505_;
wire _28506_;
wire _28507_;
wire _28508_;
wire _28509_;
wire _28510_;
wire _28511_;
wire _28512_;
wire _28513_;
wire _28514_;
wire _28515_;
wire _28516_;
wire _28517_;
wire _28518_;
wire _28519_;
wire _28520_;
wire _28521_;
wire _28522_;
wire _28523_;
wire _28524_;
wire _28525_;
wire _28526_;
wire _28527_;
wire _28528_;
wire _28529_;
wire _28530_;
wire _28531_;
wire _28532_;
wire _28533_;
wire _28534_;
wire _28535_;
wire _28536_;
wire _28537_;
wire _28538_;
wire _28539_;
wire _28540_;
wire _28541_;
wire _28542_;
wire _28543_;
wire _28544_;
wire _28545_;
wire _28546_;
wire _28547_;
wire _28548_;
wire _28549_;
wire _28550_;
wire _28551_;
wire _28552_;
wire _28553_;
wire _28554_;
wire _28555_;
wire _28556_;
wire _28557_;
wire _28558_;
wire _28559_;
wire _28560_;
wire _28561_;
wire _28562_;
wire _28563_;
wire _28564_;
wire _28565_;
wire _28566_;
wire _28567_;
wire _28568_;
wire _28569_;
wire _28570_;
wire _28571_;
wire _28572_;
wire _28573_;
wire _28574_;
wire _28575_;
wire _28576_;
wire _28577_;
wire _28578_;
wire _28579_;
wire _28580_;
wire _28581_;
wire _28582_;
wire _28583_;
wire _28584_;
wire _28585_;
wire _28586_;
wire _28587_;
wire _28588_;
wire _28589_;
wire _28590_;
wire _28591_;
wire _28592_;
wire _28593_;
wire _28594_;
wire _28595_;
wire _28596_;
wire _28597_;
wire _28598_;
wire _28599_;
wire _28600_;
wire _28601_;
wire _28602_;
wire _28603_;
wire _28604_;
wire _28605_;
wire _28606_;
wire _28607_;
wire _28608_;
wire _28609_;
wire _28610_;
wire _28611_;
wire _28612_;
wire _28613_;
wire _28614_;
wire _28615_;
wire _28616_;
wire _28617_;
wire _28618_;
wire _28619_;
wire _28620_;
wire _28621_;
wire _28622_;
wire _28623_;
wire _28624_;
wire _28625_;
wire _28626_;
wire _28627_;
wire _28628_;
wire _28629_;
wire _28630_;
wire _28631_;
wire _28632_;
wire _28633_;
wire _28634_;
wire _28635_;
wire _28636_;
wire _28637_;
wire _28638_;
wire _28639_;
wire _28640_;
wire _28641_;
wire _28642_;
wire _28643_;
wire _28644_;
wire _28645_;
wire _28646_;
wire _28647_;
wire _28648_;
wire _28649_;
wire _28650_;
wire _28651_;
wire _28652_;
wire _28653_;
wire _28654_;
wire _28655_;
wire _28656_;
wire _28657_;
wire _28658_;
wire _28659_;
wire _28660_;
wire _28661_;
wire _28662_;
wire _28663_;
wire _28664_;
wire _28665_;
wire _28666_;
wire _28667_;
wire _28668_;
wire _28669_;
wire _28670_;
wire _28671_;
wire _28672_;
wire _28673_;
wire _28674_;
wire _28675_;
wire _28676_;
wire _28677_;
wire _28678_;
wire _28679_;
wire _28680_;
wire _28681_;
wire _28682_;
wire _28683_;
wire _28684_;
wire _28685_;
wire _28686_;
wire _28687_;
wire _28688_;
wire _28689_;
wire _28690_;
wire _28691_;
wire _28692_;
wire _28693_;
wire _28694_;
wire _28695_;
wire _28696_;
wire _28697_;
wire _28698_;
wire _28699_;
wire _28700_;
wire _28701_;
wire _28702_;
wire _28703_;
wire _28704_;
wire _28705_;
wire _28706_;
wire _28707_;
wire _28708_;
wire _28709_;
wire _28710_;
wire _28711_;
wire _28712_;
wire _28713_;
wire _28714_;
wire _28715_;
wire _28716_;
wire _28717_;
wire _28718_;
wire _28719_;
wire _28720_;
wire _28721_;
wire _28722_;
wire _28723_;
wire _28724_;
wire _28725_;
wire _28726_;
wire _28727_;
wire _28728_;
wire _28729_;
wire _28730_;
wire _28731_;
wire _28732_;
wire _28733_;
wire _28734_;
wire _28735_;
wire _28736_;
wire _28737_;
wire _28738_;
wire _28739_;
wire _28740_;
wire _28741_;
wire _28742_;
wire _28743_;
wire _28744_;
wire _28745_;
wire _28746_;
wire _28747_;
wire _28748_;
wire _28749_;
wire _28750_;
wire _28751_;
wire _28752_;
wire _28753_;
wire _28754_;
wire _28755_;
wire _28756_;
wire _28757_;
wire _28758_;
wire _28759_;
wire _28760_;
wire _28761_;
wire _28762_;
wire _28763_;
wire _28764_;
wire _28765_;
wire _28766_;
wire _28767_;
wire _28768_;
wire _28769_;
wire _28770_;
wire _28771_;
wire _28772_;
wire _28773_;
wire _28774_;
wire _28775_;
wire _28776_;
wire _28777_;
wire _28778_;
wire _28779_;
wire _28780_;
wire _28781_;
wire _28782_;
wire _28783_;
wire _28784_;
wire _28785_;
wire _28786_;
wire _28787_;
wire _28788_;
wire _28789_;
wire _28790_;
wire _28791_;
wire _28792_;
wire _28793_;
wire _28794_;
wire _28795_;
wire _28796_;
wire _28797_;
wire _28798_;
wire _28799_;
wire _28800_;
wire _28801_;
wire _28802_;
wire _28803_;
wire _28804_;
wire _28805_;
wire _28806_;
wire _28807_;
wire _28808_;
wire _28809_;
wire _28810_;
wire _28811_;
wire _28812_;
wire _28813_;
wire _28814_;
wire _28815_;
wire _28816_;
wire _28817_;
wire _28818_;
wire _28819_;
wire _28820_;
wire _28821_;
wire _28822_;
wire _28823_;
wire _28824_;
wire _28825_;
wire _28826_;
wire _28827_;
wire _28828_;
wire _28829_;
wire _28830_;
wire _28831_;
wire _28832_;
wire _28833_;
wire _28834_;
wire _28835_;
wire _28836_;
wire _28837_;
wire _28838_;
wire _28839_;
wire _28840_;
wire _28841_;
wire _28842_;
wire _28843_;
wire _28844_;
wire _28845_;
wire _28846_;
wire _28847_;
wire _28848_;
wire _28849_;
wire _28850_;
wire _28851_;
wire _28852_;
wire _28853_;
wire _28854_;
wire _28855_;
wire _28856_;
wire _28857_;
wire _28858_;
wire _28859_;
wire _28860_;
wire _28861_;
wire _28862_;
wire _28863_;
wire _28864_;
wire _28865_;
wire _28866_;
wire _28867_;
wire _28868_;
wire _28869_;
wire _28870_;
wire _28871_;
wire _28872_;
wire _28873_;
wire _28874_;
wire _28875_;
wire _28876_;
wire _28877_;
wire _28878_;
wire _28879_;
wire _28880_;
wire _28881_;
wire _28882_;
wire _28883_;
wire _28884_;
wire _28885_;
wire _28886_;
wire _28887_;
wire _28888_;
wire _28889_;
wire _28890_;
wire _28891_;
wire _28892_;
wire _28893_;
wire _28894_;
wire _28895_;
wire _28896_;
wire _28897_;
wire _28898_;
wire _28899_;
wire _28900_;
wire _28901_;
wire _28902_;
wire _28903_;
wire _28904_;
wire _28905_;
wire _28906_;
wire _28907_;
wire _28908_;
wire _28909_;
wire _28910_;
wire _28911_;
wire _28912_;
wire _28913_;
wire _28914_;
wire _28915_;
wire _28916_;
wire _28917_;
wire _28918_;
wire _28919_;
wire _28920_;
wire _28921_;
wire _28922_;
wire _28923_;
wire _28924_;
wire _28925_;
wire _28926_;
wire _28927_;
wire _28928_;
wire _28929_;
wire _28930_;
wire _28931_;
wire _28932_;
wire _28933_;
wire _28934_;
wire _28935_;
wire _28936_;
wire _28937_;
wire _28938_;
wire _28939_;
wire _28940_;
wire _28941_;
wire _28942_;
wire _28943_;
wire _28944_;
wire _28945_;
wire _28946_;
wire _28947_;
wire _28948_;
wire _28949_;
wire _28950_;
wire _28951_;
wire _28952_;
wire _28953_;
wire _28954_;
wire _28955_;
wire _28956_;
wire _28957_;
wire _28958_;
wire _28959_;
wire _28960_;
wire _28961_;
wire _28962_;
wire _28963_;
wire _28964_;
wire _28965_;
wire _28966_;
wire _28967_;
wire _28968_;
wire _28969_;
wire _28970_;
wire _28971_;
wire _28972_;
wire _28973_;
wire _28974_;
wire _28975_;
wire _28976_;
wire _28977_;
wire _28978_;
wire _28979_;
wire _28980_;
wire _28981_;
wire _28982_;
wire _28983_;
wire _28984_;
wire _28985_;
wire _28986_;
wire _28987_;
wire _28988_;
wire _28989_;
wire _28990_;
wire zeroWire;
wire oneWire;
assign zeroWire = 1'b0 /*49979*/;
assign oneWire = 1'b1 /*49979*/;
assign _67_ = ~D[0] /*49593*/;
assign _65_ = R_0[63] | _67_ /*49590*/;
assign _66_ = R_0[63] ^ _67_ /*49592*/;
assign _0_ = ~_66_ /*49591*/;
assign _74_ = ~D[1] /*49589*/;
assign _71_ = R_0[64] & _74_ /*49585*/;
assign _72_ = R_0[64] ^ _74_ /*49588*/;
assign _73_ = _65_ & _72_ /*49586*/;
assign _70_ = _71_ | _73_ /*49584*/;
assign _1_ = _65_ ^ _72_ /*49587*/;
assign _79_ = ~D[2] /*49583*/;
assign _76_ = R_0[65] & _79_ /*49579*/;
assign _77_ = R_0[65] ^ _79_ /*49582*/;
assign _78_ = _70_ & _77_ /*49580*/;
assign _75_ = _76_ | _78_ /*49578*/;
assign _2_ = _70_ ^ _77_ /*49581*/;
assign _84_ = ~D[3] /*49577*/;
assign _81_ = R_0[66] & _84_ /*49573*/;
assign _82_ = R_0[66] ^ _84_ /*49576*/;
assign _83_ = _75_ & _82_ /*49574*/;
assign _80_ = _81_ | _83_ /*49572*/;
assign _3_ = _75_ ^ _82_ /*49575*/;
assign _89_ = ~D[4] /*49571*/;
assign _86_ = R_0[67] & _89_ /*49567*/;
assign _87_ = R_0[67] ^ _89_ /*49570*/;
assign _88_ = _80_ & _87_ /*49568*/;
assign _85_ = _86_ | _88_ /*49566*/;
assign _4_ = _80_ ^ _87_ /*49569*/;
assign _94_ = ~D[5] /*49565*/;
assign _91_ = R_0[68] & _94_ /*49561*/;
assign _92_ = R_0[68] ^ _94_ /*49564*/;
assign _93_ = _85_ & _92_ /*49562*/;
assign _90_ = _91_ | _93_ /*49560*/;
assign _5_ = _85_ ^ _92_ /*49563*/;
assign _99_ = ~D[6] /*49559*/;
assign _96_ = R_0[69] & _99_ /*49555*/;
assign _97_ = R_0[69] ^ _99_ /*49558*/;
assign _98_ = _90_ & _97_ /*49556*/;
assign _95_ = _96_ | _98_ /*49554*/;
assign _6_ = _90_ ^ _97_ /*49557*/;
assign _104_ = ~D[7] /*49553*/;
assign _101_ = R_0[70] & _104_ /*49549*/;
assign _102_ = R_0[70] ^ _104_ /*49552*/;
assign _103_ = _95_ & _102_ /*49550*/;
assign _100_ = _101_ | _103_ /*49548*/;
assign _7_ = _95_ ^ _102_ /*49551*/;
assign _109_ = ~D[8] /*49547*/;
assign _106_ = R_0[71] & _109_ /*49543*/;
assign _107_ = R_0[71] ^ _109_ /*49546*/;
assign _108_ = _100_ & _107_ /*49544*/;
assign _105_ = _106_ | _108_ /*49542*/;
assign _8_ = _100_ ^ _107_ /*49545*/;
assign _114_ = ~D[9] /*49541*/;
assign _111_ = R_0[72] & _114_ /*49537*/;
assign _112_ = R_0[72] ^ _114_ /*49540*/;
assign _113_ = _105_ & _112_ /*49538*/;
assign _110_ = _111_ | _113_ /*49536*/;
assign _9_ = _105_ ^ _112_ /*49539*/;
assign _119_ = ~D[10] /*49535*/;
assign _116_ = R_0[73] & _119_ /*49531*/;
assign _117_ = R_0[73] ^ _119_ /*49534*/;
assign _118_ = _110_ & _117_ /*49532*/;
assign _115_ = _116_ | _118_ /*49530*/;
assign _10_ = _110_ ^ _117_ /*49533*/;
assign _124_ = ~D[11] /*49529*/;
assign _121_ = R_0[74] & _124_ /*49525*/;
assign _122_ = R_0[74] ^ _124_ /*49528*/;
assign _123_ = _115_ & _122_ /*49526*/;
assign _120_ = _121_ | _123_ /*49524*/;
assign _11_ = _115_ ^ _122_ /*49527*/;
assign _129_ = ~D[12] /*49523*/;
assign _126_ = R_0[75] & _129_ /*49519*/;
assign _127_ = R_0[75] ^ _129_ /*49522*/;
assign _128_ = _120_ & _127_ /*49520*/;
assign _125_ = _126_ | _128_ /*49518*/;
assign _12_ = _120_ ^ _127_ /*49521*/;
assign _134_ = ~D[13] /*49517*/;
assign _131_ = R_0[76] & _134_ /*49513*/;
assign _132_ = R_0[76] ^ _134_ /*49516*/;
assign _133_ = _125_ & _132_ /*49514*/;
assign _130_ = _131_ | _133_ /*49512*/;
assign _13_ = _125_ ^ _132_ /*49515*/;
assign _139_ = ~D[14] /*49511*/;
assign _136_ = R_0[77] & _139_ /*49507*/;
assign _137_ = R_0[77] ^ _139_ /*49510*/;
assign _138_ = _130_ & _137_ /*49508*/;
assign _135_ = _136_ | _138_ /*49506*/;
assign _14_ = _130_ ^ _137_ /*49509*/;
assign _144_ = ~D[15] /*49505*/;
assign _141_ = R_0[78] & _144_ /*49501*/;
assign _142_ = R_0[78] ^ _144_ /*49504*/;
assign _143_ = _135_ & _142_ /*49502*/;
assign _140_ = _141_ | _143_ /*49500*/;
assign _15_ = _135_ ^ _142_ /*49503*/;
assign _149_ = ~D[16] /*49499*/;
assign _146_ = R_0[79] & _149_ /*49495*/;
assign _147_ = R_0[79] ^ _149_ /*49498*/;
assign _148_ = _140_ & _147_ /*49496*/;
assign _145_ = _146_ | _148_ /*49494*/;
assign _16_ = _140_ ^ _147_ /*49497*/;
assign _154_ = ~D[17] /*49493*/;
assign _151_ = R_0[80] & _154_ /*49489*/;
assign _152_ = R_0[80] ^ _154_ /*49492*/;
assign _153_ = _145_ & _152_ /*49490*/;
assign _150_ = _151_ | _153_ /*49488*/;
assign _17_ = _145_ ^ _152_ /*49491*/;
assign _159_ = ~D[18] /*49487*/;
assign _156_ = R_0[81] & _159_ /*49483*/;
assign _157_ = R_0[81] ^ _159_ /*49486*/;
assign _158_ = _150_ & _157_ /*49484*/;
assign _155_ = _156_ | _158_ /*49482*/;
assign _18_ = _150_ ^ _157_ /*49485*/;
assign _164_ = ~D[19] /*49481*/;
assign _161_ = R_0[82] & _164_ /*49477*/;
assign _162_ = R_0[82] ^ _164_ /*49480*/;
assign _163_ = _155_ & _162_ /*49478*/;
assign _160_ = _161_ | _163_ /*49476*/;
assign _19_ = _155_ ^ _162_ /*49479*/;
assign _169_ = ~D[20] /*49475*/;
assign _166_ = R_0[83] & _169_ /*49471*/;
assign _167_ = R_0[83] ^ _169_ /*49474*/;
assign _168_ = _160_ & _167_ /*49472*/;
assign _165_ = _166_ | _168_ /*49470*/;
assign _20_ = _160_ ^ _167_ /*49473*/;
assign _174_ = ~D[21] /*49469*/;
assign _171_ = R_0[84] & _174_ /*49465*/;
assign _172_ = R_0[84] ^ _174_ /*49468*/;
assign _173_ = _165_ & _172_ /*49466*/;
assign _170_ = _171_ | _173_ /*49464*/;
assign _21_ = _165_ ^ _172_ /*49467*/;
assign _179_ = ~D[22] /*49463*/;
assign _176_ = R_0[85] & _179_ /*49459*/;
assign _177_ = R_0[85] ^ _179_ /*49462*/;
assign _178_ = _170_ & _177_ /*49460*/;
assign _175_ = _176_ | _178_ /*49458*/;
assign _22_ = _170_ ^ _177_ /*49461*/;
assign _184_ = ~D[23] /*49457*/;
assign _181_ = R_0[86] & _184_ /*49453*/;
assign _182_ = R_0[86] ^ _184_ /*49456*/;
assign _183_ = _175_ & _182_ /*49454*/;
assign _180_ = _181_ | _183_ /*49452*/;
assign _23_ = _175_ ^ _182_ /*49455*/;
assign _189_ = ~D[24] /*49451*/;
assign _186_ = R_0[87] & _189_ /*49447*/;
assign _187_ = R_0[87] ^ _189_ /*49450*/;
assign _188_ = _180_ & _187_ /*49448*/;
assign _185_ = _186_ | _188_ /*49446*/;
assign _24_ = _180_ ^ _187_ /*49449*/;
assign _194_ = ~D[25] /*49445*/;
assign _191_ = R_0[88] & _194_ /*49441*/;
assign _192_ = R_0[88] ^ _194_ /*49444*/;
assign _193_ = _185_ & _192_ /*49442*/;
assign _190_ = _191_ | _193_ /*49440*/;
assign _25_ = _185_ ^ _192_ /*49443*/;
assign _199_ = ~D[26] /*49439*/;
assign _196_ = R_0[89] & _199_ /*49435*/;
assign _197_ = R_0[89] ^ _199_ /*49438*/;
assign _198_ = _190_ & _197_ /*49436*/;
assign _195_ = _196_ | _198_ /*49434*/;
assign _26_ = _190_ ^ _197_ /*49437*/;
assign _204_ = ~D[27] /*49433*/;
assign _201_ = R_0[90] & _204_ /*49429*/;
assign _202_ = R_0[90] ^ _204_ /*49432*/;
assign _203_ = _195_ & _202_ /*49430*/;
assign _200_ = _201_ | _203_ /*49428*/;
assign _27_ = _195_ ^ _202_ /*49431*/;
assign _209_ = ~D[28] /*49427*/;
assign _206_ = R_0[91] & _209_ /*49423*/;
assign _207_ = R_0[91] ^ _209_ /*49426*/;
assign _208_ = _200_ & _207_ /*49424*/;
assign _205_ = _206_ | _208_ /*49422*/;
assign _28_ = _200_ ^ _207_ /*49425*/;
assign _214_ = ~D[29] /*49421*/;
assign _211_ = R_0[92] & _214_ /*49417*/;
assign _212_ = R_0[92] ^ _214_ /*49420*/;
assign _213_ = _205_ & _212_ /*49418*/;
assign _210_ = _211_ | _213_ /*49416*/;
assign _29_ = _205_ ^ _212_ /*49419*/;
assign _219_ = ~D[30] /*49415*/;
assign _216_ = R_0[93] & _219_ /*49411*/;
assign _217_ = R_0[93] ^ _219_ /*49414*/;
assign _218_ = _210_ & _217_ /*49412*/;
assign _215_ = _216_ | _218_ /*49410*/;
assign _30_ = _210_ ^ _217_ /*49413*/;
assign _224_ = ~D[31] /*49409*/;
assign _221_ = R_0[94] & _224_ /*49405*/;
assign _222_ = R_0[94] ^ _224_ /*49408*/;
assign _223_ = _215_ & _222_ /*49406*/;
assign _220_ = _221_ | _223_ /*49404*/;
assign _31_ = _215_ ^ _222_ /*49407*/;
assign _229_ = ~D[32] /*49403*/;
assign _226_ = R_0[95] & _229_ /*49399*/;
assign _227_ = R_0[95] ^ _229_ /*49402*/;
assign _228_ = _220_ & _227_ /*49400*/;
assign _225_ = _226_ | _228_ /*49398*/;
assign _32_ = _220_ ^ _227_ /*49401*/;
assign _234_ = ~D[33] /*49397*/;
assign _231_ = R_0[96] & _234_ /*49393*/;
assign _232_ = R_0[96] ^ _234_ /*49396*/;
assign _233_ = _225_ & _232_ /*49394*/;
assign _230_ = _231_ | _233_ /*49392*/;
assign _33_ = _225_ ^ _232_ /*49395*/;
assign _239_ = ~D[34] /*49391*/;
assign _236_ = R_0[97] & _239_ /*49387*/;
assign _237_ = R_0[97] ^ _239_ /*49390*/;
assign _238_ = _230_ & _237_ /*49388*/;
assign _235_ = _236_ | _238_ /*49386*/;
assign _34_ = _230_ ^ _237_ /*49389*/;
assign _244_ = ~D[35] /*49385*/;
assign _241_ = R_0[98] & _244_ /*49381*/;
assign _242_ = R_0[98] ^ _244_ /*49384*/;
assign _243_ = _235_ & _242_ /*49382*/;
assign _240_ = _241_ | _243_ /*49380*/;
assign _35_ = _235_ ^ _242_ /*49383*/;
assign _249_ = ~D[36] /*49379*/;
assign _246_ = R_0[99] & _249_ /*49375*/;
assign _247_ = R_0[99] ^ _249_ /*49378*/;
assign _248_ = _240_ & _247_ /*49376*/;
assign _245_ = _246_ | _248_ /*49374*/;
assign _36_ = _240_ ^ _247_ /*49377*/;
assign _254_ = ~D[37] /*49373*/;
assign _251_ = R_0[100] & _254_ /*49369*/;
assign _252_ = R_0[100] ^ _254_ /*49372*/;
assign _253_ = _245_ & _252_ /*49370*/;
assign _250_ = _251_ | _253_ /*49368*/;
assign _37_ = _245_ ^ _252_ /*49371*/;
assign _259_ = ~D[38] /*49367*/;
assign _256_ = R_0[101] & _259_ /*49363*/;
assign _257_ = R_0[101] ^ _259_ /*49366*/;
assign _258_ = _250_ & _257_ /*49364*/;
assign _255_ = _256_ | _258_ /*49362*/;
assign _38_ = _250_ ^ _257_ /*49365*/;
assign _264_ = ~D[39] /*49361*/;
assign _261_ = R_0[102] & _264_ /*49357*/;
assign _262_ = R_0[102] ^ _264_ /*49360*/;
assign _263_ = _255_ & _262_ /*49358*/;
assign _260_ = _261_ | _263_ /*49356*/;
assign _39_ = _255_ ^ _262_ /*49359*/;
assign _269_ = ~D[40] /*49355*/;
assign _266_ = R_0[103] & _269_ /*49351*/;
assign _267_ = R_0[103] ^ _269_ /*49354*/;
assign _268_ = _260_ & _267_ /*49352*/;
assign _265_ = _266_ | _268_ /*49350*/;
assign _40_ = _260_ ^ _267_ /*49353*/;
assign _274_ = ~D[41] /*49349*/;
assign _271_ = R_0[104] & _274_ /*49345*/;
assign _272_ = R_0[104] ^ _274_ /*49348*/;
assign _273_ = _265_ & _272_ /*49346*/;
assign _270_ = _271_ | _273_ /*49344*/;
assign _41_ = _265_ ^ _272_ /*49347*/;
assign _279_ = ~D[42] /*49343*/;
assign _276_ = R_0[105] & _279_ /*49339*/;
assign _277_ = R_0[105] ^ _279_ /*49342*/;
assign _278_ = _270_ & _277_ /*49340*/;
assign _275_ = _276_ | _278_ /*49338*/;
assign _42_ = _270_ ^ _277_ /*49341*/;
assign _284_ = ~D[43] /*49337*/;
assign _281_ = R_0[106] & _284_ /*49333*/;
assign _282_ = R_0[106] ^ _284_ /*49336*/;
assign _283_ = _275_ & _282_ /*49334*/;
assign _280_ = _281_ | _283_ /*49332*/;
assign _43_ = _275_ ^ _282_ /*49335*/;
assign _289_ = ~D[44] /*49331*/;
assign _286_ = R_0[107] & _289_ /*49327*/;
assign _287_ = R_0[107] ^ _289_ /*49330*/;
assign _288_ = _280_ & _287_ /*49328*/;
assign _285_ = _286_ | _288_ /*49326*/;
assign _44_ = _280_ ^ _287_ /*49329*/;
assign _294_ = ~D[45] /*49325*/;
assign _291_ = R_0[108] & _294_ /*49321*/;
assign _292_ = R_0[108] ^ _294_ /*49324*/;
assign _293_ = _285_ & _292_ /*49322*/;
assign _290_ = _291_ | _293_ /*49320*/;
assign _45_ = _285_ ^ _292_ /*49323*/;
assign _299_ = ~D[46] /*49319*/;
assign _296_ = R_0[109] & _299_ /*49315*/;
assign _297_ = R_0[109] ^ _299_ /*49318*/;
assign _298_ = _290_ & _297_ /*49316*/;
assign _295_ = _296_ | _298_ /*49314*/;
assign _46_ = _290_ ^ _297_ /*49317*/;
assign _304_ = ~D[47] /*49313*/;
assign _301_ = R_0[110] & _304_ /*49309*/;
assign _302_ = R_0[110] ^ _304_ /*49312*/;
assign _303_ = _295_ & _302_ /*49310*/;
assign _300_ = _301_ | _303_ /*49308*/;
assign _47_ = _295_ ^ _302_ /*49311*/;
assign _309_ = ~D[48] /*49307*/;
assign _306_ = R_0[111] & _309_ /*49303*/;
assign _307_ = R_0[111] ^ _309_ /*49306*/;
assign _308_ = _300_ & _307_ /*49304*/;
assign _305_ = _306_ | _308_ /*49302*/;
assign _48_ = _300_ ^ _307_ /*49305*/;
assign _314_ = ~D[49] /*49301*/;
assign _311_ = R_0[112] & _314_ /*49297*/;
assign _312_ = R_0[112] ^ _314_ /*49300*/;
assign _313_ = _305_ & _312_ /*49298*/;
assign _310_ = _311_ | _313_ /*49296*/;
assign _49_ = _305_ ^ _312_ /*49299*/;
assign _319_ = ~D[50] /*49295*/;
assign _316_ = R_0[113] & _319_ /*49291*/;
assign _317_ = R_0[113] ^ _319_ /*49294*/;
assign _318_ = _310_ & _317_ /*49292*/;
assign _315_ = _316_ | _318_ /*49290*/;
assign _50_ = _310_ ^ _317_ /*49293*/;
assign _324_ = ~D[51] /*49289*/;
assign _321_ = R_0[114] & _324_ /*49285*/;
assign _322_ = R_0[114] ^ _324_ /*49288*/;
assign _323_ = _315_ & _322_ /*49286*/;
assign _320_ = _321_ | _323_ /*49284*/;
assign _51_ = _315_ ^ _322_ /*49287*/;
assign _329_ = ~D[52] /*49283*/;
assign _326_ = R_0[115] & _329_ /*49279*/;
assign _327_ = R_0[115] ^ _329_ /*49282*/;
assign _328_ = _320_ & _327_ /*49280*/;
assign _325_ = _326_ | _328_ /*49278*/;
assign _52_ = _320_ ^ _327_ /*49281*/;
assign _334_ = ~D[53] /*49277*/;
assign _331_ = R_0[116] & _334_ /*49273*/;
assign _332_ = R_0[116] ^ _334_ /*49276*/;
assign _333_ = _325_ & _332_ /*49274*/;
assign _330_ = _331_ | _333_ /*49272*/;
assign _53_ = _325_ ^ _332_ /*49275*/;
assign _339_ = ~D[54] /*49271*/;
assign _336_ = R_0[117] & _339_ /*49267*/;
assign _337_ = R_0[117] ^ _339_ /*49270*/;
assign _338_ = _330_ & _337_ /*49268*/;
assign _335_ = _336_ | _338_ /*49266*/;
assign _54_ = _330_ ^ _337_ /*49269*/;
assign _344_ = ~D[55] /*49265*/;
assign _341_ = R_0[118] & _344_ /*49261*/;
assign _342_ = R_0[118] ^ _344_ /*49264*/;
assign _343_ = _335_ & _342_ /*49262*/;
assign _340_ = _341_ | _343_ /*49260*/;
assign _55_ = _335_ ^ _342_ /*49263*/;
assign _349_ = ~D[56] /*49259*/;
assign _346_ = R_0[119] & _349_ /*49255*/;
assign _347_ = R_0[119] ^ _349_ /*49258*/;
assign _348_ = _340_ & _347_ /*49256*/;
assign _345_ = _346_ | _348_ /*49254*/;
assign _56_ = _340_ ^ _347_ /*49257*/;
assign _354_ = ~D[57] /*49253*/;
assign _351_ = R_0[120] & _354_ /*49249*/;
assign _352_ = R_0[120] ^ _354_ /*49252*/;
assign _353_ = _345_ & _352_ /*49250*/;
assign _350_ = _351_ | _353_ /*49248*/;
assign _57_ = _345_ ^ _352_ /*49251*/;
assign _359_ = ~D[58] /*49247*/;
assign _356_ = R_0[121] & _359_ /*49243*/;
assign _357_ = R_0[121] ^ _359_ /*49246*/;
assign _358_ = _350_ & _357_ /*49244*/;
assign _355_ = _356_ | _358_ /*49242*/;
assign _58_ = _350_ ^ _357_ /*49245*/;
assign _364_ = ~D[59] /*49241*/;
assign _361_ = R_0[122] & _364_ /*49237*/;
assign _362_ = R_0[122] ^ _364_ /*49240*/;
assign _363_ = _355_ & _362_ /*49238*/;
assign _360_ = _361_ | _363_ /*49236*/;
assign _59_ = _355_ ^ _362_ /*49239*/;
assign _369_ = ~D[60] /*49235*/;
assign _366_ = R_0[123] & _369_ /*49231*/;
assign _367_ = R_0[123] ^ _369_ /*49234*/;
assign _368_ = _360_ & _367_ /*49232*/;
assign _365_ = _366_ | _368_ /*49230*/;
assign _60_ = _360_ ^ _367_ /*49233*/;
assign _374_ = ~D[61] /*49229*/;
assign _371_ = R_0[124] & _374_ /*49225*/;
assign _372_ = R_0[124] ^ _374_ /*49228*/;
assign _373_ = _365_ & _372_ /*49226*/;
assign _370_ = _371_ | _373_ /*49224*/;
assign _61_ = _365_ ^ _372_ /*49227*/;
assign _379_ = ~D[62] /*49223*/;
assign _376_ = R_0[125] & _379_ /*49219*/;
assign _377_ = R_0[125] ^ _379_ /*49222*/;
assign _378_ = _370_ & _377_ /*49220*/;
assign _375_ = _376_ | _378_ /*49218*/;
assign _62_ = _370_ ^ _377_ /*49221*/;
assign _380_ = zeroWire & oneWire /*49213*/;
assign _381_ = zeroWire ^ oneWire /*49216*/;
assign _382_ = _375_ & _381_ /*49214*/;
assign Q[63] = _380_ | _382_ /*49212*/;
assign _63_ = _375_ ^ _381_ /*49215*/;
assign _454_ = D[0] ^ Q[63] /*48826*/;
assign _451_ = R_0[62] & _454_ /*48822*/;
assign _452_ = R_0[62] ^ _454_ /*48825*/;
assign _453_ = Q[63] & _452_ /*48823*/;
assign _450_ = _451_ | _453_ /*48821*/;
assign _385_ = Q[63] ^ _452_ /*48824*/;
assign _459_ = D[1] ^ Q[63] /*48820*/;
assign _456_ = _0_ & _459_ /*48816*/;
assign _457_ = _0_ ^ _459_ /*48819*/;
assign _458_ = _450_ & _457_ /*48817*/;
assign _455_ = _456_ | _458_ /*48815*/;
assign _386_ = _450_ ^ _457_ /*48818*/;
assign _464_ = D[2] ^ Q[63] /*48814*/;
assign _461_ = _1_ & _464_ /*48810*/;
assign _462_ = _1_ ^ _464_ /*48813*/;
assign _463_ = _455_ & _462_ /*48811*/;
assign _460_ = _461_ | _463_ /*48809*/;
assign _387_ = _455_ ^ _462_ /*48812*/;
assign _469_ = D[3] ^ Q[63] /*48808*/;
assign _466_ = _2_ & _469_ /*48804*/;
assign _467_ = _2_ ^ _469_ /*48807*/;
assign _468_ = _460_ & _467_ /*48805*/;
assign _465_ = _466_ | _468_ /*48803*/;
assign _388_ = _460_ ^ _467_ /*48806*/;
assign _474_ = D[4] ^ Q[63] /*48802*/;
assign _471_ = _3_ & _474_ /*48798*/;
assign _472_ = _3_ ^ _474_ /*48801*/;
assign _473_ = _465_ & _472_ /*48799*/;
assign _470_ = _471_ | _473_ /*48797*/;
assign _389_ = _465_ ^ _472_ /*48800*/;
assign _479_ = D[5] ^ Q[63] /*48796*/;
assign _476_ = _4_ & _479_ /*48792*/;
assign _477_ = _4_ ^ _479_ /*48795*/;
assign _478_ = _470_ & _477_ /*48793*/;
assign _475_ = _476_ | _478_ /*48791*/;
assign _390_ = _470_ ^ _477_ /*48794*/;
assign _484_ = D[6] ^ Q[63] /*48790*/;
assign _481_ = _5_ & _484_ /*48786*/;
assign _482_ = _5_ ^ _484_ /*48789*/;
assign _483_ = _475_ & _482_ /*48787*/;
assign _480_ = _481_ | _483_ /*48785*/;
assign _391_ = _475_ ^ _482_ /*48788*/;
assign _489_ = D[7] ^ Q[63] /*48784*/;
assign _486_ = _6_ & _489_ /*48780*/;
assign _487_ = _6_ ^ _489_ /*48783*/;
assign _488_ = _480_ & _487_ /*48781*/;
assign _485_ = _486_ | _488_ /*48779*/;
assign _392_ = _480_ ^ _487_ /*48782*/;
assign _494_ = D[8] ^ Q[63] /*48778*/;
assign _491_ = _7_ & _494_ /*48774*/;
assign _492_ = _7_ ^ _494_ /*48777*/;
assign _493_ = _485_ & _492_ /*48775*/;
assign _490_ = _491_ | _493_ /*48773*/;
assign _393_ = _485_ ^ _492_ /*48776*/;
assign _499_ = D[9] ^ Q[63] /*48772*/;
assign _496_ = _8_ & _499_ /*48768*/;
assign _497_ = _8_ ^ _499_ /*48771*/;
assign _498_ = _490_ & _497_ /*48769*/;
assign _495_ = _496_ | _498_ /*48767*/;
assign _394_ = _490_ ^ _497_ /*48770*/;
assign _504_ = D[10] ^ Q[63] /*48766*/;
assign _501_ = _9_ & _504_ /*48762*/;
assign _502_ = _9_ ^ _504_ /*48765*/;
assign _503_ = _495_ & _502_ /*48763*/;
assign _500_ = _501_ | _503_ /*48761*/;
assign _395_ = _495_ ^ _502_ /*48764*/;
assign _509_ = D[11] ^ Q[63] /*48760*/;
assign _506_ = _10_ & _509_ /*48756*/;
assign _507_ = _10_ ^ _509_ /*48759*/;
assign _508_ = _500_ & _507_ /*48757*/;
assign _505_ = _506_ | _508_ /*48755*/;
assign _396_ = _500_ ^ _507_ /*48758*/;
assign _514_ = D[12] ^ Q[63] /*48754*/;
assign _511_ = _11_ & _514_ /*48750*/;
assign _512_ = _11_ ^ _514_ /*48753*/;
assign _513_ = _505_ & _512_ /*48751*/;
assign _510_ = _511_ | _513_ /*48749*/;
assign _397_ = _505_ ^ _512_ /*48752*/;
assign _519_ = D[13] ^ Q[63] /*48748*/;
assign _516_ = _12_ & _519_ /*48744*/;
assign _517_ = _12_ ^ _519_ /*48747*/;
assign _518_ = _510_ & _517_ /*48745*/;
assign _515_ = _516_ | _518_ /*48743*/;
assign _398_ = _510_ ^ _517_ /*48746*/;
assign _524_ = D[14] ^ Q[63] /*48742*/;
assign _521_ = _13_ & _524_ /*48738*/;
assign _522_ = _13_ ^ _524_ /*48741*/;
assign _523_ = _515_ & _522_ /*48739*/;
assign _520_ = _521_ | _523_ /*48737*/;
assign _399_ = _515_ ^ _522_ /*48740*/;
assign _529_ = D[15] ^ Q[63] /*48736*/;
assign _526_ = _14_ & _529_ /*48732*/;
assign _527_ = _14_ ^ _529_ /*48735*/;
assign _528_ = _520_ & _527_ /*48733*/;
assign _525_ = _526_ | _528_ /*48731*/;
assign _400_ = _520_ ^ _527_ /*48734*/;
assign _534_ = D[16] ^ Q[63] /*48730*/;
assign _531_ = _15_ & _534_ /*48726*/;
assign _532_ = _15_ ^ _534_ /*48729*/;
assign _533_ = _525_ & _532_ /*48727*/;
assign _530_ = _531_ | _533_ /*48725*/;
assign _401_ = _525_ ^ _532_ /*48728*/;
assign _539_ = D[17] ^ Q[63] /*48724*/;
assign _536_ = _16_ & _539_ /*48720*/;
assign _537_ = _16_ ^ _539_ /*48723*/;
assign _538_ = _530_ & _537_ /*48721*/;
assign _535_ = _536_ | _538_ /*48719*/;
assign _402_ = _530_ ^ _537_ /*48722*/;
assign _544_ = D[18] ^ Q[63] /*48718*/;
assign _541_ = _17_ & _544_ /*48714*/;
assign _542_ = _17_ ^ _544_ /*48717*/;
assign _543_ = _535_ & _542_ /*48715*/;
assign _540_ = _541_ | _543_ /*48713*/;
assign _403_ = _535_ ^ _542_ /*48716*/;
assign _549_ = D[19] ^ Q[63] /*48712*/;
assign _546_ = _18_ & _549_ /*48708*/;
assign _547_ = _18_ ^ _549_ /*48711*/;
assign _548_ = _540_ & _547_ /*48709*/;
assign _545_ = _546_ | _548_ /*48707*/;
assign _404_ = _540_ ^ _547_ /*48710*/;
assign _554_ = D[20] ^ Q[63] /*48706*/;
assign _551_ = _19_ & _554_ /*48702*/;
assign _552_ = _19_ ^ _554_ /*48705*/;
assign _553_ = _545_ & _552_ /*48703*/;
assign _550_ = _551_ | _553_ /*48701*/;
assign _405_ = _545_ ^ _552_ /*48704*/;
assign _559_ = D[21] ^ Q[63] /*48700*/;
assign _556_ = _20_ & _559_ /*48696*/;
assign _557_ = _20_ ^ _559_ /*48699*/;
assign _558_ = _550_ & _557_ /*48697*/;
assign _555_ = _556_ | _558_ /*48695*/;
assign _406_ = _550_ ^ _557_ /*48698*/;
assign _564_ = D[22] ^ Q[63] /*48694*/;
assign _561_ = _21_ & _564_ /*48690*/;
assign _562_ = _21_ ^ _564_ /*48693*/;
assign _563_ = _555_ & _562_ /*48691*/;
assign _560_ = _561_ | _563_ /*48689*/;
assign _407_ = _555_ ^ _562_ /*48692*/;
assign _569_ = D[23] ^ Q[63] /*48688*/;
assign _566_ = _22_ & _569_ /*48684*/;
assign _567_ = _22_ ^ _569_ /*48687*/;
assign _568_ = _560_ & _567_ /*48685*/;
assign _565_ = _566_ | _568_ /*48683*/;
assign _408_ = _560_ ^ _567_ /*48686*/;
assign _574_ = D[24] ^ Q[63] /*48682*/;
assign _571_ = _23_ & _574_ /*48678*/;
assign _572_ = _23_ ^ _574_ /*48681*/;
assign _573_ = _565_ & _572_ /*48679*/;
assign _570_ = _571_ | _573_ /*48677*/;
assign _409_ = _565_ ^ _572_ /*48680*/;
assign _579_ = D[25] ^ Q[63] /*48676*/;
assign _576_ = _24_ & _579_ /*48672*/;
assign _577_ = _24_ ^ _579_ /*48675*/;
assign _578_ = _570_ & _577_ /*48673*/;
assign _575_ = _576_ | _578_ /*48671*/;
assign _410_ = _570_ ^ _577_ /*48674*/;
assign _584_ = D[26] ^ Q[63] /*48670*/;
assign _581_ = _25_ & _584_ /*48666*/;
assign _582_ = _25_ ^ _584_ /*48669*/;
assign _583_ = _575_ & _582_ /*48667*/;
assign _580_ = _581_ | _583_ /*48665*/;
assign _411_ = _575_ ^ _582_ /*48668*/;
assign _589_ = D[27] ^ Q[63] /*48664*/;
assign _586_ = _26_ & _589_ /*48660*/;
assign _587_ = _26_ ^ _589_ /*48663*/;
assign _588_ = _580_ & _587_ /*48661*/;
assign _585_ = _586_ | _588_ /*48659*/;
assign _412_ = _580_ ^ _587_ /*48662*/;
assign _594_ = D[28] ^ Q[63] /*48658*/;
assign _591_ = _27_ & _594_ /*48654*/;
assign _592_ = _27_ ^ _594_ /*48657*/;
assign _593_ = _585_ & _592_ /*48655*/;
assign _590_ = _591_ | _593_ /*48653*/;
assign _413_ = _585_ ^ _592_ /*48656*/;
assign _599_ = D[29] ^ Q[63] /*48652*/;
assign _596_ = _28_ & _599_ /*48648*/;
assign _597_ = _28_ ^ _599_ /*48651*/;
assign _598_ = _590_ & _597_ /*48649*/;
assign _595_ = _596_ | _598_ /*48647*/;
assign _414_ = _590_ ^ _597_ /*48650*/;
assign _604_ = D[30] ^ Q[63] /*48646*/;
assign _601_ = _29_ & _604_ /*48642*/;
assign _602_ = _29_ ^ _604_ /*48645*/;
assign _603_ = _595_ & _602_ /*48643*/;
assign _600_ = _601_ | _603_ /*48641*/;
assign _415_ = _595_ ^ _602_ /*48644*/;
assign _609_ = D[31] ^ Q[63] /*48640*/;
assign _606_ = _30_ & _609_ /*48636*/;
assign _607_ = _30_ ^ _609_ /*48639*/;
assign _608_ = _600_ & _607_ /*48637*/;
assign _605_ = _606_ | _608_ /*48635*/;
assign _416_ = _600_ ^ _607_ /*48638*/;
assign _614_ = D[32] ^ Q[63] /*48634*/;
assign _611_ = _31_ & _614_ /*48630*/;
assign _612_ = _31_ ^ _614_ /*48633*/;
assign _613_ = _605_ & _612_ /*48631*/;
assign _610_ = _611_ | _613_ /*48629*/;
assign _417_ = _605_ ^ _612_ /*48632*/;
assign _619_ = D[33] ^ Q[63] /*48628*/;
assign _616_ = _32_ & _619_ /*48624*/;
assign _617_ = _32_ ^ _619_ /*48627*/;
assign _618_ = _610_ & _617_ /*48625*/;
assign _615_ = _616_ | _618_ /*48623*/;
assign _418_ = _610_ ^ _617_ /*48626*/;
assign _624_ = D[34] ^ Q[63] /*48622*/;
assign _621_ = _33_ & _624_ /*48618*/;
assign _622_ = _33_ ^ _624_ /*48621*/;
assign _623_ = _615_ & _622_ /*48619*/;
assign _620_ = _621_ | _623_ /*48617*/;
assign _419_ = _615_ ^ _622_ /*48620*/;
assign _629_ = D[35] ^ Q[63] /*48616*/;
assign _626_ = _34_ & _629_ /*48612*/;
assign _627_ = _34_ ^ _629_ /*48615*/;
assign _628_ = _620_ & _627_ /*48613*/;
assign _625_ = _626_ | _628_ /*48611*/;
assign _420_ = _620_ ^ _627_ /*48614*/;
assign _634_ = D[36] ^ Q[63] /*48610*/;
assign _631_ = _35_ & _634_ /*48606*/;
assign _632_ = _35_ ^ _634_ /*48609*/;
assign _633_ = _625_ & _632_ /*48607*/;
assign _630_ = _631_ | _633_ /*48605*/;
assign _421_ = _625_ ^ _632_ /*48608*/;
assign _639_ = D[37] ^ Q[63] /*48604*/;
assign _636_ = _36_ & _639_ /*48600*/;
assign _637_ = _36_ ^ _639_ /*48603*/;
assign _638_ = _630_ & _637_ /*48601*/;
assign _635_ = _636_ | _638_ /*48599*/;
assign _422_ = _630_ ^ _637_ /*48602*/;
assign _644_ = D[38] ^ Q[63] /*48598*/;
assign _641_ = _37_ & _644_ /*48594*/;
assign _642_ = _37_ ^ _644_ /*48597*/;
assign _643_ = _635_ & _642_ /*48595*/;
assign _640_ = _641_ | _643_ /*48593*/;
assign _423_ = _635_ ^ _642_ /*48596*/;
assign _649_ = D[39] ^ Q[63] /*48592*/;
assign _646_ = _38_ & _649_ /*48588*/;
assign _647_ = _38_ ^ _649_ /*48591*/;
assign _648_ = _640_ & _647_ /*48589*/;
assign _645_ = _646_ | _648_ /*48587*/;
assign _424_ = _640_ ^ _647_ /*48590*/;
assign _654_ = D[40] ^ Q[63] /*48586*/;
assign _651_ = _39_ & _654_ /*48582*/;
assign _652_ = _39_ ^ _654_ /*48585*/;
assign _653_ = _645_ & _652_ /*48583*/;
assign _650_ = _651_ | _653_ /*48581*/;
assign _425_ = _645_ ^ _652_ /*48584*/;
assign _659_ = D[41] ^ Q[63] /*48580*/;
assign _656_ = _40_ & _659_ /*48576*/;
assign _657_ = _40_ ^ _659_ /*48579*/;
assign _658_ = _650_ & _657_ /*48577*/;
assign _655_ = _656_ | _658_ /*48575*/;
assign _426_ = _650_ ^ _657_ /*48578*/;
assign _664_ = D[42] ^ Q[63] /*48574*/;
assign _661_ = _41_ & _664_ /*48570*/;
assign _662_ = _41_ ^ _664_ /*48573*/;
assign _663_ = _655_ & _662_ /*48571*/;
assign _660_ = _661_ | _663_ /*48569*/;
assign _427_ = _655_ ^ _662_ /*48572*/;
assign _669_ = D[43] ^ Q[63] /*48568*/;
assign _666_ = _42_ & _669_ /*48564*/;
assign _667_ = _42_ ^ _669_ /*48567*/;
assign _668_ = _660_ & _667_ /*48565*/;
assign _665_ = _666_ | _668_ /*48563*/;
assign _428_ = _660_ ^ _667_ /*48566*/;
assign _674_ = D[44] ^ Q[63] /*48562*/;
assign _671_ = _43_ & _674_ /*48558*/;
assign _672_ = _43_ ^ _674_ /*48561*/;
assign _673_ = _665_ & _672_ /*48559*/;
assign _670_ = _671_ | _673_ /*48557*/;
assign _429_ = _665_ ^ _672_ /*48560*/;
assign _679_ = D[45] ^ Q[63] /*48556*/;
assign _676_ = _44_ & _679_ /*48552*/;
assign _677_ = _44_ ^ _679_ /*48555*/;
assign _678_ = _670_ & _677_ /*48553*/;
assign _675_ = _676_ | _678_ /*48551*/;
assign _430_ = _670_ ^ _677_ /*48554*/;
assign _684_ = D[46] ^ Q[63] /*48550*/;
assign _681_ = _45_ & _684_ /*48546*/;
assign _682_ = _45_ ^ _684_ /*48549*/;
assign _683_ = _675_ & _682_ /*48547*/;
assign _680_ = _681_ | _683_ /*48545*/;
assign _431_ = _675_ ^ _682_ /*48548*/;
assign _689_ = D[47] ^ Q[63] /*48544*/;
assign _686_ = _46_ & _689_ /*48540*/;
assign _687_ = _46_ ^ _689_ /*48543*/;
assign _688_ = _680_ & _687_ /*48541*/;
assign _685_ = _686_ | _688_ /*48539*/;
assign _432_ = _680_ ^ _687_ /*48542*/;
assign _694_ = D[48] ^ Q[63] /*48538*/;
assign _691_ = _47_ & _694_ /*48534*/;
assign _692_ = _47_ ^ _694_ /*48537*/;
assign _693_ = _685_ & _692_ /*48535*/;
assign _690_ = _691_ | _693_ /*48533*/;
assign _433_ = _685_ ^ _692_ /*48536*/;
assign _699_ = D[49] ^ Q[63] /*48532*/;
assign _696_ = _48_ & _699_ /*48528*/;
assign _697_ = _48_ ^ _699_ /*48531*/;
assign _698_ = _690_ & _697_ /*48529*/;
assign _695_ = _696_ | _698_ /*48527*/;
assign _434_ = _690_ ^ _697_ /*48530*/;
assign _704_ = D[50] ^ Q[63] /*48526*/;
assign _701_ = _49_ & _704_ /*48522*/;
assign _702_ = _49_ ^ _704_ /*48525*/;
assign _703_ = _695_ & _702_ /*48523*/;
assign _700_ = _701_ | _703_ /*48521*/;
assign _435_ = _695_ ^ _702_ /*48524*/;
assign _709_ = D[51] ^ Q[63] /*48520*/;
assign _706_ = _50_ & _709_ /*48516*/;
assign _707_ = _50_ ^ _709_ /*48519*/;
assign _708_ = _700_ & _707_ /*48517*/;
assign _705_ = _706_ | _708_ /*48515*/;
assign _436_ = _700_ ^ _707_ /*48518*/;
assign _714_ = D[52] ^ Q[63] /*48514*/;
assign _711_ = _51_ & _714_ /*48510*/;
assign _712_ = _51_ ^ _714_ /*48513*/;
assign _713_ = _705_ & _712_ /*48511*/;
assign _710_ = _711_ | _713_ /*48509*/;
assign _437_ = _705_ ^ _712_ /*48512*/;
assign _719_ = D[53] ^ Q[63] /*48508*/;
assign _716_ = _52_ & _719_ /*48504*/;
assign _717_ = _52_ ^ _719_ /*48507*/;
assign _718_ = _710_ & _717_ /*48505*/;
assign _715_ = _716_ | _718_ /*48503*/;
assign _438_ = _710_ ^ _717_ /*48506*/;
assign _724_ = D[54] ^ Q[63] /*48502*/;
assign _721_ = _53_ & _724_ /*48498*/;
assign _722_ = _53_ ^ _724_ /*48501*/;
assign _723_ = _715_ & _722_ /*48499*/;
assign _720_ = _721_ | _723_ /*48497*/;
assign _439_ = _715_ ^ _722_ /*48500*/;
assign _729_ = D[55] ^ Q[63] /*48496*/;
assign _726_ = _54_ & _729_ /*48492*/;
assign _727_ = _54_ ^ _729_ /*48495*/;
assign _728_ = _720_ & _727_ /*48493*/;
assign _725_ = _726_ | _728_ /*48491*/;
assign _440_ = _720_ ^ _727_ /*48494*/;
assign _734_ = D[56] ^ Q[63] /*48490*/;
assign _731_ = _55_ & _734_ /*48486*/;
assign _732_ = _55_ ^ _734_ /*48489*/;
assign _733_ = _725_ & _732_ /*48487*/;
assign _730_ = _731_ | _733_ /*48485*/;
assign _441_ = _725_ ^ _732_ /*48488*/;
assign _739_ = D[57] ^ Q[63] /*48484*/;
assign _736_ = _56_ & _739_ /*48480*/;
assign _737_ = _56_ ^ _739_ /*48483*/;
assign _738_ = _730_ & _737_ /*48481*/;
assign _735_ = _736_ | _738_ /*48479*/;
assign _442_ = _730_ ^ _737_ /*48482*/;
assign _744_ = D[58] ^ Q[63] /*48478*/;
assign _741_ = _57_ & _744_ /*48474*/;
assign _742_ = _57_ ^ _744_ /*48477*/;
assign _743_ = _735_ & _742_ /*48475*/;
assign _740_ = _741_ | _743_ /*48473*/;
assign _443_ = _735_ ^ _742_ /*48476*/;
assign _749_ = D[59] ^ Q[63] /*48472*/;
assign _746_ = _58_ & _749_ /*48468*/;
assign _747_ = _58_ ^ _749_ /*48471*/;
assign _748_ = _740_ & _747_ /*48469*/;
assign _745_ = _746_ | _748_ /*48467*/;
assign _444_ = _740_ ^ _747_ /*48470*/;
assign _754_ = D[60] ^ Q[63] /*48466*/;
assign _751_ = _59_ & _754_ /*48462*/;
assign _752_ = _59_ ^ _754_ /*48465*/;
assign _753_ = _745_ & _752_ /*48463*/;
assign _750_ = _751_ | _753_ /*48461*/;
assign _445_ = _745_ ^ _752_ /*48464*/;
assign _759_ = D[61] ^ Q[63] /*48460*/;
assign _756_ = _60_ & _759_ /*48456*/;
assign _757_ = _60_ ^ _759_ /*48459*/;
assign _758_ = _750_ & _757_ /*48457*/;
assign _755_ = _756_ | _758_ /*48455*/;
assign _446_ = _750_ ^ _757_ /*48458*/;
assign _764_ = D[62] ^ Q[63] /*48454*/;
assign _761_ = _61_ & _764_ /*48450*/;
assign _762_ = _61_ ^ _764_ /*48453*/;
assign _763_ = _755_ & _762_ /*48451*/;
assign _760_ = _761_ | _763_ /*48449*/;
assign _447_ = _755_ ^ _762_ /*48452*/;
assign _768_ = zeroWire ^ Q[63] /*48448*/;
assign _765_ = _62_ & _768_ /*48444*/;
assign _766_ = _62_ ^ _768_ /*48447*/;
assign _767_ = _760_ & _766_ /*48445*/;
assign Q[62] = _765_ | _767_ /*48443*/;
assign _448_ = _760_ ^ _766_ /*48446*/;
assign _839_ = D[0] ^ Q[62] /*48057*/;
assign _836_ = R_0[61] & _839_ /*48053*/;
assign _837_ = R_0[61] ^ _839_ /*48056*/;
assign _838_ = Q[62] & _837_ /*48054*/;
assign _835_ = _836_ | _838_ /*48052*/;
assign _770_ = Q[62] ^ _837_ /*48055*/;
assign _844_ = D[1] ^ Q[62] /*48051*/;
assign _841_ = _385_ & _844_ /*48047*/;
assign _842_ = _385_ ^ _844_ /*48050*/;
assign _843_ = _835_ & _842_ /*48048*/;
assign _840_ = _841_ | _843_ /*48046*/;
assign _771_ = _835_ ^ _842_ /*48049*/;
assign _849_ = D[2] ^ Q[62] /*48045*/;
assign _846_ = _386_ & _849_ /*48041*/;
assign _847_ = _386_ ^ _849_ /*48044*/;
assign _848_ = _840_ & _847_ /*48042*/;
assign _845_ = _846_ | _848_ /*48040*/;
assign _772_ = _840_ ^ _847_ /*48043*/;
assign _854_ = D[3] ^ Q[62] /*48039*/;
assign _851_ = _387_ & _854_ /*48035*/;
assign _852_ = _387_ ^ _854_ /*48038*/;
assign _853_ = _845_ & _852_ /*48036*/;
assign _850_ = _851_ | _853_ /*48034*/;
assign _773_ = _845_ ^ _852_ /*48037*/;
assign _859_ = D[4] ^ Q[62] /*48033*/;
assign _856_ = _388_ & _859_ /*48029*/;
assign _857_ = _388_ ^ _859_ /*48032*/;
assign _858_ = _850_ & _857_ /*48030*/;
assign _855_ = _856_ | _858_ /*48028*/;
assign _774_ = _850_ ^ _857_ /*48031*/;
assign _864_ = D[5] ^ Q[62] /*48027*/;
assign _861_ = _389_ & _864_ /*48023*/;
assign _862_ = _389_ ^ _864_ /*48026*/;
assign _863_ = _855_ & _862_ /*48024*/;
assign _860_ = _861_ | _863_ /*48022*/;
assign _775_ = _855_ ^ _862_ /*48025*/;
assign _869_ = D[6] ^ Q[62] /*48021*/;
assign _866_ = _390_ & _869_ /*48017*/;
assign _867_ = _390_ ^ _869_ /*48020*/;
assign _868_ = _860_ & _867_ /*48018*/;
assign _865_ = _866_ | _868_ /*48016*/;
assign _776_ = _860_ ^ _867_ /*48019*/;
assign _874_ = D[7] ^ Q[62] /*48015*/;
assign _871_ = _391_ & _874_ /*48011*/;
assign _872_ = _391_ ^ _874_ /*48014*/;
assign _873_ = _865_ & _872_ /*48012*/;
assign _870_ = _871_ | _873_ /*48010*/;
assign _777_ = _865_ ^ _872_ /*48013*/;
assign _879_ = D[8] ^ Q[62] /*48009*/;
assign _876_ = _392_ & _879_ /*48005*/;
assign _877_ = _392_ ^ _879_ /*48008*/;
assign _878_ = _870_ & _877_ /*48006*/;
assign _875_ = _876_ | _878_ /*48004*/;
assign _778_ = _870_ ^ _877_ /*48007*/;
assign _884_ = D[9] ^ Q[62] /*48003*/;
assign _881_ = _393_ & _884_ /*47999*/;
assign _882_ = _393_ ^ _884_ /*48002*/;
assign _883_ = _875_ & _882_ /*48000*/;
assign _880_ = _881_ | _883_ /*47998*/;
assign _779_ = _875_ ^ _882_ /*48001*/;
assign _889_ = D[10] ^ Q[62] /*47997*/;
assign _886_ = _394_ & _889_ /*47993*/;
assign _887_ = _394_ ^ _889_ /*47996*/;
assign _888_ = _880_ & _887_ /*47994*/;
assign _885_ = _886_ | _888_ /*47992*/;
assign _780_ = _880_ ^ _887_ /*47995*/;
assign _894_ = D[11] ^ Q[62] /*47991*/;
assign _891_ = _395_ & _894_ /*47987*/;
assign _892_ = _395_ ^ _894_ /*47990*/;
assign _893_ = _885_ & _892_ /*47988*/;
assign _890_ = _891_ | _893_ /*47986*/;
assign _781_ = _885_ ^ _892_ /*47989*/;
assign _899_ = D[12] ^ Q[62] /*47985*/;
assign _896_ = _396_ & _899_ /*47981*/;
assign _897_ = _396_ ^ _899_ /*47984*/;
assign _898_ = _890_ & _897_ /*47982*/;
assign _895_ = _896_ | _898_ /*47980*/;
assign _782_ = _890_ ^ _897_ /*47983*/;
assign _904_ = D[13] ^ Q[62] /*47979*/;
assign _901_ = _397_ & _904_ /*47975*/;
assign _902_ = _397_ ^ _904_ /*47978*/;
assign _903_ = _895_ & _902_ /*47976*/;
assign _900_ = _901_ | _903_ /*47974*/;
assign _783_ = _895_ ^ _902_ /*47977*/;
assign _909_ = D[14] ^ Q[62] /*47973*/;
assign _906_ = _398_ & _909_ /*47969*/;
assign _907_ = _398_ ^ _909_ /*47972*/;
assign _908_ = _900_ & _907_ /*47970*/;
assign _905_ = _906_ | _908_ /*47968*/;
assign _784_ = _900_ ^ _907_ /*47971*/;
assign _914_ = D[15] ^ Q[62] /*47967*/;
assign _911_ = _399_ & _914_ /*47963*/;
assign _912_ = _399_ ^ _914_ /*47966*/;
assign _913_ = _905_ & _912_ /*47964*/;
assign _910_ = _911_ | _913_ /*47962*/;
assign _785_ = _905_ ^ _912_ /*47965*/;
assign _919_ = D[16] ^ Q[62] /*47961*/;
assign _916_ = _400_ & _919_ /*47957*/;
assign _917_ = _400_ ^ _919_ /*47960*/;
assign _918_ = _910_ & _917_ /*47958*/;
assign _915_ = _916_ | _918_ /*47956*/;
assign _786_ = _910_ ^ _917_ /*47959*/;
assign _924_ = D[17] ^ Q[62] /*47955*/;
assign _921_ = _401_ & _924_ /*47951*/;
assign _922_ = _401_ ^ _924_ /*47954*/;
assign _923_ = _915_ & _922_ /*47952*/;
assign _920_ = _921_ | _923_ /*47950*/;
assign _787_ = _915_ ^ _922_ /*47953*/;
assign _929_ = D[18] ^ Q[62] /*47949*/;
assign _926_ = _402_ & _929_ /*47945*/;
assign _927_ = _402_ ^ _929_ /*47948*/;
assign _928_ = _920_ & _927_ /*47946*/;
assign _925_ = _926_ | _928_ /*47944*/;
assign _788_ = _920_ ^ _927_ /*47947*/;
assign _934_ = D[19] ^ Q[62] /*47943*/;
assign _931_ = _403_ & _934_ /*47939*/;
assign _932_ = _403_ ^ _934_ /*47942*/;
assign _933_ = _925_ & _932_ /*47940*/;
assign _930_ = _931_ | _933_ /*47938*/;
assign _789_ = _925_ ^ _932_ /*47941*/;
assign _939_ = D[20] ^ Q[62] /*47937*/;
assign _936_ = _404_ & _939_ /*47933*/;
assign _937_ = _404_ ^ _939_ /*47936*/;
assign _938_ = _930_ & _937_ /*47934*/;
assign _935_ = _936_ | _938_ /*47932*/;
assign _790_ = _930_ ^ _937_ /*47935*/;
assign _944_ = D[21] ^ Q[62] /*47931*/;
assign _941_ = _405_ & _944_ /*47927*/;
assign _942_ = _405_ ^ _944_ /*47930*/;
assign _943_ = _935_ & _942_ /*47928*/;
assign _940_ = _941_ | _943_ /*47926*/;
assign _791_ = _935_ ^ _942_ /*47929*/;
assign _949_ = D[22] ^ Q[62] /*47925*/;
assign _946_ = _406_ & _949_ /*47921*/;
assign _947_ = _406_ ^ _949_ /*47924*/;
assign _948_ = _940_ & _947_ /*47922*/;
assign _945_ = _946_ | _948_ /*47920*/;
assign _792_ = _940_ ^ _947_ /*47923*/;
assign _954_ = D[23] ^ Q[62] /*47919*/;
assign _951_ = _407_ & _954_ /*47915*/;
assign _952_ = _407_ ^ _954_ /*47918*/;
assign _953_ = _945_ & _952_ /*47916*/;
assign _950_ = _951_ | _953_ /*47914*/;
assign _793_ = _945_ ^ _952_ /*47917*/;
assign _959_ = D[24] ^ Q[62] /*47913*/;
assign _956_ = _408_ & _959_ /*47909*/;
assign _957_ = _408_ ^ _959_ /*47912*/;
assign _958_ = _950_ & _957_ /*47910*/;
assign _955_ = _956_ | _958_ /*47908*/;
assign _794_ = _950_ ^ _957_ /*47911*/;
assign _964_ = D[25] ^ Q[62] /*47907*/;
assign _961_ = _409_ & _964_ /*47903*/;
assign _962_ = _409_ ^ _964_ /*47906*/;
assign _963_ = _955_ & _962_ /*47904*/;
assign _960_ = _961_ | _963_ /*47902*/;
assign _795_ = _955_ ^ _962_ /*47905*/;
assign _969_ = D[26] ^ Q[62] /*47901*/;
assign _966_ = _410_ & _969_ /*47897*/;
assign _967_ = _410_ ^ _969_ /*47900*/;
assign _968_ = _960_ & _967_ /*47898*/;
assign _965_ = _966_ | _968_ /*47896*/;
assign _796_ = _960_ ^ _967_ /*47899*/;
assign _974_ = D[27] ^ Q[62] /*47895*/;
assign _971_ = _411_ & _974_ /*47891*/;
assign _972_ = _411_ ^ _974_ /*47894*/;
assign _973_ = _965_ & _972_ /*47892*/;
assign _970_ = _971_ | _973_ /*47890*/;
assign _797_ = _965_ ^ _972_ /*47893*/;
assign _979_ = D[28] ^ Q[62] /*47889*/;
assign _976_ = _412_ & _979_ /*47885*/;
assign _977_ = _412_ ^ _979_ /*47888*/;
assign _978_ = _970_ & _977_ /*47886*/;
assign _975_ = _976_ | _978_ /*47884*/;
assign _798_ = _970_ ^ _977_ /*47887*/;
assign _984_ = D[29] ^ Q[62] /*47883*/;
assign _981_ = _413_ & _984_ /*47879*/;
assign _982_ = _413_ ^ _984_ /*47882*/;
assign _983_ = _975_ & _982_ /*47880*/;
assign _980_ = _981_ | _983_ /*47878*/;
assign _799_ = _975_ ^ _982_ /*47881*/;
assign _989_ = D[30] ^ Q[62] /*47877*/;
assign _986_ = _414_ & _989_ /*47873*/;
assign _987_ = _414_ ^ _989_ /*47876*/;
assign _988_ = _980_ & _987_ /*47874*/;
assign _985_ = _986_ | _988_ /*47872*/;
assign _800_ = _980_ ^ _987_ /*47875*/;
assign _994_ = D[31] ^ Q[62] /*47871*/;
assign _991_ = _415_ & _994_ /*47867*/;
assign _992_ = _415_ ^ _994_ /*47870*/;
assign _993_ = _985_ & _992_ /*47868*/;
assign _990_ = _991_ | _993_ /*47866*/;
assign _801_ = _985_ ^ _992_ /*47869*/;
assign _999_ = D[32] ^ Q[62] /*47865*/;
assign _996_ = _416_ & _999_ /*47861*/;
assign _997_ = _416_ ^ _999_ /*47864*/;
assign _998_ = _990_ & _997_ /*47862*/;
assign _995_ = _996_ | _998_ /*47860*/;
assign _802_ = _990_ ^ _997_ /*47863*/;
assign _1004_ = D[33] ^ Q[62] /*47859*/;
assign _1001_ = _417_ & _1004_ /*47855*/;
assign _1002_ = _417_ ^ _1004_ /*47858*/;
assign _1003_ = _995_ & _1002_ /*47856*/;
assign _1000_ = _1001_ | _1003_ /*47854*/;
assign _803_ = _995_ ^ _1002_ /*47857*/;
assign _1009_ = D[34] ^ Q[62] /*47853*/;
assign _1006_ = _418_ & _1009_ /*47849*/;
assign _1007_ = _418_ ^ _1009_ /*47852*/;
assign _1008_ = _1000_ & _1007_ /*47850*/;
assign _1005_ = _1006_ | _1008_ /*47848*/;
assign _804_ = _1000_ ^ _1007_ /*47851*/;
assign _1014_ = D[35] ^ Q[62] /*47847*/;
assign _1011_ = _419_ & _1014_ /*47843*/;
assign _1012_ = _419_ ^ _1014_ /*47846*/;
assign _1013_ = _1005_ & _1012_ /*47844*/;
assign _1010_ = _1011_ | _1013_ /*47842*/;
assign _805_ = _1005_ ^ _1012_ /*47845*/;
assign _1019_ = D[36] ^ Q[62] /*47841*/;
assign _1016_ = _420_ & _1019_ /*47837*/;
assign _1017_ = _420_ ^ _1019_ /*47840*/;
assign _1018_ = _1010_ & _1017_ /*47838*/;
assign _1015_ = _1016_ | _1018_ /*47836*/;
assign _806_ = _1010_ ^ _1017_ /*47839*/;
assign _1024_ = D[37] ^ Q[62] /*47835*/;
assign _1021_ = _421_ & _1024_ /*47831*/;
assign _1022_ = _421_ ^ _1024_ /*47834*/;
assign _1023_ = _1015_ & _1022_ /*47832*/;
assign _1020_ = _1021_ | _1023_ /*47830*/;
assign _807_ = _1015_ ^ _1022_ /*47833*/;
assign _1029_ = D[38] ^ Q[62] /*47829*/;
assign _1026_ = _422_ & _1029_ /*47825*/;
assign _1027_ = _422_ ^ _1029_ /*47828*/;
assign _1028_ = _1020_ & _1027_ /*47826*/;
assign _1025_ = _1026_ | _1028_ /*47824*/;
assign _808_ = _1020_ ^ _1027_ /*47827*/;
assign _1034_ = D[39] ^ Q[62] /*47823*/;
assign _1031_ = _423_ & _1034_ /*47819*/;
assign _1032_ = _423_ ^ _1034_ /*47822*/;
assign _1033_ = _1025_ & _1032_ /*47820*/;
assign _1030_ = _1031_ | _1033_ /*47818*/;
assign _809_ = _1025_ ^ _1032_ /*47821*/;
assign _1039_ = D[40] ^ Q[62] /*47817*/;
assign _1036_ = _424_ & _1039_ /*47813*/;
assign _1037_ = _424_ ^ _1039_ /*47816*/;
assign _1038_ = _1030_ & _1037_ /*47814*/;
assign _1035_ = _1036_ | _1038_ /*47812*/;
assign _810_ = _1030_ ^ _1037_ /*47815*/;
assign _1044_ = D[41] ^ Q[62] /*47811*/;
assign _1041_ = _425_ & _1044_ /*47807*/;
assign _1042_ = _425_ ^ _1044_ /*47810*/;
assign _1043_ = _1035_ & _1042_ /*47808*/;
assign _1040_ = _1041_ | _1043_ /*47806*/;
assign _811_ = _1035_ ^ _1042_ /*47809*/;
assign _1049_ = D[42] ^ Q[62] /*47805*/;
assign _1046_ = _426_ & _1049_ /*47801*/;
assign _1047_ = _426_ ^ _1049_ /*47804*/;
assign _1048_ = _1040_ & _1047_ /*47802*/;
assign _1045_ = _1046_ | _1048_ /*47800*/;
assign _812_ = _1040_ ^ _1047_ /*47803*/;
assign _1054_ = D[43] ^ Q[62] /*47799*/;
assign _1051_ = _427_ & _1054_ /*47795*/;
assign _1052_ = _427_ ^ _1054_ /*47798*/;
assign _1053_ = _1045_ & _1052_ /*47796*/;
assign _1050_ = _1051_ | _1053_ /*47794*/;
assign _813_ = _1045_ ^ _1052_ /*47797*/;
assign _1059_ = D[44] ^ Q[62] /*47793*/;
assign _1056_ = _428_ & _1059_ /*47789*/;
assign _1057_ = _428_ ^ _1059_ /*47792*/;
assign _1058_ = _1050_ & _1057_ /*47790*/;
assign _1055_ = _1056_ | _1058_ /*47788*/;
assign _814_ = _1050_ ^ _1057_ /*47791*/;
assign _1064_ = D[45] ^ Q[62] /*47787*/;
assign _1061_ = _429_ & _1064_ /*47783*/;
assign _1062_ = _429_ ^ _1064_ /*47786*/;
assign _1063_ = _1055_ & _1062_ /*47784*/;
assign _1060_ = _1061_ | _1063_ /*47782*/;
assign _815_ = _1055_ ^ _1062_ /*47785*/;
assign _1069_ = D[46] ^ Q[62] /*47781*/;
assign _1066_ = _430_ & _1069_ /*47777*/;
assign _1067_ = _430_ ^ _1069_ /*47780*/;
assign _1068_ = _1060_ & _1067_ /*47778*/;
assign _1065_ = _1066_ | _1068_ /*47776*/;
assign _816_ = _1060_ ^ _1067_ /*47779*/;
assign _1074_ = D[47] ^ Q[62] /*47775*/;
assign _1071_ = _431_ & _1074_ /*47771*/;
assign _1072_ = _431_ ^ _1074_ /*47774*/;
assign _1073_ = _1065_ & _1072_ /*47772*/;
assign _1070_ = _1071_ | _1073_ /*47770*/;
assign _817_ = _1065_ ^ _1072_ /*47773*/;
assign _1079_ = D[48] ^ Q[62] /*47769*/;
assign _1076_ = _432_ & _1079_ /*47765*/;
assign _1077_ = _432_ ^ _1079_ /*47768*/;
assign _1078_ = _1070_ & _1077_ /*47766*/;
assign _1075_ = _1076_ | _1078_ /*47764*/;
assign _818_ = _1070_ ^ _1077_ /*47767*/;
assign _1084_ = D[49] ^ Q[62] /*47763*/;
assign _1081_ = _433_ & _1084_ /*47759*/;
assign _1082_ = _433_ ^ _1084_ /*47762*/;
assign _1083_ = _1075_ & _1082_ /*47760*/;
assign _1080_ = _1081_ | _1083_ /*47758*/;
assign _819_ = _1075_ ^ _1082_ /*47761*/;
assign _1089_ = D[50] ^ Q[62] /*47757*/;
assign _1086_ = _434_ & _1089_ /*47753*/;
assign _1087_ = _434_ ^ _1089_ /*47756*/;
assign _1088_ = _1080_ & _1087_ /*47754*/;
assign _1085_ = _1086_ | _1088_ /*47752*/;
assign _820_ = _1080_ ^ _1087_ /*47755*/;
assign _1094_ = D[51] ^ Q[62] /*47751*/;
assign _1091_ = _435_ & _1094_ /*47747*/;
assign _1092_ = _435_ ^ _1094_ /*47750*/;
assign _1093_ = _1085_ & _1092_ /*47748*/;
assign _1090_ = _1091_ | _1093_ /*47746*/;
assign _821_ = _1085_ ^ _1092_ /*47749*/;
assign _1099_ = D[52] ^ Q[62] /*47745*/;
assign _1096_ = _436_ & _1099_ /*47741*/;
assign _1097_ = _436_ ^ _1099_ /*47744*/;
assign _1098_ = _1090_ & _1097_ /*47742*/;
assign _1095_ = _1096_ | _1098_ /*47740*/;
assign _822_ = _1090_ ^ _1097_ /*47743*/;
assign _1104_ = D[53] ^ Q[62] /*47739*/;
assign _1101_ = _437_ & _1104_ /*47735*/;
assign _1102_ = _437_ ^ _1104_ /*47738*/;
assign _1103_ = _1095_ & _1102_ /*47736*/;
assign _1100_ = _1101_ | _1103_ /*47734*/;
assign _823_ = _1095_ ^ _1102_ /*47737*/;
assign _1109_ = D[54] ^ Q[62] /*47733*/;
assign _1106_ = _438_ & _1109_ /*47729*/;
assign _1107_ = _438_ ^ _1109_ /*47732*/;
assign _1108_ = _1100_ & _1107_ /*47730*/;
assign _1105_ = _1106_ | _1108_ /*47728*/;
assign _824_ = _1100_ ^ _1107_ /*47731*/;
assign _1114_ = D[55] ^ Q[62] /*47727*/;
assign _1111_ = _439_ & _1114_ /*47723*/;
assign _1112_ = _439_ ^ _1114_ /*47726*/;
assign _1113_ = _1105_ & _1112_ /*47724*/;
assign _1110_ = _1111_ | _1113_ /*47722*/;
assign _825_ = _1105_ ^ _1112_ /*47725*/;
assign _1119_ = D[56] ^ Q[62] /*47721*/;
assign _1116_ = _440_ & _1119_ /*47717*/;
assign _1117_ = _440_ ^ _1119_ /*47720*/;
assign _1118_ = _1110_ & _1117_ /*47718*/;
assign _1115_ = _1116_ | _1118_ /*47716*/;
assign _826_ = _1110_ ^ _1117_ /*47719*/;
assign _1124_ = D[57] ^ Q[62] /*47715*/;
assign _1121_ = _441_ & _1124_ /*47711*/;
assign _1122_ = _441_ ^ _1124_ /*47714*/;
assign _1123_ = _1115_ & _1122_ /*47712*/;
assign _1120_ = _1121_ | _1123_ /*47710*/;
assign _827_ = _1115_ ^ _1122_ /*47713*/;
assign _1129_ = D[58] ^ Q[62] /*47709*/;
assign _1126_ = _442_ & _1129_ /*47705*/;
assign _1127_ = _442_ ^ _1129_ /*47708*/;
assign _1128_ = _1120_ & _1127_ /*47706*/;
assign _1125_ = _1126_ | _1128_ /*47704*/;
assign _828_ = _1120_ ^ _1127_ /*47707*/;
assign _1134_ = D[59] ^ Q[62] /*47703*/;
assign _1131_ = _443_ & _1134_ /*47699*/;
assign _1132_ = _443_ ^ _1134_ /*47702*/;
assign _1133_ = _1125_ & _1132_ /*47700*/;
assign _1130_ = _1131_ | _1133_ /*47698*/;
assign _829_ = _1125_ ^ _1132_ /*47701*/;
assign _1139_ = D[60] ^ Q[62] /*47697*/;
assign _1136_ = _444_ & _1139_ /*47693*/;
assign _1137_ = _444_ ^ _1139_ /*47696*/;
assign _1138_ = _1130_ & _1137_ /*47694*/;
assign _1135_ = _1136_ | _1138_ /*47692*/;
assign _830_ = _1130_ ^ _1137_ /*47695*/;
assign _1144_ = D[61] ^ Q[62] /*47691*/;
assign _1141_ = _445_ & _1144_ /*47687*/;
assign _1142_ = _445_ ^ _1144_ /*47690*/;
assign _1143_ = _1135_ & _1142_ /*47688*/;
assign _1140_ = _1141_ | _1143_ /*47686*/;
assign _831_ = _1135_ ^ _1142_ /*47689*/;
assign _1149_ = D[62] ^ Q[62] /*47685*/;
assign _1146_ = _446_ & _1149_ /*47681*/;
assign _1147_ = _446_ ^ _1149_ /*47684*/;
assign _1148_ = _1140_ & _1147_ /*47682*/;
assign _1145_ = _1146_ | _1148_ /*47680*/;
assign _832_ = _1140_ ^ _1147_ /*47683*/;
assign _1153_ = zeroWire ^ Q[62] /*47679*/;
assign _1150_ = _447_ & _1153_ /*47675*/;
assign _1151_ = _447_ ^ _1153_ /*47678*/;
assign _1152_ = _1145_ & _1151_ /*47676*/;
assign Q[61] = _1150_ | _1152_ /*47674*/;
assign _833_ = _1145_ ^ _1151_ /*47677*/;
assign _1224_ = D[0] ^ Q[61] /*47288*/;
assign _1221_ = R_0[60] & _1224_ /*47284*/;
assign _1222_ = R_0[60] ^ _1224_ /*47287*/;
assign _1223_ = Q[61] & _1222_ /*47285*/;
assign _1220_ = _1221_ | _1223_ /*47283*/;
assign _1155_ = Q[61] ^ _1222_ /*47286*/;
assign _1229_ = D[1] ^ Q[61] /*47282*/;
assign _1226_ = _770_ & _1229_ /*47278*/;
assign _1227_ = _770_ ^ _1229_ /*47281*/;
assign _1228_ = _1220_ & _1227_ /*47279*/;
assign _1225_ = _1226_ | _1228_ /*47277*/;
assign _1156_ = _1220_ ^ _1227_ /*47280*/;
assign _1234_ = D[2] ^ Q[61] /*47276*/;
assign _1231_ = _771_ & _1234_ /*47272*/;
assign _1232_ = _771_ ^ _1234_ /*47275*/;
assign _1233_ = _1225_ & _1232_ /*47273*/;
assign _1230_ = _1231_ | _1233_ /*47271*/;
assign _1157_ = _1225_ ^ _1232_ /*47274*/;
assign _1239_ = D[3] ^ Q[61] /*47270*/;
assign _1236_ = _772_ & _1239_ /*47266*/;
assign _1237_ = _772_ ^ _1239_ /*47269*/;
assign _1238_ = _1230_ & _1237_ /*47267*/;
assign _1235_ = _1236_ | _1238_ /*47265*/;
assign _1158_ = _1230_ ^ _1237_ /*47268*/;
assign _1244_ = D[4] ^ Q[61] /*47264*/;
assign _1241_ = _773_ & _1244_ /*47260*/;
assign _1242_ = _773_ ^ _1244_ /*47263*/;
assign _1243_ = _1235_ & _1242_ /*47261*/;
assign _1240_ = _1241_ | _1243_ /*47259*/;
assign _1159_ = _1235_ ^ _1242_ /*47262*/;
assign _1249_ = D[5] ^ Q[61] /*47258*/;
assign _1246_ = _774_ & _1249_ /*47254*/;
assign _1247_ = _774_ ^ _1249_ /*47257*/;
assign _1248_ = _1240_ & _1247_ /*47255*/;
assign _1245_ = _1246_ | _1248_ /*47253*/;
assign _1160_ = _1240_ ^ _1247_ /*47256*/;
assign _1254_ = D[6] ^ Q[61] /*47252*/;
assign _1251_ = _775_ & _1254_ /*47248*/;
assign _1252_ = _775_ ^ _1254_ /*47251*/;
assign _1253_ = _1245_ & _1252_ /*47249*/;
assign _1250_ = _1251_ | _1253_ /*47247*/;
assign _1161_ = _1245_ ^ _1252_ /*47250*/;
assign _1259_ = D[7] ^ Q[61] /*47246*/;
assign _1256_ = _776_ & _1259_ /*47242*/;
assign _1257_ = _776_ ^ _1259_ /*47245*/;
assign _1258_ = _1250_ & _1257_ /*47243*/;
assign _1255_ = _1256_ | _1258_ /*47241*/;
assign _1162_ = _1250_ ^ _1257_ /*47244*/;
assign _1264_ = D[8] ^ Q[61] /*47240*/;
assign _1261_ = _777_ & _1264_ /*47236*/;
assign _1262_ = _777_ ^ _1264_ /*47239*/;
assign _1263_ = _1255_ & _1262_ /*47237*/;
assign _1260_ = _1261_ | _1263_ /*47235*/;
assign _1163_ = _1255_ ^ _1262_ /*47238*/;
assign _1269_ = D[9] ^ Q[61] /*47234*/;
assign _1266_ = _778_ & _1269_ /*47230*/;
assign _1267_ = _778_ ^ _1269_ /*47233*/;
assign _1268_ = _1260_ & _1267_ /*47231*/;
assign _1265_ = _1266_ | _1268_ /*47229*/;
assign _1164_ = _1260_ ^ _1267_ /*47232*/;
assign _1274_ = D[10] ^ Q[61] /*47228*/;
assign _1271_ = _779_ & _1274_ /*47224*/;
assign _1272_ = _779_ ^ _1274_ /*47227*/;
assign _1273_ = _1265_ & _1272_ /*47225*/;
assign _1270_ = _1271_ | _1273_ /*47223*/;
assign _1165_ = _1265_ ^ _1272_ /*47226*/;
assign _1279_ = D[11] ^ Q[61] /*47222*/;
assign _1276_ = _780_ & _1279_ /*47218*/;
assign _1277_ = _780_ ^ _1279_ /*47221*/;
assign _1278_ = _1270_ & _1277_ /*47219*/;
assign _1275_ = _1276_ | _1278_ /*47217*/;
assign _1166_ = _1270_ ^ _1277_ /*47220*/;
assign _1284_ = D[12] ^ Q[61] /*47216*/;
assign _1281_ = _781_ & _1284_ /*47212*/;
assign _1282_ = _781_ ^ _1284_ /*47215*/;
assign _1283_ = _1275_ & _1282_ /*47213*/;
assign _1280_ = _1281_ | _1283_ /*47211*/;
assign _1167_ = _1275_ ^ _1282_ /*47214*/;
assign _1289_ = D[13] ^ Q[61] /*47210*/;
assign _1286_ = _782_ & _1289_ /*47206*/;
assign _1287_ = _782_ ^ _1289_ /*47209*/;
assign _1288_ = _1280_ & _1287_ /*47207*/;
assign _1285_ = _1286_ | _1288_ /*47205*/;
assign _1168_ = _1280_ ^ _1287_ /*47208*/;
assign _1294_ = D[14] ^ Q[61] /*47204*/;
assign _1291_ = _783_ & _1294_ /*47200*/;
assign _1292_ = _783_ ^ _1294_ /*47203*/;
assign _1293_ = _1285_ & _1292_ /*47201*/;
assign _1290_ = _1291_ | _1293_ /*47199*/;
assign _1169_ = _1285_ ^ _1292_ /*47202*/;
assign _1299_ = D[15] ^ Q[61] /*47198*/;
assign _1296_ = _784_ & _1299_ /*47194*/;
assign _1297_ = _784_ ^ _1299_ /*47197*/;
assign _1298_ = _1290_ & _1297_ /*47195*/;
assign _1295_ = _1296_ | _1298_ /*47193*/;
assign _1170_ = _1290_ ^ _1297_ /*47196*/;
assign _1304_ = D[16] ^ Q[61] /*47192*/;
assign _1301_ = _785_ & _1304_ /*47188*/;
assign _1302_ = _785_ ^ _1304_ /*47191*/;
assign _1303_ = _1295_ & _1302_ /*47189*/;
assign _1300_ = _1301_ | _1303_ /*47187*/;
assign _1171_ = _1295_ ^ _1302_ /*47190*/;
assign _1309_ = D[17] ^ Q[61] /*47186*/;
assign _1306_ = _786_ & _1309_ /*47182*/;
assign _1307_ = _786_ ^ _1309_ /*47185*/;
assign _1308_ = _1300_ & _1307_ /*47183*/;
assign _1305_ = _1306_ | _1308_ /*47181*/;
assign _1172_ = _1300_ ^ _1307_ /*47184*/;
assign _1314_ = D[18] ^ Q[61] /*47180*/;
assign _1311_ = _787_ & _1314_ /*47176*/;
assign _1312_ = _787_ ^ _1314_ /*47179*/;
assign _1313_ = _1305_ & _1312_ /*47177*/;
assign _1310_ = _1311_ | _1313_ /*47175*/;
assign _1173_ = _1305_ ^ _1312_ /*47178*/;
assign _1319_ = D[19] ^ Q[61] /*47174*/;
assign _1316_ = _788_ & _1319_ /*47170*/;
assign _1317_ = _788_ ^ _1319_ /*47173*/;
assign _1318_ = _1310_ & _1317_ /*47171*/;
assign _1315_ = _1316_ | _1318_ /*47169*/;
assign _1174_ = _1310_ ^ _1317_ /*47172*/;
assign _1324_ = D[20] ^ Q[61] /*47168*/;
assign _1321_ = _789_ & _1324_ /*47164*/;
assign _1322_ = _789_ ^ _1324_ /*47167*/;
assign _1323_ = _1315_ & _1322_ /*47165*/;
assign _1320_ = _1321_ | _1323_ /*47163*/;
assign _1175_ = _1315_ ^ _1322_ /*47166*/;
assign _1329_ = D[21] ^ Q[61] /*47162*/;
assign _1326_ = _790_ & _1329_ /*47158*/;
assign _1327_ = _790_ ^ _1329_ /*47161*/;
assign _1328_ = _1320_ & _1327_ /*47159*/;
assign _1325_ = _1326_ | _1328_ /*47157*/;
assign _1176_ = _1320_ ^ _1327_ /*47160*/;
assign _1334_ = D[22] ^ Q[61] /*47156*/;
assign _1331_ = _791_ & _1334_ /*47152*/;
assign _1332_ = _791_ ^ _1334_ /*47155*/;
assign _1333_ = _1325_ & _1332_ /*47153*/;
assign _1330_ = _1331_ | _1333_ /*47151*/;
assign _1177_ = _1325_ ^ _1332_ /*47154*/;
assign _1339_ = D[23] ^ Q[61] /*47150*/;
assign _1336_ = _792_ & _1339_ /*47146*/;
assign _1337_ = _792_ ^ _1339_ /*47149*/;
assign _1338_ = _1330_ & _1337_ /*47147*/;
assign _1335_ = _1336_ | _1338_ /*47145*/;
assign _1178_ = _1330_ ^ _1337_ /*47148*/;
assign _1344_ = D[24] ^ Q[61] /*47144*/;
assign _1341_ = _793_ & _1344_ /*47140*/;
assign _1342_ = _793_ ^ _1344_ /*47143*/;
assign _1343_ = _1335_ & _1342_ /*47141*/;
assign _1340_ = _1341_ | _1343_ /*47139*/;
assign _1179_ = _1335_ ^ _1342_ /*47142*/;
assign _1349_ = D[25] ^ Q[61] /*47138*/;
assign _1346_ = _794_ & _1349_ /*47134*/;
assign _1347_ = _794_ ^ _1349_ /*47137*/;
assign _1348_ = _1340_ & _1347_ /*47135*/;
assign _1345_ = _1346_ | _1348_ /*47133*/;
assign _1180_ = _1340_ ^ _1347_ /*47136*/;
assign _1354_ = D[26] ^ Q[61] /*47132*/;
assign _1351_ = _795_ & _1354_ /*47128*/;
assign _1352_ = _795_ ^ _1354_ /*47131*/;
assign _1353_ = _1345_ & _1352_ /*47129*/;
assign _1350_ = _1351_ | _1353_ /*47127*/;
assign _1181_ = _1345_ ^ _1352_ /*47130*/;
assign _1359_ = D[27] ^ Q[61] /*47126*/;
assign _1356_ = _796_ & _1359_ /*47122*/;
assign _1357_ = _796_ ^ _1359_ /*47125*/;
assign _1358_ = _1350_ & _1357_ /*47123*/;
assign _1355_ = _1356_ | _1358_ /*47121*/;
assign _1182_ = _1350_ ^ _1357_ /*47124*/;
assign _1364_ = D[28] ^ Q[61] /*47120*/;
assign _1361_ = _797_ & _1364_ /*47116*/;
assign _1362_ = _797_ ^ _1364_ /*47119*/;
assign _1363_ = _1355_ & _1362_ /*47117*/;
assign _1360_ = _1361_ | _1363_ /*47115*/;
assign _1183_ = _1355_ ^ _1362_ /*47118*/;
assign _1369_ = D[29] ^ Q[61] /*47114*/;
assign _1366_ = _798_ & _1369_ /*47110*/;
assign _1367_ = _798_ ^ _1369_ /*47113*/;
assign _1368_ = _1360_ & _1367_ /*47111*/;
assign _1365_ = _1366_ | _1368_ /*47109*/;
assign _1184_ = _1360_ ^ _1367_ /*47112*/;
assign _1374_ = D[30] ^ Q[61] /*47108*/;
assign _1371_ = _799_ & _1374_ /*47104*/;
assign _1372_ = _799_ ^ _1374_ /*47107*/;
assign _1373_ = _1365_ & _1372_ /*47105*/;
assign _1370_ = _1371_ | _1373_ /*47103*/;
assign _1185_ = _1365_ ^ _1372_ /*47106*/;
assign _1379_ = D[31] ^ Q[61] /*47102*/;
assign _1376_ = _800_ & _1379_ /*47098*/;
assign _1377_ = _800_ ^ _1379_ /*47101*/;
assign _1378_ = _1370_ & _1377_ /*47099*/;
assign _1375_ = _1376_ | _1378_ /*47097*/;
assign _1186_ = _1370_ ^ _1377_ /*47100*/;
assign _1384_ = D[32] ^ Q[61] /*47096*/;
assign _1381_ = _801_ & _1384_ /*47092*/;
assign _1382_ = _801_ ^ _1384_ /*47095*/;
assign _1383_ = _1375_ & _1382_ /*47093*/;
assign _1380_ = _1381_ | _1383_ /*47091*/;
assign _1187_ = _1375_ ^ _1382_ /*47094*/;
assign _1389_ = D[33] ^ Q[61] /*47090*/;
assign _1386_ = _802_ & _1389_ /*47086*/;
assign _1387_ = _802_ ^ _1389_ /*47089*/;
assign _1388_ = _1380_ & _1387_ /*47087*/;
assign _1385_ = _1386_ | _1388_ /*47085*/;
assign _1188_ = _1380_ ^ _1387_ /*47088*/;
assign _1394_ = D[34] ^ Q[61] /*47084*/;
assign _1391_ = _803_ & _1394_ /*47080*/;
assign _1392_ = _803_ ^ _1394_ /*47083*/;
assign _1393_ = _1385_ & _1392_ /*47081*/;
assign _1390_ = _1391_ | _1393_ /*47079*/;
assign _1189_ = _1385_ ^ _1392_ /*47082*/;
assign _1399_ = D[35] ^ Q[61] /*47078*/;
assign _1396_ = _804_ & _1399_ /*47074*/;
assign _1397_ = _804_ ^ _1399_ /*47077*/;
assign _1398_ = _1390_ & _1397_ /*47075*/;
assign _1395_ = _1396_ | _1398_ /*47073*/;
assign _1190_ = _1390_ ^ _1397_ /*47076*/;
assign _1404_ = D[36] ^ Q[61] /*47072*/;
assign _1401_ = _805_ & _1404_ /*47068*/;
assign _1402_ = _805_ ^ _1404_ /*47071*/;
assign _1403_ = _1395_ & _1402_ /*47069*/;
assign _1400_ = _1401_ | _1403_ /*47067*/;
assign _1191_ = _1395_ ^ _1402_ /*47070*/;
assign _1409_ = D[37] ^ Q[61] /*47066*/;
assign _1406_ = _806_ & _1409_ /*47062*/;
assign _1407_ = _806_ ^ _1409_ /*47065*/;
assign _1408_ = _1400_ & _1407_ /*47063*/;
assign _1405_ = _1406_ | _1408_ /*47061*/;
assign _1192_ = _1400_ ^ _1407_ /*47064*/;
assign _1414_ = D[38] ^ Q[61] /*47060*/;
assign _1411_ = _807_ & _1414_ /*47056*/;
assign _1412_ = _807_ ^ _1414_ /*47059*/;
assign _1413_ = _1405_ & _1412_ /*47057*/;
assign _1410_ = _1411_ | _1413_ /*47055*/;
assign _1193_ = _1405_ ^ _1412_ /*47058*/;
assign _1419_ = D[39] ^ Q[61] /*47054*/;
assign _1416_ = _808_ & _1419_ /*47050*/;
assign _1417_ = _808_ ^ _1419_ /*47053*/;
assign _1418_ = _1410_ & _1417_ /*47051*/;
assign _1415_ = _1416_ | _1418_ /*47049*/;
assign _1194_ = _1410_ ^ _1417_ /*47052*/;
assign _1424_ = D[40] ^ Q[61] /*47048*/;
assign _1421_ = _809_ & _1424_ /*47044*/;
assign _1422_ = _809_ ^ _1424_ /*47047*/;
assign _1423_ = _1415_ & _1422_ /*47045*/;
assign _1420_ = _1421_ | _1423_ /*47043*/;
assign _1195_ = _1415_ ^ _1422_ /*47046*/;
assign _1429_ = D[41] ^ Q[61] /*47042*/;
assign _1426_ = _810_ & _1429_ /*47038*/;
assign _1427_ = _810_ ^ _1429_ /*47041*/;
assign _1428_ = _1420_ & _1427_ /*47039*/;
assign _1425_ = _1426_ | _1428_ /*47037*/;
assign _1196_ = _1420_ ^ _1427_ /*47040*/;
assign _1434_ = D[42] ^ Q[61] /*47036*/;
assign _1431_ = _811_ & _1434_ /*47032*/;
assign _1432_ = _811_ ^ _1434_ /*47035*/;
assign _1433_ = _1425_ & _1432_ /*47033*/;
assign _1430_ = _1431_ | _1433_ /*47031*/;
assign _1197_ = _1425_ ^ _1432_ /*47034*/;
assign _1439_ = D[43] ^ Q[61] /*47030*/;
assign _1436_ = _812_ & _1439_ /*47026*/;
assign _1437_ = _812_ ^ _1439_ /*47029*/;
assign _1438_ = _1430_ & _1437_ /*47027*/;
assign _1435_ = _1436_ | _1438_ /*47025*/;
assign _1198_ = _1430_ ^ _1437_ /*47028*/;
assign _1444_ = D[44] ^ Q[61] /*47024*/;
assign _1441_ = _813_ & _1444_ /*47020*/;
assign _1442_ = _813_ ^ _1444_ /*47023*/;
assign _1443_ = _1435_ & _1442_ /*47021*/;
assign _1440_ = _1441_ | _1443_ /*47019*/;
assign _1199_ = _1435_ ^ _1442_ /*47022*/;
assign _1449_ = D[45] ^ Q[61] /*47018*/;
assign _1446_ = _814_ & _1449_ /*47014*/;
assign _1447_ = _814_ ^ _1449_ /*47017*/;
assign _1448_ = _1440_ & _1447_ /*47015*/;
assign _1445_ = _1446_ | _1448_ /*47013*/;
assign _1200_ = _1440_ ^ _1447_ /*47016*/;
assign _1454_ = D[46] ^ Q[61] /*47012*/;
assign _1451_ = _815_ & _1454_ /*47008*/;
assign _1452_ = _815_ ^ _1454_ /*47011*/;
assign _1453_ = _1445_ & _1452_ /*47009*/;
assign _1450_ = _1451_ | _1453_ /*47007*/;
assign _1201_ = _1445_ ^ _1452_ /*47010*/;
assign _1459_ = D[47] ^ Q[61] /*47006*/;
assign _1456_ = _816_ & _1459_ /*47002*/;
assign _1457_ = _816_ ^ _1459_ /*47005*/;
assign _1458_ = _1450_ & _1457_ /*47003*/;
assign _1455_ = _1456_ | _1458_ /*47001*/;
assign _1202_ = _1450_ ^ _1457_ /*47004*/;
assign _1464_ = D[48] ^ Q[61] /*47000*/;
assign _1461_ = _817_ & _1464_ /*46996*/;
assign _1462_ = _817_ ^ _1464_ /*46999*/;
assign _1463_ = _1455_ & _1462_ /*46997*/;
assign _1460_ = _1461_ | _1463_ /*46995*/;
assign _1203_ = _1455_ ^ _1462_ /*46998*/;
assign _1469_ = D[49] ^ Q[61] /*46994*/;
assign _1466_ = _818_ & _1469_ /*46990*/;
assign _1467_ = _818_ ^ _1469_ /*46993*/;
assign _1468_ = _1460_ & _1467_ /*46991*/;
assign _1465_ = _1466_ | _1468_ /*46989*/;
assign _1204_ = _1460_ ^ _1467_ /*46992*/;
assign _1474_ = D[50] ^ Q[61] /*46988*/;
assign _1471_ = _819_ & _1474_ /*46984*/;
assign _1472_ = _819_ ^ _1474_ /*46987*/;
assign _1473_ = _1465_ & _1472_ /*46985*/;
assign _1470_ = _1471_ | _1473_ /*46983*/;
assign _1205_ = _1465_ ^ _1472_ /*46986*/;
assign _1479_ = D[51] ^ Q[61] /*46982*/;
assign _1476_ = _820_ & _1479_ /*46978*/;
assign _1477_ = _820_ ^ _1479_ /*46981*/;
assign _1478_ = _1470_ & _1477_ /*46979*/;
assign _1475_ = _1476_ | _1478_ /*46977*/;
assign _1206_ = _1470_ ^ _1477_ /*46980*/;
assign _1484_ = D[52] ^ Q[61] /*46976*/;
assign _1481_ = _821_ & _1484_ /*46972*/;
assign _1482_ = _821_ ^ _1484_ /*46975*/;
assign _1483_ = _1475_ & _1482_ /*46973*/;
assign _1480_ = _1481_ | _1483_ /*46971*/;
assign _1207_ = _1475_ ^ _1482_ /*46974*/;
assign _1489_ = D[53] ^ Q[61] /*46970*/;
assign _1486_ = _822_ & _1489_ /*46966*/;
assign _1487_ = _822_ ^ _1489_ /*46969*/;
assign _1488_ = _1480_ & _1487_ /*46967*/;
assign _1485_ = _1486_ | _1488_ /*46965*/;
assign _1208_ = _1480_ ^ _1487_ /*46968*/;
assign _1494_ = D[54] ^ Q[61] /*46964*/;
assign _1491_ = _823_ & _1494_ /*46960*/;
assign _1492_ = _823_ ^ _1494_ /*46963*/;
assign _1493_ = _1485_ & _1492_ /*46961*/;
assign _1490_ = _1491_ | _1493_ /*46959*/;
assign _1209_ = _1485_ ^ _1492_ /*46962*/;
assign _1499_ = D[55] ^ Q[61] /*46958*/;
assign _1496_ = _824_ & _1499_ /*46954*/;
assign _1497_ = _824_ ^ _1499_ /*46957*/;
assign _1498_ = _1490_ & _1497_ /*46955*/;
assign _1495_ = _1496_ | _1498_ /*46953*/;
assign _1210_ = _1490_ ^ _1497_ /*46956*/;
assign _1504_ = D[56] ^ Q[61] /*46952*/;
assign _1501_ = _825_ & _1504_ /*46948*/;
assign _1502_ = _825_ ^ _1504_ /*46951*/;
assign _1503_ = _1495_ & _1502_ /*46949*/;
assign _1500_ = _1501_ | _1503_ /*46947*/;
assign _1211_ = _1495_ ^ _1502_ /*46950*/;
assign _1509_ = D[57] ^ Q[61] /*46946*/;
assign _1506_ = _826_ & _1509_ /*46942*/;
assign _1507_ = _826_ ^ _1509_ /*46945*/;
assign _1508_ = _1500_ & _1507_ /*46943*/;
assign _1505_ = _1506_ | _1508_ /*46941*/;
assign _1212_ = _1500_ ^ _1507_ /*46944*/;
assign _1514_ = D[58] ^ Q[61] /*46940*/;
assign _1511_ = _827_ & _1514_ /*46936*/;
assign _1512_ = _827_ ^ _1514_ /*46939*/;
assign _1513_ = _1505_ & _1512_ /*46937*/;
assign _1510_ = _1511_ | _1513_ /*46935*/;
assign _1213_ = _1505_ ^ _1512_ /*46938*/;
assign _1519_ = D[59] ^ Q[61] /*46934*/;
assign _1516_ = _828_ & _1519_ /*46930*/;
assign _1517_ = _828_ ^ _1519_ /*46933*/;
assign _1518_ = _1510_ & _1517_ /*46931*/;
assign _1515_ = _1516_ | _1518_ /*46929*/;
assign _1214_ = _1510_ ^ _1517_ /*46932*/;
assign _1524_ = D[60] ^ Q[61] /*46928*/;
assign _1521_ = _829_ & _1524_ /*46924*/;
assign _1522_ = _829_ ^ _1524_ /*46927*/;
assign _1523_ = _1515_ & _1522_ /*46925*/;
assign _1520_ = _1521_ | _1523_ /*46923*/;
assign _1215_ = _1515_ ^ _1522_ /*46926*/;
assign _1529_ = D[61] ^ Q[61] /*46922*/;
assign _1526_ = _830_ & _1529_ /*46918*/;
assign _1527_ = _830_ ^ _1529_ /*46921*/;
assign _1528_ = _1520_ & _1527_ /*46919*/;
assign _1525_ = _1526_ | _1528_ /*46917*/;
assign _1216_ = _1520_ ^ _1527_ /*46920*/;
assign _1534_ = D[62] ^ Q[61] /*46916*/;
assign _1531_ = _831_ & _1534_ /*46912*/;
assign _1532_ = _831_ ^ _1534_ /*46915*/;
assign _1533_ = _1525_ & _1532_ /*46913*/;
assign _1530_ = _1531_ | _1533_ /*46911*/;
assign _1217_ = _1525_ ^ _1532_ /*46914*/;
assign _1538_ = zeroWire ^ Q[61] /*46910*/;
assign _1535_ = _832_ & _1538_ /*46906*/;
assign _1536_ = _832_ ^ _1538_ /*46909*/;
assign _1537_ = _1530_ & _1536_ /*46907*/;
assign Q[60] = _1535_ | _1537_ /*46905*/;
assign _1218_ = _1530_ ^ _1536_ /*46908*/;
assign _1609_ = D[0] ^ Q[60] /*46519*/;
assign _1606_ = R_0[59] & _1609_ /*46515*/;
assign _1607_ = R_0[59] ^ _1609_ /*46518*/;
assign _1608_ = Q[60] & _1607_ /*46516*/;
assign _1605_ = _1606_ | _1608_ /*46514*/;
assign _1540_ = Q[60] ^ _1607_ /*46517*/;
assign _1614_ = D[1] ^ Q[60] /*46513*/;
assign _1611_ = _1155_ & _1614_ /*46509*/;
assign _1612_ = _1155_ ^ _1614_ /*46512*/;
assign _1613_ = _1605_ & _1612_ /*46510*/;
assign _1610_ = _1611_ | _1613_ /*46508*/;
assign _1541_ = _1605_ ^ _1612_ /*46511*/;
assign _1619_ = D[2] ^ Q[60] /*46507*/;
assign _1616_ = _1156_ & _1619_ /*46503*/;
assign _1617_ = _1156_ ^ _1619_ /*46506*/;
assign _1618_ = _1610_ & _1617_ /*46504*/;
assign _1615_ = _1616_ | _1618_ /*46502*/;
assign _1542_ = _1610_ ^ _1617_ /*46505*/;
assign _1624_ = D[3] ^ Q[60] /*46501*/;
assign _1621_ = _1157_ & _1624_ /*46497*/;
assign _1622_ = _1157_ ^ _1624_ /*46500*/;
assign _1623_ = _1615_ & _1622_ /*46498*/;
assign _1620_ = _1621_ | _1623_ /*46496*/;
assign _1543_ = _1615_ ^ _1622_ /*46499*/;
assign _1629_ = D[4] ^ Q[60] /*46495*/;
assign _1626_ = _1158_ & _1629_ /*46491*/;
assign _1627_ = _1158_ ^ _1629_ /*46494*/;
assign _1628_ = _1620_ & _1627_ /*46492*/;
assign _1625_ = _1626_ | _1628_ /*46490*/;
assign _1544_ = _1620_ ^ _1627_ /*46493*/;
assign _1634_ = D[5] ^ Q[60] /*46489*/;
assign _1631_ = _1159_ & _1634_ /*46485*/;
assign _1632_ = _1159_ ^ _1634_ /*46488*/;
assign _1633_ = _1625_ & _1632_ /*46486*/;
assign _1630_ = _1631_ | _1633_ /*46484*/;
assign _1545_ = _1625_ ^ _1632_ /*46487*/;
assign _1639_ = D[6] ^ Q[60] /*46483*/;
assign _1636_ = _1160_ & _1639_ /*46479*/;
assign _1637_ = _1160_ ^ _1639_ /*46482*/;
assign _1638_ = _1630_ & _1637_ /*46480*/;
assign _1635_ = _1636_ | _1638_ /*46478*/;
assign _1546_ = _1630_ ^ _1637_ /*46481*/;
assign _1644_ = D[7] ^ Q[60] /*46477*/;
assign _1641_ = _1161_ & _1644_ /*46473*/;
assign _1642_ = _1161_ ^ _1644_ /*46476*/;
assign _1643_ = _1635_ & _1642_ /*46474*/;
assign _1640_ = _1641_ | _1643_ /*46472*/;
assign _1547_ = _1635_ ^ _1642_ /*46475*/;
assign _1649_ = D[8] ^ Q[60] /*46471*/;
assign _1646_ = _1162_ & _1649_ /*46467*/;
assign _1647_ = _1162_ ^ _1649_ /*46470*/;
assign _1648_ = _1640_ & _1647_ /*46468*/;
assign _1645_ = _1646_ | _1648_ /*46466*/;
assign _1548_ = _1640_ ^ _1647_ /*46469*/;
assign _1654_ = D[9] ^ Q[60] /*46465*/;
assign _1651_ = _1163_ & _1654_ /*46461*/;
assign _1652_ = _1163_ ^ _1654_ /*46464*/;
assign _1653_ = _1645_ & _1652_ /*46462*/;
assign _1650_ = _1651_ | _1653_ /*46460*/;
assign _1549_ = _1645_ ^ _1652_ /*46463*/;
assign _1659_ = D[10] ^ Q[60] /*46459*/;
assign _1656_ = _1164_ & _1659_ /*46455*/;
assign _1657_ = _1164_ ^ _1659_ /*46458*/;
assign _1658_ = _1650_ & _1657_ /*46456*/;
assign _1655_ = _1656_ | _1658_ /*46454*/;
assign _1550_ = _1650_ ^ _1657_ /*46457*/;
assign _1664_ = D[11] ^ Q[60] /*46453*/;
assign _1661_ = _1165_ & _1664_ /*46449*/;
assign _1662_ = _1165_ ^ _1664_ /*46452*/;
assign _1663_ = _1655_ & _1662_ /*46450*/;
assign _1660_ = _1661_ | _1663_ /*46448*/;
assign _1551_ = _1655_ ^ _1662_ /*46451*/;
assign _1669_ = D[12] ^ Q[60] /*46447*/;
assign _1666_ = _1166_ & _1669_ /*46443*/;
assign _1667_ = _1166_ ^ _1669_ /*46446*/;
assign _1668_ = _1660_ & _1667_ /*46444*/;
assign _1665_ = _1666_ | _1668_ /*46442*/;
assign _1552_ = _1660_ ^ _1667_ /*46445*/;
assign _1674_ = D[13] ^ Q[60] /*46441*/;
assign _1671_ = _1167_ & _1674_ /*46437*/;
assign _1672_ = _1167_ ^ _1674_ /*46440*/;
assign _1673_ = _1665_ & _1672_ /*46438*/;
assign _1670_ = _1671_ | _1673_ /*46436*/;
assign _1553_ = _1665_ ^ _1672_ /*46439*/;
assign _1679_ = D[14] ^ Q[60] /*46435*/;
assign _1676_ = _1168_ & _1679_ /*46431*/;
assign _1677_ = _1168_ ^ _1679_ /*46434*/;
assign _1678_ = _1670_ & _1677_ /*46432*/;
assign _1675_ = _1676_ | _1678_ /*46430*/;
assign _1554_ = _1670_ ^ _1677_ /*46433*/;
assign _1684_ = D[15] ^ Q[60] /*46429*/;
assign _1681_ = _1169_ & _1684_ /*46425*/;
assign _1682_ = _1169_ ^ _1684_ /*46428*/;
assign _1683_ = _1675_ & _1682_ /*46426*/;
assign _1680_ = _1681_ | _1683_ /*46424*/;
assign _1555_ = _1675_ ^ _1682_ /*46427*/;
assign _1689_ = D[16] ^ Q[60] /*46423*/;
assign _1686_ = _1170_ & _1689_ /*46419*/;
assign _1687_ = _1170_ ^ _1689_ /*46422*/;
assign _1688_ = _1680_ & _1687_ /*46420*/;
assign _1685_ = _1686_ | _1688_ /*46418*/;
assign _1556_ = _1680_ ^ _1687_ /*46421*/;
assign _1694_ = D[17] ^ Q[60] /*46417*/;
assign _1691_ = _1171_ & _1694_ /*46413*/;
assign _1692_ = _1171_ ^ _1694_ /*46416*/;
assign _1693_ = _1685_ & _1692_ /*46414*/;
assign _1690_ = _1691_ | _1693_ /*46412*/;
assign _1557_ = _1685_ ^ _1692_ /*46415*/;
assign _1699_ = D[18] ^ Q[60] /*46411*/;
assign _1696_ = _1172_ & _1699_ /*46407*/;
assign _1697_ = _1172_ ^ _1699_ /*46410*/;
assign _1698_ = _1690_ & _1697_ /*46408*/;
assign _1695_ = _1696_ | _1698_ /*46406*/;
assign _1558_ = _1690_ ^ _1697_ /*46409*/;
assign _1704_ = D[19] ^ Q[60] /*46405*/;
assign _1701_ = _1173_ & _1704_ /*46401*/;
assign _1702_ = _1173_ ^ _1704_ /*46404*/;
assign _1703_ = _1695_ & _1702_ /*46402*/;
assign _1700_ = _1701_ | _1703_ /*46400*/;
assign _1559_ = _1695_ ^ _1702_ /*46403*/;
assign _1709_ = D[20] ^ Q[60] /*46399*/;
assign _1706_ = _1174_ & _1709_ /*46395*/;
assign _1707_ = _1174_ ^ _1709_ /*46398*/;
assign _1708_ = _1700_ & _1707_ /*46396*/;
assign _1705_ = _1706_ | _1708_ /*46394*/;
assign _1560_ = _1700_ ^ _1707_ /*46397*/;
assign _1714_ = D[21] ^ Q[60] /*46393*/;
assign _1711_ = _1175_ & _1714_ /*46389*/;
assign _1712_ = _1175_ ^ _1714_ /*46392*/;
assign _1713_ = _1705_ & _1712_ /*46390*/;
assign _1710_ = _1711_ | _1713_ /*46388*/;
assign _1561_ = _1705_ ^ _1712_ /*46391*/;
assign _1719_ = D[22] ^ Q[60] /*46387*/;
assign _1716_ = _1176_ & _1719_ /*46383*/;
assign _1717_ = _1176_ ^ _1719_ /*46386*/;
assign _1718_ = _1710_ & _1717_ /*46384*/;
assign _1715_ = _1716_ | _1718_ /*46382*/;
assign _1562_ = _1710_ ^ _1717_ /*46385*/;
assign _1724_ = D[23] ^ Q[60] /*46381*/;
assign _1721_ = _1177_ & _1724_ /*46377*/;
assign _1722_ = _1177_ ^ _1724_ /*46380*/;
assign _1723_ = _1715_ & _1722_ /*46378*/;
assign _1720_ = _1721_ | _1723_ /*46376*/;
assign _1563_ = _1715_ ^ _1722_ /*46379*/;
assign _1729_ = D[24] ^ Q[60] /*46375*/;
assign _1726_ = _1178_ & _1729_ /*46371*/;
assign _1727_ = _1178_ ^ _1729_ /*46374*/;
assign _1728_ = _1720_ & _1727_ /*46372*/;
assign _1725_ = _1726_ | _1728_ /*46370*/;
assign _1564_ = _1720_ ^ _1727_ /*46373*/;
assign _1734_ = D[25] ^ Q[60] /*46369*/;
assign _1731_ = _1179_ & _1734_ /*46365*/;
assign _1732_ = _1179_ ^ _1734_ /*46368*/;
assign _1733_ = _1725_ & _1732_ /*46366*/;
assign _1730_ = _1731_ | _1733_ /*46364*/;
assign _1565_ = _1725_ ^ _1732_ /*46367*/;
assign _1739_ = D[26] ^ Q[60] /*46363*/;
assign _1736_ = _1180_ & _1739_ /*46359*/;
assign _1737_ = _1180_ ^ _1739_ /*46362*/;
assign _1738_ = _1730_ & _1737_ /*46360*/;
assign _1735_ = _1736_ | _1738_ /*46358*/;
assign _1566_ = _1730_ ^ _1737_ /*46361*/;
assign _1744_ = D[27] ^ Q[60] /*46357*/;
assign _1741_ = _1181_ & _1744_ /*46353*/;
assign _1742_ = _1181_ ^ _1744_ /*46356*/;
assign _1743_ = _1735_ & _1742_ /*46354*/;
assign _1740_ = _1741_ | _1743_ /*46352*/;
assign _1567_ = _1735_ ^ _1742_ /*46355*/;
assign _1749_ = D[28] ^ Q[60] /*46351*/;
assign _1746_ = _1182_ & _1749_ /*46347*/;
assign _1747_ = _1182_ ^ _1749_ /*46350*/;
assign _1748_ = _1740_ & _1747_ /*46348*/;
assign _1745_ = _1746_ | _1748_ /*46346*/;
assign _1568_ = _1740_ ^ _1747_ /*46349*/;
assign _1754_ = D[29] ^ Q[60] /*46345*/;
assign _1751_ = _1183_ & _1754_ /*46341*/;
assign _1752_ = _1183_ ^ _1754_ /*46344*/;
assign _1753_ = _1745_ & _1752_ /*46342*/;
assign _1750_ = _1751_ | _1753_ /*46340*/;
assign _1569_ = _1745_ ^ _1752_ /*46343*/;
assign _1759_ = D[30] ^ Q[60] /*46339*/;
assign _1756_ = _1184_ & _1759_ /*46335*/;
assign _1757_ = _1184_ ^ _1759_ /*46338*/;
assign _1758_ = _1750_ & _1757_ /*46336*/;
assign _1755_ = _1756_ | _1758_ /*46334*/;
assign _1570_ = _1750_ ^ _1757_ /*46337*/;
assign _1764_ = D[31] ^ Q[60] /*46333*/;
assign _1761_ = _1185_ & _1764_ /*46329*/;
assign _1762_ = _1185_ ^ _1764_ /*46332*/;
assign _1763_ = _1755_ & _1762_ /*46330*/;
assign _1760_ = _1761_ | _1763_ /*46328*/;
assign _1571_ = _1755_ ^ _1762_ /*46331*/;
assign _1769_ = D[32] ^ Q[60] /*46327*/;
assign _1766_ = _1186_ & _1769_ /*46323*/;
assign _1767_ = _1186_ ^ _1769_ /*46326*/;
assign _1768_ = _1760_ & _1767_ /*46324*/;
assign _1765_ = _1766_ | _1768_ /*46322*/;
assign _1572_ = _1760_ ^ _1767_ /*46325*/;
assign _1774_ = D[33] ^ Q[60] /*46321*/;
assign _1771_ = _1187_ & _1774_ /*46317*/;
assign _1772_ = _1187_ ^ _1774_ /*46320*/;
assign _1773_ = _1765_ & _1772_ /*46318*/;
assign _1770_ = _1771_ | _1773_ /*46316*/;
assign _1573_ = _1765_ ^ _1772_ /*46319*/;
assign _1779_ = D[34] ^ Q[60] /*46315*/;
assign _1776_ = _1188_ & _1779_ /*46311*/;
assign _1777_ = _1188_ ^ _1779_ /*46314*/;
assign _1778_ = _1770_ & _1777_ /*46312*/;
assign _1775_ = _1776_ | _1778_ /*46310*/;
assign _1574_ = _1770_ ^ _1777_ /*46313*/;
assign _1784_ = D[35] ^ Q[60] /*46309*/;
assign _1781_ = _1189_ & _1784_ /*46305*/;
assign _1782_ = _1189_ ^ _1784_ /*46308*/;
assign _1783_ = _1775_ & _1782_ /*46306*/;
assign _1780_ = _1781_ | _1783_ /*46304*/;
assign _1575_ = _1775_ ^ _1782_ /*46307*/;
assign _1789_ = D[36] ^ Q[60] /*46303*/;
assign _1786_ = _1190_ & _1789_ /*46299*/;
assign _1787_ = _1190_ ^ _1789_ /*46302*/;
assign _1788_ = _1780_ & _1787_ /*46300*/;
assign _1785_ = _1786_ | _1788_ /*46298*/;
assign _1576_ = _1780_ ^ _1787_ /*46301*/;
assign _1794_ = D[37] ^ Q[60] /*46297*/;
assign _1791_ = _1191_ & _1794_ /*46293*/;
assign _1792_ = _1191_ ^ _1794_ /*46296*/;
assign _1793_ = _1785_ & _1792_ /*46294*/;
assign _1790_ = _1791_ | _1793_ /*46292*/;
assign _1577_ = _1785_ ^ _1792_ /*46295*/;
assign _1799_ = D[38] ^ Q[60] /*46291*/;
assign _1796_ = _1192_ & _1799_ /*46287*/;
assign _1797_ = _1192_ ^ _1799_ /*46290*/;
assign _1798_ = _1790_ & _1797_ /*46288*/;
assign _1795_ = _1796_ | _1798_ /*46286*/;
assign _1578_ = _1790_ ^ _1797_ /*46289*/;
assign _1804_ = D[39] ^ Q[60] /*46285*/;
assign _1801_ = _1193_ & _1804_ /*46281*/;
assign _1802_ = _1193_ ^ _1804_ /*46284*/;
assign _1803_ = _1795_ & _1802_ /*46282*/;
assign _1800_ = _1801_ | _1803_ /*46280*/;
assign _1579_ = _1795_ ^ _1802_ /*46283*/;
assign _1809_ = D[40] ^ Q[60] /*46279*/;
assign _1806_ = _1194_ & _1809_ /*46275*/;
assign _1807_ = _1194_ ^ _1809_ /*46278*/;
assign _1808_ = _1800_ & _1807_ /*46276*/;
assign _1805_ = _1806_ | _1808_ /*46274*/;
assign _1580_ = _1800_ ^ _1807_ /*46277*/;
assign _1814_ = D[41] ^ Q[60] /*46273*/;
assign _1811_ = _1195_ & _1814_ /*46269*/;
assign _1812_ = _1195_ ^ _1814_ /*46272*/;
assign _1813_ = _1805_ & _1812_ /*46270*/;
assign _1810_ = _1811_ | _1813_ /*46268*/;
assign _1581_ = _1805_ ^ _1812_ /*46271*/;
assign _1819_ = D[42] ^ Q[60] /*46267*/;
assign _1816_ = _1196_ & _1819_ /*46263*/;
assign _1817_ = _1196_ ^ _1819_ /*46266*/;
assign _1818_ = _1810_ & _1817_ /*46264*/;
assign _1815_ = _1816_ | _1818_ /*46262*/;
assign _1582_ = _1810_ ^ _1817_ /*46265*/;
assign _1824_ = D[43] ^ Q[60] /*46261*/;
assign _1821_ = _1197_ & _1824_ /*46257*/;
assign _1822_ = _1197_ ^ _1824_ /*46260*/;
assign _1823_ = _1815_ & _1822_ /*46258*/;
assign _1820_ = _1821_ | _1823_ /*46256*/;
assign _1583_ = _1815_ ^ _1822_ /*46259*/;
assign _1829_ = D[44] ^ Q[60] /*46255*/;
assign _1826_ = _1198_ & _1829_ /*46251*/;
assign _1827_ = _1198_ ^ _1829_ /*46254*/;
assign _1828_ = _1820_ & _1827_ /*46252*/;
assign _1825_ = _1826_ | _1828_ /*46250*/;
assign _1584_ = _1820_ ^ _1827_ /*46253*/;
assign _1834_ = D[45] ^ Q[60] /*46249*/;
assign _1831_ = _1199_ & _1834_ /*46245*/;
assign _1832_ = _1199_ ^ _1834_ /*46248*/;
assign _1833_ = _1825_ & _1832_ /*46246*/;
assign _1830_ = _1831_ | _1833_ /*46244*/;
assign _1585_ = _1825_ ^ _1832_ /*46247*/;
assign _1839_ = D[46] ^ Q[60] /*46243*/;
assign _1836_ = _1200_ & _1839_ /*46239*/;
assign _1837_ = _1200_ ^ _1839_ /*46242*/;
assign _1838_ = _1830_ & _1837_ /*46240*/;
assign _1835_ = _1836_ | _1838_ /*46238*/;
assign _1586_ = _1830_ ^ _1837_ /*46241*/;
assign _1844_ = D[47] ^ Q[60] /*46237*/;
assign _1841_ = _1201_ & _1844_ /*46233*/;
assign _1842_ = _1201_ ^ _1844_ /*46236*/;
assign _1843_ = _1835_ & _1842_ /*46234*/;
assign _1840_ = _1841_ | _1843_ /*46232*/;
assign _1587_ = _1835_ ^ _1842_ /*46235*/;
assign _1849_ = D[48] ^ Q[60] /*46231*/;
assign _1846_ = _1202_ & _1849_ /*46227*/;
assign _1847_ = _1202_ ^ _1849_ /*46230*/;
assign _1848_ = _1840_ & _1847_ /*46228*/;
assign _1845_ = _1846_ | _1848_ /*46226*/;
assign _1588_ = _1840_ ^ _1847_ /*46229*/;
assign _1854_ = D[49] ^ Q[60] /*46225*/;
assign _1851_ = _1203_ & _1854_ /*46221*/;
assign _1852_ = _1203_ ^ _1854_ /*46224*/;
assign _1853_ = _1845_ & _1852_ /*46222*/;
assign _1850_ = _1851_ | _1853_ /*46220*/;
assign _1589_ = _1845_ ^ _1852_ /*46223*/;
assign _1859_ = D[50] ^ Q[60] /*46219*/;
assign _1856_ = _1204_ & _1859_ /*46215*/;
assign _1857_ = _1204_ ^ _1859_ /*46218*/;
assign _1858_ = _1850_ & _1857_ /*46216*/;
assign _1855_ = _1856_ | _1858_ /*46214*/;
assign _1590_ = _1850_ ^ _1857_ /*46217*/;
assign _1864_ = D[51] ^ Q[60] /*46213*/;
assign _1861_ = _1205_ & _1864_ /*46209*/;
assign _1862_ = _1205_ ^ _1864_ /*46212*/;
assign _1863_ = _1855_ & _1862_ /*46210*/;
assign _1860_ = _1861_ | _1863_ /*46208*/;
assign _1591_ = _1855_ ^ _1862_ /*46211*/;
assign _1869_ = D[52] ^ Q[60] /*46207*/;
assign _1866_ = _1206_ & _1869_ /*46203*/;
assign _1867_ = _1206_ ^ _1869_ /*46206*/;
assign _1868_ = _1860_ & _1867_ /*46204*/;
assign _1865_ = _1866_ | _1868_ /*46202*/;
assign _1592_ = _1860_ ^ _1867_ /*46205*/;
assign _1874_ = D[53] ^ Q[60] /*46201*/;
assign _1871_ = _1207_ & _1874_ /*46197*/;
assign _1872_ = _1207_ ^ _1874_ /*46200*/;
assign _1873_ = _1865_ & _1872_ /*46198*/;
assign _1870_ = _1871_ | _1873_ /*46196*/;
assign _1593_ = _1865_ ^ _1872_ /*46199*/;
assign _1879_ = D[54] ^ Q[60] /*46195*/;
assign _1876_ = _1208_ & _1879_ /*46191*/;
assign _1877_ = _1208_ ^ _1879_ /*46194*/;
assign _1878_ = _1870_ & _1877_ /*46192*/;
assign _1875_ = _1876_ | _1878_ /*46190*/;
assign _1594_ = _1870_ ^ _1877_ /*46193*/;
assign _1884_ = D[55] ^ Q[60] /*46189*/;
assign _1881_ = _1209_ & _1884_ /*46185*/;
assign _1882_ = _1209_ ^ _1884_ /*46188*/;
assign _1883_ = _1875_ & _1882_ /*46186*/;
assign _1880_ = _1881_ | _1883_ /*46184*/;
assign _1595_ = _1875_ ^ _1882_ /*46187*/;
assign _1889_ = D[56] ^ Q[60] /*46183*/;
assign _1886_ = _1210_ & _1889_ /*46179*/;
assign _1887_ = _1210_ ^ _1889_ /*46182*/;
assign _1888_ = _1880_ & _1887_ /*46180*/;
assign _1885_ = _1886_ | _1888_ /*46178*/;
assign _1596_ = _1880_ ^ _1887_ /*46181*/;
assign _1894_ = D[57] ^ Q[60] /*46177*/;
assign _1891_ = _1211_ & _1894_ /*46173*/;
assign _1892_ = _1211_ ^ _1894_ /*46176*/;
assign _1893_ = _1885_ & _1892_ /*46174*/;
assign _1890_ = _1891_ | _1893_ /*46172*/;
assign _1597_ = _1885_ ^ _1892_ /*46175*/;
assign _1899_ = D[58] ^ Q[60] /*46171*/;
assign _1896_ = _1212_ & _1899_ /*46167*/;
assign _1897_ = _1212_ ^ _1899_ /*46170*/;
assign _1898_ = _1890_ & _1897_ /*46168*/;
assign _1895_ = _1896_ | _1898_ /*46166*/;
assign _1598_ = _1890_ ^ _1897_ /*46169*/;
assign _1904_ = D[59] ^ Q[60] /*46165*/;
assign _1901_ = _1213_ & _1904_ /*46161*/;
assign _1902_ = _1213_ ^ _1904_ /*46164*/;
assign _1903_ = _1895_ & _1902_ /*46162*/;
assign _1900_ = _1901_ | _1903_ /*46160*/;
assign _1599_ = _1895_ ^ _1902_ /*46163*/;
assign _1909_ = D[60] ^ Q[60] /*46159*/;
assign _1906_ = _1214_ & _1909_ /*46155*/;
assign _1907_ = _1214_ ^ _1909_ /*46158*/;
assign _1908_ = _1900_ & _1907_ /*46156*/;
assign _1905_ = _1906_ | _1908_ /*46154*/;
assign _1600_ = _1900_ ^ _1907_ /*46157*/;
assign _1914_ = D[61] ^ Q[60] /*46153*/;
assign _1911_ = _1215_ & _1914_ /*46149*/;
assign _1912_ = _1215_ ^ _1914_ /*46152*/;
assign _1913_ = _1905_ & _1912_ /*46150*/;
assign _1910_ = _1911_ | _1913_ /*46148*/;
assign _1601_ = _1905_ ^ _1912_ /*46151*/;
assign _1919_ = D[62] ^ Q[60] /*46147*/;
assign _1916_ = _1216_ & _1919_ /*46143*/;
assign _1917_ = _1216_ ^ _1919_ /*46146*/;
assign _1918_ = _1910_ & _1917_ /*46144*/;
assign _1915_ = _1916_ | _1918_ /*46142*/;
assign _1602_ = _1910_ ^ _1917_ /*46145*/;
assign _1923_ = zeroWire ^ Q[60] /*46141*/;
assign _1920_ = _1217_ & _1923_ /*46137*/;
assign _1921_ = _1217_ ^ _1923_ /*46140*/;
assign _1922_ = _1915_ & _1921_ /*46138*/;
assign Q[59] = _1920_ | _1922_ /*46136*/;
assign _1603_ = _1915_ ^ _1921_ /*46139*/;
assign _1994_ = D[0] ^ Q[59] /*45750*/;
assign _1991_ = R_0[58] & _1994_ /*45746*/;
assign _1992_ = R_0[58] ^ _1994_ /*45749*/;
assign _1993_ = Q[59] & _1992_ /*45747*/;
assign _1990_ = _1991_ | _1993_ /*45745*/;
assign _1925_ = Q[59] ^ _1992_ /*45748*/;
assign _1999_ = D[1] ^ Q[59] /*45744*/;
assign _1996_ = _1540_ & _1999_ /*45740*/;
assign _1997_ = _1540_ ^ _1999_ /*45743*/;
assign _1998_ = _1990_ & _1997_ /*45741*/;
assign _1995_ = _1996_ | _1998_ /*45739*/;
assign _1926_ = _1990_ ^ _1997_ /*45742*/;
assign _2004_ = D[2] ^ Q[59] /*45738*/;
assign _2001_ = _1541_ & _2004_ /*45734*/;
assign _2002_ = _1541_ ^ _2004_ /*45737*/;
assign _2003_ = _1995_ & _2002_ /*45735*/;
assign _2000_ = _2001_ | _2003_ /*45733*/;
assign _1927_ = _1995_ ^ _2002_ /*45736*/;
assign _2009_ = D[3] ^ Q[59] /*45732*/;
assign _2006_ = _1542_ & _2009_ /*45728*/;
assign _2007_ = _1542_ ^ _2009_ /*45731*/;
assign _2008_ = _2000_ & _2007_ /*45729*/;
assign _2005_ = _2006_ | _2008_ /*45727*/;
assign _1928_ = _2000_ ^ _2007_ /*45730*/;
assign _2014_ = D[4] ^ Q[59] /*45726*/;
assign _2011_ = _1543_ & _2014_ /*45722*/;
assign _2012_ = _1543_ ^ _2014_ /*45725*/;
assign _2013_ = _2005_ & _2012_ /*45723*/;
assign _2010_ = _2011_ | _2013_ /*45721*/;
assign _1929_ = _2005_ ^ _2012_ /*45724*/;
assign _2019_ = D[5] ^ Q[59] /*45720*/;
assign _2016_ = _1544_ & _2019_ /*45716*/;
assign _2017_ = _1544_ ^ _2019_ /*45719*/;
assign _2018_ = _2010_ & _2017_ /*45717*/;
assign _2015_ = _2016_ | _2018_ /*45715*/;
assign _1930_ = _2010_ ^ _2017_ /*45718*/;
assign _2024_ = D[6] ^ Q[59] /*45714*/;
assign _2021_ = _1545_ & _2024_ /*45710*/;
assign _2022_ = _1545_ ^ _2024_ /*45713*/;
assign _2023_ = _2015_ & _2022_ /*45711*/;
assign _2020_ = _2021_ | _2023_ /*45709*/;
assign _1931_ = _2015_ ^ _2022_ /*45712*/;
assign _2029_ = D[7] ^ Q[59] /*45708*/;
assign _2026_ = _1546_ & _2029_ /*45704*/;
assign _2027_ = _1546_ ^ _2029_ /*45707*/;
assign _2028_ = _2020_ & _2027_ /*45705*/;
assign _2025_ = _2026_ | _2028_ /*45703*/;
assign _1932_ = _2020_ ^ _2027_ /*45706*/;
assign _2034_ = D[8] ^ Q[59] /*45702*/;
assign _2031_ = _1547_ & _2034_ /*45698*/;
assign _2032_ = _1547_ ^ _2034_ /*45701*/;
assign _2033_ = _2025_ & _2032_ /*45699*/;
assign _2030_ = _2031_ | _2033_ /*45697*/;
assign _1933_ = _2025_ ^ _2032_ /*45700*/;
assign _2039_ = D[9] ^ Q[59] /*45696*/;
assign _2036_ = _1548_ & _2039_ /*45692*/;
assign _2037_ = _1548_ ^ _2039_ /*45695*/;
assign _2038_ = _2030_ & _2037_ /*45693*/;
assign _2035_ = _2036_ | _2038_ /*45691*/;
assign _1934_ = _2030_ ^ _2037_ /*45694*/;
assign _2044_ = D[10] ^ Q[59] /*45690*/;
assign _2041_ = _1549_ & _2044_ /*45686*/;
assign _2042_ = _1549_ ^ _2044_ /*45689*/;
assign _2043_ = _2035_ & _2042_ /*45687*/;
assign _2040_ = _2041_ | _2043_ /*45685*/;
assign _1935_ = _2035_ ^ _2042_ /*45688*/;
assign _2049_ = D[11] ^ Q[59] /*45684*/;
assign _2046_ = _1550_ & _2049_ /*45680*/;
assign _2047_ = _1550_ ^ _2049_ /*45683*/;
assign _2048_ = _2040_ & _2047_ /*45681*/;
assign _2045_ = _2046_ | _2048_ /*45679*/;
assign _1936_ = _2040_ ^ _2047_ /*45682*/;
assign _2054_ = D[12] ^ Q[59] /*45678*/;
assign _2051_ = _1551_ & _2054_ /*45674*/;
assign _2052_ = _1551_ ^ _2054_ /*45677*/;
assign _2053_ = _2045_ & _2052_ /*45675*/;
assign _2050_ = _2051_ | _2053_ /*45673*/;
assign _1937_ = _2045_ ^ _2052_ /*45676*/;
assign _2059_ = D[13] ^ Q[59] /*45672*/;
assign _2056_ = _1552_ & _2059_ /*45668*/;
assign _2057_ = _1552_ ^ _2059_ /*45671*/;
assign _2058_ = _2050_ & _2057_ /*45669*/;
assign _2055_ = _2056_ | _2058_ /*45667*/;
assign _1938_ = _2050_ ^ _2057_ /*45670*/;
assign _2064_ = D[14] ^ Q[59] /*45666*/;
assign _2061_ = _1553_ & _2064_ /*45662*/;
assign _2062_ = _1553_ ^ _2064_ /*45665*/;
assign _2063_ = _2055_ & _2062_ /*45663*/;
assign _2060_ = _2061_ | _2063_ /*45661*/;
assign _1939_ = _2055_ ^ _2062_ /*45664*/;
assign _2069_ = D[15] ^ Q[59] /*45660*/;
assign _2066_ = _1554_ & _2069_ /*45656*/;
assign _2067_ = _1554_ ^ _2069_ /*45659*/;
assign _2068_ = _2060_ & _2067_ /*45657*/;
assign _2065_ = _2066_ | _2068_ /*45655*/;
assign _1940_ = _2060_ ^ _2067_ /*45658*/;
assign _2074_ = D[16] ^ Q[59] /*45654*/;
assign _2071_ = _1555_ & _2074_ /*45650*/;
assign _2072_ = _1555_ ^ _2074_ /*45653*/;
assign _2073_ = _2065_ & _2072_ /*45651*/;
assign _2070_ = _2071_ | _2073_ /*45649*/;
assign _1941_ = _2065_ ^ _2072_ /*45652*/;
assign _2079_ = D[17] ^ Q[59] /*45648*/;
assign _2076_ = _1556_ & _2079_ /*45644*/;
assign _2077_ = _1556_ ^ _2079_ /*45647*/;
assign _2078_ = _2070_ & _2077_ /*45645*/;
assign _2075_ = _2076_ | _2078_ /*45643*/;
assign _1942_ = _2070_ ^ _2077_ /*45646*/;
assign _2084_ = D[18] ^ Q[59] /*45642*/;
assign _2081_ = _1557_ & _2084_ /*45638*/;
assign _2082_ = _1557_ ^ _2084_ /*45641*/;
assign _2083_ = _2075_ & _2082_ /*45639*/;
assign _2080_ = _2081_ | _2083_ /*45637*/;
assign _1943_ = _2075_ ^ _2082_ /*45640*/;
assign _2089_ = D[19] ^ Q[59] /*45636*/;
assign _2086_ = _1558_ & _2089_ /*45632*/;
assign _2087_ = _1558_ ^ _2089_ /*45635*/;
assign _2088_ = _2080_ & _2087_ /*45633*/;
assign _2085_ = _2086_ | _2088_ /*45631*/;
assign _1944_ = _2080_ ^ _2087_ /*45634*/;
assign _2094_ = D[20] ^ Q[59] /*45630*/;
assign _2091_ = _1559_ & _2094_ /*45626*/;
assign _2092_ = _1559_ ^ _2094_ /*45629*/;
assign _2093_ = _2085_ & _2092_ /*45627*/;
assign _2090_ = _2091_ | _2093_ /*45625*/;
assign _1945_ = _2085_ ^ _2092_ /*45628*/;
assign _2099_ = D[21] ^ Q[59] /*45624*/;
assign _2096_ = _1560_ & _2099_ /*45620*/;
assign _2097_ = _1560_ ^ _2099_ /*45623*/;
assign _2098_ = _2090_ & _2097_ /*45621*/;
assign _2095_ = _2096_ | _2098_ /*45619*/;
assign _1946_ = _2090_ ^ _2097_ /*45622*/;
assign _2104_ = D[22] ^ Q[59] /*45618*/;
assign _2101_ = _1561_ & _2104_ /*45614*/;
assign _2102_ = _1561_ ^ _2104_ /*45617*/;
assign _2103_ = _2095_ & _2102_ /*45615*/;
assign _2100_ = _2101_ | _2103_ /*45613*/;
assign _1947_ = _2095_ ^ _2102_ /*45616*/;
assign _2109_ = D[23] ^ Q[59] /*45612*/;
assign _2106_ = _1562_ & _2109_ /*45608*/;
assign _2107_ = _1562_ ^ _2109_ /*45611*/;
assign _2108_ = _2100_ & _2107_ /*45609*/;
assign _2105_ = _2106_ | _2108_ /*45607*/;
assign _1948_ = _2100_ ^ _2107_ /*45610*/;
assign _2114_ = D[24] ^ Q[59] /*45606*/;
assign _2111_ = _1563_ & _2114_ /*45602*/;
assign _2112_ = _1563_ ^ _2114_ /*45605*/;
assign _2113_ = _2105_ & _2112_ /*45603*/;
assign _2110_ = _2111_ | _2113_ /*45601*/;
assign _1949_ = _2105_ ^ _2112_ /*45604*/;
assign _2119_ = D[25] ^ Q[59] /*45600*/;
assign _2116_ = _1564_ & _2119_ /*45596*/;
assign _2117_ = _1564_ ^ _2119_ /*45599*/;
assign _2118_ = _2110_ & _2117_ /*45597*/;
assign _2115_ = _2116_ | _2118_ /*45595*/;
assign _1950_ = _2110_ ^ _2117_ /*45598*/;
assign _2124_ = D[26] ^ Q[59] /*45594*/;
assign _2121_ = _1565_ & _2124_ /*45590*/;
assign _2122_ = _1565_ ^ _2124_ /*45593*/;
assign _2123_ = _2115_ & _2122_ /*45591*/;
assign _2120_ = _2121_ | _2123_ /*45589*/;
assign _1951_ = _2115_ ^ _2122_ /*45592*/;
assign _2129_ = D[27] ^ Q[59] /*45588*/;
assign _2126_ = _1566_ & _2129_ /*45584*/;
assign _2127_ = _1566_ ^ _2129_ /*45587*/;
assign _2128_ = _2120_ & _2127_ /*45585*/;
assign _2125_ = _2126_ | _2128_ /*45583*/;
assign _1952_ = _2120_ ^ _2127_ /*45586*/;
assign _2134_ = D[28] ^ Q[59] /*45582*/;
assign _2131_ = _1567_ & _2134_ /*45578*/;
assign _2132_ = _1567_ ^ _2134_ /*45581*/;
assign _2133_ = _2125_ & _2132_ /*45579*/;
assign _2130_ = _2131_ | _2133_ /*45577*/;
assign _1953_ = _2125_ ^ _2132_ /*45580*/;
assign _2139_ = D[29] ^ Q[59] /*45576*/;
assign _2136_ = _1568_ & _2139_ /*45572*/;
assign _2137_ = _1568_ ^ _2139_ /*45575*/;
assign _2138_ = _2130_ & _2137_ /*45573*/;
assign _2135_ = _2136_ | _2138_ /*45571*/;
assign _1954_ = _2130_ ^ _2137_ /*45574*/;
assign _2144_ = D[30] ^ Q[59] /*45570*/;
assign _2141_ = _1569_ & _2144_ /*45566*/;
assign _2142_ = _1569_ ^ _2144_ /*45569*/;
assign _2143_ = _2135_ & _2142_ /*45567*/;
assign _2140_ = _2141_ | _2143_ /*45565*/;
assign _1955_ = _2135_ ^ _2142_ /*45568*/;
assign _2149_ = D[31] ^ Q[59] /*45564*/;
assign _2146_ = _1570_ & _2149_ /*45560*/;
assign _2147_ = _1570_ ^ _2149_ /*45563*/;
assign _2148_ = _2140_ & _2147_ /*45561*/;
assign _2145_ = _2146_ | _2148_ /*45559*/;
assign _1956_ = _2140_ ^ _2147_ /*45562*/;
assign _2154_ = D[32] ^ Q[59] /*45558*/;
assign _2151_ = _1571_ & _2154_ /*45554*/;
assign _2152_ = _1571_ ^ _2154_ /*45557*/;
assign _2153_ = _2145_ & _2152_ /*45555*/;
assign _2150_ = _2151_ | _2153_ /*45553*/;
assign _1957_ = _2145_ ^ _2152_ /*45556*/;
assign _2159_ = D[33] ^ Q[59] /*45552*/;
assign _2156_ = _1572_ & _2159_ /*45548*/;
assign _2157_ = _1572_ ^ _2159_ /*45551*/;
assign _2158_ = _2150_ & _2157_ /*45549*/;
assign _2155_ = _2156_ | _2158_ /*45547*/;
assign _1958_ = _2150_ ^ _2157_ /*45550*/;
assign _2164_ = D[34] ^ Q[59] /*45546*/;
assign _2161_ = _1573_ & _2164_ /*45542*/;
assign _2162_ = _1573_ ^ _2164_ /*45545*/;
assign _2163_ = _2155_ & _2162_ /*45543*/;
assign _2160_ = _2161_ | _2163_ /*45541*/;
assign _1959_ = _2155_ ^ _2162_ /*45544*/;
assign _2169_ = D[35] ^ Q[59] /*45540*/;
assign _2166_ = _1574_ & _2169_ /*45536*/;
assign _2167_ = _1574_ ^ _2169_ /*45539*/;
assign _2168_ = _2160_ & _2167_ /*45537*/;
assign _2165_ = _2166_ | _2168_ /*45535*/;
assign _1960_ = _2160_ ^ _2167_ /*45538*/;
assign _2174_ = D[36] ^ Q[59] /*45534*/;
assign _2171_ = _1575_ & _2174_ /*45530*/;
assign _2172_ = _1575_ ^ _2174_ /*45533*/;
assign _2173_ = _2165_ & _2172_ /*45531*/;
assign _2170_ = _2171_ | _2173_ /*45529*/;
assign _1961_ = _2165_ ^ _2172_ /*45532*/;
assign _2179_ = D[37] ^ Q[59] /*45528*/;
assign _2176_ = _1576_ & _2179_ /*45524*/;
assign _2177_ = _1576_ ^ _2179_ /*45527*/;
assign _2178_ = _2170_ & _2177_ /*45525*/;
assign _2175_ = _2176_ | _2178_ /*45523*/;
assign _1962_ = _2170_ ^ _2177_ /*45526*/;
assign _2184_ = D[38] ^ Q[59] /*45522*/;
assign _2181_ = _1577_ & _2184_ /*45518*/;
assign _2182_ = _1577_ ^ _2184_ /*45521*/;
assign _2183_ = _2175_ & _2182_ /*45519*/;
assign _2180_ = _2181_ | _2183_ /*45517*/;
assign _1963_ = _2175_ ^ _2182_ /*45520*/;
assign _2189_ = D[39] ^ Q[59] /*45516*/;
assign _2186_ = _1578_ & _2189_ /*45512*/;
assign _2187_ = _1578_ ^ _2189_ /*45515*/;
assign _2188_ = _2180_ & _2187_ /*45513*/;
assign _2185_ = _2186_ | _2188_ /*45511*/;
assign _1964_ = _2180_ ^ _2187_ /*45514*/;
assign _2194_ = D[40] ^ Q[59] /*45510*/;
assign _2191_ = _1579_ & _2194_ /*45506*/;
assign _2192_ = _1579_ ^ _2194_ /*45509*/;
assign _2193_ = _2185_ & _2192_ /*45507*/;
assign _2190_ = _2191_ | _2193_ /*45505*/;
assign _1965_ = _2185_ ^ _2192_ /*45508*/;
assign _2199_ = D[41] ^ Q[59] /*45504*/;
assign _2196_ = _1580_ & _2199_ /*45500*/;
assign _2197_ = _1580_ ^ _2199_ /*45503*/;
assign _2198_ = _2190_ & _2197_ /*45501*/;
assign _2195_ = _2196_ | _2198_ /*45499*/;
assign _1966_ = _2190_ ^ _2197_ /*45502*/;
assign _2204_ = D[42] ^ Q[59] /*45498*/;
assign _2201_ = _1581_ & _2204_ /*45494*/;
assign _2202_ = _1581_ ^ _2204_ /*45497*/;
assign _2203_ = _2195_ & _2202_ /*45495*/;
assign _2200_ = _2201_ | _2203_ /*45493*/;
assign _1967_ = _2195_ ^ _2202_ /*45496*/;
assign _2209_ = D[43] ^ Q[59] /*45492*/;
assign _2206_ = _1582_ & _2209_ /*45488*/;
assign _2207_ = _1582_ ^ _2209_ /*45491*/;
assign _2208_ = _2200_ & _2207_ /*45489*/;
assign _2205_ = _2206_ | _2208_ /*45487*/;
assign _1968_ = _2200_ ^ _2207_ /*45490*/;
assign _2214_ = D[44] ^ Q[59] /*45486*/;
assign _2211_ = _1583_ & _2214_ /*45482*/;
assign _2212_ = _1583_ ^ _2214_ /*45485*/;
assign _2213_ = _2205_ & _2212_ /*45483*/;
assign _2210_ = _2211_ | _2213_ /*45481*/;
assign _1969_ = _2205_ ^ _2212_ /*45484*/;
assign _2219_ = D[45] ^ Q[59] /*45480*/;
assign _2216_ = _1584_ & _2219_ /*45476*/;
assign _2217_ = _1584_ ^ _2219_ /*45479*/;
assign _2218_ = _2210_ & _2217_ /*45477*/;
assign _2215_ = _2216_ | _2218_ /*45475*/;
assign _1970_ = _2210_ ^ _2217_ /*45478*/;
assign _2224_ = D[46] ^ Q[59] /*45474*/;
assign _2221_ = _1585_ & _2224_ /*45470*/;
assign _2222_ = _1585_ ^ _2224_ /*45473*/;
assign _2223_ = _2215_ & _2222_ /*45471*/;
assign _2220_ = _2221_ | _2223_ /*45469*/;
assign _1971_ = _2215_ ^ _2222_ /*45472*/;
assign _2229_ = D[47] ^ Q[59] /*45468*/;
assign _2226_ = _1586_ & _2229_ /*45464*/;
assign _2227_ = _1586_ ^ _2229_ /*45467*/;
assign _2228_ = _2220_ & _2227_ /*45465*/;
assign _2225_ = _2226_ | _2228_ /*45463*/;
assign _1972_ = _2220_ ^ _2227_ /*45466*/;
assign _2234_ = D[48] ^ Q[59] /*45462*/;
assign _2231_ = _1587_ & _2234_ /*45458*/;
assign _2232_ = _1587_ ^ _2234_ /*45461*/;
assign _2233_ = _2225_ & _2232_ /*45459*/;
assign _2230_ = _2231_ | _2233_ /*45457*/;
assign _1973_ = _2225_ ^ _2232_ /*45460*/;
assign _2239_ = D[49] ^ Q[59] /*45456*/;
assign _2236_ = _1588_ & _2239_ /*45452*/;
assign _2237_ = _1588_ ^ _2239_ /*45455*/;
assign _2238_ = _2230_ & _2237_ /*45453*/;
assign _2235_ = _2236_ | _2238_ /*45451*/;
assign _1974_ = _2230_ ^ _2237_ /*45454*/;
assign _2244_ = D[50] ^ Q[59] /*45450*/;
assign _2241_ = _1589_ & _2244_ /*45446*/;
assign _2242_ = _1589_ ^ _2244_ /*45449*/;
assign _2243_ = _2235_ & _2242_ /*45447*/;
assign _2240_ = _2241_ | _2243_ /*45445*/;
assign _1975_ = _2235_ ^ _2242_ /*45448*/;
assign _2249_ = D[51] ^ Q[59] /*45444*/;
assign _2246_ = _1590_ & _2249_ /*45440*/;
assign _2247_ = _1590_ ^ _2249_ /*45443*/;
assign _2248_ = _2240_ & _2247_ /*45441*/;
assign _2245_ = _2246_ | _2248_ /*45439*/;
assign _1976_ = _2240_ ^ _2247_ /*45442*/;
assign _2254_ = D[52] ^ Q[59] /*45438*/;
assign _2251_ = _1591_ & _2254_ /*45434*/;
assign _2252_ = _1591_ ^ _2254_ /*45437*/;
assign _2253_ = _2245_ & _2252_ /*45435*/;
assign _2250_ = _2251_ | _2253_ /*45433*/;
assign _1977_ = _2245_ ^ _2252_ /*45436*/;
assign _2259_ = D[53] ^ Q[59] /*45432*/;
assign _2256_ = _1592_ & _2259_ /*45428*/;
assign _2257_ = _1592_ ^ _2259_ /*45431*/;
assign _2258_ = _2250_ & _2257_ /*45429*/;
assign _2255_ = _2256_ | _2258_ /*45427*/;
assign _1978_ = _2250_ ^ _2257_ /*45430*/;
assign _2264_ = D[54] ^ Q[59] /*45426*/;
assign _2261_ = _1593_ & _2264_ /*45422*/;
assign _2262_ = _1593_ ^ _2264_ /*45425*/;
assign _2263_ = _2255_ & _2262_ /*45423*/;
assign _2260_ = _2261_ | _2263_ /*45421*/;
assign _1979_ = _2255_ ^ _2262_ /*45424*/;
assign _2269_ = D[55] ^ Q[59] /*45420*/;
assign _2266_ = _1594_ & _2269_ /*45416*/;
assign _2267_ = _1594_ ^ _2269_ /*45419*/;
assign _2268_ = _2260_ & _2267_ /*45417*/;
assign _2265_ = _2266_ | _2268_ /*45415*/;
assign _1980_ = _2260_ ^ _2267_ /*45418*/;
assign _2274_ = D[56] ^ Q[59] /*45414*/;
assign _2271_ = _1595_ & _2274_ /*45410*/;
assign _2272_ = _1595_ ^ _2274_ /*45413*/;
assign _2273_ = _2265_ & _2272_ /*45411*/;
assign _2270_ = _2271_ | _2273_ /*45409*/;
assign _1981_ = _2265_ ^ _2272_ /*45412*/;
assign _2279_ = D[57] ^ Q[59] /*45408*/;
assign _2276_ = _1596_ & _2279_ /*45404*/;
assign _2277_ = _1596_ ^ _2279_ /*45407*/;
assign _2278_ = _2270_ & _2277_ /*45405*/;
assign _2275_ = _2276_ | _2278_ /*45403*/;
assign _1982_ = _2270_ ^ _2277_ /*45406*/;
assign _2284_ = D[58] ^ Q[59] /*45402*/;
assign _2281_ = _1597_ & _2284_ /*45398*/;
assign _2282_ = _1597_ ^ _2284_ /*45401*/;
assign _2283_ = _2275_ & _2282_ /*45399*/;
assign _2280_ = _2281_ | _2283_ /*45397*/;
assign _1983_ = _2275_ ^ _2282_ /*45400*/;
assign _2289_ = D[59] ^ Q[59] /*45396*/;
assign _2286_ = _1598_ & _2289_ /*45392*/;
assign _2287_ = _1598_ ^ _2289_ /*45395*/;
assign _2288_ = _2280_ & _2287_ /*45393*/;
assign _2285_ = _2286_ | _2288_ /*45391*/;
assign _1984_ = _2280_ ^ _2287_ /*45394*/;
assign _2294_ = D[60] ^ Q[59] /*45390*/;
assign _2291_ = _1599_ & _2294_ /*45386*/;
assign _2292_ = _1599_ ^ _2294_ /*45389*/;
assign _2293_ = _2285_ & _2292_ /*45387*/;
assign _2290_ = _2291_ | _2293_ /*45385*/;
assign _1985_ = _2285_ ^ _2292_ /*45388*/;
assign _2299_ = D[61] ^ Q[59] /*45384*/;
assign _2296_ = _1600_ & _2299_ /*45380*/;
assign _2297_ = _1600_ ^ _2299_ /*45383*/;
assign _2298_ = _2290_ & _2297_ /*45381*/;
assign _2295_ = _2296_ | _2298_ /*45379*/;
assign _1986_ = _2290_ ^ _2297_ /*45382*/;
assign _2304_ = D[62] ^ Q[59] /*45378*/;
assign _2301_ = _1601_ & _2304_ /*45374*/;
assign _2302_ = _1601_ ^ _2304_ /*45377*/;
assign _2303_ = _2295_ & _2302_ /*45375*/;
assign _2300_ = _2301_ | _2303_ /*45373*/;
assign _1987_ = _2295_ ^ _2302_ /*45376*/;
assign _2308_ = zeroWire ^ Q[59] /*45372*/;
assign _2305_ = _1602_ & _2308_ /*45368*/;
assign _2306_ = _1602_ ^ _2308_ /*45371*/;
assign _2307_ = _2300_ & _2306_ /*45369*/;
assign Q[58] = _2305_ | _2307_ /*45367*/;
assign _1988_ = _2300_ ^ _2306_ /*45370*/;
assign _2379_ = D[0] ^ Q[58] /*44981*/;
assign _2376_ = R_0[57] & _2379_ /*44977*/;
assign _2377_ = R_0[57] ^ _2379_ /*44980*/;
assign _2378_ = Q[58] & _2377_ /*44978*/;
assign _2375_ = _2376_ | _2378_ /*44976*/;
assign _2310_ = Q[58] ^ _2377_ /*44979*/;
assign _2384_ = D[1] ^ Q[58] /*44975*/;
assign _2381_ = _1925_ & _2384_ /*44971*/;
assign _2382_ = _1925_ ^ _2384_ /*44974*/;
assign _2383_ = _2375_ & _2382_ /*44972*/;
assign _2380_ = _2381_ | _2383_ /*44970*/;
assign _2311_ = _2375_ ^ _2382_ /*44973*/;
assign _2389_ = D[2] ^ Q[58] /*44969*/;
assign _2386_ = _1926_ & _2389_ /*44965*/;
assign _2387_ = _1926_ ^ _2389_ /*44968*/;
assign _2388_ = _2380_ & _2387_ /*44966*/;
assign _2385_ = _2386_ | _2388_ /*44964*/;
assign _2312_ = _2380_ ^ _2387_ /*44967*/;
assign _2394_ = D[3] ^ Q[58] /*44963*/;
assign _2391_ = _1927_ & _2394_ /*44959*/;
assign _2392_ = _1927_ ^ _2394_ /*44962*/;
assign _2393_ = _2385_ & _2392_ /*44960*/;
assign _2390_ = _2391_ | _2393_ /*44958*/;
assign _2313_ = _2385_ ^ _2392_ /*44961*/;
assign _2399_ = D[4] ^ Q[58] /*44957*/;
assign _2396_ = _1928_ & _2399_ /*44953*/;
assign _2397_ = _1928_ ^ _2399_ /*44956*/;
assign _2398_ = _2390_ & _2397_ /*44954*/;
assign _2395_ = _2396_ | _2398_ /*44952*/;
assign _2314_ = _2390_ ^ _2397_ /*44955*/;
assign _2404_ = D[5] ^ Q[58] /*44951*/;
assign _2401_ = _1929_ & _2404_ /*44947*/;
assign _2402_ = _1929_ ^ _2404_ /*44950*/;
assign _2403_ = _2395_ & _2402_ /*44948*/;
assign _2400_ = _2401_ | _2403_ /*44946*/;
assign _2315_ = _2395_ ^ _2402_ /*44949*/;
assign _2409_ = D[6] ^ Q[58] /*44945*/;
assign _2406_ = _1930_ & _2409_ /*44941*/;
assign _2407_ = _1930_ ^ _2409_ /*44944*/;
assign _2408_ = _2400_ & _2407_ /*44942*/;
assign _2405_ = _2406_ | _2408_ /*44940*/;
assign _2316_ = _2400_ ^ _2407_ /*44943*/;
assign _2414_ = D[7] ^ Q[58] /*44939*/;
assign _2411_ = _1931_ & _2414_ /*44935*/;
assign _2412_ = _1931_ ^ _2414_ /*44938*/;
assign _2413_ = _2405_ & _2412_ /*44936*/;
assign _2410_ = _2411_ | _2413_ /*44934*/;
assign _2317_ = _2405_ ^ _2412_ /*44937*/;
assign _2419_ = D[8] ^ Q[58] /*44933*/;
assign _2416_ = _1932_ & _2419_ /*44929*/;
assign _2417_ = _1932_ ^ _2419_ /*44932*/;
assign _2418_ = _2410_ & _2417_ /*44930*/;
assign _2415_ = _2416_ | _2418_ /*44928*/;
assign _2318_ = _2410_ ^ _2417_ /*44931*/;
assign _2424_ = D[9] ^ Q[58] /*44927*/;
assign _2421_ = _1933_ & _2424_ /*44923*/;
assign _2422_ = _1933_ ^ _2424_ /*44926*/;
assign _2423_ = _2415_ & _2422_ /*44924*/;
assign _2420_ = _2421_ | _2423_ /*44922*/;
assign _2319_ = _2415_ ^ _2422_ /*44925*/;
assign _2429_ = D[10] ^ Q[58] /*44921*/;
assign _2426_ = _1934_ & _2429_ /*44917*/;
assign _2427_ = _1934_ ^ _2429_ /*44920*/;
assign _2428_ = _2420_ & _2427_ /*44918*/;
assign _2425_ = _2426_ | _2428_ /*44916*/;
assign _2320_ = _2420_ ^ _2427_ /*44919*/;
assign _2434_ = D[11] ^ Q[58] /*44915*/;
assign _2431_ = _1935_ & _2434_ /*44911*/;
assign _2432_ = _1935_ ^ _2434_ /*44914*/;
assign _2433_ = _2425_ & _2432_ /*44912*/;
assign _2430_ = _2431_ | _2433_ /*44910*/;
assign _2321_ = _2425_ ^ _2432_ /*44913*/;
assign _2439_ = D[12] ^ Q[58] /*44909*/;
assign _2436_ = _1936_ & _2439_ /*44905*/;
assign _2437_ = _1936_ ^ _2439_ /*44908*/;
assign _2438_ = _2430_ & _2437_ /*44906*/;
assign _2435_ = _2436_ | _2438_ /*44904*/;
assign _2322_ = _2430_ ^ _2437_ /*44907*/;
assign _2444_ = D[13] ^ Q[58] /*44903*/;
assign _2441_ = _1937_ & _2444_ /*44899*/;
assign _2442_ = _1937_ ^ _2444_ /*44902*/;
assign _2443_ = _2435_ & _2442_ /*44900*/;
assign _2440_ = _2441_ | _2443_ /*44898*/;
assign _2323_ = _2435_ ^ _2442_ /*44901*/;
assign _2449_ = D[14] ^ Q[58] /*44897*/;
assign _2446_ = _1938_ & _2449_ /*44893*/;
assign _2447_ = _1938_ ^ _2449_ /*44896*/;
assign _2448_ = _2440_ & _2447_ /*44894*/;
assign _2445_ = _2446_ | _2448_ /*44892*/;
assign _2324_ = _2440_ ^ _2447_ /*44895*/;
assign _2454_ = D[15] ^ Q[58] /*44891*/;
assign _2451_ = _1939_ & _2454_ /*44887*/;
assign _2452_ = _1939_ ^ _2454_ /*44890*/;
assign _2453_ = _2445_ & _2452_ /*44888*/;
assign _2450_ = _2451_ | _2453_ /*44886*/;
assign _2325_ = _2445_ ^ _2452_ /*44889*/;
assign _2459_ = D[16] ^ Q[58] /*44885*/;
assign _2456_ = _1940_ & _2459_ /*44881*/;
assign _2457_ = _1940_ ^ _2459_ /*44884*/;
assign _2458_ = _2450_ & _2457_ /*44882*/;
assign _2455_ = _2456_ | _2458_ /*44880*/;
assign _2326_ = _2450_ ^ _2457_ /*44883*/;
assign _2464_ = D[17] ^ Q[58] /*44879*/;
assign _2461_ = _1941_ & _2464_ /*44875*/;
assign _2462_ = _1941_ ^ _2464_ /*44878*/;
assign _2463_ = _2455_ & _2462_ /*44876*/;
assign _2460_ = _2461_ | _2463_ /*44874*/;
assign _2327_ = _2455_ ^ _2462_ /*44877*/;
assign _2469_ = D[18] ^ Q[58] /*44873*/;
assign _2466_ = _1942_ & _2469_ /*44869*/;
assign _2467_ = _1942_ ^ _2469_ /*44872*/;
assign _2468_ = _2460_ & _2467_ /*44870*/;
assign _2465_ = _2466_ | _2468_ /*44868*/;
assign _2328_ = _2460_ ^ _2467_ /*44871*/;
assign _2474_ = D[19] ^ Q[58] /*44867*/;
assign _2471_ = _1943_ & _2474_ /*44863*/;
assign _2472_ = _1943_ ^ _2474_ /*44866*/;
assign _2473_ = _2465_ & _2472_ /*44864*/;
assign _2470_ = _2471_ | _2473_ /*44862*/;
assign _2329_ = _2465_ ^ _2472_ /*44865*/;
assign _2479_ = D[20] ^ Q[58] /*44861*/;
assign _2476_ = _1944_ & _2479_ /*44857*/;
assign _2477_ = _1944_ ^ _2479_ /*44860*/;
assign _2478_ = _2470_ & _2477_ /*44858*/;
assign _2475_ = _2476_ | _2478_ /*44856*/;
assign _2330_ = _2470_ ^ _2477_ /*44859*/;
assign _2484_ = D[21] ^ Q[58] /*44855*/;
assign _2481_ = _1945_ & _2484_ /*44851*/;
assign _2482_ = _1945_ ^ _2484_ /*44854*/;
assign _2483_ = _2475_ & _2482_ /*44852*/;
assign _2480_ = _2481_ | _2483_ /*44850*/;
assign _2331_ = _2475_ ^ _2482_ /*44853*/;
assign _2489_ = D[22] ^ Q[58] /*44849*/;
assign _2486_ = _1946_ & _2489_ /*44845*/;
assign _2487_ = _1946_ ^ _2489_ /*44848*/;
assign _2488_ = _2480_ & _2487_ /*44846*/;
assign _2485_ = _2486_ | _2488_ /*44844*/;
assign _2332_ = _2480_ ^ _2487_ /*44847*/;
assign _2494_ = D[23] ^ Q[58] /*44843*/;
assign _2491_ = _1947_ & _2494_ /*44839*/;
assign _2492_ = _1947_ ^ _2494_ /*44842*/;
assign _2493_ = _2485_ & _2492_ /*44840*/;
assign _2490_ = _2491_ | _2493_ /*44838*/;
assign _2333_ = _2485_ ^ _2492_ /*44841*/;
assign _2499_ = D[24] ^ Q[58] /*44837*/;
assign _2496_ = _1948_ & _2499_ /*44833*/;
assign _2497_ = _1948_ ^ _2499_ /*44836*/;
assign _2498_ = _2490_ & _2497_ /*44834*/;
assign _2495_ = _2496_ | _2498_ /*44832*/;
assign _2334_ = _2490_ ^ _2497_ /*44835*/;
assign _2504_ = D[25] ^ Q[58] /*44831*/;
assign _2501_ = _1949_ & _2504_ /*44827*/;
assign _2502_ = _1949_ ^ _2504_ /*44830*/;
assign _2503_ = _2495_ & _2502_ /*44828*/;
assign _2500_ = _2501_ | _2503_ /*44826*/;
assign _2335_ = _2495_ ^ _2502_ /*44829*/;
assign _2509_ = D[26] ^ Q[58] /*44825*/;
assign _2506_ = _1950_ & _2509_ /*44821*/;
assign _2507_ = _1950_ ^ _2509_ /*44824*/;
assign _2508_ = _2500_ & _2507_ /*44822*/;
assign _2505_ = _2506_ | _2508_ /*44820*/;
assign _2336_ = _2500_ ^ _2507_ /*44823*/;
assign _2514_ = D[27] ^ Q[58] /*44819*/;
assign _2511_ = _1951_ & _2514_ /*44815*/;
assign _2512_ = _1951_ ^ _2514_ /*44818*/;
assign _2513_ = _2505_ & _2512_ /*44816*/;
assign _2510_ = _2511_ | _2513_ /*44814*/;
assign _2337_ = _2505_ ^ _2512_ /*44817*/;
assign _2519_ = D[28] ^ Q[58] /*44813*/;
assign _2516_ = _1952_ & _2519_ /*44809*/;
assign _2517_ = _1952_ ^ _2519_ /*44812*/;
assign _2518_ = _2510_ & _2517_ /*44810*/;
assign _2515_ = _2516_ | _2518_ /*44808*/;
assign _2338_ = _2510_ ^ _2517_ /*44811*/;
assign _2524_ = D[29] ^ Q[58] /*44807*/;
assign _2521_ = _1953_ & _2524_ /*44803*/;
assign _2522_ = _1953_ ^ _2524_ /*44806*/;
assign _2523_ = _2515_ & _2522_ /*44804*/;
assign _2520_ = _2521_ | _2523_ /*44802*/;
assign _2339_ = _2515_ ^ _2522_ /*44805*/;
assign _2529_ = D[30] ^ Q[58] /*44801*/;
assign _2526_ = _1954_ & _2529_ /*44797*/;
assign _2527_ = _1954_ ^ _2529_ /*44800*/;
assign _2528_ = _2520_ & _2527_ /*44798*/;
assign _2525_ = _2526_ | _2528_ /*44796*/;
assign _2340_ = _2520_ ^ _2527_ /*44799*/;
assign _2534_ = D[31] ^ Q[58] /*44795*/;
assign _2531_ = _1955_ & _2534_ /*44791*/;
assign _2532_ = _1955_ ^ _2534_ /*44794*/;
assign _2533_ = _2525_ & _2532_ /*44792*/;
assign _2530_ = _2531_ | _2533_ /*44790*/;
assign _2341_ = _2525_ ^ _2532_ /*44793*/;
assign _2539_ = D[32] ^ Q[58] /*44789*/;
assign _2536_ = _1956_ & _2539_ /*44785*/;
assign _2537_ = _1956_ ^ _2539_ /*44788*/;
assign _2538_ = _2530_ & _2537_ /*44786*/;
assign _2535_ = _2536_ | _2538_ /*44784*/;
assign _2342_ = _2530_ ^ _2537_ /*44787*/;
assign _2544_ = D[33] ^ Q[58] /*44783*/;
assign _2541_ = _1957_ & _2544_ /*44779*/;
assign _2542_ = _1957_ ^ _2544_ /*44782*/;
assign _2543_ = _2535_ & _2542_ /*44780*/;
assign _2540_ = _2541_ | _2543_ /*44778*/;
assign _2343_ = _2535_ ^ _2542_ /*44781*/;
assign _2549_ = D[34] ^ Q[58] /*44777*/;
assign _2546_ = _1958_ & _2549_ /*44773*/;
assign _2547_ = _1958_ ^ _2549_ /*44776*/;
assign _2548_ = _2540_ & _2547_ /*44774*/;
assign _2545_ = _2546_ | _2548_ /*44772*/;
assign _2344_ = _2540_ ^ _2547_ /*44775*/;
assign _2554_ = D[35] ^ Q[58] /*44771*/;
assign _2551_ = _1959_ & _2554_ /*44767*/;
assign _2552_ = _1959_ ^ _2554_ /*44770*/;
assign _2553_ = _2545_ & _2552_ /*44768*/;
assign _2550_ = _2551_ | _2553_ /*44766*/;
assign _2345_ = _2545_ ^ _2552_ /*44769*/;
assign _2559_ = D[36] ^ Q[58] /*44765*/;
assign _2556_ = _1960_ & _2559_ /*44761*/;
assign _2557_ = _1960_ ^ _2559_ /*44764*/;
assign _2558_ = _2550_ & _2557_ /*44762*/;
assign _2555_ = _2556_ | _2558_ /*44760*/;
assign _2346_ = _2550_ ^ _2557_ /*44763*/;
assign _2564_ = D[37] ^ Q[58] /*44759*/;
assign _2561_ = _1961_ & _2564_ /*44755*/;
assign _2562_ = _1961_ ^ _2564_ /*44758*/;
assign _2563_ = _2555_ & _2562_ /*44756*/;
assign _2560_ = _2561_ | _2563_ /*44754*/;
assign _2347_ = _2555_ ^ _2562_ /*44757*/;
assign _2569_ = D[38] ^ Q[58] /*44753*/;
assign _2566_ = _1962_ & _2569_ /*44749*/;
assign _2567_ = _1962_ ^ _2569_ /*44752*/;
assign _2568_ = _2560_ & _2567_ /*44750*/;
assign _2565_ = _2566_ | _2568_ /*44748*/;
assign _2348_ = _2560_ ^ _2567_ /*44751*/;
assign _2574_ = D[39] ^ Q[58] /*44747*/;
assign _2571_ = _1963_ & _2574_ /*44743*/;
assign _2572_ = _1963_ ^ _2574_ /*44746*/;
assign _2573_ = _2565_ & _2572_ /*44744*/;
assign _2570_ = _2571_ | _2573_ /*44742*/;
assign _2349_ = _2565_ ^ _2572_ /*44745*/;
assign _2579_ = D[40] ^ Q[58] /*44741*/;
assign _2576_ = _1964_ & _2579_ /*44737*/;
assign _2577_ = _1964_ ^ _2579_ /*44740*/;
assign _2578_ = _2570_ & _2577_ /*44738*/;
assign _2575_ = _2576_ | _2578_ /*44736*/;
assign _2350_ = _2570_ ^ _2577_ /*44739*/;
assign _2584_ = D[41] ^ Q[58] /*44735*/;
assign _2581_ = _1965_ & _2584_ /*44731*/;
assign _2582_ = _1965_ ^ _2584_ /*44734*/;
assign _2583_ = _2575_ & _2582_ /*44732*/;
assign _2580_ = _2581_ | _2583_ /*44730*/;
assign _2351_ = _2575_ ^ _2582_ /*44733*/;
assign _2589_ = D[42] ^ Q[58] /*44729*/;
assign _2586_ = _1966_ & _2589_ /*44725*/;
assign _2587_ = _1966_ ^ _2589_ /*44728*/;
assign _2588_ = _2580_ & _2587_ /*44726*/;
assign _2585_ = _2586_ | _2588_ /*44724*/;
assign _2352_ = _2580_ ^ _2587_ /*44727*/;
assign _2594_ = D[43] ^ Q[58] /*44723*/;
assign _2591_ = _1967_ & _2594_ /*44719*/;
assign _2592_ = _1967_ ^ _2594_ /*44722*/;
assign _2593_ = _2585_ & _2592_ /*44720*/;
assign _2590_ = _2591_ | _2593_ /*44718*/;
assign _2353_ = _2585_ ^ _2592_ /*44721*/;
assign _2599_ = D[44] ^ Q[58] /*44717*/;
assign _2596_ = _1968_ & _2599_ /*44713*/;
assign _2597_ = _1968_ ^ _2599_ /*44716*/;
assign _2598_ = _2590_ & _2597_ /*44714*/;
assign _2595_ = _2596_ | _2598_ /*44712*/;
assign _2354_ = _2590_ ^ _2597_ /*44715*/;
assign _2604_ = D[45] ^ Q[58] /*44711*/;
assign _2601_ = _1969_ & _2604_ /*44707*/;
assign _2602_ = _1969_ ^ _2604_ /*44710*/;
assign _2603_ = _2595_ & _2602_ /*44708*/;
assign _2600_ = _2601_ | _2603_ /*44706*/;
assign _2355_ = _2595_ ^ _2602_ /*44709*/;
assign _2609_ = D[46] ^ Q[58] /*44705*/;
assign _2606_ = _1970_ & _2609_ /*44701*/;
assign _2607_ = _1970_ ^ _2609_ /*44704*/;
assign _2608_ = _2600_ & _2607_ /*44702*/;
assign _2605_ = _2606_ | _2608_ /*44700*/;
assign _2356_ = _2600_ ^ _2607_ /*44703*/;
assign _2614_ = D[47] ^ Q[58] /*44699*/;
assign _2611_ = _1971_ & _2614_ /*44695*/;
assign _2612_ = _1971_ ^ _2614_ /*44698*/;
assign _2613_ = _2605_ & _2612_ /*44696*/;
assign _2610_ = _2611_ | _2613_ /*44694*/;
assign _2357_ = _2605_ ^ _2612_ /*44697*/;
assign _2619_ = D[48] ^ Q[58] /*44693*/;
assign _2616_ = _1972_ & _2619_ /*44689*/;
assign _2617_ = _1972_ ^ _2619_ /*44692*/;
assign _2618_ = _2610_ & _2617_ /*44690*/;
assign _2615_ = _2616_ | _2618_ /*44688*/;
assign _2358_ = _2610_ ^ _2617_ /*44691*/;
assign _2624_ = D[49] ^ Q[58] /*44687*/;
assign _2621_ = _1973_ & _2624_ /*44683*/;
assign _2622_ = _1973_ ^ _2624_ /*44686*/;
assign _2623_ = _2615_ & _2622_ /*44684*/;
assign _2620_ = _2621_ | _2623_ /*44682*/;
assign _2359_ = _2615_ ^ _2622_ /*44685*/;
assign _2629_ = D[50] ^ Q[58] /*44681*/;
assign _2626_ = _1974_ & _2629_ /*44677*/;
assign _2627_ = _1974_ ^ _2629_ /*44680*/;
assign _2628_ = _2620_ & _2627_ /*44678*/;
assign _2625_ = _2626_ | _2628_ /*44676*/;
assign _2360_ = _2620_ ^ _2627_ /*44679*/;
assign _2634_ = D[51] ^ Q[58] /*44675*/;
assign _2631_ = _1975_ & _2634_ /*44671*/;
assign _2632_ = _1975_ ^ _2634_ /*44674*/;
assign _2633_ = _2625_ & _2632_ /*44672*/;
assign _2630_ = _2631_ | _2633_ /*44670*/;
assign _2361_ = _2625_ ^ _2632_ /*44673*/;
assign _2639_ = D[52] ^ Q[58] /*44669*/;
assign _2636_ = _1976_ & _2639_ /*44665*/;
assign _2637_ = _1976_ ^ _2639_ /*44668*/;
assign _2638_ = _2630_ & _2637_ /*44666*/;
assign _2635_ = _2636_ | _2638_ /*44664*/;
assign _2362_ = _2630_ ^ _2637_ /*44667*/;
assign _2644_ = D[53] ^ Q[58] /*44663*/;
assign _2641_ = _1977_ & _2644_ /*44659*/;
assign _2642_ = _1977_ ^ _2644_ /*44662*/;
assign _2643_ = _2635_ & _2642_ /*44660*/;
assign _2640_ = _2641_ | _2643_ /*44658*/;
assign _2363_ = _2635_ ^ _2642_ /*44661*/;
assign _2649_ = D[54] ^ Q[58] /*44657*/;
assign _2646_ = _1978_ & _2649_ /*44653*/;
assign _2647_ = _1978_ ^ _2649_ /*44656*/;
assign _2648_ = _2640_ & _2647_ /*44654*/;
assign _2645_ = _2646_ | _2648_ /*44652*/;
assign _2364_ = _2640_ ^ _2647_ /*44655*/;
assign _2654_ = D[55] ^ Q[58] /*44651*/;
assign _2651_ = _1979_ & _2654_ /*44647*/;
assign _2652_ = _1979_ ^ _2654_ /*44650*/;
assign _2653_ = _2645_ & _2652_ /*44648*/;
assign _2650_ = _2651_ | _2653_ /*44646*/;
assign _2365_ = _2645_ ^ _2652_ /*44649*/;
assign _2659_ = D[56] ^ Q[58] /*44645*/;
assign _2656_ = _1980_ & _2659_ /*44641*/;
assign _2657_ = _1980_ ^ _2659_ /*44644*/;
assign _2658_ = _2650_ & _2657_ /*44642*/;
assign _2655_ = _2656_ | _2658_ /*44640*/;
assign _2366_ = _2650_ ^ _2657_ /*44643*/;
assign _2664_ = D[57] ^ Q[58] /*44639*/;
assign _2661_ = _1981_ & _2664_ /*44635*/;
assign _2662_ = _1981_ ^ _2664_ /*44638*/;
assign _2663_ = _2655_ & _2662_ /*44636*/;
assign _2660_ = _2661_ | _2663_ /*44634*/;
assign _2367_ = _2655_ ^ _2662_ /*44637*/;
assign _2669_ = D[58] ^ Q[58] /*44633*/;
assign _2666_ = _1982_ & _2669_ /*44629*/;
assign _2667_ = _1982_ ^ _2669_ /*44632*/;
assign _2668_ = _2660_ & _2667_ /*44630*/;
assign _2665_ = _2666_ | _2668_ /*44628*/;
assign _2368_ = _2660_ ^ _2667_ /*44631*/;
assign _2674_ = D[59] ^ Q[58] /*44627*/;
assign _2671_ = _1983_ & _2674_ /*44623*/;
assign _2672_ = _1983_ ^ _2674_ /*44626*/;
assign _2673_ = _2665_ & _2672_ /*44624*/;
assign _2670_ = _2671_ | _2673_ /*44622*/;
assign _2369_ = _2665_ ^ _2672_ /*44625*/;
assign _2679_ = D[60] ^ Q[58] /*44621*/;
assign _2676_ = _1984_ & _2679_ /*44617*/;
assign _2677_ = _1984_ ^ _2679_ /*44620*/;
assign _2678_ = _2670_ & _2677_ /*44618*/;
assign _2675_ = _2676_ | _2678_ /*44616*/;
assign _2370_ = _2670_ ^ _2677_ /*44619*/;
assign _2684_ = D[61] ^ Q[58] /*44615*/;
assign _2681_ = _1985_ & _2684_ /*44611*/;
assign _2682_ = _1985_ ^ _2684_ /*44614*/;
assign _2683_ = _2675_ & _2682_ /*44612*/;
assign _2680_ = _2681_ | _2683_ /*44610*/;
assign _2371_ = _2675_ ^ _2682_ /*44613*/;
assign _2689_ = D[62] ^ Q[58] /*44609*/;
assign _2686_ = _1986_ & _2689_ /*44605*/;
assign _2687_ = _1986_ ^ _2689_ /*44608*/;
assign _2688_ = _2680_ & _2687_ /*44606*/;
assign _2685_ = _2686_ | _2688_ /*44604*/;
assign _2372_ = _2680_ ^ _2687_ /*44607*/;
assign _2693_ = zeroWire ^ Q[58] /*44603*/;
assign _2690_ = _1987_ & _2693_ /*44599*/;
assign _2691_ = _1987_ ^ _2693_ /*44602*/;
assign _2692_ = _2685_ & _2691_ /*44600*/;
assign Q[57] = _2690_ | _2692_ /*44598*/;
assign _2373_ = _2685_ ^ _2691_ /*44601*/;
assign _2764_ = D[0] ^ Q[57] /*44212*/;
assign _2761_ = R_0[56] & _2764_ /*44208*/;
assign _2762_ = R_0[56] ^ _2764_ /*44211*/;
assign _2763_ = Q[57] & _2762_ /*44209*/;
assign _2760_ = _2761_ | _2763_ /*44207*/;
assign _2695_ = Q[57] ^ _2762_ /*44210*/;
assign _2769_ = D[1] ^ Q[57] /*44206*/;
assign _2766_ = _2310_ & _2769_ /*44202*/;
assign _2767_ = _2310_ ^ _2769_ /*44205*/;
assign _2768_ = _2760_ & _2767_ /*44203*/;
assign _2765_ = _2766_ | _2768_ /*44201*/;
assign _2696_ = _2760_ ^ _2767_ /*44204*/;
assign _2774_ = D[2] ^ Q[57] /*44200*/;
assign _2771_ = _2311_ & _2774_ /*44196*/;
assign _2772_ = _2311_ ^ _2774_ /*44199*/;
assign _2773_ = _2765_ & _2772_ /*44197*/;
assign _2770_ = _2771_ | _2773_ /*44195*/;
assign _2697_ = _2765_ ^ _2772_ /*44198*/;
assign _2779_ = D[3] ^ Q[57] /*44194*/;
assign _2776_ = _2312_ & _2779_ /*44190*/;
assign _2777_ = _2312_ ^ _2779_ /*44193*/;
assign _2778_ = _2770_ & _2777_ /*44191*/;
assign _2775_ = _2776_ | _2778_ /*44189*/;
assign _2698_ = _2770_ ^ _2777_ /*44192*/;
assign _2784_ = D[4] ^ Q[57] /*44188*/;
assign _2781_ = _2313_ & _2784_ /*44184*/;
assign _2782_ = _2313_ ^ _2784_ /*44187*/;
assign _2783_ = _2775_ & _2782_ /*44185*/;
assign _2780_ = _2781_ | _2783_ /*44183*/;
assign _2699_ = _2775_ ^ _2782_ /*44186*/;
assign _2789_ = D[5] ^ Q[57] /*44182*/;
assign _2786_ = _2314_ & _2789_ /*44178*/;
assign _2787_ = _2314_ ^ _2789_ /*44181*/;
assign _2788_ = _2780_ & _2787_ /*44179*/;
assign _2785_ = _2786_ | _2788_ /*44177*/;
assign _2700_ = _2780_ ^ _2787_ /*44180*/;
assign _2794_ = D[6] ^ Q[57] /*44176*/;
assign _2791_ = _2315_ & _2794_ /*44172*/;
assign _2792_ = _2315_ ^ _2794_ /*44175*/;
assign _2793_ = _2785_ & _2792_ /*44173*/;
assign _2790_ = _2791_ | _2793_ /*44171*/;
assign _2701_ = _2785_ ^ _2792_ /*44174*/;
assign _2799_ = D[7] ^ Q[57] /*44170*/;
assign _2796_ = _2316_ & _2799_ /*44166*/;
assign _2797_ = _2316_ ^ _2799_ /*44169*/;
assign _2798_ = _2790_ & _2797_ /*44167*/;
assign _2795_ = _2796_ | _2798_ /*44165*/;
assign _2702_ = _2790_ ^ _2797_ /*44168*/;
assign _2804_ = D[8] ^ Q[57] /*44164*/;
assign _2801_ = _2317_ & _2804_ /*44160*/;
assign _2802_ = _2317_ ^ _2804_ /*44163*/;
assign _2803_ = _2795_ & _2802_ /*44161*/;
assign _2800_ = _2801_ | _2803_ /*44159*/;
assign _2703_ = _2795_ ^ _2802_ /*44162*/;
assign _2809_ = D[9] ^ Q[57] /*44158*/;
assign _2806_ = _2318_ & _2809_ /*44154*/;
assign _2807_ = _2318_ ^ _2809_ /*44157*/;
assign _2808_ = _2800_ & _2807_ /*44155*/;
assign _2805_ = _2806_ | _2808_ /*44153*/;
assign _2704_ = _2800_ ^ _2807_ /*44156*/;
assign _2814_ = D[10] ^ Q[57] /*44152*/;
assign _2811_ = _2319_ & _2814_ /*44148*/;
assign _2812_ = _2319_ ^ _2814_ /*44151*/;
assign _2813_ = _2805_ & _2812_ /*44149*/;
assign _2810_ = _2811_ | _2813_ /*44147*/;
assign _2705_ = _2805_ ^ _2812_ /*44150*/;
assign _2819_ = D[11] ^ Q[57] /*44146*/;
assign _2816_ = _2320_ & _2819_ /*44142*/;
assign _2817_ = _2320_ ^ _2819_ /*44145*/;
assign _2818_ = _2810_ & _2817_ /*44143*/;
assign _2815_ = _2816_ | _2818_ /*44141*/;
assign _2706_ = _2810_ ^ _2817_ /*44144*/;
assign _2824_ = D[12] ^ Q[57] /*44140*/;
assign _2821_ = _2321_ & _2824_ /*44136*/;
assign _2822_ = _2321_ ^ _2824_ /*44139*/;
assign _2823_ = _2815_ & _2822_ /*44137*/;
assign _2820_ = _2821_ | _2823_ /*44135*/;
assign _2707_ = _2815_ ^ _2822_ /*44138*/;
assign _2829_ = D[13] ^ Q[57] /*44134*/;
assign _2826_ = _2322_ & _2829_ /*44130*/;
assign _2827_ = _2322_ ^ _2829_ /*44133*/;
assign _2828_ = _2820_ & _2827_ /*44131*/;
assign _2825_ = _2826_ | _2828_ /*44129*/;
assign _2708_ = _2820_ ^ _2827_ /*44132*/;
assign _2834_ = D[14] ^ Q[57] /*44128*/;
assign _2831_ = _2323_ & _2834_ /*44124*/;
assign _2832_ = _2323_ ^ _2834_ /*44127*/;
assign _2833_ = _2825_ & _2832_ /*44125*/;
assign _2830_ = _2831_ | _2833_ /*44123*/;
assign _2709_ = _2825_ ^ _2832_ /*44126*/;
assign _2839_ = D[15] ^ Q[57] /*44122*/;
assign _2836_ = _2324_ & _2839_ /*44118*/;
assign _2837_ = _2324_ ^ _2839_ /*44121*/;
assign _2838_ = _2830_ & _2837_ /*44119*/;
assign _2835_ = _2836_ | _2838_ /*44117*/;
assign _2710_ = _2830_ ^ _2837_ /*44120*/;
assign _2844_ = D[16] ^ Q[57] /*44116*/;
assign _2841_ = _2325_ & _2844_ /*44112*/;
assign _2842_ = _2325_ ^ _2844_ /*44115*/;
assign _2843_ = _2835_ & _2842_ /*44113*/;
assign _2840_ = _2841_ | _2843_ /*44111*/;
assign _2711_ = _2835_ ^ _2842_ /*44114*/;
assign _2849_ = D[17] ^ Q[57] /*44110*/;
assign _2846_ = _2326_ & _2849_ /*44106*/;
assign _2847_ = _2326_ ^ _2849_ /*44109*/;
assign _2848_ = _2840_ & _2847_ /*44107*/;
assign _2845_ = _2846_ | _2848_ /*44105*/;
assign _2712_ = _2840_ ^ _2847_ /*44108*/;
assign _2854_ = D[18] ^ Q[57] /*44104*/;
assign _2851_ = _2327_ & _2854_ /*44100*/;
assign _2852_ = _2327_ ^ _2854_ /*44103*/;
assign _2853_ = _2845_ & _2852_ /*44101*/;
assign _2850_ = _2851_ | _2853_ /*44099*/;
assign _2713_ = _2845_ ^ _2852_ /*44102*/;
assign _2859_ = D[19] ^ Q[57] /*44098*/;
assign _2856_ = _2328_ & _2859_ /*44094*/;
assign _2857_ = _2328_ ^ _2859_ /*44097*/;
assign _2858_ = _2850_ & _2857_ /*44095*/;
assign _2855_ = _2856_ | _2858_ /*44093*/;
assign _2714_ = _2850_ ^ _2857_ /*44096*/;
assign _2864_ = D[20] ^ Q[57] /*44092*/;
assign _2861_ = _2329_ & _2864_ /*44088*/;
assign _2862_ = _2329_ ^ _2864_ /*44091*/;
assign _2863_ = _2855_ & _2862_ /*44089*/;
assign _2860_ = _2861_ | _2863_ /*44087*/;
assign _2715_ = _2855_ ^ _2862_ /*44090*/;
assign _2869_ = D[21] ^ Q[57] /*44086*/;
assign _2866_ = _2330_ & _2869_ /*44082*/;
assign _2867_ = _2330_ ^ _2869_ /*44085*/;
assign _2868_ = _2860_ & _2867_ /*44083*/;
assign _2865_ = _2866_ | _2868_ /*44081*/;
assign _2716_ = _2860_ ^ _2867_ /*44084*/;
assign _2874_ = D[22] ^ Q[57] /*44080*/;
assign _2871_ = _2331_ & _2874_ /*44076*/;
assign _2872_ = _2331_ ^ _2874_ /*44079*/;
assign _2873_ = _2865_ & _2872_ /*44077*/;
assign _2870_ = _2871_ | _2873_ /*44075*/;
assign _2717_ = _2865_ ^ _2872_ /*44078*/;
assign _2879_ = D[23] ^ Q[57] /*44074*/;
assign _2876_ = _2332_ & _2879_ /*44070*/;
assign _2877_ = _2332_ ^ _2879_ /*44073*/;
assign _2878_ = _2870_ & _2877_ /*44071*/;
assign _2875_ = _2876_ | _2878_ /*44069*/;
assign _2718_ = _2870_ ^ _2877_ /*44072*/;
assign _2884_ = D[24] ^ Q[57] /*44068*/;
assign _2881_ = _2333_ & _2884_ /*44064*/;
assign _2882_ = _2333_ ^ _2884_ /*44067*/;
assign _2883_ = _2875_ & _2882_ /*44065*/;
assign _2880_ = _2881_ | _2883_ /*44063*/;
assign _2719_ = _2875_ ^ _2882_ /*44066*/;
assign _2889_ = D[25] ^ Q[57] /*44062*/;
assign _2886_ = _2334_ & _2889_ /*44058*/;
assign _2887_ = _2334_ ^ _2889_ /*44061*/;
assign _2888_ = _2880_ & _2887_ /*44059*/;
assign _2885_ = _2886_ | _2888_ /*44057*/;
assign _2720_ = _2880_ ^ _2887_ /*44060*/;
assign _2894_ = D[26] ^ Q[57] /*44056*/;
assign _2891_ = _2335_ & _2894_ /*44052*/;
assign _2892_ = _2335_ ^ _2894_ /*44055*/;
assign _2893_ = _2885_ & _2892_ /*44053*/;
assign _2890_ = _2891_ | _2893_ /*44051*/;
assign _2721_ = _2885_ ^ _2892_ /*44054*/;
assign _2899_ = D[27] ^ Q[57] /*44050*/;
assign _2896_ = _2336_ & _2899_ /*44046*/;
assign _2897_ = _2336_ ^ _2899_ /*44049*/;
assign _2898_ = _2890_ & _2897_ /*44047*/;
assign _2895_ = _2896_ | _2898_ /*44045*/;
assign _2722_ = _2890_ ^ _2897_ /*44048*/;
assign _2904_ = D[28] ^ Q[57] /*44044*/;
assign _2901_ = _2337_ & _2904_ /*44040*/;
assign _2902_ = _2337_ ^ _2904_ /*44043*/;
assign _2903_ = _2895_ & _2902_ /*44041*/;
assign _2900_ = _2901_ | _2903_ /*44039*/;
assign _2723_ = _2895_ ^ _2902_ /*44042*/;
assign _2909_ = D[29] ^ Q[57] /*44038*/;
assign _2906_ = _2338_ & _2909_ /*44034*/;
assign _2907_ = _2338_ ^ _2909_ /*44037*/;
assign _2908_ = _2900_ & _2907_ /*44035*/;
assign _2905_ = _2906_ | _2908_ /*44033*/;
assign _2724_ = _2900_ ^ _2907_ /*44036*/;
assign _2914_ = D[30] ^ Q[57] /*44032*/;
assign _2911_ = _2339_ & _2914_ /*44028*/;
assign _2912_ = _2339_ ^ _2914_ /*44031*/;
assign _2913_ = _2905_ & _2912_ /*44029*/;
assign _2910_ = _2911_ | _2913_ /*44027*/;
assign _2725_ = _2905_ ^ _2912_ /*44030*/;
assign _2919_ = D[31] ^ Q[57] /*44026*/;
assign _2916_ = _2340_ & _2919_ /*44022*/;
assign _2917_ = _2340_ ^ _2919_ /*44025*/;
assign _2918_ = _2910_ & _2917_ /*44023*/;
assign _2915_ = _2916_ | _2918_ /*44021*/;
assign _2726_ = _2910_ ^ _2917_ /*44024*/;
assign _2924_ = D[32] ^ Q[57] /*44020*/;
assign _2921_ = _2341_ & _2924_ /*44016*/;
assign _2922_ = _2341_ ^ _2924_ /*44019*/;
assign _2923_ = _2915_ & _2922_ /*44017*/;
assign _2920_ = _2921_ | _2923_ /*44015*/;
assign _2727_ = _2915_ ^ _2922_ /*44018*/;
assign _2929_ = D[33] ^ Q[57] /*44014*/;
assign _2926_ = _2342_ & _2929_ /*44010*/;
assign _2927_ = _2342_ ^ _2929_ /*44013*/;
assign _2928_ = _2920_ & _2927_ /*44011*/;
assign _2925_ = _2926_ | _2928_ /*44009*/;
assign _2728_ = _2920_ ^ _2927_ /*44012*/;
assign _2934_ = D[34] ^ Q[57] /*44008*/;
assign _2931_ = _2343_ & _2934_ /*44004*/;
assign _2932_ = _2343_ ^ _2934_ /*44007*/;
assign _2933_ = _2925_ & _2932_ /*44005*/;
assign _2930_ = _2931_ | _2933_ /*44003*/;
assign _2729_ = _2925_ ^ _2932_ /*44006*/;
assign _2939_ = D[35] ^ Q[57] /*44002*/;
assign _2936_ = _2344_ & _2939_ /*43998*/;
assign _2937_ = _2344_ ^ _2939_ /*44001*/;
assign _2938_ = _2930_ & _2937_ /*43999*/;
assign _2935_ = _2936_ | _2938_ /*43997*/;
assign _2730_ = _2930_ ^ _2937_ /*44000*/;
assign _2944_ = D[36] ^ Q[57] /*43996*/;
assign _2941_ = _2345_ & _2944_ /*43992*/;
assign _2942_ = _2345_ ^ _2944_ /*43995*/;
assign _2943_ = _2935_ & _2942_ /*43993*/;
assign _2940_ = _2941_ | _2943_ /*43991*/;
assign _2731_ = _2935_ ^ _2942_ /*43994*/;
assign _2949_ = D[37] ^ Q[57] /*43990*/;
assign _2946_ = _2346_ & _2949_ /*43986*/;
assign _2947_ = _2346_ ^ _2949_ /*43989*/;
assign _2948_ = _2940_ & _2947_ /*43987*/;
assign _2945_ = _2946_ | _2948_ /*43985*/;
assign _2732_ = _2940_ ^ _2947_ /*43988*/;
assign _2954_ = D[38] ^ Q[57] /*43984*/;
assign _2951_ = _2347_ & _2954_ /*43980*/;
assign _2952_ = _2347_ ^ _2954_ /*43983*/;
assign _2953_ = _2945_ & _2952_ /*43981*/;
assign _2950_ = _2951_ | _2953_ /*43979*/;
assign _2733_ = _2945_ ^ _2952_ /*43982*/;
assign _2959_ = D[39] ^ Q[57] /*43978*/;
assign _2956_ = _2348_ & _2959_ /*43974*/;
assign _2957_ = _2348_ ^ _2959_ /*43977*/;
assign _2958_ = _2950_ & _2957_ /*43975*/;
assign _2955_ = _2956_ | _2958_ /*43973*/;
assign _2734_ = _2950_ ^ _2957_ /*43976*/;
assign _2964_ = D[40] ^ Q[57] /*43972*/;
assign _2961_ = _2349_ & _2964_ /*43968*/;
assign _2962_ = _2349_ ^ _2964_ /*43971*/;
assign _2963_ = _2955_ & _2962_ /*43969*/;
assign _2960_ = _2961_ | _2963_ /*43967*/;
assign _2735_ = _2955_ ^ _2962_ /*43970*/;
assign _2969_ = D[41] ^ Q[57] /*43966*/;
assign _2966_ = _2350_ & _2969_ /*43962*/;
assign _2967_ = _2350_ ^ _2969_ /*43965*/;
assign _2968_ = _2960_ & _2967_ /*43963*/;
assign _2965_ = _2966_ | _2968_ /*43961*/;
assign _2736_ = _2960_ ^ _2967_ /*43964*/;
assign _2974_ = D[42] ^ Q[57] /*43960*/;
assign _2971_ = _2351_ & _2974_ /*43956*/;
assign _2972_ = _2351_ ^ _2974_ /*43959*/;
assign _2973_ = _2965_ & _2972_ /*43957*/;
assign _2970_ = _2971_ | _2973_ /*43955*/;
assign _2737_ = _2965_ ^ _2972_ /*43958*/;
assign _2979_ = D[43] ^ Q[57] /*43954*/;
assign _2976_ = _2352_ & _2979_ /*43950*/;
assign _2977_ = _2352_ ^ _2979_ /*43953*/;
assign _2978_ = _2970_ & _2977_ /*43951*/;
assign _2975_ = _2976_ | _2978_ /*43949*/;
assign _2738_ = _2970_ ^ _2977_ /*43952*/;
assign _2984_ = D[44] ^ Q[57] /*43948*/;
assign _2981_ = _2353_ & _2984_ /*43944*/;
assign _2982_ = _2353_ ^ _2984_ /*43947*/;
assign _2983_ = _2975_ & _2982_ /*43945*/;
assign _2980_ = _2981_ | _2983_ /*43943*/;
assign _2739_ = _2975_ ^ _2982_ /*43946*/;
assign _2989_ = D[45] ^ Q[57] /*43942*/;
assign _2986_ = _2354_ & _2989_ /*43938*/;
assign _2987_ = _2354_ ^ _2989_ /*43941*/;
assign _2988_ = _2980_ & _2987_ /*43939*/;
assign _2985_ = _2986_ | _2988_ /*43937*/;
assign _2740_ = _2980_ ^ _2987_ /*43940*/;
assign _2994_ = D[46] ^ Q[57] /*43936*/;
assign _2991_ = _2355_ & _2994_ /*43932*/;
assign _2992_ = _2355_ ^ _2994_ /*43935*/;
assign _2993_ = _2985_ & _2992_ /*43933*/;
assign _2990_ = _2991_ | _2993_ /*43931*/;
assign _2741_ = _2985_ ^ _2992_ /*43934*/;
assign _2999_ = D[47] ^ Q[57] /*43930*/;
assign _2996_ = _2356_ & _2999_ /*43926*/;
assign _2997_ = _2356_ ^ _2999_ /*43929*/;
assign _2998_ = _2990_ & _2997_ /*43927*/;
assign _2995_ = _2996_ | _2998_ /*43925*/;
assign _2742_ = _2990_ ^ _2997_ /*43928*/;
assign _3004_ = D[48] ^ Q[57] /*43924*/;
assign _3001_ = _2357_ & _3004_ /*43920*/;
assign _3002_ = _2357_ ^ _3004_ /*43923*/;
assign _3003_ = _2995_ & _3002_ /*43921*/;
assign _3000_ = _3001_ | _3003_ /*43919*/;
assign _2743_ = _2995_ ^ _3002_ /*43922*/;
assign _3009_ = D[49] ^ Q[57] /*43918*/;
assign _3006_ = _2358_ & _3009_ /*43914*/;
assign _3007_ = _2358_ ^ _3009_ /*43917*/;
assign _3008_ = _3000_ & _3007_ /*43915*/;
assign _3005_ = _3006_ | _3008_ /*43913*/;
assign _2744_ = _3000_ ^ _3007_ /*43916*/;
assign _3014_ = D[50] ^ Q[57] /*43912*/;
assign _3011_ = _2359_ & _3014_ /*43908*/;
assign _3012_ = _2359_ ^ _3014_ /*43911*/;
assign _3013_ = _3005_ & _3012_ /*43909*/;
assign _3010_ = _3011_ | _3013_ /*43907*/;
assign _2745_ = _3005_ ^ _3012_ /*43910*/;
assign _3019_ = D[51] ^ Q[57] /*43906*/;
assign _3016_ = _2360_ & _3019_ /*43902*/;
assign _3017_ = _2360_ ^ _3019_ /*43905*/;
assign _3018_ = _3010_ & _3017_ /*43903*/;
assign _3015_ = _3016_ | _3018_ /*43901*/;
assign _2746_ = _3010_ ^ _3017_ /*43904*/;
assign _3024_ = D[52] ^ Q[57] /*43900*/;
assign _3021_ = _2361_ & _3024_ /*43896*/;
assign _3022_ = _2361_ ^ _3024_ /*43899*/;
assign _3023_ = _3015_ & _3022_ /*43897*/;
assign _3020_ = _3021_ | _3023_ /*43895*/;
assign _2747_ = _3015_ ^ _3022_ /*43898*/;
assign _3029_ = D[53] ^ Q[57] /*43894*/;
assign _3026_ = _2362_ & _3029_ /*43890*/;
assign _3027_ = _2362_ ^ _3029_ /*43893*/;
assign _3028_ = _3020_ & _3027_ /*43891*/;
assign _3025_ = _3026_ | _3028_ /*43889*/;
assign _2748_ = _3020_ ^ _3027_ /*43892*/;
assign _3034_ = D[54] ^ Q[57] /*43888*/;
assign _3031_ = _2363_ & _3034_ /*43884*/;
assign _3032_ = _2363_ ^ _3034_ /*43887*/;
assign _3033_ = _3025_ & _3032_ /*43885*/;
assign _3030_ = _3031_ | _3033_ /*43883*/;
assign _2749_ = _3025_ ^ _3032_ /*43886*/;
assign _3039_ = D[55] ^ Q[57] /*43882*/;
assign _3036_ = _2364_ & _3039_ /*43878*/;
assign _3037_ = _2364_ ^ _3039_ /*43881*/;
assign _3038_ = _3030_ & _3037_ /*43879*/;
assign _3035_ = _3036_ | _3038_ /*43877*/;
assign _2750_ = _3030_ ^ _3037_ /*43880*/;
assign _3044_ = D[56] ^ Q[57] /*43876*/;
assign _3041_ = _2365_ & _3044_ /*43872*/;
assign _3042_ = _2365_ ^ _3044_ /*43875*/;
assign _3043_ = _3035_ & _3042_ /*43873*/;
assign _3040_ = _3041_ | _3043_ /*43871*/;
assign _2751_ = _3035_ ^ _3042_ /*43874*/;
assign _3049_ = D[57] ^ Q[57] /*43870*/;
assign _3046_ = _2366_ & _3049_ /*43866*/;
assign _3047_ = _2366_ ^ _3049_ /*43869*/;
assign _3048_ = _3040_ & _3047_ /*43867*/;
assign _3045_ = _3046_ | _3048_ /*43865*/;
assign _2752_ = _3040_ ^ _3047_ /*43868*/;
assign _3054_ = D[58] ^ Q[57] /*43864*/;
assign _3051_ = _2367_ & _3054_ /*43860*/;
assign _3052_ = _2367_ ^ _3054_ /*43863*/;
assign _3053_ = _3045_ & _3052_ /*43861*/;
assign _3050_ = _3051_ | _3053_ /*43859*/;
assign _2753_ = _3045_ ^ _3052_ /*43862*/;
assign _3059_ = D[59] ^ Q[57] /*43858*/;
assign _3056_ = _2368_ & _3059_ /*43854*/;
assign _3057_ = _2368_ ^ _3059_ /*43857*/;
assign _3058_ = _3050_ & _3057_ /*43855*/;
assign _3055_ = _3056_ | _3058_ /*43853*/;
assign _2754_ = _3050_ ^ _3057_ /*43856*/;
assign _3064_ = D[60] ^ Q[57] /*43852*/;
assign _3061_ = _2369_ & _3064_ /*43848*/;
assign _3062_ = _2369_ ^ _3064_ /*43851*/;
assign _3063_ = _3055_ & _3062_ /*43849*/;
assign _3060_ = _3061_ | _3063_ /*43847*/;
assign _2755_ = _3055_ ^ _3062_ /*43850*/;
assign _3069_ = D[61] ^ Q[57] /*43846*/;
assign _3066_ = _2370_ & _3069_ /*43842*/;
assign _3067_ = _2370_ ^ _3069_ /*43845*/;
assign _3068_ = _3060_ & _3067_ /*43843*/;
assign _3065_ = _3066_ | _3068_ /*43841*/;
assign _2756_ = _3060_ ^ _3067_ /*43844*/;
assign _3074_ = D[62] ^ Q[57] /*43840*/;
assign _3071_ = _2371_ & _3074_ /*43836*/;
assign _3072_ = _2371_ ^ _3074_ /*43839*/;
assign _3073_ = _3065_ & _3072_ /*43837*/;
assign _3070_ = _3071_ | _3073_ /*43835*/;
assign _2757_ = _3065_ ^ _3072_ /*43838*/;
assign _3078_ = zeroWire ^ Q[57] /*43834*/;
assign _3075_ = _2372_ & _3078_ /*43830*/;
assign _3076_ = _2372_ ^ _3078_ /*43833*/;
assign _3077_ = _3070_ & _3076_ /*43831*/;
assign Q[56] = _3075_ | _3077_ /*43829*/;
assign _2758_ = _3070_ ^ _3076_ /*43832*/;
assign _3149_ = D[0] ^ Q[56] /*43443*/;
assign _3146_ = R_0[55] & _3149_ /*43439*/;
assign _3147_ = R_0[55] ^ _3149_ /*43442*/;
assign _3148_ = Q[56] & _3147_ /*43440*/;
assign _3145_ = _3146_ | _3148_ /*43438*/;
assign _3080_ = Q[56] ^ _3147_ /*43441*/;
assign _3154_ = D[1] ^ Q[56] /*43437*/;
assign _3151_ = _2695_ & _3154_ /*43433*/;
assign _3152_ = _2695_ ^ _3154_ /*43436*/;
assign _3153_ = _3145_ & _3152_ /*43434*/;
assign _3150_ = _3151_ | _3153_ /*43432*/;
assign _3081_ = _3145_ ^ _3152_ /*43435*/;
assign _3159_ = D[2] ^ Q[56] /*43431*/;
assign _3156_ = _2696_ & _3159_ /*43427*/;
assign _3157_ = _2696_ ^ _3159_ /*43430*/;
assign _3158_ = _3150_ & _3157_ /*43428*/;
assign _3155_ = _3156_ | _3158_ /*43426*/;
assign _3082_ = _3150_ ^ _3157_ /*43429*/;
assign _3164_ = D[3] ^ Q[56] /*43425*/;
assign _3161_ = _2697_ & _3164_ /*43421*/;
assign _3162_ = _2697_ ^ _3164_ /*43424*/;
assign _3163_ = _3155_ & _3162_ /*43422*/;
assign _3160_ = _3161_ | _3163_ /*43420*/;
assign _3083_ = _3155_ ^ _3162_ /*43423*/;
assign _3169_ = D[4] ^ Q[56] /*43419*/;
assign _3166_ = _2698_ & _3169_ /*43415*/;
assign _3167_ = _2698_ ^ _3169_ /*43418*/;
assign _3168_ = _3160_ & _3167_ /*43416*/;
assign _3165_ = _3166_ | _3168_ /*43414*/;
assign _3084_ = _3160_ ^ _3167_ /*43417*/;
assign _3174_ = D[5] ^ Q[56] /*43413*/;
assign _3171_ = _2699_ & _3174_ /*43409*/;
assign _3172_ = _2699_ ^ _3174_ /*43412*/;
assign _3173_ = _3165_ & _3172_ /*43410*/;
assign _3170_ = _3171_ | _3173_ /*43408*/;
assign _3085_ = _3165_ ^ _3172_ /*43411*/;
assign _3179_ = D[6] ^ Q[56] /*43407*/;
assign _3176_ = _2700_ & _3179_ /*43403*/;
assign _3177_ = _2700_ ^ _3179_ /*43406*/;
assign _3178_ = _3170_ & _3177_ /*43404*/;
assign _3175_ = _3176_ | _3178_ /*43402*/;
assign _3086_ = _3170_ ^ _3177_ /*43405*/;
assign _3184_ = D[7] ^ Q[56] /*43401*/;
assign _3181_ = _2701_ & _3184_ /*43397*/;
assign _3182_ = _2701_ ^ _3184_ /*43400*/;
assign _3183_ = _3175_ & _3182_ /*43398*/;
assign _3180_ = _3181_ | _3183_ /*43396*/;
assign _3087_ = _3175_ ^ _3182_ /*43399*/;
assign _3189_ = D[8] ^ Q[56] /*43395*/;
assign _3186_ = _2702_ & _3189_ /*43391*/;
assign _3187_ = _2702_ ^ _3189_ /*43394*/;
assign _3188_ = _3180_ & _3187_ /*43392*/;
assign _3185_ = _3186_ | _3188_ /*43390*/;
assign _3088_ = _3180_ ^ _3187_ /*43393*/;
assign _3194_ = D[9] ^ Q[56] /*43389*/;
assign _3191_ = _2703_ & _3194_ /*43385*/;
assign _3192_ = _2703_ ^ _3194_ /*43388*/;
assign _3193_ = _3185_ & _3192_ /*43386*/;
assign _3190_ = _3191_ | _3193_ /*43384*/;
assign _3089_ = _3185_ ^ _3192_ /*43387*/;
assign _3199_ = D[10] ^ Q[56] /*43383*/;
assign _3196_ = _2704_ & _3199_ /*43379*/;
assign _3197_ = _2704_ ^ _3199_ /*43382*/;
assign _3198_ = _3190_ & _3197_ /*43380*/;
assign _3195_ = _3196_ | _3198_ /*43378*/;
assign _3090_ = _3190_ ^ _3197_ /*43381*/;
assign _3204_ = D[11] ^ Q[56] /*43377*/;
assign _3201_ = _2705_ & _3204_ /*43373*/;
assign _3202_ = _2705_ ^ _3204_ /*43376*/;
assign _3203_ = _3195_ & _3202_ /*43374*/;
assign _3200_ = _3201_ | _3203_ /*43372*/;
assign _3091_ = _3195_ ^ _3202_ /*43375*/;
assign _3209_ = D[12] ^ Q[56] /*43371*/;
assign _3206_ = _2706_ & _3209_ /*43367*/;
assign _3207_ = _2706_ ^ _3209_ /*43370*/;
assign _3208_ = _3200_ & _3207_ /*43368*/;
assign _3205_ = _3206_ | _3208_ /*43366*/;
assign _3092_ = _3200_ ^ _3207_ /*43369*/;
assign _3214_ = D[13] ^ Q[56] /*43365*/;
assign _3211_ = _2707_ & _3214_ /*43361*/;
assign _3212_ = _2707_ ^ _3214_ /*43364*/;
assign _3213_ = _3205_ & _3212_ /*43362*/;
assign _3210_ = _3211_ | _3213_ /*43360*/;
assign _3093_ = _3205_ ^ _3212_ /*43363*/;
assign _3219_ = D[14] ^ Q[56] /*43359*/;
assign _3216_ = _2708_ & _3219_ /*43355*/;
assign _3217_ = _2708_ ^ _3219_ /*43358*/;
assign _3218_ = _3210_ & _3217_ /*43356*/;
assign _3215_ = _3216_ | _3218_ /*43354*/;
assign _3094_ = _3210_ ^ _3217_ /*43357*/;
assign _3224_ = D[15] ^ Q[56] /*43353*/;
assign _3221_ = _2709_ & _3224_ /*43349*/;
assign _3222_ = _2709_ ^ _3224_ /*43352*/;
assign _3223_ = _3215_ & _3222_ /*43350*/;
assign _3220_ = _3221_ | _3223_ /*43348*/;
assign _3095_ = _3215_ ^ _3222_ /*43351*/;
assign _3229_ = D[16] ^ Q[56] /*43347*/;
assign _3226_ = _2710_ & _3229_ /*43343*/;
assign _3227_ = _2710_ ^ _3229_ /*43346*/;
assign _3228_ = _3220_ & _3227_ /*43344*/;
assign _3225_ = _3226_ | _3228_ /*43342*/;
assign _3096_ = _3220_ ^ _3227_ /*43345*/;
assign _3234_ = D[17] ^ Q[56] /*43341*/;
assign _3231_ = _2711_ & _3234_ /*43337*/;
assign _3232_ = _2711_ ^ _3234_ /*43340*/;
assign _3233_ = _3225_ & _3232_ /*43338*/;
assign _3230_ = _3231_ | _3233_ /*43336*/;
assign _3097_ = _3225_ ^ _3232_ /*43339*/;
assign _3239_ = D[18] ^ Q[56] /*43335*/;
assign _3236_ = _2712_ & _3239_ /*43331*/;
assign _3237_ = _2712_ ^ _3239_ /*43334*/;
assign _3238_ = _3230_ & _3237_ /*43332*/;
assign _3235_ = _3236_ | _3238_ /*43330*/;
assign _3098_ = _3230_ ^ _3237_ /*43333*/;
assign _3244_ = D[19] ^ Q[56] /*43329*/;
assign _3241_ = _2713_ & _3244_ /*43325*/;
assign _3242_ = _2713_ ^ _3244_ /*43328*/;
assign _3243_ = _3235_ & _3242_ /*43326*/;
assign _3240_ = _3241_ | _3243_ /*43324*/;
assign _3099_ = _3235_ ^ _3242_ /*43327*/;
assign _3249_ = D[20] ^ Q[56] /*43323*/;
assign _3246_ = _2714_ & _3249_ /*43319*/;
assign _3247_ = _2714_ ^ _3249_ /*43322*/;
assign _3248_ = _3240_ & _3247_ /*43320*/;
assign _3245_ = _3246_ | _3248_ /*43318*/;
assign _3100_ = _3240_ ^ _3247_ /*43321*/;
assign _3254_ = D[21] ^ Q[56] /*43317*/;
assign _3251_ = _2715_ & _3254_ /*43313*/;
assign _3252_ = _2715_ ^ _3254_ /*43316*/;
assign _3253_ = _3245_ & _3252_ /*43314*/;
assign _3250_ = _3251_ | _3253_ /*43312*/;
assign _3101_ = _3245_ ^ _3252_ /*43315*/;
assign _3259_ = D[22] ^ Q[56] /*43311*/;
assign _3256_ = _2716_ & _3259_ /*43307*/;
assign _3257_ = _2716_ ^ _3259_ /*43310*/;
assign _3258_ = _3250_ & _3257_ /*43308*/;
assign _3255_ = _3256_ | _3258_ /*43306*/;
assign _3102_ = _3250_ ^ _3257_ /*43309*/;
assign _3264_ = D[23] ^ Q[56] /*43305*/;
assign _3261_ = _2717_ & _3264_ /*43301*/;
assign _3262_ = _2717_ ^ _3264_ /*43304*/;
assign _3263_ = _3255_ & _3262_ /*43302*/;
assign _3260_ = _3261_ | _3263_ /*43300*/;
assign _3103_ = _3255_ ^ _3262_ /*43303*/;
assign _3269_ = D[24] ^ Q[56] /*43299*/;
assign _3266_ = _2718_ & _3269_ /*43295*/;
assign _3267_ = _2718_ ^ _3269_ /*43298*/;
assign _3268_ = _3260_ & _3267_ /*43296*/;
assign _3265_ = _3266_ | _3268_ /*43294*/;
assign _3104_ = _3260_ ^ _3267_ /*43297*/;
assign _3274_ = D[25] ^ Q[56] /*43293*/;
assign _3271_ = _2719_ & _3274_ /*43289*/;
assign _3272_ = _2719_ ^ _3274_ /*43292*/;
assign _3273_ = _3265_ & _3272_ /*43290*/;
assign _3270_ = _3271_ | _3273_ /*43288*/;
assign _3105_ = _3265_ ^ _3272_ /*43291*/;
assign _3279_ = D[26] ^ Q[56] /*43287*/;
assign _3276_ = _2720_ & _3279_ /*43283*/;
assign _3277_ = _2720_ ^ _3279_ /*43286*/;
assign _3278_ = _3270_ & _3277_ /*43284*/;
assign _3275_ = _3276_ | _3278_ /*43282*/;
assign _3106_ = _3270_ ^ _3277_ /*43285*/;
assign _3284_ = D[27] ^ Q[56] /*43281*/;
assign _3281_ = _2721_ & _3284_ /*43277*/;
assign _3282_ = _2721_ ^ _3284_ /*43280*/;
assign _3283_ = _3275_ & _3282_ /*43278*/;
assign _3280_ = _3281_ | _3283_ /*43276*/;
assign _3107_ = _3275_ ^ _3282_ /*43279*/;
assign _3289_ = D[28] ^ Q[56] /*43275*/;
assign _3286_ = _2722_ & _3289_ /*43271*/;
assign _3287_ = _2722_ ^ _3289_ /*43274*/;
assign _3288_ = _3280_ & _3287_ /*43272*/;
assign _3285_ = _3286_ | _3288_ /*43270*/;
assign _3108_ = _3280_ ^ _3287_ /*43273*/;
assign _3294_ = D[29] ^ Q[56] /*43269*/;
assign _3291_ = _2723_ & _3294_ /*43265*/;
assign _3292_ = _2723_ ^ _3294_ /*43268*/;
assign _3293_ = _3285_ & _3292_ /*43266*/;
assign _3290_ = _3291_ | _3293_ /*43264*/;
assign _3109_ = _3285_ ^ _3292_ /*43267*/;
assign _3299_ = D[30] ^ Q[56] /*43263*/;
assign _3296_ = _2724_ & _3299_ /*43259*/;
assign _3297_ = _2724_ ^ _3299_ /*43262*/;
assign _3298_ = _3290_ & _3297_ /*43260*/;
assign _3295_ = _3296_ | _3298_ /*43258*/;
assign _3110_ = _3290_ ^ _3297_ /*43261*/;
assign _3304_ = D[31] ^ Q[56] /*43257*/;
assign _3301_ = _2725_ & _3304_ /*43253*/;
assign _3302_ = _2725_ ^ _3304_ /*43256*/;
assign _3303_ = _3295_ & _3302_ /*43254*/;
assign _3300_ = _3301_ | _3303_ /*43252*/;
assign _3111_ = _3295_ ^ _3302_ /*43255*/;
assign _3309_ = D[32] ^ Q[56] /*43251*/;
assign _3306_ = _2726_ & _3309_ /*43247*/;
assign _3307_ = _2726_ ^ _3309_ /*43250*/;
assign _3308_ = _3300_ & _3307_ /*43248*/;
assign _3305_ = _3306_ | _3308_ /*43246*/;
assign _3112_ = _3300_ ^ _3307_ /*43249*/;
assign _3314_ = D[33] ^ Q[56] /*43245*/;
assign _3311_ = _2727_ & _3314_ /*43241*/;
assign _3312_ = _2727_ ^ _3314_ /*43244*/;
assign _3313_ = _3305_ & _3312_ /*43242*/;
assign _3310_ = _3311_ | _3313_ /*43240*/;
assign _3113_ = _3305_ ^ _3312_ /*43243*/;
assign _3319_ = D[34] ^ Q[56] /*43239*/;
assign _3316_ = _2728_ & _3319_ /*43235*/;
assign _3317_ = _2728_ ^ _3319_ /*43238*/;
assign _3318_ = _3310_ & _3317_ /*43236*/;
assign _3315_ = _3316_ | _3318_ /*43234*/;
assign _3114_ = _3310_ ^ _3317_ /*43237*/;
assign _3324_ = D[35] ^ Q[56] /*43233*/;
assign _3321_ = _2729_ & _3324_ /*43229*/;
assign _3322_ = _2729_ ^ _3324_ /*43232*/;
assign _3323_ = _3315_ & _3322_ /*43230*/;
assign _3320_ = _3321_ | _3323_ /*43228*/;
assign _3115_ = _3315_ ^ _3322_ /*43231*/;
assign _3329_ = D[36] ^ Q[56] /*43227*/;
assign _3326_ = _2730_ & _3329_ /*43223*/;
assign _3327_ = _2730_ ^ _3329_ /*43226*/;
assign _3328_ = _3320_ & _3327_ /*43224*/;
assign _3325_ = _3326_ | _3328_ /*43222*/;
assign _3116_ = _3320_ ^ _3327_ /*43225*/;
assign _3334_ = D[37] ^ Q[56] /*43221*/;
assign _3331_ = _2731_ & _3334_ /*43217*/;
assign _3332_ = _2731_ ^ _3334_ /*43220*/;
assign _3333_ = _3325_ & _3332_ /*43218*/;
assign _3330_ = _3331_ | _3333_ /*43216*/;
assign _3117_ = _3325_ ^ _3332_ /*43219*/;
assign _3339_ = D[38] ^ Q[56] /*43215*/;
assign _3336_ = _2732_ & _3339_ /*43211*/;
assign _3337_ = _2732_ ^ _3339_ /*43214*/;
assign _3338_ = _3330_ & _3337_ /*43212*/;
assign _3335_ = _3336_ | _3338_ /*43210*/;
assign _3118_ = _3330_ ^ _3337_ /*43213*/;
assign _3344_ = D[39] ^ Q[56] /*43209*/;
assign _3341_ = _2733_ & _3344_ /*43205*/;
assign _3342_ = _2733_ ^ _3344_ /*43208*/;
assign _3343_ = _3335_ & _3342_ /*43206*/;
assign _3340_ = _3341_ | _3343_ /*43204*/;
assign _3119_ = _3335_ ^ _3342_ /*43207*/;
assign _3349_ = D[40] ^ Q[56] /*43203*/;
assign _3346_ = _2734_ & _3349_ /*43199*/;
assign _3347_ = _2734_ ^ _3349_ /*43202*/;
assign _3348_ = _3340_ & _3347_ /*43200*/;
assign _3345_ = _3346_ | _3348_ /*43198*/;
assign _3120_ = _3340_ ^ _3347_ /*43201*/;
assign _3354_ = D[41] ^ Q[56] /*43197*/;
assign _3351_ = _2735_ & _3354_ /*43193*/;
assign _3352_ = _2735_ ^ _3354_ /*43196*/;
assign _3353_ = _3345_ & _3352_ /*43194*/;
assign _3350_ = _3351_ | _3353_ /*43192*/;
assign _3121_ = _3345_ ^ _3352_ /*43195*/;
assign _3359_ = D[42] ^ Q[56] /*43191*/;
assign _3356_ = _2736_ & _3359_ /*43187*/;
assign _3357_ = _2736_ ^ _3359_ /*43190*/;
assign _3358_ = _3350_ & _3357_ /*43188*/;
assign _3355_ = _3356_ | _3358_ /*43186*/;
assign _3122_ = _3350_ ^ _3357_ /*43189*/;
assign _3364_ = D[43] ^ Q[56] /*43185*/;
assign _3361_ = _2737_ & _3364_ /*43181*/;
assign _3362_ = _2737_ ^ _3364_ /*43184*/;
assign _3363_ = _3355_ & _3362_ /*43182*/;
assign _3360_ = _3361_ | _3363_ /*43180*/;
assign _3123_ = _3355_ ^ _3362_ /*43183*/;
assign _3369_ = D[44] ^ Q[56] /*43179*/;
assign _3366_ = _2738_ & _3369_ /*43175*/;
assign _3367_ = _2738_ ^ _3369_ /*43178*/;
assign _3368_ = _3360_ & _3367_ /*43176*/;
assign _3365_ = _3366_ | _3368_ /*43174*/;
assign _3124_ = _3360_ ^ _3367_ /*43177*/;
assign _3374_ = D[45] ^ Q[56] /*43173*/;
assign _3371_ = _2739_ & _3374_ /*43169*/;
assign _3372_ = _2739_ ^ _3374_ /*43172*/;
assign _3373_ = _3365_ & _3372_ /*43170*/;
assign _3370_ = _3371_ | _3373_ /*43168*/;
assign _3125_ = _3365_ ^ _3372_ /*43171*/;
assign _3379_ = D[46] ^ Q[56] /*43167*/;
assign _3376_ = _2740_ & _3379_ /*43163*/;
assign _3377_ = _2740_ ^ _3379_ /*43166*/;
assign _3378_ = _3370_ & _3377_ /*43164*/;
assign _3375_ = _3376_ | _3378_ /*43162*/;
assign _3126_ = _3370_ ^ _3377_ /*43165*/;
assign _3384_ = D[47] ^ Q[56] /*43161*/;
assign _3381_ = _2741_ & _3384_ /*43157*/;
assign _3382_ = _2741_ ^ _3384_ /*43160*/;
assign _3383_ = _3375_ & _3382_ /*43158*/;
assign _3380_ = _3381_ | _3383_ /*43156*/;
assign _3127_ = _3375_ ^ _3382_ /*43159*/;
assign _3389_ = D[48] ^ Q[56] /*43155*/;
assign _3386_ = _2742_ & _3389_ /*43151*/;
assign _3387_ = _2742_ ^ _3389_ /*43154*/;
assign _3388_ = _3380_ & _3387_ /*43152*/;
assign _3385_ = _3386_ | _3388_ /*43150*/;
assign _3128_ = _3380_ ^ _3387_ /*43153*/;
assign _3394_ = D[49] ^ Q[56] /*43149*/;
assign _3391_ = _2743_ & _3394_ /*43145*/;
assign _3392_ = _2743_ ^ _3394_ /*43148*/;
assign _3393_ = _3385_ & _3392_ /*43146*/;
assign _3390_ = _3391_ | _3393_ /*43144*/;
assign _3129_ = _3385_ ^ _3392_ /*43147*/;
assign _3399_ = D[50] ^ Q[56] /*43143*/;
assign _3396_ = _2744_ & _3399_ /*43139*/;
assign _3397_ = _2744_ ^ _3399_ /*43142*/;
assign _3398_ = _3390_ & _3397_ /*43140*/;
assign _3395_ = _3396_ | _3398_ /*43138*/;
assign _3130_ = _3390_ ^ _3397_ /*43141*/;
assign _3404_ = D[51] ^ Q[56] /*43137*/;
assign _3401_ = _2745_ & _3404_ /*43133*/;
assign _3402_ = _2745_ ^ _3404_ /*43136*/;
assign _3403_ = _3395_ & _3402_ /*43134*/;
assign _3400_ = _3401_ | _3403_ /*43132*/;
assign _3131_ = _3395_ ^ _3402_ /*43135*/;
assign _3409_ = D[52] ^ Q[56] /*43131*/;
assign _3406_ = _2746_ & _3409_ /*43127*/;
assign _3407_ = _2746_ ^ _3409_ /*43130*/;
assign _3408_ = _3400_ & _3407_ /*43128*/;
assign _3405_ = _3406_ | _3408_ /*43126*/;
assign _3132_ = _3400_ ^ _3407_ /*43129*/;
assign _3414_ = D[53] ^ Q[56] /*43125*/;
assign _3411_ = _2747_ & _3414_ /*43121*/;
assign _3412_ = _2747_ ^ _3414_ /*43124*/;
assign _3413_ = _3405_ & _3412_ /*43122*/;
assign _3410_ = _3411_ | _3413_ /*43120*/;
assign _3133_ = _3405_ ^ _3412_ /*43123*/;
assign _3419_ = D[54] ^ Q[56] /*43119*/;
assign _3416_ = _2748_ & _3419_ /*43115*/;
assign _3417_ = _2748_ ^ _3419_ /*43118*/;
assign _3418_ = _3410_ & _3417_ /*43116*/;
assign _3415_ = _3416_ | _3418_ /*43114*/;
assign _3134_ = _3410_ ^ _3417_ /*43117*/;
assign _3424_ = D[55] ^ Q[56] /*43113*/;
assign _3421_ = _2749_ & _3424_ /*43109*/;
assign _3422_ = _2749_ ^ _3424_ /*43112*/;
assign _3423_ = _3415_ & _3422_ /*43110*/;
assign _3420_ = _3421_ | _3423_ /*43108*/;
assign _3135_ = _3415_ ^ _3422_ /*43111*/;
assign _3429_ = D[56] ^ Q[56] /*43107*/;
assign _3426_ = _2750_ & _3429_ /*43103*/;
assign _3427_ = _2750_ ^ _3429_ /*43106*/;
assign _3428_ = _3420_ & _3427_ /*43104*/;
assign _3425_ = _3426_ | _3428_ /*43102*/;
assign _3136_ = _3420_ ^ _3427_ /*43105*/;
assign _3434_ = D[57] ^ Q[56] /*43101*/;
assign _3431_ = _2751_ & _3434_ /*43097*/;
assign _3432_ = _2751_ ^ _3434_ /*43100*/;
assign _3433_ = _3425_ & _3432_ /*43098*/;
assign _3430_ = _3431_ | _3433_ /*43096*/;
assign _3137_ = _3425_ ^ _3432_ /*43099*/;
assign _3439_ = D[58] ^ Q[56] /*43095*/;
assign _3436_ = _2752_ & _3439_ /*43091*/;
assign _3437_ = _2752_ ^ _3439_ /*43094*/;
assign _3438_ = _3430_ & _3437_ /*43092*/;
assign _3435_ = _3436_ | _3438_ /*43090*/;
assign _3138_ = _3430_ ^ _3437_ /*43093*/;
assign _3444_ = D[59] ^ Q[56] /*43089*/;
assign _3441_ = _2753_ & _3444_ /*43085*/;
assign _3442_ = _2753_ ^ _3444_ /*43088*/;
assign _3443_ = _3435_ & _3442_ /*43086*/;
assign _3440_ = _3441_ | _3443_ /*43084*/;
assign _3139_ = _3435_ ^ _3442_ /*43087*/;
assign _3449_ = D[60] ^ Q[56] /*43083*/;
assign _3446_ = _2754_ & _3449_ /*43079*/;
assign _3447_ = _2754_ ^ _3449_ /*43082*/;
assign _3448_ = _3440_ & _3447_ /*43080*/;
assign _3445_ = _3446_ | _3448_ /*43078*/;
assign _3140_ = _3440_ ^ _3447_ /*43081*/;
assign _3454_ = D[61] ^ Q[56] /*43077*/;
assign _3451_ = _2755_ & _3454_ /*43073*/;
assign _3452_ = _2755_ ^ _3454_ /*43076*/;
assign _3453_ = _3445_ & _3452_ /*43074*/;
assign _3450_ = _3451_ | _3453_ /*43072*/;
assign _3141_ = _3445_ ^ _3452_ /*43075*/;
assign _3459_ = D[62] ^ Q[56] /*43071*/;
assign _3456_ = _2756_ & _3459_ /*43067*/;
assign _3457_ = _2756_ ^ _3459_ /*43070*/;
assign _3458_ = _3450_ & _3457_ /*43068*/;
assign _3455_ = _3456_ | _3458_ /*43066*/;
assign _3142_ = _3450_ ^ _3457_ /*43069*/;
assign _3463_ = zeroWire ^ Q[56] /*43065*/;
assign _3460_ = _2757_ & _3463_ /*43061*/;
assign _3461_ = _2757_ ^ _3463_ /*43064*/;
assign _3462_ = _3455_ & _3461_ /*43062*/;
assign Q[55] = _3460_ | _3462_ /*43060*/;
assign _3143_ = _3455_ ^ _3461_ /*43063*/;
assign _3534_ = D[0] ^ Q[55] /*42674*/;
assign _3531_ = R_0[54] & _3534_ /*42670*/;
assign _3532_ = R_0[54] ^ _3534_ /*42673*/;
assign _3533_ = Q[55] & _3532_ /*42671*/;
assign _3530_ = _3531_ | _3533_ /*42669*/;
assign _3465_ = Q[55] ^ _3532_ /*42672*/;
assign _3539_ = D[1] ^ Q[55] /*42668*/;
assign _3536_ = _3080_ & _3539_ /*42664*/;
assign _3537_ = _3080_ ^ _3539_ /*42667*/;
assign _3538_ = _3530_ & _3537_ /*42665*/;
assign _3535_ = _3536_ | _3538_ /*42663*/;
assign _3466_ = _3530_ ^ _3537_ /*42666*/;
assign _3544_ = D[2] ^ Q[55] /*42662*/;
assign _3541_ = _3081_ & _3544_ /*42658*/;
assign _3542_ = _3081_ ^ _3544_ /*42661*/;
assign _3543_ = _3535_ & _3542_ /*42659*/;
assign _3540_ = _3541_ | _3543_ /*42657*/;
assign _3467_ = _3535_ ^ _3542_ /*42660*/;
assign _3549_ = D[3] ^ Q[55] /*42656*/;
assign _3546_ = _3082_ & _3549_ /*42652*/;
assign _3547_ = _3082_ ^ _3549_ /*42655*/;
assign _3548_ = _3540_ & _3547_ /*42653*/;
assign _3545_ = _3546_ | _3548_ /*42651*/;
assign _3468_ = _3540_ ^ _3547_ /*42654*/;
assign _3554_ = D[4] ^ Q[55] /*42650*/;
assign _3551_ = _3083_ & _3554_ /*42646*/;
assign _3552_ = _3083_ ^ _3554_ /*42649*/;
assign _3553_ = _3545_ & _3552_ /*42647*/;
assign _3550_ = _3551_ | _3553_ /*42645*/;
assign _3469_ = _3545_ ^ _3552_ /*42648*/;
assign _3559_ = D[5] ^ Q[55] /*42644*/;
assign _3556_ = _3084_ & _3559_ /*42640*/;
assign _3557_ = _3084_ ^ _3559_ /*42643*/;
assign _3558_ = _3550_ & _3557_ /*42641*/;
assign _3555_ = _3556_ | _3558_ /*42639*/;
assign _3470_ = _3550_ ^ _3557_ /*42642*/;
assign _3564_ = D[6] ^ Q[55] /*42638*/;
assign _3561_ = _3085_ & _3564_ /*42634*/;
assign _3562_ = _3085_ ^ _3564_ /*42637*/;
assign _3563_ = _3555_ & _3562_ /*42635*/;
assign _3560_ = _3561_ | _3563_ /*42633*/;
assign _3471_ = _3555_ ^ _3562_ /*42636*/;
assign _3569_ = D[7] ^ Q[55] /*42632*/;
assign _3566_ = _3086_ & _3569_ /*42628*/;
assign _3567_ = _3086_ ^ _3569_ /*42631*/;
assign _3568_ = _3560_ & _3567_ /*42629*/;
assign _3565_ = _3566_ | _3568_ /*42627*/;
assign _3472_ = _3560_ ^ _3567_ /*42630*/;
assign _3574_ = D[8] ^ Q[55] /*42626*/;
assign _3571_ = _3087_ & _3574_ /*42622*/;
assign _3572_ = _3087_ ^ _3574_ /*42625*/;
assign _3573_ = _3565_ & _3572_ /*42623*/;
assign _3570_ = _3571_ | _3573_ /*42621*/;
assign _3473_ = _3565_ ^ _3572_ /*42624*/;
assign _3579_ = D[9] ^ Q[55] /*42620*/;
assign _3576_ = _3088_ & _3579_ /*42616*/;
assign _3577_ = _3088_ ^ _3579_ /*42619*/;
assign _3578_ = _3570_ & _3577_ /*42617*/;
assign _3575_ = _3576_ | _3578_ /*42615*/;
assign _3474_ = _3570_ ^ _3577_ /*42618*/;
assign _3584_ = D[10] ^ Q[55] /*42614*/;
assign _3581_ = _3089_ & _3584_ /*42610*/;
assign _3582_ = _3089_ ^ _3584_ /*42613*/;
assign _3583_ = _3575_ & _3582_ /*42611*/;
assign _3580_ = _3581_ | _3583_ /*42609*/;
assign _3475_ = _3575_ ^ _3582_ /*42612*/;
assign _3589_ = D[11] ^ Q[55] /*42608*/;
assign _3586_ = _3090_ & _3589_ /*42604*/;
assign _3587_ = _3090_ ^ _3589_ /*42607*/;
assign _3588_ = _3580_ & _3587_ /*42605*/;
assign _3585_ = _3586_ | _3588_ /*42603*/;
assign _3476_ = _3580_ ^ _3587_ /*42606*/;
assign _3594_ = D[12] ^ Q[55] /*42602*/;
assign _3591_ = _3091_ & _3594_ /*42598*/;
assign _3592_ = _3091_ ^ _3594_ /*42601*/;
assign _3593_ = _3585_ & _3592_ /*42599*/;
assign _3590_ = _3591_ | _3593_ /*42597*/;
assign _3477_ = _3585_ ^ _3592_ /*42600*/;
assign _3599_ = D[13] ^ Q[55] /*42596*/;
assign _3596_ = _3092_ & _3599_ /*42592*/;
assign _3597_ = _3092_ ^ _3599_ /*42595*/;
assign _3598_ = _3590_ & _3597_ /*42593*/;
assign _3595_ = _3596_ | _3598_ /*42591*/;
assign _3478_ = _3590_ ^ _3597_ /*42594*/;
assign _3604_ = D[14] ^ Q[55] /*42590*/;
assign _3601_ = _3093_ & _3604_ /*42586*/;
assign _3602_ = _3093_ ^ _3604_ /*42589*/;
assign _3603_ = _3595_ & _3602_ /*42587*/;
assign _3600_ = _3601_ | _3603_ /*42585*/;
assign _3479_ = _3595_ ^ _3602_ /*42588*/;
assign _3609_ = D[15] ^ Q[55] /*42584*/;
assign _3606_ = _3094_ & _3609_ /*42580*/;
assign _3607_ = _3094_ ^ _3609_ /*42583*/;
assign _3608_ = _3600_ & _3607_ /*42581*/;
assign _3605_ = _3606_ | _3608_ /*42579*/;
assign _3480_ = _3600_ ^ _3607_ /*42582*/;
assign _3614_ = D[16] ^ Q[55] /*42578*/;
assign _3611_ = _3095_ & _3614_ /*42574*/;
assign _3612_ = _3095_ ^ _3614_ /*42577*/;
assign _3613_ = _3605_ & _3612_ /*42575*/;
assign _3610_ = _3611_ | _3613_ /*42573*/;
assign _3481_ = _3605_ ^ _3612_ /*42576*/;
assign _3619_ = D[17] ^ Q[55] /*42572*/;
assign _3616_ = _3096_ & _3619_ /*42568*/;
assign _3617_ = _3096_ ^ _3619_ /*42571*/;
assign _3618_ = _3610_ & _3617_ /*42569*/;
assign _3615_ = _3616_ | _3618_ /*42567*/;
assign _3482_ = _3610_ ^ _3617_ /*42570*/;
assign _3624_ = D[18] ^ Q[55] /*42566*/;
assign _3621_ = _3097_ & _3624_ /*42562*/;
assign _3622_ = _3097_ ^ _3624_ /*42565*/;
assign _3623_ = _3615_ & _3622_ /*42563*/;
assign _3620_ = _3621_ | _3623_ /*42561*/;
assign _3483_ = _3615_ ^ _3622_ /*42564*/;
assign _3629_ = D[19] ^ Q[55] /*42560*/;
assign _3626_ = _3098_ & _3629_ /*42556*/;
assign _3627_ = _3098_ ^ _3629_ /*42559*/;
assign _3628_ = _3620_ & _3627_ /*42557*/;
assign _3625_ = _3626_ | _3628_ /*42555*/;
assign _3484_ = _3620_ ^ _3627_ /*42558*/;
assign _3634_ = D[20] ^ Q[55] /*42554*/;
assign _3631_ = _3099_ & _3634_ /*42550*/;
assign _3632_ = _3099_ ^ _3634_ /*42553*/;
assign _3633_ = _3625_ & _3632_ /*42551*/;
assign _3630_ = _3631_ | _3633_ /*42549*/;
assign _3485_ = _3625_ ^ _3632_ /*42552*/;
assign _3639_ = D[21] ^ Q[55] /*42548*/;
assign _3636_ = _3100_ & _3639_ /*42544*/;
assign _3637_ = _3100_ ^ _3639_ /*42547*/;
assign _3638_ = _3630_ & _3637_ /*42545*/;
assign _3635_ = _3636_ | _3638_ /*42543*/;
assign _3486_ = _3630_ ^ _3637_ /*42546*/;
assign _3644_ = D[22] ^ Q[55] /*42542*/;
assign _3641_ = _3101_ & _3644_ /*42538*/;
assign _3642_ = _3101_ ^ _3644_ /*42541*/;
assign _3643_ = _3635_ & _3642_ /*42539*/;
assign _3640_ = _3641_ | _3643_ /*42537*/;
assign _3487_ = _3635_ ^ _3642_ /*42540*/;
assign _3649_ = D[23] ^ Q[55] /*42536*/;
assign _3646_ = _3102_ & _3649_ /*42532*/;
assign _3647_ = _3102_ ^ _3649_ /*42535*/;
assign _3648_ = _3640_ & _3647_ /*42533*/;
assign _3645_ = _3646_ | _3648_ /*42531*/;
assign _3488_ = _3640_ ^ _3647_ /*42534*/;
assign _3654_ = D[24] ^ Q[55] /*42530*/;
assign _3651_ = _3103_ & _3654_ /*42526*/;
assign _3652_ = _3103_ ^ _3654_ /*42529*/;
assign _3653_ = _3645_ & _3652_ /*42527*/;
assign _3650_ = _3651_ | _3653_ /*42525*/;
assign _3489_ = _3645_ ^ _3652_ /*42528*/;
assign _3659_ = D[25] ^ Q[55] /*42524*/;
assign _3656_ = _3104_ & _3659_ /*42520*/;
assign _3657_ = _3104_ ^ _3659_ /*42523*/;
assign _3658_ = _3650_ & _3657_ /*42521*/;
assign _3655_ = _3656_ | _3658_ /*42519*/;
assign _3490_ = _3650_ ^ _3657_ /*42522*/;
assign _3664_ = D[26] ^ Q[55] /*42518*/;
assign _3661_ = _3105_ & _3664_ /*42514*/;
assign _3662_ = _3105_ ^ _3664_ /*42517*/;
assign _3663_ = _3655_ & _3662_ /*42515*/;
assign _3660_ = _3661_ | _3663_ /*42513*/;
assign _3491_ = _3655_ ^ _3662_ /*42516*/;
assign _3669_ = D[27] ^ Q[55] /*42512*/;
assign _3666_ = _3106_ & _3669_ /*42508*/;
assign _3667_ = _3106_ ^ _3669_ /*42511*/;
assign _3668_ = _3660_ & _3667_ /*42509*/;
assign _3665_ = _3666_ | _3668_ /*42507*/;
assign _3492_ = _3660_ ^ _3667_ /*42510*/;
assign _3674_ = D[28] ^ Q[55] /*42506*/;
assign _3671_ = _3107_ & _3674_ /*42502*/;
assign _3672_ = _3107_ ^ _3674_ /*42505*/;
assign _3673_ = _3665_ & _3672_ /*42503*/;
assign _3670_ = _3671_ | _3673_ /*42501*/;
assign _3493_ = _3665_ ^ _3672_ /*42504*/;
assign _3679_ = D[29] ^ Q[55] /*42500*/;
assign _3676_ = _3108_ & _3679_ /*42496*/;
assign _3677_ = _3108_ ^ _3679_ /*42499*/;
assign _3678_ = _3670_ & _3677_ /*42497*/;
assign _3675_ = _3676_ | _3678_ /*42495*/;
assign _3494_ = _3670_ ^ _3677_ /*42498*/;
assign _3684_ = D[30] ^ Q[55] /*42494*/;
assign _3681_ = _3109_ & _3684_ /*42490*/;
assign _3682_ = _3109_ ^ _3684_ /*42493*/;
assign _3683_ = _3675_ & _3682_ /*42491*/;
assign _3680_ = _3681_ | _3683_ /*42489*/;
assign _3495_ = _3675_ ^ _3682_ /*42492*/;
assign _3689_ = D[31] ^ Q[55] /*42488*/;
assign _3686_ = _3110_ & _3689_ /*42484*/;
assign _3687_ = _3110_ ^ _3689_ /*42487*/;
assign _3688_ = _3680_ & _3687_ /*42485*/;
assign _3685_ = _3686_ | _3688_ /*42483*/;
assign _3496_ = _3680_ ^ _3687_ /*42486*/;
assign _3694_ = D[32] ^ Q[55] /*42482*/;
assign _3691_ = _3111_ & _3694_ /*42478*/;
assign _3692_ = _3111_ ^ _3694_ /*42481*/;
assign _3693_ = _3685_ & _3692_ /*42479*/;
assign _3690_ = _3691_ | _3693_ /*42477*/;
assign _3497_ = _3685_ ^ _3692_ /*42480*/;
assign _3699_ = D[33] ^ Q[55] /*42476*/;
assign _3696_ = _3112_ & _3699_ /*42472*/;
assign _3697_ = _3112_ ^ _3699_ /*42475*/;
assign _3698_ = _3690_ & _3697_ /*42473*/;
assign _3695_ = _3696_ | _3698_ /*42471*/;
assign _3498_ = _3690_ ^ _3697_ /*42474*/;
assign _3704_ = D[34] ^ Q[55] /*42470*/;
assign _3701_ = _3113_ & _3704_ /*42466*/;
assign _3702_ = _3113_ ^ _3704_ /*42469*/;
assign _3703_ = _3695_ & _3702_ /*42467*/;
assign _3700_ = _3701_ | _3703_ /*42465*/;
assign _3499_ = _3695_ ^ _3702_ /*42468*/;
assign _3709_ = D[35] ^ Q[55] /*42464*/;
assign _3706_ = _3114_ & _3709_ /*42460*/;
assign _3707_ = _3114_ ^ _3709_ /*42463*/;
assign _3708_ = _3700_ & _3707_ /*42461*/;
assign _3705_ = _3706_ | _3708_ /*42459*/;
assign _3500_ = _3700_ ^ _3707_ /*42462*/;
assign _3714_ = D[36] ^ Q[55] /*42458*/;
assign _3711_ = _3115_ & _3714_ /*42454*/;
assign _3712_ = _3115_ ^ _3714_ /*42457*/;
assign _3713_ = _3705_ & _3712_ /*42455*/;
assign _3710_ = _3711_ | _3713_ /*42453*/;
assign _3501_ = _3705_ ^ _3712_ /*42456*/;
assign _3719_ = D[37] ^ Q[55] /*42452*/;
assign _3716_ = _3116_ & _3719_ /*42448*/;
assign _3717_ = _3116_ ^ _3719_ /*42451*/;
assign _3718_ = _3710_ & _3717_ /*42449*/;
assign _3715_ = _3716_ | _3718_ /*42447*/;
assign _3502_ = _3710_ ^ _3717_ /*42450*/;
assign _3724_ = D[38] ^ Q[55] /*42446*/;
assign _3721_ = _3117_ & _3724_ /*42442*/;
assign _3722_ = _3117_ ^ _3724_ /*42445*/;
assign _3723_ = _3715_ & _3722_ /*42443*/;
assign _3720_ = _3721_ | _3723_ /*42441*/;
assign _3503_ = _3715_ ^ _3722_ /*42444*/;
assign _3729_ = D[39] ^ Q[55] /*42440*/;
assign _3726_ = _3118_ & _3729_ /*42436*/;
assign _3727_ = _3118_ ^ _3729_ /*42439*/;
assign _3728_ = _3720_ & _3727_ /*42437*/;
assign _3725_ = _3726_ | _3728_ /*42435*/;
assign _3504_ = _3720_ ^ _3727_ /*42438*/;
assign _3734_ = D[40] ^ Q[55] /*42434*/;
assign _3731_ = _3119_ & _3734_ /*42430*/;
assign _3732_ = _3119_ ^ _3734_ /*42433*/;
assign _3733_ = _3725_ & _3732_ /*42431*/;
assign _3730_ = _3731_ | _3733_ /*42429*/;
assign _3505_ = _3725_ ^ _3732_ /*42432*/;
assign _3739_ = D[41] ^ Q[55] /*42428*/;
assign _3736_ = _3120_ & _3739_ /*42424*/;
assign _3737_ = _3120_ ^ _3739_ /*42427*/;
assign _3738_ = _3730_ & _3737_ /*42425*/;
assign _3735_ = _3736_ | _3738_ /*42423*/;
assign _3506_ = _3730_ ^ _3737_ /*42426*/;
assign _3744_ = D[42] ^ Q[55] /*42422*/;
assign _3741_ = _3121_ & _3744_ /*42418*/;
assign _3742_ = _3121_ ^ _3744_ /*42421*/;
assign _3743_ = _3735_ & _3742_ /*42419*/;
assign _3740_ = _3741_ | _3743_ /*42417*/;
assign _3507_ = _3735_ ^ _3742_ /*42420*/;
assign _3749_ = D[43] ^ Q[55] /*42416*/;
assign _3746_ = _3122_ & _3749_ /*42412*/;
assign _3747_ = _3122_ ^ _3749_ /*42415*/;
assign _3748_ = _3740_ & _3747_ /*42413*/;
assign _3745_ = _3746_ | _3748_ /*42411*/;
assign _3508_ = _3740_ ^ _3747_ /*42414*/;
assign _3754_ = D[44] ^ Q[55] /*42410*/;
assign _3751_ = _3123_ & _3754_ /*42406*/;
assign _3752_ = _3123_ ^ _3754_ /*42409*/;
assign _3753_ = _3745_ & _3752_ /*42407*/;
assign _3750_ = _3751_ | _3753_ /*42405*/;
assign _3509_ = _3745_ ^ _3752_ /*42408*/;
assign _3759_ = D[45] ^ Q[55] /*42404*/;
assign _3756_ = _3124_ & _3759_ /*42400*/;
assign _3757_ = _3124_ ^ _3759_ /*42403*/;
assign _3758_ = _3750_ & _3757_ /*42401*/;
assign _3755_ = _3756_ | _3758_ /*42399*/;
assign _3510_ = _3750_ ^ _3757_ /*42402*/;
assign _3764_ = D[46] ^ Q[55] /*42398*/;
assign _3761_ = _3125_ & _3764_ /*42394*/;
assign _3762_ = _3125_ ^ _3764_ /*42397*/;
assign _3763_ = _3755_ & _3762_ /*42395*/;
assign _3760_ = _3761_ | _3763_ /*42393*/;
assign _3511_ = _3755_ ^ _3762_ /*42396*/;
assign _3769_ = D[47] ^ Q[55] /*42392*/;
assign _3766_ = _3126_ & _3769_ /*42388*/;
assign _3767_ = _3126_ ^ _3769_ /*42391*/;
assign _3768_ = _3760_ & _3767_ /*42389*/;
assign _3765_ = _3766_ | _3768_ /*42387*/;
assign _3512_ = _3760_ ^ _3767_ /*42390*/;
assign _3774_ = D[48] ^ Q[55] /*42386*/;
assign _3771_ = _3127_ & _3774_ /*42382*/;
assign _3772_ = _3127_ ^ _3774_ /*42385*/;
assign _3773_ = _3765_ & _3772_ /*42383*/;
assign _3770_ = _3771_ | _3773_ /*42381*/;
assign _3513_ = _3765_ ^ _3772_ /*42384*/;
assign _3779_ = D[49] ^ Q[55] /*42380*/;
assign _3776_ = _3128_ & _3779_ /*42376*/;
assign _3777_ = _3128_ ^ _3779_ /*42379*/;
assign _3778_ = _3770_ & _3777_ /*42377*/;
assign _3775_ = _3776_ | _3778_ /*42375*/;
assign _3514_ = _3770_ ^ _3777_ /*42378*/;
assign _3784_ = D[50] ^ Q[55] /*42374*/;
assign _3781_ = _3129_ & _3784_ /*42370*/;
assign _3782_ = _3129_ ^ _3784_ /*42373*/;
assign _3783_ = _3775_ & _3782_ /*42371*/;
assign _3780_ = _3781_ | _3783_ /*42369*/;
assign _3515_ = _3775_ ^ _3782_ /*42372*/;
assign _3789_ = D[51] ^ Q[55] /*42368*/;
assign _3786_ = _3130_ & _3789_ /*42364*/;
assign _3787_ = _3130_ ^ _3789_ /*42367*/;
assign _3788_ = _3780_ & _3787_ /*42365*/;
assign _3785_ = _3786_ | _3788_ /*42363*/;
assign _3516_ = _3780_ ^ _3787_ /*42366*/;
assign _3794_ = D[52] ^ Q[55] /*42362*/;
assign _3791_ = _3131_ & _3794_ /*42358*/;
assign _3792_ = _3131_ ^ _3794_ /*42361*/;
assign _3793_ = _3785_ & _3792_ /*42359*/;
assign _3790_ = _3791_ | _3793_ /*42357*/;
assign _3517_ = _3785_ ^ _3792_ /*42360*/;
assign _3799_ = D[53] ^ Q[55] /*42356*/;
assign _3796_ = _3132_ & _3799_ /*42352*/;
assign _3797_ = _3132_ ^ _3799_ /*42355*/;
assign _3798_ = _3790_ & _3797_ /*42353*/;
assign _3795_ = _3796_ | _3798_ /*42351*/;
assign _3518_ = _3790_ ^ _3797_ /*42354*/;
assign _3804_ = D[54] ^ Q[55] /*42350*/;
assign _3801_ = _3133_ & _3804_ /*42346*/;
assign _3802_ = _3133_ ^ _3804_ /*42349*/;
assign _3803_ = _3795_ & _3802_ /*42347*/;
assign _3800_ = _3801_ | _3803_ /*42345*/;
assign _3519_ = _3795_ ^ _3802_ /*42348*/;
assign _3809_ = D[55] ^ Q[55] /*42344*/;
assign _3806_ = _3134_ & _3809_ /*42340*/;
assign _3807_ = _3134_ ^ _3809_ /*42343*/;
assign _3808_ = _3800_ & _3807_ /*42341*/;
assign _3805_ = _3806_ | _3808_ /*42339*/;
assign _3520_ = _3800_ ^ _3807_ /*42342*/;
assign _3814_ = D[56] ^ Q[55] /*42338*/;
assign _3811_ = _3135_ & _3814_ /*42334*/;
assign _3812_ = _3135_ ^ _3814_ /*42337*/;
assign _3813_ = _3805_ & _3812_ /*42335*/;
assign _3810_ = _3811_ | _3813_ /*42333*/;
assign _3521_ = _3805_ ^ _3812_ /*42336*/;
assign _3819_ = D[57] ^ Q[55] /*42332*/;
assign _3816_ = _3136_ & _3819_ /*42328*/;
assign _3817_ = _3136_ ^ _3819_ /*42331*/;
assign _3818_ = _3810_ & _3817_ /*42329*/;
assign _3815_ = _3816_ | _3818_ /*42327*/;
assign _3522_ = _3810_ ^ _3817_ /*42330*/;
assign _3824_ = D[58] ^ Q[55] /*42326*/;
assign _3821_ = _3137_ & _3824_ /*42322*/;
assign _3822_ = _3137_ ^ _3824_ /*42325*/;
assign _3823_ = _3815_ & _3822_ /*42323*/;
assign _3820_ = _3821_ | _3823_ /*42321*/;
assign _3523_ = _3815_ ^ _3822_ /*42324*/;
assign _3829_ = D[59] ^ Q[55] /*42320*/;
assign _3826_ = _3138_ & _3829_ /*42316*/;
assign _3827_ = _3138_ ^ _3829_ /*42319*/;
assign _3828_ = _3820_ & _3827_ /*42317*/;
assign _3825_ = _3826_ | _3828_ /*42315*/;
assign _3524_ = _3820_ ^ _3827_ /*42318*/;
assign _3834_ = D[60] ^ Q[55] /*42314*/;
assign _3831_ = _3139_ & _3834_ /*42310*/;
assign _3832_ = _3139_ ^ _3834_ /*42313*/;
assign _3833_ = _3825_ & _3832_ /*42311*/;
assign _3830_ = _3831_ | _3833_ /*42309*/;
assign _3525_ = _3825_ ^ _3832_ /*42312*/;
assign _3839_ = D[61] ^ Q[55] /*42308*/;
assign _3836_ = _3140_ & _3839_ /*42304*/;
assign _3837_ = _3140_ ^ _3839_ /*42307*/;
assign _3838_ = _3830_ & _3837_ /*42305*/;
assign _3835_ = _3836_ | _3838_ /*42303*/;
assign _3526_ = _3830_ ^ _3837_ /*42306*/;
assign _3844_ = D[62] ^ Q[55] /*42302*/;
assign _3841_ = _3141_ & _3844_ /*42298*/;
assign _3842_ = _3141_ ^ _3844_ /*42301*/;
assign _3843_ = _3835_ & _3842_ /*42299*/;
assign _3840_ = _3841_ | _3843_ /*42297*/;
assign _3527_ = _3835_ ^ _3842_ /*42300*/;
assign _3848_ = zeroWire ^ Q[55] /*42296*/;
assign _3845_ = _3142_ & _3848_ /*42292*/;
assign _3846_ = _3142_ ^ _3848_ /*42295*/;
assign _3847_ = _3840_ & _3846_ /*42293*/;
assign Q[54] = _3845_ | _3847_ /*42291*/;
assign _3528_ = _3840_ ^ _3846_ /*42294*/;
assign _3919_ = D[0] ^ Q[54] /*41905*/;
assign _3916_ = R_0[53] & _3919_ /*41901*/;
assign _3917_ = R_0[53] ^ _3919_ /*41904*/;
assign _3918_ = Q[54] & _3917_ /*41902*/;
assign _3915_ = _3916_ | _3918_ /*41900*/;
assign _3850_ = Q[54] ^ _3917_ /*41903*/;
assign _3924_ = D[1] ^ Q[54] /*41899*/;
assign _3921_ = _3465_ & _3924_ /*41895*/;
assign _3922_ = _3465_ ^ _3924_ /*41898*/;
assign _3923_ = _3915_ & _3922_ /*41896*/;
assign _3920_ = _3921_ | _3923_ /*41894*/;
assign _3851_ = _3915_ ^ _3922_ /*41897*/;
assign _3929_ = D[2] ^ Q[54] /*41893*/;
assign _3926_ = _3466_ & _3929_ /*41889*/;
assign _3927_ = _3466_ ^ _3929_ /*41892*/;
assign _3928_ = _3920_ & _3927_ /*41890*/;
assign _3925_ = _3926_ | _3928_ /*41888*/;
assign _3852_ = _3920_ ^ _3927_ /*41891*/;
assign _3934_ = D[3] ^ Q[54] /*41887*/;
assign _3931_ = _3467_ & _3934_ /*41883*/;
assign _3932_ = _3467_ ^ _3934_ /*41886*/;
assign _3933_ = _3925_ & _3932_ /*41884*/;
assign _3930_ = _3931_ | _3933_ /*41882*/;
assign _3853_ = _3925_ ^ _3932_ /*41885*/;
assign _3939_ = D[4] ^ Q[54] /*41881*/;
assign _3936_ = _3468_ & _3939_ /*41877*/;
assign _3937_ = _3468_ ^ _3939_ /*41880*/;
assign _3938_ = _3930_ & _3937_ /*41878*/;
assign _3935_ = _3936_ | _3938_ /*41876*/;
assign _3854_ = _3930_ ^ _3937_ /*41879*/;
assign _3944_ = D[5] ^ Q[54] /*41875*/;
assign _3941_ = _3469_ & _3944_ /*41871*/;
assign _3942_ = _3469_ ^ _3944_ /*41874*/;
assign _3943_ = _3935_ & _3942_ /*41872*/;
assign _3940_ = _3941_ | _3943_ /*41870*/;
assign _3855_ = _3935_ ^ _3942_ /*41873*/;
assign _3949_ = D[6] ^ Q[54] /*41869*/;
assign _3946_ = _3470_ & _3949_ /*41865*/;
assign _3947_ = _3470_ ^ _3949_ /*41868*/;
assign _3948_ = _3940_ & _3947_ /*41866*/;
assign _3945_ = _3946_ | _3948_ /*41864*/;
assign _3856_ = _3940_ ^ _3947_ /*41867*/;
assign _3954_ = D[7] ^ Q[54] /*41863*/;
assign _3951_ = _3471_ & _3954_ /*41859*/;
assign _3952_ = _3471_ ^ _3954_ /*41862*/;
assign _3953_ = _3945_ & _3952_ /*41860*/;
assign _3950_ = _3951_ | _3953_ /*41858*/;
assign _3857_ = _3945_ ^ _3952_ /*41861*/;
assign _3959_ = D[8] ^ Q[54] /*41857*/;
assign _3956_ = _3472_ & _3959_ /*41853*/;
assign _3957_ = _3472_ ^ _3959_ /*41856*/;
assign _3958_ = _3950_ & _3957_ /*41854*/;
assign _3955_ = _3956_ | _3958_ /*41852*/;
assign _3858_ = _3950_ ^ _3957_ /*41855*/;
assign _3964_ = D[9] ^ Q[54] /*41851*/;
assign _3961_ = _3473_ & _3964_ /*41847*/;
assign _3962_ = _3473_ ^ _3964_ /*41850*/;
assign _3963_ = _3955_ & _3962_ /*41848*/;
assign _3960_ = _3961_ | _3963_ /*41846*/;
assign _3859_ = _3955_ ^ _3962_ /*41849*/;
assign _3969_ = D[10] ^ Q[54] /*41845*/;
assign _3966_ = _3474_ & _3969_ /*41841*/;
assign _3967_ = _3474_ ^ _3969_ /*41844*/;
assign _3968_ = _3960_ & _3967_ /*41842*/;
assign _3965_ = _3966_ | _3968_ /*41840*/;
assign _3860_ = _3960_ ^ _3967_ /*41843*/;
assign _3974_ = D[11] ^ Q[54] /*41839*/;
assign _3971_ = _3475_ & _3974_ /*41835*/;
assign _3972_ = _3475_ ^ _3974_ /*41838*/;
assign _3973_ = _3965_ & _3972_ /*41836*/;
assign _3970_ = _3971_ | _3973_ /*41834*/;
assign _3861_ = _3965_ ^ _3972_ /*41837*/;
assign _3979_ = D[12] ^ Q[54] /*41833*/;
assign _3976_ = _3476_ & _3979_ /*41829*/;
assign _3977_ = _3476_ ^ _3979_ /*41832*/;
assign _3978_ = _3970_ & _3977_ /*41830*/;
assign _3975_ = _3976_ | _3978_ /*41828*/;
assign _3862_ = _3970_ ^ _3977_ /*41831*/;
assign _3984_ = D[13] ^ Q[54] /*41827*/;
assign _3981_ = _3477_ & _3984_ /*41823*/;
assign _3982_ = _3477_ ^ _3984_ /*41826*/;
assign _3983_ = _3975_ & _3982_ /*41824*/;
assign _3980_ = _3981_ | _3983_ /*41822*/;
assign _3863_ = _3975_ ^ _3982_ /*41825*/;
assign _3989_ = D[14] ^ Q[54] /*41821*/;
assign _3986_ = _3478_ & _3989_ /*41817*/;
assign _3987_ = _3478_ ^ _3989_ /*41820*/;
assign _3988_ = _3980_ & _3987_ /*41818*/;
assign _3985_ = _3986_ | _3988_ /*41816*/;
assign _3864_ = _3980_ ^ _3987_ /*41819*/;
assign _3994_ = D[15] ^ Q[54] /*41815*/;
assign _3991_ = _3479_ & _3994_ /*41811*/;
assign _3992_ = _3479_ ^ _3994_ /*41814*/;
assign _3993_ = _3985_ & _3992_ /*41812*/;
assign _3990_ = _3991_ | _3993_ /*41810*/;
assign _3865_ = _3985_ ^ _3992_ /*41813*/;
assign _3999_ = D[16] ^ Q[54] /*41809*/;
assign _3996_ = _3480_ & _3999_ /*41805*/;
assign _3997_ = _3480_ ^ _3999_ /*41808*/;
assign _3998_ = _3990_ & _3997_ /*41806*/;
assign _3995_ = _3996_ | _3998_ /*41804*/;
assign _3866_ = _3990_ ^ _3997_ /*41807*/;
assign _4004_ = D[17] ^ Q[54] /*41803*/;
assign _4001_ = _3481_ & _4004_ /*41799*/;
assign _4002_ = _3481_ ^ _4004_ /*41802*/;
assign _4003_ = _3995_ & _4002_ /*41800*/;
assign _4000_ = _4001_ | _4003_ /*41798*/;
assign _3867_ = _3995_ ^ _4002_ /*41801*/;
assign _4009_ = D[18] ^ Q[54] /*41797*/;
assign _4006_ = _3482_ & _4009_ /*41793*/;
assign _4007_ = _3482_ ^ _4009_ /*41796*/;
assign _4008_ = _4000_ & _4007_ /*41794*/;
assign _4005_ = _4006_ | _4008_ /*41792*/;
assign _3868_ = _4000_ ^ _4007_ /*41795*/;
assign _4014_ = D[19] ^ Q[54] /*41791*/;
assign _4011_ = _3483_ & _4014_ /*41787*/;
assign _4012_ = _3483_ ^ _4014_ /*41790*/;
assign _4013_ = _4005_ & _4012_ /*41788*/;
assign _4010_ = _4011_ | _4013_ /*41786*/;
assign _3869_ = _4005_ ^ _4012_ /*41789*/;
assign _4019_ = D[20] ^ Q[54] /*41785*/;
assign _4016_ = _3484_ & _4019_ /*41781*/;
assign _4017_ = _3484_ ^ _4019_ /*41784*/;
assign _4018_ = _4010_ & _4017_ /*41782*/;
assign _4015_ = _4016_ | _4018_ /*41780*/;
assign _3870_ = _4010_ ^ _4017_ /*41783*/;
assign _4024_ = D[21] ^ Q[54] /*41779*/;
assign _4021_ = _3485_ & _4024_ /*41775*/;
assign _4022_ = _3485_ ^ _4024_ /*41778*/;
assign _4023_ = _4015_ & _4022_ /*41776*/;
assign _4020_ = _4021_ | _4023_ /*41774*/;
assign _3871_ = _4015_ ^ _4022_ /*41777*/;
assign _4029_ = D[22] ^ Q[54] /*41773*/;
assign _4026_ = _3486_ & _4029_ /*41769*/;
assign _4027_ = _3486_ ^ _4029_ /*41772*/;
assign _4028_ = _4020_ & _4027_ /*41770*/;
assign _4025_ = _4026_ | _4028_ /*41768*/;
assign _3872_ = _4020_ ^ _4027_ /*41771*/;
assign _4034_ = D[23] ^ Q[54] /*41767*/;
assign _4031_ = _3487_ & _4034_ /*41763*/;
assign _4032_ = _3487_ ^ _4034_ /*41766*/;
assign _4033_ = _4025_ & _4032_ /*41764*/;
assign _4030_ = _4031_ | _4033_ /*41762*/;
assign _3873_ = _4025_ ^ _4032_ /*41765*/;
assign _4039_ = D[24] ^ Q[54] /*41761*/;
assign _4036_ = _3488_ & _4039_ /*41757*/;
assign _4037_ = _3488_ ^ _4039_ /*41760*/;
assign _4038_ = _4030_ & _4037_ /*41758*/;
assign _4035_ = _4036_ | _4038_ /*41756*/;
assign _3874_ = _4030_ ^ _4037_ /*41759*/;
assign _4044_ = D[25] ^ Q[54] /*41755*/;
assign _4041_ = _3489_ & _4044_ /*41751*/;
assign _4042_ = _3489_ ^ _4044_ /*41754*/;
assign _4043_ = _4035_ & _4042_ /*41752*/;
assign _4040_ = _4041_ | _4043_ /*41750*/;
assign _3875_ = _4035_ ^ _4042_ /*41753*/;
assign _4049_ = D[26] ^ Q[54] /*41749*/;
assign _4046_ = _3490_ & _4049_ /*41745*/;
assign _4047_ = _3490_ ^ _4049_ /*41748*/;
assign _4048_ = _4040_ & _4047_ /*41746*/;
assign _4045_ = _4046_ | _4048_ /*41744*/;
assign _3876_ = _4040_ ^ _4047_ /*41747*/;
assign _4054_ = D[27] ^ Q[54] /*41743*/;
assign _4051_ = _3491_ & _4054_ /*41739*/;
assign _4052_ = _3491_ ^ _4054_ /*41742*/;
assign _4053_ = _4045_ & _4052_ /*41740*/;
assign _4050_ = _4051_ | _4053_ /*41738*/;
assign _3877_ = _4045_ ^ _4052_ /*41741*/;
assign _4059_ = D[28] ^ Q[54] /*41737*/;
assign _4056_ = _3492_ & _4059_ /*41733*/;
assign _4057_ = _3492_ ^ _4059_ /*41736*/;
assign _4058_ = _4050_ & _4057_ /*41734*/;
assign _4055_ = _4056_ | _4058_ /*41732*/;
assign _3878_ = _4050_ ^ _4057_ /*41735*/;
assign _4064_ = D[29] ^ Q[54] /*41731*/;
assign _4061_ = _3493_ & _4064_ /*41727*/;
assign _4062_ = _3493_ ^ _4064_ /*41730*/;
assign _4063_ = _4055_ & _4062_ /*41728*/;
assign _4060_ = _4061_ | _4063_ /*41726*/;
assign _3879_ = _4055_ ^ _4062_ /*41729*/;
assign _4069_ = D[30] ^ Q[54] /*41725*/;
assign _4066_ = _3494_ & _4069_ /*41721*/;
assign _4067_ = _3494_ ^ _4069_ /*41724*/;
assign _4068_ = _4060_ & _4067_ /*41722*/;
assign _4065_ = _4066_ | _4068_ /*41720*/;
assign _3880_ = _4060_ ^ _4067_ /*41723*/;
assign _4074_ = D[31] ^ Q[54] /*41719*/;
assign _4071_ = _3495_ & _4074_ /*41715*/;
assign _4072_ = _3495_ ^ _4074_ /*41718*/;
assign _4073_ = _4065_ & _4072_ /*41716*/;
assign _4070_ = _4071_ | _4073_ /*41714*/;
assign _3881_ = _4065_ ^ _4072_ /*41717*/;
assign _4079_ = D[32] ^ Q[54] /*41713*/;
assign _4076_ = _3496_ & _4079_ /*41709*/;
assign _4077_ = _3496_ ^ _4079_ /*41712*/;
assign _4078_ = _4070_ & _4077_ /*41710*/;
assign _4075_ = _4076_ | _4078_ /*41708*/;
assign _3882_ = _4070_ ^ _4077_ /*41711*/;
assign _4084_ = D[33] ^ Q[54] /*41707*/;
assign _4081_ = _3497_ & _4084_ /*41703*/;
assign _4082_ = _3497_ ^ _4084_ /*41706*/;
assign _4083_ = _4075_ & _4082_ /*41704*/;
assign _4080_ = _4081_ | _4083_ /*41702*/;
assign _3883_ = _4075_ ^ _4082_ /*41705*/;
assign _4089_ = D[34] ^ Q[54] /*41701*/;
assign _4086_ = _3498_ & _4089_ /*41697*/;
assign _4087_ = _3498_ ^ _4089_ /*41700*/;
assign _4088_ = _4080_ & _4087_ /*41698*/;
assign _4085_ = _4086_ | _4088_ /*41696*/;
assign _3884_ = _4080_ ^ _4087_ /*41699*/;
assign _4094_ = D[35] ^ Q[54] /*41695*/;
assign _4091_ = _3499_ & _4094_ /*41691*/;
assign _4092_ = _3499_ ^ _4094_ /*41694*/;
assign _4093_ = _4085_ & _4092_ /*41692*/;
assign _4090_ = _4091_ | _4093_ /*41690*/;
assign _3885_ = _4085_ ^ _4092_ /*41693*/;
assign _4099_ = D[36] ^ Q[54] /*41689*/;
assign _4096_ = _3500_ & _4099_ /*41685*/;
assign _4097_ = _3500_ ^ _4099_ /*41688*/;
assign _4098_ = _4090_ & _4097_ /*41686*/;
assign _4095_ = _4096_ | _4098_ /*41684*/;
assign _3886_ = _4090_ ^ _4097_ /*41687*/;
assign _4104_ = D[37] ^ Q[54] /*41683*/;
assign _4101_ = _3501_ & _4104_ /*41679*/;
assign _4102_ = _3501_ ^ _4104_ /*41682*/;
assign _4103_ = _4095_ & _4102_ /*41680*/;
assign _4100_ = _4101_ | _4103_ /*41678*/;
assign _3887_ = _4095_ ^ _4102_ /*41681*/;
assign _4109_ = D[38] ^ Q[54] /*41677*/;
assign _4106_ = _3502_ & _4109_ /*41673*/;
assign _4107_ = _3502_ ^ _4109_ /*41676*/;
assign _4108_ = _4100_ & _4107_ /*41674*/;
assign _4105_ = _4106_ | _4108_ /*41672*/;
assign _3888_ = _4100_ ^ _4107_ /*41675*/;
assign _4114_ = D[39] ^ Q[54] /*41671*/;
assign _4111_ = _3503_ & _4114_ /*41667*/;
assign _4112_ = _3503_ ^ _4114_ /*41670*/;
assign _4113_ = _4105_ & _4112_ /*41668*/;
assign _4110_ = _4111_ | _4113_ /*41666*/;
assign _3889_ = _4105_ ^ _4112_ /*41669*/;
assign _4119_ = D[40] ^ Q[54] /*41665*/;
assign _4116_ = _3504_ & _4119_ /*41661*/;
assign _4117_ = _3504_ ^ _4119_ /*41664*/;
assign _4118_ = _4110_ & _4117_ /*41662*/;
assign _4115_ = _4116_ | _4118_ /*41660*/;
assign _3890_ = _4110_ ^ _4117_ /*41663*/;
assign _4124_ = D[41] ^ Q[54] /*41659*/;
assign _4121_ = _3505_ & _4124_ /*41655*/;
assign _4122_ = _3505_ ^ _4124_ /*41658*/;
assign _4123_ = _4115_ & _4122_ /*41656*/;
assign _4120_ = _4121_ | _4123_ /*41654*/;
assign _3891_ = _4115_ ^ _4122_ /*41657*/;
assign _4129_ = D[42] ^ Q[54] /*41653*/;
assign _4126_ = _3506_ & _4129_ /*41649*/;
assign _4127_ = _3506_ ^ _4129_ /*41652*/;
assign _4128_ = _4120_ & _4127_ /*41650*/;
assign _4125_ = _4126_ | _4128_ /*41648*/;
assign _3892_ = _4120_ ^ _4127_ /*41651*/;
assign _4134_ = D[43] ^ Q[54] /*41647*/;
assign _4131_ = _3507_ & _4134_ /*41643*/;
assign _4132_ = _3507_ ^ _4134_ /*41646*/;
assign _4133_ = _4125_ & _4132_ /*41644*/;
assign _4130_ = _4131_ | _4133_ /*41642*/;
assign _3893_ = _4125_ ^ _4132_ /*41645*/;
assign _4139_ = D[44] ^ Q[54] /*41641*/;
assign _4136_ = _3508_ & _4139_ /*41637*/;
assign _4137_ = _3508_ ^ _4139_ /*41640*/;
assign _4138_ = _4130_ & _4137_ /*41638*/;
assign _4135_ = _4136_ | _4138_ /*41636*/;
assign _3894_ = _4130_ ^ _4137_ /*41639*/;
assign _4144_ = D[45] ^ Q[54] /*41635*/;
assign _4141_ = _3509_ & _4144_ /*41631*/;
assign _4142_ = _3509_ ^ _4144_ /*41634*/;
assign _4143_ = _4135_ & _4142_ /*41632*/;
assign _4140_ = _4141_ | _4143_ /*41630*/;
assign _3895_ = _4135_ ^ _4142_ /*41633*/;
assign _4149_ = D[46] ^ Q[54] /*41629*/;
assign _4146_ = _3510_ & _4149_ /*41625*/;
assign _4147_ = _3510_ ^ _4149_ /*41628*/;
assign _4148_ = _4140_ & _4147_ /*41626*/;
assign _4145_ = _4146_ | _4148_ /*41624*/;
assign _3896_ = _4140_ ^ _4147_ /*41627*/;
assign _4154_ = D[47] ^ Q[54] /*41623*/;
assign _4151_ = _3511_ & _4154_ /*41619*/;
assign _4152_ = _3511_ ^ _4154_ /*41622*/;
assign _4153_ = _4145_ & _4152_ /*41620*/;
assign _4150_ = _4151_ | _4153_ /*41618*/;
assign _3897_ = _4145_ ^ _4152_ /*41621*/;
assign _4159_ = D[48] ^ Q[54] /*41617*/;
assign _4156_ = _3512_ & _4159_ /*41613*/;
assign _4157_ = _3512_ ^ _4159_ /*41616*/;
assign _4158_ = _4150_ & _4157_ /*41614*/;
assign _4155_ = _4156_ | _4158_ /*41612*/;
assign _3898_ = _4150_ ^ _4157_ /*41615*/;
assign _4164_ = D[49] ^ Q[54] /*41611*/;
assign _4161_ = _3513_ & _4164_ /*41607*/;
assign _4162_ = _3513_ ^ _4164_ /*41610*/;
assign _4163_ = _4155_ & _4162_ /*41608*/;
assign _4160_ = _4161_ | _4163_ /*41606*/;
assign _3899_ = _4155_ ^ _4162_ /*41609*/;
assign _4169_ = D[50] ^ Q[54] /*41605*/;
assign _4166_ = _3514_ & _4169_ /*41601*/;
assign _4167_ = _3514_ ^ _4169_ /*41604*/;
assign _4168_ = _4160_ & _4167_ /*41602*/;
assign _4165_ = _4166_ | _4168_ /*41600*/;
assign _3900_ = _4160_ ^ _4167_ /*41603*/;
assign _4174_ = D[51] ^ Q[54] /*41599*/;
assign _4171_ = _3515_ & _4174_ /*41595*/;
assign _4172_ = _3515_ ^ _4174_ /*41598*/;
assign _4173_ = _4165_ & _4172_ /*41596*/;
assign _4170_ = _4171_ | _4173_ /*41594*/;
assign _3901_ = _4165_ ^ _4172_ /*41597*/;
assign _4179_ = D[52] ^ Q[54] /*41593*/;
assign _4176_ = _3516_ & _4179_ /*41589*/;
assign _4177_ = _3516_ ^ _4179_ /*41592*/;
assign _4178_ = _4170_ & _4177_ /*41590*/;
assign _4175_ = _4176_ | _4178_ /*41588*/;
assign _3902_ = _4170_ ^ _4177_ /*41591*/;
assign _4184_ = D[53] ^ Q[54] /*41587*/;
assign _4181_ = _3517_ & _4184_ /*41583*/;
assign _4182_ = _3517_ ^ _4184_ /*41586*/;
assign _4183_ = _4175_ & _4182_ /*41584*/;
assign _4180_ = _4181_ | _4183_ /*41582*/;
assign _3903_ = _4175_ ^ _4182_ /*41585*/;
assign _4189_ = D[54] ^ Q[54] /*41581*/;
assign _4186_ = _3518_ & _4189_ /*41577*/;
assign _4187_ = _3518_ ^ _4189_ /*41580*/;
assign _4188_ = _4180_ & _4187_ /*41578*/;
assign _4185_ = _4186_ | _4188_ /*41576*/;
assign _3904_ = _4180_ ^ _4187_ /*41579*/;
assign _4194_ = D[55] ^ Q[54] /*41575*/;
assign _4191_ = _3519_ & _4194_ /*41571*/;
assign _4192_ = _3519_ ^ _4194_ /*41574*/;
assign _4193_ = _4185_ & _4192_ /*41572*/;
assign _4190_ = _4191_ | _4193_ /*41570*/;
assign _3905_ = _4185_ ^ _4192_ /*41573*/;
assign _4199_ = D[56] ^ Q[54] /*41569*/;
assign _4196_ = _3520_ & _4199_ /*41565*/;
assign _4197_ = _3520_ ^ _4199_ /*41568*/;
assign _4198_ = _4190_ & _4197_ /*41566*/;
assign _4195_ = _4196_ | _4198_ /*41564*/;
assign _3906_ = _4190_ ^ _4197_ /*41567*/;
assign _4204_ = D[57] ^ Q[54] /*41563*/;
assign _4201_ = _3521_ & _4204_ /*41559*/;
assign _4202_ = _3521_ ^ _4204_ /*41562*/;
assign _4203_ = _4195_ & _4202_ /*41560*/;
assign _4200_ = _4201_ | _4203_ /*41558*/;
assign _3907_ = _4195_ ^ _4202_ /*41561*/;
assign _4209_ = D[58] ^ Q[54] /*41557*/;
assign _4206_ = _3522_ & _4209_ /*41553*/;
assign _4207_ = _3522_ ^ _4209_ /*41556*/;
assign _4208_ = _4200_ & _4207_ /*41554*/;
assign _4205_ = _4206_ | _4208_ /*41552*/;
assign _3908_ = _4200_ ^ _4207_ /*41555*/;
assign _4214_ = D[59] ^ Q[54] /*41551*/;
assign _4211_ = _3523_ & _4214_ /*41547*/;
assign _4212_ = _3523_ ^ _4214_ /*41550*/;
assign _4213_ = _4205_ & _4212_ /*41548*/;
assign _4210_ = _4211_ | _4213_ /*41546*/;
assign _3909_ = _4205_ ^ _4212_ /*41549*/;
assign _4219_ = D[60] ^ Q[54] /*41545*/;
assign _4216_ = _3524_ & _4219_ /*41541*/;
assign _4217_ = _3524_ ^ _4219_ /*41544*/;
assign _4218_ = _4210_ & _4217_ /*41542*/;
assign _4215_ = _4216_ | _4218_ /*41540*/;
assign _3910_ = _4210_ ^ _4217_ /*41543*/;
assign _4224_ = D[61] ^ Q[54] /*41539*/;
assign _4221_ = _3525_ & _4224_ /*41535*/;
assign _4222_ = _3525_ ^ _4224_ /*41538*/;
assign _4223_ = _4215_ & _4222_ /*41536*/;
assign _4220_ = _4221_ | _4223_ /*41534*/;
assign _3911_ = _4215_ ^ _4222_ /*41537*/;
assign _4229_ = D[62] ^ Q[54] /*41533*/;
assign _4226_ = _3526_ & _4229_ /*41529*/;
assign _4227_ = _3526_ ^ _4229_ /*41532*/;
assign _4228_ = _4220_ & _4227_ /*41530*/;
assign _4225_ = _4226_ | _4228_ /*41528*/;
assign _3912_ = _4220_ ^ _4227_ /*41531*/;
assign _4233_ = zeroWire ^ Q[54] /*41527*/;
assign _4230_ = _3527_ & _4233_ /*41523*/;
assign _4231_ = _3527_ ^ _4233_ /*41526*/;
assign _4232_ = _4225_ & _4231_ /*41524*/;
assign Q[53] = _4230_ | _4232_ /*41522*/;
assign _3913_ = _4225_ ^ _4231_ /*41525*/;
assign _4304_ = D[0] ^ Q[53] /*41136*/;
assign _4301_ = R_0[52] & _4304_ /*41132*/;
assign _4302_ = R_0[52] ^ _4304_ /*41135*/;
assign _4303_ = Q[53] & _4302_ /*41133*/;
assign _4300_ = _4301_ | _4303_ /*41131*/;
assign _4235_ = Q[53] ^ _4302_ /*41134*/;
assign _4309_ = D[1] ^ Q[53] /*41130*/;
assign _4306_ = _3850_ & _4309_ /*41126*/;
assign _4307_ = _3850_ ^ _4309_ /*41129*/;
assign _4308_ = _4300_ & _4307_ /*41127*/;
assign _4305_ = _4306_ | _4308_ /*41125*/;
assign _4236_ = _4300_ ^ _4307_ /*41128*/;
assign _4314_ = D[2] ^ Q[53] /*41124*/;
assign _4311_ = _3851_ & _4314_ /*41120*/;
assign _4312_ = _3851_ ^ _4314_ /*41123*/;
assign _4313_ = _4305_ & _4312_ /*41121*/;
assign _4310_ = _4311_ | _4313_ /*41119*/;
assign _4237_ = _4305_ ^ _4312_ /*41122*/;
assign _4319_ = D[3] ^ Q[53] /*41118*/;
assign _4316_ = _3852_ & _4319_ /*41114*/;
assign _4317_ = _3852_ ^ _4319_ /*41117*/;
assign _4318_ = _4310_ & _4317_ /*41115*/;
assign _4315_ = _4316_ | _4318_ /*41113*/;
assign _4238_ = _4310_ ^ _4317_ /*41116*/;
assign _4324_ = D[4] ^ Q[53] /*41112*/;
assign _4321_ = _3853_ & _4324_ /*41108*/;
assign _4322_ = _3853_ ^ _4324_ /*41111*/;
assign _4323_ = _4315_ & _4322_ /*41109*/;
assign _4320_ = _4321_ | _4323_ /*41107*/;
assign _4239_ = _4315_ ^ _4322_ /*41110*/;
assign _4329_ = D[5] ^ Q[53] /*41106*/;
assign _4326_ = _3854_ & _4329_ /*41102*/;
assign _4327_ = _3854_ ^ _4329_ /*41105*/;
assign _4328_ = _4320_ & _4327_ /*41103*/;
assign _4325_ = _4326_ | _4328_ /*41101*/;
assign _4240_ = _4320_ ^ _4327_ /*41104*/;
assign _4334_ = D[6] ^ Q[53] /*41100*/;
assign _4331_ = _3855_ & _4334_ /*41096*/;
assign _4332_ = _3855_ ^ _4334_ /*41099*/;
assign _4333_ = _4325_ & _4332_ /*41097*/;
assign _4330_ = _4331_ | _4333_ /*41095*/;
assign _4241_ = _4325_ ^ _4332_ /*41098*/;
assign _4339_ = D[7] ^ Q[53] /*41094*/;
assign _4336_ = _3856_ & _4339_ /*41090*/;
assign _4337_ = _3856_ ^ _4339_ /*41093*/;
assign _4338_ = _4330_ & _4337_ /*41091*/;
assign _4335_ = _4336_ | _4338_ /*41089*/;
assign _4242_ = _4330_ ^ _4337_ /*41092*/;
assign _4344_ = D[8] ^ Q[53] /*41088*/;
assign _4341_ = _3857_ & _4344_ /*41084*/;
assign _4342_ = _3857_ ^ _4344_ /*41087*/;
assign _4343_ = _4335_ & _4342_ /*41085*/;
assign _4340_ = _4341_ | _4343_ /*41083*/;
assign _4243_ = _4335_ ^ _4342_ /*41086*/;
assign _4349_ = D[9] ^ Q[53] /*41082*/;
assign _4346_ = _3858_ & _4349_ /*41078*/;
assign _4347_ = _3858_ ^ _4349_ /*41081*/;
assign _4348_ = _4340_ & _4347_ /*41079*/;
assign _4345_ = _4346_ | _4348_ /*41077*/;
assign _4244_ = _4340_ ^ _4347_ /*41080*/;
assign _4354_ = D[10] ^ Q[53] /*41076*/;
assign _4351_ = _3859_ & _4354_ /*41072*/;
assign _4352_ = _3859_ ^ _4354_ /*41075*/;
assign _4353_ = _4345_ & _4352_ /*41073*/;
assign _4350_ = _4351_ | _4353_ /*41071*/;
assign _4245_ = _4345_ ^ _4352_ /*41074*/;
assign _4359_ = D[11] ^ Q[53] /*41070*/;
assign _4356_ = _3860_ & _4359_ /*41066*/;
assign _4357_ = _3860_ ^ _4359_ /*41069*/;
assign _4358_ = _4350_ & _4357_ /*41067*/;
assign _4355_ = _4356_ | _4358_ /*41065*/;
assign _4246_ = _4350_ ^ _4357_ /*41068*/;
assign _4364_ = D[12] ^ Q[53] /*41064*/;
assign _4361_ = _3861_ & _4364_ /*41060*/;
assign _4362_ = _3861_ ^ _4364_ /*41063*/;
assign _4363_ = _4355_ & _4362_ /*41061*/;
assign _4360_ = _4361_ | _4363_ /*41059*/;
assign _4247_ = _4355_ ^ _4362_ /*41062*/;
assign _4369_ = D[13] ^ Q[53] /*41058*/;
assign _4366_ = _3862_ & _4369_ /*41054*/;
assign _4367_ = _3862_ ^ _4369_ /*41057*/;
assign _4368_ = _4360_ & _4367_ /*41055*/;
assign _4365_ = _4366_ | _4368_ /*41053*/;
assign _4248_ = _4360_ ^ _4367_ /*41056*/;
assign _4374_ = D[14] ^ Q[53] /*41052*/;
assign _4371_ = _3863_ & _4374_ /*41048*/;
assign _4372_ = _3863_ ^ _4374_ /*41051*/;
assign _4373_ = _4365_ & _4372_ /*41049*/;
assign _4370_ = _4371_ | _4373_ /*41047*/;
assign _4249_ = _4365_ ^ _4372_ /*41050*/;
assign _4379_ = D[15] ^ Q[53] /*41046*/;
assign _4376_ = _3864_ & _4379_ /*41042*/;
assign _4377_ = _3864_ ^ _4379_ /*41045*/;
assign _4378_ = _4370_ & _4377_ /*41043*/;
assign _4375_ = _4376_ | _4378_ /*41041*/;
assign _4250_ = _4370_ ^ _4377_ /*41044*/;
assign _4384_ = D[16] ^ Q[53] /*41040*/;
assign _4381_ = _3865_ & _4384_ /*41036*/;
assign _4382_ = _3865_ ^ _4384_ /*41039*/;
assign _4383_ = _4375_ & _4382_ /*41037*/;
assign _4380_ = _4381_ | _4383_ /*41035*/;
assign _4251_ = _4375_ ^ _4382_ /*41038*/;
assign _4389_ = D[17] ^ Q[53] /*41034*/;
assign _4386_ = _3866_ & _4389_ /*41030*/;
assign _4387_ = _3866_ ^ _4389_ /*41033*/;
assign _4388_ = _4380_ & _4387_ /*41031*/;
assign _4385_ = _4386_ | _4388_ /*41029*/;
assign _4252_ = _4380_ ^ _4387_ /*41032*/;
assign _4394_ = D[18] ^ Q[53] /*41028*/;
assign _4391_ = _3867_ & _4394_ /*41024*/;
assign _4392_ = _3867_ ^ _4394_ /*41027*/;
assign _4393_ = _4385_ & _4392_ /*41025*/;
assign _4390_ = _4391_ | _4393_ /*41023*/;
assign _4253_ = _4385_ ^ _4392_ /*41026*/;
assign _4399_ = D[19] ^ Q[53] /*41022*/;
assign _4396_ = _3868_ & _4399_ /*41018*/;
assign _4397_ = _3868_ ^ _4399_ /*41021*/;
assign _4398_ = _4390_ & _4397_ /*41019*/;
assign _4395_ = _4396_ | _4398_ /*41017*/;
assign _4254_ = _4390_ ^ _4397_ /*41020*/;
assign _4404_ = D[20] ^ Q[53] /*41016*/;
assign _4401_ = _3869_ & _4404_ /*41012*/;
assign _4402_ = _3869_ ^ _4404_ /*41015*/;
assign _4403_ = _4395_ & _4402_ /*41013*/;
assign _4400_ = _4401_ | _4403_ /*41011*/;
assign _4255_ = _4395_ ^ _4402_ /*41014*/;
assign _4409_ = D[21] ^ Q[53] /*41010*/;
assign _4406_ = _3870_ & _4409_ /*41006*/;
assign _4407_ = _3870_ ^ _4409_ /*41009*/;
assign _4408_ = _4400_ & _4407_ /*41007*/;
assign _4405_ = _4406_ | _4408_ /*41005*/;
assign _4256_ = _4400_ ^ _4407_ /*41008*/;
assign _4414_ = D[22] ^ Q[53] /*41004*/;
assign _4411_ = _3871_ & _4414_ /*41000*/;
assign _4412_ = _3871_ ^ _4414_ /*41003*/;
assign _4413_ = _4405_ & _4412_ /*41001*/;
assign _4410_ = _4411_ | _4413_ /*40999*/;
assign _4257_ = _4405_ ^ _4412_ /*41002*/;
assign _4419_ = D[23] ^ Q[53] /*40998*/;
assign _4416_ = _3872_ & _4419_ /*40994*/;
assign _4417_ = _3872_ ^ _4419_ /*40997*/;
assign _4418_ = _4410_ & _4417_ /*40995*/;
assign _4415_ = _4416_ | _4418_ /*40993*/;
assign _4258_ = _4410_ ^ _4417_ /*40996*/;
assign _4424_ = D[24] ^ Q[53] /*40992*/;
assign _4421_ = _3873_ & _4424_ /*40988*/;
assign _4422_ = _3873_ ^ _4424_ /*40991*/;
assign _4423_ = _4415_ & _4422_ /*40989*/;
assign _4420_ = _4421_ | _4423_ /*40987*/;
assign _4259_ = _4415_ ^ _4422_ /*40990*/;
assign _4429_ = D[25] ^ Q[53] /*40986*/;
assign _4426_ = _3874_ & _4429_ /*40982*/;
assign _4427_ = _3874_ ^ _4429_ /*40985*/;
assign _4428_ = _4420_ & _4427_ /*40983*/;
assign _4425_ = _4426_ | _4428_ /*40981*/;
assign _4260_ = _4420_ ^ _4427_ /*40984*/;
assign _4434_ = D[26] ^ Q[53] /*40980*/;
assign _4431_ = _3875_ & _4434_ /*40976*/;
assign _4432_ = _3875_ ^ _4434_ /*40979*/;
assign _4433_ = _4425_ & _4432_ /*40977*/;
assign _4430_ = _4431_ | _4433_ /*40975*/;
assign _4261_ = _4425_ ^ _4432_ /*40978*/;
assign _4439_ = D[27] ^ Q[53] /*40974*/;
assign _4436_ = _3876_ & _4439_ /*40970*/;
assign _4437_ = _3876_ ^ _4439_ /*40973*/;
assign _4438_ = _4430_ & _4437_ /*40971*/;
assign _4435_ = _4436_ | _4438_ /*40969*/;
assign _4262_ = _4430_ ^ _4437_ /*40972*/;
assign _4444_ = D[28] ^ Q[53] /*40968*/;
assign _4441_ = _3877_ & _4444_ /*40964*/;
assign _4442_ = _3877_ ^ _4444_ /*40967*/;
assign _4443_ = _4435_ & _4442_ /*40965*/;
assign _4440_ = _4441_ | _4443_ /*40963*/;
assign _4263_ = _4435_ ^ _4442_ /*40966*/;
assign _4449_ = D[29] ^ Q[53] /*40962*/;
assign _4446_ = _3878_ & _4449_ /*40958*/;
assign _4447_ = _3878_ ^ _4449_ /*40961*/;
assign _4448_ = _4440_ & _4447_ /*40959*/;
assign _4445_ = _4446_ | _4448_ /*40957*/;
assign _4264_ = _4440_ ^ _4447_ /*40960*/;
assign _4454_ = D[30] ^ Q[53] /*40956*/;
assign _4451_ = _3879_ & _4454_ /*40952*/;
assign _4452_ = _3879_ ^ _4454_ /*40955*/;
assign _4453_ = _4445_ & _4452_ /*40953*/;
assign _4450_ = _4451_ | _4453_ /*40951*/;
assign _4265_ = _4445_ ^ _4452_ /*40954*/;
assign _4459_ = D[31] ^ Q[53] /*40950*/;
assign _4456_ = _3880_ & _4459_ /*40946*/;
assign _4457_ = _3880_ ^ _4459_ /*40949*/;
assign _4458_ = _4450_ & _4457_ /*40947*/;
assign _4455_ = _4456_ | _4458_ /*40945*/;
assign _4266_ = _4450_ ^ _4457_ /*40948*/;
assign _4464_ = D[32] ^ Q[53] /*40944*/;
assign _4461_ = _3881_ & _4464_ /*40940*/;
assign _4462_ = _3881_ ^ _4464_ /*40943*/;
assign _4463_ = _4455_ & _4462_ /*40941*/;
assign _4460_ = _4461_ | _4463_ /*40939*/;
assign _4267_ = _4455_ ^ _4462_ /*40942*/;
assign _4469_ = D[33] ^ Q[53] /*40938*/;
assign _4466_ = _3882_ & _4469_ /*40934*/;
assign _4467_ = _3882_ ^ _4469_ /*40937*/;
assign _4468_ = _4460_ & _4467_ /*40935*/;
assign _4465_ = _4466_ | _4468_ /*40933*/;
assign _4268_ = _4460_ ^ _4467_ /*40936*/;
assign _4474_ = D[34] ^ Q[53] /*40932*/;
assign _4471_ = _3883_ & _4474_ /*40928*/;
assign _4472_ = _3883_ ^ _4474_ /*40931*/;
assign _4473_ = _4465_ & _4472_ /*40929*/;
assign _4470_ = _4471_ | _4473_ /*40927*/;
assign _4269_ = _4465_ ^ _4472_ /*40930*/;
assign _4479_ = D[35] ^ Q[53] /*40926*/;
assign _4476_ = _3884_ & _4479_ /*40922*/;
assign _4477_ = _3884_ ^ _4479_ /*40925*/;
assign _4478_ = _4470_ & _4477_ /*40923*/;
assign _4475_ = _4476_ | _4478_ /*40921*/;
assign _4270_ = _4470_ ^ _4477_ /*40924*/;
assign _4484_ = D[36] ^ Q[53] /*40920*/;
assign _4481_ = _3885_ & _4484_ /*40916*/;
assign _4482_ = _3885_ ^ _4484_ /*40919*/;
assign _4483_ = _4475_ & _4482_ /*40917*/;
assign _4480_ = _4481_ | _4483_ /*40915*/;
assign _4271_ = _4475_ ^ _4482_ /*40918*/;
assign _4489_ = D[37] ^ Q[53] /*40914*/;
assign _4486_ = _3886_ & _4489_ /*40910*/;
assign _4487_ = _3886_ ^ _4489_ /*40913*/;
assign _4488_ = _4480_ & _4487_ /*40911*/;
assign _4485_ = _4486_ | _4488_ /*40909*/;
assign _4272_ = _4480_ ^ _4487_ /*40912*/;
assign _4494_ = D[38] ^ Q[53] /*40908*/;
assign _4491_ = _3887_ & _4494_ /*40904*/;
assign _4492_ = _3887_ ^ _4494_ /*40907*/;
assign _4493_ = _4485_ & _4492_ /*40905*/;
assign _4490_ = _4491_ | _4493_ /*40903*/;
assign _4273_ = _4485_ ^ _4492_ /*40906*/;
assign _4499_ = D[39] ^ Q[53] /*40902*/;
assign _4496_ = _3888_ & _4499_ /*40898*/;
assign _4497_ = _3888_ ^ _4499_ /*40901*/;
assign _4498_ = _4490_ & _4497_ /*40899*/;
assign _4495_ = _4496_ | _4498_ /*40897*/;
assign _4274_ = _4490_ ^ _4497_ /*40900*/;
assign _4504_ = D[40] ^ Q[53] /*40896*/;
assign _4501_ = _3889_ & _4504_ /*40892*/;
assign _4502_ = _3889_ ^ _4504_ /*40895*/;
assign _4503_ = _4495_ & _4502_ /*40893*/;
assign _4500_ = _4501_ | _4503_ /*40891*/;
assign _4275_ = _4495_ ^ _4502_ /*40894*/;
assign _4509_ = D[41] ^ Q[53] /*40890*/;
assign _4506_ = _3890_ & _4509_ /*40886*/;
assign _4507_ = _3890_ ^ _4509_ /*40889*/;
assign _4508_ = _4500_ & _4507_ /*40887*/;
assign _4505_ = _4506_ | _4508_ /*40885*/;
assign _4276_ = _4500_ ^ _4507_ /*40888*/;
assign _4514_ = D[42] ^ Q[53] /*40884*/;
assign _4511_ = _3891_ & _4514_ /*40880*/;
assign _4512_ = _3891_ ^ _4514_ /*40883*/;
assign _4513_ = _4505_ & _4512_ /*40881*/;
assign _4510_ = _4511_ | _4513_ /*40879*/;
assign _4277_ = _4505_ ^ _4512_ /*40882*/;
assign _4519_ = D[43] ^ Q[53] /*40878*/;
assign _4516_ = _3892_ & _4519_ /*40874*/;
assign _4517_ = _3892_ ^ _4519_ /*40877*/;
assign _4518_ = _4510_ & _4517_ /*40875*/;
assign _4515_ = _4516_ | _4518_ /*40873*/;
assign _4278_ = _4510_ ^ _4517_ /*40876*/;
assign _4524_ = D[44] ^ Q[53] /*40872*/;
assign _4521_ = _3893_ & _4524_ /*40868*/;
assign _4522_ = _3893_ ^ _4524_ /*40871*/;
assign _4523_ = _4515_ & _4522_ /*40869*/;
assign _4520_ = _4521_ | _4523_ /*40867*/;
assign _4279_ = _4515_ ^ _4522_ /*40870*/;
assign _4529_ = D[45] ^ Q[53] /*40866*/;
assign _4526_ = _3894_ & _4529_ /*40862*/;
assign _4527_ = _3894_ ^ _4529_ /*40865*/;
assign _4528_ = _4520_ & _4527_ /*40863*/;
assign _4525_ = _4526_ | _4528_ /*40861*/;
assign _4280_ = _4520_ ^ _4527_ /*40864*/;
assign _4534_ = D[46] ^ Q[53] /*40860*/;
assign _4531_ = _3895_ & _4534_ /*40856*/;
assign _4532_ = _3895_ ^ _4534_ /*40859*/;
assign _4533_ = _4525_ & _4532_ /*40857*/;
assign _4530_ = _4531_ | _4533_ /*40855*/;
assign _4281_ = _4525_ ^ _4532_ /*40858*/;
assign _4539_ = D[47] ^ Q[53] /*40854*/;
assign _4536_ = _3896_ & _4539_ /*40850*/;
assign _4537_ = _3896_ ^ _4539_ /*40853*/;
assign _4538_ = _4530_ & _4537_ /*40851*/;
assign _4535_ = _4536_ | _4538_ /*40849*/;
assign _4282_ = _4530_ ^ _4537_ /*40852*/;
assign _4544_ = D[48] ^ Q[53] /*40848*/;
assign _4541_ = _3897_ & _4544_ /*40844*/;
assign _4542_ = _3897_ ^ _4544_ /*40847*/;
assign _4543_ = _4535_ & _4542_ /*40845*/;
assign _4540_ = _4541_ | _4543_ /*40843*/;
assign _4283_ = _4535_ ^ _4542_ /*40846*/;
assign _4549_ = D[49] ^ Q[53] /*40842*/;
assign _4546_ = _3898_ & _4549_ /*40838*/;
assign _4547_ = _3898_ ^ _4549_ /*40841*/;
assign _4548_ = _4540_ & _4547_ /*40839*/;
assign _4545_ = _4546_ | _4548_ /*40837*/;
assign _4284_ = _4540_ ^ _4547_ /*40840*/;
assign _4554_ = D[50] ^ Q[53] /*40836*/;
assign _4551_ = _3899_ & _4554_ /*40832*/;
assign _4552_ = _3899_ ^ _4554_ /*40835*/;
assign _4553_ = _4545_ & _4552_ /*40833*/;
assign _4550_ = _4551_ | _4553_ /*40831*/;
assign _4285_ = _4545_ ^ _4552_ /*40834*/;
assign _4559_ = D[51] ^ Q[53] /*40830*/;
assign _4556_ = _3900_ & _4559_ /*40826*/;
assign _4557_ = _3900_ ^ _4559_ /*40829*/;
assign _4558_ = _4550_ & _4557_ /*40827*/;
assign _4555_ = _4556_ | _4558_ /*40825*/;
assign _4286_ = _4550_ ^ _4557_ /*40828*/;
assign _4564_ = D[52] ^ Q[53] /*40824*/;
assign _4561_ = _3901_ & _4564_ /*40820*/;
assign _4562_ = _3901_ ^ _4564_ /*40823*/;
assign _4563_ = _4555_ & _4562_ /*40821*/;
assign _4560_ = _4561_ | _4563_ /*40819*/;
assign _4287_ = _4555_ ^ _4562_ /*40822*/;
assign _4569_ = D[53] ^ Q[53] /*40818*/;
assign _4566_ = _3902_ & _4569_ /*40814*/;
assign _4567_ = _3902_ ^ _4569_ /*40817*/;
assign _4568_ = _4560_ & _4567_ /*40815*/;
assign _4565_ = _4566_ | _4568_ /*40813*/;
assign _4288_ = _4560_ ^ _4567_ /*40816*/;
assign _4574_ = D[54] ^ Q[53] /*40812*/;
assign _4571_ = _3903_ & _4574_ /*40808*/;
assign _4572_ = _3903_ ^ _4574_ /*40811*/;
assign _4573_ = _4565_ & _4572_ /*40809*/;
assign _4570_ = _4571_ | _4573_ /*40807*/;
assign _4289_ = _4565_ ^ _4572_ /*40810*/;
assign _4579_ = D[55] ^ Q[53] /*40806*/;
assign _4576_ = _3904_ & _4579_ /*40802*/;
assign _4577_ = _3904_ ^ _4579_ /*40805*/;
assign _4578_ = _4570_ & _4577_ /*40803*/;
assign _4575_ = _4576_ | _4578_ /*40801*/;
assign _4290_ = _4570_ ^ _4577_ /*40804*/;
assign _4584_ = D[56] ^ Q[53] /*40800*/;
assign _4581_ = _3905_ & _4584_ /*40796*/;
assign _4582_ = _3905_ ^ _4584_ /*40799*/;
assign _4583_ = _4575_ & _4582_ /*40797*/;
assign _4580_ = _4581_ | _4583_ /*40795*/;
assign _4291_ = _4575_ ^ _4582_ /*40798*/;
assign _4589_ = D[57] ^ Q[53] /*40794*/;
assign _4586_ = _3906_ & _4589_ /*40790*/;
assign _4587_ = _3906_ ^ _4589_ /*40793*/;
assign _4588_ = _4580_ & _4587_ /*40791*/;
assign _4585_ = _4586_ | _4588_ /*40789*/;
assign _4292_ = _4580_ ^ _4587_ /*40792*/;
assign _4594_ = D[58] ^ Q[53] /*40788*/;
assign _4591_ = _3907_ & _4594_ /*40784*/;
assign _4592_ = _3907_ ^ _4594_ /*40787*/;
assign _4593_ = _4585_ & _4592_ /*40785*/;
assign _4590_ = _4591_ | _4593_ /*40783*/;
assign _4293_ = _4585_ ^ _4592_ /*40786*/;
assign _4599_ = D[59] ^ Q[53] /*40782*/;
assign _4596_ = _3908_ & _4599_ /*40778*/;
assign _4597_ = _3908_ ^ _4599_ /*40781*/;
assign _4598_ = _4590_ & _4597_ /*40779*/;
assign _4595_ = _4596_ | _4598_ /*40777*/;
assign _4294_ = _4590_ ^ _4597_ /*40780*/;
assign _4604_ = D[60] ^ Q[53] /*40776*/;
assign _4601_ = _3909_ & _4604_ /*40772*/;
assign _4602_ = _3909_ ^ _4604_ /*40775*/;
assign _4603_ = _4595_ & _4602_ /*40773*/;
assign _4600_ = _4601_ | _4603_ /*40771*/;
assign _4295_ = _4595_ ^ _4602_ /*40774*/;
assign _4609_ = D[61] ^ Q[53] /*40770*/;
assign _4606_ = _3910_ & _4609_ /*40766*/;
assign _4607_ = _3910_ ^ _4609_ /*40769*/;
assign _4608_ = _4600_ & _4607_ /*40767*/;
assign _4605_ = _4606_ | _4608_ /*40765*/;
assign _4296_ = _4600_ ^ _4607_ /*40768*/;
assign _4614_ = D[62] ^ Q[53] /*40764*/;
assign _4611_ = _3911_ & _4614_ /*40760*/;
assign _4612_ = _3911_ ^ _4614_ /*40763*/;
assign _4613_ = _4605_ & _4612_ /*40761*/;
assign _4610_ = _4611_ | _4613_ /*40759*/;
assign _4297_ = _4605_ ^ _4612_ /*40762*/;
assign _4618_ = zeroWire ^ Q[53] /*40758*/;
assign _4615_ = _3912_ & _4618_ /*40754*/;
assign _4616_ = _3912_ ^ _4618_ /*40757*/;
assign _4617_ = _4610_ & _4616_ /*40755*/;
assign Q[52] = _4615_ | _4617_ /*40753*/;
assign _4298_ = _4610_ ^ _4616_ /*40756*/;
assign _4689_ = D[0] ^ Q[52] /*40367*/;
assign _4686_ = R_0[51] & _4689_ /*40363*/;
assign _4687_ = R_0[51] ^ _4689_ /*40366*/;
assign _4688_ = Q[52] & _4687_ /*40364*/;
assign _4685_ = _4686_ | _4688_ /*40362*/;
assign _4620_ = Q[52] ^ _4687_ /*40365*/;
assign _4694_ = D[1] ^ Q[52] /*40361*/;
assign _4691_ = _4235_ & _4694_ /*40357*/;
assign _4692_ = _4235_ ^ _4694_ /*40360*/;
assign _4693_ = _4685_ & _4692_ /*40358*/;
assign _4690_ = _4691_ | _4693_ /*40356*/;
assign _4621_ = _4685_ ^ _4692_ /*40359*/;
assign _4699_ = D[2] ^ Q[52] /*40355*/;
assign _4696_ = _4236_ & _4699_ /*40351*/;
assign _4697_ = _4236_ ^ _4699_ /*40354*/;
assign _4698_ = _4690_ & _4697_ /*40352*/;
assign _4695_ = _4696_ | _4698_ /*40350*/;
assign _4622_ = _4690_ ^ _4697_ /*40353*/;
assign _4704_ = D[3] ^ Q[52] /*40349*/;
assign _4701_ = _4237_ & _4704_ /*40345*/;
assign _4702_ = _4237_ ^ _4704_ /*40348*/;
assign _4703_ = _4695_ & _4702_ /*40346*/;
assign _4700_ = _4701_ | _4703_ /*40344*/;
assign _4623_ = _4695_ ^ _4702_ /*40347*/;
assign _4709_ = D[4] ^ Q[52] /*40343*/;
assign _4706_ = _4238_ & _4709_ /*40339*/;
assign _4707_ = _4238_ ^ _4709_ /*40342*/;
assign _4708_ = _4700_ & _4707_ /*40340*/;
assign _4705_ = _4706_ | _4708_ /*40338*/;
assign _4624_ = _4700_ ^ _4707_ /*40341*/;
assign _4714_ = D[5] ^ Q[52] /*40337*/;
assign _4711_ = _4239_ & _4714_ /*40333*/;
assign _4712_ = _4239_ ^ _4714_ /*40336*/;
assign _4713_ = _4705_ & _4712_ /*40334*/;
assign _4710_ = _4711_ | _4713_ /*40332*/;
assign _4625_ = _4705_ ^ _4712_ /*40335*/;
assign _4719_ = D[6] ^ Q[52] /*40331*/;
assign _4716_ = _4240_ & _4719_ /*40327*/;
assign _4717_ = _4240_ ^ _4719_ /*40330*/;
assign _4718_ = _4710_ & _4717_ /*40328*/;
assign _4715_ = _4716_ | _4718_ /*40326*/;
assign _4626_ = _4710_ ^ _4717_ /*40329*/;
assign _4724_ = D[7] ^ Q[52] /*40325*/;
assign _4721_ = _4241_ & _4724_ /*40321*/;
assign _4722_ = _4241_ ^ _4724_ /*40324*/;
assign _4723_ = _4715_ & _4722_ /*40322*/;
assign _4720_ = _4721_ | _4723_ /*40320*/;
assign _4627_ = _4715_ ^ _4722_ /*40323*/;
assign _4729_ = D[8] ^ Q[52] /*40319*/;
assign _4726_ = _4242_ & _4729_ /*40315*/;
assign _4727_ = _4242_ ^ _4729_ /*40318*/;
assign _4728_ = _4720_ & _4727_ /*40316*/;
assign _4725_ = _4726_ | _4728_ /*40314*/;
assign _4628_ = _4720_ ^ _4727_ /*40317*/;
assign _4734_ = D[9] ^ Q[52] /*40313*/;
assign _4731_ = _4243_ & _4734_ /*40309*/;
assign _4732_ = _4243_ ^ _4734_ /*40312*/;
assign _4733_ = _4725_ & _4732_ /*40310*/;
assign _4730_ = _4731_ | _4733_ /*40308*/;
assign _4629_ = _4725_ ^ _4732_ /*40311*/;
assign _4739_ = D[10] ^ Q[52] /*40307*/;
assign _4736_ = _4244_ & _4739_ /*40303*/;
assign _4737_ = _4244_ ^ _4739_ /*40306*/;
assign _4738_ = _4730_ & _4737_ /*40304*/;
assign _4735_ = _4736_ | _4738_ /*40302*/;
assign _4630_ = _4730_ ^ _4737_ /*40305*/;
assign _4744_ = D[11] ^ Q[52] /*40301*/;
assign _4741_ = _4245_ & _4744_ /*40297*/;
assign _4742_ = _4245_ ^ _4744_ /*40300*/;
assign _4743_ = _4735_ & _4742_ /*40298*/;
assign _4740_ = _4741_ | _4743_ /*40296*/;
assign _4631_ = _4735_ ^ _4742_ /*40299*/;
assign _4749_ = D[12] ^ Q[52] /*40295*/;
assign _4746_ = _4246_ & _4749_ /*40291*/;
assign _4747_ = _4246_ ^ _4749_ /*40294*/;
assign _4748_ = _4740_ & _4747_ /*40292*/;
assign _4745_ = _4746_ | _4748_ /*40290*/;
assign _4632_ = _4740_ ^ _4747_ /*40293*/;
assign _4754_ = D[13] ^ Q[52] /*40289*/;
assign _4751_ = _4247_ & _4754_ /*40285*/;
assign _4752_ = _4247_ ^ _4754_ /*40288*/;
assign _4753_ = _4745_ & _4752_ /*40286*/;
assign _4750_ = _4751_ | _4753_ /*40284*/;
assign _4633_ = _4745_ ^ _4752_ /*40287*/;
assign _4759_ = D[14] ^ Q[52] /*40283*/;
assign _4756_ = _4248_ & _4759_ /*40279*/;
assign _4757_ = _4248_ ^ _4759_ /*40282*/;
assign _4758_ = _4750_ & _4757_ /*40280*/;
assign _4755_ = _4756_ | _4758_ /*40278*/;
assign _4634_ = _4750_ ^ _4757_ /*40281*/;
assign _4764_ = D[15] ^ Q[52] /*40277*/;
assign _4761_ = _4249_ & _4764_ /*40273*/;
assign _4762_ = _4249_ ^ _4764_ /*40276*/;
assign _4763_ = _4755_ & _4762_ /*40274*/;
assign _4760_ = _4761_ | _4763_ /*40272*/;
assign _4635_ = _4755_ ^ _4762_ /*40275*/;
assign _4769_ = D[16] ^ Q[52] /*40271*/;
assign _4766_ = _4250_ & _4769_ /*40267*/;
assign _4767_ = _4250_ ^ _4769_ /*40270*/;
assign _4768_ = _4760_ & _4767_ /*40268*/;
assign _4765_ = _4766_ | _4768_ /*40266*/;
assign _4636_ = _4760_ ^ _4767_ /*40269*/;
assign _4774_ = D[17] ^ Q[52] /*40265*/;
assign _4771_ = _4251_ & _4774_ /*40261*/;
assign _4772_ = _4251_ ^ _4774_ /*40264*/;
assign _4773_ = _4765_ & _4772_ /*40262*/;
assign _4770_ = _4771_ | _4773_ /*40260*/;
assign _4637_ = _4765_ ^ _4772_ /*40263*/;
assign _4779_ = D[18] ^ Q[52] /*40259*/;
assign _4776_ = _4252_ & _4779_ /*40255*/;
assign _4777_ = _4252_ ^ _4779_ /*40258*/;
assign _4778_ = _4770_ & _4777_ /*40256*/;
assign _4775_ = _4776_ | _4778_ /*40254*/;
assign _4638_ = _4770_ ^ _4777_ /*40257*/;
assign _4784_ = D[19] ^ Q[52] /*40253*/;
assign _4781_ = _4253_ & _4784_ /*40249*/;
assign _4782_ = _4253_ ^ _4784_ /*40252*/;
assign _4783_ = _4775_ & _4782_ /*40250*/;
assign _4780_ = _4781_ | _4783_ /*40248*/;
assign _4639_ = _4775_ ^ _4782_ /*40251*/;
assign _4789_ = D[20] ^ Q[52] /*40247*/;
assign _4786_ = _4254_ & _4789_ /*40243*/;
assign _4787_ = _4254_ ^ _4789_ /*40246*/;
assign _4788_ = _4780_ & _4787_ /*40244*/;
assign _4785_ = _4786_ | _4788_ /*40242*/;
assign _4640_ = _4780_ ^ _4787_ /*40245*/;
assign _4794_ = D[21] ^ Q[52] /*40241*/;
assign _4791_ = _4255_ & _4794_ /*40237*/;
assign _4792_ = _4255_ ^ _4794_ /*40240*/;
assign _4793_ = _4785_ & _4792_ /*40238*/;
assign _4790_ = _4791_ | _4793_ /*40236*/;
assign _4641_ = _4785_ ^ _4792_ /*40239*/;
assign _4799_ = D[22] ^ Q[52] /*40235*/;
assign _4796_ = _4256_ & _4799_ /*40231*/;
assign _4797_ = _4256_ ^ _4799_ /*40234*/;
assign _4798_ = _4790_ & _4797_ /*40232*/;
assign _4795_ = _4796_ | _4798_ /*40230*/;
assign _4642_ = _4790_ ^ _4797_ /*40233*/;
assign _4804_ = D[23] ^ Q[52] /*40229*/;
assign _4801_ = _4257_ & _4804_ /*40225*/;
assign _4802_ = _4257_ ^ _4804_ /*40228*/;
assign _4803_ = _4795_ & _4802_ /*40226*/;
assign _4800_ = _4801_ | _4803_ /*40224*/;
assign _4643_ = _4795_ ^ _4802_ /*40227*/;
assign _4809_ = D[24] ^ Q[52] /*40223*/;
assign _4806_ = _4258_ & _4809_ /*40219*/;
assign _4807_ = _4258_ ^ _4809_ /*40222*/;
assign _4808_ = _4800_ & _4807_ /*40220*/;
assign _4805_ = _4806_ | _4808_ /*40218*/;
assign _4644_ = _4800_ ^ _4807_ /*40221*/;
assign _4814_ = D[25] ^ Q[52] /*40217*/;
assign _4811_ = _4259_ & _4814_ /*40213*/;
assign _4812_ = _4259_ ^ _4814_ /*40216*/;
assign _4813_ = _4805_ & _4812_ /*40214*/;
assign _4810_ = _4811_ | _4813_ /*40212*/;
assign _4645_ = _4805_ ^ _4812_ /*40215*/;
assign _4819_ = D[26] ^ Q[52] /*40211*/;
assign _4816_ = _4260_ & _4819_ /*40207*/;
assign _4817_ = _4260_ ^ _4819_ /*40210*/;
assign _4818_ = _4810_ & _4817_ /*40208*/;
assign _4815_ = _4816_ | _4818_ /*40206*/;
assign _4646_ = _4810_ ^ _4817_ /*40209*/;
assign _4824_ = D[27] ^ Q[52] /*40205*/;
assign _4821_ = _4261_ & _4824_ /*40201*/;
assign _4822_ = _4261_ ^ _4824_ /*40204*/;
assign _4823_ = _4815_ & _4822_ /*40202*/;
assign _4820_ = _4821_ | _4823_ /*40200*/;
assign _4647_ = _4815_ ^ _4822_ /*40203*/;
assign _4829_ = D[28] ^ Q[52] /*40199*/;
assign _4826_ = _4262_ & _4829_ /*40195*/;
assign _4827_ = _4262_ ^ _4829_ /*40198*/;
assign _4828_ = _4820_ & _4827_ /*40196*/;
assign _4825_ = _4826_ | _4828_ /*40194*/;
assign _4648_ = _4820_ ^ _4827_ /*40197*/;
assign _4834_ = D[29] ^ Q[52] /*40193*/;
assign _4831_ = _4263_ & _4834_ /*40189*/;
assign _4832_ = _4263_ ^ _4834_ /*40192*/;
assign _4833_ = _4825_ & _4832_ /*40190*/;
assign _4830_ = _4831_ | _4833_ /*40188*/;
assign _4649_ = _4825_ ^ _4832_ /*40191*/;
assign _4839_ = D[30] ^ Q[52] /*40187*/;
assign _4836_ = _4264_ & _4839_ /*40183*/;
assign _4837_ = _4264_ ^ _4839_ /*40186*/;
assign _4838_ = _4830_ & _4837_ /*40184*/;
assign _4835_ = _4836_ | _4838_ /*40182*/;
assign _4650_ = _4830_ ^ _4837_ /*40185*/;
assign _4844_ = D[31] ^ Q[52] /*40181*/;
assign _4841_ = _4265_ & _4844_ /*40177*/;
assign _4842_ = _4265_ ^ _4844_ /*40180*/;
assign _4843_ = _4835_ & _4842_ /*40178*/;
assign _4840_ = _4841_ | _4843_ /*40176*/;
assign _4651_ = _4835_ ^ _4842_ /*40179*/;
assign _4849_ = D[32] ^ Q[52] /*40175*/;
assign _4846_ = _4266_ & _4849_ /*40171*/;
assign _4847_ = _4266_ ^ _4849_ /*40174*/;
assign _4848_ = _4840_ & _4847_ /*40172*/;
assign _4845_ = _4846_ | _4848_ /*40170*/;
assign _4652_ = _4840_ ^ _4847_ /*40173*/;
assign _4854_ = D[33] ^ Q[52] /*40169*/;
assign _4851_ = _4267_ & _4854_ /*40165*/;
assign _4852_ = _4267_ ^ _4854_ /*40168*/;
assign _4853_ = _4845_ & _4852_ /*40166*/;
assign _4850_ = _4851_ | _4853_ /*40164*/;
assign _4653_ = _4845_ ^ _4852_ /*40167*/;
assign _4859_ = D[34] ^ Q[52] /*40163*/;
assign _4856_ = _4268_ & _4859_ /*40159*/;
assign _4857_ = _4268_ ^ _4859_ /*40162*/;
assign _4858_ = _4850_ & _4857_ /*40160*/;
assign _4855_ = _4856_ | _4858_ /*40158*/;
assign _4654_ = _4850_ ^ _4857_ /*40161*/;
assign _4864_ = D[35] ^ Q[52] /*40157*/;
assign _4861_ = _4269_ & _4864_ /*40153*/;
assign _4862_ = _4269_ ^ _4864_ /*40156*/;
assign _4863_ = _4855_ & _4862_ /*40154*/;
assign _4860_ = _4861_ | _4863_ /*40152*/;
assign _4655_ = _4855_ ^ _4862_ /*40155*/;
assign _4869_ = D[36] ^ Q[52] /*40151*/;
assign _4866_ = _4270_ & _4869_ /*40147*/;
assign _4867_ = _4270_ ^ _4869_ /*40150*/;
assign _4868_ = _4860_ & _4867_ /*40148*/;
assign _4865_ = _4866_ | _4868_ /*40146*/;
assign _4656_ = _4860_ ^ _4867_ /*40149*/;
assign _4874_ = D[37] ^ Q[52] /*40145*/;
assign _4871_ = _4271_ & _4874_ /*40141*/;
assign _4872_ = _4271_ ^ _4874_ /*40144*/;
assign _4873_ = _4865_ & _4872_ /*40142*/;
assign _4870_ = _4871_ | _4873_ /*40140*/;
assign _4657_ = _4865_ ^ _4872_ /*40143*/;
assign _4879_ = D[38] ^ Q[52] /*40139*/;
assign _4876_ = _4272_ & _4879_ /*40135*/;
assign _4877_ = _4272_ ^ _4879_ /*40138*/;
assign _4878_ = _4870_ & _4877_ /*40136*/;
assign _4875_ = _4876_ | _4878_ /*40134*/;
assign _4658_ = _4870_ ^ _4877_ /*40137*/;
assign _4884_ = D[39] ^ Q[52] /*40133*/;
assign _4881_ = _4273_ & _4884_ /*40129*/;
assign _4882_ = _4273_ ^ _4884_ /*40132*/;
assign _4883_ = _4875_ & _4882_ /*40130*/;
assign _4880_ = _4881_ | _4883_ /*40128*/;
assign _4659_ = _4875_ ^ _4882_ /*40131*/;
assign _4889_ = D[40] ^ Q[52] /*40127*/;
assign _4886_ = _4274_ & _4889_ /*40123*/;
assign _4887_ = _4274_ ^ _4889_ /*40126*/;
assign _4888_ = _4880_ & _4887_ /*40124*/;
assign _4885_ = _4886_ | _4888_ /*40122*/;
assign _4660_ = _4880_ ^ _4887_ /*40125*/;
assign _4894_ = D[41] ^ Q[52] /*40121*/;
assign _4891_ = _4275_ & _4894_ /*40117*/;
assign _4892_ = _4275_ ^ _4894_ /*40120*/;
assign _4893_ = _4885_ & _4892_ /*40118*/;
assign _4890_ = _4891_ | _4893_ /*40116*/;
assign _4661_ = _4885_ ^ _4892_ /*40119*/;
assign _4899_ = D[42] ^ Q[52] /*40115*/;
assign _4896_ = _4276_ & _4899_ /*40111*/;
assign _4897_ = _4276_ ^ _4899_ /*40114*/;
assign _4898_ = _4890_ & _4897_ /*40112*/;
assign _4895_ = _4896_ | _4898_ /*40110*/;
assign _4662_ = _4890_ ^ _4897_ /*40113*/;
assign _4904_ = D[43] ^ Q[52] /*40109*/;
assign _4901_ = _4277_ & _4904_ /*40105*/;
assign _4902_ = _4277_ ^ _4904_ /*40108*/;
assign _4903_ = _4895_ & _4902_ /*40106*/;
assign _4900_ = _4901_ | _4903_ /*40104*/;
assign _4663_ = _4895_ ^ _4902_ /*40107*/;
assign _4909_ = D[44] ^ Q[52] /*40103*/;
assign _4906_ = _4278_ & _4909_ /*40099*/;
assign _4907_ = _4278_ ^ _4909_ /*40102*/;
assign _4908_ = _4900_ & _4907_ /*40100*/;
assign _4905_ = _4906_ | _4908_ /*40098*/;
assign _4664_ = _4900_ ^ _4907_ /*40101*/;
assign _4914_ = D[45] ^ Q[52] /*40097*/;
assign _4911_ = _4279_ & _4914_ /*40093*/;
assign _4912_ = _4279_ ^ _4914_ /*40096*/;
assign _4913_ = _4905_ & _4912_ /*40094*/;
assign _4910_ = _4911_ | _4913_ /*40092*/;
assign _4665_ = _4905_ ^ _4912_ /*40095*/;
assign _4919_ = D[46] ^ Q[52] /*40091*/;
assign _4916_ = _4280_ & _4919_ /*40087*/;
assign _4917_ = _4280_ ^ _4919_ /*40090*/;
assign _4918_ = _4910_ & _4917_ /*40088*/;
assign _4915_ = _4916_ | _4918_ /*40086*/;
assign _4666_ = _4910_ ^ _4917_ /*40089*/;
assign _4924_ = D[47] ^ Q[52] /*40085*/;
assign _4921_ = _4281_ & _4924_ /*40081*/;
assign _4922_ = _4281_ ^ _4924_ /*40084*/;
assign _4923_ = _4915_ & _4922_ /*40082*/;
assign _4920_ = _4921_ | _4923_ /*40080*/;
assign _4667_ = _4915_ ^ _4922_ /*40083*/;
assign _4929_ = D[48] ^ Q[52] /*40079*/;
assign _4926_ = _4282_ & _4929_ /*40075*/;
assign _4927_ = _4282_ ^ _4929_ /*40078*/;
assign _4928_ = _4920_ & _4927_ /*40076*/;
assign _4925_ = _4926_ | _4928_ /*40074*/;
assign _4668_ = _4920_ ^ _4927_ /*40077*/;
assign _4934_ = D[49] ^ Q[52] /*40073*/;
assign _4931_ = _4283_ & _4934_ /*40069*/;
assign _4932_ = _4283_ ^ _4934_ /*40072*/;
assign _4933_ = _4925_ & _4932_ /*40070*/;
assign _4930_ = _4931_ | _4933_ /*40068*/;
assign _4669_ = _4925_ ^ _4932_ /*40071*/;
assign _4939_ = D[50] ^ Q[52] /*40067*/;
assign _4936_ = _4284_ & _4939_ /*40063*/;
assign _4937_ = _4284_ ^ _4939_ /*40066*/;
assign _4938_ = _4930_ & _4937_ /*40064*/;
assign _4935_ = _4936_ | _4938_ /*40062*/;
assign _4670_ = _4930_ ^ _4937_ /*40065*/;
assign _4944_ = D[51] ^ Q[52] /*40061*/;
assign _4941_ = _4285_ & _4944_ /*40057*/;
assign _4942_ = _4285_ ^ _4944_ /*40060*/;
assign _4943_ = _4935_ & _4942_ /*40058*/;
assign _4940_ = _4941_ | _4943_ /*40056*/;
assign _4671_ = _4935_ ^ _4942_ /*40059*/;
assign _4949_ = D[52] ^ Q[52] /*40055*/;
assign _4946_ = _4286_ & _4949_ /*40051*/;
assign _4947_ = _4286_ ^ _4949_ /*40054*/;
assign _4948_ = _4940_ & _4947_ /*40052*/;
assign _4945_ = _4946_ | _4948_ /*40050*/;
assign _4672_ = _4940_ ^ _4947_ /*40053*/;
assign _4954_ = D[53] ^ Q[52] /*40049*/;
assign _4951_ = _4287_ & _4954_ /*40045*/;
assign _4952_ = _4287_ ^ _4954_ /*40048*/;
assign _4953_ = _4945_ & _4952_ /*40046*/;
assign _4950_ = _4951_ | _4953_ /*40044*/;
assign _4673_ = _4945_ ^ _4952_ /*40047*/;
assign _4959_ = D[54] ^ Q[52] /*40043*/;
assign _4956_ = _4288_ & _4959_ /*40039*/;
assign _4957_ = _4288_ ^ _4959_ /*40042*/;
assign _4958_ = _4950_ & _4957_ /*40040*/;
assign _4955_ = _4956_ | _4958_ /*40038*/;
assign _4674_ = _4950_ ^ _4957_ /*40041*/;
assign _4964_ = D[55] ^ Q[52] /*40037*/;
assign _4961_ = _4289_ & _4964_ /*40033*/;
assign _4962_ = _4289_ ^ _4964_ /*40036*/;
assign _4963_ = _4955_ & _4962_ /*40034*/;
assign _4960_ = _4961_ | _4963_ /*40032*/;
assign _4675_ = _4955_ ^ _4962_ /*40035*/;
assign _4969_ = D[56] ^ Q[52] /*40031*/;
assign _4966_ = _4290_ & _4969_ /*40027*/;
assign _4967_ = _4290_ ^ _4969_ /*40030*/;
assign _4968_ = _4960_ & _4967_ /*40028*/;
assign _4965_ = _4966_ | _4968_ /*40026*/;
assign _4676_ = _4960_ ^ _4967_ /*40029*/;
assign _4974_ = D[57] ^ Q[52] /*40025*/;
assign _4971_ = _4291_ & _4974_ /*40021*/;
assign _4972_ = _4291_ ^ _4974_ /*40024*/;
assign _4973_ = _4965_ & _4972_ /*40022*/;
assign _4970_ = _4971_ | _4973_ /*40020*/;
assign _4677_ = _4965_ ^ _4972_ /*40023*/;
assign _4979_ = D[58] ^ Q[52] /*40019*/;
assign _4976_ = _4292_ & _4979_ /*40015*/;
assign _4977_ = _4292_ ^ _4979_ /*40018*/;
assign _4978_ = _4970_ & _4977_ /*40016*/;
assign _4975_ = _4976_ | _4978_ /*40014*/;
assign _4678_ = _4970_ ^ _4977_ /*40017*/;
assign _4984_ = D[59] ^ Q[52] /*40013*/;
assign _4981_ = _4293_ & _4984_ /*40009*/;
assign _4982_ = _4293_ ^ _4984_ /*40012*/;
assign _4983_ = _4975_ & _4982_ /*40010*/;
assign _4980_ = _4981_ | _4983_ /*40008*/;
assign _4679_ = _4975_ ^ _4982_ /*40011*/;
assign _4989_ = D[60] ^ Q[52] /*40007*/;
assign _4986_ = _4294_ & _4989_ /*40003*/;
assign _4987_ = _4294_ ^ _4989_ /*40006*/;
assign _4988_ = _4980_ & _4987_ /*40004*/;
assign _4985_ = _4986_ | _4988_ /*40002*/;
assign _4680_ = _4980_ ^ _4987_ /*40005*/;
assign _4994_ = D[61] ^ Q[52] /*40001*/;
assign _4991_ = _4295_ & _4994_ /*39997*/;
assign _4992_ = _4295_ ^ _4994_ /*40000*/;
assign _4993_ = _4985_ & _4992_ /*39998*/;
assign _4990_ = _4991_ | _4993_ /*39996*/;
assign _4681_ = _4985_ ^ _4992_ /*39999*/;
assign _4999_ = D[62] ^ Q[52] /*39995*/;
assign _4996_ = _4296_ & _4999_ /*39991*/;
assign _4997_ = _4296_ ^ _4999_ /*39994*/;
assign _4998_ = _4990_ & _4997_ /*39992*/;
assign _4995_ = _4996_ | _4998_ /*39990*/;
assign _4682_ = _4990_ ^ _4997_ /*39993*/;
assign _5003_ = zeroWire ^ Q[52] /*39989*/;
assign _5000_ = _4297_ & _5003_ /*39985*/;
assign _5001_ = _4297_ ^ _5003_ /*39988*/;
assign _5002_ = _4995_ & _5001_ /*39986*/;
assign Q[51] = _5000_ | _5002_ /*39984*/;
assign _4683_ = _4995_ ^ _5001_ /*39987*/;
assign _5074_ = D[0] ^ Q[51] /*39598*/;
assign _5071_ = R_0[50] & _5074_ /*39594*/;
assign _5072_ = R_0[50] ^ _5074_ /*39597*/;
assign _5073_ = Q[51] & _5072_ /*39595*/;
assign _5070_ = _5071_ | _5073_ /*39593*/;
assign _5005_ = Q[51] ^ _5072_ /*39596*/;
assign _5079_ = D[1] ^ Q[51] /*39592*/;
assign _5076_ = _4620_ & _5079_ /*39588*/;
assign _5077_ = _4620_ ^ _5079_ /*39591*/;
assign _5078_ = _5070_ & _5077_ /*39589*/;
assign _5075_ = _5076_ | _5078_ /*39587*/;
assign _5006_ = _5070_ ^ _5077_ /*39590*/;
assign _5084_ = D[2] ^ Q[51] /*39586*/;
assign _5081_ = _4621_ & _5084_ /*39582*/;
assign _5082_ = _4621_ ^ _5084_ /*39585*/;
assign _5083_ = _5075_ & _5082_ /*39583*/;
assign _5080_ = _5081_ | _5083_ /*39581*/;
assign _5007_ = _5075_ ^ _5082_ /*39584*/;
assign _5089_ = D[3] ^ Q[51] /*39580*/;
assign _5086_ = _4622_ & _5089_ /*39576*/;
assign _5087_ = _4622_ ^ _5089_ /*39579*/;
assign _5088_ = _5080_ & _5087_ /*39577*/;
assign _5085_ = _5086_ | _5088_ /*39575*/;
assign _5008_ = _5080_ ^ _5087_ /*39578*/;
assign _5094_ = D[4] ^ Q[51] /*39574*/;
assign _5091_ = _4623_ & _5094_ /*39570*/;
assign _5092_ = _4623_ ^ _5094_ /*39573*/;
assign _5093_ = _5085_ & _5092_ /*39571*/;
assign _5090_ = _5091_ | _5093_ /*39569*/;
assign _5009_ = _5085_ ^ _5092_ /*39572*/;
assign _5099_ = D[5] ^ Q[51] /*39568*/;
assign _5096_ = _4624_ & _5099_ /*39564*/;
assign _5097_ = _4624_ ^ _5099_ /*39567*/;
assign _5098_ = _5090_ & _5097_ /*39565*/;
assign _5095_ = _5096_ | _5098_ /*39563*/;
assign _5010_ = _5090_ ^ _5097_ /*39566*/;
assign _5104_ = D[6] ^ Q[51] /*39562*/;
assign _5101_ = _4625_ & _5104_ /*39558*/;
assign _5102_ = _4625_ ^ _5104_ /*39561*/;
assign _5103_ = _5095_ & _5102_ /*39559*/;
assign _5100_ = _5101_ | _5103_ /*39557*/;
assign _5011_ = _5095_ ^ _5102_ /*39560*/;
assign _5109_ = D[7] ^ Q[51] /*39556*/;
assign _5106_ = _4626_ & _5109_ /*39552*/;
assign _5107_ = _4626_ ^ _5109_ /*39555*/;
assign _5108_ = _5100_ & _5107_ /*39553*/;
assign _5105_ = _5106_ | _5108_ /*39551*/;
assign _5012_ = _5100_ ^ _5107_ /*39554*/;
assign _5114_ = D[8] ^ Q[51] /*39550*/;
assign _5111_ = _4627_ & _5114_ /*39546*/;
assign _5112_ = _4627_ ^ _5114_ /*39549*/;
assign _5113_ = _5105_ & _5112_ /*39547*/;
assign _5110_ = _5111_ | _5113_ /*39545*/;
assign _5013_ = _5105_ ^ _5112_ /*39548*/;
assign _5119_ = D[9] ^ Q[51] /*39544*/;
assign _5116_ = _4628_ & _5119_ /*39540*/;
assign _5117_ = _4628_ ^ _5119_ /*39543*/;
assign _5118_ = _5110_ & _5117_ /*39541*/;
assign _5115_ = _5116_ | _5118_ /*39539*/;
assign _5014_ = _5110_ ^ _5117_ /*39542*/;
assign _5124_ = D[10] ^ Q[51] /*39538*/;
assign _5121_ = _4629_ & _5124_ /*39534*/;
assign _5122_ = _4629_ ^ _5124_ /*39537*/;
assign _5123_ = _5115_ & _5122_ /*39535*/;
assign _5120_ = _5121_ | _5123_ /*39533*/;
assign _5015_ = _5115_ ^ _5122_ /*39536*/;
assign _5129_ = D[11] ^ Q[51] /*39532*/;
assign _5126_ = _4630_ & _5129_ /*39528*/;
assign _5127_ = _4630_ ^ _5129_ /*39531*/;
assign _5128_ = _5120_ & _5127_ /*39529*/;
assign _5125_ = _5126_ | _5128_ /*39527*/;
assign _5016_ = _5120_ ^ _5127_ /*39530*/;
assign _5134_ = D[12] ^ Q[51] /*39526*/;
assign _5131_ = _4631_ & _5134_ /*39522*/;
assign _5132_ = _4631_ ^ _5134_ /*39525*/;
assign _5133_ = _5125_ & _5132_ /*39523*/;
assign _5130_ = _5131_ | _5133_ /*39521*/;
assign _5017_ = _5125_ ^ _5132_ /*39524*/;
assign _5139_ = D[13] ^ Q[51] /*39520*/;
assign _5136_ = _4632_ & _5139_ /*39516*/;
assign _5137_ = _4632_ ^ _5139_ /*39519*/;
assign _5138_ = _5130_ & _5137_ /*39517*/;
assign _5135_ = _5136_ | _5138_ /*39515*/;
assign _5018_ = _5130_ ^ _5137_ /*39518*/;
assign _5144_ = D[14] ^ Q[51] /*39514*/;
assign _5141_ = _4633_ & _5144_ /*39510*/;
assign _5142_ = _4633_ ^ _5144_ /*39513*/;
assign _5143_ = _5135_ & _5142_ /*39511*/;
assign _5140_ = _5141_ | _5143_ /*39509*/;
assign _5019_ = _5135_ ^ _5142_ /*39512*/;
assign _5149_ = D[15] ^ Q[51] /*39508*/;
assign _5146_ = _4634_ & _5149_ /*39504*/;
assign _5147_ = _4634_ ^ _5149_ /*39507*/;
assign _5148_ = _5140_ & _5147_ /*39505*/;
assign _5145_ = _5146_ | _5148_ /*39503*/;
assign _5020_ = _5140_ ^ _5147_ /*39506*/;
assign _5154_ = D[16] ^ Q[51] /*39502*/;
assign _5151_ = _4635_ & _5154_ /*39498*/;
assign _5152_ = _4635_ ^ _5154_ /*39501*/;
assign _5153_ = _5145_ & _5152_ /*39499*/;
assign _5150_ = _5151_ | _5153_ /*39497*/;
assign _5021_ = _5145_ ^ _5152_ /*39500*/;
assign _5159_ = D[17] ^ Q[51] /*39496*/;
assign _5156_ = _4636_ & _5159_ /*39492*/;
assign _5157_ = _4636_ ^ _5159_ /*39495*/;
assign _5158_ = _5150_ & _5157_ /*39493*/;
assign _5155_ = _5156_ | _5158_ /*39491*/;
assign _5022_ = _5150_ ^ _5157_ /*39494*/;
assign _5164_ = D[18] ^ Q[51] /*39490*/;
assign _5161_ = _4637_ & _5164_ /*39486*/;
assign _5162_ = _4637_ ^ _5164_ /*39489*/;
assign _5163_ = _5155_ & _5162_ /*39487*/;
assign _5160_ = _5161_ | _5163_ /*39485*/;
assign _5023_ = _5155_ ^ _5162_ /*39488*/;
assign _5169_ = D[19] ^ Q[51] /*39484*/;
assign _5166_ = _4638_ & _5169_ /*39480*/;
assign _5167_ = _4638_ ^ _5169_ /*39483*/;
assign _5168_ = _5160_ & _5167_ /*39481*/;
assign _5165_ = _5166_ | _5168_ /*39479*/;
assign _5024_ = _5160_ ^ _5167_ /*39482*/;
assign _5174_ = D[20] ^ Q[51] /*39478*/;
assign _5171_ = _4639_ & _5174_ /*39474*/;
assign _5172_ = _4639_ ^ _5174_ /*39477*/;
assign _5173_ = _5165_ & _5172_ /*39475*/;
assign _5170_ = _5171_ | _5173_ /*39473*/;
assign _5025_ = _5165_ ^ _5172_ /*39476*/;
assign _5179_ = D[21] ^ Q[51] /*39472*/;
assign _5176_ = _4640_ & _5179_ /*39468*/;
assign _5177_ = _4640_ ^ _5179_ /*39471*/;
assign _5178_ = _5170_ & _5177_ /*39469*/;
assign _5175_ = _5176_ | _5178_ /*39467*/;
assign _5026_ = _5170_ ^ _5177_ /*39470*/;
assign _5184_ = D[22] ^ Q[51] /*39466*/;
assign _5181_ = _4641_ & _5184_ /*39462*/;
assign _5182_ = _4641_ ^ _5184_ /*39465*/;
assign _5183_ = _5175_ & _5182_ /*39463*/;
assign _5180_ = _5181_ | _5183_ /*39461*/;
assign _5027_ = _5175_ ^ _5182_ /*39464*/;
assign _5189_ = D[23] ^ Q[51] /*39460*/;
assign _5186_ = _4642_ & _5189_ /*39456*/;
assign _5187_ = _4642_ ^ _5189_ /*39459*/;
assign _5188_ = _5180_ & _5187_ /*39457*/;
assign _5185_ = _5186_ | _5188_ /*39455*/;
assign _5028_ = _5180_ ^ _5187_ /*39458*/;
assign _5194_ = D[24] ^ Q[51] /*39454*/;
assign _5191_ = _4643_ & _5194_ /*39450*/;
assign _5192_ = _4643_ ^ _5194_ /*39453*/;
assign _5193_ = _5185_ & _5192_ /*39451*/;
assign _5190_ = _5191_ | _5193_ /*39449*/;
assign _5029_ = _5185_ ^ _5192_ /*39452*/;
assign _5199_ = D[25] ^ Q[51] /*39448*/;
assign _5196_ = _4644_ & _5199_ /*39444*/;
assign _5197_ = _4644_ ^ _5199_ /*39447*/;
assign _5198_ = _5190_ & _5197_ /*39445*/;
assign _5195_ = _5196_ | _5198_ /*39443*/;
assign _5030_ = _5190_ ^ _5197_ /*39446*/;
assign _5204_ = D[26] ^ Q[51] /*39442*/;
assign _5201_ = _4645_ & _5204_ /*39438*/;
assign _5202_ = _4645_ ^ _5204_ /*39441*/;
assign _5203_ = _5195_ & _5202_ /*39439*/;
assign _5200_ = _5201_ | _5203_ /*39437*/;
assign _5031_ = _5195_ ^ _5202_ /*39440*/;
assign _5209_ = D[27] ^ Q[51] /*39436*/;
assign _5206_ = _4646_ & _5209_ /*39432*/;
assign _5207_ = _4646_ ^ _5209_ /*39435*/;
assign _5208_ = _5200_ & _5207_ /*39433*/;
assign _5205_ = _5206_ | _5208_ /*39431*/;
assign _5032_ = _5200_ ^ _5207_ /*39434*/;
assign _5214_ = D[28] ^ Q[51] /*39430*/;
assign _5211_ = _4647_ & _5214_ /*39426*/;
assign _5212_ = _4647_ ^ _5214_ /*39429*/;
assign _5213_ = _5205_ & _5212_ /*39427*/;
assign _5210_ = _5211_ | _5213_ /*39425*/;
assign _5033_ = _5205_ ^ _5212_ /*39428*/;
assign _5219_ = D[29] ^ Q[51] /*39424*/;
assign _5216_ = _4648_ & _5219_ /*39420*/;
assign _5217_ = _4648_ ^ _5219_ /*39423*/;
assign _5218_ = _5210_ & _5217_ /*39421*/;
assign _5215_ = _5216_ | _5218_ /*39419*/;
assign _5034_ = _5210_ ^ _5217_ /*39422*/;
assign _5224_ = D[30] ^ Q[51] /*39418*/;
assign _5221_ = _4649_ & _5224_ /*39414*/;
assign _5222_ = _4649_ ^ _5224_ /*39417*/;
assign _5223_ = _5215_ & _5222_ /*39415*/;
assign _5220_ = _5221_ | _5223_ /*39413*/;
assign _5035_ = _5215_ ^ _5222_ /*39416*/;
assign _5229_ = D[31] ^ Q[51] /*39412*/;
assign _5226_ = _4650_ & _5229_ /*39408*/;
assign _5227_ = _4650_ ^ _5229_ /*39411*/;
assign _5228_ = _5220_ & _5227_ /*39409*/;
assign _5225_ = _5226_ | _5228_ /*39407*/;
assign _5036_ = _5220_ ^ _5227_ /*39410*/;
assign _5234_ = D[32] ^ Q[51] /*39406*/;
assign _5231_ = _4651_ & _5234_ /*39402*/;
assign _5232_ = _4651_ ^ _5234_ /*39405*/;
assign _5233_ = _5225_ & _5232_ /*39403*/;
assign _5230_ = _5231_ | _5233_ /*39401*/;
assign _5037_ = _5225_ ^ _5232_ /*39404*/;
assign _5239_ = D[33] ^ Q[51] /*39400*/;
assign _5236_ = _4652_ & _5239_ /*39396*/;
assign _5237_ = _4652_ ^ _5239_ /*39399*/;
assign _5238_ = _5230_ & _5237_ /*39397*/;
assign _5235_ = _5236_ | _5238_ /*39395*/;
assign _5038_ = _5230_ ^ _5237_ /*39398*/;
assign _5244_ = D[34] ^ Q[51] /*39394*/;
assign _5241_ = _4653_ & _5244_ /*39390*/;
assign _5242_ = _4653_ ^ _5244_ /*39393*/;
assign _5243_ = _5235_ & _5242_ /*39391*/;
assign _5240_ = _5241_ | _5243_ /*39389*/;
assign _5039_ = _5235_ ^ _5242_ /*39392*/;
assign _5249_ = D[35] ^ Q[51] /*39388*/;
assign _5246_ = _4654_ & _5249_ /*39384*/;
assign _5247_ = _4654_ ^ _5249_ /*39387*/;
assign _5248_ = _5240_ & _5247_ /*39385*/;
assign _5245_ = _5246_ | _5248_ /*39383*/;
assign _5040_ = _5240_ ^ _5247_ /*39386*/;
assign _5254_ = D[36] ^ Q[51] /*39382*/;
assign _5251_ = _4655_ & _5254_ /*39378*/;
assign _5252_ = _4655_ ^ _5254_ /*39381*/;
assign _5253_ = _5245_ & _5252_ /*39379*/;
assign _5250_ = _5251_ | _5253_ /*39377*/;
assign _5041_ = _5245_ ^ _5252_ /*39380*/;
assign _5259_ = D[37] ^ Q[51] /*39376*/;
assign _5256_ = _4656_ & _5259_ /*39372*/;
assign _5257_ = _4656_ ^ _5259_ /*39375*/;
assign _5258_ = _5250_ & _5257_ /*39373*/;
assign _5255_ = _5256_ | _5258_ /*39371*/;
assign _5042_ = _5250_ ^ _5257_ /*39374*/;
assign _5264_ = D[38] ^ Q[51] /*39370*/;
assign _5261_ = _4657_ & _5264_ /*39366*/;
assign _5262_ = _4657_ ^ _5264_ /*39369*/;
assign _5263_ = _5255_ & _5262_ /*39367*/;
assign _5260_ = _5261_ | _5263_ /*39365*/;
assign _5043_ = _5255_ ^ _5262_ /*39368*/;
assign _5269_ = D[39] ^ Q[51] /*39364*/;
assign _5266_ = _4658_ & _5269_ /*39360*/;
assign _5267_ = _4658_ ^ _5269_ /*39363*/;
assign _5268_ = _5260_ & _5267_ /*39361*/;
assign _5265_ = _5266_ | _5268_ /*39359*/;
assign _5044_ = _5260_ ^ _5267_ /*39362*/;
assign _5274_ = D[40] ^ Q[51] /*39358*/;
assign _5271_ = _4659_ & _5274_ /*39354*/;
assign _5272_ = _4659_ ^ _5274_ /*39357*/;
assign _5273_ = _5265_ & _5272_ /*39355*/;
assign _5270_ = _5271_ | _5273_ /*39353*/;
assign _5045_ = _5265_ ^ _5272_ /*39356*/;
assign _5279_ = D[41] ^ Q[51] /*39352*/;
assign _5276_ = _4660_ & _5279_ /*39348*/;
assign _5277_ = _4660_ ^ _5279_ /*39351*/;
assign _5278_ = _5270_ & _5277_ /*39349*/;
assign _5275_ = _5276_ | _5278_ /*39347*/;
assign _5046_ = _5270_ ^ _5277_ /*39350*/;
assign _5284_ = D[42] ^ Q[51] /*39346*/;
assign _5281_ = _4661_ & _5284_ /*39342*/;
assign _5282_ = _4661_ ^ _5284_ /*39345*/;
assign _5283_ = _5275_ & _5282_ /*39343*/;
assign _5280_ = _5281_ | _5283_ /*39341*/;
assign _5047_ = _5275_ ^ _5282_ /*39344*/;
assign _5289_ = D[43] ^ Q[51] /*39340*/;
assign _5286_ = _4662_ & _5289_ /*39336*/;
assign _5287_ = _4662_ ^ _5289_ /*39339*/;
assign _5288_ = _5280_ & _5287_ /*39337*/;
assign _5285_ = _5286_ | _5288_ /*39335*/;
assign _5048_ = _5280_ ^ _5287_ /*39338*/;
assign _5294_ = D[44] ^ Q[51] /*39334*/;
assign _5291_ = _4663_ & _5294_ /*39330*/;
assign _5292_ = _4663_ ^ _5294_ /*39333*/;
assign _5293_ = _5285_ & _5292_ /*39331*/;
assign _5290_ = _5291_ | _5293_ /*39329*/;
assign _5049_ = _5285_ ^ _5292_ /*39332*/;
assign _5299_ = D[45] ^ Q[51] /*39328*/;
assign _5296_ = _4664_ & _5299_ /*39324*/;
assign _5297_ = _4664_ ^ _5299_ /*39327*/;
assign _5298_ = _5290_ & _5297_ /*39325*/;
assign _5295_ = _5296_ | _5298_ /*39323*/;
assign _5050_ = _5290_ ^ _5297_ /*39326*/;
assign _5304_ = D[46] ^ Q[51] /*39322*/;
assign _5301_ = _4665_ & _5304_ /*39318*/;
assign _5302_ = _4665_ ^ _5304_ /*39321*/;
assign _5303_ = _5295_ & _5302_ /*39319*/;
assign _5300_ = _5301_ | _5303_ /*39317*/;
assign _5051_ = _5295_ ^ _5302_ /*39320*/;
assign _5309_ = D[47] ^ Q[51] /*39316*/;
assign _5306_ = _4666_ & _5309_ /*39312*/;
assign _5307_ = _4666_ ^ _5309_ /*39315*/;
assign _5308_ = _5300_ & _5307_ /*39313*/;
assign _5305_ = _5306_ | _5308_ /*39311*/;
assign _5052_ = _5300_ ^ _5307_ /*39314*/;
assign _5314_ = D[48] ^ Q[51] /*39310*/;
assign _5311_ = _4667_ & _5314_ /*39306*/;
assign _5312_ = _4667_ ^ _5314_ /*39309*/;
assign _5313_ = _5305_ & _5312_ /*39307*/;
assign _5310_ = _5311_ | _5313_ /*39305*/;
assign _5053_ = _5305_ ^ _5312_ /*39308*/;
assign _5319_ = D[49] ^ Q[51] /*39304*/;
assign _5316_ = _4668_ & _5319_ /*39300*/;
assign _5317_ = _4668_ ^ _5319_ /*39303*/;
assign _5318_ = _5310_ & _5317_ /*39301*/;
assign _5315_ = _5316_ | _5318_ /*39299*/;
assign _5054_ = _5310_ ^ _5317_ /*39302*/;
assign _5324_ = D[50] ^ Q[51] /*39298*/;
assign _5321_ = _4669_ & _5324_ /*39294*/;
assign _5322_ = _4669_ ^ _5324_ /*39297*/;
assign _5323_ = _5315_ & _5322_ /*39295*/;
assign _5320_ = _5321_ | _5323_ /*39293*/;
assign _5055_ = _5315_ ^ _5322_ /*39296*/;
assign _5329_ = D[51] ^ Q[51] /*39292*/;
assign _5326_ = _4670_ & _5329_ /*39288*/;
assign _5327_ = _4670_ ^ _5329_ /*39291*/;
assign _5328_ = _5320_ & _5327_ /*39289*/;
assign _5325_ = _5326_ | _5328_ /*39287*/;
assign _5056_ = _5320_ ^ _5327_ /*39290*/;
assign _5334_ = D[52] ^ Q[51] /*39286*/;
assign _5331_ = _4671_ & _5334_ /*39282*/;
assign _5332_ = _4671_ ^ _5334_ /*39285*/;
assign _5333_ = _5325_ & _5332_ /*39283*/;
assign _5330_ = _5331_ | _5333_ /*39281*/;
assign _5057_ = _5325_ ^ _5332_ /*39284*/;
assign _5339_ = D[53] ^ Q[51] /*39280*/;
assign _5336_ = _4672_ & _5339_ /*39276*/;
assign _5337_ = _4672_ ^ _5339_ /*39279*/;
assign _5338_ = _5330_ & _5337_ /*39277*/;
assign _5335_ = _5336_ | _5338_ /*39275*/;
assign _5058_ = _5330_ ^ _5337_ /*39278*/;
assign _5344_ = D[54] ^ Q[51] /*39274*/;
assign _5341_ = _4673_ & _5344_ /*39270*/;
assign _5342_ = _4673_ ^ _5344_ /*39273*/;
assign _5343_ = _5335_ & _5342_ /*39271*/;
assign _5340_ = _5341_ | _5343_ /*39269*/;
assign _5059_ = _5335_ ^ _5342_ /*39272*/;
assign _5349_ = D[55] ^ Q[51] /*39268*/;
assign _5346_ = _4674_ & _5349_ /*39264*/;
assign _5347_ = _4674_ ^ _5349_ /*39267*/;
assign _5348_ = _5340_ & _5347_ /*39265*/;
assign _5345_ = _5346_ | _5348_ /*39263*/;
assign _5060_ = _5340_ ^ _5347_ /*39266*/;
assign _5354_ = D[56] ^ Q[51] /*39262*/;
assign _5351_ = _4675_ & _5354_ /*39258*/;
assign _5352_ = _4675_ ^ _5354_ /*39261*/;
assign _5353_ = _5345_ & _5352_ /*39259*/;
assign _5350_ = _5351_ | _5353_ /*39257*/;
assign _5061_ = _5345_ ^ _5352_ /*39260*/;
assign _5359_ = D[57] ^ Q[51] /*39256*/;
assign _5356_ = _4676_ & _5359_ /*39252*/;
assign _5357_ = _4676_ ^ _5359_ /*39255*/;
assign _5358_ = _5350_ & _5357_ /*39253*/;
assign _5355_ = _5356_ | _5358_ /*39251*/;
assign _5062_ = _5350_ ^ _5357_ /*39254*/;
assign _5364_ = D[58] ^ Q[51] /*39250*/;
assign _5361_ = _4677_ & _5364_ /*39246*/;
assign _5362_ = _4677_ ^ _5364_ /*39249*/;
assign _5363_ = _5355_ & _5362_ /*39247*/;
assign _5360_ = _5361_ | _5363_ /*39245*/;
assign _5063_ = _5355_ ^ _5362_ /*39248*/;
assign _5369_ = D[59] ^ Q[51] /*39244*/;
assign _5366_ = _4678_ & _5369_ /*39240*/;
assign _5367_ = _4678_ ^ _5369_ /*39243*/;
assign _5368_ = _5360_ & _5367_ /*39241*/;
assign _5365_ = _5366_ | _5368_ /*39239*/;
assign _5064_ = _5360_ ^ _5367_ /*39242*/;
assign _5374_ = D[60] ^ Q[51] /*39238*/;
assign _5371_ = _4679_ & _5374_ /*39234*/;
assign _5372_ = _4679_ ^ _5374_ /*39237*/;
assign _5373_ = _5365_ & _5372_ /*39235*/;
assign _5370_ = _5371_ | _5373_ /*39233*/;
assign _5065_ = _5365_ ^ _5372_ /*39236*/;
assign _5379_ = D[61] ^ Q[51] /*39232*/;
assign _5376_ = _4680_ & _5379_ /*39228*/;
assign _5377_ = _4680_ ^ _5379_ /*39231*/;
assign _5378_ = _5370_ & _5377_ /*39229*/;
assign _5375_ = _5376_ | _5378_ /*39227*/;
assign _5066_ = _5370_ ^ _5377_ /*39230*/;
assign _5384_ = D[62] ^ Q[51] /*39226*/;
assign _5381_ = _4681_ & _5384_ /*39222*/;
assign _5382_ = _4681_ ^ _5384_ /*39225*/;
assign _5383_ = _5375_ & _5382_ /*39223*/;
assign _5380_ = _5381_ | _5383_ /*39221*/;
assign _5067_ = _5375_ ^ _5382_ /*39224*/;
assign _5388_ = zeroWire ^ Q[51] /*39220*/;
assign _5385_ = _4682_ & _5388_ /*39216*/;
assign _5386_ = _4682_ ^ _5388_ /*39219*/;
assign _5387_ = _5380_ & _5386_ /*39217*/;
assign Q[50] = _5385_ | _5387_ /*39215*/;
assign _5068_ = _5380_ ^ _5386_ /*39218*/;
assign _5459_ = D[0] ^ Q[50] /*38829*/;
assign _5456_ = R_0[49] & _5459_ /*38825*/;
assign _5457_ = R_0[49] ^ _5459_ /*38828*/;
assign _5458_ = Q[50] & _5457_ /*38826*/;
assign _5455_ = _5456_ | _5458_ /*38824*/;
assign _5390_ = Q[50] ^ _5457_ /*38827*/;
assign _5464_ = D[1] ^ Q[50] /*38823*/;
assign _5461_ = _5005_ & _5464_ /*38819*/;
assign _5462_ = _5005_ ^ _5464_ /*38822*/;
assign _5463_ = _5455_ & _5462_ /*38820*/;
assign _5460_ = _5461_ | _5463_ /*38818*/;
assign _5391_ = _5455_ ^ _5462_ /*38821*/;
assign _5469_ = D[2] ^ Q[50] /*38817*/;
assign _5466_ = _5006_ & _5469_ /*38813*/;
assign _5467_ = _5006_ ^ _5469_ /*38816*/;
assign _5468_ = _5460_ & _5467_ /*38814*/;
assign _5465_ = _5466_ | _5468_ /*38812*/;
assign _5392_ = _5460_ ^ _5467_ /*38815*/;
assign _5474_ = D[3] ^ Q[50] /*38811*/;
assign _5471_ = _5007_ & _5474_ /*38807*/;
assign _5472_ = _5007_ ^ _5474_ /*38810*/;
assign _5473_ = _5465_ & _5472_ /*38808*/;
assign _5470_ = _5471_ | _5473_ /*38806*/;
assign _5393_ = _5465_ ^ _5472_ /*38809*/;
assign _5479_ = D[4] ^ Q[50] /*38805*/;
assign _5476_ = _5008_ & _5479_ /*38801*/;
assign _5477_ = _5008_ ^ _5479_ /*38804*/;
assign _5478_ = _5470_ & _5477_ /*38802*/;
assign _5475_ = _5476_ | _5478_ /*38800*/;
assign _5394_ = _5470_ ^ _5477_ /*38803*/;
assign _5484_ = D[5] ^ Q[50] /*38799*/;
assign _5481_ = _5009_ & _5484_ /*38795*/;
assign _5482_ = _5009_ ^ _5484_ /*38798*/;
assign _5483_ = _5475_ & _5482_ /*38796*/;
assign _5480_ = _5481_ | _5483_ /*38794*/;
assign _5395_ = _5475_ ^ _5482_ /*38797*/;
assign _5489_ = D[6] ^ Q[50] /*38793*/;
assign _5486_ = _5010_ & _5489_ /*38789*/;
assign _5487_ = _5010_ ^ _5489_ /*38792*/;
assign _5488_ = _5480_ & _5487_ /*38790*/;
assign _5485_ = _5486_ | _5488_ /*38788*/;
assign _5396_ = _5480_ ^ _5487_ /*38791*/;
assign _5494_ = D[7] ^ Q[50] /*38787*/;
assign _5491_ = _5011_ & _5494_ /*38783*/;
assign _5492_ = _5011_ ^ _5494_ /*38786*/;
assign _5493_ = _5485_ & _5492_ /*38784*/;
assign _5490_ = _5491_ | _5493_ /*38782*/;
assign _5397_ = _5485_ ^ _5492_ /*38785*/;
assign _5499_ = D[8] ^ Q[50] /*38781*/;
assign _5496_ = _5012_ & _5499_ /*38777*/;
assign _5497_ = _5012_ ^ _5499_ /*38780*/;
assign _5498_ = _5490_ & _5497_ /*38778*/;
assign _5495_ = _5496_ | _5498_ /*38776*/;
assign _5398_ = _5490_ ^ _5497_ /*38779*/;
assign _5504_ = D[9] ^ Q[50] /*38775*/;
assign _5501_ = _5013_ & _5504_ /*38771*/;
assign _5502_ = _5013_ ^ _5504_ /*38774*/;
assign _5503_ = _5495_ & _5502_ /*38772*/;
assign _5500_ = _5501_ | _5503_ /*38770*/;
assign _5399_ = _5495_ ^ _5502_ /*38773*/;
assign _5509_ = D[10] ^ Q[50] /*38769*/;
assign _5506_ = _5014_ & _5509_ /*38765*/;
assign _5507_ = _5014_ ^ _5509_ /*38768*/;
assign _5508_ = _5500_ & _5507_ /*38766*/;
assign _5505_ = _5506_ | _5508_ /*38764*/;
assign _5400_ = _5500_ ^ _5507_ /*38767*/;
assign _5514_ = D[11] ^ Q[50] /*38763*/;
assign _5511_ = _5015_ & _5514_ /*38759*/;
assign _5512_ = _5015_ ^ _5514_ /*38762*/;
assign _5513_ = _5505_ & _5512_ /*38760*/;
assign _5510_ = _5511_ | _5513_ /*38758*/;
assign _5401_ = _5505_ ^ _5512_ /*38761*/;
assign _5519_ = D[12] ^ Q[50] /*38757*/;
assign _5516_ = _5016_ & _5519_ /*38753*/;
assign _5517_ = _5016_ ^ _5519_ /*38756*/;
assign _5518_ = _5510_ & _5517_ /*38754*/;
assign _5515_ = _5516_ | _5518_ /*38752*/;
assign _5402_ = _5510_ ^ _5517_ /*38755*/;
assign _5524_ = D[13] ^ Q[50] /*38751*/;
assign _5521_ = _5017_ & _5524_ /*38747*/;
assign _5522_ = _5017_ ^ _5524_ /*38750*/;
assign _5523_ = _5515_ & _5522_ /*38748*/;
assign _5520_ = _5521_ | _5523_ /*38746*/;
assign _5403_ = _5515_ ^ _5522_ /*38749*/;
assign _5529_ = D[14] ^ Q[50] /*38745*/;
assign _5526_ = _5018_ & _5529_ /*38741*/;
assign _5527_ = _5018_ ^ _5529_ /*38744*/;
assign _5528_ = _5520_ & _5527_ /*38742*/;
assign _5525_ = _5526_ | _5528_ /*38740*/;
assign _5404_ = _5520_ ^ _5527_ /*38743*/;
assign _5534_ = D[15] ^ Q[50] /*38739*/;
assign _5531_ = _5019_ & _5534_ /*38735*/;
assign _5532_ = _5019_ ^ _5534_ /*38738*/;
assign _5533_ = _5525_ & _5532_ /*38736*/;
assign _5530_ = _5531_ | _5533_ /*38734*/;
assign _5405_ = _5525_ ^ _5532_ /*38737*/;
assign _5539_ = D[16] ^ Q[50] /*38733*/;
assign _5536_ = _5020_ & _5539_ /*38729*/;
assign _5537_ = _5020_ ^ _5539_ /*38732*/;
assign _5538_ = _5530_ & _5537_ /*38730*/;
assign _5535_ = _5536_ | _5538_ /*38728*/;
assign _5406_ = _5530_ ^ _5537_ /*38731*/;
assign _5544_ = D[17] ^ Q[50] /*38727*/;
assign _5541_ = _5021_ & _5544_ /*38723*/;
assign _5542_ = _5021_ ^ _5544_ /*38726*/;
assign _5543_ = _5535_ & _5542_ /*38724*/;
assign _5540_ = _5541_ | _5543_ /*38722*/;
assign _5407_ = _5535_ ^ _5542_ /*38725*/;
assign _5549_ = D[18] ^ Q[50] /*38721*/;
assign _5546_ = _5022_ & _5549_ /*38717*/;
assign _5547_ = _5022_ ^ _5549_ /*38720*/;
assign _5548_ = _5540_ & _5547_ /*38718*/;
assign _5545_ = _5546_ | _5548_ /*38716*/;
assign _5408_ = _5540_ ^ _5547_ /*38719*/;
assign _5554_ = D[19] ^ Q[50] /*38715*/;
assign _5551_ = _5023_ & _5554_ /*38711*/;
assign _5552_ = _5023_ ^ _5554_ /*38714*/;
assign _5553_ = _5545_ & _5552_ /*38712*/;
assign _5550_ = _5551_ | _5553_ /*38710*/;
assign _5409_ = _5545_ ^ _5552_ /*38713*/;
assign _5559_ = D[20] ^ Q[50] /*38709*/;
assign _5556_ = _5024_ & _5559_ /*38705*/;
assign _5557_ = _5024_ ^ _5559_ /*38708*/;
assign _5558_ = _5550_ & _5557_ /*38706*/;
assign _5555_ = _5556_ | _5558_ /*38704*/;
assign _5410_ = _5550_ ^ _5557_ /*38707*/;
assign _5564_ = D[21] ^ Q[50] /*38703*/;
assign _5561_ = _5025_ & _5564_ /*38699*/;
assign _5562_ = _5025_ ^ _5564_ /*38702*/;
assign _5563_ = _5555_ & _5562_ /*38700*/;
assign _5560_ = _5561_ | _5563_ /*38698*/;
assign _5411_ = _5555_ ^ _5562_ /*38701*/;
assign _5569_ = D[22] ^ Q[50] /*38697*/;
assign _5566_ = _5026_ & _5569_ /*38693*/;
assign _5567_ = _5026_ ^ _5569_ /*38696*/;
assign _5568_ = _5560_ & _5567_ /*38694*/;
assign _5565_ = _5566_ | _5568_ /*38692*/;
assign _5412_ = _5560_ ^ _5567_ /*38695*/;
assign _5574_ = D[23] ^ Q[50] /*38691*/;
assign _5571_ = _5027_ & _5574_ /*38687*/;
assign _5572_ = _5027_ ^ _5574_ /*38690*/;
assign _5573_ = _5565_ & _5572_ /*38688*/;
assign _5570_ = _5571_ | _5573_ /*38686*/;
assign _5413_ = _5565_ ^ _5572_ /*38689*/;
assign _5579_ = D[24] ^ Q[50] /*38685*/;
assign _5576_ = _5028_ & _5579_ /*38681*/;
assign _5577_ = _5028_ ^ _5579_ /*38684*/;
assign _5578_ = _5570_ & _5577_ /*38682*/;
assign _5575_ = _5576_ | _5578_ /*38680*/;
assign _5414_ = _5570_ ^ _5577_ /*38683*/;
assign _5584_ = D[25] ^ Q[50] /*38679*/;
assign _5581_ = _5029_ & _5584_ /*38675*/;
assign _5582_ = _5029_ ^ _5584_ /*38678*/;
assign _5583_ = _5575_ & _5582_ /*38676*/;
assign _5580_ = _5581_ | _5583_ /*38674*/;
assign _5415_ = _5575_ ^ _5582_ /*38677*/;
assign _5589_ = D[26] ^ Q[50] /*38673*/;
assign _5586_ = _5030_ & _5589_ /*38669*/;
assign _5587_ = _5030_ ^ _5589_ /*38672*/;
assign _5588_ = _5580_ & _5587_ /*38670*/;
assign _5585_ = _5586_ | _5588_ /*38668*/;
assign _5416_ = _5580_ ^ _5587_ /*38671*/;
assign _5594_ = D[27] ^ Q[50] /*38667*/;
assign _5591_ = _5031_ & _5594_ /*38663*/;
assign _5592_ = _5031_ ^ _5594_ /*38666*/;
assign _5593_ = _5585_ & _5592_ /*38664*/;
assign _5590_ = _5591_ | _5593_ /*38662*/;
assign _5417_ = _5585_ ^ _5592_ /*38665*/;
assign _5599_ = D[28] ^ Q[50] /*38661*/;
assign _5596_ = _5032_ & _5599_ /*38657*/;
assign _5597_ = _5032_ ^ _5599_ /*38660*/;
assign _5598_ = _5590_ & _5597_ /*38658*/;
assign _5595_ = _5596_ | _5598_ /*38656*/;
assign _5418_ = _5590_ ^ _5597_ /*38659*/;
assign _5604_ = D[29] ^ Q[50] /*38655*/;
assign _5601_ = _5033_ & _5604_ /*38651*/;
assign _5602_ = _5033_ ^ _5604_ /*38654*/;
assign _5603_ = _5595_ & _5602_ /*38652*/;
assign _5600_ = _5601_ | _5603_ /*38650*/;
assign _5419_ = _5595_ ^ _5602_ /*38653*/;
assign _5609_ = D[30] ^ Q[50] /*38649*/;
assign _5606_ = _5034_ & _5609_ /*38645*/;
assign _5607_ = _5034_ ^ _5609_ /*38648*/;
assign _5608_ = _5600_ & _5607_ /*38646*/;
assign _5605_ = _5606_ | _5608_ /*38644*/;
assign _5420_ = _5600_ ^ _5607_ /*38647*/;
assign _5614_ = D[31] ^ Q[50] /*38643*/;
assign _5611_ = _5035_ & _5614_ /*38639*/;
assign _5612_ = _5035_ ^ _5614_ /*38642*/;
assign _5613_ = _5605_ & _5612_ /*38640*/;
assign _5610_ = _5611_ | _5613_ /*38638*/;
assign _5421_ = _5605_ ^ _5612_ /*38641*/;
assign _5619_ = D[32] ^ Q[50] /*38637*/;
assign _5616_ = _5036_ & _5619_ /*38633*/;
assign _5617_ = _5036_ ^ _5619_ /*38636*/;
assign _5618_ = _5610_ & _5617_ /*38634*/;
assign _5615_ = _5616_ | _5618_ /*38632*/;
assign _5422_ = _5610_ ^ _5617_ /*38635*/;
assign _5624_ = D[33] ^ Q[50] /*38631*/;
assign _5621_ = _5037_ & _5624_ /*38627*/;
assign _5622_ = _5037_ ^ _5624_ /*38630*/;
assign _5623_ = _5615_ & _5622_ /*38628*/;
assign _5620_ = _5621_ | _5623_ /*38626*/;
assign _5423_ = _5615_ ^ _5622_ /*38629*/;
assign _5629_ = D[34] ^ Q[50] /*38625*/;
assign _5626_ = _5038_ & _5629_ /*38621*/;
assign _5627_ = _5038_ ^ _5629_ /*38624*/;
assign _5628_ = _5620_ & _5627_ /*38622*/;
assign _5625_ = _5626_ | _5628_ /*38620*/;
assign _5424_ = _5620_ ^ _5627_ /*38623*/;
assign _5634_ = D[35] ^ Q[50] /*38619*/;
assign _5631_ = _5039_ & _5634_ /*38615*/;
assign _5632_ = _5039_ ^ _5634_ /*38618*/;
assign _5633_ = _5625_ & _5632_ /*38616*/;
assign _5630_ = _5631_ | _5633_ /*38614*/;
assign _5425_ = _5625_ ^ _5632_ /*38617*/;
assign _5639_ = D[36] ^ Q[50] /*38613*/;
assign _5636_ = _5040_ & _5639_ /*38609*/;
assign _5637_ = _5040_ ^ _5639_ /*38612*/;
assign _5638_ = _5630_ & _5637_ /*38610*/;
assign _5635_ = _5636_ | _5638_ /*38608*/;
assign _5426_ = _5630_ ^ _5637_ /*38611*/;
assign _5644_ = D[37] ^ Q[50] /*38607*/;
assign _5641_ = _5041_ & _5644_ /*38603*/;
assign _5642_ = _5041_ ^ _5644_ /*38606*/;
assign _5643_ = _5635_ & _5642_ /*38604*/;
assign _5640_ = _5641_ | _5643_ /*38602*/;
assign _5427_ = _5635_ ^ _5642_ /*38605*/;
assign _5649_ = D[38] ^ Q[50] /*38601*/;
assign _5646_ = _5042_ & _5649_ /*38597*/;
assign _5647_ = _5042_ ^ _5649_ /*38600*/;
assign _5648_ = _5640_ & _5647_ /*38598*/;
assign _5645_ = _5646_ | _5648_ /*38596*/;
assign _5428_ = _5640_ ^ _5647_ /*38599*/;
assign _5654_ = D[39] ^ Q[50] /*38595*/;
assign _5651_ = _5043_ & _5654_ /*38591*/;
assign _5652_ = _5043_ ^ _5654_ /*38594*/;
assign _5653_ = _5645_ & _5652_ /*38592*/;
assign _5650_ = _5651_ | _5653_ /*38590*/;
assign _5429_ = _5645_ ^ _5652_ /*38593*/;
assign _5659_ = D[40] ^ Q[50] /*38589*/;
assign _5656_ = _5044_ & _5659_ /*38585*/;
assign _5657_ = _5044_ ^ _5659_ /*38588*/;
assign _5658_ = _5650_ & _5657_ /*38586*/;
assign _5655_ = _5656_ | _5658_ /*38584*/;
assign _5430_ = _5650_ ^ _5657_ /*38587*/;
assign _5664_ = D[41] ^ Q[50] /*38583*/;
assign _5661_ = _5045_ & _5664_ /*38579*/;
assign _5662_ = _5045_ ^ _5664_ /*38582*/;
assign _5663_ = _5655_ & _5662_ /*38580*/;
assign _5660_ = _5661_ | _5663_ /*38578*/;
assign _5431_ = _5655_ ^ _5662_ /*38581*/;
assign _5669_ = D[42] ^ Q[50] /*38577*/;
assign _5666_ = _5046_ & _5669_ /*38573*/;
assign _5667_ = _5046_ ^ _5669_ /*38576*/;
assign _5668_ = _5660_ & _5667_ /*38574*/;
assign _5665_ = _5666_ | _5668_ /*38572*/;
assign _5432_ = _5660_ ^ _5667_ /*38575*/;
assign _5674_ = D[43] ^ Q[50] /*38571*/;
assign _5671_ = _5047_ & _5674_ /*38567*/;
assign _5672_ = _5047_ ^ _5674_ /*38570*/;
assign _5673_ = _5665_ & _5672_ /*38568*/;
assign _5670_ = _5671_ | _5673_ /*38566*/;
assign _5433_ = _5665_ ^ _5672_ /*38569*/;
assign _5679_ = D[44] ^ Q[50] /*38565*/;
assign _5676_ = _5048_ & _5679_ /*38561*/;
assign _5677_ = _5048_ ^ _5679_ /*38564*/;
assign _5678_ = _5670_ & _5677_ /*38562*/;
assign _5675_ = _5676_ | _5678_ /*38560*/;
assign _5434_ = _5670_ ^ _5677_ /*38563*/;
assign _5684_ = D[45] ^ Q[50] /*38559*/;
assign _5681_ = _5049_ & _5684_ /*38555*/;
assign _5682_ = _5049_ ^ _5684_ /*38558*/;
assign _5683_ = _5675_ & _5682_ /*38556*/;
assign _5680_ = _5681_ | _5683_ /*38554*/;
assign _5435_ = _5675_ ^ _5682_ /*38557*/;
assign _5689_ = D[46] ^ Q[50] /*38553*/;
assign _5686_ = _5050_ & _5689_ /*38549*/;
assign _5687_ = _5050_ ^ _5689_ /*38552*/;
assign _5688_ = _5680_ & _5687_ /*38550*/;
assign _5685_ = _5686_ | _5688_ /*38548*/;
assign _5436_ = _5680_ ^ _5687_ /*38551*/;
assign _5694_ = D[47] ^ Q[50] /*38547*/;
assign _5691_ = _5051_ & _5694_ /*38543*/;
assign _5692_ = _5051_ ^ _5694_ /*38546*/;
assign _5693_ = _5685_ & _5692_ /*38544*/;
assign _5690_ = _5691_ | _5693_ /*38542*/;
assign _5437_ = _5685_ ^ _5692_ /*38545*/;
assign _5699_ = D[48] ^ Q[50] /*38541*/;
assign _5696_ = _5052_ & _5699_ /*38537*/;
assign _5697_ = _5052_ ^ _5699_ /*38540*/;
assign _5698_ = _5690_ & _5697_ /*38538*/;
assign _5695_ = _5696_ | _5698_ /*38536*/;
assign _5438_ = _5690_ ^ _5697_ /*38539*/;
assign _5704_ = D[49] ^ Q[50] /*38535*/;
assign _5701_ = _5053_ & _5704_ /*38531*/;
assign _5702_ = _5053_ ^ _5704_ /*38534*/;
assign _5703_ = _5695_ & _5702_ /*38532*/;
assign _5700_ = _5701_ | _5703_ /*38530*/;
assign _5439_ = _5695_ ^ _5702_ /*38533*/;
assign _5709_ = D[50] ^ Q[50] /*38529*/;
assign _5706_ = _5054_ & _5709_ /*38525*/;
assign _5707_ = _5054_ ^ _5709_ /*38528*/;
assign _5708_ = _5700_ & _5707_ /*38526*/;
assign _5705_ = _5706_ | _5708_ /*38524*/;
assign _5440_ = _5700_ ^ _5707_ /*38527*/;
assign _5714_ = D[51] ^ Q[50] /*38523*/;
assign _5711_ = _5055_ & _5714_ /*38519*/;
assign _5712_ = _5055_ ^ _5714_ /*38522*/;
assign _5713_ = _5705_ & _5712_ /*38520*/;
assign _5710_ = _5711_ | _5713_ /*38518*/;
assign _5441_ = _5705_ ^ _5712_ /*38521*/;
assign _5719_ = D[52] ^ Q[50] /*38517*/;
assign _5716_ = _5056_ & _5719_ /*38513*/;
assign _5717_ = _5056_ ^ _5719_ /*38516*/;
assign _5718_ = _5710_ & _5717_ /*38514*/;
assign _5715_ = _5716_ | _5718_ /*38512*/;
assign _5442_ = _5710_ ^ _5717_ /*38515*/;
assign _5724_ = D[53] ^ Q[50] /*38511*/;
assign _5721_ = _5057_ & _5724_ /*38507*/;
assign _5722_ = _5057_ ^ _5724_ /*38510*/;
assign _5723_ = _5715_ & _5722_ /*38508*/;
assign _5720_ = _5721_ | _5723_ /*38506*/;
assign _5443_ = _5715_ ^ _5722_ /*38509*/;
assign _5729_ = D[54] ^ Q[50] /*38505*/;
assign _5726_ = _5058_ & _5729_ /*38501*/;
assign _5727_ = _5058_ ^ _5729_ /*38504*/;
assign _5728_ = _5720_ & _5727_ /*38502*/;
assign _5725_ = _5726_ | _5728_ /*38500*/;
assign _5444_ = _5720_ ^ _5727_ /*38503*/;
assign _5734_ = D[55] ^ Q[50] /*38499*/;
assign _5731_ = _5059_ & _5734_ /*38495*/;
assign _5732_ = _5059_ ^ _5734_ /*38498*/;
assign _5733_ = _5725_ & _5732_ /*38496*/;
assign _5730_ = _5731_ | _5733_ /*38494*/;
assign _5445_ = _5725_ ^ _5732_ /*38497*/;
assign _5739_ = D[56] ^ Q[50] /*38493*/;
assign _5736_ = _5060_ & _5739_ /*38489*/;
assign _5737_ = _5060_ ^ _5739_ /*38492*/;
assign _5738_ = _5730_ & _5737_ /*38490*/;
assign _5735_ = _5736_ | _5738_ /*38488*/;
assign _5446_ = _5730_ ^ _5737_ /*38491*/;
assign _5744_ = D[57] ^ Q[50] /*38487*/;
assign _5741_ = _5061_ & _5744_ /*38483*/;
assign _5742_ = _5061_ ^ _5744_ /*38486*/;
assign _5743_ = _5735_ & _5742_ /*38484*/;
assign _5740_ = _5741_ | _5743_ /*38482*/;
assign _5447_ = _5735_ ^ _5742_ /*38485*/;
assign _5749_ = D[58] ^ Q[50] /*38481*/;
assign _5746_ = _5062_ & _5749_ /*38477*/;
assign _5747_ = _5062_ ^ _5749_ /*38480*/;
assign _5748_ = _5740_ & _5747_ /*38478*/;
assign _5745_ = _5746_ | _5748_ /*38476*/;
assign _5448_ = _5740_ ^ _5747_ /*38479*/;
assign _5754_ = D[59] ^ Q[50] /*38475*/;
assign _5751_ = _5063_ & _5754_ /*38471*/;
assign _5752_ = _5063_ ^ _5754_ /*38474*/;
assign _5753_ = _5745_ & _5752_ /*38472*/;
assign _5750_ = _5751_ | _5753_ /*38470*/;
assign _5449_ = _5745_ ^ _5752_ /*38473*/;
assign _5759_ = D[60] ^ Q[50] /*38469*/;
assign _5756_ = _5064_ & _5759_ /*38465*/;
assign _5757_ = _5064_ ^ _5759_ /*38468*/;
assign _5758_ = _5750_ & _5757_ /*38466*/;
assign _5755_ = _5756_ | _5758_ /*38464*/;
assign _5450_ = _5750_ ^ _5757_ /*38467*/;
assign _5764_ = D[61] ^ Q[50] /*38463*/;
assign _5761_ = _5065_ & _5764_ /*38459*/;
assign _5762_ = _5065_ ^ _5764_ /*38462*/;
assign _5763_ = _5755_ & _5762_ /*38460*/;
assign _5760_ = _5761_ | _5763_ /*38458*/;
assign _5451_ = _5755_ ^ _5762_ /*38461*/;
assign _5769_ = D[62] ^ Q[50] /*38457*/;
assign _5766_ = _5066_ & _5769_ /*38453*/;
assign _5767_ = _5066_ ^ _5769_ /*38456*/;
assign _5768_ = _5760_ & _5767_ /*38454*/;
assign _5765_ = _5766_ | _5768_ /*38452*/;
assign _5452_ = _5760_ ^ _5767_ /*38455*/;
assign _5773_ = zeroWire ^ Q[50] /*38451*/;
assign _5770_ = _5067_ & _5773_ /*38447*/;
assign _5771_ = _5067_ ^ _5773_ /*38450*/;
assign _5772_ = _5765_ & _5771_ /*38448*/;
assign Q[49] = _5770_ | _5772_ /*38446*/;
assign _5453_ = _5765_ ^ _5771_ /*38449*/;
assign _5844_ = D[0] ^ Q[49] /*38060*/;
assign _5841_ = R_0[48] & _5844_ /*38056*/;
assign _5842_ = R_0[48] ^ _5844_ /*38059*/;
assign _5843_ = Q[49] & _5842_ /*38057*/;
assign _5840_ = _5841_ | _5843_ /*38055*/;
assign _5775_ = Q[49] ^ _5842_ /*38058*/;
assign _5849_ = D[1] ^ Q[49] /*38054*/;
assign _5846_ = _5390_ & _5849_ /*38050*/;
assign _5847_ = _5390_ ^ _5849_ /*38053*/;
assign _5848_ = _5840_ & _5847_ /*38051*/;
assign _5845_ = _5846_ | _5848_ /*38049*/;
assign _5776_ = _5840_ ^ _5847_ /*38052*/;
assign _5854_ = D[2] ^ Q[49] /*38048*/;
assign _5851_ = _5391_ & _5854_ /*38044*/;
assign _5852_ = _5391_ ^ _5854_ /*38047*/;
assign _5853_ = _5845_ & _5852_ /*38045*/;
assign _5850_ = _5851_ | _5853_ /*38043*/;
assign _5777_ = _5845_ ^ _5852_ /*38046*/;
assign _5859_ = D[3] ^ Q[49] /*38042*/;
assign _5856_ = _5392_ & _5859_ /*38038*/;
assign _5857_ = _5392_ ^ _5859_ /*38041*/;
assign _5858_ = _5850_ & _5857_ /*38039*/;
assign _5855_ = _5856_ | _5858_ /*38037*/;
assign _5778_ = _5850_ ^ _5857_ /*38040*/;
assign _5864_ = D[4] ^ Q[49] /*38036*/;
assign _5861_ = _5393_ & _5864_ /*38032*/;
assign _5862_ = _5393_ ^ _5864_ /*38035*/;
assign _5863_ = _5855_ & _5862_ /*38033*/;
assign _5860_ = _5861_ | _5863_ /*38031*/;
assign _5779_ = _5855_ ^ _5862_ /*38034*/;
assign _5869_ = D[5] ^ Q[49] /*38030*/;
assign _5866_ = _5394_ & _5869_ /*38026*/;
assign _5867_ = _5394_ ^ _5869_ /*38029*/;
assign _5868_ = _5860_ & _5867_ /*38027*/;
assign _5865_ = _5866_ | _5868_ /*38025*/;
assign _5780_ = _5860_ ^ _5867_ /*38028*/;
assign _5874_ = D[6] ^ Q[49] /*38024*/;
assign _5871_ = _5395_ & _5874_ /*38020*/;
assign _5872_ = _5395_ ^ _5874_ /*38023*/;
assign _5873_ = _5865_ & _5872_ /*38021*/;
assign _5870_ = _5871_ | _5873_ /*38019*/;
assign _5781_ = _5865_ ^ _5872_ /*38022*/;
assign _5879_ = D[7] ^ Q[49] /*38018*/;
assign _5876_ = _5396_ & _5879_ /*38014*/;
assign _5877_ = _5396_ ^ _5879_ /*38017*/;
assign _5878_ = _5870_ & _5877_ /*38015*/;
assign _5875_ = _5876_ | _5878_ /*38013*/;
assign _5782_ = _5870_ ^ _5877_ /*38016*/;
assign _5884_ = D[8] ^ Q[49] /*38012*/;
assign _5881_ = _5397_ & _5884_ /*38008*/;
assign _5882_ = _5397_ ^ _5884_ /*38011*/;
assign _5883_ = _5875_ & _5882_ /*38009*/;
assign _5880_ = _5881_ | _5883_ /*38007*/;
assign _5783_ = _5875_ ^ _5882_ /*38010*/;
assign _5889_ = D[9] ^ Q[49] /*38006*/;
assign _5886_ = _5398_ & _5889_ /*38002*/;
assign _5887_ = _5398_ ^ _5889_ /*38005*/;
assign _5888_ = _5880_ & _5887_ /*38003*/;
assign _5885_ = _5886_ | _5888_ /*38001*/;
assign _5784_ = _5880_ ^ _5887_ /*38004*/;
assign _5894_ = D[10] ^ Q[49] /*38000*/;
assign _5891_ = _5399_ & _5894_ /*37996*/;
assign _5892_ = _5399_ ^ _5894_ /*37999*/;
assign _5893_ = _5885_ & _5892_ /*37997*/;
assign _5890_ = _5891_ | _5893_ /*37995*/;
assign _5785_ = _5885_ ^ _5892_ /*37998*/;
assign _5899_ = D[11] ^ Q[49] /*37994*/;
assign _5896_ = _5400_ & _5899_ /*37990*/;
assign _5897_ = _5400_ ^ _5899_ /*37993*/;
assign _5898_ = _5890_ & _5897_ /*37991*/;
assign _5895_ = _5896_ | _5898_ /*37989*/;
assign _5786_ = _5890_ ^ _5897_ /*37992*/;
assign _5904_ = D[12] ^ Q[49] /*37988*/;
assign _5901_ = _5401_ & _5904_ /*37984*/;
assign _5902_ = _5401_ ^ _5904_ /*37987*/;
assign _5903_ = _5895_ & _5902_ /*37985*/;
assign _5900_ = _5901_ | _5903_ /*37983*/;
assign _5787_ = _5895_ ^ _5902_ /*37986*/;
assign _5909_ = D[13] ^ Q[49] /*37982*/;
assign _5906_ = _5402_ & _5909_ /*37978*/;
assign _5907_ = _5402_ ^ _5909_ /*37981*/;
assign _5908_ = _5900_ & _5907_ /*37979*/;
assign _5905_ = _5906_ | _5908_ /*37977*/;
assign _5788_ = _5900_ ^ _5907_ /*37980*/;
assign _5914_ = D[14] ^ Q[49] /*37976*/;
assign _5911_ = _5403_ & _5914_ /*37972*/;
assign _5912_ = _5403_ ^ _5914_ /*37975*/;
assign _5913_ = _5905_ & _5912_ /*37973*/;
assign _5910_ = _5911_ | _5913_ /*37971*/;
assign _5789_ = _5905_ ^ _5912_ /*37974*/;
assign _5919_ = D[15] ^ Q[49] /*37970*/;
assign _5916_ = _5404_ & _5919_ /*37966*/;
assign _5917_ = _5404_ ^ _5919_ /*37969*/;
assign _5918_ = _5910_ & _5917_ /*37967*/;
assign _5915_ = _5916_ | _5918_ /*37965*/;
assign _5790_ = _5910_ ^ _5917_ /*37968*/;
assign _5924_ = D[16] ^ Q[49] /*37964*/;
assign _5921_ = _5405_ & _5924_ /*37960*/;
assign _5922_ = _5405_ ^ _5924_ /*37963*/;
assign _5923_ = _5915_ & _5922_ /*37961*/;
assign _5920_ = _5921_ | _5923_ /*37959*/;
assign _5791_ = _5915_ ^ _5922_ /*37962*/;
assign _5929_ = D[17] ^ Q[49] /*37958*/;
assign _5926_ = _5406_ & _5929_ /*37954*/;
assign _5927_ = _5406_ ^ _5929_ /*37957*/;
assign _5928_ = _5920_ & _5927_ /*37955*/;
assign _5925_ = _5926_ | _5928_ /*37953*/;
assign _5792_ = _5920_ ^ _5927_ /*37956*/;
assign _5934_ = D[18] ^ Q[49] /*37952*/;
assign _5931_ = _5407_ & _5934_ /*37948*/;
assign _5932_ = _5407_ ^ _5934_ /*37951*/;
assign _5933_ = _5925_ & _5932_ /*37949*/;
assign _5930_ = _5931_ | _5933_ /*37947*/;
assign _5793_ = _5925_ ^ _5932_ /*37950*/;
assign _5939_ = D[19] ^ Q[49] /*37946*/;
assign _5936_ = _5408_ & _5939_ /*37942*/;
assign _5937_ = _5408_ ^ _5939_ /*37945*/;
assign _5938_ = _5930_ & _5937_ /*37943*/;
assign _5935_ = _5936_ | _5938_ /*37941*/;
assign _5794_ = _5930_ ^ _5937_ /*37944*/;
assign _5944_ = D[20] ^ Q[49] /*37940*/;
assign _5941_ = _5409_ & _5944_ /*37936*/;
assign _5942_ = _5409_ ^ _5944_ /*37939*/;
assign _5943_ = _5935_ & _5942_ /*37937*/;
assign _5940_ = _5941_ | _5943_ /*37935*/;
assign _5795_ = _5935_ ^ _5942_ /*37938*/;
assign _5949_ = D[21] ^ Q[49] /*37934*/;
assign _5946_ = _5410_ & _5949_ /*37930*/;
assign _5947_ = _5410_ ^ _5949_ /*37933*/;
assign _5948_ = _5940_ & _5947_ /*37931*/;
assign _5945_ = _5946_ | _5948_ /*37929*/;
assign _5796_ = _5940_ ^ _5947_ /*37932*/;
assign _5954_ = D[22] ^ Q[49] /*37928*/;
assign _5951_ = _5411_ & _5954_ /*37924*/;
assign _5952_ = _5411_ ^ _5954_ /*37927*/;
assign _5953_ = _5945_ & _5952_ /*37925*/;
assign _5950_ = _5951_ | _5953_ /*37923*/;
assign _5797_ = _5945_ ^ _5952_ /*37926*/;
assign _5959_ = D[23] ^ Q[49] /*37922*/;
assign _5956_ = _5412_ & _5959_ /*37918*/;
assign _5957_ = _5412_ ^ _5959_ /*37921*/;
assign _5958_ = _5950_ & _5957_ /*37919*/;
assign _5955_ = _5956_ | _5958_ /*37917*/;
assign _5798_ = _5950_ ^ _5957_ /*37920*/;
assign _5964_ = D[24] ^ Q[49] /*37916*/;
assign _5961_ = _5413_ & _5964_ /*37912*/;
assign _5962_ = _5413_ ^ _5964_ /*37915*/;
assign _5963_ = _5955_ & _5962_ /*37913*/;
assign _5960_ = _5961_ | _5963_ /*37911*/;
assign _5799_ = _5955_ ^ _5962_ /*37914*/;
assign _5969_ = D[25] ^ Q[49] /*37910*/;
assign _5966_ = _5414_ & _5969_ /*37906*/;
assign _5967_ = _5414_ ^ _5969_ /*37909*/;
assign _5968_ = _5960_ & _5967_ /*37907*/;
assign _5965_ = _5966_ | _5968_ /*37905*/;
assign _5800_ = _5960_ ^ _5967_ /*37908*/;
assign _5974_ = D[26] ^ Q[49] /*37904*/;
assign _5971_ = _5415_ & _5974_ /*37900*/;
assign _5972_ = _5415_ ^ _5974_ /*37903*/;
assign _5973_ = _5965_ & _5972_ /*37901*/;
assign _5970_ = _5971_ | _5973_ /*37899*/;
assign _5801_ = _5965_ ^ _5972_ /*37902*/;
assign _5979_ = D[27] ^ Q[49] /*37898*/;
assign _5976_ = _5416_ & _5979_ /*37894*/;
assign _5977_ = _5416_ ^ _5979_ /*37897*/;
assign _5978_ = _5970_ & _5977_ /*37895*/;
assign _5975_ = _5976_ | _5978_ /*37893*/;
assign _5802_ = _5970_ ^ _5977_ /*37896*/;
assign _5984_ = D[28] ^ Q[49] /*37892*/;
assign _5981_ = _5417_ & _5984_ /*37888*/;
assign _5982_ = _5417_ ^ _5984_ /*37891*/;
assign _5983_ = _5975_ & _5982_ /*37889*/;
assign _5980_ = _5981_ | _5983_ /*37887*/;
assign _5803_ = _5975_ ^ _5982_ /*37890*/;
assign _5989_ = D[29] ^ Q[49] /*37886*/;
assign _5986_ = _5418_ & _5989_ /*37882*/;
assign _5987_ = _5418_ ^ _5989_ /*37885*/;
assign _5988_ = _5980_ & _5987_ /*37883*/;
assign _5985_ = _5986_ | _5988_ /*37881*/;
assign _5804_ = _5980_ ^ _5987_ /*37884*/;
assign _5994_ = D[30] ^ Q[49] /*37880*/;
assign _5991_ = _5419_ & _5994_ /*37876*/;
assign _5992_ = _5419_ ^ _5994_ /*37879*/;
assign _5993_ = _5985_ & _5992_ /*37877*/;
assign _5990_ = _5991_ | _5993_ /*37875*/;
assign _5805_ = _5985_ ^ _5992_ /*37878*/;
assign _5999_ = D[31] ^ Q[49] /*37874*/;
assign _5996_ = _5420_ & _5999_ /*37870*/;
assign _5997_ = _5420_ ^ _5999_ /*37873*/;
assign _5998_ = _5990_ & _5997_ /*37871*/;
assign _5995_ = _5996_ | _5998_ /*37869*/;
assign _5806_ = _5990_ ^ _5997_ /*37872*/;
assign _6004_ = D[32] ^ Q[49] /*37868*/;
assign _6001_ = _5421_ & _6004_ /*37864*/;
assign _6002_ = _5421_ ^ _6004_ /*37867*/;
assign _6003_ = _5995_ & _6002_ /*37865*/;
assign _6000_ = _6001_ | _6003_ /*37863*/;
assign _5807_ = _5995_ ^ _6002_ /*37866*/;
assign _6009_ = D[33] ^ Q[49] /*37862*/;
assign _6006_ = _5422_ & _6009_ /*37858*/;
assign _6007_ = _5422_ ^ _6009_ /*37861*/;
assign _6008_ = _6000_ & _6007_ /*37859*/;
assign _6005_ = _6006_ | _6008_ /*37857*/;
assign _5808_ = _6000_ ^ _6007_ /*37860*/;
assign _6014_ = D[34] ^ Q[49] /*37856*/;
assign _6011_ = _5423_ & _6014_ /*37852*/;
assign _6012_ = _5423_ ^ _6014_ /*37855*/;
assign _6013_ = _6005_ & _6012_ /*37853*/;
assign _6010_ = _6011_ | _6013_ /*37851*/;
assign _5809_ = _6005_ ^ _6012_ /*37854*/;
assign _6019_ = D[35] ^ Q[49] /*37850*/;
assign _6016_ = _5424_ & _6019_ /*37846*/;
assign _6017_ = _5424_ ^ _6019_ /*37849*/;
assign _6018_ = _6010_ & _6017_ /*37847*/;
assign _6015_ = _6016_ | _6018_ /*37845*/;
assign _5810_ = _6010_ ^ _6017_ /*37848*/;
assign _6024_ = D[36] ^ Q[49] /*37844*/;
assign _6021_ = _5425_ & _6024_ /*37840*/;
assign _6022_ = _5425_ ^ _6024_ /*37843*/;
assign _6023_ = _6015_ & _6022_ /*37841*/;
assign _6020_ = _6021_ | _6023_ /*37839*/;
assign _5811_ = _6015_ ^ _6022_ /*37842*/;
assign _6029_ = D[37] ^ Q[49] /*37838*/;
assign _6026_ = _5426_ & _6029_ /*37834*/;
assign _6027_ = _5426_ ^ _6029_ /*37837*/;
assign _6028_ = _6020_ & _6027_ /*37835*/;
assign _6025_ = _6026_ | _6028_ /*37833*/;
assign _5812_ = _6020_ ^ _6027_ /*37836*/;
assign _6034_ = D[38] ^ Q[49] /*37832*/;
assign _6031_ = _5427_ & _6034_ /*37828*/;
assign _6032_ = _5427_ ^ _6034_ /*37831*/;
assign _6033_ = _6025_ & _6032_ /*37829*/;
assign _6030_ = _6031_ | _6033_ /*37827*/;
assign _5813_ = _6025_ ^ _6032_ /*37830*/;
assign _6039_ = D[39] ^ Q[49] /*37826*/;
assign _6036_ = _5428_ & _6039_ /*37822*/;
assign _6037_ = _5428_ ^ _6039_ /*37825*/;
assign _6038_ = _6030_ & _6037_ /*37823*/;
assign _6035_ = _6036_ | _6038_ /*37821*/;
assign _5814_ = _6030_ ^ _6037_ /*37824*/;
assign _6044_ = D[40] ^ Q[49] /*37820*/;
assign _6041_ = _5429_ & _6044_ /*37816*/;
assign _6042_ = _5429_ ^ _6044_ /*37819*/;
assign _6043_ = _6035_ & _6042_ /*37817*/;
assign _6040_ = _6041_ | _6043_ /*37815*/;
assign _5815_ = _6035_ ^ _6042_ /*37818*/;
assign _6049_ = D[41] ^ Q[49] /*37814*/;
assign _6046_ = _5430_ & _6049_ /*37810*/;
assign _6047_ = _5430_ ^ _6049_ /*37813*/;
assign _6048_ = _6040_ & _6047_ /*37811*/;
assign _6045_ = _6046_ | _6048_ /*37809*/;
assign _5816_ = _6040_ ^ _6047_ /*37812*/;
assign _6054_ = D[42] ^ Q[49] /*37808*/;
assign _6051_ = _5431_ & _6054_ /*37804*/;
assign _6052_ = _5431_ ^ _6054_ /*37807*/;
assign _6053_ = _6045_ & _6052_ /*37805*/;
assign _6050_ = _6051_ | _6053_ /*37803*/;
assign _5817_ = _6045_ ^ _6052_ /*37806*/;
assign _6059_ = D[43] ^ Q[49] /*37802*/;
assign _6056_ = _5432_ & _6059_ /*37798*/;
assign _6057_ = _5432_ ^ _6059_ /*37801*/;
assign _6058_ = _6050_ & _6057_ /*37799*/;
assign _6055_ = _6056_ | _6058_ /*37797*/;
assign _5818_ = _6050_ ^ _6057_ /*37800*/;
assign _6064_ = D[44] ^ Q[49] /*37796*/;
assign _6061_ = _5433_ & _6064_ /*37792*/;
assign _6062_ = _5433_ ^ _6064_ /*37795*/;
assign _6063_ = _6055_ & _6062_ /*37793*/;
assign _6060_ = _6061_ | _6063_ /*37791*/;
assign _5819_ = _6055_ ^ _6062_ /*37794*/;
assign _6069_ = D[45] ^ Q[49] /*37790*/;
assign _6066_ = _5434_ & _6069_ /*37786*/;
assign _6067_ = _5434_ ^ _6069_ /*37789*/;
assign _6068_ = _6060_ & _6067_ /*37787*/;
assign _6065_ = _6066_ | _6068_ /*37785*/;
assign _5820_ = _6060_ ^ _6067_ /*37788*/;
assign _6074_ = D[46] ^ Q[49] /*37784*/;
assign _6071_ = _5435_ & _6074_ /*37780*/;
assign _6072_ = _5435_ ^ _6074_ /*37783*/;
assign _6073_ = _6065_ & _6072_ /*37781*/;
assign _6070_ = _6071_ | _6073_ /*37779*/;
assign _5821_ = _6065_ ^ _6072_ /*37782*/;
assign _6079_ = D[47] ^ Q[49] /*37778*/;
assign _6076_ = _5436_ & _6079_ /*37774*/;
assign _6077_ = _5436_ ^ _6079_ /*37777*/;
assign _6078_ = _6070_ & _6077_ /*37775*/;
assign _6075_ = _6076_ | _6078_ /*37773*/;
assign _5822_ = _6070_ ^ _6077_ /*37776*/;
assign _6084_ = D[48] ^ Q[49] /*37772*/;
assign _6081_ = _5437_ & _6084_ /*37768*/;
assign _6082_ = _5437_ ^ _6084_ /*37771*/;
assign _6083_ = _6075_ & _6082_ /*37769*/;
assign _6080_ = _6081_ | _6083_ /*37767*/;
assign _5823_ = _6075_ ^ _6082_ /*37770*/;
assign _6089_ = D[49] ^ Q[49] /*37766*/;
assign _6086_ = _5438_ & _6089_ /*37762*/;
assign _6087_ = _5438_ ^ _6089_ /*37765*/;
assign _6088_ = _6080_ & _6087_ /*37763*/;
assign _6085_ = _6086_ | _6088_ /*37761*/;
assign _5824_ = _6080_ ^ _6087_ /*37764*/;
assign _6094_ = D[50] ^ Q[49] /*37760*/;
assign _6091_ = _5439_ & _6094_ /*37756*/;
assign _6092_ = _5439_ ^ _6094_ /*37759*/;
assign _6093_ = _6085_ & _6092_ /*37757*/;
assign _6090_ = _6091_ | _6093_ /*37755*/;
assign _5825_ = _6085_ ^ _6092_ /*37758*/;
assign _6099_ = D[51] ^ Q[49] /*37754*/;
assign _6096_ = _5440_ & _6099_ /*37750*/;
assign _6097_ = _5440_ ^ _6099_ /*37753*/;
assign _6098_ = _6090_ & _6097_ /*37751*/;
assign _6095_ = _6096_ | _6098_ /*37749*/;
assign _5826_ = _6090_ ^ _6097_ /*37752*/;
assign _6104_ = D[52] ^ Q[49] /*37748*/;
assign _6101_ = _5441_ & _6104_ /*37744*/;
assign _6102_ = _5441_ ^ _6104_ /*37747*/;
assign _6103_ = _6095_ & _6102_ /*37745*/;
assign _6100_ = _6101_ | _6103_ /*37743*/;
assign _5827_ = _6095_ ^ _6102_ /*37746*/;
assign _6109_ = D[53] ^ Q[49] /*37742*/;
assign _6106_ = _5442_ & _6109_ /*37738*/;
assign _6107_ = _5442_ ^ _6109_ /*37741*/;
assign _6108_ = _6100_ & _6107_ /*37739*/;
assign _6105_ = _6106_ | _6108_ /*37737*/;
assign _5828_ = _6100_ ^ _6107_ /*37740*/;
assign _6114_ = D[54] ^ Q[49] /*37736*/;
assign _6111_ = _5443_ & _6114_ /*37732*/;
assign _6112_ = _5443_ ^ _6114_ /*37735*/;
assign _6113_ = _6105_ & _6112_ /*37733*/;
assign _6110_ = _6111_ | _6113_ /*37731*/;
assign _5829_ = _6105_ ^ _6112_ /*37734*/;
assign _6119_ = D[55] ^ Q[49] /*37730*/;
assign _6116_ = _5444_ & _6119_ /*37726*/;
assign _6117_ = _5444_ ^ _6119_ /*37729*/;
assign _6118_ = _6110_ & _6117_ /*37727*/;
assign _6115_ = _6116_ | _6118_ /*37725*/;
assign _5830_ = _6110_ ^ _6117_ /*37728*/;
assign _6124_ = D[56] ^ Q[49] /*37724*/;
assign _6121_ = _5445_ & _6124_ /*37720*/;
assign _6122_ = _5445_ ^ _6124_ /*37723*/;
assign _6123_ = _6115_ & _6122_ /*37721*/;
assign _6120_ = _6121_ | _6123_ /*37719*/;
assign _5831_ = _6115_ ^ _6122_ /*37722*/;
assign _6129_ = D[57] ^ Q[49] /*37718*/;
assign _6126_ = _5446_ & _6129_ /*37714*/;
assign _6127_ = _5446_ ^ _6129_ /*37717*/;
assign _6128_ = _6120_ & _6127_ /*37715*/;
assign _6125_ = _6126_ | _6128_ /*37713*/;
assign _5832_ = _6120_ ^ _6127_ /*37716*/;
assign _6134_ = D[58] ^ Q[49] /*37712*/;
assign _6131_ = _5447_ & _6134_ /*37708*/;
assign _6132_ = _5447_ ^ _6134_ /*37711*/;
assign _6133_ = _6125_ & _6132_ /*37709*/;
assign _6130_ = _6131_ | _6133_ /*37707*/;
assign _5833_ = _6125_ ^ _6132_ /*37710*/;
assign _6139_ = D[59] ^ Q[49] /*37706*/;
assign _6136_ = _5448_ & _6139_ /*37702*/;
assign _6137_ = _5448_ ^ _6139_ /*37705*/;
assign _6138_ = _6130_ & _6137_ /*37703*/;
assign _6135_ = _6136_ | _6138_ /*37701*/;
assign _5834_ = _6130_ ^ _6137_ /*37704*/;
assign _6144_ = D[60] ^ Q[49] /*37700*/;
assign _6141_ = _5449_ & _6144_ /*37696*/;
assign _6142_ = _5449_ ^ _6144_ /*37699*/;
assign _6143_ = _6135_ & _6142_ /*37697*/;
assign _6140_ = _6141_ | _6143_ /*37695*/;
assign _5835_ = _6135_ ^ _6142_ /*37698*/;
assign _6149_ = D[61] ^ Q[49] /*37694*/;
assign _6146_ = _5450_ & _6149_ /*37690*/;
assign _6147_ = _5450_ ^ _6149_ /*37693*/;
assign _6148_ = _6140_ & _6147_ /*37691*/;
assign _6145_ = _6146_ | _6148_ /*37689*/;
assign _5836_ = _6140_ ^ _6147_ /*37692*/;
assign _6154_ = D[62] ^ Q[49] /*37688*/;
assign _6151_ = _5451_ & _6154_ /*37684*/;
assign _6152_ = _5451_ ^ _6154_ /*37687*/;
assign _6153_ = _6145_ & _6152_ /*37685*/;
assign _6150_ = _6151_ | _6153_ /*37683*/;
assign _5837_ = _6145_ ^ _6152_ /*37686*/;
assign _6158_ = zeroWire ^ Q[49] /*37682*/;
assign _6155_ = _5452_ & _6158_ /*37678*/;
assign _6156_ = _5452_ ^ _6158_ /*37681*/;
assign _6157_ = _6150_ & _6156_ /*37679*/;
assign Q[48] = _6155_ | _6157_ /*37677*/;
assign _5838_ = _6150_ ^ _6156_ /*37680*/;
assign _6229_ = D[0] ^ Q[48] /*37291*/;
assign _6226_ = R_0[47] & _6229_ /*37287*/;
assign _6227_ = R_0[47] ^ _6229_ /*37290*/;
assign _6228_ = Q[48] & _6227_ /*37288*/;
assign _6225_ = _6226_ | _6228_ /*37286*/;
assign _6160_ = Q[48] ^ _6227_ /*37289*/;
assign _6234_ = D[1] ^ Q[48] /*37285*/;
assign _6231_ = _5775_ & _6234_ /*37281*/;
assign _6232_ = _5775_ ^ _6234_ /*37284*/;
assign _6233_ = _6225_ & _6232_ /*37282*/;
assign _6230_ = _6231_ | _6233_ /*37280*/;
assign _6161_ = _6225_ ^ _6232_ /*37283*/;
assign _6239_ = D[2] ^ Q[48] /*37279*/;
assign _6236_ = _5776_ & _6239_ /*37275*/;
assign _6237_ = _5776_ ^ _6239_ /*37278*/;
assign _6238_ = _6230_ & _6237_ /*37276*/;
assign _6235_ = _6236_ | _6238_ /*37274*/;
assign _6162_ = _6230_ ^ _6237_ /*37277*/;
assign _6244_ = D[3] ^ Q[48] /*37273*/;
assign _6241_ = _5777_ & _6244_ /*37269*/;
assign _6242_ = _5777_ ^ _6244_ /*37272*/;
assign _6243_ = _6235_ & _6242_ /*37270*/;
assign _6240_ = _6241_ | _6243_ /*37268*/;
assign _6163_ = _6235_ ^ _6242_ /*37271*/;
assign _6249_ = D[4] ^ Q[48] /*37267*/;
assign _6246_ = _5778_ & _6249_ /*37263*/;
assign _6247_ = _5778_ ^ _6249_ /*37266*/;
assign _6248_ = _6240_ & _6247_ /*37264*/;
assign _6245_ = _6246_ | _6248_ /*37262*/;
assign _6164_ = _6240_ ^ _6247_ /*37265*/;
assign _6254_ = D[5] ^ Q[48] /*37261*/;
assign _6251_ = _5779_ & _6254_ /*37257*/;
assign _6252_ = _5779_ ^ _6254_ /*37260*/;
assign _6253_ = _6245_ & _6252_ /*37258*/;
assign _6250_ = _6251_ | _6253_ /*37256*/;
assign _6165_ = _6245_ ^ _6252_ /*37259*/;
assign _6259_ = D[6] ^ Q[48] /*37255*/;
assign _6256_ = _5780_ & _6259_ /*37251*/;
assign _6257_ = _5780_ ^ _6259_ /*37254*/;
assign _6258_ = _6250_ & _6257_ /*37252*/;
assign _6255_ = _6256_ | _6258_ /*37250*/;
assign _6166_ = _6250_ ^ _6257_ /*37253*/;
assign _6264_ = D[7] ^ Q[48] /*37249*/;
assign _6261_ = _5781_ & _6264_ /*37245*/;
assign _6262_ = _5781_ ^ _6264_ /*37248*/;
assign _6263_ = _6255_ & _6262_ /*37246*/;
assign _6260_ = _6261_ | _6263_ /*37244*/;
assign _6167_ = _6255_ ^ _6262_ /*37247*/;
assign _6269_ = D[8] ^ Q[48] /*37243*/;
assign _6266_ = _5782_ & _6269_ /*37239*/;
assign _6267_ = _5782_ ^ _6269_ /*37242*/;
assign _6268_ = _6260_ & _6267_ /*37240*/;
assign _6265_ = _6266_ | _6268_ /*37238*/;
assign _6168_ = _6260_ ^ _6267_ /*37241*/;
assign _6274_ = D[9] ^ Q[48] /*37237*/;
assign _6271_ = _5783_ & _6274_ /*37233*/;
assign _6272_ = _5783_ ^ _6274_ /*37236*/;
assign _6273_ = _6265_ & _6272_ /*37234*/;
assign _6270_ = _6271_ | _6273_ /*37232*/;
assign _6169_ = _6265_ ^ _6272_ /*37235*/;
assign _6279_ = D[10] ^ Q[48] /*37231*/;
assign _6276_ = _5784_ & _6279_ /*37227*/;
assign _6277_ = _5784_ ^ _6279_ /*37230*/;
assign _6278_ = _6270_ & _6277_ /*37228*/;
assign _6275_ = _6276_ | _6278_ /*37226*/;
assign _6170_ = _6270_ ^ _6277_ /*37229*/;
assign _6284_ = D[11] ^ Q[48] /*37225*/;
assign _6281_ = _5785_ & _6284_ /*37221*/;
assign _6282_ = _5785_ ^ _6284_ /*37224*/;
assign _6283_ = _6275_ & _6282_ /*37222*/;
assign _6280_ = _6281_ | _6283_ /*37220*/;
assign _6171_ = _6275_ ^ _6282_ /*37223*/;
assign _6289_ = D[12] ^ Q[48] /*37219*/;
assign _6286_ = _5786_ & _6289_ /*37215*/;
assign _6287_ = _5786_ ^ _6289_ /*37218*/;
assign _6288_ = _6280_ & _6287_ /*37216*/;
assign _6285_ = _6286_ | _6288_ /*37214*/;
assign _6172_ = _6280_ ^ _6287_ /*37217*/;
assign _6294_ = D[13] ^ Q[48] /*37213*/;
assign _6291_ = _5787_ & _6294_ /*37209*/;
assign _6292_ = _5787_ ^ _6294_ /*37212*/;
assign _6293_ = _6285_ & _6292_ /*37210*/;
assign _6290_ = _6291_ | _6293_ /*37208*/;
assign _6173_ = _6285_ ^ _6292_ /*37211*/;
assign _6299_ = D[14] ^ Q[48] /*37207*/;
assign _6296_ = _5788_ & _6299_ /*37203*/;
assign _6297_ = _5788_ ^ _6299_ /*37206*/;
assign _6298_ = _6290_ & _6297_ /*37204*/;
assign _6295_ = _6296_ | _6298_ /*37202*/;
assign _6174_ = _6290_ ^ _6297_ /*37205*/;
assign _6304_ = D[15] ^ Q[48] /*37201*/;
assign _6301_ = _5789_ & _6304_ /*37197*/;
assign _6302_ = _5789_ ^ _6304_ /*37200*/;
assign _6303_ = _6295_ & _6302_ /*37198*/;
assign _6300_ = _6301_ | _6303_ /*37196*/;
assign _6175_ = _6295_ ^ _6302_ /*37199*/;
assign _6309_ = D[16] ^ Q[48] /*37195*/;
assign _6306_ = _5790_ & _6309_ /*37191*/;
assign _6307_ = _5790_ ^ _6309_ /*37194*/;
assign _6308_ = _6300_ & _6307_ /*37192*/;
assign _6305_ = _6306_ | _6308_ /*37190*/;
assign _6176_ = _6300_ ^ _6307_ /*37193*/;
assign _6314_ = D[17] ^ Q[48] /*37189*/;
assign _6311_ = _5791_ & _6314_ /*37185*/;
assign _6312_ = _5791_ ^ _6314_ /*37188*/;
assign _6313_ = _6305_ & _6312_ /*37186*/;
assign _6310_ = _6311_ | _6313_ /*37184*/;
assign _6177_ = _6305_ ^ _6312_ /*37187*/;
assign _6319_ = D[18] ^ Q[48] /*37183*/;
assign _6316_ = _5792_ & _6319_ /*37179*/;
assign _6317_ = _5792_ ^ _6319_ /*37182*/;
assign _6318_ = _6310_ & _6317_ /*37180*/;
assign _6315_ = _6316_ | _6318_ /*37178*/;
assign _6178_ = _6310_ ^ _6317_ /*37181*/;
assign _6324_ = D[19] ^ Q[48] /*37177*/;
assign _6321_ = _5793_ & _6324_ /*37173*/;
assign _6322_ = _5793_ ^ _6324_ /*37176*/;
assign _6323_ = _6315_ & _6322_ /*37174*/;
assign _6320_ = _6321_ | _6323_ /*37172*/;
assign _6179_ = _6315_ ^ _6322_ /*37175*/;
assign _6329_ = D[20] ^ Q[48] /*37171*/;
assign _6326_ = _5794_ & _6329_ /*37167*/;
assign _6327_ = _5794_ ^ _6329_ /*37170*/;
assign _6328_ = _6320_ & _6327_ /*37168*/;
assign _6325_ = _6326_ | _6328_ /*37166*/;
assign _6180_ = _6320_ ^ _6327_ /*37169*/;
assign _6334_ = D[21] ^ Q[48] /*37165*/;
assign _6331_ = _5795_ & _6334_ /*37161*/;
assign _6332_ = _5795_ ^ _6334_ /*37164*/;
assign _6333_ = _6325_ & _6332_ /*37162*/;
assign _6330_ = _6331_ | _6333_ /*37160*/;
assign _6181_ = _6325_ ^ _6332_ /*37163*/;
assign _6339_ = D[22] ^ Q[48] /*37159*/;
assign _6336_ = _5796_ & _6339_ /*37155*/;
assign _6337_ = _5796_ ^ _6339_ /*37158*/;
assign _6338_ = _6330_ & _6337_ /*37156*/;
assign _6335_ = _6336_ | _6338_ /*37154*/;
assign _6182_ = _6330_ ^ _6337_ /*37157*/;
assign _6344_ = D[23] ^ Q[48] /*37153*/;
assign _6341_ = _5797_ & _6344_ /*37149*/;
assign _6342_ = _5797_ ^ _6344_ /*37152*/;
assign _6343_ = _6335_ & _6342_ /*37150*/;
assign _6340_ = _6341_ | _6343_ /*37148*/;
assign _6183_ = _6335_ ^ _6342_ /*37151*/;
assign _6349_ = D[24] ^ Q[48] /*37147*/;
assign _6346_ = _5798_ & _6349_ /*37143*/;
assign _6347_ = _5798_ ^ _6349_ /*37146*/;
assign _6348_ = _6340_ & _6347_ /*37144*/;
assign _6345_ = _6346_ | _6348_ /*37142*/;
assign _6184_ = _6340_ ^ _6347_ /*37145*/;
assign _6354_ = D[25] ^ Q[48] /*37141*/;
assign _6351_ = _5799_ & _6354_ /*37137*/;
assign _6352_ = _5799_ ^ _6354_ /*37140*/;
assign _6353_ = _6345_ & _6352_ /*37138*/;
assign _6350_ = _6351_ | _6353_ /*37136*/;
assign _6185_ = _6345_ ^ _6352_ /*37139*/;
assign _6359_ = D[26] ^ Q[48] /*37135*/;
assign _6356_ = _5800_ & _6359_ /*37131*/;
assign _6357_ = _5800_ ^ _6359_ /*37134*/;
assign _6358_ = _6350_ & _6357_ /*37132*/;
assign _6355_ = _6356_ | _6358_ /*37130*/;
assign _6186_ = _6350_ ^ _6357_ /*37133*/;
assign _6364_ = D[27] ^ Q[48] /*37129*/;
assign _6361_ = _5801_ & _6364_ /*37125*/;
assign _6362_ = _5801_ ^ _6364_ /*37128*/;
assign _6363_ = _6355_ & _6362_ /*37126*/;
assign _6360_ = _6361_ | _6363_ /*37124*/;
assign _6187_ = _6355_ ^ _6362_ /*37127*/;
assign _6369_ = D[28] ^ Q[48] /*37123*/;
assign _6366_ = _5802_ & _6369_ /*37119*/;
assign _6367_ = _5802_ ^ _6369_ /*37122*/;
assign _6368_ = _6360_ & _6367_ /*37120*/;
assign _6365_ = _6366_ | _6368_ /*37118*/;
assign _6188_ = _6360_ ^ _6367_ /*37121*/;
assign _6374_ = D[29] ^ Q[48] /*37117*/;
assign _6371_ = _5803_ & _6374_ /*37113*/;
assign _6372_ = _5803_ ^ _6374_ /*37116*/;
assign _6373_ = _6365_ & _6372_ /*37114*/;
assign _6370_ = _6371_ | _6373_ /*37112*/;
assign _6189_ = _6365_ ^ _6372_ /*37115*/;
assign _6379_ = D[30] ^ Q[48] /*37111*/;
assign _6376_ = _5804_ & _6379_ /*37107*/;
assign _6377_ = _5804_ ^ _6379_ /*37110*/;
assign _6378_ = _6370_ & _6377_ /*37108*/;
assign _6375_ = _6376_ | _6378_ /*37106*/;
assign _6190_ = _6370_ ^ _6377_ /*37109*/;
assign _6384_ = D[31] ^ Q[48] /*37105*/;
assign _6381_ = _5805_ & _6384_ /*37101*/;
assign _6382_ = _5805_ ^ _6384_ /*37104*/;
assign _6383_ = _6375_ & _6382_ /*37102*/;
assign _6380_ = _6381_ | _6383_ /*37100*/;
assign _6191_ = _6375_ ^ _6382_ /*37103*/;
assign _6389_ = D[32] ^ Q[48] /*37099*/;
assign _6386_ = _5806_ & _6389_ /*37095*/;
assign _6387_ = _5806_ ^ _6389_ /*37098*/;
assign _6388_ = _6380_ & _6387_ /*37096*/;
assign _6385_ = _6386_ | _6388_ /*37094*/;
assign _6192_ = _6380_ ^ _6387_ /*37097*/;
assign _6394_ = D[33] ^ Q[48] /*37093*/;
assign _6391_ = _5807_ & _6394_ /*37089*/;
assign _6392_ = _5807_ ^ _6394_ /*37092*/;
assign _6393_ = _6385_ & _6392_ /*37090*/;
assign _6390_ = _6391_ | _6393_ /*37088*/;
assign _6193_ = _6385_ ^ _6392_ /*37091*/;
assign _6399_ = D[34] ^ Q[48] /*37087*/;
assign _6396_ = _5808_ & _6399_ /*37083*/;
assign _6397_ = _5808_ ^ _6399_ /*37086*/;
assign _6398_ = _6390_ & _6397_ /*37084*/;
assign _6395_ = _6396_ | _6398_ /*37082*/;
assign _6194_ = _6390_ ^ _6397_ /*37085*/;
assign _6404_ = D[35] ^ Q[48] /*37081*/;
assign _6401_ = _5809_ & _6404_ /*37077*/;
assign _6402_ = _5809_ ^ _6404_ /*37080*/;
assign _6403_ = _6395_ & _6402_ /*37078*/;
assign _6400_ = _6401_ | _6403_ /*37076*/;
assign _6195_ = _6395_ ^ _6402_ /*37079*/;
assign _6409_ = D[36] ^ Q[48] /*37075*/;
assign _6406_ = _5810_ & _6409_ /*37071*/;
assign _6407_ = _5810_ ^ _6409_ /*37074*/;
assign _6408_ = _6400_ & _6407_ /*37072*/;
assign _6405_ = _6406_ | _6408_ /*37070*/;
assign _6196_ = _6400_ ^ _6407_ /*37073*/;
assign _6414_ = D[37] ^ Q[48] /*37069*/;
assign _6411_ = _5811_ & _6414_ /*37065*/;
assign _6412_ = _5811_ ^ _6414_ /*37068*/;
assign _6413_ = _6405_ & _6412_ /*37066*/;
assign _6410_ = _6411_ | _6413_ /*37064*/;
assign _6197_ = _6405_ ^ _6412_ /*37067*/;
assign _6419_ = D[38] ^ Q[48] /*37063*/;
assign _6416_ = _5812_ & _6419_ /*37059*/;
assign _6417_ = _5812_ ^ _6419_ /*37062*/;
assign _6418_ = _6410_ & _6417_ /*37060*/;
assign _6415_ = _6416_ | _6418_ /*37058*/;
assign _6198_ = _6410_ ^ _6417_ /*37061*/;
assign _6424_ = D[39] ^ Q[48] /*37057*/;
assign _6421_ = _5813_ & _6424_ /*37053*/;
assign _6422_ = _5813_ ^ _6424_ /*37056*/;
assign _6423_ = _6415_ & _6422_ /*37054*/;
assign _6420_ = _6421_ | _6423_ /*37052*/;
assign _6199_ = _6415_ ^ _6422_ /*37055*/;
assign _6429_ = D[40] ^ Q[48] /*37051*/;
assign _6426_ = _5814_ & _6429_ /*37047*/;
assign _6427_ = _5814_ ^ _6429_ /*37050*/;
assign _6428_ = _6420_ & _6427_ /*37048*/;
assign _6425_ = _6426_ | _6428_ /*37046*/;
assign _6200_ = _6420_ ^ _6427_ /*37049*/;
assign _6434_ = D[41] ^ Q[48] /*37045*/;
assign _6431_ = _5815_ & _6434_ /*37041*/;
assign _6432_ = _5815_ ^ _6434_ /*37044*/;
assign _6433_ = _6425_ & _6432_ /*37042*/;
assign _6430_ = _6431_ | _6433_ /*37040*/;
assign _6201_ = _6425_ ^ _6432_ /*37043*/;
assign _6439_ = D[42] ^ Q[48] /*37039*/;
assign _6436_ = _5816_ & _6439_ /*37035*/;
assign _6437_ = _5816_ ^ _6439_ /*37038*/;
assign _6438_ = _6430_ & _6437_ /*37036*/;
assign _6435_ = _6436_ | _6438_ /*37034*/;
assign _6202_ = _6430_ ^ _6437_ /*37037*/;
assign _6444_ = D[43] ^ Q[48] /*37033*/;
assign _6441_ = _5817_ & _6444_ /*37029*/;
assign _6442_ = _5817_ ^ _6444_ /*37032*/;
assign _6443_ = _6435_ & _6442_ /*37030*/;
assign _6440_ = _6441_ | _6443_ /*37028*/;
assign _6203_ = _6435_ ^ _6442_ /*37031*/;
assign _6449_ = D[44] ^ Q[48] /*37027*/;
assign _6446_ = _5818_ & _6449_ /*37023*/;
assign _6447_ = _5818_ ^ _6449_ /*37026*/;
assign _6448_ = _6440_ & _6447_ /*37024*/;
assign _6445_ = _6446_ | _6448_ /*37022*/;
assign _6204_ = _6440_ ^ _6447_ /*37025*/;
assign _6454_ = D[45] ^ Q[48] /*37021*/;
assign _6451_ = _5819_ & _6454_ /*37017*/;
assign _6452_ = _5819_ ^ _6454_ /*37020*/;
assign _6453_ = _6445_ & _6452_ /*37018*/;
assign _6450_ = _6451_ | _6453_ /*37016*/;
assign _6205_ = _6445_ ^ _6452_ /*37019*/;
assign _6459_ = D[46] ^ Q[48] /*37015*/;
assign _6456_ = _5820_ & _6459_ /*37011*/;
assign _6457_ = _5820_ ^ _6459_ /*37014*/;
assign _6458_ = _6450_ & _6457_ /*37012*/;
assign _6455_ = _6456_ | _6458_ /*37010*/;
assign _6206_ = _6450_ ^ _6457_ /*37013*/;
assign _6464_ = D[47] ^ Q[48] /*37009*/;
assign _6461_ = _5821_ & _6464_ /*37005*/;
assign _6462_ = _5821_ ^ _6464_ /*37008*/;
assign _6463_ = _6455_ & _6462_ /*37006*/;
assign _6460_ = _6461_ | _6463_ /*37004*/;
assign _6207_ = _6455_ ^ _6462_ /*37007*/;
assign _6469_ = D[48] ^ Q[48] /*37003*/;
assign _6466_ = _5822_ & _6469_ /*36999*/;
assign _6467_ = _5822_ ^ _6469_ /*37002*/;
assign _6468_ = _6460_ & _6467_ /*37000*/;
assign _6465_ = _6466_ | _6468_ /*36998*/;
assign _6208_ = _6460_ ^ _6467_ /*37001*/;
assign _6474_ = D[49] ^ Q[48] /*36997*/;
assign _6471_ = _5823_ & _6474_ /*36993*/;
assign _6472_ = _5823_ ^ _6474_ /*36996*/;
assign _6473_ = _6465_ & _6472_ /*36994*/;
assign _6470_ = _6471_ | _6473_ /*36992*/;
assign _6209_ = _6465_ ^ _6472_ /*36995*/;
assign _6479_ = D[50] ^ Q[48] /*36991*/;
assign _6476_ = _5824_ & _6479_ /*36987*/;
assign _6477_ = _5824_ ^ _6479_ /*36990*/;
assign _6478_ = _6470_ & _6477_ /*36988*/;
assign _6475_ = _6476_ | _6478_ /*36986*/;
assign _6210_ = _6470_ ^ _6477_ /*36989*/;
assign _6484_ = D[51] ^ Q[48] /*36985*/;
assign _6481_ = _5825_ & _6484_ /*36981*/;
assign _6482_ = _5825_ ^ _6484_ /*36984*/;
assign _6483_ = _6475_ & _6482_ /*36982*/;
assign _6480_ = _6481_ | _6483_ /*36980*/;
assign _6211_ = _6475_ ^ _6482_ /*36983*/;
assign _6489_ = D[52] ^ Q[48] /*36979*/;
assign _6486_ = _5826_ & _6489_ /*36975*/;
assign _6487_ = _5826_ ^ _6489_ /*36978*/;
assign _6488_ = _6480_ & _6487_ /*36976*/;
assign _6485_ = _6486_ | _6488_ /*36974*/;
assign _6212_ = _6480_ ^ _6487_ /*36977*/;
assign _6494_ = D[53] ^ Q[48] /*36973*/;
assign _6491_ = _5827_ & _6494_ /*36969*/;
assign _6492_ = _5827_ ^ _6494_ /*36972*/;
assign _6493_ = _6485_ & _6492_ /*36970*/;
assign _6490_ = _6491_ | _6493_ /*36968*/;
assign _6213_ = _6485_ ^ _6492_ /*36971*/;
assign _6499_ = D[54] ^ Q[48] /*36967*/;
assign _6496_ = _5828_ & _6499_ /*36963*/;
assign _6497_ = _5828_ ^ _6499_ /*36966*/;
assign _6498_ = _6490_ & _6497_ /*36964*/;
assign _6495_ = _6496_ | _6498_ /*36962*/;
assign _6214_ = _6490_ ^ _6497_ /*36965*/;
assign _6504_ = D[55] ^ Q[48] /*36961*/;
assign _6501_ = _5829_ & _6504_ /*36957*/;
assign _6502_ = _5829_ ^ _6504_ /*36960*/;
assign _6503_ = _6495_ & _6502_ /*36958*/;
assign _6500_ = _6501_ | _6503_ /*36956*/;
assign _6215_ = _6495_ ^ _6502_ /*36959*/;
assign _6509_ = D[56] ^ Q[48] /*36955*/;
assign _6506_ = _5830_ & _6509_ /*36951*/;
assign _6507_ = _5830_ ^ _6509_ /*36954*/;
assign _6508_ = _6500_ & _6507_ /*36952*/;
assign _6505_ = _6506_ | _6508_ /*36950*/;
assign _6216_ = _6500_ ^ _6507_ /*36953*/;
assign _6514_ = D[57] ^ Q[48] /*36949*/;
assign _6511_ = _5831_ & _6514_ /*36945*/;
assign _6512_ = _5831_ ^ _6514_ /*36948*/;
assign _6513_ = _6505_ & _6512_ /*36946*/;
assign _6510_ = _6511_ | _6513_ /*36944*/;
assign _6217_ = _6505_ ^ _6512_ /*36947*/;
assign _6519_ = D[58] ^ Q[48] /*36943*/;
assign _6516_ = _5832_ & _6519_ /*36939*/;
assign _6517_ = _5832_ ^ _6519_ /*36942*/;
assign _6518_ = _6510_ & _6517_ /*36940*/;
assign _6515_ = _6516_ | _6518_ /*36938*/;
assign _6218_ = _6510_ ^ _6517_ /*36941*/;
assign _6524_ = D[59] ^ Q[48] /*36937*/;
assign _6521_ = _5833_ & _6524_ /*36933*/;
assign _6522_ = _5833_ ^ _6524_ /*36936*/;
assign _6523_ = _6515_ & _6522_ /*36934*/;
assign _6520_ = _6521_ | _6523_ /*36932*/;
assign _6219_ = _6515_ ^ _6522_ /*36935*/;
assign _6529_ = D[60] ^ Q[48] /*36931*/;
assign _6526_ = _5834_ & _6529_ /*36927*/;
assign _6527_ = _5834_ ^ _6529_ /*36930*/;
assign _6528_ = _6520_ & _6527_ /*36928*/;
assign _6525_ = _6526_ | _6528_ /*36926*/;
assign _6220_ = _6520_ ^ _6527_ /*36929*/;
assign _6534_ = D[61] ^ Q[48] /*36925*/;
assign _6531_ = _5835_ & _6534_ /*36921*/;
assign _6532_ = _5835_ ^ _6534_ /*36924*/;
assign _6533_ = _6525_ & _6532_ /*36922*/;
assign _6530_ = _6531_ | _6533_ /*36920*/;
assign _6221_ = _6525_ ^ _6532_ /*36923*/;
assign _6539_ = D[62] ^ Q[48] /*36919*/;
assign _6536_ = _5836_ & _6539_ /*36915*/;
assign _6537_ = _5836_ ^ _6539_ /*36918*/;
assign _6538_ = _6530_ & _6537_ /*36916*/;
assign _6535_ = _6536_ | _6538_ /*36914*/;
assign _6222_ = _6530_ ^ _6537_ /*36917*/;
assign _6543_ = zeroWire ^ Q[48] /*36913*/;
assign _6540_ = _5837_ & _6543_ /*36909*/;
assign _6541_ = _5837_ ^ _6543_ /*36912*/;
assign _6542_ = _6535_ & _6541_ /*36910*/;
assign Q[47] = _6540_ | _6542_ /*36908*/;
assign _6223_ = _6535_ ^ _6541_ /*36911*/;
assign _6614_ = D[0] ^ Q[47] /*36522*/;
assign _6611_ = R_0[46] & _6614_ /*36518*/;
assign _6612_ = R_0[46] ^ _6614_ /*36521*/;
assign _6613_ = Q[47] & _6612_ /*36519*/;
assign _6610_ = _6611_ | _6613_ /*36517*/;
assign _6545_ = Q[47] ^ _6612_ /*36520*/;
assign _6619_ = D[1] ^ Q[47] /*36516*/;
assign _6616_ = _6160_ & _6619_ /*36512*/;
assign _6617_ = _6160_ ^ _6619_ /*36515*/;
assign _6618_ = _6610_ & _6617_ /*36513*/;
assign _6615_ = _6616_ | _6618_ /*36511*/;
assign _6546_ = _6610_ ^ _6617_ /*36514*/;
assign _6624_ = D[2] ^ Q[47] /*36510*/;
assign _6621_ = _6161_ & _6624_ /*36506*/;
assign _6622_ = _6161_ ^ _6624_ /*36509*/;
assign _6623_ = _6615_ & _6622_ /*36507*/;
assign _6620_ = _6621_ | _6623_ /*36505*/;
assign _6547_ = _6615_ ^ _6622_ /*36508*/;
assign _6629_ = D[3] ^ Q[47] /*36504*/;
assign _6626_ = _6162_ & _6629_ /*36500*/;
assign _6627_ = _6162_ ^ _6629_ /*36503*/;
assign _6628_ = _6620_ & _6627_ /*36501*/;
assign _6625_ = _6626_ | _6628_ /*36499*/;
assign _6548_ = _6620_ ^ _6627_ /*36502*/;
assign _6634_ = D[4] ^ Q[47] /*36498*/;
assign _6631_ = _6163_ & _6634_ /*36494*/;
assign _6632_ = _6163_ ^ _6634_ /*36497*/;
assign _6633_ = _6625_ & _6632_ /*36495*/;
assign _6630_ = _6631_ | _6633_ /*36493*/;
assign _6549_ = _6625_ ^ _6632_ /*36496*/;
assign _6639_ = D[5] ^ Q[47] /*36492*/;
assign _6636_ = _6164_ & _6639_ /*36488*/;
assign _6637_ = _6164_ ^ _6639_ /*36491*/;
assign _6638_ = _6630_ & _6637_ /*36489*/;
assign _6635_ = _6636_ | _6638_ /*36487*/;
assign _6550_ = _6630_ ^ _6637_ /*36490*/;
assign _6644_ = D[6] ^ Q[47] /*36486*/;
assign _6641_ = _6165_ & _6644_ /*36482*/;
assign _6642_ = _6165_ ^ _6644_ /*36485*/;
assign _6643_ = _6635_ & _6642_ /*36483*/;
assign _6640_ = _6641_ | _6643_ /*36481*/;
assign _6551_ = _6635_ ^ _6642_ /*36484*/;
assign _6649_ = D[7] ^ Q[47] /*36480*/;
assign _6646_ = _6166_ & _6649_ /*36476*/;
assign _6647_ = _6166_ ^ _6649_ /*36479*/;
assign _6648_ = _6640_ & _6647_ /*36477*/;
assign _6645_ = _6646_ | _6648_ /*36475*/;
assign _6552_ = _6640_ ^ _6647_ /*36478*/;
assign _6654_ = D[8] ^ Q[47] /*36474*/;
assign _6651_ = _6167_ & _6654_ /*36470*/;
assign _6652_ = _6167_ ^ _6654_ /*36473*/;
assign _6653_ = _6645_ & _6652_ /*36471*/;
assign _6650_ = _6651_ | _6653_ /*36469*/;
assign _6553_ = _6645_ ^ _6652_ /*36472*/;
assign _6659_ = D[9] ^ Q[47] /*36468*/;
assign _6656_ = _6168_ & _6659_ /*36464*/;
assign _6657_ = _6168_ ^ _6659_ /*36467*/;
assign _6658_ = _6650_ & _6657_ /*36465*/;
assign _6655_ = _6656_ | _6658_ /*36463*/;
assign _6554_ = _6650_ ^ _6657_ /*36466*/;
assign _6664_ = D[10] ^ Q[47] /*36462*/;
assign _6661_ = _6169_ & _6664_ /*36458*/;
assign _6662_ = _6169_ ^ _6664_ /*36461*/;
assign _6663_ = _6655_ & _6662_ /*36459*/;
assign _6660_ = _6661_ | _6663_ /*36457*/;
assign _6555_ = _6655_ ^ _6662_ /*36460*/;
assign _6669_ = D[11] ^ Q[47] /*36456*/;
assign _6666_ = _6170_ & _6669_ /*36452*/;
assign _6667_ = _6170_ ^ _6669_ /*36455*/;
assign _6668_ = _6660_ & _6667_ /*36453*/;
assign _6665_ = _6666_ | _6668_ /*36451*/;
assign _6556_ = _6660_ ^ _6667_ /*36454*/;
assign _6674_ = D[12] ^ Q[47] /*36450*/;
assign _6671_ = _6171_ & _6674_ /*36446*/;
assign _6672_ = _6171_ ^ _6674_ /*36449*/;
assign _6673_ = _6665_ & _6672_ /*36447*/;
assign _6670_ = _6671_ | _6673_ /*36445*/;
assign _6557_ = _6665_ ^ _6672_ /*36448*/;
assign _6679_ = D[13] ^ Q[47] /*36444*/;
assign _6676_ = _6172_ & _6679_ /*36440*/;
assign _6677_ = _6172_ ^ _6679_ /*36443*/;
assign _6678_ = _6670_ & _6677_ /*36441*/;
assign _6675_ = _6676_ | _6678_ /*36439*/;
assign _6558_ = _6670_ ^ _6677_ /*36442*/;
assign _6684_ = D[14] ^ Q[47] /*36438*/;
assign _6681_ = _6173_ & _6684_ /*36434*/;
assign _6682_ = _6173_ ^ _6684_ /*36437*/;
assign _6683_ = _6675_ & _6682_ /*36435*/;
assign _6680_ = _6681_ | _6683_ /*36433*/;
assign _6559_ = _6675_ ^ _6682_ /*36436*/;
assign _6689_ = D[15] ^ Q[47] /*36432*/;
assign _6686_ = _6174_ & _6689_ /*36428*/;
assign _6687_ = _6174_ ^ _6689_ /*36431*/;
assign _6688_ = _6680_ & _6687_ /*36429*/;
assign _6685_ = _6686_ | _6688_ /*36427*/;
assign _6560_ = _6680_ ^ _6687_ /*36430*/;
assign _6694_ = D[16] ^ Q[47] /*36426*/;
assign _6691_ = _6175_ & _6694_ /*36422*/;
assign _6692_ = _6175_ ^ _6694_ /*36425*/;
assign _6693_ = _6685_ & _6692_ /*36423*/;
assign _6690_ = _6691_ | _6693_ /*36421*/;
assign _6561_ = _6685_ ^ _6692_ /*36424*/;
assign _6699_ = D[17] ^ Q[47] /*36420*/;
assign _6696_ = _6176_ & _6699_ /*36416*/;
assign _6697_ = _6176_ ^ _6699_ /*36419*/;
assign _6698_ = _6690_ & _6697_ /*36417*/;
assign _6695_ = _6696_ | _6698_ /*36415*/;
assign _6562_ = _6690_ ^ _6697_ /*36418*/;
assign _6704_ = D[18] ^ Q[47] /*36414*/;
assign _6701_ = _6177_ & _6704_ /*36410*/;
assign _6702_ = _6177_ ^ _6704_ /*36413*/;
assign _6703_ = _6695_ & _6702_ /*36411*/;
assign _6700_ = _6701_ | _6703_ /*36409*/;
assign _6563_ = _6695_ ^ _6702_ /*36412*/;
assign _6709_ = D[19] ^ Q[47] /*36408*/;
assign _6706_ = _6178_ & _6709_ /*36404*/;
assign _6707_ = _6178_ ^ _6709_ /*36407*/;
assign _6708_ = _6700_ & _6707_ /*36405*/;
assign _6705_ = _6706_ | _6708_ /*36403*/;
assign _6564_ = _6700_ ^ _6707_ /*36406*/;
assign _6714_ = D[20] ^ Q[47] /*36402*/;
assign _6711_ = _6179_ & _6714_ /*36398*/;
assign _6712_ = _6179_ ^ _6714_ /*36401*/;
assign _6713_ = _6705_ & _6712_ /*36399*/;
assign _6710_ = _6711_ | _6713_ /*36397*/;
assign _6565_ = _6705_ ^ _6712_ /*36400*/;
assign _6719_ = D[21] ^ Q[47] /*36396*/;
assign _6716_ = _6180_ & _6719_ /*36392*/;
assign _6717_ = _6180_ ^ _6719_ /*36395*/;
assign _6718_ = _6710_ & _6717_ /*36393*/;
assign _6715_ = _6716_ | _6718_ /*36391*/;
assign _6566_ = _6710_ ^ _6717_ /*36394*/;
assign _6724_ = D[22] ^ Q[47] /*36390*/;
assign _6721_ = _6181_ & _6724_ /*36386*/;
assign _6722_ = _6181_ ^ _6724_ /*36389*/;
assign _6723_ = _6715_ & _6722_ /*36387*/;
assign _6720_ = _6721_ | _6723_ /*36385*/;
assign _6567_ = _6715_ ^ _6722_ /*36388*/;
assign _6729_ = D[23] ^ Q[47] /*36384*/;
assign _6726_ = _6182_ & _6729_ /*36380*/;
assign _6727_ = _6182_ ^ _6729_ /*36383*/;
assign _6728_ = _6720_ & _6727_ /*36381*/;
assign _6725_ = _6726_ | _6728_ /*36379*/;
assign _6568_ = _6720_ ^ _6727_ /*36382*/;
assign _6734_ = D[24] ^ Q[47] /*36378*/;
assign _6731_ = _6183_ & _6734_ /*36374*/;
assign _6732_ = _6183_ ^ _6734_ /*36377*/;
assign _6733_ = _6725_ & _6732_ /*36375*/;
assign _6730_ = _6731_ | _6733_ /*36373*/;
assign _6569_ = _6725_ ^ _6732_ /*36376*/;
assign _6739_ = D[25] ^ Q[47] /*36372*/;
assign _6736_ = _6184_ & _6739_ /*36368*/;
assign _6737_ = _6184_ ^ _6739_ /*36371*/;
assign _6738_ = _6730_ & _6737_ /*36369*/;
assign _6735_ = _6736_ | _6738_ /*36367*/;
assign _6570_ = _6730_ ^ _6737_ /*36370*/;
assign _6744_ = D[26] ^ Q[47] /*36366*/;
assign _6741_ = _6185_ & _6744_ /*36362*/;
assign _6742_ = _6185_ ^ _6744_ /*36365*/;
assign _6743_ = _6735_ & _6742_ /*36363*/;
assign _6740_ = _6741_ | _6743_ /*36361*/;
assign _6571_ = _6735_ ^ _6742_ /*36364*/;
assign _6749_ = D[27] ^ Q[47] /*36360*/;
assign _6746_ = _6186_ & _6749_ /*36356*/;
assign _6747_ = _6186_ ^ _6749_ /*36359*/;
assign _6748_ = _6740_ & _6747_ /*36357*/;
assign _6745_ = _6746_ | _6748_ /*36355*/;
assign _6572_ = _6740_ ^ _6747_ /*36358*/;
assign _6754_ = D[28] ^ Q[47] /*36354*/;
assign _6751_ = _6187_ & _6754_ /*36350*/;
assign _6752_ = _6187_ ^ _6754_ /*36353*/;
assign _6753_ = _6745_ & _6752_ /*36351*/;
assign _6750_ = _6751_ | _6753_ /*36349*/;
assign _6573_ = _6745_ ^ _6752_ /*36352*/;
assign _6759_ = D[29] ^ Q[47] /*36348*/;
assign _6756_ = _6188_ & _6759_ /*36344*/;
assign _6757_ = _6188_ ^ _6759_ /*36347*/;
assign _6758_ = _6750_ & _6757_ /*36345*/;
assign _6755_ = _6756_ | _6758_ /*36343*/;
assign _6574_ = _6750_ ^ _6757_ /*36346*/;
assign _6764_ = D[30] ^ Q[47] /*36342*/;
assign _6761_ = _6189_ & _6764_ /*36338*/;
assign _6762_ = _6189_ ^ _6764_ /*36341*/;
assign _6763_ = _6755_ & _6762_ /*36339*/;
assign _6760_ = _6761_ | _6763_ /*36337*/;
assign _6575_ = _6755_ ^ _6762_ /*36340*/;
assign _6769_ = D[31] ^ Q[47] /*36336*/;
assign _6766_ = _6190_ & _6769_ /*36332*/;
assign _6767_ = _6190_ ^ _6769_ /*36335*/;
assign _6768_ = _6760_ & _6767_ /*36333*/;
assign _6765_ = _6766_ | _6768_ /*36331*/;
assign _6576_ = _6760_ ^ _6767_ /*36334*/;
assign _6774_ = D[32] ^ Q[47] /*36330*/;
assign _6771_ = _6191_ & _6774_ /*36326*/;
assign _6772_ = _6191_ ^ _6774_ /*36329*/;
assign _6773_ = _6765_ & _6772_ /*36327*/;
assign _6770_ = _6771_ | _6773_ /*36325*/;
assign _6577_ = _6765_ ^ _6772_ /*36328*/;
assign _6779_ = D[33] ^ Q[47] /*36324*/;
assign _6776_ = _6192_ & _6779_ /*36320*/;
assign _6777_ = _6192_ ^ _6779_ /*36323*/;
assign _6778_ = _6770_ & _6777_ /*36321*/;
assign _6775_ = _6776_ | _6778_ /*36319*/;
assign _6578_ = _6770_ ^ _6777_ /*36322*/;
assign _6784_ = D[34] ^ Q[47] /*36318*/;
assign _6781_ = _6193_ & _6784_ /*36314*/;
assign _6782_ = _6193_ ^ _6784_ /*36317*/;
assign _6783_ = _6775_ & _6782_ /*36315*/;
assign _6780_ = _6781_ | _6783_ /*36313*/;
assign _6579_ = _6775_ ^ _6782_ /*36316*/;
assign _6789_ = D[35] ^ Q[47] /*36312*/;
assign _6786_ = _6194_ & _6789_ /*36308*/;
assign _6787_ = _6194_ ^ _6789_ /*36311*/;
assign _6788_ = _6780_ & _6787_ /*36309*/;
assign _6785_ = _6786_ | _6788_ /*36307*/;
assign _6580_ = _6780_ ^ _6787_ /*36310*/;
assign _6794_ = D[36] ^ Q[47] /*36306*/;
assign _6791_ = _6195_ & _6794_ /*36302*/;
assign _6792_ = _6195_ ^ _6794_ /*36305*/;
assign _6793_ = _6785_ & _6792_ /*36303*/;
assign _6790_ = _6791_ | _6793_ /*36301*/;
assign _6581_ = _6785_ ^ _6792_ /*36304*/;
assign _6799_ = D[37] ^ Q[47] /*36300*/;
assign _6796_ = _6196_ & _6799_ /*36296*/;
assign _6797_ = _6196_ ^ _6799_ /*36299*/;
assign _6798_ = _6790_ & _6797_ /*36297*/;
assign _6795_ = _6796_ | _6798_ /*36295*/;
assign _6582_ = _6790_ ^ _6797_ /*36298*/;
assign _6804_ = D[38] ^ Q[47] /*36294*/;
assign _6801_ = _6197_ & _6804_ /*36290*/;
assign _6802_ = _6197_ ^ _6804_ /*36293*/;
assign _6803_ = _6795_ & _6802_ /*36291*/;
assign _6800_ = _6801_ | _6803_ /*36289*/;
assign _6583_ = _6795_ ^ _6802_ /*36292*/;
assign _6809_ = D[39] ^ Q[47] /*36288*/;
assign _6806_ = _6198_ & _6809_ /*36284*/;
assign _6807_ = _6198_ ^ _6809_ /*36287*/;
assign _6808_ = _6800_ & _6807_ /*36285*/;
assign _6805_ = _6806_ | _6808_ /*36283*/;
assign _6584_ = _6800_ ^ _6807_ /*36286*/;
assign _6814_ = D[40] ^ Q[47] /*36282*/;
assign _6811_ = _6199_ & _6814_ /*36278*/;
assign _6812_ = _6199_ ^ _6814_ /*36281*/;
assign _6813_ = _6805_ & _6812_ /*36279*/;
assign _6810_ = _6811_ | _6813_ /*36277*/;
assign _6585_ = _6805_ ^ _6812_ /*36280*/;
assign _6819_ = D[41] ^ Q[47] /*36276*/;
assign _6816_ = _6200_ & _6819_ /*36272*/;
assign _6817_ = _6200_ ^ _6819_ /*36275*/;
assign _6818_ = _6810_ & _6817_ /*36273*/;
assign _6815_ = _6816_ | _6818_ /*36271*/;
assign _6586_ = _6810_ ^ _6817_ /*36274*/;
assign _6824_ = D[42] ^ Q[47] /*36270*/;
assign _6821_ = _6201_ & _6824_ /*36266*/;
assign _6822_ = _6201_ ^ _6824_ /*36269*/;
assign _6823_ = _6815_ & _6822_ /*36267*/;
assign _6820_ = _6821_ | _6823_ /*36265*/;
assign _6587_ = _6815_ ^ _6822_ /*36268*/;
assign _6829_ = D[43] ^ Q[47] /*36264*/;
assign _6826_ = _6202_ & _6829_ /*36260*/;
assign _6827_ = _6202_ ^ _6829_ /*36263*/;
assign _6828_ = _6820_ & _6827_ /*36261*/;
assign _6825_ = _6826_ | _6828_ /*36259*/;
assign _6588_ = _6820_ ^ _6827_ /*36262*/;
assign _6834_ = D[44] ^ Q[47] /*36258*/;
assign _6831_ = _6203_ & _6834_ /*36254*/;
assign _6832_ = _6203_ ^ _6834_ /*36257*/;
assign _6833_ = _6825_ & _6832_ /*36255*/;
assign _6830_ = _6831_ | _6833_ /*36253*/;
assign _6589_ = _6825_ ^ _6832_ /*36256*/;
assign _6839_ = D[45] ^ Q[47] /*36252*/;
assign _6836_ = _6204_ & _6839_ /*36248*/;
assign _6837_ = _6204_ ^ _6839_ /*36251*/;
assign _6838_ = _6830_ & _6837_ /*36249*/;
assign _6835_ = _6836_ | _6838_ /*36247*/;
assign _6590_ = _6830_ ^ _6837_ /*36250*/;
assign _6844_ = D[46] ^ Q[47] /*36246*/;
assign _6841_ = _6205_ & _6844_ /*36242*/;
assign _6842_ = _6205_ ^ _6844_ /*36245*/;
assign _6843_ = _6835_ & _6842_ /*36243*/;
assign _6840_ = _6841_ | _6843_ /*36241*/;
assign _6591_ = _6835_ ^ _6842_ /*36244*/;
assign _6849_ = D[47] ^ Q[47] /*36240*/;
assign _6846_ = _6206_ & _6849_ /*36236*/;
assign _6847_ = _6206_ ^ _6849_ /*36239*/;
assign _6848_ = _6840_ & _6847_ /*36237*/;
assign _6845_ = _6846_ | _6848_ /*36235*/;
assign _6592_ = _6840_ ^ _6847_ /*36238*/;
assign _6854_ = D[48] ^ Q[47] /*36234*/;
assign _6851_ = _6207_ & _6854_ /*36230*/;
assign _6852_ = _6207_ ^ _6854_ /*36233*/;
assign _6853_ = _6845_ & _6852_ /*36231*/;
assign _6850_ = _6851_ | _6853_ /*36229*/;
assign _6593_ = _6845_ ^ _6852_ /*36232*/;
assign _6859_ = D[49] ^ Q[47] /*36228*/;
assign _6856_ = _6208_ & _6859_ /*36224*/;
assign _6857_ = _6208_ ^ _6859_ /*36227*/;
assign _6858_ = _6850_ & _6857_ /*36225*/;
assign _6855_ = _6856_ | _6858_ /*36223*/;
assign _6594_ = _6850_ ^ _6857_ /*36226*/;
assign _6864_ = D[50] ^ Q[47] /*36222*/;
assign _6861_ = _6209_ & _6864_ /*36218*/;
assign _6862_ = _6209_ ^ _6864_ /*36221*/;
assign _6863_ = _6855_ & _6862_ /*36219*/;
assign _6860_ = _6861_ | _6863_ /*36217*/;
assign _6595_ = _6855_ ^ _6862_ /*36220*/;
assign _6869_ = D[51] ^ Q[47] /*36216*/;
assign _6866_ = _6210_ & _6869_ /*36212*/;
assign _6867_ = _6210_ ^ _6869_ /*36215*/;
assign _6868_ = _6860_ & _6867_ /*36213*/;
assign _6865_ = _6866_ | _6868_ /*36211*/;
assign _6596_ = _6860_ ^ _6867_ /*36214*/;
assign _6874_ = D[52] ^ Q[47] /*36210*/;
assign _6871_ = _6211_ & _6874_ /*36206*/;
assign _6872_ = _6211_ ^ _6874_ /*36209*/;
assign _6873_ = _6865_ & _6872_ /*36207*/;
assign _6870_ = _6871_ | _6873_ /*36205*/;
assign _6597_ = _6865_ ^ _6872_ /*36208*/;
assign _6879_ = D[53] ^ Q[47] /*36204*/;
assign _6876_ = _6212_ & _6879_ /*36200*/;
assign _6877_ = _6212_ ^ _6879_ /*36203*/;
assign _6878_ = _6870_ & _6877_ /*36201*/;
assign _6875_ = _6876_ | _6878_ /*36199*/;
assign _6598_ = _6870_ ^ _6877_ /*36202*/;
assign _6884_ = D[54] ^ Q[47] /*36198*/;
assign _6881_ = _6213_ & _6884_ /*36194*/;
assign _6882_ = _6213_ ^ _6884_ /*36197*/;
assign _6883_ = _6875_ & _6882_ /*36195*/;
assign _6880_ = _6881_ | _6883_ /*36193*/;
assign _6599_ = _6875_ ^ _6882_ /*36196*/;
assign _6889_ = D[55] ^ Q[47] /*36192*/;
assign _6886_ = _6214_ & _6889_ /*36188*/;
assign _6887_ = _6214_ ^ _6889_ /*36191*/;
assign _6888_ = _6880_ & _6887_ /*36189*/;
assign _6885_ = _6886_ | _6888_ /*36187*/;
assign _6600_ = _6880_ ^ _6887_ /*36190*/;
assign _6894_ = D[56] ^ Q[47] /*36186*/;
assign _6891_ = _6215_ & _6894_ /*36182*/;
assign _6892_ = _6215_ ^ _6894_ /*36185*/;
assign _6893_ = _6885_ & _6892_ /*36183*/;
assign _6890_ = _6891_ | _6893_ /*36181*/;
assign _6601_ = _6885_ ^ _6892_ /*36184*/;
assign _6899_ = D[57] ^ Q[47] /*36180*/;
assign _6896_ = _6216_ & _6899_ /*36176*/;
assign _6897_ = _6216_ ^ _6899_ /*36179*/;
assign _6898_ = _6890_ & _6897_ /*36177*/;
assign _6895_ = _6896_ | _6898_ /*36175*/;
assign _6602_ = _6890_ ^ _6897_ /*36178*/;
assign _6904_ = D[58] ^ Q[47] /*36174*/;
assign _6901_ = _6217_ & _6904_ /*36170*/;
assign _6902_ = _6217_ ^ _6904_ /*36173*/;
assign _6903_ = _6895_ & _6902_ /*36171*/;
assign _6900_ = _6901_ | _6903_ /*36169*/;
assign _6603_ = _6895_ ^ _6902_ /*36172*/;
assign _6909_ = D[59] ^ Q[47] /*36168*/;
assign _6906_ = _6218_ & _6909_ /*36164*/;
assign _6907_ = _6218_ ^ _6909_ /*36167*/;
assign _6908_ = _6900_ & _6907_ /*36165*/;
assign _6905_ = _6906_ | _6908_ /*36163*/;
assign _6604_ = _6900_ ^ _6907_ /*36166*/;
assign _6914_ = D[60] ^ Q[47] /*36162*/;
assign _6911_ = _6219_ & _6914_ /*36158*/;
assign _6912_ = _6219_ ^ _6914_ /*36161*/;
assign _6913_ = _6905_ & _6912_ /*36159*/;
assign _6910_ = _6911_ | _6913_ /*36157*/;
assign _6605_ = _6905_ ^ _6912_ /*36160*/;
assign _6919_ = D[61] ^ Q[47] /*36156*/;
assign _6916_ = _6220_ & _6919_ /*36152*/;
assign _6917_ = _6220_ ^ _6919_ /*36155*/;
assign _6918_ = _6910_ & _6917_ /*36153*/;
assign _6915_ = _6916_ | _6918_ /*36151*/;
assign _6606_ = _6910_ ^ _6917_ /*36154*/;
assign _6924_ = D[62] ^ Q[47] /*36150*/;
assign _6921_ = _6221_ & _6924_ /*36146*/;
assign _6922_ = _6221_ ^ _6924_ /*36149*/;
assign _6923_ = _6915_ & _6922_ /*36147*/;
assign _6920_ = _6921_ | _6923_ /*36145*/;
assign _6607_ = _6915_ ^ _6922_ /*36148*/;
assign _6928_ = zeroWire ^ Q[47] /*36144*/;
assign _6925_ = _6222_ & _6928_ /*36140*/;
assign _6926_ = _6222_ ^ _6928_ /*36143*/;
assign _6927_ = _6920_ & _6926_ /*36141*/;
assign Q[46] = _6925_ | _6927_ /*36139*/;
assign _6608_ = _6920_ ^ _6926_ /*36142*/;
assign _6999_ = D[0] ^ Q[46] /*35753*/;
assign _6996_ = R_0[45] & _6999_ /*35749*/;
assign _6997_ = R_0[45] ^ _6999_ /*35752*/;
assign _6998_ = Q[46] & _6997_ /*35750*/;
assign _6995_ = _6996_ | _6998_ /*35748*/;
assign _6930_ = Q[46] ^ _6997_ /*35751*/;
assign _7004_ = D[1] ^ Q[46] /*35747*/;
assign _7001_ = _6545_ & _7004_ /*35743*/;
assign _7002_ = _6545_ ^ _7004_ /*35746*/;
assign _7003_ = _6995_ & _7002_ /*35744*/;
assign _7000_ = _7001_ | _7003_ /*35742*/;
assign _6931_ = _6995_ ^ _7002_ /*35745*/;
assign _7009_ = D[2] ^ Q[46] /*35741*/;
assign _7006_ = _6546_ & _7009_ /*35737*/;
assign _7007_ = _6546_ ^ _7009_ /*35740*/;
assign _7008_ = _7000_ & _7007_ /*35738*/;
assign _7005_ = _7006_ | _7008_ /*35736*/;
assign _6932_ = _7000_ ^ _7007_ /*35739*/;
assign _7014_ = D[3] ^ Q[46] /*35735*/;
assign _7011_ = _6547_ & _7014_ /*35731*/;
assign _7012_ = _6547_ ^ _7014_ /*35734*/;
assign _7013_ = _7005_ & _7012_ /*35732*/;
assign _7010_ = _7011_ | _7013_ /*35730*/;
assign _6933_ = _7005_ ^ _7012_ /*35733*/;
assign _7019_ = D[4] ^ Q[46] /*35729*/;
assign _7016_ = _6548_ & _7019_ /*35725*/;
assign _7017_ = _6548_ ^ _7019_ /*35728*/;
assign _7018_ = _7010_ & _7017_ /*35726*/;
assign _7015_ = _7016_ | _7018_ /*35724*/;
assign _6934_ = _7010_ ^ _7017_ /*35727*/;
assign _7024_ = D[5] ^ Q[46] /*35723*/;
assign _7021_ = _6549_ & _7024_ /*35719*/;
assign _7022_ = _6549_ ^ _7024_ /*35722*/;
assign _7023_ = _7015_ & _7022_ /*35720*/;
assign _7020_ = _7021_ | _7023_ /*35718*/;
assign _6935_ = _7015_ ^ _7022_ /*35721*/;
assign _7029_ = D[6] ^ Q[46] /*35717*/;
assign _7026_ = _6550_ & _7029_ /*35713*/;
assign _7027_ = _6550_ ^ _7029_ /*35716*/;
assign _7028_ = _7020_ & _7027_ /*35714*/;
assign _7025_ = _7026_ | _7028_ /*35712*/;
assign _6936_ = _7020_ ^ _7027_ /*35715*/;
assign _7034_ = D[7] ^ Q[46] /*35711*/;
assign _7031_ = _6551_ & _7034_ /*35707*/;
assign _7032_ = _6551_ ^ _7034_ /*35710*/;
assign _7033_ = _7025_ & _7032_ /*35708*/;
assign _7030_ = _7031_ | _7033_ /*35706*/;
assign _6937_ = _7025_ ^ _7032_ /*35709*/;
assign _7039_ = D[8] ^ Q[46] /*35705*/;
assign _7036_ = _6552_ & _7039_ /*35701*/;
assign _7037_ = _6552_ ^ _7039_ /*35704*/;
assign _7038_ = _7030_ & _7037_ /*35702*/;
assign _7035_ = _7036_ | _7038_ /*35700*/;
assign _6938_ = _7030_ ^ _7037_ /*35703*/;
assign _7044_ = D[9] ^ Q[46] /*35699*/;
assign _7041_ = _6553_ & _7044_ /*35695*/;
assign _7042_ = _6553_ ^ _7044_ /*35698*/;
assign _7043_ = _7035_ & _7042_ /*35696*/;
assign _7040_ = _7041_ | _7043_ /*35694*/;
assign _6939_ = _7035_ ^ _7042_ /*35697*/;
assign _7049_ = D[10] ^ Q[46] /*35693*/;
assign _7046_ = _6554_ & _7049_ /*35689*/;
assign _7047_ = _6554_ ^ _7049_ /*35692*/;
assign _7048_ = _7040_ & _7047_ /*35690*/;
assign _7045_ = _7046_ | _7048_ /*35688*/;
assign _6940_ = _7040_ ^ _7047_ /*35691*/;
assign _7054_ = D[11] ^ Q[46] /*35687*/;
assign _7051_ = _6555_ & _7054_ /*35683*/;
assign _7052_ = _6555_ ^ _7054_ /*35686*/;
assign _7053_ = _7045_ & _7052_ /*35684*/;
assign _7050_ = _7051_ | _7053_ /*35682*/;
assign _6941_ = _7045_ ^ _7052_ /*35685*/;
assign _7059_ = D[12] ^ Q[46] /*35681*/;
assign _7056_ = _6556_ & _7059_ /*35677*/;
assign _7057_ = _6556_ ^ _7059_ /*35680*/;
assign _7058_ = _7050_ & _7057_ /*35678*/;
assign _7055_ = _7056_ | _7058_ /*35676*/;
assign _6942_ = _7050_ ^ _7057_ /*35679*/;
assign _7064_ = D[13] ^ Q[46] /*35675*/;
assign _7061_ = _6557_ & _7064_ /*35671*/;
assign _7062_ = _6557_ ^ _7064_ /*35674*/;
assign _7063_ = _7055_ & _7062_ /*35672*/;
assign _7060_ = _7061_ | _7063_ /*35670*/;
assign _6943_ = _7055_ ^ _7062_ /*35673*/;
assign _7069_ = D[14] ^ Q[46] /*35669*/;
assign _7066_ = _6558_ & _7069_ /*35665*/;
assign _7067_ = _6558_ ^ _7069_ /*35668*/;
assign _7068_ = _7060_ & _7067_ /*35666*/;
assign _7065_ = _7066_ | _7068_ /*35664*/;
assign _6944_ = _7060_ ^ _7067_ /*35667*/;
assign _7074_ = D[15] ^ Q[46] /*35663*/;
assign _7071_ = _6559_ & _7074_ /*35659*/;
assign _7072_ = _6559_ ^ _7074_ /*35662*/;
assign _7073_ = _7065_ & _7072_ /*35660*/;
assign _7070_ = _7071_ | _7073_ /*35658*/;
assign _6945_ = _7065_ ^ _7072_ /*35661*/;
assign _7079_ = D[16] ^ Q[46] /*35657*/;
assign _7076_ = _6560_ & _7079_ /*35653*/;
assign _7077_ = _6560_ ^ _7079_ /*35656*/;
assign _7078_ = _7070_ & _7077_ /*35654*/;
assign _7075_ = _7076_ | _7078_ /*35652*/;
assign _6946_ = _7070_ ^ _7077_ /*35655*/;
assign _7084_ = D[17] ^ Q[46] /*35651*/;
assign _7081_ = _6561_ & _7084_ /*35647*/;
assign _7082_ = _6561_ ^ _7084_ /*35650*/;
assign _7083_ = _7075_ & _7082_ /*35648*/;
assign _7080_ = _7081_ | _7083_ /*35646*/;
assign _6947_ = _7075_ ^ _7082_ /*35649*/;
assign _7089_ = D[18] ^ Q[46] /*35645*/;
assign _7086_ = _6562_ & _7089_ /*35641*/;
assign _7087_ = _6562_ ^ _7089_ /*35644*/;
assign _7088_ = _7080_ & _7087_ /*35642*/;
assign _7085_ = _7086_ | _7088_ /*35640*/;
assign _6948_ = _7080_ ^ _7087_ /*35643*/;
assign _7094_ = D[19] ^ Q[46] /*35639*/;
assign _7091_ = _6563_ & _7094_ /*35635*/;
assign _7092_ = _6563_ ^ _7094_ /*35638*/;
assign _7093_ = _7085_ & _7092_ /*35636*/;
assign _7090_ = _7091_ | _7093_ /*35634*/;
assign _6949_ = _7085_ ^ _7092_ /*35637*/;
assign _7099_ = D[20] ^ Q[46] /*35633*/;
assign _7096_ = _6564_ & _7099_ /*35629*/;
assign _7097_ = _6564_ ^ _7099_ /*35632*/;
assign _7098_ = _7090_ & _7097_ /*35630*/;
assign _7095_ = _7096_ | _7098_ /*35628*/;
assign _6950_ = _7090_ ^ _7097_ /*35631*/;
assign _7104_ = D[21] ^ Q[46] /*35627*/;
assign _7101_ = _6565_ & _7104_ /*35623*/;
assign _7102_ = _6565_ ^ _7104_ /*35626*/;
assign _7103_ = _7095_ & _7102_ /*35624*/;
assign _7100_ = _7101_ | _7103_ /*35622*/;
assign _6951_ = _7095_ ^ _7102_ /*35625*/;
assign _7109_ = D[22] ^ Q[46] /*35621*/;
assign _7106_ = _6566_ & _7109_ /*35617*/;
assign _7107_ = _6566_ ^ _7109_ /*35620*/;
assign _7108_ = _7100_ & _7107_ /*35618*/;
assign _7105_ = _7106_ | _7108_ /*35616*/;
assign _6952_ = _7100_ ^ _7107_ /*35619*/;
assign _7114_ = D[23] ^ Q[46] /*35615*/;
assign _7111_ = _6567_ & _7114_ /*35611*/;
assign _7112_ = _6567_ ^ _7114_ /*35614*/;
assign _7113_ = _7105_ & _7112_ /*35612*/;
assign _7110_ = _7111_ | _7113_ /*35610*/;
assign _6953_ = _7105_ ^ _7112_ /*35613*/;
assign _7119_ = D[24] ^ Q[46] /*35609*/;
assign _7116_ = _6568_ & _7119_ /*35605*/;
assign _7117_ = _6568_ ^ _7119_ /*35608*/;
assign _7118_ = _7110_ & _7117_ /*35606*/;
assign _7115_ = _7116_ | _7118_ /*35604*/;
assign _6954_ = _7110_ ^ _7117_ /*35607*/;
assign _7124_ = D[25] ^ Q[46] /*35603*/;
assign _7121_ = _6569_ & _7124_ /*35599*/;
assign _7122_ = _6569_ ^ _7124_ /*35602*/;
assign _7123_ = _7115_ & _7122_ /*35600*/;
assign _7120_ = _7121_ | _7123_ /*35598*/;
assign _6955_ = _7115_ ^ _7122_ /*35601*/;
assign _7129_ = D[26] ^ Q[46] /*35597*/;
assign _7126_ = _6570_ & _7129_ /*35593*/;
assign _7127_ = _6570_ ^ _7129_ /*35596*/;
assign _7128_ = _7120_ & _7127_ /*35594*/;
assign _7125_ = _7126_ | _7128_ /*35592*/;
assign _6956_ = _7120_ ^ _7127_ /*35595*/;
assign _7134_ = D[27] ^ Q[46] /*35591*/;
assign _7131_ = _6571_ & _7134_ /*35587*/;
assign _7132_ = _6571_ ^ _7134_ /*35590*/;
assign _7133_ = _7125_ & _7132_ /*35588*/;
assign _7130_ = _7131_ | _7133_ /*35586*/;
assign _6957_ = _7125_ ^ _7132_ /*35589*/;
assign _7139_ = D[28] ^ Q[46] /*35585*/;
assign _7136_ = _6572_ & _7139_ /*35581*/;
assign _7137_ = _6572_ ^ _7139_ /*35584*/;
assign _7138_ = _7130_ & _7137_ /*35582*/;
assign _7135_ = _7136_ | _7138_ /*35580*/;
assign _6958_ = _7130_ ^ _7137_ /*35583*/;
assign _7144_ = D[29] ^ Q[46] /*35579*/;
assign _7141_ = _6573_ & _7144_ /*35575*/;
assign _7142_ = _6573_ ^ _7144_ /*35578*/;
assign _7143_ = _7135_ & _7142_ /*35576*/;
assign _7140_ = _7141_ | _7143_ /*35574*/;
assign _6959_ = _7135_ ^ _7142_ /*35577*/;
assign _7149_ = D[30] ^ Q[46] /*35573*/;
assign _7146_ = _6574_ & _7149_ /*35569*/;
assign _7147_ = _6574_ ^ _7149_ /*35572*/;
assign _7148_ = _7140_ & _7147_ /*35570*/;
assign _7145_ = _7146_ | _7148_ /*35568*/;
assign _6960_ = _7140_ ^ _7147_ /*35571*/;
assign _7154_ = D[31] ^ Q[46] /*35567*/;
assign _7151_ = _6575_ & _7154_ /*35563*/;
assign _7152_ = _6575_ ^ _7154_ /*35566*/;
assign _7153_ = _7145_ & _7152_ /*35564*/;
assign _7150_ = _7151_ | _7153_ /*35562*/;
assign _6961_ = _7145_ ^ _7152_ /*35565*/;
assign _7159_ = D[32] ^ Q[46] /*35561*/;
assign _7156_ = _6576_ & _7159_ /*35557*/;
assign _7157_ = _6576_ ^ _7159_ /*35560*/;
assign _7158_ = _7150_ & _7157_ /*35558*/;
assign _7155_ = _7156_ | _7158_ /*35556*/;
assign _6962_ = _7150_ ^ _7157_ /*35559*/;
assign _7164_ = D[33] ^ Q[46] /*35555*/;
assign _7161_ = _6577_ & _7164_ /*35551*/;
assign _7162_ = _6577_ ^ _7164_ /*35554*/;
assign _7163_ = _7155_ & _7162_ /*35552*/;
assign _7160_ = _7161_ | _7163_ /*35550*/;
assign _6963_ = _7155_ ^ _7162_ /*35553*/;
assign _7169_ = D[34] ^ Q[46] /*35549*/;
assign _7166_ = _6578_ & _7169_ /*35545*/;
assign _7167_ = _6578_ ^ _7169_ /*35548*/;
assign _7168_ = _7160_ & _7167_ /*35546*/;
assign _7165_ = _7166_ | _7168_ /*35544*/;
assign _6964_ = _7160_ ^ _7167_ /*35547*/;
assign _7174_ = D[35] ^ Q[46] /*35543*/;
assign _7171_ = _6579_ & _7174_ /*35539*/;
assign _7172_ = _6579_ ^ _7174_ /*35542*/;
assign _7173_ = _7165_ & _7172_ /*35540*/;
assign _7170_ = _7171_ | _7173_ /*35538*/;
assign _6965_ = _7165_ ^ _7172_ /*35541*/;
assign _7179_ = D[36] ^ Q[46] /*35537*/;
assign _7176_ = _6580_ & _7179_ /*35533*/;
assign _7177_ = _6580_ ^ _7179_ /*35536*/;
assign _7178_ = _7170_ & _7177_ /*35534*/;
assign _7175_ = _7176_ | _7178_ /*35532*/;
assign _6966_ = _7170_ ^ _7177_ /*35535*/;
assign _7184_ = D[37] ^ Q[46] /*35531*/;
assign _7181_ = _6581_ & _7184_ /*35527*/;
assign _7182_ = _6581_ ^ _7184_ /*35530*/;
assign _7183_ = _7175_ & _7182_ /*35528*/;
assign _7180_ = _7181_ | _7183_ /*35526*/;
assign _6967_ = _7175_ ^ _7182_ /*35529*/;
assign _7189_ = D[38] ^ Q[46] /*35525*/;
assign _7186_ = _6582_ & _7189_ /*35521*/;
assign _7187_ = _6582_ ^ _7189_ /*35524*/;
assign _7188_ = _7180_ & _7187_ /*35522*/;
assign _7185_ = _7186_ | _7188_ /*35520*/;
assign _6968_ = _7180_ ^ _7187_ /*35523*/;
assign _7194_ = D[39] ^ Q[46] /*35519*/;
assign _7191_ = _6583_ & _7194_ /*35515*/;
assign _7192_ = _6583_ ^ _7194_ /*35518*/;
assign _7193_ = _7185_ & _7192_ /*35516*/;
assign _7190_ = _7191_ | _7193_ /*35514*/;
assign _6969_ = _7185_ ^ _7192_ /*35517*/;
assign _7199_ = D[40] ^ Q[46] /*35513*/;
assign _7196_ = _6584_ & _7199_ /*35509*/;
assign _7197_ = _6584_ ^ _7199_ /*35512*/;
assign _7198_ = _7190_ & _7197_ /*35510*/;
assign _7195_ = _7196_ | _7198_ /*35508*/;
assign _6970_ = _7190_ ^ _7197_ /*35511*/;
assign _7204_ = D[41] ^ Q[46] /*35507*/;
assign _7201_ = _6585_ & _7204_ /*35503*/;
assign _7202_ = _6585_ ^ _7204_ /*35506*/;
assign _7203_ = _7195_ & _7202_ /*35504*/;
assign _7200_ = _7201_ | _7203_ /*35502*/;
assign _6971_ = _7195_ ^ _7202_ /*35505*/;
assign _7209_ = D[42] ^ Q[46] /*35501*/;
assign _7206_ = _6586_ & _7209_ /*35497*/;
assign _7207_ = _6586_ ^ _7209_ /*35500*/;
assign _7208_ = _7200_ & _7207_ /*35498*/;
assign _7205_ = _7206_ | _7208_ /*35496*/;
assign _6972_ = _7200_ ^ _7207_ /*35499*/;
assign _7214_ = D[43] ^ Q[46] /*35495*/;
assign _7211_ = _6587_ & _7214_ /*35491*/;
assign _7212_ = _6587_ ^ _7214_ /*35494*/;
assign _7213_ = _7205_ & _7212_ /*35492*/;
assign _7210_ = _7211_ | _7213_ /*35490*/;
assign _6973_ = _7205_ ^ _7212_ /*35493*/;
assign _7219_ = D[44] ^ Q[46] /*35489*/;
assign _7216_ = _6588_ & _7219_ /*35485*/;
assign _7217_ = _6588_ ^ _7219_ /*35488*/;
assign _7218_ = _7210_ & _7217_ /*35486*/;
assign _7215_ = _7216_ | _7218_ /*35484*/;
assign _6974_ = _7210_ ^ _7217_ /*35487*/;
assign _7224_ = D[45] ^ Q[46] /*35483*/;
assign _7221_ = _6589_ & _7224_ /*35479*/;
assign _7222_ = _6589_ ^ _7224_ /*35482*/;
assign _7223_ = _7215_ & _7222_ /*35480*/;
assign _7220_ = _7221_ | _7223_ /*35478*/;
assign _6975_ = _7215_ ^ _7222_ /*35481*/;
assign _7229_ = D[46] ^ Q[46] /*35477*/;
assign _7226_ = _6590_ & _7229_ /*35473*/;
assign _7227_ = _6590_ ^ _7229_ /*35476*/;
assign _7228_ = _7220_ & _7227_ /*35474*/;
assign _7225_ = _7226_ | _7228_ /*35472*/;
assign _6976_ = _7220_ ^ _7227_ /*35475*/;
assign _7234_ = D[47] ^ Q[46] /*35471*/;
assign _7231_ = _6591_ & _7234_ /*35467*/;
assign _7232_ = _6591_ ^ _7234_ /*35470*/;
assign _7233_ = _7225_ & _7232_ /*35468*/;
assign _7230_ = _7231_ | _7233_ /*35466*/;
assign _6977_ = _7225_ ^ _7232_ /*35469*/;
assign _7239_ = D[48] ^ Q[46] /*35465*/;
assign _7236_ = _6592_ & _7239_ /*35461*/;
assign _7237_ = _6592_ ^ _7239_ /*35464*/;
assign _7238_ = _7230_ & _7237_ /*35462*/;
assign _7235_ = _7236_ | _7238_ /*35460*/;
assign _6978_ = _7230_ ^ _7237_ /*35463*/;
assign _7244_ = D[49] ^ Q[46] /*35459*/;
assign _7241_ = _6593_ & _7244_ /*35455*/;
assign _7242_ = _6593_ ^ _7244_ /*35458*/;
assign _7243_ = _7235_ & _7242_ /*35456*/;
assign _7240_ = _7241_ | _7243_ /*35454*/;
assign _6979_ = _7235_ ^ _7242_ /*35457*/;
assign _7249_ = D[50] ^ Q[46] /*35453*/;
assign _7246_ = _6594_ & _7249_ /*35449*/;
assign _7247_ = _6594_ ^ _7249_ /*35452*/;
assign _7248_ = _7240_ & _7247_ /*35450*/;
assign _7245_ = _7246_ | _7248_ /*35448*/;
assign _6980_ = _7240_ ^ _7247_ /*35451*/;
assign _7254_ = D[51] ^ Q[46] /*35447*/;
assign _7251_ = _6595_ & _7254_ /*35443*/;
assign _7252_ = _6595_ ^ _7254_ /*35446*/;
assign _7253_ = _7245_ & _7252_ /*35444*/;
assign _7250_ = _7251_ | _7253_ /*35442*/;
assign _6981_ = _7245_ ^ _7252_ /*35445*/;
assign _7259_ = D[52] ^ Q[46] /*35441*/;
assign _7256_ = _6596_ & _7259_ /*35437*/;
assign _7257_ = _6596_ ^ _7259_ /*35440*/;
assign _7258_ = _7250_ & _7257_ /*35438*/;
assign _7255_ = _7256_ | _7258_ /*35436*/;
assign _6982_ = _7250_ ^ _7257_ /*35439*/;
assign _7264_ = D[53] ^ Q[46] /*35435*/;
assign _7261_ = _6597_ & _7264_ /*35431*/;
assign _7262_ = _6597_ ^ _7264_ /*35434*/;
assign _7263_ = _7255_ & _7262_ /*35432*/;
assign _7260_ = _7261_ | _7263_ /*35430*/;
assign _6983_ = _7255_ ^ _7262_ /*35433*/;
assign _7269_ = D[54] ^ Q[46] /*35429*/;
assign _7266_ = _6598_ & _7269_ /*35425*/;
assign _7267_ = _6598_ ^ _7269_ /*35428*/;
assign _7268_ = _7260_ & _7267_ /*35426*/;
assign _7265_ = _7266_ | _7268_ /*35424*/;
assign _6984_ = _7260_ ^ _7267_ /*35427*/;
assign _7274_ = D[55] ^ Q[46] /*35423*/;
assign _7271_ = _6599_ & _7274_ /*35419*/;
assign _7272_ = _6599_ ^ _7274_ /*35422*/;
assign _7273_ = _7265_ & _7272_ /*35420*/;
assign _7270_ = _7271_ | _7273_ /*35418*/;
assign _6985_ = _7265_ ^ _7272_ /*35421*/;
assign _7279_ = D[56] ^ Q[46] /*35417*/;
assign _7276_ = _6600_ & _7279_ /*35413*/;
assign _7277_ = _6600_ ^ _7279_ /*35416*/;
assign _7278_ = _7270_ & _7277_ /*35414*/;
assign _7275_ = _7276_ | _7278_ /*35412*/;
assign _6986_ = _7270_ ^ _7277_ /*35415*/;
assign _7284_ = D[57] ^ Q[46] /*35411*/;
assign _7281_ = _6601_ & _7284_ /*35407*/;
assign _7282_ = _6601_ ^ _7284_ /*35410*/;
assign _7283_ = _7275_ & _7282_ /*35408*/;
assign _7280_ = _7281_ | _7283_ /*35406*/;
assign _6987_ = _7275_ ^ _7282_ /*35409*/;
assign _7289_ = D[58] ^ Q[46] /*35405*/;
assign _7286_ = _6602_ & _7289_ /*35401*/;
assign _7287_ = _6602_ ^ _7289_ /*35404*/;
assign _7288_ = _7280_ & _7287_ /*35402*/;
assign _7285_ = _7286_ | _7288_ /*35400*/;
assign _6988_ = _7280_ ^ _7287_ /*35403*/;
assign _7294_ = D[59] ^ Q[46] /*35399*/;
assign _7291_ = _6603_ & _7294_ /*35395*/;
assign _7292_ = _6603_ ^ _7294_ /*35398*/;
assign _7293_ = _7285_ & _7292_ /*35396*/;
assign _7290_ = _7291_ | _7293_ /*35394*/;
assign _6989_ = _7285_ ^ _7292_ /*35397*/;
assign _7299_ = D[60] ^ Q[46] /*35393*/;
assign _7296_ = _6604_ & _7299_ /*35389*/;
assign _7297_ = _6604_ ^ _7299_ /*35392*/;
assign _7298_ = _7290_ & _7297_ /*35390*/;
assign _7295_ = _7296_ | _7298_ /*35388*/;
assign _6990_ = _7290_ ^ _7297_ /*35391*/;
assign _7304_ = D[61] ^ Q[46] /*35387*/;
assign _7301_ = _6605_ & _7304_ /*35383*/;
assign _7302_ = _6605_ ^ _7304_ /*35386*/;
assign _7303_ = _7295_ & _7302_ /*35384*/;
assign _7300_ = _7301_ | _7303_ /*35382*/;
assign _6991_ = _7295_ ^ _7302_ /*35385*/;
assign _7309_ = D[62] ^ Q[46] /*35381*/;
assign _7306_ = _6606_ & _7309_ /*35377*/;
assign _7307_ = _6606_ ^ _7309_ /*35380*/;
assign _7308_ = _7300_ & _7307_ /*35378*/;
assign _7305_ = _7306_ | _7308_ /*35376*/;
assign _6992_ = _7300_ ^ _7307_ /*35379*/;
assign _7313_ = zeroWire ^ Q[46] /*35375*/;
assign _7310_ = _6607_ & _7313_ /*35371*/;
assign _7311_ = _6607_ ^ _7313_ /*35374*/;
assign _7312_ = _7305_ & _7311_ /*35372*/;
assign Q[45] = _7310_ | _7312_ /*35370*/;
assign _6993_ = _7305_ ^ _7311_ /*35373*/;
assign _7384_ = D[0] ^ Q[45] /*34984*/;
assign _7381_ = R_0[44] & _7384_ /*34980*/;
assign _7382_ = R_0[44] ^ _7384_ /*34983*/;
assign _7383_ = Q[45] & _7382_ /*34981*/;
assign _7380_ = _7381_ | _7383_ /*34979*/;
assign _7315_ = Q[45] ^ _7382_ /*34982*/;
assign _7389_ = D[1] ^ Q[45] /*34978*/;
assign _7386_ = _6930_ & _7389_ /*34974*/;
assign _7387_ = _6930_ ^ _7389_ /*34977*/;
assign _7388_ = _7380_ & _7387_ /*34975*/;
assign _7385_ = _7386_ | _7388_ /*34973*/;
assign _7316_ = _7380_ ^ _7387_ /*34976*/;
assign _7394_ = D[2] ^ Q[45] /*34972*/;
assign _7391_ = _6931_ & _7394_ /*34968*/;
assign _7392_ = _6931_ ^ _7394_ /*34971*/;
assign _7393_ = _7385_ & _7392_ /*34969*/;
assign _7390_ = _7391_ | _7393_ /*34967*/;
assign _7317_ = _7385_ ^ _7392_ /*34970*/;
assign _7399_ = D[3] ^ Q[45] /*34966*/;
assign _7396_ = _6932_ & _7399_ /*34962*/;
assign _7397_ = _6932_ ^ _7399_ /*34965*/;
assign _7398_ = _7390_ & _7397_ /*34963*/;
assign _7395_ = _7396_ | _7398_ /*34961*/;
assign _7318_ = _7390_ ^ _7397_ /*34964*/;
assign _7404_ = D[4] ^ Q[45] /*34960*/;
assign _7401_ = _6933_ & _7404_ /*34956*/;
assign _7402_ = _6933_ ^ _7404_ /*34959*/;
assign _7403_ = _7395_ & _7402_ /*34957*/;
assign _7400_ = _7401_ | _7403_ /*34955*/;
assign _7319_ = _7395_ ^ _7402_ /*34958*/;
assign _7409_ = D[5] ^ Q[45] /*34954*/;
assign _7406_ = _6934_ & _7409_ /*34950*/;
assign _7407_ = _6934_ ^ _7409_ /*34953*/;
assign _7408_ = _7400_ & _7407_ /*34951*/;
assign _7405_ = _7406_ | _7408_ /*34949*/;
assign _7320_ = _7400_ ^ _7407_ /*34952*/;
assign _7414_ = D[6] ^ Q[45] /*34948*/;
assign _7411_ = _6935_ & _7414_ /*34944*/;
assign _7412_ = _6935_ ^ _7414_ /*34947*/;
assign _7413_ = _7405_ & _7412_ /*34945*/;
assign _7410_ = _7411_ | _7413_ /*34943*/;
assign _7321_ = _7405_ ^ _7412_ /*34946*/;
assign _7419_ = D[7] ^ Q[45] /*34942*/;
assign _7416_ = _6936_ & _7419_ /*34938*/;
assign _7417_ = _6936_ ^ _7419_ /*34941*/;
assign _7418_ = _7410_ & _7417_ /*34939*/;
assign _7415_ = _7416_ | _7418_ /*34937*/;
assign _7322_ = _7410_ ^ _7417_ /*34940*/;
assign _7424_ = D[8] ^ Q[45] /*34936*/;
assign _7421_ = _6937_ & _7424_ /*34932*/;
assign _7422_ = _6937_ ^ _7424_ /*34935*/;
assign _7423_ = _7415_ & _7422_ /*34933*/;
assign _7420_ = _7421_ | _7423_ /*34931*/;
assign _7323_ = _7415_ ^ _7422_ /*34934*/;
assign _7429_ = D[9] ^ Q[45] /*34930*/;
assign _7426_ = _6938_ & _7429_ /*34926*/;
assign _7427_ = _6938_ ^ _7429_ /*34929*/;
assign _7428_ = _7420_ & _7427_ /*34927*/;
assign _7425_ = _7426_ | _7428_ /*34925*/;
assign _7324_ = _7420_ ^ _7427_ /*34928*/;
assign _7434_ = D[10] ^ Q[45] /*34924*/;
assign _7431_ = _6939_ & _7434_ /*34920*/;
assign _7432_ = _6939_ ^ _7434_ /*34923*/;
assign _7433_ = _7425_ & _7432_ /*34921*/;
assign _7430_ = _7431_ | _7433_ /*34919*/;
assign _7325_ = _7425_ ^ _7432_ /*34922*/;
assign _7439_ = D[11] ^ Q[45] /*34918*/;
assign _7436_ = _6940_ & _7439_ /*34914*/;
assign _7437_ = _6940_ ^ _7439_ /*34917*/;
assign _7438_ = _7430_ & _7437_ /*34915*/;
assign _7435_ = _7436_ | _7438_ /*34913*/;
assign _7326_ = _7430_ ^ _7437_ /*34916*/;
assign _7444_ = D[12] ^ Q[45] /*34912*/;
assign _7441_ = _6941_ & _7444_ /*34908*/;
assign _7442_ = _6941_ ^ _7444_ /*34911*/;
assign _7443_ = _7435_ & _7442_ /*34909*/;
assign _7440_ = _7441_ | _7443_ /*34907*/;
assign _7327_ = _7435_ ^ _7442_ /*34910*/;
assign _7449_ = D[13] ^ Q[45] /*34906*/;
assign _7446_ = _6942_ & _7449_ /*34902*/;
assign _7447_ = _6942_ ^ _7449_ /*34905*/;
assign _7448_ = _7440_ & _7447_ /*34903*/;
assign _7445_ = _7446_ | _7448_ /*34901*/;
assign _7328_ = _7440_ ^ _7447_ /*34904*/;
assign _7454_ = D[14] ^ Q[45] /*34900*/;
assign _7451_ = _6943_ & _7454_ /*34896*/;
assign _7452_ = _6943_ ^ _7454_ /*34899*/;
assign _7453_ = _7445_ & _7452_ /*34897*/;
assign _7450_ = _7451_ | _7453_ /*34895*/;
assign _7329_ = _7445_ ^ _7452_ /*34898*/;
assign _7459_ = D[15] ^ Q[45] /*34894*/;
assign _7456_ = _6944_ & _7459_ /*34890*/;
assign _7457_ = _6944_ ^ _7459_ /*34893*/;
assign _7458_ = _7450_ & _7457_ /*34891*/;
assign _7455_ = _7456_ | _7458_ /*34889*/;
assign _7330_ = _7450_ ^ _7457_ /*34892*/;
assign _7464_ = D[16] ^ Q[45] /*34888*/;
assign _7461_ = _6945_ & _7464_ /*34884*/;
assign _7462_ = _6945_ ^ _7464_ /*34887*/;
assign _7463_ = _7455_ & _7462_ /*34885*/;
assign _7460_ = _7461_ | _7463_ /*34883*/;
assign _7331_ = _7455_ ^ _7462_ /*34886*/;
assign _7469_ = D[17] ^ Q[45] /*34882*/;
assign _7466_ = _6946_ & _7469_ /*34878*/;
assign _7467_ = _6946_ ^ _7469_ /*34881*/;
assign _7468_ = _7460_ & _7467_ /*34879*/;
assign _7465_ = _7466_ | _7468_ /*34877*/;
assign _7332_ = _7460_ ^ _7467_ /*34880*/;
assign _7474_ = D[18] ^ Q[45] /*34876*/;
assign _7471_ = _6947_ & _7474_ /*34872*/;
assign _7472_ = _6947_ ^ _7474_ /*34875*/;
assign _7473_ = _7465_ & _7472_ /*34873*/;
assign _7470_ = _7471_ | _7473_ /*34871*/;
assign _7333_ = _7465_ ^ _7472_ /*34874*/;
assign _7479_ = D[19] ^ Q[45] /*34870*/;
assign _7476_ = _6948_ & _7479_ /*34866*/;
assign _7477_ = _6948_ ^ _7479_ /*34869*/;
assign _7478_ = _7470_ & _7477_ /*34867*/;
assign _7475_ = _7476_ | _7478_ /*34865*/;
assign _7334_ = _7470_ ^ _7477_ /*34868*/;
assign _7484_ = D[20] ^ Q[45] /*34864*/;
assign _7481_ = _6949_ & _7484_ /*34860*/;
assign _7482_ = _6949_ ^ _7484_ /*34863*/;
assign _7483_ = _7475_ & _7482_ /*34861*/;
assign _7480_ = _7481_ | _7483_ /*34859*/;
assign _7335_ = _7475_ ^ _7482_ /*34862*/;
assign _7489_ = D[21] ^ Q[45] /*34858*/;
assign _7486_ = _6950_ & _7489_ /*34854*/;
assign _7487_ = _6950_ ^ _7489_ /*34857*/;
assign _7488_ = _7480_ & _7487_ /*34855*/;
assign _7485_ = _7486_ | _7488_ /*34853*/;
assign _7336_ = _7480_ ^ _7487_ /*34856*/;
assign _7494_ = D[22] ^ Q[45] /*34852*/;
assign _7491_ = _6951_ & _7494_ /*34848*/;
assign _7492_ = _6951_ ^ _7494_ /*34851*/;
assign _7493_ = _7485_ & _7492_ /*34849*/;
assign _7490_ = _7491_ | _7493_ /*34847*/;
assign _7337_ = _7485_ ^ _7492_ /*34850*/;
assign _7499_ = D[23] ^ Q[45] /*34846*/;
assign _7496_ = _6952_ & _7499_ /*34842*/;
assign _7497_ = _6952_ ^ _7499_ /*34845*/;
assign _7498_ = _7490_ & _7497_ /*34843*/;
assign _7495_ = _7496_ | _7498_ /*34841*/;
assign _7338_ = _7490_ ^ _7497_ /*34844*/;
assign _7504_ = D[24] ^ Q[45] /*34840*/;
assign _7501_ = _6953_ & _7504_ /*34836*/;
assign _7502_ = _6953_ ^ _7504_ /*34839*/;
assign _7503_ = _7495_ & _7502_ /*34837*/;
assign _7500_ = _7501_ | _7503_ /*34835*/;
assign _7339_ = _7495_ ^ _7502_ /*34838*/;
assign _7509_ = D[25] ^ Q[45] /*34834*/;
assign _7506_ = _6954_ & _7509_ /*34830*/;
assign _7507_ = _6954_ ^ _7509_ /*34833*/;
assign _7508_ = _7500_ & _7507_ /*34831*/;
assign _7505_ = _7506_ | _7508_ /*34829*/;
assign _7340_ = _7500_ ^ _7507_ /*34832*/;
assign _7514_ = D[26] ^ Q[45] /*34828*/;
assign _7511_ = _6955_ & _7514_ /*34824*/;
assign _7512_ = _6955_ ^ _7514_ /*34827*/;
assign _7513_ = _7505_ & _7512_ /*34825*/;
assign _7510_ = _7511_ | _7513_ /*34823*/;
assign _7341_ = _7505_ ^ _7512_ /*34826*/;
assign _7519_ = D[27] ^ Q[45] /*34822*/;
assign _7516_ = _6956_ & _7519_ /*34818*/;
assign _7517_ = _6956_ ^ _7519_ /*34821*/;
assign _7518_ = _7510_ & _7517_ /*34819*/;
assign _7515_ = _7516_ | _7518_ /*34817*/;
assign _7342_ = _7510_ ^ _7517_ /*34820*/;
assign _7524_ = D[28] ^ Q[45] /*34816*/;
assign _7521_ = _6957_ & _7524_ /*34812*/;
assign _7522_ = _6957_ ^ _7524_ /*34815*/;
assign _7523_ = _7515_ & _7522_ /*34813*/;
assign _7520_ = _7521_ | _7523_ /*34811*/;
assign _7343_ = _7515_ ^ _7522_ /*34814*/;
assign _7529_ = D[29] ^ Q[45] /*34810*/;
assign _7526_ = _6958_ & _7529_ /*34806*/;
assign _7527_ = _6958_ ^ _7529_ /*34809*/;
assign _7528_ = _7520_ & _7527_ /*34807*/;
assign _7525_ = _7526_ | _7528_ /*34805*/;
assign _7344_ = _7520_ ^ _7527_ /*34808*/;
assign _7534_ = D[30] ^ Q[45] /*34804*/;
assign _7531_ = _6959_ & _7534_ /*34800*/;
assign _7532_ = _6959_ ^ _7534_ /*34803*/;
assign _7533_ = _7525_ & _7532_ /*34801*/;
assign _7530_ = _7531_ | _7533_ /*34799*/;
assign _7345_ = _7525_ ^ _7532_ /*34802*/;
assign _7539_ = D[31] ^ Q[45] /*34798*/;
assign _7536_ = _6960_ & _7539_ /*34794*/;
assign _7537_ = _6960_ ^ _7539_ /*34797*/;
assign _7538_ = _7530_ & _7537_ /*34795*/;
assign _7535_ = _7536_ | _7538_ /*34793*/;
assign _7346_ = _7530_ ^ _7537_ /*34796*/;
assign _7544_ = D[32] ^ Q[45] /*34792*/;
assign _7541_ = _6961_ & _7544_ /*34788*/;
assign _7542_ = _6961_ ^ _7544_ /*34791*/;
assign _7543_ = _7535_ & _7542_ /*34789*/;
assign _7540_ = _7541_ | _7543_ /*34787*/;
assign _7347_ = _7535_ ^ _7542_ /*34790*/;
assign _7549_ = D[33] ^ Q[45] /*34786*/;
assign _7546_ = _6962_ & _7549_ /*34782*/;
assign _7547_ = _6962_ ^ _7549_ /*34785*/;
assign _7548_ = _7540_ & _7547_ /*34783*/;
assign _7545_ = _7546_ | _7548_ /*34781*/;
assign _7348_ = _7540_ ^ _7547_ /*34784*/;
assign _7554_ = D[34] ^ Q[45] /*34780*/;
assign _7551_ = _6963_ & _7554_ /*34776*/;
assign _7552_ = _6963_ ^ _7554_ /*34779*/;
assign _7553_ = _7545_ & _7552_ /*34777*/;
assign _7550_ = _7551_ | _7553_ /*34775*/;
assign _7349_ = _7545_ ^ _7552_ /*34778*/;
assign _7559_ = D[35] ^ Q[45] /*34774*/;
assign _7556_ = _6964_ & _7559_ /*34770*/;
assign _7557_ = _6964_ ^ _7559_ /*34773*/;
assign _7558_ = _7550_ & _7557_ /*34771*/;
assign _7555_ = _7556_ | _7558_ /*34769*/;
assign _7350_ = _7550_ ^ _7557_ /*34772*/;
assign _7564_ = D[36] ^ Q[45] /*34768*/;
assign _7561_ = _6965_ & _7564_ /*34764*/;
assign _7562_ = _6965_ ^ _7564_ /*34767*/;
assign _7563_ = _7555_ & _7562_ /*34765*/;
assign _7560_ = _7561_ | _7563_ /*34763*/;
assign _7351_ = _7555_ ^ _7562_ /*34766*/;
assign _7569_ = D[37] ^ Q[45] /*34762*/;
assign _7566_ = _6966_ & _7569_ /*34758*/;
assign _7567_ = _6966_ ^ _7569_ /*34761*/;
assign _7568_ = _7560_ & _7567_ /*34759*/;
assign _7565_ = _7566_ | _7568_ /*34757*/;
assign _7352_ = _7560_ ^ _7567_ /*34760*/;
assign _7574_ = D[38] ^ Q[45] /*34756*/;
assign _7571_ = _6967_ & _7574_ /*34752*/;
assign _7572_ = _6967_ ^ _7574_ /*34755*/;
assign _7573_ = _7565_ & _7572_ /*34753*/;
assign _7570_ = _7571_ | _7573_ /*34751*/;
assign _7353_ = _7565_ ^ _7572_ /*34754*/;
assign _7579_ = D[39] ^ Q[45] /*34750*/;
assign _7576_ = _6968_ & _7579_ /*34746*/;
assign _7577_ = _6968_ ^ _7579_ /*34749*/;
assign _7578_ = _7570_ & _7577_ /*34747*/;
assign _7575_ = _7576_ | _7578_ /*34745*/;
assign _7354_ = _7570_ ^ _7577_ /*34748*/;
assign _7584_ = D[40] ^ Q[45] /*34744*/;
assign _7581_ = _6969_ & _7584_ /*34740*/;
assign _7582_ = _6969_ ^ _7584_ /*34743*/;
assign _7583_ = _7575_ & _7582_ /*34741*/;
assign _7580_ = _7581_ | _7583_ /*34739*/;
assign _7355_ = _7575_ ^ _7582_ /*34742*/;
assign _7589_ = D[41] ^ Q[45] /*34738*/;
assign _7586_ = _6970_ & _7589_ /*34734*/;
assign _7587_ = _6970_ ^ _7589_ /*34737*/;
assign _7588_ = _7580_ & _7587_ /*34735*/;
assign _7585_ = _7586_ | _7588_ /*34733*/;
assign _7356_ = _7580_ ^ _7587_ /*34736*/;
assign _7594_ = D[42] ^ Q[45] /*34732*/;
assign _7591_ = _6971_ & _7594_ /*34728*/;
assign _7592_ = _6971_ ^ _7594_ /*34731*/;
assign _7593_ = _7585_ & _7592_ /*34729*/;
assign _7590_ = _7591_ | _7593_ /*34727*/;
assign _7357_ = _7585_ ^ _7592_ /*34730*/;
assign _7599_ = D[43] ^ Q[45] /*34726*/;
assign _7596_ = _6972_ & _7599_ /*34722*/;
assign _7597_ = _6972_ ^ _7599_ /*34725*/;
assign _7598_ = _7590_ & _7597_ /*34723*/;
assign _7595_ = _7596_ | _7598_ /*34721*/;
assign _7358_ = _7590_ ^ _7597_ /*34724*/;
assign _7604_ = D[44] ^ Q[45] /*34720*/;
assign _7601_ = _6973_ & _7604_ /*34716*/;
assign _7602_ = _6973_ ^ _7604_ /*34719*/;
assign _7603_ = _7595_ & _7602_ /*34717*/;
assign _7600_ = _7601_ | _7603_ /*34715*/;
assign _7359_ = _7595_ ^ _7602_ /*34718*/;
assign _7609_ = D[45] ^ Q[45] /*34714*/;
assign _7606_ = _6974_ & _7609_ /*34710*/;
assign _7607_ = _6974_ ^ _7609_ /*34713*/;
assign _7608_ = _7600_ & _7607_ /*34711*/;
assign _7605_ = _7606_ | _7608_ /*34709*/;
assign _7360_ = _7600_ ^ _7607_ /*34712*/;
assign _7614_ = D[46] ^ Q[45] /*34708*/;
assign _7611_ = _6975_ & _7614_ /*34704*/;
assign _7612_ = _6975_ ^ _7614_ /*34707*/;
assign _7613_ = _7605_ & _7612_ /*34705*/;
assign _7610_ = _7611_ | _7613_ /*34703*/;
assign _7361_ = _7605_ ^ _7612_ /*34706*/;
assign _7619_ = D[47] ^ Q[45] /*34702*/;
assign _7616_ = _6976_ & _7619_ /*34698*/;
assign _7617_ = _6976_ ^ _7619_ /*34701*/;
assign _7618_ = _7610_ & _7617_ /*34699*/;
assign _7615_ = _7616_ | _7618_ /*34697*/;
assign _7362_ = _7610_ ^ _7617_ /*34700*/;
assign _7624_ = D[48] ^ Q[45] /*34696*/;
assign _7621_ = _6977_ & _7624_ /*34692*/;
assign _7622_ = _6977_ ^ _7624_ /*34695*/;
assign _7623_ = _7615_ & _7622_ /*34693*/;
assign _7620_ = _7621_ | _7623_ /*34691*/;
assign _7363_ = _7615_ ^ _7622_ /*34694*/;
assign _7629_ = D[49] ^ Q[45] /*34690*/;
assign _7626_ = _6978_ & _7629_ /*34686*/;
assign _7627_ = _6978_ ^ _7629_ /*34689*/;
assign _7628_ = _7620_ & _7627_ /*34687*/;
assign _7625_ = _7626_ | _7628_ /*34685*/;
assign _7364_ = _7620_ ^ _7627_ /*34688*/;
assign _7634_ = D[50] ^ Q[45] /*34684*/;
assign _7631_ = _6979_ & _7634_ /*34680*/;
assign _7632_ = _6979_ ^ _7634_ /*34683*/;
assign _7633_ = _7625_ & _7632_ /*34681*/;
assign _7630_ = _7631_ | _7633_ /*34679*/;
assign _7365_ = _7625_ ^ _7632_ /*34682*/;
assign _7639_ = D[51] ^ Q[45] /*34678*/;
assign _7636_ = _6980_ & _7639_ /*34674*/;
assign _7637_ = _6980_ ^ _7639_ /*34677*/;
assign _7638_ = _7630_ & _7637_ /*34675*/;
assign _7635_ = _7636_ | _7638_ /*34673*/;
assign _7366_ = _7630_ ^ _7637_ /*34676*/;
assign _7644_ = D[52] ^ Q[45] /*34672*/;
assign _7641_ = _6981_ & _7644_ /*34668*/;
assign _7642_ = _6981_ ^ _7644_ /*34671*/;
assign _7643_ = _7635_ & _7642_ /*34669*/;
assign _7640_ = _7641_ | _7643_ /*34667*/;
assign _7367_ = _7635_ ^ _7642_ /*34670*/;
assign _7649_ = D[53] ^ Q[45] /*34666*/;
assign _7646_ = _6982_ & _7649_ /*34662*/;
assign _7647_ = _6982_ ^ _7649_ /*34665*/;
assign _7648_ = _7640_ & _7647_ /*34663*/;
assign _7645_ = _7646_ | _7648_ /*34661*/;
assign _7368_ = _7640_ ^ _7647_ /*34664*/;
assign _7654_ = D[54] ^ Q[45] /*34660*/;
assign _7651_ = _6983_ & _7654_ /*34656*/;
assign _7652_ = _6983_ ^ _7654_ /*34659*/;
assign _7653_ = _7645_ & _7652_ /*34657*/;
assign _7650_ = _7651_ | _7653_ /*34655*/;
assign _7369_ = _7645_ ^ _7652_ /*34658*/;
assign _7659_ = D[55] ^ Q[45] /*34654*/;
assign _7656_ = _6984_ & _7659_ /*34650*/;
assign _7657_ = _6984_ ^ _7659_ /*34653*/;
assign _7658_ = _7650_ & _7657_ /*34651*/;
assign _7655_ = _7656_ | _7658_ /*34649*/;
assign _7370_ = _7650_ ^ _7657_ /*34652*/;
assign _7664_ = D[56] ^ Q[45] /*34648*/;
assign _7661_ = _6985_ & _7664_ /*34644*/;
assign _7662_ = _6985_ ^ _7664_ /*34647*/;
assign _7663_ = _7655_ & _7662_ /*34645*/;
assign _7660_ = _7661_ | _7663_ /*34643*/;
assign _7371_ = _7655_ ^ _7662_ /*34646*/;
assign _7669_ = D[57] ^ Q[45] /*34642*/;
assign _7666_ = _6986_ & _7669_ /*34638*/;
assign _7667_ = _6986_ ^ _7669_ /*34641*/;
assign _7668_ = _7660_ & _7667_ /*34639*/;
assign _7665_ = _7666_ | _7668_ /*34637*/;
assign _7372_ = _7660_ ^ _7667_ /*34640*/;
assign _7674_ = D[58] ^ Q[45] /*34636*/;
assign _7671_ = _6987_ & _7674_ /*34632*/;
assign _7672_ = _6987_ ^ _7674_ /*34635*/;
assign _7673_ = _7665_ & _7672_ /*34633*/;
assign _7670_ = _7671_ | _7673_ /*34631*/;
assign _7373_ = _7665_ ^ _7672_ /*34634*/;
assign _7679_ = D[59] ^ Q[45] /*34630*/;
assign _7676_ = _6988_ & _7679_ /*34626*/;
assign _7677_ = _6988_ ^ _7679_ /*34629*/;
assign _7678_ = _7670_ & _7677_ /*34627*/;
assign _7675_ = _7676_ | _7678_ /*34625*/;
assign _7374_ = _7670_ ^ _7677_ /*34628*/;
assign _7684_ = D[60] ^ Q[45] /*34624*/;
assign _7681_ = _6989_ & _7684_ /*34620*/;
assign _7682_ = _6989_ ^ _7684_ /*34623*/;
assign _7683_ = _7675_ & _7682_ /*34621*/;
assign _7680_ = _7681_ | _7683_ /*34619*/;
assign _7375_ = _7675_ ^ _7682_ /*34622*/;
assign _7689_ = D[61] ^ Q[45] /*34618*/;
assign _7686_ = _6990_ & _7689_ /*34614*/;
assign _7687_ = _6990_ ^ _7689_ /*34617*/;
assign _7688_ = _7680_ & _7687_ /*34615*/;
assign _7685_ = _7686_ | _7688_ /*34613*/;
assign _7376_ = _7680_ ^ _7687_ /*34616*/;
assign _7694_ = D[62] ^ Q[45] /*34612*/;
assign _7691_ = _6991_ & _7694_ /*34608*/;
assign _7692_ = _6991_ ^ _7694_ /*34611*/;
assign _7693_ = _7685_ & _7692_ /*34609*/;
assign _7690_ = _7691_ | _7693_ /*34607*/;
assign _7377_ = _7685_ ^ _7692_ /*34610*/;
assign _7698_ = zeroWire ^ Q[45] /*34606*/;
assign _7695_ = _6992_ & _7698_ /*34602*/;
assign _7696_ = _6992_ ^ _7698_ /*34605*/;
assign _7697_ = _7690_ & _7696_ /*34603*/;
assign Q[44] = _7695_ | _7697_ /*34601*/;
assign _7378_ = _7690_ ^ _7696_ /*34604*/;
assign _7769_ = D[0] ^ Q[44] /*34215*/;
assign _7766_ = R_0[43] & _7769_ /*34211*/;
assign _7767_ = R_0[43] ^ _7769_ /*34214*/;
assign _7768_ = Q[44] & _7767_ /*34212*/;
assign _7765_ = _7766_ | _7768_ /*34210*/;
assign _7700_ = Q[44] ^ _7767_ /*34213*/;
assign _7774_ = D[1] ^ Q[44] /*34209*/;
assign _7771_ = _7315_ & _7774_ /*34205*/;
assign _7772_ = _7315_ ^ _7774_ /*34208*/;
assign _7773_ = _7765_ & _7772_ /*34206*/;
assign _7770_ = _7771_ | _7773_ /*34204*/;
assign _7701_ = _7765_ ^ _7772_ /*34207*/;
assign _7779_ = D[2] ^ Q[44] /*34203*/;
assign _7776_ = _7316_ & _7779_ /*34199*/;
assign _7777_ = _7316_ ^ _7779_ /*34202*/;
assign _7778_ = _7770_ & _7777_ /*34200*/;
assign _7775_ = _7776_ | _7778_ /*34198*/;
assign _7702_ = _7770_ ^ _7777_ /*34201*/;
assign _7784_ = D[3] ^ Q[44] /*34197*/;
assign _7781_ = _7317_ & _7784_ /*34193*/;
assign _7782_ = _7317_ ^ _7784_ /*34196*/;
assign _7783_ = _7775_ & _7782_ /*34194*/;
assign _7780_ = _7781_ | _7783_ /*34192*/;
assign _7703_ = _7775_ ^ _7782_ /*34195*/;
assign _7789_ = D[4] ^ Q[44] /*34191*/;
assign _7786_ = _7318_ & _7789_ /*34187*/;
assign _7787_ = _7318_ ^ _7789_ /*34190*/;
assign _7788_ = _7780_ & _7787_ /*34188*/;
assign _7785_ = _7786_ | _7788_ /*34186*/;
assign _7704_ = _7780_ ^ _7787_ /*34189*/;
assign _7794_ = D[5] ^ Q[44] /*34185*/;
assign _7791_ = _7319_ & _7794_ /*34181*/;
assign _7792_ = _7319_ ^ _7794_ /*34184*/;
assign _7793_ = _7785_ & _7792_ /*34182*/;
assign _7790_ = _7791_ | _7793_ /*34180*/;
assign _7705_ = _7785_ ^ _7792_ /*34183*/;
assign _7799_ = D[6] ^ Q[44] /*34179*/;
assign _7796_ = _7320_ & _7799_ /*34175*/;
assign _7797_ = _7320_ ^ _7799_ /*34178*/;
assign _7798_ = _7790_ & _7797_ /*34176*/;
assign _7795_ = _7796_ | _7798_ /*34174*/;
assign _7706_ = _7790_ ^ _7797_ /*34177*/;
assign _7804_ = D[7] ^ Q[44] /*34173*/;
assign _7801_ = _7321_ & _7804_ /*34169*/;
assign _7802_ = _7321_ ^ _7804_ /*34172*/;
assign _7803_ = _7795_ & _7802_ /*34170*/;
assign _7800_ = _7801_ | _7803_ /*34168*/;
assign _7707_ = _7795_ ^ _7802_ /*34171*/;
assign _7809_ = D[8] ^ Q[44] /*34167*/;
assign _7806_ = _7322_ & _7809_ /*34163*/;
assign _7807_ = _7322_ ^ _7809_ /*34166*/;
assign _7808_ = _7800_ & _7807_ /*34164*/;
assign _7805_ = _7806_ | _7808_ /*34162*/;
assign _7708_ = _7800_ ^ _7807_ /*34165*/;
assign _7814_ = D[9] ^ Q[44] /*34161*/;
assign _7811_ = _7323_ & _7814_ /*34157*/;
assign _7812_ = _7323_ ^ _7814_ /*34160*/;
assign _7813_ = _7805_ & _7812_ /*34158*/;
assign _7810_ = _7811_ | _7813_ /*34156*/;
assign _7709_ = _7805_ ^ _7812_ /*34159*/;
assign _7819_ = D[10] ^ Q[44] /*34155*/;
assign _7816_ = _7324_ & _7819_ /*34151*/;
assign _7817_ = _7324_ ^ _7819_ /*34154*/;
assign _7818_ = _7810_ & _7817_ /*34152*/;
assign _7815_ = _7816_ | _7818_ /*34150*/;
assign _7710_ = _7810_ ^ _7817_ /*34153*/;
assign _7824_ = D[11] ^ Q[44] /*34149*/;
assign _7821_ = _7325_ & _7824_ /*34145*/;
assign _7822_ = _7325_ ^ _7824_ /*34148*/;
assign _7823_ = _7815_ & _7822_ /*34146*/;
assign _7820_ = _7821_ | _7823_ /*34144*/;
assign _7711_ = _7815_ ^ _7822_ /*34147*/;
assign _7829_ = D[12] ^ Q[44] /*34143*/;
assign _7826_ = _7326_ & _7829_ /*34139*/;
assign _7827_ = _7326_ ^ _7829_ /*34142*/;
assign _7828_ = _7820_ & _7827_ /*34140*/;
assign _7825_ = _7826_ | _7828_ /*34138*/;
assign _7712_ = _7820_ ^ _7827_ /*34141*/;
assign _7834_ = D[13] ^ Q[44] /*34137*/;
assign _7831_ = _7327_ & _7834_ /*34133*/;
assign _7832_ = _7327_ ^ _7834_ /*34136*/;
assign _7833_ = _7825_ & _7832_ /*34134*/;
assign _7830_ = _7831_ | _7833_ /*34132*/;
assign _7713_ = _7825_ ^ _7832_ /*34135*/;
assign _7839_ = D[14] ^ Q[44] /*34131*/;
assign _7836_ = _7328_ & _7839_ /*34127*/;
assign _7837_ = _7328_ ^ _7839_ /*34130*/;
assign _7838_ = _7830_ & _7837_ /*34128*/;
assign _7835_ = _7836_ | _7838_ /*34126*/;
assign _7714_ = _7830_ ^ _7837_ /*34129*/;
assign _7844_ = D[15] ^ Q[44] /*34125*/;
assign _7841_ = _7329_ & _7844_ /*34121*/;
assign _7842_ = _7329_ ^ _7844_ /*34124*/;
assign _7843_ = _7835_ & _7842_ /*34122*/;
assign _7840_ = _7841_ | _7843_ /*34120*/;
assign _7715_ = _7835_ ^ _7842_ /*34123*/;
assign _7849_ = D[16] ^ Q[44] /*34119*/;
assign _7846_ = _7330_ & _7849_ /*34115*/;
assign _7847_ = _7330_ ^ _7849_ /*34118*/;
assign _7848_ = _7840_ & _7847_ /*34116*/;
assign _7845_ = _7846_ | _7848_ /*34114*/;
assign _7716_ = _7840_ ^ _7847_ /*34117*/;
assign _7854_ = D[17] ^ Q[44] /*34113*/;
assign _7851_ = _7331_ & _7854_ /*34109*/;
assign _7852_ = _7331_ ^ _7854_ /*34112*/;
assign _7853_ = _7845_ & _7852_ /*34110*/;
assign _7850_ = _7851_ | _7853_ /*34108*/;
assign _7717_ = _7845_ ^ _7852_ /*34111*/;
assign _7859_ = D[18] ^ Q[44] /*34107*/;
assign _7856_ = _7332_ & _7859_ /*34103*/;
assign _7857_ = _7332_ ^ _7859_ /*34106*/;
assign _7858_ = _7850_ & _7857_ /*34104*/;
assign _7855_ = _7856_ | _7858_ /*34102*/;
assign _7718_ = _7850_ ^ _7857_ /*34105*/;
assign _7864_ = D[19] ^ Q[44] /*34101*/;
assign _7861_ = _7333_ & _7864_ /*34097*/;
assign _7862_ = _7333_ ^ _7864_ /*34100*/;
assign _7863_ = _7855_ & _7862_ /*34098*/;
assign _7860_ = _7861_ | _7863_ /*34096*/;
assign _7719_ = _7855_ ^ _7862_ /*34099*/;
assign _7869_ = D[20] ^ Q[44] /*34095*/;
assign _7866_ = _7334_ & _7869_ /*34091*/;
assign _7867_ = _7334_ ^ _7869_ /*34094*/;
assign _7868_ = _7860_ & _7867_ /*34092*/;
assign _7865_ = _7866_ | _7868_ /*34090*/;
assign _7720_ = _7860_ ^ _7867_ /*34093*/;
assign _7874_ = D[21] ^ Q[44] /*34089*/;
assign _7871_ = _7335_ & _7874_ /*34085*/;
assign _7872_ = _7335_ ^ _7874_ /*34088*/;
assign _7873_ = _7865_ & _7872_ /*34086*/;
assign _7870_ = _7871_ | _7873_ /*34084*/;
assign _7721_ = _7865_ ^ _7872_ /*34087*/;
assign _7879_ = D[22] ^ Q[44] /*34083*/;
assign _7876_ = _7336_ & _7879_ /*34079*/;
assign _7877_ = _7336_ ^ _7879_ /*34082*/;
assign _7878_ = _7870_ & _7877_ /*34080*/;
assign _7875_ = _7876_ | _7878_ /*34078*/;
assign _7722_ = _7870_ ^ _7877_ /*34081*/;
assign _7884_ = D[23] ^ Q[44] /*34077*/;
assign _7881_ = _7337_ & _7884_ /*34073*/;
assign _7882_ = _7337_ ^ _7884_ /*34076*/;
assign _7883_ = _7875_ & _7882_ /*34074*/;
assign _7880_ = _7881_ | _7883_ /*34072*/;
assign _7723_ = _7875_ ^ _7882_ /*34075*/;
assign _7889_ = D[24] ^ Q[44] /*34071*/;
assign _7886_ = _7338_ & _7889_ /*34067*/;
assign _7887_ = _7338_ ^ _7889_ /*34070*/;
assign _7888_ = _7880_ & _7887_ /*34068*/;
assign _7885_ = _7886_ | _7888_ /*34066*/;
assign _7724_ = _7880_ ^ _7887_ /*34069*/;
assign _7894_ = D[25] ^ Q[44] /*34065*/;
assign _7891_ = _7339_ & _7894_ /*34061*/;
assign _7892_ = _7339_ ^ _7894_ /*34064*/;
assign _7893_ = _7885_ & _7892_ /*34062*/;
assign _7890_ = _7891_ | _7893_ /*34060*/;
assign _7725_ = _7885_ ^ _7892_ /*34063*/;
assign _7899_ = D[26] ^ Q[44] /*34059*/;
assign _7896_ = _7340_ & _7899_ /*34055*/;
assign _7897_ = _7340_ ^ _7899_ /*34058*/;
assign _7898_ = _7890_ & _7897_ /*34056*/;
assign _7895_ = _7896_ | _7898_ /*34054*/;
assign _7726_ = _7890_ ^ _7897_ /*34057*/;
assign _7904_ = D[27] ^ Q[44] /*34053*/;
assign _7901_ = _7341_ & _7904_ /*34049*/;
assign _7902_ = _7341_ ^ _7904_ /*34052*/;
assign _7903_ = _7895_ & _7902_ /*34050*/;
assign _7900_ = _7901_ | _7903_ /*34048*/;
assign _7727_ = _7895_ ^ _7902_ /*34051*/;
assign _7909_ = D[28] ^ Q[44] /*34047*/;
assign _7906_ = _7342_ & _7909_ /*34043*/;
assign _7907_ = _7342_ ^ _7909_ /*34046*/;
assign _7908_ = _7900_ & _7907_ /*34044*/;
assign _7905_ = _7906_ | _7908_ /*34042*/;
assign _7728_ = _7900_ ^ _7907_ /*34045*/;
assign _7914_ = D[29] ^ Q[44] /*34041*/;
assign _7911_ = _7343_ & _7914_ /*34037*/;
assign _7912_ = _7343_ ^ _7914_ /*34040*/;
assign _7913_ = _7905_ & _7912_ /*34038*/;
assign _7910_ = _7911_ | _7913_ /*34036*/;
assign _7729_ = _7905_ ^ _7912_ /*34039*/;
assign _7919_ = D[30] ^ Q[44] /*34035*/;
assign _7916_ = _7344_ & _7919_ /*34031*/;
assign _7917_ = _7344_ ^ _7919_ /*34034*/;
assign _7918_ = _7910_ & _7917_ /*34032*/;
assign _7915_ = _7916_ | _7918_ /*34030*/;
assign _7730_ = _7910_ ^ _7917_ /*34033*/;
assign _7924_ = D[31] ^ Q[44] /*34029*/;
assign _7921_ = _7345_ & _7924_ /*34025*/;
assign _7922_ = _7345_ ^ _7924_ /*34028*/;
assign _7923_ = _7915_ & _7922_ /*34026*/;
assign _7920_ = _7921_ | _7923_ /*34024*/;
assign _7731_ = _7915_ ^ _7922_ /*34027*/;
assign _7929_ = D[32] ^ Q[44] /*34023*/;
assign _7926_ = _7346_ & _7929_ /*34019*/;
assign _7927_ = _7346_ ^ _7929_ /*34022*/;
assign _7928_ = _7920_ & _7927_ /*34020*/;
assign _7925_ = _7926_ | _7928_ /*34018*/;
assign _7732_ = _7920_ ^ _7927_ /*34021*/;
assign _7934_ = D[33] ^ Q[44] /*34017*/;
assign _7931_ = _7347_ & _7934_ /*34013*/;
assign _7932_ = _7347_ ^ _7934_ /*34016*/;
assign _7933_ = _7925_ & _7932_ /*34014*/;
assign _7930_ = _7931_ | _7933_ /*34012*/;
assign _7733_ = _7925_ ^ _7932_ /*34015*/;
assign _7939_ = D[34] ^ Q[44] /*34011*/;
assign _7936_ = _7348_ & _7939_ /*34007*/;
assign _7937_ = _7348_ ^ _7939_ /*34010*/;
assign _7938_ = _7930_ & _7937_ /*34008*/;
assign _7935_ = _7936_ | _7938_ /*34006*/;
assign _7734_ = _7930_ ^ _7937_ /*34009*/;
assign _7944_ = D[35] ^ Q[44] /*34005*/;
assign _7941_ = _7349_ & _7944_ /*34001*/;
assign _7942_ = _7349_ ^ _7944_ /*34004*/;
assign _7943_ = _7935_ & _7942_ /*34002*/;
assign _7940_ = _7941_ | _7943_ /*34000*/;
assign _7735_ = _7935_ ^ _7942_ /*34003*/;
assign _7949_ = D[36] ^ Q[44] /*33999*/;
assign _7946_ = _7350_ & _7949_ /*33995*/;
assign _7947_ = _7350_ ^ _7949_ /*33998*/;
assign _7948_ = _7940_ & _7947_ /*33996*/;
assign _7945_ = _7946_ | _7948_ /*33994*/;
assign _7736_ = _7940_ ^ _7947_ /*33997*/;
assign _7954_ = D[37] ^ Q[44] /*33993*/;
assign _7951_ = _7351_ & _7954_ /*33989*/;
assign _7952_ = _7351_ ^ _7954_ /*33992*/;
assign _7953_ = _7945_ & _7952_ /*33990*/;
assign _7950_ = _7951_ | _7953_ /*33988*/;
assign _7737_ = _7945_ ^ _7952_ /*33991*/;
assign _7959_ = D[38] ^ Q[44] /*33987*/;
assign _7956_ = _7352_ & _7959_ /*33983*/;
assign _7957_ = _7352_ ^ _7959_ /*33986*/;
assign _7958_ = _7950_ & _7957_ /*33984*/;
assign _7955_ = _7956_ | _7958_ /*33982*/;
assign _7738_ = _7950_ ^ _7957_ /*33985*/;
assign _7964_ = D[39] ^ Q[44] /*33981*/;
assign _7961_ = _7353_ & _7964_ /*33977*/;
assign _7962_ = _7353_ ^ _7964_ /*33980*/;
assign _7963_ = _7955_ & _7962_ /*33978*/;
assign _7960_ = _7961_ | _7963_ /*33976*/;
assign _7739_ = _7955_ ^ _7962_ /*33979*/;
assign _7969_ = D[40] ^ Q[44] /*33975*/;
assign _7966_ = _7354_ & _7969_ /*33971*/;
assign _7967_ = _7354_ ^ _7969_ /*33974*/;
assign _7968_ = _7960_ & _7967_ /*33972*/;
assign _7965_ = _7966_ | _7968_ /*33970*/;
assign _7740_ = _7960_ ^ _7967_ /*33973*/;
assign _7974_ = D[41] ^ Q[44] /*33969*/;
assign _7971_ = _7355_ & _7974_ /*33965*/;
assign _7972_ = _7355_ ^ _7974_ /*33968*/;
assign _7973_ = _7965_ & _7972_ /*33966*/;
assign _7970_ = _7971_ | _7973_ /*33964*/;
assign _7741_ = _7965_ ^ _7972_ /*33967*/;
assign _7979_ = D[42] ^ Q[44] /*33963*/;
assign _7976_ = _7356_ & _7979_ /*33959*/;
assign _7977_ = _7356_ ^ _7979_ /*33962*/;
assign _7978_ = _7970_ & _7977_ /*33960*/;
assign _7975_ = _7976_ | _7978_ /*33958*/;
assign _7742_ = _7970_ ^ _7977_ /*33961*/;
assign _7984_ = D[43] ^ Q[44] /*33957*/;
assign _7981_ = _7357_ & _7984_ /*33953*/;
assign _7982_ = _7357_ ^ _7984_ /*33956*/;
assign _7983_ = _7975_ & _7982_ /*33954*/;
assign _7980_ = _7981_ | _7983_ /*33952*/;
assign _7743_ = _7975_ ^ _7982_ /*33955*/;
assign _7989_ = D[44] ^ Q[44] /*33951*/;
assign _7986_ = _7358_ & _7989_ /*33947*/;
assign _7987_ = _7358_ ^ _7989_ /*33950*/;
assign _7988_ = _7980_ & _7987_ /*33948*/;
assign _7985_ = _7986_ | _7988_ /*33946*/;
assign _7744_ = _7980_ ^ _7987_ /*33949*/;
assign _7994_ = D[45] ^ Q[44] /*33945*/;
assign _7991_ = _7359_ & _7994_ /*33941*/;
assign _7992_ = _7359_ ^ _7994_ /*33944*/;
assign _7993_ = _7985_ & _7992_ /*33942*/;
assign _7990_ = _7991_ | _7993_ /*33940*/;
assign _7745_ = _7985_ ^ _7992_ /*33943*/;
assign _7999_ = D[46] ^ Q[44] /*33939*/;
assign _7996_ = _7360_ & _7999_ /*33935*/;
assign _7997_ = _7360_ ^ _7999_ /*33938*/;
assign _7998_ = _7990_ & _7997_ /*33936*/;
assign _7995_ = _7996_ | _7998_ /*33934*/;
assign _7746_ = _7990_ ^ _7997_ /*33937*/;
assign _8004_ = D[47] ^ Q[44] /*33933*/;
assign _8001_ = _7361_ & _8004_ /*33929*/;
assign _8002_ = _7361_ ^ _8004_ /*33932*/;
assign _8003_ = _7995_ & _8002_ /*33930*/;
assign _8000_ = _8001_ | _8003_ /*33928*/;
assign _7747_ = _7995_ ^ _8002_ /*33931*/;
assign _8009_ = D[48] ^ Q[44] /*33927*/;
assign _8006_ = _7362_ & _8009_ /*33923*/;
assign _8007_ = _7362_ ^ _8009_ /*33926*/;
assign _8008_ = _8000_ & _8007_ /*33924*/;
assign _8005_ = _8006_ | _8008_ /*33922*/;
assign _7748_ = _8000_ ^ _8007_ /*33925*/;
assign _8014_ = D[49] ^ Q[44] /*33921*/;
assign _8011_ = _7363_ & _8014_ /*33917*/;
assign _8012_ = _7363_ ^ _8014_ /*33920*/;
assign _8013_ = _8005_ & _8012_ /*33918*/;
assign _8010_ = _8011_ | _8013_ /*33916*/;
assign _7749_ = _8005_ ^ _8012_ /*33919*/;
assign _8019_ = D[50] ^ Q[44] /*33915*/;
assign _8016_ = _7364_ & _8019_ /*33911*/;
assign _8017_ = _7364_ ^ _8019_ /*33914*/;
assign _8018_ = _8010_ & _8017_ /*33912*/;
assign _8015_ = _8016_ | _8018_ /*33910*/;
assign _7750_ = _8010_ ^ _8017_ /*33913*/;
assign _8024_ = D[51] ^ Q[44] /*33909*/;
assign _8021_ = _7365_ & _8024_ /*33905*/;
assign _8022_ = _7365_ ^ _8024_ /*33908*/;
assign _8023_ = _8015_ & _8022_ /*33906*/;
assign _8020_ = _8021_ | _8023_ /*33904*/;
assign _7751_ = _8015_ ^ _8022_ /*33907*/;
assign _8029_ = D[52] ^ Q[44] /*33903*/;
assign _8026_ = _7366_ & _8029_ /*33899*/;
assign _8027_ = _7366_ ^ _8029_ /*33902*/;
assign _8028_ = _8020_ & _8027_ /*33900*/;
assign _8025_ = _8026_ | _8028_ /*33898*/;
assign _7752_ = _8020_ ^ _8027_ /*33901*/;
assign _8034_ = D[53] ^ Q[44] /*33897*/;
assign _8031_ = _7367_ & _8034_ /*33893*/;
assign _8032_ = _7367_ ^ _8034_ /*33896*/;
assign _8033_ = _8025_ & _8032_ /*33894*/;
assign _8030_ = _8031_ | _8033_ /*33892*/;
assign _7753_ = _8025_ ^ _8032_ /*33895*/;
assign _8039_ = D[54] ^ Q[44] /*33891*/;
assign _8036_ = _7368_ & _8039_ /*33887*/;
assign _8037_ = _7368_ ^ _8039_ /*33890*/;
assign _8038_ = _8030_ & _8037_ /*33888*/;
assign _8035_ = _8036_ | _8038_ /*33886*/;
assign _7754_ = _8030_ ^ _8037_ /*33889*/;
assign _8044_ = D[55] ^ Q[44] /*33885*/;
assign _8041_ = _7369_ & _8044_ /*33881*/;
assign _8042_ = _7369_ ^ _8044_ /*33884*/;
assign _8043_ = _8035_ & _8042_ /*33882*/;
assign _8040_ = _8041_ | _8043_ /*33880*/;
assign _7755_ = _8035_ ^ _8042_ /*33883*/;
assign _8049_ = D[56] ^ Q[44] /*33879*/;
assign _8046_ = _7370_ & _8049_ /*33875*/;
assign _8047_ = _7370_ ^ _8049_ /*33878*/;
assign _8048_ = _8040_ & _8047_ /*33876*/;
assign _8045_ = _8046_ | _8048_ /*33874*/;
assign _7756_ = _8040_ ^ _8047_ /*33877*/;
assign _8054_ = D[57] ^ Q[44] /*33873*/;
assign _8051_ = _7371_ & _8054_ /*33869*/;
assign _8052_ = _7371_ ^ _8054_ /*33872*/;
assign _8053_ = _8045_ & _8052_ /*33870*/;
assign _8050_ = _8051_ | _8053_ /*33868*/;
assign _7757_ = _8045_ ^ _8052_ /*33871*/;
assign _8059_ = D[58] ^ Q[44] /*33867*/;
assign _8056_ = _7372_ & _8059_ /*33863*/;
assign _8057_ = _7372_ ^ _8059_ /*33866*/;
assign _8058_ = _8050_ & _8057_ /*33864*/;
assign _8055_ = _8056_ | _8058_ /*33862*/;
assign _7758_ = _8050_ ^ _8057_ /*33865*/;
assign _8064_ = D[59] ^ Q[44] /*33861*/;
assign _8061_ = _7373_ & _8064_ /*33857*/;
assign _8062_ = _7373_ ^ _8064_ /*33860*/;
assign _8063_ = _8055_ & _8062_ /*33858*/;
assign _8060_ = _8061_ | _8063_ /*33856*/;
assign _7759_ = _8055_ ^ _8062_ /*33859*/;
assign _8069_ = D[60] ^ Q[44] /*33855*/;
assign _8066_ = _7374_ & _8069_ /*33851*/;
assign _8067_ = _7374_ ^ _8069_ /*33854*/;
assign _8068_ = _8060_ & _8067_ /*33852*/;
assign _8065_ = _8066_ | _8068_ /*33850*/;
assign _7760_ = _8060_ ^ _8067_ /*33853*/;
assign _8074_ = D[61] ^ Q[44] /*33849*/;
assign _8071_ = _7375_ & _8074_ /*33845*/;
assign _8072_ = _7375_ ^ _8074_ /*33848*/;
assign _8073_ = _8065_ & _8072_ /*33846*/;
assign _8070_ = _8071_ | _8073_ /*33844*/;
assign _7761_ = _8065_ ^ _8072_ /*33847*/;
assign _8079_ = D[62] ^ Q[44] /*33843*/;
assign _8076_ = _7376_ & _8079_ /*33839*/;
assign _8077_ = _7376_ ^ _8079_ /*33842*/;
assign _8078_ = _8070_ & _8077_ /*33840*/;
assign _8075_ = _8076_ | _8078_ /*33838*/;
assign _7762_ = _8070_ ^ _8077_ /*33841*/;
assign _8083_ = zeroWire ^ Q[44] /*33837*/;
assign _8080_ = _7377_ & _8083_ /*33833*/;
assign _8081_ = _7377_ ^ _8083_ /*33836*/;
assign _8082_ = _8075_ & _8081_ /*33834*/;
assign Q[43] = _8080_ | _8082_ /*33832*/;
assign _7763_ = _8075_ ^ _8081_ /*33835*/;
assign _8154_ = D[0] ^ Q[43] /*33446*/;
assign _8151_ = R_0[42] & _8154_ /*33442*/;
assign _8152_ = R_0[42] ^ _8154_ /*33445*/;
assign _8153_ = Q[43] & _8152_ /*33443*/;
assign _8150_ = _8151_ | _8153_ /*33441*/;
assign _8085_ = Q[43] ^ _8152_ /*33444*/;
assign _8159_ = D[1] ^ Q[43] /*33440*/;
assign _8156_ = _7700_ & _8159_ /*33436*/;
assign _8157_ = _7700_ ^ _8159_ /*33439*/;
assign _8158_ = _8150_ & _8157_ /*33437*/;
assign _8155_ = _8156_ | _8158_ /*33435*/;
assign _8086_ = _8150_ ^ _8157_ /*33438*/;
assign _8164_ = D[2] ^ Q[43] /*33434*/;
assign _8161_ = _7701_ & _8164_ /*33430*/;
assign _8162_ = _7701_ ^ _8164_ /*33433*/;
assign _8163_ = _8155_ & _8162_ /*33431*/;
assign _8160_ = _8161_ | _8163_ /*33429*/;
assign _8087_ = _8155_ ^ _8162_ /*33432*/;
assign _8169_ = D[3] ^ Q[43] /*33428*/;
assign _8166_ = _7702_ & _8169_ /*33424*/;
assign _8167_ = _7702_ ^ _8169_ /*33427*/;
assign _8168_ = _8160_ & _8167_ /*33425*/;
assign _8165_ = _8166_ | _8168_ /*33423*/;
assign _8088_ = _8160_ ^ _8167_ /*33426*/;
assign _8174_ = D[4] ^ Q[43] /*33422*/;
assign _8171_ = _7703_ & _8174_ /*33418*/;
assign _8172_ = _7703_ ^ _8174_ /*33421*/;
assign _8173_ = _8165_ & _8172_ /*33419*/;
assign _8170_ = _8171_ | _8173_ /*33417*/;
assign _8089_ = _8165_ ^ _8172_ /*33420*/;
assign _8179_ = D[5] ^ Q[43] /*33416*/;
assign _8176_ = _7704_ & _8179_ /*33412*/;
assign _8177_ = _7704_ ^ _8179_ /*33415*/;
assign _8178_ = _8170_ & _8177_ /*33413*/;
assign _8175_ = _8176_ | _8178_ /*33411*/;
assign _8090_ = _8170_ ^ _8177_ /*33414*/;
assign _8184_ = D[6] ^ Q[43] /*33410*/;
assign _8181_ = _7705_ & _8184_ /*33406*/;
assign _8182_ = _7705_ ^ _8184_ /*33409*/;
assign _8183_ = _8175_ & _8182_ /*33407*/;
assign _8180_ = _8181_ | _8183_ /*33405*/;
assign _8091_ = _8175_ ^ _8182_ /*33408*/;
assign _8189_ = D[7] ^ Q[43] /*33404*/;
assign _8186_ = _7706_ & _8189_ /*33400*/;
assign _8187_ = _7706_ ^ _8189_ /*33403*/;
assign _8188_ = _8180_ & _8187_ /*33401*/;
assign _8185_ = _8186_ | _8188_ /*33399*/;
assign _8092_ = _8180_ ^ _8187_ /*33402*/;
assign _8194_ = D[8] ^ Q[43] /*33398*/;
assign _8191_ = _7707_ & _8194_ /*33394*/;
assign _8192_ = _7707_ ^ _8194_ /*33397*/;
assign _8193_ = _8185_ & _8192_ /*33395*/;
assign _8190_ = _8191_ | _8193_ /*33393*/;
assign _8093_ = _8185_ ^ _8192_ /*33396*/;
assign _8199_ = D[9] ^ Q[43] /*33392*/;
assign _8196_ = _7708_ & _8199_ /*33388*/;
assign _8197_ = _7708_ ^ _8199_ /*33391*/;
assign _8198_ = _8190_ & _8197_ /*33389*/;
assign _8195_ = _8196_ | _8198_ /*33387*/;
assign _8094_ = _8190_ ^ _8197_ /*33390*/;
assign _8204_ = D[10] ^ Q[43] /*33386*/;
assign _8201_ = _7709_ & _8204_ /*33382*/;
assign _8202_ = _7709_ ^ _8204_ /*33385*/;
assign _8203_ = _8195_ & _8202_ /*33383*/;
assign _8200_ = _8201_ | _8203_ /*33381*/;
assign _8095_ = _8195_ ^ _8202_ /*33384*/;
assign _8209_ = D[11] ^ Q[43] /*33380*/;
assign _8206_ = _7710_ & _8209_ /*33376*/;
assign _8207_ = _7710_ ^ _8209_ /*33379*/;
assign _8208_ = _8200_ & _8207_ /*33377*/;
assign _8205_ = _8206_ | _8208_ /*33375*/;
assign _8096_ = _8200_ ^ _8207_ /*33378*/;
assign _8214_ = D[12] ^ Q[43] /*33374*/;
assign _8211_ = _7711_ & _8214_ /*33370*/;
assign _8212_ = _7711_ ^ _8214_ /*33373*/;
assign _8213_ = _8205_ & _8212_ /*33371*/;
assign _8210_ = _8211_ | _8213_ /*33369*/;
assign _8097_ = _8205_ ^ _8212_ /*33372*/;
assign _8219_ = D[13] ^ Q[43] /*33368*/;
assign _8216_ = _7712_ & _8219_ /*33364*/;
assign _8217_ = _7712_ ^ _8219_ /*33367*/;
assign _8218_ = _8210_ & _8217_ /*33365*/;
assign _8215_ = _8216_ | _8218_ /*33363*/;
assign _8098_ = _8210_ ^ _8217_ /*33366*/;
assign _8224_ = D[14] ^ Q[43] /*33362*/;
assign _8221_ = _7713_ & _8224_ /*33358*/;
assign _8222_ = _7713_ ^ _8224_ /*33361*/;
assign _8223_ = _8215_ & _8222_ /*33359*/;
assign _8220_ = _8221_ | _8223_ /*33357*/;
assign _8099_ = _8215_ ^ _8222_ /*33360*/;
assign _8229_ = D[15] ^ Q[43] /*33356*/;
assign _8226_ = _7714_ & _8229_ /*33352*/;
assign _8227_ = _7714_ ^ _8229_ /*33355*/;
assign _8228_ = _8220_ & _8227_ /*33353*/;
assign _8225_ = _8226_ | _8228_ /*33351*/;
assign _8100_ = _8220_ ^ _8227_ /*33354*/;
assign _8234_ = D[16] ^ Q[43] /*33350*/;
assign _8231_ = _7715_ & _8234_ /*33346*/;
assign _8232_ = _7715_ ^ _8234_ /*33349*/;
assign _8233_ = _8225_ & _8232_ /*33347*/;
assign _8230_ = _8231_ | _8233_ /*33345*/;
assign _8101_ = _8225_ ^ _8232_ /*33348*/;
assign _8239_ = D[17] ^ Q[43] /*33344*/;
assign _8236_ = _7716_ & _8239_ /*33340*/;
assign _8237_ = _7716_ ^ _8239_ /*33343*/;
assign _8238_ = _8230_ & _8237_ /*33341*/;
assign _8235_ = _8236_ | _8238_ /*33339*/;
assign _8102_ = _8230_ ^ _8237_ /*33342*/;
assign _8244_ = D[18] ^ Q[43] /*33338*/;
assign _8241_ = _7717_ & _8244_ /*33334*/;
assign _8242_ = _7717_ ^ _8244_ /*33337*/;
assign _8243_ = _8235_ & _8242_ /*33335*/;
assign _8240_ = _8241_ | _8243_ /*33333*/;
assign _8103_ = _8235_ ^ _8242_ /*33336*/;
assign _8249_ = D[19] ^ Q[43] /*33332*/;
assign _8246_ = _7718_ & _8249_ /*33328*/;
assign _8247_ = _7718_ ^ _8249_ /*33331*/;
assign _8248_ = _8240_ & _8247_ /*33329*/;
assign _8245_ = _8246_ | _8248_ /*33327*/;
assign _8104_ = _8240_ ^ _8247_ /*33330*/;
assign _8254_ = D[20] ^ Q[43] /*33326*/;
assign _8251_ = _7719_ & _8254_ /*33322*/;
assign _8252_ = _7719_ ^ _8254_ /*33325*/;
assign _8253_ = _8245_ & _8252_ /*33323*/;
assign _8250_ = _8251_ | _8253_ /*33321*/;
assign _8105_ = _8245_ ^ _8252_ /*33324*/;
assign _8259_ = D[21] ^ Q[43] /*33320*/;
assign _8256_ = _7720_ & _8259_ /*33316*/;
assign _8257_ = _7720_ ^ _8259_ /*33319*/;
assign _8258_ = _8250_ & _8257_ /*33317*/;
assign _8255_ = _8256_ | _8258_ /*33315*/;
assign _8106_ = _8250_ ^ _8257_ /*33318*/;
assign _8264_ = D[22] ^ Q[43] /*33314*/;
assign _8261_ = _7721_ & _8264_ /*33310*/;
assign _8262_ = _7721_ ^ _8264_ /*33313*/;
assign _8263_ = _8255_ & _8262_ /*33311*/;
assign _8260_ = _8261_ | _8263_ /*33309*/;
assign _8107_ = _8255_ ^ _8262_ /*33312*/;
assign _8269_ = D[23] ^ Q[43] /*33308*/;
assign _8266_ = _7722_ & _8269_ /*33304*/;
assign _8267_ = _7722_ ^ _8269_ /*33307*/;
assign _8268_ = _8260_ & _8267_ /*33305*/;
assign _8265_ = _8266_ | _8268_ /*33303*/;
assign _8108_ = _8260_ ^ _8267_ /*33306*/;
assign _8274_ = D[24] ^ Q[43] /*33302*/;
assign _8271_ = _7723_ & _8274_ /*33298*/;
assign _8272_ = _7723_ ^ _8274_ /*33301*/;
assign _8273_ = _8265_ & _8272_ /*33299*/;
assign _8270_ = _8271_ | _8273_ /*33297*/;
assign _8109_ = _8265_ ^ _8272_ /*33300*/;
assign _8279_ = D[25] ^ Q[43] /*33296*/;
assign _8276_ = _7724_ & _8279_ /*33292*/;
assign _8277_ = _7724_ ^ _8279_ /*33295*/;
assign _8278_ = _8270_ & _8277_ /*33293*/;
assign _8275_ = _8276_ | _8278_ /*33291*/;
assign _8110_ = _8270_ ^ _8277_ /*33294*/;
assign _8284_ = D[26] ^ Q[43] /*33290*/;
assign _8281_ = _7725_ & _8284_ /*33286*/;
assign _8282_ = _7725_ ^ _8284_ /*33289*/;
assign _8283_ = _8275_ & _8282_ /*33287*/;
assign _8280_ = _8281_ | _8283_ /*33285*/;
assign _8111_ = _8275_ ^ _8282_ /*33288*/;
assign _8289_ = D[27] ^ Q[43] /*33284*/;
assign _8286_ = _7726_ & _8289_ /*33280*/;
assign _8287_ = _7726_ ^ _8289_ /*33283*/;
assign _8288_ = _8280_ & _8287_ /*33281*/;
assign _8285_ = _8286_ | _8288_ /*33279*/;
assign _8112_ = _8280_ ^ _8287_ /*33282*/;
assign _8294_ = D[28] ^ Q[43] /*33278*/;
assign _8291_ = _7727_ & _8294_ /*33274*/;
assign _8292_ = _7727_ ^ _8294_ /*33277*/;
assign _8293_ = _8285_ & _8292_ /*33275*/;
assign _8290_ = _8291_ | _8293_ /*33273*/;
assign _8113_ = _8285_ ^ _8292_ /*33276*/;
assign _8299_ = D[29] ^ Q[43] /*33272*/;
assign _8296_ = _7728_ & _8299_ /*33268*/;
assign _8297_ = _7728_ ^ _8299_ /*33271*/;
assign _8298_ = _8290_ & _8297_ /*33269*/;
assign _8295_ = _8296_ | _8298_ /*33267*/;
assign _8114_ = _8290_ ^ _8297_ /*33270*/;
assign _8304_ = D[30] ^ Q[43] /*33266*/;
assign _8301_ = _7729_ & _8304_ /*33262*/;
assign _8302_ = _7729_ ^ _8304_ /*33265*/;
assign _8303_ = _8295_ & _8302_ /*33263*/;
assign _8300_ = _8301_ | _8303_ /*33261*/;
assign _8115_ = _8295_ ^ _8302_ /*33264*/;
assign _8309_ = D[31] ^ Q[43] /*33260*/;
assign _8306_ = _7730_ & _8309_ /*33256*/;
assign _8307_ = _7730_ ^ _8309_ /*33259*/;
assign _8308_ = _8300_ & _8307_ /*33257*/;
assign _8305_ = _8306_ | _8308_ /*33255*/;
assign _8116_ = _8300_ ^ _8307_ /*33258*/;
assign _8314_ = D[32] ^ Q[43] /*33254*/;
assign _8311_ = _7731_ & _8314_ /*33250*/;
assign _8312_ = _7731_ ^ _8314_ /*33253*/;
assign _8313_ = _8305_ & _8312_ /*33251*/;
assign _8310_ = _8311_ | _8313_ /*33249*/;
assign _8117_ = _8305_ ^ _8312_ /*33252*/;
assign _8319_ = D[33] ^ Q[43] /*33248*/;
assign _8316_ = _7732_ & _8319_ /*33244*/;
assign _8317_ = _7732_ ^ _8319_ /*33247*/;
assign _8318_ = _8310_ & _8317_ /*33245*/;
assign _8315_ = _8316_ | _8318_ /*33243*/;
assign _8118_ = _8310_ ^ _8317_ /*33246*/;
assign _8324_ = D[34] ^ Q[43] /*33242*/;
assign _8321_ = _7733_ & _8324_ /*33238*/;
assign _8322_ = _7733_ ^ _8324_ /*33241*/;
assign _8323_ = _8315_ & _8322_ /*33239*/;
assign _8320_ = _8321_ | _8323_ /*33237*/;
assign _8119_ = _8315_ ^ _8322_ /*33240*/;
assign _8329_ = D[35] ^ Q[43] /*33236*/;
assign _8326_ = _7734_ & _8329_ /*33232*/;
assign _8327_ = _7734_ ^ _8329_ /*33235*/;
assign _8328_ = _8320_ & _8327_ /*33233*/;
assign _8325_ = _8326_ | _8328_ /*33231*/;
assign _8120_ = _8320_ ^ _8327_ /*33234*/;
assign _8334_ = D[36] ^ Q[43] /*33230*/;
assign _8331_ = _7735_ & _8334_ /*33226*/;
assign _8332_ = _7735_ ^ _8334_ /*33229*/;
assign _8333_ = _8325_ & _8332_ /*33227*/;
assign _8330_ = _8331_ | _8333_ /*33225*/;
assign _8121_ = _8325_ ^ _8332_ /*33228*/;
assign _8339_ = D[37] ^ Q[43] /*33224*/;
assign _8336_ = _7736_ & _8339_ /*33220*/;
assign _8337_ = _7736_ ^ _8339_ /*33223*/;
assign _8338_ = _8330_ & _8337_ /*33221*/;
assign _8335_ = _8336_ | _8338_ /*33219*/;
assign _8122_ = _8330_ ^ _8337_ /*33222*/;
assign _8344_ = D[38] ^ Q[43] /*33218*/;
assign _8341_ = _7737_ & _8344_ /*33214*/;
assign _8342_ = _7737_ ^ _8344_ /*33217*/;
assign _8343_ = _8335_ & _8342_ /*33215*/;
assign _8340_ = _8341_ | _8343_ /*33213*/;
assign _8123_ = _8335_ ^ _8342_ /*33216*/;
assign _8349_ = D[39] ^ Q[43] /*33212*/;
assign _8346_ = _7738_ & _8349_ /*33208*/;
assign _8347_ = _7738_ ^ _8349_ /*33211*/;
assign _8348_ = _8340_ & _8347_ /*33209*/;
assign _8345_ = _8346_ | _8348_ /*33207*/;
assign _8124_ = _8340_ ^ _8347_ /*33210*/;
assign _8354_ = D[40] ^ Q[43] /*33206*/;
assign _8351_ = _7739_ & _8354_ /*33202*/;
assign _8352_ = _7739_ ^ _8354_ /*33205*/;
assign _8353_ = _8345_ & _8352_ /*33203*/;
assign _8350_ = _8351_ | _8353_ /*33201*/;
assign _8125_ = _8345_ ^ _8352_ /*33204*/;
assign _8359_ = D[41] ^ Q[43] /*33200*/;
assign _8356_ = _7740_ & _8359_ /*33196*/;
assign _8357_ = _7740_ ^ _8359_ /*33199*/;
assign _8358_ = _8350_ & _8357_ /*33197*/;
assign _8355_ = _8356_ | _8358_ /*33195*/;
assign _8126_ = _8350_ ^ _8357_ /*33198*/;
assign _8364_ = D[42] ^ Q[43] /*33194*/;
assign _8361_ = _7741_ & _8364_ /*33190*/;
assign _8362_ = _7741_ ^ _8364_ /*33193*/;
assign _8363_ = _8355_ & _8362_ /*33191*/;
assign _8360_ = _8361_ | _8363_ /*33189*/;
assign _8127_ = _8355_ ^ _8362_ /*33192*/;
assign _8369_ = D[43] ^ Q[43] /*33188*/;
assign _8366_ = _7742_ & _8369_ /*33184*/;
assign _8367_ = _7742_ ^ _8369_ /*33187*/;
assign _8368_ = _8360_ & _8367_ /*33185*/;
assign _8365_ = _8366_ | _8368_ /*33183*/;
assign _8128_ = _8360_ ^ _8367_ /*33186*/;
assign _8374_ = D[44] ^ Q[43] /*33182*/;
assign _8371_ = _7743_ & _8374_ /*33178*/;
assign _8372_ = _7743_ ^ _8374_ /*33181*/;
assign _8373_ = _8365_ & _8372_ /*33179*/;
assign _8370_ = _8371_ | _8373_ /*33177*/;
assign _8129_ = _8365_ ^ _8372_ /*33180*/;
assign _8379_ = D[45] ^ Q[43] /*33176*/;
assign _8376_ = _7744_ & _8379_ /*33172*/;
assign _8377_ = _7744_ ^ _8379_ /*33175*/;
assign _8378_ = _8370_ & _8377_ /*33173*/;
assign _8375_ = _8376_ | _8378_ /*33171*/;
assign _8130_ = _8370_ ^ _8377_ /*33174*/;
assign _8384_ = D[46] ^ Q[43] /*33170*/;
assign _8381_ = _7745_ & _8384_ /*33166*/;
assign _8382_ = _7745_ ^ _8384_ /*33169*/;
assign _8383_ = _8375_ & _8382_ /*33167*/;
assign _8380_ = _8381_ | _8383_ /*33165*/;
assign _8131_ = _8375_ ^ _8382_ /*33168*/;
assign _8389_ = D[47] ^ Q[43] /*33164*/;
assign _8386_ = _7746_ & _8389_ /*33160*/;
assign _8387_ = _7746_ ^ _8389_ /*33163*/;
assign _8388_ = _8380_ & _8387_ /*33161*/;
assign _8385_ = _8386_ | _8388_ /*33159*/;
assign _8132_ = _8380_ ^ _8387_ /*33162*/;
assign _8394_ = D[48] ^ Q[43] /*33158*/;
assign _8391_ = _7747_ & _8394_ /*33154*/;
assign _8392_ = _7747_ ^ _8394_ /*33157*/;
assign _8393_ = _8385_ & _8392_ /*33155*/;
assign _8390_ = _8391_ | _8393_ /*33153*/;
assign _8133_ = _8385_ ^ _8392_ /*33156*/;
assign _8399_ = D[49] ^ Q[43] /*33152*/;
assign _8396_ = _7748_ & _8399_ /*33148*/;
assign _8397_ = _7748_ ^ _8399_ /*33151*/;
assign _8398_ = _8390_ & _8397_ /*33149*/;
assign _8395_ = _8396_ | _8398_ /*33147*/;
assign _8134_ = _8390_ ^ _8397_ /*33150*/;
assign _8404_ = D[50] ^ Q[43] /*33146*/;
assign _8401_ = _7749_ & _8404_ /*33142*/;
assign _8402_ = _7749_ ^ _8404_ /*33145*/;
assign _8403_ = _8395_ & _8402_ /*33143*/;
assign _8400_ = _8401_ | _8403_ /*33141*/;
assign _8135_ = _8395_ ^ _8402_ /*33144*/;
assign _8409_ = D[51] ^ Q[43] /*33140*/;
assign _8406_ = _7750_ & _8409_ /*33136*/;
assign _8407_ = _7750_ ^ _8409_ /*33139*/;
assign _8408_ = _8400_ & _8407_ /*33137*/;
assign _8405_ = _8406_ | _8408_ /*33135*/;
assign _8136_ = _8400_ ^ _8407_ /*33138*/;
assign _8414_ = D[52] ^ Q[43] /*33134*/;
assign _8411_ = _7751_ & _8414_ /*33130*/;
assign _8412_ = _7751_ ^ _8414_ /*33133*/;
assign _8413_ = _8405_ & _8412_ /*33131*/;
assign _8410_ = _8411_ | _8413_ /*33129*/;
assign _8137_ = _8405_ ^ _8412_ /*33132*/;
assign _8419_ = D[53] ^ Q[43] /*33128*/;
assign _8416_ = _7752_ & _8419_ /*33124*/;
assign _8417_ = _7752_ ^ _8419_ /*33127*/;
assign _8418_ = _8410_ & _8417_ /*33125*/;
assign _8415_ = _8416_ | _8418_ /*33123*/;
assign _8138_ = _8410_ ^ _8417_ /*33126*/;
assign _8424_ = D[54] ^ Q[43] /*33122*/;
assign _8421_ = _7753_ & _8424_ /*33118*/;
assign _8422_ = _7753_ ^ _8424_ /*33121*/;
assign _8423_ = _8415_ & _8422_ /*33119*/;
assign _8420_ = _8421_ | _8423_ /*33117*/;
assign _8139_ = _8415_ ^ _8422_ /*33120*/;
assign _8429_ = D[55] ^ Q[43] /*33116*/;
assign _8426_ = _7754_ & _8429_ /*33112*/;
assign _8427_ = _7754_ ^ _8429_ /*33115*/;
assign _8428_ = _8420_ & _8427_ /*33113*/;
assign _8425_ = _8426_ | _8428_ /*33111*/;
assign _8140_ = _8420_ ^ _8427_ /*33114*/;
assign _8434_ = D[56] ^ Q[43] /*33110*/;
assign _8431_ = _7755_ & _8434_ /*33106*/;
assign _8432_ = _7755_ ^ _8434_ /*33109*/;
assign _8433_ = _8425_ & _8432_ /*33107*/;
assign _8430_ = _8431_ | _8433_ /*33105*/;
assign _8141_ = _8425_ ^ _8432_ /*33108*/;
assign _8439_ = D[57] ^ Q[43] /*33104*/;
assign _8436_ = _7756_ & _8439_ /*33100*/;
assign _8437_ = _7756_ ^ _8439_ /*33103*/;
assign _8438_ = _8430_ & _8437_ /*33101*/;
assign _8435_ = _8436_ | _8438_ /*33099*/;
assign _8142_ = _8430_ ^ _8437_ /*33102*/;
assign _8444_ = D[58] ^ Q[43] /*33098*/;
assign _8441_ = _7757_ & _8444_ /*33094*/;
assign _8442_ = _7757_ ^ _8444_ /*33097*/;
assign _8443_ = _8435_ & _8442_ /*33095*/;
assign _8440_ = _8441_ | _8443_ /*33093*/;
assign _8143_ = _8435_ ^ _8442_ /*33096*/;
assign _8449_ = D[59] ^ Q[43] /*33092*/;
assign _8446_ = _7758_ & _8449_ /*33088*/;
assign _8447_ = _7758_ ^ _8449_ /*33091*/;
assign _8448_ = _8440_ & _8447_ /*33089*/;
assign _8445_ = _8446_ | _8448_ /*33087*/;
assign _8144_ = _8440_ ^ _8447_ /*33090*/;
assign _8454_ = D[60] ^ Q[43] /*33086*/;
assign _8451_ = _7759_ & _8454_ /*33082*/;
assign _8452_ = _7759_ ^ _8454_ /*33085*/;
assign _8453_ = _8445_ & _8452_ /*33083*/;
assign _8450_ = _8451_ | _8453_ /*33081*/;
assign _8145_ = _8445_ ^ _8452_ /*33084*/;
assign _8459_ = D[61] ^ Q[43] /*33080*/;
assign _8456_ = _7760_ & _8459_ /*33076*/;
assign _8457_ = _7760_ ^ _8459_ /*33079*/;
assign _8458_ = _8450_ & _8457_ /*33077*/;
assign _8455_ = _8456_ | _8458_ /*33075*/;
assign _8146_ = _8450_ ^ _8457_ /*33078*/;
assign _8464_ = D[62] ^ Q[43] /*33074*/;
assign _8461_ = _7761_ & _8464_ /*33070*/;
assign _8462_ = _7761_ ^ _8464_ /*33073*/;
assign _8463_ = _8455_ & _8462_ /*33071*/;
assign _8460_ = _8461_ | _8463_ /*33069*/;
assign _8147_ = _8455_ ^ _8462_ /*33072*/;
assign _8468_ = zeroWire ^ Q[43] /*33068*/;
assign _8465_ = _7762_ & _8468_ /*33064*/;
assign _8466_ = _7762_ ^ _8468_ /*33067*/;
assign _8467_ = _8460_ & _8466_ /*33065*/;
assign Q[42] = _8465_ | _8467_ /*33063*/;
assign _8148_ = _8460_ ^ _8466_ /*33066*/;
assign _8539_ = D[0] ^ Q[42] /*32677*/;
assign _8536_ = R_0[41] & _8539_ /*32673*/;
assign _8537_ = R_0[41] ^ _8539_ /*32676*/;
assign _8538_ = Q[42] & _8537_ /*32674*/;
assign _8535_ = _8536_ | _8538_ /*32672*/;
assign _8470_ = Q[42] ^ _8537_ /*32675*/;
assign _8544_ = D[1] ^ Q[42] /*32671*/;
assign _8541_ = _8085_ & _8544_ /*32667*/;
assign _8542_ = _8085_ ^ _8544_ /*32670*/;
assign _8543_ = _8535_ & _8542_ /*32668*/;
assign _8540_ = _8541_ | _8543_ /*32666*/;
assign _8471_ = _8535_ ^ _8542_ /*32669*/;
assign _8549_ = D[2] ^ Q[42] /*32665*/;
assign _8546_ = _8086_ & _8549_ /*32661*/;
assign _8547_ = _8086_ ^ _8549_ /*32664*/;
assign _8548_ = _8540_ & _8547_ /*32662*/;
assign _8545_ = _8546_ | _8548_ /*32660*/;
assign _8472_ = _8540_ ^ _8547_ /*32663*/;
assign _8554_ = D[3] ^ Q[42] /*32659*/;
assign _8551_ = _8087_ & _8554_ /*32655*/;
assign _8552_ = _8087_ ^ _8554_ /*32658*/;
assign _8553_ = _8545_ & _8552_ /*32656*/;
assign _8550_ = _8551_ | _8553_ /*32654*/;
assign _8473_ = _8545_ ^ _8552_ /*32657*/;
assign _8559_ = D[4] ^ Q[42] /*32653*/;
assign _8556_ = _8088_ & _8559_ /*32649*/;
assign _8557_ = _8088_ ^ _8559_ /*32652*/;
assign _8558_ = _8550_ & _8557_ /*32650*/;
assign _8555_ = _8556_ | _8558_ /*32648*/;
assign _8474_ = _8550_ ^ _8557_ /*32651*/;
assign _8564_ = D[5] ^ Q[42] /*32647*/;
assign _8561_ = _8089_ & _8564_ /*32643*/;
assign _8562_ = _8089_ ^ _8564_ /*32646*/;
assign _8563_ = _8555_ & _8562_ /*32644*/;
assign _8560_ = _8561_ | _8563_ /*32642*/;
assign _8475_ = _8555_ ^ _8562_ /*32645*/;
assign _8569_ = D[6] ^ Q[42] /*32641*/;
assign _8566_ = _8090_ & _8569_ /*32637*/;
assign _8567_ = _8090_ ^ _8569_ /*32640*/;
assign _8568_ = _8560_ & _8567_ /*32638*/;
assign _8565_ = _8566_ | _8568_ /*32636*/;
assign _8476_ = _8560_ ^ _8567_ /*32639*/;
assign _8574_ = D[7] ^ Q[42] /*32635*/;
assign _8571_ = _8091_ & _8574_ /*32631*/;
assign _8572_ = _8091_ ^ _8574_ /*32634*/;
assign _8573_ = _8565_ & _8572_ /*32632*/;
assign _8570_ = _8571_ | _8573_ /*32630*/;
assign _8477_ = _8565_ ^ _8572_ /*32633*/;
assign _8579_ = D[8] ^ Q[42] /*32629*/;
assign _8576_ = _8092_ & _8579_ /*32625*/;
assign _8577_ = _8092_ ^ _8579_ /*32628*/;
assign _8578_ = _8570_ & _8577_ /*32626*/;
assign _8575_ = _8576_ | _8578_ /*32624*/;
assign _8478_ = _8570_ ^ _8577_ /*32627*/;
assign _8584_ = D[9] ^ Q[42] /*32623*/;
assign _8581_ = _8093_ & _8584_ /*32619*/;
assign _8582_ = _8093_ ^ _8584_ /*32622*/;
assign _8583_ = _8575_ & _8582_ /*32620*/;
assign _8580_ = _8581_ | _8583_ /*32618*/;
assign _8479_ = _8575_ ^ _8582_ /*32621*/;
assign _8589_ = D[10] ^ Q[42] /*32617*/;
assign _8586_ = _8094_ & _8589_ /*32613*/;
assign _8587_ = _8094_ ^ _8589_ /*32616*/;
assign _8588_ = _8580_ & _8587_ /*32614*/;
assign _8585_ = _8586_ | _8588_ /*32612*/;
assign _8480_ = _8580_ ^ _8587_ /*32615*/;
assign _8594_ = D[11] ^ Q[42] /*32611*/;
assign _8591_ = _8095_ & _8594_ /*32607*/;
assign _8592_ = _8095_ ^ _8594_ /*32610*/;
assign _8593_ = _8585_ & _8592_ /*32608*/;
assign _8590_ = _8591_ | _8593_ /*32606*/;
assign _8481_ = _8585_ ^ _8592_ /*32609*/;
assign _8599_ = D[12] ^ Q[42] /*32605*/;
assign _8596_ = _8096_ & _8599_ /*32601*/;
assign _8597_ = _8096_ ^ _8599_ /*32604*/;
assign _8598_ = _8590_ & _8597_ /*32602*/;
assign _8595_ = _8596_ | _8598_ /*32600*/;
assign _8482_ = _8590_ ^ _8597_ /*32603*/;
assign _8604_ = D[13] ^ Q[42] /*32599*/;
assign _8601_ = _8097_ & _8604_ /*32595*/;
assign _8602_ = _8097_ ^ _8604_ /*32598*/;
assign _8603_ = _8595_ & _8602_ /*32596*/;
assign _8600_ = _8601_ | _8603_ /*32594*/;
assign _8483_ = _8595_ ^ _8602_ /*32597*/;
assign _8609_ = D[14] ^ Q[42] /*32593*/;
assign _8606_ = _8098_ & _8609_ /*32589*/;
assign _8607_ = _8098_ ^ _8609_ /*32592*/;
assign _8608_ = _8600_ & _8607_ /*32590*/;
assign _8605_ = _8606_ | _8608_ /*32588*/;
assign _8484_ = _8600_ ^ _8607_ /*32591*/;
assign _8614_ = D[15] ^ Q[42] /*32587*/;
assign _8611_ = _8099_ & _8614_ /*32583*/;
assign _8612_ = _8099_ ^ _8614_ /*32586*/;
assign _8613_ = _8605_ & _8612_ /*32584*/;
assign _8610_ = _8611_ | _8613_ /*32582*/;
assign _8485_ = _8605_ ^ _8612_ /*32585*/;
assign _8619_ = D[16] ^ Q[42] /*32581*/;
assign _8616_ = _8100_ & _8619_ /*32577*/;
assign _8617_ = _8100_ ^ _8619_ /*32580*/;
assign _8618_ = _8610_ & _8617_ /*32578*/;
assign _8615_ = _8616_ | _8618_ /*32576*/;
assign _8486_ = _8610_ ^ _8617_ /*32579*/;
assign _8624_ = D[17] ^ Q[42] /*32575*/;
assign _8621_ = _8101_ & _8624_ /*32571*/;
assign _8622_ = _8101_ ^ _8624_ /*32574*/;
assign _8623_ = _8615_ & _8622_ /*32572*/;
assign _8620_ = _8621_ | _8623_ /*32570*/;
assign _8487_ = _8615_ ^ _8622_ /*32573*/;
assign _8629_ = D[18] ^ Q[42] /*32569*/;
assign _8626_ = _8102_ & _8629_ /*32565*/;
assign _8627_ = _8102_ ^ _8629_ /*32568*/;
assign _8628_ = _8620_ & _8627_ /*32566*/;
assign _8625_ = _8626_ | _8628_ /*32564*/;
assign _8488_ = _8620_ ^ _8627_ /*32567*/;
assign _8634_ = D[19] ^ Q[42] /*32563*/;
assign _8631_ = _8103_ & _8634_ /*32559*/;
assign _8632_ = _8103_ ^ _8634_ /*32562*/;
assign _8633_ = _8625_ & _8632_ /*32560*/;
assign _8630_ = _8631_ | _8633_ /*32558*/;
assign _8489_ = _8625_ ^ _8632_ /*32561*/;
assign _8639_ = D[20] ^ Q[42] /*32557*/;
assign _8636_ = _8104_ & _8639_ /*32553*/;
assign _8637_ = _8104_ ^ _8639_ /*32556*/;
assign _8638_ = _8630_ & _8637_ /*32554*/;
assign _8635_ = _8636_ | _8638_ /*32552*/;
assign _8490_ = _8630_ ^ _8637_ /*32555*/;
assign _8644_ = D[21] ^ Q[42] /*32551*/;
assign _8641_ = _8105_ & _8644_ /*32547*/;
assign _8642_ = _8105_ ^ _8644_ /*32550*/;
assign _8643_ = _8635_ & _8642_ /*32548*/;
assign _8640_ = _8641_ | _8643_ /*32546*/;
assign _8491_ = _8635_ ^ _8642_ /*32549*/;
assign _8649_ = D[22] ^ Q[42] /*32545*/;
assign _8646_ = _8106_ & _8649_ /*32541*/;
assign _8647_ = _8106_ ^ _8649_ /*32544*/;
assign _8648_ = _8640_ & _8647_ /*32542*/;
assign _8645_ = _8646_ | _8648_ /*32540*/;
assign _8492_ = _8640_ ^ _8647_ /*32543*/;
assign _8654_ = D[23] ^ Q[42] /*32539*/;
assign _8651_ = _8107_ & _8654_ /*32535*/;
assign _8652_ = _8107_ ^ _8654_ /*32538*/;
assign _8653_ = _8645_ & _8652_ /*32536*/;
assign _8650_ = _8651_ | _8653_ /*32534*/;
assign _8493_ = _8645_ ^ _8652_ /*32537*/;
assign _8659_ = D[24] ^ Q[42] /*32533*/;
assign _8656_ = _8108_ & _8659_ /*32529*/;
assign _8657_ = _8108_ ^ _8659_ /*32532*/;
assign _8658_ = _8650_ & _8657_ /*32530*/;
assign _8655_ = _8656_ | _8658_ /*32528*/;
assign _8494_ = _8650_ ^ _8657_ /*32531*/;
assign _8664_ = D[25] ^ Q[42] /*32527*/;
assign _8661_ = _8109_ & _8664_ /*32523*/;
assign _8662_ = _8109_ ^ _8664_ /*32526*/;
assign _8663_ = _8655_ & _8662_ /*32524*/;
assign _8660_ = _8661_ | _8663_ /*32522*/;
assign _8495_ = _8655_ ^ _8662_ /*32525*/;
assign _8669_ = D[26] ^ Q[42] /*32521*/;
assign _8666_ = _8110_ & _8669_ /*32517*/;
assign _8667_ = _8110_ ^ _8669_ /*32520*/;
assign _8668_ = _8660_ & _8667_ /*32518*/;
assign _8665_ = _8666_ | _8668_ /*32516*/;
assign _8496_ = _8660_ ^ _8667_ /*32519*/;
assign _8674_ = D[27] ^ Q[42] /*32515*/;
assign _8671_ = _8111_ & _8674_ /*32511*/;
assign _8672_ = _8111_ ^ _8674_ /*32514*/;
assign _8673_ = _8665_ & _8672_ /*32512*/;
assign _8670_ = _8671_ | _8673_ /*32510*/;
assign _8497_ = _8665_ ^ _8672_ /*32513*/;
assign _8679_ = D[28] ^ Q[42] /*32509*/;
assign _8676_ = _8112_ & _8679_ /*32505*/;
assign _8677_ = _8112_ ^ _8679_ /*32508*/;
assign _8678_ = _8670_ & _8677_ /*32506*/;
assign _8675_ = _8676_ | _8678_ /*32504*/;
assign _8498_ = _8670_ ^ _8677_ /*32507*/;
assign _8684_ = D[29] ^ Q[42] /*32503*/;
assign _8681_ = _8113_ & _8684_ /*32499*/;
assign _8682_ = _8113_ ^ _8684_ /*32502*/;
assign _8683_ = _8675_ & _8682_ /*32500*/;
assign _8680_ = _8681_ | _8683_ /*32498*/;
assign _8499_ = _8675_ ^ _8682_ /*32501*/;
assign _8689_ = D[30] ^ Q[42] /*32497*/;
assign _8686_ = _8114_ & _8689_ /*32493*/;
assign _8687_ = _8114_ ^ _8689_ /*32496*/;
assign _8688_ = _8680_ & _8687_ /*32494*/;
assign _8685_ = _8686_ | _8688_ /*32492*/;
assign _8500_ = _8680_ ^ _8687_ /*32495*/;
assign _8694_ = D[31] ^ Q[42] /*32491*/;
assign _8691_ = _8115_ & _8694_ /*32487*/;
assign _8692_ = _8115_ ^ _8694_ /*32490*/;
assign _8693_ = _8685_ & _8692_ /*32488*/;
assign _8690_ = _8691_ | _8693_ /*32486*/;
assign _8501_ = _8685_ ^ _8692_ /*32489*/;
assign _8699_ = D[32] ^ Q[42] /*32485*/;
assign _8696_ = _8116_ & _8699_ /*32481*/;
assign _8697_ = _8116_ ^ _8699_ /*32484*/;
assign _8698_ = _8690_ & _8697_ /*32482*/;
assign _8695_ = _8696_ | _8698_ /*32480*/;
assign _8502_ = _8690_ ^ _8697_ /*32483*/;
assign _8704_ = D[33] ^ Q[42] /*32479*/;
assign _8701_ = _8117_ & _8704_ /*32475*/;
assign _8702_ = _8117_ ^ _8704_ /*32478*/;
assign _8703_ = _8695_ & _8702_ /*32476*/;
assign _8700_ = _8701_ | _8703_ /*32474*/;
assign _8503_ = _8695_ ^ _8702_ /*32477*/;
assign _8709_ = D[34] ^ Q[42] /*32473*/;
assign _8706_ = _8118_ & _8709_ /*32469*/;
assign _8707_ = _8118_ ^ _8709_ /*32472*/;
assign _8708_ = _8700_ & _8707_ /*32470*/;
assign _8705_ = _8706_ | _8708_ /*32468*/;
assign _8504_ = _8700_ ^ _8707_ /*32471*/;
assign _8714_ = D[35] ^ Q[42] /*32467*/;
assign _8711_ = _8119_ & _8714_ /*32463*/;
assign _8712_ = _8119_ ^ _8714_ /*32466*/;
assign _8713_ = _8705_ & _8712_ /*32464*/;
assign _8710_ = _8711_ | _8713_ /*32462*/;
assign _8505_ = _8705_ ^ _8712_ /*32465*/;
assign _8719_ = D[36] ^ Q[42] /*32461*/;
assign _8716_ = _8120_ & _8719_ /*32457*/;
assign _8717_ = _8120_ ^ _8719_ /*32460*/;
assign _8718_ = _8710_ & _8717_ /*32458*/;
assign _8715_ = _8716_ | _8718_ /*32456*/;
assign _8506_ = _8710_ ^ _8717_ /*32459*/;
assign _8724_ = D[37] ^ Q[42] /*32455*/;
assign _8721_ = _8121_ & _8724_ /*32451*/;
assign _8722_ = _8121_ ^ _8724_ /*32454*/;
assign _8723_ = _8715_ & _8722_ /*32452*/;
assign _8720_ = _8721_ | _8723_ /*32450*/;
assign _8507_ = _8715_ ^ _8722_ /*32453*/;
assign _8729_ = D[38] ^ Q[42] /*32449*/;
assign _8726_ = _8122_ & _8729_ /*32445*/;
assign _8727_ = _8122_ ^ _8729_ /*32448*/;
assign _8728_ = _8720_ & _8727_ /*32446*/;
assign _8725_ = _8726_ | _8728_ /*32444*/;
assign _8508_ = _8720_ ^ _8727_ /*32447*/;
assign _8734_ = D[39] ^ Q[42] /*32443*/;
assign _8731_ = _8123_ & _8734_ /*32439*/;
assign _8732_ = _8123_ ^ _8734_ /*32442*/;
assign _8733_ = _8725_ & _8732_ /*32440*/;
assign _8730_ = _8731_ | _8733_ /*32438*/;
assign _8509_ = _8725_ ^ _8732_ /*32441*/;
assign _8739_ = D[40] ^ Q[42] /*32437*/;
assign _8736_ = _8124_ & _8739_ /*32433*/;
assign _8737_ = _8124_ ^ _8739_ /*32436*/;
assign _8738_ = _8730_ & _8737_ /*32434*/;
assign _8735_ = _8736_ | _8738_ /*32432*/;
assign _8510_ = _8730_ ^ _8737_ /*32435*/;
assign _8744_ = D[41] ^ Q[42] /*32431*/;
assign _8741_ = _8125_ & _8744_ /*32427*/;
assign _8742_ = _8125_ ^ _8744_ /*32430*/;
assign _8743_ = _8735_ & _8742_ /*32428*/;
assign _8740_ = _8741_ | _8743_ /*32426*/;
assign _8511_ = _8735_ ^ _8742_ /*32429*/;
assign _8749_ = D[42] ^ Q[42] /*32425*/;
assign _8746_ = _8126_ & _8749_ /*32421*/;
assign _8747_ = _8126_ ^ _8749_ /*32424*/;
assign _8748_ = _8740_ & _8747_ /*32422*/;
assign _8745_ = _8746_ | _8748_ /*32420*/;
assign _8512_ = _8740_ ^ _8747_ /*32423*/;
assign _8754_ = D[43] ^ Q[42] /*32419*/;
assign _8751_ = _8127_ & _8754_ /*32415*/;
assign _8752_ = _8127_ ^ _8754_ /*32418*/;
assign _8753_ = _8745_ & _8752_ /*32416*/;
assign _8750_ = _8751_ | _8753_ /*32414*/;
assign _8513_ = _8745_ ^ _8752_ /*32417*/;
assign _8759_ = D[44] ^ Q[42] /*32413*/;
assign _8756_ = _8128_ & _8759_ /*32409*/;
assign _8757_ = _8128_ ^ _8759_ /*32412*/;
assign _8758_ = _8750_ & _8757_ /*32410*/;
assign _8755_ = _8756_ | _8758_ /*32408*/;
assign _8514_ = _8750_ ^ _8757_ /*32411*/;
assign _8764_ = D[45] ^ Q[42] /*32407*/;
assign _8761_ = _8129_ & _8764_ /*32403*/;
assign _8762_ = _8129_ ^ _8764_ /*32406*/;
assign _8763_ = _8755_ & _8762_ /*32404*/;
assign _8760_ = _8761_ | _8763_ /*32402*/;
assign _8515_ = _8755_ ^ _8762_ /*32405*/;
assign _8769_ = D[46] ^ Q[42] /*32401*/;
assign _8766_ = _8130_ & _8769_ /*32397*/;
assign _8767_ = _8130_ ^ _8769_ /*32400*/;
assign _8768_ = _8760_ & _8767_ /*32398*/;
assign _8765_ = _8766_ | _8768_ /*32396*/;
assign _8516_ = _8760_ ^ _8767_ /*32399*/;
assign _8774_ = D[47] ^ Q[42] /*32395*/;
assign _8771_ = _8131_ & _8774_ /*32391*/;
assign _8772_ = _8131_ ^ _8774_ /*32394*/;
assign _8773_ = _8765_ & _8772_ /*32392*/;
assign _8770_ = _8771_ | _8773_ /*32390*/;
assign _8517_ = _8765_ ^ _8772_ /*32393*/;
assign _8779_ = D[48] ^ Q[42] /*32389*/;
assign _8776_ = _8132_ & _8779_ /*32385*/;
assign _8777_ = _8132_ ^ _8779_ /*32388*/;
assign _8778_ = _8770_ & _8777_ /*32386*/;
assign _8775_ = _8776_ | _8778_ /*32384*/;
assign _8518_ = _8770_ ^ _8777_ /*32387*/;
assign _8784_ = D[49] ^ Q[42] /*32383*/;
assign _8781_ = _8133_ & _8784_ /*32379*/;
assign _8782_ = _8133_ ^ _8784_ /*32382*/;
assign _8783_ = _8775_ & _8782_ /*32380*/;
assign _8780_ = _8781_ | _8783_ /*32378*/;
assign _8519_ = _8775_ ^ _8782_ /*32381*/;
assign _8789_ = D[50] ^ Q[42] /*32377*/;
assign _8786_ = _8134_ & _8789_ /*32373*/;
assign _8787_ = _8134_ ^ _8789_ /*32376*/;
assign _8788_ = _8780_ & _8787_ /*32374*/;
assign _8785_ = _8786_ | _8788_ /*32372*/;
assign _8520_ = _8780_ ^ _8787_ /*32375*/;
assign _8794_ = D[51] ^ Q[42] /*32371*/;
assign _8791_ = _8135_ & _8794_ /*32367*/;
assign _8792_ = _8135_ ^ _8794_ /*32370*/;
assign _8793_ = _8785_ & _8792_ /*32368*/;
assign _8790_ = _8791_ | _8793_ /*32366*/;
assign _8521_ = _8785_ ^ _8792_ /*32369*/;
assign _8799_ = D[52] ^ Q[42] /*32365*/;
assign _8796_ = _8136_ & _8799_ /*32361*/;
assign _8797_ = _8136_ ^ _8799_ /*32364*/;
assign _8798_ = _8790_ & _8797_ /*32362*/;
assign _8795_ = _8796_ | _8798_ /*32360*/;
assign _8522_ = _8790_ ^ _8797_ /*32363*/;
assign _8804_ = D[53] ^ Q[42] /*32359*/;
assign _8801_ = _8137_ & _8804_ /*32355*/;
assign _8802_ = _8137_ ^ _8804_ /*32358*/;
assign _8803_ = _8795_ & _8802_ /*32356*/;
assign _8800_ = _8801_ | _8803_ /*32354*/;
assign _8523_ = _8795_ ^ _8802_ /*32357*/;
assign _8809_ = D[54] ^ Q[42] /*32353*/;
assign _8806_ = _8138_ & _8809_ /*32349*/;
assign _8807_ = _8138_ ^ _8809_ /*32352*/;
assign _8808_ = _8800_ & _8807_ /*32350*/;
assign _8805_ = _8806_ | _8808_ /*32348*/;
assign _8524_ = _8800_ ^ _8807_ /*32351*/;
assign _8814_ = D[55] ^ Q[42] /*32347*/;
assign _8811_ = _8139_ & _8814_ /*32343*/;
assign _8812_ = _8139_ ^ _8814_ /*32346*/;
assign _8813_ = _8805_ & _8812_ /*32344*/;
assign _8810_ = _8811_ | _8813_ /*32342*/;
assign _8525_ = _8805_ ^ _8812_ /*32345*/;
assign _8819_ = D[56] ^ Q[42] /*32341*/;
assign _8816_ = _8140_ & _8819_ /*32337*/;
assign _8817_ = _8140_ ^ _8819_ /*32340*/;
assign _8818_ = _8810_ & _8817_ /*32338*/;
assign _8815_ = _8816_ | _8818_ /*32336*/;
assign _8526_ = _8810_ ^ _8817_ /*32339*/;
assign _8824_ = D[57] ^ Q[42] /*32335*/;
assign _8821_ = _8141_ & _8824_ /*32331*/;
assign _8822_ = _8141_ ^ _8824_ /*32334*/;
assign _8823_ = _8815_ & _8822_ /*32332*/;
assign _8820_ = _8821_ | _8823_ /*32330*/;
assign _8527_ = _8815_ ^ _8822_ /*32333*/;
assign _8829_ = D[58] ^ Q[42] /*32329*/;
assign _8826_ = _8142_ & _8829_ /*32325*/;
assign _8827_ = _8142_ ^ _8829_ /*32328*/;
assign _8828_ = _8820_ & _8827_ /*32326*/;
assign _8825_ = _8826_ | _8828_ /*32324*/;
assign _8528_ = _8820_ ^ _8827_ /*32327*/;
assign _8834_ = D[59] ^ Q[42] /*32323*/;
assign _8831_ = _8143_ & _8834_ /*32319*/;
assign _8832_ = _8143_ ^ _8834_ /*32322*/;
assign _8833_ = _8825_ & _8832_ /*32320*/;
assign _8830_ = _8831_ | _8833_ /*32318*/;
assign _8529_ = _8825_ ^ _8832_ /*32321*/;
assign _8839_ = D[60] ^ Q[42] /*32317*/;
assign _8836_ = _8144_ & _8839_ /*32313*/;
assign _8837_ = _8144_ ^ _8839_ /*32316*/;
assign _8838_ = _8830_ & _8837_ /*32314*/;
assign _8835_ = _8836_ | _8838_ /*32312*/;
assign _8530_ = _8830_ ^ _8837_ /*32315*/;
assign _8844_ = D[61] ^ Q[42] /*32311*/;
assign _8841_ = _8145_ & _8844_ /*32307*/;
assign _8842_ = _8145_ ^ _8844_ /*32310*/;
assign _8843_ = _8835_ & _8842_ /*32308*/;
assign _8840_ = _8841_ | _8843_ /*32306*/;
assign _8531_ = _8835_ ^ _8842_ /*32309*/;
assign _8849_ = D[62] ^ Q[42] /*32305*/;
assign _8846_ = _8146_ & _8849_ /*32301*/;
assign _8847_ = _8146_ ^ _8849_ /*32304*/;
assign _8848_ = _8840_ & _8847_ /*32302*/;
assign _8845_ = _8846_ | _8848_ /*32300*/;
assign _8532_ = _8840_ ^ _8847_ /*32303*/;
assign _8853_ = zeroWire ^ Q[42] /*32299*/;
assign _8850_ = _8147_ & _8853_ /*32295*/;
assign _8851_ = _8147_ ^ _8853_ /*32298*/;
assign _8852_ = _8845_ & _8851_ /*32296*/;
assign Q[41] = _8850_ | _8852_ /*32294*/;
assign _8533_ = _8845_ ^ _8851_ /*32297*/;
assign _8924_ = D[0] ^ Q[41] /*31908*/;
assign _8921_ = R_0[40] & _8924_ /*31904*/;
assign _8922_ = R_0[40] ^ _8924_ /*31907*/;
assign _8923_ = Q[41] & _8922_ /*31905*/;
assign _8920_ = _8921_ | _8923_ /*31903*/;
assign _8855_ = Q[41] ^ _8922_ /*31906*/;
assign _8929_ = D[1] ^ Q[41] /*31902*/;
assign _8926_ = _8470_ & _8929_ /*31898*/;
assign _8927_ = _8470_ ^ _8929_ /*31901*/;
assign _8928_ = _8920_ & _8927_ /*31899*/;
assign _8925_ = _8926_ | _8928_ /*31897*/;
assign _8856_ = _8920_ ^ _8927_ /*31900*/;
assign _8934_ = D[2] ^ Q[41] /*31896*/;
assign _8931_ = _8471_ & _8934_ /*31892*/;
assign _8932_ = _8471_ ^ _8934_ /*31895*/;
assign _8933_ = _8925_ & _8932_ /*31893*/;
assign _8930_ = _8931_ | _8933_ /*31891*/;
assign _8857_ = _8925_ ^ _8932_ /*31894*/;
assign _8939_ = D[3] ^ Q[41] /*31890*/;
assign _8936_ = _8472_ & _8939_ /*31886*/;
assign _8937_ = _8472_ ^ _8939_ /*31889*/;
assign _8938_ = _8930_ & _8937_ /*31887*/;
assign _8935_ = _8936_ | _8938_ /*31885*/;
assign _8858_ = _8930_ ^ _8937_ /*31888*/;
assign _8944_ = D[4] ^ Q[41] /*31884*/;
assign _8941_ = _8473_ & _8944_ /*31880*/;
assign _8942_ = _8473_ ^ _8944_ /*31883*/;
assign _8943_ = _8935_ & _8942_ /*31881*/;
assign _8940_ = _8941_ | _8943_ /*31879*/;
assign _8859_ = _8935_ ^ _8942_ /*31882*/;
assign _8949_ = D[5] ^ Q[41] /*31878*/;
assign _8946_ = _8474_ & _8949_ /*31874*/;
assign _8947_ = _8474_ ^ _8949_ /*31877*/;
assign _8948_ = _8940_ & _8947_ /*31875*/;
assign _8945_ = _8946_ | _8948_ /*31873*/;
assign _8860_ = _8940_ ^ _8947_ /*31876*/;
assign _8954_ = D[6] ^ Q[41] /*31872*/;
assign _8951_ = _8475_ & _8954_ /*31868*/;
assign _8952_ = _8475_ ^ _8954_ /*31871*/;
assign _8953_ = _8945_ & _8952_ /*31869*/;
assign _8950_ = _8951_ | _8953_ /*31867*/;
assign _8861_ = _8945_ ^ _8952_ /*31870*/;
assign _8959_ = D[7] ^ Q[41] /*31866*/;
assign _8956_ = _8476_ & _8959_ /*31862*/;
assign _8957_ = _8476_ ^ _8959_ /*31865*/;
assign _8958_ = _8950_ & _8957_ /*31863*/;
assign _8955_ = _8956_ | _8958_ /*31861*/;
assign _8862_ = _8950_ ^ _8957_ /*31864*/;
assign _8964_ = D[8] ^ Q[41] /*31860*/;
assign _8961_ = _8477_ & _8964_ /*31856*/;
assign _8962_ = _8477_ ^ _8964_ /*31859*/;
assign _8963_ = _8955_ & _8962_ /*31857*/;
assign _8960_ = _8961_ | _8963_ /*31855*/;
assign _8863_ = _8955_ ^ _8962_ /*31858*/;
assign _8969_ = D[9] ^ Q[41] /*31854*/;
assign _8966_ = _8478_ & _8969_ /*31850*/;
assign _8967_ = _8478_ ^ _8969_ /*31853*/;
assign _8968_ = _8960_ & _8967_ /*31851*/;
assign _8965_ = _8966_ | _8968_ /*31849*/;
assign _8864_ = _8960_ ^ _8967_ /*31852*/;
assign _8974_ = D[10] ^ Q[41] /*31848*/;
assign _8971_ = _8479_ & _8974_ /*31844*/;
assign _8972_ = _8479_ ^ _8974_ /*31847*/;
assign _8973_ = _8965_ & _8972_ /*31845*/;
assign _8970_ = _8971_ | _8973_ /*31843*/;
assign _8865_ = _8965_ ^ _8972_ /*31846*/;
assign _8979_ = D[11] ^ Q[41] /*31842*/;
assign _8976_ = _8480_ & _8979_ /*31838*/;
assign _8977_ = _8480_ ^ _8979_ /*31841*/;
assign _8978_ = _8970_ & _8977_ /*31839*/;
assign _8975_ = _8976_ | _8978_ /*31837*/;
assign _8866_ = _8970_ ^ _8977_ /*31840*/;
assign _8984_ = D[12] ^ Q[41] /*31836*/;
assign _8981_ = _8481_ & _8984_ /*31832*/;
assign _8982_ = _8481_ ^ _8984_ /*31835*/;
assign _8983_ = _8975_ & _8982_ /*31833*/;
assign _8980_ = _8981_ | _8983_ /*31831*/;
assign _8867_ = _8975_ ^ _8982_ /*31834*/;
assign _8989_ = D[13] ^ Q[41] /*31830*/;
assign _8986_ = _8482_ & _8989_ /*31826*/;
assign _8987_ = _8482_ ^ _8989_ /*31829*/;
assign _8988_ = _8980_ & _8987_ /*31827*/;
assign _8985_ = _8986_ | _8988_ /*31825*/;
assign _8868_ = _8980_ ^ _8987_ /*31828*/;
assign _8994_ = D[14] ^ Q[41] /*31824*/;
assign _8991_ = _8483_ & _8994_ /*31820*/;
assign _8992_ = _8483_ ^ _8994_ /*31823*/;
assign _8993_ = _8985_ & _8992_ /*31821*/;
assign _8990_ = _8991_ | _8993_ /*31819*/;
assign _8869_ = _8985_ ^ _8992_ /*31822*/;
assign _8999_ = D[15] ^ Q[41] /*31818*/;
assign _8996_ = _8484_ & _8999_ /*31814*/;
assign _8997_ = _8484_ ^ _8999_ /*31817*/;
assign _8998_ = _8990_ & _8997_ /*31815*/;
assign _8995_ = _8996_ | _8998_ /*31813*/;
assign _8870_ = _8990_ ^ _8997_ /*31816*/;
assign _9004_ = D[16] ^ Q[41] /*31812*/;
assign _9001_ = _8485_ & _9004_ /*31808*/;
assign _9002_ = _8485_ ^ _9004_ /*31811*/;
assign _9003_ = _8995_ & _9002_ /*31809*/;
assign _9000_ = _9001_ | _9003_ /*31807*/;
assign _8871_ = _8995_ ^ _9002_ /*31810*/;
assign _9009_ = D[17] ^ Q[41] /*31806*/;
assign _9006_ = _8486_ & _9009_ /*31802*/;
assign _9007_ = _8486_ ^ _9009_ /*31805*/;
assign _9008_ = _9000_ & _9007_ /*31803*/;
assign _9005_ = _9006_ | _9008_ /*31801*/;
assign _8872_ = _9000_ ^ _9007_ /*31804*/;
assign _9014_ = D[18] ^ Q[41] /*31800*/;
assign _9011_ = _8487_ & _9014_ /*31796*/;
assign _9012_ = _8487_ ^ _9014_ /*31799*/;
assign _9013_ = _9005_ & _9012_ /*31797*/;
assign _9010_ = _9011_ | _9013_ /*31795*/;
assign _8873_ = _9005_ ^ _9012_ /*31798*/;
assign _9019_ = D[19] ^ Q[41] /*31794*/;
assign _9016_ = _8488_ & _9019_ /*31790*/;
assign _9017_ = _8488_ ^ _9019_ /*31793*/;
assign _9018_ = _9010_ & _9017_ /*31791*/;
assign _9015_ = _9016_ | _9018_ /*31789*/;
assign _8874_ = _9010_ ^ _9017_ /*31792*/;
assign _9024_ = D[20] ^ Q[41] /*31788*/;
assign _9021_ = _8489_ & _9024_ /*31784*/;
assign _9022_ = _8489_ ^ _9024_ /*31787*/;
assign _9023_ = _9015_ & _9022_ /*31785*/;
assign _9020_ = _9021_ | _9023_ /*31783*/;
assign _8875_ = _9015_ ^ _9022_ /*31786*/;
assign _9029_ = D[21] ^ Q[41] /*31782*/;
assign _9026_ = _8490_ & _9029_ /*31778*/;
assign _9027_ = _8490_ ^ _9029_ /*31781*/;
assign _9028_ = _9020_ & _9027_ /*31779*/;
assign _9025_ = _9026_ | _9028_ /*31777*/;
assign _8876_ = _9020_ ^ _9027_ /*31780*/;
assign _9034_ = D[22] ^ Q[41] /*31776*/;
assign _9031_ = _8491_ & _9034_ /*31772*/;
assign _9032_ = _8491_ ^ _9034_ /*31775*/;
assign _9033_ = _9025_ & _9032_ /*31773*/;
assign _9030_ = _9031_ | _9033_ /*31771*/;
assign _8877_ = _9025_ ^ _9032_ /*31774*/;
assign _9039_ = D[23] ^ Q[41] /*31770*/;
assign _9036_ = _8492_ & _9039_ /*31766*/;
assign _9037_ = _8492_ ^ _9039_ /*31769*/;
assign _9038_ = _9030_ & _9037_ /*31767*/;
assign _9035_ = _9036_ | _9038_ /*31765*/;
assign _8878_ = _9030_ ^ _9037_ /*31768*/;
assign _9044_ = D[24] ^ Q[41] /*31764*/;
assign _9041_ = _8493_ & _9044_ /*31760*/;
assign _9042_ = _8493_ ^ _9044_ /*31763*/;
assign _9043_ = _9035_ & _9042_ /*31761*/;
assign _9040_ = _9041_ | _9043_ /*31759*/;
assign _8879_ = _9035_ ^ _9042_ /*31762*/;
assign _9049_ = D[25] ^ Q[41] /*31758*/;
assign _9046_ = _8494_ & _9049_ /*31754*/;
assign _9047_ = _8494_ ^ _9049_ /*31757*/;
assign _9048_ = _9040_ & _9047_ /*31755*/;
assign _9045_ = _9046_ | _9048_ /*31753*/;
assign _8880_ = _9040_ ^ _9047_ /*31756*/;
assign _9054_ = D[26] ^ Q[41] /*31752*/;
assign _9051_ = _8495_ & _9054_ /*31748*/;
assign _9052_ = _8495_ ^ _9054_ /*31751*/;
assign _9053_ = _9045_ & _9052_ /*31749*/;
assign _9050_ = _9051_ | _9053_ /*31747*/;
assign _8881_ = _9045_ ^ _9052_ /*31750*/;
assign _9059_ = D[27] ^ Q[41] /*31746*/;
assign _9056_ = _8496_ & _9059_ /*31742*/;
assign _9057_ = _8496_ ^ _9059_ /*31745*/;
assign _9058_ = _9050_ & _9057_ /*31743*/;
assign _9055_ = _9056_ | _9058_ /*31741*/;
assign _8882_ = _9050_ ^ _9057_ /*31744*/;
assign _9064_ = D[28] ^ Q[41] /*31740*/;
assign _9061_ = _8497_ & _9064_ /*31736*/;
assign _9062_ = _8497_ ^ _9064_ /*31739*/;
assign _9063_ = _9055_ & _9062_ /*31737*/;
assign _9060_ = _9061_ | _9063_ /*31735*/;
assign _8883_ = _9055_ ^ _9062_ /*31738*/;
assign _9069_ = D[29] ^ Q[41] /*31734*/;
assign _9066_ = _8498_ & _9069_ /*31730*/;
assign _9067_ = _8498_ ^ _9069_ /*31733*/;
assign _9068_ = _9060_ & _9067_ /*31731*/;
assign _9065_ = _9066_ | _9068_ /*31729*/;
assign _8884_ = _9060_ ^ _9067_ /*31732*/;
assign _9074_ = D[30] ^ Q[41] /*31728*/;
assign _9071_ = _8499_ & _9074_ /*31724*/;
assign _9072_ = _8499_ ^ _9074_ /*31727*/;
assign _9073_ = _9065_ & _9072_ /*31725*/;
assign _9070_ = _9071_ | _9073_ /*31723*/;
assign _8885_ = _9065_ ^ _9072_ /*31726*/;
assign _9079_ = D[31] ^ Q[41] /*31722*/;
assign _9076_ = _8500_ & _9079_ /*31718*/;
assign _9077_ = _8500_ ^ _9079_ /*31721*/;
assign _9078_ = _9070_ & _9077_ /*31719*/;
assign _9075_ = _9076_ | _9078_ /*31717*/;
assign _8886_ = _9070_ ^ _9077_ /*31720*/;
assign _9084_ = D[32] ^ Q[41] /*31716*/;
assign _9081_ = _8501_ & _9084_ /*31712*/;
assign _9082_ = _8501_ ^ _9084_ /*31715*/;
assign _9083_ = _9075_ & _9082_ /*31713*/;
assign _9080_ = _9081_ | _9083_ /*31711*/;
assign _8887_ = _9075_ ^ _9082_ /*31714*/;
assign _9089_ = D[33] ^ Q[41] /*31710*/;
assign _9086_ = _8502_ & _9089_ /*31706*/;
assign _9087_ = _8502_ ^ _9089_ /*31709*/;
assign _9088_ = _9080_ & _9087_ /*31707*/;
assign _9085_ = _9086_ | _9088_ /*31705*/;
assign _8888_ = _9080_ ^ _9087_ /*31708*/;
assign _9094_ = D[34] ^ Q[41] /*31704*/;
assign _9091_ = _8503_ & _9094_ /*31700*/;
assign _9092_ = _8503_ ^ _9094_ /*31703*/;
assign _9093_ = _9085_ & _9092_ /*31701*/;
assign _9090_ = _9091_ | _9093_ /*31699*/;
assign _8889_ = _9085_ ^ _9092_ /*31702*/;
assign _9099_ = D[35] ^ Q[41] /*31698*/;
assign _9096_ = _8504_ & _9099_ /*31694*/;
assign _9097_ = _8504_ ^ _9099_ /*31697*/;
assign _9098_ = _9090_ & _9097_ /*31695*/;
assign _9095_ = _9096_ | _9098_ /*31693*/;
assign _8890_ = _9090_ ^ _9097_ /*31696*/;
assign _9104_ = D[36] ^ Q[41] /*31692*/;
assign _9101_ = _8505_ & _9104_ /*31688*/;
assign _9102_ = _8505_ ^ _9104_ /*31691*/;
assign _9103_ = _9095_ & _9102_ /*31689*/;
assign _9100_ = _9101_ | _9103_ /*31687*/;
assign _8891_ = _9095_ ^ _9102_ /*31690*/;
assign _9109_ = D[37] ^ Q[41] /*31686*/;
assign _9106_ = _8506_ & _9109_ /*31682*/;
assign _9107_ = _8506_ ^ _9109_ /*31685*/;
assign _9108_ = _9100_ & _9107_ /*31683*/;
assign _9105_ = _9106_ | _9108_ /*31681*/;
assign _8892_ = _9100_ ^ _9107_ /*31684*/;
assign _9114_ = D[38] ^ Q[41] /*31680*/;
assign _9111_ = _8507_ & _9114_ /*31676*/;
assign _9112_ = _8507_ ^ _9114_ /*31679*/;
assign _9113_ = _9105_ & _9112_ /*31677*/;
assign _9110_ = _9111_ | _9113_ /*31675*/;
assign _8893_ = _9105_ ^ _9112_ /*31678*/;
assign _9119_ = D[39] ^ Q[41] /*31674*/;
assign _9116_ = _8508_ & _9119_ /*31670*/;
assign _9117_ = _8508_ ^ _9119_ /*31673*/;
assign _9118_ = _9110_ & _9117_ /*31671*/;
assign _9115_ = _9116_ | _9118_ /*31669*/;
assign _8894_ = _9110_ ^ _9117_ /*31672*/;
assign _9124_ = D[40] ^ Q[41] /*31668*/;
assign _9121_ = _8509_ & _9124_ /*31664*/;
assign _9122_ = _8509_ ^ _9124_ /*31667*/;
assign _9123_ = _9115_ & _9122_ /*31665*/;
assign _9120_ = _9121_ | _9123_ /*31663*/;
assign _8895_ = _9115_ ^ _9122_ /*31666*/;
assign _9129_ = D[41] ^ Q[41] /*31662*/;
assign _9126_ = _8510_ & _9129_ /*31658*/;
assign _9127_ = _8510_ ^ _9129_ /*31661*/;
assign _9128_ = _9120_ & _9127_ /*31659*/;
assign _9125_ = _9126_ | _9128_ /*31657*/;
assign _8896_ = _9120_ ^ _9127_ /*31660*/;
assign _9134_ = D[42] ^ Q[41] /*31656*/;
assign _9131_ = _8511_ & _9134_ /*31652*/;
assign _9132_ = _8511_ ^ _9134_ /*31655*/;
assign _9133_ = _9125_ & _9132_ /*31653*/;
assign _9130_ = _9131_ | _9133_ /*31651*/;
assign _8897_ = _9125_ ^ _9132_ /*31654*/;
assign _9139_ = D[43] ^ Q[41] /*31650*/;
assign _9136_ = _8512_ & _9139_ /*31646*/;
assign _9137_ = _8512_ ^ _9139_ /*31649*/;
assign _9138_ = _9130_ & _9137_ /*31647*/;
assign _9135_ = _9136_ | _9138_ /*31645*/;
assign _8898_ = _9130_ ^ _9137_ /*31648*/;
assign _9144_ = D[44] ^ Q[41] /*31644*/;
assign _9141_ = _8513_ & _9144_ /*31640*/;
assign _9142_ = _8513_ ^ _9144_ /*31643*/;
assign _9143_ = _9135_ & _9142_ /*31641*/;
assign _9140_ = _9141_ | _9143_ /*31639*/;
assign _8899_ = _9135_ ^ _9142_ /*31642*/;
assign _9149_ = D[45] ^ Q[41] /*31638*/;
assign _9146_ = _8514_ & _9149_ /*31634*/;
assign _9147_ = _8514_ ^ _9149_ /*31637*/;
assign _9148_ = _9140_ & _9147_ /*31635*/;
assign _9145_ = _9146_ | _9148_ /*31633*/;
assign _8900_ = _9140_ ^ _9147_ /*31636*/;
assign _9154_ = D[46] ^ Q[41] /*31632*/;
assign _9151_ = _8515_ & _9154_ /*31628*/;
assign _9152_ = _8515_ ^ _9154_ /*31631*/;
assign _9153_ = _9145_ & _9152_ /*31629*/;
assign _9150_ = _9151_ | _9153_ /*31627*/;
assign _8901_ = _9145_ ^ _9152_ /*31630*/;
assign _9159_ = D[47] ^ Q[41] /*31626*/;
assign _9156_ = _8516_ & _9159_ /*31622*/;
assign _9157_ = _8516_ ^ _9159_ /*31625*/;
assign _9158_ = _9150_ & _9157_ /*31623*/;
assign _9155_ = _9156_ | _9158_ /*31621*/;
assign _8902_ = _9150_ ^ _9157_ /*31624*/;
assign _9164_ = D[48] ^ Q[41] /*31620*/;
assign _9161_ = _8517_ & _9164_ /*31616*/;
assign _9162_ = _8517_ ^ _9164_ /*31619*/;
assign _9163_ = _9155_ & _9162_ /*31617*/;
assign _9160_ = _9161_ | _9163_ /*31615*/;
assign _8903_ = _9155_ ^ _9162_ /*31618*/;
assign _9169_ = D[49] ^ Q[41] /*31614*/;
assign _9166_ = _8518_ & _9169_ /*31610*/;
assign _9167_ = _8518_ ^ _9169_ /*31613*/;
assign _9168_ = _9160_ & _9167_ /*31611*/;
assign _9165_ = _9166_ | _9168_ /*31609*/;
assign _8904_ = _9160_ ^ _9167_ /*31612*/;
assign _9174_ = D[50] ^ Q[41] /*31608*/;
assign _9171_ = _8519_ & _9174_ /*31604*/;
assign _9172_ = _8519_ ^ _9174_ /*31607*/;
assign _9173_ = _9165_ & _9172_ /*31605*/;
assign _9170_ = _9171_ | _9173_ /*31603*/;
assign _8905_ = _9165_ ^ _9172_ /*31606*/;
assign _9179_ = D[51] ^ Q[41] /*31602*/;
assign _9176_ = _8520_ & _9179_ /*31598*/;
assign _9177_ = _8520_ ^ _9179_ /*31601*/;
assign _9178_ = _9170_ & _9177_ /*31599*/;
assign _9175_ = _9176_ | _9178_ /*31597*/;
assign _8906_ = _9170_ ^ _9177_ /*31600*/;
assign _9184_ = D[52] ^ Q[41] /*31596*/;
assign _9181_ = _8521_ & _9184_ /*31592*/;
assign _9182_ = _8521_ ^ _9184_ /*31595*/;
assign _9183_ = _9175_ & _9182_ /*31593*/;
assign _9180_ = _9181_ | _9183_ /*31591*/;
assign _8907_ = _9175_ ^ _9182_ /*31594*/;
assign _9189_ = D[53] ^ Q[41] /*31590*/;
assign _9186_ = _8522_ & _9189_ /*31586*/;
assign _9187_ = _8522_ ^ _9189_ /*31589*/;
assign _9188_ = _9180_ & _9187_ /*31587*/;
assign _9185_ = _9186_ | _9188_ /*31585*/;
assign _8908_ = _9180_ ^ _9187_ /*31588*/;
assign _9194_ = D[54] ^ Q[41] /*31584*/;
assign _9191_ = _8523_ & _9194_ /*31580*/;
assign _9192_ = _8523_ ^ _9194_ /*31583*/;
assign _9193_ = _9185_ & _9192_ /*31581*/;
assign _9190_ = _9191_ | _9193_ /*31579*/;
assign _8909_ = _9185_ ^ _9192_ /*31582*/;
assign _9199_ = D[55] ^ Q[41] /*31578*/;
assign _9196_ = _8524_ & _9199_ /*31574*/;
assign _9197_ = _8524_ ^ _9199_ /*31577*/;
assign _9198_ = _9190_ & _9197_ /*31575*/;
assign _9195_ = _9196_ | _9198_ /*31573*/;
assign _8910_ = _9190_ ^ _9197_ /*31576*/;
assign _9204_ = D[56] ^ Q[41] /*31572*/;
assign _9201_ = _8525_ & _9204_ /*31568*/;
assign _9202_ = _8525_ ^ _9204_ /*31571*/;
assign _9203_ = _9195_ & _9202_ /*31569*/;
assign _9200_ = _9201_ | _9203_ /*31567*/;
assign _8911_ = _9195_ ^ _9202_ /*31570*/;
assign _9209_ = D[57] ^ Q[41] /*31566*/;
assign _9206_ = _8526_ & _9209_ /*31562*/;
assign _9207_ = _8526_ ^ _9209_ /*31565*/;
assign _9208_ = _9200_ & _9207_ /*31563*/;
assign _9205_ = _9206_ | _9208_ /*31561*/;
assign _8912_ = _9200_ ^ _9207_ /*31564*/;
assign _9214_ = D[58] ^ Q[41] /*31560*/;
assign _9211_ = _8527_ & _9214_ /*31556*/;
assign _9212_ = _8527_ ^ _9214_ /*31559*/;
assign _9213_ = _9205_ & _9212_ /*31557*/;
assign _9210_ = _9211_ | _9213_ /*31555*/;
assign _8913_ = _9205_ ^ _9212_ /*31558*/;
assign _9219_ = D[59] ^ Q[41] /*31554*/;
assign _9216_ = _8528_ & _9219_ /*31550*/;
assign _9217_ = _8528_ ^ _9219_ /*31553*/;
assign _9218_ = _9210_ & _9217_ /*31551*/;
assign _9215_ = _9216_ | _9218_ /*31549*/;
assign _8914_ = _9210_ ^ _9217_ /*31552*/;
assign _9224_ = D[60] ^ Q[41] /*31548*/;
assign _9221_ = _8529_ & _9224_ /*31544*/;
assign _9222_ = _8529_ ^ _9224_ /*31547*/;
assign _9223_ = _9215_ & _9222_ /*31545*/;
assign _9220_ = _9221_ | _9223_ /*31543*/;
assign _8915_ = _9215_ ^ _9222_ /*31546*/;
assign _9229_ = D[61] ^ Q[41] /*31542*/;
assign _9226_ = _8530_ & _9229_ /*31538*/;
assign _9227_ = _8530_ ^ _9229_ /*31541*/;
assign _9228_ = _9220_ & _9227_ /*31539*/;
assign _9225_ = _9226_ | _9228_ /*31537*/;
assign _8916_ = _9220_ ^ _9227_ /*31540*/;
assign _9234_ = D[62] ^ Q[41] /*31536*/;
assign _9231_ = _8531_ & _9234_ /*31532*/;
assign _9232_ = _8531_ ^ _9234_ /*31535*/;
assign _9233_ = _9225_ & _9232_ /*31533*/;
assign _9230_ = _9231_ | _9233_ /*31531*/;
assign _8917_ = _9225_ ^ _9232_ /*31534*/;
assign _9238_ = zeroWire ^ Q[41] /*31530*/;
assign _9235_ = _8532_ & _9238_ /*31526*/;
assign _9236_ = _8532_ ^ _9238_ /*31529*/;
assign _9237_ = _9230_ & _9236_ /*31527*/;
assign Q[40] = _9235_ | _9237_ /*31525*/;
assign _8918_ = _9230_ ^ _9236_ /*31528*/;
assign _9309_ = D[0] ^ Q[40] /*31139*/;
assign _9306_ = R_0[39] & _9309_ /*31135*/;
assign _9307_ = R_0[39] ^ _9309_ /*31138*/;
assign _9308_ = Q[40] & _9307_ /*31136*/;
assign _9305_ = _9306_ | _9308_ /*31134*/;
assign _9240_ = Q[40] ^ _9307_ /*31137*/;
assign _9314_ = D[1] ^ Q[40] /*31133*/;
assign _9311_ = _8855_ & _9314_ /*31129*/;
assign _9312_ = _8855_ ^ _9314_ /*31132*/;
assign _9313_ = _9305_ & _9312_ /*31130*/;
assign _9310_ = _9311_ | _9313_ /*31128*/;
assign _9241_ = _9305_ ^ _9312_ /*31131*/;
assign _9319_ = D[2] ^ Q[40] /*31127*/;
assign _9316_ = _8856_ & _9319_ /*31123*/;
assign _9317_ = _8856_ ^ _9319_ /*31126*/;
assign _9318_ = _9310_ & _9317_ /*31124*/;
assign _9315_ = _9316_ | _9318_ /*31122*/;
assign _9242_ = _9310_ ^ _9317_ /*31125*/;
assign _9324_ = D[3] ^ Q[40] /*31121*/;
assign _9321_ = _8857_ & _9324_ /*31117*/;
assign _9322_ = _8857_ ^ _9324_ /*31120*/;
assign _9323_ = _9315_ & _9322_ /*31118*/;
assign _9320_ = _9321_ | _9323_ /*31116*/;
assign _9243_ = _9315_ ^ _9322_ /*31119*/;
assign _9329_ = D[4] ^ Q[40] /*31115*/;
assign _9326_ = _8858_ & _9329_ /*31111*/;
assign _9327_ = _8858_ ^ _9329_ /*31114*/;
assign _9328_ = _9320_ & _9327_ /*31112*/;
assign _9325_ = _9326_ | _9328_ /*31110*/;
assign _9244_ = _9320_ ^ _9327_ /*31113*/;
assign _9334_ = D[5] ^ Q[40] /*31109*/;
assign _9331_ = _8859_ & _9334_ /*31105*/;
assign _9332_ = _8859_ ^ _9334_ /*31108*/;
assign _9333_ = _9325_ & _9332_ /*31106*/;
assign _9330_ = _9331_ | _9333_ /*31104*/;
assign _9245_ = _9325_ ^ _9332_ /*31107*/;
assign _9339_ = D[6] ^ Q[40] /*31103*/;
assign _9336_ = _8860_ & _9339_ /*31099*/;
assign _9337_ = _8860_ ^ _9339_ /*31102*/;
assign _9338_ = _9330_ & _9337_ /*31100*/;
assign _9335_ = _9336_ | _9338_ /*31098*/;
assign _9246_ = _9330_ ^ _9337_ /*31101*/;
assign _9344_ = D[7] ^ Q[40] /*31097*/;
assign _9341_ = _8861_ & _9344_ /*31093*/;
assign _9342_ = _8861_ ^ _9344_ /*31096*/;
assign _9343_ = _9335_ & _9342_ /*31094*/;
assign _9340_ = _9341_ | _9343_ /*31092*/;
assign _9247_ = _9335_ ^ _9342_ /*31095*/;
assign _9349_ = D[8] ^ Q[40] /*31091*/;
assign _9346_ = _8862_ & _9349_ /*31087*/;
assign _9347_ = _8862_ ^ _9349_ /*31090*/;
assign _9348_ = _9340_ & _9347_ /*31088*/;
assign _9345_ = _9346_ | _9348_ /*31086*/;
assign _9248_ = _9340_ ^ _9347_ /*31089*/;
assign _9354_ = D[9] ^ Q[40] /*31085*/;
assign _9351_ = _8863_ & _9354_ /*31081*/;
assign _9352_ = _8863_ ^ _9354_ /*31084*/;
assign _9353_ = _9345_ & _9352_ /*31082*/;
assign _9350_ = _9351_ | _9353_ /*31080*/;
assign _9249_ = _9345_ ^ _9352_ /*31083*/;
assign _9359_ = D[10] ^ Q[40] /*31079*/;
assign _9356_ = _8864_ & _9359_ /*31075*/;
assign _9357_ = _8864_ ^ _9359_ /*31078*/;
assign _9358_ = _9350_ & _9357_ /*31076*/;
assign _9355_ = _9356_ | _9358_ /*31074*/;
assign _9250_ = _9350_ ^ _9357_ /*31077*/;
assign _9364_ = D[11] ^ Q[40] /*31073*/;
assign _9361_ = _8865_ & _9364_ /*31069*/;
assign _9362_ = _8865_ ^ _9364_ /*31072*/;
assign _9363_ = _9355_ & _9362_ /*31070*/;
assign _9360_ = _9361_ | _9363_ /*31068*/;
assign _9251_ = _9355_ ^ _9362_ /*31071*/;
assign _9369_ = D[12] ^ Q[40] /*31067*/;
assign _9366_ = _8866_ & _9369_ /*31063*/;
assign _9367_ = _8866_ ^ _9369_ /*31066*/;
assign _9368_ = _9360_ & _9367_ /*31064*/;
assign _9365_ = _9366_ | _9368_ /*31062*/;
assign _9252_ = _9360_ ^ _9367_ /*31065*/;
assign _9374_ = D[13] ^ Q[40] /*31061*/;
assign _9371_ = _8867_ & _9374_ /*31057*/;
assign _9372_ = _8867_ ^ _9374_ /*31060*/;
assign _9373_ = _9365_ & _9372_ /*31058*/;
assign _9370_ = _9371_ | _9373_ /*31056*/;
assign _9253_ = _9365_ ^ _9372_ /*31059*/;
assign _9379_ = D[14] ^ Q[40] /*31055*/;
assign _9376_ = _8868_ & _9379_ /*31051*/;
assign _9377_ = _8868_ ^ _9379_ /*31054*/;
assign _9378_ = _9370_ & _9377_ /*31052*/;
assign _9375_ = _9376_ | _9378_ /*31050*/;
assign _9254_ = _9370_ ^ _9377_ /*31053*/;
assign _9384_ = D[15] ^ Q[40] /*31049*/;
assign _9381_ = _8869_ & _9384_ /*31045*/;
assign _9382_ = _8869_ ^ _9384_ /*31048*/;
assign _9383_ = _9375_ & _9382_ /*31046*/;
assign _9380_ = _9381_ | _9383_ /*31044*/;
assign _9255_ = _9375_ ^ _9382_ /*31047*/;
assign _9389_ = D[16] ^ Q[40] /*31043*/;
assign _9386_ = _8870_ & _9389_ /*31039*/;
assign _9387_ = _8870_ ^ _9389_ /*31042*/;
assign _9388_ = _9380_ & _9387_ /*31040*/;
assign _9385_ = _9386_ | _9388_ /*31038*/;
assign _9256_ = _9380_ ^ _9387_ /*31041*/;
assign _9394_ = D[17] ^ Q[40] /*31037*/;
assign _9391_ = _8871_ & _9394_ /*31033*/;
assign _9392_ = _8871_ ^ _9394_ /*31036*/;
assign _9393_ = _9385_ & _9392_ /*31034*/;
assign _9390_ = _9391_ | _9393_ /*31032*/;
assign _9257_ = _9385_ ^ _9392_ /*31035*/;
assign _9399_ = D[18] ^ Q[40] /*31031*/;
assign _9396_ = _8872_ & _9399_ /*31027*/;
assign _9397_ = _8872_ ^ _9399_ /*31030*/;
assign _9398_ = _9390_ & _9397_ /*31028*/;
assign _9395_ = _9396_ | _9398_ /*31026*/;
assign _9258_ = _9390_ ^ _9397_ /*31029*/;
assign _9404_ = D[19] ^ Q[40] /*31025*/;
assign _9401_ = _8873_ & _9404_ /*31021*/;
assign _9402_ = _8873_ ^ _9404_ /*31024*/;
assign _9403_ = _9395_ & _9402_ /*31022*/;
assign _9400_ = _9401_ | _9403_ /*31020*/;
assign _9259_ = _9395_ ^ _9402_ /*31023*/;
assign _9409_ = D[20] ^ Q[40] /*31019*/;
assign _9406_ = _8874_ & _9409_ /*31015*/;
assign _9407_ = _8874_ ^ _9409_ /*31018*/;
assign _9408_ = _9400_ & _9407_ /*31016*/;
assign _9405_ = _9406_ | _9408_ /*31014*/;
assign _9260_ = _9400_ ^ _9407_ /*31017*/;
assign _9414_ = D[21] ^ Q[40] /*31013*/;
assign _9411_ = _8875_ & _9414_ /*31009*/;
assign _9412_ = _8875_ ^ _9414_ /*31012*/;
assign _9413_ = _9405_ & _9412_ /*31010*/;
assign _9410_ = _9411_ | _9413_ /*31008*/;
assign _9261_ = _9405_ ^ _9412_ /*31011*/;
assign _9419_ = D[22] ^ Q[40] /*31007*/;
assign _9416_ = _8876_ & _9419_ /*31003*/;
assign _9417_ = _8876_ ^ _9419_ /*31006*/;
assign _9418_ = _9410_ & _9417_ /*31004*/;
assign _9415_ = _9416_ | _9418_ /*31002*/;
assign _9262_ = _9410_ ^ _9417_ /*31005*/;
assign _9424_ = D[23] ^ Q[40] /*31001*/;
assign _9421_ = _8877_ & _9424_ /*30997*/;
assign _9422_ = _8877_ ^ _9424_ /*31000*/;
assign _9423_ = _9415_ & _9422_ /*30998*/;
assign _9420_ = _9421_ | _9423_ /*30996*/;
assign _9263_ = _9415_ ^ _9422_ /*30999*/;
assign _9429_ = D[24] ^ Q[40] /*30995*/;
assign _9426_ = _8878_ & _9429_ /*30991*/;
assign _9427_ = _8878_ ^ _9429_ /*30994*/;
assign _9428_ = _9420_ & _9427_ /*30992*/;
assign _9425_ = _9426_ | _9428_ /*30990*/;
assign _9264_ = _9420_ ^ _9427_ /*30993*/;
assign _9434_ = D[25] ^ Q[40] /*30989*/;
assign _9431_ = _8879_ & _9434_ /*30985*/;
assign _9432_ = _8879_ ^ _9434_ /*30988*/;
assign _9433_ = _9425_ & _9432_ /*30986*/;
assign _9430_ = _9431_ | _9433_ /*30984*/;
assign _9265_ = _9425_ ^ _9432_ /*30987*/;
assign _9439_ = D[26] ^ Q[40] /*30983*/;
assign _9436_ = _8880_ & _9439_ /*30979*/;
assign _9437_ = _8880_ ^ _9439_ /*30982*/;
assign _9438_ = _9430_ & _9437_ /*30980*/;
assign _9435_ = _9436_ | _9438_ /*30978*/;
assign _9266_ = _9430_ ^ _9437_ /*30981*/;
assign _9444_ = D[27] ^ Q[40] /*30977*/;
assign _9441_ = _8881_ & _9444_ /*30973*/;
assign _9442_ = _8881_ ^ _9444_ /*30976*/;
assign _9443_ = _9435_ & _9442_ /*30974*/;
assign _9440_ = _9441_ | _9443_ /*30972*/;
assign _9267_ = _9435_ ^ _9442_ /*30975*/;
assign _9449_ = D[28] ^ Q[40] /*30971*/;
assign _9446_ = _8882_ & _9449_ /*30967*/;
assign _9447_ = _8882_ ^ _9449_ /*30970*/;
assign _9448_ = _9440_ & _9447_ /*30968*/;
assign _9445_ = _9446_ | _9448_ /*30966*/;
assign _9268_ = _9440_ ^ _9447_ /*30969*/;
assign _9454_ = D[29] ^ Q[40] /*30965*/;
assign _9451_ = _8883_ & _9454_ /*30961*/;
assign _9452_ = _8883_ ^ _9454_ /*30964*/;
assign _9453_ = _9445_ & _9452_ /*30962*/;
assign _9450_ = _9451_ | _9453_ /*30960*/;
assign _9269_ = _9445_ ^ _9452_ /*30963*/;
assign _9459_ = D[30] ^ Q[40] /*30959*/;
assign _9456_ = _8884_ & _9459_ /*30955*/;
assign _9457_ = _8884_ ^ _9459_ /*30958*/;
assign _9458_ = _9450_ & _9457_ /*30956*/;
assign _9455_ = _9456_ | _9458_ /*30954*/;
assign _9270_ = _9450_ ^ _9457_ /*30957*/;
assign _9464_ = D[31] ^ Q[40] /*30953*/;
assign _9461_ = _8885_ & _9464_ /*30949*/;
assign _9462_ = _8885_ ^ _9464_ /*30952*/;
assign _9463_ = _9455_ & _9462_ /*30950*/;
assign _9460_ = _9461_ | _9463_ /*30948*/;
assign _9271_ = _9455_ ^ _9462_ /*30951*/;
assign _9469_ = D[32] ^ Q[40] /*30947*/;
assign _9466_ = _8886_ & _9469_ /*30943*/;
assign _9467_ = _8886_ ^ _9469_ /*30946*/;
assign _9468_ = _9460_ & _9467_ /*30944*/;
assign _9465_ = _9466_ | _9468_ /*30942*/;
assign _9272_ = _9460_ ^ _9467_ /*30945*/;
assign _9474_ = D[33] ^ Q[40] /*30941*/;
assign _9471_ = _8887_ & _9474_ /*30937*/;
assign _9472_ = _8887_ ^ _9474_ /*30940*/;
assign _9473_ = _9465_ & _9472_ /*30938*/;
assign _9470_ = _9471_ | _9473_ /*30936*/;
assign _9273_ = _9465_ ^ _9472_ /*30939*/;
assign _9479_ = D[34] ^ Q[40] /*30935*/;
assign _9476_ = _8888_ & _9479_ /*30931*/;
assign _9477_ = _8888_ ^ _9479_ /*30934*/;
assign _9478_ = _9470_ & _9477_ /*30932*/;
assign _9475_ = _9476_ | _9478_ /*30930*/;
assign _9274_ = _9470_ ^ _9477_ /*30933*/;
assign _9484_ = D[35] ^ Q[40] /*30929*/;
assign _9481_ = _8889_ & _9484_ /*30925*/;
assign _9482_ = _8889_ ^ _9484_ /*30928*/;
assign _9483_ = _9475_ & _9482_ /*30926*/;
assign _9480_ = _9481_ | _9483_ /*30924*/;
assign _9275_ = _9475_ ^ _9482_ /*30927*/;
assign _9489_ = D[36] ^ Q[40] /*30923*/;
assign _9486_ = _8890_ & _9489_ /*30919*/;
assign _9487_ = _8890_ ^ _9489_ /*30922*/;
assign _9488_ = _9480_ & _9487_ /*30920*/;
assign _9485_ = _9486_ | _9488_ /*30918*/;
assign _9276_ = _9480_ ^ _9487_ /*30921*/;
assign _9494_ = D[37] ^ Q[40] /*30917*/;
assign _9491_ = _8891_ & _9494_ /*30913*/;
assign _9492_ = _8891_ ^ _9494_ /*30916*/;
assign _9493_ = _9485_ & _9492_ /*30914*/;
assign _9490_ = _9491_ | _9493_ /*30912*/;
assign _9277_ = _9485_ ^ _9492_ /*30915*/;
assign _9499_ = D[38] ^ Q[40] /*30911*/;
assign _9496_ = _8892_ & _9499_ /*30907*/;
assign _9497_ = _8892_ ^ _9499_ /*30910*/;
assign _9498_ = _9490_ & _9497_ /*30908*/;
assign _9495_ = _9496_ | _9498_ /*30906*/;
assign _9278_ = _9490_ ^ _9497_ /*30909*/;
assign _9504_ = D[39] ^ Q[40] /*30905*/;
assign _9501_ = _8893_ & _9504_ /*30901*/;
assign _9502_ = _8893_ ^ _9504_ /*30904*/;
assign _9503_ = _9495_ & _9502_ /*30902*/;
assign _9500_ = _9501_ | _9503_ /*30900*/;
assign _9279_ = _9495_ ^ _9502_ /*30903*/;
assign _9509_ = D[40] ^ Q[40] /*30899*/;
assign _9506_ = _8894_ & _9509_ /*30895*/;
assign _9507_ = _8894_ ^ _9509_ /*30898*/;
assign _9508_ = _9500_ & _9507_ /*30896*/;
assign _9505_ = _9506_ | _9508_ /*30894*/;
assign _9280_ = _9500_ ^ _9507_ /*30897*/;
assign _9514_ = D[41] ^ Q[40] /*30893*/;
assign _9511_ = _8895_ & _9514_ /*30889*/;
assign _9512_ = _8895_ ^ _9514_ /*30892*/;
assign _9513_ = _9505_ & _9512_ /*30890*/;
assign _9510_ = _9511_ | _9513_ /*30888*/;
assign _9281_ = _9505_ ^ _9512_ /*30891*/;
assign _9519_ = D[42] ^ Q[40] /*30887*/;
assign _9516_ = _8896_ & _9519_ /*30883*/;
assign _9517_ = _8896_ ^ _9519_ /*30886*/;
assign _9518_ = _9510_ & _9517_ /*30884*/;
assign _9515_ = _9516_ | _9518_ /*30882*/;
assign _9282_ = _9510_ ^ _9517_ /*30885*/;
assign _9524_ = D[43] ^ Q[40] /*30881*/;
assign _9521_ = _8897_ & _9524_ /*30877*/;
assign _9522_ = _8897_ ^ _9524_ /*30880*/;
assign _9523_ = _9515_ & _9522_ /*30878*/;
assign _9520_ = _9521_ | _9523_ /*30876*/;
assign _9283_ = _9515_ ^ _9522_ /*30879*/;
assign _9529_ = D[44] ^ Q[40] /*30875*/;
assign _9526_ = _8898_ & _9529_ /*30871*/;
assign _9527_ = _8898_ ^ _9529_ /*30874*/;
assign _9528_ = _9520_ & _9527_ /*30872*/;
assign _9525_ = _9526_ | _9528_ /*30870*/;
assign _9284_ = _9520_ ^ _9527_ /*30873*/;
assign _9534_ = D[45] ^ Q[40] /*30869*/;
assign _9531_ = _8899_ & _9534_ /*30865*/;
assign _9532_ = _8899_ ^ _9534_ /*30868*/;
assign _9533_ = _9525_ & _9532_ /*30866*/;
assign _9530_ = _9531_ | _9533_ /*30864*/;
assign _9285_ = _9525_ ^ _9532_ /*30867*/;
assign _9539_ = D[46] ^ Q[40] /*30863*/;
assign _9536_ = _8900_ & _9539_ /*30859*/;
assign _9537_ = _8900_ ^ _9539_ /*30862*/;
assign _9538_ = _9530_ & _9537_ /*30860*/;
assign _9535_ = _9536_ | _9538_ /*30858*/;
assign _9286_ = _9530_ ^ _9537_ /*30861*/;
assign _9544_ = D[47] ^ Q[40] /*30857*/;
assign _9541_ = _8901_ & _9544_ /*30853*/;
assign _9542_ = _8901_ ^ _9544_ /*30856*/;
assign _9543_ = _9535_ & _9542_ /*30854*/;
assign _9540_ = _9541_ | _9543_ /*30852*/;
assign _9287_ = _9535_ ^ _9542_ /*30855*/;
assign _9549_ = D[48] ^ Q[40] /*30851*/;
assign _9546_ = _8902_ & _9549_ /*30847*/;
assign _9547_ = _8902_ ^ _9549_ /*30850*/;
assign _9548_ = _9540_ & _9547_ /*30848*/;
assign _9545_ = _9546_ | _9548_ /*30846*/;
assign _9288_ = _9540_ ^ _9547_ /*30849*/;
assign _9554_ = D[49] ^ Q[40] /*30845*/;
assign _9551_ = _8903_ & _9554_ /*30841*/;
assign _9552_ = _8903_ ^ _9554_ /*30844*/;
assign _9553_ = _9545_ & _9552_ /*30842*/;
assign _9550_ = _9551_ | _9553_ /*30840*/;
assign _9289_ = _9545_ ^ _9552_ /*30843*/;
assign _9559_ = D[50] ^ Q[40] /*30839*/;
assign _9556_ = _8904_ & _9559_ /*30835*/;
assign _9557_ = _8904_ ^ _9559_ /*30838*/;
assign _9558_ = _9550_ & _9557_ /*30836*/;
assign _9555_ = _9556_ | _9558_ /*30834*/;
assign _9290_ = _9550_ ^ _9557_ /*30837*/;
assign _9564_ = D[51] ^ Q[40] /*30833*/;
assign _9561_ = _8905_ & _9564_ /*30829*/;
assign _9562_ = _8905_ ^ _9564_ /*30832*/;
assign _9563_ = _9555_ & _9562_ /*30830*/;
assign _9560_ = _9561_ | _9563_ /*30828*/;
assign _9291_ = _9555_ ^ _9562_ /*30831*/;
assign _9569_ = D[52] ^ Q[40] /*30827*/;
assign _9566_ = _8906_ & _9569_ /*30823*/;
assign _9567_ = _8906_ ^ _9569_ /*30826*/;
assign _9568_ = _9560_ & _9567_ /*30824*/;
assign _9565_ = _9566_ | _9568_ /*30822*/;
assign _9292_ = _9560_ ^ _9567_ /*30825*/;
assign _9574_ = D[53] ^ Q[40] /*30821*/;
assign _9571_ = _8907_ & _9574_ /*30817*/;
assign _9572_ = _8907_ ^ _9574_ /*30820*/;
assign _9573_ = _9565_ & _9572_ /*30818*/;
assign _9570_ = _9571_ | _9573_ /*30816*/;
assign _9293_ = _9565_ ^ _9572_ /*30819*/;
assign _9579_ = D[54] ^ Q[40] /*30815*/;
assign _9576_ = _8908_ & _9579_ /*30811*/;
assign _9577_ = _8908_ ^ _9579_ /*30814*/;
assign _9578_ = _9570_ & _9577_ /*30812*/;
assign _9575_ = _9576_ | _9578_ /*30810*/;
assign _9294_ = _9570_ ^ _9577_ /*30813*/;
assign _9584_ = D[55] ^ Q[40] /*30809*/;
assign _9581_ = _8909_ & _9584_ /*30805*/;
assign _9582_ = _8909_ ^ _9584_ /*30808*/;
assign _9583_ = _9575_ & _9582_ /*30806*/;
assign _9580_ = _9581_ | _9583_ /*30804*/;
assign _9295_ = _9575_ ^ _9582_ /*30807*/;
assign _9589_ = D[56] ^ Q[40] /*30803*/;
assign _9586_ = _8910_ & _9589_ /*30799*/;
assign _9587_ = _8910_ ^ _9589_ /*30802*/;
assign _9588_ = _9580_ & _9587_ /*30800*/;
assign _9585_ = _9586_ | _9588_ /*30798*/;
assign _9296_ = _9580_ ^ _9587_ /*30801*/;
assign _9594_ = D[57] ^ Q[40] /*30797*/;
assign _9591_ = _8911_ & _9594_ /*30793*/;
assign _9592_ = _8911_ ^ _9594_ /*30796*/;
assign _9593_ = _9585_ & _9592_ /*30794*/;
assign _9590_ = _9591_ | _9593_ /*30792*/;
assign _9297_ = _9585_ ^ _9592_ /*30795*/;
assign _9599_ = D[58] ^ Q[40] /*30791*/;
assign _9596_ = _8912_ & _9599_ /*30787*/;
assign _9597_ = _8912_ ^ _9599_ /*30790*/;
assign _9598_ = _9590_ & _9597_ /*30788*/;
assign _9595_ = _9596_ | _9598_ /*30786*/;
assign _9298_ = _9590_ ^ _9597_ /*30789*/;
assign _9604_ = D[59] ^ Q[40] /*30785*/;
assign _9601_ = _8913_ & _9604_ /*30781*/;
assign _9602_ = _8913_ ^ _9604_ /*30784*/;
assign _9603_ = _9595_ & _9602_ /*30782*/;
assign _9600_ = _9601_ | _9603_ /*30780*/;
assign _9299_ = _9595_ ^ _9602_ /*30783*/;
assign _9609_ = D[60] ^ Q[40] /*30779*/;
assign _9606_ = _8914_ & _9609_ /*30775*/;
assign _9607_ = _8914_ ^ _9609_ /*30778*/;
assign _9608_ = _9600_ & _9607_ /*30776*/;
assign _9605_ = _9606_ | _9608_ /*30774*/;
assign _9300_ = _9600_ ^ _9607_ /*30777*/;
assign _9614_ = D[61] ^ Q[40] /*30773*/;
assign _9611_ = _8915_ & _9614_ /*30769*/;
assign _9612_ = _8915_ ^ _9614_ /*30772*/;
assign _9613_ = _9605_ & _9612_ /*30770*/;
assign _9610_ = _9611_ | _9613_ /*30768*/;
assign _9301_ = _9605_ ^ _9612_ /*30771*/;
assign _9619_ = D[62] ^ Q[40] /*30767*/;
assign _9616_ = _8916_ & _9619_ /*30763*/;
assign _9617_ = _8916_ ^ _9619_ /*30766*/;
assign _9618_ = _9610_ & _9617_ /*30764*/;
assign _9615_ = _9616_ | _9618_ /*30762*/;
assign _9302_ = _9610_ ^ _9617_ /*30765*/;
assign _9623_ = zeroWire ^ Q[40] /*30761*/;
assign _9620_ = _8917_ & _9623_ /*30757*/;
assign _9621_ = _8917_ ^ _9623_ /*30760*/;
assign _9622_ = _9615_ & _9621_ /*30758*/;
assign Q[39] = _9620_ | _9622_ /*30756*/;
assign _9303_ = _9615_ ^ _9621_ /*30759*/;
assign _9694_ = D[0] ^ Q[39] /*30370*/;
assign _9691_ = R_0[38] & _9694_ /*30366*/;
assign _9692_ = R_0[38] ^ _9694_ /*30369*/;
assign _9693_ = Q[39] & _9692_ /*30367*/;
assign _9690_ = _9691_ | _9693_ /*30365*/;
assign _9625_ = Q[39] ^ _9692_ /*30368*/;
assign _9699_ = D[1] ^ Q[39] /*30364*/;
assign _9696_ = _9240_ & _9699_ /*30360*/;
assign _9697_ = _9240_ ^ _9699_ /*30363*/;
assign _9698_ = _9690_ & _9697_ /*30361*/;
assign _9695_ = _9696_ | _9698_ /*30359*/;
assign _9626_ = _9690_ ^ _9697_ /*30362*/;
assign _9704_ = D[2] ^ Q[39] /*30358*/;
assign _9701_ = _9241_ & _9704_ /*30354*/;
assign _9702_ = _9241_ ^ _9704_ /*30357*/;
assign _9703_ = _9695_ & _9702_ /*30355*/;
assign _9700_ = _9701_ | _9703_ /*30353*/;
assign _9627_ = _9695_ ^ _9702_ /*30356*/;
assign _9709_ = D[3] ^ Q[39] /*30352*/;
assign _9706_ = _9242_ & _9709_ /*30348*/;
assign _9707_ = _9242_ ^ _9709_ /*30351*/;
assign _9708_ = _9700_ & _9707_ /*30349*/;
assign _9705_ = _9706_ | _9708_ /*30347*/;
assign _9628_ = _9700_ ^ _9707_ /*30350*/;
assign _9714_ = D[4] ^ Q[39] /*30346*/;
assign _9711_ = _9243_ & _9714_ /*30342*/;
assign _9712_ = _9243_ ^ _9714_ /*30345*/;
assign _9713_ = _9705_ & _9712_ /*30343*/;
assign _9710_ = _9711_ | _9713_ /*30341*/;
assign _9629_ = _9705_ ^ _9712_ /*30344*/;
assign _9719_ = D[5] ^ Q[39] /*30340*/;
assign _9716_ = _9244_ & _9719_ /*30336*/;
assign _9717_ = _9244_ ^ _9719_ /*30339*/;
assign _9718_ = _9710_ & _9717_ /*30337*/;
assign _9715_ = _9716_ | _9718_ /*30335*/;
assign _9630_ = _9710_ ^ _9717_ /*30338*/;
assign _9724_ = D[6] ^ Q[39] /*30334*/;
assign _9721_ = _9245_ & _9724_ /*30330*/;
assign _9722_ = _9245_ ^ _9724_ /*30333*/;
assign _9723_ = _9715_ & _9722_ /*30331*/;
assign _9720_ = _9721_ | _9723_ /*30329*/;
assign _9631_ = _9715_ ^ _9722_ /*30332*/;
assign _9729_ = D[7] ^ Q[39] /*30328*/;
assign _9726_ = _9246_ & _9729_ /*30324*/;
assign _9727_ = _9246_ ^ _9729_ /*30327*/;
assign _9728_ = _9720_ & _9727_ /*30325*/;
assign _9725_ = _9726_ | _9728_ /*30323*/;
assign _9632_ = _9720_ ^ _9727_ /*30326*/;
assign _9734_ = D[8] ^ Q[39] /*30322*/;
assign _9731_ = _9247_ & _9734_ /*30318*/;
assign _9732_ = _9247_ ^ _9734_ /*30321*/;
assign _9733_ = _9725_ & _9732_ /*30319*/;
assign _9730_ = _9731_ | _9733_ /*30317*/;
assign _9633_ = _9725_ ^ _9732_ /*30320*/;
assign _9739_ = D[9] ^ Q[39] /*30316*/;
assign _9736_ = _9248_ & _9739_ /*30312*/;
assign _9737_ = _9248_ ^ _9739_ /*30315*/;
assign _9738_ = _9730_ & _9737_ /*30313*/;
assign _9735_ = _9736_ | _9738_ /*30311*/;
assign _9634_ = _9730_ ^ _9737_ /*30314*/;
assign _9744_ = D[10] ^ Q[39] /*30310*/;
assign _9741_ = _9249_ & _9744_ /*30306*/;
assign _9742_ = _9249_ ^ _9744_ /*30309*/;
assign _9743_ = _9735_ & _9742_ /*30307*/;
assign _9740_ = _9741_ | _9743_ /*30305*/;
assign _9635_ = _9735_ ^ _9742_ /*30308*/;
assign _9749_ = D[11] ^ Q[39] /*30304*/;
assign _9746_ = _9250_ & _9749_ /*30300*/;
assign _9747_ = _9250_ ^ _9749_ /*30303*/;
assign _9748_ = _9740_ & _9747_ /*30301*/;
assign _9745_ = _9746_ | _9748_ /*30299*/;
assign _9636_ = _9740_ ^ _9747_ /*30302*/;
assign _9754_ = D[12] ^ Q[39] /*30298*/;
assign _9751_ = _9251_ & _9754_ /*30294*/;
assign _9752_ = _9251_ ^ _9754_ /*30297*/;
assign _9753_ = _9745_ & _9752_ /*30295*/;
assign _9750_ = _9751_ | _9753_ /*30293*/;
assign _9637_ = _9745_ ^ _9752_ /*30296*/;
assign _9759_ = D[13] ^ Q[39] /*30292*/;
assign _9756_ = _9252_ & _9759_ /*30288*/;
assign _9757_ = _9252_ ^ _9759_ /*30291*/;
assign _9758_ = _9750_ & _9757_ /*30289*/;
assign _9755_ = _9756_ | _9758_ /*30287*/;
assign _9638_ = _9750_ ^ _9757_ /*30290*/;
assign _9764_ = D[14] ^ Q[39] /*30286*/;
assign _9761_ = _9253_ & _9764_ /*30282*/;
assign _9762_ = _9253_ ^ _9764_ /*30285*/;
assign _9763_ = _9755_ & _9762_ /*30283*/;
assign _9760_ = _9761_ | _9763_ /*30281*/;
assign _9639_ = _9755_ ^ _9762_ /*30284*/;
assign _9769_ = D[15] ^ Q[39] /*30280*/;
assign _9766_ = _9254_ & _9769_ /*30276*/;
assign _9767_ = _9254_ ^ _9769_ /*30279*/;
assign _9768_ = _9760_ & _9767_ /*30277*/;
assign _9765_ = _9766_ | _9768_ /*30275*/;
assign _9640_ = _9760_ ^ _9767_ /*30278*/;
assign _9774_ = D[16] ^ Q[39] /*30274*/;
assign _9771_ = _9255_ & _9774_ /*30270*/;
assign _9772_ = _9255_ ^ _9774_ /*30273*/;
assign _9773_ = _9765_ & _9772_ /*30271*/;
assign _9770_ = _9771_ | _9773_ /*30269*/;
assign _9641_ = _9765_ ^ _9772_ /*30272*/;
assign _9779_ = D[17] ^ Q[39] /*30268*/;
assign _9776_ = _9256_ & _9779_ /*30264*/;
assign _9777_ = _9256_ ^ _9779_ /*30267*/;
assign _9778_ = _9770_ & _9777_ /*30265*/;
assign _9775_ = _9776_ | _9778_ /*30263*/;
assign _9642_ = _9770_ ^ _9777_ /*30266*/;
assign _9784_ = D[18] ^ Q[39] /*30262*/;
assign _9781_ = _9257_ & _9784_ /*30258*/;
assign _9782_ = _9257_ ^ _9784_ /*30261*/;
assign _9783_ = _9775_ & _9782_ /*30259*/;
assign _9780_ = _9781_ | _9783_ /*30257*/;
assign _9643_ = _9775_ ^ _9782_ /*30260*/;
assign _9789_ = D[19] ^ Q[39] /*30256*/;
assign _9786_ = _9258_ & _9789_ /*30252*/;
assign _9787_ = _9258_ ^ _9789_ /*30255*/;
assign _9788_ = _9780_ & _9787_ /*30253*/;
assign _9785_ = _9786_ | _9788_ /*30251*/;
assign _9644_ = _9780_ ^ _9787_ /*30254*/;
assign _9794_ = D[20] ^ Q[39] /*30250*/;
assign _9791_ = _9259_ & _9794_ /*30246*/;
assign _9792_ = _9259_ ^ _9794_ /*30249*/;
assign _9793_ = _9785_ & _9792_ /*30247*/;
assign _9790_ = _9791_ | _9793_ /*30245*/;
assign _9645_ = _9785_ ^ _9792_ /*30248*/;
assign _9799_ = D[21] ^ Q[39] /*30244*/;
assign _9796_ = _9260_ & _9799_ /*30240*/;
assign _9797_ = _9260_ ^ _9799_ /*30243*/;
assign _9798_ = _9790_ & _9797_ /*30241*/;
assign _9795_ = _9796_ | _9798_ /*30239*/;
assign _9646_ = _9790_ ^ _9797_ /*30242*/;
assign _9804_ = D[22] ^ Q[39] /*30238*/;
assign _9801_ = _9261_ & _9804_ /*30234*/;
assign _9802_ = _9261_ ^ _9804_ /*30237*/;
assign _9803_ = _9795_ & _9802_ /*30235*/;
assign _9800_ = _9801_ | _9803_ /*30233*/;
assign _9647_ = _9795_ ^ _9802_ /*30236*/;
assign _9809_ = D[23] ^ Q[39] /*30232*/;
assign _9806_ = _9262_ & _9809_ /*30228*/;
assign _9807_ = _9262_ ^ _9809_ /*30231*/;
assign _9808_ = _9800_ & _9807_ /*30229*/;
assign _9805_ = _9806_ | _9808_ /*30227*/;
assign _9648_ = _9800_ ^ _9807_ /*30230*/;
assign _9814_ = D[24] ^ Q[39] /*30226*/;
assign _9811_ = _9263_ & _9814_ /*30222*/;
assign _9812_ = _9263_ ^ _9814_ /*30225*/;
assign _9813_ = _9805_ & _9812_ /*30223*/;
assign _9810_ = _9811_ | _9813_ /*30221*/;
assign _9649_ = _9805_ ^ _9812_ /*30224*/;
assign _9819_ = D[25] ^ Q[39] /*30220*/;
assign _9816_ = _9264_ & _9819_ /*30216*/;
assign _9817_ = _9264_ ^ _9819_ /*30219*/;
assign _9818_ = _9810_ & _9817_ /*30217*/;
assign _9815_ = _9816_ | _9818_ /*30215*/;
assign _9650_ = _9810_ ^ _9817_ /*30218*/;
assign _9824_ = D[26] ^ Q[39] /*30214*/;
assign _9821_ = _9265_ & _9824_ /*30210*/;
assign _9822_ = _9265_ ^ _9824_ /*30213*/;
assign _9823_ = _9815_ & _9822_ /*30211*/;
assign _9820_ = _9821_ | _9823_ /*30209*/;
assign _9651_ = _9815_ ^ _9822_ /*30212*/;
assign _9829_ = D[27] ^ Q[39] /*30208*/;
assign _9826_ = _9266_ & _9829_ /*30204*/;
assign _9827_ = _9266_ ^ _9829_ /*30207*/;
assign _9828_ = _9820_ & _9827_ /*30205*/;
assign _9825_ = _9826_ | _9828_ /*30203*/;
assign _9652_ = _9820_ ^ _9827_ /*30206*/;
assign _9834_ = D[28] ^ Q[39] /*30202*/;
assign _9831_ = _9267_ & _9834_ /*30198*/;
assign _9832_ = _9267_ ^ _9834_ /*30201*/;
assign _9833_ = _9825_ & _9832_ /*30199*/;
assign _9830_ = _9831_ | _9833_ /*30197*/;
assign _9653_ = _9825_ ^ _9832_ /*30200*/;
assign _9839_ = D[29] ^ Q[39] /*30196*/;
assign _9836_ = _9268_ & _9839_ /*30192*/;
assign _9837_ = _9268_ ^ _9839_ /*30195*/;
assign _9838_ = _9830_ & _9837_ /*30193*/;
assign _9835_ = _9836_ | _9838_ /*30191*/;
assign _9654_ = _9830_ ^ _9837_ /*30194*/;
assign _9844_ = D[30] ^ Q[39] /*30190*/;
assign _9841_ = _9269_ & _9844_ /*30186*/;
assign _9842_ = _9269_ ^ _9844_ /*30189*/;
assign _9843_ = _9835_ & _9842_ /*30187*/;
assign _9840_ = _9841_ | _9843_ /*30185*/;
assign _9655_ = _9835_ ^ _9842_ /*30188*/;
assign _9849_ = D[31] ^ Q[39] /*30184*/;
assign _9846_ = _9270_ & _9849_ /*30180*/;
assign _9847_ = _9270_ ^ _9849_ /*30183*/;
assign _9848_ = _9840_ & _9847_ /*30181*/;
assign _9845_ = _9846_ | _9848_ /*30179*/;
assign _9656_ = _9840_ ^ _9847_ /*30182*/;
assign _9854_ = D[32] ^ Q[39] /*30178*/;
assign _9851_ = _9271_ & _9854_ /*30174*/;
assign _9852_ = _9271_ ^ _9854_ /*30177*/;
assign _9853_ = _9845_ & _9852_ /*30175*/;
assign _9850_ = _9851_ | _9853_ /*30173*/;
assign _9657_ = _9845_ ^ _9852_ /*30176*/;
assign _9859_ = D[33] ^ Q[39] /*30172*/;
assign _9856_ = _9272_ & _9859_ /*30168*/;
assign _9857_ = _9272_ ^ _9859_ /*30171*/;
assign _9858_ = _9850_ & _9857_ /*30169*/;
assign _9855_ = _9856_ | _9858_ /*30167*/;
assign _9658_ = _9850_ ^ _9857_ /*30170*/;
assign _9864_ = D[34] ^ Q[39] /*30166*/;
assign _9861_ = _9273_ & _9864_ /*30162*/;
assign _9862_ = _9273_ ^ _9864_ /*30165*/;
assign _9863_ = _9855_ & _9862_ /*30163*/;
assign _9860_ = _9861_ | _9863_ /*30161*/;
assign _9659_ = _9855_ ^ _9862_ /*30164*/;
assign _9869_ = D[35] ^ Q[39] /*30160*/;
assign _9866_ = _9274_ & _9869_ /*30156*/;
assign _9867_ = _9274_ ^ _9869_ /*30159*/;
assign _9868_ = _9860_ & _9867_ /*30157*/;
assign _9865_ = _9866_ | _9868_ /*30155*/;
assign _9660_ = _9860_ ^ _9867_ /*30158*/;
assign _9874_ = D[36] ^ Q[39] /*30154*/;
assign _9871_ = _9275_ & _9874_ /*30150*/;
assign _9872_ = _9275_ ^ _9874_ /*30153*/;
assign _9873_ = _9865_ & _9872_ /*30151*/;
assign _9870_ = _9871_ | _9873_ /*30149*/;
assign _9661_ = _9865_ ^ _9872_ /*30152*/;
assign _9879_ = D[37] ^ Q[39] /*30148*/;
assign _9876_ = _9276_ & _9879_ /*30144*/;
assign _9877_ = _9276_ ^ _9879_ /*30147*/;
assign _9878_ = _9870_ & _9877_ /*30145*/;
assign _9875_ = _9876_ | _9878_ /*30143*/;
assign _9662_ = _9870_ ^ _9877_ /*30146*/;
assign _9884_ = D[38] ^ Q[39] /*30142*/;
assign _9881_ = _9277_ & _9884_ /*30138*/;
assign _9882_ = _9277_ ^ _9884_ /*30141*/;
assign _9883_ = _9875_ & _9882_ /*30139*/;
assign _9880_ = _9881_ | _9883_ /*30137*/;
assign _9663_ = _9875_ ^ _9882_ /*30140*/;
assign _9889_ = D[39] ^ Q[39] /*30136*/;
assign _9886_ = _9278_ & _9889_ /*30132*/;
assign _9887_ = _9278_ ^ _9889_ /*30135*/;
assign _9888_ = _9880_ & _9887_ /*30133*/;
assign _9885_ = _9886_ | _9888_ /*30131*/;
assign _9664_ = _9880_ ^ _9887_ /*30134*/;
assign _9894_ = D[40] ^ Q[39] /*30130*/;
assign _9891_ = _9279_ & _9894_ /*30126*/;
assign _9892_ = _9279_ ^ _9894_ /*30129*/;
assign _9893_ = _9885_ & _9892_ /*30127*/;
assign _9890_ = _9891_ | _9893_ /*30125*/;
assign _9665_ = _9885_ ^ _9892_ /*30128*/;
assign _9899_ = D[41] ^ Q[39] /*30124*/;
assign _9896_ = _9280_ & _9899_ /*30120*/;
assign _9897_ = _9280_ ^ _9899_ /*30123*/;
assign _9898_ = _9890_ & _9897_ /*30121*/;
assign _9895_ = _9896_ | _9898_ /*30119*/;
assign _9666_ = _9890_ ^ _9897_ /*30122*/;
assign _9904_ = D[42] ^ Q[39] /*30118*/;
assign _9901_ = _9281_ & _9904_ /*30114*/;
assign _9902_ = _9281_ ^ _9904_ /*30117*/;
assign _9903_ = _9895_ & _9902_ /*30115*/;
assign _9900_ = _9901_ | _9903_ /*30113*/;
assign _9667_ = _9895_ ^ _9902_ /*30116*/;
assign _9909_ = D[43] ^ Q[39] /*30112*/;
assign _9906_ = _9282_ & _9909_ /*30108*/;
assign _9907_ = _9282_ ^ _9909_ /*30111*/;
assign _9908_ = _9900_ & _9907_ /*30109*/;
assign _9905_ = _9906_ | _9908_ /*30107*/;
assign _9668_ = _9900_ ^ _9907_ /*30110*/;
assign _9914_ = D[44] ^ Q[39] /*30106*/;
assign _9911_ = _9283_ & _9914_ /*30102*/;
assign _9912_ = _9283_ ^ _9914_ /*30105*/;
assign _9913_ = _9905_ & _9912_ /*30103*/;
assign _9910_ = _9911_ | _9913_ /*30101*/;
assign _9669_ = _9905_ ^ _9912_ /*30104*/;
assign _9919_ = D[45] ^ Q[39] /*30100*/;
assign _9916_ = _9284_ & _9919_ /*30096*/;
assign _9917_ = _9284_ ^ _9919_ /*30099*/;
assign _9918_ = _9910_ & _9917_ /*30097*/;
assign _9915_ = _9916_ | _9918_ /*30095*/;
assign _9670_ = _9910_ ^ _9917_ /*30098*/;
assign _9924_ = D[46] ^ Q[39] /*30094*/;
assign _9921_ = _9285_ & _9924_ /*30090*/;
assign _9922_ = _9285_ ^ _9924_ /*30093*/;
assign _9923_ = _9915_ & _9922_ /*30091*/;
assign _9920_ = _9921_ | _9923_ /*30089*/;
assign _9671_ = _9915_ ^ _9922_ /*30092*/;
assign _9929_ = D[47] ^ Q[39] /*30088*/;
assign _9926_ = _9286_ & _9929_ /*30084*/;
assign _9927_ = _9286_ ^ _9929_ /*30087*/;
assign _9928_ = _9920_ & _9927_ /*30085*/;
assign _9925_ = _9926_ | _9928_ /*30083*/;
assign _9672_ = _9920_ ^ _9927_ /*30086*/;
assign _9934_ = D[48] ^ Q[39] /*30082*/;
assign _9931_ = _9287_ & _9934_ /*30078*/;
assign _9932_ = _9287_ ^ _9934_ /*30081*/;
assign _9933_ = _9925_ & _9932_ /*30079*/;
assign _9930_ = _9931_ | _9933_ /*30077*/;
assign _9673_ = _9925_ ^ _9932_ /*30080*/;
assign _9939_ = D[49] ^ Q[39] /*30076*/;
assign _9936_ = _9288_ & _9939_ /*30072*/;
assign _9937_ = _9288_ ^ _9939_ /*30075*/;
assign _9938_ = _9930_ & _9937_ /*30073*/;
assign _9935_ = _9936_ | _9938_ /*30071*/;
assign _9674_ = _9930_ ^ _9937_ /*30074*/;
assign _9944_ = D[50] ^ Q[39] /*30070*/;
assign _9941_ = _9289_ & _9944_ /*30066*/;
assign _9942_ = _9289_ ^ _9944_ /*30069*/;
assign _9943_ = _9935_ & _9942_ /*30067*/;
assign _9940_ = _9941_ | _9943_ /*30065*/;
assign _9675_ = _9935_ ^ _9942_ /*30068*/;
assign _9949_ = D[51] ^ Q[39] /*30064*/;
assign _9946_ = _9290_ & _9949_ /*30060*/;
assign _9947_ = _9290_ ^ _9949_ /*30063*/;
assign _9948_ = _9940_ & _9947_ /*30061*/;
assign _9945_ = _9946_ | _9948_ /*30059*/;
assign _9676_ = _9940_ ^ _9947_ /*30062*/;
assign _9954_ = D[52] ^ Q[39] /*30058*/;
assign _9951_ = _9291_ & _9954_ /*30054*/;
assign _9952_ = _9291_ ^ _9954_ /*30057*/;
assign _9953_ = _9945_ & _9952_ /*30055*/;
assign _9950_ = _9951_ | _9953_ /*30053*/;
assign _9677_ = _9945_ ^ _9952_ /*30056*/;
assign _9959_ = D[53] ^ Q[39] /*30052*/;
assign _9956_ = _9292_ & _9959_ /*30048*/;
assign _9957_ = _9292_ ^ _9959_ /*30051*/;
assign _9958_ = _9950_ & _9957_ /*30049*/;
assign _9955_ = _9956_ | _9958_ /*30047*/;
assign _9678_ = _9950_ ^ _9957_ /*30050*/;
assign _9964_ = D[54] ^ Q[39] /*30046*/;
assign _9961_ = _9293_ & _9964_ /*30042*/;
assign _9962_ = _9293_ ^ _9964_ /*30045*/;
assign _9963_ = _9955_ & _9962_ /*30043*/;
assign _9960_ = _9961_ | _9963_ /*30041*/;
assign _9679_ = _9955_ ^ _9962_ /*30044*/;
assign _9969_ = D[55] ^ Q[39] /*30040*/;
assign _9966_ = _9294_ & _9969_ /*30036*/;
assign _9967_ = _9294_ ^ _9969_ /*30039*/;
assign _9968_ = _9960_ & _9967_ /*30037*/;
assign _9965_ = _9966_ | _9968_ /*30035*/;
assign _9680_ = _9960_ ^ _9967_ /*30038*/;
assign _9974_ = D[56] ^ Q[39] /*30034*/;
assign _9971_ = _9295_ & _9974_ /*30030*/;
assign _9972_ = _9295_ ^ _9974_ /*30033*/;
assign _9973_ = _9965_ & _9972_ /*30031*/;
assign _9970_ = _9971_ | _9973_ /*30029*/;
assign _9681_ = _9965_ ^ _9972_ /*30032*/;
assign _9979_ = D[57] ^ Q[39] /*30028*/;
assign _9976_ = _9296_ & _9979_ /*30024*/;
assign _9977_ = _9296_ ^ _9979_ /*30027*/;
assign _9978_ = _9970_ & _9977_ /*30025*/;
assign _9975_ = _9976_ | _9978_ /*30023*/;
assign _9682_ = _9970_ ^ _9977_ /*30026*/;
assign _9984_ = D[58] ^ Q[39] /*30022*/;
assign _9981_ = _9297_ & _9984_ /*30018*/;
assign _9982_ = _9297_ ^ _9984_ /*30021*/;
assign _9983_ = _9975_ & _9982_ /*30019*/;
assign _9980_ = _9981_ | _9983_ /*30017*/;
assign _9683_ = _9975_ ^ _9982_ /*30020*/;
assign _9989_ = D[59] ^ Q[39] /*30016*/;
assign _9986_ = _9298_ & _9989_ /*30012*/;
assign _9987_ = _9298_ ^ _9989_ /*30015*/;
assign _9988_ = _9980_ & _9987_ /*30013*/;
assign _9985_ = _9986_ | _9988_ /*30011*/;
assign _9684_ = _9980_ ^ _9987_ /*30014*/;
assign _9994_ = D[60] ^ Q[39] /*30010*/;
assign _9991_ = _9299_ & _9994_ /*30006*/;
assign _9992_ = _9299_ ^ _9994_ /*30009*/;
assign _9993_ = _9985_ & _9992_ /*30007*/;
assign _9990_ = _9991_ | _9993_ /*30005*/;
assign _9685_ = _9985_ ^ _9992_ /*30008*/;
assign _9999_ = D[61] ^ Q[39] /*30004*/;
assign _9996_ = _9300_ & _9999_ /*30000*/;
assign _9997_ = _9300_ ^ _9999_ /*30003*/;
assign _9998_ = _9990_ & _9997_ /*30001*/;
assign _9995_ = _9996_ | _9998_ /*29999*/;
assign _9686_ = _9990_ ^ _9997_ /*30002*/;
assign _10004_ = D[62] ^ Q[39] /*29998*/;
assign _10001_ = _9301_ & _10004_ /*29994*/;
assign _10002_ = _9301_ ^ _10004_ /*29997*/;
assign _10003_ = _9995_ & _10002_ /*29995*/;
assign _10000_ = _10001_ | _10003_ /*29993*/;
assign _9687_ = _9995_ ^ _10002_ /*29996*/;
assign _10008_ = zeroWire ^ Q[39] /*29992*/;
assign _10005_ = _9302_ & _10008_ /*29988*/;
assign _10006_ = _9302_ ^ _10008_ /*29991*/;
assign _10007_ = _10000_ & _10006_ /*29989*/;
assign Q[38] = _10005_ | _10007_ /*29987*/;
assign _9688_ = _10000_ ^ _10006_ /*29990*/;
assign _10079_ = D[0] ^ Q[38] /*29601*/;
assign _10076_ = R_0[37] & _10079_ /*29597*/;
assign _10077_ = R_0[37] ^ _10079_ /*29600*/;
assign _10078_ = Q[38] & _10077_ /*29598*/;
assign _10075_ = _10076_ | _10078_ /*29596*/;
assign _10010_ = Q[38] ^ _10077_ /*29599*/;
assign _10084_ = D[1] ^ Q[38] /*29595*/;
assign _10081_ = _9625_ & _10084_ /*29591*/;
assign _10082_ = _9625_ ^ _10084_ /*29594*/;
assign _10083_ = _10075_ & _10082_ /*29592*/;
assign _10080_ = _10081_ | _10083_ /*29590*/;
assign _10011_ = _10075_ ^ _10082_ /*29593*/;
assign _10089_ = D[2] ^ Q[38] /*29589*/;
assign _10086_ = _9626_ & _10089_ /*29585*/;
assign _10087_ = _9626_ ^ _10089_ /*29588*/;
assign _10088_ = _10080_ & _10087_ /*29586*/;
assign _10085_ = _10086_ | _10088_ /*29584*/;
assign _10012_ = _10080_ ^ _10087_ /*29587*/;
assign _10094_ = D[3] ^ Q[38] /*29583*/;
assign _10091_ = _9627_ & _10094_ /*29579*/;
assign _10092_ = _9627_ ^ _10094_ /*29582*/;
assign _10093_ = _10085_ & _10092_ /*29580*/;
assign _10090_ = _10091_ | _10093_ /*29578*/;
assign _10013_ = _10085_ ^ _10092_ /*29581*/;
assign _10099_ = D[4] ^ Q[38] /*29577*/;
assign _10096_ = _9628_ & _10099_ /*29573*/;
assign _10097_ = _9628_ ^ _10099_ /*29576*/;
assign _10098_ = _10090_ & _10097_ /*29574*/;
assign _10095_ = _10096_ | _10098_ /*29572*/;
assign _10014_ = _10090_ ^ _10097_ /*29575*/;
assign _10104_ = D[5] ^ Q[38] /*29571*/;
assign _10101_ = _9629_ & _10104_ /*29567*/;
assign _10102_ = _9629_ ^ _10104_ /*29570*/;
assign _10103_ = _10095_ & _10102_ /*29568*/;
assign _10100_ = _10101_ | _10103_ /*29566*/;
assign _10015_ = _10095_ ^ _10102_ /*29569*/;
assign _10109_ = D[6] ^ Q[38] /*29565*/;
assign _10106_ = _9630_ & _10109_ /*29561*/;
assign _10107_ = _9630_ ^ _10109_ /*29564*/;
assign _10108_ = _10100_ & _10107_ /*29562*/;
assign _10105_ = _10106_ | _10108_ /*29560*/;
assign _10016_ = _10100_ ^ _10107_ /*29563*/;
assign _10114_ = D[7] ^ Q[38] /*29559*/;
assign _10111_ = _9631_ & _10114_ /*29555*/;
assign _10112_ = _9631_ ^ _10114_ /*29558*/;
assign _10113_ = _10105_ & _10112_ /*29556*/;
assign _10110_ = _10111_ | _10113_ /*29554*/;
assign _10017_ = _10105_ ^ _10112_ /*29557*/;
assign _10119_ = D[8] ^ Q[38] /*29553*/;
assign _10116_ = _9632_ & _10119_ /*29549*/;
assign _10117_ = _9632_ ^ _10119_ /*29552*/;
assign _10118_ = _10110_ & _10117_ /*29550*/;
assign _10115_ = _10116_ | _10118_ /*29548*/;
assign _10018_ = _10110_ ^ _10117_ /*29551*/;
assign _10124_ = D[9] ^ Q[38] /*29547*/;
assign _10121_ = _9633_ & _10124_ /*29543*/;
assign _10122_ = _9633_ ^ _10124_ /*29546*/;
assign _10123_ = _10115_ & _10122_ /*29544*/;
assign _10120_ = _10121_ | _10123_ /*29542*/;
assign _10019_ = _10115_ ^ _10122_ /*29545*/;
assign _10129_ = D[10] ^ Q[38] /*29541*/;
assign _10126_ = _9634_ & _10129_ /*29537*/;
assign _10127_ = _9634_ ^ _10129_ /*29540*/;
assign _10128_ = _10120_ & _10127_ /*29538*/;
assign _10125_ = _10126_ | _10128_ /*29536*/;
assign _10020_ = _10120_ ^ _10127_ /*29539*/;
assign _10134_ = D[11] ^ Q[38] /*29535*/;
assign _10131_ = _9635_ & _10134_ /*29531*/;
assign _10132_ = _9635_ ^ _10134_ /*29534*/;
assign _10133_ = _10125_ & _10132_ /*29532*/;
assign _10130_ = _10131_ | _10133_ /*29530*/;
assign _10021_ = _10125_ ^ _10132_ /*29533*/;
assign _10139_ = D[12] ^ Q[38] /*29529*/;
assign _10136_ = _9636_ & _10139_ /*29525*/;
assign _10137_ = _9636_ ^ _10139_ /*29528*/;
assign _10138_ = _10130_ & _10137_ /*29526*/;
assign _10135_ = _10136_ | _10138_ /*29524*/;
assign _10022_ = _10130_ ^ _10137_ /*29527*/;
assign _10144_ = D[13] ^ Q[38] /*29523*/;
assign _10141_ = _9637_ & _10144_ /*29519*/;
assign _10142_ = _9637_ ^ _10144_ /*29522*/;
assign _10143_ = _10135_ & _10142_ /*29520*/;
assign _10140_ = _10141_ | _10143_ /*29518*/;
assign _10023_ = _10135_ ^ _10142_ /*29521*/;
assign _10149_ = D[14] ^ Q[38] /*29517*/;
assign _10146_ = _9638_ & _10149_ /*29513*/;
assign _10147_ = _9638_ ^ _10149_ /*29516*/;
assign _10148_ = _10140_ & _10147_ /*29514*/;
assign _10145_ = _10146_ | _10148_ /*29512*/;
assign _10024_ = _10140_ ^ _10147_ /*29515*/;
assign _10154_ = D[15] ^ Q[38] /*29511*/;
assign _10151_ = _9639_ & _10154_ /*29507*/;
assign _10152_ = _9639_ ^ _10154_ /*29510*/;
assign _10153_ = _10145_ & _10152_ /*29508*/;
assign _10150_ = _10151_ | _10153_ /*29506*/;
assign _10025_ = _10145_ ^ _10152_ /*29509*/;
assign _10159_ = D[16] ^ Q[38] /*29505*/;
assign _10156_ = _9640_ & _10159_ /*29501*/;
assign _10157_ = _9640_ ^ _10159_ /*29504*/;
assign _10158_ = _10150_ & _10157_ /*29502*/;
assign _10155_ = _10156_ | _10158_ /*29500*/;
assign _10026_ = _10150_ ^ _10157_ /*29503*/;
assign _10164_ = D[17] ^ Q[38] /*29499*/;
assign _10161_ = _9641_ & _10164_ /*29495*/;
assign _10162_ = _9641_ ^ _10164_ /*29498*/;
assign _10163_ = _10155_ & _10162_ /*29496*/;
assign _10160_ = _10161_ | _10163_ /*29494*/;
assign _10027_ = _10155_ ^ _10162_ /*29497*/;
assign _10169_ = D[18] ^ Q[38] /*29493*/;
assign _10166_ = _9642_ & _10169_ /*29489*/;
assign _10167_ = _9642_ ^ _10169_ /*29492*/;
assign _10168_ = _10160_ & _10167_ /*29490*/;
assign _10165_ = _10166_ | _10168_ /*29488*/;
assign _10028_ = _10160_ ^ _10167_ /*29491*/;
assign _10174_ = D[19] ^ Q[38] /*29487*/;
assign _10171_ = _9643_ & _10174_ /*29483*/;
assign _10172_ = _9643_ ^ _10174_ /*29486*/;
assign _10173_ = _10165_ & _10172_ /*29484*/;
assign _10170_ = _10171_ | _10173_ /*29482*/;
assign _10029_ = _10165_ ^ _10172_ /*29485*/;
assign _10179_ = D[20] ^ Q[38] /*29481*/;
assign _10176_ = _9644_ & _10179_ /*29477*/;
assign _10177_ = _9644_ ^ _10179_ /*29480*/;
assign _10178_ = _10170_ & _10177_ /*29478*/;
assign _10175_ = _10176_ | _10178_ /*29476*/;
assign _10030_ = _10170_ ^ _10177_ /*29479*/;
assign _10184_ = D[21] ^ Q[38] /*29475*/;
assign _10181_ = _9645_ & _10184_ /*29471*/;
assign _10182_ = _9645_ ^ _10184_ /*29474*/;
assign _10183_ = _10175_ & _10182_ /*29472*/;
assign _10180_ = _10181_ | _10183_ /*29470*/;
assign _10031_ = _10175_ ^ _10182_ /*29473*/;
assign _10189_ = D[22] ^ Q[38] /*29469*/;
assign _10186_ = _9646_ & _10189_ /*29465*/;
assign _10187_ = _9646_ ^ _10189_ /*29468*/;
assign _10188_ = _10180_ & _10187_ /*29466*/;
assign _10185_ = _10186_ | _10188_ /*29464*/;
assign _10032_ = _10180_ ^ _10187_ /*29467*/;
assign _10194_ = D[23] ^ Q[38] /*29463*/;
assign _10191_ = _9647_ & _10194_ /*29459*/;
assign _10192_ = _9647_ ^ _10194_ /*29462*/;
assign _10193_ = _10185_ & _10192_ /*29460*/;
assign _10190_ = _10191_ | _10193_ /*29458*/;
assign _10033_ = _10185_ ^ _10192_ /*29461*/;
assign _10199_ = D[24] ^ Q[38] /*29457*/;
assign _10196_ = _9648_ & _10199_ /*29453*/;
assign _10197_ = _9648_ ^ _10199_ /*29456*/;
assign _10198_ = _10190_ & _10197_ /*29454*/;
assign _10195_ = _10196_ | _10198_ /*29452*/;
assign _10034_ = _10190_ ^ _10197_ /*29455*/;
assign _10204_ = D[25] ^ Q[38] /*29451*/;
assign _10201_ = _9649_ & _10204_ /*29447*/;
assign _10202_ = _9649_ ^ _10204_ /*29450*/;
assign _10203_ = _10195_ & _10202_ /*29448*/;
assign _10200_ = _10201_ | _10203_ /*29446*/;
assign _10035_ = _10195_ ^ _10202_ /*29449*/;
assign _10209_ = D[26] ^ Q[38] /*29445*/;
assign _10206_ = _9650_ & _10209_ /*29441*/;
assign _10207_ = _9650_ ^ _10209_ /*29444*/;
assign _10208_ = _10200_ & _10207_ /*29442*/;
assign _10205_ = _10206_ | _10208_ /*29440*/;
assign _10036_ = _10200_ ^ _10207_ /*29443*/;
assign _10214_ = D[27] ^ Q[38] /*29439*/;
assign _10211_ = _9651_ & _10214_ /*29435*/;
assign _10212_ = _9651_ ^ _10214_ /*29438*/;
assign _10213_ = _10205_ & _10212_ /*29436*/;
assign _10210_ = _10211_ | _10213_ /*29434*/;
assign _10037_ = _10205_ ^ _10212_ /*29437*/;
assign _10219_ = D[28] ^ Q[38] /*29433*/;
assign _10216_ = _9652_ & _10219_ /*29429*/;
assign _10217_ = _9652_ ^ _10219_ /*29432*/;
assign _10218_ = _10210_ & _10217_ /*29430*/;
assign _10215_ = _10216_ | _10218_ /*29428*/;
assign _10038_ = _10210_ ^ _10217_ /*29431*/;
assign _10224_ = D[29] ^ Q[38] /*29427*/;
assign _10221_ = _9653_ & _10224_ /*29423*/;
assign _10222_ = _9653_ ^ _10224_ /*29426*/;
assign _10223_ = _10215_ & _10222_ /*29424*/;
assign _10220_ = _10221_ | _10223_ /*29422*/;
assign _10039_ = _10215_ ^ _10222_ /*29425*/;
assign _10229_ = D[30] ^ Q[38] /*29421*/;
assign _10226_ = _9654_ & _10229_ /*29417*/;
assign _10227_ = _9654_ ^ _10229_ /*29420*/;
assign _10228_ = _10220_ & _10227_ /*29418*/;
assign _10225_ = _10226_ | _10228_ /*29416*/;
assign _10040_ = _10220_ ^ _10227_ /*29419*/;
assign _10234_ = D[31] ^ Q[38] /*29415*/;
assign _10231_ = _9655_ & _10234_ /*29411*/;
assign _10232_ = _9655_ ^ _10234_ /*29414*/;
assign _10233_ = _10225_ & _10232_ /*29412*/;
assign _10230_ = _10231_ | _10233_ /*29410*/;
assign _10041_ = _10225_ ^ _10232_ /*29413*/;
assign _10239_ = D[32] ^ Q[38] /*29409*/;
assign _10236_ = _9656_ & _10239_ /*29405*/;
assign _10237_ = _9656_ ^ _10239_ /*29408*/;
assign _10238_ = _10230_ & _10237_ /*29406*/;
assign _10235_ = _10236_ | _10238_ /*29404*/;
assign _10042_ = _10230_ ^ _10237_ /*29407*/;
assign _10244_ = D[33] ^ Q[38] /*29403*/;
assign _10241_ = _9657_ & _10244_ /*29399*/;
assign _10242_ = _9657_ ^ _10244_ /*29402*/;
assign _10243_ = _10235_ & _10242_ /*29400*/;
assign _10240_ = _10241_ | _10243_ /*29398*/;
assign _10043_ = _10235_ ^ _10242_ /*29401*/;
assign _10249_ = D[34] ^ Q[38] /*29397*/;
assign _10246_ = _9658_ & _10249_ /*29393*/;
assign _10247_ = _9658_ ^ _10249_ /*29396*/;
assign _10248_ = _10240_ & _10247_ /*29394*/;
assign _10245_ = _10246_ | _10248_ /*29392*/;
assign _10044_ = _10240_ ^ _10247_ /*29395*/;
assign _10254_ = D[35] ^ Q[38] /*29391*/;
assign _10251_ = _9659_ & _10254_ /*29387*/;
assign _10252_ = _9659_ ^ _10254_ /*29390*/;
assign _10253_ = _10245_ & _10252_ /*29388*/;
assign _10250_ = _10251_ | _10253_ /*29386*/;
assign _10045_ = _10245_ ^ _10252_ /*29389*/;
assign _10259_ = D[36] ^ Q[38] /*29385*/;
assign _10256_ = _9660_ & _10259_ /*29381*/;
assign _10257_ = _9660_ ^ _10259_ /*29384*/;
assign _10258_ = _10250_ & _10257_ /*29382*/;
assign _10255_ = _10256_ | _10258_ /*29380*/;
assign _10046_ = _10250_ ^ _10257_ /*29383*/;
assign _10264_ = D[37] ^ Q[38] /*29379*/;
assign _10261_ = _9661_ & _10264_ /*29375*/;
assign _10262_ = _9661_ ^ _10264_ /*29378*/;
assign _10263_ = _10255_ & _10262_ /*29376*/;
assign _10260_ = _10261_ | _10263_ /*29374*/;
assign _10047_ = _10255_ ^ _10262_ /*29377*/;
assign _10269_ = D[38] ^ Q[38] /*29373*/;
assign _10266_ = _9662_ & _10269_ /*29369*/;
assign _10267_ = _9662_ ^ _10269_ /*29372*/;
assign _10268_ = _10260_ & _10267_ /*29370*/;
assign _10265_ = _10266_ | _10268_ /*29368*/;
assign _10048_ = _10260_ ^ _10267_ /*29371*/;
assign _10274_ = D[39] ^ Q[38] /*29367*/;
assign _10271_ = _9663_ & _10274_ /*29363*/;
assign _10272_ = _9663_ ^ _10274_ /*29366*/;
assign _10273_ = _10265_ & _10272_ /*29364*/;
assign _10270_ = _10271_ | _10273_ /*29362*/;
assign _10049_ = _10265_ ^ _10272_ /*29365*/;
assign _10279_ = D[40] ^ Q[38] /*29361*/;
assign _10276_ = _9664_ & _10279_ /*29357*/;
assign _10277_ = _9664_ ^ _10279_ /*29360*/;
assign _10278_ = _10270_ & _10277_ /*29358*/;
assign _10275_ = _10276_ | _10278_ /*29356*/;
assign _10050_ = _10270_ ^ _10277_ /*29359*/;
assign _10284_ = D[41] ^ Q[38] /*29355*/;
assign _10281_ = _9665_ & _10284_ /*29351*/;
assign _10282_ = _9665_ ^ _10284_ /*29354*/;
assign _10283_ = _10275_ & _10282_ /*29352*/;
assign _10280_ = _10281_ | _10283_ /*29350*/;
assign _10051_ = _10275_ ^ _10282_ /*29353*/;
assign _10289_ = D[42] ^ Q[38] /*29349*/;
assign _10286_ = _9666_ & _10289_ /*29345*/;
assign _10287_ = _9666_ ^ _10289_ /*29348*/;
assign _10288_ = _10280_ & _10287_ /*29346*/;
assign _10285_ = _10286_ | _10288_ /*29344*/;
assign _10052_ = _10280_ ^ _10287_ /*29347*/;
assign _10294_ = D[43] ^ Q[38] /*29343*/;
assign _10291_ = _9667_ & _10294_ /*29339*/;
assign _10292_ = _9667_ ^ _10294_ /*29342*/;
assign _10293_ = _10285_ & _10292_ /*29340*/;
assign _10290_ = _10291_ | _10293_ /*29338*/;
assign _10053_ = _10285_ ^ _10292_ /*29341*/;
assign _10299_ = D[44] ^ Q[38] /*29337*/;
assign _10296_ = _9668_ & _10299_ /*29333*/;
assign _10297_ = _9668_ ^ _10299_ /*29336*/;
assign _10298_ = _10290_ & _10297_ /*29334*/;
assign _10295_ = _10296_ | _10298_ /*29332*/;
assign _10054_ = _10290_ ^ _10297_ /*29335*/;
assign _10304_ = D[45] ^ Q[38] /*29331*/;
assign _10301_ = _9669_ & _10304_ /*29327*/;
assign _10302_ = _9669_ ^ _10304_ /*29330*/;
assign _10303_ = _10295_ & _10302_ /*29328*/;
assign _10300_ = _10301_ | _10303_ /*29326*/;
assign _10055_ = _10295_ ^ _10302_ /*29329*/;
assign _10309_ = D[46] ^ Q[38] /*29325*/;
assign _10306_ = _9670_ & _10309_ /*29321*/;
assign _10307_ = _9670_ ^ _10309_ /*29324*/;
assign _10308_ = _10300_ & _10307_ /*29322*/;
assign _10305_ = _10306_ | _10308_ /*29320*/;
assign _10056_ = _10300_ ^ _10307_ /*29323*/;
assign _10314_ = D[47] ^ Q[38] /*29319*/;
assign _10311_ = _9671_ & _10314_ /*29315*/;
assign _10312_ = _9671_ ^ _10314_ /*29318*/;
assign _10313_ = _10305_ & _10312_ /*29316*/;
assign _10310_ = _10311_ | _10313_ /*29314*/;
assign _10057_ = _10305_ ^ _10312_ /*29317*/;
assign _10319_ = D[48] ^ Q[38] /*29313*/;
assign _10316_ = _9672_ & _10319_ /*29309*/;
assign _10317_ = _9672_ ^ _10319_ /*29312*/;
assign _10318_ = _10310_ & _10317_ /*29310*/;
assign _10315_ = _10316_ | _10318_ /*29308*/;
assign _10058_ = _10310_ ^ _10317_ /*29311*/;
assign _10324_ = D[49] ^ Q[38] /*29307*/;
assign _10321_ = _9673_ & _10324_ /*29303*/;
assign _10322_ = _9673_ ^ _10324_ /*29306*/;
assign _10323_ = _10315_ & _10322_ /*29304*/;
assign _10320_ = _10321_ | _10323_ /*29302*/;
assign _10059_ = _10315_ ^ _10322_ /*29305*/;
assign _10329_ = D[50] ^ Q[38] /*29301*/;
assign _10326_ = _9674_ & _10329_ /*29297*/;
assign _10327_ = _9674_ ^ _10329_ /*29300*/;
assign _10328_ = _10320_ & _10327_ /*29298*/;
assign _10325_ = _10326_ | _10328_ /*29296*/;
assign _10060_ = _10320_ ^ _10327_ /*29299*/;
assign _10334_ = D[51] ^ Q[38] /*29295*/;
assign _10331_ = _9675_ & _10334_ /*29291*/;
assign _10332_ = _9675_ ^ _10334_ /*29294*/;
assign _10333_ = _10325_ & _10332_ /*29292*/;
assign _10330_ = _10331_ | _10333_ /*29290*/;
assign _10061_ = _10325_ ^ _10332_ /*29293*/;
assign _10339_ = D[52] ^ Q[38] /*29289*/;
assign _10336_ = _9676_ & _10339_ /*29285*/;
assign _10337_ = _9676_ ^ _10339_ /*29288*/;
assign _10338_ = _10330_ & _10337_ /*29286*/;
assign _10335_ = _10336_ | _10338_ /*29284*/;
assign _10062_ = _10330_ ^ _10337_ /*29287*/;
assign _10344_ = D[53] ^ Q[38] /*29283*/;
assign _10341_ = _9677_ & _10344_ /*29279*/;
assign _10342_ = _9677_ ^ _10344_ /*29282*/;
assign _10343_ = _10335_ & _10342_ /*29280*/;
assign _10340_ = _10341_ | _10343_ /*29278*/;
assign _10063_ = _10335_ ^ _10342_ /*29281*/;
assign _10349_ = D[54] ^ Q[38] /*29277*/;
assign _10346_ = _9678_ & _10349_ /*29273*/;
assign _10347_ = _9678_ ^ _10349_ /*29276*/;
assign _10348_ = _10340_ & _10347_ /*29274*/;
assign _10345_ = _10346_ | _10348_ /*29272*/;
assign _10064_ = _10340_ ^ _10347_ /*29275*/;
assign _10354_ = D[55] ^ Q[38] /*29271*/;
assign _10351_ = _9679_ & _10354_ /*29267*/;
assign _10352_ = _9679_ ^ _10354_ /*29270*/;
assign _10353_ = _10345_ & _10352_ /*29268*/;
assign _10350_ = _10351_ | _10353_ /*29266*/;
assign _10065_ = _10345_ ^ _10352_ /*29269*/;
assign _10359_ = D[56] ^ Q[38] /*29265*/;
assign _10356_ = _9680_ & _10359_ /*29261*/;
assign _10357_ = _9680_ ^ _10359_ /*29264*/;
assign _10358_ = _10350_ & _10357_ /*29262*/;
assign _10355_ = _10356_ | _10358_ /*29260*/;
assign _10066_ = _10350_ ^ _10357_ /*29263*/;
assign _10364_ = D[57] ^ Q[38] /*29259*/;
assign _10361_ = _9681_ & _10364_ /*29255*/;
assign _10362_ = _9681_ ^ _10364_ /*29258*/;
assign _10363_ = _10355_ & _10362_ /*29256*/;
assign _10360_ = _10361_ | _10363_ /*29254*/;
assign _10067_ = _10355_ ^ _10362_ /*29257*/;
assign _10369_ = D[58] ^ Q[38] /*29253*/;
assign _10366_ = _9682_ & _10369_ /*29249*/;
assign _10367_ = _9682_ ^ _10369_ /*29252*/;
assign _10368_ = _10360_ & _10367_ /*29250*/;
assign _10365_ = _10366_ | _10368_ /*29248*/;
assign _10068_ = _10360_ ^ _10367_ /*29251*/;
assign _10374_ = D[59] ^ Q[38] /*29247*/;
assign _10371_ = _9683_ & _10374_ /*29243*/;
assign _10372_ = _9683_ ^ _10374_ /*29246*/;
assign _10373_ = _10365_ & _10372_ /*29244*/;
assign _10370_ = _10371_ | _10373_ /*29242*/;
assign _10069_ = _10365_ ^ _10372_ /*29245*/;
assign _10379_ = D[60] ^ Q[38] /*29241*/;
assign _10376_ = _9684_ & _10379_ /*29237*/;
assign _10377_ = _9684_ ^ _10379_ /*29240*/;
assign _10378_ = _10370_ & _10377_ /*29238*/;
assign _10375_ = _10376_ | _10378_ /*29236*/;
assign _10070_ = _10370_ ^ _10377_ /*29239*/;
assign _10384_ = D[61] ^ Q[38] /*29235*/;
assign _10381_ = _9685_ & _10384_ /*29231*/;
assign _10382_ = _9685_ ^ _10384_ /*29234*/;
assign _10383_ = _10375_ & _10382_ /*29232*/;
assign _10380_ = _10381_ | _10383_ /*29230*/;
assign _10071_ = _10375_ ^ _10382_ /*29233*/;
assign _10389_ = D[62] ^ Q[38] /*29229*/;
assign _10386_ = _9686_ & _10389_ /*29225*/;
assign _10387_ = _9686_ ^ _10389_ /*29228*/;
assign _10388_ = _10380_ & _10387_ /*29226*/;
assign _10385_ = _10386_ | _10388_ /*29224*/;
assign _10072_ = _10380_ ^ _10387_ /*29227*/;
assign _10393_ = zeroWire ^ Q[38] /*29223*/;
assign _10390_ = _9687_ & _10393_ /*29219*/;
assign _10391_ = _9687_ ^ _10393_ /*29222*/;
assign _10392_ = _10385_ & _10391_ /*29220*/;
assign Q[37] = _10390_ | _10392_ /*29218*/;
assign _10073_ = _10385_ ^ _10391_ /*29221*/;
assign _10464_ = D[0] ^ Q[37] /*28832*/;
assign _10461_ = R_0[36] & _10464_ /*28828*/;
assign _10462_ = R_0[36] ^ _10464_ /*28831*/;
assign _10463_ = Q[37] & _10462_ /*28829*/;
assign _10460_ = _10461_ | _10463_ /*28827*/;
assign _10395_ = Q[37] ^ _10462_ /*28830*/;
assign _10469_ = D[1] ^ Q[37] /*28826*/;
assign _10466_ = _10010_ & _10469_ /*28822*/;
assign _10467_ = _10010_ ^ _10469_ /*28825*/;
assign _10468_ = _10460_ & _10467_ /*28823*/;
assign _10465_ = _10466_ | _10468_ /*28821*/;
assign _10396_ = _10460_ ^ _10467_ /*28824*/;
assign _10474_ = D[2] ^ Q[37] /*28820*/;
assign _10471_ = _10011_ & _10474_ /*28816*/;
assign _10472_ = _10011_ ^ _10474_ /*28819*/;
assign _10473_ = _10465_ & _10472_ /*28817*/;
assign _10470_ = _10471_ | _10473_ /*28815*/;
assign _10397_ = _10465_ ^ _10472_ /*28818*/;
assign _10479_ = D[3] ^ Q[37] /*28814*/;
assign _10476_ = _10012_ & _10479_ /*28810*/;
assign _10477_ = _10012_ ^ _10479_ /*28813*/;
assign _10478_ = _10470_ & _10477_ /*28811*/;
assign _10475_ = _10476_ | _10478_ /*28809*/;
assign _10398_ = _10470_ ^ _10477_ /*28812*/;
assign _10484_ = D[4] ^ Q[37] /*28808*/;
assign _10481_ = _10013_ & _10484_ /*28804*/;
assign _10482_ = _10013_ ^ _10484_ /*28807*/;
assign _10483_ = _10475_ & _10482_ /*28805*/;
assign _10480_ = _10481_ | _10483_ /*28803*/;
assign _10399_ = _10475_ ^ _10482_ /*28806*/;
assign _10489_ = D[5] ^ Q[37] /*28802*/;
assign _10486_ = _10014_ & _10489_ /*28798*/;
assign _10487_ = _10014_ ^ _10489_ /*28801*/;
assign _10488_ = _10480_ & _10487_ /*28799*/;
assign _10485_ = _10486_ | _10488_ /*28797*/;
assign _10400_ = _10480_ ^ _10487_ /*28800*/;
assign _10494_ = D[6] ^ Q[37] /*28796*/;
assign _10491_ = _10015_ & _10494_ /*28792*/;
assign _10492_ = _10015_ ^ _10494_ /*28795*/;
assign _10493_ = _10485_ & _10492_ /*28793*/;
assign _10490_ = _10491_ | _10493_ /*28791*/;
assign _10401_ = _10485_ ^ _10492_ /*28794*/;
assign _10499_ = D[7] ^ Q[37] /*28790*/;
assign _10496_ = _10016_ & _10499_ /*28786*/;
assign _10497_ = _10016_ ^ _10499_ /*28789*/;
assign _10498_ = _10490_ & _10497_ /*28787*/;
assign _10495_ = _10496_ | _10498_ /*28785*/;
assign _10402_ = _10490_ ^ _10497_ /*28788*/;
assign _10504_ = D[8] ^ Q[37] /*28784*/;
assign _10501_ = _10017_ & _10504_ /*28780*/;
assign _10502_ = _10017_ ^ _10504_ /*28783*/;
assign _10503_ = _10495_ & _10502_ /*28781*/;
assign _10500_ = _10501_ | _10503_ /*28779*/;
assign _10403_ = _10495_ ^ _10502_ /*28782*/;
assign _10509_ = D[9] ^ Q[37] /*28778*/;
assign _10506_ = _10018_ & _10509_ /*28774*/;
assign _10507_ = _10018_ ^ _10509_ /*28777*/;
assign _10508_ = _10500_ & _10507_ /*28775*/;
assign _10505_ = _10506_ | _10508_ /*28773*/;
assign _10404_ = _10500_ ^ _10507_ /*28776*/;
assign _10514_ = D[10] ^ Q[37] /*28772*/;
assign _10511_ = _10019_ & _10514_ /*28768*/;
assign _10512_ = _10019_ ^ _10514_ /*28771*/;
assign _10513_ = _10505_ & _10512_ /*28769*/;
assign _10510_ = _10511_ | _10513_ /*28767*/;
assign _10405_ = _10505_ ^ _10512_ /*28770*/;
assign _10519_ = D[11] ^ Q[37] /*28766*/;
assign _10516_ = _10020_ & _10519_ /*28762*/;
assign _10517_ = _10020_ ^ _10519_ /*28765*/;
assign _10518_ = _10510_ & _10517_ /*28763*/;
assign _10515_ = _10516_ | _10518_ /*28761*/;
assign _10406_ = _10510_ ^ _10517_ /*28764*/;
assign _10524_ = D[12] ^ Q[37] /*28760*/;
assign _10521_ = _10021_ & _10524_ /*28756*/;
assign _10522_ = _10021_ ^ _10524_ /*28759*/;
assign _10523_ = _10515_ & _10522_ /*28757*/;
assign _10520_ = _10521_ | _10523_ /*28755*/;
assign _10407_ = _10515_ ^ _10522_ /*28758*/;
assign _10529_ = D[13] ^ Q[37] /*28754*/;
assign _10526_ = _10022_ & _10529_ /*28750*/;
assign _10527_ = _10022_ ^ _10529_ /*28753*/;
assign _10528_ = _10520_ & _10527_ /*28751*/;
assign _10525_ = _10526_ | _10528_ /*28749*/;
assign _10408_ = _10520_ ^ _10527_ /*28752*/;
assign _10534_ = D[14] ^ Q[37] /*28748*/;
assign _10531_ = _10023_ & _10534_ /*28744*/;
assign _10532_ = _10023_ ^ _10534_ /*28747*/;
assign _10533_ = _10525_ & _10532_ /*28745*/;
assign _10530_ = _10531_ | _10533_ /*28743*/;
assign _10409_ = _10525_ ^ _10532_ /*28746*/;
assign _10539_ = D[15] ^ Q[37] /*28742*/;
assign _10536_ = _10024_ & _10539_ /*28738*/;
assign _10537_ = _10024_ ^ _10539_ /*28741*/;
assign _10538_ = _10530_ & _10537_ /*28739*/;
assign _10535_ = _10536_ | _10538_ /*28737*/;
assign _10410_ = _10530_ ^ _10537_ /*28740*/;
assign _10544_ = D[16] ^ Q[37] /*28736*/;
assign _10541_ = _10025_ & _10544_ /*28732*/;
assign _10542_ = _10025_ ^ _10544_ /*28735*/;
assign _10543_ = _10535_ & _10542_ /*28733*/;
assign _10540_ = _10541_ | _10543_ /*28731*/;
assign _10411_ = _10535_ ^ _10542_ /*28734*/;
assign _10549_ = D[17] ^ Q[37] /*28730*/;
assign _10546_ = _10026_ & _10549_ /*28726*/;
assign _10547_ = _10026_ ^ _10549_ /*28729*/;
assign _10548_ = _10540_ & _10547_ /*28727*/;
assign _10545_ = _10546_ | _10548_ /*28725*/;
assign _10412_ = _10540_ ^ _10547_ /*28728*/;
assign _10554_ = D[18] ^ Q[37] /*28724*/;
assign _10551_ = _10027_ & _10554_ /*28720*/;
assign _10552_ = _10027_ ^ _10554_ /*28723*/;
assign _10553_ = _10545_ & _10552_ /*28721*/;
assign _10550_ = _10551_ | _10553_ /*28719*/;
assign _10413_ = _10545_ ^ _10552_ /*28722*/;
assign _10559_ = D[19] ^ Q[37] /*28718*/;
assign _10556_ = _10028_ & _10559_ /*28714*/;
assign _10557_ = _10028_ ^ _10559_ /*28717*/;
assign _10558_ = _10550_ & _10557_ /*28715*/;
assign _10555_ = _10556_ | _10558_ /*28713*/;
assign _10414_ = _10550_ ^ _10557_ /*28716*/;
assign _10564_ = D[20] ^ Q[37] /*28712*/;
assign _10561_ = _10029_ & _10564_ /*28708*/;
assign _10562_ = _10029_ ^ _10564_ /*28711*/;
assign _10563_ = _10555_ & _10562_ /*28709*/;
assign _10560_ = _10561_ | _10563_ /*28707*/;
assign _10415_ = _10555_ ^ _10562_ /*28710*/;
assign _10569_ = D[21] ^ Q[37] /*28706*/;
assign _10566_ = _10030_ & _10569_ /*28702*/;
assign _10567_ = _10030_ ^ _10569_ /*28705*/;
assign _10568_ = _10560_ & _10567_ /*28703*/;
assign _10565_ = _10566_ | _10568_ /*28701*/;
assign _10416_ = _10560_ ^ _10567_ /*28704*/;
assign _10574_ = D[22] ^ Q[37] /*28700*/;
assign _10571_ = _10031_ & _10574_ /*28696*/;
assign _10572_ = _10031_ ^ _10574_ /*28699*/;
assign _10573_ = _10565_ & _10572_ /*28697*/;
assign _10570_ = _10571_ | _10573_ /*28695*/;
assign _10417_ = _10565_ ^ _10572_ /*28698*/;
assign _10579_ = D[23] ^ Q[37] /*28694*/;
assign _10576_ = _10032_ & _10579_ /*28690*/;
assign _10577_ = _10032_ ^ _10579_ /*28693*/;
assign _10578_ = _10570_ & _10577_ /*28691*/;
assign _10575_ = _10576_ | _10578_ /*28689*/;
assign _10418_ = _10570_ ^ _10577_ /*28692*/;
assign _10584_ = D[24] ^ Q[37] /*28688*/;
assign _10581_ = _10033_ & _10584_ /*28684*/;
assign _10582_ = _10033_ ^ _10584_ /*28687*/;
assign _10583_ = _10575_ & _10582_ /*28685*/;
assign _10580_ = _10581_ | _10583_ /*28683*/;
assign _10419_ = _10575_ ^ _10582_ /*28686*/;
assign _10589_ = D[25] ^ Q[37] /*28682*/;
assign _10586_ = _10034_ & _10589_ /*28678*/;
assign _10587_ = _10034_ ^ _10589_ /*28681*/;
assign _10588_ = _10580_ & _10587_ /*28679*/;
assign _10585_ = _10586_ | _10588_ /*28677*/;
assign _10420_ = _10580_ ^ _10587_ /*28680*/;
assign _10594_ = D[26] ^ Q[37] /*28676*/;
assign _10591_ = _10035_ & _10594_ /*28672*/;
assign _10592_ = _10035_ ^ _10594_ /*28675*/;
assign _10593_ = _10585_ & _10592_ /*28673*/;
assign _10590_ = _10591_ | _10593_ /*28671*/;
assign _10421_ = _10585_ ^ _10592_ /*28674*/;
assign _10599_ = D[27] ^ Q[37] /*28670*/;
assign _10596_ = _10036_ & _10599_ /*28666*/;
assign _10597_ = _10036_ ^ _10599_ /*28669*/;
assign _10598_ = _10590_ & _10597_ /*28667*/;
assign _10595_ = _10596_ | _10598_ /*28665*/;
assign _10422_ = _10590_ ^ _10597_ /*28668*/;
assign _10604_ = D[28] ^ Q[37] /*28664*/;
assign _10601_ = _10037_ & _10604_ /*28660*/;
assign _10602_ = _10037_ ^ _10604_ /*28663*/;
assign _10603_ = _10595_ & _10602_ /*28661*/;
assign _10600_ = _10601_ | _10603_ /*28659*/;
assign _10423_ = _10595_ ^ _10602_ /*28662*/;
assign _10609_ = D[29] ^ Q[37] /*28658*/;
assign _10606_ = _10038_ & _10609_ /*28654*/;
assign _10607_ = _10038_ ^ _10609_ /*28657*/;
assign _10608_ = _10600_ & _10607_ /*28655*/;
assign _10605_ = _10606_ | _10608_ /*28653*/;
assign _10424_ = _10600_ ^ _10607_ /*28656*/;
assign _10614_ = D[30] ^ Q[37] /*28652*/;
assign _10611_ = _10039_ & _10614_ /*28648*/;
assign _10612_ = _10039_ ^ _10614_ /*28651*/;
assign _10613_ = _10605_ & _10612_ /*28649*/;
assign _10610_ = _10611_ | _10613_ /*28647*/;
assign _10425_ = _10605_ ^ _10612_ /*28650*/;
assign _10619_ = D[31] ^ Q[37] /*28646*/;
assign _10616_ = _10040_ & _10619_ /*28642*/;
assign _10617_ = _10040_ ^ _10619_ /*28645*/;
assign _10618_ = _10610_ & _10617_ /*28643*/;
assign _10615_ = _10616_ | _10618_ /*28641*/;
assign _10426_ = _10610_ ^ _10617_ /*28644*/;
assign _10624_ = D[32] ^ Q[37] /*28640*/;
assign _10621_ = _10041_ & _10624_ /*28636*/;
assign _10622_ = _10041_ ^ _10624_ /*28639*/;
assign _10623_ = _10615_ & _10622_ /*28637*/;
assign _10620_ = _10621_ | _10623_ /*28635*/;
assign _10427_ = _10615_ ^ _10622_ /*28638*/;
assign _10629_ = D[33] ^ Q[37] /*28634*/;
assign _10626_ = _10042_ & _10629_ /*28630*/;
assign _10627_ = _10042_ ^ _10629_ /*28633*/;
assign _10628_ = _10620_ & _10627_ /*28631*/;
assign _10625_ = _10626_ | _10628_ /*28629*/;
assign _10428_ = _10620_ ^ _10627_ /*28632*/;
assign _10634_ = D[34] ^ Q[37] /*28628*/;
assign _10631_ = _10043_ & _10634_ /*28624*/;
assign _10632_ = _10043_ ^ _10634_ /*28627*/;
assign _10633_ = _10625_ & _10632_ /*28625*/;
assign _10630_ = _10631_ | _10633_ /*28623*/;
assign _10429_ = _10625_ ^ _10632_ /*28626*/;
assign _10639_ = D[35] ^ Q[37] /*28622*/;
assign _10636_ = _10044_ & _10639_ /*28618*/;
assign _10637_ = _10044_ ^ _10639_ /*28621*/;
assign _10638_ = _10630_ & _10637_ /*28619*/;
assign _10635_ = _10636_ | _10638_ /*28617*/;
assign _10430_ = _10630_ ^ _10637_ /*28620*/;
assign _10644_ = D[36] ^ Q[37] /*28616*/;
assign _10641_ = _10045_ & _10644_ /*28612*/;
assign _10642_ = _10045_ ^ _10644_ /*28615*/;
assign _10643_ = _10635_ & _10642_ /*28613*/;
assign _10640_ = _10641_ | _10643_ /*28611*/;
assign _10431_ = _10635_ ^ _10642_ /*28614*/;
assign _10649_ = D[37] ^ Q[37] /*28610*/;
assign _10646_ = _10046_ & _10649_ /*28606*/;
assign _10647_ = _10046_ ^ _10649_ /*28609*/;
assign _10648_ = _10640_ & _10647_ /*28607*/;
assign _10645_ = _10646_ | _10648_ /*28605*/;
assign _10432_ = _10640_ ^ _10647_ /*28608*/;
assign _10654_ = D[38] ^ Q[37] /*28604*/;
assign _10651_ = _10047_ & _10654_ /*28600*/;
assign _10652_ = _10047_ ^ _10654_ /*28603*/;
assign _10653_ = _10645_ & _10652_ /*28601*/;
assign _10650_ = _10651_ | _10653_ /*28599*/;
assign _10433_ = _10645_ ^ _10652_ /*28602*/;
assign _10659_ = D[39] ^ Q[37] /*28598*/;
assign _10656_ = _10048_ & _10659_ /*28594*/;
assign _10657_ = _10048_ ^ _10659_ /*28597*/;
assign _10658_ = _10650_ & _10657_ /*28595*/;
assign _10655_ = _10656_ | _10658_ /*28593*/;
assign _10434_ = _10650_ ^ _10657_ /*28596*/;
assign _10664_ = D[40] ^ Q[37] /*28592*/;
assign _10661_ = _10049_ & _10664_ /*28588*/;
assign _10662_ = _10049_ ^ _10664_ /*28591*/;
assign _10663_ = _10655_ & _10662_ /*28589*/;
assign _10660_ = _10661_ | _10663_ /*28587*/;
assign _10435_ = _10655_ ^ _10662_ /*28590*/;
assign _10669_ = D[41] ^ Q[37] /*28586*/;
assign _10666_ = _10050_ & _10669_ /*28582*/;
assign _10667_ = _10050_ ^ _10669_ /*28585*/;
assign _10668_ = _10660_ & _10667_ /*28583*/;
assign _10665_ = _10666_ | _10668_ /*28581*/;
assign _10436_ = _10660_ ^ _10667_ /*28584*/;
assign _10674_ = D[42] ^ Q[37] /*28580*/;
assign _10671_ = _10051_ & _10674_ /*28576*/;
assign _10672_ = _10051_ ^ _10674_ /*28579*/;
assign _10673_ = _10665_ & _10672_ /*28577*/;
assign _10670_ = _10671_ | _10673_ /*28575*/;
assign _10437_ = _10665_ ^ _10672_ /*28578*/;
assign _10679_ = D[43] ^ Q[37] /*28574*/;
assign _10676_ = _10052_ & _10679_ /*28570*/;
assign _10677_ = _10052_ ^ _10679_ /*28573*/;
assign _10678_ = _10670_ & _10677_ /*28571*/;
assign _10675_ = _10676_ | _10678_ /*28569*/;
assign _10438_ = _10670_ ^ _10677_ /*28572*/;
assign _10684_ = D[44] ^ Q[37] /*28568*/;
assign _10681_ = _10053_ & _10684_ /*28564*/;
assign _10682_ = _10053_ ^ _10684_ /*28567*/;
assign _10683_ = _10675_ & _10682_ /*28565*/;
assign _10680_ = _10681_ | _10683_ /*28563*/;
assign _10439_ = _10675_ ^ _10682_ /*28566*/;
assign _10689_ = D[45] ^ Q[37] /*28562*/;
assign _10686_ = _10054_ & _10689_ /*28558*/;
assign _10687_ = _10054_ ^ _10689_ /*28561*/;
assign _10688_ = _10680_ & _10687_ /*28559*/;
assign _10685_ = _10686_ | _10688_ /*28557*/;
assign _10440_ = _10680_ ^ _10687_ /*28560*/;
assign _10694_ = D[46] ^ Q[37] /*28556*/;
assign _10691_ = _10055_ & _10694_ /*28552*/;
assign _10692_ = _10055_ ^ _10694_ /*28555*/;
assign _10693_ = _10685_ & _10692_ /*28553*/;
assign _10690_ = _10691_ | _10693_ /*28551*/;
assign _10441_ = _10685_ ^ _10692_ /*28554*/;
assign _10699_ = D[47] ^ Q[37] /*28550*/;
assign _10696_ = _10056_ & _10699_ /*28546*/;
assign _10697_ = _10056_ ^ _10699_ /*28549*/;
assign _10698_ = _10690_ & _10697_ /*28547*/;
assign _10695_ = _10696_ | _10698_ /*28545*/;
assign _10442_ = _10690_ ^ _10697_ /*28548*/;
assign _10704_ = D[48] ^ Q[37] /*28544*/;
assign _10701_ = _10057_ & _10704_ /*28540*/;
assign _10702_ = _10057_ ^ _10704_ /*28543*/;
assign _10703_ = _10695_ & _10702_ /*28541*/;
assign _10700_ = _10701_ | _10703_ /*28539*/;
assign _10443_ = _10695_ ^ _10702_ /*28542*/;
assign _10709_ = D[49] ^ Q[37] /*28538*/;
assign _10706_ = _10058_ & _10709_ /*28534*/;
assign _10707_ = _10058_ ^ _10709_ /*28537*/;
assign _10708_ = _10700_ & _10707_ /*28535*/;
assign _10705_ = _10706_ | _10708_ /*28533*/;
assign _10444_ = _10700_ ^ _10707_ /*28536*/;
assign _10714_ = D[50] ^ Q[37] /*28532*/;
assign _10711_ = _10059_ & _10714_ /*28528*/;
assign _10712_ = _10059_ ^ _10714_ /*28531*/;
assign _10713_ = _10705_ & _10712_ /*28529*/;
assign _10710_ = _10711_ | _10713_ /*28527*/;
assign _10445_ = _10705_ ^ _10712_ /*28530*/;
assign _10719_ = D[51] ^ Q[37] /*28526*/;
assign _10716_ = _10060_ & _10719_ /*28522*/;
assign _10717_ = _10060_ ^ _10719_ /*28525*/;
assign _10718_ = _10710_ & _10717_ /*28523*/;
assign _10715_ = _10716_ | _10718_ /*28521*/;
assign _10446_ = _10710_ ^ _10717_ /*28524*/;
assign _10724_ = D[52] ^ Q[37] /*28520*/;
assign _10721_ = _10061_ & _10724_ /*28516*/;
assign _10722_ = _10061_ ^ _10724_ /*28519*/;
assign _10723_ = _10715_ & _10722_ /*28517*/;
assign _10720_ = _10721_ | _10723_ /*28515*/;
assign _10447_ = _10715_ ^ _10722_ /*28518*/;
assign _10729_ = D[53] ^ Q[37] /*28514*/;
assign _10726_ = _10062_ & _10729_ /*28510*/;
assign _10727_ = _10062_ ^ _10729_ /*28513*/;
assign _10728_ = _10720_ & _10727_ /*28511*/;
assign _10725_ = _10726_ | _10728_ /*28509*/;
assign _10448_ = _10720_ ^ _10727_ /*28512*/;
assign _10734_ = D[54] ^ Q[37] /*28508*/;
assign _10731_ = _10063_ & _10734_ /*28504*/;
assign _10732_ = _10063_ ^ _10734_ /*28507*/;
assign _10733_ = _10725_ & _10732_ /*28505*/;
assign _10730_ = _10731_ | _10733_ /*28503*/;
assign _10449_ = _10725_ ^ _10732_ /*28506*/;
assign _10739_ = D[55] ^ Q[37] /*28502*/;
assign _10736_ = _10064_ & _10739_ /*28498*/;
assign _10737_ = _10064_ ^ _10739_ /*28501*/;
assign _10738_ = _10730_ & _10737_ /*28499*/;
assign _10735_ = _10736_ | _10738_ /*28497*/;
assign _10450_ = _10730_ ^ _10737_ /*28500*/;
assign _10744_ = D[56] ^ Q[37] /*28496*/;
assign _10741_ = _10065_ & _10744_ /*28492*/;
assign _10742_ = _10065_ ^ _10744_ /*28495*/;
assign _10743_ = _10735_ & _10742_ /*28493*/;
assign _10740_ = _10741_ | _10743_ /*28491*/;
assign _10451_ = _10735_ ^ _10742_ /*28494*/;
assign _10749_ = D[57] ^ Q[37] /*28490*/;
assign _10746_ = _10066_ & _10749_ /*28486*/;
assign _10747_ = _10066_ ^ _10749_ /*28489*/;
assign _10748_ = _10740_ & _10747_ /*28487*/;
assign _10745_ = _10746_ | _10748_ /*28485*/;
assign _10452_ = _10740_ ^ _10747_ /*28488*/;
assign _10754_ = D[58] ^ Q[37] /*28484*/;
assign _10751_ = _10067_ & _10754_ /*28480*/;
assign _10752_ = _10067_ ^ _10754_ /*28483*/;
assign _10753_ = _10745_ & _10752_ /*28481*/;
assign _10750_ = _10751_ | _10753_ /*28479*/;
assign _10453_ = _10745_ ^ _10752_ /*28482*/;
assign _10759_ = D[59] ^ Q[37] /*28478*/;
assign _10756_ = _10068_ & _10759_ /*28474*/;
assign _10757_ = _10068_ ^ _10759_ /*28477*/;
assign _10758_ = _10750_ & _10757_ /*28475*/;
assign _10755_ = _10756_ | _10758_ /*28473*/;
assign _10454_ = _10750_ ^ _10757_ /*28476*/;
assign _10764_ = D[60] ^ Q[37] /*28472*/;
assign _10761_ = _10069_ & _10764_ /*28468*/;
assign _10762_ = _10069_ ^ _10764_ /*28471*/;
assign _10763_ = _10755_ & _10762_ /*28469*/;
assign _10760_ = _10761_ | _10763_ /*28467*/;
assign _10455_ = _10755_ ^ _10762_ /*28470*/;
assign _10769_ = D[61] ^ Q[37] /*28466*/;
assign _10766_ = _10070_ & _10769_ /*28462*/;
assign _10767_ = _10070_ ^ _10769_ /*28465*/;
assign _10768_ = _10760_ & _10767_ /*28463*/;
assign _10765_ = _10766_ | _10768_ /*28461*/;
assign _10456_ = _10760_ ^ _10767_ /*28464*/;
assign _10774_ = D[62] ^ Q[37] /*28460*/;
assign _10771_ = _10071_ & _10774_ /*28456*/;
assign _10772_ = _10071_ ^ _10774_ /*28459*/;
assign _10773_ = _10765_ & _10772_ /*28457*/;
assign _10770_ = _10771_ | _10773_ /*28455*/;
assign _10457_ = _10765_ ^ _10772_ /*28458*/;
assign _10778_ = zeroWire ^ Q[37] /*28454*/;
assign _10775_ = _10072_ & _10778_ /*28450*/;
assign _10776_ = _10072_ ^ _10778_ /*28453*/;
assign _10777_ = _10770_ & _10776_ /*28451*/;
assign Q[36] = _10775_ | _10777_ /*28449*/;
assign _10458_ = _10770_ ^ _10776_ /*28452*/;
assign _10849_ = D[0] ^ Q[36] /*28063*/;
assign _10846_ = R_0[35] & _10849_ /*28059*/;
assign _10847_ = R_0[35] ^ _10849_ /*28062*/;
assign _10848_ = Q[36] & _10847_ /*28060*/;
assign _10845_ = _10846_ | _10848_ /*28058*/;
assign _10780_ = Q[36] ^ _10847_ /*28061*/;
assign _10854_ = D[1] ^ Q[36] /*28057*/;
assign _10851_ = _10395_ & _10854_ /*28053*/;
assign _10852_ = _10395_ ^ _10854_ /*28056*/;
assign _10853_ = _10845_ & _10852_ /*28054*/;
assign _10850_ = _10851_ | _10853_ /*28052*/;
assign _10781_ = _10845_ ^ _10852_ /*28055*/;
assign _10859_ = D[2] ^ Q[36] /*28051*/;
assign _10856_ = _10396_ & _10859_ /*28047*/;
assign _10857_ = _10396_ ^ _10859_ /*28050*/;
assign _10858_ = _10850_ & _10857_ /*28048*/;
assign _10855_ = _10856_ | _10858_ /*28046*/;
assign _10782_ = _10850_ ^ _10857_ /*28049*/;
assign _10864_ = D[3] ^ Q[36] /*28045*/;
assign _10861_ = _10397_ & _10864_ /*28041*/;
assign _10862_ = _10397_ ^ _10864_ /*28044*/;
assign _10863_ = _10855_ & _10862_ /*28042*/;
assign _10860_ = _10861_ | _10863_ /*28040*/;
assign _10783_ = _10855_ ^ _10862_ /*28043*/;
assign _10869_ = D[4] ^ Q[36] /*28039*/;
assign _10866_ = _10398_ & _10869_ /*28035*/;
assign _10867_ = _10398_ ^ _10869_ /*28038*/;
assign _10868_ = _10860_ & _10867_ /*28036*/;
assign _10865_ = _10866_ | _10868_ /*28034*/;
assign _10784_ = _10860_ ^ _10867_ /*28037*/;
assign _10874_ = D[5] ^ Q[36] /*28033*/;
assign _10871_ = _10399_ & _10874_ /*28029*/;
assign _10872_ = _10399_ ^ _10874_ /*28032*/;
assign _10873_ = _10865_ & _10872_ /*28030*/;
assign _10870_ = _10871_ | _10873_ /*28028*/;
assign _10785_ = _10865_ ^ _10872_ /*28031*/;
assign _10879_ = D[6] ^ Q[36] /*28027*/;
assign _10876_ = _10400_ & _10879_ /*28023*/;
assign _10877_ = _10400_ ^ _10879_ /*28026*/;
assign _10878_ = _10870_ & _10877_ /*28024*/;
assign _10875_ = _10876_ | _10878_ /*28022*/;
assign _10786_ = _10870_ ^ _10877_ /*28025*/;
assign _10884_ = D[7] ^ Q[36] /*28021*/;
assign _10881_ = _10401_ & _10884_ /*28017*/;
assign _10882_ = _10401_ ^ _10884_ /*28020*/;
assign _10883_ = _10875_ & _10882_ /*28018*/;
assign _10880_ = _10881_ | _10883_ /*28016*/;
assign _10787_ = _10875_ ^ _10882_ /*28019*/;
assign _10889_ = D[8] ^ Q[36] /*28015*/;
assign _10886_ = _10402_ & _10889_ /*28011*/;
assign _10887_ = _10402_ ^ _10889_ /*28014*/;
assign _10888_ = _10880_ & _10887_ /*28012*/;
assign _10885_ = _10886_ | _10888_ /*28010*/;
assign _10788_ = _10880_ ^ _10887_ /*28013*/;
assign _10894_ = D[9] ^ Q[36] /*28009*/;
assign _10891_ = _10403_ & _10894_ /*28005*/;
assign _10892_ = _10403_ ^ _10894_ /*28008*/;
assign _10893_ = _10885_ & _10892_ /*28006*/;
assign _10890_ = _10891_ | _10893_ /*28004*/;
assign _10789_ = _10885_ ^ _10892_ /*28007*/;
assign _10899_ = D[10] ^ Q[36] /*28003*/;
assign _10896_ = _10404_ & _10899_ /*27999*/;
assign _10897_ = _10404_ ^ _10899_ /*28002*/;
assign _10898_ = _10890_ & _10897_ /*28000*/;
assign _10895_ = _10896_ | _10898_ /*27998*/;
assign _10790_ = _10890_ ^ _10897_ /*28001*/;
assign _10904_ = D[11] ^ Q[36] /*27997*/;
assign _10901_ = _10405_ & _10904_ /*27993*/;
assign _10902_ = _10405_ ^ _10904_ /*27996*/;
assign _10903_ = _10895_ & _10902_ /*27994*/;
assign _10900_ = _10901_ | _10903_ /*27992*/;
assign _10791_ = _10895_ ^ _10902_ /*27995*/;
assign _10909_ = D[12] ^ Q[36] /*27991*/;
assign _10906_ = _10406_ & _10909_ /*27987*/;
assign _10907_ = _10406_ ^ _10909_ /*27990*/;
assign _10908_ = _10900_ & _10907_ /*27988*/;
assign _10905_ = _10906_ | _10908_ /*27986*/;
assign _10792_ = _10900_ ^ _10907_ /*27989*/;
assign _10914_ = D[13] ^ Q[36] /*27985*/;
assign _10911_ = _10407_ & _10914_ /*27981*/;
assign _10912_ = _10407_ ^ _10914_ /*27984*/;
assign _10913_ = _10905_ & _10912_ /*27982*/;
assign _10910_ = _10911_ | _10913_ /*27980*/;
assign _10793_ = _10905_ ^ _10912_ /*27983*/;
assign _10919_ = D[14] ^ Q[36] /*27979*/;
assign _10916_ = _10408_ & _10919_ /*27975*/;
assign _10917_ = _10408_ ^ _10919_ /*27978*/;
assign _10918_ = _10910_ & _10917_ /*27976*/;
assign _10915_ = _10916_ | _10918_ /*27974*/;
assign _10794_ = _10910_ ^ _10917_ /*27977*/;
assign _10924_ = D[15] ^ Q[36] /*27973*/;
assign _10921_ = _10409_ & _10924_ /*27969*/;
assign _10922_ = _10409_ ^ _10924_ /*27972*/;
assign _10923_ = _10915_ & _10922_ /*27970*/;
assign _10920_ = _10921_ | _10923_ /*27968*/;
assign _10795_ = _10915_ ^ _10922_ /*27971*/;
assign _10929_ = D[16] ^ Q[36] /*27967*/;
assign _10926_ = _10410_ & _10929_ /*27963*/;
assign _10927_ = _10410_ ^ _10929_ /*27966*/;
assign _10928_ = _10920_ & _10927_ /*27964*/;
assign _10925_ = _10926_ | _10928_ /*27962*/;
assign _10796_ = _10920_ ^ _10927_ /*27965*/;
assign _10934_ = D[17] ^ Q[36] /*27961*/;
assign _10931_ = _10411_ & _10934_ /*27957*/;
assign _10932_ = _10411_ ^ _10934_ /*27960*/;
assign _10933_ = _10925_ & _10932_ /*27958*/;
assign _10930_ = _10931_ | _10933_ /*27956*/;
assign _10797_ = _10925_ ^ _10932_ /*27959*/;
assign _10939_ = D[18] ^ Q[36] /*27955*/;
assign _10936_ = _10412_ & _10939_ /*27951*/;
assign _10937_ = _10412_ ^ _10939_ /*27954*/;
assign _10938_ = _10930_ & _10937_ /*27952*/;
assign _10935_ = _10936_ | _10938_ /*27950*/;
assign _10798_ = _10930_ ^ _10937_ /*27953*/;
assign _10944_ = D[19] ^ Q[36] /*27949*/;
assign _10941_ = _10413_ & _10944_ /*27945*/;
assign _10942_ = _10413_ ^ _10944_ /*27948*/;
assign _10943_ = _10935_ & _10942_ /*27946*/;
assign _10940_ = _10941_ | _10943_ /*27944*/;
assign _10799_ = _10935_ ^ _10942_ /*27947*/;
assign _10949_ = D[20] ^ Q[36] /*27943*/;
assign _10946_ = _10414_ & _10949_ /*27939*/;
assign _10947_ = _10414_ ^ _10949_ /*27942*/;
assign _10948_ = _10940_ & _10947_ /*27940*/;
assign _10945_ = _10946_ | _10948_ /*27938*/;
assign _10800_ = _10940_ ^ _10947_ /*27941*/;
assign _10954_ = D[21] ^ Q[36] /*27937*/;
assign _10951_ = _10415_ & _10954_ /*27933*/;
assign _10952_ = _10415_ ^ _10954_ /*27936*/;
assign _10953_ = _10945_ & _10952_ /*27934*/;
assign _10950_ = _10951_ | _10953_ /*27932*/;
assign _10801_ = _10945_ ^ _10952_ /*27935*/;
assign _10959_ = D[22] ^ Q[36] /*27931*/;
assign _10956_ = _10416_ & _10959_ /*27927*/;
assign _10957_ = _10416_ ^ _10959_ /*27930*/;
assign _10958_ = _10950_ & _10957_ /*27928*/;
assign _10955_ = _10956_ | _10958_ /*27926*/;
assign _10802_ = _10950_ ^ _10957_ /*27929*/;
assign _10964_ = D[23] ^ Q[36] /*27925*/;
assign _10961_ = _10417_ & _10964_ /*27921*/;
assign _10962_ = _10417_ ^ _10964_ /*27924*/;
assign _10963_ = _10955_ & _10962_ /*27922*/;
assign _10960_ = _10961_ | _10963_ /*27920*/;
assign _10803_ = _10955_ ^ _10962_ /*27923*/;
assign _10969_ = D[24] ^ Q[36] /*27919*/;
assign _10966_ = _10418_ & _10969_ /*27915*/;
assign _10967_ = _10418_ ^ _10969_ /*27918*/;
assign _10968_ = _10960_ & _10967_ /*27916*/;
assign _10965_ = _10966_ | _10968_ /*27914*/;
assign _10804_ = _10960_ ^ _10967_ /*27917*/;
assign _10974_ = D[25] ^ Q[36] /*27913*/;
assign _10971_ = _10419_ & _10974_ /*27909*/;
assign _10972_ = _10419_ ^ _10974_ /*27912*/;
assign _10973_ = _10965_ & _10972_ /*27910*/;
assign _10970_ = _10971_ | _10973_ /*27908*/;
assign _10805_ = _10965_ ^ _10972_ /*27911*/;
assign _10979_ = D[26] ^ Q[36] /*27907*/;
assign _10976_ = _10420_ & _10979_ /*27903*/;
assign _10977_ = _10420_ ^ _10979_ /*27906*/;
assign _10978_ = _10970_ & _10977_ /*27904*/;
assign _10975_ = _10976_ | _10978_ /*27902*/;
assign _10806_ = _10970_ ^ _10977_ /*27905*/;
assign _10984_ = D[27] ^ Q[36] /*27901*/;
assign _10981_ = _10421_ & _10984_ /*27897*/;
assign _10982_ = _10421_ ^ _10984_ /*27900*/;
assign _10983_ = _10975_ & _10982_ /*27898*/;
assign _10980_ = _10981_ | _10983_ /*27896*/;
assign _10807_ = _10975_ ^ _10982_ /*27899*/;
assign _10989_ = D[28] ^ Q[36] /*27895*/;
assign _10986_ = _10422_ & _10989_ /*27891*/;
assign _10987_ = _10422_ ^ _10989_ /*27894*/;
assign _10988_ = _10980_ & _10987_ /*27892*/;
assign _10985_ = _10986_ | _10988_ /*27890*/;
assign _10808_ = _10980_ ^ _10987_ /*27893*/;
assign _10994_ = D[29] ^ Q[36] /*27889*/;
assign _10991_ = _10423_ & _10994_ /*27885*/;
assign _10992_ = _10423_ ^ _10994_ /*27888*/;
assign _10993_ = _10985_ & _10992_ /*27886*/;
assign _10990_ = _10991_ | _10993_ /*27884*/;
assign _10809_ = _10985_ ^ _10992_ /*27887*/;
assign _10999_ = D[30] ^ Q[36] /*27883*/;
assign _10996_ = _10424_ & _10999_ /*27879*/;
assign _10997_ = _10424_ ^ _10999_ /*27882*/;
assign _10998_ = _10990_ & _10997_ /*27880*/;
assign _10995_ = _10996_ | _10998_ /*27878*/;
assign _10810_ = _10990_ ^ _10997_ /*27881*/;
assign _11004_ = D[31] ^ Q[36] /*27877*/;
assign _11001_ = _10425_ & _11004_ /*27873*/;
assign _11002_ = _10425_ ^ _11004_ /*27876*/;
assign _11003_ = _10995_ & _11002_ /*27874*/;
assign _11000_ = _11001_ | _11003_ /*27872*/;
assign _10811_ = _10995_ ^ _11002_ /*27875*/;
assign _11009_ = D[32] ^ Q[36] /*27871*/;
assign _11006_ = _10426_ & _11009_ /*27867*/;
assign _11007_ = _10426_ ^ _11009_ /*27870*/;
assign _11008_ = _11000_ & _11007_ /*27868*/;
assign _11005_ = _11006_ | _11008_ /*27866*/;
assign _10812_ = _11000_ ^ _11007_ /*27869*/;
assign _11014_ = D[33] ^ Q[36] /*27865*/;
assign _11011_ = _10427_ & _11014_ /*27861*/;
assign _11012_ = _10427_ ^ _11014_ /*27864*/;
assign _11013_ = _11005_ & _11012_ /*27862*/;
assign _11010_ = _11011_ | _11013_ /*27860*/;
assign _10813_ = _11005_ ^ _11012_ /*27863*/;
assign _11019_ = D[34] ^ Q[36] /*27859*/;
assign _11016_ = _10428_ & _11019_ /*27855*/;
assign _11017_ = _10428_ ^ _11019_ /*27858*/;
assign _11018_ = _11010_ & _11017_ /*27856*/;
assign _11015_ = _11016_ | _11018_ /*27854*/;
assign _10814_ = _11010_ ^ _11017_ /*27857*/;
assign _11024_ = D[35] ^ Q[36] /*27853*/;
assign _11021_ = _10429_ & _11024_ /*27849*/;
assign _11022_ = _10429_ ^ _11024_ /*27852*/;
assign _11023_ = _11015_ & _11022_ /*27850*/;
assign _11020_ = _11021_ | _11023_ /*27848*/;
assign _10815_ = _11015_ ^ _11022_ /*27851*/;
assign _11029_ = D[36] ^ Q[36] /*27847*/;
assign _11026_ = _10430_ & _11029_ /*27843*/;
assign _11027_ = _10430_ ^ _11029_ /*27846*/;
assign _11028_ = _11020_ & _11027_ /*27844*/;
assign _11025_ = _11026_ | _11028_ /*27842*/;
assign _10816_ = _11020_ ^ _11027_ /*27845*/;
assign _11034_ = D[37] ^ Q[36] /*27841*/;
assign _11031_ = _10431_ & _11034_ /*27837*/;
assign _11032_ = _10431_ ^ _11034_ /*27840*/;
assign _11033_ = _11025_ & _11032_ /*27838*/;
assign _11030_ = _11031_ | _11033_ /*27836*/;
assign _10817_ = _11025_ ^ _11032_ /*27839*/;
assign _11039_ = D[38] ^ Q[36] /*27835*/;
assign _11036_ = _10432_ & _11039_ /*27831*/;
assign _11037_ = _10432_ ^ _11039_ /*27834*/;
assign _11038_ = _11030_ & _11037_ /*27832*/;
assign _11035_ = _11036_ | _11038_ /*27830*/;
assign _10818_ = _11030_ ^ _11037_ /*27833*/;
assign _11044_ = D[39] ^ Q[36] /*27829*/;
assign _11041_ = _10433_ & _11044_ /*27825*/;
assign _11042_ = _10433_ ^ _11044_ /*27828*/;
assign _11043_ = _11035_ & _11042_ /*27826*/;
assign _11040_ = _11041_ | _11043_ /*27824*/;
assign _10819_ = _11035_ ^ _11042_ /*27827*/;
assign _11049_ = D[40] ^ Q[36] /*27823*/;
assign _11046_ = _10434_ & _11049_ /*27819*/;
assign _11047_ = _10434_ ^ _11049_ /*27822*/;
assign _11048_ = _11040_ & _11047_ /*27820*/;
assign _11045_ = _11046_ | _11048_ /*27818*/;
assign _10820_ = _11040_ ^ _11047_ /*27821*/;
assign _11054_ = D[41] ^ Q[36] /*27817*/;
assign _11051_ = _10435_ & _11054_ /*27813*/;
assign _11052_ = _10435_ ^ _11054_ /*27816*/;
assign _11053_ = _11045_ & _11052_ /*27814*/;
assign _11050_ = _11051_ | _11053_ /*27812*/;
assign _10821_ = _11045_ ^ _11052_ /*27815*/;
assign _11059_ = D[42] ^ Q[36] /*27811*/;
assign _11056_ = _10436_ & _11059_ /*27807*/;
assign _11057_ = _10436_ ^ _11059_ /*27810*/;
assign _11058_ = _11050_ & _11057_ /*27808*/;
assign _11055_ = _11056_ | _11058_ /*27806*/;
assign _10822_ = _11050_ ^ _11057_ /*27809*/;
assign _11064_ = D[43] ^ Q[36] /*27805*/;
assign _11061_ = _10437_ & _11064_ /*27801*/;
assign _11062_ = _10437_ ^ _11064_ /*27804*/;
assign _11063_ = _11055_ & _11062_ /*27802*/;
assign _11060_ = _11061_ | _11063_ /*27800*/;
assign _10823_ = _11055_ ^ _11062_ /*27803*/;
assign _11069_ = D[44] ^ Q[36] /*27799*/;
assign _11066_ = _10438_ & _11069_ /*27795*/;
assign _11067_ = _10438_ ^ _11069_ /*27798*/;
assign _11068_ = _11060_ & _11067_ /*27796*/;
assign _11065_ = _11066_ | _11068_ /*27794*/;
assign _10824_ = _11060_ ^ _11067_ /*27797*/;
assign _11074_ = D[45] ^ Q[36] /*27793*/;
assign _11071_ = _10439_ & _11074_ /*27789*/;
assign _11072_ = _10439_ ^ _11074_ /*27792*/;
assign _11073_ = _11065_ & _11072_ /*27790*/;
assign _11070_ = _11071_ | _11073_ /*27788*/;
assign _10825_ = _11065_ ^ _11072_ /*27791*/;
assign _11079_ = D[46] ^ Q[36] /*27787*/;
assign _11076_ = _10440_ & _11079_ /*27783*/;
assign _11077_ = _10440_ ^ _11079_ /*27786*/;
assign _11078_ = _11070_ & _11077_ /*27784*/;
assign _11075_ = _11076_ | _11078_ /*27782*/;
assign _10826_ = _11070_ ^ _11077_ /*27785*/;
assign _11084_ = D[47] ^ Q[36] /*27781*/;
assign _11081_ = _10441_ & _11084_ /*27777*/;
assign _11082_ = _10441_ ^ _11084_ /*27780*/;
assign _11083_ = _11075_ & _11082_ /*27778*/;
assign _11080_ = _11081_ | _11083_ /*27776*/;
assign _10827_ = _11075_ ^ _11082_ /*27779*/;
assign _11089_ = D[48] ^ Q[36] /*27775*/;
assign _11086_ = _10442_ & _11089_ /*27771*/;
assign _11087_ = _10442_ ^ _11089_ /*27774*/;
assign _11088_ = _11080_ & _11087_ /*27772*/;
assign _11085_ = _11086_ | _11088_ /*27770*/;
assign _10828_ = _11080_ ^ _11087_ /*27773*/;
assign _11094_ = D[49] ^ Q[36] /*27769*/;
assign _11091_ = _10443_ & _11094_ /*27765*/;
assign _11092_ = _10443_ ^ _11094_ /*27768*/;
assign _11093_ = _11085_ & _11092_ /*27766*/;
assign _11090_ = _11091_ | _11093_ /*27764*/;
assign _10829_ = _11085_ ^ _11092_ /*27767*/;
assign _11099_ = D[50] ^ Q[36] /*27763*/;
assign _11096_ = _10444_ & _11099_ /*27759*/;
assign _11097_ = _10444_ ^ _11099_ /*27762*/;
assign _11098_ = _11090_ & _11097_ /*27760*/;
assign _11095_ = _11096_ | _11098_ /*27758*/;
assign _10830_ = _11090_ ^ _11097_ /*27761*/;
assign _11104_ = D[51] ^ Q[36] /*27757*/;
assign _11101_ = _10445_ & _11104_ /*27753*/;
assign _11102_ = _10445_ ^ _11104_ /*27756*/;
assign _11103_ = _11095_ & _11102_ /*27754*/;
assign _11100_ = _11101_ | _11103_ /*27752*/;
assign _10831_ = _11095_ ^ _11102_ /*27755*/;
assign _11109_ = D[52] ^ Q[36] /*27751*/;
assign _11106_ = _10446_ & _11109_ /*27747*/;
assign _11107_ = _10446_ ^ _11109_ /*27750*/;
assign _11108_ = _11100_ & _11107_ /*27748*/;
assign _11105_ = _11106_ | _11108_ /*27746*/;
assign _10832_ = _11100_ ^ _11107_ /*27749*/;
assign _11114_ = D[53] ^ Q[36] /*27745*/;
assign _11111_ = _10447_ & _11114_ /*27741*/;
assign _11112_ = _10447_ ^ _11114_ /*27744*/;
assign _11113_ = _11105_ & _11112_ /*27742*/;
assign _11110_ = _11111_ | _11113_ /*27740*/;
assign _10833_ = _11105_ ^ _11112_ /*27743*/;
assign _11119_ = D[54] ^ Q[36] /*27739*/;
assign _11116_ = _10448_ & _11119_ /*27735*/;
assign _11117_ = _10448_ ^ _11119_ /*27738*/;
assign _11118_ = _11110_ & _11117_ /*27736*/;
assign _11115_ = _11116_ | _11118_ /*27734*/;
assign _10834_ = _11110_ ^ _11117_ /*27737*/;
assign _11124_ = D[55] ^ Q[36] /*27733*/;
assign _11121_ = _10449_ & _11124_ /*27729*/;
assign _11122_ = _10449_ ^ _11124_ /*27732*/;
assign _11123_ = _11115_ & _11122_ /*27730*/;
assign _11120_ = _11121_ | _11123_ /*27728*/;
assign _10835_ = _11115_ ^ _11122_ /*27731*/;
assign _11129_ = D[56] ^ Q[36] /*27727*/;
assign _11126_ = _10450_ & _11129_ /*27723*/;
assign _11127_ = _10450_ ^ _11129_ /*27726*/;
assign _11128_ = _11120_ & _11127_ /*27724*/;
assign _11125_ = _11126_ | _11128_ /*27722*/;
assign _10836_ = _11120_ ^ _11127_ /*27725*/;
assign _11134_ = D[57] ^ Q[36] /*27721*/;
assign _11131_ = _10451_ & _11134_ /*27717*/;
assign _11132_ = _10451_ ^ _11134_ /*27720*/;
assign _11133_ = _11125_ & _11132_ /*27718*/;
assign _11130_ = _11131_ | _11133_ /*27716*/;
assign _10837_ = _11125_ ^ _11132_ /*27719*/;
assign _11139_ = D[58] ^ Q[36] /*27715*/;
assign _11136_ = _10452_ & _11139_ /*27711*/;
assign _11137_ = _10452_ ^ _11139_ /*27714*/;
assign _11138_ = _11130_ & _11137_ /*27712*/;
assign _11135_ = _11136_ | _11138_ /*27710*/;
assign _10838_ = _11130_ ^ _11137_ /*27713*/;
assign _11144_ = D[59] ^ Q[36] /*27709*/;
assign _11141_ = _10453_ & _11144_ /*27705*/;
assign _11142_ = _10453_ ^ _11144_ /*27708*/;
assign _11143_ = _11135_ & _11142_ /*27706*/;
assign _11140_ = _11141_ | _11143_ /*27704*/;
assign _10839_ = _11135_ ^ _11142_ /*27707*/;
assign _11149_ = D[60] ^ Q[36] /*27703*/;
assign _11146_ = _10454_ & _11149_ /*27699*/;
assign _11147_ = _10454_ ^ _11149_ /*27702*/;
assign _11148_ = _11140_ & _11147_ /*27700*/;
assign _11145_ = _11146_ | _11148_ /*27698*/;
assign _10840_ = _11140_ ^ _11147_ /*27701*/;
assign _11154_ = D[61] ^ Q[36] /*27697*/;
assign _11151_ = _10455_ & _11154_ /*27693*/;
assign _11152_ = _10455_ ^ _11154_ /*27696*/;
assign _11153_ = _11145_ & _11152_ /*27694*/;
assign _11150_ = _11151_ | _11153_ /*27692*/;
assign _10841_ = _11145_ ^ _11152_ /*27695*/;
assign _11159_ = D[62] ^ Q[36] /*27691*/;
assign _11156_ = _10456_ & _11159_ /*27687*/;
assign _11157_ = _10456_ ^ _11159_ /*27690*/;
assign _11158_ = _11150_ & _11157_ /*27688*/;
assign _11155_ = _11156_ | _11158_ /*27686*/;
assign _10842_ = _11150_ ^ _11157_ /*27689*/;
assign _11163_ = zeroWire ^ Q[36] /*27685*/;
assign _11160_ = _10457_ & _11163_ /*27681*/;
assign _11161_ = _10457_ ^ _11163_ /*27684*/;
assign _11162_ = _11155_ & _11161_ /*27682*/;
assign Q[35] = _11160_ | _11162_ /*27680*/;
assign _10843_ = _11155_ ^ _11161_ /*27683*/;
assign _11234_ = D[0] ^ Q[35] /*27294*/;
assign _11231_ = R_0[34] & _11234_ /*27290*/;
assign _11232_ = R_0[34] ^ _11234_ /*27293*/;
assign _11233_ = Q[35] & _11232_ /*27291*/;
assign _11230_ = _11231_ | _11233_ /*27289*/;
assign _11165_ = Q[35] ^ _11232_ /*27292*/;
assign _11239_ = D[1] ^ Q[35] /*27288*/;
assign _11236_ = _10780_ & _11239_ /*27284*/;
assign _11237_ = _10780_ ^ _11239_ /*27287*/;
assign _11238_ = _11230_ & _11237_ /*27285*/;
assign _11235_ = _11236_ | _11238_ /*27283*/;
assign _11166_ = _11230_ ^ _11237_ /*27286*/;
assign _11244_ = D[2] ^ Q[35] /*27282*/;
assign _11241_ = _10781_ & _11244_ /*27278*/;
assign _11242_ = _10781_ ^ _11244_ /*27281*/;
assign _11243_ = _11235_ & _11242_ /*27279*/;
assign _11240_ = _11241_ | _11243_ /*27277*/;
assign _11167_ = _11235_ ^ _11242_ /*27280*/;
assign _11249_ = D[3] ^ Q[35] /*27276*/;
assign _11246_ = _10782_ & _11249_ /*27272*/;
assign _11247_ = _10782_ ^ _11249_ /*27275*/;
assign _11248_ = _11240_ & _11247_ /*27273*/;
assign _11245_ = _11246_ | _11248_ /*27271*/;
assign _11168_ = _11240_ ^ _11247_ /*27274*/;
assign _11254_ = D[4] ^ Q[35] /*27270*/;
assign _11251_ = _10783_ & _11254_ /*27266*/;
assign _11252_ = _10783_ ^ _11254_ /*27269*/;
assign _11253_ = _11245_ & _11252_ /*27267*/;
assign _11250_ = _11251_ | _11253_ /*27265*/;
assign _11169_ = _11245_ ^ _11252_ /*27268*/;
assign _11259_ = D[5] ^ Q[35] /*27264*/;
assign _11256_ = _10784_ & _11259_ /*27260*/;
assign _11257_ = _10784_ ^ _11259_ /*27263*/;
assign _11258_ = _11250_ & _11257_ /*27261*/;
assign _11255_ = _11256_ | _11258_ /*27259*/;
assign _11170_ = _11250_ ^ _11257_ /*27262*/;
assign _11264_ = D[6] ^ Q[35] /*27258*/;
assign _11261_ = _10785_ & _11264_ /*27254*/;
assign _11262_ = _10785_ ^ _11264_ /*27257*/;
assign _11263_ = _11255_ & _11262_ /*27255*/;
assign _11260_ = _11261_ | _11263_ /*27253*/;
assign _11171_ = _11255_ ^ _11262_ /*27256*/;
assign _11269_ = D[7] ^ Q[35] /*27252*/;
assign _11266_ = _10786_ & _11269_ /*27248*/;
assign _11267_ = _10786_ ^ _11269_ /*27251*/;
assign _11268_ = _11260_ & _11267_ /*27249*/;
assign _11265_ = _11266_ | _11268_ /*27247*/;
assign _11172_ = _11260_ ^ _11267_ /*27250*/;
assign _11274_ = D[8] ^ Q[35] /*27246*/;
assign _11271_ = _10787_ & _11274_ /*27242*/;
assign _11272_ = _10787_ ^ _11274_ /*27245*/;
assign _11273_ = _11265_ & _11272_ /*27243*/;
assign _11270_ = _11271_ | _11273_ /*27241*/;
assign _11173_ = _11265_ ^ _11272_ /*27244*/;
assign _11279_ = D[9] ^ Q[35] /*27240*/;
assign _11276_ = _10788_ & _11279_ /*27236*/;
assign _11277_ = _10788_ ^ _11279_ /*27239*/;
assign _11278_ = _11270_ & _11277_ /*27237*/;
assign _11275_ = _11276_ | _11278_ /*27235*/;
assign _11174_ = _11270_ ^ _11277_ /*27238*/;
assign _11284_ = D[10] ^ Q[35] /*27234*/;
assign _11281_ = _10789_ & _11284_ /*27230*/;
assign _11282_ = _10789_ ^ _11284_ /*27233*/;
assign _11283_ = _11275_ & _11282_ /*27231*/;
assign _11280_ = _11281_ | _11283_ /*27229*/;
assign _11175_ = _11275_ ^ _11282_ /*27232*/;
assign _11289_ = D[11] ^ Q[35] /*27228*/;
assign _11286_ = _10790_ & _11289_ /*27224*/;
assign _11287_ = _10790_ ^ _11289_ /*27227*/;
assign _11288_ = _11280_ & _11287_ /*27225*/;
assign _11285_ = _11286_ | _11288_ /*27223*/;
assign _11176_ = _11280_ ^ _11287_ /*27226*/;
assign _11294_ = D[12] ^ Q[35] /*27222*/;
assign _11291_ = _10791_ & _11294_ /*27218*/;
assign _11292_ = _10791_ ^ _11294_ /*27221*/;
assign _11293_ = _11285_ & _11292_ /*27219*/;
assign _11290_ = _11291_ | _11293_ /*27217*/;
assign _11177_ = _11285_ ^ _11292_ /*27220*/;
assign _11299_ = D[13] ^ Q[35] /*27216*/;
assign _11296_ = _10792_ & _11299_ /*27212*/;
assign _11297_ = _10792_ ^ _11299_ /*27215*/;
assign _11298_ = _11290_ & _11297_ /*27213*/;
assign _11295_ = _11296_ | _11298_ /*27211*/;
assign _11178_ = _11290_ ^ _11297_ /*27214*/;
assign _11304_ = D[14] ^ Q[35] /*27210*/;
assign _11301_ = _10793_ & _11304_ /*27206*/;
assign _11302_ = _10793_ ^ _11304_ /*27209*/;
assign _11303_ = _11295_ & _11302_ /*27207*/;
assign _11300_ = _11301_ | _11303_ /*27205*/;
assign _11179_ = _11295_ ^ _11302_ /*27208*/;
assign _11309_ = D[15] ^ Q[35] /*27204*/;
assign _11306_ = _10794_ & _11309_ /*27200*/;
assign _11307_ = _10794_ ^ _11309_ /*27203*/;
assign _11308_ = _11300_ & _11307_ /*27201*/;
assign _11305_ = _11306_ | _11308_ /*27199*/;
assign _11180_ = _11300_ ^ _11307_ /*27202*/;
assign _11314_ = D[16] ^ Q[35] /*27198*/;
assign _11311_ = _10795_ & _11314_ /*27194*/;
assign _11312_ = _10795_ ^ _11314_ /*27197*/;
assign _11313_ = _11305_ & _11312_ /*27195*/;
assign _11310_ = _11311_ | _11313_ /*27193*/;
assign _11181_ = _11305_ ^ _11312_ /*27196*/;
assign _11319_ = D[17] ^ Q[35] /*27192*/;
assign _11316_ = _10796_ & _11319_ /*27188*/;
assign _11317_ = _10796_ ^ _11319_ /*27191*/;
assign _11318_ = _11310_ & _11317_ /*27189*/;
assign _11315_ = _11316_ | _11318_ /*27187*/;
assign _11182_ = _11310_ ^ _11317_ /*27190*/;
assign _11324_ = D[18] ^ Q[35] /*27186*/;
assign _11321_ = _10797_ & _11324_ /*27182*/;
assign _11322_ = _10797_ ^ _11324_ /*27185*/;
assign _11323_ = _11315_ & _11322_ /*27183*/;
assign _11320_ = _11321_ | _11323_ /*27181*/;
assign _11183_ = _11315_ ^ _11322_ /*27184*/;
assign _11329_ = D[19] ^ Q[35] /*27180*/;
assign _11326_ = _10798_ & _11329_ /*27176*/;
assign _11327_ = _10798_ ^ _11329_ /*27179*/;
assign _11328_ = _11320_ & _11327_ /*27177*/;
assign _11325_ = _11326_ | _11328_ /*27175*/;
assign _11184_ = _11320_ ^ _11327_ /*27178*/;
assign _11334_ = D[20] ^ Q[35] /*27174*/;
assign _11331_ = _10799_ & _11334_ /*27170*/;
assign _11332_ = _10799_ ^ _11334_ /*27173*/;
assign _11333_ = _11325_ & _11332_ /*27171*/;
assign _11330_ = _11331_ | _11333_ /*27169*/;
assign _11185_ = _11325_ ^ _11332_ /*27172*/;
assign _11339_ = D[21] ^ Q[35] /*27168*/;
assign _11336_ = _10800_ & _11339_ /*27164*/;
assign _11337_ = _10800_ ^ _11339_ /*27167*/;
assign _11338_ = _11330_ & _11337_ /*27165*/;
assign _11335_ = _11336_ | _11338_ /*27163*/;
assign _11186_ = _11330_ ^ _11337_ /*27166*/;
assign _11344_ = D[22] ^ Q[35] /*27162*/;
assign _11341_ = _10801_ & _11344_ /*27158*/;
assign _11342_ = _10801_ ^ _11344_ /*27161*/;
assign _11343_ = _11335_ & _11342_ /*27159*/;
assign _11340_ = _11341_ | _11343_ /*27157*/;
assign _11187_ = _11335_ ^ _11342_ /*27160*/;
assign _11349_ = D[23] ^ Q[35] /*27156*/;
assign _11346_ = _10802_ & _11349_ /*27152*/;
assign _11347_ = _10802_ ^ _11349_ /*27155*/;
assign _11348_ = _11340_ & _11347_ /*27153*/;
assign _11345_ = _11346_ | _11348_ /*27151*/;
assign _11188_ = _11340_ ^ _11347_ /*27154*/;
assign _11354_ = D[24] ^ Q[35] /*27150*/;
assign _11351_ = _10803_ & _11354_ /*27146*/;
assign _11352_ = _10803_ ^ _11354_ /*27149*/;
assign _11353_ = _11345_ & _11352_ /*27147*/;
assign _11350_ = _11351_ | _11353_ /*27145*/;
assign _11189_ = _11345_ ^ _11352_ /*27148*/;
assign _11359_ = D[25] ^ Q[35] /*27144*/;
assign _11356_ = _10804_ & _11359_ /*27140*/;
assign _11357_ = _10804_ ^ _11359_ /*27143*/;
assign _11358_ = _11350_ & _11357_ /*27141*/;
assign _11355_ = _11356_ | _11358_ /*27139*/;
assign _11190_ = _11350_ ^ _11357_ /*27142*/;
assign _11364_ = D[26] ^ Q[35] /*27138*/;
assign _11361_ = _10805_ & _11364_ /*27134*/;
assign _11362_ = _10805_ ^ _11364_ /*27137*/;
assign _11363_ = _11355_ & _11362_ /*27135*/;
assign _11360_ = _11361_ | _11363_ /*27133*/;
assign _11191_ = _11355_ ^ _11362_ /*27136*/;
assign _11369_ = D[27] ^ Q[35] /*27132*/;
assign _11366_ = _10806_ & _11369_ /*27128*/;
assign _11367_ = _10806_ ^ _11369_ /*27131*/;
assign _11368_ = _11360_ & _11367_ /*27129*/;
assign _11365_ = _11366_ | _11368_ /*27127*/;
assign _11192_ = _11360_ ^ _11367_ /*27130*/;
assign _11374_ = D[28] ^ Q[35] /*27126*/;
assign _11371_ = _10807_ & _11374_ /*27122*/;
assign _11372_ = _10807_ ^ _11374_ /*27125*/;
assign _11373_ = _11365_ & _11372_ /*27123*/;
assign _11370_ = _11371_ | _11373_ /*27121*/;
assign _11193_ = _11365_ ^ _11372_ /*27124*/;
assign _11379_ = D[29] ^ Q[35] /*27120*/;
assign _11376_ = _10808_ & _11379_ /*27116*/;
assign _11377_ = _10808_ ^ _11379_ /*27119*/;
assign _11378_ = _11370_ & _11377_ /*27117*/;
assign _11375_ = _11376_ | _11378_ /*27115*/;
assign _11194_ = _11370_ ^ _11377_ /*27118*/;
assign _11384_ = D[30] ^ Q[35] /*27114*/;
assign _11381_ = _10809_ & _11384_ /*27110*/;
assign _11382_ = _10809_ ^ _11384_ /*27113*/;
assign _11383_ = _11375_ & _11382_ /*27111*/;
assign _11380_ = _11381_ | _11383_ /*27109*/;
assign _11195_ = _11375_ ^ _11382_ /*27112*/;
assign _11389_ = D[31] ^ Q[35] /*27108*/;
assign _11386_ = _10810_ & _11389_ /*27104*/;
assign _11387_ = _10810_ ^ _11389_ /*27107*/;
assign _11388_ = _11380_ & _11387_ /*27105*/;
assign _11385_ = _11386_ | _11388_ /*27103*/;
assign _11196_ = _11380_ ^ _11387_ /*27106*/;
assign _11394_ = D[32] ^ Q[35] /*27102*/;
assign _11391_ = _10811_ & _11394_ /*27098*/;
assign _11392_ = _10811_ ^ _11394_ /*27101*/;
assign _11393_ = _11385_ & _11392_ /*27099*/;
assign _11390_ = _11391_ | _11393_ /*27097*/;
assign _11197_ = _11385_ ^ _11392_ /*27100*/;
assign _11399_ = D[33] ^ Q[35] /*27096*/;
assign _11396_ = _10812_ & _11399_ /*27092*/;
assign _11397_ = _10812_ ^ _11399_ /*27095*/;
assign _11398_ = _11390_ & _11397_ /*27093*/;
assign _11395_ = _11396_ | _11398_ /*27091*/;
assign _11198_ = _11390_ ^ _11397_ /*27094*/;
assign _11404_ = D[34] ^ Q[35] /*27090*/;
assign _11401_ = _10813_ & _11404_ /*27086*/;
assign _11402_ = _10813_ ^ _11404_ /*27089*/;
assign _11403_ = _11395_ & _11402_ /*27087*/;
assign _11400_ = _11401_ | _11403_ /*27085*/;
assign _11199_ = _11395_ ^ _11402_ /*27088*/;
assign _11409_ = D[35] ^ Q[35] /*27084*/;
assign _11406_ = _10814_ & _11409_ /*27080*/;
assign _11407_ = _10814_ ^ _11409_ /*27083*/;
assign _11408_ = _11400_ & _11407_ /*27081*/;
assign _11405_ = _11406_ | _11408_ /*27079*/;
assign _11200_ = _11400_ ^ _11407_ /*27082*/;
assign _11414_ = D[36] ^ Q[35] /*27078*/;
assign _11411_ = _10815_ & _11414_ /*27074*/;
assign _11412_ = _10815_ ^ _11414_ /*27077*/;
assign _11413_ = _11405_ & _11412_ /*27075*/;
assign _11410_ = _11411_ | _11413_ /*27073*/;
assign _11201_ = _11405_ ^ _11412_ /*27076*/;
assign _11419_ = D[37] ^ Q[35] /*27072*/;
assign _11416_ = _10816_ & _11419_ /*27068*/;
assign _11417_ = _10816_ ^ _11419_ /*27071*/;
assign _11418_ = _11410_ & _11417_ /*27069*/;
assign _11415_ = _11416_ | _11418_ /*27067*/;
assign _11202_ = _11410_ ^ _11417_ /*27070*/;
assign _11424_ = D[38] ^ Q[35] /*27066*/;
assign _11421_ = _10817_ & _11424_ /*27062*/;
assign _11422_ = _10817_ ^ _11424_ /*27065*/;
assign _11423_ = _11415_ & _11422_ /*27063*/;
assign _11420_ = _11421_ | _11423_ /*27061*/;
assign _11203_ = _11415_ ^ _11422_ /*27064*/;
assign _11429_ = D[39] ^ Q[35] /*27060*/;
assign _11426_ = _10818_ & _11429_ /*27056*/;
assign _11427_ = _10818_ ^ _11429_ /*27059*/;
assign _11428_ = _11420_ & _11427_ /*27057*/;
assign _11425_ = _11426_ | _11428_ /*27055*/;
assign _11204_ = _11420_ ^ _11427_ /*27058*/;
assign _11434_ = D[40] ^ Q[35] /*27054*/;
assign _11431_ = _10819_ & _11434_ /*27050*/;
assign _11432_ = _10819_ ^ _11434_ /*27053*/;
assign _11433_ = _11425_ & _11432_ /*27051*/;
assign _11430_ = _11431_ | _11433_ /*27049*/;
assign _11205_ = _11425_ ^ _11432_ /*27052*/;
assign _11439_ = D[41] ^ Q[35] /*27048*/;
assign _11436_ = _10820_ & _11439_ /*27044*/;
assign _11437_ = _10820_ ^ _11439_ /*27047*/;
assign _11438_ = _11430_ & _11437_ /*27045*/;
assign _11435_ = _11436_ | _11438_ /*27043*/;
assign _11206_ = _11430_ ^ _11437_ /*27046*/;
assign _11444_ = D[42] ^ Q[35] /*27042*/;
assign _11441_ = _10821_ & _11444_ /*27038*/;
assign _11442_ = _10821_ ^ _11444_ /*27041*/;
assign _11443_ = _11435_ & _11442_ /*27039*/;
assign _11440_ = _11441_ | _11443_ /*27037*/;
assign _11207_ = _11435_ ^ _11442_ /*27040*/;
assign _11449_ = D[43] ^ Q[35] /*27036*/;
assign _11446_ = _10822_ & _11449_ /*27032*/;
assign _11447_ = _10822_ ^ _11449_ /*27035*/;
assign _11448_ = _11440_ & _11447_ /*27033*/;
assign _11445_ = _11446_ | _11448_ /*27031*/;
assign _11208_ = _11440_ ^ _11447_ /*27034*/;
assign _11454_ = D[44] ^ Q[35] /*27030*/;
assign _11451_ = _10823_ & _11454_ /*27026*/;
assign _11452_ = _10823_ ^ _11454_ /*27029*/;
assign _11453_ = _11445_ & _11452_ /*27027*/;
assign _11450_ = _11451_ | _11453_ /*27025*/;
assign _11209_ = _11445_ ^ _11452_ /*27028*/;
assign _11459_ = D[45] ^ Q[35] /*27024*/;
assign _11456_ = _10824_ & _11459_ /*27020*/;
assign _11457_ = _10824_ ^ _11459_ /*27023*/;
assign _11458_ = _11450_ & _11457_ /*27021*/;
assign _11455_ = _11456_ | _11458_ /*27019*/;
assign _11210_ = _11450_ ^ _11457_ /*27022*/;
assign _11464_ = D[46] ^ Q[35] /*27018*/;
assign _11461_ = _10825_ & _11464_ /*27014*/;
assign _11462_ = _10825_ ^ _11464_ /*27017*/;
assign _11463_ = _11455_ & _11462_ /*27015*/;
assign _11460_ = _11461_ | _11463_ /*27013*/;
assign _11211_ = _11455_ ^ _11462_ /*27016*/;
assign _11469_ = D[47] ^ Q[35] /*27012*/;
assign _11466_ = _10826_ & _11469_ /*27008*/;
assign _11467_ = _10826_ ^ _11469_ /*27011*/;
assign _11468_ = _11460_ & _11467_ /*27009*/;
assign _11465_ = _11466_ | _11468_ /*27007*/;
assign _11212_ = _11460_ ^ _11467_ /*27010*/;
assign _11474_ = D[48] ^ Q[35] /*27006*/;
assign _11471_ = _10827_ & _11474_ /*27002*/;
assign _11472_ = _10827_ ^ _11474_ /*27005*/;
assign _11473_ = _11465_ & _11472_ /*27003*/;
assign _11470_ = _11471_ | _11473_ /*27001*/;
assign _11213_ = _11465_ ^ _11472_ /*27004*/;
assign _11479_ = D[49] ^ Q[35] /*27000*/;
assign _11476_ = _10828_ & _11479_ /*26996*/;
assign _11477_ = _10828_ ^ _11479_ /*26999*/;
assign _11478_ = _11470_ & _11477_ /*26997*/;
assign _11475_ = _11476_ | _11478_ /*26995*/;
assign _11214_ = _11470_ ^ _11477_ /*26998*/;
assign _11484_ = D[50] ^ Q[35] /*26994*/;
assign _11481_ = _10829_ & _11484_ /*26990*/;
assign _11482_ = _10829_ ^ _11484_ /*26993*/;
assign _11483_ = _11475_ & _11482_ /*26991*/;
assign _11480_ = _11481_ | _11483_ /*26989*/;
assign _11215_ = _11475_ ^ _11482_ /*26992*/;
assign _11489_ = D[51] ^ Q[35] /*26988*/;
assign _11486_ = _10830_ & _11489_ /*26984*/;
assign _11487_ = _10830_ ^ _11489_ /*26987*/;
assign _11488_ = _11480_ & _11487_ /*26985*/;
assign _11485_ = _11486_ | _11488_ /*26983*/;
assign _11216_ = _11480_ ^ _11487_ /*26986*/;
assign _11494_ = D[52] ^ Q[35] /*26982*/;
assign _11491_ = _10831_ & _11494_ /*26978*/;
assign _11492_ = _10831_ ^ _11494_ /*26981*/;
assign _11493_ = _11485_ & _11492_ /*26979*/;
assign _11490_ = _11491_ | _11493_ /*26977*/;
assign _11217_ = _11485_ ^ _11492_ /*26980*/;
assign _11499_ = D[53] ^ Q[35] /*26976*/;
assign _11496_ = _10832_ & _11499_ /*26972*/;
assign _11497_ = _10832_ ^ _11499_ /*26975*/;
assign _11498_ = _11490_ & _11497_ /*26973*/;
assign _11495_ = _11496_ | _11498_ /*26971*/;
assign _11218_ = _11490_ ^ _11497_ /*26974*/;
assign _11504_ = D[54] ^ Q[35] /*26970*/;
assign _11501_ = _10833_ & _11504_ /*26966*/;
assign _11502_ = _10833_ ^ _11504_ /*26969*/;
assign _11503_ = _11495_ & _11502_ /*26967*/;
assign _11500_ = _11501_ | _11503_ /*26965*/;
assign _11219_ = _11495_ ^ _11502_ /*26968*/;
assign _11509_ = D[55] ^ Q[35] /*26964*/;
assign _11506_ = _10834_ & _11509_ /*26960*/;
assign _11507_ = _10834_ ^ _11509_ /*26963*/;
assign _11508_ = _11500_ & _11507_ /*26961*/;
assign _11505_ = _11506_ | _11508_ /*26959*/;
assign _11220_ = _11500_ ^ _11507_ /*26962*/;
assign _11514_ = D[56] ^ Q[35] /*26958*/;
assign _11511_ = _10835_ & _11514_ /*26954*/;
assign _11512_ = _10835_ ^ _11514_ /*26957*/;
assign _11513_ = _11505_ & _11512_ /*26955*/;
assign _11510_ = _11511_ | _11513_ /*26953*/;
assign _11221_ = _11505_ ^ _11512_ /*26956*/;
assign _11519_ = D[57] ^ Q[35] /*26952*/;
assign _11516_ = _10836_ & _11519_ /*26948*/;
assign _11517_ = _10836_ ^ _11519_ /*26951*/;
assign _11518_ = _11510_ & _11517_ /*26949*/;
assign _11515_ = _11516_ | _11518_ /*26947*/;
assign _11222_ = _11510_ ^ _11517_ /*26950*/;
assign _11524_ = D[58] ^ Q[35] /*26946*/;
assign _11521_ = _10837_ & _11524_ /*26942*/;
assign _11522_ = _10837_ ^ _11524_ /*26945*/;
assign _11523_ = _11515_ & _11522_ /*26943*/;
assign _11520_ = _11521_ | _11523_ /*26941*/;
assign _11223_ = _11515_ ^ _11522_ /*26944*/;
assign _11529_ = D[59] ^ Q[35] /*26940*/;
assign _11526_ = _10838_ & _11529_ /*26936*/;
assign _11527_ = _10838_ ^ _11529_ /*26939*/;
assign _11528_ = _11520_ & _11527_ /*26937*/;
assign _11525_ = _11526_ | _11528_ /*26935*/;
assign _11224_ = _11520_ ^ _11527_ /*26938*/;
assign _11534_ = D[60] ^ Q[35] /*26934*/;
assign _11531_ = _10839_ & _11534_ /*26930*/;
assign _11532_ = _10839_ ^ _11534_ /*26933*/;
assign _11533_ = _11525_ & _11532_ /*26931*/;
assign _11530_ = _11531_ | _11533_ /*26929*/;
assign _11225_ = _11525_ ^ _11532_ /*26932*/;
assign _11539_ = D[61] ^ Q[35] /*26928*/;
assign _11536_ = _10840_ & _11539_ /*26924*/;
assign _11537_ = _10840_ ^ _11539_ /*26927*/;
assign _11538_ = _11530_ & _11537_ /*26925*/;
assign _11535_ = _11536_ | _11538_ /*26923*/;
assign _11226_ = _11530_ ^ _11537_ /*26926*/;
assign _11544_ = D[62] ^ Q[35] /*26922*/;
assign _11541_ = _10841_ & _11544_ /*26918*/;
assign _11542_ = _10841_ ^ _11544_ /*26921*/;
assign _11543_ = _11535_ & _11542_ /*26919*/;
assign _11540_ = _11541_ | _11543_ /*26917*/;
assign _11227_ = _11535_ ^ _11542_ /*26920*/;
assign _11548_ = zeroWire ^ Q[35] /*26916*/;
assign _11545_ = _10842_ & _11548_ /*26912*/;
assign _11546_ = _10842_ ^ _11548_ /*26915*/;
assign _11547_ = _11540_ & _11546_ /*26913*/;
assign Q[34] = _11545_ | _11547_ /*26911*/;
assign _11228_ = _11540_ ^ _11546_ /*26914*/;
assign _11619_ = D[0] ^ Q[34] /*26525*/;
assign _11616_ = R_0[33] & _11619_ /*26521*/;
assign _11617_ = R_0[33] ^ _11619_ /*26524*/;
assign _11618_ = Q[34] & _11617_ /*26522*/;
assign _11615_ = _11616_ | _11618_ /*26520*/;
assign _11550_ = Q[34] ^ _11617_ /*26523*/;
assign _11624_ = D[1] ^ Q[34] /*26519*/;
assign _11621_ = _11165_ & _11624_ /*26515*/;
assign _11622_ = _11165_ ^ _11624_ /*26518*/;
assign _11623_ = _11615_ & _11622_ /*26516*/;
assign _11620_ = _11621_ | _11623_ /*26514*/;
assign _11551_ = _11615_ ^ _11622_ /*26517*/;
assign _11629_ = D[2] ^ Q[34] /*26513*/;
assign _11626_ = _11166_ & _11629_ /*26509*/;
assign _11627_ = _11166_ ^ _11629_ /*26512*/;
assign _11628_ = _11620_ & _11627_ /*26510*/;
assign _11625_ = _11626_ | _11628_ /*26508*/;
assign _11552_ = _11620_ ^ _11627_ /*26511*/;
assign _11634_ = D[3] ^ Q[34] /*26507*/;
assign _11631_ = _11167_ & _11634_ /*26503*/;
assign _11632_ = _11167_ ^ _11634_ /*26506*/;
assign _11633_ = _11625_ & _11632_ /*26504*/;
assign _11630_ = _11631_ | _11633_ /*26502*/;
assign _11553_ = _11625_ ^ _11632_ /*26505*/;
assign _11639_ = D[4] ^ Q[34] /*26501*/;
assign _11636_ = _11168_ & _11639_ /*26497*/;
assign _11637_ = _11168_ ^ _11639_ /*26500*/;
assign _11638_ = _11630_ & _11637_ /*26498*/;
assign _11635_ = _11636_ | _11638_ /*26496*/;
assign _11554_ = _11630_ ^ _11637_ /*26499*/;
assign _11644_ = D[5] ^ Q[34] /*26495*/;
assign _11641_ = _11169_ & _11644_ /*26491*/;
assign _11642_ = _11169_ ^ _11644_ /*26494*/;
assign _11643_ = _11635_ & _11642_ /*26492*/;
assign _11640_ = _11641_ | _11643_ /*26490*/;
assign _11555_ = _11635_ ^ _11642_ /*26493*/;
assign _11649_ = D[6] ^ Q[34] /*26489*/;
assign _11646_ = _11170_ & _11649_ /*26485*/;
assign _11647_ = _11170_ ^ _11649_ /*26488*/;
assign _11648_ = _11640_ & _11647_ /*26486*/;
assign _11645_ = _11646_ | _11648_ /*26484*/;
assign _11556_ = _11640_ ^ _11647_ /*26487*/;
assign _11654_ = D[7] ^ Q[34] /*26483*/;
assign _11651_ = _11171_ & _11654_ /*26479*/;
assign _11652_ = _11171_ ^ _11654_ /*26482*/;
assign _11653_ = _11645_ & _11652_ /*26480*/;
assign _11650_ = _11651_ | _11653_ /*26478*/;
assign _11557_ = _11645_ ^ _11652_ /*26481*/;
assign _11659_ = D[8] ^ Q[34] /*26477*/;
assign _11656_ = _11172_ & _11659_ /*26473*/;
assign _11657_ = _11172_ ^ _11659_ /*26476*/;
assign _11658_ = _11650_ & _11657_ /*26474*/;
assign _11655_ = _11656_ | _11658_ /*26472*/;
assign _11558_ = _11650_ ^ _11657_ /*26475*/;
assign _11664_ = D[9] ^ Q[34] /*26471*/;
assign _11661_ = _11173_ & _11664_ /*26467*/;
assign _11662_ = _11173_ ^ _11664_ /*26470*/;
assign _11663_ = _11655_ & _11662_ /*26468*/;
assign _11660_ = _11661_ | _11663_ /*26466*/;
assign _11559_ = _11655_ ^ _11662_ /*26469*/;
assign _11669_ = D[10] ^ Q[34] /*26465*/;
assign _11666_ = _11174_ & _11669_ /*26461*/;
assign _11667_ = _11174_ ^ _11669_ /*26464*/;
assign _11668_ = _11660_ & _11667_ /*26462*/;
assign _11665_ = _11666_ | _11668_ /*26460*/;
assign _11560_ = _11660_ ^ _11667_ /*26463*/;
assign _11674_ = D[11] ^ Q[34] /*26459*/;
assign _11671_ = _11175_ & _11674_ /*26455*/;
assign _11672_ = _11175_ ^ _11674_ /*26458*/;
assign _11673_ = _11665_ & _11672_ /*26456*/;
assign _11670_ = _11671_ | _11673_ /*26454*/;
assign _11561_ = _11665_ ^ _11672_ /*26457*/;
assign _11679_ = D[12] ^ Q[34] /*26453*/;
assign _11676_ = _11176_ & _11679_ /*26449*/;
assign _11677_ = _11176_ ^ _11679_ /*26452*/;
assign _11678_ = _11670_ & _11677_ /*26450*/;
assign _11675_ = _11676_ | _11678_ /*26448*/;
assign _11562_ = _11670_ ^ _11677_ /*26451*/;
assign _11684_ = D[13] ^ Q[34] /*26447*/;
assign _11681_ = _11177_ & _11684_ /*26443*/;
assign _11682_ = _11177_ ^ _11684_ /*26446*/;
assign _11683_ = _11675_ & _11682_ /*26444*/;
assign _11680_ = _11681_ | _11683_ /*26442*/;
assign _11563_ = _11675_ ^ _11682_ /*26445*/;
assign _11689_ = D[14] ^ Q[34] /*26441*/;
assign _11686_ = _11178_ & _11689_ /*26437*/;
assign _11687_ = _11178_ ^ _11689_ /*26440*/;
assign _11688_ = _11680_ & _11687_ /*26438*/;
assign _11685_ = _11686_ | _11688_ /*26436*/;
assign _11564_ = _11680_ ^ _11687_ /*26439*/;
assign _11694_ = D[15] ^ Q[34] /*26435*/;
assign _11691_ = _11179_ & _11694_ /*26431*/;
assign _11692_ = _11179_ ^ _11694_ /*26434*/;
assign _11693_ = _11685_ & _11692_ /*26432*/;
assign _11690_ = _11691_ | _11693_ /*26430*/;
assign _11565_ = _11685_ ^ _11692_ /*26433*/;
assign _11699_ = D[16] ^ Q[34] /*26429*/;
assign _11696_ = _11180_ & _11699_ /*26425*/;
assign _11697_ = _11180_ ^ _11699_ /*26428*/;
assign _11698_ = _11690_ & _11697_ /*26426*/;
assign _11695_ = _11696_ | _11698_ /*26424*/;
assign _11566_ = _11690_ ^ _11697_ /*26427*/;
assign _11704_ = D[17] ^ Q[34] /*26423*/;
assign _11701_ = _11181_ & _11704_ /*26419*/;
assign _11702_ = _11181_ ^ _11704_ /*26422*/;
assign _11703_ = _11695_ & _11702_ /*26420*/;
assign _11700_ = _11701_ | _11703_ /*26418*/;
assign _11567_ = _11695_ ^ _11702_ /*26421*/;
assign _11709_ = D[18] ^ Q[34] /*26417*/;
assign _11706_ = _11182_ & _11709_ /*26413*/;
assign _11707_ = _11182_ ^ _11709_ /*26416*/;
assign _11708_ = _11700_ & _11707_ /*26414*/;
assign _11705_ = _11706_ | _11708_ /*26412*/;
assign _11568_ = _11700_ ^ _11707_ /*26415*/;
assign _11714_ = D[19] ^ Q[34] /*26411*/;
assign _11711_ = _11183_ & _11714_ /*26407*/;
assign _11712_ = _11183_ ^ _11714_ /*26410*/;
assign _11713_ = _11705_ & _11712_ /*26408*/;
assign _11710_ = _11711_ | _11713_ /*26406*/;
assign _11569_ = _11705_ ^ _11712_ /*26409*/;
assign _11719_ = D[20] ^ Q[34] /*26405*/;
assign _11716_ = _11184_ & _11719_ /*26401*/;
assign _11717_ = _11184_ ^ _11719_ /*26404*/;
assign _11718_ = _11710_ & _11717_ /*26402*/;
assign _11715_ = _11716_ | _11718_ /*26400*/;
assign _11570_ = _11710_ ^ _11717_ /*26403*/;
assign _11724_ = D[21] ^ Q[34] /*26399*/;
assign _11721_ = _11185_ & _11724_ /*26395*/;
assign _11722_ = _11185_ ^ _11724_ /*26398*/;
assign _11723_ = _11715_ & _11722_ /*26396*/;
assign _11720_ = _11721_ | _11723_ /*26394*/;
assign _11571_ = _11715_ ^ _11722_ /*26397*/;
assign _11729_ = D[22] ^ Q[34] /*26393*/;
assign _11726_ = _11186_ & _11729_ /*26389*/;
assign _11727_ = _11186_ ^ _11729_ /*26392*/;
assign _11728_ = _11720_ & _11727_ /*26390*/;
assign _11725_ = _11726_ | _11728_ /*26388*/;
assign _11572_ = _11720_ ^ _11727_ /*26391*/;
assign _11734_ = D[23] ^ Q[34] /*26387*/;
assign _11731_ = _11187_ & _11734_ /*26383*/;
assign _11732_ = _11187_ ^ _11734_ /*26386*/;
assign _11733_ = _11725_ & _11732_ /*26384*/;
assign _11730_ = _11731_ | _11733_ /*26382*/;
assign _11573_ = _11725_ ^ _11732_ /*26385*/;
assign _11739_ = D[24] ^ Q[34] /*26381*/;
assign _11736_ = _11188_ & _11739_ /*26377*/;
assign _11737_ = _11188_ ^ _11739_ /*26380*/;
assign _11738_ = _11730_ & _11737_ /*26378*/;
assign _11735_ = _11736_ | _11738_ /*26376*/;
assign _11574_ = _11730_ ^ _11737_ /*26379*/;
assign _11744_ = D[25] ^ Q[34] /*26375*/;
assign _11741_ = _11189_ & _11744_ /*26371*/;
assign _11742_ = _11189_ ^ _11744_ /*26374*/;
assign _11743_ = _11735_ & _11742_ /*26372*/;
assign _11740_ = _11741_ | _11743_ /*26370*/;
assign _11575_ = _11735_ ^ _11742_ /*26373*/;
assign _11749_ = D[26] ^ Q[34] /*26369*/;
assign _11746_ = _11190_ & _11749_ /*26365*/;
assign _11747_ = _11190_ ^ _11749_ /*26368*/;
assign _11748_ = _11740_ & _11747_ /*26366*/;
assign _11745_ = _11746_ | _11748_ /*26364*/;
assign _11576_ = _11740_ ^ _11747_ /*26367*/;
assign _11754_ = D[27] ^ Q[34] /*26363*/;
assign _11751_ = _11191_ & _11754_ /*26359*/;
assign _11752_ = _11191_ ^ _11754_ /*26362*/;
assign _11753_ = _11745_ & _11752_ /*26360*/;
assign _11750_ = _11751_ | _11753_ /*26358*/;
assign _11577_ = _11745_ ^ _11752_ /*26361*/;
assign _11759_ = D[28] ^ Q[34] /*26357*/;
assign _11756_ = _11192_ & _11759_ /*26353*/;
assign _11757_ = _11192_ ^ _11759_ /*26356*/;
assign _11758_ = _11750_ & _11757_ /*26354*/;
assign _11755_ = _11756_ | _11758_ /*26352*/;
assign _11578_ = _11750_ ^ _11757_ /*26355*/;
assign _11764_ = D[29] ^ Q[34] /*26351*/;
assign _11761_ = _11193_ & _11764_ /*26347*/;
assign _11762_ = _11193_ ^ _11764_ /*26350*/;
assign _11763_ = _11755_ & _11762_ /*26348*/;
assign _11760_ = _11761_ | _11763_ /*26346*/;
assign _11579_ = _11755_ ^ _11762_ /*26349*/;
assign _11769_ = D[30] ^ Q[34] /*26345*/;
assign _11766_ = _11194_ & _11769_ /*26341*/;
assign _11767_ = _11194_ ^ _11769_ /*26344*/;
assign _11768_ = _11760_ & _11767_ /*26342*/;
assign _11765_ = _11766_ | _11768_ /*26340*/;
assign _11580_ = _11760_ ^ _11767_ /*26343*/;
assign _11774_ = D[31] ^ Q[34] /*26339*/;
assign _11771_ = _11195_ & _11774_ /*26335*/;
assign _11772_ = _11195_ ^ _11774_ /*26338*/;
assign _11773_ = _11765_ & _11772_ /*26336*/;
assign _11770_ = _11771_ | _11773_ /*26334*/;
assign _11581_ = _11765_ ^ _11772_ /*26337*/;
assign _11779_ = D[32] ^ Q[34] /*26333*/;
assign _11776_ = _11196_ & _11779_ /*26329*/;
assign _11777_ = _11196_ ^ _11779_ /*26332*/;
assign _11778_ = _11770_ & _11777_ /*26330*/;
assign _11775_ = _11776_ | _11778_ /*26328*/;
assign _11582_ = _11770_ ^ _11777_ /*26331*/;
assign _11784_ = D[33] ^ Q[34] /*26327*/;
assign _11781_ = _11197_ & _11784_ /*26323*/;
assign _11782_ = _11197_ ^ _11784_ /*26326*/;
assign _11783_ = _11775_ & _11782_ /*26324*/;
assign _11780_ = _11781_ | _11783_ /*26322*/;
assign _11583_ = _11775_ ^ _11782_ /*26325*/;
assign _11789_ = D[34] ^ Q[34] /*26321*/;
assign _11786_ = _11198_ & _11789_ /*26317*/;
assign _11787_ = _11198_ ^ _11789_ /*26320*/;
assign _11788_ = _11780_ & _11787_ /*26318*/;
assign _11785_ = _11786_ | _11788_ /*26316*/;
assign _11584_ = _11780_ ^ _11787_ /*26319*/;
assign _11794_ = D[35] ^ Q[34] /*26315*/;
assign _11791_ = _11199_ & _11794_ /*26311*/;
assign _11792_ = _11199_ ^ _11794_ /*26314*/;
assign _11793_ = _11785_ & _11792_ /*26312*/;
assign _11790_ = _11791_ | _11793_ /*26310*/;
assign _11585_ = _11785_ ^ _11792_ /*26313*/;
assign _11799_ = D[36] ^ Q[34] /*26309*/;
assign _11796_ = _11200_ & _11799_ /*26305*/;
assign _11797_ = _11200_ ^ _11799_ /*26308*/;
assign _11798_ = _11790_ & _11797_ /*26306*/;
assign _11795_ = _11796_ | _11798_ /*26304*/;
assign _11586_ = _11790_ ^ _11797_ /*26307*/;
assign _11804_ = D[37] ^ Q[34] /*26303*/;
assign _11801_ = _11201_ & _11804_ /*26299*/;
assign _11802_ = _11201_ ^ _11804_ /*26302*/;
assign _11803_ = _11795_ & _11802_ /*26300*/;
assign _11800_ = _11801_ | _11803_ /*26298*/;
assign _11587_ = _11795_ ^ _11802_ /*26301*/;
assign _11809_ = D[38] ^ Q[34] /*26297*/;
assign _11806_ = _11202_ & _11809_ /*26293*/;
assign _11807_ = _11202_ ^ _11809_ /*26296*/;
assign _11808_ = _11800_ & _11807_ /*26294*/;
assign _11805_ = _11806_ | _11808_ /*26292*/;
assign _11588_ = _11800_ ^ _11807_ /*26295*/;
assign _11814_ = D[39] ^ Q[34] /*26291*/;
assign _11811_ = _11203_ & _11814_ /*26287*/;
assign _11812_ = _11203_ ^ _11814_ /*26290*/;
assign _11813_ = _11805_ & _11812_ /*26288*/;
assign _11810_ = _11811_ | _11813_ /*26286*/;
assign _11589_ = _11805_ ^ _11812_ /*26289*/;
assign _11819_ = D[40] ^ Q[34] /*26285*/;
assign _11816_ = _11204_ & _11819_ /*26281*/;
assign _11817_ = _11204_ ^ _11819_ /*26284*/;
assign _11818_ = _11810_ & _11817_ /*26282*/;
assign _11815_ = _11816_ | _11818_ /*26280*/;
assign _11590_ = _11810_ ^ _11817_ /*26283*/;
assign _11824_ = D[41] ^ Q[34] /*26279*/;
assign _11821_ = _11205_ & _11824_ /*26275*/;
assign _11822_ = _11205_ ^ _11824_ /*26278*/;
assign _11823_ = _11815_ & _11822_ /*26276*/;
assign _11820_ = _11821_ | _11823_ /*26274*/;
assign _11591_ = _11815_ ^ _11822_ /*26277*/;
assign _11829_ = D[42] ^ Q[34] /*26273*/;
assign _11826_ = _11206_ & _11829_ /*26269*/;
assign _11827_ = _11206_ ^ _11829_ /*26272*/;
assign _11828_ = _11820_ & _11827_ /*26270*/;
assign _11825_ = _11826_ | _11828_ /*26268*/;
assign _11592_ = _11820_ ^ _11827_ /*26271*/;
assign _11834_ = D[43] ^ Q[34] /*26267*/;
assign _11831_ = _11207_ & _11834_ /*26263*/;
assign _11832_ = _11207_ ^ _11834_ /*26266*/;
assign _11833_ = _11825_ & _11832_ /*26264*/;
assign _11830_ = _11831_ | _11833_ /*26262*/;
assign _11593_ = _11825_ ^ _11832_ /*26265*/;
assign _11839_ = D[44] ^ Q[34] /*26261*/;
assign _11836_ = _11208_ & _11839_ /*26257*/;
assign _11837_ = _11208_ ^ _11839_ /*26260*/;
assign _11838_ = _11830_ & _11837_ /*26258*/;
assign _11835_ = _11836_ | _11838_ /*26256*/;
assign _11594_ = _11830_ ^ _11837_ /*26259*/;
assign _11844_ = D[45] ^ Q[34] /*26255*/;
assign _11841_ = _11209_ & _11844_ /*26251*/;
assign _11842_ = _11209_ ^ _11844_ /*26254*/;
assign _11843_ = _11835_ & _11842_ /*26252*/;
assign _11840_ = _11841_ | _11843_ /*26250*/;
assign _11595_ = _11835_ ^ _11842_ /*26253*/;
assign _11849_ = D[46] ^ Q[34] /*26249*/;
assign _11846_ = _11210_ & _11849_ /*26245*/;
assign _11847_ = _11210_ ^ _11849_ /*26248*/;
assign _11848_ = _11840_ & _11847_ /*26246*/;
assign _11845_ = _11846_ | _11848_ /*26244*/;
assign _11596_ = _11840_ ^ _11847_ /*26247*/;
assign _11854_ = D[47] ^ Q[34] /*26243*/;
assign _11851_ = _11211_ & _11854_ /*26239*/;
assign _11852_ = _11211_ ^ _11854_ /*26242*/;
assign _11853_ = _11845_ & _11852_ /*26240*/;
assign _11850_ = _11851_ | _11853_ /*26238*/;
assign _11597_ = _11845_ ^ _11852_ /*26241*/;
assign _11859_ = D[48] ^ Q[34] /*26237*/;
assign _11856_ = _11212_ & _11859_ /*26233*/;
assign _11857_ = _11212_ ^ _11859_ /*26236*/;
assign _11858_ = _11850_ & _11857_ /*26234*/;
assign _11855_ = _11856_ | _11858_ /*26232*/;
assign _11598_ = _11850_ ^ _11857_ /*26235*/;
assign _11864_ = D[49] ^ Q[34] /*26231*/;
assign _11861_ = _11213_ & _11864_ /*26227*/;
assign _11862_ = _11213_ ^ _11864_ /*26230*/;
assign _11863_ = _11855_ & _11862_ /*26228*/;
assign _11860_ = _11861_ | _11863_ /*26226*/;
assign _11599_ = _11855_ ^ _11862_ /*26229*/;
assign _11869_ = D[50] ^ Q[34] /*26225*/;
assign _11866_ = _11214_ & _11869_ /*26221*/;
assign _11867_ = _11214_ ^ _11869_ /*26224*/;
assign _11868_ = _11860_ & _11867_ /*26222*/;
assign _11865_ = _11866_ | _11868_ /*26220*/;
assign _11600_ = _11860_ ^ _11867_ /*26223*/;
assign _11874_ = D[51] ^ Q[34] /*26219*/;
assign _11871_ = _11215_ & _11874_ /*26215*/;
assign _11872_ = _11215_ ^ _11874_ /*26218*/;
assign _11873_ = _11865_ & _11872_ /*26216*/;
assign _11870_ = _11871_ | _11873_ /*26214*/;
assign _11601_ = _11865_ ^ _11872_ /*26217*/;
assign _11879_ = D[52] ^ Q[34] /*26213*/;
assign _11876_ = _11216_ & _11879_ /*26209*/;
assign _11877_ = _11216_ ^ _11879_ /*26212*/;
assign _11878_ = _11870_ & _11877_ /*26210*/;
assign _11875_ = _11876_ | _11878_ /*26208*/;
assign _11602_ = _11870_ ^ _11877_ /*26211*/;
assign _11884_ = D[53] ^ Q[34] /*26207*/;
assign _11881_ = _11217_ & _11884_ /*26203*/;
assign _11882_ = _11217_ ^ _11884_ /*26206*/;
assign _11883_ = _11875_ & _11882_ /*26204*/;
assign _11880_ = _11881_ | _11883_ /*26202*/;
assign _11603_ = _11875_ ^ _11882_ /*26205*/;
assign _11889_ = D[54] ^ Q[34] /*26201*/;
assign _11886_ = _11218_ & _11889_ /*26197*/;
assign _11887_ = _11218_ ^ _11889_ /*26200*/;
assign _11888_ = _11880_ & _11887_ /*26198*/;
assign _11885_ = _11886_ | _11888_ /*26196*/;
assign _11604_ = _11880_ ^ _11887_ /*26199*/;
assign _11894_ = D[55] ^ Q[34] /*26195*/;
assign _11891_ = _11219_ & _11894_ /*26191*/;
assign _11892_ = _11219_ ^ _11894_ /*26194*/;
assign _11893_ = _11885_ & _11892_ /*26192*/;
assign _11890_ = _11891_ | _11893_ /*26190*/;
assign _11605_ = _11885_ ^ _11892_ /*26193*/;
assign _11899_ = D[56] ^ Q[34] /*26189*/;
assign _11896_ = _11220_ & _11899_ /*26185*/;
assign _11897_ = _11220_ ^ _11899_ /*26188*/;
assign _11898_ = _11890_ & _11897_ /*26186*/;
assign _11895_ = _11896_ | _11898_ /*26184*/;
assign _11606_ = _11890_ ^ _11897_ /*26187*/;
assign _11904_ = D[57] ^ Q[34] /*26183*/;
assign _11901_ = _11221_ & _11904_ /*26179*/;
assign _11902_ = _11221_ ^ _11904_ /*26182*/;
assign _11903_ = _11895_ & _11902_ /*26180*/;
assign _11900_ = _11901_ | _11903_ /*26178*/;
assign _11607_ = _11895_ ^ _11902_ /*26181*/;
assign _11909_ = D[58] ^ Q[34] /*26177*/;
assign _11906_ = _11222_ & _11909_ /*26173*/;
assign _11907_ = _11222_ ^ _11909_ /*26176*/;
assign _11908_ = _11900_ & _11907_ /*26174*/;
assign _11905_ = _11906_ | _11908_ /*26172*/;
assign _11608_ = _11900_ ^ _11907_ /*26175*/;
assign _11914_ = D[59] ^ Q[34] /*26171*/;
assign _11911_ = _11223_ & _11914_ /*26167*/;
assign _11912_ = _11223_ ^ _11914_ /*26170*/;
assign _11913_ = _11905_ & _11912_ /*26168*/;
assign _11910_ = _11911_ | _11913_ /*26166*/;
assign _11609_ = _11905_ ^ _11912_ /*26169*/;
assign _11919_ = D[60] ^ Q[34] /*26165*/;
assign _11916_ = _11224_ & _11919_ /*26161*/;
assign _11917_ = _11224_ ^ _11919_ /*26164*/;
assign _11918_ = _11910_ & _11917_ /*26162*/;
assign _11915_ = _11916_ | _11918_ /*26160*/;
assign _11610_ = _11910_ ^ _11917_ /*26163*/;
assign _11924_ = D[61] ^ Q[34] /*26159*/;
assign _11921_ = _11225_ & _11924_ /*26155*/;
assign _11922_ = _11225_ ^ _11924_ /*26158*/;
assign _11923_ = _11915_ & _11922_ /*26156*/;
assign _11920_ = _11921_ | _11923_ /*26154*/;
assign _11611_ = _11915_ ^ _11922_ /*26157*/;
assign _11929_ = D[62] ^ Q[34] /*26153*/;
assign _11926_ = _11226_ & _11929_ /*26149*/;
assign _11927_ = _11226_ ^ _11929_ /*26152*/;
assign _11928_ = _11920_ & _11927_ /*26150*/;
assign _11925_ = _11926_ | _11928_ /*26148*/;
assign _11612_ = _11920_ ^ _11927_ /*26151*/;
assign _11933_ = zeroWire ^ Q[34] /*26147*/;
assign _11930_ = _11227_ & _11933_ /*26143*/;
assign _11931_ = _11227_ ^ _11933_ /*26146*/;
assign _11932_ = _11925_ & _11931_ /*26144*/;
assign Q[33] = _11930_ | _11932_ /*26142*/;
assign _11613_ = _11925_ ^ _11931_ /*26145*/;
assign _12004_ = D[0] ^ Q[33] /*25756*/;
assign _12001_ = R_0[32] & _12004_ /*25752*/;
assign _12002_ = R_0[32] ^ _12004_ /*25755*/;
assign _12003_ = Q[33] & _12002_ /*25753*/;
assign _12000_ = _12001_ | _12003_ /*25751*/;
assign _11935_ = Q[33] ^ _12002_ /*25754*/;
assign _12009_ = D[1] ^ Q[33] /*25750*/;
assign _12006_ = _11550_ & _12009_ /*25746*/;
assign _12007_ = _11550_ ^ _12009_ /*25749*/;
assign _12008_ = _12000_ & _12007_ /*25747*/;
assign _12005_ = _12006_ | _12008_ /*25745*/;
assign _11936_ = _12000_ ^ _12007_ /*25748*/;
assign _12014_ = D[2] ^ Q[33] /*25744*/;
assign _12011_ = _11551_ & _12014_ /*25740*/;
assign _12012_ = _11551_ ^ _12014_ /*25743*/;
assign _12013_ = _12005_ & _12012_ /*25741*/;
assign _12010_ = _12011_ | _12013_ /*25739*/;
assign _11937_ = _12005_ ^ _12012_ /*25742*/;
assign _12019_ = D[3] ^ Q[33] /*25738*/;
assign _12016_ = _11552_ & _12019_ /*25734*/;
assign _12017_ = _11552_ ^ _12019_ /*25737*/;
assign _12018_ = _12010_ & _12017_ /*25735*/;
assign _12015_ = _12016_ | _12018_ /*25733*/;
assign _11938_ = _12010_ ^ _12017_ /*25736*/;
assign _12024_ = D[4] ^ Q[33] /*25732*/;
assign _12021_ = _11553_ & _12024_ /*25728*/;
assign _12022_ = _11553_ ^ _12024_ /*25731*/;
assign _12023_ = _12015_ & _12022_ /*25729*/;
assign _12020_ = _12021_ | _12023_ /*25727*/;
assign _11939_ = _12015_ ^ _12022_ /*25730*/;
assign _12029_ = D[5] ^ Q[33] /*25726*/;
assign _12026_ = _11554_ & _12029_ /*25722*/;
assign _12027_ = _11554_ ^ _12029_ /*25725*/;
assign _12028_ = _12020_ & _12027_ /*25723*/;
assign _12025_ = _12026_ | _12028_ /*25721*/;
assign _11940_ = _12020_ ^ _12027_ /*25724*/;
assign _12034_ = D[6] ^ Q[33] /*25720*/;
assign _12031_ = _11555_ & _12034_ /*25716*/;
assign _12032_ = _11555_ ^ _12034_ /*25719*/;
assign _12033_ = _12025_ & _12032_ /*25717*/;
assign _12030_ = _12031_ | _12033_ /*25715*/;
assign _11941_ = _12025_ ^ _12032_ /*25718*/;
assign _12039_ = D[7] ^ Q[33] /*25714*/;
assign _12036_ = _11556_ & _12039_ /*25710*/;
assign _12037_ = _11556_ ^ _12039_ /*25713*/;
assign _12038_ = _12030_ & _12037_ /*25711*/;
assign _12035_ = _12036_ | _12038_ /*25709*/;
assign _11942_ = _12030_ ^ _12037_ /*25712*/;
assign _12044_ = D[8] ^ Q[33] /*25708*/;
assign _12041_ = _11557_ & _12044_ /*25704*/;
assign _12042_ = _11557_ ^ _12044_ /*25707*/;
assign _12043_ = _12035_ & _12042_ /*25705*/;
assign _12040_ = _12041_ | _12043_ /*25703*/;
assign _11943_ = _12035_ ^ _12042_ /*25706*/;
assign _12049_ = D[9] ^ Q[33] /*25702*/;
assign _12046_ = _11558_ & _12049_ /*25698*/;
assign _12047_ = _11558_ ^ _12049_ /*25701*/;
assign _12048_ = _12040_ & _12047_ /*25699*/;
assign _12045_ = _12046_ | _12048_ /*25697*/;
assign _11944_ = _12040_ ^ _12047_ /*25700*/;
assign _12054_ = D[10] ^ Q[33] /*25696*/;
assign _12051_ = _11559_ & _12054_ /*25692*/;
assign _12052_ = _11559_ ^ _12054_ /*25695*/;
assign _12053_ = _12045_ & _12052_ /*25693*/;
assign _12050_ = _12051_ | _12053_ /*25691*/;
assign _11945_ = _12045_ ^ _12052_ /*25694*/;
assign _12059_ = D[11] ^ Q[33] /*25690*/;
assign _12056_ = _11560_ & _12059_ /*25686*/;
assign _12057_ = _11560_ ^ _12059_ /*25689*/;
assign _12058_ = _12050_ & _12057_ /*25687*/;
assign _12055_ = _12056_ | _12058_ /*25685*/;
assign _11946_ = _12050_ ^ _12057_ /*25688*/;
assign _12064_ = D[12] ^ Q[33] /*25684*/;
assign _12061_ = _11561_ & _12064_ /*25680*/;
assign _12062_ = _11561_ ^ _12064_ /*25683*/;
assign _12063_ = _12055_ & _12062_ /*25681*/;
assign _12060_ = _12061_ | _12063_ /*25679*/;
assign _11947_ = _12055_ ^ _12062_ /*25682*/;
assign _12069_ = D[13] ^ Q[33] /*25678*/;
assign _12066_ = _11562_ & _12069_ /*25674*/;
assign _12067_ = _11562_ ^ _12069_ /*25677*/;
assign _12068_ = _12060_ & _12067_ /*25675*/;
assign _12065_ = _12066_ | _12068_ /*25673*/;
assign _11948_ = _12060_ ^ _12067_ /*25676*/;
assign _12074_ = D[14] ^ Q[33] /*25672*/;
assign _12071_ = _11563_ & _12074_ /*25668*/;
assign _12072_ = _11563_ ^ _12074_ /*25671*/;
assign _12073_ = _12065_ & _12072_ /*25669*/;
assign _12070_ = _12071_ | _12073_ /*25667*/;
assign _11949_ = _12065_ ^ _12072_ /*25670*/;
assign _12079_ = D[15] ^ Q[33] /*25666*/;
assign _12076_ = _11564_ & _12079_ /*25662*/;
assign _12077_ = _11564_ ^ _12079_ /*25665*/;
assign _12078_ = _12070_ & _12077_ /*25663*/;
assign _12075_ = _12076_ | _12078_ /*25661*/;
assign _11950_ = _12070_ ^ _12077_ /*25664*/;
assign _12084_ = D[16] ^ Q[33] /*25660*/;
assign _12081_ = _11565_ & _12084_ /*25656*/;
assign _12082_ = _11565_ ^ _12084_ /*25659*/;
assign _12083_ = _12075_ & _12082_ /*25657*/;
assign _12080_ = _12081_ | _12083_ /*25655*/;
assign _11951_ = _12075_ ^ _12082_ /*25658*/;
assign _12089_ = D[17] ^ Q[33] /*25654*/;
assign _12086_ = _11566_ & _12089_ /*25650*/;
assign _12087_ = _11566_ ^ _12089_ /*25653*/;
assign _12088_ = _12080_ & _12087_ /*25651*/;
assign _12085_ = _12086_ | _12088_ /*25649*/;
assign _11952_ = _12080_ ^ _12087_ /*25652*/;
assign _12094_ = D[18] ^ Q[33] /*25648*/;
assign _12091_ = _11567_ & _12094_ /*25644*/;
assign _12092_ = _11567_ ^ _12094_ /*25647*/;
assign _12093_ = _12085_ & _12092_ /*25645*/;
assign _12090_ = _12091_ | _12093_ /*25643*/;
assign _11953_ = _12085_ ^ _12092_ /*25646*/;
assign _12099_ = D[19] ^ Q[33] /*25642*/;
assign _12096_ = _11568_ & _12099_ /*25638*/;
assign _12097_ = _11568_ ^ _12099_ /*25641*/;
assign _12098_ = _12090_ & _12097_ /*25639*/;
assign _12095_ = _12096_ | _12098_ /*25637*/;
assign _11954_ = _12090_ ^ _12097_ /*25640*/;
assign _12104_ = D[20] ^ Q[33] /*25636*/;
assign _12101_ = _11569_ & _12104_ /*25632*/;
assign _12102_ = _11569_ ^ _12104_ /*25635*/;
assign _12103_ = _12095_ & _12102_ /*25633*/;
assign _12100_ = _12101_ | _12103_ /*25631*/;
assign _11955_ = _12095_ ^ _12102_ /*25634*/;
assign _12109_ = D[21] ^ Q[33] /*25630*/;
assign _12106_ = _11570_ & _12109_ /*25626*/;
assign _12107_ = _11570_ ^ _12109_ /*25629*/;
assign _12108_ = _12100_ & _12107_ /*25627*/;
assign _12105_ = _12106_ | _12108_ /*25625*/;
assign _11956_ = _12100_ ^ _12107_ /*25628*/;
assign _12114_ = D[22] ^ Q[33] /*25624*/;
assign _12111_ = _11571_ & _12114_ /*25620*/;
assign _12112_ = _11571_ ^ _12114_ /*25623*/;
assign _12113_ = _12105_ & _12112_ /*25621*/;
assign _12110_ = _12111_ | _12113_ /*25619*/;
assign _11957_ = _12105_ ^ _12112_ /*25622*/;
assign _12119_ = D[23] ^ Q[33] /*25618*/;
assign _12116_ = _11572_ & _12119_ /*25614*/;
assign _12117_ = _11572_ ^ _12119_ /*25617*/;
assign _12118_ = _12110_ & _12117_ /*25615*/;
assign _12115_ = _12116_ | _12118_ /*25613*/;
assign _11958_ = _12110_ ^ _12117_ /*25616*/;
assign _12124_ = D[24] ^ Q[33] /*25612*/;
assign _12121_ = _11573_ & _12124_ /*25608*/;
assign _12122_ = _11573_ ^ _12124_ /*25611*/;
assign _12123_ = _12115_ & _12122_ /*25609*/;
assign _12120_ = _12121_ | _12123_ /*25607*/;
assign _11959_ = _12115_ ^ _12122_ /*25610*/;
assign _12129_ = D[25] ^ Q[33] /*25606*/;
assign _12126_ = _11574_ & _12129_ /*25602*/;
assign _12127_ = _11574_ ^ _12129_ /*25605*/;
assign _12128_ = _12120_ & _12127_ /*25603*/;
assign _12125_ = _12126_ | _12128_ /*25601*/;
assign _11960_ = _12120_ ^ _12127_ /*25604*/;
assign _12134_ = D[26] ^ Q[33] /*25600*/;
assign _12131_ = _11575_ & _12134_ /*25596*/;
assign _12132_ = _11575_ ^ _12134_ /*25599*/;
assign _12133_ = _12125_ & _12132_ /*25597*/;
assign _12130_ = _12131_ | _12133_ /*25595*/;
assign _11961_ = _12125_ ^ _12132_ /*25598*/;
assign _12139_ = D[27] ^ Q[33] /*25594*/;
assign _12136_ = _11576_ & _12139_ /*25590*/;
assign _12137_ = _11576_ ^ _12139_ /*25593*/;
assign _12138_ = _12130_ & _12137_ /*25591*/;
assign _12135_ = _12136_ | _12138_ /*25589*/;
assign _11962_ = _12130_ ^ _12137_ /*25592*/;
assign _12144_ = D[28] ^ Q[33] /*25588*/;
assign _12141_ = _11577_ & _12144_ /*25584*/;
assign _12142_ = _11577_ ^ _12144_ /*25587*/;
assign _12143_ = _12135_ & _12142_ /*25585*/;
assign _12140_ = _12141_ | _12143_ /*25583*/;
assign _11963_ = _12135_ ^ _12142_ /*25586*/;
assign _12149_ = D[29] ^ Q[33] /*25582*/;
assign _12146_ = _11578_ & _12149_ /*25578*/;
assign _12147_ = _11578_ ^ _12149_ /*25581*/;
assign _12148_ = _12140_ & _12147_ /*25579*/;
assign _12145_ = _12146_ | _12148_ /*25577*/;
assign _11964_ = _12140_ ^ _12147_ /*25580*/;
assign _12154_ = D[30] ^ Q[33] /*25576*/;
assign _12151_ = _11579_ & _12154_ /*25572*/;
assign _12152_ = _11579_ ^ _12154_ /*25575*/;
assign _12153_ = _12145_ & _12152_ /*25573*/;
assign _12150_ = _12151_ | _12153_ /*25571*/;
assign _11965_ = _12145_ ^ _12152_ /*25574*/;
assign _12159_ = D[31] ^ Q[33] /*25570*/;
assign _12156_ = _11580_ & _12159_ /*25566*/;
assign _12157_ = _11580_ ^ _12159_ /*25569*/;
assign _12158_ = _12150_ & _12157_ /*25567*/;
assign _12155_ = _12156_ | _12158_ /*25565*/;
assign _11966_ = _12150_ ^ _12157_ /*25568*/;
assign _12164_ = D[32] ^ Q[33] /*25564*/;
assign _12161_ = _11581_ & _12164_ /*25560*/;
assign _12162_ = _11581_ ^ _12164_ /*25563*/;
assign _12163_ = _12155_ & _12162_ /*25561*/;
assign _12160_ = _12161_ | _12163_ /*25559*/;
assign _11967_ = _12155_ ^ _12162_ /*25562*/;
assign _12169_ = D[33] ^ Q[33] /*25558*/;
assign _12166_ = _11582_ & _12169_ /*25554*/;
assign _12167_ = _11582_ ^ _12169_ /*25557*/;
assign _12168_ = _12160_ & _12167_ /*25555*/;
assign _12165_ = _12166_ | _12168_ /*25553*/;
assign _11968_ = _12160_ ^ _12167_ /*25556*/;
assign _12174_ = D[34] ^ Q[33] /*25552*/;
assign _12171_ = _11583_ & _12174_ /*25548*/;
assign _12172_ = _11583_ ^ _12174_ /*25551*/;
assign _12173_ = _12165_ & _12172_ /*25549*/;
assign _12170_ = _12171_ | _12173_ /*25547*/;
assign _11969_ = _12165_ ^ _12172_ /*25550*/;
assign _12179_ = D[35] ^ Q[33] /*25546*/;
assign _12176_ = _11584_ & _12179_ /*25542*/;
assign _12177_ = _11584_ ^ _12179_ /*25545*/;
assign _12178_ = _12170_ & _12177_ /*25543*/;
assign _12175_ = _12176_ | _12178_ /*25541*/;
assign _11970_ = _12170_ ^ _12177_ /*25544*/;
assign _12184_ = D[36] ^ Q[33] /*25540*/;
assign _12181_ = _11585_ & _12184_ /*25536*/;
assign _12182_ = _11585_ ^ _12184_ /*25539*/;
assign _12183_ = _12175_ & _12182_ /*25537*/;
assign _12180_ = _12181_ | _12183_ /*25535*/;
assign _11971_ = _12175_ ^ _12182_ /*25538*/;
assign _12189_ = D[37] ^ Q[33] /*25534*/;
assign _12186_ = _11586_ & _12189_ /*25530*/;
assign _12187_ = _11586_ ^ _12189_ /*25533*/;
assign _12188_ = _12180_ & _12187_ /*25531*/;
assign _12185_ = _12186_ | _12188_ /*25529*/;
assign _11972_ = _12180_ ^ _12187_ /*25532*/;
assign _12194_ = D[38] ^ Q[33] /*25528*/;
assign _12191_ = _11587_ & _12194_ /*25524*/;
assign _12192_ = _11587_ ^ _12194_ /*25527*/;
assign _12193_ = _12185_ & _12192_ /*25525*/;
assign _12190_ = _12191_ | _12193_ /*25523*/;
assign _11973_ = _12185_ ^ _12192_ /*25526*/;
assign _12199_ = D[39] ^ Q[33] /*25522*/;
assign _12196_ = _11588_ & _12199_ /*25518*/;
assign _12197_ = _11588_ ^ _12199_ /*25521*/;
assign _12198_ = _12190_ & _12197_ /*25519*/;
assign _12195_ = _12196_ | _12198_ /*25517*/;
assign _11974_ = _12190_ ^ _12197_ /*25520*/;
assign _12204_ = D[40] ^ Q[33] /*25516*/;
assign _12201_ = _11589_ & _12204_ /*25512*/;
assign _12202_ = _11589_ ^ _12204_ /*25515*/;
assign _12203_ = _12195_ & _12202_ /*25513*/;
assign _12200_ = _12201_ | _12203_ /*25511*/;
assign _11975_ = _12195_ ^ _12202_ /*25514*/;
assign _12209_ = D[41] ^ Q[33] /*25510*/;
assign _12206_ = _11590_ & _12209_ /*25506*/;
assign _12207_ = _11590_ ^ _12209_ /*25509*/;
assign _12208_ = _12200_ & _12207_ /*25507*/;
assign _12205_ = _12206_ | _12208_ /*25505*/;
assign _11976_ = _12200_ ^ _12207_ /*25508*/;
assign _12214_ = D[42] ^ Q[33] /*25504*/;
assign _12211_ = _11591_ & _12214_ /*25500*/;
assign _12212_ = _11591_ ^ _12214_ /*25503*/;
assign _12213_ = _12205_ & _12212_ /*25501*/;
assign _12210_ = _12211_ | _12213_ /*25499*/;
assign _11977_ = _12205_ ^ _12212_ /*25502*/;
assign _12219_ = D[43] ^ Q[33] /*25498*/;
assign _12216_ = _11592_ & _12219_ /*25494*/;
assign _12217_ = _11592_ ^ _12219_ /*25497*/;
assign _12218_ = _12210_ & _12217_ /*25495*/;
assign _12215_ = _12216_ | _12218_ /*25493*/;
assign _11978_ = _12210_ ^ _12217_ /*25496*/;
assign _12224_ = D[44] ^ Q[33] /*25492*/;
assign _12221_ = _11593_ & _12224_ /*25488*/;
assign _12222_ = _11593_ ^ _12224_ /*25491*/;
assign _12223_ = _12215_ & _12222_ /*25489*/;
assign _12220_ = _12221_ | _12223_ /*25487*/;
assign _11979_ = _12215_ ^ _12222_ /*25490*/;
assign _12229_ = D[45] ^ Q[33] /*25486*/;
assign _12226_ = _11594_ & _12229_ /*25482*/;
assign _12227_ = _11594_ ^ _12229_ /*25485*/;
assign _12228_ = _12220_ & _12227_ /*25483*/;
assign _12225_ = _12226_ | _12228_ /*25481*/;
assign _11980_ = _12220_ ^ _12227_ /*25484*/;
assign _12234_ = D[46] ^ Q[33] /*25480*/;
assign _12231_ = _11595_ & _12234_ /*25476*/;
assign _12232_ = _11595_ ^ _12234_ /*25479*/;
assign _12233_ = _12225_ & _12232_ /*25477*/;
assign _12230_ = _12231_ | _12233_ /*25475*/;
assign _11981_ = _12225_ ^ _12232_ /*25478*/;
assign _12239_ = D[47] ^ Q[33] /*25474*/;
assign _12236_ = _11596_ & _12239_ /*25470*/;
assign _12237_ = _11596_ ^ _12239_ /*25473*/;
assign _12238_ = _12230_ & _12237_ /*25471*/;
assign _12235_ = _12236_ | _12238_ /*25469*/;
assign _11982_ = _12230_ ^ _12237_ /*25472*/;
assign _12244_ = D[48] ^ Q[33] /*25468*/;
assign _12241_ = _11597_ & _12244_ /*25464*/;
assign _12242_ = _11597_ ^ _12244_ /*25467*/;
assign _12243_ = _12235_ & _12242_ /*25465*/;
assign _12240_ = _12241_ | _12243_ /*25463*/;
assign _11983_ = _12235_ ^ _12242_ /*25466*/;
assign _12249_ = D[49] ^ Q[33] /*25462*/;
assign _12246_ = _11598_ & _12249_ /*25458*/;
assign _12247_ = _11598_ ^ _12249_ /*25461*/;
assign _12248_ = _12240_ & _12247_ /*25459*/;
assign _12245_ = _12246_ | _12248_ /*25457*/;
assign _11984_ = _12240_ ^ _12247_ /*25460*/;
assign _12254_ = D[50] ^ Q[33] /*25456*/;
assign _12251_ = _11599_ & _12254_ /*25452*/;
assign _12252_ = _11599_ ^ _12254_ /*25455*/;
assign _12253_ = _12245_ & _12252_ /*25453*/;
assign _12250_ = _12251_ | _12253_ /*25451*/;
assign _11985_ = _12245_ ^ _12252_ /*25454*/;
assign _12259_ = D[51] ^ Q[33] /*25450*/;
assign _12256_ = _11600_ & _12259_ /*25446*/;
assign _12257_ = _11600_ ^ _12259_ /*25449*/;
assign _12258_ = _12250_ & _12257_ /*25447*/;
assign _12255_ = _12256_ | _12258_ /*25445*/;
assign _11986_ = _12250_ ^ _12257_ /*25448*/;
assign _12264_ = D[52] ^ Q[33] /*25444*/;
assign _12261_ = _11601_ & _12264_ /*25440*/;
assign _12262_ = _11601_ ^ _12264_ /*25443*/;
assign _12263_ = _12255_ & _12262_ /*25441*/;
assign _12260_ = _12261_ | _12263_ /*25439*/;
assign _11987_ = _12255_ ^ _12262_ /*25442*/;
assign _12269_ = D[53] ^ Q[33] /*25438*/;
assign _12266_ = _11602_ & _12269_ /*25434*/;
assign _12267_ = _11602_ ^ _12269_ /*25437*/;
assign _12268_ = _12260_ & _12267_ /*25435*/;
assign _12265_ = _12266_ | _12268_ /*25433*/;
assign _11988_ = _12260_ ^ _12267_ /*25436*/;
assign _12274_ = D[54] ^ Q[33] /*25432*/;
assign _12271_ = _11603_ & _12274_ /*25428*/;
assign _12272_ = _11603_ ^ _12274_ /*25431*/;
assign _12273_ = _12265_ & _12272_ /*25429*/;
assign _12270_ = _12271_ | _12273_ /*25427*/;
assign _11989_ = _12265_ ^ _12272_ /*25430*/;
assign _12279_ = D[55] ^ Q[33] /*25426*/;
assign _12276_ = _11604_ & _12279_ /*25422*/;
assign _12277_ = _11604_ ^ _12279_ /*25425*/;
assign _12278_ = _12270_ & _12277_ /*25423*/;
assign _12275_ = _12276_ | _12278_ /*25421*/;
assign _11990_ = _12270_ ^ _12277_ /*25424*/;
assign _12284_ = D[56] ^ Q[33] /*25420*/;
assign _12281_ = _11605_ & _12284_ /*25416*/;
assign _12282_ = _11605_ ^ _12284_ /*25419*/;
assign _12283_ = _12275_ & _12282_ /*25417*/;
assign _12280_ = _12281_ | _12283_ /*25415*/;
assign _11991_ = _12275_ ^ _12282_ /*25418*/;
assign _12289_ = D[57] ^ Q[33] /*25414*/;
assign _12286_ = _11606_ & _12289_ /*25410*/;
assign _12287_ = _11606_ ^ _12289_ /*25413*/;
assign _12288_ = _12280_ & _12287_ /*25411*/;
assign _12285_ = _12286_ | _12288_ /*25409*/;
assign _11992_ = _12280_ ^ _12287_ /*25412*/;
assign _12294_ = D[58] ^ Q[33] /*25408*/;
assign _12291_ = _11607_ & _12294_ /*25404*/;
assign _12292_ = _11607_ ^ _12294_ /*25407*/;
assign _12293_ = _12285_ & _12292_ /*25405*/;
assign _12290_ = _12291_ | _12293_ /*25403*/;
assign _11993_ = _12285_ ^ _12292_ /*25406*/;
assign _12299_ = D[59] ^ Q[33] /*25402*/;
assign _12296_ = _11608_ & _12299_ /*25398*/;
assign _12297_ = _11608_ ^ _12299_ /*25401*/;
assign _12298_ = _12290_ & _12297_ /*25399*/;
assign _12295_ = _12296_ | _12298_ /*25397*/;
assign _11994_ = _12290_ ^ _12297_ /*25400*/;
assign _12304_ = D[60] ^ Q[33] /*25396*/;
assign _12301_ = _11609_ & _12304_ /*25392*/;
assign _12302_ = _11609_ ^ _12304_ /*25395*/;
assign _12303_ = _12295_ & _12302_ /*25393*/;
assign _12300_ = _12301_ | _12303_ /*25391*/;
assign _11995_ = _12295_ ^ _12302_ /*25394*/;
assign _12309_ = D[61] ^ Q[33] /*25390*/;
assign _12306_ = _11610_ & _12309_ /*25386*/;
assign _12307_ = _11610_ ^ _12309_ /*25389*/;
assign _12308_ = _12300_ & _12307_ /*25387*/;
assign _12305_ = _12306_ | _12308_ /*25385*/;
assign _11996_ = _12300_ ^ _12307_ /*25388*/;
assign _12314_ = D[62] ^ Q[33] /*25384*/;
assign _12311_ = _11611_ & _12314_ /*25380*/;
assign _12312_ = _11611_ ^ _12314_ /*25383*/;
assign _12313_ = _12305_ & _12312_ /*25381*/;
assign _12310_ = _12311_ | _12313_ /*25379*/;
assign _11997_ = _12305_ ^ _12312_ /*25382*/;
assign _12318_ = zeroWire ^ Q[33] /*25378*/;
assign _12315_ = _11612_ & _12318_ /*25374*/;
assign _12316_ = _11612_ ^ _12318_ /*25377*/;
assign _12317_ = _12310_ & _12316_ /*25375*/;
assign Q[32] = _12315_ | _12317_ /*25373*/;
assign _11998_ = _12310_ ^ _12316_ /*25376*/;
assign _12389_ = D[0] ^ Q[32] /*24987*/;
assign _12386_ = R_0[31] & _12389_ /*24983*/;
assign _12387_ = R_0[31] ^ _12389_ /*24986*/;
assign _12388_ = Q[32] & _12387_ /*24984*/;
assign _12385_ = _12386_ | _12388_ /*24982*/;
assign _12320_ = Q[32] ^ _12387_ /*24985*/;
assign _12394_ = D[1] ^ Q[32] /*24981*/;
assign _12391_ = _11935_ & _12394_ /*24977*/;
assign _12392_ = _11935_ ^ _12394_ /*24980*/;
assign _12393_ = _12385_ & _12392_ /*24978*/;
assign _12390_ = _12391_ | _12393_ /*24976*/;
assign _12321_ = _12385_ ^ _12392_ /*24979*/;
assign _12399_ = D[2] ^ Q[32] /*24975*/;
assign _12396_ = _11936_ & _12399_ /*24971*/;
assign _12397_ = _11936_ ^ _12399_ /*24974*/;
assign _12398_ = _12390_ & _12397_ /*24972*/;
assign _12395_ = _12396_ | _12398_ /*24970*/;
assign _12322_ = _12390_ ^ _12397_ /*24973*/;
assign _12404_ = D[3] ^ Q[32] /*24969*/;
assign _12401_ = _11937_ & _12404_ /*24965*/;
assign _12402_ = _11937_ ^ _12404_ /*24968*/;
assign _12403_ = _12395_ & _12402_ /*24966*/;
assign _12400_ = _12401_ | _12403_ /*24964*/;
assign _12323_ = _12395_ ^ _12402_ /*24967*/;
assign _12409_ = D[4] ^ Q[32] /*24963*/;
assign _12406_ = _11938_ & _12409_ /*24959*/;
assign _12407_ = _11938_ ^ _12409_ /*24962*/;
assign _12408_ = _12400_ & _12407_ /*24960*/;
assign _12405_ = _12406_ | _12408_ /*24958*/;
assign _12324_ = _12400_ ^ _12407_ /*24961*/;
assign _12414_ = D[5] ^ Q[32] /*24957*/;
assign _12411_ = _11939_ & _12414_ /*24953*/;
assign _12412_ = _11939_ ^ _12414_ /*24956*/;
assign _12413_ = _12405_ & _12412_ /*24954*/;
assign _12410_ = _12411_ | _12413_ /*24952*/;
assign _12325_ = _12405_ ^ _12412_ /*24955*/;
assign _12419_ = D[6] ^ Q[32] /*24951*/;
assign _12416_ = _11940_ & _12419_ /*24947*/;
assign _12417_ = _11940_ ^ _12419_ /*24950*/;
assign _12418_ = _12410_ & _12417_ /*24948*/;
assign _12415_ = _12416_ | _12418_ /*24946*/;
assign _12326_ = _12410_ ^ _12417_ /*24949*/;
assign _12424_ = D[7] ^ Q[32] /*24945*/;
assign _12421_ = _11941_ & _12424_ /*24941*/;
assign _12422_ = _11941_ ^ _12424_ /*24944*/;
assign _12423_ = _12415_ & _12422_ /*24942*/;
assign _12420_ = _12421_ | _12423_ /*24940*/;
assign _12327_ = _12415_ ^ _12422_ /*24943*/;
assign _12429_ = D[8] ^ Q[32] /*24939*/;
assign _12426_ = _11942_ & _12429_ /*24935*/;
assign _12427_ = _11942_ ^ _12429_ /*24938*/;
assign _12428_ = _12420_ & _12427_ /*24936*/;
assign _12425_ = _12426_ | _12428_ /*24934*/;
assign _12328_ = _12420_ ^ _12427_ /*24937*/;
assign _12434_ = D[9] ^ Q[32] /*24933*/;
assign _12431_ = _11943_ & _12434_ /*24929*/;
assign _12432_ = _11943_ ^ _12434_ /*24932*/;
assign _12433_ = _12425_ & _12432_ /*24930*/;
assign _12430_ = _12431_ | _12433_ /*24928*/;
assign _12329_ = _12425_ ^ _12432_ /*24931*/;
assign _12439_ = D[10] ^ Q[32] /*24927*/;
assign _12436_ = _11944_ & _12439_ /*24923*/;
assign _12437_ = _11944_ ^ _12439_ /*24926*/;
assign _12438_ = _12430_ & _12437_ /*24924*/;
assign _12435_ = _12436_ | _12438_ /*24922*/;
assign _12330_ = _12430_ ^ _12437_ /*24925*/;
assign _12444_ = D[11] ^ Q[32] /*24921*/;
assign _12441_ = _11945_ & _12444_ /*24917*/;
assign _12442_ = _11945_ ^ _12444_ /*24920*/;
assign _12443_ = _12435_ & _12442_ /*24918*/;
assign _12440_ = _12441_ | _12443_ /*24916*/;
assign _12331_ = _12435_ ^ _12442_ /*24919*/;
assign _12449_ = D[12] ^ Q[32] /*24915*/;
assign _12446_ = _11946_ & _12449_ /*24911*/;
assign _12447_ = _11946_ ^ _12449_ /*24914*/;
assign _12448_ = _12440_ & _12447_ /*24912*/;
assign _12445_ = _12446_ | _12448_ /*24910*/;
assign _12332_ = _12440_ ^ _12447_ /*24913*/;
assign _12454_ = D[13] ^ Q[32] /*24909*/;
assign _12451_ = _11947_ & _12454_ /*24905*/;
assign _12452_ = _11947_ ^ _12454_ /*24908*/;
assign _12453_ = _12445_ & _12452_ /*24906*/;
assign _12450_ = _12451_ | _12453_ /*24904*/;
assign _12333_ = _12445_ ^ _12452_ /*24907*/;
assign _12459_ = D[14] ^ Q[32] /*24903*/;
assign _12456_ = _11948_ & _12459_ /*24899*/;
assign _12457_ = _11948_ ^ _12459_ /*24902*/;
assign _12458_ = _12450_ & _12457_ /*24900*/;
assign _12455_ = _12456_ | _12458_ /*24898*/;
assign _12334_ = _12450_ ^ _12457_ /*24901*/;
assign _12464_ = D[15] ^ Q[32] /*24897*/;
assign _12461_ = _11949_ & _12464_ /*24893*/;
assign _12462_ = _11949_ ^ _12464_ /*24896*/;
assign _12463_ = _12455_ & _12462_ /*24894*/;
assign _12460_ = _12461_ | _12463_ /*24892*/;
assign _12335_ = _12455_ ^ _12462_ /*24895*/;
assign _12469_ = D[16] ^ Q[32] /*24891*/;
assign _12466_ = _11950_ & _12469_ /*24887*/;
assign _12467_ = _11950_ ^ _12469_ /*24890*/;
assign _12468_ = _12460_ & _12467_ /*24888*/;
assign _12465_ = _12466_ | _12468_ /*24886*/;
assign _12336_ = _12460_ ^ _12467_ /*24889*/;
assign _12474_ = D[17] ^ Q[32] /*24885*/;
assign _12471_ = _11951_ & _12474_ /*24881*/;
assign _12472_ = _11951_ ^ _12474_ /*24884*/;
assign _12473_ = _12465_ & _12472_ /*24882*/;
assign _12470_ = _12471_ | _12473_ /*24880*/;
assign _12337_ = _12465_ ^ _12472_ /*24883*/;
assign _12479_ = D[18] ^ Q[32] /*24879*/;
assign _12476_ = _11952_ & _12479_ /*24875*/;
assign _12477_ = _11952_ ^ _12479_ /*24878*/;
assign _12478_ = _12470_ & _12477_ /*24876*/;
assign _12475_ = _12476_ | _12478_ /*24874*/;
assign _12338_ = _12470_ ^ _12477_ /*24877*/;
assign _12484_ = D[19] ^ Q[32] /*24873*/;
assign _12481_ = _11953_ & _12484_ /*24869*/;
assign _12482_ = _11953_ ^ _12484_ /*24872*/;
assign _12483_ = _12475_ & _12482_ /*24870*/;
assign _12480_ = _12481_ | _12483_ /*24868*/;
assign _12339_ = _12475_ ^ _12482_ /*24871*/;
assign _12489_ = D[20] ^ Q[32] /*24867*/;
assign _12486_ = _11954_ & _12489_ /*24863*/;
assign _12487_ = _11954_ ^ _12489_ /*24866*/;
assign _12488_ = _12480_ & _12487_ /*24864*/;
assign _12485_ = _12486_ | _12488_ /*24862*/;
assign _12340_ = _12480_ ^ _12487_ /*24865*/;
assign _12494_ = D[21] ^ Q[32] /*24861*/;
assign _12491_ = _11955_ & _12494_ /*24857*/;
assign _12492_ = _11955_ ^ _12494_ /*24860*/;
assign _12493_ = _12485_ & _12492_ /*24858*/;
assign _12490_ = _12491_ | _12493_ /*24856*/;
assign _12341_ = _12485_ ^ _12492_ /*24859*/;
assign _12499_ = D[22] ^ Q[32] /*24855*/;
assign _12496_ = _11956_ & _12499_ /*24851*/;
assign _12497_ = _11956_ ^ _12499_ /*24854*/;
assign _12498_ = _12490_ & _12497_ /*24852*/;
assign _12495_ = _12496_ | _12498_ /*24850*/;
assign _12342_ = _12490_ ^ _12497_ /*24853*/;
assign _12504_ = D[23] ^ Q[32] /*24849*/;
assign _12501_ = _11957_ & _12504_ /*24845*/;
assign _12502_ = _11957_ ^ _12504_ /*24848*/;
assign _12503_ = _12495_ & _12502_ /*24846*/;
assign _12500_ = _12501_ | _12503_ /*24844*/;
assign _12343_ = _12495_ ^ _12502_ /*24847*/;
assign _12509_ = D[24] ^ Q[32] /*24843*/;
assign _12506_ = _11958_ & _12509_ /*24839*/;
assign _12507_ = _11958_ ^ _12509_ /*24842*/;
assign _12508_ = _12500_ & _12507_ /*24840*/;
assign _12505_ = _12506_ | _12508_ /*24838*/;
assign _12344_ = _12500_ ^ _12507_ /*24841*/;
assign _12514_ = D[25] ^ Q[32] /*24837*/;
assign _12511_ = _11959_ & _12514_ /*24833*/;
assign _12512_ = _11959_ ^ _12514_ /*24836*/;
assign _12513_ = _12505_ & _12512_ /*24834*/;
assign _12510_ = _12511_ | _12513_ /*24832*/;
assign _12345_ = _12505_ ^ _12512_ /*24835*/;
assign _12519_ = D[26] ^ Q[32] /*24831*/;
assign _12516_ = _11960_ & _12519_ /*24827*/;
assign _12517_ = _11960_ ^ _12519_ /*24830*/;
assign _12518_ = _12510_ & _12517_ /*24828*/;
assign _12515_ = _12516_ | _12518_ /*24826*/;
assign _12346_ = _12510_ ^ _12517_ /*24829*/;
assign _12524_ = D[27] ^ Q[32] /*24825*/;
assign _12521_ = _11961_ & _12524_ /*24821*/;
assign _12522_ = _11961_ ^ _12524_ /*24824*/;
assign _12523_ = _12515_ & _12522_ /*24822*/;
assign _12520_ = _12521_ | _12523_ /*24820*/;
assign _12347_ = _12515_ ^ _12522_ /*24823*/;
assign _12529_ = D[28] ^ Q[32] /*24819*/;
assign _12526_ = _11962_ & _12529_ /*24815*/;
assign _12527_ = _11962_ ^ _12529_ /*24818*/;
assign _12528_ = _12520_ & _12527_ /*24816*/;
assign _12525_ = _12526_ | _12528_ /*24814*/;
assign _12348_ = _12520_ ^ _12527_ /*24817*/;
assign _12534_ = D[29] ^ Q[32] /*24813*/;
assign _12531_ = _11963_ & _12534_ /*24809*/;
assign _12532_ = _11963_ ^ _12534_ /*24812*/;
assign _12533_ = _12525_ & _12532_ /*24810*/;
assign _12530_ = _12531_ | _12533_ /*24808*/;
assign _12349_ = _12525_ ^ _12532_ /*24811*/;
assign _12539_ = D[30] ^ Q[32] /*24807*/;
assign _12536_ = _11964_ & _12539_ /*24803*/;
assign _12537_ = _11964_ ^ _12539_ /*24806*/;
assign _12538_ = _12530_ & _12537_ /*24804*/;
assign _12535_ = _12536_ | _12538_ /*24802*/;
assign _12350_ = _12530_ ^ _12537_ /*24805*/;
assign _12544_ = D[31] ^ Q[32] /*24801*/;
assign _12541_ = _11965_ & _12544_ /*24797*/;
assign _12542_ = _11965_ ^ _12544_ /*24800*/;
assign _12543_ = _12535_ & _12542_ /*24798*/;
assign _12540_ = _12541_ | _12543_ /*24796*/;
assign _12351_ = _12535_ ^ _12542_ /*24799*/;
assign _12549_ = D[32] ^ Q[32] /*24795*/;
assign _12546_ = _11966_ & _12549_ /*24791*/;
assign _12547_ = _11966_ ^ _12549_ /*24794*/;
assign _12548_ = _12540_ & _12547_ /*24792*/;
assign _12545_ = _12546_ | _12548_ /*24790*/;
assign _12352_ = _12540_ ^ _12547_ /*24793*/;
assign _12554_ = D[33] ^ Q[32] /*24789*/;
assign _12551_ = _11967_ & _12554_ /*24785*/;
assign _12552_ = _11967_ ^ _12554_ /*24788*/;
assign _12553_ = _12545_ & _12552_ /*24786*/;
assign _12550_ = _12551_ | _12553_ /*24784*/;
assign _12353_ = _12545_ ^ _12552_ /*24787*/;
assign _12559_ = D[34] ^ Q[32] /*24783*/;
assign _12556_ = _11968_ & _12559_ /*24779*/;
assign _12557_ = _11968_ ^ _12559_ /*24782*/;
assign _12558_ = _12550_ & _12557_ /*24780*/;
assign _12555_ = _12556_ | _12558_ /*24778*/;
assign _12354_ = _12550_ ^ _12557_ /*24781*/;
assign _12564_ = D[35] ^ Q[32] /*24777*/;
assign _12561_ = _11969_ & _12564_ /*24773*/;
assign _12562_ = _11969_ ^ _12564_ /*24776*/;
assign _12563_ = _12555_ & _12562_ /*24774*/;
assign _12560_ = _12561_ | _12563_ /*24772*/;
assign _12355_ = _12555_ ^ _12562_ /*24775*/;
assign _12569_ = D[36] ^ Q[32] /*24771*/;
assign _12566_ = _11970_ & _12569_ /*24767*/;
assign _12567_ = _11970_ ^ _12569_ /*24770*/;
assign _12568_ = _12560_ & _12567_ /*24768*/;
assign _12565_ = _12566_ | _12568_ /*24766*/;
assign _12356_ = _12560_ ^ _12567_ /*24769*/;
assign _12574_ = D[37] ^ Q[32] /*24765*/;
assign _12571_ = _11971_ & _12574_ /*24761*/;
assign _12572_ = _11971_ ^ _12574_ /*24764*/;
assign _12573_ = _12565_ & _12572_ /*24762*/;
assign _12570_ = _12571_ | _12573_ /*24760*/;
assign _12357_ = _12565_ ^ _12572_ /*24763*/;
assign _12579_ = D[38] ^ Q[32] /*24759*/;
assign _12576_ = _11972_ & _12579_ /*24755*/;
assign _12577_ = _11972_ ^ _12579_ /*24758*/;
assign _12578_ = _12570_ & _12577_ /*24756*/;
assign _12575_ = _12576_ | _12578_ /*24754*/;
assign _12358_ = _12570_ ^ _12577_ /*24757*/;
assign _12584_ = D[39] ^ Q[32] /*24753*/;
assign _12581_ = _11973_ & _12584_ /*24749*/;
assign _12582_ = _11973_ ^ _12584_ /*24752*/;
assign _12583_ = _12575_ & _12582_ /*24750*/;
assign _12580_ = _12581_ | _12583_ /*24748*/;
assign _12359_ = _12575_ ^ _12582_ /*24751*/;
assign _12589_ = D[40] ^ Q[32] /*24747*/;
assign _12586_ = _11974_ & _12589_ /*24743*/;
assign _12587_ = _11974_ ^ _12589_ /*24746*/;
assign _12588_ = _12580_ & _12587_ /*24744*/;
assign _12585_ = _12586_ | _12588_ /*24742*/;
assign _12360_ = _12580_ ^ _12587_ /*24745*/;
assign _12594_ = D[41] ^ Q[32] /*24741*/;
assign _12591_ = _11975_ & _12594_ /*24737*/;
assign _12592_ = _11975_ ^ _12594_ /*24740*/;
assign _12593_ = _12585_ & _12592_ /*24738*/;
assign _12590_ = _12591_ | _12593_ /*24736*/;
assign _12361_ = _12585_ ^ _12592_ /*24739*/;
assign _12599_ = D[42] ^ Q[32] /*24735*/;
assign _12596_ = _11976_ & _12599_ /*24731*/;
assign _12597_ = _11976_ ^ _12599_ /*24734*/;
assign _12598_ = _12590_ & _12597_ /*24732*/;
assign _12595_ = _12596_ | _12598_ /*24730*/;
assign _12362_ = _12590_ ^ _12597_ /*24733*/;
assign _12604_ = D[43] ^ Q[32] /*24729*/;
assign _12601_ = _11977_ & _12604_ /*24725*/;
assign _12602_ = _11977_ ^ _12604_ /*24728*/;
assign _12603_ = _12595_ & _12602_ /*24726*/;
assign _12600_ = _12601_ | _12603_ /*24724*/;
assign _12363_ = _12595_ ^ _12602_ /*24727*/;
assign _12609_ = D[44] ^ Q[32] /*24723*/;
assign _12606_ = _11978_ & _12609_ /*24719*/;
assign _12607_ = _11978_ ^ _12609_ /*24722*/;
assign _12608_ = _12600_ & _12607_ /*24720*/;
assign _12605_ = _12606_ | _12608_ /*24718*/;
assign _12364_ = _12600_ ^ _12607_ /*24721*/;
assign _12614_ = D[45] ^ Q[32] /*24717*/;
assign _12611_ = _11979_ & _12614_ /*24713*/;
assign _12612_ = _11979_ ^ _12614_ /*24716*/;
assign _12613_ = _12605_ & _12612_ /*24714*/;
assign _12610_ = _12611_ | _12613_ /*24712*/;
assign _12365_ = _12605_ ^ _12612_ /*24715*/;
assign _12619_ = D[46] ^ Q[32] /*24711*/;
assign _12616_ = _11980_ & _12619_ /*24707*/;
assign _12617_ = _11980_ ^ _12619_ /*24710*/;
assign _12618_ = _12610_ & _12617_ /*24708*/;
assign _12615_ = _12616_ | _12618_ /*24706*/;
assign _12366_ = _12610_ ^ _12617_ /*24709*/;
assign _12624_ = D[47] ^ Q[32] /*24705*/;
assign _12621_ = _11981_ & _12624_ /*24701*/;
assign _12622_ = _11981_ ^ _12624_ /*24704*/;
assign _12623_ = _12615_ & _12622_ /*24702*/;
assign _12620_ = _12621_ | _12623_ /*24700*/;
assign _12367_ = _12615_ ^ _12622_ /*24703*/;
assign _12629_ = D[48] ^ Q[32] /*24699*/;
assign _12626_ = _11982_ & _12629_ /*24695*/;
assign _12627_ = _11982_ ^ _12629_ /*24698*/;
assign _12628_ = _12620_ & _12627_ /*24696*/;
assign _12625_ = _12626_ | _12628_ /*24694*/;
assign _12368_ = _12620_ ^ _12627_ /*24697*/;
assign _12634_ = D[49] ^ Q[32] /*24693*/;
assign _12631_ = _11983_ & _12634_ /*24689*/;
assign _12632_ = _11983_ ^ _12634_ /*24692*/;
assign _12633_ = _12625_ & _12632_ /*24690*/;
assign _12630_ = _12631_ | _12633_ /*24688*/;
assign _12369_ = _12625_ ^ _12632_ /*24691*/;
assign _12639_ = D[50] ^ Q[32] /*24687*/;
assign _12636_ = _11984_ & _12639_ /*24683*/;
assign _12637_ = _11984_ ^ _12639_ /*24686*/;
assign _12638_ = _12630_ & _12637_ /*24684*/;
assign _12635_ = _12636_ | _12638_ /*24682*/;
assign _12370_ = _12630_ ^ _12637_ /*24685*/;
assign _12644_ = D[51] ^ Q[32] /*24681*/;
assign _12641_ = _11985_ & _12644_ /*24677*/;
assign _12642_ = _11985_ ^ _12644_ /*24680*/;
assign _12643_ = _12635_ & _12642_ /*24678*/;
assign _12640_ = _12641_ | _12643_ /*24676*/;
assign _12371_ = _12635_ ^ _12642_ /*24679*/;
assign _12649_ = D[52] ^ Q[32] /*24675*/;
assign _12646_ = _11986_ & _12649_ /*24671*/;
assign _12647_ = _11986_ ^ _12649_ /*24674*/;
assign _12648_ = _12640_ & _12647_ /*24672*/;
assign _12645_ = _12646_ | _12648_ /*24670*/;
assign _12372_ = _12640_ ^ _12647_ /*24673*/;
assign _12654_ = D[53] ^ Q[32] /*24669*/;
assign _12651_ = _11987_ & _12654_ /*24665*/;
assign _12652_ = _11987_ ^ _12654_ /*24668*/;
assign _12653_ = _12645_ & _12652_ /*24666*/;
assign _12650_ = _12651_ | _12653_ /*24664*/;
assign _12373_ = _12645_ ^ _12652_ /*24667*/;
assign _12659_ = D[54] ^ Q[32] /*24663*/;
assign _12656_ = _11988_ & _12659_ /*24659*/;
assign _12657_ = _11988_ ^ _12659_ /*24662*/;
assign _12658_ = _12650_ & _12657_ /*24660*/;
assign _12655_ = _12656_ | _12658_ /*24658*/;
assign _12374_ = _12650_ ^ _12657_ /*24661*/;
assign _12664_ = D[55] ^ Q[32] /*24657*/;
assign _12661_ = _11989_ & _12664_ /*24653*/;
assign _12662_ = _11989_ ^ _12664_ /*24656*/;
assign _12663_ = _12655_ & _12662_ /*24654*/;
assign _12660_ = _12661_ | _12663_ /*24652*/;
assign _12375_ = _12655_ ^ _12662_ /*24655*/;
assign _12669_ = D[56] ^ Q[32] /*24651*/;
assign _12666_ = _11990_ & _12669_ /*24647*/;
assign _12667_ = _11990_ ^ _12669_ /*24650*/;
assign _12668_ = _12660_ & _12667_ /*24648*/;
assign _12665_ = _12666_ | _12668_ /*24646*/;
assign _12376_ = _12660_ ^ _12667_ /*24649*/;
assign _12674_ = D[57] ^ Q[32] /*24645*/;
assign _12671_ = _11991_ & _12674_ /*24641*/;
assign _12672_ = _11991_ ^ _12674_ /*24644*/;
assign _12673_ = _12665_ & _12672_ /*24642*/;
assign _12670_ = _12671_ | _12673_ /*24640*/;
assign _12377_ = _12665_ ^ _12672_ /*24643*/;
assign _12679_ = D[58] ^ Q[32] /*24639*/;
assign _12676_ = _11992_ & _12679_ /*24635*/;
assign _12677_ = _11992_ ^ _12679_ /*24638*/;
assign _12678_ = _12670_ & _12677_ /*24636*/;
assign _12675_ = _12676_ | _12678_ /*24634*/;
assign _12378_ = _12670_ ^ _12677_ /*24637*/;
assign _12684_ = D[59] ^ Q[32] /*24633*/;
assign _12681_ = _11993_ & _12684_ /*24629*/;
assign _12682_ = _11993_ ^ _12684_ /*24632*/;
assign _12683_ = _12675_ & _12682_ /*24630*/;
assign _12680_ = _12681_ | _12683_ /*24628*/;
assign _12379_ = _12675_ ^ _12682_ /*24631*/;
assign _12689_ = D[60] ^ Q[32] /*24627*/;
assign _12686_ = _11994_ & _12689_ /*24623*/;
assign _12687_ = _11994_ ^ _12689_ /*24626*/;
assign _12688_ = _12680_ & _12687_ /*24624*/;
assign _12685_ = _12686_ | _12688_ /*24622*/;
assign _12380_ = _12680_ ^ _12687_ /*24625*/;
assign _12694_ = D[61] ^ Q[32] /*24621*/;
assign _12691_ = _11995_ & _12694_ /*24617*/;
assign _12692_ = _11995_ ^ _12694_ /*24620*/;
assign _12693_ = _12685_ & _12692_ /*24618*/;
assign _12690_ = _12691_ | _12693_ /*24616*/;
assign _12381_ = _12685_ ^ _12692_ /*24619*/;
assign _12699_ = D[62] ^ Q[32] /*24615*/;
assign _12696_ = _11996_ & _12699_ /*24611*/;
assign _12697_ = _11996_ ^ _12699_ /*24614*/;
assign _12698_ = _12690_ & _12697_ /*24612*/;
assign _12695_ = _12696_ | _12698_ /*24610*/;
assign _12382_ = _12690_ ^ _12697_ /*24613*/;
assign _12703_ = zeroWire ^ Q[32] /*24609*/;
assign _12700_ = _11997_ & _12703_ /*24605*/;
assign _12701_ = _11997_ ^ _12703_ /*24608*/;
assign _12702_ = _12695_ & _12701_ /*24606*/;
assign Q[31] = _12700_ | _12702_ /*24604*/;
assign _12383_ = _12695_ ^ _12701_ /*24607*/;
assign _12774_ = D[0] ^ Q[31] /*24218*/;
assign _12771_ = R_0[30] & _12774_ /*24214*/;
assign _12772_ = R_0[30] ^ _12774_ /*24217*/;
assign _12773_ = Q[31] & _12772_ /*24215*/;
assign _12770_ = _12771_ | _12773_ /*24213*/;
assign _12705_ = Q[31] ^ _12772_ /*24216*/;
assign _12779_ = D[1] ^ Q[31] /*24212*/;
assign _12776_ = _12320_ & _12779_ /*24208*/;
assign _12777_ = _12320_ ^ _12779_ /*24211*/;
assign _12778_ = _12770_ & _12777_ /*24209*/;
assign _12775_ = _12776_ | _12778_ /*24207*/;
assign _12706_ = _12770_ ^ _12777_ /*24210*/;
assign _12784_ = D[2] ^ Q[31] /*24206*/;
assign _12781_ = _12321_ & _12784_ /*24202*/;
assign _12782_ = _12321_ ^ _12784_ /*24205*/;
assign _12783_ = _12775_ & _12782_ /*24203*/;
assign _12780_ = _12781_ | _12783_ /*24201*/;
assign _12707_ = _12775_ ^ _12782_ /*24204*/;
assign _12789_ = D[3] ^ Q[31] /*24200*/;
assign _12786_ = _12322_ & _12789_ /*24196*/;
assign _12787_ = _12322_ ^ _12789_ /*24199*/;
assign _12788_ = _12780_ & _12787_ /*24197*/;
assign _12785_ = _12786_ | _12788_ /*24195*/;
assign _12708_ = _12780_ ^ _12787_ /*24198*/;
assign _12794_ = D[4] ^ Q[31] /*24194*/;
assign _12791_ = _12323_ & _12794_ /*24190*/;
assign _12792_ = _12323_ ^ _12794_ /*24193*/;
assign _12793_ = _12785_ & _12792_ /*24191*/;
assign _12790_ = _12791_ | _12793_ /*24189*/;
assign _12709_ = _12785_ ^ _12792_ /*24192*/;
assign _12799_ = D[5] ^ Q[31] /*24188*/;
assign _12796_ = _12324_ & _12799_ /*24184*/;
assign _12797_ = _12324_ ^ _12799_ /*24187*/;
assign _12798_ = _12790_ & _12797_ /*24185*/;
assign _12795_ = _12796_ | _12798_ /*24183*/;
assign _12710_ = _12790_ ^ _12797_ /*24186*/;
assign _12804_ = D[6] ^ Q[31] /*24182*/;
assign _12801_ = _12325_ & _12804_ /*24178*/;
assign _12802_ = _12325_ ^ _12804_ /*24181*/;
assign _12803_ = _12795_ & _12802_ /*24179*/;
assign _12800_ = _12801_ | _12803_ /*24177*/;
assign _12711_ = _12795_ ^ _12802_ /*24180*/;
assign _12809_ = D[7] ^ Q[31] /*24176*/;
assign _12806_ = _12326_ & _12809_ /*24172*/;
assign _12807_ = _12326_ ^ _12809_ /*24175*/;
assign _12808_ = _12800_ & _12807_ /*24173*/;
assign _12805_ = _12806_ | _12808_ /*24171*/;
assign _12712_ = _12800_ ^ _12807_ /*24174*/;
assign _12814_ = D[8] ^ Q[31] /*24170*/;
assign _12811_ = _12327_ & _12814_ /*24166*/;
assign _12812_ = _12327_ ^ _12814_ /*24169*/;
assign _12813_ = _12805_ & _12812_ /*24167*/;
assign _12810_ = _12811_ | _12813_ /*24165*/;
assign _12713_ = _12805_ ^ _12812_ /*24168*/;
assign _12819_ = D[9] ^ Q[31] /*24164*/;
assign _12816_ = _12328_ & _12819_ /*24160*/;
assign _12817_ = _12328_ ^ _12819_ /*24163*/;
assign _12818_ = _12810_ & _12817_ /*24161*/;
assign _12815_ = _12816_ | _12818_ /*24159*/;
assign _12714_ = _12810_ ^ _12817_ /*24162*/;
assign _12824_ = D[10] ^ Q[31] /*24158*/;
assign _12821_ = _12329_ & _12824_ /*24154*/;
assign _12822_ = _12329_ ^ _12824_ /*24157*/;
assign _12823_ = _12815_ & _12822_ /*24155*/;
assign _12820_ = _12821_ | _12823_ /*24153*/;
assign _12715_ = _12815_ ^ _12822_ /*24156*/;
assign _12829_ = D[11] ^ Q[31] /*24152*/;
assign _12826_ = _12330_ & _12829_ /*24148*/;
assign _12827_ = _12330_ ^ _12829_ /*24151*/;
assign _12828_ = _12820_ & _12827_ /*24149*/;
assign _12825_ = _12826_ | _12828_ /*24147*/;
assign _12716_ = _12820_ ^ _12827_ /*24150*/;
assign _12834_ = D[12] ^ Q[31] /*24146*/;
assign _12831_ = _12331_ & _12834_ /*24142*/;
assign _12832_ = _12331_ ^ _12834_ /*24145*/;
assign _12833_ = _12825_ & _12832_ /*24143*/;
assign _12830_ = _12831_ | _12833_ /*24141*/;
assign _12717_ = _12825_ ^ _12832_ /*24144*/;
assign _12839_ = D[13] ^ Q[31] /*24140*/;
assign _12836_ = _12332_ & _12839_ /*24136*/;
assign _12837_ = _12332_ ^ _12839_ /*24139*/;
assign _12838_ = _12830_ & _12837_ /*24137*/;
assign _12835_ = _12836_ | _12838_ /*24135*/;
assign _12718_ = _12830_ ^ _12837_ /*24138*/;
assign _12844_ = D[14] ^ Q[31] /*24134*/;
assign _12841_ = _12333_ & _12844_ /*24130*/;
assign _12842_ = _12333_ ^ _12844_ /*24133*/;
assign _12843_ = _12835_ & _12842_ /*24131*/;
assign _12840_ = _12841_ | _12843_ /*24129*/;
assign _12719_ = _12835_ ^ _12842_ /*24132*/;
assign _12849_ = D[15] ^ Q[31] /*24128*/;
assign _12846_ = _12334_ & _12849_ /*24124*/;
assign _12847_ = _12334_ ^ _12849_ /*24127*/;
assign _12848_ = _12840_ & _12847_ /*24125*/;
assign _12845_ = _12846_ | _12848_ /*24123*/;
assign _12720_ = _12840_ ^ _12847_ /*24126*/;
assign _12854_ = D[16] ^ Q[31] /*24122*/;
assign _12851_ = _12335_ & _12854_ /*24118*/;
assign _12852_ = _12335_ ^ _12854_ /*24121*/;
assign _12853_ = _12845_ & _12852_ /*24119*/;
assign _12850_ = _12851_ | _12853_ /*24117*/;
assign _12721_ = _12845_ ^ _12852_ /*24120*/;
assign _12859_ = D[17] ^ Q[31] /*24116*/;
assign _12856_ = _12336_ & _12859_ /*24112*/;
assign _12857_ = _12336_ ^ _12859_ /*24115*/;
assign _12858_ = _12850_ & _12857_ /*24113*/;
assign _12855_ = _12856_ | _12858_ /*24111*/;
assign _12722_ = _12850_ ^ _12857_ /*24114*/;
assign _12864_ = D[18] ^ Q[31] /*24110*/;
assign _12861_ = _12337_ & _12864_ /*24106*/;
assign _12862_ = _12337_ ^ _12864_ /*24109*/;
assign _12863_ = _12855_ & _12862_ /*24107*/;
assign _12860_ = _12861_ | _12863_ /*24105*/;
assign _12723_ = _12855_ ^ _12862_ /*24108*/;
assign _12869_ = D[19] ^ Q[31] /*24104*/;
assign _12866_ = _12338_ & _12869_ /*24100*/;
assign _12867_ = _12338_ ^ _12869_ /*24103*/;
assign _12868_ = _12860_ & _12867_ /*24101*/;
assign _12865_ = _12866_ | _12868_ /*24099*/;
assign _12724_ = _12860_ ^ _12867_ /*24102*/;
assign _12874_ = D[20] ^ Q[31] /*24098*/;
assign _12871_ = _12339_ & _12874_ /*24094*/;
assign _12872_ = _12339_ ^ _12874_ /*24097*/;
assign _12873_ = _12865_ & _12872_ /*24095*/;
assign _12870_ = _12871_ | _12873_ /*24093*/;
assign _12725_ = _12865_ ^ _12872_ /*24096*/;
assign _12879_ = D[21] ^ Q[31] /*24092*/;
assign _12876_ = _12340_ & _12879_ /*24088*/;
assign _12877_ = _12340_ ^ _12879_ /*24091*/;
assign _12878_ = _12870_ & _12877_ /*24089*/;
assign _12875_ = _12876_ | _12878_ /*24087*/;
assign _12726_ = _12870_ ^ _12877_ /*24090*/;
assign _12884_ = D[22] ^ Q[31] /*24086*/;
assign _12881_ = _12341_ & _12884_ /*24082*/;
assign _12882_ = _12341_ ^ _12884_ /*24085*/;
assign _12883_ = _12875_ & _12882_ /*24083*/;
assign _12880_ = _12881_ | _12883_ /*24081*/;
assign _12727_ = _12875_ ^ _12882_ /*24084*/;
assign _12889_ = D[23] ^ Q[31] /*24080*/;
assign _12886_ = _12342_ & _12889_ /*24076*/;
assign _12887_ = _12342_ ^ _12889_ /*24079*/;
assign _12888_ = _12880_ & _12887_ /*24077*/;
assign _12885_ = _12886_ | _12888_ /*24075*/;
assign _12728_ = _12880_ ^ _12887_ /*24078*/;
assign _12894_ = D[24] ^ Q[31] /*24074*/;
assign _12891_ = _12343_ & _12894_ /*24070*/;
assign _12892_ = _12343_ ^ _12894_ /*24073*/;
assign _12893_ = _12885_ & _12892_ /*24071*/;
assign _12890_ = _12891_ | _12893_ /*24069*/;
assign _12729_ = _12885_ ^ _12892_ /*24072*/;
assign _12899_ = D[25] ^ Q[31] /*24068*/;
assign _12896_ = _12344_ & _12899_ /*24064*/;
assign _12897_ = _12344_ ^ _12899_ /*24067*/;
assign _12898_ = _12890_ & _12897_ /*24065*/;
assign _12895_ = _12896_ | _12898_ /*24063*/;
assign _12730_ = _12890_ ^ _12897_ /*24066*/;
assign _12904_ = D[26] ^ Q[31] /*24062*/;
assign _12901_ = _12345_ & _12904_ /*24058*/;
assign _12902_ = _12345_ ^ _12904_ /*24061*/;
assign _12903_ = _12895_ & _12902_ /*24059*/;
assign _12900_ = _12901_ | _12903_ /*24057*/;
assign _12731_ = _12895_ ^ _12902_ /*24060*/;
assign _12909_ = D[27] ^ Q[31] /*24056*/;
assign _12906_ = _12346_ & _12909_ /*24052*/;
assign _12907_ = _12346_ ^ _12909_ /*24055*/;
assign _12908_ = _12900_ & _12907_ /*24053*/;
assign _12905_ = _12906_ | _12908_ /*24051*/;
assign _12732_ = _12900_ ^ _12907_ /*24054*/;
assign _12914_ = D[28] ^ Q[31] /*24050*/;
assign _12911_ = _12347_ & _12914_ /*24046*/;
assign _12912_ = _12347_ ^ _12914_ /*24049*/;
assign _12913_ = _12905_ & _12912_ /*24047*/;
assign _12910_ = _12911_ | _12913_ /*24045*/;
assign _12733_ = _12905_ ^ _12912_ /*24048*/;
assign _12919_ = D[29] ^ Q[31] /*24044*/;
assign _12916_ = _12348_ & _12919_ /*24040*/;
assign _12917_ = _12348_ ^ _12919_ /*24043*/;
assign _12918_ = _12910_ & _12917_ /*24041*/;
assign _12915_ = _12916_ | _12918_ /*24039*/;
assign _12734_ = _12910_ ^ _12917_ /*24042*/;
assign _12924_ = D[30] ^ Q[31] /*24038*/;
assign _12921_ = _12349_ & _12924_ /*24034*/;
assign _12922_ = _12349_ ^ _12924_ /*24037*/;
assign _12923_ = _12915_ & _12922_ /*24035*/;
assign _12920_ = _12921_ | _12923_ /*24033*/;
assign _12735_ = _12915_ ^ _12922_ /*24036*/;
assign _12929_ = D[31] ^ Q[31] /*24032*/;
assign _12926_ = _12350_ & _12929_ /*24028*/;
assign _12927_ = _12350_ ^ _12929_ /*24031*/;
assign _12928_ = _12920_ & _12927_ /*24029*/;
assign _12925_ = _12926_ | _12928_ /*24027*/;
assign _12736_ = _12920_ ^ _12927_ /*24030*/;
assign _12934_ = D[32] ^ Q[31] /*24026*/;
assign _12931_ = _12351_ & _12934_ /*24022*/;
assign _12932_ = _12351_ ^ _12934_ /*24025*/;
assign _12933_ = _12925_ & _12932_ /*24023*/;
assign _12930_ = _12931_ | _12933_ /*24021*/;
assign _12737_ = _12925_ ^ _12932_ /*24024*/;
assign _12939_ = D[33] ^ Q[31] /*24020*/;
assign _12936_ = _12352_ & _12939_ /*24016*/;
assign _12937_ = _12352_ ^ _12939_ /*24019*/;
assign _12938_ = _12930_ & _12937_ /*24017*/;
assign _12935_ = _12936_ | _12938_ /*24015*/;
assign _12738_ = _12930_ ^ _12937_ /*24018*/;
assign _12944_ = D[34] ^ Q[31] /*24014*/;
assign _12941_ = _12353_ & _12944_ /*24010*/;
assign _12942_ = _12353_ ^ _12944_ /*24013*/;
assign _12943_ = _12935_ & _12942_ /*24011*/;
assign _12940_ = _12941_ | _12943_ /*24009*/;
assign _12739_ = _12935_ ^ _12942_ /*24012*/;
assign _12949_ = D[35] ^ Q[31] /*24008*/;
assign _12946_ = _12354_ & _12949_ /*24004*/;
assign _12947_ = _12354_ ^ _12949_ /*24007*/;
assign _12948_ = _12940_ & _12947_ /*24005*/;
assign _12945_ = _12946_ | _12948_ /*24003*/;
assign _12740_ = _12940_ ^ _12947_ /*24006*/;
assign _12954_ = D[36] ^ Q[31] /*24002*/;
assign _12951_ = _12355_ & _12954_ /*23998*/;
assign _12952_ = _12355_ ^ _12954_ /*24001*/;
assign _12953_ = _12945_ & _12952_ /*23999*/;
assign _12950_ = _12951_ | _12953_ /*23997*/;
assign _12741_ = _12945_ ^ _12952_ /*24000*/;
assign _12959_ = D[37] ^ Q[31] /*23996*/;
assign _12956_ = _12356_ & _12959_ /*23992*/;
assign _12957_ = _12356_ ^ _12959_ /*23995*/;
assign _12958_ = _12950_ & _12957_ /*23993*/;
assign _12955_ = _12956_ | _12958_ /*23991*/;
assign _12742_ = _12950_ ^ _12957_ /*23994*/;
assign _12964_ = D[38] ^ Q[31] /*23990*/;
assign _12961_ = _12357_ & _12964_ /*23986*/;
assign _12962_ = _12357_ ^ _12964_ /*23989*/;
assign _12963_ = _12955_ & _12962_ /*23987*/;
assign _12960_ = _12961_ | _12963_ /*23985*/;
assign _12743_ = _12955_ ^ _12962_ /*23988*/;
assign _12969_ = D[39] ^ Q[31] /*23984*/;
assign _12966_ = _12358_ & _12969_ /*23980*/;
assign _12967_ = _12358_ ^ _12969_ /*23983*/;
assign _12968_ = _12960_ & _12967_ /*23981*/;
assign _12965_ = _12966_ | _12968_ /*23979*/;
assign _12744_ = _12960_ ^ _12967_ /*23982*/;
assign _12974_ = D[40] ^ Q[31] /*23978*/;
assign _12971_ = _12359_ & _12974_ /*23974*/;
assign _12972_ = _12359_ ^ _12974_ /*23977*/;
assign _12973_ = _12965_ & _12972_ /*23975*/;
assign _12970_ = _12971_ | _12973_ /*23973*/;
assign _12745_ = _12965_ ^ _12972_ /*23976*/;
assign _12979_ = D[41] ^ Q[31] /*23972*/;
assign _12976_ = _12360_ & _12979_ /*23968*/;
assign _12977_ = _12360_ ^ _12979_ /*23971*/;
assign _12978_ = _12970_ & _12977_ /*23969*/;
assign _12975_ = _12976_ | _12978_ /*23967*/;
assign _12746_ = _12970_ ^ _12977_ /*23970*/;
assign _12984_ = D[42] ^ Q[31] /*23966*/;
assign _12981_ = _12361_ & _12984_ /*23962*/;
assign _12982_ = _12361_ ^ _12984_ /*23965*/;
assign _12983_ = _12975_ & _12982_ /*23963*/;
assign _12980_ = _12981_ | _12983_ /*23961*/;
assign _12747_ = _12975_ ^ _12982_ /*23964*/;
assign _12989_ = D[43] ^ Q[31] /*23960*/;
assign _12986_ = _12362_ & _12989_ /*23956*/;
assign _12987_ = _12362_ ^ _12989_ /*23959*/;
assign _12988_ = _12980_ & _12987_ /*23957*/;
assign _12985_ = _12986_ | _12988_ /*23955*/;
assign _12748_ = _12980_ ^ _12987_ /*23958*/;
assign _12994_ = D[44] ^ Q[31] /*23954*/;
assign _12991_ = _12363_ & _12994_ /*23950*/;
assign _12992_ = _12363_ ^ _12994_ /*23953*/;
assign _12993_ = _12985_ & _12992_ /*23951*/;
assign _12990_ = _12991_ | _12993_ /*23949*/;
assign _12749_ = _12985_ ^ _12992_ /*23952*/;
assign _12999_ = D[45] ^ Q[31] /*23948*/;
assign _12996_ = _12364_ & _12999_ /*23944*/;
assign _12997_ = _12364_ ^ _12999_ /*23947*/;
assign _12998_ = _12990_ & _12997_ /*23945*/;
assign _12995_ = _12996_ | _12998_ /*23943*/;
assign _12750_ = _12990_ ^ _12997_ /*23946*/;
assign _13004_ = D[46] ^ Q[31] /*23942*/;
assign _13001_ = _12365_ & _13004_ /*23938*/;
assign _13002_ = _12365_ ^ _13004_ /*23941*/;
assign _13003_ = _12995_ & _13002_ /*23939*/;
assign _13000_ = _13001_ | _13003_ /*23937*/;
assign _12751_ = _12995_ ^ _13002_ /*23940*/;
assign _13009_ = D[47] ^ Q[31] /*23936*/;
assign _13006_ = _12366_ & _13009_ /*23932*/;
assign _13007_ = _12366_ ^ _13009_ /*23935*/;
assign _13008_ = _13000_ & _13007_ /*23933*/;
assign _13005_ = _13006_ | _13008_ /*23931*/;
assign _12752_ = _13000_ ^ _13007_ /*23934*/;
assign _13014_ = D[48] ^ Q[31] /*23930*/;
assign _13011_ = _12367_ & _13014_ /*23926*/;
assign _13012_ = _12367_ ^ _13014_ /*23929*/;
assign _13013_ = _13005_ & _13012_ /*23927*/;
assign _13010_ = _13011_ | _13013_ /*23925*/;
assign _12753_ = _13005_ ^ _13012_ /*23928*/;
assign _13019_ = D[49] ^ Q[31] /*23924*/;
assign _13016_ = _12368_ & _13019_ /*23920*/;
assign _13017_ = _12368_ ^ _13019_ /*23923*/;
assign _13018_ = _13010_ & _13017_ /*23921*/;
assign _13015_ = _13016_ | _13018_ /*23919*/;
assign _12754_ = _13010_ ^ _13017_ /*23922*/;
assign _13024_ = D[50] ^ Q[31] /*23918*/;
assign _13021_ = _12369_ & _13024_ /*23914*/;
assign _13022_ = _12369_ ^ _13024_ /*23917*/;
assign _13023_ = _13015_ & _13022_ /*23915*/;
assign _13020_ = _13021_ | _13023_ /*23913*/;
assign _12755_ = _13015_ ^ _13022_ /*23916*/;
assign _13029_ = D[51] ^ Q[31] /*23912*/;
assign _13026_ = _12370_ & _13029_ /*23908*/;
assign _13027_ = _12370_ ^ _13029_ /*23911*/;
assign _13028_ = _13020_ & _13027_ /*23909*/;
assign _13025_ = _13026_ | _13028_ /*23907*/;
assign _12756_ = _13020_ ^ _13027_ /*23910*/;
assign _13034_ = D[52] ^ Q[31] /*23906*/;
assign _13031_ = _12371_ & _13034_ /*23902*/;
assign _13032_ = _12371_ ^ _13034_ /*23905*/;
assign _13033_ = _13025_ & _13032_ /*23903*/;
assign _13030_ = _13031_ | _13033_ /*23901*/;
assign _12757_ = _13025_ ^ _13032_ /*23904*/;
assign _13039_ = D[53] ^ Q[31] /*23900*/;
assign _13036_ = _12372_ & _13039_ /*23896*/;
assign _13037_ = _12372_ ^ _13039_ /*23899*/;
assign _13038_ = _13030_ & _13037_ /*23897*/;
assign _13035_ = _13036_ | _13038_ /*23895*/;
assign _12758_ = _13030_ ^ _13037_ /*23898*/;
assign _13044_ = D[54] ^ Q[31] /*23894*/;
assign _13041_ = _12373_ & _13044_ /*23890*/;
assign _13042_ = _12373_ ^ _13044_ /*23893*/;
assign _13043_ = _13035_ & _13042_ /*23891*/;
assign _13040_ = _13041_ | _13043_ /*23889*/;
assign _12759_ = _13035_ ^ _13042_ /*23892*/;
assign _13049_ = D[55] ^ Q[31] /*23888*/;
assign _13046_ = _12374_ & _13049_ /*23884*/;
assign _13047_ = _12374_ ^ _13049_ /*23887*/;
assign _13048_ = _13040_ & _13047_ /*23885*/;
assign _13045_ = _13046_ | _13048_ /*23883*/;
assign _12760_ = _13040_ ^ _13047_ /*23886*/;
assign _13054_ = D[56] ^ Q[31] /*23882*/;
assign _13051_ = _12375_ & _13054_ /*23878*/;
assign _13052_ = _12375_ ^ _13054_ /*23881*/;
assign _13053_ = _13045_ & _13052_ /*23879*/;
assign _13050_ = _13051_ | _13053_ /*23877*/;
assign _12761_ = _13045_ ^ _13052_ /*23880*/;
assign _13059_ = D[57] ^ Q[31] /*23876*/;
assign _13056_ = _12376_ & _13059_ /*23872*/;
assign _13057_ = _12376_ ^ _13059_ /*23875*/;
assign _13058_ = _13050_ & _13057_ /*23873*/;
assign _13055_ = _13056_ | _13058_ /*23871*/;
assign _12762_ = _13050_ ^ _13057_ /*23874*/;
assign _13064_ = D[58] ^ Q[31] /*23870*/;
assign _13061_ = _12377_ & _13064_ /*23866*/;
assign _13062_ = _12377_ ^ _13064_ /*23869*/;
assign _13063_ = _13055_ & _13062_ /*23867*/;
assign _13060_ = _13061_ | _13063_ /*23865*/;
assign _12763_ = _13055_ ^ _13062_ /*23868*/;
assign _13069_ = D[59] ^ Q[31] /*23864*/;
assign _13066_ = _12378_ & _13069_ /*23860*/;
assign _13067_ = _12378_ ^ _13069_ /*23863*/;
assign _13068_ = _13060_ & _13067_ /*23861*/;
assign _13065_ = _13066_ | _13068_ /*23859*/;
assign _12764_ = _13060_ ^ _13067_ /*23862*/;
assign _13074_ = D[60] ^ Q[31] /*23858*/;
assign _13071_ = _12379_ & _13074_ /*23854*/;
assign _13072_ = _12379_ ^ _13074_ /*23857*/;
assign _13073_ = _13065_ & _13072_ /*23855*/;
assign _13070_ = _13071_ | _13073_ /*23853*/;
assign _12765_ = _13065_ ^ _13072_ /*23856*/;
assign _13079_ = D[61] ^ Q[31] /*23852*/;
assign _13076_ = _12380_ & _13079_ /*23848*/;
assign _13077_ = _12380_ ^ _13079_ /*23851*/;
assign _13078_ = _13070_ & _13077_ /*23849*/;
assign _13075_ = _13076_ | _13078_ /*23847*/;
assign _12766_ = _13070_ ^ _13077_ /*23850*/;
assign _13084_ = D[62] ^ Q[31] /*23846*/;
assign _13081_ = _12381_ & _13084_ /*23842*/;
assign _13082_ = _12381_ ^ _13084_ /*23845*/;
assign _13083_ = _13075_ & _13082_ /*23843*/;
assign _13080_ = _13081_ | _13083_ /*23841*/;
assign _12767_ = _13075_ ^ _13082_ /*23844*/;
assign _13088_ = zeroWire ^ Q[31] /*23840*/;
assign _13085_ = _12382_ & _13088_ /*23836*/;
assign _13086_ = _12382_ ^ _13088_ /*23839*/;
assign _13087_ = _13080_ & _13086_ /*23837*/;
assign Q[30] = _13085_ | _13087_ /*23835*/;
assign _12768_ = _13080_ ^ _13086_ /*23838*/;
assign _13159_ = D[0] ^ Q[30] /*23449*/;
assign _13156_ = R_0[29] & _13159_ /*23445*/;
assign _13157_ = R_0[29] ^ _13159_ /*23448*/;
assign _13158_ = Q[30] & _13157_ /*23446*/;
assign _13155_ = _13156_ | _13158_ /*23444*/;
assign _13090_ = Q[30] ^ _13157_ /*23447*/;
assign _13164_ = D[1] ^ Q[30] /*23443*/;
assign _13161_ = _12705_ & _13164_ /*23439*/;
assign _13162_ = _12705_ ^ _13164_ /*23442*/;
assign _13163_ = _13155_ & _13162_ /*23440*/;
assign _13160_ = _13161_ | _13163_ /*23438*/;
assign _13091_ = _13155_ ^ _13162_ /*23441*/;
assign _13169_ = D[2] ^ Q[30] /*23437*/;
assign _13166_ = _12706_ & _13169_ /*23433*/;
assign _13167_ = _12706_ ^ _13169_ /*23436*/;
assign _13168_ = _13160_ & _13167_ /*23434*/;
assign _13165_ = _13166_ | _13168_ /*23432*/;
assign _13092_ = _13160_ ^ _13167_ /*23435*/;
assign _13174_ = D[3] ^ Q[30] /*23431*/;
assign _13171_ = _12707_ & _13174_ /*23427*/;
assign _13172_ = _12707_ ^ _13174_ /*23430*/;
assign _13173_ = _13165_ & _13172_ /*23428*/;
assign _13170_ = _13171_ | _13173_ /*23426*/;
assign _13093_ = _13165_ ^ _13172_ /*23429*/;
assign _13179_ = D[4] ^ Q[30] /*23425*/;
assign _13176_ = _12708_ & _13179_ /*23421*/;
assign _13177_ = _12708_ ^ _13179_ /*23424*/;
assign _13178_ = _13170_ & _13177_ /*23422*/;
assign _13175_ = _13176_ | _13178_ /*23420*/;
assign _13094_ = _13170_ ^ _13177_ /*23423*/;
assign _13184_ = D[5] ^ Q[30] /*23419*/;
assign _13181_ = _12709_ & _13184_ /*23415*/;
assign _13182_ = _12709_ ^ _13184_ /*23418*/;
assign _13183_ = _13175_ & _13182_ /*23416*/;
assign _13180_ = _13181_ | _13183_ /*23414*/;
assign _13095_ = _13175_ ^ _13182_ /*23417*/;
assign _13189_ = D[6] ^ Q[30] /*23413*/;
assign _13186_ = _12710_ & _13189_ /*23409*/;
assign _13187_ = _12710_ ^ _13189_ /*23412*/;
assign _13188_ = _13180_ & _13187_ /*23410*/;
assign _13185_ = _13186_ | _13188_ /*23408*/;
assign _13096_ = _13180_ ^ _13187_ /*23411*/;
assign _13194_ = D[7] ^ Q[30] /*23407*/;
assign _13191_ = _12711_ & _13194_ /*23403*/;
assign _13192_ = _12711_ ^ _13194_ /*23406*/;
assign _13193_ = _13185_ & _13192_ /*23404*/;
assign _13190_ = _13191_ | _13193_ /*23402*/;
assign _13097_ = _13185_ ^ _13192_ /*23405*/;
assign _13199_ = D[8] ^ Q[30] /*23401*/;
assign _13196_ = _12712_ & _13199_ /*23397*/;
assign _13197_ = _12712_ ^ _13199_ /*23400*/;
assign _13198_ = _13190_ & _13197_ /*23398*/;
assign _13195_ = _13196_ | _13198_ /*23396*/;
assign _13098_ = _13190_ ^ _13197_ /*23399*/;
assign _13204_ = D[9] ^ Q[30] /*23395*/;
assign _13201_ = _12713_ & _13204_ /*23391*/;
assign _13202_ = _12713_ ^ _13204_ /*23394*/;
assign _13203_ = _13195_ & _13202_ /*23392*/;
assign _13200_ = _13201_ | _13203_ /*23390*/;
assign _13099_ = _13195_ ^ _13202_ /*23393*/;
assign _13209_ = D[10] ^ Q[30] /*23389*/;
assign _13206_ = _12714_ & _13209_ /*23385*/;
assign _13207_ = _12714_ ^ _13209_ /*23388*/;
assign _13208_ = _13200_ & _13207_ /*23386*/;
assign _13205_ = _13206_ | _13208_ /*23384*/;
assign _13100_ = _13200_ ^ _13207_ /*23387*/;
assign _13214_ = D[11] ^ Q[30] /*23383*/;
assign _13211_ = _12715_ & _13214_ /*23379*/;
assign _13212_ = _12715_ ^ _13214_ /*23382*/;
assign _13213_ = _13205_ & _13212_ /*23380*/;
assign _13210_ = _13211_ | _13213_ /*23378*/;
assign _13101_ = _13205_ ^ _13212_ /*23381*/;
assign _13219_ = D[12] ^ Q[30] /*23377*/;
assign _13216_ = _12716_ & _13219_ /*23373*/;
assign _13217_ = _12716_ ^ _13219_ /*23376*/;
assign _13218_ = _13210_ & _13217_ /*23374*/;
assign _13215_ = _13216_ | _13218_ /*23372*/;
assign _13102_ = _13210_ ^ _13217_ /*23375*/;
assign _13224_ = D[13] ^ Q[30] /*23371*/;
assign _13221_ = _12717_ & _13224_ /*23367*/;
assign _13222_ = _12717_ ^ _13224_ /*23370*/;
assign _13223_ = _13215_ & _13222_ /*23368*/;
assign _13220_ = _13221_ | _13223_ /*23366*/;
assign _13103_ = _13215_ ^ _13222_ /*23369*/;
assign _13229_ = D[14] ^ Q[30] /*23365*/;
assign _13226_ = _12718_ & _13229_ /*23361*/;
assign _13227_ = _12718_ ^ _13229_ /*23364*/;
assign _13228_ = _13220_ & _13227_ /*23362*/;
assign _13225_ = _13226_ | _13228_ /*23360*/;
assign _13104_ = _13220_ ^ _13227_ /*23363*/;
assign _13234_ = D[15] ^ Q[30] /*23359*/;
assign _13231_ = _12719_ & _13234_ /*23355*/;
assign _13232_ = _12719_ ^ _13234_ /*23358*/;
assign _13233_ = _13225_ & _13232_ /*23356*/;
assign _13230_ = _13231_ | _13233_ /*23354*/;
assign _13105_ = _13225_ ^ _13232_ /*23357*/;
assign _13239_ = D[16] ^ Q[30] /*23353*/;
assign _13236_ = _12720_ & _13239_ /*23349*/;
assign _13237_ = _12720_ ^ _13239_ /*23352*/;
assign _13238_ = _13230_ & _13237_ /*23350*/;
assign _13235_ = _13236_ | _13238_ /*23348*/;
assign _13106_ = _13230_ ^ _13237_ /*23351*/;
assign _13244_ = D[17] ^ Q[30] /*23347*/;
assign _13241_ = _12721_ & _13244_ /*23343*/;
assign _13242_ = _12721_ ^ _13244_ /*23346*/;
assign _13243_ = _13235_ & _13242_ /*23344*/;
assign _13240_ = _13241_ | _13243_ /*23342*/;
assign _13107_ = _13235_ ^ _13242_ /*23345*/;
assign _13249_ = D[18] ^ Q[30] /*23341*/;
assign _13246_ = _12722_ & _13249_ /*23337*/;
assign _13247_ = _12722_ ^ _13249_ /*23340*/;
assign _13248_ = _13240_ & _13247_ /*23338*/;
assign _13245_ = _13246_ | _13248_ /*23336*/;
assign _13108_ = _13240_ ^ _13247_ /*23339*/;
assign _13254_ = D[19] ^ Q[30] /*23335*/;
assign _13251_ = _12723_ & _13254_ /*23331*/;
assign _13252_ = _12723_ ^ _13254_ /*23334*/;
assign _13253_ = _13245_ & _13252_ /*23332*/;
assign _13250_ = _13251_ | _13253_ /*23330*/;
assign _13109_ = _13245_ ^ _13252_ /*23333*/;
assign _13259_ = D[20] ^ Q[30] /*23329*/;
assign _13256_ = _12724_ & _13259_ /*23325*/;
assign _13257_ = _12724_ ^ _13259_ /*23328*/;
assign _13258_ = _13250_ & _13257_ /*23326*/;
assign _13255_ = _13256_ | _13258_ /*23324*/;
assign _13110_ = _13250_ ^ _13257_ /*23327*/;
assign _13264_ = D[21] ^ Q[30] /*23323*/;
assign _13261_ = _12725_ & _13264_ /*23319*/;
assign _13262_ = _12725_ ^ _13264_ /*23322*/;
assign _13263_ = _13255_ & _13262_ /*23320*/;
assign _13260_ = _13261_ | _13263_ /*23318*/;
assign _13111_ = _13255_ ^ _13262_ /*23321*/;
assign _13269_ = D[22] ^ Q[30] /*23317*/;
assign _13266_ = _12726_ & _13269_ /*23313*/;
assign _13267_ = _12726_ ^ _13269_ /*23316*/;
assign _13268_ = _13260_ & _13267_ /*23314*/;
assign _13265_ = _13266_ | _13268_ /*23312*/;
assign _13112_ = _13260_ ^ _13267_ /*23315*/;
assign _13274_ = D[23] ^ Q[30] /*23311*/;
assign _13271_ = _12727_ & _13274_ /*23307*/;
assign _13272_ = _12727_ ^ _13274_ /*23310*/;
assign _13273_ = _13265_ & _13272_ /*23308*/;
assign _13270_ = _13271_ | _13273_ /*23306*/;
assign _13113_ = _13265_ ^ _13272_ /*23309*/;
assign _13279_ = D[24] ^ Q[30] /*23305*/;
assign _13276_ = _12728_ & _13279_ /*23301*/;
assign _13277_ = _12728_ ^ _13279_ /*23304*/;
assign _13278_ = _13270_ & _13277_ /*23302*/;
assign _13275_ = _13276_ | _13278_ /*23300*/;
assign _13114_ = _13270_ ^ _13277_ /*23303*/;
assign _13284_ = D[25] ^ Q[30] /*23299*/;
assign _13281_ = _12729_ & _13284_ /*23295*/;
assign _13282_ = _12729_ ^ _13284_ /*23298*/;
assign _13283_ = _13275_ & _13282_ /*23296*/;
assign _13280_ = _13281_ | _13283_ /*23294*/;
assign _13115_ = _13275_ ^ _13282_ /*23297*/;
assign _13289_ = D[26] ^ Q[30] /*23293*/;
assign _13286_ = _12730_ & _13289_ /*23289*/;
assign _13287_ = _12730_ ^ _13289_ /*23292*/;
assign _13288_ = _13280_ & _13287_ /*23290*/;
assign _13285_ = _13286_ | _13288_ /*23288*/;
assign _13116_ = _13280_ ^ _13287_ /*23291*/;
assign _13294_ = D[27] ^ Q[30] /*23287*/;
assign _13291_ = _12731_ & _13294_ /*23283*/;
assign _13292_ = _12731_ ^ _13294_ /*23286*/;
assign _13293_ = _13285_ & _13292_ /*23284*/;
assign _13290_ = _13291_ | _13293_ /*23282*/;
assign _13117_ = _13285_ ^ _13292_ /*23285*/;
assign _13299_ = D[28] ^ Q[30] /*23281*/;
assign _13296_ = _12732_ & _13299_ /*23277*/;
assign _13297_ = _12732_ ^ _13299_ /*23280*/;
assign _13298_ = _13290_ & _13297_ /*23278*/;
assign _13295_ = _13296_ | _13298_ /*23276*/;
assign _13118_ = _13290_ ^ _13297_ /*23279*/;
assign _13304_ = D[29] ^ Q[30] /*23275*/;
assign _13301_ = _12733_ & _13304_ /*23271*/;
assign _13302_ = _12733_ ^ _13304_ /*23274*/;
assign _13303_ = _13295_ & _13302_ /*23272*/;
assign _13300_ = _13301_ | _13303_ /*23270*/;
assign _13119_ = _13295_ ^ _13302_ /*23273*/;
assign _13309_ = D[30] ^ Q[30] /*23269*/;
assign _13306_ = _12734_ & _13309_ /*23265*/;
assign _13307_ = _12734_ ^ _13309_ /*23268*/;
assign _13308_ = _13300_ & _13307_ /*23266*/;
assign _13305_ = _13306_ | _13308_ /*23264*/;
assign _13120_ = _13300_ ^ _13307_ /*23267*/;
assign _13314_ = D[31] ^ Q[30] /*23263*/;
assign _13311_ = _12735_ & _13314_ /*23259*/;
assign _13312_ = _12735_ ^ _13314_ /*23262*/;
assign _13313_ = _13305_ & _13312_ /*23260*/;
assign _13310_ = _13311_ | _13313_ /*23258*/;
assign _13121_ = _13305_ ^ _13312_ /*23261*/;
assign _13319_ = D[32] ^ Q[30] /*23257*/;
assign _13316_ = _12736_ & _13319_ /*23253*/;
assign _13317_ = _12736_ ^ _13319_ /*23256*/;
assign _13318_ = _13310_ & _13317_ /*23254*/;
assign _13315_ = _13316_ | _13318_ /*23252*/;
assign _13122_ = _13310_ ^ _13317_ /*23255*/;
assign _13324_ = D[33] ^ Q[30] /*23251*/;
assign _13321_ = _12737_ & _13324_ /*23247*/;
assign _13322_ = _12737_ ^ _13324_ /*23250*/;
assign _13323_ = _13315_ & _13322_ /*23248*/;
assign _13320_ = _13321_ | _13323_ /*23246*/;
assign _13123_ = _13315_ ^ _13322_ /*23249*/;
assign _13329_ = D[34] ^ Q[30] /*23245*/;
assign _13326_ = _12738_ & _13329_ /*23241*/;
assign _13327_ = _12738_ ^ _13329_ /*23244*/;
assign _13328_ = _13320_ & _13327_ /*23242*/;
assign _13325_ = _13326_ | _13328_ /*23240*/;
assign _13124_ = _13320_ ^ _13327_ /*23243*/;
assign _13334_ = D[35] ^ Q[30] /*23239*/;
assign _13331_ = _12739_ & _13334_ /*23235*/;
assign _13332_ = _12739_ ^ _13334_ /*23238*/;
assign _13333_ = _13325_ & _13332_ /*23236*/;
assign _13330_ = _13331_ | _13333_ /*23234*/;
assign _13125_ = _13325_ ^ _13332_ /*23237*/;
assign _13339_ = D[36] ^ Q[30] /*23233*/;
assign _13336_ = _12740_ & _13339_ /*23229*/;
assign _13337_ = _12740_ ^ _13339_ /*23232*/;
assign _13338_ = _13330_ & _13337_ /*23230*/;
assign _13335_ = _13336_ | _13338_ /*23228*/;
assign _13126_ = _13330_ ^ _13337_ /*23231*/;
assign _13344_ = D[37] ^ Q[30] /*23227*/;
assign _13341_ = _12741_ & _13344_ /*23223*/;
assign _13342_ = _12741_ ^ _13344_ /*23226*/;
assign _13343_ = _13335_ & _13342_ /*23224*/;
assign _13340_ = _13341_ | _13343_ /*23222*/;
assign _13127_ = _13335_ ^ _13342_ /*23225*/;
assign _13349_ = D[38] ^ Q[30] /*23221*/;
assign _13346_ = _12742_ & _13349_ /*23217*/;
assign _13347_ = _12742_ ^ _13349_ /*23220*/;
assign _13348_ = _13340_ & _13347_ /*23218*/;
assign _13345_ = _13346_ | _13348_ /*23216*/;
assign _13128_ = _13340_ ^ _13347_ /*23219*/;
assign _13354_ = D[39] ^ Q[30] /*23215*/;
assign _13351_ = _12743_ & _13354_ /*23211*/;
assign _13352_ = _12743_ ^ _13354_ /*23214*/;
assign _13353_ = _13345_ & _13352_ /*23212*/;
assign _13350_ = _13351_ | _13353_ /*23210*/;
assign _13129_ = _13345_ ^ _13352_ /*23213*/;
assign _13359_ = D[40] ^ Q[30] /*23209*/;
assign _13356_ = _12744_ & _13359_ /*23205*/;
assign _13357_ = _12744_ ^ _13359_ /*23208*/;
assign _13358_ = _13350_ & _13357_ /*23206*/;
assign _13355_ = _13356_ | _13358_ /*23204*/;
assign _13130_ = _13350_ ^ _13357_ /*23207*/;
assign _13364_ = D[41] ^ Q[30] /*23203*/;
assign _13361_ = _12745_ & _13364_ /*23199*/;
assign _13362_ = _12745_ ^ _13364_ /*23202*/;
assign _13363_ = _13355_ & _13362_ /*23200*/;
assign _13360_ = _13361_ | _13363_ /*23198*/;
assign _13131_ = _13355_ ^ _13362_ /*23201*/;
assign _13369_ = D[42] ^ Q[30] /*23197*/;
assign _13366_ = _12746_ & _13369_ /*23193*/;
assign _13367_ = _12746_ ^ _13369_ /*23196*/;
assign _13368_ = _13360_ & _13367_ /*23194*/;
assign _13365_ = _13366_ | _13368_ /*23192*/;
assign _13132_ = _13360_ ^ _13367_ /*23195*/;
assign _13374_ = D[43] ^ Q[30] /*23191*/;
assign _13371_ = _12747_ & _13374_ /*23187*/;
assign _13372_ = _12747_ ^ _13374_ /*23190*/;
assign _13373_ = _13365_ & _13372_ /*23188*/;
assign _13370_ = _13371_ | _13373_ /*23186*/;
assign _13133_ = _13365_ ^ _13372_ /*23189*/;
assign _13379_ = D[44] ^ Q[30] /*23185*/;
assign _13376_ = _12748_ & _13379_ /*23181*/;
assign _13377_ = _12748_ ^ _13379_ /*23184*/;
assign _13378_ = _13370_ & _13377_ /*23182*/;
assign _13375_ = _13376_ | _13378_ /*23180*/;
assign _13134_ = _13370_ ^ _13377_ /*23183*/;
assign _13384_ = D[45] ^ Q[30] /*23179*/;
assign _13381_ = _12749_ & _13384_ /*23175*/;
assign _13382_ = _12749_ ^ _13384_ /*23178*/;
assign _13383_ = _13375_ & _13382_ /*23176*/;
assign _13380_ = _13381_ | _13383_ /*23174*/;
assign _13135_ = _13375_ ^ _13382_ /*23177*/;
assign _13389_ = D[46] ^ Q[30] /*23173*/;
assign _13386_ = _12750_ & _13389_ /*23169*/;
assign _13387_ = _12750_ ^ _13389_ /*23172*/;
assign _13388_ = _13380_ & _13387_ /*23170*/;
assign _13385_ = _13386_ | _13388_ /*23168*/;
assign _13136_ = _13380_ ^ _13387_ /*23171*/;
assign _13394_ = D[47] ^ Q[30] /*23167*/;
assign _13391_ = _12751_ & _13394_ /*23163*/;
assign _13392_ = _12751_ ^ _13394_ /*23166*/;
assign _13393_ = _13385_ & _13392_ /*23164*/;
assign _13390_ = _13391_ | _13393_ /*23162*/;
assign _13137_ = _13385_ ^ _13392_ /*23165*/;
assign _13399_ = D[48] ^ Q[30] /*23161*/;
assign _13396_ = _12752_ & _13399_ /*23157*/;
assign _13397_ = _12752_ ^ _13399_ /*23160*/;
assign _13398_ = _13390_ & _13397_ /*23158*/;
assign _13395_ = _13396_ | _13398_ /*23156*/;
assign _13138_ = _13390_ ^ _13397_ /*23159*/;
assign _13404_ = D[49] ^ Q[30] /*23155*/;
assign _13401_ = _12753_ & _13404_ /*23151*/;
assign _13402_ = _12753_ ^ _13404_ /*23154*/;
assign _13403_ = _13395_ & _13402_ /*23152*/;
assign _13400_ = _13401_ | _13403_ /*23150*/;
assign _13139_ = _13395_ ^ _13402_ /*23153*/;
assign _13409_ = D[50] ^ Q[30] /*23149*/;
assign _13406_ = _12754_ & _13409_ /*23145*/;
assign _13407_ = _12754_ ^ _13409_ /*23148*/;
assign _13408_ = _13400_ & _13407_ /*23146*/;
assign _13405_ = _13406_ | _13408_ /*23144*/;
assign _13140_ = _13400_ ^ _13407_ /*23147*/;
assign _13414_ = D[51] ^ Q[30] /*23143*/;
assign _13411_ = _12755_ & _13414_ /*23139*/;
assign _13412_ = _12755_ ^ _13414_ /*23142*/;
assign _13413_ = _13405_ & _13412_ /*23140*/;
assign _13410_ = _13411_ | _13413_ /*23138*/;
assign _13141_ = _13405_ ^ _13412_ /*23141*/;
assign _13419_ = D[52] ^ Q[30] /*23137*/;
assign _13416_ = _12756_ & _13419_ /*23133*/;
assign _13417_ = _12756_ ^ _13419_ /*23136*/;
assign _13418_ = _13410_ & _13417_ /*23134*/;
assign _13415_ = _13416_ | _13418_ /*23132*/;
assign _13142_ = _13410_ ^ _13417_ /*23135*/;
assign _13424_ = D[53] ^ Q[30] /*23131*/;
assign _13421_ = _12757_ & _13424_ /*23127*/;
assign _13422_ = _12757_ ^ _13424_ /*23130*/;
assign _13423_ = _13415_ & _13422_ /*23128*/;
assign _13420_ = _13421_ | _13423_ /*23126*/;
assign _13143_ = _13415_ ^ _13422_ /*23129*/;
assign _13429_ = D[54] ^ Q[30] /*23125*/;
assign _13426_ = _12758_ & _13429_ /*23121*/;
assign _13427_ = _12758_ ^ _13429_ /*23124*/;
assign _13428_ = _13420_ & _13427_ /*23122*/;
assign _13425_ = _13426_ | _13428_ /*23120*/;
assign _13144_ = _13420_ ^ _13427_ /*23123*/;
assign _13434_ = D[55] ^ Q[30] /*23119*/;
assign _13431_ = _12759_ & _13434_ /*23115*/;
assign _13432_ = _12759_ ^ _13434_ /*23118*/;
assign _13433_ = _13425_ & _13432_ /*23116*/;
assign _13430_ = _13431_ | _13433_ /*23114*/;
assign _13145_ = _13425_ ^ _13432_ /*23117*/;
assign _13439_ = D[56] ^ Q[30] /*23113*/;
assign _13436_ = _12760_ & _13439_ /*23109*/;
assign _13437_ = _12760_ ^ _13439_ /*23112*/;
assign _13438_ = _13430_ & _13437_ /*23110*/;
assign _13435_ = _13436_ | _13438_ /*23108*/;
assign _13146_ = _13430_ ^ _13437_ /*23111*/;
assign _13444_ = D[57] ^ Q[30] /*23107*/;
assign _13441_ = _12761_ & _13444_ /*23103*/;
assign _13442_ = _12761_ ^ _13444_ /*23106*/;
assign _13443_ = _13435_ & _13442_ /*23104*/;
assign _13440_ = _13441_ | _13443_ /*23102*/;
assign _13147_ = _13435_ ^ _13442_ /*23105*/;
assign _13449_ = D[58] ^ Q[30] /*23101*/;
assign _13446_ = _12762_ & _13449_ /*23097*/;
assign _13447_ = _12762_ ^ _13449_ /*23100*/;
assign _13448_ = _13440_ & _13447_ /*23098*/;
assign _13445_ = _13446_ | _13448_ /*23096*/;
assign _13148_ = _13440_ ^ _13447_ /*23099*/;
assign _13454_ = D[59] ^ Q[30] /*23095*/;
assign _13451_ = _12763_ & _13454_ /*23091*/;
assign _13452_ = _12763_ ^ _13454_ /*23094*/;
assign _13453_ = _13445_ & _13452_ /*23092*/;
assign _13450_ = _13451_ | _13453_ /*23090*/;
assign _13149_ = _13445_ ^ _13452_ /*23093*/;
assign _13459_ = D[60] ^ Q[30] /*23089*/;
assign _13456_ = _12764_ & _13459_ /*23085*/;
assign _13457_ = _12764_ ^ _13459_ /*23088*/;
assign _13458_ = _13450_ & _13457_ /*23086*/;
assign _13455_ = _13456_ | _13458_ /*23084*/;
assign _13150_ = _13450_ ^ _13457_ /*23087*/;
assign _13464_ = D[61] ^ Q[30] /*23083*/;
assign _13461_ = _12765_ & _13464_ /*23079*/;
assign _13462_ = _12765_ ^ _13464_ /*23082*/;
assign _13463_ = _13455_ & _13462_ /*23080*/;
assign _13460_ = _13461_ | _13463_ /*23078*/;
assign _13151_ = _13455_ ^ _13462_ /*23081*/;
assign _13469_ = D[62] ^ Q[30] /*23077*/;
assign _13466_ = _12766_ & _13469_ /*23073*/;
assign _13467_ = _12766_ ^ _13469_ /*23076*/;
assign _13468_ = _13460_ & _13467_ /*23074*/;
assign _13465_ = _13466_ | _13468_ /*23072*/;
assign _13152_ = _13460_ ^ _13467_ /*23075*/;
assign _13473_ = zeroWire ^ Q[30] /*23071*/;
assign _13470_ = _12767_ & _13473_ /*23067*/;
assign _13471_ = _12767_ ^ _13473_ /*23070*/;
assign _13472_ = _13465_ & _13471_ /*23068*/;
assign Q[29] = _13470_ | _13472_ /*23066*/;
assign _13153_ = _13465_ ^ _13471_ /*23069*/;
assign _13544_ = D[0] ^ Q[29] /*22680*/;
assign _13541_ = R_0[28] & _13544_ /*22676*/;
assign _13542_ = R_0[28] ^ _13544_ /*22679*/;
assign _13543_ = Q[29] & _13542_ /*22677*/;
assign _13540_ = _13541_ | _13543_ /*22675*/;
assign _13475_ = Q[29] ^ _13542_ /*22678*/;
assign _13549_ = D[1] ^ Q[29] /*22674*/;
assign _13546_ = _13090_ & _13549_ /*22670*/;
assign _13547_ = _13090_ ^ _13549_ /*22673*/;
assign _13548_ = _13540_ & _13547_ /*22671*/;
assign _13545_ = _13546_ | _13548_ /*22669*/;
assign _13476_ = _13540_ ^ _13547_ /*22672*/;
assign _13554_ = D[2] ^ Q[29] /*22668*/;
assign _13551_ = _13091_ & _13554_ /*22664*/;
assign _13552_ = _13091_ ^ _13554_ /*22667*/;
assign _13553_ = _13545_ & _13552_ /*22665*/;
assign _13550_ = _13551_ | _13553_ /*22663*/;
assign _13477_ = _13545_ ^ _13552_ /*22666*/;
assign _13559_ = D[3] ^ Q[29] /*22662*/;
assign _13556_ = _13092_ & _13559_ /*22658*/;
assign _13557_ = _13092_ ^ _13559_ /*22661*/;
assign _13558_ = _13550_ & _13557_ /*22659*/;
assign _13555_ = _13556_ | _13558_ /*22657*/;
assign _13478_ = _13550_ ^ _13557_ /*22660*/;
assign _13564_ = D[4] ^ Q[29] /*22656*/;
assign _13561_ = _13093_ & _13564_ /*22652*/;
assign _13562_ = _13093_ ^ _13564_ /*22655*/;
assign _13563_ = _13555_ & _13562_ /*22653*/;
assign _13560_ = _13561_ | _13563_ /*22651*/;
assign _13479_ = _13555_ ^ _13562_ /*22654*/;
assign _13569_ = D[5] ^ Q[29] /*22650*/;
assign _13566_ = _13094_ & _13569_ /*22646*/;
assign _13567_ = _13094_ ^ _13569_ /*22649*/;
assign _13568_ = _13560_ & _13567_ /*22647*/;
assign _13565_ = _13566_ | _13568_ /*22645*/;
assign _13480_ = _13560_ ^ _13567_ /*22648*/;
assign _13574_ = D[6] ^ Q[29] /*22644*/;
assign _13571_ = _13095_ & _13574_ /*22640*/;
assign _13572_ = _13095_ ^ _13574_ /*22643*/;
assign _13573_ = _13565_ & _13572_ /*22641*/;
assign _13570_ = _13571_ | _13573_ /*22639*/;
assign _13481_ = _13565_ ^ _13572_ /*22642*/;
assign _13579_ = D[7] ^ Q[29] /*22638*/;
assign _13576_ = _13096_ & _13579_ /*22634*/;
assign _13577_ = _13096_ ^ _13579_ /*22637*/;
assign _13578_ = _13570_ & _13577_ /*22635*/;
assign _13575_ = _13576_ | _13578_ /*22633*/;
assign _13482_ = _13570_ ^ _13577_ /*22636*/;
assign _13584_ = D[8] ^ Q[29] /*22632*/;
assign _13581_ = _13097_ & _13584_ /*22628*/;
assign _13582_ = _13097_ ^ _13584_ /*22631*/;
assign _13583_ = _13575_ & _13582_ /*22629*/;
assign _13580_ = _13581_ | _13583_ /*22627*/;
assign _13483_ = _13575_ ^ _13582_ /*22630*/;
assign _13589_ = D[9] ^ Q[29] /*22626*/;
assign _13586_ = _13098_ & _13589_ /*22622*/;
assign _13587_ = _13098_ ^ _13589_ /*22625*/;
assign _13588_ = _13580_ & _13587_ /*22623*/;
assign _13585_ = _13586_ | _13588_ /*22621*/;
assign _13484_ = _13580_ ^ _13587_ /*22624*/;
assign _13594_ = D[10] ^ Q[29] /*22620*/;
assign _13591_ = _13099_ & _13594_ /*22616*/;
assign _13592_ = _13099_ ^ _13594_ /*22619*/;
assign _13593_ = _13585_ & _13592_ /*22617*/;
assign _13590_ = _13591_ | _13593_ /*22615*/;
assign _13485_ = _13585_ ^ _13592_ /*22618*/;
assign _13599_ = D[11] ^ Q[29] /*22614*/;
assign _13596_ = _13100_ & _13599_ /*22610*/;
assign _13597_ = _13100_ ^ _13599_ /*22613*/;
assign _13598_ = _13590_ & _13597_ /*22611*/;
assign _13595_ = _13596_ | _13598_ /*22609*/;
assign _13486_ = _13590_ ^ _13597_ /*22612*/;
assign _13604_ = D[12] ^ Q[29] /*22608*/;
assign _13601_ = _13101_ & _13604_ /*22604*/;
assign _13602_ = _13101_ ^ _13604_ /*22607*/;
assign _13603_ = _13595_ & _13602_ /*22605*/;
assign _13600_ = _13601_ | _13603_ /*22603*/;
assign _13487_ = _13595_ ^ _13602_ /*22606*/;
assign _13609_ = D[13] ^ Q[29] /*22602*/;
assign _13606_ = _13102_ & _13609_ /*22598*/;
assign _13607_ = _13102_ ^ _13609_ /*22601*/;
assign _13608_ = _13600_ & _13607_ /*22599*/;
assign _13605_ = _13606_ | _13608_ /*22597*/;
assign _13488_ = _13600_ ^ _13607_ /*22600*/;
assign _13614_ = D[14] ^ Q[29] /*22596*/;
assign _13611_ = _13103_ & _13614_ /*22592*/;
assign _13612_ = _13103_ ^ _13614_ /*22595*/;
assign _13613_ = _13605_ & _13612_ /*22593*/;
assign _13610_ = _13611_ | _13613_ /*22591*/;
assign _13489_ = _13605_ ^ _13612_ /*22594*/;
assign _13619_ = D[15] ^ Q[29] /*22590*/;
assign _13616_ = _13104_ & _13619_ /*22586*/;
assign _13617_ = _13104_ ^ _13619_ /*22589*/;
assign _13618_ = _13610_ & _13617_ /*22587*/;
assign _13615_ = _13616_ | _13618_ /*22585*/;
assign _13490_ = _13610_ ^ _13617_ /*22588*/;
assign _13624_ = D[16] ^ Q[29] /*22584*/;
assign _13621_ = _13105_ & _13624_ /*22580*/;
assign _13622_ = _13105_ ^ _13624_ /*22583*/;
assign _13623_ = _13615_ & _13622_ /*22581*/;
assign _13620_ = _13621_ | _13623_ /*22579*/;
assign _13491_ = _13615_ ^ _13622_ /*22582*/;
assign _13629_ = D[17] ^ Q[29] /*22578*/;
assign _13626_ = _13106_ & _13629_ /*22574*/;
assign _13627_ = _13106_ ^ _13629_ /*22577*/;
assign _13628_ = _13620_ & _13627_ /*22575*/;
assign _13625_ = _13626_ | _13628_ /*22573*/;
assign _13492_ = _13620_ ^ _13627_ /*22576*/;
assign _13634_ = D[18] ^ Q[29] /*22572*/;
assign _13631_ = _13107_ & _13634_ /*22568*/;
assign _13632_ = _13107_ ^ _13634_ /*22571*/;
assign _13633_ = _13625_ & _13632_ /*22569*/;
assign _13630_ = _13631_ | _13633_ /*22567*/;
assign _13493_ = _13625_ ^ _13632_ /*22570*/;
assign _13639_ = D[19] ^ Q[29] /*22566*/;
assign _13636_ = _13108_ & _13639_ /*22562*/;
assign _13637_ = _13108_ ^ _13639_ /*22565*/;
assign _13638_ = _13630_ & _13637_ /*22563*/;
assign _13635_ = _13636_ | _13638_ /*22561*/;
assign _13494_ = _13630_ ^ _13637_ /*22564*/;
assign _13644_ = D[20] ^ Q[29] /*22560*/;
assign _13641_ = _13109_ & _13644_ /*22556*/;
assign _13642_ = _13109_ ^ _13644_ /*22559*/;
assign _13643_ = _13635_ & _13642_ /*22557*/;
assign _13640_ = _13641_ | _13643_ /*22555*/;
assign _13495_ = _13635_ ^ _13642_ /*22558*/;
assign _13649_ = D[21] ^ Q[29] /*22554*/;
assign _13646_ = _13110_ & _13649_ /*22550*/;
assign _13647_ = _13110_ ^ _13649_ /*22553*/;
assign _13648_ = _13640_ & _13647_ /*22551*/;
assign _13645_ = _13646_ | _13648_ /*22549*/;
assign _13496_ = _13640_ ^ _13647_ /*22552*/;
assign _13654_ = D[22] ^ Q[29] /*22548*/;
assign _13651_ = _13111_ & _13654_ /*22544*/;
assign _13652_ = _13111_ ^ _13654_ /*22547*/;
assign _13653_ = _13645_ & _13652_ /*22545*/;
assign _13650_ = _13651_ | _13653_ /*22543*/;
assign _13497_ = _13645_ ^ _13652_ /*22546*/;
assign _13659_ = D[23] ^ Q[29] /*22542*/;
assign _13656_ = _13112_ & _13659_ /*22538*/;
assign _13657_ = _13112_ ^ _13659_ /*22541*/;
assign _13658_ = _13650_ & _13657_ /*22539*/;
assign _13655_ = _13656_ | _13658_ /*22537*/;
assign _13498_ = _13650_ ^ _13657_ /*22540*/;
assign _13664_ = D[24] ^ Q[29] /*22536*/;
assign _13661_ = _13113_ & _13664_ /*22532*/;
assign _13662_ = _13113_ ^ _13664_ /*22535*/;
assign _13663_ = _13655_ & _13662_ /*22533*/;
assign _13660_ = _13661_ | _13663_ /*22531*/;
assign _13499_ = _13655_ ^ _13662_ /*22534*/;
assign _13669_ = D[25] ^ Q[29] /*22530*/;
assign _13666_ = _13114_ & _13669_ /*22526*/;
assign _13667_ = _13114_ ^ _13669_ /*22529*/;
assign _13668_ = _13660_ & _13667_ /*22527*/;
assign _13665_ = _13666_ | _13668_ /*22525*/;
assign _13500_ = _13660_ ^ _13667_ /*22528*/;
assign _13674_ = D[26] ^ Q[29] /*22524*/;
assign _13671_ = _13115_ & _13674_ /*22520*/;
assign _13672_ = _13115_ ^ _13674_ /*22523*/;
assign _13673_ = _13665_ & _13672_ /*22521*/;
assign _13670_ = _13671_ | _13673_ /*22519*/;
assign _13501_ = _13665_ ^ _13672_ /*22522*/;
assign _13679_ = D[27] ^ Q[29] /*22518*/;
assign _13676_ = _13116_ & _13679_ /*22514*/;
assign _13677_ = _13116_ ^ _13679_ /*22517*/;
assign _13678_ = _13670_ & _13677_ /*22515*/;
assign _13675_ = _13676_ | _13678_ /*22513*/;
assign _13502_ = _13670_ ^ _13677_ /*22516*/;
assign _13684_ = D[28] ^ Q[29] /*22512*/;
assign _13681_ = _13117_ & _13684_ /*22508*/;
assign _13682_ = _13117_ ^ _13684_ /*22511*/;
assign _13683_ = _13675_ & _13682_ /*22509*/;
assign _13680_ = _13681_ | _13683_ /*22507*/;
assign _13503_ = _13675_ ^ _13682_ /*22510*/;
assign _13689_ = D[29] ^ Q[29] /*22506*/;
assign _13686_ = _13118_ & _13689_ /*22502*/;
assign _13687_ = _13118_ ^ _13689_ /*22505*/;
assign _13688_ = _13680_ & _13687_ /*22503*/;
assign _13685_ = _13686_ | _13688_ /*22501*/;
assign _13504_ = _13680_ ^ _13687_ /*22504*/;
assign _13694_ = D[30] ^ Q[29] /*22500*/;
assign _13691_ = _13119_ & _13694_ /*22496*/;
assign _13692_ = _13119_ ^ _13694_ /*22499*/;
assign _13693_ = _13685_ & _13692_ /*22497*/;
assign _13690_ = _13691_ | _13693_ /*22495*/;
assign _13505_ = _13685_ ^ _13692_ /*22498*/;
assign _13699_ = D[31] ^ Q[29] /*22494*/;
assign _13696_ = _13120_ & _13699_ /*22490*/;
assign _13697_ = _13120_ ^ _13699_ /*22493*/;
assign _13698_ = _13690_ & _13697_ /*22491*/;
assign _13695_ = _13696_ | _13698_ /*22489*/;
assign _13506_ = _13690_ ^ _13697_ /*22492*/;
assign _13704_ = D[32] ^ Q[29] /*22488*/;
assign _13701_ = _13121_ & _13704_ /*22484*/;
assign _13702_ = _13121_ ^ _13704_ /*22487*/;
assign _13703_ = _13695_ & _13702_ /*22485*/;
assign _13700_ = _13701_ | _13703_ /*22483*/;
assign _13507_ = _13695_ ^ _13702_ /*22486*/;
assign _13709_ = D[33] ^ Q[29] /*22482*/;
assign _13706_ = _13122_ & _13709_ /*22478*/;
assign _13707_ = _13122_ ^ _13709_ /*22481*/;
assign _13708_ = _13700_ & _13707_ /*22479*/;
assign _13705_ = _13706_ | _13708_ /*22477*/;
assign _13508_ = _13700_ ^ _13707_ /*22480*/;
assign _13714_ = D[34] ^ Q[29] /*22476*/;
assign _13711_ = _13123_ & _13714_ /*22472*/;
assign _13712_ = _13123_ ^ _13714_ /*22475*/;
assign _13713_ = _13705_ & _13712_ /*22473*/;
assign _13710_ = _13711_ | _13713_ /*22471*/;
assign _13509_ = _13705_ ^ _13712_ /*22474*/;
assign _13719_ = D[35] ^ Q[29] /*22470*/;
assign _13716_ = _13124_ & _13719_ /*22466*/;
assign _13717_ = _13124_ ^ _13719_ /*22469*/;
assign _13718_ = _13710_ & _13717_ /*22467*/;
assign _13715_ = _13716_ | _13718_ /*22465*/;
assign _13510_ = _13710_ ^ _13717_ /*22468*/;
assign _13724_ = D[36] ^ Q[29] /*22464*/;
assign _13721_ = _13125_ & _13724_ /*22460*/;
assign _13722_ = _13125_ ^ _13724_ /*22463*/;
assign _13723_ = _13715_ & _13722_ /*22461*/;
assign _13720_ = _13721_ | _13723_ /*22459*/;
assign _13511_ = _13715_ ^ _13722_ /*22462*/;
assign _13729_ = D[37] ^ Q[29] /*22458*/;
assign _13726_ = _13126_ & _13729_ /*22454*/;
assign _13727_ = _13126_ ^ _13729_ /*22457*/;
assign _13728_ = _13720_ & _13727_ /*22455*/;
assign _13725_ = _13726_ | _13728_ /*22453*/;
assign _13512_ = _13720_ ^ _13727_ /*22456*/;
assign _13734_ = D[38] ^ Q[29] /*22452*/;
assign _13731_ = _13127_ & _13734_ /*22448*/;
assign _13732_ = _13127_ ^ _13734_ /*22451*/;
assign _13733_ = _13725_ & _13732_ /*22449*/;
assign _13730_ = _13731_ | _13733_ /*22447*/;
assign _13513_ = _13725_ ^ _13732_ /*22450*/;
assign _13739_ = D[39] ^ Q[29] /*22446*/;
assign _13736_ = _13128_ & _13739_ /*22442*/;
assign _13737_ = _13128_ ^ _13739_ /*22445*/;
assign _13738_ = _13730_ & _13737_ /*22443*/;
assign _13735_ = _13736_ | _13738_ /*22441*/;
assign _13514_ = _13730_ ^ _13737_ /*22444*/;
assign _13744_ = D[40] ^ Q[29] /*22440*/;
assign _13741_ = _13129_ & _13744_ /*22436*/;
assign _13742_ = _13129_ ^ _13744_ /*22439*/;
assign _13743_ = _13735_ & _13742_ /*22437*/;
assign _13740_ = _13741_ | _13743_ /*22435*/;
assign _13515_ = _13735_ ^ _13742_ /*22438*/;
assign _13749_ = D[41] ^ Q[29] /*22434*/;
assign _13746_ = _13130_ & _13749_ /*22430*/;
assign _13747_ = _13130_ ^ _13749_ /*22433*/;
assign _13748_ = _13740_ & _13747_ /*22431*/;
assign _13745_ = _13746_ | _13748_ /*22429*/;
assign _13516_ = _13740_ ^ _13747_ /*22432*/;
assign _13754_ = D[42] ^ Q[29] /*22428*/;
assign _13751_ = _13131_ & _13754_ /*22424*/;
assign _13752_ = _13131_ ^ _13754_ /*22427*/;
assign _13753_ = _13745_ & _13752_ /*22425*/;
assign _13750_ = _13751_ | _13753_ /*22423*/;
assign _13517_ = _13745_ ^ _13752_ /*22426*/;
assign _13759_ = D[43] ^ Q[29] /*22422*/;
assign _13756_ = _13132_ & _13759_ /*22418*/;
assign _13757_ = _13132_ ^ _13759_ /*22421*/;
assign _13758_ = _13750_ & _13757_ /*22419*/;
assign _13755_ = _13756_ | _13758_ /*22417*/;
assign _13518_ = _13750_ ^ _13757_ /*22420*/;
assign _13764_ = D[44] ^ Q[29] /*22416*/;
assign _13761_ = _13133_ & _13764_ /*22412*/;
assign _13762_ = _13133_ ^ _13764_ /*22415*/;
assign _13763_ = _13755_ & _13762_ /*22413*/;
assign _13760_ = _13761_ | _13763_ /*22411*/;
assign _13519_ = _13755_ ^ _13762_ /*22414*/;
assign _13769_ = D[45] ^ Q[29] /*22410*/;
assign _13766_ = _13134_ & _13769_ /*22406*/;
assign _13767_ = _13134_ ^ _13769_ /*22409*/;
assign _13768_ = _13760_ & _13767_ /*22407*/;
assign _13765_ = _13766_ | _13768_ /*22405*/;
assign _13520_ = _13760_ ^ _13767_ /*22408*/;
assign _13774_ = D[46] ^ Q[29] /*22404*/;
assign _13771_ = _13135_ & _13774_ /*22400*/;
assign _13772_ = _13135_ ^ _13774_ /*22403*/;
assign _13773_ = _13765_ & _13772_ /*22401*/;
assign _13770_ = _13771_ | _13773_ /*22399*/;
assign _13521_ = _13765_ ^ _13772_ /*22402*/;
assign _13779_ = D[47] ^ Q[29] /*22398*/;
assign _13776_ = _13136_ & _13779_ /*22394*/;
assign _13777_ = _13136_ ^ _13779_ /*22397*/;
assign _13778_ = _13770_ & _13777_ /*22395*/;
assign _13775_ = _13776_ | _13778_ /*22393*/;
assign _13522_ = _13770_ ^ _13777_ /*22396*/;
assign _13784_ = D[48] ^ Q[29] /*22392*/;
assign _13781_ = _13137_ & _13784_ /*22388*/;
assign _13782_ = _13137_ ^ _13784_ /*22391*/;
assign _13783_ = _13775_ & _13782_ /*22389*/;
assign _13780_ = _13781_ | _13783_ /*22387*/;
assign _13523_ = _13775_ ^ _13782_ /*22390*/;
assign _13789_ = D[49] ^ Q[29] /*22386*/;
assign _13786_ = _13138_ & _13789_ /*22382*/;
assign _13787_ = _13138_ ^ _13789_ /*22385*/;
assign _13788_ = _13780_ & _13787_ /*22383*/;
assign _13785_ = _13786_ | _13788_ /*22381*/;
assign _13524_ = _13780_ ^ _13787_ /*22384*/;
assign _13794_ = D[50] ^ Q[29] /*22380*/;
assign _13791_ = _13139_ & _13794_ /*22376*/;
assign _13792_ = _13139_ ^ _13794_ /*22379*/;
assign _13793_ = _13785_ & _13792_ /*22377*/;
assign _13790_ = _13791_ | _13793_ /*22375*/;
assign _13525_ = _13785_ ^ _13792_ /*22378*/;
assign _13799_ = D[51] ^ Q[29] /*22374*/;
assign _13796_ = _13140_ & _13799_ /*22370*/;
assign _13797_ = _13140_ ^ _13799_ /*22373*/;
assign _13798_ = _13790_ & _13797_ /*22371*/;
assign _13795_ = _13796_ | _13798_ /*22369*/;
assign _13526_ = _13790_ ^ _13797_ /*22372*/;
assign _13804_ = D[52] ^ Q[29] /*22368*/;
assign _13801_ = _13141_ & _13804_ /*22364*/;
assign _13802_ = _13141_ ^ _13804_ /*22367*/;
assign _13803_ = _13795_ & _13802_ /*22365*/;
assign _13800_ = _13801_ | _13803_ /*22363*/;
assign _13527_ = _13795_ ^ _13802_ /*22366*/;
assign _13809_ = D[53] ^ Q[29] /*22362*/;
assign _13806_ = _13142_ & _13809_ /*22358*/;
assign _13807_ = _13142_ ^ _13809_ /*22361*/;
assign _13808_ = _13800_ & _13807_ /*22359*/;
assign _13805_ = _13806_ | _13808_ /*22357*/;
assign _13528_ = _13800_ ^ _13807_ /*22360*/;
assign _13814_ = D[54] ^ Q[29] /*22356*/;
assign _13811_ = _13143_ & _13814_ /*22352*/;
assign _13812_ = _13143_ ^ _13814_ /*22355*/;
assign _13813_ = _13805_ & _13812_ /*22353*/;
assign _13810_ = _13811_ | _13813_ /*22351*/;
assign _13529_ = _13805_ ^ _13812_ /*22354*/;
assign _13819_ = D[55] ^ Q[29] /*22350*/;
assign _13816_ = _13144_ & _13819_ /*22346*/;
assign _13817_ = _13144_ ^ _13819_ /*22349*/;
assign _13818_ = _13810_ & _13817_ /*22347*/;
assign _13815_ = _13816_ | _13818_ /*22345*/;
assign _13530_ = _13810_ ^ _13817_ /*22348*/;
assign _13824_ = D[56] ^ Q[29] /*22344*/;
assign _13821_ = _13145_ & _13824_ /*22340*/;
assign _13822_ = _13145_ ^ _13824_ /*22343*/;
assign _13823_ = _13815_ & _13822_ /*22341*/;
assign _13820_ = _13821_ | _13823_ /*22339*/;
assign _13531_ = _13815_ ^ _13822_ /*22342*/;
assign _13829_ = D[57] ^ Q[29] /*22338*/;
assign _13826_ = _13146_ & _13829_ /*22334*/;
assign _13827_ = _13146_ ^ _13829_ /*22337*/;
assign _13828_ = _13820_ & _13827_ /*22335*/;
assign _13825_ = _13826_ | _13828_ /*22333*/;
assign _13532_ = _13820_ ^ _13827_ /*22336*/;
assign _13834_ = D[58] ^ Q[29] /*22332*/;
assign _13831_ = _13147_ & _13834_ /*22328*/;
assign _13832_ = _13147_ ^ _13834_ /*22331*/;
assign _13833_ = _13825_ & _13832_ /*22329*/;
assign _13830_ = _13831_ | _13833_ /*22327*/;
assign _13533_ = _13825_ ^ _13832_ /*22330*/;
assign _13839_ = D[59] ^ Q[29] /*22326*/;
assign _13836_ = _13148_ & _13839_ /*22322*/;
assign _13837_ = _13148_ ^ _13839_ /*22325*/;
assign _13838_ = _13830_ & _13837_ /*22323*/;
assign _13835_ = _13836_ | _13838_ /*22321*/;
assign _13534_ = _13830_ ^ _13837_ /*22324*/;
assign _13844_ = D[60] ^ Q[29] /*22320*/;
assign _13841_ = _13149_ & _13844_ /*22316*/;
assign _13842_ = _13149_ ^ _13844_ /*22319*/;
assign _13843_ = _13835_ & _13842_ /*22317*/;
assign _13840_ = _13841_ | _13843_ /*22315*/;
assign _13535_ = _13835_ ^ _13842_ /*22318*/;
assign _13849_ = D[61] ^ Q[29] /*22314*/;
assign _13846_ = _13150_ & _13849_ /*22310*/;
assign _13847_ = _13150_ ^ _13849_ /*22313*/;
assign _13848_ = _13840_ & _13847_ /*22311*/;
assign _13845_ = _13846_ | _13848_ /*22309*/;
assign _13536_ = _13840_ ^ _13847_ /*22312*/;
assign _13854_ = D[62] ^ Q[29] /*22308*/;
assign _13851_ = _13151_ & _13854_ /*22304*/;
assign _13852_ = _13151_ ^ _13854_ /*22307*/;
assign _13853_ = _13845_ & _13852_ /*22305*/;
assign _13850_ = _13851_ | _13853_ /*22303*/;
assign _13537_ = _13845_ ^ _13852_ /*22306*/;
assign _13858_ = zeroWire ^ Q[29] /*22302*/;
assign _13855_ = _13152_ & _13858_ /*22298*/;
assign _13856_ = _13152_ ^ _13858_ /*22301*/;
assign _13857_ = _13850_ & _13856_ /*22299*/;
assign Q[28] = _13855_ | _13857_ /*22297*/;
assign _13538_ = _13850_ ^ _13856_ /*22300*/;
assign _13929_ = D[0] ^ Q[28] /*21911*/;
assign _13926_ = R_0[27] & _13929_ /*21907*/;
assign _13927_ = R_0[27] ^ _13929_ /*21910*/;
assign _13928_ = Q[28] & _13927_ /*21908*/;
assign _13925_ = _13926_ | _13928_ /*21906*/;
assign _13860_ = Q[28] ^ _13927_ /*21909*/;
assign _13934_ = D[1] ^ Q[28] /*21905*/;
assign _13931_ = _13475_ & _13934_ /*21901*/;
assign _13932_ = _13475_ ^ _13934_ /*21904*/;
assign _13933_ = _13925_ & _13932_ /*21902*/;
assign _13930_ = _13931_ | _13933_ /*21900*/;
assign _13861_ = _13925_ ^ _13932_ /*21903*/;
assign _13939_ = D[2] ^ Q[28] /*21899*/;
assign _13936_ = _13476_ & _13939_ /*21895*/;
assign _13937_ = _13476_ ^ _13939_ /*21898*/;
assign _13938_ = _13930_ & _13937_ /*21896*/;
assign _13935_ = _13936_ | _13938_ /*21894*/;
assign _13862_ = _13930_ ^ _13937_ /*21897*/;
assign _13944_ = D[3] ^ Q[28] /*21893*/;
assign _13941_ = _13477_ & _13944_ /*21889*/;
assign _13942_ = _13477_ ^ _13944_ /*21892*/;
assign _13943_ = _13935_ & _13942_ /*21890*/;
assign _13940_ = _13941_ | _13943_ /*21888*/;
assign _13863_ = _13935_ ^ _13942_ /*21891*/;
assign _13949_ = D[4] ^ Q[28] /*21887*/;
assign _13946_ = _13478_ & _13949_ /*21883*/;
assign _13947_ = _13478_ ^ _13949_ /*21886*/;
assign _13948_ = _13940_ & _13947_ /*21884*/;
assign _13945_ = _13946_ | _13948_ /*21882*/;
assign _13864_ = _13940_ ^ _13947_ /*21885*/;
assign _13954_ = D[5] ^ Q[28] /*21881*/;
assign _13951_ = _13479_ & _13954_ /*21877*/;
assign _13952_ = _13479_ ^ _13954_ /*21880*/;
assign _13953_ = _13945_ & _13952_ /*21878*/;
assign _13950_ = _13951_ | _13953_ /*21876*/;
assign _13865_ = _13945_ ^ _13952_ /*21879*/;
assign _13959_ = D[6] ^ Q[28] /*21875*/;
assign _13956_ = _13480_ & _13959_ /*21871*/;
assign _13957_ = _13480_ ^ _13959_ /*21874*/;
assign _13958_ = _13950_ & _13957_ /*21872*/;
assign _13955_ = _13956_ | _13958_ /*21870*/;
assign _13866_ = _13950_ ^ _13957_ /*21873*/;
assign _13964_ = D[7] ^ Q[28] /*21869*/;
assign _13961_ = _13481_ & _13964_ /*21865*/;
assign _13962_ = _13481_ ^ _13964_ /*21868*/;
assign _13963_ = _13955_ & _13962_ /*21866*/;
assign _13960_ = _13961_ | _13963_ /*21864*/;
assign _13867_ = _13955_ ^ _13962_ /*21867*/;
assign _13969_ = D[8] ^ Q[28] /*21863*/;
assign _13966_ = _13482_ & _13969_ /*21859*/;
assign _13967_ = _13482_ ^ _13969_ /*21862*/;
assign _13968_ = _13960_ & _13967_ /*21860*/;
assign _13965_ = _13966_ | _13968_ /*21858*/;
assign _13868_ = _13960_ ^ _13967_ /*21861*/;
assign _13974_ = D[9] ^ Q[28] /*21857*/;
assign _13971_ = _13483_ & _13974_ /*21853*/;
assign _13972_ = _13483_ ^ _13974_ /*21856*/;
assign _13973_ = _13965_ & _13972_ /*21854*/;
assign _13970_ = _13971_ | _13973_ /*21852*/;
assign _13869_ = _13965_ ^ _13972_ /*21855*/;
assign _13979_ = D[10] ^ Q[28] /*21851*/;
assign _13976_ = _13484_ & _13979_ /*21847*/;
assign _13977_ = _13484_ ^ _13979_ /*21850*/;
assign _13978_ = _13970_ & _13977_ /*21848*/;
assign _13975_ = _13976_ | _13978_ /*21846*/;
assign _13870_ = _13970_ ^ _13977_ /*21849*/;
assign _13984_ = D[11] ^ Q[28] /*21845*/;
assign _13981_ = _13485_ & _13984_ /*21841*/;
assign _13982_ = _13485_ ^ _13984_ /*21844*/;
assign _13983_ = _13975_ & _13982_ /*21842*/;
assign _13980_ = _13981_ | _13983_ /*21840*/;
assign _13871_ = _13975_ ^ _13982_ /*21843*/;
assign _13989_ = D[12] ^ Q[28] /*21839*/;
assign _13986_ = _13486_ & _13989_ /*21835*/;
assign _13987_ = _13486_ ^ _13989_ /*21838*/;
assign _13988_ = _13980_ & _13987_ /*21836*/;
assign _13985_ = _13986_ | _13988_ /*21834*/;
assign _13872_ = _13980_ ^ _13987_ /*21837*/;
assign _13994_ = D[13] ^ Q[28] /*21833*/;
assign _13991_ = _13487_ & _13994_ /*21829*/;
assign _13992_ = _13487_ ^ _13994_ /*21832*/;
assign _13993_ = _13985_ & _13992_ /*21830*/;
assign _13990_ = _13991_ | _13993_ /*21828*/;
assign _13873_ = _13985_ ^ _13992_ /*21831*/;
assign _13999_ = D[14] ^ Q[28] /*21827*/;
assign _13996_ = _13488_ & _13999_ /*21823*/;
assign _13997_ = _13488_ ^ _13999_ /*21826*/;
assign _13998_ = _13990_ & _13997_ /*21824*/;
assign _13995_ = _13996_ | _13998_ /*21822*/;
assign _13874_ = _13990_ ^ _13997_ /*21825*/;
assign _14004_ = D[15] ^ Q[28] /*21821*/;
assign _14001_ = _13489_ & _14004_ /*21817*/;
assign _14002_ = _13489_ ^ _14004_ /*21820*/;
assign _14003_ = _13995_ & _14002_ /*21818*/;
assign _14000_ = _14001_ | _14003_ /*21816*/;
assign _13875_ = _13995_ ^ _14002_ /*21819*/;
assign _14009_ = D[16] ^ Q[28] /*21815*/;
assign _14006_ = _13490_ & _14009_ /*21811*/;
assign _14007_ = _13490_ ^ _14009_ /*21814*/;
assign _14008_ = _14000_ & _14007_ /*21812*/;
assign _14005_ = _14006_ | _14008_ /*21810*/;
assign _13876_ = _14000_ ^ _14007_ /*21813*/;
assign _14014_ = D[17] ^ Q[28] /*21809*/;
assign _14011_ = _13491_ & _14014_ /*21805*/;
assign _14012_ = _13491_ ^ _14014_ /*21808*/;
assign _14013_ = _14005_ & _14012_ /*21806*/;
assign _14010_ = _14011_ | _14013_ /*21804*/;
assign _13877_ = _14005_ ^ _14012_ /*21807*/;
assign _14019_ = D[18] ^ Q[28] /*21803*/;
assign _14016_ = _13492_ & _14019_ /*21799*/;
assign _14017_ = _13492_ ^ _14019_ /*21802*/;
assign _14018_ = _14010_ & _14017_ /*21800*/;
assign _14015_ = _14016_ | _14018_ /*21798*/;
assign _13878_ = _14010_ ^ _14017_ /*21801*/;
assign _14024_ = D[19] ^ Q[28] /*21797*/;
assign _14021_ = _13493_ & _14024_ /*21793*/;
assign _14022_ = _13493_ ^ _14024_ /*21796*/;
assign _14023_ = _14015_ & _14022_ /*21794*/;
assign _14020_ = _14021_ | _14023_ /*21792*/;
assign _13879_ = _14015_ ^ _14022_ /*21795*/;
assign _14029_ = D[20] ^ Q[28] /*21791*/;
assign _14026_ = _13494_ & _14029_ /*21787*/;
assign _14027_ = _13494_ ^ _14029_ /*21790*/;
assign _14028_ = _14020_ & _14027_ /*21788*/;
assign _14025_ = _14026_ | _14028_ /*21786*/;
assign _13880_ = _14020_ ^ _14027_ /*21789*/;
assign _14034_ = D[21] ^ Q[28] /*21785*/;
assign _14031_ = _13495_ & _14034_ /*21781*/;
assign _14032_ = _13495_ ^ _14034_ /*21784*/;
assign _14033_ = _14025_ & _14032_ /*21782*/;
assign _14030_ = _14031_ | _14033_ /*21780*/;
assign _13881_ = _14025_ ^ _14032_ /*21783*/;
assign _14039_ = D[22] ^ Q[28] /*21779*/;
assign _14036_ = _13496_ & _14039_ /*21775*/;
assign _14037_ = _13496_ ^ _14039_ /*21778*/;
assign _14038_ = _14030_ & _14037_ /*21776*/;
assign _14035_ = _14036_ | _14038_ /*21774*/;
assign _13882_ = _14030_ ^ _14037_ /*21777*/;
assign _14044_ = D[23] ^ Q[28] /*21773*/;
assign _14041_ = _13497_ & _14044_ /*21769*/;
assign _14042_ = _13497_ ^ _14044_ /*21772*/;
assign _14043_ = _14035_ & _14042_ /*21770*/;
assign _14040_ = _14041_ | _14043_ /*21768*/;
assign _13883_ = _14035_ ^ _14042_ /*21771*/;
assign _14049_ = D[24] ^ Q[28] /*21767*/;
assign _14046_ = _13498_ & _14049_ /*21763*/;
assign _14047_ = _13498_ ^ _14049_ /*21766*/;
assign _14048_ = _14040_ & _14047_ /*21764*/;
assign _14045_ = _14046_ | _14048_ /*21762*/;
assign _13884_ = _14040_ ^ _14047_ /*21765*/;
assign _14054_ = D[25] ^ Q[28] /*21761*/;
assign _14051_ = _13499_ & _14054_ /*21757*/;
assign _14052_ = _13499_ ^ _14054_ /*21760*/;
assign _14053_ = _14045_ & _14052_ /*21758*/;
assign _14050_ = _14051_ | _14053_ /*21756*/;
assign _13885_ = _14045_ ^ _14052_ /*21759*/;
assign _14059_ = D[26] ^ Q[28] /*21755*/;
assign _14056_ = _13500_ & _14059_ /*21751*/;
assign _14057_ = _13500_ ^ _14059_ /*21754*/;
assign _14058_ = _14050_ & _14057_ /*21752*/;
assign _14055_ = _14056_ | _14058_ /*21750*/;
assign _13886_ = _14050_ ^ _14057_ /*21753*/;
assign _14064_ = D[27] ^ Q[28] /*21749*/;
assign _14061_ = _13501_ & _14064_ /*21745*/;
assign _14062_ = _13501_ ^ _14064_ /*21748*/;
assign _14063_ = _14055_ & _14062_ /*21746*/;
assign _14060_ = _14061_ | _14063_ /*21744*/;
assign _13887_ = _14055_ ^ _14062_ /*21747*/;
assign _14069_ = D[28] ^ Q[28] /*21743*/;
assign _14066_ = _13502_ & _14069_ /*21739*/;
assign _14067_ = _13502_ ^ _14069_ /*21742*/;
assign _14068_ = _14060_ & _14067_ /*21740*/;
assign _14065_ = _14066_ | _14068_ /*21738*/;
assign _13888_ = _14060_ ^ _14067_ /*21741*/;
assign _14074_ = D[29] ^ Q[28] /*21737*/;
assign _14071_ = _13503_ & _14074_ /*21733*/;
assign _14072_ = _13503_ ^ _14074_ /*21736*/;
assign _14073_ = _14065_ & _14072_ /*21734*/;
assign _14070_ = _14071_ | _14073_ /*21732*/;
assign _13889_ = _14065_ ^ _14072_ /*21735*/;
assign _14079_ = D[30] ^ Q[28] /*21731*/;
assign _14076_ = _13504_ & _14079_ /*21727*/;
assign _14077_ = _13504_ ^ _14079_ /*21730*/;
assign _14078_ = _14070_ & _14077_ /*21728*/;
assign _14075_ = _14076_ | _14078_ /*21726*/;
assign _13890_ = _14070_ ^ _14077_ /*21729*/;
assign _14084_ = D[31] ^ Q[28] /*21725*/;
assign _14081_ = _13505_ & _14084_ /*21721*/;
assign _14082_ = _13505_ ^ _14084_ /*21724*/;
assign _14083_ = _14075_ & _14082_ /*21722*/;
assign _14080_ = _14081_ | _14083_ /*21720*/;
assign _13891_ = _14075_ ^ _14082_ /*21723*/;
assign _14089_ = D[32] ^ Q[28] /*21719*/;
assign _14086_ = _13506_ & _14089_ /*21715*/;
assign _14087_ = _13506_ ^ _14089_ /*21718*/;
assign _14088_ = _14080_ & _14087_ /*21716*/;
assign _14085_ = _14086_ | _14088_ /*21714*/;
assign _13892_ = _14080_ ^ _14087_ /*21717*/;
assign _14094_ = D[33] ^ Q[28] /*21713*/;
assign _14091_ = _13507_ & _14094_ /*21709*/;
assign _14092_ = _13507_ ^ _14094_ /*21712*/;
assign _14093_ = _14085_ & _14092_ /*21710*/;
assign _14090_ = _14091_ | _14093_ /*21708*/;
assign _13893_ = _14085_ ^ _14092_ /*21711*/;
assign _14099_ = D[34] ^ Q[28] /*21707*/;
assign _14096_ = _13508_ & _14099_ /*21703*/;
assign _14097_ = _13508_ ^ _14099_ /*21706*/;
assign _14098_ = _14090_ & _14097_ /*21704*/;
assign _14095_ = _14096_ | _14098_ /*21702*/;
assign _13894_ = _14090_ ^ _14097_ /*21705*/;
assign _14104_ = D[35] ^ Q[28] /*21701*/;
assign _14101_ = _13509_ & _14104_ /*21697*/;
assign _14102_ = _13509_ ^ _14104_ /*21700*/;
assign _14103_ = _14095_ & _14102_ /*21698*/;
assign _14100_ = _14101_ | _14103_ /*21696*/;
assign _13895_ = _14095_ ^ _14102_ /*21699*/;
assign _14109_ = D[36] ^ Q[28] /*21695*/;
assign _14106_ = _13510_ & _14109_ /*21691*/;
assign _14107_ = _13510_ ^ _14109_ /*21694*/;
assign _14108_ = _14100_ & _14107_ /*21692*/;
assign _14105_ = _14106_ | _14108_ /*21690*/;
assign _13896_ = _14100_ ^ _14107_ /*21693*/;
assign _14114_ = D[37] ^ Q[28] /*21689*/;
assign _14111_ = _13511_ & _14114_ /*21685*/;
assign _14112_ = _13511_ ^ _14114_ /*21688*/;
assign _14113_ = _14105_ & _14112_ /*21686*/;
assign _14110_ = _14111_ | _14113_ /*21684*/;
assign _13897_ = _14105_ ^ _14112_ /*21687*/;
assign _14119_ = D[38] ^ Q[28] /*21683*/;
assign _14116_ = _13512_ & _14119_ /*21679*/;
assign _14117_ = _13512_ ^ _14119_ /*21682*/;
assign _14118_ = _14110_ & _14117_ /*21680*/;
assign _14115_ = _14116_ | _14118_ /*21678*/;
assign _13898_ = _14110_ ^ _14117_ /*21681*/;
assign _14124_ = D[39] ^ Q[28] /*21677*/;
assign _14121_ = _13513_ & _14124_ /*21673*/;
assign _14122_ = _13513_ ^ _14124_ /*21676*/;
assign _14123_ = _14115_ & _14122_ /*21674*/;
assign _14120_ = _14121_ | _14123_ /*21672*/;
assign _13899_ = _14115_ ^ _14122_ /*21675*/;
assign _14129_ = D[40] ^ Q[28] /*21671*/;
assign _14126_ = _13514_ & _14129_ /*21667*/;
assign _14127_ = _13514_ ^ _14129_ /*21670*/;
assign _14128_ = _14120_ & _14127_ /*21668*/;
assign _14125_ = _14126_ | _14128_ /*21666*/;
assign _13900_ = _14120_ ^ _14127_ /*21669*/;
assign _14134_ = D[41] ^ Q[28] /*21665*/;
assign _14131_ = _13515_ & _14134_ /*21661*/;
assign _14132_ = _13515_ ^ _14134_ /*21664*/;
assign _14133_ = _14125_ & _14132_ /*21662*/;
assign _14130_ = _14131_ | _14133_ /*21660*/;
assign _13901_ = _14125_ ^ _14132_ /*21663*/;
assign _14139_ = D[42] ^ Q[28] /*21659*/;
assign _14136_ = _13516_ & _14139_ /*21655*/;
assign _14137_ = _13516_ ^ _14139_ /*21658*/;
assign _14138_ = _14130_ & _14137_ /*21656*/;
assign _14135_ = _14136_ | _14138_ /*21654*/;
assign _13902_ = _14130_ ^ _14137_ /*21657*/;
assign _14144_ = D[43] ^ Q[28] /*21653*/;
assign _14141_ = _13517_ & _14144_ /*21649*/;
assign _14142_ = _13517_ ^ _14144_ /*21652*/;
assign _14143_ = _14135_ & _14142_ /*21650*/;
assign _14140_ = _14141_ | _14143_ /*21648*/;
assign _13903_ = _14135_ ^ _14142_ /*21651*/;
assign _14149_ = D[44] ^ Q[28] /*21647*/;
assign _14146_ = _13518_ & _14149_ /*21643*/;
assign _14147_ = _13518_ ^ _14149_ /*21646*/;
assign _14148_ = _14140_ & _14147_ /*21644*/;
assign _14145_ = _14146_ | _14148_ /*21642*/;
assign _13904_ = _14140_ ^ _14147_ /*21645*/;
assign _14154_ = D[45] ^ Q[28] /*21641*/;
assign _14151_ = _13519_ & _14154_ /*21637*/;
assign _14152_ = _13519_ ^ _14154_ /*21640*/;
assign _14153_ = _14145_ & _14152_ /*21638*/;
assign _14150_ = _14151_ | _14153_ /*21636*/;
assign _13905_ = _14145_ ^ _14152_ /*21639*/;
assign _14159_ = D[46] ^ Q[28] /*21635*/;
assign _14156_ = _13520_ & _14159_ /*21631*/;
assign _14157_ = _13520_ ^ _14159_ /*21634*/;
assign _14158_ = _14150_ & _14157_ /*21632*/;
assign _14155_ = _14156_ | _14158_ /*21630*/;
assign _13906_ = _14150_ ^ _14157_ /*21633*/;
assign _14164_ = D[47] ^ Q[28] /*21629*/;
assign _14161_ = _13521_ & _14164_ /*21625*/;
assign _14162_ = _13521_ ^ _14164_ /*21628*/;
assign _14163_ = _14155_ & _14162_ /*21626*/;
assign _14160_ = _14161_ | _14163_ /*21624*/;
assign _13907_ = _14155_ ^ _14162_ /*21627*/;
assign _14169_ = D[48] ^ Q[28] /*21623*/;
assign _14166_ = _13522_ & _14169_ /*21619*/;
assign _14167_ = _13522_ ^ _14169_ /*21622*/;
assign _14168_ = _14160_ & _14167_ /*21620*/;
assign _14165_ = _14166_ | _14168_ /*21618*/;
assign _13908_ = _14160_ ^ _14167_ /*21621*/;
assign _14174_ = D[49] ^ Q[28] /*21617*/;
assign _14171_ = _13523_ & _14174_ /*21613*/;
assign _14172_ = _13523_ ^ _14174_ /*21616*/;
assign _14173_ = _14165_ & _14172_ /*21614*/;
assign _14170_ = _14171_ | _14173_ /*21612*/;
assign _13909_ = _14165_ ^ _14172_ /*21615*/;
assign _14179_ = D[50] ^ Q[28] /*21611*/;
assign _14176_ = _13524_ & _14179_ /*21607*/;
assign _14177_ = _13524_ ^ _14179_ /*21610*/;
assign _14178_ = _14170_ & _14177_ /*21608*/;
assign _14175_ = _14176_ | _14178_ /*21606*/;
assign _13910_ = _14170_ ^ _14177_ /*21609*/;
assign _14184_ = D[51] ^ Q[28] /*21605*/;
assign _14181_ = _13525_ & _14184_ /*21601*/;
assign _14182_ = _13525_ ^ _14184_ /*21604*/;
assign _14183_ = _14175_ & _14182_ /*21602*/;
assign _14180_ = _14181_ | _14183_ /*21600*/;
assign _13911_ = _14175_ ^ _14182_ /*21603*/;
assign _14189_ = D[52] ^ Q[28] /*21599*/;
assign _14186_ = _13526_ & _14189_ /*21595*/;
assign _14187_ = _13526_ ^ _14189_ /*21598*/;
assign _14188_ = _14180_ & _14187_ /*21596*/;
assign _14185_ = _14186_ | _14188_ /*21594*/;
assign _13912_ = _14180_ ^ _14187_ /*21597*/;
assign _14194_ = D[53] ^ Q[28] /*21593*/;
assign _14191_ = _13527_ & _14194_ /*21589*/;
assign _14192_ = _13527_ ^ _14194_ /*21592*/;
assign _14193_ = _14185_ & _14192_ /*21590*/;
assign _14190_ = _14191_ | _14193_ /*21588*/;
assign _13913_ = _14185_ ^ _14192_ /*21591*/;
assign _14199_ = D[54] ^ Q[28] /*21587*/;
assign _14196_ = _13528_ & _14199_ /*21583*/;
assign _14197_ = _13528_ ^ _14199_ /*21586*/;
assign _14198_ = _14190_ & _14197_ /*21584*/;
assign _14195_ = _14196_ | _14198_ /*21582*/;
assign _13914_ = _14190_ ^ _14197_ /*21585*/;
assign _14204_ = D[55] ^ Q[28] /*21581*/;
assign _14201_ = _13529_ & _14204_ /*21577*/;
assign _14202_ = _13529_ ^ _14204_ /*21580*/;
assign _14203_ = _14195_ & _14202_ /*21578*/;
assign _14200_ = _14201_ | _14203_ /*21576*/;
assign _13915_ = _14195_ ^ _14202_ /*21579*/;
assign _14209_ = D[56] ^ Q[28] /*21575*/;
assign _14206_ = _13530_ & _14209_ /*21571*/;
assign _14207_ = _13530_ ^ _14209_ /*21574*/;
assign _14208_ = _14200_ & _14207_ /*21572*/;
assign _14205_ = _14206_ | _14208_ /*21570*/;
assign _13916_ = _14200_ ^ _14207_ /*21573*/;
assign _14214_ = D[57] ^ Q[28] /*21569*/;
assign _14211_ = _13531_ & _14214_ /*21565*/;
assign _14212_ = _13531_ ^ _14214_ /*21568*/;
assign _14213_ = _14205_ & _14212_ /*21566*/;
assign _14210_ = _14211_ | _14213_ /*21564*/;
assign _13917_ = _14205_ ^ _14212_ /*21567*/;
assign _14219_ = D[58] ^ Q[28] /*21563*/;
assign _14216_ = _13532_ & _14219_ /*21559*/;
assign _14217_ = _13532_ ^ _14219_ /*21562*/;
assign _14218_ = _14210_ & _14217_ /*21560*/;
assign _14215_ = _14216_ | _14218_ /*21558*/;
assign _13918_ = _14210_ ^ _14217_ /*21561*/;
assign _14224_ = D[59] ^ Q[28] /*21557*/;
assign _14221_ = _13533_ & _14224_ /*21553*/;
assign _14222_ = _13533_ ^ _14224_ /*21556*/;
assign _14223_ = _14215_ & _14222_ /*21554*/;
assign _14220_ = _14221_ | _14223_ /*21552*/;
assign _13919_ = _14215_ ^ _14222_ /*21555*/;
assign _14229_ = D[60] ^ Q[28] /*21551*/;
assign _14226_ = _13534_ & _14229_ /*21547*/;
assign _14227_ = _13534_ ^ _14229_ /*21550*/;
assign _14228_ = _14220_ & _14227_ /*21548*/;
assign _14225_ = _14226_ | _14228_ /*21546*/;
assign _13920_ = _14220_ ^ _14227_ /*21549*/;
assign _14234_ = D[61] ^ Q[28] /*21545*/;
assign _14231_ = _13535_ & _14234_ /*21541*/;
assign _14232_ = _13535_ ^ _14234_ /*21544*/;
assign _14233_ = _14225_ & _14232_ /*21542*/;
assign _14230_ = _14231_ | _14233_ /*21540*/;
assign _13921_ = _14225_ ^ _14232_ /*21543*/;
assign _14239_ = D[62] ^ Q[28] /*21539*/;
assign _14236_ = _13536_ & _14239_ /*21535*/;
assign _14237_ = _13536_ ^ _14239_ /*21538*/;
assign _14238_ = _14230_ & _14237_ /*21536*/;
assign _14235_ = _14236_ | _14238_ /*21534*/;
assign _13922_ = _14230_ ^ _14237_ /*21537*/;
assign _14243_ = zeroWire ^ Q[28] /*21533*/;
assign _14240_ = _13537_ & _14243_ /*21529*/;
assign _14241_ = _13537_ ^ _14243_ /*21532*/;
assign _14242_ = _14235_ & _14241_ /*21530*/;
assign Q[27] = _14240_ | _14242_ /*21528*/;
assign _13923_ = _14235_ ^ _14241_ /*21531*/;
assign _14314_ = D[0] ^ Q[27] /*21142*/;
assign _14311_ = R_0[26] & _14314_ /*21138*/;
assign _14312_ = R_0[26] ^ _14314_ /*21141*/;
assign _14313_ = Q[27] & _14312_ /*21139*/;
assign _14310_ = _14311_ | _14313_ /*21137*/;
assign _14245_ = Q[27] ^ _14312_ /*21140*/;
assign _14319_ = D[1] ^ Q[27] /*21136*/;
assign _14316_ = _13860_ & _14319_ /*21132*/;
assign _14317_ = _13860_ ^ _14319_ /*21135*/;
assign _14318_ = _14310_ & _14317_ /*21133*/;
assign _14315_ = _14316_ | _14318_ /*21131*/;
assign _14246_ = _14310_ ^ _14317_ /*21134*/;
assign _14324_ = D[2] ^ Q[27] /*21130*/;
assign _14321_ = _13861_ & _14324_ /*21126*/;
assign _14322_ = _13861_ ^ _14324_ /*21129*/;
assign _14323_ = _14315_ & _14322_ /*21127*/;
assign _14320_ = _14321_ | _14323_ /*21125*/;
assign _14247_ = _14315_ ^ _14322_ /*21128*/;
assign _14329_ = D[3] ^ Q[27] /*21124*/;
assign _14326_ = _13862_ & _14329_ /*21120*/;
assign _14327_ = _13862_ ^ _14329_ /*21123*/;
assign _14328_ = _14320_ & _14327_ /*21121*/;
assign _14325_ = _14326_ | _14328_ /*21119*/;
assign _14248_ = _14320_ ^ _14327_ /*21122*/;
assign _14334_ = D[4] ^ Q[27] /*21118*/;
assign _14331_ = _13863_ & _14334_ /*21114*/;
assign _14332_ = _13863_ ^ _14334_ /*21117*/;
assign _14333_ = _14325_ & _14332_ /*21115*/;
assign _14330_ = _14331_ | _14333_ /*21113*/;
assign _14249_ = _14325_ ^ _14332_ /*21116*/;
assign _14339_ = D[5] ^ Q[27] /*21112*/;
assign _14336_ = _13864_ & _14339_ /*21108*/;
assign _14337_ = _13864_ ^ _14339_ /*21111*/;
assign _14338_ = _14330_ & _14337_ /*21109*/;
assign _14335_ = _14336_ | _14338_ /*21107*/;
assign _14250_ = _14330_ ^ _14337_ /*21110*/;
assign _14344_ = D[6] ^ Q[27] /*21106*/;
assign _14341_ = _13865_ & _14344_ /*21102*/;
assign _14342_ = _13865_ ^ _14344_ /*21105*/;
assign _14343_ = _14335_ & _14342_ /*21103*/;
assign _14340_ = _14341_ | _14343_ /*21101*/;
assign _14251_ = _14335_ ^ _14342_ /*21104*/;
assign _14349_ = D[7] ^ Q[27] /*21100*/;
assign _14346_ = _13866_ & _14349_ /*21096*/;
assign _14347_ = _13866_ ^ _14349_ /*21099*/;
assign _14348_ = _14340_ & _14347_ /*21097*/;
assign _14345_ = _14346_ | _14348_ /*21095*/;
assign _14252_ = _14340_ ^ _14347_ /*21098*/;
assign _14354_ = D[8] ^ Q[27] /*21094*/;
assign _14351_ = _13867_ & _14354_ /*21090*/;
assign _14352_ = _13867_ ^ _14354_ /*21093*/;
assign _14353_ = _14345_ & _14352_ /*21091*/;
assign _14350_ = _14351_ | _14353_ /*21089*/;
assign _14253_ = _14345_ ^ _14352_ /*21092*/;
assign _14359_ = D[9] ^ Q[27] /*21088*/;
assign _14356_ = _13868_ & _14359_ /*21084*/;
assign _14357_ = _13868_ ^ _14359_ /*21087*/;
assign _14358_ = _14350_ & _14357_ /*21085*/;
assign _14355_ = _14356_ | _14358_ /*21083*/;
assign _14254_ = _14350_ ^ _14357_ /*21086*/;
assign _14364_ = D[10] ^ Q[27] /*21082*/;
assign _14361_ = _13869_ & _14364_ /*21078*/;
assign _14362_ = _13869_ ^ _14364_ /*21081*/;
assign _14363_ = _14355_ & _14362_ /*21079*/;
assign _14360_ = _14361_ | _14363_ /*21077*/;
assign _14255_ = _14355_ ^ _14362_ /*21080*/;
assign _14369_ = D[11] ^ Q[27] /*21076*/;
assign _14366_ = _13870_ & _14369_ /*21072*/;
assign _14367_ = _13870_ ^ _14369_ /*21075*/;
assign _14368_ = _14360_ & _14367_ /*21073*/;
assign _14365_ = _14366_ | _14368_ /*21071*/;
assign _14256_ = _14360_ ^ _14367_ /*21074*/;
assign _14374_ = D[12] ^ Q[27] /*21070*/;
assign _14371_ = _13871_ & _14374_ /*21066*/;
assign _14372_ = _13871_ ^ _14374_ /*21069*/;
assign _14373_ = _14365_ & _14372_ /*21067*/;
assign _14370_ = _14371_ | _14373_ /*21065*/;
assign _14257_ = _14365_ ^ _14372_ /*21068*/;
assign _14379_ = D[13] ^ Q[27] /*21064*/;
assign _14376_ = _13872_ & _14379_ /*21060*/;
assign _14377_ = _13872_ ^ _14379_ /*21063*/;
assign _14378_ = _14370_ & _14377_ /*21061*/;
assign _14375_ = _14376_ | _14378_ /*21059*/;
assign _14258_ = _14370_ ^ _14377_ /*21062*/;
assign _14384_ = D[14] ^ Q[27] /*21058*/;
assign _14381_ = _13873_ & _14384_ /*21054*/;
assign _14382_ = _13873_ ^ _14384_ /*21057*/;
assign _14383_ = _14375_ & _14382_ /*21055*/;
assign _14380_ = _14381_ | _14383_ /*21053*/;
assign _14259_ = _14375_ ^ _14382_ /*21056*/;
assign _14389_ = D[15] ^ Q[27] /*21052*/;
assign _14386_ = _13874_ & _14389_ /*21048*/;
assign _14387_ = _13874_ ^ _14389_ /*21051*/;
assign _14388_ = _14380_ & _14387_ /*21049*/;
assign _14385_ = _14386_ | _14388_ /*21047*/;
assign _14260_ = _14380_ ^ _14387_ /*21050*/;
assign _14394_ = D[16] ^ Q[27] /*21046*/;
assign _14391_ = _13875_ & _14394_ /*21042*/;
assign _14392_ = _13875_ ^ _14394_ /*21045*/;
assign _14393_ = _14385_ & _14392_ /*21043*/;
assign _14390_ = _14391_ | _14393_ /*21041*/;
assign _14261_ = _14385_ ^ _14392_ /*21044*/;
assign _14399_ = D[17] ^ Q[27] /*21040*/;
assign _14396_ = _13876_ & _14399_ /*21036*/;
assign _14397_ = _13876_ ^ _14399_ /*21039*/;
assign _14398_ = _14390_ & _14397_ /*21037*/;
assign _14395_ = _14396_ | _14398_ /*21035*/;
assign _14262_ = _14390_ ^ _14397_ /*21038*/;
assign _14404_ = D[18] ^ Q[27] /*21034*/;
assign _14401_ = _13877_ & _14404_ /*21030*/;
assign _14402_ = _13877_ ^ _14404_ /*21033*/;
assign _14403_ = _14395_ & _14402_ /*21031*/;
assign _14400_ = _14401_ | _14403_ /*21029*/;
assign _14263_ = _14395_ ^ _14402_ /*21032*/;
assign _14409_ = D[19] ^ Q[27] /*21028*/;
assign _14406_ = _13878_ & _14409_ /*21024*/;
assign _14407_ = _13878_ ^ _14409_ /*21027*/;
assign _14408_ = _14400_ & _14407_ /*21025*/;
assign _14405_ = _14406_ | _14408_ /*21023*/;
assign _14264_ = _14400_ ^ _14407_ /*21026*/;
assign _14414_ = D[20] ^ Q[27] /*21022*/;
assign _14411_ = _13879_ & _14414_ /*21018*/;
assign _14412_ = _13879_ ^ _14414_ /*21021*/;
assign _14413_ = _14405_ & _14412_ /*21019*/;
assign _14410_ = _14411_ | _14413_ /*21017*/;
assign _14265_ = _14405_ ^ _14412_ /*21020*/;
assign _14419_ = D[21] ^ Q[27] /*21016*/;
assign _14416_ = _13880_ & _14419_ /*21012*/;
assign _14417_ = _13880_ ^ _14419_ /*21015*/;
assign _14418_ = _14410_ & _14417_ /*21013*/;
assign _14415_ = _14416_ | _14418_ /*21011*/;
assign _14266_ = _14410_ ^ _14417_ /*21014*/;
assign _14424_ = D[22] ^ Q[27] /*21010*/;
assign _14421_ = _13881_ & _14424_ /*21006*/;
assign _14422_ = _13881_ ^ _14424_ /*21009*/;
assign _14423_ = _14415_ & _14422_ /*21007*/;
assign _14420_ = _14421_ | _14423_ /*21005*/;
assign _14267_ = _14415_ ^ _14422_ /*21008*/;
assign _14429_ = D[23] ^ Q[27] /*21004*/;
assign _14426_ = _13882_ & _14429_ /*21000*/;
assign _14427_ = _13882_ ^ _14429_ /*21003*/;
assign _14428_ = _14420_ & _14427_ /*21001*/;
assign _14425_ = _14426_ | _14428_ /*20999*/;
assign _14268_ = _14420_ ^ _14427_ /*21002*/;
assign _14434_ = D[24] ^ Q[27] /*20998*/;
assign _14431_ = _13883_ & _14434_ /*20994*/;
assign _14432_ = _13883_ ^ _14434_ /*20997*/;
assign _14433_ = _14425_ & _14432_ /*20995*/;
assign _14430_ = _14431_ | _14433_ /*20993*/;
assign _14269_ = _14425_ ^ _14432_ /*20996*/;
assign _14439_ = D[25] ^ Q[27] /*20992*/;
assign _14436_ = _13884_ & _14439_ /*20988*/;
assign _14437_ = _13884_ ^ _14439_ /*20991*/;
assign _14438_ = _14430_ & _14437_ /*20989*/;
assign _14435_ = _14436_ | _14438_ /*20987*/;
assign _14270_ = _14430_ ^ _14437_ /*20990*/;
assign _14444_ = D[26] ^ Q[27] /*20986*/;
assign _14441_ = _13885_ & _14444_ /*20982*/;
assign _14442_ = _13885_ ^ _14444_ /*20985*/;
assign _14443_ = _14435_ & _14442_ /*20983*/;
assign _14440_ = _14441_ | _14443_ /*20981*/;
assign _14271_ = _14435_ ^ _14442_ /*20984*/;
assign _14449_ = D[27] ^ Q[27] /*20980*/;
assign _14446_ = _13886_ & _14449_ /*20976*/;
assign _14447_ = _13886_ ^ _14449_ /*20979*/;
assign _14448_ = _14440_ & _14447_ /*20977*/;
assign _14445_ = _14446_ | _14448_ /*20975*/;
assign _14272_ = _14440_ ^ _14447_ /*20978*/;
assign _14454_ = D[28] ^ Q[27] /*20974*/;
assign _14451_ = _13887_ & _14454_ /*20970*/;
assign _14452_ = _13887_ ^ _14454_ /*20973*/;
assign _14453_ = _14445_ & _14452_ /*20971*/;
assign _14450_ = _14451_ | _14453_ /*20969*/;
assign _14273_ = _14445_ ^ _14452_ /*20972*/;
assign _14459_ = D[29] ^ Q[27] /*20968*/;
assign _14456_ = _13888_ & _14459_ /*20964*/;
assign _14457_ = _13888_ ^ _14459_ /*20967*/;
assign _14458_ = _14450_ & _14457_ /*20965*/;
assign _14455_ = _14456_ | _14458_ /*20963*/;
assign _14274_ = _14450_ ^ _14457_ /*20966*/;
assign _14464_ = D[30] ^ Q[27] /*20962*/;
assign _14461_ = _13889_ & _14464_ /*20958*/;
assign _14462_ = _13889_ ^ _14464_ /*20961*/;
assign _14463_ = _14455_ & _14462_ /*20959*/;
assign _14460_ = _14461_ | _14463_ /*20957*/;
assign _14275_ = _14455_ ^ _14462_ /*20960*/;
assign _14469_ = D[31] ^ Q[27] /*20956*/;
assign _14466_ = _13890_ & _14469_ /*20952*/;
assign _14467_ = _13890_ ^ _14469_ /*20955*/;
assign _14468_ = _14460_ & _14467_ /*20953*/;
assign _14465_ = _14466_ | _14468_ /*20951*/;
assign _14276_ = _14460_ ^ _14467_ /*20954*/;
assign _14474_ = D[32] ^ Q[27] /*20950*/;
assign _14471_ = _13891_ & _14474_ /*20946*/;
assign _14472_ = _13891_ ^ _14474_ /*20949*/;
assign _14473_ = _14465_ & _14472_ /*20947*/;
assign _14470_ = _14471_ | _14473_ /*20945*/;
assign _14277_ = _14465_ ^ _14472_ /*20948*/;
assign _14479_ = D[33] ^ Q[27] /*20944*/;
assign _14476_ = _13892_ & _14479_ /*20940*/;
assign _14477_ = _13892_ ^ _14479_ /*20943*/;
assign _14478_ = _14470_ & _14477_ /*20941*/;
assign _14475_ = _14476_ | _14478_ /*20939*/;
assign _14278_ = _14470_ ^ _14477_ /*20942*/;
assign _14484_ = D[34] ^ Q[27] /*20938*/;
assign _14481_ = _13893_ & _14484_ /*20934*/;
assign _14482_ = _13893_ ^ _14484_ /*20937*/;
assign _14483_ = _14475_ & _14482_ /*20935*/;
assign _14480_ = _14481_ | _14483_ /*20933*/;
assign _14279_ = _14475_ ^ _14482_ /*20936*/;
assign _14489_ = D[35] ^ Q[27] /*20932*/;
assign _14486_ = _13894_ & _14489_ /*20928*/;
assign _14487_ = _13894_ ^ _14489_ /*20931*/;
assign _14488_ = _14480_ & _14487_ /*20929*/;
assign _14485_ = _14486_ | _14488_ /*20927*/;
assign _14280_ = _14480_ ^ _14487_ /*20930*/;
assign _14494_ = D[36] ^ Q[27] /*20926*/;
assign _14491_ = _13895_ & _14494_ /*20922*/;
assign _14492_ = _13895_ ^ _14494_ /*20925*/;
assign _14493_ = _14485_ & _14492_ /*20923*/;
assign _14490_ = _14491_ | _14493_ /*20921*/;
assign _14281_ = _14485_ ^ _14492_ /*20924*/;
assign _14499_ = D[37] ^ Q[27] /*20920*/;
assign _14496_ = _13896_ & _14499_ /*20916*/;
assign _14497_ = _13896_ ^ _14499_ /*20919*/;
assign _14498_ = _14490_ & _14497_ /*20917*/;
assign _14495_ = _14496_ | _14498_ /*20915*/;
assign _14282_ = _14490_ ^ _14497_ /*20918*/;
assign _14504_ = D[38] ^ Q[27] /*20914*/;
assign _14501_ = _13897_ & _14504_ /*20910*/;
assign _14502_ = _13897_ ^ _14504_ /*20913*/;
assign _14503_ = _14495_ & _14502_ /*20911*/;
assign _14500_ = _14501_ | _14503_ /*20909*/;
assign _14283_ = _14495_ ^ _14502_ /*20912*/;
assign _14509_ = D[39] ^ Q[27] /*20908*/;
assign _14506_ = _13898_ & _14509_ /*20904*/;
assign _14507_ = _13898_ ^ _14509_ /*20907*/;
assign _14508_ = _14500_ & _14507_ /*20905*/;
assign _14505_ = _14506_ | _14508_ /*20903*/;
assign _14284_ = _14500_ ^ _14507_ /*20906*/;
assign _14514_ = D[40] ^ Q[27] /*20902*/;
assign _14511_ = _13899_ & _14514_ /*20898*/;
assign _14512_ = _13899_ ^ _14514_ /*20901*/;
assign _14513_ = _14505_ & _14512_ /*20899*/;
assign _14510_ = _14511_ | _14513_ /*20897*/;
assign _14285_ = _14505_ ^ _14512_ /*20900*/;
assign _14519_ = D[41] ^ Q[27] /*20896*/;
assign _14516_ = _13900_ & _14519_ /*20892*/;
assign _14517_ = _13900_ ^ _14519_ /*20895*/;
assign _14518_ = _14510_ & _14517_ /*20893*/;
assign _14515_ = _14516_ | _14518_ /*20891*/;
assign _14286_ = _14510_ ^ _14517_ /*20894*/;
assign _14524_ = D[42] ^ Q[27] /*20890*/;
assign _14521_ = _13901_ & _14524_ /*20886*/;
assign _14522_ = _13901_ ^ _14524_ /*20889*/;
assign _14523_ = _14515_ & _14522_ /*20887*/;
assign _14520_ = _14521_ | _14523_ /*20885*/;
assign _14287_ = _14515_ ^ _14522_ /*20888*/;
assign _14529_ = D[43] ^ Q[27] /*20884*/;
assign _14526_ = _13902_ & _14529_ /*20880*/;
assign _14527_ = _13902_ ^ _14529_ /*20883*/;
assign _14528_ = _14520_ & _14527_ /*20881*/;
assign _14525_ = _14526_ | _14528_ /*20879*/;
assign _14288_ = _14520_ ^ _14527_ /*20882*/;
assign _14534_ = D[44] ^ Q[27] /*20878*/;
assign _14531_ = _13903_ & _14534_ /*20874*/;
assign _14532_ = _13903_ ^ _14534_ /*20877*/;
assign _14533_ = _14525_ & _14532_ /*20875*/;
assign _14530_ = _14531_ | _14533_ /*20873*/;
assign _14289_ = _14525_ ^ _14532_ /*20876*/;
assign _14539_ = D[45] ^ Q[27] /*20872*/;
assign _14536_ = _13904_ & _14539_ /*20868*/;
assign _14537_ = _13904_ ^ _14539_ /*20871*/;
assign _14538_ = _14530_ & _14537_ /*20869*/;
assign _14535_ = _14536_ | _14538_ /*20867*/;
assign _14290_ = _14530_ ^ _14537_ /*20870*/;
assign _14544_ = D[46] ^ Q[27] /*20866*/;
assign _14541_ = _13905_ & _14544_ /*20862*/;
assign _14542_ = _13905_ ^ _14544_ /*20865*/;
assign _14543_ = _14535_ & _14542_ /*20863*/;
assign _14540_ = _14541_ | _14543_ /*20861*/;
assign _14291_ = _14535_ ^ _14542_ /*20864*/;
assign _14549_ = D[47] ^ Q[27] /*20860*/;
assign _14546_ = _13906_ & _14549_ /*20856*/;
assign _14547_ = _13906_ ^ _14549_ /*20859*/;
assign _14548_ = _14540_ & _14547_ /*20857*/;
assign _14545_ = _14546_ | _14548_ /*20855*/;
assign _14292_ = _14540_ ^ _14547_ /*20858*/;
assign _14554_ = D[48] ^ Q[27] /*20854*/;
assign _14551_ = _13907_ & _14554_ /*20850*/;
assign _14552_ = _13907_ ^ _14554_ /*20853*/;
assign _14553_ = _14545_ & _14552_ /*20851*/;
assign _14550_ = _14551_ | _14553_ /*20849*/;
assign _14293_ = _14545_ ^ _14552_ /*20852*/;
assign _14559_ = D[49] ^ Q[27] /*20848*/;
assign _14556_ = _13908_ & _14559_ /*20844*/;
assign _14557_ = _13908_ ^ _14559_ /*20847*/;
assign _14558_ = _14550_ & _14557_ /*20845*/;
assign _14555_ = _14556_ | _14558_ /*20843*/;
assign _14294_ = _14550_ ^ _14557_ /*20846*/;
assign _14564_ = D[50] ^ Q[27] /*20842*/;
assign _14561_ = _13909_ & _14564_ /*20838*/;
assign _14562_ = _13909_ ^ _14564_ /*20841*/;
assign _14563_ = _14555_ & _14562_ /*20839*/;
assign _14560_ = _14561_ | _14563_ /*20837*/;
assign _14295_ = _14555_ ^ _14562_ /*20840*/;
assign _14569_ = D[51] ^ Q[27] /*20836*/;
assign _14566_ = _13910_ & _14569_ /*20832*/;
assign _14567_ = _13910_ ^ _14569_ /*20835*/;
assign _14568_ = _14560_ & _14567_ /*20833*/;
assign _14565_ = _14566_ | _14568_ /*20831*/;
assign _14296_ = _14560_ ^ _14567_ /*20834*/;
assign _14574_ = D[52] ^ Q[27] /*20830*/;
assign _14571_ = _13911_ & _14574_ /*20826*/;
assign _14572_ = _13911_ ^ _14574_ /*20829*/;
assign _14573_ = _14565_ & _14572_ /*20827*/;
assign _14570_ = _14571_ | _14573_ /*20825*/;
assign _14297_ = _14565_ ^ _14572_ /*20828*/;
assign _14579_ = D[53] ^ Q[27] /*20824*/;
assign _14576_ = _13912_ & _14579_ /*20820*/;
assign _14577_ = _13912_ ^ _14579_ /*20823*/;
assign _14578_ = _14570_ & _14577_ /*20821*/;
assign _14575_ = _14576_ | _14578_ /*20819*/;
assign _14298_ = _14570_ ^ _14577_ /*20822*/;
assign _14584_ = D[54] ^ Q[27] /*20818*/;
assign _14581_ = _13913_ & _14584_ /*20814*/;
assign _14582_ = _13913_ ^ _14584_ /*20817*/;
assign _14583_ = _14575_ & _14582_ /*20815*/;
assign _14580_ = _14581_ | _14583_ /*20813*/;
assign _14299_ = _14575_ ^ _14582_ /*20816*/;
assign _14589_ = D[55] ^ Q[27] /*20812*/;
assign _14586_ = _13914_ & _14589_ /*20808*/;
assign _14587_ = _13914_ ^ _14589_ /*20811*/;
assign _14588_ = _14580_ & _14587_ /*20809*/;
assign _14585_ = _14586_ | _14588_ /*20807*/;
assign _14300_ = _14580_ ^ _14587_ /*20810*/;
assign _14594_ = D[56] ^ Q[27] /*20806*/;
assign _14591_ = _13915_ & _14594_ /*20802*/;
assign _14592_ = _13915_ ^ _14594_ /*20805*/;
assign _14593_ = _14585_ & _14592_ /*20803*/;
assign _14590_ = _14591_ | _14593_ /*20801*/;
assign _14301_ = _14585_ ^ _14592_ /*20804*/;
assign _14599_ = D[57] ^ Q[27] /*20800*/;
assign _14596_ = _13916_ & _14599_ /*20796*/;
assign _14597_ = _13916_ ^ _14599_ /*20799*/;
assign _14598_ = _14590_ & _14597_ /*20797*/;
assign _14595_ = _14596_ | _14598_ /*20795*/;
assign _14302_ = _14590_ ^ _14597_ /*20798*/;
assign _14604_ = D[58] ^ Q[27] /*20794*/;
assign _14601_ = _13917_ & _14604_ /*20790*/;
assign _14602_ = _13917_ ^ _14604_ /*20793*/;
assign _14603_ = _14595_ & _14602_ /*20791*/;
assign _14600_ = _14601_ | _14603_ /*20789*/;
assign _14303_ = _14595_ ^ _14602_ /*20792*/;
assign _14609_ = D[59] ^ Q[27] /*20788*/;
assign _14606_ = _13918_ & _14609_ /*20784*/;
assign _14607_ = _13918_ ^ _14609_ /*20787*/;
assign _14608_ = _14600_ & _14607_ /*20785*/;
assign _14605_ = _14606_ | _14608_ /*20783*/;
assign _14304_ = _14600_ ^ _14607_ /*20786*/;
assign _14614_ = D[60] ^ Q[27] /*20782*/;
assign _14611_ = _13919_ & _14614_ /*20778*/;
assign _14612_ = _13919_ ^ _14614_ /*20781*/;
assign _14613_ = _14605_ & _14612_ /*20779*/;
assign _14610_ = _14611_ | _14613_ /*20777*/;
assign _14305_ = _14605_ ^ _14612_ /*20780*/;
assign _14619_ = D[61] ^ Q[27] /*20776*/;
assign _14616_ = _13920_ & _14619_ /*20772*/;
assign _14617_ = _13920_ ^ _14619_ /*20775*/;
assign _14618_ = _14610_ & _14617_ /*20773*/;
assign _14615_ = _14616_ | _14618_ /*20771*/;
assign _14306_ = _14610_ ^ _14617_ /*20774*/;
assign _14624_ = D[62] ^ Q[27] /*20770*/;
assign _14621_ = _13921_ & _14624_ /*20766*/;
assign _14622_ = _13921_ ^ _14624_ /*20769*/;
assign _14623_ = _14615_ & _14622_ /*20767*/;
assign _14620_ = _14621_ | _14623_ /*20765*/;
assign _14307_ = _14615_ ^ _14622_ /*20768*/;
assign _14628_ = zeroWire ^ Q[27] /*20764*/;
assign _14625_ = _13922_ & _14628_ /*20760*/;
assign _14626_ = _13922_ ^ _14628_ /*20763*/;
assign _14627_ = _14620_ & _14626_ /*20761*/;
assign Q[26] = _14625_ | _14627_ /*20759*/;
assign _14308_ = _14620_ ^ _14626_ /*20762*/;
assign _14699_ = D[0] ^ Q[26] /*20373*/;
assign _14696_ = R_0[25] & _14699_ /*20369*/;
assign _14697_ = R_0[25] ^ _14699_ /*20372*/;
assign _14698_ = Q[26] & _14697_ /*20370*/;
assign _14695_ = _14696_ | _14698_ /*20368*/;
assign _14630_ = Q[26] ^ _14697_ /*20371*/;
assign _14704_ = D[1] ^ Q[26] /*20367*/;
assign _14701_ = _14245_ & _14704_ /*20363*/;
assign _14702_ = _14245_ ^ _14704_ /*20366*/;
assign _14703_ = _14695_ & _14702_ /*20364*/;
assign _14700_ = _14701_ | _14703_ /*20362*/;
assign _14631_ = _14695_ ^ _14702_ /*20365*/;
assign _14709_ = D[2] ^ Q[26] /*20361*/;
assign _14706_ = _14246_ & _14709_ /*20357*/;
assign _14707_ = _14246_ ^ _14709_ /*20360*/;
assign _14708_ = _14700_ & _14707_ /*20358*/;
assign _14705_ = _14706_ | _14708_ /*20356*/;
assign _14632_ = _14700_ ^ _14707_ /*20359*/;
assign _14714_ = D[3] ^ Q[26] /*20355*/;
assign _14711_ = _14247_ & _14714_ /*20351*/;
assign _14712_ = _14247_ ^ _14714_ /*20354*/;
assign _14713_ = _14705_ & _14712_ /*20352*/;
assign _14710_ = _14711_ | _14713_ /*20350*/;
assign _14633_ = _14705_ ^ _14712_ /*20353*/;
assign _14719_ = D[4] ^ Q[26] /*20349*/;
assign _14716_ = _14248_ & _14719_ /*20345*/;
assign _14717_ = _14248_ ^ _14719_ /*20348*/;
assign _14718_ = _14710_ & _14717_ /*20346*/;
assign _14715_ = _14716_ | _14718_ /*20344*/;
assign _14634_ = _14710_ ^ _14717_ /*20347*/;
assign _14724_ = D[5] ^ Q[26] /*20343*/;
assign _14721_ = _14249_ & _14724_ /*20339*/;
assign _14722_ = _14249_ ^ _14724_ /*20342*/;
assign _14723_ = _14715_ & _14722_ /*20340*/;
assign _14720_ = _14721_ | _14723_ /*20338*/;
assign _14635_ = _14715_ ^ _14722_ /*20341*/;
assign _14729_ = D[6] ^ Q[26] /*20337*/;
assign _14726_ = _14250_ & _14729_ /*20333*/;
assign _14727_ = _14250_ ^ _14729_ /*20336*/;
assign _14728_ = _14720_ & _14727_ /*20334*/;
assign _14725_ = _14726_ | _14728_ /*20332*/;
assign _14636_ = _14720_ ^ _14727_ /*20335*/;
assign _14734_ = D[7] ^ Q[26] /*20331*/;
assign _14731_ = _14251_ & _14734_ /*20327*/;
assign _14732_ = _14251_ ^ _14734_ /*20330*/;
assign _14733_ = _14725_ & _14732_ /*20328*/;
assign _14730_ = _14731_ | _14733_ /*20326*/;
assign _14637_ = _14725_ ^ _14732_ /*20329*/;
assign _14739_ = D[8] ^ Q[26] /*20325*/;
assign _14736_ = _14252_ & _14739_ /*20321*/;
assign _14737_ = _14252_ ^ _14739_ /*20324*/;
assign _14738_ = _14730_ & _14737_ /*20322*/;
assign _14735_ = _14736_ | _14738_ /*20320*/;
assign _14638_ = _14730_ ^ _14737_ /*20323*/;
assign _14744_ = D[9] ^ Q[26] /*20319*/;
assign _14741_ = _14253_ & _14744_ /*20315*/;
assign _14742_ = _14253_ ^ _14744_ /*20318*/;
assign _14743_ = _14735_ & _14742_ /*20316*/;
assign _14740_ = _14741_ | _14743_ /*20314*/;
assign _14639_ = _14735_ ^ _14742_ /*20317*/;
assign _14749_ = D[10] ^ Q[26] /*20313*/;
assign _14746_ = _14254_ & _14749_ /*20309*/;
assign _14747_ = _14254_ ^ _14749_ /*20312*/;
assign _14748_ = _14740_ & _14747_ /*20310*/;
assign _14745_ = _14746_ | _14748_ /*20308*/;
assign _14640_ = _14740_ ^ _14747_ /*20311*/;
assign _14754_ = D[11] ^ Q[26] /*20307*/;
assign _14751_ = _14255_ & _14754_ /*20303*/;
assign _14752_ = _14255_ ^ _14754_ /*20306*/;
assign _14753_ = _14745_ & _14752_ /*20304*/;
assign _14750_ = _14751_ | _14753_ /*20302*/;
assign _14641_ = _14745_ ^ _14752_ /*20305*/;
assign _14759_ = D[12] ^ Q[26] /*20301*/;
assign _14756_ = _14256_ & _14759_ /*20297*/;
assign _14757_ = _14256_ ^ _14759_ /*20300*/;
assign _14758_ = _14750_ & _14757_ /*20298*/;
assign _14755_ = _14756_ | _14758_ /*20296*/;
assign _14642_ = _14750_ ^ _14757_ /*20299*/;
assign _14764_ = D[13] ^ Q[26] /*20295*/;
assign _14761_ = _14257_ & _14764_ /*20291*/;
assign _14762_ = _14257_ ^ _14764_ /*20294*/;
assign _14763_ = _14755_ & _14762_ /*20292*/;
assign _14760_ = _14761_ | _14763_ /*20290*/;
assign _14643_ = _14755_ ^ _14762_ /*20293*/;
assign _14769_ = D[14] ^ Q[26] /*20289*/;
assign _14766_ = _14258_ & _14769_ /*20285*/;
assign _14767_ = _14258_ ^ _14769_ /*20288*/;
assign _14768_ = _14760_ & _14767_ /*20286*/;
assign _14765_ = _14766_ | _14768_ /*20284*/;
assign _14644_ = _14760_ ^ _14767_ /*20287*/;
assign _14774_ = D[15] ^ Q[26] /*20283*/;
assign _14771_ = _14259_ & _14774_ /*20279*/;
assign _14772_ = _14259_ ^ _14774_ /*20282*/;
assign _14773_ = _14765_ & _14772_ /*20280*/;
assign _14770_ = _14771_ | _14773_ /*20278*/;
assign _14645_ = _14765_ ^ _14772_ /*20281*/;
assign _14779_ = D[16] ^ Q[26] /*20277*/;
assign _14776_ = _14260_ & _14779_ /*20273*/;
assign _14777_ = _14260_ ^ _14779_ /*20276*/;
assign _14778_ = _14770_ & _14777_ /*20274*/;
assign _14775_ = _14776_ | _14778_ /*20272*/;
assign _14646_ = _14770_ ^ _14777_ /*20275*/;
assign _14784_ = D[17] ^ Q[26] /*20271*/;
assign _14781_ = _14261_ & _14784_ /*20267*/;
assign _14782_ = _14261_ ^ _14784_ /*20270*/;
assign _14783_ = _14775_ & _14782_ /*20268*/;
assign _14780_ = _14781_ | _14783_ /*20266*/;
assign _14647_ = _14775_ ^ _14782_ /*20269*/;
assign _14789_ = D[18] ^ Q[26] /*20265*/;
assign _14786_ = _14262_ & _14789_ /*20261*/;
assign _14787_ = _14262_ ^ _14789_ /*20264*/;
assign _14788_ = _14780_ & _14787_ /*20262*/;
assign _14785_ = _14786_ | _14788_ /*20260*/;
assign _14648_ = _14780_ ^ _14787_ /*20263*/;
assign _14794_ = D[19] ^ Q[26] /*20259*/;
assign _14791_ = _14263_ & _14794_ /*20255*/;
assign _14792_ = _14263_ ^ _14794_ /*20258*/;
assign _14793_ = _14785_ & _14792_ /*20256*/;
assign _14790_ = _14791_ | _14793_ /*20254*/;
assign _14649_ = _14785_ ^ _14792_ /*20257*/;
assign _14799_ = D[20] ^ Q[26] /*20253*/;
assign _14796_ = _14264_ & _14799_ /*20249*/;
assign _14797_ = _14264_ ^ _14799_ /*20252*/;
assign _14798_ = _14790_ & _14797_ /*20250*/;
assign _14795_ = _14796_ | _14798_ /*20248*/;
assign _14650_ = _14790_ ^ _14797_ /*20251*/;
assign _14804_ = D[21] ^ Q[26] /*20247*/;
assign _14801_ = _14265_ & _14804_ /*20243*/;
assign _14802_ = _14265_ ^ _14804_ /*20246*/;
assign _14803_ = _14795_ & _14802_ /*20244*/;
assign _14800_ = _14801_ | _14803_ /*20242*/;
assign _14651_ = _14795_ ^ _14802_ /*20245*/;
assign _14809_ = D[22] ^ Q[26] /*20241*/;
assign _14806_ = _14266_ & _14809_ /*20237*/;
assign _14807_ = _14266_ ^ _14809_ /*20240*/;
assign _14808_ = _14800_ & _14807_ /*20238*/;
assign _14805_ = _14806_ | _14808_ /*20236*/;
assign _14652_ = _14800_ ^ _14807_ /*20239*/;
assign _14814_ = D[23] ^ Q[26] /*20235*/;
assign _14811_ = _14267_ & _14814_ /*20231*/;
assign _14812_ = _14267_ ^ _14814_ /*20234*/;
assign _14813_ = _14805_ & _14812_ /*20232*/;
assign _14810_ = _14811_ | _14813_ /*20230*/;
assign _14653_ = _14805_ ^ _14812_ /*20233*/;
assign _14819_ = D[24] ^ Q[26] /*20229*/;
assign _14816_ = _14268_ & _14819_ /*20225*/;
assign _14817_ = _14268_ ^ _14819_ /*20228*/;
assign _14818_ = _14810_ & _14817_ /*20226*/;
assign _14815_ = _14816_ | _14818_ /*20224*/;
assign _14654_ = _14810_ ^ _14817_ /*20227*/;
assign _14824_ = D[25] ^ Q[26] /*20223*/;
assign _14821_ = _14269_ & _14824_ /*20219*/;
assign _14822_ = _14269_ ^ _14824_ /*20222*/;
assign _14823_ = _14815_ & _14822_ /*20220*/;
assign _14820_ = _14821_ | _14823_ /*20218*/;
assign _14655_ = _14815_ ^ _14822_ /*20221*/;
assign _14829_ = D[26] ^ Q[26] /*20217*/;
assign _14826_ = _14270_ & _14829_ /*20213*/;
assign _14827_ = _14270_ ^ _14829_ /*20216*/;
assign _14828_ = _14820_ & _14827_ /*20214*/;
assign _14825_ = _14826_ | _14828_ /*20212*/;
assign _14656_ = _14820_ ^ _14827_ /*20215*/;
assign _14834_ = D[27] ^ Q[26] /*20211*/;
assign _14831_ = _14271_ & _14834_ /*20207*/;
assign _14832_ = _14271_ ^ _14834_ /*20210*/;
assign _14833_ = _14825_ & _14832_ /*20208*/;
assign _14830_ = _14831_ | _14833_ /*20206*/;
assign _14657_ = _14825_ ^ _14832_ /*20209*/;
assign _14839_ = D[28] ^ Q[26] /*20205*/;
assign _14836_ = _14272_ & _14839_ /*20201*/;
assign _14837_ = _14272_ ^ _14839_ /*20204*/;
assign _14838_ = _14830_ & _14837_ /*20202*/;
assign _14835_ = _14836_ | _14838_ /*20200*/;
assign _14658_ = _14830_ ^ _14837_ /*20203*/;
assign _14844_ = D[29] ^ Q[26] /*20199*/;
assign _14841_ = _14273_ & _14844_ /*20195*/;
assign _14842_ = _14273_ ^ _14844_ /*20198*/;
assign _14843_ = _14835_ & _14842_ /*20196*/;
assign _14840_ = _14841_ | _14843_ /*20194*/;
assign _14659_ = _14835_ ^ _14842_ /*20197*/;
assign _14849_ = D[30] ^ Q[26] /*20193*/;
assign _14846_ = _14274_ & _14849_ /*20189*/;
assign _14847_ = _14274_ ^ _14849_ /*20192*/;
assign _14848_ = _14840_ & _14847_ /*20190*/;
assign _14845_ = _14846_ | _14848_ /*20188*/;
assign _14660_ = _14840_ ^ _14847_ /*20191*/;
assign _14854_ = D[31] ^ Q[26] /*20187*/;
assign _14851_ = _14275_ & _14854_ /*20183*/;
assign _14852_ = _14275_ ^ _14854_ /*20186*/;
assign _14853_ = _14845_ & _14852_ /*20184*/;
assign _14850_ = _14851_ | _14853_ /*20182*/;
assign _14661_ = _14845_ ^ _14852_ /*20185*/;
assign _14859_ = D[32] ^ Q[26] /*20181*/;
assign _14856_ = _14276_ & _14859_ /*20177*/;
assign _14857_ = _14276_ ^ _14859_ /*20180*/;
assign _14858_ = _14850_ & _14857_ /*20178*/;
assign _14855_ = _14856_ | _14858_ /*20176*/;
assign _14662_ = _14850_ ^ _14857_ /*20179*/;
assign _14864_ = D[33] ^ Q[26] /*20175*/;
assign _14861_ = _14277_ & _14864_ /*20171*/;
assign _14862_ = _14277_ ^ _14864_ /*20174*/;
assign _14863_ = _14855_ & _14862_ /*20172*/;
assign _14860_ = _14861_ | _14863_ /*20170*/;
assign _14663_ = _14855_ ^ _14862_ /*20173*/;
assign _14869_ = D[34] ^ Q[26] /*20169*/;
assign _14866_ = _14278_ & _14869_ /*20165*/;
assign _14867_ = _14278_ ^ _14869_ /*20168*/;
assign _14868_ = _14860_ & _14867_ /*20166*/;
assign _14865_ = _14866_ | _14868_ /*20164*/;
assign _14664_ = _14860_ ^ _14867_ /*20167*/;
assign _14874_ = D[35] ^ Q[26] /*20163*/;
assign _14871_ = _14279_ & _14874_ /*20159*/;
assign _14872_ = _14279_ ^ _14874_ /*20162*/;
assign _14873_ = _14865_ & _14872_ /*20160*/;
assign _14870_ = _14871_ | _14873_ /*20158*/;
assign _14665_ = _14865_ ^ _14872_ /*20161*/;
assign _14879_ = D[36] ^ Q[26] /*20157*/;
assign _14876_ = _14280_ & _14879_ /*20153*/;
assign _14877_ = _14280_ ^ _14879_ /*20156*/;
assign _14878_ = _14870_ & _14877_ /*20154*/;
assign _14875_ = _14876_ | _14878_ /*20152*/;
assign _14666_ = _14870_ ^ _14877_ /*20155*/;
assign _14884_ = D[37] ^ Q[26] /*20151*/;
assign _14881_ = _14281_ & _14884_ /*20147*/;
assign _14882_ = _14281_ ^ _14884_ /*20150*/;
assign _14883_ = _14875_ & _14882_ /*20148*/;
assign _14880_ = _14881_ | _14883_ /*20146*/;
assign _14667_ = _14875_ ^ _14882_ /*20149*/;
assign _14889_ = D[38] ^ Q[26] /*20145*/;
assign _14886_ = _14282_ & _14889_ /*20141*/;
assign _14887_ = _14282_ ^ _14889_ /*20144*/;
assign _14888_ = _14880_ & _14887_ /*20142*/;
assign _14885_ = _14886_ | _14888_ /*20140*/;
assign _14668_ = _14880_ ^ _14887_ /*20143*/;
assign _14894_ = D[39] ^ Q[26] /*20139*/;
assign _14891_ = _14283_ & _14894_ /*20135*/;
assign _14892_ = _14283_ ^ _14894_ /*20138*/;
assign _14893_ = _14885_ & _14892_ /*20136*/;
assign _14890_ = _14891_ | _14893_ /*20134*/;
assign _14669_ = _14885_ ^ _14892_ /*20137*/;
assign _14899_ = D[40] ^ Q[26] /*20133*/;
assign _14896_ = _14284_ & _14899_ /*20129*/;
assign _14897_ = _14284_ ^ _14899_ /*20132*/;
assign _14898_ = _14890_ & _14897_ /*20130*/;
assign _14895_ = _14896_ | _14898_ /*20128*/;
assign _14670_ = _14890_ ^ _14897_ /*20131*/;
assign _14904_ = D[41] ^ Q[26] /*20127*/;
assign _14901_ = _14285_ & _14904_ /*20123*/;
assign _14902_ = _14285_ ^ _14904_ /*20126*/;
assign _14903_ = _14895_ & _14902_ /*20124*/;
assign _14900_ = _14901_ | _14903_ /*20122*/;
assign _14671_ = _14895_ ^ _14902_ /*20125*/;
assign _14909_ = D[42] ^ Q[26] /*20121*/;
assign _14906_ = _14286_ & _14909_ /*20117*/;
assign _14907_ = _14286_ ^ _14909_ /*20120*/;
assign _14908_ = _14900_ & _14907_ /*20118*/;
assign _14905_ = _14906_ | _14908_ /*20116*/;
assign _14672_ = _14900_ ^ _14907_ /*20119*/;
assign _14914_ = D[43] ^ Q[26] /*20115*/;
assign _14911_ = _14287_ & _14914_ /*20111*/;
assign _14912_ = _14287_ ^ _14914_ /*20114*/;
assign _14913_ = _14905_ & _14912_ /*20112*/;
assign _14910_ = _14911_ | _14913_ /*20110*/;
assign _14673_ = _14905_ ^ _14912_ /*20113*/;
assign _14919_ = D[44] ^ Q[26] /*20109*/;
assign _14916_ = _14288_ & _14919_ /*20105*/;
assign _14917_ = _14288_ ^ _14919_ /*20108*/;
assign _14918_ = _14910_ & _14917_ /*20106*/;
assign _14915_ = _14916_ | _14918_ /*20104*/;
assign _14674_ = _14910_ ^ _14917_ /*20107*/;
assign _14924_ = D[45] ^ Q[26] /*20103*/;
assign _14921_ = _14289_ & _14924_ /*20099*/;
assign _14922_ = _14289_ ^ _14924_ /*20102*/;
assign _14923_ = _14915_ & _14922_ /*20100*/;
assign _14920_ = _14921_ | _14923_ /*20098*/;
assign _14675_ = _14915_ ^ _14922_ /*20101*/;
assign _14929_ = D[46] ^ Q[26] /*20097*/;
assign _14926_ = _14290_ & _14929_ /*20093*/;
assign _14927_ = _14290_ ^ _14929_ /*20096*/;
assign _14928_ = _14920_ & _14927_ /*20094*/;
assign _14925_ = _14926_ | _14928_ /*20092*/;
assign _14676_ = _14920_ ^ _14927_ /*20095*/;
assign _14934_ = D[47] ^ Q[26] /*20091*/;
assign _14931_ = _14291_ & _14934_ /*20087*/;
assign _14932_ = _14291_ ^ _14934_ /*20090*/;
assign _14933_ = _14925_ & _14932_ /*20088*/;
assign _14930_ = _14931_ | _14933_ /*20086*/;
assign _14677_ = _14925_ ^ _14932_ /*20089*/;
assign _14939_ = D[48] ^ Q[26] /*20085*/;
assign _14936_ = _14292_ & _14939_ /*20081*/;
assign _14937_ = _14292_ ^ _14939_ /*20084*/;
assign _14938_ = _14930_ & _14937_ /*20082*/;
assign _14935_ = _14936_ | _14938_ /*20080*/;
assign _14678_ = _14930_ ^ _14937_ /*20083*/;
assign _14944_ = D[49] ^ Q[26] /*20079*/;
assign _14941_ = _14293_ & _14944_ /*20075*/;
assign _14942_ = _14293_ ^ _14944_ /*20078*/;
assign _14943_ = _14935_ & _14942_ /*20076*/;
assign _14940_ = _14941_ | _14943_ /*20074*/;
assign _14679_ = _14935_ ^ _14942_ /*20077*/;
assign _14949_ = D[50] ^ Q[26] /*20073*/;
assign _14946_ = _14294_ & _14949_ /*20069*/;
assign _14947_ = _14294_ ^ _14949_ /*20072*/;
assign _14948_ = _14940_ & _14947_ /*20070*/;
assign _14945_ = _14946_ | _14948_ /*20068*/;
assign _14680_ = _14940_ ^ _14947_ /*20071*/;
assign _14954_ = D[51] ^ Q[26] /*20067*/;
assign _14951_ = _14295_ & _14954_ /*20063*/;
assign _14952_ = _14295_ ^ _14954_ /*20066*/;
assign _14953_ = _14945_ & _14952_ /*20064*/;
assign _14950_ = _14951_ | _14953_ /*20062*/;
assign _14681_ = _14945_ ^ _14952_ /*20065*/;
assign _14959_ = D[52] ^ Q[26] /*20061*/;
assign _14956_ = _14296_ & _14959_ /*20057*/;
assign _14957_ = _14296_ ^ _14959_ /*20060*/;
assign _14958_ = _14950_ & _14957_ /*20058*/;
assign _14955_ = _14956_ | _14958_ /*20056*/;
assign _14682_ = _14950_ ^ _14957_ /*20059*/;
assign _14964_ = D[53] ^ Q[26] /*20055*/;
assign _14961_ = _14297_ & _14964_ /*20051*/;
assign _14962_ = _14297_ ^ _14964_ /*20054*/;
assign _14963_ = _14955_ & _14962_ /*20052*/;
assign _14960_ = _14961_ | _14963_ /*20050*/;
assign _14683_ = _14955_ ^ _14962_ /*20053*/;
assign _14969_ = D[54] ^ Q[26] /*20049*/;
assign _14966_ = _14298_ & _14969_ /*20045*/;
assign _14967_ = _14298_ ^ _14969_ /*20048*/;
assign _14968_ = _14960_ & _14967_ /*20046*/;
assign _14965_ = _14966_ | _14968_ /*20044*/;
assign _14684_ = _14960_ ^ _14967_ /*20047*/;
assign _14974_ = D[55] ^ Q[26] /*20043*/;
assign _14971_ = _14299_ & _14974_ /*20039*/;
assign _14972_ = _14299_ ^ _14974_ /*20042*/;
assign _14973_ = _14965_ & _14972_ /*20040*/;
assign _14970_ = _14971_ | _14973_ /*20038*/;
assign _14685_ = _14965_ ^ _14972_ /*20041*/;
assign _14979_ = D[56] ^ Q[26] /*20037*/;
assign _14976_ = _14300_ & _14979_ /*20033*/;
assign _14977_ = _14300_ ^ _14979_ /*20036*/;
assign _14978_ = _14970_ & _14977_ /*20034*/;
assign _14975_ = _14976_ | _14978_ /*20032*/;
assign _14686_ = _14970_ ^ _14977_ /*20035*/;
assign _14984_ = D[57] ^ Q[26] /*20031*/;
assign _14981_ = _14301_ & _14984_ /*20027*/;
assign _14982_ = _14301_ ^ _14984_ /*20030*/;
assign _14983_ = _14975_ & _14982_ /*20028*/;
assign _14980_ = _14981_ | _14983_ /*20026*/;
assign _14687_ = _14975_ ^ _14982_ /*20029*/;
assign _14989_ = D[58] ^ Q[26] /*20025*/;
assign _14986_ = _14302_ & _14989_ /*20021*/;
assign _14987_ = _14302_ ^ _14989_ /*20024*/;
assign _14988_ = _14980_ & _14987_ /*20022*/;
assign _14985_ = _14986_ | _14988_ /*20020*/;
assign _14688_ = _14980_ ^ _14987_ /*20023*/;
assign _14994_ = D[59] ^ Q[26] /*20019*/;
assign _14991_ = _14303_ & _14994_ /*20015*/;
assign _14992_ = _14303_ ^ _14994_ /*20018*/;
assign _14993_ = _14985_ & _14992_ /*20016*/;
assign _14990_ = _14991_ | _14993_ /*20014*/;
assign _14689_ = _14985_ ^ _14992_ /*20017*/;
assign _14999_ = D[60] ^ Q[26] /*20013*/;
assign _14996_ = _14304_ & _14999_ /*20009*/;
assign _14997_ = _14304_ ^ _14999_ /*20012*/;
assign _14998_ = _14990_ & _14997_ /*20010*/;
assign _14995_ = _14996_ | _14998_ /*20008*/;
assign _14690_ = _14990_ ^ _14997_ /*20011*/;
assign _15004_ = D[61] ^ Q[26] /*20007*/;
assign _15001_ = _14305_ & _15004_ /*20003*/;
assign _15002_ = _14305_ ^ _15004_ /*20006*/;
assign _15003_ = _14995_ & _15002_ /*20004*/;
assign _15000_ = _15001_ | _15003_ /*20002*/;
assign _14691_ = _14995_ ^ _15002_ /*20005*/;
assign _15009_ = D[62] ^ Q[26] /*20001*/;
assign _15006_ = _14306_ & _15009_ /*19997*/;
assign _15007_ = _14306_ ^ _15009_ /*20000*/;
assign _15008_ = _15000_ & _15007_ /*19998*/;
assign _15005_ = _15006_ | _15008_ /*19996*/;
assign _14692_ = _15000_ ^ _15007_ /*19999*/;
assign _15013_ = zeroWire ^ Q[26] /*19995*/;
assign _15010_ = _14307_ & _15013_ /*19991*/;
assign _15011_ = _14307_ ^ _15013_ /*19994*/;
assign _15012_ = _15005_ & _15011_ /*19992*/;
assign Q[25] = _15010_ | _15012_ /*19990*/;
assign _14693_ = _15005_ ^ _15011_ /*19993*/;
assign _15084_ = D[0] ^ Q[25] /*19604*/;
assign _15081_ = R_0[24] & _15084_ /*19600*/;
assign _15082_ = R_0[24] ^ _15084_ /*19603*/;
assign _15083_ = Q[25] & _15082_ /*19601*/;
assign _15080_ = _15081_ | _15083_ /*19599*/;
assign _15015_ = Q[25] ^ _15082_ /*19602*/;
assign _15089_ = D[1] ^ Q[25] /*19598*/;
assign _15086_ = _14630_ & _15089_ /*19594*/;
assign _15087_ = _14630_ ^ _15089_ /*19597*/;
assign _15088_ = _15080_ & _15087_ /*19595*/;
assign _15085_ = _15086_ | _15088_ /*19593*/;
assign _15016_ = _15080_ ^ _15087_ /*19596*/;
assign _15094_ = D[2] ^ Q[25] /*19592*/;
assign _15091_ = _14631_ & _15094_ /*19588*/;
assign _15092_ = _14631_ ^ _15094_ /*19591*/;
assign _15093_ = _15085_ & _15092_ /*19589*/;
assign _15090_ = _15091_ | _15093_ /*19587*/;
assign _15017_ = _15085_ ^ _15092_ /*19590*/;
assign _15099_ = D[3] ^ Q[25] /*19586*/;
assign _15096_ = _14632_ & _15099_ /*19582*/;
assign _15097_ = _14632_ ^ _15099_ /*19585*/;
assign _15098_ = _15090_ & _15097_ /*19583*/;
assign _15095_ = _15096_ | _15098_ /*19581*/;
assign _15018_ = _15090_ ^ _15097_ /*19584*/;
assign _15104_ = D[4] ^ Q[25] /*19580*/;
assign _15101_ = _14633_ & _15104_ /*19576*/;
assign _15102_ = _14633_ ^ _15104_ /*19579*/;
assign _15103_ = _15095_ & _15102_ /*19577*/;
assign _15100_ = _15101_ | _15103_ /*19575*/;
assign _15019_ = _15095_ ^ _15102_ /*19578*/;
assign _15109_ = D[5] ^ Q[25] /*19574*/;
assign _15106_ = _14634_ & _15109_ /*19570*/;
assign _15107_ = _14634_ ^ _15109_ /*19573*/;
assign _15108_ = _15100_ & _15107_ /*19571*/;
assign _15105_ = _15106_ | _15108_ /*19569*/;
assign _15020_ = _15100_ ^ _15107_ /*19572*/;
assign _15114_ = D[6] ^ Q[25] /*19568*/;
assign _15111_ = _14635_ & _15114_ /*19564*/;
assign _15112_ = _14635_ ^ _15114_ /*19567*/;
assign _15113_ = _15105_ & _15112_ /*19565*/;
assign _15110_ = _15111_ | _15113_ /*19563*/;
assign _15021_ = _15105_ ^ _15112_ /*19566*/;
assign _15119_ = D[7] ^ Q[25] /*19562*/;
assign _15116_ = _14636_ & _15119_ /*19558*/;
assign _15117_ = _14636_ ^ _15119_ /*19561*/;
assign _15118_ = _15110_ & _15117_ /*19559*/;
assign _15115_ = _15116_ | _15118_ /*19557*/;
assign _15022_ = _15110_ ^ _15117_ /*19560*/;
assign _15124_ = D[8] ^ Q[25] /*19556*/;
assign _15121_ = _14637_ & _15124_ /*19552*/;
assign _15122_ = _14637_ ^ _15124_ /*19555*/;
assign _15123_ = _15115_ & _15122_ /*19553*/;
assign _15120_ = _15121_ | _15123_ /*19551*/;
assign _15023_ = _15115_ ^ _15122_ /*19554*/;
assign _15129_ = D[9] ^ Q[25] /*19550*/;
assign _15126_ = _14638_ & _15129_ /*19546*/;
assign _15127_ = _14638_ ^ _15129_ /*19549*/;
assign _15128_ = _15120_ & _15127_ /*19547*/;
assign _15125_ = _15126_ | _15128_ /*19545*/;
assign _15024_ = _15120_ ^ _15127_ /*19548*/;
assign _15134_ = D[10] ^ Q[25] /*19544*/;
assign _15131_ = _14639_ & _15134_ /*19540*/;
assign _15132_ = _14639_ ^ _15134_ /*19543*/;
assign _15133_ = _15125_ & _15132_ /*19541*/;
assign _15130_ = _15131_ | _15133_ /*19539*/;
assign _15025_ = _15125_ ^ _15132_ /*19542*/;
assign _15139_ = D[11] ^ Q[25] /*19538*/;
assign _15136_ = _14640_ & _15139_ /*19534*/;
assign _15137_ = _14640_ ^ _15139_ /*19537*/;
assign _15138_ = _15130_ & _15137_ /*19535*/;
assign _15135_ = _15136_ | _15138_ /*19533*/;
assign _15026_ = _15130_ ^ _15137_ /*19536*/;
assign _15144_ = D[12] ^ Q[25] /*19532*/;
assign _15141_ = _14641_ & _15144_ /*19528*/;
assign _15142_ = _14641_ ^ _15144_ /*19531*/;
assign _15143_ = _15135_ & _15142_ /*19529*/;
assign _15140_ = _15141_ | _15143_ /*19527*/;
assign _15027_ = _15135_ ^ _15142_ /*19530*/;
assign _15149_ = D[13] ^ Q[25] /*19526*/;
assign _15146_ = _14642_ & _15149_ /*19522*/;
assign _15147_ = _14642_ ^ _15149_ /*19525*/;
assign _15148_ = _15140_ & _15147_ /*19523*/;
assign _15145_ = _15146_ | _15148_ /*19521*/;
assign _15028_ = _15140_ ^ _15147_ /*19524*/;
assign _15154_ = D[14] ^ Q[25] /*19520*/;
assign _15151_ = _14643_ & _15154_ /*19516*/;
assign _15152_ = _14643_ ^ _15154_ /*19519*/;
assign _15153_ = _15145_ & _15152_ /*19517*/;
assign _15150_ = _15151_ | _15153_ /*19515*/;
assign _15029_ = _15145_ ^ _15152_ /*19518*/;
assign _15159_ = D[15] ^ Q[25] /*19514*/;
assign _15156_ = _14644_ & _15159_ /*19510*/;
assign _15157_ = _14644_ ^ _15159_ /*19513*/;
assign _15158_ = _15150_ & _15157_ /*19511*/;
assign _15155_ = _15156_ | _15158_ /*19509*/;
assign _15030_ = _15150_ ^ _15157_ /*19512*/;
assign _15164_ = D[16] ^ Q[25] /*19508*/;
assign _15161_ = _14645_ & _15164_ /*19504*/;
assign _15162_ = _14645_ ^ _15164_ /*19507*/;
assign _15163_ = _15155_ & _15162_ /*19505*/;
assign _15160_ = _15161_ | _15163_ /*19503*/;
assign _15031_ = _15155_ ^ _15162_ /*19506*/;
assign _15169_ = D[17] ^ Q[25] /*19502*/;
assign _15166_ = _14646_ & _15169_ /*19498*/;
assign _15167_ = _14646_ ^ _15169_ /*19501*/;
assign _15168_ = _15160_ & _15167_ /*19499*/;
assign _15165_ = _15166_ | _15168_ /*19497*/;
assign _15032_ = _15160_ ^ _15167_ /*19500*/;
assign _15174_ = D[18] ^ Q[25] /*19496*/;
assign _15171_ = _14647_ & _15174_ /*19492*/;
assign _15172_ = _14647_ ^ _15174_ /*19495*/;
assign _15173_ = _15165_ & _15172_ /*19493*/;
assign _15170_ = _15171_ | _15173_ /*19491*/;
assign _15033_ = _15165_ ^ _15172_ /*19494*/;
assign _15179_ = D[19] ^ Q[25] /*19490*/;
assign _15176_ = _14648_ & _15179_ /*19486*/;
assign _15177_ = _14648_ ^ _15179_ /*19489*/;
assign _15178_ = _15170_ & _15177_ /*19487*/;
assign _15175_ = _15176_ | _15178_ /*19485*/;
assign _15034_ = _15170_ ^ _15177_ /*19488*/;
assign _15184_ = D[20] ^ Q[25] /*19484*/;
assign _15181_ = _14649_ & _15184_ /*19480*/;
assign _15182_ = _14649_ ^ _15184_ /*19483*/;
assign _15183_ = _15175_ & _15182_ /*19481*/;
assign _15180_ = _15181_ | _15183_ /*19479*/;
assign _15035_ = _15175_ ^ _15182_ /*19482*/;
assign _15189_ = D[21] ^ Q[25] /*19478*/;
assign _15186_ = _14650_ & _15189_ /*19474*/;
assign _15187_ = _14650_ ^ _15189_ /*19477*/;
assign _15188_ = _15180_ & _15187_ /*19475*/;
assign _15185_ = _15186_ | _15188_ /*19473*/;
assign _15036_ = _15180_ ^ _15187_ /*19476*/;
assign _15194_ = D[22] ^ Q[25] /*19472*/;
assign _15191_ = _14651_ & _15194_ /*19468*/;
assign _15192_ = _14651_ ^ _15194_ /*19471*/;
assign _15193_ = _15185_ & _15192_ /*19469*/;
assign _15190_ = _15191_ | _15193_ /*19467*/;
assign _15037_ = _15185_ ^ _15192_ /*19470*/;
assign _15199_ = D[23] ^ Q[25] /*19466*/;
assign _15196_ = _14652_ & _15199_ /*19462*/;
assign _15197_ = _14652_ ^ _15199_ /*19465*/;
assign _15198_ = _15190_ & _15197_ /*19463*/;
assign _15195_ = _15196_ | _15198_ /*19461*/;
assign _15038_ = _15190_ ^ _15197_ /*19464*/;
assign _15204_ = D[24] ^ Q[25] /*19460*/;
assign _15201_ = _14653_ & _15204_ /*19456*/;
assign _15202_ = _14653_ ^ _15204_ /*19459*/;
assign _15203_ = _15195_ & _15202_ /*19457*/;
assign _15200_ = _15201_ | _15203_ /*19455*/;
assign _15039_ = _15195_ ^ _15202_ /*19458*/;
assign _15209_ = D[25] ^ Q[25] /*19454*/;
assign _15206_ = _14654_ & _15209_ /*19450*/;
assign _15207_ = _14654_ ^ _15209_ /*19453*/;
assign _15208_ = _15200_ & _15207_ /*19451*/;
assign _15205_ = _15206_ | _15208_ /*19449*/;
assign _15040_ = _15200_ ^ _15207_ /*19452*/;
assign _15214_ = D[26] ^ Q[25] /*19448*/;
assign _15211_ = _14655_ & _15214_ /*19444*/;
assign _15212_ = _14655_ ^ _15214_ /*19447*/;
assign _15213_ = _15205_ & _15212_ /*19445*/;
assign _15210_ = _15211_ | _15213_ /*19443*/;
assign _15041_ = _15205_ ^ _15212_ /*19446*/;
assign _15219_ = D[27] ^ Q[25] /*19442*/;
assign _15216_ = _14656_ & _15219_ /*19438*/;
assign _15217_ = _14656_ ^ _15219_ /*19441*/;
assign _15218_ = _15210_ & _15217_ /*19439*/;
assign _15215_ = _15216_ | _15218_ /*19437*/;
assign _15042_ = _15210_ ^ _15217_ /*19440*/;
assign _15224_ = D[28] ^ Q[25] /*19436*/;
assign _15221_ = _14657_ & _15224_ /*19432*/;
assign _15222_ = _14657_ ^ _15224_ /*19435*/;
assign _15223_ = _15215_ & _15222_ /*19433*/;
assign _15220_ = _15221_ | _15223_ /*19431*/;
assign _15043_ = _15215_ ^ _15222_ /*19434*/;
assign _15229_ = D[29] ^ Q[25] /*19430*/;
assign _15226_ = _14658_ & _15229_ /*19426*/;
assign _15227_ = _14658_ ^ _15229_ /*19429*/;
assign _15228_ = _15220_ & _15227_ /*19427*/;
assign _15225_ = _15226_ | _15228_ /*19425*/;
assign _15044_ = _15220_ ^ _15227_ /*19428*/;
assign _15234_ = D[30] ^ Q[25] /*19424*/;
assign _15231_ = _14659_ & _15234_ /*19420*/;
assign _15232_ = _14659_ ^ _15234_ /*19423*/;
assign _15233_ = _15225_ & _15232_ /*19421*/;
assign _15230_ = _15231_ | _15233_ /*19419*/;
assign _15045_ = _15225_ ^ _15232_ /*19422*/;
assign _15239_ = D[31] ^ Q[25] /*19418*/;
assign _15236_ = _14660_ & _15239_ /*19414*/;
assign _15237_ = _14660_ ^ _15239_ /*19417*/;
assign _15238_ = _15230_ & _15237_ /*19415*/;
assign _15235_ = _15236_ | _15238_ /*19413*/;
assign _15046_ = _15230_ ^ _15237_ /*19416*/;
assign _15244_ = D[32] ^ Q[25] /*19412*/;
assign _15241_ = _14661_ & _15244_ /*19408*/;
assign _15242_ = _14661_ ^ _15244_ /*19411*/;
assign _15243_ = _15235_ & _15242_ /*19409*/;
assign _15240_ = _15241_ | _15243_ /*19407*/;
assign _15047_ = _15235_ ^ _15242_ /*19410*/;
assign _15249_ = D[33] ^ Q[25] /*19406*/;
assign _15246_ = _14662_ & _15249_ /*19402*/;
assign _15247_ = _14662_ ^ _15249_ /*19405*/;
assign _15248_ = _15240_ & _15247_ /*19403*/;
assign _15245_ = _15246_ | _15248_ /*19401*/;
assign _15048_ = _15240_ ^ _15247_ /*19404*/;
assign _15254_ = D[34] ^ Q[25] /*19400*/;
assign _15251_ = _14663_ & _15254_ /*19396*/;
assign _15252_ = _14663_ ^ _15254_ /*19399*/;
assign _15253_ = _15245_ & _15252_ /*19397*/;
assign _15250_ = _15251_ | _15253_ /*19395*/;
assign _15049_ = _15245_ ^ _15252_ /*19398*/;
assign _15259_ = D[35] ^ Q[25] /*19394*/;
assign _15256_ = _14664_ & _15259_ /*19390*/;
assign _15257_ = _14664_ ^ _15259_ /*19393*/;
assign _15258_ = _15250_ & _15257_ /*19391*/;
assign _15255_ = _15256_ | _15258_ /*19389*/;
assign _15050_ = _15250_ ^ _15257_ /*19392*/;
assign _15264_ = D[36] ^ Q[25] /*19388*/;
assign _15261_ = _14665_ & _15264_ /*19384*/;
assign _15262_ = _14665_ ^ _15264_ /*19387*/;
assign _15263_ = _15255_ & _15262_ /*19385*/;
assign _15260_ = _15261_ | _15263_ /*19383*/;
assign _15051_ = _15255_ ^ _15262_ /*19386*/;
assign _15269_ = D[37] ^ Q[25] /*19382*/;
assign _15266_ = _14666_ & _15269_ /*19378*/;
assign _15267_ = _14666_ ^ _15269_ /*19381*/;
assign _15268_ = _15260_ & _15267_ /*19379*/;
assign _15265_ = _15266_ | _15268_ /*19377*/;
assign _15052_ = _15260_ ^ _15267_ /*19380*/;
assign _15274_ = D[38] ^ Q[25] /*19376*/;
assign _15271_ = _14667_ & _15274_ /*19372*/;
assign _15272_ = _14667_ ^ _15274_ /*19375*/;
assign _15273_ = _15265_ & _15272_ /*19373*/;
assign _15270_ = _15271_ | _15273_ /*19371*/;
assign _15053_ = _15265_ ^ _15272_ /*19374*/;
assign _15279_ = D[39] ^ Q[25] /*19370*/;
assign _15276_ = _14668_ & _15279_ /*19366*/;
assign _15277_ = _14668_ ^ _15279_ /*19369*/;
assign _15278_ = _15270_ & _15277_ /*19367*/;
assign _15275_ = _15276_ | _15278_ /*19365*/;
assign _15054_ = _15270_ ^ _15277_ /*19368*/;
assign _15284_ = D[40] ^ Q[25] /*19364*/;
assign _15281_ = _14669_ & _15284_ /*19360*/;
assign _15282_ = _14669_ ^ _15284_ /*19363*/;
assign _15283_ = _15275_ & _15282_ /*19361*/;
assign _15280_ = _15281_ | _15283_ /*19359*/;
assign _15055_ = _15275_ ^ _15282_ /*19362*/;
assign _15289_ = D[41] ^ Q[25] /*19358*/;
assign _15286_ = _14670_ & _15289_ /*19354*/;
assign _15287_ = _14670_ ^ _15289_ /*19357*/;
assign _15288_ = _15280_ & _15287_ /*19355*/;
assign _15285_ = _15286_ | _15288_ /*19353*/;
assign _15056_ = _15280_ ^ _15287_ /*19356*/;
assign _15294_ = D[42] ^ Q[25] /*19352*/;
assign _15291_ = _14671_ & _15294_ /*19348*/;
assign _15292_ = _14671_ ^ _15294_ /*19351*/;
assign _15293_ = _15285_ & _15292_ /*19349*/;
assign _15290_ = _15291_ | _15293_ /*19347*/;
assign _15057_ = _15285_ ^ _15292_ /*19350*/;
assign _15299_ = D[43] ^ Q[25] /*19346*/;
assign _15296_ = _14672_ & _15299_ /*19342*/;
assign _15297_ = _14672_ ^ _15299_ /*19345*/;
assign _15298_ = _15290_ & _15297_ /*19343*/;
assign _15295_ = _15296_ | _15298_ /*19341*/;
assign _15058_ = _15290_ ^ _15297_ /*19344*/;
assign _15304_ = D[44] ^ Q[25] /*19340*/;
assign _15301_ = _14673_ & _15304_ /*19336*/;
assign _15302_ = _14673_ ^ _15304_ /*19339*/;
assign _15303_ = _15295_ & _15302_ /*19337*/;
assign _15300_ = _15301_ | _15303_ /*19335*/;
assign _15059_ = _15295_ ^ _15302_ /*19338*/;
assign _15309_ = D[45] ^ Q[25] /*19334*/;
assign _15306_ = _14674_ & _15309_ /*19330*/;
assign _15307_ = _14674_ ^ _15309_ /*19333*/;
assign _15308_ = _15300_ & _15307_ /*19331*/;
assign _15305_ = _15306_ | _15308_ /*19329*/;
assign _15060_ = _15300_ ^ _15307_ /*19332*/;
assign _15314_ = D[46] ^ Q[25] /*19328*/;
assign _15311_ = _14675_ & _15314_ /*19324*/;
assign _15312_ = _14675_ ^ _15314_ /*19327*/;
assign _15313_ = _15305_ & _15312_ /*19325*/;
assign _15310_ = _15311_ | _15313_ /*19323*/;
assign _15061_ = _15305_ ^ _15312_ /*19326*/;
assign _15319_ = D[47] ^ Q[25] /*19322*/;
assign _15316_ = _14676_ & _15319_ /*19318*/;
assign _15317_ = _14676_ ^ _15319_ /*19321*/;
assign _15318_ = _15310_ & _15317_ /*19319*/;
assign _15315_ = _15316_ | _15318_ /*19317*/;
assign _15062_ = _15310_ ^ _15317_ /*19320*/;
assign _15324_ = D[48] ^ Q[25] /*19316*/;
assign _15321_ = _14677_ & _15324_ /*19312*/;
assign _15322_ = _14677_ ^ _15324_ /*19315*/;
assign _15323_ = _15315_ & _15322_ /*19313*/;
assign _15320_ = _15321_ | _15323_ /*19311*/;
assign _15063_ = _15315_ ^ _15322_ /*19314*/;
assign _15329_ = D[49] ^ Q[25] /*19310*/;
assign _15326_ = _14678_ & _15329_ /*19306*/;
assign _15327_ = _14678_ ^ _15329_ /*19309*/;
assign _15328_ = _15320_ & _15327_ /*19307*/;
assign _15325_ = _15326_ | _15328_ /*19305*/;
assign _15064_ = _15320_ ^ _15327_ /*19308*/;
assign _15334_ = D[50] ^ Q[25] /*19304*/;
assign _15331_ = _14679_ & _15334_ /*19300*/;
assign _15332_ = _14679_ ^ _15334_ /*19303*/;
assign _15333_ = _15325_ & _15332_ /*19301*/;
assign _15330_ = _15331_ | _15333_ /*19299*/;
assign _15065_ = _15325_ ^ _15332_ /*19302*/;
assign _15339_ = D[51] ^ Q[25] /*19298*/;
assign _15336_ = _14680_ & _15339_ /*19294*/;
assign _15337_ = _14680_ ^ _15339_ /*19297*/;
assign _15338_ = _15330_ & _15337_ /*19295*/;
assign _15335_ = _15336_ | _15338_ /*19293*/;
assign _15066_ = _15330_ ^ _15337_ /*19296*/;
assign _15344_ = D[52] ^ Q[25] /*19292*/;
assign _15341_ = _14681_ & _15344_ /*19288*/;
assign _15342_ = _14681_ ^ _15344_ /*19291*/;
assign _15343_ = _15335_ & _15342_ /*19289*/;
assign _15340_ = _15341_ | _15343_ /*19287*/;
assign _15067_ = _15335_ ^ _15342_ /*19290*/;
assign _15349_ = D[53] ^ Q[25] /*19286*/;
assign _15346_ = _14682_ & _15349_ /*19282*/;
assign _15347_ = _14682_ ^ _15349_ /*19285*/;
assign _15348_ = _15340_ & _15347_ /*19283*/;
assign _15345_ = _15346_ | _15348_ /*19281*/;
assign _15068_ = _15340_ ^ _15347_ /*19284*/;
assign _15354_ = D[54] ^ Q[25] /*19280*/;
assign _15351_ = _14683_ & _15354_ /*19276*/;
assign _15352_ = _14683_ ^ _15354_ /*19279*/;
assign _15353_ = _15345_ & _15352_ /*19277*/;
assign _15350_ = _15351_ | _15353_ /*19275*/;
assign _15069_ = _15345_ ^ _15352_ /*19278*/;
assign _15359_ = D[55] ^ Q[25] /*19274*/;
assign _15356_ = _14684_ & _15359_ /*19270*/;
assign _15357_ = _14684_ ^ _15359_ /*19273*/;
assign _15358_ = _15350_ & _15357_ /*19271*/;
assign _15355_ = _15356_ | _15358_ /*19269*/;
assign _15070_ = _15350_ ^ _15357_ /*19272*/;
assign _15364_ = D[56] ^ Q[25] /*19268*/;
assign _15361_ = _14685_ & _15364_ /*19264*/;
assign _15362_ = _14685_ ^ _15364_ /*19267*/;
assign _15363_ = _15355_ & _15362_ /*19265*/;
assign _15360_ = _15361_ | _15363_ /*19263*/;
assign _15071_ = _15355_ ^ _15362_ /*19266*/;
assign _15369_ = D[57] ^ Q[25] /*19262*/;
assign _15366_ = _14686_ & _15369_ /*19258*/;
assign _15367_ = _14686_ ^ _15369_ /*19261*/;
assign _15368_ = _15360_ & _15367_ /*19259*/;
assign _15365_ = _15366_ | _15368_ /*19257*/;
assign _15072_ = _15360_ ^ _15367_ /*19260*/;
assign _15374_ = D[58] ^ Q[25] /*19256*/;
assign _15371_ = _14687_ & _15374_ /*19252*/;
assign _15372_ = _14687_ ^ _15374_ /*19255*/;
assign _15373_ = _15365_ & _15372_ /*19253*/;
assign _15370_ = _15371_ | _15373_ /*19251*/;
assign _15073_ = _15365_ ^ _15372_ /*19254*/;
assign _15379_ = D[59] ^ Q[25] /*19250*/;
assign _15376_ = _14688_ & _15379_ /*19246*/;
assign _15377_ = _14688_ ^ _15379_ /*19249*/;
assign _15378_ = _15370_ & _15377_ /*19247*/;
assign _15375_ = _15376_ | _15378_ /*19245*/;
assign _15074_ = _15370_ ^ _15377_ /*19248*/;
assign _15384_ = D[60] ^ Q[25] /*19244*/;
assign _15381_ = _14689_ & _15384_ /*19240*/;
assign _15382_ = _14689_ ^ _15384_ /*19243*/;
assign _15383_ = _15375_ & _15382_ /*19241*/;
assign _15380_ = _15381_ | _15383_ /*19239*/;
assign _15075_ = _15375_ ^ _15382_ /*19242*/;
assign _15389_ = D[61] ^ Q[25] /*19238*/;
assign _15386_ = _14690_ & _15389_ /*19234*/;
assign _15387_ = _14690_ ^ _15389_ /*19237*/;
assign _15388_ = _15380_ & _15387_ /*19235*/;
assign _15385_ = _15386_ | _15388_ /*19233*/;
assign _15076_ = _15380_ ^ _15387_ /*19236*/;
assign _15394_ = D[62] ^ Q[25] /*19232*/;
assign _15391_ = _14691_ & _15394_ /*19228*/;
assign _15392_ = _14691_ ^ _15394_ /*19231*/;
assign _15393_ = _15385_ & _15392_ /*19229*/;
assign _15390_ = _15391_ | _15393_ /*19227*/;
assign _15077_ = _15385_ ^ _15392_ /*19230*/;
assign _15398_ = zeroWire ^ Q[25] /*19226*/;
assign _15395_ = _14692_ & _15398_ /*19222*/;
assign _15396_ = _14692_ ^ _15398_ /*19225*/;
assign _15397_ = _15390_ & _15396_ /*19223*/;
assign Q[24] = _15395_ | _15397_ /*19221*/;
assign _15078_ = _15390_ ^ _15396_ /*19224*/;
assign _15469_ = D[0] ^ Q[24] /*18835*/;
assign _15466_ = R_0[23] & _15469_ /*18831*/;
assign _15467_ = R_0[23] ^ _15469_ /*18834*/;
assign _15468_ = Q[24] & _15467_ /*18832*/;
assign _15465_ = _15466_ | _15468_ /*18830*/;
assign _15400_ = Q[24] ^ _15467_ /*18833*/;
assign _15474_ = D[1] ^ Q[24] /*18829*/;
assign _15471_ = _15015_ & _15474_ /*18825*/;
assign _15472_ = _15015_ ^ _15474_ /*18828*/;
assign _15473_ = _15465_ & _15472_ /*18826*/;
assign _15470_ = _15471_ | _15473_ /*18824*/;
assign _15401_ = _15465_ ^ _15472_ /*18827*/;
assign _15479_ = D[2] ^ Q[24] /*18823*/;
assign _15476_ = _15016_ & _15479_ /*18819*/;
assign _15477_ = _15016_ ^ _15479_ /*18822*/;
assign _15478_ = _15470_ & _15477_ /*18820*/;
assign _15475_ = _15476_ | _15478_ /*18818*/;
assign _15402_ = _15470_ ^ _15477_ /*18821*/;
assign _15484_ = D[3] ^ Q[24] /*18817*/;
assign _15481_ = _15017_ & _15484_ /*18813*/;
assign _15482_ = _15017_ ^ _15484_ /*18816*/;
assign _15483_ = _15475_ & _15482_ /*18814*/;
assign _15480_ = _15481_ | _15483_ /*18812*/;
assign _15403_ = _15475_ ^ _15482_ /*18815*/;
assign _15489_ = D[4] ^ Q[24] /*18811*/;
assign _15486_ = _15018_ & _15489_ /*18807*/;
assign _15487_ = _15018_ ^ _15489_ /*18810*/;
assign _15488_ = _15480_ & _15487_ /*18808*/;
assign _15485_ = _15486_ | _15488_ /*18806*/;
assign _15404_ = _15480_ ^ _15487_ /*18809*/;
assign _15494_ = D[5] ^ Q[24] /*18805*/;
assign _15491_ = _15019_ & _15494_ /*18801*/;
assign _15492_ = _15019_ ^ _15494_ /*18804*/;
assign _15493_ = _15485_ & _15492_ /*18802*/;
assign _15490_ = _15491_ | _15493_ /*18800*/;
assign _15405_ = _15485_ ^ _15492_ /*18803*/;
assign _15499_ = D[6] ^ Q[24] /*18799*/;
assign _15496_ = _15020_ & _15499_ /*18795*/;
assign _15497_ = _15020_ ^ _15499_ /*18798*/;
assign _15498_ = _15490_ & _15497_ /*18796*/;
assign _15495_ = _15496_ | _15498_ /*18794*/;
assign _15406_ = _15490_ ^ _15497_ /*18797*/;
assign _15504_ = D[7] ^ Q[24] /*18793*/;
assign _15501_ = _15021_ & _15504_ /*18789*/;
assign _15502_ = _15021_ ^ _15504_ /*18792*/;
assign _15503_ = _15495_ & _15502_ /*18790*/;
assign _15500_ = _15501_ | _15503_ /*18788*/;
assign _15407_ = _15495_ ^ _15502_ /*18791*/;
assign _15509_ = D[8] ^ Q[24] /*18787*/;
assign _15506_ = _15022_ & _15509_ /*18783*/;
assign _15507_ = _15022_ ^ _15509_ /*18786*/;
assign _15508_ = _15500_ & _15507_ /*18784*/;
assign _15505_ = _15506_ | _15508_ /*18782*/;
assign _15408_ = _15500_ ^ _15507_ /*18785*/;
assign _15514_ = D[9] ^ Q[24] /*18781*/;
assign _15511_ = _15023_ & _15514_ /*18777*/;
assign _15512_ = _15023_ ^ _15514_ /*18780*/;
assign _15513_ = _15505_ & _15512_ /*18778*/;
assign _15510_ = _15511_ | _15513_ /*18776*/;
assign _15409_ = _15505_ ^ _15512_ /*18779*/;
assign _15519_ = D[10] ^ Q[24] /*18775*/;
assign _15516_ = _15024_ & _15519_ /*18771*/;
assign _15517_ = _15024_ ^ _15519_ /*18774*/;
assign _15518_ = _15510_ & _15517_ /*18772*/;
assign _15515_ = _15516_ | _15518_ /*18770*/;
assign _15410_ = _15510_ ^ _15517_ /*18773*/;
assign _15524_ = D[11] ^ Q[24] /*18769*/;
assign _15521_ = _15025_ & _15524_ /*18765*/;
assign _15522_ = _15025_ ^ _15524_ /*18768*/;
assign _15523_ = _15515_ & _15522_ /*18766*/;
assign _15520_ = _15521_ | _15523_ /*18764*/;
assign _15411_ = _15515_ ^ _15522_ /*18767*/;
assign _15529_ = D[12] ^ Q[24] /*18763*/;
assign _15526_ = _15026_ & _15529_ /*18759*/;
assign _15527_ = _15026_ ^ _15529_ /*18762*/;
assign _15528_ = _15520_ & _15527_ /*18760*/;
assign _15525_ = _15526_ | _15528_ /*18758*/;
assign _15412_ = _15520_ ^ _15527_ /*18761*/;
assign _15534_ = D[13] ^ Q[24] /*18757*/;
assign _15531_ = _15027_ & _15534_ /*18753*/;
assign _15532_ = _15027_ ^ _15534_ /*18756*/;
assign _15533_ = _15525_ & _15532_ /*18754*/;
assign _15530_ = _15531_ | _15533_ /*18752*/;
assign _15413_ = _15525_ ^ _15532_ /*18755*/;
assign _15539_ = D[14] ^ Q[24] /*18751*/;
assign _15536_ = _15028_ & _15539_ /*18747*/;
assign _15537_ = _15028_ ^ _15539_ /*18750*/;
assign _15538_ = _15530_ & _15537_ /*18748*/;
assign _15535_ = _15536_ | _15538_ /*18746*/;
assign _15414_ = _15530_ ^ _15537_ /*18749*/;
assign _15544_ = D[15] ^ Q[24] /*18745*/;
assign _15541_ = _15029_ & _15544_ /*18741*/;
assign _15542_ = _15029_ ^ _15544_ /*18744*/;
assign _15543_ = _15535_ & _15542_ /*18742*/;
assign _15540_ = _15541_ | _15543_ /*18740*/;
assign _15415_ = _15535_ ^ _15542_ /*18743*/;
assign _15549_ = D[16] ^ Q[24] /*18739*/;
assign _15546_ = _15030_ & _15549_ /*18735*/;
assign _15547_ = _15030_ ^ _15549_ /*18738*/;
assign _15548_ = _15540_ & _15547_ /*18736*/;
assign _15545_ = _15546_ | _15548_ /*18734*/;
assign _15416_ = _15540_ ^ _15547_ /*18737*/;
assign _15554_ = D[17] ^ Q[24] /*18733*/;
assign _15551_ = _15031_ & _15554_ /*18729*/;
assign _15552_ = _15031_ ^ _15554_ /*18732*/;
assign _15553_ = _15545_ & _15552_ /*18730*/;
assign _15550_ = _15551_ | _15553_ /*18728*/;
assign _15417_ = _15545_ ^ _15552_ /*18731*/;
assign _15559_ = D[18] ^ Q[24] /*18727*/;
assign _15556_ = _15032_ & _15559_ /*18723*/;
assign _15557_ = _15032_ ^ _15559_ /*18726*/;
assign _15558_ = _15550_ & _15557_ /*18724*/;
assign _15555_ = _15556_ | _15558_ /*18722*/;
assign _15418_ = _15550_ ^ _15557_ /*18725*/;
assign _15564_ = D[19] ^ Q[24] /*18721*/;
assign _15561_ = _15033_ & _15564_ /*18717*/;
assign _15562_ = _15033_ ^ _15564_ /*18720*/;
assign _15563_ = _15555_ & _15562_ /*18718*/;
assign _15560_ = _15561_ | _15563_ /*18716*/;
assign _15419_ = _15555_ ^ _15562_ /*18719*/;
assign _15569_ = D[20] ^ Q[24] /*18715*/;
assign _15566_ = _15034_ & _15569_ /*18711*/;
assign _15567_ = _15034_ ^ _15569_ /*18714*/;
assign _15568_ = _15560_ & _15567_ /*18712*/;
assign _15565_ = _15566_ | _15568_ /*18710*/;
assign _15420_ = _15560_ ^ _15567_ /*18713*/;
assign _15574_ = D[21] ^ Q[24] /*18709*/;
assign _15571_ = _15035_ & _15574_ /*18705*/;
assign _15572_ = _15035_ ^ _15574_ /*18708*/;
assign _15573_ = _15565_ & _15572_ /*18706*/;
assign _15570_ = _15571_ | _15573_ /*18704*/;
assign _15421_ = _15565_ ^ _15572_ /*18707*/;
assign _15579_ = D[22] ^ Q[24] /*18703*/;
assign _15576_ = _15036_ & _15579_ /*18699*/;
assign _15577_ = _15036_ ^ _15579_ /*18702*/;
assign _15578_ = _15570_ & _15577_ /*18700*/;
assign _15575_ = _15576_ | _15578_ /*18698*/;
assign _15422_ = _15570_ ^ _15577_ /*18701*/;
assign _15584_ = D[23] ^ Q[24] /*18697*/;
assign _15581_ = _15037_ & _15584_ /*18693*/;
assign _15582_ = _15037_ ^ _15584_ /*18696*/;
assign _15583_ = _15575_ & _15582_ /*18694*/;
assign _15580_ = _15581_ | _15583_ /*18692*/;
assign _15423_ = _15575_ ^ _15582_ /*18695*/;
assign _15589_ = D[24] ^ Q[24] /*18691*/;
assign _15586_ = _15038_ & _15589_ /*18687*/;
assign _15587_ = _15038_ ^ _15589_ /*18690*/;
assign _15588_ = _15580_ & _15587_ /*18688*/;
assign _15585_ = _15586_ | _15588_ /*18686*/;
assign _15424_ = _15580_ ^ _15587_ /*18689*/;
assign _15594_ = D[25] ^ Q[24] /*18685*/;
assign _15591_ = _15039_ & _15594_ /*18681*/;
assign _15592_ = _15039_ ^ _15594_ /*18684*/;
assign _15593_ = _15585_ & _15592_ /*18682*/;
assign _15590_ = _15591_ | _15593_ /*18680*/;
assign _15425_ = _15585_ ^ _15592_ /*18683*/;
assign _15599_ = D[26] ^ Q[24] /*18679*/;
assign _15596_ = _15040_ & _15599_ /*18675*/;
assign _15597_ = _15040_ ^ _15599_ /*18678*/;
assign _15598_ = _15590_ & _15597_ /*18676*/;
assign _15595_ = _15596_ | _15598_ /*18674*/;
assign _15426_ = _15590_ ^ _15597_ /*18677*/;
assign _15604_ = D[27] ^ Q[24] /*18673*/;
assign _15601_ = _15041_ & _15604_ /*18669*/;
assign _15602_ = _15041_ ^ _15604_ /*18672*/;
assign _15603_ = _15595_ & _15602_ /*18670*/;
assign _15600_ = _15601_ | _15603_ /*18668*/;
assign _15427_ = _15595_ ^ _15602_ /*18671*/;
assign _15609_ = D[28] ^ Q[24] /*18667*/;
assign _15606_ = _15042_ & _15609_ /*18663*/;
assign _15607_ = _15042_ ^ _15609_ /*18666*/;
assign _15608_ = _15600_ & _15607_ /*18664*/;
assign _15605_ = _15606_ | _15608_ /*18662*/;
assign _15428_ = _15600_ ^ _15607_ /*18665*/;
assign _15614_ = D[29] ^ Q[24] /*18661*/;
assign _15611_ = _15043_ & _15614_ /*18657*/;
assign _15612_ = _15043_ ^ _15614_ /*18660*/;
assign _15613_ = _15605_ & _15612_ /*18658*/;
assign _15610_ = _15611_ | _15613_ /*18656*/;
assign _15429_ = _15605_ ^ _15612_ /*18659*/;
assign _15619_ = D[30] ^ Q[24] /*18655*/;
assign _15616_ = _15044_ & _15619_ /*18651*/;
assign _15617_ = _15044_ ^ _15619_ /*18654*/;
assign _15618_ = _15610_ & _15617_ /*18652*/;
assign _15615_ = _15616_ | _15618_ /*18650*/;
assign _15430_ = _15610_ ^ _15617_ /*18653*/;
assign _15624_ = D[31] ^ Q[24] /*18649*/;
assign _15621_ = _15045_ & _15624_ /*18645*/;
assign _15622_ = _15045_ ^ _15624_ /*18648*/;
assign _15623_ = _15615_ & _15622_ /*18646*/;
assign _15620_ = _15621_ | _15623_ /*18644*/;
assign _15431_ = _15615_ ^ _15622_ /*18647*/;
assign _15629_ = D[32] ^ Q[24] /*18643*/;
assign _15626_ = _15046_ & _15629_ /*18639*/;
assign _15627_ = _15046_ ^ _15629_ /*18642*/;
assign _15628_ = _15620_ & _15627_ /*18640*/;
assign _15625_ = _15626_ | _15628_ /*18638*/;
assign _15432_ = _15620_ ^ _15627_ /*18641*/;
assign _15634_ = D[33] ^ Q[24] /*18637*/;
assign _15631_ = _15047_ & _15634_ /*18633*/;
assign _15632_ = _15047_ ^ _15634_ /*18636*/;
assign _15633_ = _15625_ & _15632_ /*18634*/;
assign _15630_ = _15631_ | _15633_ /*18632*/;
assign _15433_ = _15625_ ^ _15632_ /*18635*/;
assign _15639_ = D[34] ^ Q[24] /*18631*/;
assign _15636_ = _15048_ & _15639_ /*18627*/;
assign _15637_ = _15048_ ^ _15639_ /*18630*/;
assign _15638_ = _15630_ & _15637_ /*18628*/;
assign _15635_ = _15636_ | _15638_ /*18626*/;
assign _15434_ = _15630_ ^ _15637_ /*18629*/;
assign _15644_ = D[35] ^ Q[24] /*18625*/;
assign _15641_ = _15049_ & _15644_ /*18621*/;
assign _15642_ = _15049_ ^ _15644_ /*18624*/;
assign _15643_ = _15635_ & _15642_ /*18622*/;
assign _15640_ = _15641_ | _15643_ /*18620*/;
assign _15435_ = _15635_ ^ _15642_ /*18623*/;
assign _15649_ = D[36] ^ Q[24] /*18619*/;
assign _15646_ = _15050_ & _15649_ /*18615*/;
assign _15647_ = _15050_ ^ _15649_ /*18618*/;
assign _15648_ = _15640_ & _15647_ /*18616*/;
assign _15645_ = _15646_ | _15648_ /*18614*/;
assign _15436_ = _15640_ ^ _15647_ /*18617*/;
assign _15654_ = D[37] ^ Q[24] /*18613*/;
assign _15651_ = _15051_ & _15654_ /*18609*/;
assign _15652_ = _15051_ ^ _15654_ /*18612*/;
assign _15653_ = _15645_ & _15652_ /*18610*/;
assign _15650_ = _15651_ | _15653_ /*18608*/;
assign _15437_ = _15645_ ^ _15652_ /*18611*/;
assign _15659_ = D[38] ^ Q[24] /*18607*/;
assign _15656_ = _15052_ & _15659_ /*18603*/;
assign _15657_ = _15052_ ^ _15659_ /*18606*/;
assign _15658_ = _15650_ & _15657_ /*18604*/;
assign _15655_ = _15656_ | _15658_ /*18602*/;
assign _15438_ = _15650_ ^ _15657_ /*18605*/;
assign _15664_ = D[39] ^ Q[24] /*18601*/;
assign _15661_ = _15053_ & _15664_ /*18597*/;
assign _15662_ = _15053_ ^ _15664_ /*18600*/;
assign _15663_ = _15655_ & _15662_ /*18598*/;
assign _15660_ = _15661_ | _15663_ /*18596*/;
assign _15439_ = _15655_ ^ _15662_ /*18599*/;
assign _15669_ = D[40] ^ Q[24] /*18595*/;
assign _15666_ = _15054_ & _15669_ /*18591*/;
assign _15667_ = _15054_ ^ _15669_ /*18594*/;
assign _15668_ = _15660_ & _15667_ /*18592*/;
assign _15665_ = _15666_ | _15668_ /*18590*/;
assign _15440_ = _15660_ ^ _15667_ /*18593*/;
assign _15674_ = D[41] ^ Q[24] /*18589*/;
assign _15671_ = _15055_ & _15674_ /*18585*/;
assign _15672_ = _15055_ ^ _15674_ /*18588*/;
assign _15673_ = _15665_ & _15672_ /*18586*/;
assign _15670_ = _15671_ | _15673_ /*18584*/;
assign _15441_ = _15665_ ^ _15672_ /*18587*/;
assign _15679_ = D[42] ^ Q[24] /*18583*/;
assign _15676_ = _15056_ & _15679_ /*18579*/;
assign _15677_ = _15056_ ^ _15679_ /*18582*/;
assign _15678_ = _15670_ & _15677_ /*18580*/;
assign _15675_ = _15676_ | _15678_ /*18578*/;
assign _15442_ = _15670_ ^ _15677_ /*18581*/;
assign _15684_ = D[43] ^ Q[24] /*18577*/;
assign _15681_ = _15057_ & _15684_ /*18573*/;
assign _15682_ = _15057_ ^ _15684_ /*18576*/;
assign _15683_ = _15675_ & _15682_ /*18574*/;
assign _15680_ = _15681_ | _15683_ /*18572*/;
assign _15443_ = _15675_ ^ _15682_ /*18575*/;
assign _15689_ = D[44] ^ Q[24] /*18571*/;
assign _15686_ = _15058_ & _15689_ /*18567*/;
assign _15687_ = _15058_ ^ _15689_ /*18570*/;
assign _15688_ = _15680_ & _15687_ /*18568*/;
assign _15685_ = _15686_ | _15688_ /*18566*/;
assign _15444_ = _15680_ ^ _15687_ /*18569*/;
assign _15694_ = D[45] ^ Q[24] /*18565*/;
assign _15691_ = _15059_ & _15694_ /*18561*/;
assign _15692_ = _15059_ ^ _15694_ /*18564*/;
assign _15693_ = _15685_ & _15692_ /*18562*/;
assign _15690_ = _15691_ | _15693_ /*18560*/;
assign _15445_ = _15685_ ^ _15692_ /*18563*/;
assign _15699_ = D[46] ^ Q[24] /*18559*/;
assign _15696_ = _15060_ & _15699_ /*18555*/;
assign _15697_ = _15060_ ^ _15699_ /*18558*/;
assign _15698_ = _15690_ & _15697_ /*18556*/;
assign _15695_ = _15696_ | _15698_ /*18554*/;
assign _15446_ = _15690_ ^ _15697_ /*18557*/;
assign _15704_ = D[47] ^ Q[24] /*18553*/;
assign _15701_ = _15061_ & _15704_ /*18549*/;
assign _15702_ = _15061_ ^ _15704_ /*18552*/;
assign _15703_ = _15695_ & _15702_ /*18550*/;
assign _15700_ = _15701_ | _15703_ /*18548*/;
assign _15447_ = _15695_ ^ _15702_ /*18551*/;
assign _15709_ = D[48] ^ Q[24] /*18547*/;
assign _15706_ = _15062_ & _15709_ /*18543*/;
assign _15707_ = _15062_ ^ _15709_ /*18546*/;
assign _15708_ = _15700_ & _15707_ /*18544*/;
assign _15705_ = _15706_ | _15708_ /*18542*/;
assign _15448_ = _15700_ ^ _15707_ /*18545*/;
assign _15714_ = D[49] ^ Q[24] /*18541*/;
assign _15711_ = _15063_ & _15714_ /*18537*/;
assign _15712_ = _15063_ ^ _15714_ /*18540*/;
assign _15713_ = _15705_ & _15712_ /*18538*/;
assign _15710_ = _15711_ | _15713_ /*18536*/;
assign _15449_ = _15705_ ^ _15712_ /*18539*/;
assign _15719_ = D[50] ^ Q[24] /*18535*/;
assign _15716_ = _15064_ & _15719_ /*18531*/;
assign _15717_ = _15064_ ^ _15719_ /*18534*/;
assign _15718_ = _15710_ & _15717_ /*18532*/;
assign _15715_ = _15716_ | _15718_ /*18530*/;
assign _15450_ = _15710_ ^ _15717_ /*18533*/;
assign _15724_ = D[51] ^ Q[24] /*18529*/;
assign _15721_ = _15065_ & _15724_ /*18525*/;
assign _15722_ = _15065_ ^ _15724_ /*18528*/;
assign _15723_ = _15715_ & _15722_ /*18526*/;
assign _15720_ = _15721_ | _15723_ /*18524*/;
assign _15451_ = _15715_ ^ _15722_ /*18527*/;
assign _15729_ = D[52] ^ Q[24] /*18523*/;
assign _15726_ = _15066_ & _15729_ /*18519*/;
assign _15727_ = _15066_ ^ _15729_ /*18522*/;
assign _15728_ = _15720_ & _15727_ /*18520*/;
assign _15725_ = _15726_ | _15728_ /*18518*/;
assign _15452_ = _15720_ ^ _15727_ /*18521*/;
assign _15734_ = D[53] ^ Q[24] /*18517*/;
assign _15731_ = _15067_ & _15734_ /*18513*/;
assign _15732_ = _15067_ ^ _15734_ /*18516*/;
assign _15733_ = _15725_ & _15732_ /*18514*/;
assign _15730_ = _15731_ | _15733_ /*18512*/;
assign _15453_ = _15725_ ^ _15732_ /*18515*/;
assign _15739_ = D[54] ^ Q[24] /*18511*/;
assign _15736_ = _15068_ & _15739_ /*18507*/;
assign _15737_ = _15068_ ^ _15739_ /*18510*/;
assign _15738_ = _15730_ & _15737_ /*18508*/;
assign _15735_ = _15736_ | _15738_ /*18506*/;
assign _15454_ = _15730_ ^ _15737_ /*18509*/;
assign _15744_ = D[55] ^ Q[24] /*18505*/;
assign _15741_ = _15069_ & _15744_ /*18501*/;
assign _15742_ = _15069_ ^ _15744_ /*18504*/;
assign _15743_ = _15735_ & _15742_ /*18502*/;
assign _15740_ = _15741_ | _15743_ /*18500*/;
assign _15455_ = _15735_ ^ _15742_ /*18503*/;
assign _15749_ = D[56] ^ Q[24] /*18499*/;
assign _15746_ = _15070_ & _15749_ /*18495*/;
assign _15747_ = _15070_ ^ _15749_ /*18498*/;
assign _15748_ = _15740_ & _15747_ /*18496*/;
assign _15745_ = _15746_ | _15748_ /*18494*/;
assign _15456_ = _15740_ ^ _15747_ /*18497*/;
assign _15754_ = D[57] ^ Q[24] /*18493*/;
assign _15751_ = _15071_ & _15754_ /*18489*/;
assign _15752_ = _15071_ ^ _15754_ /*18492*/;
assign _15753_ = _15745_ & _15752_ /*18490*/;
assign _15750_ = _15751_ | _15753_ /*18488*/;
assign _15457_ = _15745_ ^ _15752_ /*18491*/;
assign _15759_ = D[58] ^ Q[24] /*18487*/;
assign _15756_ = _15072_ & _15759_ /*18483*/;
assign _15757_ = _15072_ ^ _15759_ /*18486*/;
assign _15758_ = _15750_ & _15757_ /*18484*/;
assign _15755_ = _15756_ | _15758_ /*18482*/;
assign _15458_ = _15750_ ^ _15757_ /*18485*/;
assign _15764_ = D[59] ^ Q[24] /*18481*/;
assign _15761_ = _15073_ & _15764_ /*18477*/;
assign _15762_ = _15073_ ^ _15764_ /*18480*/;
assign _15763_ = _15755_ & _15762_ /*18478*/;
assign _15760_ = _15761_ | _15763_ /*18476*/;
assign _15459_ = _15755_ ^ _15762_ /*18479*/;
assign _15769_ = D[60] ^ Q[24] /*18475*/;
assign _15766_ = _15074_ & _15769_ /*18471*/;
assign _15767_ = _15074_ ^ _15769_ /*18474*/;
assign _15768_ = _15760_ & _15767_ /*18472*/;
assign _15765_ = _15766_ | _15768_ /*18470*/;
assign _15460_ = _15760_ ^ _15767_ /*18473*/;
assign _15774_ = D[61] ^ Q[24] /*18469*/;
assign _15771_ = _15075_ & _15774_ /*18465*/;
assign _15772_ = _15075_ ^ _15774_ /*18468*/;
assign _15773_ = _15765_ & _15772_ /*18466*/;
assign _15770_ = _15771_ | _15773_ /*18464*/;
assign _15461_ = _15765_ ^ _15772_ /*18467*/;
assign _15779_ = D[62] ^ Q[24] /*18463*/;
assign _15776_ = _15076_ & _15779_ /*18459*/;
assign _15777_ = _15076_ ^ _15779_ /*18462*/;
assign _15778_ = _15770_ & _15777_ /*18460*/;
assign _15775_ = _15776_ | _15778_ /*18458*/;
assign _15462_ = _15770_ ^ _15777_ /*18461*/;
assign _15783_ = zeroWire ^ Q[24] /*18457*/;
assign _15780_ = _15077_ & _15783_ /*18453*/;
assign _15781_ = _15077_ ^ _15783_ /*18456*/;
assign _15782_ = _15775_ & _15781_ /*18454*/;
assign Q[23] = _15780_ | _15782_ /*18452*/;
assign _15463_ = _15775_ ^ _15781_ /*18455*/;
assign _15854_ = D[0] ^ Q[23] /*18066*/;
assign _15851_ = R_0[22] & _15854_ /*18062*/;
assign _15852_ = R_0[22] ^ _15854_ /*18065*/;
assign _15853_ = Q[23] & _15852_ /*18063*/;
assign _15850_ = _15851_ | _15853_ /*18061*/;
assign _15785_ = Q[23] ^ _15852_ /*18064*/;
assign _15859_ = D[1] ^ Q[23] /*18060*/;
assign _15856_ = _15400_ & _15859_ /*18056*/;
assign _15857_ = _15400_ ^ _15859_ /*18059*/;
assign _15858_ = _15850_ & _15857_ /*18057*/;
assign _15855_ = _15856_ | _15858_ /*18055*/;
assign _15786_ = _15850_ ^ _15857_ /*18058*/;
assign _15864_ = D[2] ^ Q[23] /*18054*/;
assign _15861_ = _15401_ & _15864_ /*18050*/;
assign _15862_ = _15401_ ^ _15864_ /*18053*/;
assign _15863_ = _15855_ & _15862_ /*18051*/;
assign _15860_ = _15861_ | _15863_ /*18049*/;
assign _15787_ = _15855_ ^ _15862_ /*18052*/;
assign _15869_ = D[3] ^ Q[23] /*18048*/;
assign _15866_ = _15402_ & _15869_ /*18044*/;
assign _15867_ = _15402_ ^ _15869_ /*18047*/;
assign _15868_ = _15860_ & _15867_ /*18045*/;
assign _15865_ = _15866_ | _15868_ /*18043*/;
assign _15788_ = _15860_ ^ _15867_ /*18046*/;
assign _15874_ = D[4] ^ Q[23] /*18042*/;
assign _15871_ = _15403_ & _15874_ /*18038*/;
assign _15872_ = _15403_ ^ _15874_ /*18041*/;
assign _15873_ = _15865_ & _15872_ /*18039*/;
assign _15870_ = _15871_ | _15873_ /*18037*/;
assign _15789_ = _15865_ ^ _15872_ /*18040*/;
assign _15879_ = D[5] ^ Q[23] /*18036*/;
assign _15876_ = _15404_ & _15879_ /*18032*/;
assign _15877_ = _15404_ ^ _15879_ /*18035*/;
assign _15878_ = _15870_ & _15877_ /*18033*/;
assign _15875_ = _15876_ | _15878_ /*18031*/;
assign _15790_ = _15870_ ^ _15877_ /*18034*/;
assign _15884_ = D[6] ^ Q[23] /*18030*/;
assign _15881_ = _15405_ & _15884_ /*18026*/;
assign _15882_ = _15405_ ^ _15884_ /*18029*/;
assign _15883_ = _15875_ & _15882_ /*18027*/;
assign _15880_ = _15881_ | _15883_ /*18025*/;
assign _15791_ = _15875_ ^ _15882_ /*18028*/;
assign _15889_ = D[7] ^ Q[23] /*18024*/;
assign _15886_ = _15406_ & _15889_ /*18020*/;
assign _15887_ = _15406_ ^ _15889_ /*18023*/;
assign _15888_ = _15880_ & _15887_ /*18021*/;
assign _15885_ = _15886_ | _15888_ /*18019*/;
assign _15792_ = _15880_ ^ _15887_ /*18022*/;
assign _15894_ = D[8] ^ Q[23] /*18018*/;
assign _15891_ = _15407_ & _15894_ /*18014*/;
assign _15892_ = _15407_ ^ _15894_ /*18017*/;
assign _15893_ = _15885_ & _15892_ /*18015*/;
assign _15890_ = _15891_ | _15893_ /*18013*/;
assign _15793_ = _15885_ ^ _15892_ /*18016*/;
assign _15899_ = D[9] ^ Q[23] /*18012*/;
assign _15896_ = _15408_ & _15899_ /*18008*/;
assign _15897_ = _15408_ ^ _15899_ /*18011*/;
assign _15898_ = _15890_ & _15897_ /*18009*/;
assign _15895_ = _15896_ | _15898_ /*18007*/;
assign _15794_ = _15890_ ^ _15897_ /*18010*/;
assign _15904_ = D[10] ^ Q[23] /*18006*/;
assign _15901_ = _15409_ & _15904_ /*18002*/;
assign _15902_ = _15409_ ^ _15904_ /*18005*/;
assign _15903_ = _15895_ & _15902_ /*18003*/;
assign _15900_ = _15901_ | _15903_ /*18001*/;
assign _15795_ = _15895_ ^ _15902_ /*18004*/;
assign _15909_ = D[11] ^ Q[23] /*18000*/;
assign _15906_ = _15410_ & _15909_ /*17996*/;
assign _15907_ = _15410_ ^ _15909_ /*17999*/;
assign _15908_ = _15900_ & _15907_ /*17997*/;
assign _15905_ = _15906_ | _15908_ /*17995*/;
assign _15796_ = _15900_ ^ _15907_ /*17998*/;
assign _15914_ = D[12] ^ Q[23] /*17994*/;
assign _15911_ = _15411_ & _15914_ /*17990*/;
assign _15912_ = _15411_ ^ _15914_ /*17993*/;
assign _15913_ = _15905_ & _15912_ /*17991*/;
assign _15910_ = _15911_ | _15913_ /*17989*/;
assign _15797_ = _15905_ ^ _15912_ /*17992*/;
assign _15919_ = D[13] ^ Q[23] /*17988*/;
assign _15916_ = _15412_ & _15919_ /*17984*/;
assign _15917_ = _15412_ ^ _15919_ /*17987*/;
assign _15918_ = _15910_ & _15917_ /*17985*/;
assign _15915_ = _15916_ | _15918_ /*17983*/;
assign _15798_ = _15910_ ^ _15917_ /*17986*/;
assign _15924_ = D[14] ^ Q[23] /*17982*/;
assign _15921_ = _15413_ & _15924_ /*17978*/;
assign _15922_ = _15413_ ^ _15924_ /*17981*/;
assign _15923_ = _15915_ & _15922_ /*17979*/;
assign _15920_ = _15921_ | _15923_ /*17977*/;
assign _15799_ = _15915_ ^ _15922_ /*17980*/;
assign _15929_ = D[15] ^ Q[23] /*17976*/;
assign _15926_ = _15414_ & _15929_ /*17972*/;
assign _15927_ = _15414_ ^ _15929_ /*17975*/;
assign _15928_ = _15920_ & _15927_ /*17973*/;
assign _15925_ = _15926_ | _15928_ /*17971*/;
assign _15800_ = _15920_ ^ _15927_ /*17974*/;
assign _15934_ = D[16] ^ Q[23] /*17970*/;
assign _15931_ = _15415_ & _15934_ /*17966*/;
assign _15932_ = _15415_ ^ _15934_ /*17969*/;
assign _15933_ = _15925_ & _15932_ /*17967*/;
assign _15930_ = _15931_ | _15933_ /*17965*/;
assign _15801_ = _15925_ ^ _15932_ /*17968*/;
assign _15939_ = D[17] ^ Q[23] /*17964*/;
assign _15936_ = _15416_ & _15939_ /*17960*/;
assign _15937_ = _15416_ ^ _15939_ /*17963*/;
assign _15938_ = _15930_ & _15937_ /*17961*/;
assign _15935_ = _15936_ | _15938_ /*17959*/;
assign _15802_ = _15930_ ^ _15937_ /*17962*/;
assign _15944_ = D[18] ^ Q[23] /*17958*/;
assign _15941_ = _15417_ & _15944_ /*17954*/;
assign _15942_ = _15417_ ^ _15944_ /*17957*/;
assign _15943_ = _15935_ & _15942_ /*17955*/;
assign _15940_ = _15941_ | _15943_ /*17953*/;
assign _15803_ = _15935_ ^ _15942_ /*17956*/;
assign _15949_ = D[19] ^ Q[23] /*17952*/;
assign _15946_ = _15418_ & _15949_ /*17948*/;
assign _15947_ = _15418_ ^ _15949_ /*17951*/;
assign _15948_ = _15940_ & _15947_ /*17949*/;
assign _15945_ = _15946_ | _15948_ /*17947*/;
assign _15804_ = _15940_ ^ _15947_ /*17950*/;
assign _15954_ = D[20] ^ Q[23] /*17946*/;
assign _15951_ = _15419_ & _15954_ /*17942*/;
assign _15952_ = _15419_ ^ _15954_ /*17945*/;
assign _15953_ = _15945_ & _15952_ /*17943*/;
assign _15950_ = _15951_ | _15953_ /*17941*/;
assign _15805_ = _15945_ ^ _15952_ /*17944*/;
assign _15959_ = D[21] ^ Q[23] /*17940*/;
assign _15956_ = _15420_ & _15959_ /*17936*/;
assign _15957_ = _15420_ ^ _15959_ /*17939*/;
assign _15958_ = _15950_ & _15957_ /*17937*/;
assign _15955_ = _15956_ | _15958_ /*17935*/;
assign _15806_ = _15950_ ^ _15957_ /*17938*/;
assign _15964_ = D[22] ^ Q[23] /*17934*/;
assign _15961_ = _15421_ & _15964_ /*17930*/;
assign _15962_ = _15421_ ^ _15964_ /*17933*/;
assign _15963_ = _15955_ & _15962_ /*17931*/;
assign _15960_ = _15961_ | _15963_ /*17929*/;
assign _15807_ = _15955_ ^ _15962_ /*17932*/;
assign _15969_ = D[23] ^ Q[23] /*17928*/;
assign _15966_ = _15422_ & _15969_ /*17924*/;
assign _15967_ = _15422_ ^ _15969_ /*17927*/;
assign _15968_ = _15960_ & _15967_ /*17925*/;
assign _15965_ = _15966_ | _15968_ /*17923*/;
assign _15808_ = _15960_ ^ _15967_ /*17926*/;
assign _15974_ = D[24] ^ Q[23] /*17922*/;
assign _15971_ = _15423_ & _15974_ /*17918*/;
assign _15972_ = _15423_ ^ _15974_ /*17921*/;
assign _15973_ = _15965_ & _15972_ /*17919*/;
assign _15970_ = _15971_ | _15973_ /*17917*/;
assign _15809_ = _15965_ ^ _15972_ /*17920*/;
assign _15979_ = D[25] ^ Q[23] /*17916*/;
assign _15976_ = _15424_ & _15979_ /*17912*/;
assign _15977_ = _15424_ ^ _15979_ /*17915*/;
assign _15978_ = _15970_ & _15977_ /*17913*/;
assign _15975_ = _15976_ | _15978_ /*17911*/;
assign _15810_ = _15970_ ^ _15977_ /*17914*/;
assign _15984_ = D[26] ^ Q[23] /*17910*/;
assign _15981_ = _15425_ & _15984_ /*17906*/;
assign _15982_ = _15425_ ^ _15984_ /*17909*/;
assign _15983_ = _15975_ & _15982_ /*17907*/;
assign _15980_ = _15981_ | _15983_ /*17905*/;
assign _15811_ = _15975_ ^ _15982_ /*17908*/;
assign _15989_ = D[27] ^ Q[23] /*17904*/;
assign _15986_ = _15426_ & _15989_ /*17900*/;
assign _15987_ = _15426_ ^ _15989_ /*17903*/;
assign _15988_ = _15980_ & _15987_ /*17901*/;
assign _15985_ = _15986_ | _15988_ /*17899*/;
assign _15812_ = _15980_ ^ _15987_ /*17902*/;
assign _15994_ = D[28] ^ Q[23] /*17898*/;
assign _15991_ = _15427_ & _15994_ /*17894*/;
assign _15992_ = _15427_ ^ _15994_ /*17897*/;
assign _15993_ = _15985_ & _15992_ /*17895*/;
assign _15990_ = _15991_ | _15993_ /*17893*/;
assign _15813_ = _15985_ ^ _15992_ /*17896*/;
assign _15999_ = D[29] ^ Q[23] /*17892*/;
assign _15996_ = _15428_ & _15999_ /*17888*/;
assign _15997_ = _15428_ ^ _15999_ /*17891*/;
assign _15998_ = _15990_ & _15997_ /*17889*/;
assign _15995_ = _15996_ | _15998_ /*17887*/;
assign _15814_ = _15990_ ^ _15997_ /*17890*/;
assign _16004_ = D[30] ^ Q[23] /*17886*/;
assign _16001_ = _15429_ & _16004_ /*17882*/;
assign _16002_ = _15429_ ^ _16004_ /*17885*/;
assign _16003_ = _15995_ & _16002_ /*17883*/;
assign _16000_ = _16001_ | _16003_ /*17881*/;
assign _15815_ = _15995_ ^ _16002_ /*17884*/;
assign _16009_ = D[31] ^ Q[23] /*17880*/;
assign _16006_ = _15430_ & _16009_ /*17876*/;
assign _16007_ = _15430_ ^ _16009_ /*17879*/;
assign _16008_ = _16000_ & _16007_ /*17877*/;
assign _16005_ = _16006_ | _16008_ /*17875*/;
assign _15816_ = _16000_ ^ _16007_ /*17878*/;
assign _16014_ = D[32] ^ Q[23] /*17874*/;
assign _16011_ = _15431_ & _16014_ /*17870*/;
assign _16012_ = _15431_ ^ _16014_ /*17873*/;
assign _16013_ = _16005_ & _16012_ /*17871*/;
assign _16010_ = _16011_ | _16013_ /*17869*/;
assign _15817_ = _16005_ ^ _16012_ /*17872*/;
assign _16019_ = D[33] ^ Q[23] /*17868*/;
assign _16016_ = _15432_ & _16019_ /*17864*/;
assign _16017_ = _15432_ ^ _16019_ /*17867*/;
assign _16018_ = _16010_ & _16017_ /*17865*/;
assign _16015_ = _16016_ | _16018_ /*17863*/;
assign _15818_ = _16010_ ^ _16017_ /*17866*/;
assign _16024_ = D[34] ^ Q[23] /*17862*/;
assign _16021_ = _15433_ & _16024_ /*17858*/;
assign _16022_ = _15433_ ^ _16024_ /*17861*/;
assign _16023_ = _16015_ & _16022_ /*17859*/;
assign _16020_ = _16021_ | _16023_ /*17857*/;
assign _15819_ = _16015_ ^ _16022_ /*17860*/;
assign _16029_ = D[35] ^ Q[23] /*17856*/;
assign _16026_ = _15434_ & _16029_ /*17852*/;
assign _16027_ = _15434_ ^ _16029_ /*17855*/;
assign _16028_ = _16020_ & _16027_ /*17853*/;
assign _16025_ = _16026_ | _16028_ /*17851*/;
assign _15820_ = _16020_ ^ _16027_ /*17854*/;
assign _16034_ = D[36] ^ Q[23] /*17850*/;
assign _16031_ = _15435_ & _16034_ /*17846*/;
assign _16032_ = _15435_ ^ _16034_ /*17849*/;
assign _16033_ = _16025_ & _16032_ /*17847*/;
assign _16030_ = _16031_ | _16033_ /*17845*/;
assign _15821_ = _16025_ ^ _16032_ /*17848*/;
assign _16039_ = D[37] ^ Q[23] /*17844*/;
assign _16036_ = _15436_ & _16039_ /*17840*/;
assign _16037_ = _15436_ ^ _16039_ /*17843*/;
assign _16038_ = _16030_ & _16037_ /*17841*/;
assign _16035_ = _16036_ | _16038_ /*17839*/;
assign _15822_ = _16030_ ^ _16037_ /*17842*/;
assign _16044_ = D[38] ^ Q[23] /*17838*/;
assign _16041_ = _15437_ & _16044_ /*17834*/;
assign _16042_ = _15437_ ^ _16044_ /*17837*/;
assign _16043_ = _16035_ & _16042_ /*17835*/;
assign _16040_ = _16041_ | _16043_ /*17833*/;
assign _15823_ = _16035_ ^ _16042_ /*17836*/;
assign _16049_ = D[39] ^ Q[23] /*17832*/;
assign _16046_ = _15438_ & _16049_ /*17828*/;
assign _16047_ = _15438_ ^ _16049_ /*17831*/;
assign _16048_ = _16040_ & _16047_ /*17829*/;
assign _16045_ = _16046_ | _16048_ /*17827*/;
assign _15824_ = _16040_ ^ _16047_ /*17830*/;
assign _16054_ = D[40] ^ Q[23] /*17826*/;
assign _16051_ = _15439_ & _16054_ /*17822*/;
assign _16052_ = _15439_ ^ _16054_ /*17825*/;
assign _16053_ = _16045_ & _16052_ /*17823*/;
assign _16050_ = _16051_ | _16053_ /*17821*/;
assign _15825_ = _16045_ ^ _16052_ /*17824*/;
assign _16059_ = D[41] ^ Q[23] /*17820*/;
assign _16056_ = _15440_ & _16059_ /*17816*/;
assign _16057_ = _15440_ ^ _16059_ /*17819*/;
assign _16058_ = _16050_ & _16057_ /*17817*/;
assign _16055_ = _16056_ | _16058_ /*17815*/;
assign _15826_ = _16050_ ^ _16057_ /*17818*/;
assign _16064_ = D[42] ^ Q[23] /*17814*/;
assign _16061_ = _15441_ & _16064_ /*17810*/;
assign _16062_ = _15441_ ^ _16064_ /*17813*/;
assign _16063_ = _16055_ & _16062_ /*17811*/;
assign _16060_ = _16061_ | _16063_ /*17809*/;
assign _15827_ = _16055_ ^ _16062_ /*17812*/;
assign _16069_ = D[43] ^ Q[23] /*17808*/;
assign _16066_ = _15442_ & _16069_ /*17804*/;
assign _16067_ = _15442_ ^ _16069_ /*17807*/;
assign _16068_ = _16060_ & _16067_ /*17805*/;
assign _16065_ = _16066_ | _16068_ /*17803*/;
assign _15828_ = _16060_ ^ _16067_ /*17806*/;
assign _16074_ = D[44] ^ Q[23] /*17802*/;
assign _16071_ = _15443_ & _16074_ /*17798*/;
assign _16072_ = _15443_ ^ _16074_ /*17801*/;
assign _16073_ = _16065_ & _16072_ /*17799*/;
assign _16070_ = _16071_ | _16073_ /*17797*/;
assign _15829_ = _16065_ ^ _16072_ /*17800*/;
assign _16079_ = D[45] ^ Q[23] /*17796*/;
assign _16076_ = _15444_ & _16079_ /*17792*/;
assign _16077_ = _15444_ ^ _16079_ /*17795*/;
assign _16078_ = _16070_ & _16077_ /*17793*/;
assign _16075_ = _16076_ | _16078_ /*17791*/;
assign _15830_ = _16070_ ^ _16077_ /*17794*/;
assign _16084_ = D[46] ^ Q[23] /*17790*/;
assign _16081_ = _15445_ & _16084_ /*17786*/;
assign _16082_ = _15445_ ^ _16084_ /*17789*/;
assign _16083_ = _16075_ & _16082_ /*17787*/;
assign _16080_ = _16081_ | _16083_ /*17785*/;
assign _15831_ = _16075_ ^ _16082_ /*17788*/;
assign _16089_ = D[47] ^ Q[23] /*17784*/;
assign _16086_ = _15446_ & _16089_ /*17780*/;
assign _16087_ = _15446_ ^ _16089_ /*17783*/;
assign _16088_ = _16080_ & _16087_ /*17781*/;
assign _16085_ = _16086_ | _16088_ /*17779*/;
assign _15832_ = _16080_ ^ _16087_ /*17782*/;
assign _16094_ = D[48] ^ Q[23] /*17778*/;
assign _16091_ = _15447_ & _16094_ /*17774*/;
assign _16092_ = _15447_ ^ _16094_ /*17777*/;
assign _16093_ = _16085_ & _16092_ /*17775*/;
assign _16090_ = _16091_ | _16093_ /*17773*/;
assign _15833_ = _16085_ ^ _16092_ /*17776*/;
assign _16099_ = D[49] ^ Q[23] /*17772*/;
assign _16096_ = _15448_ & _16099_ /*17768*/;
assign _16097_ = _15448_ ^ _16099_ /*17771*/;
assign _16098_ = _16090_ & _16097_ /*17769*/;
assign _16095_ = _16096_ | _16098_ /*17767*/;
assign _15834_ = _16090_ ^ _16097_ /*17770*/;
assign _16104_ = D[50] ^ Q[23] /*17766*/;
assign _16101_ = _15449_ & _16104_ /*17762*/;
assign _16102_ = _15449_ ^ _16104_ /*17765*/;
assign _16103_ = _16095_ & _16102_ /*17763*/;
assign _16100_ = _16101_ | _16103_ /*17761*/;
assign _15835_ = _16095_ ^ _16102_ /*17764*/;
assign _16109_ = D[51] ^ Q[23] /*17760*/;
assign _16106_ = _15450_ & _16109_ /*17756*/;
assign _16107_ = _15450_ ^ _16109_ /*17759*/;
assign _16108_ = _16100_ & _16107_ /*17757*/;
assign _16105_ = _16106_ | _16108_ /*17755*/;
assign _15836_ = _16100_ ^ _16107_ /*17758*/;
assign _16114_ = D[52] ^ Q[23] /*17754*/;
assign _16111_ = _15451_ & _16114_ /*17750*/;
assign _16112_ = _15451_ ^ _16114_ /*17753*/;
assign _16113_ = _16105_ & _16112_ /*17751*/;
assign _16110_ = _16111_ | _16113_ /*17749*/;
assign _15837_ = _16105_ ^ _16112_ /*17752*/;
assign _16119_ = D[53] ^ Q[23] /*17748*/;
assign _16116_ = _15452_ & _16119_ /*17744*/;
assign _16117_ = _15452_ ^ _16119_ /*17747*/;
assign _16118_ = _16110_ & _16117_ /*17745*/;
assign _16115_ = _16116_ | _16118_ /*17743*/;
assign _15838_ = _16110_ ^ _16117_ /*17746*/;
assign _16124_ = D[54] ^ Q[23] /*17742*/;
assign _16121_ = _15453_ & _16124_ /*17738*/;
assign _16122_ = _15453_ ^ _16124_ /*17741*/;
assign _16123_ = _16115_ & _16122_ /*17739*/;
assign _16120_ = _16121_ | _16123_ /*17737*/;
assign _15839_ = _16115_ ^ _16122_ /*17740*/;
assign _16129_ = D[55] ^ Q[23] /*17736*/;
assign _16126_ = _15454_ & _16129_ /*17732*/;
assign _16127_ = _15454_ ^ _16129_ /*17735*/;
assign _16128_ = _16120_ & _16127_ /*17733*/;
assign _16125_ = _16126_ | _16128_ /*17731*/;
assign _15840_ = _16120_ ^ _16127_ /*17734*/;
assign _16134_ = D[56] ^ Q[23] /*17730*/;
assign _16131_ = _15455_ & _16134_ /*17726*/;
assign _16132_ = _15455_ ^ _16134_ /*17729*/;
assign _16133_ = _16125_ & _16132_ /*17727*/;
assign _16130_ = _16131_ | _16133_ /*17725*/;
assign _15841_ = _16125_ ^ _16132_ /*17728*/;
assign _16139_ = D[57] ^ Q[23] /*17724*/;
assign _16136_ = _15456_ & _16139_ /*17720*/;
assign _16137_ = _15456_ ^ _16139_ /*17723*/;
assign _16138_ = _16130_ & _16137_ /*17721*/;
assign _16135_ = _16136_ | _16138_ /*17719*/;
assign _15842_ = _16130_ ^ _16137_ /*17722*/;
assign _16144_ = D[58] ^ Q[23] /*17718*/;
assign _16141_ = _15457_ & _16144_ /*17714*/;
assign _16142_ = _15457_ ^ _16144_ /*17717*/;
assign _16143_ = _16135_ & _16142_ /*17715*/;
assign _16140_ = _16141_ | _16143_ /*17713*/;
assign _15843_ = _16135_ ^ _16142_ /*17716*/;
assign _16149_ = D[59] ^ Q[23] /*17712*/;
assign _16146_ = _15458_ & _16149_ /*17708*/;
assign _16147_ = _15458_ ^ _16149_ /*17711*/;
assign _16148_ = _16140_ & _16147_ /*17709*/;
assign _16145_ = _16146_ | _16148_ /*17707*/;
assign _15844_ = _16140_ ^ _16147_ /*17710*/;
assign _16154_ = D[60] ^ Q[23] /*17706*/;
assign _16151_ = _15459_ & _16154_ /*17702*/;
assign _16152_ = _15459_ ^ _16154_ /*17705*/;
assign _16153_ = _16145_ & _16152_ /*17703*/;
assign _16150_ = _16151_ | _16153_ /*17701*/;
assign _15845_ = _16145_ ^ _16152_ /*17704*/;
assign _16159_ = D[61] ^ Q[23] /*17700*/;
assign _16156_ = _15460_ & _16159_ /*17696*/;
assign _16157_ = _15460_ ^ _16159_ /*17699*/;
assign _16158_ = _16150_ & _16157_ /*17697*/;
assign _16155_ = _16156_ | _16158_ /*17695*/;
assign _15846_ = _16150_ ^ _16157_ /*17698*/;
assign _16164_ = D[62] ^ Q[23] /*17694*/;
assign _16161_ = _15461_ & _16164_ /*17690*/;
assign _16162_ = _15461_ ^ _16164_ /*17693*/;
assign _16163_ = _16155_ & _16162_ /*17691*/;
assign _16160_ = _16161_ | _16163_ /*17689*/;
assign _15847_ = _16155_ ^ _16162_ /*17692*/;
assign _16168_ = zeroWire ^ Q[23] /*17688*/;
assign _16165_ = _15462_ & _16168_ /*17684*/;
assign _16166_ = _15462_ ^ _16168_ /*17687*/;
assign _16167_ = _16160_ & _16166_ /*17685*/;
assign Q[22] = _16165_ | _16167_ /*17683*/;
assign _15848_ = _16160_ ^ _16166_ /*17686*/;
assign _16239_ = D[0] ^ Q[22] /*17297*/;
assign _16236_ = R_0[21] & _16239_ /*17293*/;
assign _16237_ = R_0[21] ^ _16239_ /*17296*/;
assign _16238_ = Q[22] & _16237_ /*17294*/;
assign _16235_ = _16236_ | _16238_ /*17292*/;
assign _16170_ = Q[22] ^ _16237_ /*17295*/;
assign _16244_ = D[1] ^ Q[22] /*17291*/;
assign _16241_ = _15785_ & _16244_ /*17287*/;
assign _16242_ = _15785_ ^ _16244_ /*17290*/;
assign _16243_ = _16235_ & _16242_ /*17288*/;
assign _16240_ = _16241_ | _16243_ /*17286*/;
assign _16171_ = _16235_ ^ _16242_ /*17289*/;
assign _16249_ = D[2] ^ Q[22] /*17285*/;
assign _16246_ = _15786_ & _16249_ /*17281*/;
assign _16247_ = _15786_ ^ _16249_ /*17284*/;
assign _16248_ = _16240_ & _16247_ /*17282*/;
assign _16245_ = _16246_ | _16248_ /*17280*/;
assign _16172_ = _16240_ ^ _16247_ /*17283*/;
assign _16254_ = D[3] ^ Q[22] /*17279*/;
assign _16251_ = _15787_ & _16254_ /*17275*/;
assign _16252_ = _15787_ ^ _16254_ /*17278*/;
assign _16253_ = _16245_ & _16252_ /*17276*/;
assign _16250_ = _16251_ | _16253_ /*17274*/;
assign _16173_ = _16245_ ^ _16252_ /*17277*/;
assign _16259_ = D[4] ^ Q[22] /*17273*/;
assign _16256_ = _15788_ & _16259_ /*17269*/;
assign _16257_ = _15788_ ^ _16259_ /*17272*/;
assign _16258_ = _16250_ & _16257_ /*17270*/;
assign _16255_ = _16256_ | _16258_ /*17268*/;
assign _16174_ = _16250_ ^ _16257_ /*17271*/;
assign _16264_ = D[5] ^ Q[22] /*17267*/;
assign _16261_ = _15789_ & _16264_ /*17263*/;
assign _16262_ = _15789_ ^ _16264_ /*17266*/;
assign _16263_ = _16255_ & _16262_ /*17264*/;
assign _16260_ = _16261_ | _16263_ /*17262*/;
assign _16175_ = _16255_ ^ _16262_ /*17265*/;
assign _16269_ = D[6] ^ Q[22] /*17261*/;
assign _16266_ = _15790_ & _16269_ /*17257*/;
assign _16267_ = _15790_ ^ _16269_ /*17260*/;
assign _16268_ = _16260_ & _16267_ /*17258*/;
assign _16265_ = _16266_ | _16268_ /*17256*/;
assign _16176_ = _16260_ ^ _16267_ /*17259*/;
assign _16274_ = D[7] ^ Q[22] /*17255*/;
assign _16271_ = _15791_ & _16274_ /*17251*/;
assign _16272_ = _15791_ ^ _16274_ /*17254*/;
assign _16273_ = _16265_ & _16272_ /*17252*/;
assign _16270_ = _16271_ | _16273_ /*17250*/;
assign _16177_ = _16265_ ^ _16272_ /*17253*/;
assign _16279_ = D[8] ^ Q[22] /*17249*/;
assign _16276_ = _15792_ & _16279_ /*17245*/;
assign _16277_ = _15792_ ^ _16279_ /*17248*/;
assign _16278_ = _16270_ & _16277_ /*17246*/;
assign _16275_ = _16276_ | _16278_ /*17244*/;
assign _16178_ = _16270_ ^ _16277_ /*17247*/;
assign _16284_ = D[9] ^ Q[22] /*17243*/;
assign _16281_ = _15793_ & _16284_ /*17239*/;
assign _16282_ = _15793_ ^ _16284_ /*17242*/;
assign _16283_ = _16275_ & _16282_ /*17240*/;
assign _16280_ = _16281_ | _16283_ /*17238*/;
assign _16179_ = _16275_ ^ _16282_ /*17241*/;
assign _16289_ = D[10] ^ Q[22] /*17237*/;
assign _16286_ = _15794_ & _16289_ /*17233*/;
assign _16287_ = _15794_ ^ _16289_ /*17236*/;
assign _16288_ = _16280_ & _16287_ /*17234*/;
assign _16285_ = _16286_ | _16288_ /*17232*/;
assign _16180_ = _16280_ ^ _16287_ /*17235*/;
assign _16294_ = D[11] ^ Q[22] /*17231*/;
assign _16291_ = _15795_ & _16294_ /*17227*/;
assign _16292_ = _15795_ ^ _16294_ /*17230*/;
assign _16293_ = _16285_ & _16292_ /*17228*/;
assign _16290_ = _16291_ | _16293_ /*17226*/;
assign _16181_ = _16285_ ^ _16292_ /*17229*/;
assign _16299_ = D[12] ^ Q[22] /*17225*/;
assign _16296_ = _15796_ & _16299_ /*17221*/;
assign _16297_ = _15796_ ^ _16299_ /*17224*/;
assign _16298_ = _16290_ & _16297_ /*17222*/;
assign _16295_ = _16296_ | _16298_ /*17220*/;
assign _16182_ = _16290_ ^ _16297_ /*17223*/;
assign _16304_ = D[13] ^ Q[22] /*17219*/;
assign _16301_ = _15797_ & _16304_ /*17215*/;
assign _16302_ = _15797_ ^ _16304_ /*17218*/;
assign _16303_ = _16295_ & _16302_ /*17216*/;
assign _16300_ = _16301_ | _16303_ /*17214*/;
assign _16183_ = _16295_ ^ _16302_ /*17217*/;
assign _16309_ = D[14] ^ Q[22] /*17213*/;
assign _16306_ = _15798_ & _16309_ /*17209*/;
assign _16307_ = _15798_ ^ _16309_ /*17212*/;
assign _16308_ = _16300_ & _16307_ /*17210*/;
assign _16305_ = _16306_ | _16308_ /*17208*/;
assign _16184_ = _16300_ ^ _16307_ /*17211*/;
assign _16314_ = D[15] ^ Q[22] /*17207*/;
assign _16311_ = _15799_ & _16314_ /*17203*/;
assign _16312_ = _15799_ ^ _16314_ /*17206*/;
assign _16313_ = _16305_ & _16312_ /*17204*/;
assign _16310_ = _16311_ | _16313_ /*17202*/;
assign _16185_ = _16305_ ^ _16312_ /*17205*/;
assign _16319_ = D[16] ^ Q[22] /*17201*/;
assign _16316_ = _15800_ & _16319_ /*17197*/;
assign _16317_ = _15800_ ^ _16319_ /*17200*/;
assign _16318_ = _16310_ & _16317_ /*17198*/;
assign _16315_ = _16316_ | _16318_ /*17196*/;
assign _16186_ = _16310_ ^ _16317_ /*17199*/;
assign _16324_ = D[17] ^ Q[22] /*17195*/;
assign _16321_ = _15801_ & _16324_ /*17191*/;
assign _16322_ = _15801_ ^ _16324_ /*17194*/;
assign _16323_ = _16315_ & _16322_ /*17192*/;
assign _16320_ = _16321_ | _16323_ /*17190*/;
assign _16187_ = _16315_ ^ _16322_ /*17193*/;
assign _16329_ = D[18] ^ Q[22] /*17189*/;
assign _16326_ = _15802_ & _16329_ /*17185*/;
assign _16327_ = _15802_ ^ _16329_ /*17188*/;
assign _16328_ = _16320_ & _16327_ /*17186*/;
assign _16325_ = _16326_ | _16328_ /*17184*/;
assign _16188_ = _16320_ ^ _16327_ /*17187*/;
assign _16334_ = D[19] ^ Q[22] /*17183*/;
assign _16331_ = _15803_ & _16334_ /*17179*/;
assign _16332_ = _15803_ ^ _16334_ /*17182*/;
assign _16333_ = _16325_ & _16332_ /*17180*/;
assign _16330_ = _16331_ | _16333_ /*17178*/;
assign _16189_ = _16325_ ^ _16332_ /*17181*/;
assign _16339_ = D[20] ^ Q[22] /*17177*/;
assign _16336_ = _15804_ & _16339_ /*17173*/;
assign _16337_ = _15804_ ^ _16339_ /*17176*/;
assign _16338_ = _16330_ & _16337_ /*17174*/;
assign _16335_ = _16336_ | _16338_ /*17172*/;
assign _16190_ = _16330_ ^ _16337_ /*17175*/;
assign _16344_ = D[21] ^ Q[22] /*17171*/;
assign _16341_ = _15805_ & _16344_ /*17167*/;
assign _16342_ = _15805_ ^ _16344_ /*17170*/;
assign _16343_ = _16335_ & _16342_ /*17168*/;
assign _16340_ = _16341_ | _16343_ /*17166*/;
assign _16191_ = _16335_ ^ _16342_ /*17169*/;
assign _16349_ = D[22] ^ Q[22] /*17165*/;
assign _16346_ = _15806_ & _16349_ /*17161*/;
assign _16347_ = _15806_ ^ _16349_ /*17164*/;
assign _16348_ = _16340_ & _16347_ /*17162*/;
assign _16345_ = _16346_ | _16348_ /*17160*/;
assign _16192_ = _16340_ ^ _16347_ /*17163*/;
assign _16354_ = D[23] ^ Q[22] /*17159*/;
assign _16351_ = _15807_ & _16354_ /*17155*/;
assign _16352_ = _15807_ ^ _16354_ /*17158*/;
assign _16353_ = _16345_ & _16352_ /*17156*/;
assign _16350_ = _16351_ | _16353_ /*17154*/;
assign _16193_ = _16345_ ^ _16352_ /*17157*/;
assign _16359_ = D[24] ^ Q[22] /*17153*/;
assign _16356_ = _15808_ & _16359_ /*17149*/;
assign _16357_ = _15808_ ^ _16359_ /*17152*/;
assign _16358_ = _16350_ & _16357_ /*17150*/;
assign _16355_ = _16356_ | _16358_ /*17148*/;
assign _16194_ = _16350_ ^ _16357_ /*17151*/;
assign _16364_ = D[25] ^ Q[22] /*17147*/;
assign _16361_ = _15809_ & _16364_ /*17143*/;
assign _16362_ = _15809_ ^ _16364_ /*17146*/;
assign _16363_ = _16355_ & _16362_ /*17144*/;
assign _16360_ = _16361_ | _16363_ /*17142*/;
assign _16195_ = _16355_ ^ _16362_ /*17145*/;
assign _16369_ = D[26] ^ Q[22] /*17141*/;
assign _16366_ = _15810_ & _16369_ /*17137*/;
assign _16367_ = _15810_ ^ _16369_ /*17140*/;
assign _16368_ = _16360_ & _16367_ /*17138*/;
assign _16365_ = _16366_ | _16368_ /*17136*/;
assign _16196_ = _16360_ ^ _16367_ /*17139*/;
assign _16374_ = D[27] ^ Q[22] /*17135*/;
assign _16371_ = _15811_ & _16374_ /*17131*/;
assign _16372_ = _15811_ ^ _16374_ /*17134*/;
assign _16373_ = _16365_ & _16372_ /*17132*/;
assign _16370_ = _16371_ | _16373_ /*17130*/;
assign _16197_ = _16365_ ^ _16372_ /*17133*/;
assign _16379_ = D[28] ^ Q[22] /*17129*/;
assign _16376_ = _15812_ & _16379_ /*17125*/;
assign _16377_ = _15812_ ^ _16379_ /*17128*/;
assign _16378_ = _16370_ & _16377_ /*17126*/;
assign _16375_ = _16376_ | _16378_ /*17124*/;
assign _16198_ = _16370_ ^ _16377_ /*17127*/;
assign _16384_ = D[29] ^ Q[22] /*17123*/;
assign _16381_ = _15813_ & _16384_ /*17119*/;
assign _16382_ = _15813_ ^ _16384_ /*17122*/;
assign _16383_ = _16375_ & _16382_ /*17120*/;
assign _16380_ = _16381_ | _16383_ /*17118*/;
assign _16199_ = _16375_ ^ _16382_ /*17121*/;
assign _16389_ = D[30] ^ Q[22] /*17117*/;
assign _16386_ = _15814_ & _16389_ /*17113*/;
assign _16387_ = _15814_ ^ _16389_ /*17116*/;
assign _16388_ = _16380_ & _16387_ /*17114*/;
assign _16385_ = _16386_ | _16388_ /*17112*/;
assign _16200_ = _16380_ ^ _16387_ /*17115*/;
assign _16394_ = D[31] ^ Q[22] /*17111*/;
assign _16391_ = _15815_ & _16394_ /*17107*/;
assign _16392_ = _15815_ ^ _16394_ /*17110*/;
assign _16393_ = _16385_ & _16392_ /*17108*/;
assign _16390_ = _16391_ | _16393_ /*17106*/;
assign _16201_ = _16385_ ^ _16392_ /*17109*/;
assign _16399_ = D[32] ^ Q[22] /*17105*/;
assign _16396_ = _15816_ & _16399_ /*17101*/;
assign _16397_ = _15816_ ^ _16399_ /*17104*/;
assign _16398_ = _16390_ & _16397_ /*17102*/;
assign _16395_ = _16396_ | _16398_ /*17100*/;
assign _16202_ = _16390_ ^ _16397_ /*17103*/;
assign _16404_ = D[33] ^ Q[22] /*17099*/;
assign _16401_ = _15817_ & _16404_ /*17095*/;
assign _16402_ = _15817_ ^ _16404_ /*17098*/;
assign _16403_ = _16395_ & _16402_ /*17096*/;
assign _16400_ = _16401_ | _16403_ /*17094*/;
assign _16203_ = _16395_ ^ _16402_ /*17097*/;
assign _16409_ = D[34] ^ Q[22] /*17093*/;
assign _16406_ = _15818_ & _16409_ /*17089*/;
assign _16407_ = _15818_ ^ _16409_ /*17092*/;
assign _16408_ = _16400_ & _16407_ /*17090*/;
assign _16405_ = _16406_ | _16408_ /*17088*/;
assign _16204_ = _16400_ ^ _16407_ /*17091*/;
assign _16414_ = D[35] ^ Q[22] /*17087*/;
assign _16411_ = _15819_ & _16414_ /*17083*/;
assign _16412_ = _15819_ ^ _16414_ /*17086*/;
assign _16413_ = _16405_ & _16412_ /*17084*/;
assign _16410_ = _16411_ | _16413_ /*17082*/;
assign _16205_ = _16405_ ^ _16412_ /*17085*/;
assign _16419_ = D[36] ^ Q[22] /*17081*/;
assign _16416_ = _15820_ & _16419_ /*17077*/;
assign _16417_ = _15820_ ^ _16419_ /*17080*/;
assign _16418_ = _16410_ & _16417_ /*17078*/;
assign _16415_ = _16416_ | _16418_ /*17076*/;
assign _16206_ = _16410_ ^ _16417_ /*17079*/;
assign _16424_ = D[37] ^ Q[22] /*17075*/;
assign _16421_ = _15821_ & _16424_ /*17071*/;
assign _16422_ = _15821_ ^ _16424_ /*17074*/;
assign _16423_ = _16415_ & _16422_ /*17072*/;
assign _16420_ = _16421_ | _16423_ /*17070*/;
assign _16207_ = _16415_ ^ _16422_ /*17073*/;
assign _16429_ = D[38] ^ Q[22] /*17069*/;
assign _16426_ = _15822_ & _16429_ /*17065*/;
assign _16427_ = _15822_ ^ _16429_ /*17068*/;
assign _16428_ = _16420_ & _16427_ /*17066*/;
assign _16425_ = _16426_ | _16428_ /*17064*/;
assign _16208_ = _16420_ ^ _16427_ /*17067*/;
assign _16434_ = D[39] ^ Q[22] /*17063*/;
assign _16431_ = _15823_ & _16434_ /*17059*/;
assign _16432_ = _15823_ ^ _16434_ /*17062*/;
assign _16433_ = _16425_ & _16432_ /*17060*/;
assign _16430_ = _16431_ | _16433_ /*17058*/;
assign _16209_ = _16425_ ^ _16432_ /*17061*/;
assign _16439_ = D[40] ^ Q[22] /*17057*/;
assign _16436_ = _15824_ & _16439_ /*17053*/;
assign _16437_ = _15824_ ^ _16439_ /*17056*/;
assign _16438_ = _16430_ & _16437_ /*17054*/;
assign _16435_ = _16436_ | _16438_ /*17052*/;
assign _16210_ = _16430_ ^ _16437_ /*17055*/;
assign _16444_ = D[41] ^ Q[22] /*17051*/;
assign _16441_ = _15825_ & _16444_ /*17047*/;
assign _16442_ = _15825_ ^ _16444_ /*17050*/;
assign _16443_ = _16435_ & _16442_ /*17048*/;
assign _16440_ = _16441_ | _16443_ /*17046*/;
assign _16211_ = _16435_ ^ _16442_ /*17049*/;
assign _16449_ = D[42] ^ Q[22] /*17045*/;
assign _16446_ = _15826_ & _16449_ /*17041*/;
assign _16447_ = _15826_ ^ _16449_ /*17044*/;
assign _16448_ = _16440_ & _16447_ /*17042*/;
assign _16445_ = _16446_ | _16448_ /*17040*/;
assign _16212_ = _16440_ ^ _16447_ /*17043*/;
assign _16454_ = D[43] ^ Q[22] /*17039*/;
assign _16451_ = _15827_ & _16454_ /*17035*/;
assign _16452_ = _15827_ ^ _16454_ /*17038*/;
assign _16453_ = _16445_ & _16452_ /*17036*/;
assign _16450_ = _16451_ | _16453_ /*17034*/;
assign _16213_ = _16445_ ^ _16452_ /*17037*/;
assign _16459_ = D[44] ^ Q[22] /*17033*/;
assign _16456_ = _15828_ & _16459_ /*17029*/;
assign _16457_ = _15828_ ^ _16459_ /*17032*/;
assign _16458_ = _16450_ & _16457_ /*17030*/;
assign _16455_ = _16456_ | _16458_ /*17028*/;
assign _16214_ = _16450_ ^ _16457_ /*17031*/;
assign _16464_ = D[45] ^ Q[22] /*17027*/;
assign _16461_ = _15829_ & _16464_ /*17023*/;
assign _16462_ = _15829_ ^ _16464_ /*17026*/;
assign _16463_ = _16455_ & _16462_ /*17024*/;
assign _16460_ = _16461_ | _16463_ /*17022*/;
assign _16215_ = _16455_ ^ _16462_ /*17025*/;
assign _16469_ = D[46] ^ Q[22] /*17021*/;
assign _16466_ = _15830_ & _16469_ /*17017*/;
assign _16467_ = _15830_ ^ _16469_ /*17020*/;
assign _16468_ = _16460_ & _16467_ /*17018*/;
assign _16465_ = _16466_ | _16468_ /*17016*/;
assign _16216_ = _16460_ ^ _16467_ /*17019*/;
assign _16474_ = D[47] ^ Q[22] /*17015*/;
assign _16471_ = _15831_ & _16474_ /*17011*/;
assign _16472_ = _15831_ ^ _16474_ /*17014*/;
assign _16473_ = _16465_ & _16472_ /*17012*/;
assign _16470_ = _16471_ | _16473_ /*17010*/;
assign _16217_ = _16465_ ^ _16472_ /*17013*/;
assign _16479_ = D[48] ^ Q[22] /*17009*/;
assign _16476_ = _15832_ & _16479_ /*17005*/;
assign _16477_ = _15832_ ^ _16479_ /*17008*/;
assign _16478_ = _16470_ & _16477_ /*17006*/;
assign _16475_ = _16476_ | _16478_ /*17004*/;
assign _16218_ = _16470_ ^ _16477_ /*17007*/;
assign _16484_ = D[49] ^ Q[22] /*17003*/;
assign _16481_ = _15833_ & _16484_ /*16999*/;
assign _16482_ = _15833_ ^ _16484_ /*17002*/;
assign _16483_ = _16475_ & _16482_ /*17000*/;
assign _16480_ = _16481_ | _16483_ /*16998*/;
assign _16219_ = _16475_ ^ _16482_ /*17001*/;
assign _16489_ = D[50] ^ Q[22] /*16997*/;
assign _16486_ = _15834_ & _16489_ /*16993*/;
assign _16487_ = _15834_ ^ _16489_ /*16996*/;
assign _16488_ = _16480_ & _16487_ /*16994*/;
assign _16485_ = _16486_ | _16488_ /*16992*/;
assign _16220_ = _16480_ ^ _16487_ /*16995*/;
assign _16494_ = D[51] ^ Q[22] /*16991*/;
assign _16491_ = _15835_ & _16494_ /*16987*/;
assign _16492_ = _15835_ ^ _16494_ /*16990*/;
assign _16493_ = _16485_ & _16492_ /*16988*/;
assign _16490_ = _16491_ | _16493_ /*16986*/;
assign _16221_ = _16485_ ^ _16492_ /*16989*/;
assign _16499_ = D[52] ^ Q[22] /*16985*/;
assign _16496_ = _15836_ & _16499_ /*16981*/;
assign _16497_ = _15836_ ^ _16499_ /*16984*/;
assign _16498_ = _16490_ & _16497_ /*16982*/;
assign _16495_ = _16496_ | _16498_ /*16980*/;
assign _16222_ = _16490_ ^ _16497_ /*16983*/;
assign _16504_ = D[53] ^ Q[22] /*16979*/;
assign _16501_ = _15837_ & _16504_ /*16975*/;
assign _16502_ = _15837_ ^ _16504_ /*16978*/;
assign _16503_ = _16495_ & _16502_ /*16976*/;
assign _16500_ = _16501_ | _16503_ /*16974*/;
assign _16223_ = _16495_ ^ _16502_ /*16977*/;
assign _16509_ = D[54] ^ Q[22] /*16973*/;
assign _16506_ = _15838_ & _16509_ /*16969*/;
assign _16507_ = _15838_ ^ _16509_ /*16972*/;
assign _16508_ = _16500_ & _16507_ /*16970*/;
assign _16505_ = _16506_ | _16508_ /*16968*/;
assign _16224_ = _16500_ ^ _16507_ /*16971*/;
assign _16514_ = D[55] ^ Q[22] /*16967*/;
assign _16511_ = _15839_ & _16514_ /*16963*/;
assign _16512_ = _15839_ ^ _16514_ /*16966*/;
assign _16513_ = _16505_ & _16512_ /*16964*/;
assign _16510_ = _16511_ | _16513_ /*16962*/;
assign _16225_ = _16505_ ^ _16512_ /*16965*/;
assign _16519_ = D[56] ^ Q[22] /*16961*/;
assign _16516_ = _15840_ & _16519_ /*16957*/;
assign _16517_ = _15840_ ^ _16519_ /*16960*/;
assign _16518_ = _16510_ & _16517_ /*16958*/;
assign _16515_ = _16516_ | _16518_ /*16956*/;
assign _16226_ = _16510_ ^ _16517_ /*16959*/;
assign _16524_ = D[57] ^ Q[22] /*16955*/;
assign _16521_ = _15841_ & _16524_ /*16951*/;
assign _16522_ = _15841_ ^ _16524_ /*16954*/;
assign _16523_ = _16515_ & _16522_ /*16952*/;
assign _16520_ = _16521_ | _16523_ /*16950*/;
assign _16227_ = _16515_ ^ _16522_ /*16953*/;
assign _16529_ = D[58] ^ Q[22] /*16949*/;
assign _16526_ = _15842_ & _16529_ /*16945*/;
assign _16527_ = _15842_ ^ _16529_ /*16948*/;
assign _16528_ = _16520_ & _16527_ /*16946*/;
assign _16525_ = _16526_ | _16528_ /*16944*/;
assign _16228_ = _16520_ ^ _16527_ /*16947*/;
assign _16534_ = D[59] ^ Q[22] /*16943*/;
assign _16531_ = _15843_ & _16534_ /*16939*/;
assign _16532_ = _15843_ ^ _16534_ /*16942*/;
assign _16533_ = _16525_ & _16532_ /*16940*/;
assign _16530_ = _16531_ | _16533_ /*16938*/;
assign _16229_ = _16525_ ^ _16532_ /*16941*/;
assign _16539_ = D[60] ^ Q[22] /*16937*/;
assign _16536_ = _15844_ & _16539_ /*16933*/;
assign _16537_ = _15844_ ^ _16539_ /*16936*/;
assign _16538_ = _16530_ & _16537_ /*16934*/;
assign _16535_ = _16536_ | _16538_ /*16932*/;
assign _16230_ = _16530_ ^ _16537_ /*16935*/;
assign _16544_ = D[61] ^ Q[22] /*16931*/;
assign _16541_ = _15845_ & _16544_ /*16927*/;
assign _16542_ = _15845_ ^ _16544_ /*16930*/;
assign _16543_ = _16535_ & _16542_ /*16928*/;
assign _16540_ = _16541_ | _16543_ /*16926*/;
assign _16231_ = _16535_ ^ _16542_ /*16929*/;
assign _16549_ = D[62] ^ Q[22] /*16925*/;
assign _16546_ = _15846_ & _16549_ /*16921*/;
assign _16547_ = _15846_ ^ _16549_ /*16924*/;
assign _16548_ = _16540_ & _16547_ /*16922*/;
assign _16545_ = _16546_ | _16548_ /*16920*/;
assign _16232_ = _16540_ ^ _16547_ /*16923*/;
assign _16553_ = zeroWire ^ Q[22] /*16919*/;
assign _16550_ = _15847_ & _16553_ /*16915*/;
assign _16551_ = _15847_ ^ _16553_ /*16918*/;
assign _16552_ = _16545_ & _16551_ /*16916*/;
assign Q[21] = _16550_ | _16552_ /*16914*/;
assign _16233_ = _16545_ ^ _16551_ /*16917*/;
assign _16624_ = D[0] ^ Q[21] /*16528*/;
assign _16621_ = R_0[20] & _16624_ /*16524*/;
assign _16622_ = R_0[20] ^ _16624_ /*16527*/;
assign _16623_ = Q[21] & _16622_ /*16525*/;
assign _16620_ = _16621_ | _16623_ /*16523*/;
assign _16555_ = Q[21] ^ _16622_ /*16526*/;
assign _16629_ = D[1] ^ Q[21] /*16522*/;
assign _16626_ = _16170_ & _16629_ /*16518*/;
assign _16627_ = _16170_ ^ _16629_ /*16521*/;
assign _16628_ = _16620_ & _16627_ /*16519*/;
assign _16625_ = _16626_ | _16628_ /*16517*/;
assign _16556_ = _16620_ ^ _16627_ /*16520*/;
assign _16634_ = D[2] ^ Q[21] /*16516*/;
assign _16631_ = _16171_ & _16634_ /*16512*/;
assign _16632_ = _16171_ ^ _16634_ /*16515*/;
assign _16633_ = _16625_ & _16632_ /*16513*/;
assign _16630_ = _16631_ | _16633_ /*16511*/;
assign _16557_ = _16625_ ^ _16632_ /*16514*/;
assign _16639_ = D[3] ^ Q[21] /*16510*/;
assign _16636_ = _16172_ & _16639_ /*16506*/;
assign _16637_ = _16172_ ^ _16639_ /*16509*/;
assign _16638_ = _16630_ & _16637_ /*16507*/;
assign _16635_ = _16636_ | _16638_ /*16505*/;
assign _16558_ = _16630_ ^ _16637_ /*16508*/;
assign _16644_ = D[4] ^ Q[21] /*16504*/;
assign _16641_ = _16173_ & _16644_ /*16500*/;
assign _16642_ = _16173_ ^ _16644_ /*16503*/;
assign _16643_ = _16635_ & _16642_ /*16501*/;
assign _16640_ = _16641_ | _16643_ /*16499*/;
assign _16559_ = _16635_ ^ _16642_ /*16502*/;
assign _16649_ = D[5] ^ Q[21] /*16498*/;
assign _16646_ = _16174_ & _16649_ /*16494*/;
assign _16647_ = _16174_ ^ _16649_ /*16497*/;
assign _16648_ = _16640_ & _16647_ /*16495*/;
assign _16645_ = _16646_ | _16648_ /*16493*/;
assign _16560_ = _16640_ ^ _16647_ /*16496*/;
assign _16654_ = D[6] ^ Q[21] /*16492*/;
assign _16651_ = _16175_ & _16654_ /*16488*/;
assign _16652_ = _16175_ ^ _16654_ /*16491*/;
assign _16653_ = _16645_ & _16652_ /*16489*/;
assign _16650_ = _16651_ | _16653_ /*16487*/;
assign _16561_ = _16645_ ^ _16652_ /*16490*/;
assign _16659_ = D[7] ^ Q[21] /*16486*/;
assign _16656_ = _16176_ & _16659_ /*16482*/;
assign _16657_ = _16176_ ^ _16659_ /*16485*/;
assign _16658_ = _16650_ & _16657_ /*16483*/;
assign _16655_ = _16656_ | _16658_ /*16481*/;
assign _16562_ = _16650_ ^ _16657_ /*16484*/;
assign _16664_ = D[8] ^ Q[21] /*16480*/;
assign _16661_ = _16177_ & _16664_ /*16476*/;
assign _16662_ = _16177_ ^ _16664_ /*16479*/;
assign _16663_ = _16655_ & _16662_ /*16477*/;
assign _16660_ = _16661_ | _16663_ /*16475*/;
assign _16563_ = _16655_ ^ _16662_ /*16478*/;
assign _16669_ = D[9] ^ Q[21] /*16474*/;
assign _16666_ = _16178_ & _16669_ /*16470*/;
assign _16667_ = _16178_ ^ _16669_ /*16473*/;
assign _16668_ = _16660_ & _16667_ /*16471*/;
assign _16665_ = _16666_ | _16668_ /*16469*/;
assign _16564_ = _16660_ ^ _16667_ /*16472*/;
assign _16674_ = D[10] ^ Q[21] /*16468*/;
assign _16671_ = _16179_ & _16674_ /*16464*/;
assign _16672_ = _16179_ ^ _16674_ /*16467*/;
assign _16673_ = _16665_ & _16672_ /*16465*/;
assign _16670_ = _16671_ | _16673_ /*16463*/;
assign _16565_ = _16665_ ^ _16672_ /*16466*/;
assign _16679_ = D[11] ^ Q[21] /*16462*/;
assign _16676_ = _16180_ & _16679_ /*16458*/;
assign _16677_ = _16180_ ^ _16679_ /*16461*/;
assign _16678_ = _16670_ & _16677_ /*16459*/;
assign _16675_ = _16676_ | _16678_ /*16457*/;
assign _16566_ = _16670_ ^ _16677_ /*16460*/;
assign _16684_ = D[12] ^ Q[21] /*16456*/;
assign _16681_ = _16181_ & _16684_ /*16452*/;
assign _16682_ = _16181_ ^ _16684_ /*16455*/;
assign _16683_ = _16675_ & _16682_ /*16453*/;
assign _16680_ = _16681_ | _16683_ /*16451*/;
assign _16567_ = _16675_ ^ _16682_ /*16454*/;
assign _16689_ = D[13] ^ Q[21] /*16450*/;
assign _16686_ = _16182_ & _16689_ /*16446*/;
assign _16687_ = _16182_ ^ _16689_ /*16449*/;
assign _16688_ = _16680_ & _16687_ /*16447*/;
assign _16685_ = _16686_ | _16688_ /*16445*/;
assign _16568_ = _16680_ ^ _16687_ /*16448*/;
assign _16694_ = D[14] ^ Q[21] /*16444*/;
assign _16691_ = _16183_ & _16694_ /*16440*/;
assign _16692_ = _16183_ ^ _16694_ /*16443*/;
assign _16693_ = _16685_ & _16692_ /*16441*/;
assign _16690_ = _16691_ | _16693_ /*16439*/;
assign _16569_ = _16685_ ^ _16692_ /*16442*/;
assign _16699_ = D[15] ^ Q[21] /*16438*/;
assign _16696_ = _16184_ & _16699_ /*16434*/;
assign _16697_ = _16184_ ^ _16699_ /*16437*/;
assign _16698_ = _16690_ & _16697_ /*16435*/;
assign _16695_ = _16696_ | _16698_ /*16433*/;
assign _16570_ = _16690_ ^ _16697_ /*16436*/;
assign _16704_ = D[16] ^ Q[21] /*16432*/;
assign _16701_ = _16185_ & _16704_ /*16428*/;
assign _16702_ = _16185_ ^ _16704_ /*16431*/;
assign _16703_ = _16695_ & _16702_ /*16429*/;
assign _16700_ = _16701_ | _16703_ /*16427*/;
assign _16571_ = _16695_ ^ _16702_ /*16430*/;
assign _16709_ = D[17] ^ Q[21] /*16426*/;
assign _16706_ = _16186_ & _16709_ /*16422*/;
assign _16707_ = _16186_ ^ _16709_ /*16425*/;
assign _16708_ = _16700_ & _16707_ /*16423*/;
assign _16705_ = _16706_ | _16708_ /*16421*/;
assign _16572_ = _16700_ ^ _16707_ /*16424*/;
assign _16714_ = D[18] ^ Q[21] /*16420*/;
assign _16711_ = _16187_ & _16714_ /*16416*/;
assign _16712_ = _16187_ ^ _16714_ /*16419*/;
assign _16713_ = _16705_ & _16712_ /*16417*/;
assign _16710_ = _16711_ | _16713_ /*16415*/;
assign _16573_ = _16705_ ^ _16712_ /*16418*/;
assign _16719_ = D[19] ^ Q[21] /*16414*/;
assign _16716_ = _16188_ & _16719_ /*16410*/;
assign _16717_ = _16188_ ^ _16719_ /*16413*/;
assign _16718_ = _16710_ & _16717_ /*16411*/;
assign _16715_ = _16716_ | _16718_ /*16409*/;
assign _16574_ = _16710_ ^ _16717_ /*16412*/;
assign _16724_ = D[20] ^ Q[21] /*16408*/;
assign _16721_ = _16189_ & _16724_ /*16404*/;
assign _16722_ = _16189_ ^ _16724_ /*16407*/;
assign _16723_ = _16715_ & _16722_ /*16405*/;
assign _16720_ = _16721_ | _16723_ /*16403*/;
assign _16575_ = _16715_ ^ _16722_ /*16406*/;
assign _16729_ = D[21] ^ Q[21] /*16402*/;
assign _16726_ = _16190_ & _16729_ /*16398*/;
assign _16727_ = _16190_ ^ _16729_ /*16401*/;
assign _16728_ = _16720_ & _16727_ /*16399*/;
assign _16725_ = _16726_ | _16728_ /*16397*/;
assign _16576_ = _16720_ ^ _16727_ /*16400*/;
assign _16734_ = D[22] ^ Q[21] /*16396*/;
assign _16731_ = _16191_ & _16734_ /*16392*/;
assign _16732_ = _16191_ ^ _16734_ /*16395*/;
assign _16733_ = _16725_ & _16732_ /*16393*/;
assign _16730_ = _16731_ | _16733_ /*16391*/;
assign _16577_ = _16725_ ^ _16732_ /*16394*/;
assign _16739_ = D[23] ^ Q[21] /*16390*/;
assign _16736_ = _16192_ & _16739_ /*16386*/;
assign _16737_ = _16192_ ^ _16739_ /*16389*/;
assign _16738_ = _16730_ & _16737_ /*16387*/;
assign _16735_ = _16736_ | _16738_ /*16385*/;
assign _16578_ = _16730_ ^ _16737_ /*16388*/;
assign _16744_ = D[24] ^ Q[21] /*16384*/;
assign _16741_ = _16193_ & _16744_ /*16380*/;
assign _16742_ = _16193_ ^ _16744_ /*16383*/;
assign _16743_ = _16735_ & _16742_ /*16381*/;
assign _16740_ = _16741_ | _16743_ /*16379*/;
assign _16579_ = _16735_ ^ _16742_ /*16382*/;
assign _16749_ = D[25] ^ Q[21] /*16378*/;
assign _16746_ = _16194_ & _16749_ /*16374*/;
assign _16747_ = _16194_ ^ _16749_ /*16377*/;
assign _16748_ = _16740_ & _16747_ /*16375*/;
assign _16745_ = _16746_ | _16748_ /*16373*/;
assign _16580_ = _16740_ ^ _16747_ /*16376*/;
assign _16754_ = D[26] ^ Q[21] /*16372*/;
assign _16751_ = _16195_ & _16754_ /*16368*/;
assign _16752_ = _16195_ ^ _16754_ /*16371*/;
assign _16753_ = _16745_ & _16752_ /*16369*/;
assign _16750_ = _16751_ | _16753_ /*16367*/;
assign _16581_ = _16745_ ^ _16752_ /*16370*/;
assign _16759_ = D[27] ^ Q[21] /*16366*/;
assign _16756_ = _16196_ & _16759_ /*16362*/;
assign _16757_ = _16196_ ^ _16759_ /*16365*/;
assign _16758_ = _16750_ & _16757_ /*16363*/;
assign _16755_ = _16756_ | _16758_ /*16361*/;
assign _16582_ = _16750_ ^ _16757_ /*16364*/;
assign _16764_ = D[28] ^ Q[21] /*16360*/;
assign _16761_ = _16197_ & _16764_ /*16356*/;
assign _16762_ = _16197_ ^ _16764_ /*16359*/;
assign _16763_ = _16755_ & _16762_ /*16357*/;
assign _16760_ = _16761_ | _16763_ /*16355*/;
assign _16583_ = _16755_ ^ _16762_ /*16358*/;
assign _16769_ = D[29] ^ Q[21] /*16354*/;
assign _16766_ = _16198_ & _16769_ /*16350*/;
assign _16767_ = _16198_ ^ _16769_ /*16353*/;
assign _16768_ = _16760_ & _16767_ /*16351*/;
assign _16765_ = _16766_ | _16768_ /*16349*/;
assign _16584_ = _16760_ ^ _16767_ /*16352*/;
assign _16774_ = D[30] ^ Q[21] /*16348*/;
assign _16771_ = _16199_ & _16774_ /*16344*/;
assign _16772_ = _16199_ ^ _16774_ /*16347*/;
assign _16773_ = _16765_ & _16772_ /*16345*/;
assign _16770_ = _16771_ | _16773_ /*16343*/;
assign _16585_ = _16765_ ^ _16772_ /*16346*/;
assign _16779_ = D[31] ^ Q[21] /*16342*/;
assign _16776_ = _16200_ & _16779_ /*16338*/;
assign _16777_ = _16200_ ^ _16779_ /*16341*/;
assign _16778_ = _16770_ & _16777_ /*16339*/;
assign _16775_ = _16776_ | _16778_ /*16337*/;
assign _16586_ = _16770_ ^ _16777_ /*16340*/;
assign _16784_ = D[32] ^ Q[21] /*16336*/;
assign _16781_ = _16201_ & _16784_ /*16332*/;
assign _16782_ = _16201_ ^ _16784_ /*16335*/;
assign _16783_ = _16775_ & _16782_ /*16333*/;
assign _16780_ = _16781_ | _16783_ /*16331*/;
assign _16587_ = _16775_ ^ _16782_ /*16334*/;
assign _16789_ = D[33] ^ Q[21] /*16330*/;
assign _16786_ = _16202_ & _16789_ /*16326*/;
assign _16787_ = _16202_ ^ _16789_ /*16329*/;
assign _16788_ = _16780_ & _16787_ /*16327*/;
assign _16785_ = _16786_ | _16788_ /*16325*/;
assign _16588_ = _16780_ ^ _16787_ /*16328*/;
assign _16794_ = D[34] ^ Q[21] /*16324*/;
assign _16791_ = _16203_ & _16794_ /*16320*/;
assign _16792_ = _16203_ ^ _16794_ /*16323*/;
assign _16793_ = _16785_ & _16792_ /*16321*/;
assign _16790_ = _16791_ | _16793_ /*16319*/;
assign _16589_ = _16785_ ^ _16792_ /*16322*/;
assign _16799_ = D[35] ^ Q[21] /*16318*/;
assign _16796_ = _16204_ & _16799_ /*16314*/;
assign _16797_ = _16204_ ^ _16799_ /*16317*/;
assign _16798_ = _16790_ & _16797_ /*16315*/;
assign _16795_ = _16796_ | _16798_ /*16313*/;
assign _16590_ = _16790_ ^ _16797_ /*16316*/;
assign _16804_ = D[36] ^ Q[21] /*16312*/;
assign _16801_ = _16205_ & _16804_ /*16308*/;
assign _16802_ = _16205_ ^ _16804_ /*16311*/;
assign _16803_ = _16795_ & _16802_ /*16309*/;
assign _16800_ = _16801_ | _16803_ /*16307*/;
assign _16591_ = _16795_ ^ _16802_ /*16310*/;
assign _16809_ = D[37] ^ Q[21] /*16306*/;
assign _16806_ = _16206_ & _16809_ /*16302*/;
assign _16807_ = _16206_ ^ _16809_ /*16305*/;
assign _16808_ = _16800_ & _16807_ /*16303*/;
assign _16805_ = _16806_ | _16808_ /*16301*/;
assign _16592_ = _16800_ ^ _16807_ /*16304*/;
assign _16814_ = D[38] ^ Q[21] /*16300*/;
assign _16811_ = _16207_ & _16814_ /*16296*/;
assign _16812_ = _16207_ ^ _16814_ /*16299*/;
assign _16813_ = _16805_ & _16812_ /*16297*/;
assign _16810_ = _16811_ | _16813_ /*16295*/;
assign _16593_ = _16805_ ^ _16812_ /*16298*/;
assign _16819_ = D[39] ^ Q[21] /*16294*/;
assign _16816_ = _16208_ & _16819_ /*16290*/;
assign _16817_ = _16208_ ^ _16819_ /*16293*/;
assign _16818_ = _16810_ & _16817_ /*16291*/;
assign _16815_ = _16816_ | _16818_ /*16289*/;
assign _16594_ = _16810_ ^ _16817_ /*16292*/;
assign _16824_ = D[40] ^ Q[21] /*16288*/;
assign _16821_ = _16209_ & _16824_ /*16284*/;
assign _16822_ = _16209_ ^ _16824_ /*16287*/;
assign _16823_ = _16815_ & _16822_ /*16285*/;
assign _16820_ = _16821_ | _16823_ /*16283*/;
assign _16595_ = _16815_ ^ _16822_ /*16286*/;
assign _16829_ = D[41] ^ Q[21] /*16282*/;
assign _16826_ = _16210_ & _16829_ /*16278*/;
assign _16827_ = _16210_ ^ _16829_ /*16281*/;
assign _16828_ = _16820_ & _16827_ /*16279*/;
assign _16825_ = _16826_ | _16828_ /*16277*/;
assign _16596_ = _16820_ ^ _16827_ /*16280*/;
assign _16834_ = D[42] ^ Q[21] /*16276*/;
assign _16831_ = _16211_ & _16834_ /*16272*/;
assign _16832_ = _16211_ ^ _16834_ /*16275*/;
assign _16833_ = _16825_ & _16832_ /*16273*/;
assign _16830_ = _16831_ | _16833_ /*16271*/;
assign _16597_ = _16825_ ^ _16832_ /*16274*/;
assign _16839_ = D[43] ^ Q[21] /*16270*/;
assign _16836_ = _16212_ & _16839_ /*16266*/;
assign _16837_ = _16212_ ^ _16839_ /*16269*/;
assign _16838_ = _16830_ & _16837_ /*16267*/;
assign _16835_ = _16836_ | _16838_ /*16265*/;
assign _16598_ = _16830_ ^ _16837_ /*16268*/;
assign _16844_ = D[44] ^ Q[21] /*16264*/;
assign _16841_ = _16213_ & _16844_ /*16260*/;
assign _16842_ = _16213_ ^ _16844_ /*16263*/;
assign _16843_ = _16835_ & _16842_ /*16261*/;
assign _16840_ = _16841_ | _16843_ /*16259*/;
assign _16599_ = _16835_ ^ _16842_ /*16262*/;
assign _16849_ = D[45] ^ Q[21] /*16258*/;
assign _16846_ = _16214_ & _16849_ /*16254*/;
assign _16847_ = _16214_ ^ _16849_ /*16257*/;
assign _16848_ = _16840_ & _16847_ /*16255*/;
assign _16845_ = _16846_ | _16848_ /*16253*/;
assign _16600_ = _16840_ ^ _16847_ /*16256*/;
assign _16854_ = D[46] ^ Q[21] /*16252*/;
assign _16851_ = _16215_ & _16854_ /*16248*/;
assign _16852_ = _16215_ ^ _16854_ /*16251*/;
assign _16853_ = _16845_ & _16852_ /*16249*/;
assign _16850_ = _16851_ | _16853_ /*16247*/;
assign _16601_ = _16845_ ^ _16852_ /*16250*/;
assign _16859_ = D[47] ^ Q[21] /*16246*/;
assign _16856_ = _16216_ & _16859_ /*16242*/;
assign _16857_ = _16216_ ^ _16859_ /*16245*/;
assign _16858_ = _16850_ & _16857_ /*16243*/;
assign _16855_ = _16856_ | _16858_ /*16241*/;
assign _16602_ = _16850_ ^ _16857_ /*16244*/;
assign _16864_ = D[48] ^ Q[21] /*16240*/;
assign _16861_ = _16217_ & _16864_ /*16236*/;
assign _16862_ = _16217_ ^ _16864_ /*16239*/;
assign _16863_ = _16855_ & _16862_ /*16237*/;
assign _16860_ = _16861_ | _16863_ /*16235*/;
assign _16603_ = _16855_ ^ _16862_ /*16238*/;
assign _16869_ = D[49] ^ Q[21] /*16234*/;
assign _16866_ = _16218_ & _16869_ /*16230*/;
assign _16867_ = _16218_ ^ _16869_ /*16233*/;
assign _16868_ = _16860_ & _16867_ /*16231*/;
assign _16865_ = _16866_ | _16868_ /*16229*/;
assign _16604_ = _16860_ ^ _16867_ /*16232*/;
assign _16874_ = D[50] ^ Q[21] /*16228*/;
assign _16871_ = _16219_ & _16874_ /*16224*/;
assign _16872_ = _16219_ ^ _16874_ /*16227*/;
assign _16873_ = _16865_ & _16872_ /*16225*/;
assign _16870_ = _16871_ | _16873_ /*16223*/;
assign _16605_ = _16865_ ^ _16872_ /*16226*/;
assign _16879_ = D[51] ^ Q[21] /*16222*/;
assign _16876_ = _16220_ & _16879_ /*16218*/;
assign _16877_ = _16220_ ^ _16879_ /*16221*/;
assign _16878_ = _16870_ & _16877_ /*16219*/;
assign _16875_ = _16876_ | _16878_ /*16217*/;
assign _16606_ = _16870_ ^ _16877_ /*16220*/;
assign _16884_ = D[52] ^ Q[21] /*16216*/;
assign _16881_ = _16221_ & _16884_ /*16212*/;
assign _16882_ = _16221_ ^ _16884_ /*16215*/;
assign _16883_ = _16875_ & _16882_ /*16213*/;
assign _16880_ = _16881_ | _16883_ /*16211*/;
assign _16607_ = _16875_ ^ _16882_ /*16214*/;
assign _16889_ = D[53] ^ Q[21] /*16210*/;
assign _16886_ = _16222_ & _16889_ /*16206*/;
assign _16887_ = _16222_ ^ _16889_ /*16209*/;
assign _16888_ = _16880_ & _16887_ /*16207*/;
assign _16885_ = _16886_ | _16888_ /*16205*/;
assign _16608_ = _16880_ ^ _16887_ /*16208*/;
assign _16894_ = D[54] ^ Q[21] /*16204*/;
assign _16891_ = _16223_ & _16894_ /*16200*/;
assign _16892_ = _16223_ ^ _16894_ /*16203*/;
assign _16893_ = _16885_ & _16892_ /*16201*/;
assign _16890_ = _16891_ | _16893_ /*16199*/;
assign _16609_ = _16885_ ^ _16892_ /*16202*/;
assign _16899_ = D[55] ^ Q[21] /*16198*/;
assign _16896_ = _16224_ & _16899_ /*16194*/;
assign _16897_ = _16224_ ^ _16899_ /*16197*/;
assign _16898_ = _16890_ & _16897_ /*16195*/;
assign _16895_ = _16896_ | _16898_ /*16193*/;
assign _16610_ = _16890_ ^ _16897_ /*16196*/;
assign _16904_ = D[56] ^ Q[21] /*16192*/;
assign _16901_ = _16225_ & _16904_ /*16188*/;
assign _16902_ = _16225_ ^ _16904_ /*16191*/;
assign _16903_ = _16895_ & _16902_ /*16189*/;
assign _16900_ = _16901_ | _16903_ /*16187*/;
assign _16611_ = _16895_ ^ _16902_ /*16190*/;
assign _16909_ = D[57] ^ Q[21] /*16186*/;
assign _16906_ = _16226_ & _16909_ /*16182*/;
assign _16907_ = _16226_ ^ _16909_ /*16185*/;
assign _16908_ = _16900_ & _16907_ /*16183*/;
assign _16905_ = _16906_ | _16908_ /*16181*/;
assign _16612_ = _16900_ ^ _16907_ /*16184*/;
assign _16914_ = D[58] ^ Q[21] /*16180*/;
assign _16911_ = _16227_ & _16914_ /*16176*/;
assign _16912_ = _16227_ ^ _16914_ /*16179*/;
assign _16913_ = _16905_ & _16912_ /*16177*/;
assign _16910_ = _16911_ | _16913_ /*16175*/;
assign _16613_ = _16905_ ^ _16912_ /*16178*/;
assign _16919_ = D[59] ^ Q[21] /*16174*/;
assign _16916_ = _16228_ & _16919_ /*16170*/;
assign _16917_ = _16228_ ^ _16919_ /*16173*/;
assign _16918_ = _16910_ & _16917_ /*16171*/;
assign _16915_ = _16916_ | _16918_ /*16169*/;
assign _16614_ = _16910_ ^ _16917_ /*16172*/;
assign _16924_ = D[60] ^ Q[21] /*16168*/;
assign _16921_ = _16229_ & _16924_ /*16164*/;
assign _16922_ = _16229_ ^ _16924_ /*16167*/;
assign _16923_ = _16915_ & _16922_ /*16165*/;
assign _16920_ = _16921_ | _16923_ /*16163*/;
assign _16615_ = _16915_ ^ _16922_ /*16166*/;
assign _16929_ = D[61] ^ Q[21] /*16162*/;
assign _16926_ = _16230_ & _16929_ /*16158*/;
assign _16927_ = _16230_ ^ _16929_ /*16161*/;
assign _16928_ = _16920_ & _16927_ /*16159*/;
assign _16925_ = _16926_ | _16928_ /*16157*/;
assign _16616_ = _16920_ ^ _16927_ /*16160*/;
assign _16934_ = D[62] ^ Q[21] /*16156*/;
assign _16931_ = _16231_ & _16934_ /*16152*/;
assign _16932_ = _16231_ ^ _16934_ /*16155*/;
assign _16933_ = _16925_ & _16932_ /*16153*/;
assign _16930_ = _16931_ | _16933_ /*16151*/;
assign _16617_ = _16925_ ^ _16932_ /*16154*/;
assign _16938_ = zeroWire ^ Q[21] /*16150*/;
assign _16935_ = _16232_ & _16938_ /*16146*/;
assign _16936_ = _16232_ ^ _16938_ /*16149*/;
assign _16937_ = _16930_ & _16936_ /*16147*/;
assign Q[20] = _16935_ | _16937_ /*16145*/;
assign _16618_ = _16930_ ^ _16936_ /*16148*/;
assign _17009_ = D[0] ^ Q[20] /*15759*/;
assign _17006_ = R_0[19] & _17009_ /*15755*/;
assign _17007_ = R_0[19] ^ _17009_ /*15758*/;
assign _17008_ = Q[20] & _17007_ /*15756*/;
assign _17005_ = _17006_ | _17008_ /*15754*/;
assign _16940_ = Q[20] ^ _17007_ /*15757*/;
assign _17014_ = D[1] ^ Q[20] /*15753*/;
assign _17011_ = _16555_ & _17014_ /*15749*/;
assign _17012_ = _16555_ ^ _17014_ /*15752*/;
assign _17013_ = _17005_ & _17012_ /*15750*/;
assign _17010_ = _17011_ | _17013_ /*15748*/;
assign _16941_ = _17005_ ^ _17012_ /*15751*/;
assign _17019_ = D[2] ^ Q[20] /*15747*/;
assign _17016_ = _16556_ & _17019_ /*15743*/;
assign _17017_ = _16556_ ^ _17019_ /*15746*/;
assign _17018_ = _17010_ & _17017_ /*15744*/;
assign _17015_ = _17016_ | _17018_ /*15742*/;
assign _16942_ = _17010_ ^ _17017_ /*15745*/;
assign _17024_ = D[3] ^ Q[20] /*15741*/;
assign _17021_ = _16557_ & _17024_ /*15737*/;
assign _17022_ = _16557_ ^ _17024_ /*15740*/;
assign _17023_ = _17015_ & _17022_ /*15738*/;
assign _17020_ = _17021_ | _17023_ /*15736*/;
assign _16943_ = _17015_ ^ _17022_ /*15739*/;
assign _17029_ = D[4] ^ Q[20] /*15735*/;
assign _17026_ = _16558_ & _17029_ /*15731*/;
assign _17027_ = _16558_ ^ _17029_ /*15734*/;
assign _17028_ = _17020_ & _17027_ /*15732*/;
assign _17025_ = _17026_ | _17028_ /*15730*/;
assign _16944_ = _17020_ ^ _17027_ /*15733*/;
assign _17034_ = D[5] ^ Q[20] /*15729*/;
assign _17031_ = _16559_ & _17034_ /*15725*/;
assign _17032_ = _16559_ ^ _17034_ /*15728*/;
assign _17033_ = _17025_ & _17032_ /*15726*/;
assign _17030_ = _17031_ | _17033_ /*15724*/;
assign _16945_ = _17025_ ^ _17032_ /*15727*/;
assign _17039_ = D[6] ^ Q[20] /*15723*/;
assign _17036_ = _16560_ & _17039_ /*15719*/;
assign _17037_ = _16560_ ^ _17039_ /*15722*/;
assign _17038_ = _17030_ & _17037_ /*15720*/;
assign _17035_ = _17036_ | _17038_ /*15718*/;
assign _16946_ = _17030_ ^ _17037_ /*15721*/;
assign _17044_ = D[7] ^ Q[20] /*15717*/;
assign _17041_ = _16561_ & _17044_ /*15713*/;
assign _17042_ = _16561_ ^ _17044_ /*15716*/;
assign _17043_ = _17035_ & _17042_ /*15714*/;
assign _17040_ = _17041_ | _17043_ /*15712*/;
assign _16947_ = _17035_ ^ _17042_ /*15715*/;
assign _17049_ = D[8] ^ Q[20] /*15711*/;
assign _17046_ = _16562_ & _17049_ /*15707*/;
assign _17047_ = _16562_ ^ _17049_ /*15710*/;
assign _17048_ = _17040_ & _17047_ /*15708*/;
assign _17045_ = _17046_ | _17048_ /*15706*/;
assign _16948_ = _17040_ ^ _17047_ /*15709*/;
assign _17054_ = D[9] ^ Q[20] /*15705*/;
assign _17051_ = _16563_ & _17054_ /*15701*/;
assign _17052_ = _16563_ ^ _17054_ /*15704*/;
assign _17053_ = _17045_ & _17052_ /*15702*/;
assign _17050_ = _17051_ | _17053_ /*15700*/;
assign _16949_ = _17045_ ^ _17052_ /*15703*/;
assign _17059_ = D[10] ^ Q[20] /*15699*/;
assign _17056_ = _16564_ & _17059_ /*15695*/;
assign _17057_ = _16564_ ^ _17059_ /*15698*/;
assign _17058_ = _17050_ & _17057_ /*15696*/;
assign _17055_ = _17056_ | _17058_ /*15694*/;
assign _16950_ = _17050_ ^ _17057_ /*15697*/;
assign _17064_ = D[11] ^ Q[20] /*15693*/;
assign _17061_ = _16565_ & _17064_ /*15689*/;
assign _17062_ = _16565_ ^ _17064_ /*15692*/;
assign _17063_ = _17055_ & _17062_ /*15690*/;
assign _17060_ = _17061_ | _17063_ /*15688*/;
assign _16951_ = _17055_ ^ _17062_ /*15691*/;
assign _17069_ = D[12] ^ Q[20] /*15687*/;
assign _17066_ = _16566_ & _17069_ /*15683*/;
assign _17067_ = _16566_ ^ _17069_ /*15686*/;
assign _17068_ = _17060_ & _17067_ /*15684*/;
assign _17065_ = _17066_ | _17068_ /*15682*/;
assign _16952_ = _17060_ ^ _17067_ /*15685*/;
assign _17074_ = D[13] ^ Q[20] /*15681*/;
assign _17071_ = _16567_ & _17074_ /*15677*/;
assign _17072_ = _16567_ ^ _17074_ /*15680*/;
assign _17073_ = _17065_ & _17072_ /*15678*/;
assign _17070_ = _17071_ | _17073_ /*15676*/;
assign _16953_ = _17065_ ^ _17072_ /*15679*/;
assign _17079_ = D[14] ^ Q[20] /*15675*/;
assign _17076_ = _16568_ & _17079_ /*15671*/;
assign _17077_ = _16568_ ^ _17079_ /*15674*/;
assign _17078_ = _17070_ & _17077_ /*15672*/;
assign _17075_ = _17076_ | _17078_ /*15670*/;
assign _16954_ = _17070_ ^ _17077_ /*15673*/;
assign _17084_ = D[15] ^ Q[20] /*15669*/;
assign _17081_ = _16569_ & _17084_ /*15665*/;
assign _17082_ = _16569_ ^ _17084_ /*15668*/;
assign _17083_ = _17075_ & _17082_ /*15666*/;
assign _17080_ = _17081_ | _17083_ /*15664*/;
assign _16955_ = _17075_ ^ _17082_ /*15667*/;
assign _17089_ = D[16] ^ Q[20] /*15663*/;
assign _17086_ = _16570_ & _17089_ /*15659*/;
assign _17087_ = _16570_ ^ _17089_ /*15662*/;
assign _17088_ = _17080_ & _17087_ /*15660*/;
assign _17085_ = _17086_ | _17088_ /*15658*/;
assign _16956_ = _17080_ ^ _17087_ /*15661*/;
assign _17094_ = D[17] ^ Q[20] /*15657*/;
assign _17091_ = _16571_ & _17094_ /*15653*/;
assign _17092_ = _16571_ ^ _17094_ /*15656*/;
assign _17093_ = _17085_ & _17092_ /*15654*/;
assign _17090_ = _17091_ | _17093_ /*15652*/;
assign _16957_ = _17085_ ^ _17092_ /*15655*/;
assign _17099_ = D[18] ^ Q[20] /*15651*/;
assign _17096_ = _16572_ & _17099_ /*15647*/;
assign _17097_ = _16572_ ^ _17099_ /*15650*/;
assign _17098_ = _17090_ & _17097_ /*15648*/;
assign _17095_ = _17096_ | _17098_ /*15646*/;
assign _16958_ = _17090_ ^ _17097_ /*15649*/;
assign _17104_ = D[19] ^ Q[20] /*15645*/;
assign _17101_ = _16573_ & _17104_ /*15641*/;
assign _17102_ = _16573_ ^ _17104_ /*15644*/;
assign _17103_ = _17095_ & _17102_ /*15642*/;
assign _17100_ = _17101_ | _17103_ /*15640*/;
assign _16959_ = _17095_ ^ _17102_ /*15643*/;
assign _17109_ = D[20] ^ Q[20] /*15639*/;
assign _17106_ = _16574_ & _17109_ /*15635*/;
assign _17107_ = _16574_ ^ _17109_ /*15638*/;
assign _17108_ = _17100_ & _17107_ /*15636*/;
assign _17105_ = _17106_ | _17108_ /*15634*/;
assign _16960_ = _17100_ ^ _17107_ /*15637*/;
assign _17114_ = D[21] ^ Q[20] /*15633*/;
assign _17111_ = _16575_ & _17114_ /*15629*/;
assign _17112_ = _16575_ ^ _17114_ /*15632*/;
assign _17113_ = _17105_ & _17112_ /*15630*/;
assign _17110_ = _17111_ | _17113_ /*15628*/;
assign _16961_ = _17105_ ^ _17112_ /*15631*/;
assign _17119_ = D[22] ^ Q[20] /*15627*/;
assign _17116_ = _16576_ & _17119_ /*15623*/;
assign _17117_ = _16576_ ^ _17119_ /*15626*/;
assign _17118_ = _17110_ & _17117_ /*15624*/;
assign _17115_ = _17116_ | _17118_ /*15622*/;
assign _16962_ = _17110_ ^ _17117_ /*15625*/;
assign _17124_ = D[23] ^ Q[20] /*15621*/;
assign _17121_ = _16577_ & _17124_ /*15617*/;
assign _17122_ = _16577_ ^ _17124_ /*15620*/;
assign _17123_ = _17115_ & _17122_ /*15618*/;
assign _17120_ = _17121_ | _17123_ /*15616*/;
assign _16963_ = _17115_ ^ _17122_ /*15619*/;
assign _17129_ = D[24] ^ Q[20] /*15615*/;
assign _17126_ = _16578_ & _17129_ /*15611*/;
assign _17127_ = _16578_ ^ _17129_ /*15614*/;
assign _17128_ = _17120_ & _17127_ /*15612*/;
assign _17125_ = _17126_ | _17128_ /*15610*/;
assign _16964_ = _17120_ ^ _17127_ /*15613*/;
assign _17134_ = D[25] ^ Q[20] /*15609*/;
assign _17131_ = _16579_ & _17134_ /*15605*/;
assign _17132_ = _16579_ ^ _17134_ /*15608*/;
assign _17133_ = _17125_ & _17132_ /*15606*/;
assign _17130_ = _17131_ | _17133_ /*15604*/;
assign _16965_ = _17125_ ^ _17132_ /*15607*/;
assign _17139_ = D[26] ^ Q[20] /*15603*/;
assign _17136_ = _16580_ & _17139_ /*15599*/;
assign _17137_ = _16580_ ^ _17139_ /*15602*/;
assign _17138_ = _17130_ & _17137_ /*15600*/;
assign _17135_ = _17136_ | _17138_ /*15598*/;
assign _16966_ = _17130_ ^ _17137_ /*15601*/;
assign _17144_ = D[27] ^ Q[20] /*15597*/;
assign _17141_ = _16581_ & _17144_ /*15593*/;
assign _17142_ = _16581_ ^ _17144_ /*15596*/;
assign _17143_ = _17135_ & _17142_ /*15594*/;
assign _17140_ = _17141_ | _17143_ /*15592*/;
assign _16967_ = _17135_ ^ _17142_ /*15595*/;
assign _17149_ = D[28] ^ Q[20] /*15591*/;
assign _17146_ = _16582_ & _17149_ /*15587*/;
assign _17147_ = _16582_ ^ _17149_ /*15590*/;
assign _17148_ = _17140_ & _17147_ /*15588*/;
assign _17145_ = _17146_ | _17148_ /*15586*/;
assign _16968_ = _17140_ ^ _17147_ /*15589*/;
assign _17154_ = D[29] ^ Q[20] /*15585*/;
assign _17151_ = _16583_ & _17154_ /*15581*/;
assign _17152_ = _16583_ ^ _17154_ /*15584*/;
assign _17153_ = _17145_ & _17152_ /*15582*/;
assign _17150_ = _17151_ | _17153_ /*15580*/;
assign _16969_ = _17145_ ^ _17152_ /*15583*/;
assign _17159_ = D[30] ^ Q[20] /*15579*/;
assign _17156_ = _16584_ & _17159_ /*15575*/;
assign _17157_ = _16584_ ^ _17159_ /*15578*/;
assign _17158_ = _17150_ & _17157_ /*15576*/;
assign _17155_ = _17156_ | _17158_ /*15574*/;
assign _16970_ = _17150_ ^ _17157_ /*15577*/;
assign _17164_ = D[31] ^ Q[20] /*15573*/;
assign _17161_ = _16585_ & _17164_ /*15569*/;
assign _17162_ = _16585_ ^ _17164_ /*15572*/;
assign _17163_ = _17155_ & _17162_ /*15570*/;
assign _17160_ = _17161_ | _17163_ /*15568*/;
assign _16971_ = _17155_ ^ _17162_ /*15571*/;
assign _17169_ = D[32] ^ Q[20] /*15567*/;
assign _17166_ = _16586_ & _17169_ /*15563*/;
assign _17167_ = _16586_ ^ _17169_ /*15566*/;
assign _17168_ = _17160_ & _17167_ /*15564*/;
assign _17165_ = _17166_ | _17168_ /*15562*/;
assign _16972_ = _17160_ ^ _17167_ /*15565*/;
assign _17174_ = D[33] ^ Q[20] /*15561*/;
assign _17171_ = _16587_ & _17174_ /*15557*/;
assign _17172_ = _16587_ ^ _17174_ /*15560*/;
assign _17173_ = _17165_ & _17172_ /*15558*/;
assign _17170_ = _17171_ | _17173_ /*15556*/;
assign _16973_ = _17165_ ^ _17172_ /*15559*/;
assign _17179_ = D[34] ^ Q[20] /*15555*/;
assign _17176_ = _16588_ & _17179_ /*15551*/;
assign _17177_ = _16588_ ^ _17179_ /*15554*/;
assign _17178_ = _17170_ & _17177_ /*15552*/;
assign _17175_ = _17176_ | _17178_ /*15550*/;
assign _16974_ = _17170_ ^ _17177_ /*15553*/;
assign _17184_ = D[35] ^ Q[20] /*15549*/;
assign _17181_ = _16589_ & _17184_ /*15545*/;
assign _17182_ = _16589_ ^ _17184_ /*15548*/;
assign _17183_ = _17175_ & _17182_ /*15546*/;
assign _17180_ = _17181_ | _17183_ /*15544*/;
assign _16975_ = _17175_ ^ _17182_ /*15547*/;
assign _17189_ = D[36] ^ Q[20] /*15543*/;
assign _17186_ = _16590_ & _17189_ /*15539*/;
assign _17187_ = _16590_ ^ _17189_ /*15542*/;
assign _17188_ = _17180_ & _17187_ /*15540*/;
assign _17185_ = _17186_ | _17188_ /*15538*/;
assign _16976_ = _17180_ ^ _17187_ /*15541*/;
assign _17194_ = D[37] ^ Q[20] /*15537*/;
assign _17191_ = _16591_ & _17194_ /*15533*/;
assign _17192_ = _16591_ ^ _17194_ /*15536*/;
assign _17193_ = _17185_ & _17192_ /*15534*/;
assign _17190_ = _17191_ | _17193_ /*15532*/;
assign _16977_ = _17185_ ^ _17192_ /*15535*/;
assign _17199_ = D[38] ^ Q[20] /*15531*/;
assign _17196_ = _16592_ & _17199_ /*15527*/;
assign _17197_ = _16592_ ^ _17199_ /*15530*/;
assign _17198_ = _17190_ & _17197_ /*15528*/;
assign _17195_ = _17196_ | _17198_ /*15526*/;
assign _16978_ = _17190_ ^ _17197_ /*15529*/;
assign _17204_ = D[39] ^ Q[20] /*15525*/;
assign _17201_ = _16593_ & _17204_ /*15521*/;
assign _17202_ = _16593_ ^ _17204_ /*15524*/;
assign _17203_ = _17195_ & _17202_ /*15522*/;
assign _17200_ = _17201_ | _17203_ /*15520*/;
assign _16979_ = _17195_ ^ _17202_ /*15523*/;
assign _17209_ = D[40] ^ Q[20] /*15519*/;
assign _17206_ = _16594_ & _17209_ /*15515*/;
assign _17207_ = _16594_ ^ _17209_ /*15518*/;
assign _17208_ = _17200_ & _17207_ /*15516*/;
assign _17205_ = _17206_ | _17208_ /*15514*/;
assign _16980_ = _17200_ ^ _17207_ /*15517*/;
assign _17214_ = D[41] ^ Q[20] /*15513*/;
assign _17211_ = _16595_ & _17214_ /*15509*/;
assign _17212_ = _16595_ ^ _17214_ /*15512*/;
assign _17213_ = _17205_ & _17212_ /*15510*/;
assign _17210_ = _17211_ | _17213_ /*15508*/;
assign _16981_ = _17205_ ^ _17212_ /*15511*/;
assign _17219_ = D[42] ^ Q[20] /*15507*/;
assign _17216_ = _16596_ & _17219_ /*15503*/;
assign _17217_ = _16596_ ^ _17219_ /*15506*/;
assign _17218_ = _17210_ & _17217_ /*15504*/;
assign _17215_ = _17216_ | _17218_ /*15502*/;
assign _16982_ = _17210_ ^ _17217_ /*15505*/;
assign _17224_ = D[43] ^ Q[20] /*15501*/;
assign _17221_ = _16597_ & _17224_ /*15497*/;
assign _17222_ = _16597_ ^ _17224_ /*15500*/;
assign _17223_ = _17215_ & _17222_ /*15498*/;
assign _17220_ = _17221_ | _17223_ /*15496*/;
assign _16983_ = _17215_ ^ _17222_ /*15499*/;
assign _17229_ = D[44] ^ Q[20] /*15495*/;
assign _17226_ = _16598_ & _17229_ /*15491*/;
assign _17227_ = _16598_ ^ _17229_ /*15494*/;
assign _17228_ = _17220_ & _17227_ /*15492*/;
assign _17225_ = _17226_ | _17228_ /*15490*/;
assign _16984_ = _17220_ ^ _17227_ /*15493*/;
assign _17234_ = D[45] ^ Q[20] /*15489*/;
assign _17231_ = _16599_ & _17234_ /*15485*/;
assign _17232_ = _16599_ ^ _17234_ /*15488*/;
assign _17233_ = _17225_ & _17232_ /*15486*/;
assign _17230_ = _17231_ | _17233_ /*15484*/;
assign _16985_ = _17225_ ^ _17232_ /*15487*/;
assign _17239_ = D[46] ^ Q[20] /*15483*/;
assign _17236_ = _16600_ & _17239_ /*15479*/;
assign _17237_ = _16600_ ^ _17239_ /*15482*/;
assign _17238_ = _17230_ & _17237_ /*15480*/;
assign _17235_ = _17236_ | _17238_ /*15478*/;
assign _16986_ = _17230_ ^ _17237_ /*15481*/;
assign _17244_ = D[47] ^ Q[20] /*15477*/;
assign _17241_ = _16601_ & _17244_ /*15473*/;
assign _17242_ = _16601_ ^ _17244_ /*15476*/;
assign _17243_ = _17235_ & _17242_ /*15474*/;
assign _17240_ = _17241_ | _17243_ /*15472*/;
assign _16987_ = _17235_ ^ _17242_ /*15475*/;
assign _17249_ = D[48] ^ Q[20] /*15471*/;
assign _17246_ = _16602_ & _17249_ /*15467*/;
assign _17247_ = _16602_ ^ _17249_ /*15470*/;
assign _17248_ = _17240_ & _17247_ /*15468*/;
assign _17245_ = _17246_ | _17248_ /*15466*/;
assign _16988_ = _17240_ ^ _17247_ /*15469*/;
assign _17254_ = D[49] ^ Q[20] /*15465*/;
assign _17251_ = _16603_ & _17254_ /*15461*/;
assign _17252_ = _16603_ ^ _17254_ /*15464*/;
assign _17253_ = _17245_ & _17252_ /*15462*/;
assign _17250_ = _17251_ | _17253_ /*15460*/;
assign _16989_ = _17245_ ^ _17252_ /*15463*/;
assign _17259_ = D[50] ^ Q[20] /*15459*/;
assign _17256_ = _16604_ & _17259_ /*15455*/;
assign _17257_ = _16604_ ^ _17259_ /*15458*/;
assign _17258_ = _17250_ & _17257_ /*15456*/;
assign _17255_ = _17256_ | _17258_ /*15454*/;
assign _16990_ = _17250_ ^ _17257_ /*15457*/;
assign _17264_ = D[51] ^ Q[20] /*15453*/;
assign _17261_ = _16605_ & _17264_ /*15449*/;
assign _17262_ = _16605_ ^ _17264_ /*15452*/;
assign _17263_ = _17255_ & _17262_ /*15450*/;
assign _17260_ = _17261_ | _17263_ /*15448*/;
assign _16991_ = _17255_ ^ _17262_ /*15451*/;
assign _17269_ = D[52] ^ Q[20] /*15447*/;
assign _17266_ = _16606_ & _17269_ /*15443*/;
assign _17267_ = _16606_ ^ _17269_ /*15446*/;
assign _17268_ = _17260_ & _17267_ /*15444*/;
assign _17265_ = _17266_ | _17268_ /*15442*/;
assign _16992_ = _17260_ ^ _17267_ /*15445*/;
assign _17274_ = D[53] ^ Q[20] /*15441*/;
assign _17271_ = _16607_ & _17274_ /*15437*/;
assign _17272_ = _16607_ ^ _17274_ /*15440*/;
assign _17273_ = _17265_ & _17272_ /*15438*/;
assign _17270_ = _17271_ | _17273_ /*15436*/;
assign _16993_ = _17265_ ^ _17272_ /*15439*/;
assign _17279_ = D[54] ^ Q[20] /*15435*/;
assign _17276_ = _16608_ & _17279_ /*15431*/;
assign _17277_ = _16608_ ^ _17279_ /*15434*/;
assign _17278_ = _17270_ & _17277_ /*15432*/;
assign _17275_ = _17276_ | _17278_ /*15430*/;
assign _16994_ = _17270_ ^ _17277_ /*15433*/;
assign _17284_ = D[55] ^ Q[20] /*15429*/;
assign _17281_ = _16609_ & _17284_ /*15425*/;
assign _17282_ = _16609_ ^ _17284_ /*15428*/;
assign _17283_ = _17275_ & _17282_ /*15426*/;
assign _17280_ = _17281_ | _17283_ /*15424*/;
assign _16995_ = _17275_ ^ _17282_ /*15427*/;
assign _17289_ = D[56] ^ Q[20] /*15423*/;
assign _17286_ = _16610_ & _17289_ /*15419*/;
assign _17287_ = _16610_ ^ _17289_ /*15422*/;
assign _17288_ = _17280_ & _17287_ /*15420*/;
assign _17285_ = _17286_ | _17288_ /*15418*/;
assign _16996_ = _17280_ ^ _17287_ /*15421*/;
assign _17294_ = D[57] ^ Q[20] /*15417*/;
assign _17291_ = _16611_ & _17294_ /*15413*/;
assign _17292_ = _16611_ ^ _17294_ /*15416*/;
assign _17293_ = _17285_ & _17292_ /*15414*/;
assign _17290_ = _17291_ | _17293_ /*15412*/;
assign _16997_ = _17285_ ^ _17292_ /*15415*/;
assign _17299_ = D[58] ^ Q[20] /*15411*/;
assign _17296_ = _16612_ & _17299_ /*15407*/;
assign _17297_ = _16612_ ^ _17299_ /*15410*/;
assign _17298_ = _17290_ & _17297_ /*15408*/;
assign _17295_ = _17296_ | _17298_ /*15406*/;
assign _16998_ = _17290_ ^ _17297_ /*15409*/;
assign _17304_ = D[59] ^ Q[20] /*15405*/;
assign _17301_ = _16613_ & _17304_ /*15401*/;
assign _17302_ = _16613_ ^ _17304_ /*15404*/;
assign _17303_ = _17295_ & _17302_ /*15402*/;
assign _17300_ = _17301_ | _17303_ /*15400*/;
assign _16999_ = _17295_ ^ _17302_ /*15403*/;
assign _17309_ = D[60] ^ Q[20] /*15399*/;
assign _17306_ = _16614_ & _17309_ /*15395*/;
assign _17307_ = _16614_ ^ _17309_ /*15398*/;
assign _17308_ = _17300_ & _17307_ /*15396*/;
assign _17305_ = _17306_ | _17308_ /*15394*/;
assign _17000_ = _17300_ ^ _17307_ /*15397*/;
assign _17314_ = D[61] ^ Q[20] /*15393*/;
assign _17311_ = _16615_ & _17314_ /*15389*/;
assign _17312_ = _16615_ ^ _17314_ /*15392*/;
assign _17313_ = _17305_ & _17312_ /*15390*/;
assign _17310_ = _17311_ | _17313_ /*15388*/;
assign _17001_ = _17305_ ^ _17312_ /*15391*/;
assign _17319_ = D[62] ^ Q[20] /*15387*/;
assign _17316_ = _16616_ & _17319_ /*15383*/;
assign _17317_ = _16616_ ^ _17319_ /*15386*/;
assign _17318_ = _17310_ & _17317_ /*15384*/;
assign _17315_ = _17316_ | _17318_ /*15382*/;
assign _17002_ = _17310_ ^ _17317_ /*15385*/;
assign _17323_ = zeroWire ^ Q[20] /*15381*/;
assign _17320_ = _16617_ & _17323_ /*15377*/;
assign _17321_ = _16617_ ^ _17323_ /*15380*/;
assign _17322_ = _17315_ & _17321_ /*15378*/;
assign Q[19] = _17320_ | _17322_ /*15376*/;
assign _17003_ = _17315_ ^ _17321_ /*15379*/;
assign _17394_ = D[0] ^ Q[19] /*14990*/;
assign _17391_ = R_0[18] & _17394_ /*14986*/;
assign _17392_ = R_0[18] ^ _17394_ /*14989*/;
assign _17393_ = Q[19] & _17392_ /*14987*/;
assign _17390_ = _17391_ | _17393_ /*14985*/;
assign _17325_ = Q[19] ^ _17392_ /*14988*/;
assign _17399_ = D[1] ^ Q[19] /*14984*/;
assign _17396_ = _16940_ & _17399_ /*14980*/;
assign _17397_ = _16940_ ^ _17399_ /*14983*/;
assign _17398_ = _17390_ & _17397_ /*14981*/;
assign _17395_ = _17396_ | _17398_ /*14979*/;
assign _17326_ = _17390_ ^ _17397_ /*14982*/;
assign _17404_ = D[2] ^ Q[19] /*14978*/;
assign _17401_ = _16941_ & _17404_ /*14974*/;
assign _17402_ = _16941_ ^ _17404_ /*14977*/;
assign _17403_ = _17395_ & _17402_ /*14975*/;
assign _17400_ = _17401_ | _17403_ /*14973*/;
assign _17327_ = _17395_ ^ _17402_ /*14976*/;
assign _17409_ = D[3] ^ Q[19] /*14972*/;
assign _17406_ = _16942_ & _17409_ /*14968*/;
assign _17407_ = _16942_ ^ _17409_ /*14971*/;
assign _17408_ = _17400_ & _17407_ /*14969*/;
assign _17405_ = _17406_ | _17408_ /*14967*/;
assign _17328_ = _17400_ ^ _17407_ /*14970*/;
assign _17414_ = D[4] ^ Q[19] /*14966*/;
assign _17411_ = _16943_ & _17414_ /*14962*/;
assign _17412_ = _16943_ ^ _17414_ /*14965*/;
assign _17413_ = _17405_ & _17412_ /*14963*/;
assign _17410_ = _17411_ | _17413_ /*14961*/;
assign _17329_ = _17405_ ^ _17412_ /*14964*/;
assign _17419_ = D[5] ^ Q[19] /*14960*/;
assign _17416_ = _16944_ & _17419_ /*14956*/;
assign _17417_ = _16944_ ^ _17419_ /*14959*/;
assign _17418_ = _17410_ & _17417_ /*14957*/;
assign _17415_ = _17416_ | _17418_ /*14955*/;
assign _17330_ = _17410_ ^ _17417_ /*14958*/;
assign _17424_ = D[6] ^ Q[19] /*14954*/;
assign _17421_ = _16945_ & _17424_ /*14950*/;
assign _17422_ = _16945_ ^ _17424_ /*14953*/;
assign _17423_ = _17415_ & _17422_ /*14951*/;
assign _17420_ = _17421_ | _17423_ /*14949*/;
assign _17331_ = _17415_ ^ _17422_ /*14952*/;
assign _17429_ = D[7] ^ Q[19] /*14948*/;
assign _17426_ = _16946_ & _17429_ /*14944*/;
assign _17427_ = _16946_ ^ _17429_ /*14947*/;
assign _17428_ = _17420_ & _17427_ /*14945*/;
assign _17425_ = _17426_ | _17428_ /*14943*/;
assign _17332_ = _17420_ ^ _17427_ /*14946*/;
assign _17434_ = D[8] ^ Q[19] /*14942*/;
assign _17431_ = _16947_ & _17434_ /*14938*/;
assign _17432_ = _16947_ ^ _17434_ /*14941*/;
assign _17433_ = _17425_ & _17432_ /*14939*/;
assign _17430_ = _17431_ | _17433_ /*14937*/;
assign _17333_ = _17425_ ^ _17432_ /*14940*/;
assign _17439_ = D[9] ^ Q[19] /*14936*/;
assign _17436_ = _16948_ & _17439_ /*14932*/;
assign _17437_ = _16948_ ^ _17439_ /*14935*/;
assign _17438_ = _17430_ & _17437_ /*14933*/;
assign _17435_ = _17436_ | _17438_ /*14931*/;
assign _17334_ = _17430_ ^ _17437_ /*14934*/;
assign _17444_ = D[10] ^ Q[19] /*14930*/;
assign _17441_ = _16949_ & _17444_ /*14926*/;
assign _17442_ = _16949_ ^ _17444_ /*14929*/;
assign _17443_ = _17435_ & _17442_ /*14927*/;
assign _17440_ = _17441_ | _17443_ /*14925*/;
assign _17335_ = _17435_ ^ _17442_ /*14928*/;
assign _17449_ = D[11] ^ Q[19] /*14924*/;
assign _17446_ = _16950_ & _17449_ /*14920*/;
assign _17447_ = _16950_ ^ _17449_ /*14923*/;
assign _17448_ = _17440_ & _17447_ /*14921*/;
assign _17445_ = _17446_ | _17448_ /*14919*/;
assign _17336_ = _17440_ ^ _17447_ /*14922*/;
assign _17454_ = D[12] ^ Q[19] /*14918*/;
assign _17451_ = _16951_ & _17454_ /*14914*/;
assign _17452_ = _16951_ ^ _17454_ /*14917*/;
assign _17453_ = _17445_ & _17452_ /*14915*/;
assign _17450_ = _17451_ | _17453_ /*14913*/;
assign _17337_ = _17445_ ^ _17452_ /*14916*/;
assign _17459_ = D[13] ^ Q[19] /*14912*/;
assign _17456_ = _16952_ & _17459_ /*14908*/;
assign _17457_ = _16952_ ^ _17459_ /*14911*/;
assign _17458_ = _17450_ & _17457_ /*14909*/;
assign _17455_ = _17456_ | _17458_ /*14907*/;
assign _17338_ = _17450_ ^ _17457_ /*14910*/;
assign _17464_ = D[14] ^ Q[19] /*14906*/;
assign _17461_ = _16953_ & _17464_ /*14902*/;
assign _17462_ = _16953_ ^ _17464_ /*14905*/;
assign _17463_ = _17455_ & _17462_ /*14903*/;
assign _17460_ = _17461_ | _17463_ /*14901*/;
assign _17339_ = _17455_ ^ _17462_ /*14904*/;
assign _17469_ = D[15] ^ Q[19] /*14900*/;
assign _17466_ = _16954_ & _17469_ /*14896*/;
assign _17467_ = _16954_ ^ _17469_ /*14899*/;
assign _17468_ = _17460_ & _17467_ /*14897*/;
assign _17465_ = _17466_ | _17468_ /*14895*/;
assign _17340_ = _17460_ ^ _17467_ /*14898*/;
assign _17474_ = D[16] ^ Q[19] /*14894*/;
assign _17471_ = _16955_ & _17474_ /*14890*/;
assign _17472_ = _16955_ ^ _17474_ /*14893*/;
assign _17473_ = _17465_ & _17472_ /*14891*/;
assign _17470_ = _17471_ | _17473_ /*14889*/;
assign _17341_ = _17465_ ^ _17472_ /*14892*/;
assign _17479_ = D[17] ^ Q[19] /*14888*/;
assign _17476_ = _16956_ & _17479_ /*14884*/;
assign _17477_ = _16956_ ^ _17479_ /*14887*/;
assign _17478_ = _17470_ & _17477_ /*14885*/;
assign _17475_ = _17476_ | _17478_ /*14883*/;
assign _17342_ = _17470_ ^ _17477_ /*14886*/;
assign _17484_ = D[18] ^ Q[19] /*14882*/;
assign _17481_ = _16957_ & _17484_ /*14878*/;
assign _17482_ = _16957_ ^ _17484_ /*14881*/;
assign _17483_ = _17475_ & _17482_ /*14879*/;
assign _17480_ = _17481_ | _17483_ /*14877*/;
assign _17343_ = _17475_ ^ _17482_ /*14880*/;
assign _17489_ = D[19] ^ Q[19] /*14876*/;
assign _17486_ = _16958_ & _17489_ /*14872*/;
assign _17487_ = _16958_ ^ _17489_ /*14875*/;
assign _17488_ = _17480_ & _17487_ /*14873*/;
assign _17485_ = _17486_ | _17488_ /*14871*/;
assign _17344_ = _17480_ ^ _17487_ /*14874*/;
assign _17494_ = D[20] ^ Q[19] /*14870*/;
assign _17491_ = _16959_ & _17494_ /*14866*/;
assign _17492_ = _16959_ ^ _17494_ /*14869*/;
assign _17493_ = _17485_ & _17492_ /*14867*/;
assign _17490_ = _17491_ | _17493_ /*14865*/;
assign _17345_ = _17485_ ^ _17492_ /*14868*/;
assign _17499_ = D[21] ^ Q[19] /*14864*/;
assign _17496_ = _16960_ & _17499_ /*14860*/;
assign _17497_ = _16960_ ^ _17499_ /*14863*/;
assign _17498_ = _17490_ & _17497_ /*14861*/;
assign _17495_ = _17496_ | _17498_ /*14859*/;
assign _17346_ = _17490_ ^ _17497_ /*14862*/;
assign _17504_ = D[22] ^ Q[19] /*14858*/;
assign _17501_ = _16961_ & _17504_ /*14854*/;
assign _17502_ = _16961_ ^ _17504_ /*14857*/;
assign _17503_ = _17495_ & _17502_ /*14855*/;
assign _17500_ = _17501_ | _17503_ /*14853*/;
assign _17347_ = _17495_ ^ _17502_ /*14856*/;
assign _17509_ = D[23] ^ Q[19] /*14852*/;
assign _17506_ = _16962_ & _17509_ /*14848*/;
assign _17507_ = _16962_ ^ _17509_ /*14851*/;
assign _17508_ = _17500_ & _17507_ /*14849*/;
assign _17505_ = _17506_ | _17508_ /*14847*/;
assign _17348_ = _17500_ ^ _17507_ /*14850*/;
assign _17514_ = D[24] ^ Q[19] /*14846*/;
assign _17511_ = _16963_ & _17514_ /*14842*/;
assign _17512_ = _16963_ ^ _17514_ /*14845*/;
assign _17513_ = _17505_ & _17512_ /*14843*/;
assign _17510_ = _17511_ | _17513_ /*14841*/;
assign _17349_ = _17505_ ^ _17512_ /*14844*/;
assign _17519_ = D[25] ^ Q[19] /*14840*/;
assign _17516_ = _16964_ & _17519_ /*14836*/;
assign _17517_ = _16964_ ^ _17519_ /*14839*/;
assign _17518_ = _17510_ & _17517_ /*14837*/;
assign _17515_ = _17516_ | _17518_ /*14835*/;
assign _17350_ = _17510_ ^ _17517_ /*14838*/;
assign _17524_ = D[26] ^ Q[19] /*14834*/;
assign _17521_ = _16965_ & _17524_ /*14830*/;
assign _17522_ = _16965_ ^ _17524_ /*14833*/;
assign _17523_ = _17515_ & _17522_ /*14831*/;
assign _17520_ = _17521_ | _17523_ /*14829*/;
assign _17351_ = _17515_ ^ _17522_ /*14832*/;
assign _17529_ = D[27] ^ Q[19] /*14828*/;
assign _17526_ = _16966_ & _17529_ /*14824*/;
assign _17527_ = _16966_ ^ _17529_ /*14827*/;
assign _17528_ = _17520_ & _17527_ /*14825*/;
assign _17525_ = _17526_ | _17528_ /*14823*/;
assign _17352_ = _17520_ ^ _17527_ /*14826*/;
assign _17534_ = D[28] ^ Q[19] /*14822*/;
assign _17531_ = _16967_ & _17534_ /*14818*/;
assign _17532_ = _16967_ ^ _17534_ /*14821*/;
assign _17533_ = _17525_ & _17532_ /*14819*/;
assign _17530_ = _17531_ | _17533_ /*14817*/;
assign _17353_ = _17525_ ^ _17532_ /*14820*/;
assign _17539_ = D[29] ^ Q[19] /*14816*/;
assign _17536_ = _16968_ & _17539_ /*14812*/;
assign _17537_ = _16968_ ^ _17539_ /*14815*/;
assign _17538_ = _17530_ & _17537_ /*14813*/;
assign _17535_ = _17536_ | _17538_ /*14811*/;
assign _17354_ = _17530_ ^ _17537_ /*14814*/;
assign _17544_ = D[30] ^ Q[19] /*14810*/;
assign _17541_ = _16969_ & _17544_ /*14806*/;
assign _17542_ = _16969_ ^ _17544_ /*14809*/;
assign _17543_ = _17535_ & _17542_ /*14807*/;
assign _17540_ = _17541_ | _17543_ /*14805*/;
assign _17355_ = _17535_ ^ _17542_ /*14808*/;
assign _17549_ = D[31] ^ Q[19] /*14804*/;
assign _17546_ = _16970_ & _17549_ /*14800*/;
assign _17547_ = _16970_ ^ _17549_ /*14803*/;
assign _17548_ = _17540_ & _17547_ /*14801*/;
assign _17545_ = _17546_ | _17548_ /*14799*/;
assign _17356_ = _17540_ ^ _17547_ /*14802*/;
assign _17554_ = D[32] ^ Q[19] /*14798*/;
assign _17551_ = _16971_ & _17554_ /*14794*/;
assign _17552_ = _16971_ ^ _17554_ /*14797*/;
assign _17553_ = _17545_ & _17552_ /*14795*/;
assign _17550_ = _17551_ | _17553_ /*14793*/;
assign _17357_ = _17545_ ^ _17552_ /*14796*/;
assign _17559_ = D[33] ^ Q[19] /*14792*/;
assign _17556_ = _16972_ & _17559_ /*14788*/;
assign _17557_ = _16972_ ^ _17559_ /*14791*/;
assign _17558_ = _17550_ & _17557_ /*14789*/;
assign _17555_ = _17556_ | _17558_ /*14787*/;
assign _17358_ = _17550_ ^ _17557_ /*14790*/;
assign _17564_ = D[34] ^ Q[19] /*14786*/;
assign _17561_ = _16973_ & _17564_ /*14782*/;
assign _17562_ = _16973_ ^ _17564_ /*14785*/;
assign _17563_ = _17555_ & _17562_ /*14783*/;
assign _17560_ = _17561_ | _17563_ /*14781*/;
assign _17359_ = _17555_ ^ _17562_ /*14784*/;
assign _17569_ = D[35] ^ Q[19] /*14780*/;
assign _17566_ = _16974_ & _17569_ /*14776*/;
assign _17567_ = _16974_ ^ _17569_ /*14779*/;
assign _17568_ = _17560_ & _17567_ /*14777*/;
assign _17565_ = _17566_ | _17568_ /*14775*/;
assign _17360_ = _17560_ ^ _17567_ /*14778*/;
assign _17574_ = D[36] ^ Q[19] /*14774*/;
assign _17571_ = _16975_ & _17574_ /*14770*/;
assign _17572_ = _16975_ ^ _17574_ /*14773*/;
assign _17573_ = _17565_ & _17572_ /*14771*/;
assign _17570_ = _17571_ | _17573_ /*14769*/;
assign _17361_ = _17565_ ^ _17572_ /*14772*/;
assign _17579_ = D[37] ^ Q[19] /*14768*/;
assign _17576_ = _16976_ & _17579_ /*14764*/;
assign _17577_ = _16976_ ^ _17579_ /*14767*/;
assign _17578_ = _17570_ & _17577_ /*14765*/;
assign _17575_ = _17576_ | _17578_ /*14763*/;
assign _17362_ = _17570_ ^ _17577_ /*14766*/;
assign _17584_ = D[38] ^ Q[19] /*14762*/;
assign _17581_ = _16977_ & _17584_ /*14758*/;
assign _17582_ = _16977_ ^ _17584_ /*14761*/;
assign _17583_ = _17575_ & _17582_ /*14759*/;
assign _17580_ = _17581_ | _17583_ /*14757*/;
assign _17363_ = _17575_ ^ _17582_ /*14760*/;
assign _17589_ = D[39] ^ Q[19] /*14756*/;
assign _17586_ = _16978_ & _17589_ /*14752*/;
assign _17587_ = _16978_ ^ _17589_ /*14755*/;
assign _17588_ = _17580_ & _17587_ /*14753*/;
assign _17585_ = _17586_ | _17588_ /*14751*/;
assign _17364_ = _17580_ ^ _17587_ /*14754*/;
assign _17594_ = D[40] ^ Q[19] /*14750*/;
assign _17591_ = _16979_ & _17594_ /*14746*/;
assign _17592_ = _16979_ ^ _17594_ /*14749*/;
assign _17593_ = _17585_ & _17592_ /*14747*/;
assign _17590_ = _17591_ | _17593_ /*14745*/;
assign _17365_ = _17585_ ^ _17592_ /*14748*/;
assign _17599_ = D[41] ^ Q[19] /*14744*/;
assign _17596_ = _16980_ & _17599_ /*14740*/;
assign _17597_ = _16980_ ^ _17599_ /*14743*/;
assign _17598_ = _17590_ & _17597_ /*14741*/;
assign _17595_ = _17596_ | _17598_ /*14739*/;
assign _17366_ = _17590_ ^ _17597_ /*14742*/;
assign _17604_ = D[42] ^ Q[19] /*14738*/;
assign _17601_ = _16981_ & _17604_ /*14734*/;
assign _17602_ = _16981_ ^ _17604_ /*14737*/;
assign _17603_ = _17595_ & _17602_ /*14735*/;
assign _17600_ = _17601_ | _17603_ /*14733*/;
assign _17367_ = _17595_ ^ _17602_ /*14736*/;
assign _17609_ = D[43] ^ Q[19] /*14732*/;
assign _17606_ = _16982_ & _17609_ /*14728*/;
assign _17607_ = _16982_ ^ _17609_ /*14731*/;
assign _17608_ = _17600_ & _17607_ /*14729*/;
assign _17605_ = _17606_ | _17608_ /*14727*/;
assign _17368_ = _17600_ ^ _17607_ /*14730*/;
assign _17614_ = D[44] ^ Q[19] /*14726*/;
assign _17611_ = _16983_ & _17614_ /*14722*/;
assign _17612_ = _16983_ ^ _17614_ /*14725*/;
assign _17613_ = _17605_ & _17612_ /*14723*/;
assign _17610_ = _17611_ | _17613_ /*14721*/;
assign _17369_ = _17605_ ^ _17612_ /*14724*/;
assign _17619_ = D[45] ^ Q[19] /*14720*/;
assign _17616_ = _16984_ & _17619_ /*14716*/;
assign _17617_ = _16984_ ^ _17619_ /*14719*/;
assign _17618_ = _17610_ & _17617_ /*14717*/;
assign _17615_ = _17616_ | _17618_ /*14715*/;
assign _17370_ = _17610_ ^ _17617_ /*14718*/;
assign _17624_ = D[46] ^ Q[19] /*14714*/;
assign _17621_ = _16985_ & _17624_ /*14710*/;
assign _17622_ = _16985_ ^ _17624_ /*14713*/;
assign _17623_ = _17615_ & _17622_ /*14711*/;
assign _17620_ = _17621_ | _17623_ /*14709*/;
assign _17371_ = _17615_ ^ _17622_ /*14712*/;
assign _17629_ = D[47] ^ Q[19] /*14708*/;
assign _17626_ = _16986_ & _17629_ /*14704*/;
assign _17627_ = _16986_ ^ _17629_ /*14707*/;
assign _17628_ = _17620_ & _17627_ /*14705*/;
assign _17625_ = _17626_ | _17628_ /*14703*/;
assign _17372_ = _17620_ ^ _17627_ /*14706*/;
assign _17634_ = D[48] ^ Q[19] /*14702*/;
assign _17631_ = _16987_ & _17634_ /*14698*/;
assign _17632_ = _16987_ ^ _17634_ /*14701*/;
assign _17633_ = _17625_ & _17632_ /*14699*/;
assign _17630_ = _17631_ | _17633_ /*14697*/;
assign _17373_ = _17625_ ^ _17632_ /*14700*/;
assign _17639_ = D[49] ^ Q[19] /*14696*/;
assign _17636_ = _16988_ & _17639_ /*14692*/;
assign _17637_ = _16988_ ^ _17639_ /*14695*/;
assign _17638_ = _17630_ & _17637_ /*14693*/;
assign _17635_ = _17636_ | _17638_ /*14691*/;
assign _17374_ = _17630_ ^ _17637_ /*14694*/;
assign _17644_ = D[50] ^ Q[19] /*14690*/;
assign _17641_ = _16989_ & _17644_ /*14686*/;
assign _17642_ = _16989_ ^ _17644_ /*14689*/;
assign _17643_ = _17635_ & _17642_ /*14687*/;
assign _17640_ = _17641_ | _17643_ /*14685*/;
assign _17375_ = _17635_ ^ _17642_ /*14688*/;
assign _17649_ = D[51] ^ Q[19] /*14684*/;
assign _17646_ = _16990_ & _17649_ /*14680*/;
assign _17647_ = _16990_ ^ _17649_ /*14683*/;
assign _17648_ = _17640_ & _17647_ /*14681*/;
assign _17645_ = _17646_ | _17648_ /*14679*/;
assign _17376_ = _17640_ ^ _17647_ /*14682*/;
assign _17654_ = D[52] ^ Q[19] /*14678*/;
assign _17651_ = _16991_ & _17654_ /*14674*/;
assign _17652_ = _16991_ ^ _17654_ /*14677*/;
assign _17653_ = _17645_ & _17652_ /*14675*/;
assign _17650_ = _17651_ | _17653_ /*14673*/;
assign _17377_ = _17645_ ^ _17652_ /*14676*/;
assign _17659_ = D[53] ^ Q[19] /*14672*/;
assign _17656_ = _16992_ & _17659_ /*14668*/;
assign _17657_ = _16992_ ^ _17659_ /*14671*/;
assign _17658_ = _17650_ & _17657_ /*14669*/;
assign _17655_ = _17656_ | _17658_ /*14667*/;
assign _17378_ = _17650_ ^ _17657_ /*14670*/;
assign _17664_ = D[54] ^ Q[19] /*14666*/;
assign _17661_ = _16993_ & _17664_ /*14662*/;
assign _17662_ = _16993_ ^ _17664_ /*14665*/;
assign _17663_ = _17655_ & _17662_ /*14663*/;
assign _17660_ = _17661_ | _17663_ /*14661*/;
assign _17379_ = _17655_ ^ _17662_ /*14664*/;
assign _17669_ = D[55] ^ Q[19] /*14660*/;
assign _17666_ = _16994_ & _17669_ /*14656*/;
assign _17667_ = _16994_ ^ _17669_ /*14659*/;
assign _17668_ = _17660_ & _17667_ /*14657*/;
assign _17665_ = _17666_ | _17668_ /*14655*/;
assign _17380_ = _17660_ ^ _17667_ /*14658*/;
assign _17674_ = D[56] ^ Q[19] /*14654*/;
assign _17671_ = _16995_ & _17674_ /*14650*/;
assign _17672_ = _16995_ ^ _17674_ /*14653*/;
assign _17673_ = _17665_ & _17672_ /*14651*/;
assign _17670_ = _17671_ | _17673_ /*14649*/;
assign _17381_ = _17665_ ^ _17672_ /*14652*/;
assign _17679_ = D[57] ^ Q[19] /*14648*/;
assign _17676_ = _16996_ & _17679_ /*14644*/;
assign _17677_ = _16996_ ^ _17679_ /*14647*/;
assign _17678_ = _17670_ & _17677_ /*14645*/;
assign _17675_ = _17676_ | _17678_ /*14643*/;
assign _17382_ = _17670_ ^ _17677_ /*14646*/;
assign _17684_ = D[58] ^ Q[19] /*14642*/;
assign _17681_ = _16997_ & _17684_ /*14638*/;
assign _17682_ = _16997_ ^ _17684_ /*14641*/;
assign _17683_ = _17675_ & _17682_ /*14639*/;
assign _17680_ = _17681_ | _17683_ /*14637*/;
assign _17383_ = _17675_ ^ _17682_ /*14640*/;
assign _17689_ = D[59] ^ Q[19] /*14636*/;
assign _17686_ = _16998_ & _17689_ /*14632*/;
assign _17687_ = _16998_ ^ _17689_ /*14635*/;
assign _17688_ = _17680_ & _17687_ /*14633*/;
assign _17685_ = _17686_ | _17688_ /*14631*/;
assign _17384_ = _17680_ ^ _17687_ /*14634*/;
assign _17694_ = D[60] ^ Q[19] /*14630*/;
assign _17691_ = _16999_ & _17694_ /*14626*/;
assign _17692_ = _16999_ ^ _17694_ /*14629*/;
assign _17693_ = _17685_ & _17692_ /*14627*/;
assign _17690_ = _17691_ | _17693_ /*14625*/;
assign _17385_ = _17685_ ^ _17692_ /*14628*/;
assign _17699_ = D[61] ^ Q[19] /*14624*/;
assign _17696_ = _17000_ & _17699_ /*14620*/;
assign _17697_ = _17000_ ^ _17699_ /*14623*/;
assign _17698_ = _17690_ & _17697_ /*14621*/;
assign _17695_ = _17696_ | _17698_ /*14619*/;
assign _17386_ = _17690_ ^ _17697_ /*14622*/;
assign _17704_ = D[62] ^ Q[19] /*14618*/;
assign _17701_ = _17001_ & _17704_ /*14614*/;
assign _17702_ = _17001_ ^ _17704_ /*14617*/;
assign _17703_ = _17695_ & _17702_ /*14615*/;
assign _17700_ = _17701_ | _17703_ /*14613*/;
assign _17387_ = _17695_ ^ _17702_ /*14616*/;
assign _17708_ = zeroWire ^ Q[19] /*14612*/;
assign _17705_ = _17002_ & _17708_ /*14608*/;
assign _17706_ = _17002_ ^ _17708_ /*14611*/;
assign _17707_ = _17700_ & _17706_ /*14609*/;
assign Q[18] = _17705_ | _17707_ /*14607*/;
assign _17388_ = _17700_ ^ _17706_ /*14610*/;
assign _17779_ = D[0] ^ Q[18] /*14221*/;
assign _17776_ = R_0[17] & _17779_ /*14217*/;
assign _17777_ = R_0[17] ^ _17779_ /*14220*/;
assign _17778_ = Q[18] & _17777_ /*14218*/;
assign _17775_ = _17776_ | _17778_ /*14216*/;
assign _17710_ = Q[18] ^ _17777_ /*14219*/;
assign _17784_ = D[1] ^ Q[18] /*14215*/;
assign _17781_ = _17325_ & _17784_ /*14211*/;
assign _17782_ = _17325_ ^ _17784_ /*14214*/;
assign _17783_ = _17775_ & _17782_ /*14212*/;
assign _17780_ = _17781_ | _17783_ /*14210*/;
assign _17711_ = _17775_ ^ _17782_ /*14213*/;
assign _17789_ = D[2] ^ Q[18] /*14209*/;
assign _17786_ = _17326_ & _17789_ /*14205*/;
assign _17787_ = _17326_ ^ _17789_ /*14208*/;
assign _17788_ = _17780_ & _17787_ /*14206*/;
assign _17785_ = _17786_ | _17788_ /*14204*/;
assign _17712_ = _17780_ ^ _17787_ /*14207*/;
assign _17794_ = D[3] ^ Q[18] /*14203*/;
assign _17791_ = _17327_ & _17794_ /*14199*/;
assign _17792_ = _17327_ ^ _17794_ /*14202*/;
assign _17793_ = _17785_ & _17792_ /*14200*/;
assign _17790_ = _17791_ | _17793_ /*14198*/;
assign _17713_ = _17785_ ^ _17792_ /*14201*/;
assign _17799_ = D[4] ^ Q[18] /*14197*/;
assign _17796_ = _17328_ & _17799_ /*14193*/;
assign _17797_ = _17328_ ^ _17799_ /*14196*/;
assign _17798_ = _17790_ & _17797_ /*14194*/;
assign _17795_ = _17796_ | _17798_ /*14192*/;
assign _17714_ = _17790_ ^ _17797_ /*14195*/;
assign _17804_ = D[5] ^ Q[18] /*14191*/;
assign _17801_ = _17329_ & _17804_ /*14187*/;
assign _17802_ = _17329_ ^ _17804_ /*14190*/;
assign _17803_ = _17795_ & _17802_ /*14188*/;
assign _17800_ = _17801_ | _17803_ /*14186*/;
assign _17715_ = _17795_ ^ _17802_ /*14189*/;
assign _17809_ = D[6] ^ Q[18] /*14185*/;
assign _17806_ = _17330_ & _17809_ /*14181*/;
assign _17807_ = _17330_ ^ _17809_ /*14184*/;
assign _17808_ = _17800_ & _17807_ /*14182*/;
assign _17805_ = _17806_ | _17808_ /*14180*/;
assign _17716_ = _17800_ ^ _17807_ /*14183*/;
assign _17814_ = D[7] ^ Q[18] /*14179*/;
assign _17811_ = _17331_ & _17814_ /*14175*/;
assign _17812_ = _17331_ ^ _17814_ /*14178*/;
assign _17813_ = _17805_ & _17812_ /*14176*/;
assign _17810_ = _17811_ | _17813_ /*14174*/;
assign _17717_ = _17805_ ^ _17812_ /*14177*/;
assign _17819_ = D[8] ^ Q[18] /*14173*/;
assign _17816_ = _17332_ & _17819_ /*14169*/;
assign _17817_ = _17332_ ^ _17819_ /*14172*/;
assign _17818_ = _17810_ & _17817_ /*14170*/;
assign _17815_ = _17816_ | _17818_ /*14168*/;
assign _17718_ = _17810_ ^ _17817_ /*14171*/;
assign _17824_ = D[9] ^ Q[18] /*14167*/;
assign _17821_ = _17333_ & _17824_ /*14163*/;
assign _17822_ = _17333_ ^ _17824_ /*14166*/;
assign _17823_ = _17815_ & _17822_ /*14164*/;
assign _17820_ = _17821_ | _17823_ /*14162*/;
assign _17719_ = _17815_ ^ _17822_ /*14165*/;
assign _17829_ = D[10] ^ Q[18] /*14161*/;
assign _17826_ = _17334_ & _17829_ /*14157*/;
assign _17827_ = _17334_ ^ _17829_ /*14160*/;
assign _17828_ = _17820_ & _17827_ /*14158*/;
assign _17825_ = _17826_ | _17828_ /*14156*/;
assign _17720_ = _17820_ ^ _17827_ /*14159*/;
assign _17834_ = D[11] ^ Q[18] /*14155*/;
assign _17831_ = _17335_ & _17834_ /*14151*/;
assign _17832_ = _17335_ ^ _17834_ /*14154*/;
assign _17833_ = _17825_ & _17832_ /*14152*/;
assign _17830_ = _17831_ | _17833_ /*14150*/;
assign _17721_ = _17825_ ^ _17832_ /*14153*/;
assign _17839_ = D[12] ^ Q[18] /*14149*/;
assign _17836_ = _17336_ & _17839_ /*14145*/;
assign _17837_ = _17336_ ^ _17839_ /*14148*/;
assign _17838_ = _17830_ & _17837_ /*14146*/;
assign _17835_ = _17836_ | _17838_ /*14144*/;
assign _17722_ = _17830_ ^ _17837_ /*14147*/;
assign _17844_ = D[13] ^ Q[18] /*14143*/;
assign _17841_ = _17337_ & _17844_ /*14139*/;
assign _17842_ = _17337_ ^ _17844_ /*14142*/;
assign _17843_ = _17835_ & _17842_ /*14140*/;
assign _17840_ = _17841_ | _17843_ /*14138*/;
assign _17723_ = _17835_ ^ _17842_ /*14141*/;
assign _17849_ = D[14] ^ Q[18] /*14137*/;
assign _17846_ = _17338_ & _17849_ /*14133*/;
assign _17847_ = _17338_ ^ _17849_ /*14136*/;
assign _17848_ = _17840_ & _17847_ /*14134*/;
assign _17845_ = _17846_ | _17848_ /*14132*/;
assign _17724_ = _17840_ ^ _17847_ /*14135*/;
assign _17854_ = D[15] ^ Q[18] /*14131*/;
assign _17851_ = _17339_ & _17854_ /*14127*/;
assign _17852_ = _17339_ ^ _17854_ /*14130*/;
assign _17853_ = _17845_ & _17852_ /*14128*/;
assign _17850_ = _17851_ | _17853_ /*14126*/;
assign _17725_ = _17845_ ^ _17852_ /*14129*/;
assign _17859_ = D[16] ^ Q[18] /*14125*/;
assign _17856_ = _17340_ & _17859_ /*14121*/;
assign _17857_ = _17340_ ^ _17859_ /*14124*/;
assign _17858_ = _17850_ & _17857_ /*14122*/;
assign _17855_ = _17856_ | _17858_ /*14120*/;
assign _17726_ = _17850_ ^ _17857_ /*14123*/;
assign _17864_ = D[17] ^ Q[18] /*14119*/;
assign _17861_ = _17341_ & _17864_ /*14115*/;
assign _17862_ = _17341_ ^ _17864_ /*14118*/;
assign _17863_ = _17855_ & _17862_ /*14116*/;
assign _17860_ = _17861_ | _17863_ /*14114*/;
assign _17727_ = _17855_ ^ _17862_ /*14117*/;
assign _17869_ = D[18] ^ Q[18] /*14113*/;
assign _17866_ = _17342_ & _17869_ /*14109*/;
assign _17867_ = _17342_ ^ _17869_ /*14112*/;
assign _17868_ = _17860_ & _17867_ /*14110*/;
assign _17865_ = _17866_ | _17868_ /*14108*/;
assign _17728_ = _17860_ ^ _17867_ /*14111*/;
assign _17874_ = D[19] ^ Q[18] /*14107*/;
assign _17871_ = _17343_ & _17874_ /*14103*/;
assign _17872_ = _17343_ ^ _17874_ /*14106*/;
assign _17873_ = _17865_ & _17872_ /*14104*/;
assign _17870_ = _17871_ | _17873_ /*14102*/;
assign _17729_ = _17865_ ^ _17872_ /*14105*/;
assign _17879_ = D[20] ^ Q[18] /*14101*/;
assign _17876_ = _17344_ & _17879_ /*14097*/;
assign _17877_ = _17344_ ^ _17879_ /*14100*/;
assign _17878_ = _17870_ & _17877_ /*14098*/;
assign _17875_ = _17876_ | _17878_ /*14096*/;
assign _17730_ = _17870_ ^ _17877_ /*14099*/;
assign _17884_ = D[21] ^ Q[18] /*14095*/;
assign _17881_ = _17345_ & _17884_ /*14091*/;
assign _17882_ = _17345_ ^ _17884_ /*14094*/;
assign _17883_ = _17875_ & _17882_ /*14092*/;
assign _17880_ = _17881_ | _17883_ /*14090*/;
assign _17731_ = _17875_ ^ _17882_ /*14093*/;
assign _17889_ = D[22] ^ Q[18] /*14089*/;
assign _17886_ = _17346_ & _17889_ /*14085*/;
assign _17887_ = _17346_ ^ _17889_ /*14088*/;
assign _17888_ = _17880_ & _17887_ /*14086*/;
assign _17885_ = _17886_ | _17888_ /*14084*/;
assign _17732_ = _17880_ ^ _17887_ /*14087*/;
assign _17894_ = D[23] ^ Q[18] /*14083*/;
assign _17891_ = _17347_ & _17894_ /*14079*/;
assign _17892_ = _17347_ ^ _17894_ /*14082*/;
assign _17893_ = _17885_ & _17892_ /*14080*/;
assign _17890_ = _17891_ | _17893_ /*14078*/;
assign _17733_ = _17885_ ^ _17892_ /*14081*/;
assign _17899_ = D[24] ^ Q[18] /*14077*/;
assign _17896_ = _17348_ & _17899_ /*14073*/;
assign _17897_ = _17348_ ^ _17899_ /*14076*/;
assign _17898_ = _17890_ & _17897_ /*14074*/;
assign _17895_ = _17896_ | _17898_ /*14072*/;
assign _17734_ = _17890_ ^ _17897_ /*14075*/;
assign _17904_ = D[25] ^ Q[18] /*14071*/;
assign _17901_ = _17349_ & _17904_ /*14067*/;
assign _17902_ = _17349_ ^ _17904_ /*14070*/;
assign _17903_ = _17895_ & _17902_ /*14068*/;
assign _17900_ = _17901_ | _17903_ /*14066*/;
assign _17735_ = _17895_ ^ _17902_ /*14069*/;
assign _17909_ = D[26] ^ Q[18] /*14065*/;
assign _17906_ = _17350_ & _17909_ /*14061*/;
assign _17907_ = _17350_ ^ _17909_ /*14064*/;
assign _17908_ = _17900_ & _17907_ /*14062*/;
assign _17905_ = _17906_ | _17908_ /*14060*/;
assign _17736_ = _17900_ ^ _17907_ /*14063*/;
assign _17914_ = D[27] ^ Q[18] /*14059*/;
assign _17911_ = _17351_ & _17914_ /*14055*/;
assign _17912_ = _17351_ ^ _17914_ /*14058*/;
assign _17913_ = _17905_ & _17912_ /*14056*/;
assign _17910_ = _17911_ | _17913_ /*14054*/;
assign _17737_ = _17905_ ^ _17912_ /*14057*/;
assign _17919_ = D[28] ^ Q[18] /*14053*/;
assign _17916_ = _17352_ & _17919_ /*14049*/;
assign _17917_ = _17352_ ^ _17919_ /*14052*/;
assign _17918_ = _17910_ & _17917_ /*14050*/;
assign _17915_ = _17916_ | _17918_ /*14048*/;
assign _17738_ = _17910_ ^ _17917_ /*14051*/;
assign _17924_ = D[29] ^ Q[18] /*14047*/;
assign _17921_ = _17353_ & _17924_ /*14043*/;
assign _17922_ = _17353_ ^ _17924_ /*14046*/;
assign _17923_ = _17915_ & _17922_ /*14044*/;
assign _17920_ = _17921_ | _17923_ /*14042*/;
assign _17739_ = _17915_ ^ _17922_ /*14045*/;
assign _17929_ = D[30] ^ Q[18] /*14041*/;
assign _17926_ = _17354_ & _17929_ /*14037*/;
assign _17927_ = _17354_ ^ _17929_ /*14040*/;
assign _17928_ = _17920_ & _17927_ /*14038*/;
assign _17925_ = _17926_ | _17928_ /*14036*/;
assign _17740_ = _17920_ ^ _17927_ /*14039*/;
assign _17934_ = D[31] ^ Q[18] /*14035*/;
assign _17931_ = _17355_ & _17934_ /*14031*/;
assign _17932_ = _17355_ ^ _17934_ /*14034*/;
assign _17933_ = _17925_ & _17932_ /*14032*/;
assign _17930_ = _17931_ | _17933_ /*14030*/;
assign _17741_ = _17925_ ^ _17932_ /*14033*/;
assign _17939_ = D[32] ^ Q[18] /*14029*/;
assign _17936_ = _17356_ & _17939_ /*14025*/;
assign _17937_ = _17356_ ^ _17939_ /*14028*/;
assign _17938_ = _17930_ & _17937_ /*14026*/;
assign _17935_ = _17936_ | _17938_ /*14024*/;
assign _17742_ = _17930_ ^ _17937_ /*14027*/;
assign _17944_ = D[33] ^ Q[18] /*14023*/;
assign _17941_ = _17357_ & _17944_ /*14019*/;
assign _17942_ = _17357_ ^ _17944_ /*14022*/;
assign _17943_ = _17935_ & _17942_ /*14020*/;
assign _17940_ = _17941_ | _17943_ /*14018*/;
assign _17743_ = _17935_ ^ _17942_ /*14021*/;
assign _17949_ = D[34] ^ Q[18] /*14017*/;
assign _17946_ = _17358_ & _17949_ /*14013*/;
assign _17947_ = _17358_ ^ _17949_ /*14016*/;
assign _17948_ = _17940_ & _17947_ /*14014*/;
assign _17945_ = _17946_ | _17948_ /*14012*/;
assign _17744_ = _17940_ ^ _17947_ /*14015*/;
assign _17954_ = D[35] ^ Q[18] /*14011*/;
assign _17951_ = _17359_ & _17954_ /*14007*/;
assign _17952_ = _17359_ ^ _17954_ /*14010*/;
assign _17953_ = _17945_ & _17952_ /*14008*/;
assign _17950_ = _17951_ | _17953_ /*14006*/;
assign _17745_ = _17945_ ^ _17952_ /*14009*/;
assign _17959_ = D[36] ^ Q[18] /*14005*/;
assign _17956_ = _17360_ & _17959_ /*14001*/;
assign _17957_ = _17360_ ^ _17959_ /*14004*/;
assign _17958_ = _17950_ & _17957_ /*14002*/;
assign _17955_ = _17956_ | _17958_ /*14000*/;
assign _17746_ = _17950_ ^ _17957_ /*14003*/;
assign _17964_ = D[37] ^ Q[18] /*13999*/;
assign _17961_ = _17361_ & _17964_ /*13995*/;
assign _17962_ = _17361_ ^ _17964_ /*13998*/;
assign _17963_ = _17955_ & _17962_ /*13996*/;
assign _17960_ = _17961_ | _17963_ /*13994*/;
assign _17747_ = _17955_ ^ _17962_ /*13997*/;
assign _17969_ = D[38] ^ Q[18] /*13993*/;
assign _17966_ = _17362_ & _17969_ /*13989*/;
assign _17967_ = _17362_ ^ _17969_ /*13992*/;
assign _17968_ = _17960_ & _17967_ /*13990*/;
assign _17965_ = _17966_ | _17968_ /*13988*/;
assign _17748_ = _17960_ ^ _17967_ /*13991*/;
assign _17974_ = D[39] ^ Q[18] /*13987*/;
assign _17971_ = _17363_ & _17974_ /*13983*/;
assign _17972_ = _17363_ ^ _17974_ /*13986*/;
assign _17973_ = _17965_ & _17972_ /*13984*/;
assign _17970_ = _17971_ | _17973_ /*13982*/;
assign _17749_ = _17965_ ^ _17972_ /*13985*/;
assign _17979_ = D[40] ^ Q[18] /*13981*/;
assign _17976_ = _17364_ & _17979_ /*13977*/;
assign _17977_ = _17364_ ^ _17979_ /*13980*/;
assign _17978_ = _17970_ & _17977_ /*13978*/;
assign _17975_ = _17976_ | _17978_ /*13976*/;
assign _17750_ = _17970_ ^ _17977_ /*13979*/;
assign _17984_ = D[41] ^ Q[18] /*13975*/;
assign _17981_ = _17365_ & _17984_ /*13971*/;
assign _17982_ = _17365_ ^ _17984_ /*13974*/;
assign _17983_ = _17975_ & _17982_ /*13972*/;
assign _17980_ = _17981_ | _17983_ /*13970*/;
assign _17751_ = _17975_ ^ _17982_ /*13973*/;
assign _17989_ = D[42] ^ Q[18] /*13969*/;
assign _17986_ = _17366_ & _17989_ /*13965*/;
assign _17987_ = _17366_ ^ _17989_ /*13968*/;
assign _17988_ = _17980_ & _17987_ /*13966*/;
assign _17985_ = _17986_ | _17988_ /*13964*/;
assign _17752_ = _17980_ ^ _17987_ /*13967*/;
assign _17994_ = D[43] ^ Q[18] /*13963*/;
assign _17991_ = _17367_ & _17994_ /*13959*/;
assign _17992_ = _17367_ ^ _17994_ /*13962*/;
assign _17993_ = _17985_ & _17992_ /*13960*/;
assign _17990_ = _17991_ | _17993_ /*13958*/;
assign _17753_ = _17985_ ^ _17992_ /*13961*/;
assign _17999_ = D[44] ^ Q[18] /*13957*/;
assign _17996_ = _17368_ & _17999_ /*13953*/;
assign _17997_ = _17368_ ^ _17999_ /*13956*/;
assign _17998_ = _17990_ & _17997_ /*13954*/;
assign _17995_ = _17996_ | _17998_ /*13952*/;
assign _17754_ = _17990_ ^ _17997_ /*13955*/;
assign _18004_ = D[45] ^ Q[18] /*13951*/;
assign _18001_ = _17369_ & _18004_ /*13947*/;
assign _18002_ = _17369_ ^ _18004_ /*13950*/;
assign _18003_ = _17995_ & _18002_ /*13948*/;
assign _18000_ = _18001_ | _18003_ /*13946*/;
assign _17755_ = _17995_ ^ _18002_ /*13949*/;
assign _18009_ = D[46] ^ Q[18] /*13945*/;
assign _18006_ = _17370_ & _18009_ /*13941*/;
assign _18007_ = _17370_ ^ _18009_ /*13944*/;
assign _18008_ = _18000_ & _18007_ /*13942*/;
assign _18005_ = _18006_ | _18008_ /*13940*/;
assign _17756_ = _18000_ ^ _18007_ /*13943*/;
assign _18014_ = D[47] ^ Q[18] /*13939*/;
assign _18011_ = _17371_ & _18014_ /*13935*/;
assign _18012_ = _17371_ ^ _18014_ /*13938*/;
assign _18013_ = _18005_ & _18012_ /*13936*/;
assign _18010_ = _18011_ | _18013_ /*13934*/;
assign _17757_ = _18005_ ^ _18012_ /*13937*/;
assign _18019_ = D[48] ^ Q[18] /*13933*/;
assign _18016_ = _17372_ & _18019_ /*13929*/;
assign _18017_ = _17372_ ^ _18019_ /*13932*/;
assign _18018_ = _18010_ & _18017_ /*13930*/;
assign _18015_ = _18016_ | _18018_ /*13928*/;
assign _17758_ = _18010_ ^ _18017_ /*13931*/;
assign _18024_ = D[49] ^ Q[18] /*13927*/;
assign _18021_ = _17373_ & _18024_ /*13923*/;
assign _18022_ = _17373_ ^ _18024_ /*13926*/;
assign _18023_ = _18015_ & _18022_ /*13924*/;
assign _18020_ = _18021_ | _18023_ /*13922*/;
assign _17759_ = _18015_ ^ _18022_ /*13925*/;
assign _18029_ = D[50] ^ Q[18] /*13921*/;
assign _18026_ = _17374_ & _18029_ /*13917*/;
assign _18027_ = _17374_ ^ _18029_ /*13920*/;
assign _18028_ = _18020_ & _18027_ /*13918*/;
assign _18025_ = _18026_ | _18028_ /*13916*/;
assign _17760_ = _18020_ ^ _18027_ /*13919*/;
assign _18034_ = D[51] ^ Q[18] /*13915*/;
assign _18031_ = _17375_ & _18034_ /*13911*/;
assign _18032_ = _17375_ ^ _18034_ /*13914*/;
assign _18033_ = _18025_ & _18032_ /*13912*/;
assign _18030_ = _18031_ | _18033_ /*13910*/;
assign _17761_ = _18025_ ^ _18032_ /*13913*/;
assign _18039_ = D[52] ^ Q[18] /*13909*/;
assign _18036_ = _17376_ & _18039_ /*13905*/;
assign _18037_ = _17376_ ^ _18039_ /*13908*/;
assign _18038_ = _18030_ & _18037_ /*13906*/;
assign _18035_ = _18036_ | _18038_ /*13904*/;
assign _17762_ = _18030_ ^ _18037_ /*13907*/;
assign _18044_ = D[53] ^ Q[18] /*13903*/;
assign _18041_ = _17377_ & _18044_ /*13899*/;
assign _18042_ = _17377_ ^ _18044_ /*13902*/;
assign _18043_ = _18035_ & _18042_ /*13900*/;
assign _18040_ = _18041_ | _18043_ /*13898*/;
assign _17763_ = _18035_ ^ _18042_ /*13901*/;
assign _18049_ = D[54] ^ Q[18] /*13897*/;
assign _18046_ = _17378_ & _18049_ /*13893*/;
assign _18047_ = _17378_ ^ _18049_ /*13896*/;
assign _18048_ = _18040_ & _18047_ /*13894*/;
assign _18045_ = _18046_ | _18048_ /*13892*/;
assign _17764_ = _18040_ ^ _18047_ /*13895*/;
assign _18054_ = D[55] ^ Q[18] /*13891*/;
assign _18051_ = _17379_ & _18054_ /*13887*/;
assign _18052_ = _17379_ ^ _18054_ /*13890*/;
assign _18053_ = _18045_ & _18052_ /*13888*/;
assign _18050_ = _18051_ | _18053_ /*13886*/;
assign _17765_ = _18045_ ^ _18052_ /*13889*/;
assign _18059_ = D[56] ^ Q[18] /*13885*/;
assign _18056_ = _17380_ & _18059_ /*13881*/;
assign _18057_ = _17380_ ^ _18059_ /*13884*/;
assign _18058_ = _18050_ & _18057_ /*13882*/;
assign _18055_ = _18056_ | _18058_ /*13880*/;
assign _17766_ = _18050_ ^ _18057_ /*13883*/;
assign _18064_ = D[57] ^ Q[18] /*13879*/;
assign _18061_ = _17381_ & _18064_ /*13875*/;
assign _18062_ = _17381_ ^ _18064_ /*13878*/;
assign _18063_ = _18055_ & _18062_ /*13876*/;
assign _18060_ = _18061_ | _18063_ /*13874*/;
assign _17767_ = _18055_ ^ _18062_ /*13877*/;
assign _18069_ = D[58] ^ Q[18] /*13873*/;
assign _18066_ = _17382_ & _18069_ /*13869*/;
assign _18067_ = _17382_ ^ _18069_ /*13872*/;
assign _18068_ = _18060_ & _18067_ /*13870*/;
assign _18065_ = _18066_ | _18068_ /*13868*/;
assign _17768_ = _18060_ ^ _18067_ /*13871*/;
assign _18074_ = D[59] ^ Q[18] /*13867*/;
assign _18071_ = _17383_ & _18074_ /*13863*/;
assign _18072_ = _17383_ ^ _18074_ /*13866*/;
assign _18073_ = _18065_ & _18072_ /*13864*/;
assign _18070_ = _18071_ | _18073_ /*13862*/;
assign _17769_ = _18065_ ^ _18072_ /*13865*/;
assign _18079_ = D[60] ^ Q[18] /*13861*/;
assign _18076_ = _17384_ & _18079_ /*13857*/;
assign _18077_ = _17384_ ^ _18079_ /*13860*/;
assign _18078_ = _18070_ & _18077_ /*13858*/;
assign _18075_ = _18076_ | _18078_ /*13856*/;
assign _17770_ = _18070_ ^ _18077_ /*13859*/;
assign _18084_ = D[61] ^ Q[18] /*13855*/;
assign _18081_ = _17385_ & _18084_ /*13851*/;
assign _18082_ = _17385_ ^ _18084_ /*13854*/;
assign _18083_ = _18075_ & _18082_ /*13852*/;
assign _18080_ = _18081_ | _18083_ /*13850*/;
assign _17771_ = _18075_ ^ _18082_ /*13853*/;
assign _18089_ = D[62] ^ Q[18] /*13849*/;
assign _18086_ = _17386_ & _18089_ /*13845*/;
assign _18087_ = _17386_ ^ _18089_ /*13848*/;
assign _18088_ = _18080_ & _18087_ /*13846*/;
assign _18085_ = _18086_ | _18088_ /*13844*/;
assign _17772_ = _18080_ ^ _18087_ /*13847*/;
assign _18093_ = zeroWire ^ Q[18] /*13843*/;
assign _18090_ = _17387_ & _18093_ /*13839*/;
assign _18091_ = _17387_ ^ _18093_ /*13842*/;
assign _18092_ = _18085_ & _18091_ /*13840*/;
assign Q[17] = _18090_ | _18092_ /*13838*/;
assign _17773_ = _18085_ ^ _18091_ /*13841*/;
assign _18164_ = D[0] ^ Q[17] /*13452*/;
assign _18161_ = R_0[16] & _18164_ /*13448*/;
assign _18162_ = R_0[16] ^ _18164_ /*13451*/;
assign _18163_ = Q[17] & _18162_ /*13449*/;
assign _18160_ = _18161_ | _18163_ /*13447*/;
assign _18095_ = Q[17] ^ _18162_ /*13450*/;
assign _18169_ = D[1] ^ Q[17] /*13446*/;
assign _18166_ = _17710_ & _18169_ /*13442*/;
assign _18167_ = _17710_ ^ _18169_ /*13445*/;
assign _18168_ = _18160_ & _18167_ /*13443*/;
assign _18165_ = _18166_ | _18168_ /*13441*/;
assign _18096_ = _18160_ ^ _18167_ /*13444*/;
assign _18174_ = D[2] ^ Q[17] /*13440*/;
assign _18171_ = _17711_ & _18174_ /*13436*/;
assign _18172_ = _17711_ ^ _18174_ /*13439*/;
assign _18173_ = _18165_ & _18172_ /*13437*/;
assign _18170_ = _18171_ | _18173_ /*13435*/;
assign _18097_ = _18165_ ^ _18172_ /*13438*/;
assign _18179_ = D[3] ^ Q[17] /*13434*/;
assign _18176_ = _17712_ & _18179_ /*13430*/;
assign _18177_ = _17712_ ^ _18179_ /*13433*/;
assign _18178_ = _18170_ & _18177_ /*13431*/;
assign _18175_ = _18176_ | _18178_ /*13429*/;
assign _18098_ = _18170_ ^ _18177_ /*13432*/;
assign _18184_ = D[4] ^ Q[17] /*13428*/;
assign _18181_ = _17713_ & _18184_ /*13424*/;
assign _18182_ = _17713_ ^ _18184_ /*13427*/;
assign _18183_ = _18175_ & _18182_ /*13425*/;
assign _18180_ = _18181_ | _18183_ /*13423*/;
assign _18099_ = _18175_ ^ _18182_ /*13426*/;
assign _18189_ = D[5] ^ Q[17] /*13422*/;
assign _18186_ = _17714_ & _18189_ /*13418*/;
assign _18187_ = _17714_ ^ _18189_ /*13421*/;
assign _18188_ = _18180_ & _18187_ /*13419*/;
assign _18185_ = _18186_ | _18188_ /*13417*/;
assign _18100_ = _18180_ ^ _18187_ /*13420*/;
assign _18194_ = D[6] ^ Q[17] /*13416*/;
assign _18191_ = _17715_ & _18194_ /*13412*/;
assign _18192_ = _17715_ ^ _18194_ /*13415*/;
assign _18193_ = _18185_ & _18192_ /*13413*/;
assign _18190_ = _18191_ | _18193_ /*13411*/;
assign _18101_ = _18185_ ^ _18192_ /*13414*/;
assign _18199_ = D[7] ^ Q[17] /*13410*/;
assign _18196_ = _17716_ & _18199_ /*13406*/;
assign _18197_ = _17716_ ^ _18199_ /*13409*/;
assign _18198_ = _18190_ & _18197_ /*13407*/;
assign _18195_ = _18196_ | _18198_ /*13405*/;
assign _18102_ = _18190_ ^ _18197_ /*13408*/;
assign _18204_ = D[8] ^ Q[17] /*13404*/;
assign _18201_ = _17717_ & _18204_ /*13400*/;
assign _18202_ = _17717_ ^ _18204_ /*13403*/;
assign _18203_ = _18195_ & _18202_ /*13401*/;
assign _18200_ = _18201_ | _18203_ /*13399*/;
assign _18103_ = _18195_ ^ _18202_ /*13402*/;
assign _18209_ = D[9] ^ Q[17] /*13398*/;
assign _18206_ = _17718_ & _18209_ /*13394*/;
assign _18207_ = _17718_ ^ _18209_ /*13397*/;
assign _18208_ = _18200_ & _18207_ /*13395*/;
assign _18205_ = _18206_ | _18208_ /*13393*/;
assign _18104_ = _18200_ ^ _18207_ /*13396*/;
assign _18214_ = D[10] ^ Q[17] /*13392*/;
assign _18211_ = _17719_ & _18214_ /*13388*/;
assign _18212_ = _17719_ ^ _18214_ /*13391*/;
assign _18213_ = _18205_ & _18212_ /*13389*/;
assign _18210_ = _18211_ | _18213_ /*13387*/;
assign _18105_ = _18205_ ^ _18212_ /*13390*/;
assign _18219_ = D[11] ^ Q[17] /*13386*/;
assign _18216_ = _17720_ & _18219_ /*13382*/;
assign _18217_ = _17720_ ^ _18219_ /*13385*/;
assign _18218_ = _18210_ & _18217_ /*13383*/;
assign _18215_ = _18216_ | _18218_ /*13381*/;
assign _18106_ = _18210_ ^ _18217_ /*13384*/;
assign _18224_ = D[12] ^ Q[17] /*13380*/;
assign _18221_ = _17721_ & _18224_ /*13376*/;
assign _18222_ = _17721_ ^ _18224_ /*13379*/;
assign _18223_ = _18215_ & _18222_ /*13377*/;
assign _18220_ = _18221_ | _18223_ /*13375*/;
assign _18107_ = _18215_ ^ _18222_ /*13378*/;
assign _18229_ = D[13] ^ Q[17] /*13374*/;
assign _18226_ = _17722_ & _18229_ /*13370*/;
assign _18227_ = _17722_ ^ _18229_ /*13373*/;
assign _18228_ = _18220_ & _18227_ /*13371*/;
assign _18225_ = _18226_ | _18228_ /*13369*/;
assign _18108_ = _18220_ ^ _18227_ /*13372*/;
assign _18234_ = D[14] ^ Q[17] /*13368*/;
assign _18231_ = _17723_ & _18234_ /*13364*/;
assign _18232_ = _17723_ ^ _18234_ /*13367*/;
assign _18233_ = _18225_ & _18232_ /*13365*/;
assign _18230_ = _18231_ | _18233_ /*13363*/;
assign _18109_ = _18225_ ^ _18232_ /*13366*/;
assign _18239_ = D[15] ^ Q[17] /*13362*/;
assign _18236_ = _17724_ & _18239_ /*13358*/;
assign _18237_ = _17724_ ^ _18239_ /*13361*/;
assign _18238_ = _18230_ & _18237_ /*13359*/;
assign _18235_ = _18236_ | _18238_ /*13357*/;
assign _18110_ = _18230_ ^ _18237_ /*13360*/;
assign _18244_ = D[16] ^ Q[17] /*13356*/;
assign _18241_ = _17725_ & _18244_ /*13352*/;
assign _18242_ = _17725_ ^ _18244_ /*13355*/;
assign _18243_ = _18235_ & _18242_ /*13353*/;
assign _18240_ = _18241_ | _18243_ /*13351*/;
assign _18111_ = _18235_ ^ _18242_ /*13354*/;
assign _18249_ = D[17] ^ Q[17] /*13350*/;
assign _18246_ = _17726_ & _18249_ /*13346*/;
assign _18247_ = _17726_ ^ _18249_ /*13349*/;
assign _18248_ = _18240_ & _18247_ /*13347*/;
assign _18245_ = _18246_ | _18248_ /*13345*/;
assign _18112_ = _18240_ ^ _18247_ /*13348*/;
assign _18254_ = D[18] ^ Q[17] /*13344*/;
assign _18251_ = _17727_ & _18254_ /*13340*/;
assign _18252_ = _17727_ ^ _18254_ /*13343*/;
assign _18253_ = _18245_ & _18252_ /*13341*/;
assign _18250_ = _18251_ | _18253_ /*13339*/;
assign _18113_ = _18245_ ^ _18252_ /*13342*/;
assign _18259_ = D[19] ^ Q[17] /*13338*/;
assign _18256_ = _17728_ & _18259_ /*13334*/;
assign _18257_ = _17728_ ^ _18259_ /*13337*/;
assign _18258_ = _18250_ & _18257_ /*13335*/;
assign _18255_ = _18256_ | _18258_ /*13333*/;
assign _18114_ = _18250_ ^ _18257_ /*13336*/;
assign _18264_ = D[20] ^ Q[17] /*13332*/;
assign _18261_ = _17729_ & _18264_ /*13328*/;
assign _18262_ = _17729_ ^ _18264_ /*13331*/;
assign _18263_ = _18255_ & _18262_ /*13329*/;
assign _18260_ = _18261_ | _18263_ /*13327*/;
assign _18115_ = _18255_ ^ _18262_ /*13330*/;
assign _18269_ = D[21] ^ Q[17] /*13326*/;
assign _18266_ = _17730_ & _18269_ /*13322*/;
assign _18267_ = _17730_ ^ _18269_ /*13325*/;
assign _18268_ = _18260_ & _18267_ /*13323*/;
assign _18265_ = _18266_ | _18268_ /*13321*/;
assign _18116_ = _18260_ ^ _18267_ /*13324*/;
assign _18274_ = D[22] ^ Q[17] /*13320*/;
assign _18271_ = _17731_ & _18274_ /*13316*/;
assign _18272_ = _17731_ ^ _18274_ /*13319*/;
assign _18273_ = _18265_ & _18272_ /*13317*/;
assign _18270_ = _18271_ | _18273_ /*13315*/;
assign _18117_ = _18265_ ^ _18272_ /*13318*/;
assign _18279_ = D[23] ^ Q[17] /*13314*/;
assign _18276_ = _17732_ & _18279_ /*13310*/;
assign _18277_ = _17732_ ^ _18279_ /*13313*/;
assign _18278_ = _18270_ & _18277_ /*13311*/;
assign _18275_ = _18276_ | _18278_ /*13309*/;
assign _18118_ = _18270_ ^ _18277_ /*13312*/;
assign _18284_ = D[24] ^ Q[17] /*13308*/;
assign _18281_ = _17733_ & _18284_ /*13304*/;
assign _18282_ = _17733_ ^ _18284_ /*13307*/;
assign _18283_ = _18275_ & _18282_ /*13305*/;
assign _18280_ = _18281_ | _18283_ /*13303*/;
assign _18119_ = _18275_ ^ _18282_ /*13306*/;
assign _18289_ = D[25] ^ Q[17] /*13302*/;
assign _18286_ = _17734_ & _18289_ /*13298*/;
assign _18287_ = _17734_ ^ _18289_ /*13301*/;
assign _18288_ = _18280_ & _18287_ /*13299*/;
assign _18285_ = _18286_ | _18288_ /*13297*/;
assign _18120_ = _18280_ ^ _18287_ /*13300*/;
assign _18294_ = D[26] ^ Q[17] /*13296*/;
assign _18291_ = _17735_ & _18294_ /*13292*/;
assign _18292_ = _17735_ ^ _18294_ /*13295*/;
assign _18293_ = _18285_ & _18292_ /*13293*/;
assign _18290_ = _18291_ | _18293_ /*13291*/;
assign _18121_ = _18285_ ^ _18292_ /*13294*/;
assign _18299_ = D[27] ^ Q[17] /*13290*/;
assign _18296_ = _17736_ & _18299_ /*13286*/;
assign _18297_ = _17736_ ^ _18299_ /*13289*/;
assign _18298_ = _18290_ & _18297_ /*13287*/;
assign _18295_ = _18296_ | _18298_ /*13285*/;
assign _18122_ = _18290_ ^ _18297_ /*13288*/;
assign _18304_ = D[28] ^ Q[17] /*13284*/;
assign _18301_ = _17737_ & _18304_ /*13280*/;
assign _18302_ = _17737_ ^ _18304_ /*13283*/;
assign _18303_ = _18295_ & _18302_ /*13281*/;
assign _18300_ = _18301_ | _18303_ /*13279*/;
assign _18123_ = _18295_ ^ _18302_ /*13282*/;
assign _18309_ = D[29] ^ Q[17] /*13278*/;
assign _18306_ = _17738_ & _18309_ /*13274*/;
assign _18307_ = _17738_ ^ _18309_ /*13277*/;
assign _18308_ = _18300_ & _18307_ /*13275*/;
assign _18305_ = _18306_ | _18308_ /*13273*/;
assign _18124_ = _18300_ ^ _18307_ /*13276*/;
assign _18314_ = D[30] ^ Q[17] /*13272*/;
assign _18311_ = _17739_ & _18314_ /*13268*/;
assign _18312_ = _17739_ ^ _18314_ /*13271*/;
assign _18313_ = _18305_ & _18312_ /*13269*/;
assign _18310_ = _18311_ | _18313_ /*13267*/;
assign _18125_ = _18305_ ^ _18312_ /*13270*/;
assign _18319_ = D[31] ^ Q[17] /*13266*/;
assign _18316_ = _17740_ & _18319_ /*13262*/;
assign _18317_ = _17740_ ^ _18319_ /*13265*/;
assign _18318_ = _18310_ & _18317_ /*13263*/;
assign _18315_ = _18316_ | _18318_ /*13261*/;
assign _18126_ = _18310_ ^ _18317_ /*13264*/;
assign _18324_ = D[32] ^ Q[17] /*13260*/;
assign _18321_ = _17741_ & _18324_ /*13256*/;
assign _18322_ = _17741_ ^ _18324_ /*13259*/;
assign _18323_ = _18315_ & _18322_ /*13257*/;
assign _18320_ = _18321_ | _18323_ /*13255*/;
assign _18127_ = _18315_ ^ _18322_ /*13258*/;
assign _18329_ = D[33] ^ Q[17] /*13254*/;
assign _18326_ = _17742_ & _18329_ /*13250*/;
assign _18327_ = _17742_ ^ _18329_ /*13253*/;
assign _18328_ = _18320_ & _18327_ /*13251*/;
assign _18325_ = _18326_ | _18328_ /*13249*/;
assign _18128_ = _18320_ ^ _18327_ /*13252*/;
assign _18334_ = D[34] ^ Q[17] /*13248*/;
assign _18331_ = _17743_ & _18334_ /*13244*/;
assign _18332_ = _17743_ ^ _18334_ /*13247*/;
assign _18333_ = _18325_ & _18332_ /*13245*/;
assign _18330_ = _18331_ | _18333_ /*13243*/;
assign _18129_ = _18325_ ^ _18332_ /*13246*/;
assign _18339_ = D[35] ^ Q[17] /*13242*/;
assign _18336_ = _17744_ & _18339_ /*13238*/;
assign _18337_ = _17744_ ^ _18339_ /*13241*/;
assign _18338_ = _18330_ & _18337_ /*13239*/;
assign _18335_ = _18336_ | _18338_ /*13237*/;
assign _18130_ = _18330_ ^ _18337_ /*13240*/;
assign _18344_ = D[36] ^ Q[17] /*13236*/;
assign _18341_ = _17745_ & _18344_ /*13232*/;
assign _18342_ = _17745_ ^ _18344_ /*13235*/;
assign _18343_ = _18335_ & _18342_ /*13233*/;
assign _18340_ = _18341_ | _18343_ /*13231*/;
assign _18131_ = _18335_ ^ _18342_ /*13234*/;
assign _18349_ = D[37] ^ Q[17] /*13230*/;
assign _18346_ = _17746_ & _18349_ /*13226*/;
assign _18347_ = _17746_ ^ _18349_ /*13229*/;
assign _18348_ = _18340_ & _18347_ /*13227*/;
assign _18345_ = _18346_ | _18348_ /*13225*/;
assign _18132_ = _18340_ ^ _18347_ /*13228*/;
assign _18354_ = D[38] ^ Q[17] /*13224*/;
assign _18351_ = _17747_ & _18354_ /*13220*/;
assign _18352_ = _17747_ ^ _18354_ /*13223*/;
assign _18353_ = _18345_ & _18352_ /*13221*/;
assign _18350_ = _18351_ | _18353_ /*13219*/;
assign _18133_ = _18345_ ^ _18352_ /*13222*/;
assign _18359_ = D[39] ^ Q[17] /*13218*/;
assign _18356_ = _17748_ & _18359_ /*13214*/;
assign _18357_ = _17748_ ^ _18359_ /*13217*/;
assign _18358_ = _18350_ & _18357_ /*13215*/;
assign _18355_ = _18356_ | _18358_ /*13213*/;
assign _18134_ = _18350_ ^ _18357_ /*13216*/;
assign _18364_ = D[40] ^ Q[17] /*13212*/;
assign _18361_ = _17749_ & _18364_ /*13208*/;
assign _18362_ = _17749_ ^ _18364_ /*13211*/;
assign _18363_ = _18355_ & _18362_ /*13209*/;
assign _18360_ = _18361_ | _18363_ /*13207*/;
assign _18135_ = _18355_ ^ _18362_ /*13210*/;
assign _18369_ = D[41] ^ Q[17] /*13206*/;
assign _18366_ = _17750_ & _18369_ /*13202*/;
assign _18367_ = _17750_ ^ _18369_ /*13205*/;
assign _18368_ = _18360_ & _18367_ /*13203*/;
assign _18365_ = _18366_ | _18368_ /*13201*/;
assign _18136_ = _18360_ ^ _18367_ /*13204*/;
assign _18374_ = D[42] ^ Q[17] /*13200*/;
assign _18371_ = _17751_ & _18374_ /*13196*/;
assign _18372_ = _17751_ ^ _18374_ /*13199*/;
assign _18373_ = _18365_ & _18372_ /*13197*/;
assign _18370_ = _18371_ | _18373_ /*13195*/;
assign _18137_ = _18365_ ^ _18372_ /*13198*/;
assign _18379_ = D[43] ^ Q[17] /*13194*/;
assign _18376_ = _17752_ & _18379_ /*13190*/;
assign _18377_ = _17752_ ^ _18379_ /*13193*/;
assign _18378_ = _18370_ & _18377_ /*13191*/;
assign _18375_ = _18376_ | _18378_ /*13189*/;
assign _18138_ = _18370_ ^ _18377_ /*13192*/;
assign _18384_ = D[44] ^ Q[17] /*13188*/;
assign _18381_ = _17753_ & _18384_ /*13184*/;
assign _18382_ = _17753_ ^ _18384_ /*13187*/;
assign _18383_ = _18375_ & _18382_ /*13185*/;
assign _18380_ = _18381_ | _18383_ /*13183*/;
assign _18139_ = _18375_ ^ _18382_ /*13186*/;
assign _18389_ = D[45] ^ Q[17] /*13182*/;
assign _18386_ = _17754_ & _18389_ /*13178*/;
assign _18387_ = _17754_ ^ _18389_ /*13181*/;
assign _18388_ = _18380_ & _18387_ /*13179*/;
assign _18385_ = _18386_ | _18388_ /*13177*/;
assign _18140_ = _18380_ ^ _18387_ /*13180*/;
assign _18394_ = D[46] ^ Q[17] /*13176*/;
assign _18391_ = _17755_ & _18394_ /*13172*/;
assign _18392_ = _17755_ ^ _18394_ /*13175*/;
assign _18393_ = _18385_ & _18392_ /*13173*/;
assign _18390_ = _18391_ | _18393_ /*13171*/;
assign _18141_ = _18385_ ^ _18392_ /*13174*/;
assign _18399_ = D[47] ^ Q[17] /*13170*/;
assign _18396_ = _17756_ & _18399_ /*13166*/;
assign _18397_ = _17756_ ^ _18399_ /*13169*/;
assign _18398_ = _18390_ & _18397_ /*13167*/;
assign _18395_ = _18396_ | _18398_ /*13165*/;
assign _18142_ = _18390_ ^ _18397_ /*13168*/;
assign _18404_ = D[48] ^ Q[17] /*13164*/;
assign _18401_ = _17757_ & _18404_ /*13160*/;
assign _18402_ = _17757_ ^ _18404_ /*13163*/;
assign _18403_ = _18395_ & _18402_ /*13161*/;
assign _18400_ = _18401_ | _18403_ /*13159*/;
assign _18143_ = _18395_ ^ _18402_ /*13162*/;
assign _18409_ = D[49] ^ Q[17] /*13158*/;
assign _18406_ = _17758_ & _18409_ /*13154*/;
assign _18407_ = _17758_ ^ _18409_ /*13157*/;
assign _18408_ = _18400_ & _18407_ /*13155*/;
assign _18405_ = _18406_ | _18408_ /*13153*/;
assign _18144_ = _18400_ ^ _18407_ /*13156*/;
assign _18414_ = D[50] ^ Q[17] /*13152*/;
assign _18411_ = _17759_ & _18414_ /*13148*/;
assign _18412_ = _17759_ ^ _18414_ /*13151*/;
assign _18413_ = _18405_ & _18412_ /*13149*/;
assign _18410_ = _18411_ | _18413_ /*13147*/;
assign _18145_ = _18405_ ^ _18412_ /*13150*/;
assign _18419_ = D[51] ^ Q[17] /*13146*/;
assign _18416_ = _17760_ & _18419_ /*13142*/;
assign _18417_ = _17760_ ^ _18419_ /*13145*/;
assign _18418_ = _18410_ & _18417_ /*13143*/;
assign _18415_ = _18416_ | _18418_ /*13141*/;
assign _18146_ = _18410_ ^ _18417_ /*13144*/;
assign _18424_ = D[52] ^ Q[17] /*13140*/;
assign _18421_ = _17761_ & _18424_ /*13136*/;
assign _18422_ = _17761_ ^ _18424_ /*13139*/;
assign _18423_ = _18415_ & _18422_ /*13137*/;
assign _18420_ = _18421_ | _18423_ /*13135*/;
assign _18147_ = _18415_ ^ _18422_ /*13138*/;
assign _18429_ = D[53] ^ Q[17] /*13134*/;
assign _18426_ = _17762_ & _18429_ /*13130*/;
assign _18427_ = _17762_ ^ _18429_ /*13133*/;
assign _18428_ = _18420_ & _18427_ /*13131*/;
assign _18425_ = _18426_ | _18428_ /*13129*/;
assign _18148_ = _18420_ ^ _18427_ /*13132*/;
assign _18434_ = D[54] ^ Q[17] /*13128*/;
assign _18431_ = _17763_ & _18434_ /*13124*/;
assign _18432_ = _17763_ ^ _18434_ /*13127*/;
assign _18433_ = _18425_ & _18432_ /*13125*/;
assign _18430_ = _18431_ | _18433_ /*13123*/;
assign _18149_ = _18425_ ^ _18432_ /*13126*/;
assign _18439_ = D[55] ^ Q[17] /*13122*/;
assign _18436_ = _17764_ & _18439_ /*13118*/;
assign _18437_ = _17764_ ^ _18439_ /*13121*/;
assign _18438_ = _18430_ & _18437_ /*13119*/;
assign _18435_ = _18436_ | _18438_ /*13117*/;
assign _18150_ = _18430_ ^ _18437_ /*13120*/;
assign _18444_ = D[56] ^ Q[17] /*13116*/;
assign _18441_ = _17765_ & _18444_ /*13112*/;
assign _18442_ = _17765_ ^ _18444_ /*13115*/;
assign _18443_ = _18435_ & _18442_ /*13113*/;
assign _18440_ = _18441_ | _18443_ /*13111*/;
assign _18151_ = _18435_ ^ _18442_ /*13114*/;
assign _18449_ = D[57] ^ Q[17] /*13110*/;
assign _18446_ = _17766_ & _18449_ /*13106*/;
assign _18447_ = _17766_ ^ _18449_ /*13109*/;
assign _18448_ = _18440_ & _18447_ /*13107*/;
assign _18445_ = _18446_ | _18448_ /*13105*/;
assign _18152_ = _18440_ ^ _18447_ /*13108*/;
assign _18454_ = D[58] ^ Q[17] /*13104*/;
assign _18451_ = _17767_ & _18454_ /*13100*/;
assign _18452_ = _17767_ ^ _18454_ /*13103*/;
assign _18453_ = _18445_ & _18452_ /*13101*/;
assign _18450_ = _18451_ | _18453_ /*13099*/;
assign _18153_ = _18445_ ^ _18452_ /*13102*/;
assign _18459_ = D[59] ^ Q[17] /*13098*/;
assign _18456_ = _17768_ & _18459_ /*13094*/;
assign _18457_ = _17768_ ^ _18459_ /*13097*/;
assign _18458_ = _18450_ & _18457_ /*13095*/;
assign _18455_ = _18456_ | _18458_ /*13093*/;
assign _18154_ = _18450_ ^ _18457_ /*13096*/;
assign _18464_ = D[60] ^ Q[17] /*13092*/;
assign _18461_ = _17769_ & _18464_ /*13088*/;
assign _18462_ = _17769_ ^ _18464_ /*13091*/;
assign _18463_ = _18455_ & _18462_ /*13089*/;
assign _18460_ = _18461_ | _18463_ /*13087*/;
assign _18155_ = _18455_ ^ _18462_ /*13090*/;
assign _18469_ = D[61] ^ Q[17] /*13086*/;
assign _18466_ = _17770_ & _18469_ /*13082*/;
assign _18467_ = _17770_ ^ _18469_ /*13085*/;
assign _18468_ = _18460_ & _18467_ /*13083*/;
assign _18465_ = _18466_ | _18468_ /*13081*/;
assign _18156_ = _18460_ ^ _18467_ /*13084*/;
assign _18474_ = D[62] ^ Q[17] /*13080*/;
assign _18471_ = _17771_ & _18474_ /*13076*/;
assign _18472_ = _17771_ ^ _18474_ /*13079*/;
assign _18473_ = _18465_ & _18472_ /*13077*/;
assign _18470_ = _18471_ | _18473_ /*13075*/;
assign _18157_ = _18465_ ^ _18472_ /*13078*/;
assign _18478_ = zeroWire ^ Q[17] /*13074*/;
assign _18475_ = _17772_ & _18478_ /*13070*/;
assign _18476_ = _17772_ ^ _18478_ /*13073*/;
assign _18477_ = _18470_ & _18476_ /*13071*/;
assign Q[16] = _18475_ | _18477_ /*13069*/;
assign _18158_ = _18470_ ^ _18476_ /*13072*/;
assign _18549_ = D[0] ^ Q[16] /*12683*/;
assign _18546_ = R_0[15] & _18549_ /*12679*/;
assign _18547_ = R_0[15] ^ _18549_ /*12682*/;
assign _18548_ = Q[16] & _18547_ /*12680*/;
assign _18545_ = _18546_ | _18548_ /*12678*/;
assign _18480_ = Q[16] ^ _18547_ /*12681*/;
assign _18554_ = D[1] ^ Q[16] /*12677*/;
assign _18551_ = _18095_ & _18554_ /*12673*/;
assign _18552_ = _18095_ ^ _18554_ /*12676*/;
assign _18553_ = _18545_ & _18552_ /*12674*/;
assign _18550_ = _18551_ | _18553_ /*12672*/;
assign _18481_ = _18545_ ^ _18552_ /*12675*/;
assign _18559_ = D[2] ^ Q[16] /*12671*/;
assign _18556_ = _18096_ & _18559_ /*12667*/;
assign _18557_ = _18096_ ^ _18559_ /*12670*/;
assign _18558_ = _18550_ & _18557_ /*12668*/;
assign _18555_ = _18556_ | _18558_ /*12666*/;
assign _18482_ = _18550_ ^ _18557_ /*12669*/;
assign _18564_ = D[3] ^ Q[16] /*12665*/;
assign _18561_ = _18097_ & _18564_ /*12661*/;
assign _18562_ = _18097_ ^ _18564_ /*12664*/;
assign _18563_ = _18555_ & _18562_ /*12662*/;
assign _18560_ = _18561_ | _18563_ /*12660*/;
assign _18483_ = _18555_ ^ _18562_ /*12663*/;
assign _18569_ = D[4] ^ Q[16] /*12659*/;
assign _18566_ = _18098_ & _18569_ /*12655*/;
assign _18567_ = _18098_ ^ _18569_ /*12658*/;
assign _18568_ = _18560_ & _18567_ /*12656*/;
assign _18565_ = _18566_ | _18568_ /*12654*/;
assign _18484_ = _18560_ ^ _18567_ /*12657*/;
assign _18574_ = D[5] ^ Q[16] /*12653*/;
assign _18571_ = _18099_ & _18574_ /*12649*/;
assign _18572_ = _18099_ ^ _18574_ /*12652*/;
assign _18573_ = _18565_ & _18572_ /*12650*/;
assign _18570_ = _18571_ | _18573_ /*12648*/;
assign _18485_ = _18565_ ^ _18572_ /*12651*/;
assign _18579_ = D[6] ^ Q[16] /*12647*/;
assign _18576_ = _18100_ & _18579_ /*12643*/;
assign _18577_ = _18100_ ^ _18579_ /*12646*/;
assign _18578_ = _18570_ & _18577_ /*12644*/;
assign _18575_ = _18576_ | _18578_ /*12642*/;
assign _18486_ = _18570_ ^ _18577_ /*12645*/;
assign _18584_ = D[7] ^ Q[16] /*12641*/;
assign _18581_ = _18101_ & _18584_ /*12637*/;
assign _18582_ = _18101_ ^ _18584_ /*12640*/;
assign _18583_ = _18575_ & _18582_ /*12638*/;
assign _18580_ = _18581_ | _18583_ /*12636*/;
assign _18487_ = _18575_ ^ _18582_ /*12639*/;
assign _18589_ = D[8] ^ Q[16] /*12635*/;
assign _18586_ = _18102_ & _18589_ /*12631*/;
assign _18587_ = _18102_ ^ _18589_ /*12634*/;
assign _18588_ = _18580_ & _18587_ /*12632*/;
assign _18585_ = _18586_ | _18588_ /*12630*/;
assign _18488_ = _18580_ ^ _18587_ /*12633*/;
assign _18594_ = D[9] ^ Q[16] /*12629*/;
assign _18591_ = _18103_ & _18594_ /*12625*/;
assign _18592_ = _18103_ ^ _18594_ /*12628*/;
assign _18593_ = _18585_ & _18592_ /*12626*/;
assign _18590_ = _18591_ | _18593_ /*12624*/;
assign _18489_ = _18585_ ^ _18592_ /*12627*/;
assign _18599_ = D[10] ^ Q[16] /*12623*/;
assign _18596_ = _18104_ & _18599_ /*12619*/;
assign _18597_ = _18104_ ^ _18599_ /*12622*/;
assign _18598_ = _18590_ & _18597_ /*12620*/;
assign _18595_ = _18596_ | _18598_ /*12618*/;
assign _18490_ = _18590_ ^ _18597_ /*12621*/;
assign _18604_ = D[11] ^ Q[16] /*12617*/;
assign _18601_ = _18105_ & _18604_ /*12613*/;
assign _18602_ = _18105_ ^ _18604_ /*12616*/;
assign _18603_ = _18595_ & _18602_ /*12614*/;
assign _18600_ = _18601_ | _18603_ /*12612*/;
assign _18491_ = _18595_ ^ _18602_ /*12615*/;
assign _18609_ = D[12] ^ Q[16] /*12611*/;
assign _18606_ = _18106_ & _18609_ /*12607*/;
assign _18607_ = _18106_ ^ _18609_ /*12610*/;
assign _18608_ = _18600_ & _18607_ /*12608*/;
assign _18605_ = _18606_ | _18608_ /*12606*/;
assign _18492_ = _18600_ ^ _18607_ /*12609*/;
assign _18614_ = D[13] ^ Q[16] /*12605*/;
assign _18611_ = _18107_ & _18614_ /*12601*/;
assign _18612_ = _18107_ ^ _18614_ /*12604*/;
assign _18613_ = _18605_ & _18612_ /*12602*/;
assign _18610_ = _18611_ | _18613_ /*12600*/;
assign _18493_ = _18605_ ^ _18612_ /*12603*/;
assign _18619_ = D[14] ^ Q[16] /*12599*/;
assign _18616_ = _18108_ & _18619_ /*12595*/;
assign _18617_ = _18108_ ^ _18619_ /*12598*/;
assign _18618_ = _18610_ & _18617_ /*12596*/;
assign _18615_ = _18616_ | _18618_ /*12594*/;
assign _18494_ = _18610_ ^ _18617_ /*12597*/;
assign _18624_ = D[15] ^ Q[16] /*12593*/;
assign _18621_ = _18109_ & _18624_ /*12589*/;
assign _18622_ = _18109_ ^ _18624_ /*12592*/;
assign _18623_ = _18615_ & _18622_ /*12590*/;
assign _18620_ = _18621_ | _18623_ /*12588*/;
assign _18495_ = _18615_ ^ _18622_ /*12591*/;
assign _18629_ = D[16] ^ Q[16] /*12587*/;
assign _18626_ = _18110_ & _18629_ /*12583*/;
assign _18627_ = _18110_ ^ _18629_ /*12586*/;
assign _18628_ = _18620_ & _18627_ /*12584*/;
assign _18625_ = _18626_ | _18628_ /*12582*/;
assign _18496_ = _18620_ ^ _18627_ /*12585*/;
assign _18634_ = D[17] ^ Q[16] /*12581*/;
assign _18631_ = _18111_ & _18634_ /*12577*/;
assign _18632_ = _18111_ ^ _18634_ /*12580*/;
assign _18633_ = _18625_ & _18632_ /*12578*/;
assign _18630_ = _18631_ | _18633_ /*12576*/;
assign _18497_ = _18625_ ^ _18632_ /*12579*/;
assign _18639_ = D[18] ^ Q[16] /*12575*/;
assign _18636_ = _18112_ & _18639_ /*12571*/;
assign _18637_ = _18112_ ^ _18639_ /*12574*/;
assign _18638_ = _18630_ & _18637_ /*12572*/;
assign _18635_ = _18636_ | _18638_ /*12570*/;
assign _18498_ = _18630_ ^ _18637_ /*12573*/;
assign _18644_ = D[19] ^ Q[16] /*12569*/;
assign _18641_ = _18113_ & _18644_ /*12565*/;
assign _18642_ = _18113_ ^ _18644_ /*12568*/;
assign _18643_ = _18635_ & _18642_ /*12566*/;
assign _18640_ = _18641_ | _18643_ /*12564*/;
assign _18499_ = _18635_ ^ _18642_ /*12567*/;
assign _18649_ = D[20] ^ Q[16] /*12563*/;
assign _18646_ = _18114_ & _18649_ /*12559*/;
assign _18647_ = _18114_ ^ _18649_ /*12562*/;
assign _18648_ = _18640_ & _18647_ /*12560*/;
assign _18645_ = _18646_ | _18648_ /*12558*/;
assign _18500_ = _18640_ ^ _18647_ /*12561*/;
assign _18654_ = D[21] ^ Q[16] /*12557*/;
assign _18651_ = _18115_ & _18654_ /*12553*/;
assign _18652_ = _18115_ ^ _18654_ /*12556*/;
assign _18653_ = _18645_ & _18652_ /*12554*/;
assign _18650_ = _18651_ | _18653_ /*12552*/;
assign _18501_ = _18645_ ^ _18652_ /*12555*/;
assign _18659_ = D[22] ^ Q[16] /*12551*/;
assign _18656_ = _18116_ & _18659_ /*12547*/;
assign _18657_ = _18116_ ^ _18659_ /*12550*/;
assign _18658_ = _18650_ & _18657_ /*12548*/;
assign _18655_ = _18656_ | _18658_ /*12546*/;
assign _18502_ = _18650_ ^ _18657_ /*12549*/;
assign _18664_ = D[23] ^ Q[16] /*12545*/;
assign _18661_ = _18117_ & _18664_ /*12541*/;
assign _18662_ = _18117_ ^ _18664_ /*12544*/;
assign _18663_ = _18655_ & _18662_ /*12542*/;
assign _18660_ = _18661_ | _18663_ /*12540*/;
assign _18503_ = _18655_ ^ _18662_ /*12543*/;
assign _18669_ = D[24] ^ Q[16] /*12539*/;
assign _18666_ = _18118_ & _18669_ /*12535*/;
assign _18667_ = _18118_ ^ _18669_ /*12538*/;
assign _18668_ = _18660_ & _18667_ /*12536*/;
assign _18665_ = _18666_ | _18668_ /*12534*/;
assign _18504_ = _18660_ ^ _18667_ /*12537*/;
assign _18674_ = D[25] ^ Q[16] /*12533*/;
assign _18671_ = _18119_ & _18674_ /*12529*/;
assign _18672_ = _18119_ ^ _18674_ /*12532*/;
assign _18673_ = _18665_ & _18672_ /*12530*/;
assign _18670_ = _18671_ | _18673_ /*12528*/;
assign _18505_ = _18665_ ^ _18672_ /*12531*/;
assign _18679_ = D[26] ^ Q[16] /*12527*/;
assign _18676_ = _18120_ & _18679_ /*12523*/;
assign _18677_ = _18120_ ^ _18679_ /*12526*/;
assign _18678_ = _18670_ & _18677_ /*12524*/;
assign _18675_ = _18676_ | _18678_ /*12522*/;
assign _18506_ = _18670_ ^ _18677_ /*12525*/;
assign _18684_ = D[27] ^ Q[16] /*12521*/;
assign _18681_ = _18121_ & _18684_ /*12517*/;
assign _18682_ = _18121_ ^ _18684_ /*12520*/;
assign _18683_ = _18675_ & _18682_ /*12518*/;
assign _18680_ = _18681_ | _18683_ /*12516*/;
assign _18507_ = _18675_ ^ _18682_ /*12519*/;
assign _18689_ = D[28] ^ Q[16] /*12515*/;
assign _18686_ = _18122_ & _18689_ /*12511*/;
assign _18687_ = _18122_ ^ _18689_ /*12514*/;
assign _18688_ = _18680_ & _18687_ /*12512*/;
assign _18685_ = _18686_ | _18688_ /*12510*/;
assign _18508_ = _18680_ ^ _18687_ /*12513*/;
assign _18694_ = D[29] ^ Q[16] /*12509*/;
assign _18691_ = _18123_ & _18694_ /*12505*/;
assign _18692_ = _18123_ ^ _18694_ /*12508*/;
assign _18693_ = _18685_ & _18692_ /*12506*/;
assign _18690_ = _18691_ | _18693_ /*12504*/;
assign _18509_ = _18685_ ^ _18692_ /*12507*/;
assign _18699_ = D[30] ^ Q[16] /*12503*/;
assign _18696_ = _18124_ & _18699_ /*12499*/;
assign _18697_ = _18124_ ^ _18699_ /*12502*/;
assign _18698_ = _18690_ & _18697_ /*12500*/;
assign _18695_ = _18696_ | _18698_ /*12498*/;
assign _18510_ = _18690_ ^ _18697_ /*12501*/;
assign _18704_ = D[31] ^ Q[16] /*12497*/;
assign _18701_ = _18125_ & _18704_ /*12493*/;
assign _18702_ = _18125_ ^ _18704_ /*12496*/;
assign _18703_ = _18695_ & _18702_ /*12494*/;
assign _18700_ = _18701_ | _18703_ /*12492*/;
assign _18511_ = _18695_ ^ _18702_ /*12495*/;
assign _18709_ = D[32] ^ Q[16] /*12491*/;
assign _18706_ = _18126_ & _18709_ /*12487*/;
assign _18707_ = _18126_ ^ _18709_ /*12490*/;
assign _18708_ = _18700_ & _18707_ /*12488*/;
assign _18705_ = _18706_ | _18708_ /*12486*/;
assign _18512_ = _18700_ ^ _18707_ /*12489*/;
assign _18714_ = D[33] ^ Q[16] /*12485*/;
assign _18711_ = _18127_ & _18714_ /*12481*/;
assign _18712_ = _18127_ ^ _18714_ /*12484*/;
assign _18713_ = _18705_ & _18712_ /*12482*/;
assign _18710_ = _18711_ | _18713_ /*12480*/;
assign _18513_ = _18705_ ^ _18712_ /*12483*/;
assign _18719_ = D[34] ^ Q[16] /*12479*/;
assign _18716_ = _18128_ & _18719_ /*12475*/;
assign _18717_ = _18128_ ^ _18719_ /*12478*/;
assign _18718_ = _18710_ & _18717_ /*12476*/;
assign _18715_ = _18716_ | _18718_ /*12474*/;
assign _18514_ = _18710_ ^ _18717_ /*12477*/;
assign _18724_ = D[35] ^ Q[16] /*12473*/;
assign _18721_ = _18129_ & _18724_ /*12469*/;
assign _18722_ = _18129_ ^ _18724_ /*12472*/;
assign _18723_ = _18715_ & _18722_ /*12470*/;
assign _18720_ = _18721_ | _18723_ /*12468*/;
assign _18515_ = _18715_ ^ _18722_ /*12471*/;
assign _18729_ = D[36] ^ Q[16] /*12467*/;
assign _18726_ = _18130_ & _18729_ /*12463*/;
assign _18727_ = _18130_ ^ _18729_ /*12466*/;
assign _18728_ = _18720_ & _18727_ /*12464*/;
assign _18725_ = _18726_ | _18728_ /*12462*/;
assign _18516_ = _18720_ ^ _18727_ /*12465*/;
assign _18734_ = D[37] ^ Q[16] /*12461*/;
assign _18731_ = _18131_ & _18734_ /*12457*/;
assign _18732_ = _18131_ ^ _18734_ /*12460*/;
assign _18733_ = _18725_ & _18732_ /*12458*/;
assign _18730_ = _18731_ | _18733_ /*12456*/;
assign _18517_ = _18725_ ^ _18732_ /*12459*/;
assign _18739_ = D[38] ^ Q[16] /*12455*/;
assign _18736_ = _18132_ & _18739_ /*12451*/;
assign _18737_ = _18132_ ^ _18739_ /*12454*/;
assign _18738_ = _18730_ & _18737_ /*12452*/;
assign _18735_ = _18736_ | _18738_ /*12450*/;
assign _18518_ = _18730_ ^ _18737_ /*12453*/;
assign _18744_ = D[39] ^ Q[16] /*12449*/;
assign _18741_ = _18133_ & _18744_ /*12445*/;
assign _18742_ = _18133_ ^ _18744_ /*12448*/;
assign _18743_ = _18735_ & _18742_ /*12446*/;
assign _18740_ = _18741_ | _18743_ /*12444*/;
assign _18519_ = _18735_ ^ _18742_ /*12447*/;
assign _18749_ = D[40] ^ Q[16] /*12443*/;
assign _18746_ = _18134_ & _18749_ /*12439*/;
assign _18747_ = _18134_ ^ _18749_ /*12442*/;
assign _18748_ = _18740_ & _18747_ /*12440*/;
assign _18745_ = _18746_ | _18748_ /*12438*/;
assign _18520_ = _18740_ ^ _18747_ /*12441*/;
assign _18754_ = D[41] ^ Q[16] /*12437*/;
assign _18751_ = _18135_ & _18754_ /*12433*/;
assign _18752_ = _18135_ ^ _18754_ /*12436*/;
assign _18753_ = _18745_ & _18752_ /*12434*/;
assign _18750_ = _18751_ | _18753_ /*12432*/;
assign _18521_ = _18745_ ^ _18752_ /*12435*/;
assign _18759_ = D[42] ^ Q[16] /*12431*/;
assign _18756_ = _18136_ & _18759_ /*12427*/;
assign _18757_ = _18136_ ^ _18759_ /*12430*/;
assign _18758_ = _18750_ & _18757_ /*12428*/;
assign _18755_ = _18756_ | _18758_ /*12426*/;
assign _18522_ = _18750_ ^ _18757_ /*12429*/;
assign _18764_ = D[43] ^ Q[16] /*12425*/;
assign _18761_ = _18137_ & _18764_ /*12421*/;
assign _18762_ = _18137_ ^ _18764_ /*12424*/;
assign _18763_ = _18755_ & _18762_ /*12422*/;
assign _18760_ = _18761_ | _18763_ /*12420*/;
assign _18523_ = _18755_ ^ _18762_ /*12423*/;
assign _18769_ = D[44] ^ Q[16] /*12419*/;
assign _18766_ = _18138_ & _18769_ /*12415*/;
assign _18767_ = _18138_ ^ _18769_ /*12418*/;
assign _18768_ = _18760_ & _18767_ /*12416*/;
assign _18765_ = _18766_ | _18768_ /*12414*/;
assign _18524_ = _18760_ ^ _18767_ /*12417*/;
assign _18774_ = D[45] ^ Q[16] /*12413*/;
assign _18771_ = _18139_ & _18774_ /*12409*/;
assign _18772_ = _18139_ ^ _18774_ /*12412*/;
assign _18773_ = _18765_ & _18772_ /*12410*/;
assign _18770_ = _18771_ | _18773_ /*12408*/;
assign _18525_ = _18765_ ^ _18772_ /*12411*/;
assign _18779_ = D[46] ^ Q[16] /*12407*/;
assign _18776_ = _18140_ & _18779_ /*12403*/;
assign _18777_ = _18140_ ^ _18779_ /*12406*/;
assign _18778_ = _18770_ & _18777_ /*12404*/;
assign _18775_ = _18776_ | _18778_ /*12402*/;
assign _18526_ = _18770_ ^ _18777_ /*12405*/;
assign _18784_ = D[47] ^ Q[16] /*12401*/;
assign _18781_ = _18141_ & _18784_ /*12397*/;
assign _18782_ = _18141_ ^ _18784_ /*12400*/;
assign _18783_ = _18775_ & _18782_ /*12398*/;
assign _18780_ = _18781_ | _18783_ /*12396*/;
assign _18527_ = _18775_ ^ _18782_ /*12399*/;
assign _18789_ = D[48] ^ Q[16] /*12395*/;
assign _18786_ = _18142_ & _18789_ /*12391*/;
assign _18787_ = _18142_ ^ _18789_ /*12394*/;
assign _18788_ = _18780_ & _18787_ /*12392*/;
assign _18785_ = _18786_ | _18788_ /*12390*/;
assign _18528_ = _18780_ ^ _18787_ /*12393*/;
assign _18794_ = D[49] ^ Q[16] /*12389*/;
assign _18791_ = _18143_ & _18794_ /*12385*/;
assign _18792_ = _18143_ ^ _18794_ /*12388*/;
assign _18793_ = _18785_ & _18792_ /*12386*/;
assign _18790_ = _18791_ | _18793_ /*12384*/;
assign _18529_ = _18785_ ^ _18792_ /*12387*/;
assign _18799_ = D[50] ^ Q[16] /*12383*/;
assign _18796_ = _18144_ & _18799_ /*12379*/;
assign _18797_ = _18144_ ^ _18799_ /*12382*/;
assign _18798_ = _18790_ & _18797_ /*12380*/;
assign _18795_ = _18796_ | _18798_ /*12378*/;
assign _18530_ = _18790_ ^ _18797_ /*12381*/;
assign _18804_ = D[51] ^ Q[16] /*12377*/;
assign _18801_ = _18145_ & _18804_ /*12373*/;
assign _18802_ = _18145_ ^ _18804_ /*12376*/;
assign _18803_ = _18795_ & _18802_ /*12374*/;
assign _18800_ = _18801_ | _18803_ /*12372*/;
assign _18531_ = _18795_ ^ _18802_ /*12375*/;
assign _18809_ = D[52] ^ Q[16] /*12371*/;
assign _18806_ = _18146_ & _18809_ /*12367*/;
assign _18807_ = _18146_ ^ _18809_ /*12370*/;
assign _18808_ = _18800_ & _18807_ /*12368*/;
assign _18805_ = _18806_ | _18808_ /*12366*/;
assign _18532_ = _18800_ ^ _18807_ /*12369*/;
assign _18814_ = D[53] ^ Q[16] /*12365*/;
assign _18811_ = _18147_ & _18814_ /*12361*/;
assign _18812_ = _18147_ ^ _18814_ /*12364*/;
assign _18813_ = _18805_ & _18812_ /*12362*/;
assign _18810_ = _18811_ | _18813_ /*12360*/;
assign _18533_ = _18805_ ^ _18812_ /*12363*/;
assign _18819_ = D[54] ^ Q[16] /*12359*/;
assign _18816_ = _18148_ & _18819_ /*12355*/;
assign _18817_ = _18148_ ^ _18819_ /*12358*/;
assign _18818_ = _18810_ & _18817_ /*12356*/;
assign _18815_ = _18816_ | _18818_ /*12354*/;
assign _18534_ = _18810_ ^ _18817_ /*12357*/;
assign _18824_ = D[55] ^ Q[16] /*12353*/;
assign _18821_ = _18149_ & _18824_ /*12349*/;
assign _18822_ = _18149_ ^ _18824_ /*12352*/;
assign _18823_ = _18815_ & _18822_ /*12350*/;
assign _18820_ = _18821_ | _18823_ /*12348*/;
assign _18535_ = _18815_ ^ _18822_ /*12351*/;
assign _18829_ = D[56] ^ Q[16] /*12347*/;
assign _18826_ = _18150_ & _18829_ /*12343*/;
assign _18827_ = _18150_ ^ _18829_ /*12346*/;
assign _18828_ = _18820_ & _18827_ /*12344*/;
assign _18825_ = _18826_ | _18828_ /*12342*/;
assign _18536_ = _18820_ ^ _18827_ /*12345*/;
assign _18834_ = D[57] ^ Q[16] /*12341*/;
assign _18831_ = _18151_ & _18834_ /*12337*/;
assign _18832_ = _18151_ ^ _18834_ /*12340*/;
assign _18833_ = _18825_ & _18832_ /*12338*/;
assign _18830_ = _18831_ | _18833_ /*12336*/;
assign _18537_ = _18825_ ^ _18832_ /*12339*/;
assign _18839_ = D[58] ^ Q[16] /*12335*/;
assign _18836_ = _18152_ & _18839_ /*12331*/;
assign _18837_ = _18152_ ^ _18839_ /*12334*/;
assign _18838_ = _18830_ & _18837_ /*12332*/;
assign _18835_ = _18836_ | _18838_ /*12330*/;
assign _18538_ = _18830_ ^ _18837_ /*12333*/;
assign _18844_ = D[59] ^ Q[16] /*12329*/;
assign _18841_ = _18153_ & _18844_ /*12325*/;
assign _18842_ = _18153_ ^ _18844_ /*12328*/;
assign _18843_ = _18835_ & _18842_ /*12326*/;
assign _18840_ = _18841_ | _18843_ /*12324*/;
assign _18539_ = _18835_ ^ _18842_ /*12327*/;
assign _18849_ = D[60] ^ Q[16] /*12323*/;
assign _18846_ = _18154_ & _18849_ /*12319*/;
assign _18847_ = _18154_ ^ _18849_ /*12322*/;
assign _18848_ = _18840_ & _18847_ /*12320*/;
assign _18845_ = _18846_ | _18848_ /*12318*/;
assign _18540_ = _18840_ ^ _18847_ /*12321*/;
assign _18854_ = D[61] ^ Q[16] /*12317*/;
assign _18851_ = _18155_ & _18854_ /*12313*/;
assign _18852_ = _18155_ ^ _18854_ /*12316*/;
assign _18853_ = _18845_ & _18852_ /*12314*/;
assign _18850_ = _18851_ | _18853_ /*12312*/;
assign _18541_ = _18845_ ^ _18852_ /*12315*/;
assign _18859_ = D[62] ^ Q[16] /*12311*/;
assign _18856_ = _18156_ & _18859_ /*12307*/;
assign _18857_ = _18156_ ^ _18859_ /*12310*/;
assign _18858_ = _18850_ & _18857_ /*12308*/;
assign _18855_ = _18856_ | _18858_ /*12306*/;
assign _18542_ = _18850_ ^ _18857_ /*12309*/;
assign _18863_ = zeroWire ^ Q[16] /*12305*/;
assign _18860_ = _18157_ & _18863_ /*12301*/;
assign _18861_ = _18157_ ^ _18863_ /*12304*/;
assign _18862_ = _18855_ & _18861_ /*12302*/;
assign Q[15] = _18860_ | _18862_ /*12300*/;
assign _18543_ = _18855_ ^ _18861_ /*12303*/;
assign _18934_ = D[0] ^ Q[15] /*11914*/;
assign _18931_ = R_0[14] & _18934_ /*11910*/;
assign _18932_ = R_0[14] ^ _18934_ /*11913*/;
assign _18933_ = Q[15] & _18932_ /*11911*/;
assign _18930_ = _18931_ | _18933_ /*11909*/;
assign _18865_ = Q[15] ^ _18932_ /*11912*/;
assign _18939_ = D[1] ^ Q[15] /*11908*/;
assign _18936_ = _18480_ & _18939_ /*11904*/;
assign _18937_ = _18480_ ^ _18939_ /*11907*/;
assign _18938_ = _18930_ & _18937_ /*11905*/;
assign _18935_ = _18936_ | _18938_ /*11903*/;
assign _18866_ = _18930_ ^ _18937_ /*11906*/;
assign _18944_ = D[2] ^ Q[15] /*11902*/;
assign _18941_ = _18481_ & _18944_ /*11898*/;
assign _18942_ = _18481_ ^ _18944_ /*11901*/;
assign _18943_ = _18935_ & _18942_ /*11899*/;
assign _18940_ = _18941_ | _18943_ /*11897*/;
assign _18867_ = _18935_ ^ _18942_ /*11900*/;
assign _18949_ = D[3] ^ Q[15] /*11896*/;
assign _18946_ = _18482_ & _18949_ /*11892*/;
assign _18947_ = _18482_ ^ _18949_ /*11895*/;
assign _18948_ = _18940_ & _18947_ /*11893*/;
assign _18945_ = _18946_ | _18948_ /*11891*/;
assign _18868_ = _18940_ ^ _18947_ /*11894*/;
assign _18954_ = D[4] ^ Q[15] /*11890*/;
assign _18951_ = _18483_ & _18954_ /*11886*/;
assign _18952_ = _18483_ ^ _18954_ /*11889*/;
assign _18953_ = _18945_ & _18952_ /*11887*/;
assign _18950_ = _18951_ | _18953_ /*11885*/;
assign _18869_ = _18945_ ^ _18952_ /*11888*/;
assign _18959_ = D[5] ^ Q[15] /*11884*/;
assign _18956_ = _18484_ & _18959_ /*11880*/;
assign _18957_ = _18484_ ^ _18959_ /*11883*/;
assign _18958_ = _18950_ & _18957_ /*11881*/;
assign _18955_ = _18956_ | _18958_ /*11879*/;
assign _18870_ = _18950_ ^ _18957_ /*11882*/;
assign _18964_ = D[6] ^ Q[15] /*11878*/;
assign _18961_ = _18485_ & _18964_ /*11874*/;
assign _18962_ = _18485_ ^ _18964_ /*11877*/;
assign _18963_ = _18955_ & _18962_ /*11875*/;
assign _18960_ = _18961_ | _18963_ /*11873*/;
assign _18871_ = _18955_ ^ _18962_ /*11876*/;
assign _18969_ = D[7] ^ Q[15] /*11872*/;
assign _18966_ = _18486_ & _18969_ /*11868*/;
assign _18967_ = _18486_ ^ _18969_ /*11871*/;
assign _18968_ = _18960_ & _18967_ /*11869*/;
assign _18965_ = _18966_ | _18968_ /*11867*/;
assign _18872_ = _18960_ ^ _18967_ /*11870*/;
assign _18974_ = D[8] ^ Q[15] /*11866*/;
assign _18971_ = _18487_ & _18974_ /*11862*/;
assign _18972_ = _18487_ ^ _18974_ /*11865*/;
assign _18973_ = _18965_ & _18972_ /*11863*/;
assign _18970_ = _18971_ | _18973_ /*11861*/;
assign _18873_ = _18965_ ^ _18972_ /*11864*/;
assign _18979_ = D[9] ^ Q[15] /*11860*/;
assign _18976_ = _18488_ & _18979_ /*11856*/;
assign _18977_ = _18488_ ^ _18979_ /*11859*/;
assign _18978_ = _18970_ & _18977_ /*11857*/;
assign _18975_ = _18976_ | _18978_ /*11855*/;
assign _18874_ = _18970_ ^ _18977_ /*11858*/;
assign _18984_ = D[10] ^ Q[15] /*11854*/;
assign _18981_ = _18489_ & _18984_ /*11850*/;
assign _18982_ = _18489_ ^ _18984_ /*11853*/;
assign _18983_ = _18975_ & _18982_ /*11851*/;
assign _18980_ = _18981_ | _18983_ /*11849*/;
assign _18875_ = _18975_ ^ _18982_ /*11852*/;
assign _18989_ = D[11] ^ Q[15] /*11848*/;
assign _18986_ = _18490_ & _18989_ /*11844*/;
assign _18987_ = _18490_ ^ _18989_ /*11847*/;
assign _18988_ = _18980_ & _18987_ /*11845*/;
assign _18985_ = _18986_ | _18988_ /*11843*/;
assign _18876_ = _18980_ ^ _18987_ /*11846*/;
assign _18994_ = D[12] ^ Q[15] /*11842*/;
assign _18991_ = _18491_ & _18994_ /*11838*/;
assign _18992_ = _18491_ ^ _18994_ /*11841*/;
assign _18993_ = _18985_ & _18992_ /*11839*/;
assign _18990_ = _18991_ | _18993_ /*11837*/;
assign _18877_ = _18985_ ^ _18992_ /*11840*/;
assign _18999_ = D[13] ^ Q[15] /*11836*/;
assign _18996_ = _18492_ & _18999_ /*11832*/;
assign _18997_ = _18492_ ^ _18999_ /*11835*/;
assign _18998_ = _18990_ & _18997_ /*11833*/;
assign _18995_ = _18996_ | _18998_ /*11831*/;
assign _18878_ = _18990_ ^ _18997_ /*11834*/;
assign _19004_ = D[14] ^ Q[15] /*11830*/;
assign _19001_ = _18493_ & _19004_ /*11826*/;
assign _19002_ = _18493_ ^ _19004_ /*11829*/;
assign _19003_ = _18995_ & _19002_ /*11827*/;
assign _19000_ = _19001_ | _19003_ /*11825*/;
assign _18879_ = _18995_ ^ _19002_ /*11828*/;
assign _19009_ = D[15] ^ Q[15] /*11824*/;
assign _19006_ = _18494_ & _19009_ /*11820*/;
assign _19007_ = _18494_ ^ _19009_ /*11823*/;
assign _19008_ = _19000_ & _19007_ /*11821*/;
assign _19005_ = _19006_ | _19008_ /*11819*/;
assign _18880_ = _19000_ ^ _19007_ /*11822*/;
assign _19014_ = D[16] ^ Q[15] /*11818*/;
assign _19011_ = _18495_ & _19014_ /*11814*/;
assign _19012_ = _18495_ ^ _19014_ /*11817*/;
assign _19013_ = _19005_ & _19012_ /*11815*/;
assign _19010_ = _19011_ | _19013_ /*11813*/;
assign _18881_ = _19005_ ^ _19012_ /*11816*/;
assign _19019_ = D[17] ^ Q[15] /*11812*/;
assign _19016_ = _18496_ & _19019_ /*11808*/;
assign _19017_ = _18496_ ^ _19019_ /*11811*/;
assign _19018_ = _19010_ & _19017_ /*11809*/;
assign _19015_ = _19016_ | _19018_ /*11807*/;
assign _18882_ = _19010_ ^ _19017_ /*11810*/;
assign _19024_ = D[18] ^ Q[15] /*11806*/;
assign _19021_ = _18497_ & _19024_ /*11802*/;
assign _19022_ = _18497_ ^ _19024_ /*11805*/;
assign _19023_ = _19015_ & _19022_ /*11803*/;
assign _19020_ = _19021_ | _19023_ /*11801*/;
assign _18883_ = _19015_ ^ _19022_ /*11804*/;
assign _19029_ = D[19] ^ Q[15] /*11800*/;
assign _19026_ = _18498_ & _19029_ /*11796*/;
assign _19027_ = _18498_ ^ _19029_ /*11799*/;
assign _19028_ = _19020_ & _19027_ /*11797*/;
assign _19025_ = _19026_ | _19028_ /*11795*/;
assign _18884_ = _19020_ ^ _19027_ /*11798*/;
assign _19034_ = D[20] ^ Q[15] /*11794*/;
assign _19031_ = _18499_ & _19034_ /*11790*/;
assign _19032_ = _18499_ ^ _19034_ /*11793*/;
assign _19033_ = _19025_ & _19032_ /*11791*/;
assign _19030_ = _19031_ | _19033_ /*11789*/;
assign _18885_ = _19025_ ^ _19032_ /*11792*/;
assign _19039_ = D[21] ^ Q[15] /*11788*/;
assign _19036_ = _18500_ & _19039_ /*11784*/;
assign _19037_ = _18500_ ^ _19039_ /*11787*/;
assign _19038_ = _19030_ & _19037_ /*11785*/;
assign _19035_ = _19036_ | _19038_ /*11783*/;
assign _18886_ = _19030_ ^ _19037_ /*11786*/;
assign _19044_ = D[22] ^ Q[15] /*11782*/;
assign _19041_ = _18501_ & _19044_ /*11778*/;
assign _19042_ = _18501_ ^ _19044_ /*11781*/;
assign _19043_ = _19035_ & _19042_ /*11779*/;
assign _19040_ = _19041_ | _19043_ /*11777*/;
assign _18887_ = _19035_ ^ _19042_ /*11780*/;
assign _19049_ = D[23] ^ Q[15] /*11776*/;
assign _19046_ = _18502_ & _19049_ /*11772*/;
assign _19047_ = _18502_ ^ _19049_ /*11775*/;
assign _19048_ = _19040_ & _19047_ /*11773*/;
assign _19045_ = _19046_ | _19048_ /*11771*/;
assign _18888_ = _19040_ ^ _19047_ /*11774*/;
assign _19054_ = D[24] ^ Q[15] /*11770*/;
assign _19051_ = _18503_ & _19054_ /*11766*/;
assign _19052_ = _18503_ ^ _19054_ /*11769*/;
assign _19053_ = _19045_ & _19052_ /*11767*/;
assign _19050_ = _19051_ | _19053_ /*11765*/;
assign _18889_ = _19045_ ^ _19052_ /*11768*/;
assign _19059_ = D[25] ^ Q[15] /*11764*/;
assign _19056_ = _18504_ & _19059_ /*11760*/;
assign _19057_ = _18504_ ^ _19059_ /*11763*/;
assign _19058_ = _19050_ & _19057_ /*11761*/;
assign _19055_ = _19056_ | _19058_ /*11759*/;
assign _18890_ = _19050_ ^ _19057_ /*11762*/;
assign _19064_ = D[26] ^ Q[15] /*11758*/;
assign _19061_ = _18505_ & _19064_ /*11754*/;
assign _19062_ = _18505_ ^ _19064_ /*11757*/;
assign _19063_ = _19055_ & _19062_ /*11755*/;
assign _19060_ = _19061_ | _19063_ /*11753*/;
assign _18891_ = _19055_ ^ _19062_ /*11756*/;
assign _19069_ = D[27] ^ Q[15] /*11752*/;
assign _19066_ = _18506_ & _19069_ /*11748*/;
assign _19067_ = _18506_ ^ _19069_ /*11751*/;
assign _19068_ = _19060_ & _19067_ /*11749*/;
assign _19065_ = _19066_ | _19068_ /*11747*/;
assign _18892_ = _19060_ ^ _19067_ /*11750*/;
assign _19074_ = D[28] ^ Q[15] /*11746*/;
assign _19071_ = _18507_ & _19074_ /*11742*/;
assign _19072_ = _18507_ ^ _19074_ /*11745*/;
assign _19073_ = _19065_ & _19072_ /*11743*/;
assign _19070_ = _19071_ | _19073_ /*11741*/;
assign _18893_ = _19065_ ^ _19072_ /*11744*/;
assign _19079_ = D[29] ^ Q[15] /*11740*/;
assign _19076_ = _18508_ & _19079_ /*11736*/;
assign _19077_ = _18508_ ^ _19079_ /*11739*/;
assign _19078_ = _19070_ & _19077_ /*11737*/;
assign _19075_ = _19076_ | _19078_ /*11735*/;
assign _18894_ = _19070_ ^ _19077_ /*11738*/;
assign _19084_ = D[30] ^ Q[15] /*11734*/;
assign _19081_ = _18509_ & _19084_ /*11730*/;
assign _19082_ = _18509_ ^ _19084_ /*11733*/;
assign _19083_ = _19075_ & _19082_ /*11731*/;
assign _19080_ = _19081_ | _19083_ /*11729*/;
assign _18895_ = _19075_ ^ _19082_ /*11732*/;
assign _19089_ = D[31] ^ Q[15] /*11728*/;
assign _19086_ = _18510_ & _19089_ /*11724*/;
assign _19087_ = _18510_ ^ _19089_ /*11727*/;
assign _19088_ = _19080_ & _19087_ /*11725*/;
assign _19085_ = _19086_ | _19088_ /*11723*/;
assign _18896_ = _19080_ ^ _19087_ /*11726*/;
assign _19094_ = D[32] ^ Q[15] /*11722*/;
assign _19091_ = _18511_ & _19094_ /*11718*/;
assign _19092_ = _18511_ ^ _19094_ /*11721*/;
assign _19093_ = _19085_ & _19092_ /*11719*/;
assign _19090_ = _19091_ | _19093_ /*11717*/;
assign _18897_ = _19085_ ^ _19092_ /*11720*/;
assign _19099_ = D[33] ^ Q[15] /*11716*/;
assign _19096_ = _18512_ & _19099_ /*11712*/;
assign _19097_ = _18512_ ^ _19099_ /*11715*/;
assign _19098_ = _19090_ & _19097_ /*11713*/;
assign _19095_ = _19096_ | _19098_ /*11711*/;
assign _18898_ = _19090_ ^ _19097_ /*11714*/;
assign _19104_ = D[34] ^ Q[15] /*11710*/;
assign _19101_ = _18513_ & _19104_ /*11706*/;
assign _19102_ = _18513_ ^ _19104_ /*11709*/;
assign _19103_ = _19095_ & _19102_ /*11707*/;
assign _19100_ = _19101_ | _19103_ /*11705*/;
assign _18899_ = _19095_ ^ _19102_ /*11708*/;
assign _19109_ = D[35] ^ Q[15] /*11704*/;
assign _19106_ = _18514_ & _19109_ /*11700*/;
assign _19107_ = _18514_ ^ _19109_ /*11703*/;
assign _19108_ = _19100_ & _19107_ /*11701*/;
assign _19105_ = _19106_ | _19108_ /*11699*/;
assign _18900_ = _19100_ ^ _19107_ /*11702*/;
assign _19114_ = D[36] ^ Q[15] /*11698*/;
assign _19111_ = _18515_ & _19114_ /*11694*/;
assign _19112_ = _18515_ ^ _19114_ /*11697*/;
assign _19113_ = _19105_ & _19112_ /*11695*/;
assign _19110_ = _19111_ | _19113_ /*11693*/;
assign _18901_ = _19105_ ^ _19112_ /*11696*/;
assign _19119_ = D[37] ^ Q[15] /*11692*/;
assign _19116_ = _18516_ & _19119_ /*11688*/;
assign _19117_ = _18516_ ^ _19119_ /*11691*/;
assign _19118_ = _19110_ & _19117_ /*11689*/;
assign _19115_ = _19116_ | _19118_ /*11687*/;
assign _18902_ = _19110_ ^ _19117_ /*11690*/;
assign _19124_ = D[38] ^ Q[15] /*11686*/;
assign _19121_ = _18517_ & _19124_ /*11682*/;
assign _19122_ = _18517_ ^ _19124_ /*11685*/;
assign _19123_ = _19115_ & _19122_ /*11683*/;
assign _19120_ = _19121_ | _19123_ /*11681*/;
assign _18903_ = _19115_ ^ _19122_ /*11684*/;
assign _19129_ = D[39] ^ Q[15] /*11680*/;
assign _19126_ = _18518_ & _19129_ /*11676*/;
assign _19127_ = _18518_ ^ _19129_ /*11679*/;
assign _19128_ = _19120_ & _19127_ /*11677*/;
assign _19125_ = _19126_ | _19128_ /*11675*/;
assign _18904_ = _19120_ ^ _19127_ /*11678*/;
assign _19134_ = D[40] ^ Q[15] /*11674*/;
assign _19131_ = _18519_ & _19134_ /*11670*/;
assign _19132_ = _18519_ ^ _19134_ /*11673*/;
assign _19133_ = _19125_ & _19132_ /*11671*/;
assign _19130_ = _19131_ | _19133_ /*11669*/;
assign _18905_ = _19125_ ^ _19132_ /*11672*/;
assign _19139_ = D[41] ^ Q[15] /*11668*/;
assign _19136_ = _18520_ & _19139_ /*11664*/;
assign _19137_ = _18520_ ^ _19139_ /*11667*/;
assign _19138_ = _19130_ & _19137_ /*11665*/;
assign _19135_ = _19136_ | _19138_ /*11663*/;
assign _18906_ = _19130_ ^ _19137_ /*11666*/;
assign _19144_ = D[42] ^ Q[15] /*11662*/;
assign _19141_ = _18521_ & _19144_ /*11658*/;
assign _19142_ = _18521_ ^ _19144_ /*11661*/;
assign _19143_ = _19135_ & _19142_ /*11659*/;
assign _19140_ = _19141_ | _19143_ /*11657*/;
assign _18907_ = _19135_ ^ _19142_ /*11660*/;
assign _19149_ = D[43] ^ Q[15] /*11656*/;
assign _19146_ = _18522_ & _19149_ /*11652*/;
assign _19147_ = _18522_ ^ _19149_ /*11655*/;
assign _19148_ = _19140_ & _19147_ /*11653*/;
assign _19145_ = _19146_ | _19148_ /*11651*/;
assign _18908_ = _19140_ ^ _19147_ /*11654*/;
assign _19154_ = D[44] ^ Q[15] /*11650*/;
assign _19151_ = _18523_ & _19154_ /*11646*/;
assign _19152_ = _18523_ ^ _19154_ /*11649*/;
assign _19153_ = _19145_ & _19152_ /*11647*/;
assign _19150_ = _19151_ | _19153_ /*11645*/;
assign _18909_ = _19145_ ^ _19152_ /*11648*/;
assign _19159_ = D[45] ^ Q[15] /*11644*/;
assign _19156_ = _18524_ & _19159_ /*11640*/;
assign _19157_ = _18524_ ^ _19159_ /*11643*/;
assign _19158_ = _19150_ & _19157_ /*11641*/;
assign _19155_ = _19156_ | _19158_ /*11639*/;
assign _18910_ = _19150_ ^ _19157_ /*11642*/;
assign _19164_ = D[46] ^ Q[15] /*11638*/;
assign _19161_ = _18525_ & _19164_ /*11634*/;
assign _19162_ = _18525_ ^ _19164_ /*11637*/;
assign _19163_ = _19155_ & _19162_ /*11635*/;
assign _19160_ = _19161_ | _19163_ /*11633*/;
assign _18911_ = _19155_ ^ _19162_ /*11636*/;
assign _19169_ = D[47] ^ Q[15] /*11632*/;
assign _19166_ = _18526_ & _19169_ /*11628*/;
assign _19167_ = _18526_ ^ _19169_ /*11631*/;
assign _19168_ = _19160_ & _19167_ /*11629*/;
assign _19165_ = _19166_ | _19168_ /*11627*/;
assign _18912_ = _19160_ ^ _19167_ /*11630*/;
assign _19174_ = D[48] ^ Q[15] /*11626*/;
assign _19171_ = _18527_ & _19174_ /*11622*/;
assign _19172_ = _18527_ ^ _19174_ /*11625*/;
assign _19173_ = _19165_ & _19172_ /*11623*/;
assign _19170_ = _19171_ | _19173_ /*11621*/;
assign _18913_ = _19165_ ^ _19172_ /*11624*/;
assign _19179_ = D[49] ^ Q[15] /*11620*/;
assign _19176_ = _18528_ & _19179_ /*11616*/;
assign _19177_ = _18528_ ^ _19179_ /*11619*/;
assign _19178_ = _19170_ & _19177_ /*11617*/;
assign _19175_ = _19176_ | _19178_ /*11615*/;
assign _18914_ = _19170_ ^ _19177_ /*11618*/;
assign _19184_ = D[50] ^ Q[15] /*11614*/;
assign _19181_ = _18529_ & _19184_ /*11610*/;
assign _19182_ = _18529_ ^ _19184_ /*11613*/;
assign _19183_ = _19175_ & _19182_ /*11611*/;
assign _19180_ = _19181_ | _19183_ /*11609*/;
assign _18915_ = _19175_ ^ _19182_ /*11612*/;
assign _19189_ = D[51] ^ Q[15] /*11608*/;
assign _19186_ = _18530_ & _19189_ /*11604*/;
assign _19187_ = _18530_ ^ _19189_ /*11607*/;
assign _19188_ = _19180_ & _19187_ /*11605*/;
assign _19185_ = _19186_ | _19188_ /*11603*/;
assign _18916_ = _19180_ ^ _19187_ /*11606*/;
assign _19194_ = D[52] ^ Q[15] /*11602*/;
assign _19191_ = _18531_ & _19194_ /*11598*/;
assign _19192_ = _18531_ ^ _19194_ /*11601*/;
assign _19193_ = _19185_ & _19192_ /*11599*/;
assign _19190_ = _19191_ | _19193_ /*11597*/;
assign _18917_ = _19185_ ^ _19192_ /*11600*/;
assign _19199_ = D[53] ^ Q[15] /*11596*/;
assign _19196_ = _18532_ & _19199_ /*11592*/;
assign _19197_ = _18532_ ^ _19199_ /*11595*/;
assign _19198_ = _19190_ & _19197_ /*11593*/;
assign _19195_ = _19196_ | _19198_ /*11591*/;
assign _18918_ = _19190_ ^ _19197_ /*11594*/;
assign _19204_ = D[54] ^ Q[15] /*11590*/;
assign _19201_ = _18533_ & _19204_ /*11586*/;
assign _19202_ = _18533_ ^ _19204_ /*11589*/;
assign _19203_ = _19195_ & _19202_ /*11587*/;
assign _19200_ = _19201_ | _19203_ /*11585*/;
assign _18919_ = _19195_ ^ _19202_ /*11588*/;
assign _19209_ = D[55] ^ Q[15] /*11584*/;
assign _19206_ = _18534_ & _19209_ /*11580*/;
assign _19207_ = _18534_ ^ _19209_ /*11583*/;
assign _19208_ = _19200_ & _19207_ /*11581*/;
assign _19205_ = _19206_ | _19208_ /*11579*/;
assign _18920_ = _19200_ ^ _19207_ /*11582*/;
assign _19214_ = D[56] ^ Q[15] /*11578*/;
assign _19211_ = _18535_ & _19214_ /*11574*/;
assign _19212_ = _18535_ ^ _19214_ /*11577*/;
assign _19213_ = _19205_ & _19212_ /*11575*/;
assign _19210_ = _19211_ | _19213_ /*11573*/;
assign _18921_ = _19205_ ^ _19212_ /*11576*/;
assign _19219_ = D[57] ^ Q[15] /*11572*/;
assign _19216_ = _18536_ & _19219_ /*11568*/;
assign _19217_ = _18536_ ^ _19219_ /*11571*/;
assign _19218_ = _19210_ & _19217_ /*11569*/;
assign _19215_ = _19216_ | _19218_ /*11567*/;
assign _18922_ = _19210_ ^ _19217_ /*11570*/;
assign _19224_ = D[58] ^ Q[15] /*11566*/;
assign _19221_ = _18537_ & _19224_ /*11562*/;
assign _19222_ = _18537_ ^ _19224_ /*11565*/;
assign _19223_ = _19215_ & _19222_ /*11563*/;
assign _19220_ = _19221_ | _19223_ /*11561*/;
assign _18923_ = _19215_ ^ _19222_ /*11564*/;
assign _19229_ = D[59] ^ Q[15] /*11560*/;
assign _19226_ = _18538_ & _19229_ /*11556*/;
assign _19227_ = _18538_ ^ _19229_ /*11559*/;
assign _19228_ = _19220_ & _19227_ /*11557*/;
assign _19225_ = _19226_ | _19228_ /*11555*/;
assign _18924_ = _19220_ ^ _19227_ /*11558*/;
assign _19234_ = D[60] ^ Q[15] /*11554*/;
assign _19231_ = _18539_ & _19234_ /*11550*/;
assign _19232_ = _18539_ ^ _19234_ /*11553*/;
assign _19233_ = _19225_ & _19232_ /*11551*/;
assign _19230_ = _19231_ | _19233_ /*11549*/;
assign _18925_ = _19225_ ^ _19232_ /*11552*/;
assign _19239_ = D[61] ^ Q[15] /*11548*/;
assign _19236_ = _18540_ & _19239_ /*11544*/;
assign _19237_ = _18540_ ^ _19239_ /*11547*/;
assign _19238_ = _19230_ & _19237_ /*11545*/;
assign _19235_ = _19236_ | _19238_ /*11543*/;
assign _18926_ = _19230_ ^ _19237_ /*11546*/;
assign _19244_ = D[62] ^ Q[15] /*11542*/;
assign _19241_ = _18541_ & _19244_ /*11538*/;
assign _19242_ = _18541_ ^ _19244_ /*11541*/;
assign _19243_ = _19235_ & _19242_ /*11539*/;
assign _19240_ = _19241_ | _19243_ /*11537*/;
assign _18927_ = _19235_ ^ _19242_ /*11540*/;
assign _19248_ = zeroWire ^ Q[15] /*11536*/;
assign _19245_ = _18542_ & _19248_ /*11532*/;
assign _19246_ = _18542_ ^ _19248_ /*11535*/;
assign _19247_ = _19240_ & _19246_ /*11533*/;
assign Q[14] = _19245_ | _19247_ /*11531*/;
assign _18928_ = _19240_ ^ _19246_ /*11534*/;
assign _19319_ = D[0] ^ Q[14] /*11145*/;
assign _19316_ = R_0[13] & _19319_ /*11141*/;
assign _19317_ = R_0[13] ^ _19319_ /*11144*/;
assign _19318_ = Q[14] & _19317_ /*11142*/;
assign _19315_ = _19316_ | _19318_ /*11140*/;
assign _19250_ = Q[14] ^ _19317_ /*11143*/;
assign _19324_ = D[1] ^ Q[14] /*11139*/;
assign _19321_ = _18865_ & _19324_ /*11135*/;
assign _19322_ = _18865_ ^ _19324_ /*11138*/;
assign _19323_ = _19315_ & _19322_ /*11136*/;
assign _19320_ = _19321_ | _19323_ /*11134*/;
assign _19251_ = _19315_ ^ _19322_ /*11137*/;
assign _19329_ = D[2] ^ Q[14] /*11133*/;
assign _19326_ = _18866_ & _19329_ /*11129*/;
assign _19327_ = _18866_ ^ _19329_ /*11132*/;
assign _19328_ = _19320_ & _19327_ /*11130*/;
assign _19325_ = _19326_ | _19328_ /*11128*/;
assign _19252_ = _19320_ ^ _19327_ /*11131*/;
assign _19334_ = D[3] ^ Q[14] /*11127*/;
assign _19331_ = _18867_ & _19334_ /*11123*/;
assign _19332_ = _18867_ ^ _19334_ /*11126*/;
assign _19333_ = _19325_ & _19332_ /*11124*/;
assign _19330_ = _19331_ | _19333_ /*11122*/;
assign _19253_ = _19325_ ^ _19332_ /*11125*/;
assign _19339_ = D[4] ^ Q[14] /*11121*/;
assign _19336_ = _18868_ & _19339_ /*11117*/;
assign _19337_ = _18868_ ^ _19339_ /*11120*/;
assign _19338_ = _19330_ & _19337_ /*11118*/;
assign _19335_ = _19336_ | _19338_ /*11116*/;
assign _19254_ = _19330_ ^ _19337_ /*11119*/;
assign _19344_ = D[5] ^ Q[14] /*11115*/;
assign _19341_ = _18869_ & _19344_ /*11111*/;
assign _19342_ = _18869_ ^ _19344_ /*11114*/;
assign _19343_ = _19335_ & _19342_ /*11112*/;
assign _19340_ = _19341_ | _19343_ /*11110*/;
assign _19255_ = _19335_ ^ _19342_ /*11113*/;
assign _19349_ = D[6] ^ Q[14] /*11109*/;
assign _19346_ = _18870_ & _19349_ /*11105*/;
assign _19347_ = _18870_ ^ _19349_ /*11108*/;
assign _19348_ = _19340_ & _19347_ /*11106*/;
assign _19345_ = _19346_ | _19348_ /*11104*/;
assign _19256_ = _19340_ ^ _19347_ /*11107*/;
assign _19354_ = D[7] ^ Q[14] /*11103*/;
assign _19351_ = _18871_ & _19354_ /*11099*/;
assign _19352_ = _18871_ ^ _19354_ /*11102*/;
assign _19353_ = _19345_ & _19352_ /*11100*/;
assign _19350_ = _19351_ | _19353_ /*11098*/;
assign _19257_ = _19345_ ^ _19352_ /*11101*/;
assign _19359_ = D[8] ^ Q[14] /*11097*/;
assign _19356_ = _18872_ & _19359_ /*11093*/;
assign _19357_ = _18872_ ^ _19359_ /*11096*/;
assign _19358_ = _19350_ & _19357_ /*11094*/;
assign _19355_ = _19356_ | _19358_ /*11092*/;
assign _19258_ = _19350_ ^ _19357_ /*11095*/;
assign _19364_ = D[9] ^ Q[14] /*11091*/;
assign _19361_ = _18873_ & _19364_ /*11087*/;
assign _19362_ = _18873_ ^ _19364_ /*11090*/;
assign _19363_ = _19355_ & _19362_ /*11088*/;
assign _19360_ = _19361_ | _19363_ /*11086*/;
assign _19259_ = _19355_ ^ _19362_ /*11089*/;
assign _19369_ = D[10] ^ Q[14] /*11085*/;
assign _19366_ = _18874_ & _19369_ /*11081*/;
assign _19367_ = _18874_ ^ _19369_ /*11084*/;
assign _19368_ = _19360_ & _19367_ /*11082*/;
assign _19365_ = _19366_ | _19368_ /*11080*/;
assign _19260_ = _19360_ ^ _19367_ /*11083*/;
assign _19374_ = D[11] ^ Q[14] /*11079*/;
assign _19371_ = _18875_ & _19374_ /*11075*/;
assign _19372_ = _18875_ ^ _19374_ /*11078*/;
assign _19373_ = _19365_ & _19372_ /*11076*/;
assign _19370_ = _19371_ | _19373_ /*11074*/;
assign _19261_ = _19365_ ^ _19372_ /*11077*/;
assign _19379_ = D[12] ^ Q[14] /*11073*/;
assign _19376_ = _18876_ & _19379_ /*11069*/;
assign _19377_ = _18876_ ^ _19379_ /*11072*/;
assign _19378_ = _19370_ & _19377_ /*11070*/;
assign _19375_ = _19376_ | _19378_ /*11068*/;
assign _19262_ = _19370_ ^ _19377_ /*11071*/;
assign _19384_ = D[13] ^ Q[14] /*11067*/;
assign _19381_ = _18877_ & _19384_ /*11063*/;
assign _19382_ = _18877_ ^ _19384_ /*11066*/;
assign _19383_ = _19375_ & _19382_ /*11064*/;
assign _19380_ = _19381_ | _19383_ /*11062*/;
assign _19263_ = _19375_ ^ _19382_ /*11065*/;
assign _19389_ = D[14] ^ Q[14] /*11061*/;
assign _19386_ = _18878_ & _19389_ /*11057*/;
assign _19387_ = _18878_ ^ _19389_ /*11060*/;
assign _19388_ = _19380_ & _19387_ /*11058*/;
assign _19385_ = _19386_ | _19388_ /*11056*/;
assign _19264_ = _19380_ ^ _19387_ /*11059*/;
assign _19394_ = D[15] ^ Q[14] /*11055*/;
assign _19391_ = _18879_ & _19394_ /*11051*/;
assign _19392_ = _18879_ ^ _19394_ /*11054*/;
assign _19393_ = _19385_ & _19392_ /*11052*/;
assign _19390_ = _19391_ | _19393_ /*11050*/;
assign _19265_ = _19385_ ^ _19392_ /*11053*/;
assign _19399_ = D[16] ^ Q[14] /*11049*/;
assign _19396_ = _18880_ & _19399_ /*11045*/;
assign _19397_ = _18880_ ^ _19399_ /*11048*/;
assign _19398_ = _19390_ & _19397_ /*11046*/;
assign _19395_ = _19396_ | _19398_ /*11044*/;
assign _19266_ = _19390_ ^ _19397_ /*11047*/;
assign _19404_ = D[17] ^ Q[14] /*11043*/;
assign _19401_ = _18881_ & _19404_ /*11039*/;
assign _19402_ = _18881_ ^ _19404_ /*11042*/;
assign _19403_ = _19395_ & _19402_ /*11040*/;
assign _19400_ = _19401_ | _19403_ /*11038*/;
assign _19267_ = _19395_ ^ _19402_ /*11041*/;
assign _19409_ = D[18] ^ Q[14] /*11037*/;
assign _19406_ = _18882_ & _19409_ /*11033*/;
assign _19407_ = _18882_ ^ _19409_ /*11036*/;
assign _19408_ = _19400_ & _19407_ /*11034*/;
assign _19405_ = _19406_ | _19408_ /*11032*/;
assign _19268_ = _19400_ ^ _19407_ /*11035*/;
assign _19414_ = D[19] ^ Q[14] /*11031*/;
assign _19411_ = _18883_ & _19414_ /*11027*/;
assign _19412_ = _18883_ ^ _19414_ /*11030*/;
assign _19413_ = _19405_ & _19412_ /*11028*/;
assign _19410_ = _19411_ | _19413_ /*11026*/;
assign _19269_ = _19405_ ^ _19412_ /*11029*/;
assign _19419_ = D[20] ^ Q[14] /*11025*/;
assign _19416_ = _18884_ & _19419_ /*11021*/;
assign _19417_ = _18884_ ^ _19419_ /*11024*/;
assign _19418_ = _19410_ & _19417_ /*11022*/;
assign _19415_ = _19416_ | _19418_ /*11020*/;
assign _19270_ = _19410_ ^ _19417_ /*11023*/;
assign _19424_ = D[21] ^ Q[14] /*11019*/;
assign _19421_ = _18885_ & _19424_ /*11015*/;
assign _19422_ = _18885_ ^ _19424_ /*11018*/;
assign _19423_ = _19415_ & _19422_ /*11016*/;
assign _19420_ = _19421_ | _19423_ /*11014*/;
assign _19271_ = _19415_ ^ _19422_ /*11017*/;
assign _19429_ = D[22] ^ Q[14] /*11013*/;
assign _19426_ = _18886_ & _19429_ /*11009*/;
assign _19427_ = _18886_ ^ _19429_ /*11012*/;
assign _19428_ = _19420_ & _19427_ /*11010*/;
assign _19425_ = _19426_ | _19428_ /*11008*/;
assign _19272_ = _19420_ ^ _19427_ /*11011*/;
assign _19434_ = D[23] ^ Q[14] /*11007*/;
assign _19431_ = _18887_ & _19434_ /*11003*/;
assign _19432_ = _18887_ ^ _19434_ /*11006*/;
assign _19433_ = _19425_ & _19432_ /*11004*/;
assign _19430_ = _19431_ | _19433_ /*11002*/;
assign _19273_ = _19425_ ^ _19432_ /*11005*/;
assign _19439_ = D[24] ^ Q[14] /*11001*/;
assign _19436_ = _18888_ & _19439_ /*10997*/;
assign _19437_ = _18888_ ^ _19439_ /*11000*/;
assign _19438_ = _19430_ & _19437_ /*10998*/;
assign _19435_ = _19436_ | _19438_ /*10996*/;
assign _19274_ = _19430_ ^ _19437_ /*10999*/;
assign _19444_ = D[25] ^ Q[14] /*10995*/;
assign _19441_ = _18889_ & _19444_ /*10991*/;
assign _19442_ = _18889_ ^ _19444_ /*10994*/;
assign _19443_ = _19435_ & _19442_ /*10992*/;
assign _19440_ = _19441_ | _19443_ /*10990*/;
assign _19275_ = _19435_ ^ _19442_ /*10993*/;
assign _19449_ = D[26] ^ Q[14] /*10989*/;
assign _19446_ = _18890_ & _19449_ /*10985*/;
assign _19447_ = _18890_ ^ _19449_ /*10988*/;
assign _19448_ = _19440_ & _19447_ /*10986*/;
assign _19445_ = _19446_ | _19448_ /*10984*/;
assign _19276_ = _19440_ ^ _19447_ /*10987*/;
assign _19454_ = D[27] ^ Q[14] /*10983*/;
assign _19451_ = _18891_ & _19454_ /*10979*/;
assign _19452_ = _18891_ ^ _19454_ /*10982*/;
assign _19453_ = _19445_ & _19452_ /*10980*/;
assign _19450_ = _19451_ | _19453_ /*10978*/;
assign _19277_ = _19445_ ^ _19452_ /*10981*/;
assign _19459_ = D[28] ^ Q[14] /*10977*/;
assign _19456_ = _18892_ & _19459_ /*10973*/;
assign _19457_ = _18892_ ^ _19459_ /*10976*/;
assign _19458_ = _19450_ & _19457_ /*10974*/;
assign _19455_ = _19456_ | _19458_ /*10972*/;
assign _19278_ = _19450_ ^ _19457_ /*10975*/;
assign _19464_ = D[29] ^ Q[14] /*10971*/;
assign _19461_ = _18893_ & _19464_ /*10967*/;
assign _19462_ = _18893_ ^ _19464_ /*10970*/;
assign _19463_ = _19455_ & _19462_ /*10968*/;
assign _19460_ = _19461_ | _19463_ /*10966*/;
assign _19279_ = _19455_ ^ _19462_ /*10969*/;
assign _19469_ = D[30] ^ Q[14] /*10965*/;
assign _19466_ = _18894_ & _19469_ /*10961*/;
assign _19467_ = _18894_ ^ _19469_ /*10964*/;
assign _19468_ = _19460_ & _19467_ /*10962*/;
assign _19465_ = _19466_ | _19468_ /*10960*/;
assign _19280_ = _19460_ ^ _19467_ /*10963*/;
assign _19474_ = D[31] ^ Q[14] /*10959*/;
assign _19471_ = _18895_ & _19474_ /*10955*/;
assign _19472_ = _18895_ ^ _19474_ /*10958*/;
assign _19473_ = _19465_ & _19472_ /*10956*/;
assign _19470_ = _19471_ | _19473_ /*10954*/;
assign _19281_ = _19465_ ^ _19472_ /*10957*/;
assign _19479_ = D[32] ^ Q[14] /*10953*/;
assign _19476_ = _18896_ & _19479_ /*10949*/;
assign _19477_ = _18896_ ^ _19479_ /*10952*/;
assign _19478_ = _19470_ & _19477_ /*10950*/;
assign _19475_ = _19476_ | _19478_ /*10948*/;
assign _19282_ = _19470_ ^ _19477_ /*10951*/;
assign _19484_ = D[33] ^ Q[14] /*10947*/;
assign _19481_ = _18897_ & _19484_ /*10943*/;
assign _19482_ = _18897_ ^ _19484_ /*10946*/;
assign _19483_ = _19475_ & _19482_ /*10944*/;
assign _19480_ = _19481_ | _19483_ /*10942*/;
assign _19283_ = _19475_ ^ _19482_ /*10945*/;
assign _19489_ = D[34] ^ Q[14] /*10941*/;
assign _19486_ = _18898_ & _19489_ /*10937*/;
assign _19487_ = _18898_ ^ _19489_ /*10940*/;
assign _19488_ = _19480_ & _19487_ /*10938*/;
assign _19485_ = _19486_ | _19488_ /*10936*/;
assign _19284_ = _19480_ ^ _19487_ /*10939*/;
assign _19494_ = D[35] ^ Q[14] /*10935*/;
assign _19491_ = _18899_ & _19494_ /*10931*/;
assign _19492_ = _18899_ ^ _19494_ /*10934*/;
assign _19493_ = _19485_ & _19492_ /*10932*/;
assign _19490_ = _19491_ | _19493_ /*10930*/;
assign _19285_ = _19485_ ^ _19492_ /*10933*/;
assign _19499_ = D[36] ^ Q[14] /*10929*/;
assign _19496_ = _18900_ & _19499_ /*10925*/;
assign _19497_ = _18900_ ^ _19499_ /*10928*/;
assign _19498_ = _19490_ & _19497_ /*10926*/;
assign _19495_ = _19496_ | _19498_ /*10924*/;
assign _19286_ = _19490_ ^ _19497_ /*10927*/;
assign _19504_ = D[37] ^ Q[14] /*10923*/;
assign _19501_ = _18901_ & _19504_ /*10919*/;
assign _19502_ = _18901_ ^ _19504_ /*10922*/;
assign _19503_ = _19495_ & _19502_ /*10920*/;
assign _19500_ = _19501_ | _19503_ /*10918*/;
assign _19287_ = _19495_ ^ _19502_ /*10921*/;
assign _19509_ = D[38] ^ Q[14] /*10917*/;
assign _19506_ = _18902_ & _19509_ /*10913*/;
assign _19507_ = _18902_ ^ _19509_ /*10916*/;
assign _19508_ = _19500_ & _19507_ /*10914*/;
assign _19505_ = _19506_ | _19508_ /*10912*/;
assign _19288_ = _19500_ ^ _19507_ /*10915*/;
assign _19514_ = D[39] ^ Q[14] /*10911*/;
assign _19511_ = _18903_ & _19514_ /*10907*/;
assign _19512_ = _18903_ ^ _19514_ /*10910*/;
assign _19513_ = _19505_ & _19512_ /*10908*/;
assign _19510_ = _19511_ | _19513_ /*10906*/;
assign _19289_ = _19505_ ^ _19512_ /*10909*/;
assign _19519_ = D[40] ^ Q[14] /*10905*/;
assign _19516_ = _18904_ & _19519_ /*10901*/;
assign _19517_ = _18904_ ^ _19519_ /*10904*/;
assign _19518_ = _19510_ & _19517_ /*10902*/;
assign _19515_ = _19516_ | _19518_ /*10900*/;
assign _19290_ = _19510_ ^ _19517_ /*10903*/;
assign _19524_ = D[41] ^ Q[14] /*10899*/;
assign _19521_ = _18905_ & _19524_ /*10895*/;
assign _19522_ = _18905_ ^ _19524_ /*10898*/;
assign _19523_ = _19515_ & _19522_ /*10896*/;
assign _19520_ = _19521_ | _19523_ /*10894*/;
assign _19291_ = _19515_ ^ _19522_ /*10897*/;
assign _19529_ = D[42] ^ Q[14] /*10893*/;
assign _19526_ = _18906_ & _19529_ /*10889*/;
assign _19527_ = _18906_ ^ _19529_ /*10892*/;
assign _19528_ = _19520_ & _19527_ /*10890*/;
assign _19525_ = _19526_ | _19528_ /*10888*/;
assign _19292_ = _19520_ ^ _19527_ /*10891*/;
assign _19534_ = D[43] ^ Q[14] /*10887*/;
assign _19531_ = _18907_ & _19534_ /*10883*/;
assign _19532_ = _18907_ ^ _19534_ /*10886*/;
assign _19533_ = _19525_ & _19532_ /*10884*/;
assign _19530_ = _19531_ | _19533_ /*10882*/;
assign _19293_ = _19525_ ^ _19532_ /*10885*/;
assign _19539_ = D[44] ^ Q[14] /*10881*/;
assign _19536_ = _18908_ & _19539_ /*10877*/;
assign _19537_ = _18908_ ^ _19539_ /*10880*/;
assign _19538_ = _19530_ & _19537_ /*10878*/;
assign _19535_ = _19536_ | _19538_ /*10876*/;
assign _19294_ = _19530_ ^ _19537_ /*10879*/;
assign _19544_ = D[45] ^ Q[14] /*10875*/;
assign _19541_ = _18909_ & _19544_ /*10871*/;
assign _19542_ = _18909_ ^ _19544_ /*10874*/;
assign _19543_ = _19535_ & _19542_ /*10872*/;
assign _19540_ = _19541_ | _19543_ /*10870*/;
assign _19295_ = _19535_ ^ _19542_ /*10873*/;
assign _19549_ = D[46] ^ Q[14] /*10869*/;
assign _19546_ = _18910_ & _19549_ /*10865*/;
assign _19547_ = _18910_ ^ _19549_ /*10868*/;
assign _19548_ = _19540_ & _19547_ /*10866*/;
assign _19545_ = _19546_ | _19548_ /*10864*/;
assign _19296_ = _19540_ ^ _19547_ /*10867*/;
assign _19554_ = D[47] ^ Q[14] /*10863*/;
assign _19551_ = _18911_ & _19554_ /*10859*/;
assign _19552_ = _18911_ ^ _19554_ /*10862*/;
assign _19553_ = _19545_ & _19552_ /*10860*/;
assign _19550_ = _19551_ | _19553_ /*10858*/;
assign _19297_ = _19545_ ^ _19552_ /*10861*/;
assign _19559_ = D[48] ^ Q[14] /*10857*/;
assign _19556_ = _18912_ & _19559_ /*10853*/;
assign _19557_ = _18912_ ^ _19559_ /*10856*/;
assign _19558_ = _19550_ & _19557_ /*10854*/;
assign _19555_ = _19556_ | _19558_ /*10852*/;
assign _19298_ = _19550_ ^ _19557_ /*10855*/;
assign _19564_ = D[49] ^ Q[14] /*10851*/;
assign _19561_ = _18913_ & _19564_ /*10847*/;
assign _19562_ = _18913_ ^ _19564_ /*10850*/;
assign _19563_ = _19555_ & _19562_ /*10848*/;
assign _19560_ = _19561_ | _19563_ /*10846*/;
assign _19299_ = _19555_ ^ _19562_ /*10849*/;
assign _19569_ = D[50] ^ Q[14] /*10845*/;
assign _19566_ = _18914_ & _19569_ /*10841*/;
assign _19567_ = _18914_ ^ _19569_ /*10844*/;
assign _19568_ = _19560_ & _19567_ /*10842*/;
assign _19565_ = _19566_ | _19568_ /*10840*/;
assign _19300_ = _19560_ ^ _19567_ /*10843*/;
assign _19574_ = D[51] ^ Q[14] /*10839*/;
assign _19571_ = _18915_ & _19574_ /*10835*/;
assign _19572_ = _18915_ ^ _19574_ /*10838*/;
assign _19573_ = _19565_ & _19572_ /*10836*/;
assign _19570_ = _19571_ | _19573_ /*10834*/;
assign _19301_ = _19565_ ^ _19572_ /*10837*/;
assign _19579_ = D[52] ^ Q[14] /*10833*/;
assign _19576_ = _18916_ & _19579_ /*10829*/;
assign _19577_ = _18916_ ^ _19579_ /*10832*/;
assign _19578_ = _19570_ & _19577_ /*10830*/;
assign _19575_ = _19576_ | _19578_ /*10828*/;
assign _19302_ = _19570_ ^ _19577_ /*10831*/;
assign _19584_ = D[53] ^ Q[14] /*10827*/;
assign _19581_ = _18917_ & _19584_ /*10823*/;
assign _19582_ = _18917_ ^ _19584_ /*10826*/;
assign _19583_ = _19575_ & _19582_ /*10824*/;
assign _19580_ = _19581_ | _19583_ /*10822*/;
assign _19303_ = _19575_ ^ _19582_ /*10825*/;
assign _19589_ = D[54] ^ Q[14] /*10821*/;
assign _19586_ = _18918_ & _19589_ /*10817*/;
assign _19587_ = _18918_ ^ _19589_ /*10820*/;
assign _19588_ = _19580_ & _19587_ /*10818*/;
assign _19585_ = _19586_ | _19588_ /*10816*/;
assign _19304_ = _19580_ ^ _19587_ /*10819*/;
assign _19594_ = D[55] ^ Q[14] /*10815*/;
assign _19591_ = _18919_ & _19594_ /*10811*/;
assign _19592_ = _18919_ ^ _19594_ /*10814*/;
assign _19593_ = _19585_ & _19592_ /*10812*/;
assign _19590_ = _19591_ | _19593_ /*10810*/;
assign _19305_ = _19585_ ^ _19592_ /*10813*/;
assign _19599_ = D[56] ^ Q[14] /*10809*/;
assign _19596_ = _18920_ & _19599_ /*10805*/;
assign _19597_ = _18920_ ^ _19599_ /*10808*/;
assign _19598_ = _19590_ & _19597_ /*10806*/;
assign _19595_ = _19596_ | _19598_ /*10804*/;
assign _19306_ = _19590_ ^ _19597_ /*10807*/;
assign _19604_ = D[57] ^ Q[14] /*10803*/;
assign _19601_ = _18921_ & _19604_ /*10799*/;
assign _19602_ = _18921_ ^ _19604_ /*10802*/;
assign _19603_ = _19595_ & _19602_ /*10800*/;
assign _19600_ = _19601_ | _19603_ /*10798*/;
assign _19307_ = _19595_ ^ _19602_ /*10801*/;
assign _19609_ = D[58] ^ Q[14] /*10797*/;
assign _19606_ = _18922_ & _19609_ /*10793*/;
assign _19607_ = _18922_ ^ _19609_ /*10796*/;
assign _19608_ = _19600_ & _19607_ /*10794*/;
assign _19605_ = _19606_ | _19608_ /*10792*/;
assign _19308_ = _19600_ ^ _19607_ /*10795*/;
assign _19614_ = D[59] ^ Q[14] /*10791*/;
assign _19611_ = _18923_ & _19614_ /*10787*/;
assign _19612_ = _18923_ ^ _19614_ /*10790*/;
assign _19613_ = _19605_ & _19612_ /*10788*/;
assign _19610_ = _19611_ | _19613_ /*10786*/;
assign _19309_ = _19605_ ^ _19612_ /*10789*/;
assign _19619_ = D[60] ^ Q[14] /*10785*/;
assign _19616_ = _18924_ & _19619_ /*10781*/;
assign _19617_ = _18924_ ^ _19619_ /*10784*/;
assign _19618_ = _19610_ & _19617_ /*10782*/;
assign _19615_ = _19616_ | _19618_ /*10780*/;
assign _19310_ = _19610_ ^ _19617_ /*10783*/;
assign _19624_ = D[61] ^ Q[14] /*10779*/;
assign _19621_ = _18925_ & _19624_ /*10775*/;
assign _19622_ = _18925_ ^ _19624_ /*10778*/;
assign _19623_ = _19615_ & _19622_ /*10776*/;
assign _19620_ = _19621_ | _19623_ /*10774*/;
assign _19311_ = _19615_ ^ _19622_ /*10777*/;
assign _19629_ = D[62] ^ Q[14] /*10773*/;
assign _19626_ = _18926_ & _19629_ /*10769*/;
assign _19627_ = _18926_ ^ _19629_ /*10772*/;
assign _19628_ = _19620_ & _19627_ /*10770*/;
assign _19625_ = _19626_ | _19628_ /*10768*/;
assign _19312_ = _19620_ ^ _19627_ /*10771*/;
assign _19633_ = zeroWire ^ Q[14] /*10767*/;
assign _19630_ = _18927_ & _19633_ /*10763*/;
assign _19631_ = _18927_ ^ _19633_ /*10766*/;
assign _19632_ = _19625_ & _19631_ /*10764*/;
assign Q[13] = _19630_ | _19632_ /*10762*/;
assign _19313_ = _19625_ ^ _19631_ /*10765*/;
assign _19704_ = D[0] ^ Q[13] /*10376*/;
assign _19701_ = R_0[12] & _19704_ /*10372*/;
assign _19702_ = R_0[12] ^ _19704_ /*10375*/;
assign _19703_ = Q[13] & _19702_ /*10373*/;
assign _19700_ = _19701_ | _19703_ /*10371*/;
assign _19635_ = Q[13] ^ _19702_ /*10374*/;
assign _19709_ = D[1] ^ Q[13] /*10370*/;
assign _19706_ = _19250_ & _19709_ /*10366*/;
assign _19707_ = _19250_ ^ _19709_ /*10369*/;
assign _19708_ = _19700_ & _19707_ /*10367*/;
assign _19705_ = _19706_ | _19708_ /*10365*/;
assign _19636_ = _19700_ ^ _19707_ /*10368*/;
assign _19714_ = D[2] ^ Q[13] /*10364*/;
assign _19711_ = _19251_ & _19714_ /*10360*/;
assign _19712_ = _19251_ ^ _19714_ /*10363*/;
assign _19713_ = _19705_ & _19712_ /*10361*/;
assign _19710_ = _19711_ | _19713_ /*10359*/;
assign _19637_ = _19705_ ^ _19712_ /*10362*/;
assign _19719_ = D[3] ^ Q[13] /*10358*/;
assign _19716_ = _19252_ & _19719_ /*10354*/;
assign _19717_ = _19252_ ^ _19719_ /*10357*/;
assign _19718_ = _19710_ & _19717_ /*10355*/;
assign _19715_ = _19716_ | _19718_ /*10353*/;
assign _19638_ = _19710_ ^ _19717_ /*10356*/;
assign _19724_ = D[4] ^ Q[13] /*10352*/;
assign _19721_ = _19253_ & _19724_ /*10348*/;
assign _19722_ = _19253_ ^ _19724_ /*10351*/;
assign _19723_ = _19715_ & _19722_ /*10349*/;
assign _19720_ = _19721_ | _19723_ /*10347*/;
assign _19639_ = _19715_ ^ _19722_ /*10350*/;
assign _19729_ = D[5] ^ Q[13] /*10346*/;
assign _19726_ = _19254_ & _19729_ /*10342*/;
assign _19727_ = _19254_ ^ _19729_ /*10345*/;
assign _19728_ = _19720_ & _19727_ /*10343*/;
assign _19725_ = _19726_ | _19728_ /*10341*/;
assign _19640_ = _19720_ ^ _19727_ /*10344*/;
assign _19734_ = D[6] ^ Q[13] /*10340*/;
assign _19731_ = _19255_ & _19734_ /*10336*/;
assign _19732_ = _19255_ ^ _19734_ /*10339*/;
assign _19733_ = _19725_ & _19732_ /*10337*/;
assign _19730_ = _19731_ | _19733_ /*10335*/;
assign _19641_ = _19725_ ^ _19732_ /*10338*/;
assign _19739_ = D[7] ^ Q[13] /*10334*/;
assign _19736_ = _19256_ & _19739_ /*10330*/;
assign _19737_ = _19256_ ^ _19739_ /*10333*/;
assign _19738_ = _19730_ & _19737_ /*10331*/;
assign _19735_ = _19736_ | _19738_ /*10329*/;
assign _19642_ = _19730_ ^ _19737_ /*10332*/;
assign _19744_ = D[8] ^ Q[13] /*10328*/;
assign _19741_ = _19257_ & _19744_ /*10324*/;
assign _19742_ = _19257_ ^ _19744_ /*10327*/;
assign _19743_ = _19735_ & _19742_ /*10325*/;
assign _19740_ = _19741_ | _19743_ /*10323*/;
assign _19643_ = _19735_ ^ _19742_ /*10326*/;
assign _19749_ = D[9] ^ Q[13] /*10322*/;
assign _19746_ = _19258_ & _19749_ /*10318*/;
assign _19747_ = _19258_ ^ _19749_ /*10321*/;
assign _19748_ = _19740_ & _19747_ /*10319*/;
assign _19745_ = _19746_ | _19748_ /*10317*/;
assign _19644_ = _19740_ ^ _19747_ /*10320*/;
assign _19754_ = D[10] ^ Q[13] /*10316*/;
assign _19751_ = _19259_ & _19754_ /*10312*/;
assign _19752_ = _19259_ ^ _19754_ /*10315*/;
assign _19753_ = _19745_ & _19752_ /*10313*/;
assign _19750_ = _19751_ | _19753_ /*10311*/;
assign _19645_ = _19745_ ^ _19752_ /*10314*/;
assign _19759_ = D[11] ^ Q[13] /*10310*/;
assign _19756_ = _19260_ & _19759_ /*10306*/;
assign _19757_ = _19260_ ^ _19759_ /*10309*/;
assign _19758_ = _19750_ & _19757_ /*10307*/;
assign _19755_ = _19756_ | _19758_ /*10305*/;
assign _19646_ = _19750_ ^ _19757_ /*10308*/;
assign _19764_ = D[12] ^ Q[13] /*10304*/;
assign _19761_ = _19261_ & _19764_ /*10300*/;
assign _19762_ = _19261_ ^ _19764_ /*10303*/;
assign _19763_ = _19755_ & _19762_ /*10301*/;
assign _19760_ = _19761_ | _19763_ /*10299*/;
assign _19647_ = _19755_ ^ _19762_ /*10302*/;
assign _19769_ = D[13] ^ Q[13] /*10298*/;
assign _19766_ = _19262_ & _19769_ /*10294*/;
assign _19767_ = _19262_ ^ _19769_ /*10297*/;
assign _19768_ = _19760_ & _19767_ /*10295*/;
assign _19765_ = _19766_ | _19768_ /*10293*/;
assign _19648_ = _19760_ ^ _19767_ /*10296*/;
assign _19774_ = D[14] ^ Q[13] /*10292*/;
assign _19771_ = _19263_ & _19774_ /*10288*/;
assign _19772_ = _19263_ ^ _19774_ /*10291*/;
assign _19773_ = _19765_ & _19772_ /*10289*/;
assign _19770_ = _19771_ | _19773_ /*10287*/;
assign _19649_ = _19765_ ^ _19772_ /*10290*/;
assign _19779_ = D[15] ^ Q[13] /*10286*/;
assign _19776_ = _19264_ & _19779_ /*10282*/;
assign _19777_ = _19264_ ^ _19779_ /*10285*/;
assign _19778_ = _19770_ & _19777_ /*10283*/;
assign _19775_ = _19776_ | _19778_ /*10281*/;
assign _19650_ = _19770_ ^ _19777_ /*10284*/;
assign _19784_ = D[16] ^ Q[13] /*10280*/;
assign _19781_ = _19265_ & _19784_ /*10276*/;
assign _19782_ = _19265_ ^ _19784_ /*10279*/;
assign _19783_ = _19775_ & _19782_ /*10277*/;
assign _19780_ = _19781_ | _19783_ /*10275*/;
assign _19651_ = _19775_ ^ _19782_ /*10278*/;
assign _19789_ = D[17] ^ Q[13] /*10274*/;
assign _19786_ = _19266_ & _19789_ /*10270*/;
assign _19787_ = _19266_ ^ _19789_ /*10273*/;
assign _19788_ = _19780_ & _19787_ /*10271*/;
assign _19785_ = _19786_ | _19788_ /*10269*/;
assign _19652_ = _19780_ ^ _19787_ /*10272*/;
assign _19794_ = D[18] ^ Q[13] /*10268*/;
assign _19791_ = _19267_ & _19794_ /*10264*/;
assign _19792_ = _19267_ ^ _19794_ /*10267*/;
assign _19793_ = _19785_ & _19792_ /*10265*/;
assign _19790_ = _19791_ | _19793_ /*10263*/;
assign _19653_ = _19785_ ^ _19792_ /*10266*/;
assign _19799_ = D[19] ^ Q[13] /*10262*/;
assign _19796_ = _19268_ & _19799_ /*10258*/;
assign _19797_ = _19268_ ^ _19799_ /*10261*/;
assign _19798_ = _19790_ & _19797_ /*10259*/;
assign _19795_ = _19796_ | _19798_ /*10257*/;
assign _19654_ = _19790_ ^ _19797_ /*10260*/;
assign _19804_ = D[20] ^ Q[13] /*10256*/;
assign _19801_ = _19269_ & _19804_ /*10252*/;
assign _19802_ = _19269_ ^ _19804_ /*10255*/;
assign _19803_ = _19795_ & _19802_ /*10253*/;
assign _19800_ = _19801_ | _19803_ /*10251*/;
assign _19655_ = _19795_ ^ _19802_ /*10254*/;
assign _19809_ = D[21] ^ Q[13] /*10250*/;
assign _19806_ = _19270_ & _19809_ /*10246*/;
assign _19807_ = _19270_ ^ _19809_ /*10249*/;
assign _19808_ = _19800_ & _19807_ /*10247*/;
assign _19805_ = _19806_ | _19808_ /*10245*/;
assign _19656_ = _19800_ ^ _19807_ /*10248*/;
assign _19814_ = D[22] ^ Q[13] /*10244*/;
assign _19811_ = _19271_ & _19814_ /*10240*/;
assign _19812_ = _19271_ ^ _19814_ /*10243*/;
assign _19813_ = _19805_ & _19812_ /*10241*/;
assign _19810_ = _19811_ | _19813_ /*10239*/;
assign _19657_ = _19805_ ^ _19812_ /*10242*/;
assign _19819_ = D[23] ^ Q[13] /*10238*/;
assign _19816_ = _19272_ & _19819_ /*10234*/;
assign _19817_ = _19272_ ^ _19819_ /*10237*/;
assign _19818_ = _19810_ & _19817_ /*10235*/;
assign _19815_ = _19816_ | _19818_ /*10233*/;
assign _19658_ = _19810_ ^ _19817_ /*10236*/;
assign _19824_ = D[24] ^ Q[13] /*10232*/;
assign _19821_ = _19273_ & _19824_ /*10228*/;
assign _19822_ = _19273_ ^ _19824_ /*10231*/;
assign _19823_ = _19815_ & _19822_ /*10229*/;
assign _19820_ = _19821_ | _19823_ /*10227*/;
assign _19659_ = _19815_ ^ _19822_ /*10230*/;
assign _19829_ = D[25] ^ Q[13] /*10226*/;
assign _19826_ = _19274_ & _19829_ /*10222*/;
assign _19827_ = _19274_ ^ _19829_ /*10225*/;
assign _19828_ = _19820_ & _19827_ /*10223*/;
assign _19825_ = _19826_ | _19828_ /*10221*/;
assign _19660_ = _19820_ ^ _19827_ /*10224*/;
assign _19834_ = D[26] ^ Q[13] /*10220*/;
assign _19831_ = _19275_ & _19834_ /*10216*/;
assign _19832_ = _19275_ ^ _19834_ /*10219*/;
assign _19833_ = _19825_ & _19832_ /*10217*/;
assign _19830_ = _19831_ | _19833_ /*10215*/;
assign _19661_ = _19825_ ^ _19832_ /*10218*/;
assign _19839_ = D[27] ^ Q[13] /*10214*/;
assign _19836_ = _19276_ & _19839_ /*10210*/;
assign _19837_ = _19276_ ^ _19839_ /*10213*/;
assign _19838_ = _19830_ & _19837_ /*10211*/;
assign _19835_ = _19836_ | _19838_ /*10209*/;
assign _19662_ = _19830_ ^ _19837_ /*10212*/;
assign _19844_ = D[28] ^ Q[13] /*10208*/;
assign _19841_ = _19277_ & _19844_ /*10204*/;
assign _19842_ = _19277_ ^ _19844_ /*10207*/;
assign _19843_ = _19835_ & _19842_ /*10205*/;
assign _19840_ = _19841_ | _19843_ /*10203*/;
assign _19663_ = _19835_ ^ _19842_ /*10206*/;
assign _19849_ = D[29] ^ Q[13] /*10202*/;
assign _19846_ = _19278_ & _19849_ /*10198*/;
assign _19847_ = _19278_ ^ _19849_ /*10201*/;
assign _19848_ = _19840_ & _19847_ /*10199*/;
assign _19845_ = _19846_ | _19848_ /*10197*/;
assign _19664_ = _19840_ ^ _19847_ /*10200*/;
assign _19854_ = D[30] ^ Q[13] /*10196*/;
assign _19851_ = _19279_ & _19854_ /*10192*/;
assign _19852_ = _19279_ ^ _19854_ /*10195*/;
assign _19853_ = _19845_ & _19852_ /*10193*/;
assign _19850_ = _19851_ | _19853_ /*10191*/;
assign _19665_ = _19845_ ^ _19852_ /*10194*/;
assign _19859_ = D[31] ^ Q[13] /*10190*/;
assign _19856_ = _19280_ & _19859_ /*10186*/;
assign _19857_ = _19280_ ^ _19859_ /*10189*/;
assign _19858_ = _19850_ & _19857_ /*10187*/;
assign _19855_ = _19856_ | _19858_ /*10185*/;
assign _19666_ = _19850_ ^ _19857_ /*10188*/;
assign _19864_ = D[32] ^ Q[13] /*10184*/;
assign _19861_ = _19281_ & _19864_ /*10180*/;
assign _19862_ = _19281_ ^ _19864_ /*10183*/;
assign _19863_ = _19855_ & _19862_ /*10181*/;
assign _19860_ = _19861_ | _19863_ /*10179*/;
assign _19667_ = _19855_ ^ _19862_ /*10182*/;
assign _19869_ = D[33] ^ Q[13] /*10178*/;
assign _19866_ = _19282_ & _19869_ /*10174*/;
assign _19867_ = _19282_ ^ _19869_ /*10177*/;
assign _19868_ = _19860_ & _19867_ /*10175*/;
assign _19865_ = _19866_ | _19868_ /*10173*/;
assign _19668_ = _19860_ ^ _19867_ /*10176*/;
assign _19874_ = D[34] ^ Q[13] /*10172*/;
assign _19871_ = _19283_ & _19874_ /*10168*/;
assign _19872_ = _19283_ ^ _19874_ /*10171*/;
assign _19873_ = _19865_ & _19872_ /*10169*/;
assign _19870_ = _19871_ | _19873_ /*10167*/;
assign _19669_ = _19865_ ^ _19872_ /*10170*/;
assign _19879_ = D[35] ^ Q[13] /*10166*/;
assign _19876_ = _19284_ & _19879_ /*10162*/;
assign _19877_ = _19284_ ^ _19879_ /*10165*/;
assign _19878_ = _19870_ & _19877_ /*10163*/;
assign _19875_ = _19876_ | _19878_ /*10161*/;
assign _19670_ = _19870_ ^ _19877_ /*10164*/;
assign _19884_ = D[36] ^ Q[13] /*10160*/;
assign _19881_ = _19285_ & _19884_ /*10156*/;
assign _19882_ = _19285_ ^ _19884_ /*10159*/;
assign _19883_ = _19875_ & _19882_ /*10157*/;
assign _19880_ = _19881_ | _19883_ /*10155*/;
assign _19671_ = _19875_ ^ _19882_ /*10158*/;
assign _19889_ = D[37] ^ Q[13] /*10154*/;
assign _19886_ = _19286_ & _19889_ /*10150*/;
assign _19887_ = _19286_ ^ _19889_ /*10153*/;
assign _19888_ = _19880_ & _19887_ /*10151*/;
assign _19885_ = _19886_ | _19888_ /*10149*/;
assign _19672_ = _19880_ ^ _19887_ /*10152*/;
assign _19894_ = D[38] ^ Q[13] /*10148*/;
assign _19891_ = _19287_ & _19894_ /*10144*/;
assign _19892_ = _19287_ ^ _19894_ /*10147*/;
assign _19893_ = _19885_ & _19892_ /*10145*/;
assign _19890_ = _19891_ | _19893_ /*10143*/;
assign _19673_ = _19885_ ^ _19892_ /*10146*/;
assign _19899_ = D[39] ^ Q[13] /*10142*/;
assign _19896_ = _19288_ & _19899_ /*10138*/;
assign _19897_ = _19288_ ^ _19899_ /*10141*/;
assign _19898_ = _19890_ & _19897_ /*10139*/;
assign _19895_ = _19896_ | _19898_ /*10137*/;
assign _19674_ = _19890_ ^ _19897_ /*10140*/;
assign _19904_ = D[40] ^ Q[13] /*10136*/;
assign _19901_ = _19289_ & _19904_ /*10132*/;
assign _19902_ = _19289_ ^ _19904_ /*10135*/;
assign _19903_ = _19895_ & _19902_ /*10133*/;
assign _19900_ = _19901_ | _19903_ /*10131*/;
assign _19675_ = _19895_ ^ _19902_ /*10134*/;
assign _19909_ = D[41] ^ Q[13] /*10130*/;
assign _19906_ = _19290_ & _19909_ /*10126*/;
assign _19907_ = _19290_ ^ _19909_ /*10129*/;
assign _19908_ = _19900_ & _19907_ /*10127*/;
assign _19905_ = _19906_ | _19908_ /*10125*/;
assign _19676_ = _19900_ ^ _19907_ /*10128*/;
assign _19914_ = D[42] ^ Q[13] /*10124*/;
assign _19911_ = _19291_ & _19914_ /*10120*/;
assign _19912_ = _19291_ ^ _19914_ /*10123*/;
assign _19913_ = _19905_ & _19912_ /*10121*/;
assign _19910_ = _19911_ | _19913_ /*10119*/;
assign _19677_ = _19905_ ^ _19912_ /*10122*/;
assign _19919_ = D[43] ^ Q[13] /*10118*/;
assign _19916_ = _19292_ & _19919_ /*10114*/;
assign _19917_ = _19292_ ^ _19919_ /*10117*/;
assign _19918_ = _19910_ & _19917_ /*10115*/;
assign _19915_ = _19916_ | _19918_ /*10113*/;
assign _19678_ = _19910_ ^ _19917_ /*10116*/;
assign _19924_ = D[44] ^ Q[13] /*10112*/;
assign _19921_ = _19293_ & _19924_ /*10108*/;
assign _19922_ = _19293_ ^ _19924_ /*10111*/;
assign _19923_ = _19915_ & _19922_ /*10109*/;
assign _19920_ = _19921_ | _19923_ /*10107*/;
assign _19679_ = _19915_ ^ _19922_ /*10110*/;
assign _19929_ = D[45] ^ Q[13] /*10106*/;
assign _19926_ = _19294_ & _19929_ /*10102*/;
assign _19927_ = _19294_ ^ _19929_ /*10105*/;
assign _19928_ = _19920_ & _19927_ /*10103*/;
assign _19925_ = _19926_ | _19928_ /*10101*/;
assign _19680_ = _19920_ ^ _19927_ /*10104*/;
assign _19934_ = D[46] ^ Q[13] /*10100*/;
assign _19931_ = _19295_ & _19934_ /*10096*/;
assign _19932_ = _19295_ ^ _19934_ /*10099*/;
assign _19933_ = _19925_ & _19932_ /*10097*/;
assign _19930_ = _19931_ | _19933_ /*10095*/;
assign _19681_ = _19925_ ^ _19932_ /*10098*/;
assign _19939_ = D[47] ^ Q[13] /*10094*/;
assign _19936_ = _19296_ & _19939_ /*10090*/;
assign _19937_ = _19296_ ^ _19939_ /*10093*/;
assign _19938_ = _19930_ & _19937_ /*10091*/;
assign _19935_ = _19936_ | _19938_ /*10089*/;
assign _19682_ = _19930_ ^ _19937_ /*10092*/;
assign _19944_ = D[48] ^ Q[13] /*10088*/;
assign _19941_ = _19297_ & _19944_ /*10084*/;
assign _19942_ = _19297_ ^ _19944_ /*10087*/;
assign _19943_ = _19935_ & _19942_ /*10085*/;
assign _19940_ = _19941_ | _19943_ /*10083*/;
assign _19683_ = _19935_ ^ _19942_ /*10086*/;
assign _19949_ = D[49] ^ Q[13] /*10082*/;
assign _19946_ = _19298_ & _19949_ /*10078*/;
assign _19947_ = _19298_ ^ _19949_ /*10081*/;
assign _19948_ = _19940_ & _19947_ /*10079*/;
assign _19945_ = _19946_ | _19948_ /*10077*/;
assign _19684_ = _19940_ ^ _19947_ /*10080*/;
assign _19954_ = D[50] ^ Q[13] /*10076*/;
assign _19951_ = _19299_ & _19954_ /*10072*/;
assign _19952_ = _19299_ ^ _19954_ /*10075*/;
assign _19953_ = _19945_ & _19952_ /*10073*/;
assign _19950_ = _19951_ | _19953_ /*10071*/;
assign _19685_ = _19945_ ^ _19952_ /*10074*/;
assign _19959_ = D[51] ^ Q[13] /*10070*/;
assign _19956_ = _19300_ & _19959_ /*10066*/;
assign _19957_ = _19300_ ^ _19959_ /*10069*/;
assign _19958_ = _19950_ & _19957_ /*10067*/;
assign _19955_ = _19956_ | _19958_ /*10065*/;
assign _19686_ = _19950_ ^ _19957_ /*10068*/;
assign _19964_ = D[52] ^ Q[13] /*10064*/;
assign _19961_ = _19301_ & _19964_ /*10060*/;
assign _19962_ = _19301_ ^ _19964_ /*10063*/;
assign _19963_ = _19955_ & _19962_ /*10061*/;
assign _19960_ = _19961_ | _19963_ /*10059*/;
assign _19687_ = _19955_ ^ _19962_ /*10062*/;
assign _19969_ = D[53] ^ Q[13] /*10058*/;
assign _19966_ = _19302_ & _19969_ /*10054*/;
assign _19967_ = _19302_ ^ _19969_ /*10057*/;
assign _19968_ = _19960_ & _19967_ /*10055*/;
assign _19965_ = _19966_ | _19968_ /*10053*/;
assign _19688_ = _19960_ ^ _19967_ /*10056*/;
assign _19974_ = D[54] ^ Q[13] /*10052*/;
assign _19971_ = _19303_ & _19974_ /*10048*/;
assign _19972_ = _19303_ ^ _19974_ /*10051*/;
assign _19973_ = _19965_ & _19972_ /*10049*/;
assign _19970_ = _19971_ | _19973_ /*10047*/;
assign _19689_ = _19965_ ^ _19972_ /*10050*/;
assign _19979_ = D[55] ^ Q[13] /*10046*/;
assign _19976_ = _19304_ & _19979_ /*10042*/;
assign _19977_ = _19304_ ^ _19979_ /*10045*/;
assign _19978_ = _19970_ & _19977_ /*10043*/;
assign _19975_ = _19976_ | _19978_ /*10041*/;
assign _19690_ = _19970_ ^ _19977_ /*10044*/;
assign _19984_ = D[56] ^ Q[13] /*10040*/;
assign _19981_ = _19305_ & _19984_ /*10036*/;
assign _19982_ = _19305_ ^ _19984_ /*10039*/;
assign _19983_ = _19975_ & _19982_ /*10037*/;
assign _19980_ = _19981_ | _19983_ /*10035*/;
assign _19691_ = _19975_ ^ _19982_ /*10038*/;
assign _19989_ = D[57] ^ Q[13] /*10034*/;
assign _19986_ = _19306_ & _19989_ /*10030*/;
assign _19987_ = _19306_ ^ _19989_ /*10033*/;
assign _19988_ = _19980_ & _19987_ /*10031*/;
assign _19985_ = _19986_ | _19988_ /*10029*/;
assign _19692_ = _19980_ ^ _19987_ /*10032*/;
assign _19994_ = D[58] ^ Q[13] /*10028*/;
assign _19991_ = _19307_ & _19994_ /*10024*/;
assign _19992_ = _19307_ ^ _19994_ /*10027*/;
assign _19993_ = _19985_ & _19992_ /*10025*/;
assign _19990_ = _19991_ | _19993_ /*10023*/;
assign _19693_ = _19985_ ^ _19992_ /*10026*/;
assign _19999_ = D[59] ^ Q[13] /*10022*/;
assign _19996_ = _19308_ & _19999_ /*10018*/;
assign _19997_ = _19308_ ^ _19999_ /*10021*/;
assign _19998_ = _19990_ & _19997_ /*10019*/;
assign _19995_ = _19996_ | _19998_ /*10017*/;
assign _19694_ = _19990_ ^ _19997_ /*10020*/;
assign _20004_ = D[60] ^ Q[13] /*10016*/;
assign _20001_ = _19309_ & _20004_ /*10012*/;
assign _20002_ = _19309_ ^ _20004_ /*10015*/;
assign _20003_ = _19995_ & _20002_ /*10013*/;
assign _20000_ = _20001_ | _20003_ /*10011*/;
assign _19695_ = _19995_ ^ _20002_ /*10014*/;
assign _20009_ = D[61] ^ Q[13] /*10010*/;
assign _20006_ = _19310_ & _20009_ /*10006*/;
assign _20007_ = _19310_ ^ _20009_ /*10009*/;
assign _20008_ = _20000_ & _20007_ /*10007*/;
assign _20005_ = _20006_ | _20008_ /*10005*/;
assign _19696_ = _20000_ ^ _20007_ /*10008*/;
assign _20014_ = D[62] ^ Q[13] /*10004*/;
assign _20011_ = _19311_ & _20014_ /*10000*/;
assign _20012_ = _19311_ ^ _20014_ /*10003*/;
assign _20013_ = _20005_ & _20012_ /*10001*/;
assign _20010_ = _20011_ | _20013_ /*9999*/;
assign _19697_ = _20005_ ^ _20012_ /*10002*/;
assign _20018_ = zeroWire ^ Q[13] /*9998*/;
assign _20015_ = _19312_ & _20018_ /*9994*/;
assign _20016_ = _19312_ ^ _20018_ /*9997*/;
assign _20017_ = _20010_ & _20016_ /*9995*/;
assign Q[12] = _20015_ | _20017_ /*9993*/;
assign _19698_ = _20010_ ^ _20016_ /*9996*/;
assign _20089_ = D[0] ^ Q[12] /*9607*/;
assign _20086_ = R_0[11] & _20089_ /*9603*/;
assign _20087_ = R_0[11] ^ _20089_ /*9606*/;
assign _20088_ = Q[12] & _20087_ /*9604*/;
assign _20085_ = _20086_ | _20088_ /*9602*/;
assign _20020_ = Q[12] ^ _20087_ /*9605*/;
assign _20094_ = D[1] ^ Q[12] /*9601*/;
assign _20091_ = _19635_ & _20094_ /*9597*/;
assign _20092_ = _19635_ ^ _20094_ /*9600*/;
assign _20093_ = _20085_ & _20092_ /*9598*/;
assign _20090_ = _20091_ | _20093_ /*9596*/;
assign _20021_ = _20085_ ^ _20092_ /*9599*/;
assign _20099_ = D[2] ^ Q[12] /*9595*/;
assign _20096_ = _19636_ & _20099_ /*9591*/;
assign _20097_ = _19636_ ^ _20099_ /*9594*/;
assign _20098_ = _20090_ & _20097_ /*9592*/;
assign _20095_ = _20096_ | _20098_ /*9590*/;
assign _20022_ = _20090_ ^ _20097_ /*9593*/;
assign _20104_ = D[3] ^ Q[12] /*9589*/;
assign _20101_ = _19637_ & _20104_ /*9585*/;
assign _20102_ = _19637_ ^ _20104_ /*9588*/;
assign _20103_ = _20095_ & _20102_ /*9586*/;
assign _20100_ = _20101_ | _20103_ /*9584*/;
assign _20023_ = _20095_ ^ _20102_ /*9587*/;
assign _20109_ = D[4] ^ Q[12] /*9583*/;
assign _20106_ = _19638_ & _20109_ /*9579*/;
assign _20107_ = _19638_ ^ _20109_ /*9582*/;
assign _20108_ = _20100_ & _20107_ /*9580*/;
assign _20105_ = _20106_ | _20108_ /*9578*/;
assign _20024_ = _20100_ ^ _20107_ /*9581*/;
assign _20114_ = D[5] ^ Q[12] /*9577*/;
assign _20111_ = _19639_ & _20114_ /*9573*/;
assign _20112_ = _19639_ ^ _20114_ /*9576*/;
assign _20113_ = _20105_ & _20112_ /*9574*/;
assign _20110_ = _20111_ | _20113_ /*9572*/;
assign _20025_ = _20105_ ^ _20112_ /*9575*/;
assign _20119_ = D[6] ^ Q[12] /*9571*/;
assign _20116_ = _19640_ & _20119_ /*9567*/;
assign _20117_ = _19640_ ^ _20119_ /*9570*/;
assign _20118_ = _20110_ & _20117_ /*9568*/;
assign _20115_ = _20116_ | _20118_ /*9566*/;
assign _20026_ = _20110_ ^ _20117_ /*9569*/;
assign _20124_ = D[7] ^ Q[12] /*9565*/;
assign _20121_ = _19641_ & _20124_ /*9561*/;
assign _20122_ = _19641_ ^ _20124_ /*9564*/;
assign _20123_ = _20115_ & _20122_ /*9562*/;
assign _20120_ = _20121_ | _20123_ /*9560*/;
assign _20027_ = _20115_ ^ _20122_ /*9563*/;
assign _20129_ = D[8] ^ Q[12] /*9559*/;
assign _20126_ = _19642_ & _20129_ /*9555*/;
assign _20127_ = _19642_ ^ _20129_ /*9558*/;
assign _20128_ = _20120_ & _20127_ /*9556*/;
assign _20125_ = _20126_ | _20128_ /*9554*/;
assign _20028_ = _20120_ ^ _20127_ /*9557*/;
assign _20134_ = D[9] ^ Q[12] /*9553*/;
assign _20131_ = _19643_ & _20134_ /*9549*/;
assign _20132_ = _19643_ ^ _20134_ /*9552*/;
assign _20133_ = _20125_ & _20132_ /*9550*/;
assign _20130_ = _20131_ | _20133_ /*9548*/;
assign _20029_ = _20125_ ^ _20132_ /*9551*/;
assign _20139_ = D[10] ^ Q[12] /*9547*/;
assign _20136_ = _19644_ & _20139_ /*9543*/;
assign _20137_ = _19644_ ^ _20139_ /*9546*/;
assign _20138_ = _20130_ & _20137_ /*9544*/;
assign _20135_ = _20136_ | _20138_ /*9542*/;
assign _20030_ = _20130_ ^ _20137_ /*9545*/;
assign _20144_ = D[11] ^ Q[12] /*9541*/;
assign _20141_ = _19645_ & _20144_ /*9537*/;
assign _20142_ = _19645_ ^ _20144_ /*9540*/;
assign _20143_ = _20135_ & _20142_ /*9538*/;
assign _20140_ = _20141_ | _20143_ /*9536*/;
assign _20031_ = _20135_ ^ _20142_ /*9539*/;
assign _20149_ = D[12] ^ Q[12] /*9535*/;
assign _20146_ = _19646_ & _20149_ /*9531*/;
assign _20147_ = _19646_ ^ _20149_ /*9534*/;
assign _20148_ = _20140_ & _20147_ /*9532*/;
assign _20145_ = _20146_ | _20148_ /*9530*/;
assign _20032_ = _20140_ ^ _20147_ /*9533*/;
assign _20154_ = D[13] ^ Q[12] /*9529*/;
assign _20151_ = _19647_ & _20154_ /*9525*/;
assign _20152_ = _19647_ ^ _20154_ /*9528*/;
assign _20153_ = _20145_ & _20152_ /*9526*/;
assign _20150_ = _20151_ | _20153_ /*9524*/;
assign _20033_ = _20145_ ^ _20152_ /*9527*/;
assign _20159_ = D[14] ^ Q[12] /*9523*/;
assign _20156_ = _19648_ & _20159_ /*9519*/;
assign _20157_ = _19648_ ^ _20159_ /*9522*/;
assign _20158_ = _20150_ & _20157_ /*9520*/;
assign _20155_ = _20156_ | _20158_ /*9518*/;
assign _20034_ = _20150_ ^ _20157_ /*9521*/;
assign _20164_ = D[15] ^ Q[12] /*9517*/;
assign _20161_ = _19649_ & _20164_ /*9513*/;
assign _20162_ = _19649_ ^ _20164_ /*9516*/;
assign _20163_ = _20155_ & _20162_ /*9514*/;
assign _20160_ = _20161_ | _20163_ /*9512*/;
assign _20035_ = _20155_ ^ _20162_ /*9515*/;
assign _20169_ = D[16] ^ Q[12] /*9511*/;
assign _20166_ = _19650_ & _20169_ /*9507*/;
assign _20167_ = _19650_ ^ _20169_ /*9510*/;
assign _20168_ = _20160_ & _20167_ /*9508*/;
assign _20165_ = _20166_ | _20168_ /*9506*/;
assign _20036_ = _20160_ ^ _20167_ /*9509*/;
assign _20174_ = D[17] ^ Q[12] /*9505*/;
assign _20171_ = _19651_ & _20174_ /*9501*/;
assign _20172_ = _19651_ ^ _20174_ /*9504*/;
assign _20173_ = _20165_ & _20172_ /*9502*/;
assign _20170_ = _20171_ | _20173_ /*9500*/;
assign _20037_ = _20165_ ^ _20172_ /*9503*/;
assign _20179_ = D[18] ^ Q[12] /*9499*/;
assign _20176_ = _19652_ & _20179_ /*9495*/;
assign _20177_ = _19652_ ^ _20179_ /*9498*/;
assign _20178_ = _20170_ & _20177_ /*9496*/;
assign _20175_ = _20176_ | _20178_ /*9494*/;
assign _20038_ = _20170_ ^ _20177_ /*9497*/;
assign _20184_ = D[19] ^ Q[12] /*9493*/;
assign _20181_ = _19653_ & _20184_ /*9489*/;
assign _20182_ = _19653_ ^ _20184_ /*9492*/;
assign _20183_ = _20175_ & _20182_ /*9490*/;
assign _20180_ = _20181_ | _20183_ /*9488*/;
assign _20039_ = _20175_ ^ _20182_ /*9491*/;
assign _20189_ = D[20] ^ Q[12] /*9487*/;
assign _20186_ = _19654_ & _20189_ /*9483*/;
assign _20187_ = _19654_ ^ _20189_ /*9486*/;
assign _20188_ = _20180_ & _20187_ /*9484*/;
assign _20185_ = _20186_ | _20188_ /*9482*/;
assign _20040_ = _20180_ ^ _20187_ /*9485*/;
assign _20194_ = D[21] ^ Q[12] /*9481*/;
assign _20191_ = _19655_ & _20194_ /*9477*/;
assign _20192_ = _19655_ ^ _20194_ /*9480*/;
assign _20193_ = _20185_ & _20192_ /*9478*/;
assign _20190_ = _20191_ | _20193_ /*9476*/;
assign _20041_ = _20185_ ^ _20192_ /*9479*/;
assign _20199_ = D[22] ^ Q[12] /*9475*/;
assign _20196_ = _19656_ & _20199_ /*9471*/;
assign _20197_ = _19656_ ^ _20199_ /*9474*/;
assign _20198_ = _20190_ & _20197_ /*9472*/;
assign _20195_ = _20196_ | _20198_ /*9470*/;
assign _20042_ = _20190_ ^ _20197_ /*9473*/;
assign _20204_ = D[23] ^ Q[12] /*9469*/;
assign _20201_ = _19657_ & _20204_ /*9465*/;
assign _20202_ = _19657_ ^ _20204_ /*9468*/;
assign _20203_ = _20195_ & _20202_ /*9466*/;
assign _20200_ = _20201_ | _20203_ /*9464*/;
assign _20043_ = _20195_ ^ _20202_ /*9467*/;
assign _20209_ = D[24] ^ Q[12] /*9463*/;
assign _20206_ = _19658_ & _20209_ /*9459*/;
assign _20207_ = _19658_ ^ _20209_ /*9462*/;
assign _20208_ = _20200_ & _20207_ /*9460*/;
assign _20205_ = _20206_ | _20208_ /*9458*/;
assign _20044_ = _20200_ ^ _20207_ /*9461*/;
assign _20214_ = D[25] ^ Q[12] /*9457*/;
assign _20211_ = _19659_ & _20214_ /*9453*/;
assign _20212_ = _19659_ ^ _20214_ /*9456*/;
assign _20213_ = _20205_ & _20212_ /*9454*/;
assign _20210_ = _20211_ | _20213_ /*9452*/;
assign _20045_ = _20205_ ^ _20212_ /*9455*/;
assign _20219_ = D[26] ^ Q[12] /*9451*/;
assign _20216_ = _19660_ & _20219_ /*9447*/;
assign _20217_ = _19660_ ^ _20219_ /*9450*/;
assign _20218_ = _20210_ & _20217_ /*9448*/;
assign _20215_ = _20216_ | _20218_ /*9446*/;
assign _20046_ = _20210_ ^ _20217_ /*9449*/;
assign _20224_ = D[27] ^ Q[12] /*9445*/;
assign _20221_ = _19661_ & _20224_ /*9441*/;
assign _20222_ = _19661_ ^ _20224_ /*9444*/;
assign _20223_ = _20215_ & _20222_ /*9442*/;
assign _20220_ = _20221_ | _20223_ /*9440*/;
assign _20047_ = _20215_ ^ _20222_ /*9443*/;
assign _20229_ = D[28] ^ Q[12] /*9439*/;
assign _20226_ = _19662_ & _20229_ /*9435*/;
assign _20227_ = _19662_ ^ _20229_ /*9438*/;
assign _20228_ = _20220_ & _20227_ /*9436*/;
assign _20225_ = _20226_ | _20228_ /*9434*/;
assign _20048_ = _20220_ ^ _20227_ /*9437*/;
assign _20234_ = D[29] ^ Q[12] /*9433*/;
assign _20231_ = _19663_ & _20234_ /*9429*/;
assign _20232_ = _19663_ ^ _20234_ /*9432*/;
assign _20233_ = _20225_ & _20232_ /*9430*/;
assign _20230_ = _20231_ | _20233_ /*9428*/;
assign _20049_ = _20225_ ^ _20232_ /*9431*/;
assign _20239_ = D[30] ^ Q[12] /*9427*/;
assign _20236_ = _19664_ & _20239_ /*9423*/;
assign _20237_ = _19664_ ^ _20239_ /*9426*/;
assign _20238_ = _20230_ & _20237_ /*9424*/;
assign _20235_ = _20236_ | _20238_ /*9422*/;
assign _20050_ = _20230_ ^ _20237_ /*9425*/;
assign _20244_ = D[31] ^ Q[12] /*9421*/;
assign _20241_ = _19665_ & _20244_ /*9417*/;
assign _20242_ = _19665_ ^ _20244_ /*9420*/;
assign _20243_ = _20235_ & _20242_ /*9418*/;
assign _20240_ = _20241_ | _20243_ /*9416*/;
assign _20051_ = _20235_ ^ _20242_ /*9419*/;
assign _20249_ = D[32] ^ Q[12] /*9415*/;
assign _20246_ = _19666_ & _20249_ /*9411*/;
assign _20247_ = _19666_ ^ _20249_ /*9414*/;
assign _20248_ = _20240_ & _20247_ /*9412*/;
assign _20245_ = _20246_ | _20248_ /*9410*/;
assign _20052_ = _20240_ ^ _20247_ /*9413*/;
assign _20254_ = D[33] ^ Q[12] /*9409*/;
assign _20251_ = _19667_ & _20254_ /*9405*/;
assign _20252_ = _19667_ ^ _20254_ /*9408*/;
assign _20253_ = _20245_ & _20252_ /*9406*/;
assign _20250_ = _20251_ | _20253_ /*9404*/;
assign _20053_ = _20245_ ^ _20252_ /*9407*/;
assign _20259_ = D[34] ^ Q[12] /*9403*/;
assign _20256_ = _19668_ & _20259_ /*9399*/;
assign _20257_ = _19668_ ^ _20259_ /*9402*/;
assign _20258_ = _20250_ & _20257_ /*9400*/;
assign _20255_ = _20256_ | _20258_ /*9398*/;
assign _20054_ = _20250_ ^ _20257_ /*9401*/;
assign _20264_ = D[35] ^ Q[12] /*9397*/;
assign _20261_ = _19669_ & _20264_ /*9393*/;
assign _20262_ = _19669_ ^ _20264_ /*9396*/;
assign _20263_ = _20255_ & _20262_ /*9394*/;
assign _20260_ = _20261_ | _20263_ /*9392*/;
assign _20055_ = _20255_ ^ _20262_ /*9395*/;
assign _20269_ = D[36] ^ Q[12] /*9391*/;
assign _20266_ = _19670_ & _20269_ /*9387*/;
assign _20267_ = _19670_ ^ _20269_ /*9390*/;
assign _20268_ = _20260_ & _20267_ /*9388*/;
assign _20265_ = _20266_ | _20268_ /*9386*/;
assign _20056_ = _20260_ ^ _20267_ /*9389*/;
assign _20274_ = D[37] ^ Q[12] /*9385*/;
assign _20271_ = _19671_ & _20274_ /*9381*/;
assign _20272_ = _19671_ ^ _20274_ /*9384*/;
assign _20273_ = _20265_ & _20272_ /*9382*/;
assign _20270_ = _20271_ | _20273_ /*9380*/;
assign _20057_ = _20265_ ^ _20272_ /*9383*/;
assign _20279_ = D[38] ^ Q[12] /*9379*/;
assign _20276_ = _19672_ & _20279_ /*9375*/;
assign _20277_ = _19672_ ^ _20279_ /*9378*/;
assign _20278_ = _20270_ & _20277_ /*9376*/;
assign _20275_ = _20276_ | _20278_ /*9374*/;
assign _20058_ = _20270_ ^ _20277_ /*9377*/;
assign _20284_ = D[39] ^ Q[12] /*9373*/;
assign _20281_ = _19673_ & _20284_ /*9369*/;
assign _20282_ = _19673_ ^ _20284_ /*9372*/;
assign _20283_ = _20275_ & _20282_ /*9370*/;
assign _20280_ = _20281_ | _20283_ /*9368*/;
assign _20059_ = _20275_ ^ _20282_ /*9371*/;
assign _20289_ = D[40] ^ Q[12] /*9367*/;
assign _20286_ = _19674_ & _20289_ /*9363*/;
assign _20287_ = _19674_ ^ _20289_ /*9366*/;
assign _20288_ = _20280_ & _20287_ /*9364*/;
assign _20285_ = _20286_ | _20288_ /*9362*/;
assign _20060_ = _20280_ ^ _20287_ /*9365*/;
assign _20294_ = D[41] ^ Q[12] /*9361*/;
assign _20291_ = _19675_ & _20294_ /*9357*/;
assign _20292_ = _19675_ ^ _20294_ /*9360*/;
assign _20293_ = _20285_ & _20292_ /*9358*/;
assign _20290_ = _20291_ | _20293_ /*9356*/;
assign _20061_ = _20285_ ^ _20292_ /*9359*/;
assign _20299_ = D[42] ^ Q[12] /*9355*/;
assign _20296_ = _19676_ & _20299_ /*9351*/;
assign _20297_ = _19676_ ^ _20299_ /*9354*/;
assign _20298_ = _20290_ & _20297_ /*9352*/;
assign _20295_ = _20296_ | _20298_ /*9350*/;
assign _20062_ = _20290_ ^ _20297_ /*9353*/;
assign _20304_ = D[43] ^ Q[12] /*9349*/;
assign _20301_ = _19677_ & _20304_ /*9345*/;
assign _20302_ = _19677_ ^ _20304_ /*9348*/;
assign _20303_ = _20295_ & _20302_ /*9346*/;
assign _20300_ = _20301_ | _20303_ /*9344*/;
assign _20063_ = _20295_ ^ _20302_ /*9347*/;
assign _20309_ = D[44] ^ Q[12] /*9343*/;
assign _20306_ = _19678_ & _20309_ /*9339*/;
assign _20307_ = _19678_ ^ _20309_ /*9342*/;
assign _20308_ = _20300_ & _20307_ /*9340*/;
assign _20305_ = _20306_ | _20308_ /*9338*/;
assign _20064_ = _20300_ ^ _20307_ /*9341*/;
assign _20314_ = D[45] ^ Q[12] /*9337*/;
assign _20311_ = _19679_ & _20314_ /*9333*/;
assign _20312_ = _19679_ ^ _20314_ /*9336*/;
assign _20313_ = _20305_ & _20312_ /*9334*/;
assign _20310_ = _20311_ | _20313_ /*9332*/;
assign _20065_ = _20305_ ^ _20312_ /*9335*/;
assign _20319_ = D[46] ^ Q[12] /*9331*/;
assign _20316_ = _19680_ & _20319_ /*9327*/;
assign _20317_ = _19680_ ^ _20319_ /*9330*/;
assign _20318_ = _20310_ & _20317_ /*9328*/;
assign _20315_ = _20316_ | _20318_ /*9326*/;
assign _20066_ = _20310_ ^ _20317_ /*9329*/;
assign _20324_ = D[47] ^ Q[12] /*9325*/;
assign _20321_ = _19681_ & _20324_ /*9321*/;
assign _20322_ = _19681_ ^ _20324_ /*9324*/;
assign _20323_ = _20315_ & _20322_ /*9322*/;
assign _20320_ = _20321_ | _20323_ /*9320*/;
assign _20067_ = _20315_ ^ _20322_ /*9323*/;
assign _20329_ = D[48] ^ Q[12] /*9319*/;
assign _20326_ = _19682_ & _20329_ /*9315*/;
assign _20327_ = _19682_ ^ _20329_ /*9318*/;
assign _20328_ = _20320_ & _20327_ /*9316*/;
assign _20325_ = _20326_ | _20328_ /*9314*/;
assign _20068_ = _20320_ ^ _20327_ /*9317*/;
assign _20334_ = D[49] ^ Q[12] /*9313*/;
assign _20331_ = _19683_ & _20334_ /*9309*/;
assign _20332_ = _19683_ ^ _20334_ /*9312*/;
assign _20333_ = _20325_ & _20332_ /*9310*/;
assign _20330_ = _20331_ | _20333_ /*9308*/;
assign _20069_ = _20325_ ^ _20332_ /*9311*/;
assign _20339_ = D[50] ^ Q[12] /*9307*/;
assign _20336_ = _19684_ & _20339_ /*9303*/;
assign _20337_ = _19684_ ^ _20339_ /*9306*/;
assign _20338_ = _20330_ & _20337_ /*9304*/;
assign _20335_ = _20336_ | _20338_ /*9302*/;
assign _20070_ = _20330_ ^ _20337_ /*9305*/;
assign _20344_ = D[51] ^ Q[12] /*9301*/;
assign _20341_ = _19685_ & _20344_ /*9297*/;
assign _20342_ = _19685_ ^ _20344_ /*9300*/;
assign _20343_ = _20335_ & _20342_ /*9298*/;
assign _20340_ = _20341_ | _20343_ /*9296*/;
assign _20071_ = _20335_ ^ _20342_ /*9299*/;
assign _20349_ = D[52] ^ Q[12] /*9295*/;
assign _20346_ = _19686_ & _20349_ /*9291*/;
assign _20347_ = _19686_ ^ _20349_ /*9294*/;
assign _20348_ = _20340_ & _20347_ /*9292*/;
assign _20345_ = _20346_ | _20348_ /*9290*/;
assign _20072_ = _20340_ ^ _20347_ /*9293*/;
assign _20354_ = D[53] ^ Q[12] /*9289*/;
assign _20351_ = _19687_ & _20354_ /*9285*/;
assign _20352_ = _19687_ ^ _20354_ /*9288*/;
assign _20353_ = _20345_ & _20352_ /*9286*/;
assign _20350_ = _20351_ | _20353_ /*9284*/;
assign _20073_ = _20345_ ^ _20352_ /*9287*/;
assign _20359_ = D[54] ^ Q[12] /*9283*/;
assign _20356_ = _19688_ & _20359_ /*9279*/;
assign _20357_ = _19688_ ^ _20359_ /*9282*/;
assign _20358_ = _20350_ & _20357_ /*9280*/;
assign _20355_ = _20356_ | _20358_ /*9278*/;
assign _20074_ = _20350_ ^ _20357_ /*9281*/;
assign _20364_ = D[55] ^ Q[12] /*9277*/;
assign _20361_ = _19689_ & _20364_ /*9273*/;
assign _20362_ = _19689_ ^ _20364_ /*9276*/;
assign _20363_ = _20355_ & _20362_ /*9274*/;
assign _20360_ = _20361_ | _20363_ /*9272*/;
assign _20075_ = _20355_ ^ _20362_ /*9275*/;
assign _20369_ = D[56] ^ Q[12] /*9271*/;
assign _20366_ = _19690_ & _20369_ /*9267*/;
assign _20367_ = _19690_ ^ _20369_ /*9270*/;
assign _20368_ = _20360_ & _20367_ /*9268*/;
assign _20365_ = _20366_ | _20368_ /*9266*/;
assign _20076_ = _20360_ ^ _20367_ /*9269*/;
assign _20374_ = D[57] ^ Q[12] /*9265*/;
assign _20371_ = _19691_ & _20374_ /*9261*/;
assign _20372_ = _19691_ ^ _20374_ /*9264*/;
assign _20373_ = _20365_ & _20372_ /*9262*/;
assign _20370_ = _20371_ | _20373_ /*9260*/;
assign _20077_ = _20365_ ^ _20372_ /*9263*/;
assign _20379_ = D[58] ^ Q[12] /*9259*/;
assign _20376_ = _19692_ & _20379_ /*9255*/;
assign _20377_ = _19692_ ^ _20379_ /*9258*/;
assign _20378_ = _20370_ & _20377_ /*9256*/;
assign _20375_ = _20376_ | _20378_ /*9254*/;
assign _20078_ = _20370_ ^ _20377_ /*9257*/;
assign _20384_ = D[59] ^ Q[12] /*9253*/;
assign _20381_ = _19693_ & _20384_ /*9249*/;
assign _20382_ = _19693_ ^ _20384_ /*9252*/;
assign _20383_ = _20375_ & _20382_ /*9250*/;
assign _20380_ = _20381_ | _20383_ /*9248*/;
assign _20079_ = _20375_ ^ _20382_ /*9251*/;
assign _20389_ = D[60] ^ Q[12] /*9247*/;
assign _20386_ = _19694_ & _20389_ /*9243*/;
assign _20387_ = _19694_ ^ _20389_ /*9246*/;
assign _20388_ = _20380_ & _20387_ /*9244*/;
assign _20385_ = _20386_ | _20388_ /*9242*/;
assign _20080_ = _20380_ ^ _20387_ /*9245*/;
assign _20394_ = D[61] ^ Q[12] /*9241*/;
assign _20391_ = _19695_ & _20394_ /*9237*/;
assign _20392_ = _19695_ ^ _20394_ /*9240*/;
assign _20393_ = _20385_ & _20392_ /*9238*/;
assign _20390_ = _20391_ | _20393_ /*9236*/;
assign _20081_ = _20385_ ^ _20392_ /*9239*/;
assign _20399_ = D[62] ^ Q[12] /*9235*/;
assign _20396_ = _19696_ & _20399_ /*9231*/;
assign _20397_ = _19696_ ^ _20399_ /*9234*/;
assign _20398_ = _20390_ & _20397_ /*9232*/;
assign _20395_ = _20396_ | _20398_ /*9230*/;
assign _20082_ = _20390_ ^ _20397_ /*9233*/;
assign _20403_ = zeroWire ^ Q[12] /*9229*/;
assign _20400_ = _19697_ & _20403_ /*9225*/;
assign _20401_ = _19697_ ^ _20403_ /*9228*/;
assign _20402_ = _20395_ & _20401_ /*9226*/;
assign Q[11] = _20400_ | _20402_ /*9224*/;
assign _20083_ = _20395_ ^ _20401_ /*9227*/;
assign _20474_ = D[0] ^ Q[11] /*8838*/;
assign _20471_ = R_0[10] & _20474_ /*8834*/;
assign _20472_ = R_0[10] ^ _20474_ /*8837*/;
assign _20473_ = Q[11] & _20472_ /*8835*/;
assign _20470_ = _20471_ | _20473_ /*8833*/;
assign _20405_ = Q[11] ^ _20472_ /*8836*/;
assign _20479_ = D[1] ^ Q[11] /*8832*/;
assign _20476_ = _20020_ & _20479_ /*8828*/;
assign _20477_ = _20020_ ^ _20479_ /*8831*/;
assign _20478_ = _20470_ & _20477_ /*8829*/;
assign _20475_ = _20476_ | _20478_ /*8827*/;
assign _20406_ = _20470_ ^ _20477_ /*8830*/;
assign _20484_ = D[2] ^ Q[11] /*8826*/;
assign _20481_ = _20021_ & _20484_ /*8822*/;
assign _20482_ = _20021_ ^ _20484_ /*8825*/;
assign _20483_ = _20475_ & _20482_ /*8823*/;
assign _20480_ = _20481_ | _20483_ /*8821*/;
assign _20407_ = _20475_ ^ _20482_ /*8824*/;
assign _20489_ = D[3] ^ Q[11] /*8820*/;
assign _20486_ = _20022_ & _20489_ /*8816*/;
assign _20487_ = _20022_ ^ _20489_ /*8819*/;
assign _20488_ = _20480_ & _20487_ /*8817*/;
assign _20485_ = _20486_ | _20488_ /*8815*/;
assign _20408_ = _20480_ ^ _20487_ /*8818*/;
assign _20494_ = D[4] ^ Q[11] /*8814*/;
assign _20491_ = _20023_ & _20494_ /*8810*/;
assign _20492_ = _20023_ ^ _20494_ /*8813*/;
assign _20493_ = _20485_ & _20492_ /*8811*/;
assign _20490_ = _20491_ | _20493_ /*8809*/;
assign _20409_ = _20485_ ^ _20492_ /*8812*/;
assign _20499_ = D[5] ^ Q[11] /*8808*/;
assign _20496_ = _20024_ & _20499_ /*8804*/;
assign _20497_ = _20024_ ^ _20499_ /*8807*/;
assign _20498_ = _20490_ & _20497_ /*8805*/;
assign _20495_ = _20496_ | _20498_ /*8803*/;
assign _20410_ = _20490_ ^ _20497_ /*8806*/;
assign _20504_ = D[6] ^ Q[11] /*8802*/;
assign _20501_ = _20025_ & _20504_ /*8798*/;
assign _20502_ = _20025_ ^ _20504_ /*8801*/;
assign _20503_ = _20495_ & _20502_ /*8799*/;
assign _20500_ = _20501_ | _20503_ /*8797*/;
assign _20411_ = _20495_ ^ _20502_ /*8800*/;
assign _20509_ = D[7] ^ Q[11] /*8796*/;
assign _20506_ = _20026_ & _20509_ /*8792*/;
assign _20507_ = _20026_ ^ _20509_ /*8795*/;
assign _20508_ = _20500_ & _20507_ /*8793*/;
assign _20505_ = _20506_ | _20508_ /*8791*/;
assign _20412_ = _20500_ ^ _20507_ /*8794*/;
assign _20514_ = D[8] ^ Q[11] /*8790*/;
assign _20511_ = _20027_ & _20514_ /*8786*/;
assign _20512_ = _20027_ ^ _20514_ /*8789*/;
assign _20513_ = _20505_ & _20512_ /*8787*/;
assign _20510_ = _20511_ | _20513_ /*8785*/;
assign _20413_ = _20505_ ^ _20512_ /*8788*/;
assign _20519_ = D[9] ^ Q[11] /*8784*/;
assign _20516_ = _20028_ & _20519_ /*8780*/;
assign _20517_ = _20028_ ^ _20519_ /*8783*/;
assign _20518_ = _20510_ & _20517_ /*8781*/;
assign _20515_ = _20516_ | _20518_ /*8779*/;
assign _20414_ = _20510_ ^ _20517_ /*8782*/;
assign _20524_ = D[10] ^ Q[11] /*8778*/;
assign _20521_ = _20029_ & _20524_ /*8774*/;
assign _20522_ = _20029_ ^ _20524_ /*8777*/;
assign _20523_ = _20515_ & _20522_ /*8775*/;
assign _20520_ = _20521_ | _20523_ /*8773*/;
assign _20415_ = _20515_ ^ _20522_ /*8776*/;
assign _20529_ = D[11] ^ Q[11] /*8772*/;
assign _20526_ = _20030_ & _20529_ /*8768*/;
assign _20527_ = _20030_ ^ _20529_ /*8771*/;
assign _20528_ = _20520_ & _20527_ /*8769*/;
assign _20525_ = _20526_ | _20528_ /*8767*/;
assign _20416_ = _20520_ ^ _20527_ /*8770*/;
assign _20534_ = D[12] ^ Q[11] /*8766*/;
assign _20531_ = _20031_ & _20534_ /*8762*/;
assign _20532_ = _20031_ ^ _20534_ /*8765*/;
assign _20533_ = _20525_ & _20532_ /*8763*/;
assign _20530_ = _20531_ | _20533_ /*8761*/;
assign _20417_ = _20525_ ^ _20532_ /*8764*/;
assign _20539_ = D[13] ^ Q[11] /*8760*/;
assign _20536_ = _20032_ & _20539_ /*8756*/;
assign _20537_ = _20032_ ^ _20539_ /*8759*/;
assign _20538_ = _20530_ & _20537_ /*8757*/;
assign _20535_ = _20536_ | _20538_ /*8755*/;
assign _20418_ = _20530_ ^ _20537_ /*8758*/;
assign _20544_ = D[14] ^ Q[11] /*8754*/;
assign _20541_ = _20033_ & _20544_ /*8750*/;
assign _20542_ = _20033_ ^ _20544_ /*8753*/;
assign _20543_ = _20535_ & _20542_ /*8751*/;
assign _20540_ = _20541_ | _20543_ /*8749*/;
assign _20419_ = _20535_ ^ _20542_ /*8752*/;
assign _20549_ = D[15] ^ Q[11] /*8748*/;
assign _20546_ = _20034_ & _20549_ /*8744*/;
assign _20547_ = _20034_ ^ _20549_ /*8747*/;
assign _20548_ = _20540_ & _20547_ /*8745*/;
assign _20545_ = _20546_ | _20548_ /*8743*/;
assign _20420_ = _20540_ ^ _20547_ /*8746*/;
assign _20554_ = D[16] ^ Q[11] /*8742*/;
assign _20551_ = _20035_ & _20554_ /*8738*/;
assign _20552_ = _20035_ ^ _20554_ /*8741*/;
assign _20553_ = _20545_ & _20552_ /*8739*/;
assign _20550_ = _20551_ | _20553_ /*8737*/;
assign _20421_ = _20545_ ^ _20552_ /*8740*/;
assign _20559_ = D[17] ^ Q[11] /*8736*/;
assign _20556_ = _20036_ & _20559_ /*8732*/;
assign _20557_ = _20036_ ^ _20559_ /*8735*/;
assign _20558_ = _20550_ & _20557_ /*8733*/;
assign _20555_ = _20556_ | _20558_ /*8731*/;
assign _20422_ = _20550_ ^ _20557_ /*8734*/;
assign _20564_ = D[18] ^ Q[11] /*8730*/;
assign _20561_ = _20037_ & _20564_ /*8726*/;
assign _20562_ = _20037_ ^ _20564_ /*8729*/;
assign _20563_ = _20555_ & _20562_ /*8727*/;
assign _20560_ = _20561_ | _20563_ /*8725*/;
assign _20423_ = _20555_ ^ _20562_ /*8728*/;
assign _20569_ = D[19] ^ Q[11] /*8724*/;
assign _20566_ = _20038_ & _20569_ /*8720*/;
assign _20567_ = _20038_ ^ _20569_ /*8723*/;
assign _20568_ = _20560_ & _20567_ /*8721*/;
assign _20565_ = _20566_ | _20568_ /*8719*/;
assign _20424_ = _20560_ ^ _20567_ /*8722*/;
assign _20574_ = D[20] ^ Q[11] /*8718*/;
assign _20571_ = _20039_ & _20574_ /*8714*/;
assign _20572_ = _20039_ ^ _20574_ /*8717*/;
assign _20573_ = _20565_ & _20572_ /*8715*/;
assign _20570_ = _20571_ | _20573_ /*8713*/;
assign _20425_ = _20565_ ^ _20572_ /*8716*/;
assign _20579_ = D[21] ^ Q[11] /*8712*/;
assign _20576_ = _20040_ & _20579_ /*8708*/;
assign _20577_ = _20040_ ^ _20579_ /*8711*/;
assign _20578_ = _20570_ & _20577_ /*8709*/;
assign _20575_ = _20576_ | _20578_ /*8707*/;
assign _20426_ = _20570_ ^ _20577_ /*8710*/;
assign _20584_ = D[22] ^ Q[11] /*8706*/;
assign _20581_ = _20041_ & _20584_ /*8702*/;
assign _20582_ = _20041_ ^ _20584_ /*8705*/;
assign _20583_ = _20575_ & _20582_ /*8703*/;
assign _20580_ = _20581_ | _20583_ /*8701*/;
assign _20427_ = _20575_ ^ _20582_ /*8704*/;
assign _20589_ = D[23] ^ Q[11] /*8700*/;
assign _20586_ = _20042_ & _20589_ /*8696*/;
assign _20587_ = _20042_ ^ _20589_ /*8699*/;
assign _20588_ = _20580_ & _20587_ /*8697*/;
assign _20585_ = _20586_ | _20588_ /*8695*/;
assign _20428_ = _20580_ ^ _20587_ /*8698*/;
assign _20594_ = D[24] ^ Q[11] /*8694*/;
assign _20591_ = _20043_ & _20594_ /*8690*/;
assign _20592_ = _20043_ ^ _20594_ /*8693*/;
assign _20593_ = _20585_ & _20592_ /*8691*/;
assign _20590_ = _20591_ | _20593_ /*8689*/;
assign _20429_ = _20585_ ^ _20592_ /*8692*/;
assign _20599_ = D[25] ^ Q[11] /*8688*/;
assign _20596_ = _20044_ & _20599_ /*8684*/;
assign _20597_ = _20044_ ^ _20599_ /*8687*/;
assign _20598_ = _20590_ & _20597_ /*8685*/;
assign _20595_ = _20596_ | _20598_ /*8683*/;
assign _20430_ = _20590_ ^ _20597_ /*8686*/;
assign _20604_ = D[26] ^ Q[11] /*8682*/;
assign _20601_ = _20045_ & _20604_ /*8678*/;
assign _20602_ = _20045_ ^ _20604_ /*8681*/;
assign _20603_ = _20595_ & _20602_ /*8679*/;
assign _20600_ = _20601_ | _20603_ /*8677*/;
assign _20431_ = _20595_ ^ _20602_ /*8680*/;
assign _20609_ = D[27] ^ Q[11] /*8676*/;
assign _20606_ = _20046_ & _20609_ /*8672*/;
assign _20607_ = _20046_ ^ _20609_ /*8675*/;
assign _20608_ = _20600_ & _20607_ /*8673*/;
assign _20605_ = _20606_ | _20608_ /*8671*/;
assign _20432_ = _20600_ ^ _20607_ /*8674*/;
assign _20614_ = D[28] ^ Q[11] /*8670*/;
assign _20611_ = _20047_ & _20614_ /*8666*/;
assign _20612_ = _20047_ ^ _20614_ /*8669*/;
assign _20613_ = _20605_ & _20612_ /*8667*/;
assign _20610_ = _20611_ | _20613_ /*8665*/;
assign _20433_ = _20605_ ^ _20612_ /*8668*/;
assign _20619_ = D[29] ^ Q[11] /*8664*/;
assign _20616_ = _20048_ & _20619_ /*8660*/;
assign _20617_ = _20048_ ^ _20619_ /*8663*/;
assign _20618_ = _20610_ & _20617_ /*8661*/;
assign _20615_ = _20616_ | _20618_ /*8659*/;
assign _20434_ = _20610_ ^ _20617_ /*8662*/;
assign _20624_ = D[30] ^ Q[11] /*8658*/;
assign _20621_ = _20049_ & _20624_ /*8654*/;
assign _20622_ = _20049_ ^ _20624_ /*8657*/;
assign _20623_ = _20615_ & _20622_ /*8655*/;
assign _20620_ = _20621_ | _20623_ /*8653*/;
assign _20435_ = _20615_ ^ _20622_ /*8656*/;
assign _20629_ = D[31] ^ Q[11] /*8652*/;
assign _20626_ = _20050_ & _20629_ /*8648*/;
assign _20627_ = _20050_ ^ _20629_ /*8651*/;
assign _20628_ = _20620_ & _20627_ /*8649*/;
assign _20625_ = _20626_ | _20628_ /*8647*/;
assign _20436_ = _20620_ ^ _20627_ /*8650*/;
assign _20634_ = D[32] ^ Q[11] /*8646*/;
assign _20631_ = _20051_ & _20634_ /*8642*/;
assign _20632_ = _20051_ ^ _20634_ /*8645*/;
assign _20633_ = _20625_ & _20632_ /*8643*/;
assign _20630_ = _20631_ | _20633_ /*8641*/;
assign _20437_ = _20625_ ^ _20632_ /*8644*/;
assign _20639_ = D[33] ^ Q[11] /*8640*/;
assign _20636_ = _20052_ & _20639_ /*8636*/;
assign _20637_ = _20052_ ^ _20639_ /*8639*/;
assign _20638_ = _20630_ & _20637_ /*8637*/;
assign _20635_ = _20636_ | _20638_ /*8635*/;
assign _20438_ = _20630_ ^ _20637_ /*8638*/;
assign _20644_ = D[34] ^ Q[11] /*8634*/;
assign _20641_ = _20053_ & _20644_ /*8630*/;
assign _20642_ = _20053_ ^ _20644_ /*8633*/;
assign _20643_ = _20635_ & _20642_ /*8631*/;
assign _20640_ = _20641_ | _20643_ /*8629*/;
assign _20439_ = _20635_ ^ _20642_ /*8632*/;
assign _20649_ = D[35] ^ Q[11] /*8628*/;
assign _20646_ = _20054_ & _20649_ /*8624*/;
assign _20647_ = _20054_ ^ _20649_ /*8627*/;
assign _20648_ = _20640_ & _20647_ /*8625*/;
assign _20645_ = _20646_ | _20648_ /*8623*/;
assign _20440_ = _20640_ ^ _20647_ /*8626*/;
assign _20654_ = D[36] ^ Q[11] /*8622*/;
assign _20651_ = _20055_ & _20654_ /*8618*/;
assign _20652_ = _20055_ ^ _20654_ /*8621*/;
assign _20653_ = _20645_ & _20652_ /*8619*/;
assign _20650_ = _20651_ | _20653_ /*8617*/;
assign _20441_ = _20645_ ^ _20652_ /*8620*/;
assign _20659_ = D[37] ^ Q[11] /*8616*/;
assign _20656_ = _20056_ & _20659_ /*8612*/;
assign _20657_ = _20056_ ^ _20659_ /*8615*/;
assign _20658_ = _20650_ & _20657_ /*8613*/;
assign _20655_ = _20656_ | _20658_ /*8611*/;
assign _20442_ = _20650_ ^ _20657_ /*8614*/;
assign _20664_ = D[38] ^ Q[11] /*8610*/;
assign _20661_ = _20057_ & _20664_ /*8606*/;
assign _20662_ = _20057_ ^ _20664_ /*8609*/;
assign _20663_ = _20655_ & _20662_ /*8607*/;
assign _20660_ = _20661_ | _20663_ /*8605*/;
assign _20443_ = _20655_ ^ _20662_ /*8608*/;
assign _20669_ = D[39] ^ Q[11] /*8604*/;
assign _20666_ = _20058_ & _20669_ /*8600*/;
assign _20667_ = _20058_ ^ _20669_ /*8603*/;
assign _20668_ = _20660_ & _20667_ /*8601*/;
assign _20665_ = _20666_ | _20668_ /*8599*/;
assign _20444_ = _20660_ ^ _20667_ /*8602*/;
assign _20674_ = D[40] ^ Q[11] /*8598*/;
assign _20671_ = _20059_ & _20674_ /*8594*/;
assign _20672_ = _20059_ ^ _20674_ /*8597*/;
assign _20673_ = _20665_ & _20672_ /*8595*/;
assign _20670_ = _20671_ | _20673_ /*8593*/;
assign _20445_ = _20665_ ^ _20672_ /*8596*/;
assign _20679_ = D[41] ^ Q[11] /*8592*/;
assign _20676_ = _20060_ & _20679_ /*8588*/;
assign _20677_ = _20060_ ^ _20679_ /*8591*/;
assign _20678_ = _20670_ & _20677_ /*8589*/;
assign _20675_ = _20676_ | _20678_ /*8587*/;
assign _20446_ = _20670_ ^ _20677_ /*8590*/;
assign _20684_ = D[42] ^ Q[11] /*8586*/;
assign _20681_ = _20061_ & _20684_ /*8582*/;
assign _20682_ = _20061_ ^ _20684_ /*8585*/;
assign _20683_ = _20675_ & _20682_ /*8583*/;
assign _20680_ = _20681_ | _20683_ /*8581*/;
assign _20447_ = _20675_ ^ _20682_ /*8584*/;
assign _20689_ = D[43] ^ Q[11] /*8580*/;
assign _20686_ = _20062_ & _20689_ /*8576*/;
assign _20687_ = _20062_ ^ _20689_ /*8579*/;
assign _20688_ = _20680_ & _20687_ /*8577*/;
assign _20685_ = _20686_ | _20688_ /*8575*/;
assign _20448_ = _20680_ ^ _20687_ /*8578*/;
assign _20694_ = D[44] ^ Q[11] /*8574*/;
assign _20691_ = _20063_ & _20694_ /*8570*/;
assign _20692_ = _20063_ ^ _20694_ /*8573*/;
assign _20693_ = _20685_ & _20692_ /*8571*/;
assign _20690_ = _20691_ | _20693_ /*8569*/;
assign _20449_ = _20685_ ^ _20692_ /*8572*/;
assign _20699_ = D[45] ^ Q[11] /*8568*/;
assign _20696_ = _20064_ & _20699_ /*8564*/;
assign _20697_ = _20064_ ^ _20699_ /*8567*/;
assign _20698_ = _20690_ & _20697_ /*8565*/;
assign _20695_ = _20696_ | _20698_ /*8563*/;
assign _20450_ = _20690_ ^ _20697_ /*8566*/;
assign _20704_ = D[46] ^ Q[11] /*8562*/;
assign _20701_ = _20065_ & _20704_ /*8558*/;
assign _20702_ = _20065_ ^ _20704_ /*8561*/;
assign _20703_ = _20695_ & _20702_ /*8559*/;
assign _20700_ = _20701_ | _20703_ /*8557*/;
assign _20451_ = _20695_ ^ _20702_ /*8560*/;
assign _20709_ = D[47] ^ Q[11] /*8556*/;
assign _20706_ = _20066_ & _20709_ /*8552*/;
assign _20707_ = _20066_ ^ _20709_ /*8555*/;
assign _20708_ = _20700_ & _20707_ /*8553*/;
assign _20705_ = _20706_ | _20708_ /*8551*/;
assign _20452_ = _20700_ ^ _20707_ /*8554*/;
assign _20714_ = D[48] ^ Q[11] /*8550*/;
assign _20711_ = _20067_ & _20714_ /*8546*/;
assign _20712_ = _20067_ ^ _20714_ /*8549*/;
assign _20713_ = _20705_ & _20712_ /*8547*/;
assign _20710_ = _20711_ | _20713_ /*8545*/;
assign _20453_ = _20705_ ^ _20712_ /*8548*/;
assign _20719_ = D[49] ^ Q[11] /*8544*/;
assign _20716_ = _20068_ & _20719_ /*8540*/;
assign _20717_ = _20068_ ^ _20719_ /*8543*/;
assign _20718_ = _20710_ & _20717_ /*8541*/;
assign _20715_ = _20716_ | _20718_ /*8539*/;
assign _20454_ = _20710_ ^ _20717_ /*8542*/;
assign _20724_ = D[50] ^ Q[11] /*8538*/;
assign _20721_ = _20069_ & _20724_ /*8534*/;
assign _20722_ = _20069_ ^ _20724_ /*8537*/;
assign _20723_ = _20715_ & _20722_ /*8535*/;
assign _20720_ = _20721_ | _20723_ /*8533*/;
assign _20455_ = _20715_ ^ _20722_ /*8536*/;
assign _20729_ = D[51] ^ Q[11] /*8532*/;
assign _20726_ = _20070_ & _20729_ /*8528*/;
assign _20727_ = _20070_ ^ _20729_ /*8531*/;
assign _20728_ = _20720_ & _20727_ /*8529*/;
assign _20725_ = _20726_ | _20728_ /*8527*/;
assign _20456_ = _20720_ ^ _20727_ /*8530*/;
assign _20734_ = D[52] ^ Q[11] /*8526*/;
assign _20731_ = _20071_ & _20734_ /*8522*/;
assign _20732_ = _20071_ ^ _20734_ /*8525*/;
assign _20733_ = _20725_ & _20732_ /*8523*/;
assign _20730_ = _20731_ | _20733_ /*8521*/;
assign _20457_ = _20725_ ^ _20732_ /*8524*/;
assign _20739_ = D[53] ^ Q[11] /*8520*/;
assign _20736_ = _20072_ & _20739_ /*8516*/;
assign _20737_ = _20072_ ^ _20739_ /*8519*/;
assign _20738_ = _20730_ & _20737_ /*8517*/;
assign _20735_ = _20736_ | _20738_ /*8515*/;
assign _20458_ = _20730_ ^ _20737_ /*8518*/;
assign _20744_ = D[54] ^ Q[11] /*8514*/;
assign _20741_ = _20073_ & _20744_ /*8510*/;
assign _20742_ = _20073_ ^ _20744_ /*8513*/;
assign _20743_ = _20735_ & _20742_ /*8511*/;
assign _20740_ = _20741_ | _20743_ /*8509*/;
assign _20459_ = _20735_ ^ _20742_ /*8512*/;
assign _20749_ = D[55] ^ Q[11] /*8508*/;
assign _20746_ = _20074_ & _20749_ /*8504*/;
assign _20747_ = _20074_ ^ _20749_ /*8507*/;
assign _20748_ = _20740_ & _20747_ /*8505*/;
assign _20745_ = _20746_ | _20748_ /*8503*/;
assign _20460_ = _20740_ ^ _20747_ /*8506*/;
assign _20754_ = D[56] ^ Q[11] /*8502*/;
assign _20751_ = _20075_ & _20754_ /*8498*/;
assign _20752_ = _20075_ ^ _20754_ /*8501*/;
assign _20753_ = _20745_ & _20752_ /*8499*/;
assign _20750_ = _20751_ | _20753_ /*8497*/;
assign _20461_ = _20745_ ^ _20752_ /*8500*/;
assign _20759_ = D[57] ^ Q[11] /*8496*/;
assign _20756_ = _20076_ & _20759_ /*8492*/;
assign _20757_ = _20076_ ^ _20759_ /*8495*/;
assign _20758_ = _20750_ & _20757_ /*8493*/;
assign _20755_ = _20756_ | _20758_ /*8491*/;
assign _20462_ = _20750_ ^ _20757_ /*8494*/;
assign _20764_ = D[58] ^ Q[11] /*8490*/;
assign _20761_ = _20077_ & _20764_ /*8486*/;
assign _20762_ = _20077_ ^ _20764_ /*8489*/;
assign _20763_ = _20755_ & _20762_ /*8487*/;
assign _20760_ = _20761_ | _20763_ /*8485*/;
assign _20463_ = _20755_ ^ _20762_ /*8488*/;
assign _20769_ = D[59] ^ Q[11] /*8484*/;
assign _20766_ = _20078_ & _20769_ /*8480*/;
assign _20767_ = _20078_ ^ _20769_ /*8483*/;
assign _20768_ = _20760_ & _20767_ /*8481*/;
assign _20765_ = _20766_ | _20768_ /*8479*/;
assign _20464_ = _20760_ ^ _20767_ /*8482*/;
assign _20774_ = D[60] ^ Q[11] /*8478*/;
assign _20771_ = _20079_ & _20774_ /*8474*/;
assign _20772_ = _20079_ ^ _20774_ /*8477*/;
assign _20773_ = _20765_ & _20772_ /*8475*/;
assign _20770_ = _20771_ | _20773_ /*8473*/;
assign _20465_ = _20765_ ^ _20772_ /*8476*/;
assign _20779_ = D[61] ^ Q[11] /*8472*/;
assign _20776_ = _20080_ & _20779_ /*8468*/;
assign _20777_ = _20080_ ^ _20779_ /*8471*/;
assign _20778_ = _20770_ & _20777_ /*8469*/;
assign _20775_ = _20776_ | _20778_ /*8467*/;
assign _20466_ = _20770_ ^ _20777_ /*8470*/;
assign _20784_ = D[62] ^ Q[11] /*8466*/;
assign _20781_ = _20081_ & _20784_ /*8462*/;
assign _20782_ = _20081_ ^ _20784_ /*8465*/;
assign _20783_ = _20775_ & _20782_ /*8463*/;
assign _20780_ = _20781_ | _20783_ /*8461*/;
assign _20467_ = _20775_ ^ _20782_ /*8464*/;
assign _20788_ = zeroWire ^ Q[11] /*8460*/;
assign _20785_ = _20082_ & _20788_ /*8456*/;
assign _20786_ = _20082_ ^ _20788_ /*8459*/;
assign _20787_ = _20780_ & _20786_ /*8457*/;
assign Q[10] = _20785_ | _20787_ /*8455*/;
assign _20468_ = _20780_ ^ _20786_ /*8458*/;
assign _20859_ = D[0] ^ Q[10] /*8069*/;
assign _20856_ = R_0[9] & _20859_ /*8065*/;
assign _20857_ = R_0[9] ^ _20859_ /*8068*/;
assign _20858_ = Q[10] & _20857_ /*8066*/;
assign _20855_ = _20856_ | _20858_ /*8064*/;
assign _20790_ = Q[10] ^ _20857_ /*8067*/;
assign _20864_ = D[1] ^ Q[10] /*8063*/;
assign _20861_ = _20405_ & _20864_ /*8059*/;
assign _20862_ = _20405_ ^ _20864_ /*8062*/;
assign _20863_ = _20855_ & _20862_ /*8060*/;
assign _20860_ = _20861_ | _20863_ /*8058*/;
assign _20791_ = _20855_ ^ _20862_ /*8061*/;
assign _20869_ = D[2] ^ Q[10] /*8057*/;
assign _20866_ = _20406_ & _20869_ /*8053*/;
assign _20867_ = _20406_ ^ _20869_ /*8056*/;
assign _20868_ = _20860_ & _20867_ /*8054*/;
assign _20865_ = _20866_ | _20868_ /*8052*/;
assign _20792_ = _20860_ ^ _20867_ /*8055*/;
assign _20874_ = D[3] ^ Q[10] /*8051*/;
assign _20871_ = _20407_ & _20874_ /*8047*/;
assign _20872_ = _20407_ ^ _20874_ /*8050*/;
assign _20873_ = _20865_ & _20872_ /*8048*/;
assign _20870_ = _20871_ | _20873_ /*8046*/;
assign _20793_ = _20865_ ^ _20872_ /*8049*/;
assign _20879_ = D[4] ^ Q[10] /*8045*/;
assign _20876_ = _20408_ & _20879_ /*8041*/;
assign _20877_ = _20408_ ^ _20879_ /*8044*/;
assign _20878_ = _20870_ & _20877_ /*8042*/;
assign _20875_ = _20876_ | _20878_ /*8040*/;
assign _20794_ = _20870_ ^ _20877_ /*8043*/;
assign _20884_ = D[5] ^ Q[10] /*8039*/;
assign _20881_ = _20409_ & _20884_ /*8035*/;
assign _20882_ = _20409_ ^ _20884_ /*8038*/;
assign _20883_ = _20875_ & _20882_ /*8036*/;
assign _20880_ = _20881_ | _20883_ /*8034*/;
assign _20795_ = _20875_ ^ _20882_ /*8037*/;
assign _20889_ = D[6] ^ Q[10] /*8033*/;
assign _20886_ = _20410_ & _20889_ /*8029*/;
assign _20887_ = _20410_ ^ _20889_ /*8032*/;
assign _20888_ = _20880_ & _20887_ /*8030*/;
assign _20885_ = _20886_ | _20888_ /*8028*/;
assign _20796_ = _20880_ ^ _20887_ /*8031*/;
assign _20894_ = D[7] ^ Q[10] /*8027*/;
assign _20891_ = _20411_ & _20894_ /*8023*/;
assign _20892_ = _20411_ ^ _20894_ /*8026*/;
assign _20893_ = _20885_ & _20892_ /*8024*/;
assign _20890_ = _20891_ | _20893_ /*8022*/;
assign _20797_ = _20885_ ^ _20892_ /*8025*/;
assign _20899_ = D[8] ^ Q[10] /*8021*/;
assign _20896_ = _20412_ & _20899_ /*8017*/;
assign _20897_ = _20412_ ^ _20899_ /*8020*/;
assign _20898_ = _20890_ & _20897_ /*8018*/;
assign _20895_ = _20896_ | _20898_ /*8016*/;
assign _20798_ = _20890_ ^ _20897_ /*8019*/;
assign _20904_ = D[9] ^ Q[10] /*8015*/;
assign _20901_ = _20413_ & _20904_ /*8011*/;
assign _20902_ = _20413_ ^ _20904_ /*8014*/;
assign _20903_ = _20895_ & _20902_ /*8012*/;
assign _20900_ = _20901_ | _20903_ /*8010*/;
assign _20799_ = _20895_ ^ _20902_ /*8013*/;
assign _20909_ = D[10] ^ Q[10] /*8009*/;
assign _20906_ = _20414_ & _20909_ /*8005*/;
assign _20907_ = _20414_ ^ _20909_ /*8008*/;
assign _20908_ = _20900_ & _20907_ /*8006*/;
assign _20905_ = _20906_ | _20908_ /*8004*/;
assign _20800_ = _20900_ ^ _20907_ /*8007*/;
assign _20914_ = D[11] ^ Q[10] /*8003*/;
assign _20911_ = _20415_ & _20914_ /*7999*/;
assign _20912_ = _20415_ ^ _20914_ /*8002*/;
assign _20913_ = _20905_ & _20912_ /*8000*/;
assign _20910_ = _20911_ | _20913_ /*7998*/;
assign _20801_ = _20905_ ^ _20912_ /*8001*/;
assign _20919_ = D[12] ^ Q[10] /*7997*/;
assign _20916_ = _20416_ & _20919_ /*7993*/;
assign _20917_ = _20416_ ^ _20919_ /*7996*/;
assign _20918_ = _20910_ & _20917_ /*7994*/;
assign _20915_ = _20916_ | _20918_ /*7992*/;
assign _20802_ = _20910_ ^ _20917_ /*7995*/;
assign _20924_ = D[13] ^ Q[10] /*7991*/;
assign _20921_ = _20417_ & _20924_ /*7987*/;
assign _20922_ = _20417_ ^ _20924_ /*7990*/;
assign _20923_ = _20915_ & _20922_ /*7988*/;
assign _20920_ = _20921_ | _20923_ /*7986*/;
assign _20803_ = _20915_ ^ _20922_ /*7989*/;
assign _20929_ = D[14] ^ Q[10] /*7985*/;
assign _20926_ = _20418_ & _20929_ /*7981*/;
assign _20927_ = _20418_ ^ _20929_ /*7984*/;
assign _20928_ = _20920_ & _20927_ /*7982*/;
assign _20925_ = _20926_ | _20928_ /*7980*/;
assign _20804_ = _20920_ ^ _20927_ /*7983*/;
assign _20934_ = D[15] ^ Q[10] /*7979*/;
assign _20931_ = _20419_ & _20934_ /*7975*/;
assign _20932_ = _20419_ ^ _20934_ /*7978*/;
assign _20933_ = _20925_ & _20932_ /*7976*/;
assign _20930_ = _20931_ | _20933_ /*7974*/;
assign _20805_ = _20925_ ^ _20932_ /*7977*/;
assign _20939_ = D[16] ^ Q[10] /*7973*/;
assign _20936_ = _20420_ & _20939_ /*7969*/;
assign _20937_ = _20420_ ^ _20939_ /*7972*/;
assign _20938_ = _20930_ & _20937_ /*7970*/;
assign _20935_ = _20936_ | _20938_ /*7968*/;
assign _20806_ = _20930_ ^ _20937_ /*7971*/;
assign _20944_ = D[17] ^ Q[10] /*7967*/;
assign _20941_ = _20421_ & _20944_ /*7963*/;
assign _20942_ = _20421_ ^ _20944_ /*7966*/;
assign _20943_ = _20935_ & _20942_ /*7964*/;
assign _20940_ = _20941_ | _20943_ /*7962*/;
assign _20807_ = _20935_ ^ _20942_ /*7965*/;
assign _20949_ = D[18] ^ Q[10] /*7961*/;
assign _20946_ = _20422_ & _20949_ /*7957*/;
assign _20947_ = _20422_ ^ _20949_ /*7960*/;
assign _20948_ = _20940_ & _20947_ /*7958*/;
assign _20945_ = _20946_ | _20948_ /*7956*/;
assign _20808_ = _20940_ ^ _20947_ /*7959*/;
assign _20954_ = D[19] ^ Q[10] /*7955*/;
assign _20951_ = _20423_ & _20954_ /*7951*/;
assign _20952_ = _20423_ ^ _20954_ /*7954*/;
assign _20953_ = _20945_ & _20952_ /*7952*/;
assign _20950_ = _20951_ | _20953_ /*7950*/;
assign _20809_ = _20945_ ^ _20952_ /*7953*/;
assign _20959_ = D[20] ^ Q[10] /*7949*/;
assign _20956_ = _20424_ & _20959_ /*7945*/;
assign _20957_ = _20424_ ^ _20959_ /*7948*/;
assign _20958_ = _20950_ & _20957_ /*7946*/;
assign _20955_ = _20956_ | _20958_ /*7944*/;
assign _20810_ = _20950_ ^ _20957_ /*7947*/;
assign _20964_ = D[21] ^ Q[10] /*7943*/;
assign _20961_ = _20425_ & _20964_ /*7939*/;
assign _20962_ = _20425_ ^ _20964_ /*7942*/;
assign _20963_ = _20955_ & _20962_ /*7940*/;
assign _20960_ = _20961_ | _20963_ /*7938*/;
assign _20811_ = _20955_ ^ _20962_ /*7941*/;
assign _20969_ = D[22] ^ Q[10] /*7937*/;
assign _20966_ = _20426_ & _20969_ /*7933*/;
assign _20967_ = _20426_ ^ _20969_ /*7936*/;
assign _20968_ = _20960_ & _20967_ /*7934*/;
assign _20965_ = _20966_ | _20968_ /*7932*/;
assign _20812_ = _20960_ ^ _20967_ /*7935*/;
assign _20974_ = D[23] ^ Q[10] /*7931*/;
assign _20971_ = _20427_ & _20974_ /*7927*/;
assign _20972_ = _20427_ ^ _20974_ /*7930*/;
assign _20973_ = _20965_ & _20972_ /*7928*/;
assign _20970_ = _20971_ | _20973_ /*7926*/;
assign _20813_ = _20965_ ^ _20972_ /*7929*/;
assign _20979_ = D[24] ^ Q[10] /*7925*/;
assign _20976_ = _20428_ & _20979_ /*7921*/;
assign _20977_ = _20428_ ^ _20979_ /*7924*/;
assign _20978_ = _20970_ & _20977_ /*7922*/;
assign _20975_ = _20976_ | _20978_ /*7920*/;
assign _20814_ = _20970_ ^ _20977_ /*7923*/;
assign _20984_ = D[25] ^ Q[10] /*7919*/;
assign _20981_ = _20429_ & _20984_ /*7915*/;
assign _20982_ = _20429_ ^ _20984_ /*7918*/;
assign _20983_ = _20975_ & _20982_ /*7916*/;
assign _20980_ = _20981_ | _20983_ /*7914*/;
assign _20815_ = _20975_ ^ _20982_ /*7917*/;
assign _20989_ = D[26] ^ Q[10] /*7913*/;
assign _20986_ = _20430_ & _20989_ /*7909*/;
assign _20987_ = _20430_ ^ _20989_ /*7912*/;
assign _20988_ = _20980_ & _20987_ /*7910*/;
assign _20985_ = _20986_ | _20988_ /*7908*/;
assign _20816_ = _20980_ ^ _20987_ /*7911*/;
assign _20994_ = D[27] ^ Q[10] /*7907*/;
assign _20991_ = _20431_ & _20994_ /*7903*/;
assign _20992_ = _20431_ ^ _20994_ /*7906*/;
assign _20993_ = _20985_ & _20992_ /*7904*/;
assign _20990_ = _20991_ | _20993_ /*7902*/;
assign _20817_ = _20985_ ^ _20992_ /*7905*/;
assign _20999_ = D[28] ^ Q[10] /*7901*/;
assign _20996_ = _20432_ & _20999_ /*7897*/;
assign _20997_ = _20432_ ^ _20999_ /*7900*/;
assign _20998_ = _20990_ & _20997_ /*7898*/;
assign _20995_ = _20996_ | _20998_ /*7896*/;
assign _20818_ = _20990_ ^ _20997_ /*7899*/;
assign _21004_ = D[29] ^ Q[10] /*7895*/;
assign _21001_ = _20433_ & _21004_ /*7891*/;
assign _21002_ = _20433_ ^ _21004_ /*7894*/;
assign _21003_ = _20995_ & _21002_ /*7892*/;
assign _21000_ = _21001_ | _21003_ /*7890*/;
assign _20819_ = _20995_ ^ _21002_ /*7893*/;
assign _21009_ = D[30] ^ Q[10] /*7889*/;
assign _21006_ = _20434_ & _21009_ /*7885*/;
assign _21007_ = _20434_ ^ _21009_ /*7888*/;
assign _21008_ = _21000_ & _21007_ /*7886*/;
assign _21005_ = _21006_ | _21008_ /*7884*/;
assign _20820_ = _21000_ ^ _21007_ /*7887*/;
assign _21014_ = D[31] ^ Q[10] /*7883*/;
assign _21011_ = _20435_ & _21014_ /*7879*/;
assign _21012_ = _20435_ ^ _21014_ /*7882*/;
assign _21013_ = _21005_ & _21012_ /*7880*/;
assign _21010_ = _21011_ | _21013_ /*7878*/;
assign _20821_ = _21005_ ^ _21012_ /*7881*/;
assign _21019_ = D[32] ^ Q[10] /*7877*/;
assign _21016_ = _20436_ & _21019_ /*7873*/;
assign _21017_ = _20436_ ^ _21019_ /*7876*/;
assign _21018_ = _21010_ & _21017_ /*7874*/;
assign _21015_ = _21016_ | _21018_ /*7872*/;
assign _20822_ = _21010_ ^ _21017_ /*7875*/;
assign _21024_ = D[33] ^ Q[10] /*7871*/;
assign _21021_ = _20437_ & _21024_ /*7867*/;
assign _21022_ = _20437_ ^ _21024_ /*7870*/;
assign _21023_ = _21015_ & _21022_ /*7868*/;
assign _21020_ = _21021_ | _21023_ /*7866*/;
assign _20823_ = _21015_ ^ _21022_ /*7869*/;
assign _21029_ = D[34] ^ Q[10] /*7865*/;
assign _21026_ = _20438_ & _21029_ /*7861*/;
assign _21027_ = _20438_ ^ _21029_ /*7864*/;
assign _21028_ = _21020_ & _21027_ /*7862*/;
assign _21025_ = _21026_ | _21028_ /*7860*/;
assign _20824_ = _21020_ ^ _21027_ /*7863*/;
assign _21034_ = D[35] ^ Q[10] /*7859*/;
assign _21031_ = _20439_ & _21034_ /*7855*/;
assign _21032_ = _20439_ ^ _21034_ /*7858*/;
assign _21033_ = _21025_ & _21032_ /*7856*/;
assign _21030_ = _21031_ | _21033_ /*7854*/;
assign _20825_ = _21025_ ^ _21032_ /*7857*/;
assign _21039_ = D[36] ^ Q[10] /*7853*/;
assign _21036_ = _20440_ & _21039_ /*7849*/;
assign _21037_ = _20440_ ^ _21039_ /*7852*/;
assign _21038_ = _21030_ & _21037_ /*7850*/;
assign _21035_ = _21036_ | _21038_ /*7848*/;
assign _20826_ = _21030_ ^ _21037_ /*7851*/;
assign _21044_ = D[37] ^ Q[10] /*7847*/;
assign _21041_ = _20441_ & _21044_ /*7843*/;
assign _21042_ = _20441_ ^ _21044_ /*7846*/;
assign _21043_ = _21035_ & _21042_ /*7844*/;
assign _21040_ = _21041_ | _21043_ /*7842*/;
assign _20827_ = _21035_ ^ _21042_ /*7845*/;
assign _21049_ = D[38] ^ Q[10] /*7841*/;
assign _21046_ = _20442_ & _21049_ /*7837*/;
assign _21047_ = _20442_ ^ _21049_ /*7840*/;
assign _21048_ = _21040_ & _21047_ /*7838*/;
assign _21045_ = _21046_ | _21048_ /*7836*/;
assign _20828_ = _21040_ ^ _21047_ /*7839*/;
assign _21054_ = D[39] ^ Q[10] /*7835*/;
assign _21051_ = _20443_ & _21054_ /*7831*/;
assign _21052_ = _20443_ ^ _21054_ /*7834*/;
assign _21053_ = _21045_ & _21052_ /*7832*/;
assign _21050_ = _21051_ | _21053_ /*7830*/;
assign _20829_ = _21045_ ^ _21052_ /*7833*/;
assign _21059_ = D[40] ^ Q[10] /*7829*/;
assign _21056_ = _20444_ & _21059_ /*7825*/;
assign _21057_ = _20444_ ^ _21059_ /*7828*/;
assign _21058_ = _21050_ & _21057_ /*7826*/;
assign _21055_ = _21056_ | _21058_ /*7824*/;
assign _20830_ = _21050_ ^ _21057_ /*7827*/;
assign _21064_ = D[41] ^ Q[10] /*7823*/;
assign _21061_ = _20445_ & _21064_ /*7819*/;
assign _21062_ = _20445_ ^ _21064_ /*7822*/;
assign _21063_ = _21055_ & _21062_ /*7820*/;
assign _21060_ = _21061_ | _21063_ /*7818*/;
assign _20831_ = _21055_ ^ _21062_ /*7821*/;
assign _21069_ = D[42] ^ Q[10] /*7817*/;
assign _21066_ = _20446_ & _21069_ /*7813*/;
assign _21067_ = _20446_ ^ _21069_ /*7816*/;
assign _21068_ = _21060_ & _21067_ /*7814*/;
assign _21065_ = _21066_ | _21068_ /*7812*/;
assign _20832_ = _21060_ ^ _21067_ /*7815*/;
assign _21074_ = D[43] ^ Q[10] /*7811*/;
assign _21071_ = _20447_ & _21074_ /*7807*/;
assign _21072_ = _20447_ ^ _21074_ /*7810*/;
assign _21073_ = _21065_ & _21072_ /*7808*/;
assign _21070_ = _21071_ | _21073_ /*7806*/;
assign _20833_ = _21065_ ^ _21072_ /*7809*/;
assign _21079_ = D[44] ^ Q[10] /*7805*/;
assign _21076_ = _20448_ & _21079_ /*7801*/;
assign _21077_ = _20448_ ^ _21079_ /*7804*/;
assign _21078_ = _21070_ & _21077_ /*7802*/;
assign _21075_ = _21076_ | _21078_ /*7800*/;
assign _20834_ = _21070_ ^ _21077_ /*7803*/;
assign _21084_ = D[45] ^ Q[10] /*7799*/;
assign _21081_ = _20449_ & _21084_ /*7795*/;
assign _21082_ = _20449_ ^ _21084_ /*7798*/;
assign _21083_ = _21075_ & _21082_ /*7796*/;
assign _21080_ = _21081_ | _21083_ /*7794*/;
assign _20835_ = _21075_ ^ _21082_ /*7797*/;
assign _21089_ = D[46] ^ Q[10] /*7793*/;
assign _21086_ = _20450_ & _21089_ /*7789*/;
assign _21087_ = _20450_ ^ _21089_ /*7792*/;
assign _21088_ = _21080_ & _21087_ /*7790*/;
assign _21085_ = _21086_ | _21088_ /*7788*/;
assign _20836_ = _21080_ ^ _21087_ /*7791*/;
assign _21094_ = D[47] ^ Q[10] /*7787*/;
assign _21091_ = _20451_ & _21094_ /*7783*/;
assign _21092_ = _20451_ ^ _21094_ /*7786*/;
assign _21093_ = _21085_ & _21092_ /*7784*/;
assign _21090_ = _21091_ | _21093_ /*7782*/;
assign _20837_ = _21085_ ^ _21092_ /*7785*/;
assign _21099_ = D[48] ^ Q[10] /*7781*/;
assign _21096_ = _20452_ & _21099_ /*7777*/;
assign _21097_ = _20452_ ^ _21099_ /*7780*/;
assign _21098_ = _21090_ & _21097_ /*7778*/;
assign _21095_ = _21096_ | _21098_ /*7776*/;
assign _20838_ = _21090_ ^ _21097_ /*7779*/;
assign _21104_ = D[49] ^ Q[10] /*7775*/;
assign _21101_ = _20453_ & _21104_ /*7771*/;
assign _21102_ = _20453_ ^ _21104_ /*7774*/;
assign _21103_ = _21095_ & _21102_ /*7772*/;
assign _21100_ = _21101_ | _21103_ /*7770*/;
assign _20839_ = _21095_ ^ _21102_ /*7773*/;
assign _21109_ = D[50] ^ Q[10] /*7769*/;
assign _21106_ = _20454_ & _21109_ /*7765*/;
assign _21107_ = _20454_ ^ _21109_ /*7768*/;
assign _21108_ = _21100_ & _21107_ /*7766*/;
assign _21105_ = _21106_ | _21108_ /*7764*/;
assign _20840_ = _21100_ ^ _21107_ /*7767*/;
assign _21114_ = D[51] ^ Q[10] /*7763*/;
assign _21111_ = _20455_ & _21114_ /*7759*/;
assign _21112_ = _20455_ ^ _21114_ /*7762*/;
assign _21113_ = _21105_ & _21112_ /*7760*/;
assign _21110_ = _21111_ | _21113_ /*7758*/;
assign _20841_ = _21105_ ^ _21112_ /*7761*/;
assign _21119_ = D[52] ^ Q[10] /*7757*/;
assign _21116_ = _20456_ & _21119_ /*7753*/;
assign _21117_ = _20456_ ^ _21119_ /*7756*/;
assign _21118_ = _21110_ & _21117_ /*7754*/;
assign _21115_ = _21116_ | _21118_ /*7752*/;
assign _20842_ = _21110_ ^ _21117_ /*7755*/;
assign _21124_ = D[53] ^ Q[10] /*7751*/;
assign _21121_ = _20457_ & _21124_ /*7747*/;
assign _21122_ = _20457_ ^ _21124_ /*7750*/;
assign _21123_ = _21115_ & _21122_ /*7748*/;
assign _21120_ = _21121_ | _21123_ /*7746*/;
assign _20843_ = _21115_ ^ _21122_ /*7749*/;
assign _21129_ = D[54] ^ Q[10] /*7745*/;
assign _21126_ = _20458_ & _21129_ /*7741*/;
assign _21127_ = _20458_ ^ _21129_ /*7744*/;
assign _21128_ = _21120_ & _21127_ /*7742*/;
assign _21125_ = _21126_ | _21128_ /*7740*/;
assign _20844_ = _21120_ ^ _21127_ /*7743*/;
assign _21134_ = D[55] ^ Q[10] /*7739*/;
assign _21131_ = _20459_ & _21134_ /*7735*/;
assign _21132_ = _20459_ ^ _21134_ /*7738*/;
assign _21133_ = _21125_ & _21132_ /*7736*/;
assign _21130_ = _21131_ | _21133_ /*7734*/;
assign _20845_ = _21125_ ^ _21132_ /*7737*/;
assign _21139_ = D[56] ^ Q[10] /*7733*/;
assign _21136_ = _20460_ & _21139_ /*7729*/;
assign _21137_ = _20460_ ^ _21139_ /*7732*/;
assign _21138_ = _21130_ & _21137_ /*7730*/;
assign _21135_ = _21136_ | _21138_ /*7728*/;
assign _20846_ = _21130_ ^ _21137_ /*7731*/;
assign _21144_ = D[57] ^ Q[10] /*7727*/;
assign _21141_ = _20461_ & _21144_ /*7723*/;
assign _21142_ = _20461_ ^ _21144_ /*7726*/;
assign _21143_ = _21135_ & _21142_ /*7724*/;
assign _21140_ = _21141_ | _21143_ /*7722*/;
assign _20847_ = _21135_ ^ _21142_ /*7725*/;
assign _21149_ = D[58] ^ Q[10] /*7721*/;
assign _21146_ = _20462_ & _21149_ /*7717*/;
assign _21147_ = _20462_ ^ _21149_ /*7720*/;
assign _21148_ = _21140_ & _21147_ /*7718*/;
assign _21145_ = _21146_ | _21148_ /*7716*/;
assign _20848_ = _21140_ ^ _21147_ /*7719*/;
assign _21154_ = D[59] ^ Q[10] /*7715*/;
assign _21151_ = _20463_ & _21154_ /*7711*/;
assign _21152_ = _20463_ ^ _21154_ /*7714*/;
assign _21153_ = _21145_ & _21152_ /*7712*/;
assign _21150_ = _21151_ | _21153_ /*7710*/;
assign _20849_ = _21145_ ^ _21152_ /*7713*/;
assign _21159_ = D[60] ^ Q[10] /*7709*/;
assign _21156_ = _20464_ & _21159_ /*7705*/;
assign _21157_ = _20464_ ^ _21159_ /*7708*/;
assign _21158_ = _21150_ & _21157_ /*7706*/;
assign _21155_ = _21156_ | _21158_ /*7704*/;
assign _20850_ = _21150_ ^ _21157_ /*7707*/;
assign _21164_ = D[61] ^ Q[10] /*7703*/;
assign _21161_ = _20465_ & _21164_ /*7699*/;
assign _21162_ = _20465_ ^ _21164_ /*7702*/;
assign _21163_ = _21155_ & _21162_ /*7700*/;
assign _21160_ = _21161_ | _21163_ /*7698*/;
assign _20851_ = _21155_ ^ _21162_ /*7701*/;
assign _21169_ = D[62] ^ Q[10] /*7697*/;
assign _21166_ = _20466_ & _21169_ /*7693*/;
assign _21167_ = _20466_ ^ _21169_ /*7696*/;
assign _21168_ = _21160_ & _21167_ /*7694*/;
assign _21165_ = _21166_ | _21168_ /*7692*/;
assign _20852_ = _21160_ ^ _21167_ /*7695*/;
assign _21173_ = zeroWire ^ Q[10] /*7691*/;
assign _21170_ = _20467_ & _21173_ /*7687*/;
assign _21171_ = _20467_ ^ _21173_ /*7690*/;
assign _21172_ = _21165_ & _21171_ /*7688*/;
assign Q[9] = _21170_ | _21172_ /*7686*/;
assign _20853_ = _21165_ ^ _21171_ /*7689*/;
assign _21244_ = D[0] ^ Q[9] /*7300*/;
assign _21241_ = R_0[8] & _21244_ /*7296*/;
assign _21242_ = R_0[8] ^ _21244_ /*7299*/;
assign _21243_ = Q[9] & _21242_ /*7297*/;
assign _21240_ = _21241_ | _21243_ /*7295*/;
assign _21175_ = Q[9] ^ _21242_ /*7298*/;
assign _21249_ = D[1] ^ Q[9] /*7294*/;
assign _21246_ = _20790_ & _21249_ /*7290*/;
assign _21247_ = _20790_ ^ _21249_ /*7293*/;
assign _21248_ = _21240_ & _21247_ /*7291*/;
assign _21245_ = _21246_ | _21248_ /*7289*/;
assign _21176_ = _21240_ ^ _21247_ /*7292*/;
assign _21254_ = D[2] ^ Q[9] /*7288*/;
assign _21251_ = _20791_ & _21254_ /*7284*/;
assign _21252_ = _20791_ ^ _21254_ /*7287*/;
assign _21253_ = _21245_ & _21252_ /*7285*/;
assign _21250_ = _21251_ | _21253_ /*7283*/;
assign _21177_ = _21245_ ^ _21252_ /*7286*/;
assign _21259_ = D[3] ^ Q[9] /*7282*/;
assign _21256_ = _20792_ & _21259_ /*7278*/;
assign _21257_ = _20792_ ^ _21259_ /*7281*/;
assign _21258_ = _21250_ & _21257_ /*7279*/;
assign _21255_ = _21256_ | _21258_ /*7277*/;
assign _21178_ = _21250_ ^ _21257_ /*7280*/;
assign _21264_ = D[4] ^ Q[9] /*7276*/;
assign _21261_ = _20793_ & _21264_ /*7272*/;
assign _21262_ = _20793_ ^ _21264_ /*7275*/;
assign _21263_ = _21255_ & _21262_ /*7273*/;
assign _21260_ = _21261_ | _21263_ /*7271*/;
assign _21179_ = _21255_ ^ _21262_ /*7274*/;
assign _21269_ = D[5] ^ Q[9] /*7270*/;
assign _21266_ = _20794_ & _21269_ /*7266*/;
assign _21267_ = _20794_ ^ _21269_ /*7269*/;
assign _21268_ = _21260_ & _21267_ /*7267*/;
assign _21265_ = _21266_ | _21268_ /*7265*/;
assign _21180_ = _21260_ ^ _21267_ /*7268*/;
assign _21274_ = D[6] ^ Q[9] /*7264*/;
assign _21271_ = _20795_ & _21274_ /*7260*/;
assign _21272_ = _20795_ ^ _21274_ /*7263*/;
assign _21273_ = _21265_ & _21272_ /*7261*/;
assign _21270_ = _21271_ | _21273_ /*7259*/;
assign _21181_ = _21265_ ^ _21272_ /*7262*/;
assign _21279_ = D[7] ^ Q[9] /*7258*/;
assign _21276_ = _20796_ & _21279_ /*7254*/;
assign _21277_ = _20796_ ^ _21279_ /*7257*/;
assign _21278_ = _21270_ & _21277_ /*7255*/;
assign _21275_ = _21276_ | _21278_ /*7253*/;
assign _21182_ = _21270_ ^ _21277_ /*7256*/;
assign _21284_ = D[8] ^ Q[9] /*7252*/;
assign _21281_ = _20797_ & _21284_ /*7248*/;
assign _21282_ = _20797_ ^ _21284_ /*7251*/;
assign _21283_ = _21275_ & _21282_ /*7249*/;
assign _21280_ = _21281_ | _21283_ /*7247*/;
assign _21183_ = _21275_ ^ _21282_ /*7250*/;
assign _21289_ = D[9] ^ Q[9] /*7246*/;
assign _21286_ = _20798_ & _21289_ /*7242*/;
assign _21287_ = _20798_ ^ _21289_ /*7245*/;
assign _21288_ = _21280_ & _21287_ /*7243*/;
assign _21285_ = _21286_ | _21288_ /*7241*/;
assign _21184_ = _21280_ ^ _21287_ /*7244*/;
assign _21294_ = D[10] ^ Q[9] /*7240*/;
assign _21291_ = _20799_ & _21294_ /*7236*/;
assign _21292_ = _20799_ ^ _21294_ /*7239*/;
assign _21293_ = _21285_ & _21292_ /*7237*/;
assign _21290_ = _21291_ | _21293_ /*7235*/;
assign _21185_ = _21285_ ^ _21292_ /*7238*/;
assign _21299_ = D[11] ^ Q[9] /*7234*/;
assign _21296_ = _20800_ & _21299_ /*7230*/;
assign _21297_ = _20800_ ^ _21299_ /*7233*/;
assign _21298_ = _21290_ & _21297_ /*7231*/;
assign _21295_ = _21296_ | _21298_ /*7229*/;
assign _21186_ = _21290_ ^ _21297_ /*7232*/;
assign _21304_ = D[12] ^ Q[9] /*7228*/;
assign _21301_ = _20801_ & _21304_ /*7224*/;
assign _21302_ = _20801_ ^ _21304_ /*7227*/;
assign _21303_ = _21295_ & _21302_ /*7225*/;
assign _21300_ = _21301_ | _21303_ /*7223*/;
assign _21187_ = _21295_ ^ _21302_ /*7226*/;
assign _21309_ = D[13] ^ Q[9] /*7222*/;
assign _21306_ = _20802_ & _21309_ /*7218*/;
assign _21307_ = _20802_ ^ _21309_ /*7221*/;
assign _21308_ = _21300_ & _21307_ /*7219*/;
assign _21305_ = _21306_ | _21308_ /*7217*/;
assign _21188_ = _21300_ ^ _21307_ /*7220*/;
assign _21314_ = D[14] ^ Q[9] /*7216*/;
assign _21311_ = _20803_ & _21314_ /*7212*/;
assign _21312_ = _20803_ ^ _21314_ /*7215*/;
assign _21313_ = _21305_ & _21312_ /*7213*/;
assign _21310_ = _21311_ | _21313_ /*7211*/;
assign _21189_ = _21305_ ^ _21312_ /*7214*/;
assign _21319_ = D[15] ^ Q[9] /*7210*/;
assign _21316_ = _20804_ & _21319_ /*7206*/;
assign _21317_ = _20804_ ^ _21319_ /*7209*/;
assign _21318_ = _21310_ & _21317_ /*7207*/;
assign _21315_ = _21316_ | _21318_ /*7205*/;
assign _21190_ = _21310_ ^ _21317_ /*7208*/;
assign _21324_ = D[16] ^ Q[9] /*7204*/;
assign _21321_ = _20805_ & _21324_ /*7200*/;
assign _21322_ = _20805_ ^ _21324_ /*7203*/;
assign _21323_ = _21315_ & _21322_ /*7201*/;
assign _21320_ = _21321_ | _21323_ /*7199*/;
assign _21191_ = _21315_ ^ _21322_ /*7202*/;
assign _21329_ = D[17] ^ Q[9] /*7198*/;
assign _21326_ = _20806_ & _21329_ /*7194*/;
assign _21327_ = _20806_ ^ _21329_ /*7197*/;
assign _21328_ = _21320_ & _21327_ /*7195*/;
assign _21325_ = _21326_ | _21328_ /*7193*/;
assign _21192_ = _21320_ ^ _21327_ /*7196*/;
assign _21334_ = D[18] ^ Q[9] /*7192*/;
assign _21331_ = _20807_ & _21334_ /*7188*/;
assign _21332_ = _20807_ ^ _21334_ /*7191*/;
assign _21333_ = _21325_ & _21332_ /*7189*/;
assign _21330_ = _21331_ | _21333_ /*7187*/;
assign _21193_ = _21325_ ^ _21332_ /*7190*/;
assign _21339_ = D[19] ^ Q[9] /*7186*/;
assign _21336_ = _20808_ & _21339_ /*7182*/;
assign _21337_ = _20808_ ^ _21339_ /*7185*/;
assign _21338_ = _21330_ & _21337_ /*7183*/;
assign _21335_ = _21336_ | _21338_ /*7181*/;
assign _21194_ = _21330_ ^ _21337_ /*7184*/;
assign _21344_ = D[20] ^ Q[9] /*7180*/;
assign _21341_ = _20809_ & _21344_ /*7176*/;
assign _21342_ = _20809_ ^ _21344_ /*7179*/;
assign _21343_ = _21335_ & _21342_ /*7177*/;
assign _21340_ = _21341_ | _21343_ /*7175*/;
assign _21195_ = _21335_ ^ _21342_ /*7178*/;
assign _21349_ = D[21] ^ Q[9] /*7174*/;
assign _21346_ = _20810_ & _21349_ /*7170*/;
assign _21347_ = _20810_ ^ _21349_ /*7173*/;
assign _21348_ = _21340_ & _21347_ /*7171*/;
assign _21345_ = _21346_ | _21348_ /*7169*/;
assign _21196_ = _21340_ ^ _21347_ /*7172*/;
assign _21354_ = D[22] ^ Q[9] /*7168*/;
assign _21351_ = _20811_ & _21354_ /*7164*/;
assign _21352_ = _20811_ ^ _21354_ /*7167*/;
assign _21353_ = _21345_ & _21352_ /*7165*/;
assign _21350_ = _21351_ | _21353_ /*7163*/;
assign _21197_ = _21345_ ^ _21352_ /*7166*/;
assign _21359_ = D[23] ^ Q[9] /*7162*/;
assign _21356_ = _20812_ & _21359_ /*7158*/;
assign _21357_ = _20812_ ^ _21359_ /*7161*/;
assign _21358_ = _21350_ & _21357_ /*7159*/;
assign _21355_ = _21356_ | _21358_ /*7157*/;
assign _21198_ = _21350_ ^ _21357_ /*7160*/;
assign _21364_ = D[24] ^ Q[9] /*7156*/;
assign _21361_ = _20813_ & _21364_ /*7152*/;
assign _21362_ = _20813_ ^ _21364_ /*7155*/;
assign _21363_ = _21355_ & _21362_ /*7153*/;
assign _21360_ = _21361_ | _21363_ /*7151*/;
assign _21199_ = _21355_ ^ _21362_ /*7154*/;
assign _21369_ = D[25] ^ Q[9] /*7150*/;
assign _21366_ = _20814_ & _21369_ /*7146*/;
assign _21367_ = _20814_ ^ _21369_ /*7149*/;
assign _21368_ = _21360_ & _21367_ /*7147*/;
assign _21365_ = _21366_ | _21368_ /*7145*/;
assign _21200_ = _21360_ ^ _21367_ /*7148*/;
assign _21374_ = D[26] ^ Q[9] /*7144*/;
assign _21371_ = _20815_ & _21374_ /*7140*/;
assign _21372_ = _20815_ ^ _21374_ /*7143*/;
assign _21373_ = _21365_ & _21372_ /*7141*/;
assign _21370_ = _21371_ | _21373_ /*7139*/;
assign _21201_ = _21365_ ^ _21372_ /*7142*/;
assign _21379_ = D[27] ^ Q[9] /*7138*/;
assign _21376_ = _20816_ & _21379_ /*7134*/;
assign _21377_ = _20816_ ^ _21379_ /*7137*/;
assign _21378_ = _21370_ & _21377_ /*7135*/;
assign _21375_ = _21376_ | _21378_ /*7133*/;
assign _21202_ = _21370_ ^ _21377_ /*7136*/;
assign _21384_ = D[28] ^ Q[9] /*7132*/;
assign _21381_ = _20817_ & _21384_ /*7128*/;
assign _21382_ = _20817_ ^ _21384_ /*7131*/;
assign _21383_ = _21375_ & _21382_ /*7129*/;
assign _21380_ = _21381_ | _21383_ /*7127*/;
assign _21203_ = _21375_ ^ _21382_ /*7130*/;
assign _21389_ = D[29] ^ Q[9] /*7126*/;
assign _21386_ = _20818_ & _21389_ /*7122*/;
assign _21387_ = _20818_ ^ _21389_ /*7125*/;
assign _21388_ = _21380_ & _21387_ /*7123*/;
assign _21385_ = _21386_ | _21388_ /*7121*/;
assign _21204_ = _21380_ ^ _21387_ /*7124*/;
assign _21394_ = D[30] ^ Q[9] /*7120*/;
assign _21391_ = _20819_ & _21394_ /*7116*/;
assign _21392_ = _20819_ ^ _21394_ /*7119*/;
assign _21393_ = _21385_ & _21392_ /*7117*/;
assign _21390_ = _21391_ | _21393_ /*7115*/;
assign _21205_ = _21385_ ^ _21392_ /*7118*/;
assign _21399_ = D[31] ^ Q[9] /*7114*/;
assign _21396_ = _20820_ & _21399_ /*7110*/;
assign _21397_ = _20820_ ^ _21399_ /*7113*/;
assign _21398_ = _21390_ & _21397_ /*7111*/;
assign _21395_ = _21396_ | _21398_ /*7109*/;
assign _21206_ = _21390_ ^ _21397_ /*7112*/;
assign _21404_ = D[32] ^ Q[9] /*7108*/;
assign _21401_ = _20821_ & _21404_ /*7104*/;
assign _21402_ = _20821_ ^ _21404_ /*7107*/;
assign _21403_ = _21395_ & _21402_ /*7105*/;
assign _21400_ = _21401_ | _21403_ /*7103*/;
assign _21207_ = _21395_ ^ _21402_ /*7106*/;
assign _21409_ = D[33] ^ Q[9] /*7102*/;
assign _21406_ = _20822_ & _21409_ /*7098*/;
assign _21407_ = _20822_ ^ _21409_ /*7101*/;
assign _21408_ = _21400_ & _21407_ /*7099*/;
assign _21405_ = _21406_ | _21408_ /*7097*/;
assign _21208_ = _21400_ ^ _21407_ /*7100*/;
assign _21414_ = D[34] ^ Q[9] /*7096*/;
assign _21411_ = _20823_ & _21414_ /*7092*/;
assign _21412_ = _20823_ ^ _21414_ /*7095*/;
assign _21413_ = _21405_ & _21412_ /*7093*/;
assign _21410_ = _21411_ | _21413_ /*7091*/;
assign _21209_ = _21405_ ^ _21412_ /*7094*/;
assign _21419_ = D[35] ^ Q[9] /*7090*/;
assign _21416_ = _20824_ & _21419_ /*7086*/;
assign _21417_ = _20824_ ^ _21419_ /*7089*/;
assign _21418_ = _21410_ & _21417_ /*7087*/;
assign _21415_ = _21416_ | _21418_ /*7085*/;
assign _21210_ = _21410_ ^ _21417_ /*7088*/;
assign _21424_ = D[36] ^ Q[9] /*7084*/;
assign _21421_ = _20825_ & _21424_ /*7080*/;
assign _21422_ = _20825_ ^ _21424_ /*7083*/;
assign _21423_ = _21415_ & _21422_ /*7081*/;
assign _21420_ = _21421_ | _21423_ /*7079*/;
assign _21211_ = _21415_ ^ _21422_ /*7082*/;
assign _21429_ = D[37] ^ Q[9] /*7078*/;
assign _21426_ = _20826_ & _21429_ /*7074*/;
assign _21427_ = _20826_ ^ _21429_ /*7077*/;
assign _21428_ = _21420_ & _21427_ /*7075*/;
assign _21425_ = _21426_ | _21428_ /*7073*/;
assign _21212_ = _21420_ ^ _21427_ /*7076*/;
assign _21434_ = D[38] ^ Q[9] /*7072*/;
assign _21431_ = _20827_ & _21434_ /*7068*/;
assign _21432_ = _20827_ ^ _21434_ /*7071*/;
assign _21433_ = _21425_ & _21432_ /*7069*/;
assign _21430_ = _21431_ | _21433_ /*7067*/;
assign _21213_ = _21425_ ^ _21432_ /*7070*/;
assign _21439_ = D[39] ^ Q[9] /*7066*/;
assign _21436_ = _20828_ & _21439_ /*7062*/;
assign _21437_ = _20828_ ^ _21439_ /*7065*/;
assign _21438_ = _21430_ & _21437_ /*7063*/;
assign _21435_ = _21436_ | _21438_ /*7061*/;
assign _21214_ = _21430_ ^ _21437_ /*7064*/;
assign _21444_ = D[40] ^ Q[9] /*7060*/;
assign _21441_ = _20829_ & _21444_ /*7056*/;
assign _21442_ = _20829_ ^ _21444_ /*7059*/;
assign _21443_ = _21435_ & _21442_ /*7057*/;
assign _21440_ = _21441_ | _21443_ /*7055*/;
assign _21215_ = _21435_ ^ _21442_ /*7058*/;
assign _21449_ = D[41] ^ Q[9] /*7054*/;
assign _21446_ = _20830_ & _21449_ /*7050*/;
assign _21447_ = _20830_ ^ _21449_ /*7053*/;
assign _21448_ = _21440_ & _21447_ /*7051*/;
assign _21445_ = _21446_ | _21448_ /*7049*/;
assign _21216_ = _21440_ ^ _21447_ /*7052*/;
assign _21454_ = D[42] ^ Q[9] /*7048*/;
assign _21451_ = _20831_ & _21454_ /*7044*/;
assign _21452_ = _20831_ ^ _21454_ /*7047*/;
assign _21453_ = _21445_ & _21452_ /*7045*/;
assign _21450_ = _21451_ | _21453_ /*7043*/;
assign _21217_ = _21445_ ^ _21452_ /*7046*/;
assign _21459_ = D[43] ^ Q[9] /*7042*/;
assign _21456_ = _20832_ & _21459_ /*7038*/;
assign _21457_ = _20832_ ^ _21459_ /*7041*/;
assign _21458_ = _21450_ & _21457_ /*7039*/;
assign _21455_ = _21456_ | _21458_ /*7037*/;
assign _21218_ = _21450_ ^ _21457_ /*7040*/;
assign _21464_ = D[44] ^ Q[9] /*7036*/;
assign _21461_ = _20833_ & _21464_ /*7032*/;
assign _21462_ = _20833_ ^ _21464_ /*7035*/;
assign _21463_ = _21455_ & _21462_ /*7033*/;
assign _21460_ = _21461_ | _21463_ /*7031*/;
assign _21219_ = _21455_ ^ _21462_ /*7034*/;
assign _21469_ = D[45] ^ Q[9] /*7030*/;
assign _21466_ = _20834_ & _21469_ /*7026*/;
assign _21467_ = _20834_ ^ _21469_ /*7029*/;
assign _21468_ = _21460_ & _21467_ /*7027*/;
assign _21465_ = _21466_ | _21468_ /*7025*/;
assign _21220_ = _21460_ ^ _21467_ /*7028*/;
assign _21474_ = D[46] ^ Q[9] /*7024*/;
assign _21471_ = _20835_ & _21474_ /*7020*/;
assign _21472_ = _20835_ ^ _21474_ /*7023*/;
assign _21473_ = _21465_ & _21472_ /*7021*/;
assign _21470_ = _21471_ | _21473_ /*7019*/;
assign _21221_ = _21465_ ^ _21472_ /*7022*/;
assign _21479_ = D[47] ^ Q[9] /*7018*/;
assign _21476_ = _20836_ & _21479_ /*7014*/;
assign _21477_ = _20836_ ^ _21479_ /*7017*/;
assign _21478_ = _21470_ & _21477_ /*7015*/;
assign _21475_ = _21476_ | _21478_ /*7013*/;
assign _21222_ = _21470_ ^ _21477_ /*7016*/;
assign _21484_ = D[48] ^ Q[9] /*7012*/;
assign _21481_ = _20837_ & _21484_ /*7008*/;
assign _21482_ = _20837_ ^ _21484_ /*7011*/;
assign _21483_ = _21475_ & _21482_ /*7009*/;
assign _21480_ = _21481_ | _21483_ /*7007*/;
assign _21223_ = _21475_ ^ _21482_ /*7010*/;
assign _21489_ = D[49] ^ Q[9] /*7006*/;
assign _21486_ = _20838_ & _21489_ /*7002*/;
assign _21487_ = _20838_ ^ _21489_ /*7005*/;
assign _21488_ = _21480_ & _21487_ /*7003*/;
assign _21485_ = _21486_ | _21488_ /*7001*/;
assign _21224_ = _21480_ ^ _21487_ /*7004*/;
assign _21494_ = D[50] ^ Q[9] /*7000*/;
assign _21491_ = _20839_ & _21494_ /*6996*/;
assign _21492_ = _20839_ ^ _21494_ /*6999*/;
assign _21493_ = _21485_ & _21492_ /*6997*/;
assign _21490_ = _21491_ | _21493_ /*6995*/;
assign _21225_ = _21485_ ^ _21492_ /*6998*/;
assign _21499_ = D[51] ^ Q[9] /*6994*/;
assign _21496_ = _20840_ & _21499_ /*6990*/;
assign _21497_ = _20840_ ^ _21499_ /*6993*/;
assign _21498_ = _21490_ & _21497_ /*6991*/;
assign _21495_ = _21496_ | _21498_ /*6989*/;
assign _21226_ = _21490_ ^ _21497_ /*6992*/;
assign _21504_ = D[52] ^ Q[9] /*6988*/;
assign _21501_ = _20841_ & _21504_ /*6984*/;
assign _21502_ = _20841_ ^ _21504_ /*6987*/;
assign _21503_ = _21495_ & _21502_ /*6985*/;
assign _21500_ = _21501_ | _21503_ /*6983*/;
assign _21227_ = _21495_ ^ _21502_ /*6986*/;
assign _21509_ = D[53] ^ Q[9] /*6982*/;
assign _21506_ = _20842_ & _21509_ /*6978*/;
assign _21507_ = _20842_ ^ _21509_ /*6981*/;
assign _21508_ = _21500_ & _21507_ /*6979*/;
assign _21505_ = _21506_ | _21508_ /*6977*/;
assign _21228_ = _21500_ ^ _21507_ /*6980*/;
assign _21514_ = D[54] ^ Q[9] /*6976*/;
assign _21511_ = _20843_ & _21514_ /*6972*/;
assign _21512_ = _20843_ ^ _21514_ /*6975*/;
assign _21513_ = _21505_ & _21512_ /*6973*/;
assign _21510_ = _21511_ | _21513_ /*6971*/;
assign _21229_ = _21505_ ^ _21512_ /*6974*/;
assign _21519_ = D[55] ^ Q[9] /*6970*/;
assign _21516_ = _20844_ & _21519_ /*6966*/;
assign _21517_ = _20844_ ^ _21519_ /*6969*/;
assign _21518_ = _21510_ & _21517_ /*6967*/;
assign _21515_ = _21516_ | _21518_ /*6965*/;
assign _21230_ = _21510_ ^ _21517_ /*6968*/;
assign _21524_ = D[56] ^ Q[9] /*6964*/;
assign _21521_ = _20845_ & _21524_ /*6960*/;
assign _21522_ = _20845_ ^ _21524_ /*6963*/;
assign _21523_ = _21515_ & _21522_ /*6961*/;
assign _21520_ = _21521_ | _21523_ /*6959*/;
assign _21231_ = _21515_ ^ _21522_ /*6962*/;
assign _21529_ = D[57] ^ Q[9] /*6958*/;
assign _21526_ = _20846_ & _21529_ /*6954*/;
assign _21527_ = _20846_ ^ _21529_ /*6957*/;
assign _21528_ = _21520_ & _21527_ /*6955*/;
assign _21525_ = _21526_ | _21528_ /*6953*/;
assign _21232_ = _21520_ ^ _21527_ /*6956*/;
assign _21534_ = D[58] ^ Q[9] /*6952*/;
assign _21531_ = _20847_ & _21534_ /*6948*/;
assign _21532_ = _20847_ ^ _21534_ /*6951*/;
assign _21533_ = _21525_ & _21532_ /*6949*/;
assign _21530_ = _21531_ | _21533_ /*6947*/;
assign _21233_ = _21525_ ^ _21532_ /*6950*/;
assign _21539_ = D[59] ^ Q[9] /*6946*/;
assign _21536_ = _20848_ & _21539_ /*6942*/;
assign _21537_ = _20848_ ^ _21539_ /*6945*/;
assign _21538_ = _21530_ & _21537_ /*6943*/;
assign _21535_ = _21536_ | _21538_ /*6941*/;
assign _21234_ = _21530_ ^ _21537_ /*6944*/;
assign _21544_ = D[60] ^ Q[9] /*6940*/;
assign _21541_ = _20849_ & _21544_ /*6936*/;
assign _21542_ = _20849_ ^ _21544_ /*6939*/;
assign _21543_ = _21535_ & _21542_ /*6937*/;
assign _21540_ = _21541_ | _21543_ /*6935*/;
assign _21235_ = _21535_ ^ _21542_ /*6938*/;
assign _21549_ = D[61] ^ Q[9] /*6934*/;
assign _21546_ = _20850_ & _21549_ /*6930*/;
assign _21547_ = _20850_ ^ _21549_ /*6933*/;
assign _21548_ = _21540_ & _21547_ /*6931*/;
assign _21545_ = _21546_ | _21548_ /*6929*/;
assign _21236_ = _21540_ ^ _21547_ /*6932*/;
assign _21554_ = D[62] ^ Q[9] /*6928*/;
assign _21551_ = _20851_ & _21554_ /*6924*/;
assign _21552_ = _20851_ ^ _21554_ /*6927*/;
assign _21553_ = _21545_ & _21552_ /*6925*/;
assign _21550_ = _21551_ | _21553_ /*6923*/;
assign _21237_ = _21545_ ^ _21552_ /*6926*/;
assign _21558_ = zeroWire ^ Q[9] /*6922*/;
assign _21555_ = _20852_ & _21558_ /*6918*/;
assign _21556_ = _20852_ ^ _21558_ /*6921*/;
assign _21557_ = _21550_ & _21556_ /*6919*/;
assign Q[8] = _21555_ | _21557_ /*6917*/;
assign _21238_ = _21550_ ^ _21556_ /*6920*/;
assign _21629_ = D[0] ^ Q[8] /*6531*/;
assign _21626_ = R_0[7] & _21629_ /*6527*/;
assign _21627_ = R_0[7] ^ _21629_ /*6530*/;
assign _21628_ = Q[8] & _21627_ /*6528*/;
assign _21625_ = _21626_ | _21628_ /*6526*/;
assign _21560_ = Q[8] ^ _21627_ /*6529*/;
assign _21634_ = D[1] ^ Q[8] /*6525*/;
assign _21631_ = _21175_ & _21634_ /*6521*/;
assign _21632_ = _21175_ ^ _21634_ /*6524*/;
assign _21633_ = _21625_ & _21632_ /*6522*/;
assign _21630_ = _21631_ | _21633_ /*6520*/;
assign _21561_ = _21625_ ^ _21632_ /*6523*/;
assign _21639_ = D[2] ^ Q[8] /*6519*/;
assign _21636_ = _21176_ & _21639_ /*6515*/;
assign _21637_ = _21176_ ^ _21639_ /*6518*/;
assign _21638_ = _21630_ & _21637_ /*6516*/;
assign _21635_ = _21636_ | _21638_ /*6514*/;
assign _21562_ = _21630_ ^ _21637_ /*6517*/;
assign _21644_ = D[3] ^ Q[8] /*6513*/;
assign _21641_ = _21177_ & _21644_ /*6509*/;
assign _21642_ = _21177_ ^ _21644_ /*6512*/;
assign _21643_ = _21635_ & _21642_ /*6510*/;
assign _21640_ = _21641_ | _21643_ /*6508*/;
assign _21563_ = _21635_ ^ _21642_ /*6511*/;
assign _21649_ = D[4] ^ Q[8] /*6507*/;
assign _21646_ = _21178_ & _21649_ /*6503*/;
assign _21647_ = _21178_ ^ _21649_ /*6506*/;
assign _21648_ = _21640_ & _21647_ /*6504*/;
assign _21645_ = _21646_ | _21648_ /*6502*/;
assign _21564_ = _21640_ ^ _21647_ /*6505*/;
assign _21654_ = D[5] ^ Q[8] /*6501*/;
assign _21651_ = _21179_ & _21654_ /*6497*/;
assign _21652_ = _21179_ ^ _21654_ /*6500*/;
assign _21653_ = _21645_ & _21652_ /*6498*/;
assign _21650_ = _21651_ | _21653_ /*6496*/;
assign _21565_ = _21645_ ^ _21652_ /*6499*/;
assign _21659_ = D[6] ^ Q[8] /*6495*/;
assign _21656_ = _21180_ & _21659_ /*6491*/;
assign _21657_ = _21180_ ^ _21659_ /*6494*/;
assign _21658_ = _21650_ & _21657_ /*6492*/;
assign _21655_ = _21656_ | _21658_ /*6490*/;
assign _21566_ = _21650_ ^ _21657_ /*6493*/;
assign _21664_ = D[7] ^ Q[8] /*6489*/;
assign _21661_ = _21181_ & _21664_ /*6485*/;
assign _21662_ = _21181_ ^ _21664_ /*6488*/;
assign _21663_ = _21655_ & _21662_ /*6486*/;
assign _21660_ = _21661_ | _21663_ /*6484*/;
assign _21567_ = _21655_ ^ _21662_ /*6487*/;
assign _21669_ = D[8] ^ Q[8] /*6483*/;
assign _21666_ = _21182_ & _21669_ /*6479*/;
assign _21667_ = _21182_ ^ _21669_ /*6482*/;
assign _21668_ = _21660_ & _21667_ /*6480*/;
assign _21665_ = _21666_ | _21668_ /*6478*/;
assign _21568_ = _21660_ ^ _21667_ /*6481*/;
assign _21674_ = D[9] ^ Q[8] /*6477*/;
assign _21671_ = _21183_ & _21674_ /*6473*/;
assign _21672_ = _21183_ ^ _21674_ /*6476*/;
assign _21673_ = _21665_ & _21672_ /*6474*/;
assign _21670_ = _21671_ | _21673_ /*6472*/;
assign _21569_ = _21665_ ^ _21672_ /*6475*/;
assign _21679_ = D[10] ^ Q[8] /*6471*/;
assign _21676_ = _21184_ & _21679_ /*6467*/;
assign _21677_ = _21184_ ^ _21679_ /*6470*/;
assign _21678_ = _21670_ & _21677_ /*6468*/;
assign _21675_ = _21676_ | _21678_ /*6466*/;
assign _21570_ = _21670_ ^ _21677_ /*6469*/;
assign _21684_ = D[11] ^ Q[8] /*6465*/;
assign _21681_ = _21185_ & _21684_ /*6461*/;
assign _21682_ = _21185_ ^ _21684_ /*6464*/;
assign _21683_ = _21675_ & _21682_ /*6462*/;
assign _21680_ = _21681_ | _21683_ /*6460*/;
assign _21571_ = _21675_ ^ _21682_ /*6463*/;
assign _21689_ = D[12] ^ Q[8] /*6459*/;
assign _21686_ = _21186_ & _21689_ /*6455*/;
assign _21687_ = _21186_ ^ _21689_ /*6458*/;
assign _21688_ = _21680_ & _21687_ /*6456*/;
assign _21685_ = _21686_ | _21688_ /*6454*/;
assign _21572_ = _21680_ ^ _21687_ /*6457*/;
assign _21694_ = D[13] ^ Q[8] /*6453*/;
assign _21691_ = _21187_ & _21694_ /*6449*/;
assign _21692_ = _21187_ ^ _21694_ /*6452*/;
assign _21693_ = _21685_ & _21692_ /*6450*/;
assign _21690_ = _21691_ | _21693_ /*6448*/;
assign _21573_ = _21685_ ^ _21692_ /*6451*/;
assign _21699_ = D[14] ^ Q[8] /*6447*/;
assign _21696_ = _21188_ & _21699_ /*6443*/;
assign _21697_ = _21188_ ^ _21699_ /*6446*/;
assign _21698_ = _21690_ & _21697_ /*6444*/;
assign _21695_ = _21696_ | _21698_ /*6442*/;
assign _21574_ = _21690_ ^ _21697_ /*6445*/;
assign _21704_ = D[15] ^ Q[8] /*6441*/;
assign _21701_ = _21189_ & _21704_ /*6437*/;
assign _21702_ = _21189_ ^ _21704_ /*6440*/;
assign _21703_ = _21695_ & _21702_ /*6438*/;
assign _21700_ = _21701_ | _21703_ /*6436*/;
assign _21575_ = _21695_ ^ _21702_ /*6439*/;
assign _21709_ = D[16] ^ Q[8] /*6435*/;
assign _21706_ = _21190_ & _21709_ /*6431*/;
assign _21707_ = _21190_ ^ _21709_ /*6434*/;
assign _21708_ = _21700_ & _21707_ /*6432*/;
assign _21705_ = _21706_ | _21708_ /*6430*/;
assign _21576_ = _21700_ ^ _21707_ /*6433*/;
assign _21714_ = D[17] ^ Q[8] /*6429*/;
assign _21711_ = _21191_ & _21714_ /*6425*/;
assign _21712_ = _21191_ ^ _21714_ /*6428*/;
assign _21713_ = _21705_ & _21712_ /*6426*/;
assign _21710_ = _21711_ | _21713_ /*6424*/;
assign _21577_ = _21705_ ^ _21712_ /*6427*/;
assign _21719_ = D[18] ^ Q[8] /*6423*/;
assign _21716_ = _21192_ & _21719_ /*6419*/;
assign _21717_ = _21192_ ^ _21719_ /*6422*/;
assign _21718_ = _21710_ & _21717_ /*6420*/;
assign _21715_ = _21716_ | _21718_ /*6418*/;
assign _21578_ = _21710_ ^ _21717_ /*6421*/;
assign _21724_ = D[19] ^ Q[8] /*6417*/;
assign _21721_ = _21193_ & _21724_ /*6413*/;
assign _21722_ = _21193_ ^ _21724_ /*6416*/;
assign _21723_ = _21715_ & _21722_ /*6414*/;
assign _21720_ = _21721_ | _21723_ /*6412*/;
assign _21579_ = _21715_ ^ _21722_ /*6415*/;
assign _21729_ = D[20] ^ Q[8] /*6411*/;
assign _21726_ = _21194_ & _21729_ /*6407*/;
assign _21727_ = _21194_ ^ _21729_ /*6410*/;
assign _21728_ = _21720_ & _21727_ /*6408*/;
assign _21725_ = _21726_ | _21728_ /*6406*/;
assign _21580_ = _21720_ ^ _21727_ /*6409*/;
assign _21734_ = D[21] ^ Q[8] /*6405*/;
assign _21731_ = _21195_ & _21734_ /*6401*/;
assign _21732_ = _21195_ ^ _21734_ /*6404*/;
assign _21733_ = _21725_ & _21732_ /*6402*/;
assign _21730_ = _21731_ | _21733_ /*6400*/;
assign _21581_ = _21725_ ^ _21732_ /*6403*/;
assign _21739_ = D[22] ^ Q[8] /*6399*/;
assign _21736_ = _21196_ & _21739_ /*6395*/;
assign _21737_ = _21196_ ^ _21739_ /*6398*/;
assign _21738_ = _21730_ & _21737_ /*6396*/;
assign _21735_ = _21736_ | _21738_ /*6394*/;
assign _21582_ = _21730_ ^ _21737_ /*6397*/;
assign _21744_ = D[23] ^ Q[8] /*6393*/;
assign _21741_ = _21197_ & _21744_ /*6389*/;
assign _21742_ = _21197_ ^ _21744_ /*6392*/;
assign _21743_ = _21735_ & _21742_ /*6390*/;
assign _21740_ = _21741_ | _21743_ /*6388*/;
assign _21583_ = _21735_ ^ _21742_ /*6391*/;
assign _21749_ = D[24] ^ Q[8] /*6387*/;
assign _21746_ = _21198_ & _21749_ /*6383*/;
assign _21747_ = _21198_ ^ _21749_ /*6386*/;
assign _21748_ = _21740_ & _21747_ /*6384*/;
assign _21745_ = _21746_ | _21748_ /*6382*/;
assign _21584_ = _21740_ ^ _21747_ /*6385*/;
assign _21754_ = D[25] ^ Q[8] /*6381*/;
assign _21751_ = _21199_ & _21754_ /*6377*/;
assign _21752_ = _21199_ ^ _21754_ /*6380*/;
assign _21753_ = _21745_ & _21752_ /*6378*/;
assign _21750_ = _21751_ | _21753_ /*6376*/;
assign _21585_ = _21745_ ^ _21752_ /*6379*/;
assign _21759_ = D[26] ^ Q[8] /*6375*/;
assign _21756_ = _21200_ & _21759_ /*6371*/;
assign _21757_ = _21200_ ^ _21759_ /*6374*/;
assign _21758_ = _21750_ & _21757_ /*6372*/;
assign _21755_ = _21756_ | _21758_ /*6370*/;
assign _21586_ = _21750_ ^ _21757_ /*6373*/;
assign _21764_ = D[27] ^ Q[8] /*6369*/;
assign _21761_ = _21201_ & _21764_ /*6365*/;
assign _21762_ = _21201_ ^ _21764_ /*6368*/;
assign _21763_ = _21755_ & _21762_ /*6366*/;
assign _21760_ = _21761_ | _21763_ /*6364*/;
assign _21587_ = _21755_ ^ _21762_ /*6367*/;
assign _21769_ = D[28] ^ Q[8] /*6363*/;
assign _21766_ = _21202_ & _21769_ /*6359*/;
assign _21767_ = _21202_ ^ _21769_ /*6362*/;
assign _21768_ = _21760_ & _21767_ /*6360*/;
assign _21765_ = _21766_ | _21768_ /*6358*/;
assign _21588_ = _21760_ ^ _21767_ /*6361*/;
assign _21774_ = D[29] ^ Q[8] /*6357*/;
assign _21771_ = _21203_ & _21774_ /*6353*/;
assign _21772_ = _21203_ ^ _21774_ /*6356*/;
assign _21773_ = _21765_ & _21772_ /*6354*/;
assign _21770_ = _21771_ | _21773_ /*6352*/;
assign _21589_ = _21765_ ^ _21772_ /*6355*/;
assign _21779_ = D[30] ^ Q[8] /*6351*/;
assign _21776_ = _21204_ & _21779_ /*6347*/;
assign _21777_ = _21204_ ^ _21779_ /*6350*/;
assign _21778_ = _21770_ & _21777_ /*6348*/;
assign _21775_ = _21776_ | _21778_ /*6346*/;
assign _21590_ = _21770_ ^ _21777_ /*6349*/;
assign _21784_ = D[31] ^ Q[8] /*6345*/;
assign _21781_ = _21205_ & _21784_ /*6341*/;
assign _21782_ = _21205_ ^ _21784_ /*6344*/;
assign _21783_ = _21775_ & _21782_ /*6342*/;
assign _21780_ = _21781_ | _21783_ /*6340*/;
assign _21591_ = _21775_ ^ _21782_ /*6343*/;
assign _21789_ = D[32] ^ Q[8] /*6339*/;
assign _21786_ = _21206_ & _21789_ /*6335*/;
assign _21787_ = _21206_ ^ _21789_ /*6338*/;
assign _21788_ = _21780_ & _21787_ /*6336*/;
assign _21785_ = _21786_ | _21788_ /*6334*/;
assign _21592_ = _21780_ ^ _21787_ /*6337*/;
assign _21794_ = D[33] ^ Q[8] /*6333*/;
assign _21791_ = _21207_ & _21794_ /*6329*/;
assign _21792_ = _21207_ ^ _21794_ /*6332*/;
assign _21793_ = _21785_ & _21792_ /*6330*/;
assign _21790_ = _21791_ | _21793_ /*6328*/;
assign _21593_ = _21785_ ^ _21792_ /*6331*/;
assign _21799_ = D[34] ^ Q[8] /*6327*/;
assign _21796_ = _21208_ & _21799_ /*6323*/;
assign _21797_ = _21208_ ^ _21799_ /*6326*/;
assign _21798_ = _21790_ & _21797_ /*6324*/;
assign _21795_ = _21796_ | _21798_ /*6322*/;
assign _21594_ = _21790_ ^ _21797_ /*6325*/;
assign _21804_ = D[35] ^ Q[8] /*6321*/;
assign _21801_ = _21209_ & _21804_ /*6317*/;
assign _21802_ = _21209_ ^ _21804_ /*6320*/;
assign _21803_ = _21795_ & _21802_ /*6318*/;
assign _21800_ = _21801_ | _21803_ /*6316*/;
assign _21595_ = _21795_ ^ _21802_ /*6319*/;
assign _21809_ = D[36] ^ Q[8] /*6315*/;
assign _21806_ = _21210_ & _21809_ /*6311*/;
assign _21807_ = _21210_ ^ _21809_ /*6314*/;
assign _21808_ = _21800_ & _21807_ /*6312*/;
assign _21805_ = _21806_ | _21808_ /*6310*/;
assign _21596_ = _21800_ ^ _21807_ /*6313*/;
assign _21814_ = D[37] ^ Q[8] /*6309*/;
assign _21811_ = _21211_ & _21814_ /*6305*/;
assign _21812_ = _21211_ ^ _21814_ /*6308*/;
assign _21813_ = _21805_ & _21812_ /*6306*/;
assign _21810_ = _21811_ | _21813_ /*6304*/;
assign _21597_ = _21805_ ^ _21812_ /*6307*/;
assign _21819_ = D[38] ^ Q[8] /*6303*/;
assign _21816_ = _21212_ & _21819_ /*6299*/;
assign _21817_ = _21212_ ^ _21819_ /*6302*/;
assign _21818_ = _21810_ & _21817_ /*6300*/;
assign _21815_ = _21816_ | _21818_ /*6298*/;
assign _21598_ = _21810_ ^ _21817_ /*6301*/;
assign _21824_ = D[39] ^ Q[8] /*6297*/;
assign _21821_ = _21213_ & _21824_ /*6293*/;
assign _21822_ = _21213_ ^ _21824_ /*6296*/;
assign _21823_ = _21815_ & _21822_ /*6294*/;
assign _21820_ = _21821_ | _21823_ /*6292*/;
assign _21599_ = _21815_ ^ _21822_ /*6295*/;
assign _21829_ = D[40] ^ Q[8] /*6291*/;
assign _21826_ = _21214_ & _21829_ /*6287*/;
assign _21827_ = _21214_ ^ _21829_ /*6290*/;
assign _21828_ = _21820_ & _21827_ /*6288*/;
assign _21825_ = _21826_ | _21828_ /*6286*/;
assign _21600_ = _21820_ ^ _21827_ /*6289*/;
assign _21834_ = D[41] ^ Q[8] /*6285*/;
assign _21831_ = _21215_ & _21834_ /*6281*/;
assign _21832_ = _21215_ ^ _21834_ /*6284*/;
assign _21833_ = _21825_ & _21832_ /*6282*/;
assign _21830_ = _21831_ | _21833_ /*6280*/;
assign _21601_ = _21825_ ^ _21832_ /*6283*/;
assign _21839_ = D[42] ^ Q[8] /*6279*/;
assign _21836_ = _21216_ & _21839_ /*6275*/;
assign _21837_ = _21216_ ^ _21839_ /*6278*/;
assign _21838_ = _21830_ & _21837_ /*6276*/;
assign _21835_ = _21836_ | _21838_ /*6274*/;
assign _21602_ = _21830_ ^ _21837_ /*6277*/;
assign _21844_ = D[43] ^ Q[8] /*6273*/;
assign _21841_ = _21217_ & _21844_ /*6269*/;
assign _21842_ = _21217_ ^ _21844_ /*6272*/;
assign _21843_ = _21835_ & _21842_ /*6270*/;
assign _21840_ = _21841_ | _21843_ /*6268*/;
assign _21603_ = _21835_ ^ _21842_ /*6271*/;
assign _21849_ = D[44] ^ Q[8] /*6267*/;
assign _21846_ = _21218_ & _21849_ /*6263*/;
assign _21847_ = _21218_ ^ _21849_ /*6266*/;
assign _21848_ = _21840_ & _21847_ /*6264*/;
assign _21845_ = _21846_ | _21848_ /*6262*/;
assign _21604_ = _21840_ ^ _21847_ /*6265*/;
assign _21854_ = D[45] ^ Q[8] /*6261*/;
assign _21851_ = _21219_ & _21854_ /*6257*/;
assign _21852_ = _21219_ ^ _21854_ /*6260*/;
assign _21853_ = _21845_ & _21852_ /*6258*/;
assign _21850_ = _21851_ | _21853_ /*6256*/;
assign _21605_ = _21845_ ^ _21852_ /*6259*/;
assign _21859_ = D[46] ^ Q[8] /*6255*/;
assign _21856_ = _21220_ & _21859_ /*6251*/;
assign _21857_ = _21220_ ^ _21859_ /*6254*/;
assign _21858_ = _21850_ & _21857_ /*6252*/;
assign _21855_ = _21856_ | _21858_ /*6250*/;
assign _21606_ = _21850_ ^ _21857_ /*6253*/;
assign _21864_ = D[47] ^ Q[8] /*6249*/;
assign _21861_ = _21221_ & _21864_ /*6245*/;
assign _21862_ = _21221_ ^ _21864_ /*6248*/;
assign _21863_ = _21855_ & _21862_ /*6246*/;
assign _21860_ = _21861_ | _21863_ /*6244*/;
assign _21607_ = _21855_ ^ _21862_ /*6247*/;
assign _21869_ = D[48] ^ Q[8] /*6243*/;
assign _21866_ = _21222_ & _21869_ /*6239*/;
assign _21867_ = _21222_ ^ _21869_ /*6242*/;
assign _21868_ = _21860_ & _21867_ /*6240*/;
assign _21865_ = _21866_ | _21868_ /*6238*/;
assign _21608_ = _21860_ ^ _21867_ /*6241*/;
assign _21874_ = D[49] ^ Q[8] /*6237*/;
assign _21871_ = _21223_ & _21874_ /*6233*/;
assign _21872_ = _21223_ ^ _21874_ /*6236*/;
assign _21873_ = _21865_ & _21872_ /*6234*/;
assign _21870_ = _21871_ | _21873_ /*6232*/;
assign _21609_ = _21865_ ^ _21872_ /*6235*/;
assign _21879_ = D[50] ^ Q[8] /*6231*/;
assign _21876_ = _21224_ & _21879_ /*6227*/;
assign _21877_ = _21224_ ^ _21879_ /*6230*/;
assign _21878_ = _21870_ & _21877_ /*6228*/;
assign _21875_ = _21876_ | _21878_ /*6226*/;
assign _21610_ = _21870_ ^ _21877_ /*6229*/;
assign _21884_ = D[51] ^ Q[8] /*6225*/;
assign _21881_ = _21225_ & _21884_ /*6221*/;
assign _21882_ = _21225_ ^ _21884_ /*6224*/;
assign _21883_ = _21875_ & _21882_ /*6222*/;
assign _21880_ = _21881_ | _21883_ /*6220*/;
assign _21611_ = _21875_ ^ _21882_ /*6223*/;
assign _21889_ = D[52] ^ Q[8] /*6219*/;
assign _21886_ = _21226_ & _21889_ /*6215*/;
assign _21887_ = _21226_ ^ _21889_ /*6218*/;
assign _21888_ = _21880_ & _21887_ /*6216*/;
assign _21885_ = _21886_ | _21888_ /*6214*/;
assign _21612_ = _21880_ ^ _21887_ /*6217*/;
assign _21894_ = D[53] ^ Q[8] /*6213*/;
assign _21891_ = _21227_ & _21894_ /*6209*/;
assign _21892_ = _21227_ ^ _21894_ /*6212*/;
assign _21893_ = _21885_ & _21892_ /*6210*/;
assign _21890_ = _21891_ | _21893_ /*6208*/;
assign _21613_ = _21885_ ^ _21892_ /*6211*/;
assign _21899_ = D[54] ^ Q[8] /*6207*/;
assign _21896_ = _21228_ & _21899_ /*6203*/;
assign _21897_ = _21228_ ^ _21899_ /*6206*/;
assign _21898_ = _21890_ & _21897_ /*6204*/;
assign _21895_ = _21896_ | _21898_ /*6202*/;
assign _21614_ = _21890_ ^ _21897_ /*6205*/;
assign _21904_ = D[55] ^ Q[8] /*6201*/;
assign _21901_ = _21229_ & _21904_ /*6197*/;
assign _21902_ = _21229_ ^ _21904_ /*6200*/;
assign _21903_ = _21895_ & _21902_ /*6198*/;
assign _21900_ = _21901_ | _21903_ /*6196*/;
assign _21615_ = _21895_ ^ _21902_ /*6199*/;
assign _21909_ = D[56] ^ Q[8] /*6195*/;
assign _21906_ = _21230_ & _21909_ /*6191*/;
assign _21907_ = _21230_ ^ _21909_ /*6194*/;
assign _21908_ = _21900_ & _21907_ /*6192*/;
assign _21905_ = _21906_ | _21908_ /*6190*/;
assign _21616_ = _21900_ ^ _21907_ /*6193*/;
assign _21914_ = D[57] ^ Q[8] /*6189*/;
assign _21911_ = _21231_ & _21914_ /*6185*/;
assign _21912_ = _21231_ ^ _21914_ /*6188*/;
assign _21913_ = _21905_ & _21912_ /*6186*/;
assign _21910_ = _21911_ | _21913_ /*6184*/;
assign _21617_ = _21905_ ^ _21912_ /*6187*/;
assign _21919_ = D[58] ^ Q[8] /*6183*/;
assign _21916_ = _21232_ & _21919_ /*6179*/;
assign _21917_ = _21232_ ^ _21919_ /*6182*/;
assign _21918_ = _21910_ & _21917_ /*6180*/;
assign _21915_ = _21916_ | _21918_ /*6178*/;
assign _21618_ = _21910_ ^ _21917_ /*6181*/;
assign _21924_ = D[59] ^ Q[8] /*6177*/;
assign _21921_ = _21233_ & _21924_ /*6173*/;
assign _21922_ = _21233_ ^ _21924_ /*6176*/;
assign _21923_ = _21915_ & _21922_ /*6174*/;
assign _21920_ = _21921_ | _21923_ /*6172*/;
assign _21619_ = _21915_ ^ _21922_ /*6175*/;
assign _21929_ = D[60] ^ Q[8] /*6171*/;
assign _21926_ = _21234_ & _21929_ /*6167*/;
assign _21927_ = _21234_ ^ _21929_ /*6170*/;
assign _21928_ = _21920_ & _21927_ /*6168*/;
assign _21925_ = _21926_ | _21928_ /*6166*/;
assign _21620_ = _21920_ ^ _21927_ /*6169*/;
assign _21934_ = D[61] ^ Q[8] /*6165*/;
assign _21931_ = _21235_ & _21934_ /*6161*/;
assign _21932_ = _21235_ ^ _21934_ /*6164*/;
assign _21933_ = _21925_ & _21932_ /*6162*/;
assign _21930_ = _21931_ | _21933_ /*6160*/;
assign _21621_ = _21925_ ^ _21932_ /*6163*/;
assign _21939_ = D[62] ^ Q[8] /*6159*/;
assign _21936_ = _21236_ & _21939_ /*6155*/;
assign _21937_ = _21236_ ^ _21939_ /*6158*/;
assign _21938_ = _21930_ & _21937_ /*6156*/;
assign _21935_ = _21936_ | _21938_ /*6154*/;
assign _21622_ = _21930_ ^ _21937_ /*6157*/;
assign _21943_ = zeroWire ^ Q[8] /*6153*/;
assign _21940_ = _21237_ & _21943_ /*6149*/;
assign _21941_ = _21237_ ^ _21943_ /*6152*/;
assign _21942_ = _21935_ & _21941_ /*6150*/;
assign Q[7] = _21940_ | _21942_ /*6148*/;
assign _21623_ = _21935_ ^ _21941_ /*6151*/;
assign _22014_ = D[0] ^ Q[7] /*5762*/;
assign _22011_ = R_0[6] & _22014_ /*5758*/;
assign _22012_ = R_0[6] ^ _22014_ /*5761*/;
assign _22013_ = Q[7] & _22012_ /*5759*/;
assign _22010_ = _22011_ | _22013_ /*5757*/;
assign _21945_ = Q[7] ^ _22012_ /*5760*/;
assign _22019_ = D[1] ^ Q[7] /*5756*/;
assign _22016_ = _21560_ & _22019_ /*5752*/;
assign _22017_ = _21560_ ^ _22019_ /*5755*/;
assign _22018_ = _22010_ & _22017_ /*5753*/;
assign _22015_ = _22016_ | _22018_ /*5751*/;
assign _21946_ = _22010_ ^ _22017_ /*5754*/;
assign _22024_ = D[2] ^ Q[7] /*5750*/;
assign _22021_ = _21561_ & _22024_ /*5746*/;
assign _22022_ = _21561_ ^ _22024_ /*5749*/;
assign _22023_ = _22015_ & _22022_ /*5747*/;
assign _22020_ = _22021_ | _22023_ /*5745*/;
assign _21947_ = _22015_ ^ _22022_ /*5748*/;
assign _22029_ = D[3] ^ Q[7] /*5744*/;
assign _22026_ = _21562_ & _22029_ /*5740*/;
assign _22027_ = _21562_ ^ _22029_ /*5743*/;
assign _22028_ = _22020_ & _22027_ /*5741*/;
assign _22025_ = _22026_ | _22028_ /*5739*/;
assign _21948_ = _22020_ ^ _22027_ /*5742*/;
assign _22034_ = D[4] ^ Q[7] /*5738*/;
assign _22031_ = _21563_ & _22034_ /*5734*/;
assign _22032_ = _21563_ ^ _22034_ /*5737*/;
assign _22033_ = _22025_ & _22032_ /*5735*/;
assign _22030_ = _22031_ | _22033_ /*5733*/;
assign _21949_ = _22025_ ^ _22032_ /*5736*/;
assign _22039_ = D[5] ^ Q[7] /*5732*/;
assign _22036_ = _21564_ & _22039_ /*5728*/;
assign _22037_ = _21564_ ^ _22039_ /*5731*/;
assign _22038_ = _22030_ & _22037_ /*5729*/;
assign _22035_ = _22036_ | _22038_ /*5727*/;
assign _21950_ = _22030_ ^ _22037_ /*5730*/;
assign _22044_ = D[6] ^ Q[7] /*5726*/;
assign _22041_ = _21565_ & _22044_ /*5722*/;
assign _22042_ = _21565_ ^ _22044_ /*5725*/;
assign _22043_ = _22035_ & _22042_ /*5723*/;
assign _22040_ = _22041_ | _22043_ /*5721*/;
assign _21951_ = _22035_ ^ _22042_ /*5724*/;
assign _22049_ = D[7] ^ Q[7] /*5720*/;
assign _22046_ = _21566_ & _22049_ /*5716*/;
assign _22047_ = _21566_ ^ _22049_ /*5719*/;
assign _22048_ = _22040_ & _22047_ /*5717*/;
assign _22045_ = _22046_ | _22048_ /*5715*/;
assign _21952_ = _22040_ ^ _22047_ /*5718*/;
assign _22054_ = D[8] ^ Q[7] /*5714*/;
assign _22051_ = _21567_ & _22054_ /*5710*/;
assign _22052_ = _21567_ ^ _22054_ /*5713*/;
assign _22053_ = _22045_ & _22052_ /*5711*/;
assign _22050_ = _22051_ | _22053_ /*5709*/;
assign _21953_ = _22045_ ^ _22052_ /*5712*/;
assign _22059_ = D[9] ^ Q[7] /*5708*/;
assign _22056_ = _21568_ & _22059_ /*5704*/;
assign _22057_ = _21568_ ^ _22059_ /*5707*/;
assign _22058_ = _22050_ & _22057_ /*5705*/;
assign _22055_ = _22056_ | _22058_ /*5703*/;
assign _21954_ = _22050_ ^ _22057_ /*5706*/;
assign _22064_ = D[10] ^ Q[7] /*5702*/;
assign _22061_ = _21569_ & _22064_ /*5698*/;
assign _22062_ = _21569_ ^ _22064_ /*5701*/;
assign _22063_ = _22055_ & _22062_ /*5699*/;
assign _22060_ = _22061_ | _22063_ /*5697*/;
assign _21955_ = _22055_ ^ _22062_ /*5700*/;
assign _22069_ = D[11] ^ Q[7] /*5696*/;
assign _22066_ = _21570_ & _22069_ /*5692*/;
assign _22067_ = _21570_ ^ _22069_ /*5695*/;
assign _22068_ = _22060_ & _22067_ /*5693*/;
assign _22065_ = _22066_ | _22068_ /*5691*/;
assign _21956_ = _22060_ ^ _22067_ /*5694*/;
assign _22074_ = D[12] ^ Q[7] /*5690*/;
assign _22071_ = _21571_ & _22074_ /*5686*/;
assign _22072_ = _21571_ ^ _22074_ /*5689*/;
assign _22073_ = _22065_ & _22072_ /*5687*/;
assign _22070_ = _22071_ | _22073_ /*5685*/;
assign _21957_ = _22065_ ^ _22072_ /*5688*/;
assign _22079_ = D[13] ^ Q[7] /*5684*/;
assign _22076_ = _21572_ & _22079_ /*5680*/;
assign _22077_ = _21572_ ^ _22079_ /*5683*/;
assign _22078_ = _22070_ & _22077_ /*5681*/;
assign _22075_ = _22076_ | _22078_ /*5679*/;
assign _21958_ = _22070_ ^ _22077_ /*5682*/;
assign _22084_ = D[14] ^ Q[7] /*5678*/;
assign _22081_ = _21573_ & _22084_ /*5674*/;
assign _22082_ = _21573_ ^ _22084_ /*5677*/;
assign _22083_ = _22075_ & _22082_ /*5675*/;
assign _22080_ = _22081_ | _22083_ /*5673*/;
assign _21959_ = _22075_ ^ _22082_ /*5676*/;
assign _22089_ = D[15] ^ Q[7] /*5672*/;
assign _22086_ = _21574_ & _22089_ /*5668*/;
assign _22087_ = _21574_ ^ _22089_ /*5671*/;
assign _22088_ = _22080_ & _22087_ /*5669*/;
assign _22085_ = _22086_ | _22088_ /*5667*/;
assign _21960_ = _22080_ ^ _22087_ /*5670*/;
assign _22094_ = D[16] ^ Q[7] /*5666*/;
assign _22091_ = _21575_ & _22094_ /*5662*/;
assign _22092_ = _21575_ ^ _22094_ /*5665*/;
assign _22093_ = _22085_ & _22092_ /*5663*/;
assign _22090_ = _22091_ | _22093_ /*5661*/;
assign _21961_ = _22085_ ^ _22092_ /*5664*/;
assign _22099_ = D[17] ^ Q[7] /*5660*/;
assign _22096_ = _21576_ & _22099_ /*5656*/;
assign _22097_ = _21576_ ^ _22099_ /*5659*/;
assign _22098_ = _22090_ & _22097_ /*5657*/;
assign _22095_ = _22096_ | _22098_ /*5655*/;
assign _21962_ = _22090_ ^ _22097_ /*5658*/;
assign _22104_ = D[18] ^ Q[7] /*5654*/;
assign _22101_ = _21577_ & _22104_ /*5650*/;
assign _22102_ = _21577_ ^ _22104_ /*5653*/;
assign _22103_ = _22095_ & _22102_ /*5651*/;
assign _22100_ = _22101_ | _22103_ /*5649*/;
assign _21963_ = _22095_ ^ _22102_ /*5652*/;
assign _22109_ = D[19] ^ Q[7] /*5648*/;
assign _22106_ = _21578_ & _22109_ /*5644*/;
assign _22107_ = _21578_ ^ _22109_ /*5647*/;
assign _22108_ = _22100_ & _22107_ /*5645*/;
assign _22105_ = _22106_ | _22108_ /*5643*/;
assign _21964_ = _22100_ ^ _22107_ /*5646*/;
assign _22114_ = D[20] ^ Q[7] /*5642*/;
assign _22111_ = _21579_ & _22114_ /*5638*/;
assign _22112_ = _21579_ ^ _22114_ /*5641*/;
assign _22113_ = _22105_ & _22112_ /*5639*/;
assign _22110_ = _22111_ | _22113_ /*5637*/;
assign _21965_ = _22105_ ^ _22112_ /*5640*/;
assign _22119_ = D[21] ^ Q[7] /*5636*/;
assign _22116_ = _21580_ & _22119_ /*5632*/;
assign _22117_ = _21580_ ^ _22119_ /*5635*/;
assign _22118_ = _22110_ & _22117_ /*5633*/;
assign _22115_ = _22116_ | _22118_ /*5631*/;
assign _21966_ = _22110_ ^ _22117_ /*5634*/;
assign _22124_ = D[22] ^ Q[7] /*5630*/;
assign _22121_ = _21581_ & _22124_ /*5626*/;
assign _22122_ = _21581_ ^ _22124_ /*5629*/;
assign _22123_ = _22115_ & _22122_ /*5627*/;
assign _22120_ = _22121_ | _22123_ /*5625*/;
assign _21967_ = _22115_ ^ _22122_ /*5628*/;
assign _22129_ = D[23] ^ Q[7] /*5624*/;
assign _22126_ = _21582_ & _22129_ /*5620*/;
assign _22127_ = _21582_ ^ _22129_ /*5623*/;
assign _22128_ = _22120_ & _22127_ /*5621*/;
assign _22125_ = _22126_ | _22128_ /*5619*/;
assign _21968_ = _22120_ ^ _22127_ /*5622*/;
assign _22134_ = D[24] ^ Q[7] /*5618*/;
assign _22131_ = _21583_ & _22134_ /*5614*/;
assign _22132_ = _21583_ ^ _22134_ /*5617*/;
assign _22133_ = _22125_ & _22132_ /*5615*/;
assign _22130_ = _22131_ | _22133_ /*5613*/;
assign _21969_ = _22125_ ^ _22132_ /*5616*/;
assign _22139_ = D[25] ^ Q[7] /*5612*/;
assign _22136_ = _21584_ & _22139_ /*5608*/;
assign _22137_ = _21584_ ^ _22139_ /*5611*/;
assign _22138_ = _22130_ & _22137_ /*5609*/;
assign _22135_ = _22136_ | _22138_ /*5607*/;
assign _21970_ = _22130_ ^ _22137_ /*5610*/;
assign _22144_ = D[26] ^ Q[7] /*5606*/;
assign _22141_ = _21585_ & _22144_ /*5602*/;
assign _22142_ = _21585_ ^ _22144_ /*5605*/;
assign _22143_ = _22135_ & _22142_ /*5603*/;
assign _22140_ = _22141_ | _22143_ /*5601*/;
assign _21971_ = _22135_ ^ _22142_ /*5604*/;
assign _22149_ = D[27] ^ Q[7] /*5600*/;
assign _22146_ = _21586_ & _22149_ /*5596*/;
assign _22147_ = _21586_ ^ _22149_ /*5599*/;
assign _22148_ = _22140_ & _22147_ /*5597*/;
assign _22145_ = _22146_ | _22148_ /*5595*/;
assign _21972_ = _22140_ ^ _22147_ /*5598*/;
assign _22154_ = D[28] ^ Q[7] /*5594*/;
assign _22151_ = _21587_ & _22154_ /*5590*/;
assign _22152_ = _21587_ ^ _22154_ /*5593*/;
assign _22153_ = _22145_ & _22152_ /*5591*/;
assign _22150_ = _22151_ | _22153_ /*5589*/;
assign _21973_ = _22145_ ^ _22152_ /*5592*/;
assign _22159_ = D[29] ^ Q[7] /*5588*/;
assign _22156_ = _21588_ & _22159_ /*5584*/;
assign _22157_ = _21588_ ^ _22159_ /*5587*/;
assign _22158_ = _22150_ & _22157_ /*5585*/;
assign _22155_ = _22156_ | _22158_ /*5583*/;
assign _21974_ = _22150_ ^ _22157_ /*5586*/;
assign _22164_ = D[30] ^ Q[7] /*5582*/;
assign _22161_ = _21589_ & _22164_ /*5578*/;
assign _22162_ = _21589_ ^ _22164_ /*5581*/;
assign _22163_ = _22155_ & _22162_ /*5579*/;
assign _22160_ = _22161_ | _22163_ /*5577*/;
assign _21975_ = _22155_ ^ _22162_ /*5580*/;
assign _22169_ = D[31] ^ Q[7] /*5576*/;
assign _22166_ = _21590_ & _22169_ /*5572*/;
assign _22167_ = _21590_ ^ _22169_ /*5575*/;
assign _22168_ = _22160_ & _22167_ /*5573*/;
assign _22165_ = _22166_ | _22168_ /*5571*/;
assign _21976_ = _22160_ ^ _22167_ /*5574*/;
assign _22174_ = D[32] ^ Q[7] /*5570*/;
assign _22171_ = _21591_ & _22174_ /*5566*/;
assign _22172_ = _21591_ ^ _22174_ /*5569*/;
assign _22173_ = _22165_ & _22172_ /*5567*/;
assign _22170_ = _22171_ | _22173_ /*5565*/;
assign _21977_ = _22165_ ^ _22172_ /*5568*/;
assign _22179_ = D[33] ^ Q[7] /*5564*/;
assign _22176_ = _21592_ & _22179_ /*5560*/;
assign _22177_ = _21592_ ^ _22179_ /*5563*/;
assign _22178_ = _22170_ & _22177_ /*5561*/;
assign _22175_ = _22176_ | _22178_ /*5559*/;
assign _21978_ = _22170_ ^ _22177_ /*5562*/;
assign _22184_ = D[34] ^ Q[7] /*5558*/;
assign _22181_ = _21593_ & _22184_ /*5554*/;
assign _22182_ = _21593_ ^ _22184_ /*5557*/;
assign _22183_ = _22175_ & _22182_ /*5555*/;
assign _22180_ = _22181_ | _22183_ /*5553*/;
assign _21979_ = _22175_ ^ _22182_ /*5556*/;
assign _22189_ = D[35] ^ Q[7] /*5552*/;
assign _22186_ = _21594_ & _22189_ /*5548*/;
assign _22187_ = _21594_ ^ _22189_ /*5551*/;
assign _22188_ = _22180_ & _22187_ /*5549*/;
assign _22185_ = _22186_ | _22188_ /*5547*/;
assign _21980_ = _22180_ ^ _22187_ /*5550*/;
assign _22194_ = D[36] ^ Q[7] /*5546*/;
assign _22191_ = _21595_ & _22194_ /*5542*/;
assign _22192_ = _21595_ ^ _22194_ /*5545*/;
assign _22193_ = _22185_ & _22192_ /*5543*/;
assign _22190_ = _22191_ | _22193_ /*5541*/;
assign _21981_ = _22185_ ^ _22192_ /*5544*/;
assign _22199_ = D[37] ^ Q[7] /*5540*/;
assign _22196_ = _21596_ & _22199_ /*5536*/;
assign _22197_ = _21596_ ^ _22199_ /*5539*/;
assign _22198_ = _22190_ & _22197_ /*5537*/;
assign _22195_ = _22196_ | _22198_ /*5535*/;
assign _21982_ = _22190_ ^ _22197_ /*5538*/;
assign _22204_ = D[38] ^ Q[7] /*5534*/;
assign _22201_ = _21597_ & _22204_ /*5530*/;
assign _22202_ = _21597_ ^ _22204_ /*5533*/;
assign _22203_ = _22195_ & _22202_ /*5531*/;
assign _22200_ = _22201_ | _22203_ /*5529*/;
assign _21983_ = _22195_ ^ _22202_ /*5532*/;
assign _22209_ = D[39] ^ Q[7] /*5528*/;
assign _22206_ = _21598_ & _22209_ /*5524*/;
assign _22207_ = _21598_ ^ _22209_ /*5527*/;
assign _22208_ = _22200_ & _22207_ /*5525*/;
assign _22205_ = _22206_ | _22208_ /*5523*/;
assign _21984_ = _22200_ ^ _22207_ /*5526*/;
assign _22214_ = D[40] ^ Q[7] /*5522*/;
assign _22211_ = _21599_ & _22214_ /*5518*/;
assign _22212_ = _21599_ ^ _22214_ /*5521*/;
assign _22213_ = _22205_ & _22212_ /*5519*/;
assign _22210_ = _22211_ | _22213_ /*5517*/;
assign _21985_ = _22205_ ^ _22212_ /*5520*/;
assign _22219_ = D[41] ^ Q[7] /*5516*/;
assign _22216_ = _21600_ & _22219_ /*5512*/;
assign _22217_ = _21600_ ^ _22219_ /*5515*/;
assign _22218_ = _22210_ & _22217_ /*5513*/;
assign _22215_ = _22216_ | _22218_ /*5511*/;
assign _21986_ = _22210_ ^ _22217_ /*5514*/;
assign _22224_ = D[42] ^ Q[7] /*5510*/;
assign _22221_ = _21601_ & _22224_ /*5506*/;
assign _22222_ = _21601_ ^ _22224_ /*5509*/;
assign _22223_ = _22215_ & _22222_ /*5507*/;
assign _22220_ = _22221_ | _22223_ /*5505*/;
assign _21987_ = _22215_ ^ _22222_ /*5508*/;
assign _22229_ = D[43] ^ Q[7] /*5504*/;
assign _22226_ = _21602_ & _22229_ /*5500*/;
assign _22227_ = _21602_ ^ _22229_ /*5503*/;
assign _22228_ = _22220_ & _22227_ /*5501*/;
assign _22225_ = _22226_ | _22228_ /*5499*/;
assign _21988_ = _22220_ ^ _22227_ /*5502*/;
assign _22234_ = D[44] ^ Q[7] /*5498*/;
assign _22231_ = _21603_ & _22234_ /*5494*/;
assign _22232_ = _21603_ ^ _22234_ /*5497*/;
assign _22233_ = _22225_ & _22232_ /*5495*/;
assign _22230_ = _22231_ | _22233_ /*5493*/;
assign _21989_ = _22225_ ^ _22232_ /*5496*/;
assign _22239_ = D[45] ^ Q[7] /*5492*/;
assign _22236_ = _21604_ & _22239_ /*5488*/;
assign _22237_ = _21604_ ^ _22239_ /*5491*/;
assign _22238_ = _22230_ & _22237_ /*5489*/;
assign _22235_ = _22236_ | _22238_ /*5487*/;
assign _21990_ = _22230_ ^ _22237_ /*5490*/;
assign _22244_ = D[46] ^ Q[7] /*5486*/;
assign _22241_ = _21605_ & _22244_ /*5482*/;
assign _22242_ = _21605_ ^ _22244_ /*5485*/;
assign _22243_ = _22235_ & _22242_ /*5483*/;
assign _22240_ = _22241_ | _22243_ /*5481*/;
assign _21991_ = _22235_ ^ _22242_ /*5484*/;
assign _22249_ = D[47] ^ Q[7] /*5480*/;
assign _22246_ = _21606_ & _22249_ /*5476*/;
assign _22247_ = _21606_ ^ _22249_ /*5479*/;
assign _22248_ = _22240_ & _22247_ /*5477*/;
assign _22245_ = _22246_ | _22248_ /*5475*/;
assign _21992_ = _22240_ ^ _22247_ /*5478*/;
assign _22254_ = D[48] ^ Q[7] /*5474*/;
assign _22251_ = _21607_ & _22254_ /*5470*/;
assign _22252_ = _21607_ ^ _22254_ /*5473*/;
assign _22253_ = _22245_ & _22252_ /*5471*/;
assign _22250_ = _22251_ | _22253_ /*5469*/;
assign _21993_ = _22245_ ^ _22252_ /*5472*/;
assign _22259_ = D[49] ^ Q[7] /*5468*/;
assign _22256_ = _21608_ & _22259_ /*5464*/;
assign _22257_ = _21608_ ^ _22259_ /*5467*/;
assign _22258_ = _22250_ & _22257_ /*5465*/;
assign _22255_ = _22256_ | _22258_ /*5463*/;
assign _21994_ = _22250_ ^ _22257_ /*5466*/;
assign _22264_ = D[50] ^ Q[7] /*5462*/;
assign _22261_ = _21609_ & _22264_ /*5458*/;
assign _22262_ = _21609_ ^ _22264_ /*5461*/;
assign _22263_ = _22255_ & _22262_ /*5459*/;
assign _22260_ = _22261_ | _22263_ /*5457*/;
assign _21995_ = _22255_ ^ _22262_ /*5460*/;
assign _22269_ = D[51] ^ Q[7] /*5456*/;
assign _22266_ = _21610_ & _22269_ /*5452*/;
assign _22267_ = _21610_ ^ _22269_ /*5455*/;
assign _22268_ = _22260_ & _22267_ /*5453*/;
assign _22265_ = _22266_ | _22268_ /*5451*/;
assign _21996_ = _22260_ ^ _22267_ /*5454*/;
assign _22274_ = D[52] ^ Q[7] /*5450*/;
assign _22271_ = _21611_ & _22274_ /*5446*/;
assign _22272_ = _21611_ ^ _22274_ /*5449*/;
assign _22273_ = _22265_ & _22272_ /*5447*/;
assign _22270_ = _22271_ | _22273_ /*5445*/;
assign _21997_ = _22265_ ^ _22272_ /*5448*/;
assign _22279_ = D[53] ^ Q[7] /*5444*/;
assign _22276_ = _21612_ & _22279_ /*5440*/;
assign _22277_ = _21612_ ^ _22279_ /*5443*/;
assign _22278_ = _22270_ & _22277_ /*5441*/;
assign _22275_ = _22276_ | _22278_ /*5439*/;
assign _21998_ = _22270_ ^ _22277_ /*5442*/;
assign _22284_ = D[54] ^ Q[7] /*5438*/;
assign _22281_ = _21613_ & _22284_ /*5434*/;
assign _22282_ = _21613_ ^ _22284_ /*5437*/;
assign _22283_ = _22275_ & _22282_ /*5435*/;
assign _22280_ = _22281_ | _22283_ /*5433*/;
assign _21999_ = _22275_ ^ _22282_ /*5436*/;
assign _22289_ = D[55] ^ Q[7] /*5432*/;
assign _22286_ = _21614_ & _22289_ /*5428*/;
assign _22287_ = _21614_ ^ _22289_ /*5431*/;
assign _22288_ = _22280_ & _22287_ /*5429*/;
assign _22285_ = _22286_ | _22288_ /*5427*/;
assign _22000_ = _22280_ ^ _22287_ /*5430*/;
assign _22294_ = D[56] ^ Q[7] /*5426*/;
assign _22291_ = _21615_ & _22294_ /*5422*/;
assign _22292_ = _21615_ ^ _22294_ /*5425*/;
assign _22293_ = _22285_ & _22292_ /*5423*/;
assign _22290_ = _22291_ | _22293_ /*5421*/;
assign _22001_ = _22285_ ^ _22292_ /*5424*/;
assign _22299_ = D[57] ^ Q[7] /*5420*/;
assign _22296_ = _21616_ & _22299_ /*5416*/;
assign _22297_ = _21616_ ^ _22299_ /*5419*/;
assign _22298_ = _22290_ & _22297_ /*5417*/;
assign _22295_ = _22296_ | _22298_ /*5415*/;
assign _22002_ = _22290_ ^ _22297_ /*5418*/;
assign _22304_ = D[58] ^ Q[7] /*5414*/;
assign _22301_ = _21617_ & _22304_ /*5410*/;
assign _22302_ = _21617_ ^ _22304_ /*5413*/;
assign _22303_ = _22295_ & _22302_ /*5411*/;
assign _22300_ = _22301_ | _22303_ /*5409*/;
assign _22003_ = _22295_ ^ _22302_ /*5412*/;
assign _22309_ = D[59] ^ Q[7] /*5408*/;
assign _22306_ = _21618_ & _22309_ /*5404*/;
assign _22307_ = _21618_ ^ _22309_ /*5407*/;
assign _22308_ = _22300_ & _22307_ /*5405*/;
assign _22305_ = _22306_ | _22308_ /*5403*/;
assign _22004_ = _22300_ ^ _22307_ /*5406*/;
assign _22314_ = D[60] ^ Q[7] /*5402*/;
assign _22311_ = _21619_ & _22314_ /*5398*/;
assign _22312_ = _21619_ ^ _22314_ /*5401*/;
assign _22313_ = _22305_ & _22312_ /*5399*/;
assign _22310_ = _22311_ | _22313_ /*5397*/;
assign _22005_ = _22305_ ^ _22312_ /*5400*/;
assign _22319_ = D[61] ^ Q[7] /*5396*/;
assign _22316_ = _21620_ & _22319_ /*5392*/;
assign _22317_ = _21620_ ^ _22319_ /*5395*/;
assign _22318_ = _22310_ & _22317_ /*5393*/;
assign _22315_ = _22316_ | _22318_ /*5391*/;
assign _22006_ = _22310_ ^ _22317_ /*5394*/;
assign _22324_ = D[62] ^ Q[7] /*5390*/;
assign _22321_ = _21621_ & _22324_ /*5386*/;
assign _22322_ = _21621_ ^ _22324_ /*5389*/;
assign _22323_ = _22315_ & _22322_ /*5387*/;
assign _22320_ = _22321_ | _22323_ /*5385*/;
assign _22007_ = _22315_ ^ _22322_ /*5388*/;
assign _22328_ = zeroWire ^ Q[7] /*5384*/;
assign _22325_ = _21622_ & _22328_ /*5380*/;
assign _22326_ = _21622_ ^ _22328_ /*5383*/;
assign _22327_ = _22320_ & _22326_ /*5381*/;
assign Q[6] = _22325_ | _22327_ /*5379*/;
assign _22008_ = _22320_ ^ _22326_ /*5382*/;
assign _22399_ = D[0] ^ Q[6] /*4993*/;
assign _22396_ = R_0[5] & _22399_ /*4989*/;
assign _22397_ = R_0[5] ^ _22399_ /*4992*/;
assign _22398_ = Q[6] & _22397_ /*4990*/;
assign _22395_ = _22396_ | _22398_ /*4988*/;
assign _22330_ = Q[6] ^ _22397_ /*4991*/;
assign _22404_ = D[1] ^ Q[6] /*4987*/;
assign _22401_ = _21945_ & _22404_ /*4983*/;
assign _22402_ = _21945_ ^ _22404_ /*4986*/;
assign _22403_ = _22395_ & _22402_ /*4984*/;
assign _22400_ = _22401_ | _22403_ /*4982*/;
assign _22331_ = _22395_ ^ _22402_ /*4985*/;
assign _22409_ = D[2] ^ Q[6] /*4981*/;
assign _22406_ = _21946_ & _22409_ /*4977*/;
assign _22407_ = _21946_ ^ _22409_ /*4980*/;
assign _22408_ = _22400_ & _22407_ /*4978*/;
assign _22405_ = _22406_ | _22408_ /*4976*/;
assign _22332_ = _22400_ ^ _22407_ /*4979*/;
assign _22414_ = D[3] ^ Q[6] /*4975*/;
assign _22411_ = _21947_ & _22414_ /*4971*/;
assign _22412_ = _21947_ ^ _22414_ /*4974*/;
assign _22413_ = _22405_ & _22412_ /*4972*/;
assign _22410_ = _22411_ | _22413_ /*4970*/;
assign _22333_ = _22405_ ^ _22412_ /*4973*/;
assign _22419_ = D[4] ^ Q[6] /*4969*/;
assign _22416_ = _21948_ & _22419_ /*4965*/;
assign _22417_ = _21948_ ^ _22419_ /*4968*/;
assign _22418_ = _22410_ & _22417_ /*4966*/;
assign _22415_ = _22416_ | _22418_ /*4964*/;
assign _22334_ = _22410_ ^ _22417_ /*4967*/;
assign _22424_ = D[5] ^ Q[6] /*4963*/;
assign _22421_ = _21949_ & _22424_ /*4959*/;
assign _22422_ = _21949_ ^ _22424_ /*4962*/;
assign _22423_ = _22415_ & _22422_ /*4960*/;
assign _22420_ = _22421_ | _22423_ /*4958*/;
assign _22335_ = _22415_ ^ _22422_ /*4961*/;
assign _22429_ = D[6] ^ Q[6] /*4957*/;
assign _22426_ = _21950_ & _22429_ /*4953*/;
assign _22427_ = _21950_ ^ _22429_ /*4956*/;
assign _22428_ = _22420_ & _22427_ /*4954*/;
assign _22425_ = _22426_ | _22428_ /*4952*/;
assign _22336_ = _22420_ ^ _22427_ /*4955*/;
assign _22434_ = D[7] ^ Q[6] /*4951*/;
assign _22431_ = _21951_ & _22434_ /*4947*/;
assign _22432_ = _21951_ ^ _22434_ /*4950*/;
assign _22433_ = _22425_ & _22432_ /*4948*/;
assign _22430_ = _22431_ | _22433_ /*4946*/;
assign _22337_ = _22425_ ^ _22432_ /*4949*/;
assign _22439_ = D[8] ^ Q[6] /*4945*/;
assign _22436_ = _21952_ & _22439_ /*4941*/;
assign _22437_ = _21952_ ^ _22439_ /*4944*/;
assign _22438_ = _22430_ & _22437_ /*4942*/;
assign _22435_ = _22436_ | _22438_ /*4940*/;
assign _22338_ = _22430_ ^ _22437_ /*4943*/;
assign _22444_ = D[9] ^ Q[6] /*4939*/;
assign _22441_ = _21953_ & _22444_ /*4935*/;
assign _22442_ = _21953_ ^ _22444_ /*4938*/;
assign _22443_ = _22435_ & _22442_ /*4936*/;
assign _22440_ = _22441_ | _22443_ /*4934*/;
assign _22339_ = _22435_ ^ _22442_ /*4937*/;
assign _22449_ = D[10] ^ Q[6] /*4933*/;
assign _22446_ = _21954_ & _22449_ /*4929*/;
assign _22447_ = _21954_ ^ _22449_ /*4932*/;
assign _22448_ = _22440_ & _22447_ /*4930*/;
assign _22445_ = _22446_ | _22448_ /*4928*/;
assign _22340_ = _22440_ ^ _22447_ /*4931*/;
assign _22454_ = D[11] ^ Q[6] /*4927*/;
assign _22451_ = _21955_ & _22454_ /*4923*/;
assign _22452_ = _21955_ ^ _22454_ /*4926*/;
assign _22453_ = _22445_ & _22452_ /*4924*/;
assign _22450_ = _22451_ | _22453_ /*4922*/;
assign _22341_ = _22445_ ^ _22452_ /*4925*/;
assign _22459_ = D[12] ^ Q[6] /*4921*/;
assign _22456_ = _21956_ & _22459_ /*4917*/;
assign _22457_ = _21956_ ^ _22459_ /*4920*/;
assign _22458_ = _22450_ & _22457_ /*4918*/;
assign _22455_ = _22456_ | _22458_ /*4916*/;
assign _22342_ = _22450_ ^ _22457_ /*4919*/;
assign _22464_ = D[13] ^ Q[6] /*4915*/;
assign _22461_ = _21957_ & _22464_ /*4911*/;
assign _22462_ = _21957_ ^ _22464_ /*4914*/;
assign _22463_ = _22455_ & _22462_ /*4912*/;
assign _22460_ = _22461_ | _22463_ /*4910*/;
assign _22343_ = _22455_ ^ _22462_ /*4913*/;
assign _22469_ = D[14] ^ Q[6] /*4909*/;
assign _22466_ = _21958_ & _22469_ /*4905*/;
assign _22467_ = _21958_ ^ _22469_ /*4908*/;
assign _22468_ = _22460_ & _22467_ /*4906*/;
assign _22465_ = _22466_ | _22468_ /*4904*/;
assign _22344_ = _22460_ ^ _22467_ /*4907*/;
assign _22474_ = D[15] ^ Q[6] /*4903*/;
assign _22471_ = _21959_ & _22474_ /*4899*/;
assign _22472_ = _21959_ ^ _22474_ /*4902*/;
assign _22473_ = _22465_ & _22472_ /*4900*/;
assign _22470_ = _22471_ | _22473_ /*4898*/;
assign _22345_ = _22465_ ^ _22472_ /*4901*/;
assign _22479_ = D[16] ^ Q[6] /*4897*/;
assign _22476_ = _21960_ & _22479_ /*4893*/;
assign _22477_ = _21960_ ^ _22479_ /*4896*/;
assign _22478_ = _22470_ & _22477_ /*4894*/;
assign _22475_ = _22476_ | _22478_ /*4892*/;
assign _22346_ = _22470_ ^ _22477_ /*4895*/;
assign _22484_ = D[17] ^ Q[6] /*4891*/;
assign _22481_ = _21961_ & _22484_ /*4887*/;
assign _22482_ = _21961_ ^ _22484_ /*4890*/;
assign _22483_ = _22475_ & _22482_ /*4888*/;
assign _22480_ = _22481_ | _22483_ /*4886*/;
assign _22347_ = _22475_ ^ _22482_ /*4889*/;
assign _22489_ = D[18] ^ Q[6] /*4885*/;
assign _22486_ = _21962_ & _22489_ /*4881*/;
assign _22487_ = _21962_ ^ _22489_ /*4884*/;
assign _22488_ = _22480_ & _22487_ /*4882*/;
assign _22485_ = _22486_ | _22488_ /*4880*/;
assign _22348_ = _22480_ ^ _22487_ /*4883*/;
assign _22494_ = D[19] ^ Q[6] /*4879*/;
assign _22491_ = _21963_ & _22494_ /*4875*/;
assign _22492_ = _21963_ ^ _22494_ /*4878*/;
assign _22493_ = _22485_ & _22492_ /*4876*/;
assign _22490_ = _22491_ | _22493_ /*4874*/;
assign _22349_ = _22485_ ^ _22492_ /*4877*/;
assign _22499_ = D[20] ^ Q[6] /*4873*/;
assign _22496_ = _21964_ & _22499_ /*4869*/;
assign _22497_ = _21964_ ^ _22499_ /*4872*/;
assign _22498_ = _22490_ & _22497_ /*4870*/;
assign _22495_ = _22496_ | _22498_ /*4868*/;
assign _22350_ = _22490_ ^ _22497_ /*4871*/;
assign _22504_ = D[21] ^ Q[6] /*4867*/;
assign _22501_ = _21965_ & _22504_ /*4863*/;
assign _22502_ = _21965_ ^ _22504_ /*4866*/;
assign _22503_ = _22495_ & _22502_ /*4864*/;
assign _22500_ = _22501_ | _22503_ /*4862*/;
assign _22351_ = _22495_ ^ _22502_ /*4865*/;
assign _22509_ = D[22] ^ Q[6] /*4861*/;
assign _22506_ = _21966_ & _22509_ /*4857*/;
assign _22507_ = _21966_ ^ _22509_ /*4860*/;
assign _22508_ = _22500_ & _22507_ /*4858*/;
assign _22505_ = _22506_ | _22508_ /*4856*/;
assign _22352_ = _22500_ ^ _22507_ /*4859*/;
assign _22514_ = D[23] ^ Q[6] /*4855*/;
assign _22511_ = _21967_ & _22514_ /*4851*/;
assign _22512_ = _21967_ ^ _22514_ /*4854*/;
assign _22513_ = _22505_ & _22512_ /*4852*/;
assign _22510_ = _22511_ | _22513_ /*4850*/;
assign _22353_ = _22505_ ^ _22512_ /*4853*/;
assign _22519_ = D[24] ^ Q[6] /*4849*/;
assign _22516_ = _21968_ & _22519_ /*4845*/;
assign _22517_ = _21968_ ^ _22519_ /*4848*/;
assign _22518_ = _22510_ & _22517_ /*4846*/;
assign _22515_ = _22516_ | _22518_ /*4844*/;
assign _22354_ = _22510_ ^ _22517_ /*4847*/;
assign _22524_ = D[25] ^ Q[6] /*4843*/;
assign _22521_ = _21969_ & _22524_ /*4839*/;
assign _22522_ = _21969_ ^ _22524_ /*4842*/;
assign _22523_ = _22515_ & _22522_ /*4840*/;
assign _22520_ = _22521_ | _22523_ /*4838*/;
assign _22355_ = _22515_ ^ _22522_ /*4841*/;
assign _22529_ = D[26] ^ Q[6] /*4837*/;
assign _22526_ = _21970_ & _22529_ /*4833*/;
assign _22527_ = _21970_ ^ _22529_ /*4836*/;
assign _22528_ = _22520_ & _22527_ /*4834*/;
assign _22525_ = _22526_ | _22528_ /*4832*/;
assign _22356_ = _22520_ ^ _22527_ /*4835*/;
assign _22534_ = D[27] ^ Q[6] /*4831*/;
assign _22531_ = _21971_ & _22534_ /*4827*/;
assign _22532_ = _21971_ ^ _22534_ /*4830*/;
assign _22533_ = _22525_ & _22532_ /*4828*/;
assign _22530_ = _22531_ | _22533_ /*4826*/;
assign _22357_ = _22525_ ^ _22532_ /*4829*/;
assign _22539_ = D[28] ^ Q[6] /*4825*/;
assign _22536_ = _21972_ & _22539_ /*4821*/;
assign _22537_ = _21972_ ^ _22539_ /*4824*/;
assign _22538_ = _22530_ & _22537_ /*4822*/;
assign _22535_ = _22536_ | _22538_ /*4820*/;
assign _22358_ = _22530_ ^ _22537_ /*4823*/;
assign _22544_ = D[29] ^ Q[6] /*4819*/;
assign _22541_ = _21973_ & _22544_ /*4815*/;
assign _22542_ = _21973_ ^ _22544_ /*4818*/;
assign _22543_ = _22535_ & _22542_ /*4816*/;
assign _22540_ = _22541_ | _22543_ /*4814*/;
assign _22359_ = _22535_ ^ _22542_ /*4817*/;
assign _22549_ = D[30] ^ Q[6] /*4813*/;
assign _22546_ = _21974_ & _22549_ /*4809*/;
assign _22547_ = _21974_ ^ _22549_ /*4812*/;
assign _22548_ = _22540_ & _22547_ /*4810*/;
assign _22545_ = _22546_ | _22548_ /*4808*/;
assign _22360_ = _22540_ ^ _22547_ /*4811*/;
assign _22554_ = D[31] ^ Q[6] /*4807*/;
assign _22551_ = _21975_ & _22554_ /*4803*/;
assign _22552_ = _21975_ ^ _22554_ /*4806*/;
assign _22553_ = _22545_ & _22552_ /*4804*/;
assign _22550_ = _22551_ | _22553_ /*4802*/;
assign _22361_ = _22545_ ^ _22552_ /*4805*/;
assign _22559_ = D[32] ^ Q[6] /*4801*/;
assign _22556_ = _21976_ & _22559_ /*4797*/;
assign _22557_ = _21976_ ^ _22559_ /*4800*/;
assign _22558_ = _22550_ & _22557_ /*4798*/;
assign _22555_ = _22556_ | _22558_ /*4796*/;
assign _22362_ = _22550_ ^ _22557_ /*4799*/;
assign _22564_ = D[33] ^ Q[6] /*4795*/;
assign _22561_ = _21977_ & _22564_ /*4791*/;
assign _22562_ = _21977_ ^ _22564_ /*4794*/;
assign _22563_ = _22555_ & _22562_ /*4792*/;
assign _22560_ = _22561_ | _22563_ /*4790*/;
assign _22363_ = _22555_ ^ _22562_ /*4793*/;
assign _22569_ = D[34] ^ Q[6] /*4789*/;
assign _22566_ = _21978_ & _22569_ /*4785*/;
assign _22567_ = _21978_ ^ _22569_ /*4788*/;
assign _22568_ = _22560_ & _22567_ /*4786*/;
assign _22565_ = _22566_ | _22568_ /*4784*/;
assign _22364_ = _22560_ ^ _22567_ /*4787*/;
assign _22574_ = D[35] ^ Q[6] /*4783*/;
assign _22571_ = _21979_ & _22574_ /*4779*/;
assign _22572_ = _21979_ ^ _22574_ /*4782*/;
assign _22573_ = _22565_ & _22572_ /*4780*/;
assign _22570_ = _22571_ | _22573_ /*4778*/;
assign _22365_ = _22565_ ^ _22572_ /*4781*/;
assign _22579_ = D[36] ^ Q[6] /*4777*/;
assign _22576_ = _21980_ & _22579_ /*4773*/;
assign _22577_ = _21980_ ^ _22579_ /*4776*/;
assign _22578_ = _22570_ & _22577_ /*4774*/;
assign _22575_ = _22576_ | _22578_ /*4772*/;
assign _22366_ = _22570_ ^ _22577_ /*4775*/;
assign _22584_ = D[37] ^ Q[6] /*4771*/;
assign _22581_ = _21981_ & _22584_ /*4767*/;
assign _22582_ = _21981_ ^ _22584_ /*4770*/;
assign _22583_ = _22575_ & _22582_ /*4768*/;
assign _22580_ = _22581_ | _22583_ /*4766*/;
assign _22367_ = _22575_ ^ _22582_ /*4769*/;
assign _22589_ = D[38] ^ Q[6] /*4765*/;
assign _22586_ = _21982_ & _22589_ /*4761*/;
assign _22587_ = _21982_ ^ _22589_ /*4764*/;
assign _22588_ = _22580_ & _22587_ /*4762*/;
assign _22585_ = _22586_ | _22588_ /*4760*/;
assign _22368_ = _22580_ ^ _22587_ /*4763*/;
assign _22594_ = D[39] ^ Q[6] /*4759*/;
assign _22591_ = _21983_ & _22594_ /*4755*/;
assign _22592_ = _21983_ ^ _22594_ /*4758*/;
assign _22593_ = _22585_ & _22592_ /*4756*/;
assign _22590_ = _22591_ | _22593_ /*4754*/;
assign _22369_ = _22585_ ^ _22592_ /*4757*/;
assign _22599_ = D[40] ^ Q[6] /*4753*/;
assign _22596_ = _21984_ & _22599_ /*4749*/;
assign _22597_ = _21984_ ^ _22599_ /*4752*/;
assign _22598_ = _22590_ & _22597_ /*4750*/;
assign _22595_ = _22596_ | _22598_ /*4748*/;
assign _22370_ = _22590_ ^ _22597_ /*4751*/;
assign _22604_ = D[41] ^ Q[6] /*4747*/;
assign _22601_ = _21985_ & _22604_ /*4743*/;
assign _22602_ = _21985_ ^ _22604_ /*4746*/;
assign _22603_ = _22595_ & _22602_ /*4744*/;
assign _22600_ = _22601_ | _22603_ /*4742*/;
assign _22371_ = _22595_ ^ _22602_ /*4745*/;
assign _22609_ = D[42] ^ Q[6] /*4741*/;
assign _22606_ = _21986_ & _22609_ /*4737*/;
assign _22607_ = _21986_ ^ _22609_ /*4740*/;
assign _22608_ = _22600_ & _22607_ /*4738*/;
assign _22605_ = _22606_ | _22608_ /*4736*/;
assign _22372_ = _22600_ ^ _22607_ /*4739*/;
assign _22614_ = D[43] ^ Q[6] /*4735*/;
assign _22611_ = _21987_ & _22614_ /*4731*/;
assign _22612_ = _21987_ ^ _22614_ /*4734*/;
assign _22613_ = _22605_ & _22612_ /*4732*/;
assign _22610_ = _22611_ | _22613_ /*4730*/;
assign _22373_ = _22605_ ^ _22612_ /*4733*/;
assign _22619_ = D[44] ^ Q[6] /*4729*/;
assign _22616_ = _21988_ & _22619_ /*4725*/;
assign _22617_ = _21988_ ^ _22619_ /*4728*/;
assign _22618_ = _22610_ & _22617_ /*4726*/;
assign _22615_ = _22616_ | _22618_ /*4724*/;
assign _22374_ = _22610_ ^ _22617_ /*4727*/;
assign _22624_ = D[45] ^ Q[6] /*4723*/;
assign _22621_ = _21989_ & _22624_ /*4719*/;
assign _22622_ = _21989_ ^ _22624_ /*4722*/;
assign _22623_ = _22615_ & _22622_ /*4720*/;
assign _22620_ = _22621_ | _22623_ /*4718*/;
assign _22375_ = _22615_ ^ _22622_ /*4721*/;
assign _22629_ = D[46] ^ Q[6] /*4717*/;
assign _22626_ = _21990_ & _22629_ /*4713*/;
assign _22627_ = _21990_ ^ _22629_ /*4716*/;
assign _22628_ = _22620_ & _22627_ /*4714*/;
assign _22625_ = _22626_ | _22628_ /*4712*/;
assign _22376_ = _22620_ ^ _22627_ /*4715*/;
assign _22634_ = D[47] ^ Q[6] /*4711*/;
assign _22631_ = _21991_ & _22634_ /*4707*/;
assign _22632_ = _21991_ ^ _22634_ /*4710*/;
assign _22633_ = _22625_ & _22632_ /*4708*/;
assign _22630_ = _22631_ | _22633_ /*4706*/;
assign _22377_ = _22625_ ^ _22632_ /*4709*/;
assign _22639_ = D[48] ^ Q[6] /*4705*/;
assign _22636_ = _21992_ & _22639_ /*4701*/;
assign _22637_ = _21992_ ^ _22639_ /*4704*/;
assign _22638_ = _22630_ & _22637_ /*4702*/;
assign _22635_ = _22636_ | _22638_ /*4700*/;
assign _22378_ = _22630_ ^ _22637_ /*4703*/;
assign _22644_ = D[49] ^ Q[6] /*4699*/;
assign _22641_ = _21993_ & _22644_ /*4695*/;
assign _22642_ = _21993_ ^ _22644_ /*4698*/;
assign _22643_ = _22635_ & _22642_ /*4696*/;
assign _22640_ = _22641_ | _22643_ /*4694*/;
assign _22379_ = _22635_ ^ _22642_ /*4697*/;
assign _22649_ = D[50] ^ Q[6] /*4693*/;
assign _22646_ = _21994_ & _22649_ /*4689*/;
assign _22647_ = _21994_ ^ _22649_ /*4692*/;
assign _22648_ = _22640_ & _22647_ /*4690*/;
assign _22645_ = _22646_ | _22648_ /*4688*/;
assign _22380_ = _22640_ ^ _22647_ /*4691*/;
assign _22654_ = D[51] ^ Q[6] /*4687*/;
assign _22651_ = _21995_ & _22654_ /*4683*/;
assign _22652_ = _21995_ ^ _22654_ /*4686*/;
assign _22653_ = _22645_ & _22652_ /*4684*/;
assign _22650_ = _22651_ | _22653_ /*4682*/;
assign _22381_ = _22645_ ^ _22652_ /*4685*/;
assign _22659_ = D[52] ^ Q[6] /*4681*/;
assign _22656_ = _21996_ & _22659_ /*4677*/;
assign _22657_ = _21996_ ^ _22659_ /*4680*/;
assign _22658_ = _22650_ & _22657_ /*4678*/;
assign _22655_ = _22656_ | _22658_ /*4676*/;
assign _22382_ = _22650_ ^ _22657_ /*4679*/;
assign _22664_ = D[53] ^ Q[6] /*4675*/;
assign _22661_ = _21997_ & _22664_ /*4671*/;
assign _22662_ = _21997_ ^ _22664_ /*4674*/;
assign _22663_ = _22655_ & _22662_ /*4672*/;
assign _22660_ = _22661_ | _22663_ /*4670*/;
assign _22383_ = _22655_ ^ _22662_ /*4673*/;
assign _22669_ = D[54] ^ Q[6] /*4669*/;
assign _22666_ = _21998_ & _22669_ /*4665*/;
assign _22667_ = _21998_ ^ _22669_ /*4668*/;
assign _22668_ = _22660_ & _22667_ /*4666*/;
assign _22665_ = _22666_ | _22668_ /*4664*/;
assign _22384_ = _22660_ ^ _22667_ /*4667*/;
assign _22674_ = D[55] ^ Q[6] /*4663*/;
assign _22671_ = _21999_ & _22674_ /*4659*/;
assign _22672_ = _21999_ ^ _22674_ /*4662*/;
assign _22673_ = _22665_ & _22672_ /*4660*/;
assign _22670_ = _22671_ | _22673_ /*4658*/;
assign _22385_ = _22665_ ^ _22672_ /*4661*/;
assign _22679_ = D[56] ^ Q[6] /*4657*/;
assign _22676_ = _22000_ & _22679_ /*4653*/;
assign _22677_ = _22000_ ^ _22679_ /*4656*/;
assign _22678_ = _22670_ & _22677_ /*4654*/;
assign _22675_ = _22676_ | _22678_ /*4652*/;
assign _22386_ = _22670_ ^ _22677_ /*4655*/;
assign _22684_ = D[57] ^ Q[6] /*4651*/;
assign _22681_ = _22001_ & _22684_ /*4647*/;
assign _22682_ = _22001_ ^ _22684_ /*4650*/;
assign _22683_ = _22675_ & _22682_ /*4648*/;
assign _22680_ = _22681_ | _22683_ /*4646*/;
assign _22387_ = _22675_ ^ _22682_ /*4649*/;
assign _22689_ = D[58] ^ Q[6] /*4645*/;
assign _22686_ = _22002_ & _22689_ /*4641*/;
assign _22687_ = _22002_ ^ _22689_ /*4644*/;
assign _22688_ = _22680_ & _22687_ /*4642*/;
assign _22685_ = _22686_ | _22688_ /*4640*/;
assign _22388_ = _22680_ ^ _22687_ /*4643*/;
assign _22694_ = D[59] ^ Q[6] /*4639*/;
assign _22691_ = _22003_ & _22694_ /*4635*/;
assign _22692_ = _22003_ ^ _22694_ /*4638*/;
assign _22693_ = _22685_ & _22692_ /*4636*/;
assign _22690_ = _22691_ | _22693_ /*4634*/;
assign _22389_ = _22685_ ^ _22692_ /*4637*/;
assign _22699_ = D[60] ^ Q[6] /*4633*/;
assign _22696_ = _22004_ & _22699_ /*4629*/;
assign _22697_ = _22004_ ^ _22699_ /*4632*/;
assign _22698_ = _22690_ & _22697_ /*4630*/;
assign _22695_ = _22696_ | _22698_ /*4628*/;
assign _22390_ = _22690_ ^ _22697_ /*4631*/;
assign _22704_ = D[61] ^ Q[6] /*4627*/;
assign _22701_ = _22005_ & _22704_ /*4623*/;
assign _22702_ = _22005_ ^ _22704_ /*4626*/;
assign _22703_ = _22695_ & _22702_ /*4624*/;
assign _22700_ = _22701_ | _22703_ /*4622*/;
assign _22391_ = _22695_ ^ _22702_ /*4625*/;
assign _22709_ = D[62] ^ Q[6] /*4621*/;
assign _22706_ = _22006_ & _22709_ /*4617*/;
assign _22707_ = _22006_ ^ _22709_ /*4620*/;
assign _22708_ = _22700_ & _22707_ /*4618*/;
assign _22705_ = _22706_ | _22708_ /*4616*/;
assign _22392_ = _22700_ ^ _22707_ /*4619*/;
assign _22713_ = zeroWire ^ Q[6] /*4615*/;
assign _22710_ = _22007_ & _22713_ /*4611*/;
assign _22711_ = _22007_ ^ _22713_ /*4614*/;
assign _22712_ = _22705_ & _22711_ /*4612*/;
assign Q[5] = _22710_ | _22712_ /*4610*/;
assign _22393_ = _22705_ ^ _22711_ /*4613*/;
assign _22784_ = D[0] ^ Q[5] /*4224*/;
assign _22781_ = R_0[4] & _22784_ /*4220*/;
assign _22782_ = R_0[4] ^ _22784_ /*4223*/;
assign _22783_ = Q[5] & _22782_ /*4221*/;
assign _22780_ = _22781_ | _22783_ /*4219*/;
assign _22715_ = Q[5] ^ _22782_ /*4222*/;
assign _22789_ = D[1] ^ Q[5] /*4218*/;
assign _22786_ = _22330_ & _22789_ /*4214*/;
assign _22787_ = _22330_ ^ _22789_ /*4217*/;
assign _22788_ = _22780_ & _22787_ /*4215*/;
assign _22785_ = _22786_ | _22788_ /*4213*/;
assign _22716_ = _22780_ ^ _22787_ /*4216*/;
assign _22794_ = D[2] ^ Q[5] /*4212*/;
assign _22791_ = _22331_ & _22794_ /*4208*/;
assign _22792_ = _22331_ ^ _22794_ /*4211*/;
assign _22793_ = _22785_ & _22792_ /*4209*/;
assign _22790_ = _22791_ | _22793_ /*4207*/;
assign _22717_ = _22785_ ^ _22792_ /*4210*/;
assign _22799_ = D[3] ^ Q[5] /*4206*/;
assign _22796_ = _22332_ & _22799_ /*4202*/;
assign _22797_ = _22332_ ^ _22799_ /*4205*/;
assign _22798_ = _22790_ & _22797_ /*4203*/;
assign _22795_ = _22796_ | _22798_ /*4201*/;
assign _22718_ = _22790_ ^ _22797_ /*4204*/;
assign _22804_ = D[4] ^ Q[5] /*4200*/;
assign _22801_ = _22333_ & _22804_ /*4196*/;
assign _22802_ = _22333_ ^ _22804_ /*4199*/;
assign _22803_ = _22795_ & _22802_ /*4197*/;
assign _22800_ = _22801_ | _22803_ /*4195*/;
assign _22719_ = _22795_ ^ _22802_ /*4198*/;
assign _22809_ = D[5] ^ Q[5] /*4194*/;
assign _22806_ = _22334_ & _22809_ /*4190*/;
assign _22807_ = _22334_ ^ _22809_ /*4193*/;
assign _22808_ = _22800_ & _22807_ /*4191*/;
assign _22805_ = _22806_ | _22808_ /*4189*/;
assign _22720_ = _22800_ ^ _22807_ /*4192*/;
assign _22814_ = D[6] ^ Q[5] /*4188*/;
assign _22811_ = _22335_ & _22814_ /*4184*/;
assign _22812_ = _22335_ ^ _22814_ /*4187*/;
assign _22813_ = _22805_ & _22812_ /*4185*/;
assign _22810_ = _22811_ | _22813_ /*4183*/;
assign _22721_ = _22805_ ^ _22812_ /*4186*/;
assign _22819_ = D[7] ^ Q[5] /*4182*/;
assign _22816_ = _22336_ & _22819_ /*4178*/;
assign _22817_ = _22336_ ^ _22819_ /*4181*/;
assign _22818_ = _22810_ & _22817_ /*4179*/;
assign _22815_ = _22816_ | _22818_ /*4177*/;
assign _22722_ = _22810_ ^ _22817_ /*4180*/;
assign _22824_ = D[8] ^ Q[5] /*4176*/;
assign _22821_ = _22337_ & _22824_ /*4172*/;
assign _22822_ = _22337_ ^ _22824_ /*4175*/;
assign _22823_ = _22815_ & _22822_ /*4173*/;
assign _22820_ = _22821_ | _22823_ /*4171*/;
assign _22723_ = _22815_ ^ _22822_ /*4174*/;
assign _22829_ = D[9] ^ Q[5] /*4170*/;
assign _22826_ = _22338_ & _22829_ /*4166*/;
assign _22827_ = _22338_ ^ _22829_ /*4169*/;
assign _22828_ = _22820_ & _22827_ /*4167*/;
assign _22825_ = _22826_ | _22828_ /*4165*/;
assign _22724_ = _22820_ ^ _22827_ /*4168*/;
assign _22834_ = D[10] ^ Q[5] /*4164*/;
assign _22831_ = _22339_ & _22834_ /*4160*/;
assign _22832_ = _22339_ ^ _22834_ /*4163*/;
assign _22833_ = _22825_ & _22832_ /*4161*/;
assign _22830_ = _22831_ | _22833_ /*4159*/;
assign _22725_ = _22825_ ^ _22832_ /*4162*/;
assign _22839_ = D[11] ^ Q[5] /*4158*/;
assign _22836_ = _22340_ & _22839_ /*4154*/;
assign _22837_ = _22340_ ^ _22839_ /*4157*/;
assign _22838_ = _22830_ & _22837_ /*4155*/;
assign _22835_ = _22836_ | _22838_ /*4153*/;
assign _22726_ = _22830_ ^ _22837_ /*4156*/;
assign _22844_ = D[12] ^ Q[5] /*4152*/;
assign _22841_ = _22341_ & _22844_ /*4148*/;
assign _22842_ = _22341_ ^ _22844_ /*4151*/;
assign _22843_ = _22835_ & _22842_ /*4149*/;
assign _22840_ = _22841_ | _22843_ /*4147*/;
assign _22727_ = _22835_ ^ _22842_ /*4150*/;
assign _22849_ = D[13] ^ Q[5] /*4146*/;
assign _22846_ = _22342_ & _22849_ /*4142*/;
assign _22847_ = _22342_ ^ _22849_ /*4145*/;
assign _22848_ = _22840_ & _22847_ /*4143*/;
assign _22845_ = _22846_ | _22848_ /*4141*/;
assign _22728_ = _22840_ ^ _22847_ /*4144*/;
assign _22854_ = D[14] ^ Q[5] /*4140*/;
assign _22851_ = _22343_ & _22854_ /*4136*/;
assign _22852_ = _22343_ ^ _22854_ /*4139*/;
assign _22853_ = _22845_ & _22852_ /*4137*/;
assign _22850_ = _22851_ | _22853_ /*4135*/;
assign _22729_ = _22845_ ^ _22852_ /*4138*/;
assign _22859_ = D[15] ^ Q[5] /*4134*/;
assign _22856_ = _22344_ & _22859_ /*4130*/;
assign _22857_ = _22344_ ^ _22859_ /*4133*/;
assign _22858_ = _22850_ & _22857_ /*4131*/;
assign _22855_ = _22856_ | _22858_ /*4129*/;
assign _22730_ = _22850_ ^ _22857_ /*4132*/;
assign _22864_ = D[16] ^ Q[5] /*4128*/;
assign _22861_ = _22345_ & _22864_ /*4124*/;
assign _22862_ = _22345_ ^ _22864_ /*4127*/;
assign _22863_ = _22855_ & _22862_ /*4125*/;
assign _22860_ = _22861_ | _22863_ /*4123*/;
assign _22731_ = _22855_ ^ _22862_ /*4126*/;
assign _22869_ = D[17] ^ Q[5] /*4122*/;
assign _22866_ = _22346_ & _22869_ /*4118*/;
assign _22867_ = _22346_ ^ _22869_ /*4121*/;
assign _22868_ = _22860_ & _22867_ /*4119*/;
assign _22865_ = _22866_ | _22868_ /*4117*/;
assign _22732_ = _22860_ ^ _22867_ /*4120*/;
assign _22874_ = D[18] ^ Q[5] /*4116*/;
assign _22871_ = _22347_ & _22874_ /*4112*/;
assign _22872_ = _22347_ ^ _22874_ /*4115*/;
assign _22873_ = _22865_ & _22872_ /*4113*/;
assign _22870_ = _22871_ | _22873_ /*4111*/;
assign _22733_ = _22865_ ^ _22872_ /*4114*/;
assign _22879_ = D[19] ^ Q[5] /*4110*/;
assign _22876_ = _22348_ & _22879_ /*4106*/;
assign _22877_ = _22348_ ^ _22879_ /*4109*/;
assign _22878_ = _22870_ & _22877_ /*4107*/;
assign _22875_ = _22876_ | _22878_ /*4105*/;
assign _22734_ = _22870_ ^ _22877_ /*4108*/;
assign _22884_ = D[20] ^ Q[5] /*4104*/;
assign _22881_ = _22349_ & _22884_ /*4100*/;
assign _22882_ = _22349_ ^ _22884_ /*4103*/;
assign _22883_ = _22875_ & _22882_ /*4101*/;
assign _22880_ = _22881_ | _22883_ /*4099*/;
assign _22735_ = _22875_ ^ _22882_ /*4102*/;
assign _22889_ = D[21] ^ Q[5] /*4098*/;
assign _22886_ = _22350_ & _22889_ /*4094*/;
assign _22887_ = _22350_ ^ _22889_ /*4097*/;
assign _22888_ = _22880_ & _22887_ /*4095*/;
assign _22885_ = _22886_ | _22888_ /*4093*/;
assign _22736_ = _22880_ ^ _22887_ /*4096*/;
assign _22894_ = D[22] ^ Q[5] /*4092*/;
assign _22891_ = _22351_ & _22894_ /*4088*/;
assign _22892_ = _22351_ ^ _22894_ /*4091*/;
assign _22893_ = _22885_ & _22892_ /*4089*/;
assign _22890_ = _22891_ | _22893_ /*4087*/;
assign _22737_ = _22885_ ^ _22892_ /*4090*/;
assign _22899_ = D[23] ^ Q[5] /*4086*/;
assign _22896_ = _22352_ & _22899_ /*4082*/;
assign _22897_ = _22352_ ^ _22899_ /*4085*/;
assign _22898_ = _22890_ & _22897_ /*4083*/;
assign _22895_ = _22896_ | _22898_ /*4081*/;
assign _22738_ = _22890_ ^ _22897_ /*4084*/;
assign _22904_ = D[24] ^ Q[5] /*4080*/;
assign _22901_ = _22353_ & _22904_ /*4076*/;
assign _22902_ = _22353_ ^ _22904_ /*4079*/;
assign _22903_ = _22895_ & _22902_ /*4077*/;
assign _22900_ = _22901_ | _22903_ /*4075*/;
assign _22739_ = _22895_ ^ _22902_ /*4078*/;
assign _22909_ = D[25] ^ Q[5] /*4074*/;
assign _22906_ = _22354_ & _22909_ /*4070*/;
assign _22907_ = _22354_ ^ _22909_ /*4073*/;
assign _22908_ = _22900_ & _22907_ /*4071*/;
assign _22905_ = _22906_ | _22908_ /*4069*/;
assign _22740_ = _22900_ ^ _22907_ /*4072*/;
assign _22914_ = D[26] ^ Q[5] /*4068*/;
assign _22911_ = _22355_ & _22914_ /*4064*/;
assign _22912_ = _22355_ ^ _22914_ /*4067*/;
assign _22913_ = _22905_ & _22912_ /*4065*/;
assign _22910_ = _22911_ | _22913_ /*4063*/;
assign _22741_ = _22905_ ^ _22912_ /*4066*/;
assign _22919_ = D[27] ^ Q[5] /*4062*/;
assign _22916_ = _22356_ & _22919_ /*4058*/;
assign _22917_ = _22356_ ^ _22919_ /*4061*/;
assign _22918_ = _22910_ & _22917_ /*4059*/;
assign _22915_ = _22916_ | _22918_ /*4057*/;
assign _22742_ = _22910_ ^ _22917_ /*4060*/;
assign _22924_ = D[28] ^ Q[5] /*4056*/;
assign _22921_ = _22357_ & _22924_ /*4052*/;
assign _22922_ = _22357_ ^ _22924_ /*4055*/;
assign _22923_ = _22915_ & _22922_ /*4053*/;
assign _22920_ = _22921_ | _22923_ /*4051*/;
assign _22743_ = _22915_ ^ _22922_ /*4054*/;
assign _22929_ = D[29] ^ Q[5] /*4050*/;
assign _22926_ = _22358_ & _22929_ /*4046*/;
assign _22927_ = _22358_ ^ _22929_ /*4049*/;
assign _22928_ = _22920_ & _22927_ /*4047*/;
assign _22925_ = _22926_ | _22928_ /*4045*/;
assign _22744_ = _22920_ ^ _22927_ /*4048*/;
assign _22934_ = D[30] ^ Q[5] /*4044*/;
assign _22931_ = _22359_ & _22934_ /*4040*/;
assign _22932_ = _22359_ ^ _22934_ /*4043*/;
assign _22933_ = _22925_ & _22932_ /*4041*/;
assign _22930_ = _22931_ | _22933_ /*4039*/;
assign _22745_ = _22925_ ^ _22932_ /*4042*/;
assign _22939_ = D[31] ^ Q[5] /*4038*/;
assign _22936_ = _22360_ & _22939_ /*4034*/;
assign _22937_ = _22360_ ^ _22939_ /*4037*/;
assign _22938_ = _22930_ & _22937_ /*4035*/;
assign _22935_ = _22936_ | _22938_ /*4033*/;
assign _22746_ = _22930_ ^ _22937_ /*4036*/;
assign _22944_ = D[32] ^ Q[5] /*4032*/;
assign _22941_ = _22361_ & _22944_ /*4028*/;
assign _22942_ = _22361_ ^ _22944_ /*4031*/;
assign _22943_ = _22935_ & _22942_ /*4029*/;
assign _22940_ = _22941_ | _22943_ /*4027*/;
assign _22747_ = _22935_ ^ _22942_ /*4030*/;
assign _22949_ = D[33] ^ Q[5] /*4026*/;
assign _22946_ = _22362_ & _22949_ /*4022*/;
assign _22947_ = _22362_ ^ _22949_ /*4025*/;
assign _22948_ = _22940_ & _22947_ /*4023*/;
assign _22945_ = _22946_ | _22948_ /*4021*/;
assign _22748_ = _22940_ ^ _22947_ /*4024*/;
assign _22954_ = D[34] ^ Q[5] /*4020*/;
assign _22951_ = _22363_ & _22954_ /*4016*/;
assign _22952_ = _22363_ ^ _22954_ /*4019*/;
assign _22953_ = _22945_ & _22952_ /*4017*/;
assign _22950_ = _22951_ | _22953_ /*4015*/;
assign _22749_ = _22945_ ^ _22952_ /*4018*/;
assign _22959_ = D[35] ^ Q[5] /*4014*/;
assign _22956_ = _22364_ & _22959_ /*4010*/;
assign _22957_ = _22364_ ^ _22959_ /*4013*/;
assign _22958_ = _22950_ & _22957_ /*4011*/;
assign _22955_ = _22956_ | _22958_ /*4009*/;
assign _22750_ = _22950_ ^ _22957_ /*4012*/;
assign _22964_ = D[36] ^ Q[5] /*4008*/;
assign _22961_ = _22365_ & _22964_ /*4004*/;
assign _22962_ = _22365_ ^ _22964_ /*4007*/;
assign _22963_ = _22955_ & _22962_ /*4005*/;
assign _22960_ = _22961_ | _22963_ /*4003*/;
assign _22751_ = _22955_ ^ _22962_ /*4006*/;
assign _22969_ = D[37] ^ Q[5] /*4002*/;
assign _22966_ = _22366_ & _22969_ /*3998*/;
assign _22967_ = _22366_ ^ _22969_ /*4001*/;
assign _22968_ = _22960_ & _22967_ /*3999*/;
assign _22965_ = _22966_ | _22968_ /*3997*/;
assign _22752_ = _22960_ ^ _22967_ /*4000*/;
assign _22974_ = D[38] ^ Q[5] /*3996*/;
assign _22971_ = _22367_ & _22974_ /*3992*/;
assign _22972_ = _22367_ ^ _22974_ /*3995*/;
assign _22973_ = _22965_ & _22972_ /*3993*/;
assign _22970_ = _22971_ | _22973_ /*3991*/;
assign _22753_ = _22965_ ^ _22972_ /*3994*/;
assign _22979_ = D[39] ^ Q[5] /*3990*/;
assign _22976_ = _22368_ & _22979_ /*3986*/;
assign _22977_ = _22368_ ^ _22979_ /*3989*/;
assign _22978_ = _22970_ & _22977_ /*3987*/;
assign _22975_ = _22976_ | _22978_ /*3985*/;
assign _22754_ = _22970_ ^ _22977_ /*3988*/;
assign _22984_ = D[40] ^ Q[5] /*3984*/;
assign _22981_ = _22369_ & _22984_ /*3980*/;
assign _22982_ = _22369_ ^ _22984_ /*3983*/;
assign _22983_ = _22975_ & _22982_ /*3981*/;
assign _22980_ = _22981_ | _22983_ /*3979*/;
assign _22755_ = _22975_ ^ _22982_ /*3982*/;
assign _22989_ = D[41] ^ Q[5] /*3978*/;
assign _22986_ = _22370_ & _22989_ /*3974*/;
assign _22987_ = _22370_ ^ _22989_ /*3977*/;
assign _22988_ = _22980_ & _22987_ /*3975*/;
assign _22985_ = _22986_ | _22988_ /*3973*/;
assign _22756_ = _22980_ ^ _22987_ /*3976*/;
assign _22994_ = D[42] ^ Q[5] /*3972*/;
assign _22991_ = _22371_ & _22994_ /*3968*/;
assign _22992_ = _22371_ ^ _22994_ /*3971*/;
assign _22993_ = _22985_ & _22992_ /*3969*/;
assign _22990_ = _22991_ | _22993_ /*3967*/;
assign _22757_ = _22985_ ^ _22992_ /*3970*/;
assign _22999_ = D[43] ^ Q[5] /*3966*/;
assign _22996_ = _22372_ & _22999_ /*3962*/;
assign _22997_ = _22372_ ^ _22999_ /*3965*/;
assign _22998_ = _22990_ & _22997_ /*3963*/;
assign _22995_ = _22996_ | _22998_ /*3961*/;
assign _22758_ = _22990_ ^ _22997_ /*3964*/;
assign _23004_ = D[44] ^ Q[5] /*3960*/;
assign _23001_ = _22373_ & _23004_ /*3956*/;
assign _23002_ = _22373_ ^ _23004_ /*3959*/;
assign _23003_ = _22995_ & _23002_ /*3957*/;
assign _23000_ = _23001_ | _23003_ /*3955*/;
assign _22759_ = _22995_ ^ _23002_ /*3958*/;
assign _23009_ = D[45] ^ Q[5] /*3954*/;
assign _23006_ = _22374_ & _23009_ /*3950*/;
assign _23007_ = _22374_ ^ _23009_ /*3953*/;
assign _23008_ = _23000_ & _23007_ /*3951*/;
assign _23005_ = _23006_ | _23008_ /*3949*/;
assign _22760_ = _23000_ ^ _23007_ /*3952*/;
assign _23014_ = D[46] ^ Q[5] /*3948*/;
assign _23011_ = _22375_ & _23014_ /*3944*/;
assign _23012_ = _22375_ ^ _23014_ /*3947*/;
assign _23013_ = _23005_ & _23012_ /*3945*/;
assign _23010_ = _23011_ | _23013_ /*3943*/;
assign _22761_ = _23005_ ^ _23012_ /*3946*/;
assign _23019_ = D[47] ^ Q[5] /*3942*/;
assign _23016_ = _22376_ & _23019_ /*3938*/;
assign _23017_ = _22376_ ^ _23019_ /*3941*/;
assign _23018_ = _23010_ & _23017_ /*3939*/;
assign _23015_ = _23016_ | _23018_ /*3937*/;
assign _22762_ = _23010_ ^ _23017_ /*3940*/;
assign _23024_ = D[48] ^ Q[5] /*3936*/;
assign _23021_ = _22377_ & _23024_ /*3932*/;
assign _23022_ = _22377_ ^ _23024_ /*3935*/;
assign _23023_ = _23015_ & _23022_ /*3933*/;
assign _23020_ = _23021_ | _23023_ /*3931*/;
assign _22763_ = _23015_ ^ _23022_ /*3934*/;
assign _23029_ = D[49] ^ Q[5] /*3930*/;
assign _23026_ = _22378_ & _23029_ /*3926*/;
assign _23027_ = _22378_ ^ _23029_ /*3929*/;
assign _23028_ = _23020_ & _23027_ /*3927*/;
assign _23025_ = _23026_ | _23028_ /*3925*/;
assign _22764_ = _23020_ ^ _23027_ /*3928*/;
assign _23034_ = D[50] ^ Q[5] /*3924*/;
assign _23031_ = _22379_ & _23034_ /*3920*/;
assign _23032_ = _22379_ ^ _23034_ /*3923*/;
assign _23033_ = _23025_ & _23032_ /*3921*/;
assign _23030_ = _23031_ | _23033_ /*3919*/;
assign _22765_ = _23025_ ^ _23032_ /*3922*/;
assign _23039_ = D[51] ^ Q[5] /*3918*/;
assign _23036_ = _22380_ & _23039_ /*3914*/;
assign _23037_ = _22380_ ^ _23039_ /*3917*/;
assign _23038_ = _23030_ & _23037_ /*3915*/;
assign _23035_ = _23036_ | _23038_ /*3913*/;
assign _22766_ = _23030_ ^ _23037_ /*3916*/;
assign _23044_ = D[52] ^ Q[5] /*3912*/;
assign _23041_ = _22381_ & _23044_ /*3908*/;
assign _23042_ = _22381_ ^ _23044_ /*3911*/;
assign _23043_ = _23035_ & _23042_ /*3909*/;
assign _23040_ = _23041_ | _23043_ /*3907*/;
assign _22767_ = _23035_ ^ _23042_ /*3910*/;
assign _23049_ = D[53] ^ Q[5] /*3906*/;
assign _23046_ = _22382_ & _23049_ /*3902*/;
assign _23047_ = _22382_ ^ _23049_ /*3905*/;
assign _23048_ = _23040_ & _23047_ /*3903*/;
assign _23045_ = _23046_ | _23048_ /*3901*/;
assign _22768_ = _23040_ ^ _23047_ /*3904*/;
assign _23054_ = D[54] ^ Q[5] /*3900*/;
assign _23051_ = _22383_ & _23054_ /*3896*/;
assign _23052_ = _22383_ ^ _23054_ /*3899*/;
assign _23053_ = _23045_ & _23052_ /*3897*/;
assign _23050_ = _23051_ | _23053_ /*3895*/;
assign _22769_ = _23045_ ^ _23052_ /*3898*/;
assign _23059_ = D[55] ^ Q[5] /*3894*/;
assign _23056_ = _22384_ & _23059_ /*3890*/;
assign _23057_ = _22384_ ^ _23059_ /*3893*/;
assign _23058_ = _23050_ & _23057_ /*3891*/;
assign _23055_ = _23056_ | _23058_ /*3889*/;
assign _22770_ = _23050_ ^ _23057_ /*3892*/;
assign _23064_ = D[56] ^ Q[5] /*3888*/;
assign _23061_ = _22385_ & _23064_ /*3884*/;
assign _23062_ = _22385_ ^ _23064_ /*3887*/;
assign _23063_ = _23055_ & _23062_ /*3885*/;
assign _23060_ = _23061_ | _23063_ /*3883*/;
assign _22771_ = _23055_ ^ _23062_ /*3886*/;
assign _23069_ = D[57] ^ Q[5] /*3882*/;
assign _23066_ = _22386_ & _23069_ /*3878*/;
assign _23067_ = _22386_ ^ _23069_ /*3881*/;
assign _23068_ = _23060_ & _23067_ /*3879*/;
assign _23065_ = _23066_ | _23068_ /*3877*/;
assign _22772_ = _23060_ ^ _23067_ /*3880*/;
assign _23074_ = D[58] ^ Q[5] /*3876*/;
assign _23071_ = _22387_ & _23074_ /*3872*/;
assign _23072_ = _22387_ ^ _23074_ /*3875*/;
assign _23073_ = _23065_ & _23072_ /*3873*/;
assign _23070_ = _23071_ | _23073_ /*3871*/;
assign _22773_ = _23065_ ^ _23072_ /*3874*/;
assign _23079_ = D[59] ^ Q[5] /*3870*/;
assign _23076_ = _22388_ & _23079_ /*3866*/;
assign _23077_ = _22388_ ^ _23079_ /*3869*/;
assign _23078_ = _23070_ & _23077_ /*3867*/;
assign _23075_ = _23076_ | _23078_ /*3865*/;
assign _22774_ = _23070_ ^ _23077_ /*3868*/;
assign _23084_ = D[60] ^ Q[5] /*3864*/;
assign _23081_ = _22389_ & _23084_ /*3860*/;
assign _23082_ = _22389_ ^ _23084_ /*3863*/;
assign _23083_ = _23075_ & _23082_ /*3861*/;
assign _23080_ = _23081_ | _23083_ /*3859*/;
assign _22775_ = _23075_ ^ _23082_ /*3862*/;
assign _23089_ = D[61] ^ Q[5] /*3858*/;
assign _23086_ = _22390_ & _23089_ /*3854*/;
assign _23087_ = _22390_ ^ _23089_ /*3857*/;
assign _23088_ = _23080_ & _23087_ /*3855*/;
assign _23085_ = _23086_ | _23088_ /*3853*/;
assign _22776_ = _23080_ ^ _23087_ /*3856*/;
assign _23094_ = D[62] ^ Q[5] /*3852*/;
assign _23091_ = _22391_ & _23094_ /*3848*/;
assign _23092_ = _22391_ ^ _23094_ /*3851*/;
assign _23093_ = _23085_ & _23092_ /*3849*/;
assign _23090_ = _23091_ | _23093_ /*3847*/;
assign _22777_ = _23085_ ^ _23092_ /*3850*/;
assign _23098_ = zeroWire ^ Q[5] /*3846*/;
assign _23095_ = _22392_ & _23098_ /*3842*/;
assign _23096_ = _22392_ ^ _23098_ /*3845*/;
assign _23097_ = _23090_ & _23096_ /*3843*/;
assign Q[4] = _23095_ | _23097_ /*3841*/;
assign _22778_ = _23090_ ^ _23096_ /*3844*/;
assign _23169_ = D[0] ^ Q[4] /*3455*/;
assign _23166_ = R_0[3] & _23169_ /*3451*/;
assign _23167_ = R_0[3] ^ _23169_ /*3454*/;
assign _23168_ = Q[4] & _23167_ /*3452*/;
assign _23165_ = _23166_ | _23168_ /*3450*/;
assign _23100_ = Q[4] ^ _23167_ /*3453*/;
assign _23174_ = D[1] ^ Q[4] /*3449*/;
assign _23171_ = _22715_ & _23174_ /*3445*/;
assign _23172_ = _22715_ ^ _23174_ /*3448*/;
assign _23173_ = _23165_ & _23172_ /*3446*/;
assign _23170_ = _23171_ | _23173_ /*3444*/;
assign _23101_ = _23165_ ^ _23172_ /*3447*/;
assign _23179_ = D[2] ^ Q[4] /*3443*/;
assign _23176_ = _22716_ & _23179_ /*3439*/;
assign _23177_ = _22716_ ^ _23179_ /*3442*/;
assign _23178_ = _23170_ & _23177_ /*3440*/;
assign _23175_ = _23176_ | _23178_ /*3438*/;
assign _23102_ = _23170_ ^ _23177_ /*3441*/;
assign _23184_ = D[3] ^ Q[4] /*3437*/;
assign _23181_ = _22717_ & _23184_ /*3433*/;
assign _23182_ = _22717_ ^ _23184_ /*3436*/;
assign _23183_ = _23175_ & _23182_ /*3434*/;
assign _23180_ = _23181_ | _23183_ /*3432*/;
assign _23103_ = _23175_ ^ _23182_ /*3435*/;
assign _23189_ = D[4] ^ Q[4] /*3431*/;
assign _23186_ = _22718_ & _23189_ /*3427*/;
assign _23187_ = _22718_ ^ _23189_ /*3430*/;
assign _23188_ = _23180_ & _23187_ /*3428*/;
assign _23185_ = _23186_ | _23188_ /*3426*/;
assign _23104_ = _23180_ ^ _23187_ /*3429*/;
assign _23194_ = D[5] ^ Q[4] /*3425*/;
assign _23191_ = _22719_ & _23194_ /*3421*/;
assign _23192_ = _22719_ ^ _23194_ /*3424*/;
assign _23193_ = _23185_ & _23192_ /*3422*/;
assign _23190_ = _23191_ | _23193_ /*3420*/;
assign _23105_ = _23185_ ^ _23192_ /*3423*/;
assign _23199_ = D[6] ^ Q[4] /*3419*/;
assign _23196_ = _22720_ & _23199_ /*3415*/;
assign _23197_ = _22720_ ^ _23199_ /*3418*/;
assign _23198_ = _23190_ & _23197_ /*3416*/;
assign _23195_ = _23196_ | _23198_ /*3414*/;
assign _23106_ = _23190_ ^ _23197_ /*3417*/;
assign _23204_ = D[7] ^ Q[4] /*3413*/;
assign _23201_ = _22721_ & _23204_ /*3409*/;
assign _23202_ = _22721_ ^ _23204_ /*3412*/;
assign _23203_ = _23195_ & _23202_ /*3410*/;
assign _23200_ = _23201_ | _23203_ /*3408*/;
assign _23107_ = _23195_ ^ _23202_ /*3411*/;
assign _23209_ = D[8] ^ Q[4] /*3407*/;
assign _23206_ = _22722_ & _23209_ /*3403*/;
assign _23207_ = _22722_ ^ _23209_ /*3406*/;
assign _23208_ = _23200_ & _23207_ /*3404*/;
assign _23205_ = _23206_ | _23208_ /*3402*/;
assign _23108_ = _23200_ ^ _23207_ /*3405*/;
assign _23214_ = D[9] ^ Q[4] /*3401*/;
assign _23211_ = _22723_ & _23214_ /*3397*/;
assign _23212_ = _22723_ ^ _23214_ /*3400*/;
assign _23213_ = _23205_ & _23212_ /*3398*/;
assign _23210_ = _23211_ | _23213_ /*3396*/;
assign _23109_ = _23205_ ^ _23212_ /*3399*/;
assign _23219_ = D[10] ^ Q[4] /*3395*/;
assign _23216_ = _22724_ & _23219_ /*3391*/;
assign _23217_ = _22724_ ^ _23219_ /*3394*/;
assign _23218_ = _23210_ & _23217_ /*3392*/;
assign _23215_ = _23216_ | _23218_ /*3390*/;
assign _23110_ = _23210_ ^ _23217_ /*3393*/;
assign _23224_ = D[11] ^ Q[4] /*3389*/;
assign _23221_ = _22725_ & _23224_ /*3385*/;
assign _23222_ = _22725_ ^ _23224_ /*3388*/;
assign _23223_ = _23215_ & _23222_ /*3386*/;
assign _23220_ = _23221_ | _23223_ /*3384*/;
assign _23111_ = _23215_ ^ _23222_ /*3387*/;
assign _23229_ = D[12] ^ Q[4] /*3383*/;
assign _23226_ = _22726_ & _23229_ /*3379*/;
assign _23227_ = _22726_ ^ _23229_ /*3382*/;
assign _23228_ = _23220_ & _23227_ /*3380*/;
assign _23225_ = _23226_ | _23228_ /*3378*/;
assign _23112_ = _23220_ ^ _23227_ /*3381*/;
assign _23234_ = D[13] ^ Q[4] /*3377*/;
assign _23231_ = _22727_ & _23234_ /*3373*/;
assign _23232_ = _22727_ ^ _23234_ /*3376*/;
assign _23233_ = _23225_ & _23232_ /*3374*/;
assign _23230_ = _23231_ | _23233_ /*3372*/;
assign _23113_ = _23225_ ^ _23232_ /*3375*/;
assign _23239_ = D[14] ^ Q[4] /*3371*/;
assign _23236_ = _22728_ & _23239_ /*3367*/;
assign _23237_ = _22728_ ^ _23239_ /*3370*/;
assign _23238_ = _23230_ & _23237_ /*3368*/;
assign _23235_ = _23236_ | _23238_ /*3366*/;
assign _23114_ = _23230_ ^ _23237_ /*3369*/;
assign _23244_ = D[15] ^ Q[4] /*3365*/;
assign _23241_ = _22729_ & _23244_ /*3361*/;
assign _23242_ = _22729_ ^ _23244_ /*3364*/;
assign _23243_ = _23235_ & _23242_ /*3362*/;
assign _23240_ = _23241_ | _23243_ /*3360*/;
assign _23115_ = _23235_ ^ _23242_ /*3363*/;
assign _23249_ = D[16] ^ Q[4] /*3359*/;
assign _23246_ = _22730_ & _23249_ /*3355*/;
assign _23247_ = _22730_ ^ _23249_ /*3358*/;
assign _23248_ = _23240_ & _23247_ /*3356*/;
assign _23245_ = _23246_ | _23248_ /*3354*/;
assign _23116_ = _23240_ ^ _23247_ /*3357*/;
assign _23254_ = D[17] ^ Q[4] /*3353*/;
assign _23251_ = _22731_ & _23254_ /*3349*/;
assign _23252_ = _22731_ ^ _23254_ /*3352*/;
assign _23253_ = _23245_ & _23252_ /*3350*/;
assign _23250_ = _23251_ | _23253_ /*3348*/;
assign _23117_ = _23245_ ^ _23252_ /*3351*/;
assign _23259_ = D[18] ^ Q[4] /*3347*/;
assign _23256_ = _22732_ & _23259_ /*3343*/;
assign _23257_ = _22732_ ^ _23259_ /*3346*/;
assign _23258_ = _23250_ & _23257_ /*3344*/;
assign _23255_ = _23256_ | _23258_ /*3342*/;
assign _23118_ = _23250_ ^ _23257_ /*3345*/;
assign _23264_ = D[19] ^ Q[4] /*3341*/;
assign _23261_ = _22733_ & _23264_ /*3337*/;
assign _23262_ = _22733_ ^ _23264_ /*3340*/;
assign _23263_ = _23255_ & _23262_ /*3338*/;
assign _23260_ = _23261_ | _23263_ /*3336*/;
assign _23119_ = _23255_ ^ _23262_ /*3339*/;
assign _23269_ = D[20] ^ Q[4] /*3335*/;
assign _23266_ = _22734_ & _23269_ /*3331*/;
assign _23267_ = _22734_ ^ _23269_ /*3334*/;
assign _23268_ = _23260_ & _23267_ /*3332*/;
assign _23265_ = _23266_ | _23268_ /*3330*/;
assign _23120_ = _23260_ ^ _23267_ /*3333*/;
assign _23274_ = D[21] ^ Q[4] /*3329*/;
assign _23271_ = _22735_ & _23274_ /*3325*/;
assign _23272_ = _22735_ ^ _23274_ /*3328*/;
assign _23273_ = _23265_ & _23272_ /*3326*/;
assign _23270_ = _23271_ | _23273_ /*3324*/;
assign _23121_ = _23265_ ^ _23272_ /*3327*/;
assign _23279_ = D[22] ^ Q[4] /*3323*/;
assign _23276_ = _22736_ & _23279_ /*3319*/;
assign _23277_ = _22736_ ^ _23279_ /*3322*/;
assign _23278_ = _23270_ & _23277_ /*3320*/;
assign _23275_ = _23276_ | _23278_ /*3318*/;
assign _23122_ = _23270_ ^ _23277_ /*3321*/;
assign _23284_ = D[23] ^ Q[4] /*3317*/;
assign _23281_ = _22737_ & _23284_ /*3313*/;
assign _23282_ = _22737_ ^ _23284_ /*3316*/;
assign _23283_ = _23275_ & _23282_ /*3314*/;
assign _23280_ = _23281_ | _23283_ /*3312*/;
assign _23123_ = _23275_ ^ _23282_ /*3315*/;
assign _23289_ = D[24] ^ Q[4] /*3311*/;
assign _23286_ = _22738_ & _23289_ /*3307*/;
assign _23287_ = _22738_ ^ _23289_ /*3310*/;
assign _23288_ = _23280_ & _23287_ /*3308*/;
assign _23285_ = _23286_ | _23288_ /*3306*/;
assign _23124_ = _23280_ ^ _23287_ /*3309*/;
assign _23294_ = D[25] ^ Q[4] /*3305*/;
assign _23291_ = _22739_ & _23294_ /*3301*/;
assign _23292_ = _22739_ ^ _23294_ /*3304*/;
assign _23293_ = _23285_ & _23292_ /*3302*/;
assign _23290_ = _23291_ | _23293_ /*3300*/;
assign _23125_ = _23285_ ^ _23292_ /*3303*/;
assign _23299_ = D[26] ^ Q[4] /*3299*/;
assign _23296_ = _22740_ & _23299_ /*3295*/;
assign _23297_ = _22740_ ^ _23299_ /*3298*/;
assign _23298_ = _23290_ & _23297_ /*3296*/;
assign _23295_ = _23296_ | _23298_ /*3294*/;
assign _23126_ = _23290_ ^ _23297_ /*3297*/;
assign _23304_ = D[27] ^ Q[4] /*3293*/;
assign _23301_ = _22741_ & _23304_ /*3289*/;
assign _23302_ = _22741_ ^ _23304_ /*3292*/;
assign _23303_ = _23295_ & _23302_ /*3290*/;
assign _23300_ = _23301_ | _23303_ /*3288*/;
assign _23127_ = _23295_ ^ _23302_ /*3291*/;
assign _23309_ = D[28] ^ Q[4] /*3287*/;
assign _23306_ = _22742_ & _23309_ /*3283*/;
assign _23307_ = _22742_ ^ _23309_ /*3286*/;
assign _23308_ = _23300_ & _23307_ /*3284*/;
assign _23305_ = _23306_ | _23308_ /*3282*/;
assign _23128_ = _23300_ ^ _23307_ /*3285*/;
assign _23314_ = D[29] ^ Q[4] /*3281*/;
assign _23311_ = _22743_ & _23314_ /*3277*/;
assign _23312_ = _22743_ ^ _23314_ /*3280*/;
assign _23313_ = _23305_ & _23312_ /*3278*/;
assign _23310_ = _23311_ | _23313_ /*3276*/;
assign _23129_ = _23305_ ^ _23312_ /*3279*/;
assign _23319_ = D[30] ^ Q[4] /*3275*/;
assign _23316_ = _22744_ & _23319_ /*3271*/;
assign _23317_ = _22744_ ^ _23319_ /*3274*/;
assign _23318_ = _23310_ & _23317_ /*3272*/;
assign _23315_ = _23316_ | _23318_ /*3270*/;
assign _23130_ = _23310_ ^ _23317_ /*3273*/;
assign _23324_ = D[31] ^ Q[4] /*3269*/;
assign _23321_ = _22745_ & _23324_ /*3265*/;
assign _23322_ = _22745_ ^ _23324_ /*3268*/;
assign _23323_ = _23315_ & _23322_ /*3266*/;
assign _23320_ = _23321_ | _23323_ /*3264*/;
assign _23131_ = _23315_ ^ _23322_ /*3267*/;
assign _23329_ = D[32] ^ Q[4] /*3263*/;
assign _23326_ = _22746_ & _23329_ /*3259*/;
assign _23327_ = _22746_ ^ _23329_ /*3262*/;
assign _23328_ = _23320_ & _23327_ /*3260*/;
assign _23325_ = _23326_ | _23328_ /*3258*/;
assign _23132_ = _23320_ ^ _23327_ /*3261*/;
assign _23334_ = D[33] ^ Q[4] /*3257*/;
assign _23331_ = _22747_ & _23334_ /*3253*/;
assign _23332_ = _22747_ ^ _23334_ /*3256*/;
assign _23333_ = _23325_ & _23332_ /*3254*/;
assign _23330_ = _23331_ | _23333_ /*3252*/;
assign _23133_ = _23325_ ^ _23332_ /*3255*/;
assign _23339_ = D[34] ^ Q[4] /*3251*/;
assign _23336_ = _22748_ & _23339_ /*3247*/;
assign _23337_ = _22748_ ^ _23339_ /*3250*/;
assign _23338_ = _23330_ & _23337_ /*3248*/;
assign _23335_ = _23336_ | _23338_ /*3246*/;
assign _23134_ = _23330_ ^ _23337_ /*3249*/;
assign _23344_ = D[35] ^ Q[4] /*3245*/;
assign _23341_ = _22749_ & _23344_ /*3241*/;
assign _23342_ = _22749_ ^ _23344_ /*3244*/;
assign _23343_ = _23335_ & _23342_ /*3242*/;
assign _23340_ = _23341_ | _23343_ /*3240*/;
assign _23135_ = _23335_ ^ _23342_ /*3243*/;
assign _23349_ = D[36] ^ Q[4] /*3239*/;
assign _23346_ = _22750_ & _23349_ /*3235*/;
assign _23347_ = _22750_ ^ _23349_ /*3238*/;
assign _23348_ = _23340_ & _23347_ /*3236*/;
assign _23345_ = _23346_ | _23348_ /*3234*/;
assign _23136_ = _23340_ ^ _23347_ /*3237*/;
assign _23354_ = D[37] ^ Q[4] /*3233*/;
assign _23351_ = _22751_ & _23354_ /*3229*/;
assign _23352_ = _22751_ ^ _23354_ /*3232*/;
assign _23353_ = _23345_ & _23352_ /*3230*/;
assign _23350_ = _23351_ | _23353_ /*3228*/;
assign _23137_ = _23345_ ^ _23352_ /*3231*/;
assign _23359_ = D[38] ^ Q[4] /*3227*/;
assign _23356_ = _22752_ & _23359_ /*3223*/;
assign _23357_ = _22752_ ^ _23359_ /*3226*/;
assign _23358_ = _23350_ & _23357_ /*3224*/;
assign _23355_ = _23356_ | _23358_ /*3222*/;
assign _23138_ = _23350_ ^ _23357_ /*3225*/;
assign _23364_ = D[39] ^ Q[4] /*3221*/;
assign _23361_ = _22753_ & _23364_ /*3217*/;
assign _23362_ = _22753_ ^ _23364_ /*3220*/;
assign _23363_ = _23355_ & _23362_ /*3218*/;
assign _23360_ = _23361_ | _23363_ /*3216*/;
assign _23139_ = _23355_ ^ _23362_ /*3219*/;
assign _23369_ = D[40] ^ Q[4] /*3215*/;
assign _23366_ = _22754_ & _23369_ /*3211*/;
assign _23367_ = _22754_ ^ _23369_ /*3214*/;
assign _23368_ = _23360_ & _23367_ /*3212*/;
assign _23365_ = _23366_ | _23368_ /*3210*/;
assign _23140_ = _23360_ ^ _23367_ /*3213*/;
assign _23374_ = D[41] ^ Q[4] /*3209*/;
assign _23371_ = _22755_ & _23374_ /*3205*/;
assign _23372_ = _22755_ ^ _23374_ /*3208*/;
assign _23373_ = _23365_ & _23372_ /*3206*/;
assign _23370_ = _23371_ | _23373_ /*3204*/;
assign _23141_ = _23365_ ^ _23372_ /*3207*/;
assign _23379_ = D[42] ^ Q[4] /*3203*/;
assign _23376_ = _22756_ & _23379_ /*3199*/;
assign _23377_ = _22756_ ^ _23379_ /*3202*/;
assign _23378_ = _23370_ & _23377_ /*3200*/;
assign _23375_ = _23376_ | _23378_ /*3198*/;
assign _23142_ = _23370_ ^ _23377_ /*3201*/;
assign _23384_ = D[43] ^ Q[4] /*3197*/;
assign _23381_ = _22757_ & _23384_ /*3193*/;
assign _23382_ = _22757_ ^ _23384_ /*3196*/;
assign _23383_ = _23375_ & _23382_ /*3194*/;
assign _23380_ = _23381_ | _23383_ /*3192*/;
assign _23143_ = _23375_ ^ _23382_ /*3195*/;
assign _23389_ = D[44] ^ Q[4] /*3191*/;
assign _23386_ = _22758_ & _23389_ /*3187*/;
assign _23387_ = _22758_ ^ _23389_ /*3190*/;
assign _23388_ = _23380_ & _23387_ /*3188*/;
assign _23385_ = _23386_ | _23388_ /*3186*/;
assign _23144_ = _23380_ ^ _23387_ /*3189*/;
assign _23394_ = D[45] ^ Q[4] /*3185*/;
assign _23391_ = _22759_ & _23394_ /*3181*/;
assign _23392_ = _22759_ ^ _23394_ /*3184*/;
assign _23393_ = _23385_ & _23392_ /*3182*/;
assign _23390_ = _23391_ | _23393_ /*3180*/;
assign _23145_ = _23385_ ^ _23392_ /*3183*/;
assign _23399_ = D[46] ^ Q[4] /*3179*/;
assign _23396_ = _22760_ & _23399_ /*3175*/;
assign _23397_ = _22760_ ^ _23399_ /*3178*/;
assign _23398_ = _23390_ & _23397_ /*3176*/;
assign _23395_ = _23396_ | _23398_ /*3174*/;
assign _23146_ = _23390_ ^ _23397_ /*3177*/;
assign _23404_ = D[47] ^ Q[4] /*3173*/;
assign _23401_ = _22761_ & _23404_ /*3169*/;
assign _23402_ = _22761_ ^ _23404_ /*3172*/;
assign _23403_ = _23395_ & _23402_ /*3170*/;
assign _23400_ = _23401_ | _23403_ /*3168*/;
assign _23147_ = _23395_ ^ _23402_ /*3171*/;
assign _23409_ = D[48] ^ Q[4] /*3167*/;
assign _23406_ = _22762_ & _23409_ /*3163*/;
assign _23407_ = _22762_ ^ _23409_ /*3166*/;
assign _23408_ = _23400_ & _23407_ /*3164*/;
assign _23405_ = _23406_ | _23408_ /*3162*/;
assign _23148_ = _23400_ ^ _23407_ /*3165*/;
assign _23414_ = D[49] ^ Q[4] /*3161*/;
assign _23411_ = _22763_ & _23414_ /*3157*/;
assign _23412_ = _22763_ ^ _23414_ /*3160*/;
assign _23413_ = _23405_ & _23412_ /*3158*/;
assign _23410_ = _23411_ | _23413_ /*3156*/;
assign _23149_ = _23405_ ^ _23412_ /*3159*/;
assign _23419_ = D[50] ^ Q[4] /*3155*/;
assign _23416_ = _22764_ & _23419_ /*3151*/;
assign _23417_ = _22764_ ^ _23419_ /*3154*/;
assign _23418_ = _23410_ & _23417_ /*3152*/;
assign _23415_ = _23416_ | _23418_ /*3150*/;
assign _23150_ = _23410_ ^ _23417_ /*3153*/;
assign _23424_ = D[51] ^ Q[4] /*3149*/;
assign _23421_ = _22765_ & _23424_ /*3145*/;
assign _23422_ = _22765_ ^ _23424_ /*3148*/;
assign _23423_ = _23415_ & _23422_ /*3146*/;
assign _23420_ = _23421_ | _23423_ /*3144*/;
assign _23151_ = _23415_ ^ _23422_ /*3147*/;
assign _23429_ = D[52] ^ Q[4] /*3143*/;
assign _23426_ = _22766_ & _23429_ /*3139*/;
assign _23427_ = _22766_ ^ _23429_ /*3142*/;
assign _23428_ = _23420_ & _23427_ /*3140*/;
assign _23425_ = _23426_ | _23428_ /*3138*/;
assign _23152_ = _23420_ ^ _23427_ /*3141*/;
assign _23434_ = D[53] ^ Q[4] /*3137*/;
assign _23431_ = _22767_ & _23434_ /*3133*/;
assign _23432_ = _22767_ ^ _23434_ /*3136*/;
assign _23433_ = _23425_ & _23432_ /*3134*/;
assign _23430_ = _23431_ | _23433_ /*3132*/;
assign _23153_ = _23425_ ^ _23432_ /*3135*/;
assign _23439_ = D[54] ^ Q[4] /*3131*/;
assign _23436_ = _22768_ & _23439_ /*3127*/;
assign _23437_ = _22768_ ^ _23439_ /*3130*/;
assign _23438_ = _23430_ & _23437_ /*3128*/;
assign _23435_ = _23436_ | _23438_ /*3126*/;
assign _23154_ = _23430_ ^ _23437_ /*3129*/;
assign _23444_ = D[55] ^ Q[4] /*3125*/;
assign _23441_ = _22769_ & _23444_ /*3121*/;
assign _23442_ = _22769_ ^ _23444_ /*3124*/;
assign _23443_ = _23435_ & _23442_ /*3122*/;
assign _23440_ = _23441_ | _23443_ /*3120*/;
assign _23155_ = _23435_ ^ _23442_ /*3123*/;
assign _23449_ = D[56] ^ Q[4] /*3119*/;
assign _23446_ = _22770_ & _23449_ /*3115*/;
assign _23447_ = _22770_ ^ _23449_ /*3118*/;
assign _23448_ = _23440_ & _23447_ /*3116*/;
assign _23445_ = _23446_ | _23448_ /*3114*/;
assign _23156_ = _23440_ ^ _23447_ /*3117*/;
assign _23454_ = D[57] ^ Q[4] /*3113*/;
assign _23451_ = _22771_ & _23454_ /*3109*/;
assign _23452_ = _22771_ ^ _23454_ /*3112*/;
assign _23453_ = _23445_ & _23452_ /*3110*/;
assign _23450_ = _23451_ | _23453_ /*3108*/;
assign _23157_ = _23445_ ^ _23452_ /*3111*/;
assign _23459_ = D[58] ^ Q[4] /*3107*/;
assign _23456_ = _22772_ & _23459_ /*3103*/;
assign _23457_ = _22772_ ^ _23459_ /*3106*/;
assign _23458_ = _23450_ & _23457_ /*3104*/;
assign _23455_ = _23456_ | _23458_ /*3102*/;
assign _23158_ = _23450_ ^ _23457_ /*3105*/;
assign _23464_ = D[59] ^ Q[4] /*3101*/;
assign _23461_ = _22773_ & _23464_ /*3097*/;
assign _23462_ = _22773_ ^ _23464_ /*3100*/;
assign _23463_ = _23455_ & _23462_ /*3098*/;
assign _23460_ = _23461_ | _23463_ /*3096*/;
assign _23159_ = _23455_ ^ _23462_ /*3099*/;
assign _23469_ = D[60] ^ Q[4] /*3095*/;
assign _23466_ = _22774_ & _23469_ /*3091*/;
assign _23467_ = _22774_ ^ _23469_ /*3094*/;
assign _23468_ = _23460_ & _23467_ /*3092*/;
assign _23465_ = _23466_ | _23468_ /*3090*/;
assign _23160_ = _23460_ ^ _23467_ /*3093*/;
assign _23474_ = D[61] ^ Q[4] /*3089*/;
assign _23471_ = _22775_ & _23474_ /*3085*/;
assign _23472_ = _22775_ ^ _23474_ /*3088*/;
assign _23473_ = _23465_ & _23472_ /*3086*/;
assign _23470_ = _23471_ | _23473_ /*3084*/;
assign _23161_ = _23465_ ^ _23472_ /*3087*/;
assign _23479_ = D[62] ^ Q[4] /*3083*/;
assign _23476_ = _22776_ & _23479_ /*3079*/;
assign _23477_ = _22776_ ^ _23479_ /*3082*/;
assign _23478_ = _23470_ & _23477_ /*3080*/;
assign _23475_ = _23476_ | _23478_ /*3078*/;
assign _23162_ = _23470_ ^ _23477_ /*3081*/;
assign _23483_ = zeroWire ^ Q[4] /*3077*/;
assign _23480_ = _22777_ & _23483_ /*3073*/;
assign _23481_ = _22777_ ^ _23483_ /*3076*/;
assign _23482_ = _23475_ & _23481_ /*3074*/;
assign Q[3] = _23480_ | _23482_ /*3072*/;
assign _23163_ = _23475_ ^ _23481_ /*3075*/;
assign _23554_ = D[0] ^ Q[3] /*2686*/;
assign _23551_ = R_0[2] & _23554_ /*2682*/;
assign _23552_ = R_0[2] ^ _23554_ /*2685*/;
assign _23553_ = Q[3] & _23552_ /*2683*/;
assign _23550_ = _23551_ | _23553_ /*2681*/;
assign _23485_ = Q[3] ^ _23552_ /*2684*/;
assign _23559_ = D[1] ^ Q[3] /*2680*/;
assign _23556_ = _23100_ & _23559_ /*2676*/;
assign _23557_ = _23100_ ^ _23559_ /*2679*/;
assign _23558_ = _23550_ & _23557_ /*2677*/;
assign _23555_ = _23556_ | _23558_ /*2675*/;
assign _23486_ = _23550_ ^ _23557_ /*2678*/;
assign _23564_ = D[2] ^ Q[3] /*2674*/;
assign _23561_ = _23101_ & _23564_ /*2670*/;
assign _23562_ = _23101_ ^ _23564_ /*2673*/;
assign _23563_ = _23555_ & _23562_ /*2671*/;
assign _23560_ = _23561_ | _23563_ /*2669*/;
assign _23487_ = _23555_ ^ _23562_ /*2672*/;
assign _23569_ = D[3] ^ Q[3] /*2668*/;
assign _23566_ = _23102_ & _23569_ /*2664*/;
assign _23567_ = _23102_ ^ _23569_ /*2667*/;
assign _23568_ = _23560_ & _23567_ /*2665*/;
assign _23565_ = _23566_ | _23568_ /*2663*/;
assign _23488_ = _23560_ ^ _23567_ /*2666*/;
assign _23574_ = D[4] ^ Q[3] /*2662*/;
assign _23571_ = _23103_ & _23574_ /*2658*/;
assign _23572_ = _23103_ ^ _23574_ /*2661*/;
assign _23573_ = _23565_ & _23572_ /*2659*/;
assign _23570_ = _23571_ | _23573_ /*2657*/;
assign _23489_ = _23565_ ^ _23572_ /*2660*/;
assign _23579_ = D[5] ^ Q[3] /*2656*/;
assign _23576_ = _23104_ & _23579_ /*2652*/;
assign _23577_ = _23104_ ^ _23579_ /*2655*/;
assign _23578_ = _23570_ & _23577_ /*2653*/;
assign _23575_ = _23576_ | _23578_ /*2651*/;
assign _23490_ = _23570_ ^ _23577_ /*2654*/;
assign _23584_ = D[6] ^ Q[3] /*2650*/;
assign _23581_ = _23105_ & _23584_ /*2646*/;
assign _23582_ = _23105_ ^ _23584_ /*2649*/;
assign _23583_ = _23575_ & _23582_ /*2647*/;
assign _23580_ = _23581_ | _23583_ /*2645*/;
assign _23491_ = _23575_ ^ _23582_ /*2648*/;
assign _23589_ = D[7] ^ Q[3] /*2644*/;
assign _23586_ = _23106_ & _23589_ /*2640*/;
assign _23587_ = _23106_ ^ _23589_ /*2643*/;
assign _23588_ = _23580_ & _23587_ /*2641*/;
assign _23585_ = _23586_ | _23588_ /*2639*/;
assign _23492_ = _23580_ ^ _23587_ /*2642*/;
assign _23594_ = D[8] ^ Q[3] /*2638*/;
assign _23591_ = _23107_ & _23594_ /*2634*/;
assign _23592_ = _23107_ ^ _23594_ /*2637*/;
assign _23593_ = _23585_ & _23592_ /*2635*/;
assign _23590_ = _23591_ | _23593_ /*2633*/;
assign _23493_ = _23585_ ^ _23592_ /*2636*/;
assign _23599_ = D[9] ^ Q[3] /*2632*/;
assign _23596_ = _23108_ & _23599_ /*2628*/;
assign _23597_ = _23108_ ^ _23599_ /*2631*/;
assign _23598_ = _23590_ & _23597_ /*2629*/;
assign _23595_ = _23596_ | _23598_ /*2627*/;
assign _23494_ = _23590_ ^ _23597_ /*2630*/;
assign _23604_ = D[10] ^ Q[3] /*2626*/;
assign _23601_ = _23109_ & _23604_ /*2622*/;
assign _23602_ = _23109_ ^ _23604_ /*2625*/;
assign _23603_ = _23595_ & _23602_ /*2623*/;
assign _23600_ = _23601_ | _23603_ /*2621*/;
assign _23495_ = _23595_ ^ _23602_ /*2624*/;
assign _23609_ = D[11] ^ Q[3] /*2620*/;
assign _23606_ = _23110_ & _23609_ /*2616*/;
assign _23607_ = _23110_ ^ _23609_ /*2619*/;
assign _23608_ = _23600_ & _23607_ /*2617*/;
assign _23605_ = _23606_ | _23608_ /*2615*/;
assign _23496_ = _23600_ ^ _23607_ /*2618*/;
assign _23614_ = D[12] ^ Q[3] /*2614*/;
assign _23611_ = _23111_ & _23614_ /*2610*/;
assign _23612_ = _23111_ ^ _23614_ /*2613*/;
assign _23613_ = _23605_ & _23612_ /*2611*/;
assign _23610_ = _23611_ | _23613_ /*2609*/;
assign _23497_ = _23605_ ^ _23612_ /*2612*/;
assign _23619_ = D[13] ^ Q[3] /*2608*/;
assign _23616_ = _23112_ & _23619_ /*2604*/;
assign _23617_ = _23112_ ^ _23619_ /*2607*/;
assign _23618_ = _23610_ & _23617_ /*2605*/;
assign _23615_ = _23616_ | _23618_ /*2603*/;
assign _23498_ = _23610_ ^ _23617_ /*2606*/;
assign _23624_ = D[14] ^ Q[3] /*2602*/;
assign _23621_ = _23113_ & _23624_ /*2598*/;
assign _23622_ = _23113_ ^ _23624_ /*2601*/;
assign _23623_ = _23615_ & _23622_ /*2599*/;
assign _23620_ = _23621_ | _23623_ /*2597*/;
assign _23499_ = _23615_ ^ _23622_ /*2600*/;
assign _23629_ = D[15] ^ Q[3] /*2596*/;
assign _23626_ = _23114_ & _23629_ /*2592*/;
assign _23627_ = _23114_ ^ _23629_ /*2595*/;
assign _23628_ = _23620_ & _23627_ /*2593*/;
assign _23625_ = _23626_ | _23628_ /*2591*/;
assign _23500_ = _23620_ ^ _23627_ /*2594*/;
assign _23634_ = D[16] ^ Q[3] /*2590*/;
assign _23631_ = _23115_ & _23634_ /*2586*/;
assign _23632_ = _23115_ ^ _23634_ /*2589*/;
assign _23633_ = _23625_ & _23632_ /*2587*/;
assign _23630_ = _23631_ | _23633_ /*2585*/;
assign _23501_ = _23625_ ^ _23632_ /*2588*/;
assign _23639_ = D[17] ^ Q[3] /*2584*/;
assign _23636_ = _23116_ & _23639_ /*2580*/;
assign _23637_ = _23116_ ^ _23639_ /*2583*/;
assign _23638_ = _23630_ & _23637_ /*2581*/;
assign _23635_ = _23636_ | _23638_ /*2579*/;
assign _23502_ = _23630_ ^ _23637_ /*2582*/;
assign _23644_ = D[18] ^ Q[3] /*2578*/;
assign _23641_ = _23117_ & _23644_ /*2574*/;
assign _23642_ = _23117_ ^ _23644_ /*2577*/;
assign _23643_ = _23635_ & _23642_ /*2575*/;
assign _23640_ = _23641_ | _23643_ /*2573*/;
assign _23503_ = _23635_ ^ _23642_ /*2576*/;
assign _23649_ = D[19] ^ Q[3] /*2572*/;
assign _23646_ = _23118_ & _23649_ /*2568*/;
assign _23647_ = _23118_ ^ _23649_ /*2571*/;
assign _23648_ = _23640_ & _23647_ /*2569*/;
assign _23645_ = _23646_ | _23648_ /*2567*/;
assign _23504_ = _23640_ ^ _23647_ /*2570*/;
assign _23654_ = D[20] ^ Q[3] /*2566*/;
assign _23651_ = _23119_ & _23654_ /*2562*/;
assign _23652_ = _23119_ ^ _23654_ /*2565*/;
assign _23653_ = _23645_ & _23652_ /*2563*/;
assign _23650_ = _23651_ | _23653_ /*2561*/;
assign _23505_ = _23645_ ^ _23652_ /*2564*/;
assign _23659_ = D[21] ^ Q[3] /*2560*/;
assign _23656_ = _23120_ & _23659_ /*2556*/;
assign _23657_ = _23120_ ^ _23659_ /*2559*/;
assign _23658_ = _23650_ & _23657_ /*2557*/;
assign _23655_ = _23656_ | _23658_ /*2555*/;
assign _23506_ = _23650_ ^ _23657_ /*2558*/;
assign _23664_ = D[22] ^ Q[3] /*2554*/;
assign _23661_ = _23121_ & _23664_ /*2550*/;
assign _23662_ = _23121_ ^ _23664_ /*2553*/;
assign _23663_ = _23655_ & _23662_ /*2551*/;
assign _23660_ = _23661_ | _23663_ /*2549*/;
assign _23507_ = _23655_ ^ _23662_ /*2552*/;
assign _23669_ = D[23] ^ Q[3] /*2548*/;
assign _23666_ = _23122_ & _23669_ /*2544*/;
assign _23667_ = _23122_ ^ _23669_ /*2547*/;
assign _23668_ = _23660_ & _23667_ /*2545*/;
assign _23665_ = _23666_ | _23668_ /*2543*/;
assign _23508_ = _23660_ ^ _23667_ /*2546*/;
assign _23674_ = D[24] ^ Q[3] /*2542*/;
assign _23671_ = _23123_ & _23674_ /*2538*/;
assign _23672_ = _23123_ ^ _23674_ /*2541*/;
assign _23673_ = _23665_ & _23672_ /*2539*/;
assign _23670_ = _23671_ | _23673_ /*2537*/;
assign _23509_ = _23665_ ^ _23672_ /*2540*/;
assign _23679_ = D[25] ^ Q[3] /*2536*/;
assign _23676_ = _23124_ & _23679_ /*2532*/;
assign _23677_ = _23124_ ^ _23679_ /*2535*/;
assign _23678_ = _23670_ & _23677_ /*2533*/;
assign _23675_ = _23676_ | _23678_ /*2531*/;
assign _23510_ = _23670_ ^ _23677_ /*2534*/;
assign _23684_ = D[26] ^ Q[3] /*2530*/;
assign _23681_ = _23125_ & _23684_ /*2526*/;
assign _23682_ = _23125_ ^ _23684_ /*2529*/;
assign _23683_ = _23675_ & _23682_ /*2527*/;
assign _23680_ = _23681_ | _23683_ /*2525*/;
assign _23511_ = _23675_ ^ _23682_ /*2528*/;
assign _23689_ = D[27] ^ Q[3] /*2524*/;
assign _23686_ = _23126_ & _23689_ /*2520*/;
assign _23687_ = _23126_ ^ _23689_ /*2523*/;
assign _23688_ = _23680_ & _23687_ /*2521*/;
assign _23685_ = _23686_ | _23688_ /*2519*/;
assign _23512_ = _23680_ ^ _23687_ /*2522*/;
assign _23694_ = D[28] ^ Q[3] /*2518*/;
assign _23691_ = _23127_ & _23694_ /*2514*/;
assign _23692_ = _23127_ ^ _23694_ /*2517*/;
assign _23693_ = _23685_ & _23692_ /*2515*/;
assign _23690_ = _23691_ | _23693_ /*2513*/;
assign _23513_ = _23685_ ^ _23692_ /*2516*/;
assign _23699_ = D[29] ^ Q[3] /*2512*/;
assign _23696_ = _23128_ & _23699_ /*2508*/;
assign _23697_ = _23128_ ^ _23699_ /*2511*/;
assign _23698_ = _23690_ & _23697_ /*2509*/;
assign _23695_ = _23696_ | _23698_ /*2507*/;
assign _23514_ = _23690_ ^ _23697_ /*2510*/;
assign _23704_ = D[30] ^ Q[3] /*2506*/;
assign _23701_ = _23129_ & _23704_ /*2502*/;
assign _23702_ = _23129_ ^ _23704_ /*2505*/;
assign _23703_ = _23695_ & _23702_ /*2503*/;
assign _23700_ = _23701_ | _23703_ /*2501*/;
assign _23515_ = _23695_ ^ _23702_ /*2504*/;
assign _23709_ = D[31] ^ Q[3] /*2500*/;
assign _23706_ = _23130_ & _23709_ /*2496*/;
assign _23707_ = _23130_ ^ _23709_ /*2499*/;
assign _23708_ = _23700_ & _23707_ /*2497*/;
assign _23705_ = _23706_ | _23708_ /*2495*/;
assign _23516_ = _23700_ ^ _23707_ /*2498*/;
assign _23714_ = D[32] ^ Q[3] /*2494*/;
assign _23711_ = _23131_ & _23714_ /*2490*/;
assign _23712_ = _23131_ ^ _23714_ /*2493*/;
assign _23713_ = _23705_ & _23712_ /*2491*/;
assign _23710_ = _23711_ | _23713_ /*2489*/;
assign _23517_ = _23705_ ^ _23712_ /*2492*/;
assign _23719_ = D[33] ^ Q[3] /*2488*/;
assign _23716_ = _23132_ & _23719_ /*2484*/;
assign _23717_ = _23132_ ^ _23719_ /*2487*/;
assign _23718_ = _23710_ & _23717_ /*2485*/;
assign _23715_ = _23716_ | _23718_ /*2483*/;
assign _23518_ = _23710_ ^ _23717_ /*2486*/;
assign _23724_ = D[34] ^ Q[3] /*2482*/;
assign _23721_ = _23133_ & _23724_ /*2478*/;
assign _23722_ = _23133_ ^ _23724_ /*2481*/;
assign _23723_ = _23715_ & _23722_ /*2479*/;
assign _23720_ = _23721_ | _23723_ /*2477*/;
assign _23519_ = _23715_ ^ _23722_ /*2480*/;
assign _23729_ = D[35] ^ Q[3] /*2476*/;
assign _23726_ = _23134_ & _23729_ /*2472*/;
assign _23727_ = _23134_ ^ _23729_ /*2475*/;
assign _23728_ = _23720_ & _23727_ /*2473*/;
assign _23725_ = _23726_ | _23728_ /*2471*/;
assign _23520_ = _23720_ ^ _23727_ /*2474*/;
assign _23734_ = D[36] ^ Q[3] /*2470*/;
assign _23731_ = _23135_ & _23734_ /*2466*/;
assign _23732_ = _23135_ ^ _23734_ /*2469*/;
assign _23733_ = _23725_ & _23732_ /*2467*/;
assign _23730_ = _23731_ | _23733_ /*2465*/;
assign _23521_ = _23725_ ^ _23732_ /*2468*/;
assign _23739_ = D[37] ^ Q[3] /*2464*/;
assign _23736_ = _23136_ & _23739_ /*2460*/;
assign _23737_ = _23136_ ^ _23739_ /*2463*/;
assign _23738_ = _23730_ & _23737_ /*2461*/;
assign _23735_ = _23736_ | _23738_ /*2459*/;
assign _23522_ = _23730_ ^ _23737_ /*2462*/;
assign _23744_ = D[38] ^ Q[3] /*2458*/;
assign _23741_ = _23137_ & _23744_ /*2454*/;
assign _23742_ = _23137_ ^ _23744_ /*2457*/;
assign _23743_ = _23735_ & _23742_ /*2455*/;
assign _23740_ = _23741_ | _23743_ /*2453*/;
assign _23523_ = _23735_ ^ _23742_ /*2456*/;
assign _23749_ = D[39] ^ Q[3] /*2452*/;
assign _23746_ = _23138_ & _23749_ /*2448*/;
assign _23747_ = _23138_ ^ _23749_ /*2451*/;
assign _23748_ = _23740_ & _23747_ /*2449*/;
assign _23745_ = _23746_ | _23748_ /*2447*/;
assign _23524_ = _23740_ ^ _23747_ /*2450*/;
assign _23754_ = D[40] ^ Q[3] /*2446*/;
assign _23751_ = _23139_ & _23754_ /*2442*/;
assign _23752_ = _23139_ ^ _23754_ /*2445*/;
assign _23753_ = _23745_ & _23752_ /*2443*/;
assign _23750_ = _23751_ | _23753_ /*2441*/;
assign _23525_ = _23745_ ^ _23752_ /*2444*/;
assign _23759_ = D[41] ^ Q[3] /*2440*/;
assign _23756_ = _23140_ & _23759_ /*2436*/;
assign _23757_ = _23140_ ^ _23759_ /*2439*/;
assign _23758_ = _23750_ & _23757_ /*2437*/;
assign _23755_ = _23756_ | _23758_ /*2435*/;
assign _23526_ = _23750_ ^ _23757_ /*2438*/;
assign _23764_ = D[42] ^ Q[3] /*2434*/;
assign _23761_ = _23141_ & _23764_ /*2430*/;
assign _23762_ = _23141_ ^ _23764_ /*2433*/;
assign _23763_ = _23755_ & _23762_ /*2431*/;
assign _23760_ = _23761_ | _23763_ /*2429*/;
assign _23527_ = _23755_ ^ _23762_ /*2432*/;
assign _23769_ = D[43] ^ Q[3] /*2428*/;
assign _23766_ = _23142_ & _23769_ /*2424*/;
assign _23767_ = _23142_ ^ _23769_ /*2427*/;
assign _23768_ = _23760_ & _23767_ /*2425*/;
assign _23765_ = _23766_ | _23768_ /*2423*/;
assign _23528_ = _23760_ ^ _23767_ /*2426*/;
assign _23774_ = D[44] ^ Q[3] /*2422*/;
assign _23771_ = _23143_ & _23774_ /*2418*/;
assign _23772_ = _23143_ ^ _23774_ /*2421*/;
assign _23773_ = _23765_ & _23772_ /*2419*/;
assign _23770_ = _23771_ | _23773_ /*2417*/;
assign _23529_ = _23765_ ^ _23772_ /*2420*/;
assign _23779_ = D[45] ^ Q[3] /*2416*/;
assign _23776_ = _23144_ & _23779_ /*2412*/;
assign _23777_ = _23144_ ^ _23779_ /*2415*/;
assign _23778_ = _23770_ & _23777_ /*2413*/;
assign _23775_ = _23776_ | _23778_ /*2411*/;
assign _23530_ = _23770_ ^ _23777_ /*2414*/;
assign _23784_ = D[46] ^ Q[3] /*2410*/;
assign _23781_ = _23145_ & _23784_ /*2406*/;
assign _23782_ = _23145_ ^ _23784_ /*2409*/;
assign _23783_ = _23775_ & _23782_ /*2407*/;
assign _23780_ = _23781_ | _23783_ /*2405*/;
assign _23531_ = _23775_ ^ _23782_ /*2408*/;
assign _23789_ = D[47] ^ Q[3] /*2404*/;
assign _23786_ = _23146_ & _23789_ /*2400*/;
assign _23787_ = _23146_ ^ _23789_ /*2403*/;
assign _23788_ = _23780_ & _23787_ /*2401*/;
assign _23785_ = _23786_ | _23788_ /*2399*/;
assign _23532_ = _23780_ ^ _23787_ /*2402*/;
assign _23794_ = D[48] ^ Q[3] /*2398*/;
assign _23791_ = _23147_ & _23794_ /*2394*/;
assign _23792_ = _23147_ ^ _23794_ /*2397*/;
assign _23793_ = _23785_ & _23792_ /*2395*/;
assign _23790_ = _23791_ | _23793_ /*2393*/;
assign _23533_ = _23785_ ^ _23792_ /*2396*/;
assign _23799_ = D[49] ^ Q[3] /*2392*/;
assign _23796_ = _23148_ & _23799_ /*2388*/;
assign _23797_ = _23148_ ^ _23799_ /*2391*/;
assign _23798_ = _23790_ & _23797_ /*2389*/;
assign _23795_ = _23796_ | _23798_ /*2387*/;
assign _23534_ = _23790_ ^ _23797_ /*2390*/;
assign _23804_ = D[50] ^ Q[3] /*2386*/;
assign _23801_ = _23149_ & _23804_ /*2382*/;
assign _23802_ = _23149_ ^ _23804_ /*2385*/;
assign _23803_ = _23795_ & _23802_ /*2383*/;
assign _23800_ = _23801_ | _23803_ /*2381*/;
assign _23535_ = _23795_ ^ _23802_ /*2384*/;
assign _23809_ = D[51] ^ Q[3] /*2380*/;
assign _23806_ = _23150_ & _23809_ /*2376*/;
assign _23807_ = _23150_ ^ _23809_ /*2379*/;
assign _23808_ = _23800_ & _23807_ /*2377*/;
assign _23805_ = _23806_ | _23808_ /*2375*/;
assign _23536_ = _23800_ ^ _23807_ /*2378*/;
assign _23814_ = D[52] ^ Q[3] /*2374*/;
assign _23811_ = _23151_ & _23814_ /*2370*/;
assign _23812_ = _23151_ ^ _23814_ /*2373*/;
assign _23813_ = _23805_ & _23812_ /*2371*/;
assign _23810_ = _23811_ | _23813_ /*2369*/;
assign _23537_ = _23805_ ^ _23812_ /*2372*/;
assign _23819_ = D[53] ^ Q[3] /*2368*/;
assign _23816_ = _23152_ & _23819_ /*2364*/;
assign _23817_ = _23152_ ^ _23819_ /*2367*/;
assign _23818_ = _23810_ & _23817_ /*2365*/;
assign _23815_ = _23816_ | _23818_ /*2363*/;
assign _23538_ = _23810_ ^ _23817_ /*2366*/;
assign _23824_ = D[54] ^ Q[3] /*2362*/;
assign _23821_ = _23153_ & _23824_ /*2358*/;
assign _23822_ = _23153_ ^ _23824_ /*2361*/;
assign _23823_ = _23815_ & _23822_ /*2359*/;
assign _23820_ = _23821_ | _23823_ /*2357*/;
assign _23539_ = _23815_ ^ _23822_ /*2360*/;
assign _23829_ = D[55] ^ Q[3] /*2356*/;
assign _23826_ = _23154_ & _23829_ /*2352*/;
assign _23827_ = _23154_ ^ _23829_ /*2355*/;
assign _23828_ = _23820_ & _23827_ /*2353*/;
assign _23825_ = _23826_ | _23828_ /*2351*/;
assign _23540_ = _23820_ ^ _23827_ /*2354*/;
assign _23834_ = D[56] ^ Q[3] /*2350*/;
assign _23831_ = _23155_ & _23834_ /*2346*/;
assign _23832_ = _23155_ ^ _23834_ /*2349*/;
assign _23833_ = _23825_ & _23832_ /*2347*/;
assign _23830_ = _23831_ | _23833_ /*2345*/;
assign _23541_ = _23825_ ^ _23832_ /*2348*/;
assign _23839_ = D[57] ^ Q[3] /*2344*/;
assign _23836_ = _23156_ & _23839_ /*2340*/;
assign _23837_ = _23156_ ^ _23839_ /*2343*/;
assign _23838_ = _23830_ & _23837_ /*2341*/;
assign _23835_ = _23836_ | _23838_ /*2339*/;
assign _23542_ = _23830_ ^ _23837_ /*2342*/;
assign _23844_ = D[58] ^ Q[3] /*2338*/;
assign _23841_ = _23157_ & _23844_ /*2334*/;
assign _23842_ = _23157_ ^ _23844_ /*2337*/;
assign _23843_ = _23835_ & _23842_ /*2335*/;
assign _23840_ = _23841_ | _23843_ /*2333*/;
assign _23543_ = _23835_ ^ _23842_ /*2336*/;
assign _23849_ = D[59] ^ Q[3] /*2332*/;
assign _23846_ = _23158_ & _23849_ /*2328*/;
assign _23847_ = _23158_ ^ _23849_ /*2331*/;
assign _23848_ = _23840_ & _23847_ /*2329*/;
assign _23845_ = _23846_ | _23848_ /*2327*/;
assign _23544_ = _23840_ ^ _23847_ /*2330*/;
assign _23854_ = D[60] ^ Q[3] /*2326*/;
assign _23851_ = _23159_ & _23854_ /*2322*/;
assign _23852_ = _23159_ ^ _23854_ /*2325*/;
assign _23853_ = _23845_ & _23852_ /*2323*/;
assign _23850_ = _23851_ | _23853_ /*2321*/;
assign _23545_ = _23845_ ^ _23852_ /*2324*/;
assign _23859_ = D[61] ^ Q[3] /*2320*/;
assign _23856_ = _23160_ & _23859_ /*2316*/;
assign _23857_ = _23160_ ^ _23859_ /*2319*/;
assign _23858_ = _23850_ & _23857_ /*2317*/;
assign _23855_ = _23856_ | _23858_ /*2315*/;
assign _23546_ = _23850_ ^ _23857_ /*2318*/;
assign _23864_ = D[62] ^ Q[3] /*2314*/;
assign _23861_ = _23161_ & _23864_ /*2310*/;
assign _23862_ = _23161_ ^ _23864_ /*2313*/;
assign _23863_ = _23855_ & _23862_ /*2311*/;
assign _23860_ = _23861_ | _23863_ /*2309*/;
assign _23547_ = _23855_ ^ _23862_ /*2312*/;
assign _23868_ = zeroWire ^ Q[3] /*2308*/;
assign _23865_ = _23162_ & _23868_ /*2304*/;
assign _23866_ = _23162_ ^ _23868_ /*2307*/;
assign _23867_ = _23860_ & _23866_ /*2305*/;
assign Q[2] = _23865_ | _23867_ /*2303*/;
assign _23548_ = _23860_ ^ _23866_ /*2306*/;
assign _23939_ = D[0] ^ Q[2] /*1917*/;
assign _23936_ = R_0[1] & _23939_ /*1913*/;
assign _23937_ = R_0[1] ^ _23939_ /*1916*/;
assign _23938_ = Q[2] & _23937_ /*1914*/;
assign _23935_ = _23936_ | _23938_ /*1912*/;
assign _23870_ = Q[2] ^ _23937_ /*1915*/;
assign _23944_ = D[1] ^ Q[2] /*1911*/;
assign _23941_ = _23485_ & _23944_ /*1907*/;
assign _23942_ = _23485_ ^ _23944_ /*1910*/;
assign _23943_ = _23935_ & _23942_ /*1908*/;
assign _23940_ = _23941_ | _23943_ /*1906*/;
assign _23871_ = _23935_ ^ _23942_ /*1909*/;
assign _23949_ = D[2] ^ Q[2] /*1905*/;
assign _23946_ = _23486_ & _23949_ /*1901*/;
assign _23947_ = _23486_ ^ _23949_ /*1904*/;
assign _23948_ = _23940_ & _23947_ /*1902*/;
assign _23945_ = _23946_ | _23948_ /*1900*/;
assign _23872_ = _23940_ ^ _23947_ /*1903*/;
assign _23954_ = D[3] ^ Q[2] /*1899*/;
assign _23951_ = _23487_ & _23954_ /*1895*/;
assign _23952_ = _23487_ ^ _23954_ /*1898*/;
assign _23953_ = _23945_ & _23952_ /*1896*/;
assign _23950_ = _23951_ | _23953_ /*1894*/;
assign _23873_ = _23945_ ^ _23952_ /*1897*/;
assign _23959_ = D[4] ^ Q[2] /*1893*/;
assign _23956_ = _23488_ & _23959_ /*1889*/;
assign _23957_ = _23488_ ^ _23959_ /*1892*/;
assign _23958_ = _23950_ & _23957_ /*1890*/;
assign _23955_ = _23956_ | _23958_ /*1888*/;
assign _23874_ = _23950_ ^ _23957_ /*1891*/;
assign _23964_ = D[5] ^ Q[2] /*1887*/;
assign _23961_ = _23489_ & _23964_ /*1883*/;
assign _23962_ = _23489_ ^ _23964_ /*1886*/;
assign _23963_ = _23955_ & _23962_ /*1884*/;
assign _23960_ = _23961_ | _23963_ /*1882*/;
assign _23875_ = _23955_ ^ _23962_ /*1885*/;
assign _23969_ = D[6] ^ Q[2] /*1881*/;
assign _23966_ = _23490_ & _23969_ /*1877*/;
assign _23967_ = _23490_ ^ _23969_ /*1880*/;
assign _23968_ = _23960_ & _23967_ /*1878*/;
assign _23965_ = _23966_ | _23968_ /*1876*/;
assign _23876_ = _23960_ ^ _23967_ /*1879*/;
assign _23974_ = D[7] ^ Q[2] /*1875*/;
assign _23971_ = _23491_ & _23974_ /*1871*/;
assign _23972_ = _23491_ ^ _23974_ /*1874*/;
assign _23973_ = _23965_ & _23972_ /*1872*/;
assign _23970_ = _23971_ | _23973_ /*1870*/;
assign _23877_ = _23965_ ^ _23972_ /*1873*/;
assign _23979_ = D[8] ^ Q[2] /*1869*/;
assign _23976_ = _23492_ & _23979_ /*1865*/;
assign _23977_ = _23492_ ^ _23979_ /*1868*/;
assign _23978_ = _23970_ & _23977_ /*1866*/;
assign _23975_ = _23976_ | _23978_ /*1864*/;
assign _23878_ = _23970_ ^ _23977_ /*1867*/;
assign _23984_ = D[9] ^ Q[2] /*1863*/;
assign _23981_ = _23493_ & _23984_ /*1859*/;
assign _23982_ = _23493_ ^ _23984_ /*1862*/;
assign _23983_ = _23975_ & _23982_ /*1860*/;
assign _23980_ = _23981_ | _23983_ /*1858*/;
assign _23879_ = _23975_ ^ _23982_ /*1861*/;
assign _23989_ = D[10] ^ Q[2] /*1857*/;
assign _23986_ = _23494_ & _23989_ /*1853*/;
assign _23987_ = _23494_ ^ _23989_ /*1856*/;
assign _23988_ = _23980_ & _23987_ /*1854*/;
assign _23985_ = _23986_ | _23988_ /*1852*/;
assign _23880_ = _23980_ ^ _23987_ /*1855*/;
assign _23994_ = D[11] ^ Q[2] /*1851*/;
assign _23991_ = _23495_ & _23994_ /*1847*/;
assign _23992_ = _23495_ ^ _23994_ /*1850*/;
assign _23993_ = _23985_ & _23992_ /*1848*/;
assign _23990_ = _23991_ | _23993_ /*1846*/;
assign _23881_ = _23985_ ^ _23992_ /*1849*/;
assign _23999_ = D[12] ^ Q[2] /*1845*/;
assign _23996_ = _23496_ & _23999_ /*1841*/;
assign _23997_ = _23496_ ^ _23999_ /*1844*/;
assign _23998_ = _23990_ & _23997_ /*1842*/;
assign _23995_ = _23996_ | _23998_ /*1840*/;
assign _23882_ = _23990_ ^ _23997_ /*1843*/;
assign _24004_ = D[13] ^ Q[2] /*1839*/;
assign _24001_ = _23497_ & _24004_ /*1835*/;
assign _24002_ = _23497_ ^ _24004_ /*1838*/;
assign _24003_ = _23995_ & _24002_ /*1836*/;
assign _24000_ = _24001_ | _24003_ /*1834*/;
assign _23883_ = _23995_ ^ _24002_ /*1837*/;
assign _24009_ = D[14] ^ Q[2] /*1833*/;
assign _24006_ = _23498_ & _24009_ /*1829*/;
assign _24007_ = _23498_ ^ _24009_ /*1832*/;
assign _24008_ = _24000_ & _24007_ /*1830*/;
assign _24005_ = _24006_ | _24008_ /*1828*/;
assign _23884_ = _24000_ ^ _24007_ /*1831*/;
assign _24014_ = D[15] ^ Q[2] /*1827*/;
assign _24011_ = _23499_ & _24014_ /*1823*/;
assign _24012_ = _23499_ ^ _24014_ /*1826*/;
assign _24013_ = _24005_ & _24012_ /*1824*/;
assign _24010_ = _24011_ | _24013_ /*1822*/;
assign _23885_ = _24005_ ^ _24012_ /*1825*/;
assign _24019_ = D[16] ^ Q[2] /*1821*/;
assign _24016_ = _23500_ & _24019_ /*1817*/;
assign _24017_ = _23500_ ^ _24019_ /*1820*/;
assign _24018_ = _24010_ & _24017_ /*1818*/;
assign _24015_ = _24016_ | _24018_ /*1816*/;
assign _23886_ = _24010_ ^ _24017_ /*1819*/;
assign _24024_ = D[17] ^ Q[2] /*1815*/;
assign _24021_ = _23501_ & _24024_ /*1811*/;
assign _24022_ = _23501_ ^ _24024_ /*1814*/;
assign _24023_ = _24015_ & _24022_ /*1812*/;
assign _24020_ = _24021_ | _24023_ /*1810*/;
assign _23887_ = _24015_ ^ _24022_ /*1813*/;
assign _24029_ = D[18] ^ Q[2] /*1809*/;
assign _24026_ = _23502_ & _24029_ /*1805*/;
assign _24027_ = _23502_ ^ _24029_ /*1808*/;
assign _24028_ = _24020_ & _24027_ /*1806*/;
assign _24025_ = _24026_ | _24028_ /*1804*/;
assign _23888_ = _24020_ ^ _24027_ /*1807*/;
assign _24034_ = D[19] ^ Q[2] /*1803*/;
assign _24031_ = _23503_ & _24034_ /*1799*/;
assign _24032_ = _23503_ ^ _24034_ /*1802*/;
assign _24033_ = _24025_ & _24032_ /*1800*/;
assign _24030_ = _24031_ | _24033_ /*1798*/;
assign _23889_ = _24025_ ^ _24032_ /*1801*/;
assign _24039_ = D[20] ^ Q[2] /*1797*/;
assign _24036_ = _23504_ & _24039_ /*1793*/;
assign _24037_ = _23504_ ^ _24039_ /*1796*/;
assign _24038_ = _24030_ & _24037_ /*1794*/;
assign _24035_ = _24036_ | _24038_ /*1792*/;
assign _23890_ = _24030_ ^ _24037_ /*1795*/;
assign _24044_ = D[21] ^ Q[2] /*1791*/;
assign _24041_ = _23505_ & _24044_ /*1787*/;
assign _24042_ = _23505_ ^ _24044_ /*1790*/;
assign _24043_ = _24035_ & _24042_ /*1788*/;
assign _24040_ = _24041_ | _24043_ /*1786*/;
assign _23891_ = _24035_ ^ _24042_ /*1789*/;
assign _24049_ = D[22] ^ Q[2] /*1785*/;
assign _24046_ = _23506_ & _24049_ /*1781*/;
assign _24047_ = _23506_ ^ _24049_ /*1784*/;
assign _24048_ = _24040_ & _24047_ /*1782*/;
assign _24045_ = _24046_ | _24048_ /*1780*/;
assign _23892_ = _24040_ ^ _24047_ /*1783*/;
assign _24054_ = D[23] ^ Q[2] /*1779*/;
assign _24051_ = _23507_ & _24054_ /*1775*/;
assign _24052_ = _23507_ ^ _24054_ /*1778*/;
assign _24053_ = _24045_ & _24052_ /*1776*/;
assign _24050_ = _24051_ | _24053_ /*1774*/;
assign _23893_ = _24045_ ^ _24052_ /*1777*/;
assign _24059_ = D[24] ^ Q[2] /*1773*/;
assign _24056_ = _23508_ & _24059_ /*1769*/;
assign _24057_ = _23508_ ^ _24059_ /*1772*/;
assign _24058_ = _24050_ & _24057_ /*1770*/;
assign _24055_ = _24056_ | _24058_ /*1768*/;
assign _23894_ = _24050_ ^ _24057_ /*1771*/;
assign _24064_ = D[25] ^ Q[2] /*1767*/;
assign _24061_ = _23509_ & _24064_ /*1763*/;
assign _24062_ = _23509_ ^ _24064_ /*1766*/;
assign _24063_ = _24055_ & _24062_ /*1764*/;
assign _24060_ = _24061_ | _24063_ /*1762*/;
assign _23895_ = _24055_ ^ _24062_ /*1765*/;
assign _24069_ = D[26] ^ Q[2] /*1761*/;
assign _24066_ = _23510_ & _24069_ /*1757*/;
assign _24067_ = _23510_ ^ _24069_ /*1760*/;
assign _24068_ = _24060_ & _24067_ /*1758*/;
assign _24065_ = _24066_ | _24068_ /*1756*/;
assign _23896_ = _24060_ ^ _24067_ /*1759*/;
assign _24074_ = D[27] ^ Q[2] /*1755*/;
assign _24071_ = _23511_ & _24074_ /*1751*/;
assign _24072_ = _23511_ ^ _24074_ /*1754*/;
assign _24073_ = _24065_ & _24072_ /*1752*/;
assign _24070_ = _24071_ | _24073_ /*1750*/;
assign _23897_ = _24065_ ^ _24072_ /*1753*/;
assign _24079_ = D[28] ^ Q[2] /*1749*/;
assign _24076_ = _23512_ & _24079_ /*1745*/;
assign _24077_ = _23512_ ^ _24079_ /*1748*/;
assign _24078_ = _24070_ & _24077_ /*1746*/;
assign _24075_ = _24076_ | _24078_ /*1744*/;
assign _23898_ = _24070_ ^ _24077_ /*1747*/;
assign _24084_ = D[29] ^ Q[2] /*1743*/;
assign _24081_ = _23513_ & _24084_ /*1739*/;
assign _24082_ = _23513_ ^ _24084_ /*1742*/;
assign _24083_ = _24075_ & _24082_ /*1740*/;
assign _24080_ = _24081_ | _24083_ /*1738*/;
assign _23899_ = _24075_ ^ _24082_ /*1741*/;
assign _24089_ = D[30] ^ Q[2] /*1737*/;
assign _24086_ = _23514_ & _24089_ /*1733*/;
assign _24087_ = _23514_ ^ _24089_ /*1736*/;
assign _24088_ = _24080_ & _24087_ /*1734*/;
assign _24085_ = _24086_ | _24088_ /*1732*/;
assign _23900_ = _24080_ ^ _24087_ /*1735*/;
assign _24094_ = D[31] ^ Q[2] /*1731*/;
assign _24091_ = _23515_ & _24094_ /*1727*/;
assign _24092_ = _23515_ ^ _24094_ /*1730*/;
assign _24093_ = _24085_ & _24092_ /*1728*/;
assign _24090_ = _24091_ | _24093_ /*1726*/;
assign _23901_ = _24085_ ^ _24092_ /*1729*/;
assign _24099_ = D[32] ^ Q[2] /*1725*/;
assign _24096_ = _23516_ & _24099_ /*1721*/;
assign _24097_ = _23516_ ^ _24099_ /*1724*/;
assign _24098_ = _24090_ & _24097_ /*1722*/;
assign _24095_ = _24096_ | _24098_ /*1720*/;
assign _23902_ = _24090_ ^ _24097_ /*1723*/;
assign _24104_ = D[33] ^ Q[2] /*1719*/;
assign _24101_ = _23517_ & _24104_ /*1715*/;
assign _24102_ = _23517_ ^ _24104_ /*1718*/;
assign _24103_ = _24095_ & _24102_ /*1716*/;
assign _24100_ = _24101_ | _24103_ /*1714*/;
assign _23903_ = _24095_ ^ _24102_ /*1717*/;
assign _24109_ = D[34] ^ Q[2] /*1713*/;
assign _24106_ = _23518_ & _24109_ /*1709*/;
assign _24107_ = _23518_ ^ _24109_ /*1712*/;
assign _24108_ = _24100_ & _24107_ /*1710*/;
assign _24105_ = _24106_ | _24108_ /*1708*/;
assign _23904_ = _24100_ ^ _24107_ /*1711*/;
assign _24114_ = D[35] ^ Q[2] /*1707*/;
assign _24111_ = _23519_ & _24114_ /*1703*/;
assign _24112_ = _23519_ ^ _24114_ /*1706*/;
assign _24113_ = _24105_ & _24112_ /*1704*/;
assign _24110_ = _24111_ | _24113_ /*1702*/;
assign _23905_ = _24105_ ^ _24112_ /*1705*/;
assign _24119_ = D[36] ^ Q[2] /*1701*/;
assign _24116_ = _23520_ & _24119_ /*1697*/;
assign _24117_ = _23520_ ^ _24119_ /*1700*/;
assign _24118_ = _24110_ & _24117_ /*1698*/;
assign _24115_ = _24116_ | _24118_ /*1696*/;
assign _23906_ = _24110_ ^ _24117_ /*1699*/;
assign _24124_ = D[37] ^ Q[2] /*1695*/;
assign _24121_ = _23521_ & _24124_ /*1691*/;
assign _24122_ = _23521_ ^ _24124_ /*1694*/;
assign _24123_ = _24115_ & _24122_ /*1692*/;
assign _24120_ = _24121_ | _24123_ /*1690*/;
assign _23907_ = _24115_ ^ _24122_ /*1693*/;
assign _24129_ = D[38] ^ Q[2] /*1689*/;
assign _24126_ = _23522_ & _24129_ /*1685*/;
assign _24127_ = _23522_ ^ _24129_ /*1688*/;
assign _24128_ = _24120_ & _24127_ /*1686*/;
assign _24125_ = _24126_ | _24128_ /*1684*/;
assign _23908_ = _24120_ ^ _24127_ /*1687*/;
assign _24134_ = D[39] ^ Q[2] /*1683*/;
assign _24131_ = _23523_ & _24134_ /*1679*/;
assign _24132_ = _23523_ ^ _24134_ /*1682*/;
assign _24133_ = _24125_ & _24132_ /*1680*/;
assign _24130_ = _24131_ | _24133_ /*1678*/;
assign _23909_ = _24125_ ^ _24132_ /*1681*/;
assign _24139_ = D[40] ^ Q[2] /*1677*/;
assign _24136_ = _23524_ & _24139_ /*1673*/;
assign _24137_ = _23524_ ^ _24139_ /*1676*/;
assign _24138_ = _24130_ & _24137_ /*1674*/;
assign _24135_ = _24136_ | _24138_ /*1672*/;
assign _23910_ = _24130_ ^ _24137_ /*1675*/;
assign _24144_ = D[41] ^ Q[2] /*1671*/;
assign _24141_ = _23525_ & _24144_ /*1667*/;
assign _24142_ = _23525_ ^ _24144_ /*1670*/;
assign _24143_ = _24135_ & _24142_ /*1668*/;
assign _24140_ = _24141_ | _24143_ /*1666*/;
assign _23911_ = _24135_ ^ _24142_ /*1669*/;
assign _24149_ = D[42] ^ Q[2] /*1665*/;
assign _24146_ = _23526_ & _24149_ /*1661*/;
assign _24147_ = _23526_ ^ _24149_ /*1664*/;
assign _24148_ = _24140_ & _24147_ /*1662*/;
assign _24145_ = _24146_ | _24148_ /*1660*/;
assign _23912_ = _24140_ ^ _24147_ /*1663*/;
assign _24154_ = D[43] ^ Q[2] /*1659*/;
assign _24151_ = _23527_ & _24154_ /*1655*/;
assign _24152_ = _23527_ ^ _24154_ /*1658*/;
assign _24153_ = _24145_ & _24152_ /*1656*/;
assign _24150_ = _24151_ | _24153_ /*1654*/;
assign _23913_ = _24145_ ^ _24152_ /*1657*/;
assign _24159_ = D[44] ^ Q[2] /*1653*/;
assign _24156_ = _23528_ & _24159_ /*1649*/;
assign _24157_ = _23528_ ^ _24159_ /*1652*/;
assign _24158_ = _24150_ & _24157_ /*1650*/;
assign _24155_ = _24156_ | _24158_ /*1648*/;
assign _23914_ = _24150_ ^ _24157_ /*1651*/;
assign _24164_ = D[45] ^ Q[2] /*1647*/;
assign _24161_ = _23529_ & _24164_ /*1643*/;
assign _24162_ = _23529_ ^ _24164_ /*1646*/;
assign _24163_ = _24155_ & _24162_ /*1644*/;
assign _24160_ = _24161_ | _24163_ /*1642*/;
assign _23915_ = _24155_ ^ _24162_ /*1645*/;
assign _24169_ = D[46] ^ Q[2] /*1641*/;
assign _24166_ = _23530_ & _24169_ /*1637*/;
assign _24167_ = _23530_ ^ _24169_ /*1640*/;
assign _24168_ = _24160_ & _24167_ /*1638*/;
assign _24165_ = _24166_ | _24168_ /*1636*/;
assign _23916_ = _24160_ ^ _24167_ /*1639*/;
assign _24174_ = D[47] ^ Q[2] /*1635*/;
assign _24171_ = _23531_ & _24174_ /*1631*/;
assign _24172_ = _23531_ ^ _24174_ /*1634*/;
assign _24173_ = _24165_ & _24172_ /*1632*/;
assign _24170_ = _24171_ | _24173_ /*1630*/;
assign _23917_ = _24165_ ^ _24172_ /*1633*/;
assign _24179_ = D[48] ^ Q[2] /*1629*/;
assign _24176_ = _23532_ & _24179_ /*1625*/;
assign _24177_ = _23532_ ^ _24179_ /*1628*/;
assign _24178_ = _24170_ & _24177_ /*1626*/;
assign _24175_ = _24176_ | _24178_ /*1624*/;
assign _23918_ = _24170_ ^ _24177_ /*1627*/;
assign _24184_ = D[49] ^ Q[2] /*1623*/;
assign _24181_ = _23533_ & _24184_ /*1619*/;
assign _24182_ = _23533_ ^ _24184_ /*1622*/;
assign _24183_ = _24175_ & _24182_ /*1620*/;
assign _24180_ = _24181_ | _24183_ /*1618*/;
assign _23919_ = _24175_ ^ _24182_ /*1621*/;
assign _24189_ = D[50] ^ Q[2] /*1617*/;
assign _24186_ = _23534_ & _24189_ /*1613*/;
assign _24187_ = _23534_ ^ _24189_ /*1616*/;
assign _24188_ = _24180_ & _24187_ /*1614*/;
assign _24185_ = _24186_ | _24188_ /*1612*/;
assign _23920_ = _24180_ ^ _24187_ /*1615*/;
assign _24194_ = D[51] ^ Q[2] /*1611*/;
assign _24191_ = _23535_ & _24194_ /*1607*/;
assign _24192_ = _23535_ ^ _24194_ /*1610*/;
assign _24193_ = _24185_ & _24192_ /*1608*/;
assign _24190_ = _24191_ | _24193_ /*1606*/;
assign _23921_ = _24185_ ^ _24192_ /*1609*/;
assign _24199_ = D[52] ^ Q[2] /*1605*/;
assign _24196_ = _23536_ & _24199_ /*1601*/;
assign _24197_ = _23536_ ^ _24199_ /*1604*/;
assign _24198_ = _24190_ & _24197_ /*1602*/;
assign _24195_ = _24196_ | _24198_ /*1600*/;
assign _23922_ = _24190_ ^ _24197_ /*1603*/;
assign _24204_ = D[53] ^ Q[2] /*1599*/;
assign _24201_ = _23537_ & _24204_ /*1595*/;
assign _24202_ = _23537_ ^ _24204_ /*1598*/;
assign _24203_ = _24195_ & _24202_ /*1596*/;
assign _24200_ = _24201_ | _24203_ /*1594*/;
assign _23923_ = _24195_ ^ _24202_ /*1597*/;
assign _24209_ = D[54] ^ Q[2] /*1593*/;
assign _24206_ = _23538_ & _24209_ /*1589*/;
assign _24207_ = _23538_ ^ _24209_ /*1592*/;
assign _24208_ = _24200_ & _24207_ /*1590*/;
assign _24205_ = _24206_ | _24208_ /*1588*/;
assign _23924_ = _24200_ ^ _24207_ /*1591*/;
assign _24214_ = D[55] ^ Q[2] /*1587*/;
assign _24211_ = _23539_ & _24214_ /*1583*/;
assign _24212_ = _23539_ ^ _24214_ /*1586*/;
assign _24213_ = _24205_ & _24212_ /*1584*/;
assign _24210_ = _24211_ | _24213_ /*1582*/;
assign _23925_ = _24205_ ^ _24212_ /*1585*/;
assign _24219_ = D[56] ^ Q[2] /*1581*/;
assign _24216_ = _23540_ & _24219_ /*1577*/;
assign _24217_ = _23540_ ^ _24219_ /*1580*/;
assign _24218_ = _24210_ & _24217_ /*1578*/;
assign _24215_ = _24216_ | _24218_ /*1576*/;
assign _23926_ = _24210_ ^ _24217_ /*1579*/;
assign _24224_ = D[57] ^ Q[2] /*1575*/;
assign _24221_ = _23541_ & _24224_ /*1571*/;
assign _24222_ = _23541_ ^ _24224_ /*1574*/;
assign _24223_ = _24215_ & _24222_ /*1572*/;
assign _24220_ = _24221_ | _24223_ /*1570*/;
assign _23927_ = _24215_ ^ _24222_ /*1573*/;
assign _24229_ = D[58] ^ Q[2] /*1569*/;
assign _24226_ = _23542_ & _24229_ /*1565*/;
assign _24227_ = _23542_ ^ _24229_ /*1568*/;
assign _24228_ = _24220_ & _24227_ /*1566*/;
assign _24225_ = _24226_ | _24228_ /*1564*/;
assign _23928_ = _24220_ ^ _24227_ /*1567*/;
assign _24234_ = D[59] ^ Q[2] /*1563*/;
assign _24231_ = _23543_ & _24234_ /*1559*/;
assign _24232_ = _23543_ ^ _24234_ /*1562*/;
assign _24233_ = _24225_ & _24232_ /*1560*/;
assign _24230_ = _24231_ | _24233_ /*1558*/;
assign _23929_ = _24225_ ^ _24232_ /*1561*/;
assign _24239_ = D[60] ^ Q[2] /*1557*/;
assign _24236_ = _23544_ & _24239_ /*1553*/;
assign _24237_ = _23544_ ^ _24239_ /*1556*/;
assign _24238_ = _24230_ & _24237_ /*1554*/;
assign _24235_ = _24236_ | _24238_ /*1552*/;
assign _23930_ = _24230_ ^ _24237_ /*1555*/;
assign _24244_ = D[61] ^ Q[2] /*1551*/;
assign _24241_ = _23545_ & _24244_ /*1547*/;
assign _24242_ = _23545_ ^ _24244_ /*1550*/;
assign _24243_ = _24235_ & _24242_ /*1548*/;
assign _24240_ = _24241_ | _24243_ /*1546*/;
assign _23931_ = _24235_ ^ _24242_ /*1549*/;
assign _24249_ = D[62] ^ Q[2] /*1545*/;
assign _24246_ = _23546_ & _24249_ /*1541*/;
assign _24247_ = _23546_ ^ _24249_ /*1544*/;
assign _24248_ = _24240_ & _24247_ /*1542*/;
assign _24245_ = _24246_ | _24248_ /*1540*/;
assign _23932_ = _24240_ ^ _24247_ /*1543*/;
assign _24253_ = zeroWire ^ Q[2] /*1539*/;
assign _24250_ = _23547_ & _24253_ /*1535*/;
assign _24251_ = _23547_ ^ _24253_ /*1538*/;
assign _24252_ = _24245_ & _24251_ /*1536*/;
assign Q[1] = _24250_ | _24252_ /*1534*/;
assign _23933_ = _24245_ ^ _24251_ /*1537*/;
assign _24324_ = D[0] ^ Q[1] /*1148*/;
assign _24321_ = R_0[0] & _24324_ /*1144*/;
assign _24322_ = R_0[0] ^ _24324_ /*1147*/;
assign _24323_ = Q[1] & _24322_ /*1145*/;
assign _24320_ = _24321_ | _24323_ /*1143*/;
assign _24255_ = Q[1] ^ _24322_ /*1146*/;
assign _24329_ = D[1] ^ Q[1] /*1142*/;
assign _24326_ = _23870_ & _24329_ /*1138*/;
assign _24327_ = _23870_ ^ _24329_ /*1141*/;
assign _24328_ = _24320_ & _24327_ /*1139*/;
assign _24325_ = _24326_ | _24328_ /*1137*/;
assign _24256_ = _24320_ ^ _24327_ /*1140*/;
assign _24334_ = D[2] ^ Q[1] /*1136*/;
assign _24331_ = _23871_ & _24334_ /*1132*/;
assign _24332_ = _23871_ ^ _24334_ /*1135*/;
assign _24333_ = _24325_ & _24332_ /*1133*/;
assign _24330_ = _24331_ | _24333_ /*1131*/;
assign _24257_ = _24325_ ^ _24332_ /*1134*/;
assign _24339_ = D[3] ^ Q[1] /*1130*/;
assign _24336_ = _23872_ & _24339_ /*1126*/;
assign _24337_ = _23872_ ^ _24339_ /*1129*/;
assign _24338_ = _24330_ & _24337_ /*1127*/;
assign _24335_ = _24336_ | _24338_ /*1125*/;
assign _24258_ = _24330_ ^ _24337_ /*1128*/;
assign _24344_ = D[4] ^ Q[1] /*1124*/;
assign _24341_ = _23873_ & _24344_ /*1120*/;
assign _24342_ = _23873_ ^ _24344_ /*1123*/;
assign _24343_ = _24335_ & _24342_ /*1121*/;
assign _24340_ = _24341_ | _24343_ /*1119*/;
assign _24259_ = _24335_ ^ _24342_ /*1122*/;
assign _24349_ = D[5] ^ Q[1] /*1118*/;
assign _24346_ = _23874_ & _24349_ /*1114*/;
assign _24347_ = _23874_ ^ _24349_ /*1117*/;
assign _24348_ = _24340_ & _24347_ /*1115*/;
assign _24345_ = _24346_ | _24348_ /*1113*/;
assign _24260_ = _24340_ ^ _24347_ /*1116*/;
assign _24354_ = D[6] ^ Q[1] /*1112*/;
assign _24351_ = _23875_ & _24354_ /*1108*/;
assign _24352_ = _23875_ ^ _24354_ /*1111*/;
assign _24353_ = _24345_ & _24352_ /*1109*/;
assign _24350_ = _24351_ | _24353_ /*1107*/;
assign _24261_ = _24345_ ^ _24352_ /*1110*/;
assign _24359_ = D[7] ^ Q[1] /*1106*/;
assign _24356_ = _23876_ & _24359_ /*1102*/;
assign _24357_ = _23876_ ^ _24359_ /*1105*/;
assign _24358_ = _24350_ & _24357_ /*1103*/;
assign _24355_ = _24356_ | _24358_ /*1101*/;
assign _24262_ = _24350_ ^ _24357_ /*1104*/;
assign _24364_ = D[8] ^ Q[1] /*1100*/;
assign _24361_ = _23877_ & _24364_ /*1096*/;
assign _24362_ = _23877_ ^ _24364_ /*1099*/;
assign _24363_ = _24355_ & _24362_ /*1097*/;
assign _24360_ = _24361_ | _24363_ /*1095*/;
assign _24263_ = _24355_ ^ _24362_ /*1098*/;
assign _24369_ = D[9] ^ Q[1] /*1094*/;
assign _24366_ = _23878_ & _24369_ /*1090*/;
assign _24367_ = _23878_ ^ _24369_ /*1093*/;
assign _24368_ = _24360_ & _24367_ /*1091*/;
assign _24365_ = _24366_ | _24368_ /*1089*/;
assign _24264_ = _24360_ ^ _24367_ /*1092*/;
assign _24374_ = D[10] ^ Q[1] /*1088*/;
assign _24371_ = _23879_ & _24374_ /*1084*/;
assign _24372_ = _23879_ ^ _24374_ /*1087*/;
assign _24373_ = _24365_ & _24372_ /*1085*/;
assign _24370_ = _24371_ | _24373_ /*1083*/;
assign _24265_ = _24365_ ^ _24372_ /*1086*/;
assign _24379_ = D[11] ^ Q[1] /*1082*/;
assign _24376_ = _23880_ & _24379_ /*1078*/;
assign _24377_ = _23880_ ^ _24379_ /*1081*/;
assign _24378_ = _24370_ & _24377_ /*1079*/;
assign _24375_ = _24376_ | _24378_ /*1077*/;
assign _24266_ = _24370_ ^ _24377_ /*1080*/;
assign _24384_ = D[12] ^ Q[1] /*1076*/;
assign _24381_ = _23881_ & _24384_ /*1072*/;
assign _24382_ = _23881_ ^ _24384_ /*1075*/;
assign _24383_ = _24375_ & _24382_ /*1073*/;
assign _24380_ = _24381_ | _24383_ /*1071*/;
assign _24267_ = _24375_ ^ _24382_ /*1074*/;
assign _24389_ = D[13] ^ Q[1] /*1070*/;
assign _24386_ = _23882_ & _24389_ /*1066*/;
assign _24387_ = _23882_ ^ _24389_ /*1069*/;
assign _24388_ = _24380_ & _24387_ /*1067*/;
assign _24385_ = _24386_ | _24388_ /*1065*/;
assign _24268_ = _24380_ ^ _24387_ /*1068*/;
assign _24394_ = D[14] ^ Q[1] /*1064*/;
assign _24391_ = _23883_ & _24394_ /*1060*/;
assign _24392_ = _23883_ ^ _24394_ /*1063*/;
assign _24393_ = _24385_ & _24392_ /*1061*/;
assign _24390_ = _24391_ | _24393_ /*1059*/;
assign _24269_ = _24385_ ^ _24392_ /*1062*/;
assign _24399_ = D[15] ^ Q[1] /*1058*/;
assign _24396_ = _23884_ & _24399_ /*1054*/;
assign _24397_ = _23884_ ^ _24399_ /*1057*/;
assign _24398_ = _24390_ & _24397_ /*1055*/;
assign _24395_ = _24396_ | _24398_ /*1053*/;
assign _24270_ = _24390_ ^ _24397_ /*1056*/;
assign _24404_ = D[16] ^ Q[1] /*1052*/;
assign _24401_ = _23885_ & _24404_ /*1048*/;
assign _24402_ = _23885_ ^ _24404_ /*1051*/;
assign _24403_ = _24395_ & _24402_ /*1049*/;
assign _24400_ = _24401_ | _24403_ /*1047*/;
assign _24271_ = _24395_ ^ _24402_ /*1050*/;
assign _24409_ = D[17] ^ Q[1] /*1046*/;
assign _24406_ = _23886_ & _24409_ /*1042*/;
assign _24407_ = _23886_ ^ _24409_ /*1045*/;
assign _24408_ = _24400_ & _24407_ /*1043*/;
assign _24405_ = _24406_ | _24408_ /*1041*/;
assign _24272_ = _24400_ ^ _24407_ /*1044*/;
assign _24414_ = D[18] ^ Q[1] /*1040*/;
assign _24411_ = _23887_ & _24414_ /*1036*/;
assign _24412_ = _23887_ ^ _24414_ /*1039*/;
assign _24413_ = _24405_ & _24412_ /*1037*/;
assign _24410_ = _24411_ | _24413_ /*1035*/;
assign _24273_ = _24405_ ^ _24412_ /*1038*/;
assign _24419_ = D[19] ^ Q[1] /*1034*/;
assign _24416_ = _23888_ & _24419_ /*1030*/;
assign _24417_ = _23888_ ^ _24419_ /*1033*/;
assign _24418_ = _24410_ & _24417_ /*1031*/;
assign _24415_ = _24416_ | _24418_ /*1029*/;
assign _24274_ = _24410_ ^ _24417_ /*1032*/;
assign _24424_ = D[20] ^ Q[1] /*1028*/;
assign _24421_ = _23889_ & _24424_ /*1024*/;
assign _24422_ = _23889_ ^ _24424_ /*1027*/;
assign _24423_ = _24415_ & _24422_ /*1025*/;
assign _24420_ = _24421_ | _24423_ /*1023*/;
assign _24275_ = _24415_ ^ _24422_ /*1026*/;
assign _24429_ = D[21] ^ Q[1] /*1022*/;
assign _24426_ = _23890_ & _24429_ /*1018*/;
assign _24427_ = _23890_ ^ _24429_ /*1021*/;
assign _24428_ = _24420_ & _24427_ /*1019*/;
assign _24425_ = _24426_ | _24428_ /*1017*/;
assign _24276_ = _24420_ ^ _24427_ /*1020*/;
assign _24434_ = D[22] ^ Q[1] /*1016*/;
assign _24431_ = _23891_ & _24434_ /*1012*/;
assign _24432_ = _23891_ ^ _24434_ /*1015*/;
assign _24433_ = _24425_ & _24432_ /*1013*/;
assign _24430_ = _24431_ | _24433_ /*1011*/;
assign _24277_ = _24425_ ^ _24432_ /*1014*/;
assign _24439_ = D[23] ^ Q[1] /*1010*/;
assign _24436_ = _23892_ & _24439_ /*1006*/;
assign _24437_ = _23892_ ^ _24439_ /*1009*/;
assign _24438_ = _24430_ & _24437_ /*1007*/;
assign _24435_ = _24436_ | _24438_ /*1005*/;
assign _24278_ = _24430_ ^ _24437_ /*1008*/;
assign _24444_ = D[24] ^ Q[1] /*1004*/;
assign _24441_ = _23893_ & _24444_ /*1000*/;
assign _24442_ = _23893_ ^ _24444_ /*1003*/;
assign _24443_ = _24435_ & _24442_ /*1001*/;
assign _24440_ = _24441_ | _24443_ /*999*/;
assign _24279_ = _24435_ ^ _24442_ /*1002*/;
assign _24449_ = D[25] ^ Q[1] /*998*/;
assign _24446_ = _23894_ & _24449_ /*994*/;
assign _24447_ = _23894_ ^ _24449_ /*997*/;
assign _24448_ = _24440_ & _24447_ /*995*/;
assign _24445_ = _24446_ | _24448_ /*993*/;
assign _24280_ = _24440_ ^ _24447_ /*996*/;
assign _24454_ = D[26] ^ Q[1] /*992*/;
assign _24451_ = _23895_ & _24454_ /*988*/;
assign _24452_ = _23895_ ^ _24454_ /*991*/;
assign _24453_ = _24445_ & _24452_ /*989*/;
assign _24450_ = _24451_ | _24453_ /*987*/;
assign _24281_ = _24445_ ^ _24452_ /*990*/;
assign _24459_ = D[27] ^ Q[1] /*986*/;
assign _24456_ = _23896_ & _24459_ /*982*/;
assign _24457_ = _23896_ ^ _24459_ /*985*/;
assign _24458_ = _24450_ & _24457_ /*983*/;
assign _24455_ = _24456_ | _24458_ /*981*/;
assign _24282_ = _24450_ ^ _24457_ /*984*/;
assign _24464_ = D[28] ^ Q[1] /*980*/;
assign _24461_ = _23897_ & _24464_ /*976*/;
assign _24462_ = _23897_ ^ _24464_ /*979*/;
assign _24463_ = _24455_ & _24462_ /*977*/;
assign _24460_ = _24461_ | _24463_ /*975*/;
assign _24283_ = _24455_ ^ _24462_ /*978*/;
assign _24469_ = D[29] ^ Q[1] /*974*/;
assign _24466_ = _23898_ & _24469_ /*970*/;
assign _24467_ = _23898_ ^ _24469_ /*973*/;
assign _24468_ = _24460_ & _24467_ /*971*/;
assign _24465_ = _24466_ | _24468_ /*969*/;
assign _24284_ = _24460_ ^ _24467_ /*972*/;
assign _24474_ = D[30] ^ Q[1] /*968*/;
assign _24471_ = _23899_ & _24474_ /*964*/;
assign _24472_ = _23899_ ^ _24474_ /*967*/;
assign _24473_ = _24465_ & _24472_ /*965*/;
assign _24470_ = _24471_ | _24473_ /*963*/;
assign _24285_ = _24465_ ^ _24472_ /*966*/;
assign _24479_ = D[31] ^ Q[1] /*962*/;
assign _24476_ = _23900_ & _24479_ /*958*/;
assign _24477_ = _23900_ ^ _24479_ /*961*/;
assign _24478_ = _24470_ & _24477_ /*959*/;
assign _24475_ = _24476_ | _24478_ /*957*/;
assign _24286_ = _24470_ ^ _24477_ /*960*/;
assign _24484_ = D[32] ^ Q[1] /*956*/;
assign _24481_ = _23901_ & _24484_ /*952*/;
assign _24482_ = _23901_ ^ _24484_ /*955*/;
assign _24483_ = _24475_ & _24482_ /*953*/;
assign _24480_ = _24481_ | _24483_ /*951*/;
assign _24287_ = _24475_ ^ _24482_ /*954*/;
assign _24489_ = D[33] ^ Q[1] /*950*/;
assign _24486_ = _23902_ & _24489_ /*946*/;
assign _24487_ = _23902_ ^ _24489_ /*949*/;
assign _24488_ = _24480_ & _24487_ /*947*/;
assign _24485_ = _24486_ | _24488_ /*945*/;
assign _24288_ = _24480_ ^ _24487_ /*948*/;
assign _24494_ = D[34] ^ Q[1] /*944*/;
assign _24491_ = _23903_ & _24494_ /*940*/;
assign _24492_ = _23903_ ^ _24494_ /*943*/;
assign _24493_ = _24485_ & _24492_ /*941*/;
assign _24490_ = _24491_ | _24493_ /*939*/;
assign _24289_ = _24485_ ^ _24492_ /*942*/;
assign _24499_ = D[35] ^ Q[1] /*938*/;
assign _24496_ = _23904_ & _24499_ /*934*/;
assign _24497_ = _23904_ ^ _24499_ /*937*/;
assign _24498_ = _24490_ & _24497_ /*935*/;
assign _24495_ = _24496_ | _24498_ /*933*/;
assign _24290_ = _24490_ ^ _24497_ /*936*/;
assign _24504_ = D[36] ^ Q[1] /*932*/;
assign _24501_ = _23905_ & _24504_ /*928*/;
assign _24502_ = _23905_ ^ _24504_ /*931*/;
assign _24503_ = _24495_ & _24502_ /*929*/;
assign _24500_ = _24501_ | _24503_ /*927*/;
assign _24291_ = _24495_ ^ _24502_ /*930*/;
assign _24509_ = D[37] ^ Q[1] /*926*/;
assign _24506_ = _23906_ & _24509_ /*922*/;
assign _24507_ = _23906_ ^ _24509_ /*925*/;
assign _24508_ = _24500_ & _24507_ /*923*/;
assign _24505_ = _24506_ | _24508_ /*921*/;
assign _24292_ = _24500_ ^ _24507_ /*924*/;
assign _24514_ = D[38] ^ Q[1] /*920*/;
assign _24511_ = _23907_ & _24514_ /*916*/;
assign _24512_ = _23907_ ^ _24514_ /*919*/;
assign _24513_ = _24505_ & _24512_ /*917*/;
assign _24510_ = _24511_ | _24513_ /*915*/;
assign _24293_ = _24505_ ^ _24512_ /*918*/;
assign _24519_ = D[39] ^ Q[1] /*914*/;
assign _24516_ = _23908_ & _24519_ /*910*/;
assign _24517_ = _23908_ ^ _24519_ /*913*/;
assign _24518_ = _24510_ & _24517_ /*911*/;
assign _24515_ = _24516_ | _24518_ /*909*/;
assign _24294_ = _24510_ ^ _24517_ /*912*/;
assign _24524_ = D[40] ^ Q[1] /*908*/;
assign _24521_ = _23909_ & _24524_ /*904*/;
assign _24522_ = _23909_ ^ _24524_ /*907*/;
assign _24523_ = _24515_ & _24522_ /*905*/;
assign _24520_ = _24521_ | _24523_ /*903*/;
assign _24295_ = _24515_ ^ _24522_ /*906*/;
assign _24529_ = D[41] ^ Q[1] /*902*/;
assign _24526_ = _23910_ & _24529_ /*898*/;
assign _24527_ = _23910_ ^ _24529_ /*901*/;
assign _24528_ = _24520_ & _24527_ /*899*/;
assign _24525_ = _24526_ | _24528_ /*897*/;
assign _24296_ = _24520_ ^ _24527_ /*900*/;
assign _24534_ = D[42] ^ Q[1] /*896*/;
assign _24531_ = _23911_ & _24534_ /*892*/;
assign _24532_ = _23911_ ^ _24534_ /*895*/;
assign _24533_ = _24525_ & _24532_ /*893*/;
assign _24530_ = _24531_ | _24533_ /*891*/;
assign _24297_ = _24525_ ^ _24532_ /*894*/;
assign _24539_ = D[43] ^ Q[1] /*890*/;
assign _24536_ = _23912_ & _24539_ /*886*/;
assign _24537_ = _23912_ ^ _24539_ /*889*/;
assign _24538_ = _24530_ & _24537_ /*887*/;
assign _24535_ = _24536_ | _24538_ /*885*/;
assign _24298_ = _24530_ ^ _24537_ /*888*/;
assign _24544_ = D[44] ^ Q[1] /*884*/;
assign _24541_ = _23913_ & _24544_ /*880*/;
assign _24542_ = _23913_ ^ _24544_ /*883*/;
assign _24543_ = _24535_ & _24542_ /*881*/;
assign _24540_ = _24541_ | _24543_ /*879*/;
assign _24299_ = _24535_ ^ _24542_ /*882*/;
assign _24549_ = D[45] ^ Q[1] /*878*/;
assign _24546_ = _23914_ & _24549_ /*874*/;
assign _24547_ = _23914_ ^ _24549_ /*877*/;
assign _24548_ = _24540_ & _24547_ /*875*/;
assign _24545_ = _24546_ | _24548_ /*873*/;
assign _24300_ = _24540_ ^ _24547_ /*876*/;
assign _24554_ = D[46] ^ Q[1] /*872*/;
assign _24551_ = _23915_ & _24554_ /*868*/;
assign _24552_ = _23915_ ^ _24554_ /*871*/;
assign _24553_ = _24545_ & _24552_ /*869*/;
assign _24550_ = _24551_ | _24553_ /*867*/;
assign _24301_ = _24545_ ^ _24552_ /*870*/;
assign _24559_ = D[47] ^ Q[1] /*866*/;
assign _24556_ = _23916_ & _24559_ /*862*/;
assign _24557_ = _23916_ ^ _24559_ /*865*/;
assign _24558_ = _24550_ & _24557_ /*863*/;
assign _24555_ = _24556_ | _24558_ /*861*/;
assign _24302_ = _24550_ ^ _24557_ /*864*/;
assign _24564_ = D[48] ^ Q[1] /*860*/;
assign _24561_ = _23917_ & _24564_ /*856*/;
assign _24562_ = _23917_ ^ _24564_ /*859*/;
assign _24563_ = _24555_ & _24562_ /*857*/;
assign _24560_ = _24561_ | _24563_ /*855*/;
assign _24303_ = _24555_ ^ _24562_ /*858*/;
assign _24569_ = D[49] ^ Q[1] /*854*/;
assign _24566_ = _23918_ & _24569_ /*850*/;
assign _24567_ = _23918_ ^ _24569_ /*853*/;
assign _24568_ = _24560_ & _24567_ /*851*/;
assign _24565_ = _24566_ | _24568_ /*849*/;
assign _24304_ = _24560_ ^ _24567_ /*852*/;
assign _24574_ = D[50] ^ Q[1] /*848*/;
assign _24571_ = _23919_ & _24574_ /*844*/;
assign _24572_ = _23919_ ^ _24574_ /*847*/;
assign _24573_ = _24565_ & _24572_ /*845*/;
assign _24570_ = _24571_ | _24573_ /*843*/;
assign _24305_ = _24565_ ^ _24572_ /*846*/;
assign _24579_ = D[51] ^ Q[1] /*842*/;
assign _24576_ = _23920_ & _24579_ /*838*/;
assign _24577_ = _23920_ ^ _24579_ /*841*/;
assign _24578_ = _24570_ & _24577_ /*839*/;
assign _24575_ = _24576_ | _24578_ /*837*/;
assign _24306_ = _24570_ ^ _24577_ /*840*/;
assign _24584_ = D[52] ^ Q[1] /*836*/;
assign _24581_ = _23921_ & _24584_ /*832*/;
assign _24582_ = _23921_ ^ _24584_ /*835*/;
assign _24583_ = _24575_ & _24582_ /*833*/;
assign _24580_ = _24581_ | _24583_ /*831*/;
assign _24307_ = _24575_ ^ _24582_ /*834*/;
assign _24589_ = D[53] ^ Q[1] /*830*/;
assign _24586_ = _23922_ & _24589_ /*826*/;
assign _24587_ = _23922_ ^ _24589_ /*829*/;
assign _24588_ = _24580_ & _24587_ /*827*/;
assign _24585_ = _24586_ | _24588_ /*825*/;
assign _24308_ = _24580_ ^ _24587_ /*828*/;
assign _24594_ = D[54] ^ Q[1] /*824*/;
assign _24591_ = _23923_ & _24594_ /*820*/;
assign _24592_ = _23923_ ^ _24594_ /*823*/;
assign _24593_ = _24585_ & _24592_ /*821*/;
assign _24590_ = _24591_ | _24593_ /*819*/;
assign _24309_ = _24585_ ^ _24592_ /*822*/;
assign _24599_ = D[55] ^ Q[1] /*818*/;
assign _24596_ = _23924_ & _24599_ /*814*/;
assign _24597_ = _23924_ ^ _24599_ /*817*/;
assign _24598_ = _24590_ & _24597_ /*815*/;
assign _24595_ = _24596_ | _24598_ /*813*/;
assign _24310_ = _24590_ ^ _24597_ /*816*/;
assign _24604_ = D[56] ^ Q[1] /*812*/;
assign _24601_ = _23925_ & _24604_ /*808*/;
assign _24602_ = _23925_ ^ _24604_ /*811*/;
assign _24603_ = _24595_ & _24602_ /*809*/;
assign _24600_ = _24601_ | _24603_ /*807*/;
assign _24311_ = _24595_ ^ _24602_ /*810*/;
assign _24609_ = D[57] ^ Q[1] /*806*/;
assign _24606_ = _23926_ & _24609_ /*802*/;
assign _24607_ = _23926_ ^ _24609_ /*805*/;
assign _24608_ = _24600_ & _24607_ /*803*/;
assign _24605_ = _24606_ | _24608_ /*801*/;
assign _24312_ = _24600_ ^ _24607_ /*804*/;
assign _24614_ = D[58] ^ Q[1] /*800*/;
assign _24611_ = _23927_ & _24614_ /*796*/;
assign _24612_ = _23927_ ^ _24614_ /*799*/;
assign _24613_ = _24605_ & _24612_ /*797*/;
assign _24610_ = _24611_ | _24613_ /*795*/;
assign _24313_ = _24605_ ^ _24612_ /*798*/;
assign _24619_ = D[59] ^ Q[1] /*794*/;
assign _24616_ = _23928_ & _24619_ /*790*/;
assign _24617_ = _23928_ ^ _24619_ /*793*/;
assign _24618_ = _24610_ & _24617_ /*791*/;
assign _24615_ = _24616_ | _24618_ /*789*/;
assign _24314_ = _24610_ ^ _24617_ /*792*/;
assign _24624_ = D[60] ^ Q[1] /*788*/;
assign _24621_ = _23929_ & _24624_ /*784*/;
assign _24622_ = _23929_ ^ _24624_ /*787*/;
assign _24623_ = _24615_ & _24622_ /*785*/;
assign _24620_ = _24621_ | _24623_ /*783*/;
assign _24315_ = _24615_ ^ _24622_ /*786*/;
assign _24629_ = D[61] ^ Q[1] /*782*/;
assign _24626_ = _23930_ & _24629_ /*778*/;
assign _24627_ = _23930_ ^ _24629_ /*781*/;
assign _24628_ = _24620_ & _24627_ /*779*/;
assign _24625_ = _24626_ | _24628_ /*777*/;
assign _24316_ = _24620_ ^ _24627_ /*780*/;
assign _24634_ = D[62] ^ Q[1] /*776*/;
assign _24631_ = _23931_ & _24634_ /*772*/;
assign _24632_ = _23931_ ^ _24634_ /*775*/;
assign _24633_ = _24625_ & _24632_ /*773*/;
assign _24630_ = _24631_ | _24633_ /*771*/;
assign _24317_ = _24625_ ^ _24632_ /*774*/;
assign _24638_ = zeroWire ^ Q[1] /*770*/;
assign _24635_ = _23932_ & _24638_ /*766*/;
assign _24636_ = _23932_ ^ _24638_ /*769*/;
assign _24637_ = _24630_ & _24636_ /*767*/;
assign Q[0] = _24635_ | _24637_ /*765*/;
assign _24318_ = _24630_ ^ _24636_ /*764*/;
assign _24640_ = ~Q[0] /*379*/;
assign _24641_ = _24640_ & D[0] /*378*/;
assign _24642_ = _24255_ & _24641_ /*376*/;
assign R_n1[0] = _24255_ ^ _24641_ /*377*/;
assign _24646_ = _24640_ & D[1] /*375*/;
assign _24648_ = _24256_ & _24646_ /*371*/;
assign _24649_ = _24256_ ^ _24646_ /*374*/;
assign _24650_ = _24642_ & _24649_ /*372*/;
assign _24647_ = _24648_ | _24650_ /*370*/;
assign R_n1[1] = _24642_ ^ _24649_ /*373*/;
assign _24651_ = _24640_ & D[2] /*369*/;
assign _24653_ = _24257_ & _24651_ /*365*/;
assign _24654_ = _24257_ ^ _24651_ /*368*/;
assign _24655_ = _24647_ & _24654_ /*366*/;
assign _24652_ = _24653_ | _24655_ /*364*/;
assign R_n1[2] = _24647_ ^ _24654_ /*367*/;
assign _24656_ = _24640_ & D[3] /*363*/;
assign _24658_ = _24258_ & _24656_ /*359*/;
assign _24659_ = _24258_ ^ _24656_ /*362*/;
assign _24660_ = _24652_ & _24659_ /*360*/;
assign _24657_ = _24658_ | _24660_ /*358*/;
assign R_n1[3] = _24652_ ^ _24659_ /*361*/;
assign _24661_ = _24640_ & D[4] /*357*/;
assign _24663_ = _24259_ & _24661_ /*353*/;
assign _24664_ = _24259_ ^ _24661_ /*356*/;
assign _24665_ = _24657_ & _24664_ /*354*/;
assign _24662_ = _24663_ | _24665_ /*352*/;
assign R_n1[4] = _24657_ ^ _24664_ /*355*/;
assign _24666_ = _24640_ & D[5] /*351*/;
assign _24668_ = _24260_ & _24666_ /*347*/;
assign _24669_ = _24260_ ^ _24666_ /*350*/;
assign _24670_ = _24662_ & _24669_ /*348*/;
assign _24667_ = _24668_ | _24670_ /*346*/;
assign R_n1[5] = _24662_ ^ _24669_ /*349*/;
assign _24671_ = _24640_ & D[6] /*345*/;
assign _24673_ = _24261_ & _24671_ /*341*/;
assign _24674_ = _24261_ ^ _24671_ /*344*/;
assign _24675_ = _24667_ & _24674_ /*342*/;
assign _24672_ = _24673_ | _24675_ /*340*/;
assign R_n1[6] = _24667_ ^ _24674_ /*343*/;
assign _24676_ = _24640_ & D[7] /*339*/;
assign _24678_ = _24262_ & _24676_ /*335*/;
assign _24679_ = _24262_ ^ _24676_ /*338*/;
assign _24680_ = _24672_ & _24679_ /*336*/;
assign _24677_ = _24678_ | _24680_ /*334*/;
assign R_n1[7] = _24672_ ^ _24679_ /*337*/;
assign _24681_ = _24640_ & D[8] /*333*/;
assign _24683_ = _24263_ & _24681_ /*329*/;
assign _24684_ = _24263_ ^ _24681_ /*332*/;
assign _24685_ = _24677_ & _24684_ /*330*/;
assign _24682_ = _24683_ | _24685_ /*328*/;
assign R_n1[8] = _24677_ ^ _24684_ /*331*/;
assign _24686_ = _24640_ & D[9] /*327*/;
assign _24688_ = _24264_ & _24686_ /*323*/;
assign _24689_ = _24264_ ^ _24686_ /*326*/;
assign _24690_ = _24682_ & _24689_ /*324*/;
assign _24687_ = _24688_ | _24690_ /*322*/;
assign R_n1[9] = _24682_ ^ _24689_ /*325*/;
assign _24691_ = _24640_ & D[10] /*321*/;
assign _24693_ = _24265_ & _24691_ /*317*/;
assign _24694_ = _24265_ ^ _24691_ /*320*/;
assign _24695_ = _24687_ & _24694_ /*318*/;
assign _24692_ = _24693_ | _24695_ /*316*/;
assign R_n1[10] = _24687_ ^ _24694_ /*319*/;
assign _24696_ = _24640_ & D[11] /*315*/;
assign _24698_ = _24266_ & _24696_ /*311*/;
assign _24699_ = _24266_ ^ _24696_ /*314*/;
assign _24700_ = _24692_ & _24699_ /*312*/;
assign _24697_ = _24698_ | _24700_ /*310*/;
assign R_n1[11] = _24692_ ^ _24699_ /*313*/;
assign _24701_ = _24640_ & D[12] /*309*/;
assign _24703_ = _24267_ & _24701_ /*305*/;
assign _24704_ = _24267_ ^ _24701_ /*308*/;
assign _24705_ = _24697_ & _24704_ /*306*/;
assign _24702_ = _24703_ | _24705_ /*304*/;
assign R_n1[12] = _24697_ ^ _24704_ /*307*/;
assign _24706_ = _24640_ & D[13] /*303*/;
assign _24708_ = _24268_ & _24706_ /*299*/;
assign _24709_ = _24268_ ^ _24706_ /*302*/;
assign _24710_ = _24702_ & _24709_ /*300*/;
assign _24707_ = _24708_ | _24710_ /*298*/;
assign R_n1[13] = _24702_ ^ _24709_ /*301*/;
assign _24711_ = _24640_ & D[14] /*297*/;
assign _24713_ = _24269_ & _24711_ /*293*/;
assign _24714_ = _24269_ ^ _24711_ /*296*/;
assign _24715_ = _24707_ & _24714_ /*294*/;
assign _24712_ = _24713_ | _24715_ /*292*/;
assign R_n1[14] = _24707_ ^ _24714_ /*295*/;
assign _24716_ = _24640_ & D[15] /*291*/;
assign _24718_ = _24270_ & _24716_ /*287*/;
assign _24719_ = _24270_ ^ _24716_ /*290*/;
assign _24720_ = _24712_ & _24719_ /*288*/;
assign _24717_ = _24718_ | _24720_ /*286*/;
assign R_n1[15] = _24712_ ^ _24719_ /*289*/;
assign _24721_ = _24640_ & D[16] /*285*/;
assign _24723_ = _24271_ & _24721_ /*281*/;
assign _24724_ = _24271_ ^ _24721_ /*284*/;
assign _24725_ = _24717_ & _24724_ /*282*/;
assign _24722_ = _24723_ | _24725_ /*280*/;
assign R_n1[16] = _24717_ ^ _24724_ /*283*/;
assign _24726_ = _24640_ & D[17] /*279*/;
assign _24728_ = _24272_ & _24726_ /*275*/;
assign _24729_ = _24272_ ^ _24726_ /*278*/;
assign _24730_ = _24722_ & _24729_ /*276*/;
assign _24727_ = _24728_ | _24730_ /*274*/;
assign R_n1[17] = _24722_ ^ _24729_ /*277*/;
assign _24731_ = _24640_ & D[18] /*273*/;
assign _24733_ = _24273_ & _24731_ /*269*/;
assign _24734_ = _24273_ ^ _24731_ /*272*/;
assign _24735_ = _24727_ & _24734_ /*270*/;
assign _24732_ = _24733_ | _24735_ /*268*/;
assign R_n1[18] = _24727_ ^ _24734_ /*271*/;
assign _24736_ = _24640_ & D[19] /*267*/;
assign _24738_ = _24274_ & _24736_ /*263*/;
assign _24739_ = _24274_ ^ _24736_ /*266*/;
assign _24740_ = _24732_ & _24739_ /*264*/;
assign _24737_ = _24738_ | _24740_ /*262*/;
assign R_n1[19] = _24732_ ^ _24739_ /*265*/;
assign _24741_ = _24640_ & D[20] /*261*/;
assign _24743_ = _24275_ & _24741_ /*257*/;
assign _24744_ = _24275_ ^ _24741_ /*260*/;
assign _24745_ = _24737_ & _24744_ /*258*/;
assign _24742_ = _24743_ | _24745_ /*256*/;
assign R_n1[20] = _24737_ ^ _24744_ /*259*/;
assign _24746_ = _24640_ & D[21] /*255*/;
assign _24748_ = _24276_ & _24746_ /*251*/;
assign _24749_ = _24276_ ^ _24746_ /*254*/;
assign _24750_ = _24742_ & _24749_ /*252*/;
assign _24747_ = _24748_ | _24750_ /*250*/;
assign R_n1[21] = _24742_ ^ _24749_ /*253*/;
assign _24751_ = _24640_ & D[22] /*249*/;
assign _24753_ = _24277_ & _24751_ /*245*/;
assign _24754_ = _24277_ ^ _24751_ /*248*/;
assign _24755_ = _24747_ & _24754_ /*246*/;
assign _24752_ = _24753_ | _24755_ /*244*/;
assign R_n1[22] = _24747_ ^ _24754_ /*247*/;
assign _24756_ = _24640_ & D[23] /*243*/;
assign _24758_ = _24278_ & _24756_ /*239*/;
assign _24759_ = _24278_ ^ _24756_ /*242*/;
assign _24760_ = _24752_ & _24759_ /*240*/;
assign _24757_ = _24758_ | _24760_ /*238*/;
assign R_n1[23] = _24752_ ^ _24759_ /*241*/;
assign _24761_ = _24640_ & D[24] /*237*/;
assign _24763_ = _24279_ & _24761_ /*233*/;
assign _24764_ = _24279_ ^ _24761_ /*236*/;
assign _24765_ = _24757_ & _24764_ /*234*/;
assign _24762_ = _24763_ | _24765_ /*232*/;
assign R_n1[24] = _24757_ ^ _24764_ /*235*/;
assign _24766_ = _24640_ & D[25] /*231*/;
assign _24768_ = _24280_ & _24766_ /*227*/;
assign _24769_ = _24280_ ^ _24766_ /*230*/;
assign _24770_ = _24762_ & _24769_ /*228*/;
assign _24767_ = _24768_ | _24770_ /*226*/;
assign R_n1[25] = _24762_ ^ _24769_ /*229*/;
assign _24771_ = _24640_ & D[26] /*225*/;
assign _24773_ = _24281_ & _24771_ /*221*/;
assign _24774_ = _24281_ ^ _24771_ /*224*/;
assign _24775_ = _24767_ & _24774_ /*222*/;
assign _24772_ = _24773_ | _24775_ /*220*/;
assign R_n1[26] = _24767_ ^ _24774_ /*223*/;
assign _24776_ = _24640_ & D[27] /*219*/;
assign _24778_ = _24282_ & _24776_ /*215*/;
assign _24779_ = _24282_ ^ _24776_ /*218*/;
assign _24780_ = _24772_ & _24779_ /*216*/;
assign _24777_ = _24778_ | _24780_ /*214*/;
assign R_n1[27] = _24772_ ^ _24779_ /*217*/;
assign _24781_ = _24640_ & D[28] /*213*/;
assign _24783_ = _24283_ & _24781_ /*209*/;
assign _24784_ = _24283_ ^ _24781_ /*212*/;
assign _24785_ = _24777_ & _24784_ /*210*/;
assign _24782_ = _24783_ | _24785_ /*208*/;
assign R_n1[28] = _24777_ ^ _24784_ /*211*/;
assign _24786_ = _24640_ & D[29] /*207*/;
assign _24788_ = _24284_ & _24786_ /*203*/;
assign _24789_ = _24284_ ^ _24786_ /*206*/;
assign _24790_ = _24782_ & _24789_ /*204*/;
assign _24787_ = _24788_ | _24790_ /*202*/;
assign R_n1[29] = _24782_ ^ _24789_ /*205*/;
assign _24791_ = _24640_ & D[30] /*201*/;
assign _24793_ = _24285_ & _24791_ /*197*/;
assign _24794_ = _24285_ ^ _24791_ /*200*/;
assign _24795_ = _24787_ & _24794_ /*198*/;
assign _24792_ = _24793_ | _24795_ /*196*/;
assign R_n1[30] = _24787_ ^ _24794_ /*199*/;
assign _24796_ = _24640_ & D[31] /*195*/;
assign _24798_ = _24286_ & _24796_ /*191*/;
assign _24799_ = _24286_ ^ _24796_ /*194*/;
assign _24800_ = _24792_ & _24799_ /*192*/;
assign _24797_ = _24798_ | _24800_ /*190*/;
assign R_n1[31] = _24792_ ^ _24799_ /*193*/;
assign _24801_ = _24640_ & D[32] /*189*/;
assign _24803_ = _24287_ & _24801_ /*185*/;
assign _24804_ = _24287_ ^ _24801_ /*188*/;
assign _24805_ = _24797_ & _24804_ /*186*/;
assign _24802_ = _24803_ | _24805_ /*184*/;
assign R_n1[32] = _24797_ ^ _24804_ /*187*/;
assign _24806_ = _24640_ & D[33] /*183*/;
assign _24808_ = _24288_ & _24806_ /*179*/;
assign _24809_ = _24288_ ^ _24806_ /*182*/;
assign _24810_ = _24802_ & _24809_ /*180*/;
assign _24807_ = _24808_ | _24810_ /*178*/;
assign R_n1[33] = _24802_ ^ _24809_ /*181*/;
assign _24811_ = _24640_ & D[34] /*177*/;
assign _24813_ = _24289_ & _24811_ /*173*/;
assign _24814_ = _24289_ ^ _24811_ /*176*/;
assign _24815_ = _24807_ & _24814_ /*174*/;
assign _24812_ = _24813_ | _24815_ /*172*/;
assign R_n1[34] = _24807_ ^ _24814_ /*175*/;
assign _24816_ = _24640_ & D[35] /*171*/;
assign _24818_ = _24290_ & _24816_ /*167*/;
assign _24819_ = _24290_ ^ _24816_ /*170*/;
assign _24820_ = _24812_ & _24819_ /*168*/;
assign _24817_ = _24818_ | _24820_ /*166*/;
assign R_n1[35] = _24812_ ^ _24819_ /*169*/;
assign _24821_ = _24640_ & D[36] /*165*/;
assign _24823_ = _24291_ & _24821_ /*161*/;
assign _24824_ = _24291_ ^ _24821_ /*164*/;
assign _24825_ = _24817_ & _24824_ /*162*/;
assign _24822_ = _24823_ | _24825_ /*160*/;
assign R_n1[36] = _24817_ ^ _24824_ /*163*/;
assign _24826_ = _24640_ & D[37] /*159*/;
assign _24828_ = _24292_ & _24826_ /*155*/;
assign _24829_ = _24292_ ^ _24826_ /*158*/;
assign _24830_ = _24822_ & _24829_ /*156*/;
assign _24827_ = _24828_ | _24830_ /*154*/;
assign R_n1[37] = _24822_ ^ _24829_ /*157*/;
assign _24831_ = _24640_ & D[38] /*153*/;
assign _24833_ = _24293_ & _24831_ /*149*/;
assign _24834_ = _24293_ ^ _24831_ /*152*/;
assign _24835_ = _24827_ & _24834_ /*150*/;
assign _24832_ = _24833_ | _24835_ /*148*/;
assign R_n1[38] = _24827_ ^ _24834_ /*151*/;
assign _24836_ = _24640_ & D[39] /*147*/;
assign _24838_ = _24294_ & _24836_ /*143*/;
assign _24839_ = _24294_ ^ _24836_ /*146*/;
assign _24840_ = _24832_ & _24839_ /*144*/;
assign _24837_ = _24838_ | _24840_ /*142*/;
assign R_n1[39] = _24832_ ^ _24839_ /*145*/;
assign _24841_ = _24640_ & D[40] /*141*/;
assign _24843_ = _24295_ & _24841_ /*137*/;
assign _24844_ = _24295_ ^ _24841_ /*140*/;
assign _24845_ = _24837_ & _24844_ /*138*/;
assign _24842_ = _24843_ | _24845_ /*136*/;
assign R_n1[40] = _24837_ ^ _24844_ /*139*/;
assign _24846_ = _24640_ & D[41] /*135*/;
assign _24848_ = _24296_ & _24846_ /*131*/;
assign _24849_ = _24296_ ^ _24846_ /*134*/;
assign _24850_ = _24842_ & _24849_ /*132*/;
assign _24847_ = _24848_ | _24850_ /*130*/;
assign R_n1[41] = _24842_ ^ _24849_ /*133*/;
assign _24851_ = _24640_ & D[42] /*129*/;
assign _24853_ = _24297_ & _24851_ /*125*/;
assign _24854_ = _24297_ ^ _24851_ /*128*/;
assign _24855_ = _24847_ & _24854_ /*126*/;
assign _24852_ = _24853_ | _24855_ /*124*/;
assign R_n1[42] = _24847_ ^ _24854_ /*127*/;
assign _24856_ = _24640_ & D[43] /*123*/;
assign _24858_ = _24298_ & _24856_ /*119*/;
assign _24859_ = _24298_ ^ _24856_ /*122*/;
assign _24860_ = _24852_ & _24859_ /*120*/;
assign _24857_ = _24858_ | _24860_ /*118*/;
assign R_n1[43] = _24852_ ^ _24859_ /*121*/;
assign _24861_ = _24640_ & D[44] /*117*/;
assign _24863_ = _24299_ & _24861_ /*113*/;
assign _24864_ = _24299_ ^ _24861_ /*116*/;
assign _24865_ = _24857_ & _24864_ /*114*/;
assign _24862_ = _24863_ | _24865_ /*112*/;
assign R_n1[44] = _24857_ ^ _24864_ /*115*/;
assign _24866_ = _24640_ & D[45] /*111*/;
assign _24868_ = _24300_ & _24866_ /*107*/;
assign _24869_ = _24300_ ^ _24866_ /*110*/;
assign _24870_ = _24862_ & _24869_ /*108*/;
assign _24867_ = _24868_ | _24870_ /*106*/;
assign R_n1[45] = _24862_ ^ _24869_ /*109*/;
assign _24871_ = _24640_ & D[46] /*105*/;
assign _24873_ = _24301_ & _24871_ /*101*/;
assign _24874_ = _24301_ ^ _24871_ /*104*/;
assign _24875_ = _24867_ & _24874_ /*102*/;
assign _24872_ = _24873_ | _24875_ /*100*/;
assign R_n1[46] = _24867_ ^ _24874_ /*103*/;
assign _24876_ = _24640_ & D[47] /*99*/;
assign _24878_ = _24302_ & _24876_ /*95*/;
assign _24879_ = _24302_ ^ _24876_ /*98*/;
assign _24880_ = _24872_ & _24879_ /*96*/;
assign _24877_ = _24878_ | _24880_ /*94*/;
assign R_n1[47] = _24872_ ^ _24879_ /*97*/;
assign _24881_ = _24640_ & D[48] /*93*/;
assign _24883_ = _24303_ & _24881_ /*89*/;
assign _24884_ = _24303_ ^ _24881_ /*92*/;
assign _24885_ = _24877_ & _24884_ /*90*/;
assign _24882_ = _24883_ | _24885_ /*88*/;
assign R_n1[48] = _24877_ ^ _24884_ /*91*/;
assign _24886_ = _24640_ & D[49] /*87*/;
assign _24888_ = _24304_ & _24886_ /*83*/;
assign _24889_ = _24304_ ^ _24886_ /*86*/;
assign _24890_ = _24882_ & _24889_ /*84*/;
assign _24887_ = _24888_ | _24890_ /*82*/;
assign R_n1[49] = _24882_ ^ _24889_ /*85*/;
assign _24891_ = _24640_ & D[50] /*81*/;
assign _24893_ = _24305_ & _24891_ /*77*/;
assign _24894_ = _24305_ ^ _24891_ /*80*/;
assign _24895_ = _24887_ & _24894_ /*78*/;
assign _24892_ = _24893_ | _24895_ /*76*/;
assign R_n1[50] = _24887_ ^ _24894_ /*79*/;
assign _24896_ = _24640_ & D[51] /*75*/;
assign _24898_ = _24306_ & _24896_ /*71*/;
assign _24899_ = _24306_ ^ _24896_ /*74*/;
assign _24900_ = _24892_ & _24899_ /*72*/;
assign _24897_ = _24898_ | _24900_ /*70*/;
assign R_n1[51] = _24892_ ^ _24899_ /*73*/;
assign _24901_ = _24640_ & D[52] /*69*/;
assign _24903_ = _24307_ & _24901_ /*65*/;
assign _24904_ = _24307_ ^ _24901_ /*68*/;
assign _24905_ = _24897_ & _24904_ /*66*/;
assign _24902_ = _24903_ | _24905_ /*64*/;
assign R_n1[52] = _24897_ ^ _24904_ /*67*/;
assign _24906_ = _24640_ & D[53] /*63*/;
assign _24908_ = _24308_ & _24906_ /*59*/;
assign _24909_ = _24308_ ^ _24906_ /*62*/;
assign _24910_ = _24902_ & _24909_ /*60*/;
assign _24907_ = _24908_ | _24910_ /*58*/;
assign R_n1[53] = _24902_ ^ _24909_ /*61*/;
assign _24911_ = _24640_ & D[54] /*57*/;
assign _24913_ = _24309_ & _24911_ /*53*/;
assign _24914_ = _24309_ ^ _24911_ /*56*/;
assign _24915_ = _24907_ & _24914_ /*54*/;
assign _24912_ = _24913_ | _24915_ /*52*/;
assign R_n1[54] = _24907_ ^ _24914_ /*55*/;
assign _24916_ = _24640_ & D[55] /*51*/;
assign _24918_ = _24310_ & _24916_ /*47*/;
assign _24919_ = _24310_ ^ _24916_ /*50*/;
assign _24920_ = _24912_ & _24919_ /*48*/;
assign _24917_ = _24918_ | _24920_ /*46*/;
assign R_n1[55] = _24912_ ^ _24919_ /*49*/;
assign _24921_ = _24640_ & D[56] /*45*/;
assign _24923_ = _24311_ & _24921_ /*41*/;
assign _24924_ = _24311_ ^ _24921_ /*44*/;
assign _24925_ = _24917_ & _24924_ /*42*/;
assign _24922_ = _24923_ | _24925_ /*40*/;
assign R_n1[56] = _24917_ ^ _24924_ /*43*/;
assign _24926_ = _24640_ & D[57] /*39*/;
assign _24928_ = _24312_ & _24926_ /*35*/;
assign _24929_ = _24312_ ^ _24926_ /*38*/;
assign _24930_ = _24922_ & _24929_ /*36*/;
assign _24927_ = _24928_ | _24930_ /*34*/;
assign R_n1[57] = _24922_ ^ _24929_ /*37*/;
assign _24931_ = _24640_ & D[58] /*33*/;
assign _24933_ = _24313_ & _24931_ /*29*/;
assign _24934_ = _24313_ ^ _24931_ /*32*/;
assign _24935_ = _24927_ & _24934_ /*30*/;
assign _24932_ = _24933_ | _24935_ /*28*/;
assign R_n1[58] = _24927_ ^ _24934_ /*31*/;
assign _24936_ = _24640_ & D[59] /*27*/;
assign _24938_ = _24314_ & _24936_ /*23*/;
assign _24939_ = _24314_ ^ _24936_ /*26*/;
assign _24940_ = _24932_ & _24939_ /*24*/;
assign _24937_ = _24938_ | _24940_ /*22*/;
assign R_n1[59] = _24932_ ^ _24939_ /*25*/;
assign _24941_ = _24640_ & D[60] /*21*/;
assign _24943_ = _24315_ & _24941_ /*17*/;
assign _24944_ = _24315_ ^ _24941_ /*20*/;
assign _24945_ = _24937_ & _24944_ /*18*/;
assign _24942_ = _24943_ | _24945_ /*16*/;
assign R_n1[60] = _24937_ ^ _24944_ /*19*/;
assign _24946_ = _24640_ & D[61] /*15*/;
assign _24948_ = _24316_ & _24946_ /*11*/;
assign _24949_ = _24316_ ^ _24946_ /*14*/;
assign _24950_ = _24942_ & _24949_ /*12*/;
assign _24947_ = _24948_ | _24950_ /*10*/;
assign R_n1[61] = _24942_ ^ _24949_ /*13*/;
assign _24951_ = _24640_ & D[62] /*9*/;
assign _24953_ = _24317_ & _24951_ /*5*/;
assign _24954_ = _24317_ ^ _24951_ /*8*/;
assign _24955_ = _24947_ & _24954_ /*6*/;
assign _24952_ = _24953_ | _24955_ /*4*/;
assign R_n1[62] = _24947_ ^ _24954_ /*7*/;
assign _24956_ = _24640_ & zeroWire /*3*/;
assign _24957_ = _24318_ ^ _24956_ /*2*/;
assign R_n1[63] = _24957_ ^ _24952_ /*1*/;
endmodule
