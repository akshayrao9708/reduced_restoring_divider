module nonresdivReduced(R_0, D, Q, R_n1);
input [5:0] R_0;
input [2:0] D;
output [3:0] Q;
output [3:0] R_n1;
wire _0_;
wire _1_;
wire _2_;
wire _3_;
wire _4_;
wire _5_;
wire _6_;
wire _7_;
wire _8_;
wire _9_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire _30_;
wire _31_;
wire _32_;
wire _33_;
wire _34_;
wire _35_;
wire _36_;
wire _37_;
wire _38_;
wire _39_;
wire _40_;
wire _41_;
wire _42_;
wire _43_;
wire _44_;
wire _45_;
wire _46_;
wire _47_;
wire _48_;
wire _49_;
wire _50_;
wire _51_;
wire _52_;
wire _53_;
wire _54_;
wire _55_;
wire _56_;
wire _57_;
wire _58_;
wire _59_;
wire _60_;
wire _61_;
wire _62_;
wire _63_;
wire _64_;
wire _65_;
wire _66_;
wire _67_;
wire _68_;
wire _69_;
wire _70_;
wire _71_;
wire _72_;
wire _73_;
wire _74_;
wire _75_;
wire _76_;
wire _77_;
wire _78_;
wire _79_;
wire _80_;
wire _81_;
wire _82_;
wire _83_;
wire _84_;
wire _85_;
wire _86_;
wire _87_;
wire _88_;
wire _89_;
wire _90_;
wire _91_;
wire _92_;
wire _93_;
wire _94_;
wire _95_;
wire _96_;
wire _97_;
wire _98_;
wire _99_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire zeroWire;
wire oneWire;
assign zeroWire = 1'b0 /*239*/;
assign oneWire = 1'b1 /*239*/;
assign _7_ = ~D[0] /*213*/;
assign _5_ = R_0[3] | _7_ /*210*/;
assign _6_ = R_0[3] ^ _7_ /*212*/;
assign _0_ = ~_6_ /*211*/;
assign _14_ = ~D[1] /*209*/;
assign _11_ = R_0[4] & _14_ /*205*/;
assign _12_ = R_0[4] ^ _14_ /*208*/;
assign _13_ = _5_ & _12_ /*206*/;
assign _10_ = _11_ | _13_ /*204*/;
assign _1_ = _5_ ^ _12_ /*207*/;
assign _19_ = ~D[2] /*203*/;
assign _16_ = R_0[5] & _19_ /*199*/;
assign _17_ = R_0[5] ^ _19_ /*202*/;
assign _18_ = _10_ & _17_ /*200*/;
assign _15_ = _16_ | _18_ /*198*/;
assign _2_ = _10_ ^ _17_ /*201*/;
assign _20_ = zeroWire & oneWire /*193*/;
assign _21_ = zeroWire ^ oneWire /*196*/;
assign _22_ = _15_ & _21_ /*194*/;
assign Q[3] = _20_ | _22_ /*192*/;
assign _3_ = _15_ ^ _21_ /*195*/;
assign _34_ = D[0] ^ Q[3] /*166*/;
assign _31_ = R_0[2] & _34_ /*162*/;
assign _32_ = R_0[2] ^ _34_ /*165*/;
assign _33_ = Q[3] & _32_ /*163*/;
assign _30_ = _31_ | _33_ /*161*/;
assign _25_ = Q[3] ^ _32_ /*164*/;
assign _39_ = D[1] ^ Q[3] /*160*/;
assign _36_ = _0_ & _39_ /*156*/;
assign _37_ = _0_ ^ _39_ /*159*/;
assign _38_ = _30_ & _37_ /*157*/;
assign _35_ = _36_ | _38_ /*155*/;
assign _26_ = _30_ ^ _37_ /*158*/;
assign _44_ = D[2] ^ Q[3] /*154*/;
assign _41_ = _1_ & _44_ /*150*/;
assign _42_ = _1_ ^ _44_ /*153*/;
assign _43_ = _35_ & _42_ /*151*/;
assign _40_ = _41_ | _43_ /*149*/;
assign _27_ = _35_ ^ _42_ /*152*/;
assign _48_ = zeroWire ^ Q[3] /*148*/;
assign _45_ = _2_ & _48_ /*144*/;
assign _46_ = _2_ ^ _48_ /*147*/;
assign _47_ = _40_ & _46_ /*145*/;
assign Q[2] = _45_ | _47_ /*143*/;
assign _28_ = _40_ ^ _46_ /*146*/;
assign _59_ = D[0] ^ Q[2] /*117*/;
assign _56_ = R_0[1] & _59_ /*113*/;
assign _57_ = R_0[1] ^ _59_ /*116*/;
assign _58_ = Q[2] & _57_ /*114*/;
assign _55_ = _56_ | _58_ /*112*/;
assign _50_ = Q[2] ^ _57_ /*115*/;
assign _64_ = D[1] ^ Q[2] /*111*/;
assign _61_ = _25_ & _64_ /*107*/;
assign _62_ = _25_ ^ _64_ /*110*/;
assign _63_ = _55_ & _62_ /*108*/;
assign _60_ = _61_ | _63_ /*106*/;
assign _51_ = _55_ ^ _62_ /*109*/;
assign _69_ = D[2] ^ Q[2] /*105*/;
assign _66_ = _26_ & _69_ /*101*/;
assign _67_ = _26_ ^ _69_ /*104*/;
assign _68_ = _60_ & _67_ /*102*/;
assign _65_ = _66_ | _68_ /*100*/;
assign _52_ = _60_ ^ _67_ /*103*/;
assign _73_ = zeroWire ^ Q[2] /*99*/;
assign _70_ = _27_ & _73_ /*95*/;
assign _71_ = _27_ ^ _73_ /*98*/;
assign _72_ = _65_ & _71_ /*96*/;
assign Q[1] = _70_ | _72_ /*94*/;
assign _53_ = _65_ ^ _71_ /*97*/;
assign _84_ = D[0] ^ Q[1] /*68*/;
assign _81_ = R_0[0] & _84_ /*64*/;
assign _82_ = R_0[0] ^ _84_ /*67*/;
assign _83_ = Q[1] & _82_ /*65*/;
assign _80_ = _81_ | _83_ /*63*/;
assign _75_ = Q[1] ^ _82_ /*66*/;
assign _89_ = D[1] ^ Q[1] /*62*/;
assign _86_ = _50_ & _89_ /*58*/;
assign _87_ = _50_ ^ _89_ /*61*/;
assign _88_ = _80_ & _87_ /*59*/;
assign _85_ = _86_ | _88_ /*57*/;
assign _76_ = _80_ ^ _87_ /*60*/;
assign _94_ = D[2] ^ Q[1] /*56*/;
assign _91_ = _51_ & _94_ /*52*/;
assign _92_ = _51_ ^ _94_ /*55*/;
assign _93_ = _85_ & _92_ /*53*/;
assign _90_ = _91_ | _93_ /*51*/;
assign _77_ = _85_ ^ _92_ /*54*/;
assign _98_ = zeroWire ^ Q[1] /*50*/;
assign _95_ = _52_ & _98_ /*46*/;
assign _96_ = _52_ ^ _98_ /*49*/;
assign _97_ = _90_ & _96_ /*47*/;
assign Q[0] = _95_ | _97_ /*45*/;
assign _78_ = _90_ ^ _96_ /*44*/;
assign _100_ = ~Q[0] /*19*/;
assign _101_ = _100_ & D[0] /*18*/;
assign _102_ = _75_ & _101_ /*16*/;
assign R_n1[0] = _75_ ^ _101_ /*17*/;
assign _106_ = _100_ & D[1] /*15*/;
assign _108_ = _76_ & _106_ /*11*/;
assign _109_ = _76_ ^ _106_ /*14*/;
assign _110_ = _102_ & _109_ /*12*/;
assign _107_ = _108_ | _110_ /*10*/;
assign R_n1[1] = _102_ ^ _109_ /*13*/;
assign _111_ = _100_ & D[2] /*9*/;
assign _113_ = _77_ & _111_ /*5*/;
assign _114_ = _77_ ^ _111_ /*8*/;
assign _115_ = _107_ & _114_ /*6*/;
assign _112_ = _113_ | _115_ /*4*/;
assign R_n1[2] = _107_ ^ _114_ /*7*/;
assign _116_ = _100_ & zeroWire /*3*/;
assign _117_ = _78_ ^ _116_ /*2*/;
assign R_n1[3] = _117_ ^ _112_ /*1*/;
endmodule
