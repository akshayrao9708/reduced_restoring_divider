module divider(R_0, D, Q, R_n1);
input [125:0] R_0;
input [62:0] D;
output [63:0] Q;
output [62:0] R_n1;
wire _0_;
wire _1_;
wire _2_;
wire _3_;
wire _4_;
wire _5_;
wire _6_;
wire _7_;
wire _8_;
wire _9_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire _30_;
wire _31_;
wire _32_;
wire _33_;
wire _34_;
wire _35_;
wire _36_;
wire _37_;
wire _38_;
wire _39_;
wire _40_;
wire _41_;
wire _42_;
wire _43_;
wire _44_;
wire _45_;
wire _46_;
wire _47_;
wire _48_;
wire _49_;
wire _50_;
wire _51_;
wire _52_;
wire _53_;
wire _54_;
wire _55_;
wire _56_;
wire _57_;
wire _58_;
wire _59_;
wire _60_;
wire _61_;
wire _62_;
wire _63_;
wire _64_;
wire _65_;
wire _66_;
wire _67_;
wire _68_;
wire _69_;
wire _70_;
wire _71_;
wire _72_;
wire _73_;
wire _74_;
wire _75_;
wire _76_;
wire _77_;
wire _78_;
wire _79_;
wire _80_;
wire _81_;
wire _82_;
wire _83_;
wire _84_;
wire _85_;
wire _86_;
wire _87_;
wire _88_;
wire _89_;
wire _90_;
wire _91_;
wire _92_;
wire _93_;
wire _94_;
wire _95_;
wire _96_;
wire _97_;
wire _98_;
wire _99_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
wire _255_;
wire _256_;
wire _257_;
wire _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire _267_;
wire _268_;
wire _269_;
wire _270_;
wire _271_;
wire _272_;
wire _273_;
wire _274_;
wire _275_;
wire _276_;
wire _277_;
wire _278_;
wire _279_;
wire _280_;
wire _281_;
wire _282_;
wire _283_;
wire _284_;
wire _285_;
wire _286_;
wire _287_;
wire _288_;
wire _289_;
wire _290_;
wire _291_;
wire _292_;
wire _293_;
wire _294_;
wire _295_;
wire _296_;
wire _297_;
wire _298_;
wire _299_;
wire _300_;
wire _301_;
wire _302_;
wire _303_;
wire _304_;
wire _305_;
wire _306_;
wire _307_;
wire _308_;
wire _309_;
wire _310_;
wire _311_;
wire _312_;
wire _313_;
wire _314_;
wire _315_;
wire _316_;
wire _317_;
wire _318_;
wire _319_;
wire _320_;
wire _321_;
wire _322_;
wire _323_;
wire _324_;
wire _325_;
wire _326_;
wire _327_;
wire _328_;
wire _329_;
wire _330_;
wire _331_;
wire _332_;
wire _333_;
wire _334_;
wire _335_;
wire _336_;
wire _337_;
wire _338_;
wire _339_;
wire _340_;
wire _341_;
wire _342_;
wire _343_;
wire _344_;
wire _345_;
wire _346_;
wire _347_;
wire _348_;
wire _349_;
wire _350_;
wire _351_;
wire _352_;
wire _353_;
wire _354_;
wire _355_;
wire _356_;
wire _357_;
wire _358_;
wire _359_;
wire _360_;
wire _361_;
wire _362_;
wire _363_;
wire _364_;
wire _365_;
wire _366_;
wire _367_;
wire _368_;
wire _369_;
wire _370_;
wire _371_;
wire _372_;
wire _373_;
wire _374_;
wire _375_;
wire _376_;
wire _377_;
wire _378_;
wire _379_;
wire _380_;
wire _381_;
wire _382_;
wire _383_;
wire _384_;
wire _385_;
wire _386_;
wire _387_;
wire _388_;
wire _389_;
wire _390_;
wire _391_;
wire _392_;
wire _393_;
wire _394_;
wire _395_;
wire _396_;
wire _397_;
wire _398_;
wire _399_;
wire _400_;
wire _401_;
wire _402_;
wire _403_;
wire _404_;
wire _405_;
wire _406_;
wire _407_;
wire _408_;
wire _409_;
wire _410_;
wire _411_;
wire _412_;
wire _413_;
wire _414_;
wire _415_;
wire _416_;
wire _417_;
wire _418_;
wire _419_;
wire _420_;
wire _421_;
wire _422_;
wire _423_;
wire _424_;
wire _425_;
wire _426_;
wire _427_;
wire _428_;
wire _429_;
wire _430_;
wire _431_;
wire _432_;
wire _433_;
wire _434_;
wire _435_;
wire _436_;
wire _437_;
wire _438_;
wire _439_;
wire _440_;
wire _441_;
wire _442_;
wire _443_;
wire _444_;
wire _445_;
wire _446_;
wire _447_;
wire _448_;
wire _449_;
wire _450_;
wire _451_;
wire _452_;
wire _453_;
wire _454_;
wire _455_;
wire _456_;
wire _457_;
wire _458_;
wire _459_;
wire _460_;
wire _461_;
wire _462_;
wire _463_;
wire _464_;
wire _465_;
wire _466_;
wire _467_;
wire _468_;
wire _469_;
wire _470_;
wire _471_;
wire _472_;
wire _473_;
wire _474_;
wire _475_;
wire _476_;
wire _477_;
wire _478_;
wire _479_;
wire _480_;
wire _481_;
wire _482_;
wire _483_;
wire _484_;
wire _485_;
wire _486_;
wire _487_;
wire _488_;
wire _489_;
wire _490_;
wire _491_;
wire _492_;
wire _493_;
wire _494_;
wire _495_;
wire _496_;
wire _497_;
wire _498_;
wire _499_;
wire _500_;
wire _501_;
wire _502_;
wire _503_;
wire _504_;
wire _505_;
wire _506_;
wire _507_;
wire _508_;
wire _509_;
wire _510_;
wire _511_;
wire _512_;
wire _513_;
wire _514_;
wire _515_;
wire _516_;
wire _517_;
wire _518_;
wire _519_;
wire _520_;
wire _521_;
wire _522_;
wire _523_;
wire _524_;
wire _525_;
wire _526_;
wire _527_;
wire _528_;
wire _529_;
wire _530_;
wire _531_;
wire _532_;
wire _533_;
wire _534_;
wire _535_;
wire _536_;
wire _537_;
wire _538_;
wire _539_;
wire _540_;
wire _541_;
wire _542_;
wire _543_;
wire _544_;
wire _545_;
wire _546_;
wire _547_;
wire _548_;
wire _549_;
wire _550_;
wire _551_;
wire _552_;
wire _553_;
wire _554_;
wire _555_;
wire _556_;
wire _557_;
wire _558_;
wire _559_;
wire _560_;
wire _561_;
wire _562_;
wire _563_;
wire _564_;
wire _565_;
wire _566_;
wire _567_;
wire _568_;
wire _569_;
wire _570_;
wire _571_;
wire _572_;
wire _573_;
wire _574_;
wire _575_;
wire _576_;
wire _577_;
wire _578_;
wire _579_;
wire _580_;
wire _581_;
wire _582_;
wire _583_;
wire _584_;
wire _585_;
wire _586_;
wire _587_;
wire _588_;
wire _589_;
wire _590_;
wire _591_;
wire _592_;
wire _593_;
wire _594_;
wire _595_;
wire _596_;
wire _597_;
wire _598_;
wire _599_;
wire _600_;
wire _601_;
wire _602_;
wire _603_;
wire _604_;
wire _605_;
wire _606_;
wire _607_;
wire _608_;
wire _609_;
wire _610_;
wire _611_;
wire _612_;
wire _613_;
wire _614_;
wire _615_;
wire _616_;
wire _617_;
wire _618_;
wire _619_;
wire _620_;
wire _621_;
wire _622_;
wire _623_;
wire _624_;
wire _625_;
wire _626_;
wire _627_;
wire _628_;
wire _629_;
wire _630_;
wire _631_;
wire _632_;
wire _633_;
wire _634_;
wire _635_;
wire _636_;
wire _637_;
wire _638_;
wire _639_;
wire _640_;
wire _641_;
wire _642_;
wire _643_;
wire _644_;
wire _645_;
wire _646_;
wire _647_;
wire _648_;
wire _649_;
wire _650_;
wire _651_;
wire _652_;
wire _653_;
wire _654_;
wire _655_;
wire _656_;
wire _657_;
wire _658_;
wire _659_;
wire _660_;
wire _661_;
wire _662_;
wire _663_;
wire _664_;
wire _665_;
wire _666_;
wire _667_;
wire _668_;
wire _669_;
wire _670_;
wire _671_;
wire _672_;
wire _673_;
wire _674_;
wire _675_;
wire _676_;
wire _677_;
wire _678_;
wire _679_;
wire _680_;
wire _681_;
wire _682_;
wire _683_;
wire _684_;
wire _685_;
wire _686_;
wire _687_;
wire _688_;
wire _689_;
wire _690_;
wire _691_;
wire _692_;
wire _693_;
wire _694_;
wire _695_;
wire _696_;
wire _697_;
wire _698_;
wire _699_;
wire _700_;
wire _701_;
wire _702_;
wire _703_;
wire _704_;
wire _705_;
wire _706_;
wire _707_;
wire _708_;
wire _709_;
wire _710_;
wire _711_;
wire _712_;
wire _713_;
wire _714_;
wire _715_;
wire _716_;
wire _717_;
wire _718_;
wire _719_;
wire _720_;
wire _721_;
wire _722_;
wire _723_;
wire _724_;
wire _725_;
wire _726_;
wire _727_;
wire _728_;
wire _729_;
wire _730_;
wire _731_;
wire _732_;
wire _733_;
wire _734_;
wire _735_;
wire _736_;
wire _737_;
wire _738_;
wire _739_;
wire _740_;
wire _741_;
wire _742_;
wire _743_;
wire _744_;
wire _745_;
wire _746_;
wire _747_;
wire _748_;
wire _749_;
wire _750_;
wire _751_;
wire _752_;
wire _753_;
wire _754_;
wire _755_;
wire _756_;
wire _757_;
wire _758_;
wire _759_;
wire _760_;
wire _761_;
wire _762_;
wire _763_;
wire _764_;
wire _765_;
wire _766_;
wire _767_;
wire _768_;
wire _769_;
wire _770_;
wire _771_;
wire _772_;
wire _773_;
wire _774_;
wire _775_;
wire _776_;
wire _777_;
wire _778_;
wire _779_;
wire _780_;
wire _781_;
wire _782_;
wire _783_;
wire _784_;
wire _785_;
wire _786_;
wire _787_;
wire _788_;
wire _789_;
wire _790_;
wire _791_;
wire _792_;
wire _793_;
wire _794_;
wire _795_;
wire _796_;
wire _797_;
wire _798_;
wire _799_;
wire _800_;
wire _801_;
wire _802_;
wire _803_;
wire _804_;
wire _805_;
wire _806_;
wire _807_;
wire _808_;
wire _809_;
wire _810_;
wire _811_;
wire _812_;
wire _813_;
wire _814_;
wire _815_;
wire _816_;
wire _817_;
wire _818_;
wire _819_;
wire _820_;
wire _821_;
wire _822_;
wire _823_;
wire _824_;
wire _825_;
wire _826_;
wire _827_;
wire _828_;
wire _829_;
wire _830_;
wire _831_;
wire _832_;
wire _833_;
wire _834_;
wire _835_;
wire _836_;
wire _837_;
wire _838_;
wire _839_;
wire _840_;
wire _841_;
wire _842_;
wire _843_;
wire _844_;
wire _845_;
wire _846_;
wire _847_;
wire _848_;
wire _849_;
wire _850_;
wire _851_;
wire _852_;
wire _853_;
wire _854_;
wire _855_;
wire _856_;
wire _857_;
wire _858_;
wire _859_;
wire _860_;
wire _861_;
wire _862_;
wire _863_;
wire _864_;
wire _865_;
wire _866_;
wire _867_;
wire _868_;
wire _869_;
wire _870_;
wire _871_;
wire _872_;
wire _873_;
wire _874_;
wire _875_;
wire _876_;
wire _877_;
wire _878_;
wire _879_;
wire _880_;
wire _881_;
wire _882_;
wire _883_;
wire _884_;
wire _885_;
wire _886_;
wire _887_;
wire _888_;
wire _889_;
wire _890_;
wire _891_;
wire _892_;
wire _893_;
wire _894_;
wire _895_;
wire _896_;
wire _897_;
wire _898_;
wire _899_;
wire _900_;
wire _901_;
wire _902_;
wire _903_;
wire _904_;
wire _905_;
wire _906_;
wire _907_;
wire _908_;
wire _909_;
wire _910_;
wire _911_;
wire _912_;
wire _913_;
wire _914_;
wire _915_;
wire _916_;
wire _917_;
wire _918_;
wire _919_;
wire _920_;
wire _921_;
wire _922_;
wire _923_;
wire _924_;
wire _925_;
wire _926_;
wire _927_;
wire _928_;
wire _929_;
wire _930_;
wire _931_;
wire _932_;
wire _933_;
wire _934_;
wire _935_;
wire _936_;
wire _937_;
wire _938_;
wire _939_;
wire _940_;
wire _941_;
wire _942_;
wire _943_;
wire _944_;
wire _945_;
wire _946_;
wire _947_;
wire _948_;
wire _949_;
wire _950_;
wire _951_;
wire _952_;
wire _953_;
wire _954_;
wire _955_;
wire _956_;
wire _957_;
wire _958_;
wire _959_;
wire _960_;
wire _961_;
wire _962_;
wire _963_;
wire _964_;
wire _965_;
wire _966_;
wire _967_;
wire _968_;
wire _969_;
wire _970_;
wire _971_;
wire _972_;
wire _973_;
wire _974_;
wire _975_;
wire _976_;
wire _977_;
wire _978_;
wire _979_;
wire _980_;
wire _981_;
wire _982_;
wire _983_;
wire _984_;
wire _985_;
wire _986_;
wire _987_;
wire _988_;
wire _989_;
wire _990_;
wire _991_;
wire _992_;
wire _993_;
wire _994_;
wire _995_;
wire _996_;
wire _997_;
wire _998_;
wire _999_;
wire _1000_;
wire _1001_;
wire _1002_;
wire _1003_;
wire _1004_;
wire _1005_;
wire _1006_;
wire _1007_;
wire _1008_;
wire _1009_;
wire _1010_;
wire _1011_;
wire _1012_;
wire _1013_;
wire _1014_;
wire _1015_;
wire _1016_;
wire _1017_;
wire _1018_;
wire _1019_;
wire _1020_;
wire _1021_;
wire _1022_;
wire _1023_;
wire _1024_;
wire _1025_;
wire _1026_;
wire _1027_;
wire _1028_;
wire _1029_;
wire _1030_;
wire _1031_;
wire _1032_;
wire _1033_;
wire _1034_;
wire _1035_;
wire _1036_;
wire _1037_;
wire _1038_;
wire _1039_;
wire _1040_;
wire _1041_;
wire _1042_;
wire _1043_;
wire _1044_;
wire _1045_;
wire _1046_;
wire _1047_;
wire _1048_;
wire _1049_;
wire _1050_;
wire _1051_;
wire _1052_;
wire _1053_;
wire _1054_;
wire _1055_;
wire _1056_;
wire _1057_;
wire _1058_;
wire _1059_;
wire _1060_;
wire _1061_;
wire _1062_;
wire _1063_;
wire _1064_;
wire _1065_;
wire _1066_;
wire _1067_;
wire _1068_;
wire _1069_;
wire _1070_;
wire _1071_;
wire _1072_;
wire _1073_;
wire _1074_;
wire _1075_;
wire _1076_;
wire _1077_;
wire _1078_;
wire _1079_;
wire _1080_;
wire _1081_;
wire _1082_;
wire _1083_;
wire _1084_;
wire _1085_;
wire _1086_;
wire _1087_;
wire _1088_;
wire _1089_;
wire _1090_;
wire _1091_;
wire _1092_;
wire _1093_;
wire _1094_;
wire _1095_;
wire _1096_;
wire _1097_;
wire _1098_;
wire _1099_;
wire _1100_;
wire _1101_;
wire _1102_;
wire _1103_;
wire _1104_;
wire _1105_;
wire _1106_;
wire _1107_;
wire _1108_;
wire _1109_;
wire _1110_;
wire _1111_;
wire _1112_;
wire _1113_;
wire _1114_;
wire _1115_;
wire _1116_;
wire _1117_;
wire _1118_;
wire _1119_;
wire _1120_;
wire _1121_;
wire _1122_;
wire _1123_;
wire _1124_;
wire _1125_;
wire _1126_;
wire _1127_;
wire _1128_;
wire _1129_;
wire _1130_;
wire _1131_;
wire _1132_;
wire _1133_;
wire _1134_;
wire _1135_;
wire _1136_;
wire _1137_;
wire _1138_;
wire _1139_;
wire _1140_;
wire _1141_;
wire _1142_;
wire _1143_;
wire _1144_;
wire _1145_;
wire _1146_;
wire _1147_;
wire _1148_;
wire _1149_;
wire _1150_;
wire _1151_;
wire _1152_;
wire _1153_;
wire _1154_;
wire _1155_;
wire _1156_;
wire _1157_;
wire _1158_;
wire _1159_;
wire _1160_;
wire _1161_;
wire _1162_;
wire _1163_;
wire _1164_;
wire _1165_;
wire _1166_;
wire _1167_;
wire _1168_;
wire _1169_;
wire _1170_;
wire _1171_;
wire _1172_;
wire _1173_;
wire _1174_;
wire _1175_;
wire _1176_;
wire _1177_;
wire _1178_;
wire _1179_;
wire _1180_;
wire _1181_;
wire _1182_;
wire _1183_;
wire _1184_;
wire _1185_;
wire _1186_;
wire _1187_;
wire _1188_;
wire _1189_;
wire _1190_;
wire _1191_;
wire _1192_;
wire _1193_;
wire _1194_;
wire _1195_;
wire _1196_;
wire _1197_;
wire _1198_;
wire _1199_;
wire _1200_;
wire _1201_;
wire _1202_;
wire _1203_;
wire _1204_;
wire _1205_;
wire _1206_;
wire _1207_;
wire _1208_;
wire _1209_;
wire _1210_;
wire _1211_;
wire _1212_;
wire _1213_;
wire _1214_;
wire _1215_;
wire _1216_;
wire _1217_;
wire _1218_;
wire _1219_;
wire _1220_;
wire _1221_;
wire _1222_;
wire _1223_;
wire _1224_;
wire _1225_;
wire _1226_;
wire _1227_;
wire _1228_;
wire _1229_;
wire _1230_;
wire _1231_;
wire _1232_;
wire _1233_;
wire _1234_;
wire _1235_;
wire _1236_;
wire _1237_;
wire _1238_;
wire _1239_;
wire _1240_;
wire _1241_;
wire _1242_;
wire _1243_;
wire _1244_;
wire _1245_;
wire _1246_;
wire _1247_;
wire _1248_;
wire _1249_;
wire _1250_;
wire _1251_;
wire _1252_;
wire _1253_;
wire _1254_;
wire _1255_;
wire _1256_;
wire _1257_;
wire _1258_;
wire _1259_;
wire _1260_;
wire _1261_;
wire _1262_;
wire _1263_;
wire _1264_;
wire _1265_;
wire _1266_;
wire _1267_;
wire _1268_;
wire _1269_;
wire _1270_;
wire _1271_;
wire _1272_;
wire _1273_;
wire _1274_;
wire _1275_;
wire _1276_;
wire _1277_;
wire _1278_;
wire _1279_;
wire _1280_;
wire _1281_;
wire _1282_;
wire _1283_;
wire _1284_;
wire _1285_;
wire _1286_;
wire _1287_;
wire _1288_;
wire _1289_;
wire _1290_;
wire _1291_;
wire _1292_;
wire _1293_;
wire _1294_;
wire _1295_;
wire _1296_;
wire _1297_;
wire _1298_;
wire _1299_;
wire _1300_;
wire _1301_;
wire _1302_;
wire _1303_;
wire _1304_;
wire _1305_;
wire _1306_;
wire _1307_;
wire _1308_;
wire _1309_;
wire _1310_;
wire _1311_;
wire _1312_;
wire _1313_;
wire _1314_;
wire _1315_;
wire _1316_;
wire _1317_;
wire _1318_;
wire _1319_;
wire _1320_;
wire _1321_;
wire _1322_;
wire _1323_;
wire _1324_;
wire _1325_;
wire _1326_;
wire _1327_;
wire _1328_;
wire _1329_;
wire _1330_;
wire _1331_;
wire _1332_;
wire _1333_;
wire _1334_;
wire _1335_;
wire _1336_;
wire _1337_;
wire _1338_;
wire _1339_;
wire _1340_;
wire _1341_;
wire _1342_;
wire _1343_;
wire _1344_;
wire _1345_;
wire _1346_;
wire _1347_;
wire _1348_;
wire _1349_;
wire _1350_;
wire _1351_;
wire _1352_;
wire _1353_;
wire _1354_;
wire _1355_;
wire _1356_;
wire _1357_;
wire _1358_;
wire _1359_;
wire _1360_;
wire _1361_;
wire _1362_;
wire _1363_;
wire _1364_;
wire _1365_;
wire _1366_;
wire _1367_;
wire _1368_;
wire _1369_;
wire _1370_;
wire _1371_;
wire _1372_;
wire _1373_;
wire _1374_;
wire _1375_;
wire _1376_;
wire _1377_;
wire _1378_;
wire _1379_;
wire _1380_;
wire _1381_;
wire _1382_;
wire _1383_;
wire _1384_;
wire _1385_;
wire _1386_;
wire _1387_;
wire _1388_;
wire _1389_;
wire _1390_;
wire _1391_;
wire _1392_;
wire _1393_;
wire _1394_;
wire _1395_;
wire _1396_;
wire _1397_;
wire _1398_;
wire _1399_;
wire _1400_;
wire _1401_;
wire _1402_;
wire _1403_;
wire _1404_;
wire _1405_;
wire _1406_;
wire _1407_;
wire _1408_;
wire _1409_;
wire _1410_;
wire _1411_;
wire _1412_;
wire _1413_;
wire _1414_;
wire _1415_;
wire _1416_;
wire _1417_;
wire _1418_;
wire _1419_;
wire _1420_;
wire _1421_;
wire _1422_;
wire _1423_;
wire _1424_;
wire _1425_;
wire _1426_;
wire _1427_;
wire _1428_;
wire _1429_;
wire _1430_;
wire _1431_;
wire _1432_;
wire _1433_;
wire _1434_;
wire _1435_;
wire _1436_;
wire _1437_;
wire _1438_;
wire _1439_;
wire _1440_;
wire _1441_;
wire _1442_;
wire _1443_;
wire _1444_;
wire _1445_;
wire _1446_;
wire _1447_;
wire _1448_;
wire _1449_;
wire _1450_;
wire _1451_;
wire _1452_;
wire _1453_;
wire _1454_;
wire _1455_;
wire _1456_;
wire _1457_;
wire _1458_;
wire _1459_;
wire _1460_;
wire _1461_;
wire _1462_;
wire _1463_;
wire _1464_;
wire _1465_;
wire _1466_;
wire _1467_;
wire _1468_;
wire _1469_;
wire _1470_;
wire _1471_;
wire _1472_;
wire _1473_;
wire _1474_;
wire _1475_;
wire _1476_;
wire _1477_;
wire _1478_;
wire _1479_;
wire _1480_;
wire _1481_;
wire _1482_;
wire _1483_;
wire _1484_;
wire _1485_;
wire _1486_;
wire _1487_;
wire _1488_;
wire _1489_;
wire _1490_;
wire _1491_;
wire _1492_;
wire _1493_;
wire _1494_;
wire _1495_;
wire _1496_;
wire _1497_;
wire _1498_;
wire _1499_;
wire _1500_;
wire _1501_;
wire _1502_;
wire _1503_;
wire _1504_;
wire _1505_;
wire _1506_;
wire _1507_;
wire _1508_;
wire _1509_;
wire _1510_;
wire _1511_;
wire _1512_;
wire _1513_;
wire _1514_;
wire _1515_;
wire _1516_;
wire _1517_;
wire _1518_;
wire _1519_;
wire _1520_;
wire _1521_;
wire _1522_;
wire _1523_;
wire _1524_;
wire _1525_;
wire _1526_;
wire _1527_;
wire _1528_;
wire _1529_;
wire _1530_;
wire _1531_;
wire _1532_;
wire _1533_;
wire _1534_;
wire _1535_;
wire _1536_;
wire _1537_;
wire _1538_;
wire _1539_;
wire _1540_;
wire _1541_;
wire _1542_;
wire _1543_;
wire _1544_;
wire _1545_;
wire _1546_;
wire _1547_;
wire _1548_;
wire _1549_;
wire _1550_;
wire _1551_;
wire _1552_;
wire _1553_;
wire _1554_;
wire _1555_;
wire _1556_;
wire _1557_;
wire _1558_;
wire _1559_;
wire _1560_;
wire _1561_;
wire _1562_;
wire _1563_;
wire _1564_;
wire _1565_;
wire _1566_;
wire _1567_;
wire _1568_;
wire _1569_;
wire _1570_;
wire _1571_;
wire _1572_;
wire _1573_;
wire _1574_;
wire _1575_;
wire _1576_;
wire _1577_;
wire _1578_;
wire _1579_;
wire _1580_;
wire _1581_;
wire _1582_;
wire _1583_;
wire _1584_;
wire _1585_;
wire _1586_;
wire _1587_;
wire _1588_;
wire _1589_;
wire _1590_;
wire _1591_;
wire _1592_;
wire _1593_;
wire _1594_;
wire _1595_;
wire _1596_;
wire _1597_;
wire _1598_;
wire _1599_;
wire _1600_;
wire _1601_;
wire _1602_;
wire _1603_;
wire _1604_;
wire _1605_;
wire _1606_;
wire _1607_;
wire _1608_;
wire _1609_;
wire _1610_;
wire _1611_;
wire _1612_;
wire _1613_;
wire _1614_;
wire _1615_;
wire _1616_;
wire _1617_;
wire _1618_;
wire _1619_;
wire _1620_;
wire _1621_;
wire _1622_;
wire _1623_;
wire _1624_;
wire _1625_;
wire _1626_;
wire _1627_;
wire _1628_;
wire _1629_;
wire _1630_;
wire _1631_;
wire _1632_;
wire _1633_;
wire _1634_;
wire _1635_;
wire _1636_;
wire _1637_;
wire _1638_;
wire _1639_;
wire _1640_;
wire _1641_;
wire _1642_;
wire _1643_;
wire _1644_;
wire _1645_;
wire _1646_;
wire _1647_;
wire _1648_;
wire _1649_;
wire _1650_;
wire _1651_;
wire _1652_;
wire _1653_;
wire _1654_;
wire _1655_;
wire _1656_;
wire _1657_;
wire _1658_;
wire _1659_;
wire _1660_;
wire _1661_;
wire _1662_;
wire _1663_;
wire _1664_;
wire _1665_;
wire _1666_;
wire _1667_;
wire _1668_;
wire _1669_;
wire _1670_;
wire _1671_;
wire _1672_;
wire _1673_;
wire _1674_;
wire _1675_;
wire _1676_;
wire _1677_;
wire _1678_;
wire _1679_;
wire _1680_;
wire _1681_;
wire _1682_;
wire _1683_;
wire _1684_;
wire _1685_;
wire _1686_;
wire _1687_;
wire _1688_;
wire _1689_;
wire _1690_;
wire _1691_;
wire _1692_;
wire _1693_;
wire _1694_;
wire _1695_;
wire _1696_;
wire _1697_;
wire _1698_;
wire _1699_;
wire _1700_;
wire _1701_;
wire _1702_;
wire _1703_;
wire _1704_;
wire _1705_;
wire _1706_;
wire _1707_;
wire _1708_;
wire _1709_;
wire _1710_;
wire _1711_;
wire _1712_;
wire _1713_;
wire _1714_;
wire _1715_;
wire _1716_;
wire _1717_;
wire _1718_;
wire _1719_;
wire _1720_;
wire _1721_;
wire _1722_;
wire _1723_;
wire _1724_;
wire _1725_;
wire _1726_;
wire _1727_;
wire _1728_;
wire _1729_;
wire _1730_;
wire _1731_;
wire _1732_;
wire _1733_;
wire _1734_;
wire _1735_;
wire _1736_;
wire _1737_;
wire _1738_;
wire _1739_;
wire _1740_;
wire _1741_;
wire _1742_;
wire _1743_;
wire _1744_;
wire _1745_;
wire _1746_;
wire _1747_;
wire _1748_;
wire _1749_;
wire _1750_;
wire _1751_;
wire _1752_;
wire _1753_;
wire _1754_;
wire _1755_;
wire _1756_;
wire _1757_;
wire _1758_;
wire _1759_;
wire _1760_;
wire _1761_;
wire _1762_;
wire _1763_;
wire _1764_;
wire _1765_;
wire _1766_;
wire _1767_;
wire _1768_;
wire _1769_;
wire _1770_;
wire _1771_;
wire _1772_;
wire _1773_;
wire _1774_;
wire _1775_;
wire _1776_;
wire _1777_;
wire _1778_;
wire _1779_;
wire _1780_;
wire _1781_;
wire _1782_;
wire _1783_;
wire _1784_;
wire _1785_;
wire _1786_;
wire _1787_;
wire _1788_;
wire _1789_;
wire _1790_;
wire _1791_;
wire _1792_;
wire _1793_;
wire _1794_;
wire _1795_;
wire _1796_;
wire _1797_;
wire _1798_;
wire _1799_;
wire _1800_;
wire _1801_;
wire _1802_;
wire _1803_;
wire _1804_;
wire _1805_;
wire _1806_;
wire _1807_;
wire _1808_;
wire _1809_;
wire _1810_;
wire _1811_;
wire _1812_;
wire _1813_;
wire _1814_;
wire _1815_;
wire _1816_;
wire _1817_;
wire _1818_;
wire _1819_;
wire _1820_;
wire _1821_;
wire _1822_;
wire _1823_;
wire _1824_;
wire _1825_;
wire _1826_;
wire _1827_;
wire _1828_;
wire _1829_;
wire _1830_;
wire _1831_;
wire _1832_;
wire _1833_;
wire _1834_;
wire _1835_;
wire _1836_;
wire _1837_;
wire _1838_;
wire _1839_;
wire _1840_;
wire _1841_;
wire _1842_;
wire _1843_;
wire _1844_;
wire _1845_;
wire _1846_;
wire _1847_;
wire _1848_;
wire _1849_;
wire _1850_;
wire _1851_;
wire _1852_;
wire _1853_;
wire _1854_;
wire _1855_;
wire _1856_;
wire _1857_;
wire _1858_;
wire _1859_;
wire _1860_;
wire _1861_;
wire _1862_;
wire _1863_;
wire _1864_;
wire _1865_;
wire _1866_;
wire _1867_;
wire _1868_;
wire _1869_;
wire _1870_;
wire _1871_;
wire _1872_;
wire _1873_;
wire _1874_;
wire _1875_;
wire _1876_;
wire _1877_;
wire _1878_;
wire _1879_;
wire _1880_;
wire _1881_;
wire _1882_;
wire _1883_;
wire _1884_;
wire _1885_;
wire _1886_;
wire _1887_;
wire _1888_;
wire _1889_;
wire _1890_;
wire _1891_;
wire _1892_;
wire _1893_;
wire _1894_;
wire _1895_;
wire _1896_;
wire _1897_;
wire _1898_;
wire _1899_;
wire _1900_;
wire _1901_;
wire _1902_;
wire _1903_;
wire _1904_;
wire _1905_;
wire _1906_;
wire _1907_;
wire _1908_;
wire _1909_;
wire _1910_;
wire _1911_;
wire _1912_;
wire _1913_;
wire _1914_;
wire _1915_;
wire _1916_;
wire _1917_;
wire _1918_;
wire _1919_;
wire _1920_;
wire _1921_;
wire _1922_;
wire _1923_;
wire _1924_;
wire _1925_;
wire _1926_;
wire _1927_;
wire _1928_;
wire _1929_;
wire _1930_;
wire _1931_;
wire _1932_;
wire _1933_;
wire _1934_;
wire _1935_;
wire _1936_;
wire _1937_;
wire _1938_;
wire _1939_;
wire _1940_;
wire _1941_;
wire _1942_;
wire _1943_;
wire _1944_;
wire _1945_;
wire _1946_;
wire _1947_;
wire _1948_;
wire _1949_;
wire _1950_;
wire _1951_;
wire _1952_;
wire _1953_;
wire _1954_;
wire _1955_;
wire _1956_;
wire _1957_;
wire _1958_;
wire _1959_;
wire _1960_;
wire _1961_;
wire _1962_;
wire _1963_;
wire _1964_;
wire _1965_;
wire _1966_;
wire _1967_;
wire _1968_;
wire _1969_;
wire _1970_;
wire _1971_;
wire _1972_;
wire _1973_;
wire _1974_;
wire _1975_;
wire _1976_;
wire _1977_;
wire _1978_;
wire _1979_;
wire _1980_;
wire _1981_;
wire _1982_;
wire _1983_;
wire _1984_;
wire _1985_;
wire _1986_;
wire _1987_;
wire _1988_;
wire _1989_;
wire _1990_;
wire _1991_;
wire _1992_;
wire _1993_;
wire _1994_;
wire _1995_;
wire _1996_;
wire _1997_;
wire _1998_;
wire _1999_;
wire _2000_;
wire _2001_;
wire _2002_;
wire _2003_;
wire _2004_;
wire _2005_;
wire _2006_;
wire _2007_;
wire _2008_;
wire _2009_;
wire _2010_;
wire _2011_;
wire _2012_;
wire _2013_;
wire _2014_;
wire _2015_;
wire _2016_;
wire _2017_;
wire _2018_;
wire _2019_;
wire _2020_;
wire _2021_;
wire _2022_;
wire _2023_;
wire _2024_;
wire _2025_;
wire _2026_;
wire _2027_;
wire _2028_;
wire _2029_;
wire _2030_;
wire _2031_;
wire _2032_;
wire _2033_;
wire _2034_;
wire _2035_;
wire _2036_;
wire _2037_;
wire _2038_;
wire _2039_;
wire _2040_;
wire _2041_;
wire _2042_;
wire _2043_;
wire _2044_;
wire _2045_;
wire _2046_;
wire _2047_;
wire _2048_;
wire _2049_;
wire _2050_;
wire _2051_;
wire _2052_;
wire _2053_;
wire _2054_;
wire _2055_;
wire _2056_;
wire _2057_;
wire _2058_;
wire _2059_;
wire _2060_;
wire _2061_;
wire _2062_;
wire _2063_;
wire _2064_;
wire _2065_;
wire _2066_;
wire _2067_;
wire _2068_;
wire _2069_;
wire _2070_;
wire _2071_;
wire _2072_;
wire _2073_;
wire _2074_;
wire _2075_;
wire _2076_;
wire _2077_;
wire _2078_;
wire _2079_;
wire _2080_;
wire _2081_;
wire _2082_;
wire _2083_;
wire _2084_;
wire _2085_;
wire _2086_;
wire _2087_;
wire _2088_;
wire _2089_;
wire _2090_;
wire _2091_;
wire _2092_;
wire _2093_;
wire _2094_;
wire _2095_;
wire _2096_;
wire _2097_;
wire _2098_;
wire _2099_;
wire _2100_;
wire _2101_;
wire _2102_;
wire _2103_;
wire _2104_;
wire _2105_;
wire _2106_;
wire _2107_;
wire _2108_;
wire _2109_;
wire _2110_;
wire _2111_;
wire _2112_;
wire _2113_;
wire _2114_;
wire _2115_;
wire _2116_;
wire _2117_;
wire _2118_;
wire _2119_;
wire _2120_;
wire _2121_;
wire _2122_;
wire _2123_;
wire _2124_;
wire _2125_;
wire _2126_;
wire _2127_;
wire _2128_;
wire _2129_;
wire _2130_;
wire _2131_;
wire _2132_;
wire _2133_;
wire _2134_;
wire _2135_;
wire _2136_;
wire _2137_;
wire _2138_;
wire _2139_;
wire _2140_;
wire _2141_;
wire _2142_;
wire _2143_;
wire _2144_;
wire _2145_;
wire _2146_;
wire _2147_;
wire _2148_;
wire _2149_;
wire _2150_;
wire _2151_;
wire _2152_;
wire _2153_;
wire _2154_;
wire _2155_;
wire _2156_;
wire _2157_;
wire _2158_;
wire _2159_;
wire _2160_;
wire _2161_;
wire _2162_;
wire _2163_;
wire _2164_;
wire _2165_;
wire _2166_;
wire _2167_;
wire _2168_;
wire _2169_;
wire _2170_;
wire _2171_;
wire _2172_;
wire _2173_;
wire _2174_;
wire _2175_;
wire _2176_;
wire _2177_;
wire _2178_;
wire _2179_;
wire _2180_;
wire _2181_;
wire _2182_;
wire _2183_;
wire _2184_;
wire _2185_;
wire _2186_;
wire _2187_;
wire _2188_;
wire _2189_;
wire _2190_;
wire _2191_;
wire _2192_;
wire _2193_;
wire _2194_;
wire _2195_;
wire _2196_;
wire _2197_;
wire _2198_;
wire _2199_;
wire _2200_;
wire _2201_;
wire _2202_;
wire _2203_;
wire _2204_;
wire _2205_;
wire _2206_;
wire _2207_;
wire _2208_;
wire _2209_;
wire _2210_;
wire _2211_;
wire _2212_;
wire _2213_;
wire _2214_;
wire _2215_;
wire _2216_;
wire _2217_;
wire _2218_;
wire _2219_;
wire _2220_;
wire _2221_;
wire _2222_;
wire _2223_;
wire _2224_;
wire _2225_;
wire _2226_;
wire _2227_;
wire _2228_;
wire _2229_;
wire _2230_;
wire _2231_;
wire _2232_;
wire _2233_;
wire _2234_;
wire _2235_;
wire _2236_;
wire _2237_;
wire _2238_;
wire _2239_;
wire _2240_;
wire _2241_;
wire _2242_;
wire _2243_;
wire _2244_;
wire _2245_;
wire _2246_;
wire _2247_;
wire _2248_;
wire _2249_;
wire _2250_;
wire _2251_;
wire _2252_;
wire _2253_;
wire _2254_;
wire _2255_;
wire _2256_;
wire _2257_;
wire _2258_;
wire _2259_;
wire _2260_;
wire _2261_;
wire _2262_;
wire _2263_;
wire _2264_;
wire _2265_;
wire _2266_;
wire _2267_;
wire _2268_;
wire _2269_;
wire _2270_;
wire _2271_;
wire _2272_;
wire _2273_;
wire _2274_;
wire _2275_;
wire _2276_;
wire _2277_;
wire _2278_;
wire _2279_;
wire _2280_;
wire _2281_;
wire _2282_;
wire _2283_;
wire _2284_;
wire _2285_;
wire _2286_;
wire _2287_;
wire _2288_;
wire _2289_;
wire _2290_;
wire _2291_;
wire _2292_;
wire _2293_;
wire _2294_;
wire _2295_;
wire _2296_;
wire _2297_;
wire _2298_;
wire _2299_;
wire _2300_;
wire _2301_;
wire _2302_;
wire _2303_;
wire _2304_;
wire _2305_;
wire _2306_;
wire _2307_;
wire _2308_;
wire _2309_;
wire _2310_;
wire _2311_;
wire _2312_;
wire _2313_;
wire _2314_;
wire _2315_;
wire _2316_;
wire _2317_;
wire _2318_;
wire _2319_;
wire _2320_;
wire _2321_;
wire _2322_;
wire _2323_;
wire _2324_;
wire _2325_;
wire _2326_;
wire _2327_;
wire _2328_;
wire _2329_;
wire _2330_;
wire _2331_;
wire _2332_;
wire _2333_;
wire _2334_;
wire _2335_;
wire _2336_;
wire _2337_;
wire _2338_;
wire _2339_;
wire _2340_;
wire _2341_;
wire _2342_;
wire _2343_;
wire _2344_;
wire _2345_;
wire _2346_;
wire _2347_;
wire _2348_;
wire _2349_;
wire _2350_;
wire _2351_;
wire _2352_;
wire _2353_;
wire _2354_;
wire _2355_;
wire _2356_;
wire _2357_;
wire _2358_;
wire _2359_;
wire _2360_;
wire _2361_;
wire _2362_;
wire _2363_;
wire _2364_;
wire _2365_;
wire _2366_;
wire _2367_;
wire _2368_;
wire _2369_;
wire _2370_;
wire _2371_;
wire _2372_;
wire _2373_;
wire _2374_;
wire _2375_;
wire _2376_;
wire _2377_;
wire _2378_;
wire _2379_;
wire _2380_;
wire _2381_;
wire _2382_;
wire _2383_;
wire _2384_;
wire _2385_;
wire _2386_;
wire _2387_;
wire _2388_;
wire _2389_;
wire _2390_;
wire _2391_;
wire _2392_;
wire _2393_;
wire _2394_;
wire _2395_;
wire _2396_;
wire _2397_;
wire _2398_;
wire _2399_;
wire _2400_;
wire _2401_;
wire _2402_;
wire _2403_;
wire _2404_;
wire _2405_;
wire _2406_;
wire _2407_;
wire _2408_;
wire _2409_;
wire _2410_;
wire _2411_;
wire _2412_;
wire _2413_;
wire _2414_;
wire _2415_;
wire _2416_;
wire _2417_;
wire _2418_;
wire _2419_;
wire _2420_;
wire _2421_;
wire _2422_;
wire _2423_;
wire _2424_;
wire _2425_;
wire _2426_;
wire _2427_;
wire _2428_;
wire _2429_;
wire _2430_;
wire _2431_;
wire _2432_;
wire _2433_;
wire _2434_;
wire _2435_;
wire _2436_;
wire _2437_;
wire _2438_;
wire _2439_;
wire _2440_;
wire _2441_;
wire _2442_;
wire _2443_;
wire _2444_;
wire _2445_;
wire _2446_;
wire _2447_;
wire _2448_;
wire _2449_;
wire _2450_;
wire _2451_;
wire _2452_;
wire _2453_;
wire _2454_;
wire _2455_;
wire _2456_;
wire _2457_;
wire _2458_;
wire _2459_;
wire _2460_;
wire _2461_;
wire _2462_;
wire _2463_;
wire _2464_;
wire _2465_;
wire _2466_;
wire _2467_;
wire _2468_;
wire _2469_;
wire _2470_;
wire _2471_;
wire _2472_;
wire _2473_;
wire _2474_;
wire _2475_;
wire _2476_;
wire _2477_;
wire _2478_;
wire _2479_;
wire _2480_;
wire _2481_;
wire _2482_;
wire _2483_;
wire _2484_;
wire _2485_;
wire _2486_;
wire _2487_;
wire _2488_;
wire _2489_;
wire _2490_;
wire _2491_;
wire _2492_;
wire _2493_;
wire _2494_;
wire _2495_;
wire _2496_;
wire _2497_;
wire _2498_;
wire _2499_;
wire _2500_;
wire _2501_;
wire _2502_;
wire _2503_;
wire _2504_;
wire _2505_;
wire _2506_;
wire _2507_;
wire _2508_;
wire _2509_;
wire _2510_;
wire _2511_;
wire _2512_;
wire _2513_;
wire _2514_;
wire _2515_;
wire _2516_;
wire _2517_;
wire _2518_;
wire _2519_;
wire _2520_;
wire _2521_;
wire _2522_;
wire _2523_;
wire _2524_;
wire _2525_;
wire _2526_;
wire _2527_;
wire _2528_;
wire _2529_;
wire _2530_;
wire _2531_;
wire _2532_;
wire _2533_;
wire _2534_;
wire _2535_;
wire _2536_;
wire _2537_;
wire _2538_;
wire _2539_;
wire _2540_;
wire _2541_;
wire _2542_;
wire _2543_;
wire _2544_;
wire _2545_;
wire _2546_;
wire _2547_;
wire _2548_;
wire _2549_;
wire _2550_;
wire _2551_;
wire _2552_;
wire _2553_;
wire _2554_;
wire _2555_;
wire _2556_;
wire _2557_;
wire _2558_;
wire _2559_;
wire _2560_;
wire _2561_;
wire _2562_;
wire _2563_;
wire _2564_;
wire _2565_;
wire _2566_;
wire _2567_;
wire _2568_;
wire _2569_;
wire _2570_;
wire _2571_;
wire _2572_;
wire _2573_;
wire _2574_;
wire _2575_;
wire _2576_;
wire _2577_;
wire _2578_;
wire _2579_;
wire _2580_;
wire _2581_;
wire _2582_;
wire _2583_;
wire _2584_;
wire _2585_;
wire _2586_;
wire _2587_;
wire _2588_;
wire _2589_;
wire _2590_;
wire _2591_;
wire _2592_;
wire _2593_;
wire _2594_;
wire _2595_;
wire _2596_;
wire _2597_;
wire _2598_;
wire _2599_;
wire _2600_;
wire _2601_;
wire _2602_;
wire _2603_;
wire _2604_;
wire _2605_;
wire _2606_;
wire _2607_;
wire _2608_;
wire _2609_;
wire _2610_;
wire _2611_;
wire _2612_;
wire _2613_;
wire _2614_;
wire _2615_;
wire _2616_;
wire _2617_;
wire _2618_;
wire _2619_;
wire _2620_;
wire _2621_;
wire _2622_;
wire _2623_;
wire _2624_;
wire _2625_;
wire _2626_;
wire _2627_;
wire _2628_;
wire _2629_;
wire _2630_;
wire _2631_;
wire _2632_;
wire _2633_;
wire _2634_;
wire _2635_;
wire _2636_;
wire _2637_;
wire _2638_;
wire _2639_;
wire _2640_;
wire _2641_;
wire _2642_;
wire _2643_;
wire _2644_;
wire _2645_;
wire _2646_;
wire _2647_;
wire _2648_;
wire _2649_;
wire _2650_;
wire _2651_;
wire _2652_;
wire _2653_;
wire _2654_;
wire _2655_;
wire _2656_;
wire _2657_;
wire _2658_;
wire _2659_;
wire _2660_;
wire _2661_;
wire _2662_;
wire _2663_;
wire _2664_;
wire _2665_;
wire _2666_;
wire _2667_;
wire _2668_;
wire _2669_;
wire _2670_;
wire _2671_;
wire _2672_;
wire _2673_;
wire _2674_;
wire _2675_;
wire _2676_;
wire _2677_;
wire _2678_;
wire _2679_;
wire _2680_;
wire _2681_;
wire _2682_;
wire _2683_;
wire _2684_;
wire _2685_;
wire _2686_;
wire _2687_;
wire _2688_;
wire _2689_;
wire _2690_;
wire _2691_;
wire _2692_;
wire _2693_;
wire _2694_;
wire _2695_;
wire _2696_;
wire _2697_;
wire _2698_;
wire _2699_;
wire _2700_;
wire _2701_;
wire _2702_;
wire _2703_;
wire _2704_;
wire _2705_;
wire _2706_;
wire _2707_;
wire _2708_;
wire _2709_;
wire _2710_;
wire _2711_;
wire _2712_;
wire _2713_;
wire _2714_;
wire _2715_;
wire _2716_;
wire _2717_;
wire _2718_;
wire _2719_;
wire _2720_;
wire _2721_;
wire _2722_;
wire _2723_;
wire _2724_;
wire _2725_;
wire _2726_;
wire _2727_;
wire _2728_;
wire _2729_;
wire _2730_;
wire _2731_;
wire _2732_;
wire _2733_;
wire _2734_;
wire _2735_;
wire _2736_;
wire _2737_;
wire _2738_;
wire _2739_;
wire _2740_;
wire _2741_;
wire _2742_;
wire _2743_;
wire _2744_;
wire _2745_;
wire _2746_;
wire _2747_;
wire _2748_;
wire _2749_;
wire _2750_;
wire _2751_;
wire _2752_;
wire _2753_;
wire _2754_;
wire _2755_;
wire _2756_;
wire _2757_;
wire _2758_;
wire _2759_;
wire _2760_;
wire _2761_;
wire _2762_;
wire _2763_;
wire _2764_;
wire _2765_;
wire _2766_;
wire _2767_;
wire _2768_;
wire _2769_;
wire _2770_;
wire _2771_;
wire _2772_;
wire _2773_;
wire _2774_;
wire _2775_;
wire _2776_;
wire _2777_;
wire _2778_;
wire _2779_;
wire _2780_;
wire _2781_;
wire _2782_;
wire _2783_;
wire _2784_;
wire _2785_;
wire _2786_;
wire _2787_;
wire _2788_;
wire _2789_;
wire _2790_;
wire _2791_;
wire _2792_;
wire _2793_;
wire _2794_;
wire _2795_;
wire _2796_;
wire _2797_;
wire _2798_;
wire _2799_;
wire _2800_;
wire _2801_;
wire _2802_;
wire _2803_;
wire _2804_;
wire _2805_;
wire _2806_;
wire _2807_;
wire _2808_;
wire _2809_;
wire _2810_;
wire _2811_;
wire _2812_;
wire _2813_;
wire _2814_;
wire _2815_;
wire _2816_;
wire _2817_;
wire _2818_;
wire _2819_;
wire _2820_;
wire _2821_;
wire _2822_;
wire _2823_;
wire _2824_;
wire _2825_;
wire _2826_;
wire _2827_;
wire _2828_;
wire _2829_;
wire _2830_;
wire _2831_;
wire _2832_;
wire _2833_;
wire _2834_;
wire _2835_;
wire _2836_;
wire _2837_;
wire _2838_;
wire _2839_;
wire _2840_;
wire _2841_;
wire _2842_;
wire _2843_;
wire _2844_;
wire _2845_;
wire _2846_;
wire _2847_;
wire _2848_;
wire _2849_;
wire _2850_;
wire _2851_;
wire _2852_;
wire _2853_;
wire _2854_;
wire _2855_;
wire _2856_;
wire _2857_;
wire _2858_;
wire _2859_;
wire _2860_;
wire _2861_;
wire _2862_;
wire _2863_;
wire _2864_;
wire _2865_;
wire _2866_;
wire _2867_;
wire _2868_;
wire _2869_;
wire _2870_;
wire _2871_;
wire _2872_;
wire _2873_;
wire _2874_;
wire _2875_;
wire _2876_;
wire _2877_;
wire _2878_;
wire _2879_;
wire _2880_;
wire _2881_;
wire _2882_;
wire _2883_;
wire _2884_;
wire _2885_;
wire _2886_;
wire _2887_;
wire _2888_;
wire _2889_;
wire _2890_;
wire _2891_;
wire _2892_;
wire _2893_;
wire _2894_;
wire _2895_;
wire _2896_;
wire _2897_;
wire _2898_;
wire _2899_;
wire _2900_;
wire _2901_;
wire _2902_;
wire _2903_;
wire _2904_;
wire _2905_;
wire _2906_;
wire _2907_;
wire _2908_;
wire _2909_;
wire _2910_;
wire _2911_;
wire _2912_;
wire _2913_;
wire _2914_;
wire _2915_;
wire _2916_;
wire _2917_;
wire _2918_;
wire _2919_;
wire _2920_;
wire _2921_;
wire _2922_;
wire _2923_;
wire _2924_;
wire _2925_;
wire _2926_;
wire _2927_;
wire _2928_;
wire _2929_;
wire _2930_;
wire _2931_;
wire _2932_;
wire _2933_;
wire _2934_;
wire _2935_;
wire _2936_;
wire _2937_;
wire _2938_;
wire _2939_;
wire _2940_;
wire _2941_;
wire _2942_;
wire _2943_;
wire _2944_;
wire _2945_;
wire _2946_;
wire _2947_;
wire _2948_;
wire _2949_;
wire _2950_;
wire _2951_;
wire _2952_;
wire _2953_;
wire _2954_;
wire _2955_;
wire _2956_;
wire _2957_;
wire _2958_;
wire _2959_;
wire _2960_;
wire _2961_;
wire _2962_;
wire _2963_;
wire _2964_;
wire _2965_;
wire _2966_;
wire _2967_;
wire _2968_;
wire _2969_;
wire _2970_;
wire _2971_;
wire _2972_;
wire _2973_;
wire _2974_;
wire _2975_;
wire _2976_;
wire _2977_;
wire _2978_;
wire _2979_;
wire _2980_;
wire _2981_;
wire _2982_;
wire _2983_;
wire _2984_;
wire _2985_;
wire _2986_;
wire _2987_;
wire _2988_;
wire _2989_;
wire _2990_;
wire _2991_;
wire _2992_;
wire _2993_;
wire _2994_;
wire _2995_;
wire _2996_;
wire _2997_;
wire _2998_;
wire _2999_;
wire _3000_;
wire _3001_;
wire _3002_;
wire _3003_;
wire _3004_;
wire _3005_;
wire _3006_;
wire _3007_;
wire _3008_;
wire _3009_;
wire _3010_;
wire _3011_;
wire _3012_;
wire _3013_;
wire _3014_;
wire _3015_;
wire _3016_;
wire _3017_;
wire _3018_;
wire _3019_;
wire _3020_;
wire _3021_;
wire _3022_;
wire _3023_;
wire _3024_;
wire _3025_;
wire _3026_;
wire _3027_;
wire _3028_;
wire _3029_;
wire _3030_;
wire _3031_;
wire _3032_;
wire _3033_;
wire _3034_;
wire _3035_;
wire _3036_;
wire _3037_;
wire _3038_;
wire _3039_;
wire _3040_;
wire _3041_;
wire _3042_;
wire _3043_;
wire _3044_;
wire _3045_;
wire _3046_;
wire _3047_;
wire _3048_;
wire _3049_;
wire _3050_;
wire _3051_;
wire _3052_;
wire _3053_;
wire _3054_;
wire _3055_;
wire _3056_;
wire _3057_;
wire _3058_;
wire _3059_;
wire _3060_;
wire _3061_;
wire _3062_;
wire _3063_;
wire _3064_;
wire _3065_;
wire _3066_;
wire _3067_;
wire _3068_;
wire _3069_;
wire _3070_;
wire _3071_;
wire _3072_;
wire _3073_;
wire _3074_;
wire _3075_;
wire _3076_;
wire _3077_;
wire _3078_;
wire _3079_;
wire _3080_;
wire _3081_;
wire _3082_;
wire _3083_;
wire _3084_;
wire _3085_;
wire _3086_;
wire _3087_;
wire _3088_;
wire _3089_;
wire _3090_;
wire _3091_;
wire _3092_;
wire _3093_;
wire _3094_;
wire _3095_;
wire _3096_;
wire _3097_;
wire _3098_;
wire _3099_;
wire _3100_;
wire _3101_;
wire _3102_;
wire _3103_;
wire _3104_;
wire _3105_;
wire _3106_;
wire _3107_;
wire _3108_;
wire _3109_;
wire _3110_;
wire _3111_;
wire _3112_;
wire _3113_;
wire _3114_;
wire _3115_;
wire _3116_;
wire _3117_;
wire _3118_;
wire _3119_;
wire _3120_;
wire _3121_;
wire _3122_;
wire _3123_;
wire _3124_;
wire _3125_;
wire _3126_;
wire _3127_;
wire _3128_;
wire _3129_;
wire _3130_;
wire _3131_;
wire _3132_;
wire _3133_;
wire _3134_;
wire _3135_;
wire _3136_;
wire _3137_;
wire _3138_;
wire _3139_;
wire _3140_;
wire _3141_;
wire _3142_;
wire _3143_;
wire _3144_;
wire _3145_;
wire _3146_;
wire _3147_;
wire _3148_;
wire _3149_;
wire _3150_;
wire _3151_;
wire _3152_;
wire _3153_;
wire _3154_;
wire _3155_;
wire _3156_;
wire _3157_;
wire _3158_;
wire _3159_;
wire _3160_;
wire _3161_;
wire _3162_;
wire _3163_;
wire _3164_;
wire _3165_;
wire _3166_;
wire _3167_;
wire _3168_;
wire _3169_;
wire _3170_;
wire _3171_;
wire _3172_;
wire _3173_;
wire _3174_;
wire _3175_;
wire _3176_;
wire _3177_;
wire _3178_;
wire _3179_;
wire _3180_;
wire _3181_;
wire _3182_;
wire _3183_;
wire _3184_;
wire _3185_;
wire _3186_;
wire _3187_;
wire _3188_;
wire _3189_;
wire _3190_;
wire _3191_;
wire _3192_;
wire _3193_;
wire _3194_;
wire _3195_;
wire _3196_;
wire _3197_;
wire _3198_;
wire _3199_;
wire _3200_;
wire _3201_;
wire _3202_;
wire _3203_;
wire _3204_;
wire _3205_;
wire _3206_;
wire _3207_;
wire _3208_;
wire _3209_;
wire _3210_;
wire _3211_;
wire _3212_;
wire _3213_;
wire _3214_;
wire _3215_;
wire _3216_;
wire _3217_;
wire _3218_;
wire _3219_;
wire _3220_;
wire _3221_;
wire _3222_;
wire _3223_;
wire _3224_;
wire _3225_;
wire _3226_;
wire _3227_;
wire _3228_;
wire _3229_;
wire _3230_;
wire _3231_;
wire _3232_;
wire _3233_;
wire _3234_;
wire _3235_;
wire _3236_;
wire _3237_;
wire _3238_;
wire _3239_;
wire _3240_;
wire _3241_;
wire _3242_;
wire _3243_;
wire _3244_;
wire _3245_;
wire _3246_;
wire _3247_;
wire _3248_;
wire _3249_;
wire _3250_;
wire _3251_;
wire _3252_;
wire _3253_;
wire _3254_;
wire _3255_;
wire _3256_;
wire _3257_;
wire _3258_;
wire _3259_;
wire _3260_;
wire _3261_;
wire _3262_;
wire _3263_;
wire _3264_;
wire _3265_;
wire _3266_;
wire _3267_;
wire _3268_;
wire _3269_;
wire _3270_;
wire _3271_;
wire _3272_;
wire _3273_;
wire _3274_;
wire _3275_;
wire _3276_;
wire _3277_;
wire _3278_;
wire _3279_;
wire _3280_;
wire _3281_;
wire _3282_;
wire _3283_;
wire _3284_;
wire _3285_;
wire _3286_;
wire _3287_;
wire _3288_;
wire _3289_;
wire _3290_;
wire _3291_;
wire _3292_;
wire _3293_;
wire _3294_;
wire _3295_;
wire _3296_;
wire _3297_;
wire _3298_;
wire _3299_;
wire _3300_;
wire _3301_;
wire _3302_;
wire _3303_;
wire _3304_;
wire _3305_;
wire _3306_;
wire _3307_;
wire _3308_;
wire _3309_;
wire _3310_;
wire _3311_;
wire _3312_;
wire _3313_;
wire _3314_;
wire _3315_;
wire _3316_;
wire _3317_;
wire _3318_;
wire _3319_;
wire _3320_;
wire _3321_;
wire _3322_;
wire _3323_;
wire _3324_;
wire _3325_;
wire _3326_;
wire _3327_;
wire _3328_;
wire _3329_;
wire _3330_;
wire _3331_;
wire _3332_;
wire _3333_;
wire _3334_;
wire _3335_;
wire _3336_;
wire _3337_;
wire _3338_;
wire _3339_;
wire _3340_;
wire _3341_;
wire _3342_;
wire _3343_;
wire _3344_;
wire _3345_;
wire _3346_;
wire _3347_;
wire _3348_;
wire _3349_;
wire _3350_;
wire _3351_;
wire _3352_;
wire _3353_;
wire _3354_;
wire _3355_;
wire _3356_;
wire _3357_;
wire _3358_;
wire _3359_;
wire _3360_;
wire _3361_;
wire _3362_;
wire _3363_;
wire _3364_;
wire _3365_;
wire _3366_;
wire _3367_;
wire _3368_;
wire _3369_;
wire _3370_;
wire _3371_;
wire _3372_;
wire _3373_;
wire _3374_;
wire _3375_;
wire _3376_;
wire _3377_;
wire _3378_;
wire _3379_;
wire _3380_;
wire _3381_;
wire _3382_;
wire _3383_;
wire _3384_;
wire _3385_;
wire _3386_;
wire _3387_;
wire _3388_;
wire _3389_;
wire _3390_;
wire _3391_;
wire _3392_;
wire _3393_;
wire _3394_;
wire _3395_;
wire _3396_;
wire _3397_;
wire _3398_;
wire _3399_;
wire _3400_;
wire _3401_;
wire _3402_;
wire _3403_;
wire _3404_;
wire _3405_;
wire _3406_;
wire _3407_;
wire _3408_;
wire _3409_;
wire _3410_;
wire _3411_;
wire _3412_;
wire _3413_;
wire _3414_;
wire _3415_;
wire _3416_;
wire _3417_;
wire _3418_;
wire _3419_;
wire _3420_;
wire _3421_;
wire _3422_;
wire _3423_;
wire _3424_;
wire _3425_;
wire _3426_;
wire _3427_;
wire _3428_;
wire _3429_;
wire _3430_;
wire _3431_;
wire _3432_;
wire _3433_;
wire _3434_;
wire _3435_;
wire _3436_;
wire _3437_;
wire _3438_;
wire _3439_;
wire _3440_;
wire _3441_;
wire _3442_;
wire _3443_;
wire _3444_;
wire _3445_;
wire _3446_;
wire _3447_;
wire _3448_;
wire _3449_;
wire _3450_;
wire _3451_;
wire _3452_;
wire _3453_;
wire _3454_;
wire _3455_;
wire _3456_;
wire _3457_;
wire _3458_;
wire _3459_;
wire _3460_;
wire _3461_;
wire _3462_;
wire _3463_;
wire _3464_;
wire _3465_;
wire _3466_;
wire _3467_;
wire _3468_;
wire _3469_;
wire _3470_;
wire _3471_;
wire _3472_;
wire _3473_;
wire _3474_;
wire _3475_;
wire _3476_;
wire _3477_;
wire _3478_;
wire _3479_;
wire _3480_;
wire _3481_;
wire _3482_;
wire _3483_;
wire _3484_;
wire _3485_;
wire _3486_;
wire _3487_;
wire _3488_;
wire _3489_;
wire _3490_;
wire _3491_;
wire _3492_;
wire _3493_;
wire _3494_;
wire _3495_;
wire _3496_;
wire _3497_;
wire _3498_;
wire _3499_;
wire _3500_;
wire _3501_;
wire _3502_;
wire _3503_;
wire _3504_;
wire _3505_;
wire _3506_;
wire _3507_;
wire _3508_;
wire _3509_;
wire _3510_;
wire _3511_;
wire _3512_;
wire _3513_;
wire _3514_;
wire _3515_;
wire _3516_;
wire _3517_;
wire _3518_;
wire _3519_;
wire _3520_;
wire _3521_;
wire _3522_;
wire _3523_;
wire _3524_;
wire _3525_;
wire _3526_;
wire _3527_;
wire _3528_;
wire _3529_;
wire _3530_;
wire _3531_;
wire _3532_;
wire _3533_;
wire _3534_;
wire _3535_;
wire _3536_;
wire _3537_;
wire _3538_;
wire _3539_;
wire _3540_;
wire _3541_;
wire _3542_;
wire _3543_;
wire _3544_;
wire _3545_;
wire _3546_;
wire _3547_;
wire _3548_;
wire _3549_;
wire _3550_;
wire _3551_;
wire _3552_;
wire _3553_;
wire _3554_;
wire _3555_;
wire _3556_;
wire _3557_;
wire _3558_;
wire _3559_;
wire _3560_;
wire _3561_;
wire _3562_;
wire _3563_;
wire _3564_;
wire _3565_;
wire _3566_;
wire _3567_;
wire _3568_;
wire _3569_;
wire _3570_;
wire _3571_;
wire _3572_;
wire _3573_;
wire _3574_;
wire _3575_;
wire _3576_;
wire _3577_;
wire _3578_;
wire _3579_;
wire _3580_;
wire _3581_;
wire _3582_;
wire _3583_;
wire _3584_;
wire _3585_;
wire _3586_;
wire _3587_;
wire _3588_;
wire _3589_;
wire _3590_;
wire _3591_;
wire _3592_;
wire _3593_;
wire _3594_;
wire _3595_;
wire _3596_;
wire _3597_;
wire _3598_;
wire _3599_;
wire _3600_;
wire _3601_;
wire _3602_;
wire _3603_;
wire _3604_;
wire _3605_;
wire _3606_;
wire _3607_;
wire _3608_;
wire _3609_;
wire _3610_;
wire _3611_;
wire _3612_;
wire _3613_;
wire _3614_;
wire _3615_;
wire _3616_;
wire _3617_;
wire _3618_;
wire _3619_;
wire _3620_;
wire _3621_;
wire _3622_;
wire _3623_;
wire _3624_;
wire _3625_;
wire _3626_;
wire _3627_;
wire _3628_;
wire _3629_;
wire _3630_;
wire _3631_;
wire _3632_;
wire _3633_;
wire _3634_;
wire _3635_;
wire _3636_;
wire _3637_;
wire _3638_;
wire _3639_;
wire _3640_;
wire _3641_;
wire _3642_;
wire _3643_;
wire _3644_;
wire _3645_;
wire _3646_;
wire _3647_;
wire _3648_;
wire _3649_;
wire _3650_;
wire _3651_;
wire _3652_;
wire _3653_;
wire _3654_;
wire _3655_;
wire _3656_;
wire _3657_;
wire _3658_;
wire _3659_;
wire _3660_;
wire _3661_;
wire _3662_;
wire _3663_;
wire _3664_;
wire _3665_;
wire _3666_;
wire _3667_;
wire _3668_;
wire _3669_;
wire _3670_;
wire _3671_;
wire _3672_;
wire _3673_;
wire _3674_;
wire _3675_;
wire _3676_;
wire _3677_;
wire _3678_;
wire _3679_;
wire _3680_;
wire _3681_;
wire _3682_;
wire _3683_;
wire _3684_;
wire _3685_;
wire _3686_;
wire _3687_;
wire _3688_;
wire _3689_;
wire _3690_;
wire _3691_;
wire _3692_;
wire _3693_;
wire _3694_;
wire _3695_;
wire _3696_;
wire _3697_;
wire _3698_;
wire _3699_;
wire _3700_;
wire _3701_;
wire _3702_;
wire _3703_;
wire _3704_;
wire _3705_;
wire _3706_;
wire _3707_;
wire _3708_;
wire _3709_;
wire _3710_;
wire _3711_;
wire _3712_;
wire _3713_;
wire _3714_;
wire _3715_;
wire _3716_;
wire _3717_;
wire _3718_;
wire _3719_;
wire _3720_;
wire _3721_;
wire _3722_;
wire _3723_;
wire _3724_;
wire _3725_;
wire _3726_;
wire _3727_;
wire _3728_;
wire _3729_;
wire _3730_;
wire _3731_;
wire _3732_;
wire _3733_;
wire _3734_;
wire _3735_;
wire _3736_;
wire _3737_;
wire _3738_;
wire _3739_;
wire _3740_;
wire _3741_;
wire _3742_;
wire _3743_;
wire _3744_;
wire _3745_;
wire _3746_;
wire _3747_;
wire _3748_;
wire _3749_;
wire _3750_;
wire _3751_;
wire _3752_;
wire _3753_;
wire _3754_;
wire _3755_;
wire _3756_;
wire _3757_;
wire _3758_;
wire _3759_;
wire _3760_;
wire _3761_;
wire _3762_;
wire _3763_;
wire _3764_;
wire _3765_;
wire _3766_;
wire _3767_;
wire _3768_;
wire _3769_;
wire _3770_;
wire _3771_;
wire _3772_;
wire _3773_;
wire _3774_;
wire _3775_;
wire _3776_;
wire _3777_;
wire _3778_;
wire _3779_;
wire _3780_;
wire _3781_;
wire _3782_;
wire _3783_;
wire _3784_;
wire _3785_;
wire _3786_;
wire _3787_;
wire _3788_;
wire _3789_;
wire _3790_;
wire _3791_;
wire _3792_;
wire _3793_;
wire _3794_;
wire _3795_;
wire _3796_;
wire _3797_;
wire _3798_;
wire _3799_;
wire _3800_;
wire _3801_;
wire _3802_;
wire _3803_;
wire _3804_;
wire _3805_;
wire _3806_;
wire _3807_;
wire _3808_;
wire _3809_;
wire _3810_;
wire _3811_;
wire _3812_;
wire _3813_;
wire _3814_;
wire _3815_;
wire _3816_;
wire _3817_;
wire _3818_;
wire _3819_;
wire _3820_;
wire _3821_;
wire _3822_;
wire _3823_;
wire _3824_;
wire _3825_;
wire _3826_;
wire _3827_;
wire _3828_;
wire _3829_;
wire _3830_;
wire _3831_;
wire _3832_;
wire _3833_;
wire _3834_;
wire _3835_;
wire _3836_;
wire _3837_;
wire _3838_;
wire _3839_;
wire _3840_;
wire _3841_;
wire _3842_;
wire _3843_;
wire _3844_;
wire _3845_;
wire _3846_;
wire _3847_;
wire _3848_;
wire _3849_;
wire _3850_;
wire _3851_;
wire _3852_;
wire _3853_;
wire _3854_;
wire _3855_;
wire _3856_;
wire _3857_;
wire _3858_;
wire _3859_;
wire _3860_;
wire _3861_;
wire _3862_;
wire _3863_;
wire _3864_;
wire _3865_;
wire _3866_;
wire _3867_;
wire _3868_;
wire _3869_;
wire _3870_;
wire _3871_;
wire _3872_;
wire _3873_;
wire _3874_;
wire _3875_;
wire _3876_;
wire _3877_;
wire _3878_;
wire _3879_;
wire _3880_;
wire _3881_;
wire _3882_;
wire _3883_;
wire _3884_;
wire _3885_;
wire _3886_;
wire _3887_;
wire _3888_;
wire _3889_;
wire _3890_;
wire _3891_;
wire _3892_;
wire _3893_;
wire _3894_;
wire _3895_;
wire _3896_;
wire _3897_;
wire _3898_;
wire _3899_;
wire _3900_;
wire _3901_;
wire _3902_;
wire _3903_;
wire _3904_;
wire _3905_;
wire _3906_;
wire _3907_;
wire _3908_;
wire _3909_;
wire _3910_;
wire _3911_;
wire _3912_;
wire _3913_;
wire _3914_;
wire _3915_;
wire _3916_;
wire _3917_;
wire _3918_;
wire _3919_;
wire _3920_;
wire _3921_;
wire _3922_;
wire _3923_;
wire _3924_;
wire _3925_;
wire _3926_;
wire _3927_;
wire _3928_;
wire _3929_;
wire _3930_;
wire _3931_;
wire _3932_;
wire _3933_;
wire _3934_;
wire _3935_;
wire _3936_;
wire _3937_;
wire _3938_;
wire _3939_;
wire _3940_;
wire _3941_;
wire _3942_;
wire _3943_;
wire _3944_;
wire _3945_;
wire _3946_;
wire _3947_;
wire _3948_;
wire _3949_;
wire _3950_;
wire _3951_;
wire _3952_;
wire _3953_;
wire _3954_;
wire _3955_;
wire _3956_;
wire _3957_;
wire _3958_;
wire _3959_;
wire _3960_;
wire _3961_;
wire _3962_;
wire _3963_;
wire _3964_;
wire _3965_;
wire _3966_;
wire _3967_;
wire _3968_;
wire _3969_;
wire _3970_;
wire _3971_;
wire _3972_;
wire _3973_;
wire _3974_;
wire _3975_;
wire _3976_;
wire _3977_;
wire _3978_;
wire _3979_;
wire _3980_;
wire _3981_;
wire _3982_;
wire _3983_;
wire _3984_;
wire _3985_;
wire _3986_;
wire _3987_;
wire _3988_;
wire _3989_;
wire _3990_;
wire _3991_;
wire _3992_;
wire _3993_;
wire _3994_;
wire _3995_;
wire _3996_;
wire _3997_;
wire _3998_;
wire _3999_;
wire _4000_;
wire _4001_;
wire _4002_;
wire _4003_;
wire _4004_;
wire _4005_;
wire _4006_;
wire _4007_;
wire _4008_;
wire _4009_;
wire _4010_;
wire _4011_;
wire _4012_;
wire _4013_;
wire _4014_;
wire _4015_;
wire _4016_;
wire _4017_;
wire _4018_;
wire _4019_;
wire _4020_;
wire _4021_;
wire _4022_;
wire _4023_;
wire _4024_;
wire _4025_;
wire _4026_;
wire _4027_;
wire _4028_;
wire _4029_;
wire _4030_;
wire _4031_;
wire _4032_;
wire _4033_;
wire _4034_;
wire _4035_;
wire _4036_;
wire _4037_;
wire _4038_;
wire _4039_;
wire _4040_;
wire _4041_;
wire _4042_;
wire _4043_;
wire _4044_;
wire _4045_;
wire _4046_;
wire _4047_;
wire _4048_;
wire _4049_;
wire _4050_;
wire _4051_;
wire _4052_;
wire _4053_;
wire _4054_;
wire _4055_;
wire _4056_;
wire _4057_;
wire _4058_;
wire _4059_;
wire _4060_;
wire _4061_;
wire _4062_;
wire _4063_;
wire _4064_;
wire _4065_;
wire _4066_;
wire _4067_;
wire _4068_;
wire _4069_;
wire _4070_;
wire _4071_;
wire _4072_;
wire _4073_;
wire _4074_;
wire _4075_;
wire _4076_;
wire _4077_;
wire _4078_;
wire _4079_;
wire _4080_;
wire _4081_;
wire _4082_;
wire _4083_;
wire _4084_;
wire _4085_;
wire _4086_;
wire _4087_;
wire _4088_;
wire _4089_;
wire _4090_;
wire _4091_;
wire _4092_;
wire _4093_;
wire _4094_;
wire _4095_;
wire _4096_;
wire _4097_;
wire _4098_;
wire _4099_;
wire _4100_;
wire _4101_;
wire _4102_;
wire _4103_;
wire _4104_;
wire _4105_;
wire _4106_;
wire _4107_;
wire _4108_;
wire _4109_;
wire _4110_;
wire _4111_;
wire _4112_;
wire _4113_;
wire _4114_;
wire _4115_;
wire _4116_;
wire _4117_;
wire _4118_;
wire _4119_;
wire _4120_;
wire _4121_;
wire _4122_;
wire _4123_;
wire _4124_;
wire _4125_;
wire _4126_;
wire _4127_;
wire _4128_;
wire _4129_;
wire _4130_;
wire _4131_;
wire _4132_;
wire _4133_;
wire _4134_;
wire _4135_;
wire _4136_;
wire _4137_;
wire _4138_;
wire _4139_;
wire _4140_;
wire _4141_;
wire _4142_;
wire _4143_;
wire _4144_;
wire _4145_;
wire _4146_;
wire _4147_;
wire _4148_;
wire _4149_;
wire _4150_;
wire _4151_;
wire _4152_;
wire _4153_;
wire _4154_;
wire _4155_;
wire _4156_;
wire _4157_;
wire _4158_;
wire _4159_;
wire _4160_;
wire _4161_;
wire _4162_;
wire _4163_;
wire _4164_;
wire _4165_;
wire _4166_;
wire _4167_;
wire _4168_;
wire _4169_;
wire _4170_;
wire _4171_;
wire _4172_;
wire _4173_;
wire _4174_;
wire _4175_;
wire _4176_;
wire _4177_;
wire _4178_;
wire _4179_;
wire _4180_;
wire _4181_;
wire _4182_;
wire _4183_;
wire _4184_;
wire _4185_;
wire _4186_;
wire _4187_;
wire _4188_;
wire _4189_;
wire _4190_;
wire _4191_;
wire _4192_;
wire _4193_;
wire _4194_;
wire _4195_;
wire _4196_;
wire _4197_;
wire _4198_;
wire _4199_;
wire _4200_;
wire _4201_;
wire _4202_;
wire _4203_;
wire _4204_;
wire _4205_;
wire _4206_;
wire _4207_;
wire _4208_;
wire _4209_;
wire _4210_;
wire _4211_;
wire _4212_;
wire _4213_;
wire _4214_;
wire _4215_;
wire _4216_;
wire _4217_;
wire _4218_;
wire _4219_;
wire _4220_;
wire _4221_;
wire _4222_;
wire _4223_;
wire _4224_;
wire _4225_;
wire _4226_;
wire _4227_;
wire _4228_;
wire _4229_;
wire _4230_;
wire _4231_;
wire _4232_;
wire _4233_;
wire _4234_;
wire _4235_;
wire _4236_;
wire _4237_;
wire _4238_;
wire _4239_;
wire _4240_;
wire _4241_;
wire _4242_;
wire _4243_;
wire _4244_;
wire _4245_;
wire _4246_;
wire _4247_;
wire _4248_;
wire _4249_;
wire _4250_;
wire _4251_;
wire _4252_;
wire _4253_;
wire _4254_;
wire _4255_;
wire _4256_;
wire _4257_;
wire _4258_;
wire _4259_;
wire _4260_;
wire _4261_;
wire _4262_;
wire _4263_;
wire _4264_;
wire _4265_;
wire _4266_;
wire _4267_;
wire _4268_;
wire _4269_;
wire _4270_;
wire _4271_;
wire _4272_;
wire _4273_;
wire _4274_;
wire _4275_;
wire _4276_;
wire _4277_;
wire _4278_;
wire _4279_;
wire _4280_;
wire _4281_;
wire _4282_;
wire _4283_;
wire _4284_;
wire _4285_;
wire _4286_;
wire _4287_;
wire _4288_;
wire _4289_;
wire _4290_;
wire _4291_;
wire _4292_;
wire _4293_;
wire _4294_;
wire _4295_;
wire _4296_;
wire _4297_;
wire _4298_;
wire _4299_;
wire _4300_;
wire _4301_;
wire _4302_;
wire _4303_;
wire _4304_;
wire _4305_;
wire _4306_;
wire _4307_;
wire _4308_;
wire _4309_;
wire _4310_;
wire _4311_;
wire _4312_;
wire _4313_;
wire _4314_;
wire _4315_;
wire _4316_;
wire _4317_;
wire _4318_;
wire _4319_;
wire _4320_;
wire _4321_;
wire _4322_;
wire _4323_;
wire _4324_;
wire _4325_;
wire _4326_;
wire _4327_;
wire _4328_;
wire _4329_;
wire _4330_;
wire _4331_;
wire _4332_;
wire _4333_;
wire _4334_;
wire _4335_;
wire _4336_;
wire _4337_;
wire _4338_;
wire _4339_;
wire _4340_;
wire _4341_;
wire _4342_;
wire _4343_;
wire _4344_;
wire _4345_;
wire _4346_;
wire _4347_;
wire _4348_;
wire _4349_;
wire _4350_;
wire _4351_;
wire _4352_;
wire _4353_;
wire _4354_;
wire _4355_;
wire _4356_;
wire _4357_;
wire _4358_;
wire _4359_;
wire _4360_;
wire _4361_;
wire _4362_;
wire _4363_;
wire _4364_;
wire _4365_;
wire _4366_;
wire _4367_;
wire _4368_;
wire _4369_;
wire _4370_;
wire _4371_;
wire _4372_;
wire _4373_;
wire _4374_;
wire _4375_;
wire _4376_;
wire _4377_;
wire _4378_;
wire _4379_;
wire _4380_;
wire _4381_;
wire _4382_;
wire _4383_;
wire _4384_;
wire _4385_;
wire _4386_;
wire _4387_;
wire _4388_;
wire _4389_;
wire _4390_;
wire _4391_;
wire _4392_;
wire _4393_;
wire _4394_;
wire _4395_;
wire _4396_;
wire _4397_;
wire _4398_;
wire _4399_;
wire _4400_;
wire _4401_;
wire _4402_;
wire _4403_;
wire _4404_;
wire _4405_;
wire _4406_;
wire _4407_;
wire _4408_;
wire _4409_;
wire _4410_;
wire _4411_;
wire _4412_;
wire _4413_;
wire _4414_;
wire _4415_;
wire _4416_;
wire _4417_;
wire _4418_;
wire _4419_;
wire _4420_;
wire _4421_;
wire _4422_;
wire _4423_;
wire _4424_;
wire _4425_;
wire _4426_;
wire _4427_;
wire _4428_;
wire _4429_;
wire _4430_;
wire _4431_;
wire _4432_;
wire _4433_;
wire _4434_;
wire _4435_;
wire _4436_;
wire _4437_;
wire _4438_;
wire _4439_;
wire _4440_;
wire _4441_;
wire _4442_;
wire _4443_;
wire _4444_;
wire _4445_;
wire _4446_;
wire _4447_;
wire _4448_;
wire _4449_;
wire _4450_;
wire _4451_;
wire _4452_;
wire _4453_;
wire _4454_;
wire _4455_;
wire _4456_;
wire _4457_;
wire _4458_;
wire _4459_;
wire _4460_;
wire _4461_;
wire _4462_;
wire _4463_;
wire _4464_;
wire _4465_;
wire _4466_;
wire _4467_;
wire _4468_;
wire _4469_;
wire _4470_;
wire _4471_;
wire _4472_;
wire _4473_;
wire _4474_;
wire _4475_;
wire _4476_;
wire _4477_;
wire _4478_;
wire _4479_;
wire _4480_;
wire _4481_;
wire _4482_;
wire _4483_;
wire _4484_;
wire _4485_;
wire _4486_;
wire _4487_;
wire _4488_;
wire _4489_;
wire _4490_;
wire _4491_;
wire _4492_;
wire _4493_;
wire _4494_;
wire _4495_;
wire _4496_;
wire _4497_;
wire _4498_;
wire _4499_;
wire _4500_;
wire _4501_;
wire _4502_;
wire _4503_;
wire _4504_;
wire _4505_;
wire _4506_;
wire _4507_;
wire _4508_;
wire _4509_;
wire _4510_;
wire _4511_;
wire _4512_;
wire _4513_;
wire _4514_;
wire _4515_;
wire _4516_;
wire _4517_;
wire _4518_;
wire _4519_;
wire _4520_;
wire _4521_;
wire _4522_;
wire _4523_;
wire _4524_;
wire _4525_;
wire _4526_;
wire _4527_;
wire _4528_;
wire _4529_;
wire _4530_;
wire _4531_;
wire _4532_;
wire _4533_;
wire _4534_;
wire _4535_;
wire _4536_;
wire _4537_;
wire _4538_;
wire _4539_;
wire _4540_;
wire _4541_;
wire _4542_;
wire _4543_;
wire _4544_;
wire _4545_;
wire _4546_;
wire _4547_;
wire _4548_;
wire _4549_;
wire _4550_;
wire _4551_;
wire _4552_;
wire _4553_;
wire _4554_;
wire _4555_;
wire _4556_;
wire _4557_;
wire _4558_;
wire _4559_;
wire _4560_;
wire _4561_;
wire _4562_;
wire _4563_;
wire _4564_;
wire _4565_;
wire _4566_;
wire _4567_;
wire _4568_;
wire _4569_;
wire _4570_;
wire _4571_;
wire _4572_;
wire _4573_;
wire _4574_;
wire _4575_;
wire _4576_;
wire _4577_;
wire _4578_;
wire _4579_;
wire _4580_;
wire _4581_;
wire _4582_;
wire _4583_;
wire _4584_;
wire _4585_;
wire _4586_;
wire _4587_;
wire _4588_;
wire _4589_;
wire _4590_;
wire _4591_;
wire _4592_;
wire _4593_;
wire _4594_;
wire _4595_;
wire _4596_;
wire _4597_;
wire _4598_;
wire _4599_;
wire _4600_;
wire _4601_;
wire _4602_;
wire _4603_;
wire _4604_;
wire _4605_;
wire _4606_;
wire _4607_;
wire _4608_;
wire _4609_;
wire _4610_;
wire _4611_;
wire _4612_;
wire _4613_;
wire _4614_;
wire _4615_;
wire _4616_;
wire _4617_;
wire _4618_;
wire _4619_;
wire _4620_;
wire _4621_;
wire _4622_;
wire _4623_;
wire _4624_;
wire _4625_;
wire _4626_;
wire _4627_;
wire _4628_;
wire _4629_;
wire _4630_;
wire _4631_;
wire _4632_;
wire _4633_;
wire _4634_;
wire _4635_;
wire _4636_;
wire _4637_;
wire _4638_;
wire _4639_;
wire _4640_;
wire _4641_;
wire _4642_;
wire _4643_;
wire _4644_;
wire _4645_;
wire _4646_;
wire _4647_;
wire _4648_;
wire _4649_;
wire _4650_;
wire _4651_;
wire _4652_;
wire _4653_;
wire _4654_;
wire _4655_;
wire _4656_;
wire _4657_;
wire _4658_;
wire _4659_;
wire _4660_;
wire _4661_;
wire _4662_;
wire _4663_;
wire _4664_;
wire _4665_;
wire _4666_;
wire _4667_;
wire _4668_;
wire _4669_;
wire _4670_;
wire _4671_;
wire _4672_;
wire _4673_;
wire _4674_;
wire _4675_;
wire _4676_;
wire _4677_;
wire _4678_;
wire _4679_;
wire _4680_;
wire _4681_;
wire _4682_;
wire _4683_;
wire _4684_;
wire _4685_;
wire _4686_;
wire _4687_;
wire _4688_;
wire _4689_;
wire _4690_;
wire _4691_;
wire _4692_;
wire _4693_;
wire _4694_;
wire _4695_;
wire _4696_;
wire _4697_;
wire _4698_;
wire _4699_;
wire _4700_;
wire _4701_;
wire _4702_;
wire _4703_;
wire _4704_;
wire _4705_;
wire _4706_;
wire _4707_;
wire _4708_;
wire _4709_;
wire _4710_;
wire _4711_;
wire _4712_;
wire _4713_;
wire _4714_;
wire _4715_;
wire _4716_;
wire _4717_;
wire _4718_;
wire _4719_;
wire _4720_;
wire _4721_;
wire _4722_;
wire _4723_;
wire _4724_;
wire _4725_;
wire _4726_;
wire _4727_;
wire _4728_;
wire _4729_;
wire _4730_;
wire _4731_;
wire _4732_;
wire _4733_;
wire _4734_;
wire _4735_;
wire _4736_;
wire _4737_;
wire _4738_;
wire _4739_;
wire _4740_;
wire _4741_;
wire _4742_;
wire _4743_;
wire _4744_;
wire _4745_;
wire _4746_;
wire _4747_;
wire _4748_;
wire _4749_;
wire _4750_;
wire _4751_;
wire _4752_;
wire _4753_;
wire _4754_;
wire _4755_;
wire _4756_;
wire _4757_;
wire _4758_;
wire _4759_;
wire _4760_;
wire _4761_;
wire _4762_;
wire _4763_;
wire _4764_;
wire _4765_;
wire _4766_;
wire _4767_;
wire _4768_;
wire _4769_;
wire _4770_;
wire _4771_;
wire _4772_;
wire _4773_;
wire _4774_;
wire _4775_;
wire _4776_;
wire _4777_;
wire _4778_;
wire _4779_;
wire _4780_;
wire _4781_;
wire _4782_;
wire _4783_;
wire _4784_;
wire _4785_;
wire _4786_;
wire _4787_;
wire _4788_;
wire _4789_;
wire _4790_;
wire _4791_;
wire _4792_;
wire _4793_;
wire _4794_;
wire _4795_;
wire _4796_;
wire _4797_;
wire _4798_;
wire _4799_;
wire _4800_;
wire _4801_;
wire _4802_;
wire _4803_;
wire _4804_;
wire _4805_;
wire _4806_;
wire _4807_;
wire _4808_;
wire _4809_;
wire _4810_;
wire _4811_;
wire _4812_;
wire _4813_;
wire _4814_;
wire _4815_;
wire _4816_;
wire _4817_;
wire _4818_;
wire _4819_;
wire _4820_;
wire _4821_;
wire _4822_;
wire _4823_;
wire _4824_;
wire _4825_;
wire _4826_;
wire _4827_;
wire _4828_;
wire _4829_;
wire _4830_;
wire _4831_;
wire _4832_;
wire _4833_;
wire _4834_;
wire _4835_;
wire _4836_;
wire _4837_;
wire _4838_;
wire _4839_;
wire _4840_;
wire _4841_;
wire _4842_;
wire _4843_;
wire _4844_;
wire _4845_;
wire _4846_;
wire _4847_;
wire _4848_;
wire _4849_;
wire _4850_;
wire _4851_;
wire _4852_;
wire _4853_;
wire _4854_;
wire _4855_;
wire _4856_;
wire _4857_;
wire _4858_;
wire _4859_;
wire _4860_;
wire _4861_;
wire _4862_;
wire _4863_;
wire _4864_;
wire _4865_;
wire _4866_;
wire _4867_;
wire _4868_;
wire _4869_;
wire _4870_;
wire _4871_;
wire _4872_;
wire _4873_;
wire _4874_;
wire _4875_;
wire _4876_;
wire _4877_;
wire _4878_;
wire _4879_;
wire _4880_;
wire _4881_;
wire _4882_;
wire _4883_;
wire _4884_;
wire _4885_;
wire _4886_;
wire _4887_;
wire _4888_;
wire _4889_;
wire _4890_;
wire _4891_;
wire _4892_;
wire _4893_;
wire _4894_;
wire _4895_;
wire _4896_;
wire _4897_;
wire _4898_;
wire _4899_;
wire _4900_;
wire _4901_;
wire _4902_;
wire _4903_;
wire _4904_;
wire _4905_;
wire _4906_;
wire _4907_;
wire _4908_;
wire _4909_;
wire _4910_;
wire _4911_;
wire _4912_;
wire _4913_;
wire _4914_;
wire _4915_;
wire _4916_;
wire _4917_;
wire _4918_;
wire _4919_;
wire _4920_;
wire _4921_;
wire _4922_;
wire _4923_;
wire _4924_;
wire _4925_;
wire _4926_;
wire _4927_;
wire _4928_;
wire _4929_;
wire _4930_;
wire _4931_;
wire _4932_;
wire _4933_;
wire _4934_;
wire _4935_;
wire _4936_;
wire _4937_;
wire _4938_;
wire _4939_;
wire _4940_;
wire _4941_;
wire _4942_;
wire _4943_;
wire _4944_;
wire _4945_;
wire _4946_;
wire _4947_;
wire _4948_;
wire _4949_;
wire _4950_;
wire _4951_;
wire _4952_;
wire _4953_;
wire _4954_;
wire _4955_;
wire _4956_;
wire _4957_;
wire _4958_;
wire _4959_;
wire _4960_;
wire _4961_;
wire _4962_;
wire _4963_;
wire _4964_;
wire _4965_;
wire _4966_;
wire _4967_;
wire _4968_;
wire _4969_;
wire _4970_;
wire _4971_;
wire _4972_;
wire _4973_;
wire _4974_;
wire _4975_;
wire _4976_;
wire _4977_;
wire _4978_;
wire _4979_;
wire _4980_;
wire _4981_;
wire _4982_;
wire _4983_;
wire _4984_;
wire _4985_;
wire _4986_;
wire _4987_;
wire _4988_;
wire _4989_;
wire _4990_;
wire _4991_;
wire _4992_;
wire _4993_;
wire _4994_;
wire _4995_;
wire _4996_;
wire _4997_;
wire _4998_;
wire _4999_;
wire _5000_;
wire _5001_;
wire _5002_;
wire _5003_;
wire _5004_;
wire _5005_;
wire _5006_;
wire _5007_;
wire _5008_;
wire _5009_;
wire _5010_;
wire _5011_;
wire _5012_;
wire _5013_;
wire _5014_;
wire _5015_;
wire _5016_;
wire _5017_;
wire _5018_;
wire _5019_;
wire _5020_;
wire _5021_;
wire _5022_;
wire _5023_;
wire _5024_;
wire _5025_;
wire _5026_;
wire _5027_;
wire _5028_;
wire _5029_;
wire _5030_;
wire _5031_;
wire _5032_;
wire _5033_;
wire _5034_;
wire _5035_;
wire _5036_;
wire _5037_;
wire _5038_;
wire _5039_;
wire _5040_;
wire _5041_;
wire _5042_;
wire _5043_;
wire _5044_;
wire _5045_;
wire _5046_;
wire _5047_;
wire _5048_;
wire _5049_;
wire _5050_;
wire _5051_;
wire _5052_;
wire _5053_;
wire _5054_;
wire _5055_;
wire _5056_;
wire _5057_;
wire _5058_;
wire _5059_;
wire _5060_;
wire _5061_;
wire _5062_;
wire _5063_;
wire _5064_;
wire _5065_;
wire _5066_;
wire _5067_;
wire _5068_;
wire _5069_;
wire _5070_;
wire _5071_;
wire _5072_;
wire _5073_;
wire _5074_;
wire _5075_;
wire _5076_;
wire _5077_;
wire _5078_;
wire _5079_;
wire _5080_;
wire _5081_;
wire _5082_;
wire _5083_;
wire _5084_;
wire _5085_;
wire _5086_;
wire _5087_;
wire _5088_;
wire _5089_;
wire _5090_;
wire _5091_;
wire _5092_;
wire _5093_;
wire _5094_;
wire _5095_;
wire _5096_;
wire _5097_;
wire _5098_;
wire _5099_;
wire _5100_;
wire _5101_;
wire _5102_;
wire _5103_;
wire _5104_;
wire _5105_;
wire _5106_;
wire _5107_;
wire _5108_;
wire _5109_;
wire _5110_;
wire _5111_;
wire _5112_;
wire _5113_;
wire _5114_;
wire _5115_;
wire _5116_;
wire _5117_;
wire _5118_;
wire _5119_;
wire _5120_;
wire _5121_;
wire _5122_;
wire _5123_;
wire _5124_;
wire _5125_;
wire _5126_;
wire _5127_;
wire _5128_;
wire _5129_;
wire _5130_;
wire _5131_;
wire _5132_;
wire _5133_;
wire _5134_;
wire _5135_;
wire _5136_;
wire _5137_;
wire _5138_;
wire _5139_;
wire _5140_;
wire _5141_;
wire _5142_;
wire _5143_;
wire _5144_;
wire _5145_;
wire _5146_;
wire _5147_;
wire _5148_;
wire _5149_;
wire _5150_;
wire _5151_;
wire _5152_;
wire _5153_;
wire _5154_;
wire _5155_;
wire _5156_;
wire _5157_;
wire _5158_;
wire _5159_;
wire _5160_;
wire _5161_;
wire _5162_;
wire _5163_;
wire _5164_;
wire _5165_;
wire _5166_;
wire _5167_;
wire _5168_;
wire _5169_;
wire _5170_;
wire _5171_;
wire _5172_;
wire _5173_;
wire _5174_;
wire _5175_;
wire _5176_;
wire _5177_;
wire _5178_;
wire _5179_;
wire _5180_;
wire _5181_;
wire _5182_;
wire _5183_;
wire _5184_;
wire _5185_;
wire _5186_;
wire _5187_;
wire _5188_;
wire _5189_;
wire _5190_;
wire _5191_;
wire _5192_;
wire _5193_;
wire _5194_;
wire _5195_;
wire _5196_;
wire _5197_;
wire _5198_;
wire _5199_;
wire _5200_;
wire _5201_;
wire _5202_;
wire _5203_;
wire _5204_;
wire _5205_;
wire _5206_;
wire _5207_;
wire _5208_;
wire _5209_;
wire _5210_;
wire _5211_;
wire _5212_;
wire _5213_;
wire _5214_;
wire _5215_;
wire _5216_;
wire _5217_;
wire _5218_;
wire _5219_;
wire _5220_;
wire _5221_;
wire _5222_;
wire _5223_;
wire _5224_;
wire _5225_;
wire _5226_;
wire _5227_;
wire _5228_;
wire _5229_;
wire _5230_;
wire _5231_;
wire _5232_;
wire _5233_;
wire _5234_;
wire _5235_;
wire _5236_;
wire _5237_;
wire _5238_;
wire _5239_;
wire _5240_;
wire _5241_;
wire _5242_;
wire _5243_;
wire _5244_;
wire _5245_;
wire _5246_;
wire _5247_;
wire _5248_;
wire _5249_;
wire _5250_;
wire _5251_;
wire _5252_;
wire _5253_;
wire _5254_;
wire _5255_;
wire _5256_;
wire _5257_;
wire _5258_;
wire _5259_;
wire _5260_;
wire _5261_;
wire _5262_;
wire _5263_;
wire _5264_;
wire _5265_;
wire _5266_;
wire _5267_;
wire _5268_;
wire _5269_;
wire _5270_;
wire _5271_;
wire _5272_;
wire _5273_;
wire _5274_;
wire _5275_;
wire _5276_;
wire _5277_;
wire _5278_;
wire _5279_;
wire _5280_;
wire _5281_;
wire _5282_;
wire _5283_;
wire _5284_;
wire _5285_;
wire _5286_;
wire _5287_;
wire _5288_;
wire _5289_;
wire _5290_;
wire _5291_;
wire _5292_;
wire _5293_;
wire _5294_;
wire _5295_;
wire _5296_;
wire _5297_;
wire _5298_;
wire _5299_;
wire _5300_;
wire _5301_;
wire _5302_;
wire _5303_;
wire _5304_;
wire _5305_;
wire _5306_;
wire _5307_;
wire _5308_;
wire _5309_;
wire _5310_;
wire _5311_;
wire _5312_;
wire _5313_;
wire _5314_;
wire _5315_;
wire _5316_;
wire _5317_;
wire _5318_;
wire _5319_;
wire _5320_;
wire _5321_;
wire _5322_;
wire _5323_;
wire _5324_;
wire _5325_;
wire _5326_;
wire _5327_;
wire _5328_;
wire _5329_;
wire _5330_;
wire _5331_;
wire _5332_;
wire _5333_;
wire _5334_;
wire _5335_;
wire _5336_;
wire _5337_;
wire _5338_;
wire _5339_;
wire _5340_;
wire _5341_;
wire _5342_;
wire _5343_;
wire _5344_;
wire _5345_;
wire _5346_;
wire _5347_;
wire _5348_;
wire _5349_;
wire _5350_;
wire _5351_;
wire _5352_;
wire _5353_;
wire _5354_;
wire _5355_;
wire _5356_;
wire _5357_;
wire _5358_;
wire _5359_;
wire _5360_;
wire _5361_;
wire _5362_;
wire _5363_;
wire _5364_;
wire _5365_;
wire _5366_;
wire _5367_;
wire _5368_;
wire _5369_;
wire _5370_;
wire _5371_;
wire _5372_;
wire _5373_;
wire _5374_;
wire _5375_;
wire _5376_;
wire _5377_;
wire _5378_;
wire _5379_;
wire _5380_;
wire _5381_;
wire _5382_;
wire _5383_;
wire _5384_;
wire _5385_;
wire _5386_;
wire _5387_;
wire _5388_;
wire _5389_;
wire _5390_;
wire _5391_;
wire _5392_;
wire _5393_;
wire _5394_;
wire _5395_;
wire _5396_;
wire _5397_;
wire _5398_;
wire _5399_;
wire _5400_;
wire _5401_;
wire _5402_;
wire _5403_;
wire _5404_;
wire _5405_;
wire _5406_;
wire _5407_;
wire _5408_;
wire _5409_;
wire _5410_;
wire _5411_;
wire _5412_;
wire _5413_;
wire _5414_;
wire _5415_;
wire _5416_;
wire _5417_;
wire _5418_;
wire _5419_;
wire _5420_;
wire _5421_;
wire _5422_;
wire _5423_;
wire _5424_;
wire _5425_;
wire _5426_;
wire _5427_;
wire _5428_;
wire _5429_;
wire _5430_;
wire _5431_;
wire _5432_;
wire _5433_;
wire _5434_;
wire _5435_;
wire _5436_;
wire _5437_;
wire _5438_;
wire _5439_;
wire _5440_;
wire _5441_;
wire _5442_;
wire _5443_;
wire _5444_;
wire _5445_;
wire _5446_;
wire _5447_;
wire _5448_;
wire _5449_;
wire _5450_;
wire _5451_;
wire _5452_;
wire _5453_;
wire _5454_;
wire _5455_;
wire _5456_;
wire _5457_;
wire _5458_;
wire _5459_;
wire _5460_;
wire _5461_;
wire _5462_;
wire _5463_;
wire _5464_;
wire _5465_;
wire _5466_;
wire _5467_;
wire _5468_;
wire _5469_;
wire _5470_;
wire _5471_;
wire _5472_;
wire _5473_;
wire _5474_;
wire _5475_;
wire _5476_;
wire _5477_;
wire _5478_;
wire _5479_;
wire _5480_;
wire _5481_;
wire _5482_;
wire _5483_;
wire _5484_;
wire _5485_;
wire _5486_;
wire _5487_;
wire _5488_;
wire _5489_;
wire _5490_;
wire _5491_;
wire _5492_;
wire _5493_;
wire _5494_;
wire _5495_;
wire _5496_;
wire _5497_;
wire _5498_;
wire _5499_;
wire _5500_;
wire _5501_;
wire _5502_;
wire _5503_;
wire _5504_;
wire _5505_;
wire _5506_;
wire _5507_;
wire _5508_;
wire _5509_;
wire _5510_;
wire _5511_;
wire _5512_;
wire _5513_;
wire _5514_;
wire _5515_;
wire _5516_;
wire _5517_;
wire _5518_;
wire _5519_;
wire _5520_;
wire _5521_;
wire _5522_;
wire _5523_;
wire _5524_;
wire _5525_;
wire _5526_;
wire _5527_;
wire _5528_;
wire _5529_;
wire _5530_;
wire _5531_;
wire _5532_;
wire _5533_;
wire _5534_;
wire _5535_;
wire _5536_;
wire _5537_;
wire _5538_;
wire _5539_;
wire _5540_;
wire _5541_;
wire _5542_;
wire _5543_;
wire _5544_;
wire _5545_;
wire _5546_;
wire _5547_;
wire _5548_;
wire _5549_;
wire _5550_;
wire _5551_;
wire _5552_;
wire _5553_;
wire _5554_;
wire _5555_;
wire _5556_;
wire _5557_;
wire _5558_;
wire _5559_;
wire _5560_;
wire _5561_;
wire _5562_;
wire _5563_;
wire _5564_;
wire _5565_;
wire _5566_;
wire _5567_;
wire _5568_;
wire _5569_;
wire _5570_;
wire _5571_;
wire _5572_;
wire _5573_;
wire _5574_;
wire _5575_;
wire _5576_;
wire _5577_;
wire _5578_;
wire _5579_;
wire _5580_;
wire _5581_;
wire _5582_;
wire _5583_;
wire _5584_;
wire _5585_;
wire _5586_;
wire _5587_;
wire _5588_;
wire _5589_;
wire _5590_;
wire _5591_;
wire _5592_;
wire _5593_;
wire _5594_;
wire _5595_;
wire _5596_;
wire _5597_;
wire _5598_;
wire _5599_;
wire _5600_;
wire _5601_;
wire _5602_;
wire _5603_;
wire _5604_;
wire _5605_;
wire _5606_;
wire _5607_;
wire _5608_;
wire _5609_;
wire _5610_;
wire _5611_;
wire _5612_;
wire _5613_;
wire _5614_;
wire _5615_;
wire _5616_;
wire _5617_;
wire _5618_;
wire _5619_;
wire _5620_;
wire _5621_;
wire _5622_;
wire _5623_;
wire _5624_;
wire _5625_;
wire _5626_;
wire _5627_;
wire _5628_;
wire _5629_;
wire _5630_;
wire _5631_;
wire _5632_;
wire _5633_;
wire _5634_;
wire _5635_;
wire _5636_;
wire _5637_;
wire _5638_;
wire _5639_;
wire _5640_;
wire _5641_;
wire _5642_;
wire _5643_;
wire _5644_;
wire _5645_;
wire _5646_;
wire _5647_;
wire _5648_;
wire _5649_;
wire _5650_;
wire _5651_;
wire _5652_;
wire _5653_;
wire _5654_;
wire _5655_;
wire _5656_;
wire _5657_;
wire _5658_;
wire _5659_;
wire _5660_;
wire _5661_;
wire _5662_;
wire _5663_;
wire _5664_;
wire _5665_;
wire _5666_;
wire _5667_;
wire _5668_;
wire _5669_;
wire _5670_;
wire _5671_;
wire _5672_;
wire _5673_;
wire _5674_;
wire _5675_;
wire _5676_;
wire _5677_;
wire _5678_;
wire _5679_;
wire _5680_;
wire _5681_;
wire _5682_;
wire _5683_;
wire _5684_;
wire _5685_;
wire _5686_;
wire _5687_;
wire _5688_;
wire _5689_;
wire _5690_;
wire _5691_;
wire _5692_;
wire _5693_;
wire _5694_;
wire _5695_;
wire _5696_;
wire _5697_;
wire _5698_;
wire _5699_;
wire _5700_;
wire _5701_;
wire _5702_;
wire _5703_;
wire _5704_;
wire _5705_;
wire _5706_;
wire _5707_;
wire _5708_;
wire _5709_;
wire _5710_;
wire _5711_;
wire _5712_;
wire _5713_;
wire _5714_;
wire _5715_;
wire _5716_;
wire _5717_;
wire _5718_;
wire _5719_;
wire _5720_;
wire _5721_;
wire _5722_;
wire _5723_;
wire _5724_;
wire _5725_;
wire _5726_;
wire _5727_;
wire _5728_;
wire _5729_;
wire _5730_;
wire _5731_;
wire _5732_;
wire _5733_;
wire _5734_;
wire _5735_;
wire _5736_;
wire _5737_;
wire _5738_;
wire _5739_;
wire _5740_;
wire _5741_;
wire _5742_;
wire _5743_;
wire _5744_;
wire _5745_;
wire _5746_;
wire _5747_;
wire _5748_;
wire _5749_;
wire _5750_;
wire _5751_;
wire _5752_;
wire _5753_;
wire _5754_;
wire _5755_;
wire _5756_;
wire _5757_;
wire _5758_;
wire _5759_;
wire _5760_;
wire _5761_;
wire _5762_;
wire _5763_;
wire _5764_;
wire _5765_;
wire _5766_;
wire _5767_;
wire _5768_;
wire _5769_;
wire _5770_;
wire _5771_;
wire _5772_;
wire _5773_;
wire _5774_;
wire _5775_;
wire _5776_;
wire _5777_;
wire _5778_;
wire _5779_;
wire _5780_;
wire _5781_;
wire _5782_;
wire _5783_;
wire _5784_;
wire _5785_;
wire _5786_;
wire _5787_;
wire _5788_;
wire _5789_;
wire _5790_;
wire _5791_;
wire _5792_;
wire _5793_;
wire _5794_;
wire _5795_;
wire _5796_;
wire _5797_;
wire _5798_;
wire _5799_;
wire _5800_;
wire _5801_;
wire _5802_;
wire _5803_;
wire _5804_;
wire _5805_;
wire _5806_;
wire _5807_;
wire _5808_;
wire _5809_;
wire _5810_;
wire _5811_;
wire _5812_;
wire _5813_;
wire _5814_;
wire _5815_;
wire _5816_;
wire _5817_;
wire _5818_;
wire _5819_;
wire _5820_;
wire _5821_;
wire _5822_;
wire _5823_;
wire _5824_;
wire _5825_;
wire _5826_;
wire _5827_;
wire _5828_;
wire _5829_;
wire _5830_;
wire _5831_;
wire _5832_;
wire _5833_;
wire _5834_;
wire _5835_;
wire _5836_;
wire _5837_;
wire _5838_;
wire _5839_;
wire _5840_;
wire _5841_;
wire _5842_;
wire _5843_;
wire _5844_;
wire _5845_;
wire _5846_;
wire _5847_;
wire _5848_;
wire _5849_;
wire _5850_;
wire _5851_;
wire _5852_;
wire _5853_;
wire _5854_;
wire _5855_;
wire _5856_;
wire _5857_;
wire _5858_;
wire _5859_;
wire _5860_;
wire _5861_;
wire _5862_;
wire _5863_;
wire _5864_;
wire _5865_;
wire _5866_;
wire _5867_;
wire _5868_;
wire _5869_;
wire _5870_;
wire _5871_;
wire _5872_;
wire _5873_;
wire _5874_;
wire _5875_;
wire _5876_;
wire _5877_;
wire _5878_;
wire _5879_;
wire _5880_;
wire _5881_;
wire _5882_;
wire _5883_;
wire _5884_;
wire _5885_;
wire _5886_;
wire _5887_;
wire _5888_;
wire _5889_;
wire _5890_;
wire _5891_;
wire _5892_;
wire _5893_;
wire _5894_;
wire _5895_;
wire _5896_;
wire _5897_;
wire _5898_;
wire _5899_;
wire _5900_;
wire _5901_;
wire _5902_;
wire _5903_;
wire _5904_;
wire _5905_;
wire _5906_;
wire _5907_;
wire _5908_;
wire _5909_;
wire _5910_;
wire _5911_;
wire _5912_;
wire _5913_;
wire _5914_;
wire _5915_;
wire _5916_;
wire _5917_;
wire _5918_;
wire _5919_;
wire _5920_;
wire _5921_;
wire _5922_;
wire _5923_;
wire _5924_;
wire _5925_;
wire _5926_;
wire _5927_;
wire _5928_;
wire _5929_;
wire _5930_;
wire _5931_;
wire _5932_;
wire _5933_;
wire _5934_;
wire _5935_;
wire _5936_;
wire _5937_;
wire _5938_;
wire _5939_;
wire _5940_;
wire _5941_;
wire _5942_;
wire _5943_;
wire _5944_;
wire _5945_;
wire _5946_;
wire _5947_;
wire _5948_;
wire _5949_;
wire _5950_;
wire _5951_;
wire _5952_;
wire _5953_;
wire _5954_;
wire _5955_;
wire _5956_;
wire _5957_;
wire _5958_;
wire _5959_;
wire _5960_;
wire _5961_;
wire _5962_;
wire _5963_;
wire _5964_;
wire _5965_;
wire _5966_;
wire _5967_;
wire _5968_;
wire _5969_;
wire _5970_;
wire _5971_;
wire _5972_;
wire _5973_;
wire _5974_;
wire _5975_;
wire _5976_;
wire _5977_;
wire _5978_;
wire _5979_;
wire _5980_;
wire _5981_;
wire _5982_;
wire _5983_;
wire _5984_;
wire _5985_;
wire _5986_;
wire _5987_;
wire _5988_;
wire _5989_;
wire _5990_;
wire _5991_;
wire _5992_;
wire _5993_;
wire _5994_;
wire _5995_;
wire _5996_;
wire _5997_;
wire _5998_;
wire _5999_;
wire _6000_;
wire _6001_;
wire _6002_;
wire _6003_;
wire _6004_;
wire _6005_;
wire _6006_;
wire _6007_;
wire _6008_;
wire _6009_;
wire _6010_;
wire _6011_;
wire _6012_;
wire _6013_;
wire _6014_;
wire _6015_;
wire _6016_;
wire _6017_;
wire _6018_;
wire _6019_;
wire _6020_;
wire _6021_;
wire _6022_;
wire _6023_;
wire _6024_;
wire _6025_;
wire _6026_;
wire _6027_;
wire _6028_;
wire _6029_;
wire _6030_;
wire _6031_;
wire _6032_;
wire _6033_;
wire _6034_;
wire _6035_;
wire _6036_;
wire _6037_;
wire _6038_;
wire _6039_;
wire _6040_;
wire _6041_;
wire _6042_;
wire _6043_;
wire _6044_;
wire _6045_;
wire _6046_;
wire _6047_;
wire _6048_;
wire _6049_;
wire _6050_;
wire _6051_;
wire _6052_;
wire _6053_;
wire _6054_;
wire _6055_;
wire _6056_;
wire _6057_;
wire _6058_;
wire _6059_;
wire _6060_;
wire _6061_;
wire _6062_;
wire _6063_;
wire _6064_;
wire _6065_;
wire _6066_;
wire _6067_;
wire _6068_;
wire _6069_;
wire _6070_;
wire _6071_;
wire _6072_;
wire _6073_;
wire _6074_;
wire _6075_;
wire _6076_;
wire _6077_;
wire _6078_;
wire _6079_;
wire _6080_;
wire _6081_;
wire _6082_;
wire _6083_;
wire _6084_;
wire _6085_;
wire _6086_;
wire _6087_;
wire _6088_;
wire _6089_;
wire _6090_;
wire _6091_;
wire _6092_;
wire _6093_;
wire _6094_;
wire _6095_;
wire _6096_;
wire _6097_;
wire _6098_;
wire _6099_;
wire _6100_;
wire _6101_;
wire _6102_;
wire _6103_;
wire _6104_;
wire _6105_;
wire _6106_;
wire _6107_;
wire _6108_;
wire _6109_;
wire _6110_;
wire _6111_;
wire _6112_;
wire _6113_;
wire _6114_;
wire _6115_;
wire _6116_;
wire _6117_;
wire _6118_;
wire _6119_;
wire _6120_;
wire _6121_;
wire _6122_;
wire _6123_;
wire _6124_;
wire _6125_;
wire _6126_;
wire _6127_;
wire _6128_;
wire _6129_;
wire _6130_;
wire _6131_;
wire _6132_;
wire _6133_;
wire _6134_;
wire _6135_;
wire _6136_;
wire _6137_;
wire _6138_;
wire _6139_;
wire _6140_;
wire _6141_;
wire _6142_;
wire _6143_;
wire _6144_;
wire _6145_;
wire _6146_;
wire _6147_;
wire _6148_;
wire _6149_;
wire _6150_;
wire _6151_;
wire _6152_;
wire _6153_;
wire _6154_;
wire _6155_;
wire _6156_;
wire _6157_;
wire _6158_;
wire _6159_;
wire _6160_;
wire _6161_;
wire _6162_;
wire _6163_;
wire _6164_;
wire _6165_;
wire _6166_;
wire _6167_;
wire _6168_;
wire _6169_;
wire _6170_;
wire _6171_;
wire _6172_;
wire _6173_;
wire _6174_;
wire _6175_;
wire _6176_;
wire _6177_;
wire _6178_;
wire _6179_;
wire _6180_;
wire _6181_;
wire _6182_;
wire _6183_;
wire _6184_;
wire _6185_;
wire _6186_;
wire _6187_;
wire _6188_;
wire _6189_;
wire _6190_;
wire _6191_;
wire _6192_;
wire _6193_;
wire _6194_;
wire _6195_;
wire _6196_;
wire _6197_;
wire _6198_;
wire _6199_;
wire _6200_;
wire _6201_;
wire _6202_;
wire _6203_;
wire _6204_;
wire _6205_;
wire _6206_;
wire _6207_;
wire _6208_;
wire _6209_;
wire _6210_;
wire _6211_;
wire _6212_;
wire _6213_;
wire _6214_;
wire _6215_;
wire _6216_;
wire _6217_;
wire _6218_;
wire _6219_;
wire _6220_;
wire _6221_;
wire _6222_;
wire _6223_;
wire _6224_;
wire _6225_;
wire _6226_;
wire _6227_;
wire _6228_;
wire _6229_;
wire _6230_;
wire _6231_;
wire _6232_;
wire _6233_;
wire _6234_;
wire _6235_;
wire _6236_;
wire _6237_;
wire _6238_;
wire _6239_;
wire _6240_;
wire _6241_;
wire _6242_;
wire _6243_;
wire _6244_;
wire _6245_;
wire _6246_;
wire _6247_;
wire _6248_;
wire _6249_;
wire _6250_;
wire _6251_;
wire _6252_;
wire _6253_;
wire _6254_;
wire _6255_;
wire _6256_;
wire _6257_;
wire _6258_;
wire _6259_;
wire _6260_;
wire _6261_;
wire _6262_;
wire _6263_;
wire _6264_;
wire _6265_;
wire _6266_;
wire _6267_;
wire _6268_;
wire _6269_;
wire _6270_;
wire _6271_;
wire _6272_;
wire _6273_;
wire _6274_;
wire _6275_;
wire _6276_;
wire _6277_;
wire _6278_;
wire _6279_;
wire _6280_;
wire _6281_;
wire _6282_;
wire _6283_;
wire _6284_;
wire _6285_;
wire _6286_;
wire _6287_;
wire _6288_;
wire _6289_;
wire _6290_;
wire _6291_;
wire _6292_;
wire _6293_;
wire _6294_;
wire _6295_;
wire _6296_;
wire _6297_;
wire _6298_;
wire _6299_;
wire _6300_;
wire _6301_;
wire _6302_;
wire _6303_;
wire _6304_;
wire _6305_;
wire _6306_;
wire _6307_;
wire _6308_;
wire _6309_;
wire _6310_;
wire _6311_;
wire _6312_;
wire _6313_;
wire _6314_;
wire _6315_;
wire _6316_;
wire _6317_;
wire _6318_;
wire _6319_;
wire _6320_;
wire _6321_;
wire _6322_;
wire _6323_;
wire _6324_;
wire _6325_;
wire _6326_;
wire _6327_;
wire _6328_;
wire _6329_;
wire _6330_;
wire _6331_;
wire _6332_;
wire _6333_;
wire _6334_;
wire _6335_;
wire _6336_;
wire _6337_;
wire _6338_;
wire _6339_;
wire _6340_;
wire _6341_;
wire _6342_;
wire _6343_;
wire _6344_;
wire _6345_;
wire _6346_;
wire _6347_;
wire _6348_;
wire _6349_;
wire _6350_;
wire _6351_;
wire _6352_;
wire _6353_;
wire _6354_;
wire _6355_;
wire _6356_;
wire _6357_;
wire _6358_;
wire _6359_;
wire _6360_;
wire _6361_;
wire _6362_;
wire _6363_;
wire _6364_;
wire _6365_;
wire _6366_;
wire _6367_;
wire _6368_;
wire _6369_;
wire _6370_;
wire _6371_;
wire _6372_;
wire _6373_;
wire _6374_;
wire _6375_;
wire _6376_;
wire _6377_;
wire _6378_;
wire _6379_;
wire _6380_;
wire _6381_;
wire _6382_;
wire _6383_;
wire _6384_;
wire _6385_;
wire _6386_;
wire _6387_;
wire _6388_;
wire _6389_;
wire _6390_;
wire _6391_;
wire _6392_;
wire _6393_;
wire _6394_;
wire _6395_;
wire _6396_;
wire _6397_;
wire _6398_;
wire _6399_;
wire _6400_;
wire _6401_;
wire _6402_;
wire _6403_;
wire _6404_;
wire _6405_;
wire _6406_;
wire _6407_;
wire _6408_;
wire _6409_;
wire _6410_;
wire _6411_;
wire _6412_;
wire _6413_;
wire _6414_;
wire _6415_;
wire _6416_;
wire _6417_;
wire _6418_;
wire _6419_;
wire _6420_;
wire _6421_;
wire _6422_;
wire _6423_;
wire _6424_;
wire _6425_;
wire _6426_;
wire _6427_;
wire _6428_;
wire _6429_;
wire _6430_;
wire _6431_;
wire _6432_;
wire _6433_;
wire _6434_;
wire _6435_;
wire _6436_;
wire _6437_;
wire _6438_;
wire _6439_;
wire _6440_;
wire _6441_;
wire _6442_;
wire _6443_;
wire _6444_;
wire _6445_;
wire _6446_;
wire _6447_;
wire _6448_;
wire _6449_;
wire _6450_;
wire _6451_;
wire _6452_;
wire _6453_;
wire _6454_;
wire _6455_;
wire _6456_;
wire _6457_;
wire _6458_;
wire _6459_;
wire _6460_;
wire _6461_;
wire _6462_;
wire _6463_;
wire _6464_;
wire _6465_;
wire _6466_;
wire _6467_;
wire _6468_;
wire _6469_;
wire _6470_;
wire _6471_;
wire _6472_;
wire _6473_;
wire _6474_;
wire _6475_;
wire _6476_;
wire _6477_;
wire _6478_;
wire _6479_;
wire _6480_;
wire _6481_;
wire _6482_;
wire _6483_;
wire _6484_;
wire _6485_;
wire _6486_;
wire _6487_;
wire _6488_;
wire _6489_;
wire _6490_;
wire _6491_;
wire _6492_;
wire _6493_;
wire _6494_;
wire _6495_;
wire _6496_;
wire _6497_;
wire _6498_;
wire _6499_;
wire _6500_;
wire _6501_;
wire _6502_;
wire _6503_;
wire _6504_;
wire _6505_;
wire _6506_;
wire _6507_;
wire _6508_;
wire _6509_;
wire _6510_;
wire _6511_;
wire _6512_;
wire _6513_;
wire _6514_;
wire _6515_;
wire _6516_;
wire _6517_;
wire _6518_;
wire _6519_;
wire _6520_;
wire _6521_;
wire _6522_;
wire _6523_;
wire _6524_;
wire _6525_;
wire _6526_;
wire _6527_;
wire _6528_;
wire _6529_;
wire _6530_;
wire _6531_;
wire _6532_;
wire _6533_;
wire _6534_;
wire _6535_;
wire _6536_;
wire _6537_;
wire _6538_;
wire _6539_;
wire _6540_;
wire _6541_;
wire _6542_;
wire _6543_;
wire _6544_;
wire _6545_;
wire _6546_;
wire _6547_;
wire _6548_;
wire _6549_;
wire _6550_;
wire _6551_;
wire _6552_;
wire _6553_;
wire _6554_;
wire _6555_;
wire _6556_;
wire _6557_;
wire _6558_;
wire _6559_;
wire _6560_;
wire _6561_;
wire _6562_;
wire _6563_;
wire _6564_;
wire _6565_;
wire _6566_;
wire _6567_;
wire _6568_;
wire _6569_;
wire _6570_;
wire _6571_;
wire _6572_;
wire _6573_;
wire _6574_;
wire _6575_;
wire _6576_;
wire _6577_;
wire _6578_;
wire _6579_;
wire _6580_;
wire _6581_;
wire _6582_;
wire _6583_;
wire _6584_;
wire _6585_;
wire _6586_;
wire _6587_;
wire _6588_;
wire _6589_;
wire _6590_;
wire _6591_;
wire _6592_;
wire _6593_;
wire _6594_;
wire _6595_;
wire _6596_;
wire _6597_;
wire _6598_;
wire _6599_;
wire _6600_;
wire _6601_;
wire _6602_;
wire _6603_;
wire _6604_;
wire _6605_;
wire _6606_;
wire _6607_;
wire _6608_;
wire _6609_;
wire _6610_;
wire _6611_;
wire _6612_;
wire _6613_;
wire _6614_;
wire _6615_;
wire _6616_;
wire _6617_;
wire _6618_;
wire _6619_;
wire _6620_;
wire _6621_;
wire _6622_;
wire _6623_;
wire _6624_;
wire _6625_;
wire _6626_;
wire _6627_;
wire _6628_;
wire _6629_;
wire _6630_;
wire _6631_;
wire _6632_;
wire _6633_;
wire _6634_;
wire _6635_;
wire _6636_;
wire _6637_;
wire _6638_;
wire _6639_;
wire _6640_;
wire _6641_;
wire _6642_;
wire _6643_;
wire _6644_;
wire _6645_;
wire _6646_;
wire _6647_;
wire _6648_;
wire _6649_;
wire _6650_;
wire _6651_;
wire _6652_;
wire _6653_;
wire _6654_;
wire _6655_;
wire _6656_;
wire _6657_;
wire _6658_;
wire _6659_;
wire _6660_;
wire _6661_;
wire _6662_;
wire _6663_;
wire _6664_;
wire _6665_;
wire _6666_;
wire _6667_;
wire _6668_;
wire _6669_;
wire _6670_;
wire _6671_;
wire _6672_;
wire _6673_;
wire _6674_;
wire _6675_;
wire _6676_;
wire _6677_;
wire _6678_;
wire _6679_;
wire _6680_;
wire _6681_;
wire _6682_;
wire _6683_;
wire _6684_;
wire _6685_;
wire _6686_;
wire _6687_;
wire _6688_;
wire _6689_;
wire _6690_;
wire _6691_;
wire _6692_;
wire _6693_;
wire _6694_;
wire _6695_;
wire _6696_;
wire _6697_;
wire _6698_;
wire _6699_;
wire _6700_;
wire _6701_;
wire _6702_;
wire _6703_;
wire _6704_;
wire _6705_;
wire _6706_;
wire _6707_;
wire _6708_;
wire _6709_;
wire _6710_;
wire _6711_;
wire _6712_;
wire _6713_;
wire _6714_;
wire _6715_;
wire _6716_;
wire _6717_;
wire _6718_;
wire _6719_;
wire _6720_;
wire _6721_;
wire _6722_;
wire _6723_;
wire _6724_;
wire _6725_;
wire _6726_;
wire _6727_;
wire _6728_;
wire _6729_;
wire _6730_;
wire _6731_;
wire _6732_;
wire _6733_;
wire _6734_;
wire _6735_;
wire _6736_;
wire _6737_;
wire _6738_;
wire _6739_;
wire _6740_;
wire _6741_;
wire _6742_;
wire _6743_;
wire _6744_;
wire _6745_;
wire _6746_;
wire _6747_;
wire _6748_;
wire _6749_;
wire _6750_;
wire _6751_;
wire _6752_;
wire _6753_;
wire _6754_;
wire _6755_;
wire _6756_;
wire _6757_;
wire _6758_;
wire _6759_;
wire _6760_;
wire _6761_;
wire _6762_;
wire _6763_;
wire _6764_;
wire _6765_;
wire _6766_;
wire _6767_;
wire _6768_;
wire _6769_;
wire _6770_;
wire _6771_;
wire _6772_;
wire _6773_;
wire _6774_;
wire _6775_;
wire _6776_;
wire _6777_;
wire _6778_;
wire _6779_;
wire _6780_;
wire _6781_;
wire _6782_;
wire _6783_;
wire _6784_;
wire _6785_;
wire _6786_;
wire _6787_;
wire _6788_;
wire _6789_;
wire _6790_;
wire _6791_;
wire _6792_;
wire _6793_;
wire _6794_;
wire _6795_;
wire _6796_;
wire _6797_;
wire _6798_;
wire _6799_;
wire _6800_;
wire _6801_;
wire _6802_;
wire _6803_;
wire _6804_;
wire _6805_;
wire _6806_;
wire _6807_;
wire _6808_;
wire _6809_;
wire _6810_;
wire _6811_;
wire _6812_;
wire _6813_;
wire _6814_;
wire _6815_;
wire _6816_;
wire _6817_;
wire _6818_;
wire _6819_;
wire _6820_;
wire _6821_;
wire _6822_;
wire _6823_;
wire _6824_;
wire _6825_;
wire _6826_;
wire _6827_;
wire _6828_;
wire _6829_;
wire _6830_;
wire _6831_;
wire _6832_;
wire _6833_;
wire _6834_;
wire _6835_;
wire _6836_;
wire _6837_;
wire _6838_;
wire _6839_;
wire _6840_;
wire _6841_;
wire _6842_;
wire _6843_;
wire _6844_;
wire _6845_;
wire _6846_;
wire _6847_;
wire _6848_;
wire _6849_;
wire _6850_;
wire _6851_;
wire _6852_;
wire _6853_;
wire _6854_;
wire _6855_;
wire _6856_;
wire _6857_;
wire _6858_;
wire _6859_;
wire _6860_;
wire _6861_;
wire _6862_;
wire _6863_;
wire _6864_;
wire _6865_;
wire _6866_;
wire _6867_;
wire _6868_;
wire _6869_;
wire _6870_;
wire _6871_;
wire _6872_;
wire _6873_;
wire _6874_;
wire _6875_;
wire _6876_;
wire _6877_;
wire _6878_;
wire _6879_;
wire _6880_;
wire _6881_;
wire _6882_;
wire _6883_;
wire _6884_;
wire _6885_;
wire _6886_;
wire _6887_;
wire _6888_;
wire _6889_;
wire _6890_;
wire _6891_;
wire _6892_;
wire _6893_;
wire _6894_;
wire _6895_;
wire _6896_;
wire _6897_;
wire _6898_;
wire _6899_;
wire _6900_;
wire _6901_;
wire _6902_;
wire _6903_;
wire _6904_;
wire _6905_;
wire _6906_;
wire _6907_;
wire _6908_;
wire _6909_;
wire _6910_;
wire _6911_;
wire _6912_;
wire _6913_;
wire _6914_;
wire _6915_;
wire _6916_;
wire _6917_;
wire _6918_;
wire _6919_;
wire _6920_;
wire _6921_;
wire _6922_;
wire _6923_;
wire _6924_;
wire _6925_;
wire _6926_;
wire _6927_;
wire _6928_;
wire _6929_;
wire _6930_;
wire _6931_;
wire _6932_;
wire _6933_;
wire _6934_;
wire _6935_;
wire _6936_;
wire _6937_;
wire _6938_;
wire _6939_;
wire _6940_;
wire _6941_;
wire _6942_;
wire _6943_;
wire _6944_;
wire _6945_;
wire _6946_;
wire _6947_;
wire _6948_;
wire _6949_;
wire _6950_;
wire _6951_;
wire _6952_;
wire _6953_;
wire _6954_;
wire _6955_;
wire _6956_;
wire _6957_;
wire _6958_;
wire _6959_;
wire _6960_;
wire _6961_;
wire _6962_;
wire _6963_;
wire _6964_;
wire _6965_;
wire _6966_;
wire _6967_;
wire _6968_;
wire _6969_;
wire _6970_;
wire _6971_;
wire _6972_;
wire _6973_;
wire _6974_;
wire _6975_;
wire _6976_;
wire _6977_;
wire _6978_;
wire _6979_;
wire _6980_;
wire _6981_;
wire _6982_;
wire _6983_;
wire _6984_;
wire _6985_;
wire _6986_;
wire _6987_;
wire _6988_;
wire _6989_;
wire _6990_;
wire _6991_;
wire _6992_;
wire _6993_;
wire _6994_;
wire _6995_;
wire _6996_;
wire _6997_;
wire _6998_;
wire _6999_;
wire _7000_;
wire _7001_;
wire _7002_;
wire _7003_;
wire _7004_;
wire _7005_;
wire _7006_;
wire _7007_;
wire _7008_;
wire _7009_;
wire _7010_;
wire _7011_;
wire _7012_;
wire _7013_;
wire _7014_;
wire _7015_;
wire _7016_;
wire _7017_;
wire _7018_;
wire _7019_;
wire _7020_;
wire _7021_;
wire _7022_;
wire _7023_;
wire _7024_;
wire _7025_;
wire _7026_;
wire _7027_;
wire _7028_;
wire _7029_;
wire _7030_;
wire _7031_;
wire _7032_;
wire _7033_;
wire _7034_;
wire _7035_;
wire _7036_;
wire _7037_;
wire _7038_;
wire _7039_;
wire _7040_;
wire _7041_;
wire _7042_;
wire _7043_;
wire _7044_;
wire _7045_;
wire _7046_;
wire _7047_;
wire _7048_;
wire _7049_;
wire _7050_;
wire _7051_;
wire _7052_;
wire _7053_;
wire _7054_;
wire _7055_;
wire _7056_;
wire _7057_;
wire _7058_;
wire _7059_;
wire _7060_;
wire _7061_;
wire _7062_;
wire _7063_;
wire _7064_;
wire _7065_;
wire _7066_;
wire _7067_;
wire _7068_;
wire _7069_;
wire _7070_;
wire _7071_;
wire _7072_;
wire _7073_;
wire _7074_;
wire _7075_;
wire _7076_;
wire _7077_;
wire _7078_;
wire _7079_;
wire _7080_;
wire _7081_;
wire _7082_;
wire _7083_;
wire _7084_;
wire _7085_;
wire _7086_;
wire _7087_;
wire _7088_;
wire _7089_;
wire _7090_;
wire _7091_;
wire _7092_;
wire _7093_;
wire _7094_;
wire _7095_;
wire _7096_;
wire _7097_;
wire _7098_;
wire _7099_;
wire _7100_;
wire _7101_;
wire _7102_;
wire _7103_;
wire _7104_;
wire _7105_;
wire _7106_;
wire _7107_;
wire _7108_;
wire _7109_;
wire _7110_;
wire _7111_;
wire _7112_;
wire _7113_;
wire _7114_;
wire _7115_;
wire _7116_;
wire _7117_;
wire _7118_;
wire _7119_;
wire _7120_;
wire _7121_;
wire _7122_;
wire _7123_;
wire _7124_;
wire _7125_;
wire _7126_;
wire _7127_;
wire _7128_;
wire _7129_;
wire _7130_;
wire _7131_;
wire _7132_;
wire _7133_;
wire _7134_;
wire _7135_;
wire _7136_;
wire _7137_;
wire _7138_;
wire _7139_;
wire _7140_;
wire _7141_;
wire _7142_;
wire _7143_;
wire _7144_;
wire _7145_;
wire _7146_;
wire _7147_;
wire _7148_;
wire _7149_;
wire _7150_;
wire _7151_;
wire _7152_;
wire _7153_;
wire _7154_;
wire _7155_;
wire _7156_;
wire _7157_;
wire _7158_;
wire _7159_;
wire _7160_;
wire _7161_;
wire _7162_;
wire _7163_;
wire _7164_;
wire _7165_;
wire _7166_;
wire _7167_;
wire _7168_;
wire _7169_;
wire _7170_;
wire _7171_;
wire _7172_;
wire _7173_;
wire _7174_;
wire _7175_;
wire _7176_;
wire _7177_;
wire _7178_;
wire _7179_;
wire _7180_;
wire _7181_;
wire _7182_;
wire _7183_;
wire _7184_;
wire _7185_;
wire _7186_;
wire _7187_;
wire _7188_;
wire _7189_;
wire _7190_;
wire _7191_;
wire _7192_;
wire _7193_;
wire _7194_;
wire _7195_;
wire _7196_;
wire _7197_;
wire _7198_;
wire _7199_;
wire _7200_;
wire _7201_;
wire _7202_;
wire _7203_;
wire _7204_;
wire _7205_;
wire _7206_;
wire _7207_;
wire _7208_;
wire _7209_;
wire _7210_;
wire _7211_;
wire _7212_;
wire _7213_;
wire _7214_;
wire _7215_;
wire _7216_;
wire _7217_;
wire _7218_;
wire _7219_;
wire _7220_;
wire _7221_;
wire _7222_;
wire _7223_;
wire _7224_;
wire _7225_;
wire _7226_;
wire _7227_;
wire _7228_;
wire _7229_;
wire _7230_;
wire _7231_;
wire _7232_;
wire _7233_;
wire _7234_;
wire _7235_;
wire _7236_;
wire _7237_;
wire _7238_;
wire _7239_;
wire _7240_;
wire _7241_;
wire _7242_;
wire _7243_;
wire _7244_;
wire _7245_;
wire _7246_;
wire _7247_;
wire _7248_;
wire _7249_;
wire _7250_;
wire _7251_;
wire _7252_;
wire _7253_;
wire _7254_;
wire _7255_;
wire _7256_;
wire _7257_;
wire _7258_;
wire _7259_;
wire _7260_;
wire _7261_;
wire _7262_;
wire _7263_;
wire _7264_;
wire _7265_;
wire _7266_;
wire _7267_;
wire _7268_;
wire _7269_;
wire _7270_;
wire _7271_;
wire _7272_;
wire _7273_;
wire _7274_;
wire _7275_;
wire _7276_;
wire _7277_;
wire _7278_;
wire _7279_;
wire _7280_;
wire _7281_;
wire _7282_;
wire _7283_;
wire _7284_;
wire _7285_;
wire _7286_;
wire _7287_;
wire _7288_;
wire _7289_;
wire _7290_;
wire _7291_;
wire _7292_;
wire _7293_;
wire _7294_;
wire _7295_;
wire _7296_;
wire _7297_;
wire _7298_;
wire _7299_;
wire _7300_;
wire _7301_;
wire _7302_;
wire _7303_;
wire _7304_;
wire _7305_;
wire _7306_;
wire _7307_;
wire _7308_;
wire _7309_;
wire _7310_;
wire _7311_;
wire _7312_;
wire _7313_;
wire _7314_;
wire _7315_;
wire _7316_;
wire _7317_;
wire _7318_;
wire _7319_;
wire _7320_;
wire _7321_;
wire _7322_;
wire _7323_;
wire _7324_;
wire _7325_;
wire _7326_;
wire _7327_;
wire _7328_;
wire _7329_;
wire _7330_;
wire _7331_;
wire _7332_;
wire _7333_;
wire _7334_;
wire _7335_;
wire _7336_;
wire _7337_;
wire _7338_;
wire _7339_;
wire _7340_;
wire _7341_;
wire _7342_;
wire _7343_;
wire _7344_;
wire _7345_;
wire _7346_;
wire _7347_;
wire _7348_;
wire _7349_;
wire _7350_;
wire _7351_;
wire _7352_;
wire _7353_;
wire _7354_;
wire _7355_;
wire _7356_;
wire _7357_;
wire _7358_;
wire _7359_;
wire _7360_;
wire _7361_;
wire _7362_;
wire _7363_;
wire _7364_;
wire _7365_;
wire _7366_;
wire _7367_;
wire _7368_;
wire _7369_;
wire _7370_;
wire _7371_;
wire _7372_;
wire _7373_;
wire _7374_;
wire _7375_;
wire _7376_;
wire _7377_;
wire _7378_;
wire _7379_;
wire _7380_;
wire _7381_;
wire _7382_;
wire _7383_;
wire _7384_;
wire _7385_;
wire _7386_;
wire _7387_;
wire _7388_;
wire _7389_;
wire _7390_;
wire _7391_;
wire _7392_;
wire _7393_;
wire _7394_;
wire _7395_;
wire _7396_;
wire _7397_;
wire _7398_;
wire _7399_;
wire _7400_;
wire _7401_;
wire _7402_;
wire _7403_;
wire _7404_;
wire _7405_;
wire _7406_;
wire _7407_;
wire _7408_;
wire _7409_;
wire _7410_;
wire _7411_;
wire _7412_;
wire _7413_;
wire _7414_;
wire _7415_;
wire _7416_;
wire _7417_;
wire _7418_;
wire _7419_;
wire _7420_;
wire _7421_;
wire _7422_;
wire _7423_;
wire _7424_;
wire _7425_;
wire _7426_;
wire _7427_;
wire _7428_;
wire _7429_;
wire _7430_;
wire _7431_;
wire _7432_;
wire _7433_;
wire _7434_;
wire _7435_;
wire _7436_;
wire _7437_;
wire _7438_;
wire _7439_;
wire _7440_;
wire _7441_;
wire _7442_;
wire _7443_;
wire _7444_;
wire _7445_;
wire _7446_;
wire _7447_;
wire _7448_;
wire _7449_;
wire _7450_;
wire _7451_;
wire _7452_;
wire _7453_;
wire _7454_;
wire _7455_;
wire _7456_;
wire _7457_;
wire _7458_;
wire _7459_;
wire _7460_;
wire _7461_;
wire _7462_;
wire _7463_;
wire _7464_;
wire _7465_;
wire _7466_;
wire _7467_;
wire _7468_;
wire _7469_;
wire _7470_;
wire _7471_;
wire _7472_;
wire _7473_;
wire _7474_;
wire _7475_;
wire _7476_;
wire _7477_;
wire _7478_;
wire _7479_;
wire _7480_;
wire _7481_;
wire _7482_;
wire _7483_;
wire _7484_;
wire _7485_;
wire _7486_;
wire _7487_;
wire _7488_;
wire _7489_;
wire _7490_;
wire _7491_;
wire _7492_;
wire _7493_;
wire _7494_;
wire _7495_;
wire _7496_;
wire _7497_;
wire _7498_;
wire _7499_;
wire _7500_;
wire _7501_;
wire _7502_;
wire _7503_;
wire _7504_;
wire _7505_;
wire _7506_;
wire _7507_;
wire _7508_;
wire _7509_;
wire _7510_;
wire _7511_;
wire _7512_;
wire _7513_;
wire _7514_;
wire _7515_;
wire _7516_;
wire _7517_;
wire _7518_;
wire _7519_;
wire _7520_;
wire _7521_;
wire _7522_;
wire _7523_;
wire _7524_;
wire _7525_;
wire _7526_;
wire _7527_;
wire _7528_;
wire _7529_;
wire _7530_;
wire _7531_;
wire _7532_;
wire _7533_;
wire _7534_;
wire _7535_;
wire _7536_;
wire _7537_;
wire _7538_;
wire _7539_;
wire _7540_;
wire _7541_;
wire _7542_;
wire _7543_;
wire _7544_;
wire _7545_;
wire _7546_;
wire _7547_;
wire _7548_;
wire _7549_;
wire _7550_;
wire _7551_;
wire _7552_;
wire _7553_;
wire _7554_;
wire _7555_;
wire _7556_;
wire _7557_;
wire _7558_;
wire _7559_;
wire _7560_;
wire _7561_;
wire _7562_;
wire _7563_;
wire _7564_;
wire _7565_;
wire _7566_;
wire _7567_;
wire _7568_;
wire _7569_;
wire _7570_;
wire _7571_;
wire _7572_;
wire _7573_;
wire _7574_;
wire _7575_;
wire _7576_;
wire _7577_;
wire _7578_;
wire _7579_;
wire _7580_;
wire _7581_;
wire _7582_;
wire _7583_;
wire _7584_;
wire _7585_;
wire _7586_;
wire _7587_;
wire _7588_;
wire _7589_;
wire _7590_;
wire _7591_;
wire _7592_;
wire _7593_;
wire _7594_;
wire _7595_;
wire _7596_;
wire _7597_;
wire _7598_;
wire _7599_;
wire _7600_;
wire _7601_;
wire _7602_;
wire _7603_;
wire _7604_;
wire _7605_;
wire _7606_;
wire _7607_;
wire _7608_;
wire _7609_;
wire _7610_;
wire _7611_;
wire _7612_;
wire _7613_;
wire _7614_;
wire _7615_;
wire _7616_;
wire _7617_;
wire _7618_;
wire _7619_;
wire _7620_;
wire _7621_;
wire _7622_;
wire _7623_;
wire _7624_;
wire _7625_;
wire _7626_;
wire _7627_;
wire _7628_;
wire _7629_;
wire _7630_;
wire _7631_;
wire _7632_;
wire _7633_;
wire _7634_;
wire _7635_;
wire _7636_;
wire _7637_;
wire _7638_;
wire _7639_;
wire _7640_;
wire _7641_;
wire _7642_;
wire _7643_;
wire _7644_;
wire _7645_;
wire _7646_;
wire _7647_;
wire _7648_;
wire _7649_;
wire _7650_;
wire _7651_;
wire _7652_;
wire _7653_;
wire _7654_;
wire _7655_;
wire _7656_;
wire _7657_;
wire _7658_;
wire _7659_;
wire _7660_;
wire _7661_;
wire _7662_;
wire _7663_;
wire _7664_;
wire _7665_;
wire _7666_;
wire _7667_;
wire _7668_;
wire _7669_;
wire _7670_;
wire _7671_;
wire _7672_;
wire _7673_;
wire _7674_;
wire _7675_;
wire _7676_;
wire _7677_;
wire _7678_;
wire _7679_;
wire _7680_;
wire _7681_;
wire _7682_;
wire _7683_;
wire _7684_;
wire _7685_;
wire _7686_;
wire _7687_;
wire _7688_;
wire _7689_;
wire _7690_;
wire _7691_;
wire _7692_;
wire _7693_;
wire _7694_;
wire _7695_;
wire _7696_;
wire _7697_;
wire _7698_;
wire _7699_;
wire _7700_;
wire _7701_;
wire _7702_;
wire _7703_;
wire _7704_;
wire _7705_;
wire _7706_;
wire _7707_;
wire _7708_;
wire _7709_;
wire _7710_;
wire _7711_;
wire _7712_;
wire _7713_;
wire _7714_;
wire _7715_;
wire _7716_;
wire _7717_;
wire _7718_;
wire _7719_;
wire _7720_;
wire _7721_;
wire _7722_;
wire _7723_;
wire _7724_;
wire _7725_;
wire _7726_;
wire _7727_;
wire _7728_;
wire _7729_;
wire _7730_;
wire _7731_;
wire _7732_;
wire _7733_;
wire _7734_;
wire _7735_;
wire _7736_;
wire _7737_;
wire _7738_;
wire _7739_;
wire _7740_;
wire _7741_;
wire _7742_;
wire _7743_;
wire _7744_;
wire _7745_;
wire _7746_;
wire _7747_;
wire _7748_;
wire _7749_;
wire _7750_;
wire _7751_;
wire _7752_;
wire _7753_;
wire _7754_;
wire _7755_;
wire _7756_;
wire _7757_;
wire _7758_;
wire _7759_;
wire _7760_;
wire _7761_;
wire _7762_;
wire _7763_;
wire _7764_;
wire _7765_;
wire _7766_;
wire _7767_;
wire _7768_;
wire _7769_;
wire _7770_;
wire _7771_;
wire _7772_;
wire _7773_;
wire _7774_;
wire _7775_;
wire _7776_;
wire _7777_;
wire _7778_;
wire _7779_;
wire _7780_;
wire _7781_;
wire _7782_;
wire _7783_;
wire _7784_;
wire _7785_;
wire _7786_;
wire _7787_;
wire _7788_;
wire _7789_;
wire _7790_;
wire _7791_;
wire _7792_;
wire _7793_;
wire _7794_;
wire _7795_;
wire _7796_;
wire _7797_;
wire _7798_;
wire _7799_;
wire _7800_;
wire _7801_;
wire _7802_;
wire _7803_;
wire _7804_;
wire _7805_;
wire _7806_;
wire _7807_;
wire _7808_;
wire _7809_;
wire _7810_;
wire _7811_;
wire _7812_;
wire _7813_;
wire _7814_;
wire _7815_;
wire _7816_;
wire _7817_;
wire _7818_;
wire _7819_;
wire _7820_;
wire _7821_;
wire _7822_;
wire _7823_;
wire _7824_;
wire _7825_;
wire _7826_;
wire _7827_;
wire _7828_;
wire _7829_;
wire _7830_;
wire _7831_;
wire _7832_;
wire _7833_;
wire _7834_;
wire _7835_;
wire _7836_;
wire _7837_;
wire _7838_;
wire _7839_;
wire _7840_;
wire _7841_;
wire _7842_;
wire _7843_;
wire _7844_;
wire _7845_;
wire _7846_;
wire _7847_;
wire _7848_;
wire _7849_;
wire _7850_;
wire _7851_;
wire _7852_;
wire _7853_;
wire _7854_;
wire _7855_;
wire _7856_;
wire _7857_;
wire _7858_;
wire _7859_;
wire _7860_;
wire _7861_;
wire _7862_;
wire _7863_;
wire _7864_;
wire _7865_;
wire _7866_;
wire _7867_;
wire _7868_;
wire _7869_;
wire _7870_;
wire _7871_;
wire _7872_;
wire _7873_;
wire _7874_;
wire _7875_;
wire _7876_;
wire _7877_;
wire _7878_;
wire _7879_;
wire _7880_;
wire _7881_;
wire _7882_;
wire _7883_;
wire _7884_;
wire _7885_;
wire _7886_;
wire _7887_;
wire _7888_;
wire _7889_;
wire _7890_;
wire _7891_;
wire _7892_;
wire _7893_;
wire _7894_;
wire _7895_;
wire _7896_;
wire _7897_;
wire _7898_;
wire _7899_;
wire _7900_;
wire _7901_;
wire _7902_;
wire _7903_;
wire _7904_;
wire _7905_;
wire _7906_;
wire _7907_;
wire _7908_;
wire _7909_;
wire _7910_;
wire _7911_;
wire _7912_;
wire _7913_;
wire _7914_;
wire _7915_;
wire _7916_;
wire _7917_;
wire _7918_;
wire _7919_;
wire _7920_;
wire _7921_;
wire _7922_;
wire _7923_;
wire _7924_;
wire _7925_;
wire _7926_;
wire _7927_;
wire _7928_;
wire _7929_;
wire _7930_;
wire _7931_;
wire _7932_;
wire _7933_;
wire _7934_;
wire _7935_;
wire _7936_;
wire _7937_;
wire _7938_;
wire _7939_;
wire _7940_;
wire _7941_;
wire _7942_;
wire _7943_;
wire _7944_;
wire _7945_;
wire _7946_;
wire _7947_;
wire _7948_;
wire _7949_;
wire _7950_;
wire _7951_;
wire _7952_;
wire _7953_;
wire _7954_;
wire _7955_;
wire _7956_;
wire _7957_;
wire _7958_;
wire _7959_;
wire _7960_;
wire _7961_;
wire _7962_;
wire _7963_;
wire _7964_;
wire _7965_;
wire _7966_;
wire _7967_;
wire _7968_;
wire _7969_;
wire _7970_;
wire _7971_;
wire _7972_;
wire _7973_;
wire _7974_;
wire _7975_;
wire _7976_;
wire _7977_;
wire _7978_;
wire _7979_;
wire _7980_;
wire _7981_;
wire _7982_;
wire _7983_;
wire _7984_;
wire _7985_;
wire _7986_;
wire _7987_;
wire _7988_;
wire _7989_;
wire _7990_;
wire _7991_;
wire _7992_;
wire _7993_;
wire _7994_;
wire _7995_;
wire _7996_;
wire _7997_;
wire _7998_;
wire _7999_;
wire _8000_;
wire _8001_;
wire _8002_;
wire _8003_;
wire _8004_;
wire _8005_;
wire _8006_;
wire _8007_;
wire _8008_;
wire _8009_;
wire _8010_;
wire _8011_;
wire _8012_;
wire _8013_;
wire _8014_;
wire _8015_;
wire _8016_;
wire _8017_;
wire _8018_;
wire _8019_;
wire _8020_;
wire _8021_;
wire _8022_;
wire _8023_;
wire _8024_;
wire _8025_;
wire _8026_;
wire _8027_;
wire _8028_;
wire _8029_;
wire _8030_;
wire _8031_;
wire _8032_;
wire _8033_;
wire _8034_;
wire _8035_;
wire _8036_;
wire _8037_;
wire _8038_;
wire _8039_;
wire _8040_;
wire _8041_;
wire _8042_;
wire _8043_;
wire _8044_;
wire _8045_;
wire _8046_;
wire _8047_;
wire _8048_;
wire _8049_;
wire _8050_;
wire _8051_;
wire _8052_;
wire _8053_;
wire _8054_;
wire _8055_;
wire _8056_;
wire _8057_;
wire _8058_;
wire _8059_;
wire _8060_;
wire _8061_;
wire _8062_;
wire _8063_;
wire _8064_;
wire _8065_;
wire _8066_;
wire _8067_;
wire _8068_;
wire _8069_;
wire _8070_;
wire _8071_;
wire _8072_;
wire _8073_;
wire _8074_;
wire _8075_;
wire _8076_;
wire _8077_;
wire _8078_;
wire _8079_;
wire _8080_;
wire _8081_;
wire _8082_;
wire _8083_;
wire _8084_;
wire _8085_;
wire _8086_;
wire _8087_;
wire _8088_;
wire _8089_;
wire _8090_;
wire _8091_;
wire _8092_;
wire _8093_;
wire _8094_;
wire _8095_;
wire _8096_;
wire _8097_;
wire _8098_;
wire _8099_;
wire _8100_;
wire _8101_;
wire _8102_;
wire _8103_;
wire _8104_;
wire _8105_;
wire _8106_;
wire _8107_;
wire _8108_;
wire _8109_;
wire _8110_;
wire _8111_;
wire _8112_;
wire _8113_;
wire _8114_;
wire _8115_;
wire _8116_;
wire _8117_;
wire _8118_;
wire _8119_;
wire _8120_;
wire _8121_;
wire _8122_;
wire _8123_;
wire _8124_;
wire _8125_;
wire _8126_;
wire _8127_;
wire _8128_;
wire _8129_;
wire _8130_;
wire _8131_;
wire _8132_;
wire _8133_;
wire _8134_;
wire _8135_;
wire _8136_;
wire _8137_;
wire _8138_;
wire _8139_;
wire _8140_;
wire _8141_;
wire _8142_;
wire _8143_;
wire _8144_;
wire _8145_;
wire _8146_;
wire _8147_;
wire _8148_;
wire _8149_;
wire _8150_;
wire _8151_;
wire _8152_;
wire _8153_;
wire _8154_;
wire _8155_;
wire _8156_;
wire _8157_;
wire _8158_;
wire _8159_;
wire _8160_;
wire _8161_;
wire _8162_;
wire _8163_;
wire _8164_;
wire _8165_;
wire _8166_;
wire _8167_;
wire _8168_;
wire _8169_;
wire _8170_;
wire _8171_;
wire _8172_;
wire _8173_;
wire _8174_;
wire _8175_;
wire _8176_;
wire _8177_;
wire _8178_;
wire _8179_;
wire _8180_;
wire _8181_;
wire _8182_;
wire _8183_;
wire _8184_;
wire _8185_;
wire _8186_;
wire _8187_;
wire _8188_;
wire _8189_;
wire _8190_;
wire _8191_;
wire _8192_;
wire _8193_;
wire _8194_;
wire _8195_;
wire _8196_;
wire _8197_;
wire _8198_;
wire _8199_;
wire _8200_;
wire _8201_;
wire _8202_;
wire _8203_;
wire _8204_;
wire _8205_;
wire _8206_;
wire _8207_;
wire _8208_;
wire _8209_;
wire _8210_;
wire _8211_;
wire _8212_;
wire _8213_;
wire _8214_;
wire _8215_;
wire _8216_;
wire _8217_;
wire _8218_;
wire _8219_;
wire _8220_;
wire _8221_;
wire _8222_;
wire _8223_;
wire _8224_;
wire _8225_;
wire _8226_;
wire _8227_;
wire _8228_;
wire _8229_;
wire _8230_;
wire _8231_;
wire _8232_;
wire _8233_;
wire _8234_;
wire _8235_;
wire _8236_;
wire _8237_;
wire _8238_;
wire _8239_;
wire _8240_;
wire _8241_;
wire _8242_;
wire _8243_;
wire _8244_;
wire _8245_;
wire _8246_;
wire _8247_;
wire _8248_;
wire _8249_;
wire _8250_;
wire _8251_;
wire _8252_;
wire _8253_;
wire _8254_;
wire _8255_;
wire _8256_;
wire _8257_;
wire _8258_;
wire _8259_;
wire _8260_;
wire _8261_;
wire _8262_;
wire _8263_;
wire _8264_;
wire _8265_;
wire _8266_;
wire _8267_;
wire _8268_;
wire _8269_;
wire _8270_;
wire _8271_;
wire _8272_;
wire _8273_;
wire _8274_;
wire _8275_;
wire _8276_;
wire _8277_;
wire _8278_;
wire _8279_;
wire _8280_;
wire _8281_;
wire _8282_;
wire _8283_;
wire _8284_;
wire _8285_;
wire _8286_;
wire _8287_;
wire _8288_;
wire _8289_;
wire _8290_;
wire _8291_;
wire _8292_;
wire _8293_;
wire _8294_;
wire _8295_;
wire _8296_;
wire _8297_;
wire _8298_;
wire _8299_;
wire _8300_;
wire _8301_;
wire _8302_;
wire _8303_;
wire _8304_;
wire _8305_;
wire _8306_;
wire _8307_;
wire _8308_;
wire _8309_;
wire _8310_;
wire _8311_;
wire _8312_;
wire _8313_;
wire _8314_;
wire _8315_;
wire _8316_;
wire _8317_;
wire _8318_;
wire _8319_;
wire _8320_;
wire _8321_;
wire _8322_;
wire _8323_;
wire _8324_;
wire _8325_;
wire _8326_;
wire _8327_;
wire _8328_;
wire _8329_;
wire _8330_;
wire _8331_;
wire _8332_;
wire _8333_;
wire _8334_;
wire _8335_;
wire _8336_;
wire _8337_;
wire _8338_;
wire _8339_;
wire _8340_;
wire _8341_;
wire _8342_;
wire _8343_;
wire _8344_;
wire _8345_;
wire _8346_;
wire _8347_;
wire _8348_;
wire _8349_;
wire _8350_;
wire _8351_;
wire _8352_;
wire _8353_;
wire _8354_;
wire _8355_;
wire _8356_;
wire _8357_;
wire _8358_;
wire _8359_;
wire _8360_;
wire _8361_;
wire _8362_;
wire _8363_;
wire _8364_;
wire _8365_;
wire _8366_;
wire _8367_;
wire _8368_;
wire _8369_;
wire _8370_;
wire _8371_;
wire _8372_;
wire _8373_;
wire _8374_;
wire _8375_;
wire _8376_;
wire _8377_;
wire _8378_;
wire _8379_;
wire _8380_;
wire _8381_;
wire _8382_;
wire _8383_;
wire _8384_;
wire _8385_;
wire _8386_;
wire _8387_;
wire _8388_;
wire _8389_;
wire _8390_;
wire _8391_;
wire _8392_;
wire _8393_;
wire _8394_;
wire _8395_;
wire _8396_;
wire _8397_;
wire _8398_;
wire _8399_;
wire _8400_;
wire _8401_;
wire _8402_;
wire _8403_;
wire _8404_;
wire _8405_;
wire _8406_;
wire _8407_;
wire _8408_;
wire _8409_;
wire _8410_;
wire _8411_;
wire _8412_;
wire _8413_;
wire _8414_;
wire _8415_;
wire _8416_;
wire _8417_;
wire _8418_;
wire _8419_;
wire _8420_;
wire _8421_;
wire _8422_;
wire _8423_;
wire _8424_;
wire _8425_;
wire _8426_;
wire _8427_;
wire _8428_;
wire _8429_;
wire _8430_;
wire _8431_;
wire _8432_;
wire _8433_;
wire _8434_;
wire _8435_;
wire _8436_;
wire _8437_;
wire _8438_;
wire _8439_;
wire _8440_;
wire _8441_;
wire _8442_;
wire _8443_;
wire _8444_;
wire _8445_;
wire _8446_;
wire _8447_;
wire _8448_;
wire _8449_;
wire _8450_;
wire _8451_;
wire _8452_;
wire _8453_;
wire _8454_;
wire _8455_;
wire _8456_;
wire _8457_;
wire _8458_;
wire _8459_;
wire _8460_;
wire _8461_;
wire _8462_;
wire _8463_;
wire _8464_;
wire _8465_;
wire _8466_;
wire _8467_;
wire _8468_;
wire _8469_;
wire _8470_;
wire _8471_;
wire _8472_;
wire _8473_;
wire _8474_;
wire _8475_;
wire _8476_;
wire _8477_;
wire _8478_;
wire _8479_;
wire _8480_;
wire _8481_;
wire _8482_;
wire _8483_;
wire _8484_;
wire _8485_;
wire _8486_;
wire _8487_;
wire _8488_;
wire _8489_;
wire _8490_;
wire _8491_;
wire _8492_;
wire _8493_;
wire _8494_;
wire _8495_;
wire _8496_;
wire _8497_;
wire _8498_;
wire _8499_;
wire _8500_;
wire _8501_;
wire _8502_;
wire _8503_;
wire _8504_;
wire _8505_;
wire _8506_;
wire _8507_;
wire _8508_;
wire _8509_;
wire _8510_;
wire _8511_;
wire _8512_;
wire _8513_;
wire _8514_;
wire _8515_;
wire _8516_;
wire _8517_;
wire _8518_;
wire _8519_;
wire _8520_;
wire _8521_;
wire _8522_;
wire _8523_;
wire _8524_;
wire _8525_;
wire _8526_;
wire _8527_;
wire _8528_;
wire _8529_;
wire _8530_;
wire _8531_;
wire _8532_;
wire _8533_;
wire _8534_;
wire _8535_;
wire _8536_;
wire _8537_;
wire _8538_;
wire _8539_;
wire _8540_;
wire _8541_;
wire _8542_;
wire _8543_;
wire _8544_;
wire _8545_;
wire _8546_;
wire _8547_;
wire _8548_;
wire _8549_;
wire _8550_;
wire _8551_;
wire _8552_;
wire _8553_;
wire _8554_;
wire _8555_;
wire _8556_;
wire _8557_;
wire _8558_;
wire _8559_;
wire _8560_;
wire _8561_;
wire _8562_;
wire _8563_;
wire _8564_;
wire _8565_;
wire _8566_;
wire _8567_;
wire _8568_;
wire _8569_;
wire _8570_;
wire _8571_;
wire _8572_;
wire _8573_;
wire _8574_;
wire _8575_;
wire _8576_;
wire _8577_;
wire _8578_;
wire _8579_;
wire _8580_;
wire _8581_;
wire _8582_;
wire _8583_;
wire _8584_;
wire _8585_;
wire _8586_;
wire _8587_;
wire _8588_;
wire _8589_;
wire _8590_;
wire _8591_;
wire _8592_;
wire _8593_;
wire _8594_;
wire _8595_;
wire _8596_;
wire _8597_;
wire _8598_;
wire _8599_;
wire _8600_;
wire _8601_;
wire _8602_;
wire _8603_;
wire _8604_;
wire _8605_;
wire _8606_;
wire _8607_;
wire _8608_;
wire _8609_;
wire _8610_;
wire _8611_;
wire _8612_;
wire _8613_;
wire _8614_;
wire _8615_;
wire _8616_;
wire _8617_;
wire _8618_;
wire _8619_;
wire _8620_;
wire _8621_;
wire _8622_;
wire _8623_;
wire _8624_;
wire _8625_;
wire _8626_;
wire _8627_;
wire _8628_;
wire _8629_;
wire _8630_;
wire _8631_;
wire _8632_;
wire _8633_;
wire _8634_;
wire _8635_;
wire _8636_;
wire _8637_;
wire _8638_;
wire _8639_;
wire _8640_;
wire _8641_;
wire _8642_;
wire _8643_;
wire _8644_;
wire _8645_;
wire _8646_;
wire _8647_;
wire _8648_;
wire _8649_;
wire _8650_;
wire _8651_;
wire _8652_;
wire _8653_;
wire _8654_;
wire _8655_;
wire _8656_;
wire _8657_;
wire _8658_;
wire _8659_;
wire _8660_;
wire _8661_;
wire _8662_;
wire _8663_;
wire _8664_;
wire _8665_;
wire _8666_;
wire _8667_;
wire _8668_;
wire _8669_;
wire _8670_;
wire _8671_;
wire _8672_;
wire _8673_;
wire _8674_;
wire _8675_;
wire _8676_;
wire _8677_;
wire _8678_;
wire _8679_;
wire _8680_;
wire _8681_;
wire _8682_;
wire _8683_;
wire _8684_;
wire _8685_;
wire _8686_;
wire _8687_;
wire _8688_;
wire _8689_;
wire _8690_;
wire _8691_;
wire _8692_;
wire _8693_;
wire _8694_;
wire _8695_;
wire _8696_;
wire _8697_;
wire _8698_;
wire _8699_;
wire _8700_;
wire _8701_;
wire _8702_;
wire _8703_;
wire _8704_;
wire _8705_;
wire _8706_;
wire _8707_;
wire _8708_;
wire _8709_;
wire _8710_;
wire _8711_;
wire _8712_;
wire _8713_;
wire _8714_;
wire _8715_;
wire _8716_;
wire _8717_;
wire _8718_;
wire _8719_;
wire _8720_;
wire _8721_;
wire _8722_;
wire _8723_;
wire _8724_;
wire _8725_;
wire _8726_;
wire _8727_;
wire _8728_;
wire _8729_;
wire _8730_;
wire _8731_;
wire _8732_;
wire _8733_;
wire _8734_;
wire _8735_;
wire _8736_;
wire _8737_;
wire _8738_;
wire _8739_;
wire _8740_;
wire _8741_;
wire _8742_;
wire _8743_;
wire _8744_;
wire _8745_;
wire _8746_;
wire _8747_;
wire _8748_;
wire _8749_;
wire _8750_;
wire _8751_;
wire _8752_;
wire _8753_;
wire _8754_;
wire _8755_;
wire _8756_;
wire _8757_;
wire _8758_;
wire _8759_;
wire _8760_;
wire _8761_;
wire _8762_;
wire _8763_;
wire _8764_;
wire _8765_;
wire _8766_;
wire _8767_;
wire _8768_;
wire _8769_;
wire _8770_;
wire _8771_;
wire _8772_;
wire _8773_;
wire _8774_;
wire _8775_;
wire _8776_;
wire _8777_;
wire _8778_;
wire _8779_;
wire _8780_;
wire _8781_;
wire _8782_;
wire _8783_;
wire _8784_;
wire _8785_;
wire _8786_;
wire _8787_;
wire _8788_;
wire _8789_;
wire _8790_;
wire _8791_;
wire _8792_;
wire _8793_;
wire _8794_;
wire _8795_;
wire _8796_;
wire _8797_;
wire _8798_;
wire _8799_;
wire _8800_;
wire _8801_;
wire _8802_;
wire _8803_;
wire _8804_;
wire _8805_;
wire _8806_;
wire _8807_;
wire _8808_;
wire _8809_;
wire _8810_;
wire _8811_;
wire _8812_;
wire _8813_;
wire _8814_;
wire _8815_;
wire _8816_;
wire _8817_;
wire _8818_;
wire _8819_;
wire _8820_;
wire _8821_;
wire _8822_;
wire _8823_;
wire _8824_;
wire _8825_;
wire _8826_;
wire _8827_;
wire _8828_;
wire _8829_;
wire _8830_;
wire _8831_;
wire _8832_;
wire _8833_;
wire _8834_;
wire _8835_;
wire _8836_;
wire _8837_;
wire _8838_;
wire _8839_;
wire _8840_;
wire _8841_;
wire _8842_;
wire _8843_;
wire _8844_;
wire _8845_;
wire _8846_;
wire _8847_;
wire _8848_;
wire _8849_;
wire _8850_;
wire _8851_;
wire _8852_;
wire _8853_;
wire _8854_;
wire _8855_;
wire _8856_;
wire _8857_;
wire _8858_;
wire _8859_;
wire _8860_;
wire _8861_;
wire _8862_;
wire _8863_;
wire _8864_;
wire _8865_;
wire _8866_;
wire _8867_;
wire _8868_;
wire _8869_;
wire _8870_;
wire _8871_;
wire _8872_;
wire _8873_;
wire _8874_;
wire _8875_;
wire _8876_;
wire _8877_;
wire _8878_;
wire _8879_;
wire _8880_;
wire _8881_;
wire _8882_;
wire _8883_;
wire _8884_;
wire _8885_;
wire _8886_;
wire _8887_;
wire _8888_;
wire _8889_;
wire _8890_;
wire _8891_;
wire _8892_;
wire _8893_;
wire _8894_;
wire _8895_;
wire _8896_;
wire _8897_;
wire _8898_;
wire _8899_;
wire _8900_;
wire _8901_;
wire _8902_;
wire _8903_;
wire _8904_;
wire _8905_;
wire _8906_;
wire _8907_;
wire _8908_;
wire _8909_;
wire _8910_;
wire _8911_;
wire _8912_;
wire _8913_;
wire _8914_;
wire _8915_;
wire _8916_;
wire _8917_;
wire _8918_;
wire _8919_;
wire _8920_;
wire _8921_;
wire _8922_;
wire _8923_;
wire _8924_;
wire _8925_;
wire _8926_;
wire _8927_;
wire _8928_;
wire _8929_;
wire _8930_;
wire _8931_;
wire _8932_;
wire _8933_;
wire _8934_;
wire _8935_;
wire _8936_;
wire _8937_;
wire _8938_;
wire _8939_;
wire _8940_;
wire _8941_;
wire _8942_;
wire _8943_;
wire _8944_;
wire _8945_;
wire _8946_;
wire _8947_;
wire _8948_;
wire _8949_;
wire _8950_;
wire _8951_;
wire _8952_;
wire _8953_;
wire _8954_;
wire _8955_;
wire _8956_;
wire _8957_;
wire _8958_;
wire _8959_;
wire _8960_;
wire _8961_;
wire _8962_;
wire _8963_;
wire _8964_;
wire _8965_;
wire _8966_;
wire _8967_;
wire _8968_;
wire _8969_;
wire _8970_;
wire _8971_;
wire _8972_;
wire _8973_;
wire _8974_;
wire _8975_;
wire _8976_;
wire _8977_;
wire _8978_;
wire _8979_;
wire _8980_;
wire _8981_;
wire _8982_;
wire _8983_;
wire _8984_;
wire _8985_;
wire _8986_;
wire _8987_;
wire _8988_;
wire _8989_;
wire _8990_;
wire _8991_;
wire _8992_;
wire _8993_;
wire _8994_;
wire _8995_;
wire _8996_;
wire _8997_;
wire _8998_;
wire _8999_;
wire _9000_;
wire _9001_;
wire _9002_;
wire _9003_;
wire _9004_;
wire _9005_;
wire _9006_;
wire _9007_;
wire _9008_;
wire _9009_;
wire _9010_;
wire _9011_;
wire _9012_;
wire _9013_;
wire _9014_;
wire _9015_;
wire _9016_;
wire _9017_;
wire _9018_;
wire _9019_;
wire _9020_;
wire _9021_;
wire _9022_;
wire _9023_;
wire _9024_;
wire _9025_;
wire _9026_;
wire _9027_;
wire _9028_;
wire _9029_;
wire _9030_;
wire _9031_;
wire _9032_;
wire _9033_;
wire _9034_;
wire _9035_;
wire _9036_;
wire _9037_;
wire _9038_;
wire _9039_;
wire _9040_;
wire _9041_;
wire _9042_;
wire _9043_;
wire _9044_;
wire _9045_;
wire _9046_;
wire _9047_;
wire _9048_;
wire _9049_;
wire _9050_;
wire _9051_;
wire _9052_;
wire _9053_;
wire _9054_;
wire _9055_;
wire _9056_;
wire _9057_;
wire _9058_;
wire _9059_;
wire _9060_;
wire _9061_;
wire _9062_;
wire _9063_;
wire _9064_;
wire _9065_;
wire _9066_;
wire _9067_;
wire _9068_;
wire _9069_;
wire _9070_;
wire _9071_;
wire _9072_;
wire _9073_;
wire _9074_;
wire _9075_;
wire _9076_;
wire _9077_;
wire _9078_;
wire _9079_;
wire _9080_;
wire _9081_;
wire _9082_;
wire _9083_;
wire _9084_;
wire _9085_;
wire _9086_;
wire _9087_;
wire _9088_;
wire _9089_;
wire _9090_;
wire _9091_;
wire _9092_;
wire _9093_;
wire _9094_;
wire _9095_;
wire _9096_;
wire _9097_;
wire _9098_;
wire _9099_;
wire _9100_;
wire _9101_;
wire _9102_;
wire _9103_;
wire _9104_;
wire _9105_;
wire _9106_;
wire _9107_;
wire _9108_;
wire _9109_;
wire _9110_;
wire _9111_;
wire _9112_;
wire _9113_;
wire _9114_;
wire _9115_;
wire _9116_;
wire _9117_;
wire _9118_;
wire _9119_;
wire _9120_;
wire _9121_;
wire _9122_;
wire _9123_;
wire _9124_;
wire _9125_;
wire _9126_;
wire _9127_;
wire _9128_;
wire _9129_;
wire _9130_;
wire _9131_;
wire _9132_;
wire _9133_;
wire _9134_;
wire _9135_;
wire _9136_;
wire _9137_;
wire _9138_;
wire _9139_;
wire _9140_;
wire _9141_;
wire _9142_;
wire _9143_;
wire _9144_;
wire _9145_;
wire _9146_;
wire _9147_;
wire _9148_;
wire _9149_;
wire _9150_;
wire _9151_;
wire _9152_;
wire _9153_;
wire _9154_;
wire _9155_;
wire _9156_;
wire _9157_;
wire _9158_;
wire _9159_;
wire _9160_;
wire _9161_;
wire _9162_;
wire _9163_;
wire _9164_;
wire _9165_;
wire _9166_;
wire _9167_;
wire _9168_;
wire _9169_;
wire _9170_;
wire _9171_;
wire _9172_;
wire _9173_;
wire _9174_;
wire _9175_;
wire _9176_;
wire _9177_;
wire _9178_;
wire _9179_;
wire _9180_;
wire _9181_;
wire _9182_;
wire _9183_;
wire _9184_;
wire _9185_;
wire _9186_;
wire _9187_;
wire _9188_;
wire _9189_;
wire _9190_;
wire _9191_;
wire _9192_;
wire _9193_;
wire _9194_;
wire _9195_;
wire _9196_;
wire _9197_;
wire _9198_;
wire _9199_;
wire _9200_;
wire _9201_;
wire _9202_;
wire _9203_;
wire _9204_;
wire _9205_;
wire _9206_;
wire _9207_;
wire _9208_;
wire _9209_;
wire _9210_;
wire _9211_;
wire _9212_;
wire _9213_;
wire _9214_;
wire _9215_;
wire _9216_;
wire _9217_;
wire _9218_;
wire _9219_;
wire _9220_;
wire _9221_;
wire _9222_;
wire _9223_;
wire _9224_;
wire _9225_;
wire _9226_;
wire _9227_;
wire _9228_;
wire _9229_;
wire _9230_;
wire _9231_;
wire _9232_;
wire _9233_;
wire _9234_;
wire _9235_;
wire _9236_;
wire _9237_;
wire _9238_;
wire _9239_;
wire _9240_;
wire _9241_;
wire _9242_;
wire _9243_;
wire _9244_;
wire _9245_;
wire _9246_;
wire _9247_;
wire _9248_;
wire _9249_;
wire _9250_;
wire _9251_;
wire _9252_;
wire _9253_;
wire _9254_;
wire _9255_;
wire _9256_;
wire _9257_;
wire _9258_;
wire _9259_;
wire _9260_;
wire _9261_;
wire _9262_;
wire _9263_;
wire _9264_;
wire _9265_;
wire _9266_;
wire _9267_;
wire _9268_;
wire _9269_;
wire _9270_;
wire _9271_;
wire _9272_;
wire _9273_;
wire _9274_;
wire _9275_;
wire _9276_;
wire _9277_;
wire _9278_;
wire _9279_;
wire _9280_;
wire _9281_;
wire _9282_;
wire _9283_;
wire _9284_;
wire _9285_;
wire _9286_;
wire _9287_;
wire _9288_;
wire _9289_;
wire _9290_;
wire _9291_;
wire _9292_;
wire _9293_;
wire _9294_;
wire _9295_;
wire _9296_;
wire _9297_;
wire _9298_;
wire _9299_;
wire _9300_;
wire _9301_;
wire _9302_;
wire _9303_;
wire _9304_;
wire _9305_;
wire _9306_;
wire _9307_;
wire _9308_;
wire _9309_;
wire _9310_;
wire _9311_;
wire _9312_;
wire _9313_;
wire _9314_;
wire _9315_;
wire _9316_;
wire _9317_;
wire _9318_;
wire _9319_;
wire _9320_;
wire _9321_;
wire _9322_;
wire _9323_;
wire _9324_;
wire _9325_;
wire _9326_;
wire _9327_;
wire _9328_;
wire _9329_;
wire _9330_;
wire _9331_;
wire _9332_;
wire _9333_;
wire _9334_;
wire _9335_;
wire _9336_;
wire _9337_;
wire _9338_;
wire _9339_;
wire _9340_;
wire _9341_;
wire _9342_;
wire _9343_;
wire _9344_;
wire _9345_;
wire _9346_;
wire _9347_;
wire _9348_;
wire _9349_;
wire _9350_;
wire _9351_;
wire _9352_;
wire _9353_;
wire _9354_;
wire _9355_;
wire _9356_;
wire _9357_;
wire _9358_;
wire _9359_;
wire _9360_;
wire _9361_;
wire _9362_;
wire _9363_;
wire _9364_;
wire _9365_;
wire _9366_;
wire _9367_;
wire _9368_;
wire _9369_;
wire _9370_;
wire _9371_;
wire _9372_;
wire _9373_;
wire _9374_;
wire _9375_;
wire _9376_;
wire _9377_;
wire _9378_;
wire _9379_;
wire _9380_;
wire _9381_;
wire _9382_;
wire _9383_;
wire _9384_;
wire _9385_;
wire _9386_;
wire _9387_;
wire _9388_;
wire _9389_;
wire _9390_;
wire _9391_;
wire _9392_;
wire _9393_;
wire _9394_;
wire _9395_;
wire _9396_;
wire _9397_;
wire _9398_;
wire _9399_;
wire _9400_;
wire _9401_;
wire _9402_;
wire _9403_;
wire _9404_;
wire _9405_;
wire _9406_;
wire _9407_;
wire _9408_;
wire _9409_;
wire _9410_;
wire _9411_;
wire _9412_;
wire _9413_;
wire _9414_;
wire _9415_;
wire _9416_;
wire _9417_;
wire _9418_;
wire _9419_;
wire _9420_;
wire _9421_;
wire _9422_;
wire _9423_;
wire _9424_;
wire _9425_;
wire _9426_;
wire _9427_;
wire _9428_;
wire _9429_;
wire _9430_;
wire _9431_;
wire _9432_;
wire _9433_;
wire _9434_;
wire _9435_;
wire _9436_;
wire _9437_;
wire _9438_;
wire _9439_;
wire _9440_;
wire _9441_;
wire _9442_;
wire _9443_;
wire _9444_;
wire _9445_;
wire _9446_;
wire _9447_;
wire _9448_;
wire _9449_;
wire _9450_;
wire _9451_;
wire _9452_;
wire _9453_;
wire _9454_;
wire _9455_;
wire _9456_;
wire _9457_;
wire _9458_;
wire _9459_;
wire _9460_;
wire _9461_;
wire _9462_;
wire _9463_;
wire _9464_;
wire _9465_;
wire _9466_;
wire _9467_;
wire _9468_;
wire _9469_;
wire _9470_;
wire _9471_;
wire _9472_;
wire _9473_;
wire _9474_;
wire _9475_;
wire _9476_;
wire _9477_;
wire _9478_;
wire _9479_;
wire _9480_;
wire _9481_;
wire _9482_;
wire _9483_;
wire _9484_;
wire _9485_;
wire _9486_;
wire _9487_;
wire _9488_;
wire _9489_;
wire _9490_;
wire _9491_;
wire _9492_;
wire _9493_;
wire _9494_;
wire _9495_;
wire _9496_;
wire _9497_;
wire _9498_;
wire _9499_;
wire _9500_;
wire _9501_;
wire _9502_;
wire _9503_;
wire _9504_;
wire _9505_;
wire _9506_;
wire _9507_;
wire _9508_;
wire _9509_;
wire _9510_;
wire _9511_;
wire _9512_;
wire _9513_;
wire _9514_;
wire _9515_;
wire _9516_;
wire _9517_;
wire _9518_;
wire _9519_;
wire _9520_;
wire _9521_;
wire _9522_;
wire _9523_;
wire _9524_;
wire _9525_;
wire _9526_;
wire _9527_;
wire _9528_;
wire _9529_;
wire _9530_;
wire _9531_;
wire _9532_;
wire _9533_;
wire _9534_;
wire _9535_;
wire _9536_;
wire _9537_;
wire _9538_;
wire _9539_;
wire _9540_;
wire _9541_;
wire _9542_;
wire _9543_;
wire _9544_;
wire _9545_;
wire _9546_;
wire _9547_;
wire _9548_;
wire _9549_;
wire _9550_;
wire _9551_;
wire _9552_;
wire _9553_;
wire _9554_;
wire _9555_;
wire _9556_;
wire _9557_;
wire _9558_;
wire _9559_;
wire _9560_;
wire _9561_;
wire _9562_;
wire _9563_;
wire _9564_;
wire _9565_;
wire _9566_;
wire _9567_;
wire _9568_;
wire _9569_;
wire _9570_;
wire _9571_;
wire _9572_;
wire _9573_;
wire _9574_;
wire _9575_;
wire _9576_;
wire _9577_;
wire _9578_;
wire _9579_;
wire _9580_;
wire _9581_;
wire _9582_;
wire _9583_;
wire _9584_;
wire _9585_;
wire _9586_;
wire _9587_;
wire _9588_;
wire _9589_;
wire _9590_;
wire _9591_;
wire _9592_;
wire _9593_;
wire _9594_;
wire _9595_;
wire _9596_;
wire _9597_;
wire _9598_;
wire _9599_;
wire _9600_;
wire _9601_;
wire _9602_;
wire _9603_;
wire _9604_;
wire _9605_;
wire _9606_;
wire _9607_;
wire _9608_;
wire _9609_;
wire _9610_;
wire _9611_;
wire _9612_;
wire _9613_;
wire _9614_;
wire _9615_;
wire _9616_;
wire _9617_;
wire _9618_;
wire _9619_;
wire _9620_;
wire _9621_;
wire _9622_;
wire _9623_;
wire _9624_;
wire _9625_;
wire _9626_;
wire _9627_;
wire _9628_;
wire _9629_;
wire _9630_;
wire _9631_;
wire _9632_;
wire _9633_;
wire _9634_;
wire _9635_;
wire _9636_;
wire _9637_;
wire _9638_;
wire _9639_;
wire _9640_;
wire _9641_;
wire _9642_;
wire _9643_;
wire _9644_;
wire _9645_;
wire _9646_;
wire _9647_;
wire _9648_;
wire _9649_;
wire _9650_;
wire _9651_;
wire _9652_;
wire _9653_;
wire _9654_;
wire _9655_;
wire _9656_;
wire _9657_;
wire _9658_;
wire _9659_;
wire _9660_;
wire _9661_;
wire _9662_;
wire _9663_;
wire _9664_;
wire _9665_;
wire _9666_;
wire _9667_;
wire _9668_;
wire _9669_;
wire _9670_;
wire _9671_;
wire _9672_;
wire _9673_;
wire _9674_;
wire _9675_;
wire _9676_;
wire _9677_;
wire _9678_;
wire _9679_;
wire _9680_;
wire _9681_;
wire _9682_;
wire _9683_;
wire _9684_;
wire _9685_;
wire _9686_;
wire _9687_;
wire _9688_;
wire _9689_;
wire _9690_;
wire _9691_;
wire _9692_;
wire _9693_;
wire _9694_;
wire _9695_;
wire _9696_;
wire _9697_;
wire _9698_;
wire _9699_;
wire _9700_;
wire _9701_;
wire _9702_;
wire _9703_;
wire _9704_;
wire _9705_;
wire _9706_;
wire _9707_;
wire _9708_;
wire _9709_;
wire _9710_;
wire _9711_;
wire _9712_;
wire _9713_;
wire _9714_;
wire _9715_;
wire _9716_;
wire _9717_;
wire _9718_;
wire _9719_;
wire _9720_;
wire _9721_;
wire _9722_;
wire _9723_;
wire _9724_;
wire _9725_;
wire _9726_;
wire _9727_;
wire _9728_;
wire _9729_;
wire _9730_;
wire _9731_;
wire _9732_;
wire _9733_;
wire _9734_;
wire _9735_;
wire _9736_;
wire _9737_;
wire _9738_;
wire _9739_;
wire _9740_;
wire _9741_;
wire _9742_;
wire _9743_;
wire _9744_;
wire _9745_;
wire _9746_;
wire _9747_;
wire _9748_;
wire _9749_;
wire _9750_;
wire _9751_;
wire _9752_;
wire _9753_;
wire _9754_;
wire _9755_;
wire _9756_;
wire _9757_;
wire _9758_;
wire _9759_;
wire _9760_;
wire _9761_;
wire _9762_;
wire _9763_;
wire _9764_;
wire _9765_;
wire _9766_;
wire _9767_;
wire _9768_;
wire _9769_;
wire _9770_;
wire _9771_;
wire _9772_;
wire _9773_;
wire _9774_;
wire _9775_;
wire _9776_;
wire _9777_;
wire _9778_;
wire _9779_;
wire _9780_;
wire _9781_;
wire _9782_;
wire _9783_;
wire _9784_;
wire _9785_;
wire _9786_;
wire _9787_;
wire _9788_;
wire _9789_;
wire _9790_;
wire _9791_;
wire _9792_;
wire _9793_;
wire _9794_;
wire _9795_;
wire _9796_;
wire _9797_;
wire _9798_;
wire _9799_;
wire _9800_;
wire _9801_;
wire _9802_;
wire _9803_;
wire _9804_;
wire _9805_;
wire _9806_;
wire _9807_;
wire _9808_;
wire _9809_;
wire _9810_;
wire _9811_;
wire _9812_;
wire _9813_;
wire _9814_;
wire _9815_;
wire _9816_;
wire _9817_;
wire _9818_;
wire _9819_;
wire _9820_;
wire _9821_;
wire _9822_;
wire _9823_;
wire _9824_;
wire _9825_;
wire _9826_;
wire _9827_;
wire _9828_;
wire _9829_;
wire _9830_;
wire _9831_;
wire _9832_;
wire _9833_;
wire _9834_;
wire _9835_;
wire _9836_;
wire _9837_;
wire _9838_;
wire _9839_;
wire _9840_;
wire _9841_;
wire _9842_;
wire _9843_;
wire _9844_;
wire _9845_;
wire _9846_;
wire _9847_;
wire _9848_;
wire _9849_;
wire _9850_;
wire _9851_;
wire _9852_;
wire _9853_;
wire _9854_;
wire _9855_;
wire _9856_;
wire _9857_;
wire _9858_;
wire _9859_;
wire _9860_;
wire _9861_;
wire _9862_;
wire _9863_;
wire _9864_;
wire _9865_;
wire _9866_;
wire _9867_;
wire _9868_;
wire _9869_;
wire _9870_;
wire _9871_;
wire _9872_;
wire _9873_;
wire _9874_;
wire _9875_;
wire _9876_;
wire _9877_;
wire _9878_;
wire _9879_;
wire _9880_;
wire _9881_;
wire _9882_;
wire _9883_;
wire _9884_;
wire _9885_;
wire _9886_;
wire _9887_;
wire _9888_;
wire _9889_;
wire _9890_;
wire _9891_;
wire _9892_;
wire _9893_;
wire _9894_;
wire _9895_;
wire _9896_;
wire _9897_;
wire _9898_;
wire _9899_;
wire _9900_;
wire _9901_;
wire _9902_;
wire _9903_;
wire _9904_;
wire _9905_;
wire _9906_;
wire _9907_;
wire _9908_;
wire _9909_;
wire _9910_;
wire _9911_;
wire _9912_;
wire _9913_;
wire _9914_;
wire _9915_;
wire _9916_;
wire _9917_;
wire _9918_;
wire _9919_;
wire _9920_;
wire _9921_;
wire _9922_;
wire _9923_;
wire _9924_;
wire _9925_;
wire _9926_;
wire _9927_;
wire _9928_;
wire _9929_;
wire _9930_;
wire _9931_;
wire _9932_;
wire _9933_;
wire _9934_;
wire _9935_;
wire _9936_;
wire _9937_;
wire _9938_;
wire _9939_;
wire _9940_;
wire _9941_;
wire _9942_;
wire _9943_;
wire _9944_;
wire _9945_;
wire _9946_;
wire _9947_;
wire _9948_;
wire _9949_;
wire _9950_;
wire _9951_;
wire _9952_;
wire _9953_;
wire _9954_;
wire _9955_;
wire _9956_;
wire _9957_;
wire _9958_;
wire _9959_;
wire _9960_;
wire _9961_;
wire _9962_;
wire _9963_;
wire _9964_;
wire _9965_;
wire _9966_;
wire _9967_;
wire _9968_;
wire _9969_;
wire _9970_;
wire _9971_;
wire _9972_;
wire _9973_;
wire _9974_;
wire _9975_;
wire _9976_;
wire _9977_;
wire _9978_;
wire _9979_;
wire _9980_;
wire _9981_;
wire _9982_;
wire _9983_;
wire _9984_;
wire _9985_;
wire _9986_;
wire _9987_;
wire _9988_;
wire _9989_;
wire _9990_;
wire _9991_;
wire _9992_;
wire _9993_;
wire _9994_;
wire _9995_;
wire _9996_;
wire _9997_;
wire _9998_;
wire _9999_;
wire _10000_;
wire _10001_;
wire _10002_;
wire _10003_;
wire _10004_;
wire _10005_;
wire _10006_;
wire _10007_;
wire _10008_;
wire _10009_;
wire _10010_;
wire _10011_;
wire _10012_;
wire _10013_;
wire _10014_;
wire _10015_;
wire _10016_;
wire _10017_;
wire _10018_;
wire _10019_;
wire _10020_;
wire _10021_;
wire _10022_;
wire _10023_;
wire _10024_;
wire _10025_;
wire _10026_;
wire _10027_;
wire _10028_;
wire _10029_;
wire _10030_;
wire _10031_;
wire _10032_;
wire _10033_;
wire _10034_;
wire _10035_;
wire _10036_;
wire _10037_;
wire _10038_;
wire _10039_;
wire _10040_;
wire _10041_;
wire _10042_;
wire _10043_;
wire _10044_;
wire _10045_;
wire _10046_;
wire _10047_;
wire _10048_;
wire _10049_;
wire _10050_;
wire _10051_;
wire _10052_;
wire _10053_;
wire _10054_;
wire _10055_;
wire _10056_;
wire _10057_;
wire _10058_;
wire _10059_;
wire _10060_;
wire _10061_;
wire _10062_;
wire _10063_;
wire _10064_;
wire _10065_;
wire _10066_;
wire _10067_;
wire _10068_;
wire _10069_;
wire _10070_;
wire _10071_;
wire _10072_;
wire _10073_;
wire _10074_;
wire _10075_;
wire _10076_;
wire _10077_;
wire _10078_;
wire _10079_;
wire _10080_;
wire _10081_;
wire _10082_;
wire _10083_;
wire _10084_;
wire _10085_;
wire _10086_;
wire _10087_;
wire _10088_;
wire _10089_;
wire _10090_;
wire _10091_;
wire _10092_;
wire _10093_;
wire _10094_;
wire _10095_;
wire _10096_;
wire _10097_;
wire _10098_;
wire _10099_;
wire _10100_;
wire _10101_;
wire _10102_;
wire _10103_;
wire _10104_;
wire _10105_;
wire _10106_;
wire _10107_;
wire _10108_;
wire _10109_;
wire _10110_;
wire _10111_;
wire _10112_;
wire _10113_;
wire _10114_;
wire _10115_;
wire _10116_;
wire _10117_;
wire _10118_;
wire _10119_;
wire _10120_;
wire _10121_;
wire _10122_;
wire _10123_;
wire _10124_;
wire _10125_;
wire _10126_;
wire _10127_;
wire _10128_;
wire _10129_;
wire _10130_;
wire _10131_;
wire _10132_;
wire _10133_;
wire _10134_;
wire _10135_;
wire _10136_;
wire _10137_;
wire _10138_;
wire _10139_;
wire _10140_;
wire _10141_;
wire _10142_;
wire _10143_;
wire _10144_;
wire _10145_;
wire _10146_;
wire _10147_;
wire _10148_;
wire _10149_;
wire _10150_;
wire _10151_;
wire _10152_;
wire _10153_;
wire _10154_;
wire _10155_;
wire _10156_;
wire _10157_;
wire _10158_;
wire _10159_;
wire _10160_;
wire _10161_;
wire _10162_;
wire _10163_;
wire _10164_;
wire _10165_;
wire _10166_;
wire _10167_;
wire _10168_;
wire _10169_;
wire _10170_;
wire _10171_;
wire _10172_;
wire _10173_;
wire _10174_;
wire _10175_;
wire _10176_;
wire _10177_;
wire _10178_;
wire _10179_;
wire _10180_;
wire _10181_;
wire _10182_;
wire _10183_;
wire _10184_;
wire _10185_;
wire _10186_;
wire _10187_;
wire _10188_;
wire _10189_;
wire _10190_;
wire _10191_;
wire _10192_;
wire _10193_;
wire _10194_;
wire _10195_;
wire _10196_;
wire _10197_;
wire _10198_;
wire _10199_;
wire _10200_;
wire _10201_;
wire _10202_;
wire _10203_;
wire _10204_;
wire _10205_;
wire _10206_;
wire _10207_;
wire _10208_;
wire _10209_;
wire _10210_;
wire _10211_;
wire _10212_;
wire _10213_;
wire _10214_;
wire _10215_;
wire _10216_;
wire _10217_;
wire _10218_;
wire _10219_;
wire _10220_;
wire _10221_;
wire _10222_;
wire _10223_;
wire _10224_;
wire _10225_;
wire _10226_;
wire _10227_;
wire _10228_;
wire _10229_;
wire _10230_;
wire _10231_;
wire _10232_;
wire _10233_;
wire _10234_;
wire _10235_;
wire _10236_;
wire _10237_;
wire _10238_;
wire _10239_;
wire _10240_;
wire _10241_;
wire _10242_;
wire _10243_;
wire _10244_;
wire _10245_;
wire _10246_;
wire _10247_;
wire _10248_;
wire _10249_;
wire _10250_;
wire _10251_;
wire _10252_;
wire _10253_;
wire _10254_;
wire _10255_;
wire _10256_;
wire _10257_;
wire _10258_;
wire _10259_;
wire _10260_;
wire _10261_;
wire _10262_;
wire _10263_;
wire _10264_;
wire _10265_;
wire _10266_;
wire _10267_;
wire _10268_;
wire _10269_;
wire _10270_;
wire _10271_;
wire _10272_;
wire _10273_;
wire _10274_;
wire _10275_;
wire _10276_;
wire _10277_;
wire _10278_;
wire _10279_;
wire _10280_;
wire _10281_;
wire _10282_;
wire _10283_;
wire _10284_;
wire _10285_;
wire _10286_;
wire _10287_;
wire _10288_;
wire _10289_;
wire _10290_;
wire _10291_;
wire _10292_;
wire _10293_;
wire _10294_;
wire _10295_;
wire _10296_;
wire _10297_;
wire _10298_;
wire _10299_;
wire _10300_;
wire _10301_;
wire _10302_;
wire _10303_;
wire _10304_;
wire _10305_;
wire _10306_;
wire _10307_;
wire _10308_;
wire _10309_;
wire _10310_;
wire _10311_;
wire _10312_;
wire _10313_;
wire _10314_;
wire _10315_;
wire _10316_;
wire _10317_;
wire _10318_;
wire _10319_;
wire _10320_;
wire _10321_;
wire _10322_;
wire _10323_;
wire _10324_;
wire _10325_;
wire _10326_;
wire _10327_;
wire _10328_;
wire _10329_;
wire _10330_;
wire _10331_;
wire _10332_;
wire _10333_;
wire _10334_;
wire _10335_;
wire _10336_;
wire _10337_;
wire _10338_;
wire _10339_;
wire _10340_;
wire _10341_;
wire _10342_;
wire _10343_;
wire _10344_;
wire _10345_;
wire _10346_;
wire _10347_;
wire _10348_;
wire _10349_;
wire _10350_;
wire _10351_;
wire _10352_;
wire _10353_;
wire _10354_;
wire _10355_;
wire _10356_;
wire _10357_;
wire _10358_;
wire _10359_;
wire _10360_;
wire _10361_;
wire _10362_;
wire _10363_;
wire _10364_;
wire _10365_;
wire _10366_;
wire _10367_;
wire _10368_;
wire _10369_;
wire _10370_;
wire _10371_;
wire _10372_;
wire _10373_;
wire _10374_;
wire _10375_;
wire _10376_;
wire _10377_;
wire _10378_;
wire _10379_;
wire _10380_;
wire _10381_;
wire _10382_;
wire _10383_;
wire _10384_;
wire _10385_;
wire _10386_;
wire _10387_;
wire _10388_;
wire _10389_;
wire _10390_;
wire _10391_;
wire _10392_;
wire _10393_;
wire _10394_;
wire _10395_;
wire _10396_;
wire _10397_;
wire _10398_;
wire _10399_;
wire _10400_;
wire _10401_;
wire _10402_;
wire _10403_;
wire _10404_;
wire _10405_;
wire _10406_;
wire _10407_;
wire _10408_;
wire _10409_;
wire _10410_;
wire _10411_;
wire _10412_;
wire _10413_;
wire _10414_;
wire _10415_;
wire _10416_;
wire _10417_;
wire _10418_;
wire _10419_;
wire _10420_;
wire _10421_;
wire _10422_;
wire _10423_;
wire _10424_;
wire _10425_;
wire _10426_;
wire _10427_;
wire _10428_;
wire _10429_;
wire _10430_;
wire _10431_;
wire _10432_;
wire _10433_;
wire _10434_;
wire _10435_;
wire _10436_;
wire _10437_;
wire _10438_;
wire _10439_;
wire _10440_;
wire _10441_;
wire _10442_;
wire _10443_;
wire _10444_;
wire _10445_;
wire _10446_;
wire _10447_;
wire _10448_;
wire _10449_;
wire _10450_;
wire _10451_;
wire _10452_;
wire _10453_;
wire _10454_;
wire _10455_;
wire _10456_;
wire _10457_;
wire _10458_;
wire _10459_;
wire _10460_;
wire _10461_;
wire _10462_;
wire _10463_;
wire _10464_;
wire _10465_;
wire _10466_;
wire _10467_;
wire _10468_;
wire _10469_;
wire _10470_;
wire _10471_;
wire _10472_;
wire _10473_;
wire _10474_;
wire _10475_;
wire _10476_;
wire _10477_;
wire _10478_;
wire _10479_;
wire _10480_;
wire _10481_;
wire _10482_;
wire _10483_;
wire _10484_;
wire _10485_;
wire _10486_;
wire _10487_;
wire _10488_;
wire _10489_;
wire _10490_;
wire _10491_;
wire _10492_;
wire _10493_;
wire _10494_;
wire _10495_;
wire _10496_;
wire _10497_;
wire _10498_;
wire _10499_;
wire _10500_;
wire _10501_;
wire _10502_;
wire _10503_;
wire _10504_;
wire _10505_;
wire _10506_;
wire _10507_;
wire _10508_;
wire _10509_;
wire _10510_;
wire _10511_;
wire _10512_;
wire _10513_;
wire _10514_;
wire _10515_;
wire _10516_;
wire _10517_;
wire _10518_;
wire _10519_;
wire _10520_;
wire _10521_;
wire _10522_;
wire _10523_;
wire _10524_;
wire _10525_;
wire _10526_;
wire _10527_;
wire _10528_;
wire _10529_;
wire _10530_;
wire _10531_;
wire _10532_;
wire _10533_;
wire _10534_;
wire _10535_;
wire _10536_;
wire _10537_;
wire _10538_;
wire _10539_;
wire _10540_;
wire _10541_;
wire _10542_;
wire _10543_;
wire _10544_;
wire _10545_;
wire _10546_;
wire _10547_;
wire _10548_;
wire _10549_;
wire _10550_;
wire _10551_;
wire _10552_;
wire _10553_;
wire _10554_;
wire _10555_;
wire _10556_;
wire _10557_;
wire _10558_;
wire _10559_;
wire _10560_;
wire _10561_;
wire _10562_;
wire _10563_;
wire _10564_;
wire _10565_;
wire _10566_;
wire _10567_;
wire _10568_;
wire _10569_;
wire _10570_;
wire _10571_;
wire _10572_;
wire _10573_;
wire _10574_;
wire _10575_;
wire _10576_;
wire _10577_;
wire _10578_;
wire _10579_;
wire _10580_;
wire _10581_;
wire _10582_;
wire _10583_;
wire _10584_;
wire _10585_;
wire _10586_;
wire _10587_;
wire _10588_;
wire _10589_;
wire _10590_;
wire _10591_;
wire _10592_;
wire _10593_;
wire _10594_;
wire _10595_;
wire _10596_;
wire _10597_;
wire _10598_;
wire _10599_;
wire _10600_;
wire _10601_;
wire _10602_;
wire _10603_;
wire _10604_;
wire _10605_;
wire _10606_;
wire _10607_;
wire _10608_;
wire _10609_;
wire _10610_;
wire _10611_;
wire _10612_;
wire _10613_;
wire _10614_;
wire _10615_;
wire _10616_;
wire _10617_;
wire _10618_;
wire _10619_;
wire _10620_;
wire _10621_;
wire _10622_;
wire _10623_;
wire _10624_;
wire _10625_;
wire _10626_;
wire _10627_;
wire _10628_;
wire _10629_;
wire _10630_;
wire _10631_;
wire _10632_;
wire _10633_;
wire _10634_;
wire _10635_;
wire _10636_;
wire _10637_;
wire _10638_;
wire _10639_;
wire _10640_;
wire _10641_;
wire _10642_;
wire _10643_;
wire _10644_;
wire _10645_;
wire _10646_;
wire _10647_;
wire _10648_;
wire _10649_;
wire _10650_;
wire _10651_;
wire _10652_;
wire _10653_;
wire _10654_;
wire _10655_;
wire _10656_;
wire _10657_;
wire _10658_;
wire _10659_;
wire _10660_;
wire _10661_;
wire _10662_;
wire _10663_;
wire _10664_;
wire _10665_;
wire _10666_;
wire _10667_;
wire _10668_;
wire _10669_;
wire _10670_;
wire _10671_;
wire _10672_;
wire _10673_;
wire _10674_;
wire _10675_;
wire _10676_;
wire _10677_;
wire _10678_;
wire _10679_;
wire _10680_;
wire _10681_;
wire _10682_;
wire _10683_;
wire _10684_;
wire _10685_;
wire _10686_;
wire _10687_;
wire _10688_;
wire _10689_;
wire _10690_;
wire _10691_;
wire _10692_;
wire _10693_;
wire _10694_;
wire _10695_;
wire _10696_;
wire _10697_;
wire _10698_;
wire _10699_;
wire _10700_;
wire _10701_;
wire _10702_;
wire _10703_;
wire _10704_;
wire _10705_;
wire _10706_;
wire _10707_;
wire _10708_;
wire _10709_;
wire _10710_;
wire _10711_;
wire _10712_;
wire _10713_;
wire _10714_;
wire _10715_;
wire _10716_;
wire _10717_;
wire _10718_;
wire _10719_;
wire _10720_;
wire _10721_;
wire _10722_;
wire _10723_;
wire _10724_;
wire _10725_;
wire _10726_;
wire _10727_;
wire _10728_;
wire _10729_;
wire _10730_;
wire _10731_;
wire _10732_;
wire _10733_;
wire _10734_;
wire _10735_;
wire _10736_;
wire _10737_;
wire _10738_;
wire _10739_;
wire _10740_;
wire _10741_;
wire _10742_;
wire _10743_;
wire _10744_;
wire _10745_;
wire _10746_;
wire _10747_;
wire _10748_;
wire _10749_;
wire _10750_;
wire _10751_;
wire _10752_;
wire _10753_;
wire _10754_;
wire _10755_;
wire _10756_;
wire _10757_;
wire _10758_;
wire _10759_;
wire _10760_;
wire _10761_;
wire _10762_;
wire _10763_;
wire _10764_;
wire _10765_;
wire _10766_;
wire _10767_;
wire _10768_;
wire _10769_;
wire _10770_;
wire _10771_;
wire _10772_;
wire _10773_;
wire _10774_;
wire _10775_;
wire _10776_;
wire _10777_;
wire _10778_;
wire _10779_;
wire _10780_;
wire _10781_;
wire _10782_;
wire _10783_;
wire _10784_;
wire _10785_;
wire _10786_;
wire _10787_;
wire _10788_;
wire _10789_;
wire _10790_;
wire _10791_;
wire _10792_;
wire _10793_;
wire _10794_;
wire _10795_;
wire _10796_;
wire _10797_;
wire _10798_;
wire _10799_;
wire _10800_;
wire _10801_;
wire _10802_;
wire _10803_;
wire _10804_;
wire _10805_;
wire _10806_;
wire _10807_;
wire _10808_;
wire _10809_;
wire _10810_;
wire _10811_;
wire _10812_;
wire _10813_;
wire _10814_;
wire _10815_;
wire _10816_;
wire _10817_;
wire _10818_;
wire _10819_;
wire _10820_;
wire _10821_;
wire _10822_;
wire _10823_;
wire _10824_;
wire _10825_;
wire _10826_;
wire _10827_;
wire _10828_;
wire _10829_;
wire _10830_;
wire _10831_;
wire _10832_;
wire _10833_;
wire _10834_;
wire _10835_;
wire _10836_;
wire _10837_;
wire _10838_;
wire _10839_;
wire _10840_;
wire _10841_;
wire _10842_;
wire _10843_;
wire _10844_;
wire _10845_;
wire _10846_;
wire _10847_;
wire _10848_;
wire _10849_;
wire _10850_;
wire _10851_;
wire _10852_;
wire _10853_;
wire _10854_;
wire _10855_;
wire _10856_;
wire _10857_;
wire _10858_;
wire _10859_;
wire _10860_;
wire _10861_;
wire _10862_;
wire _10863_;
wire _10864_;
wire _10865_;
wire _10866_;
wire _10867_;
wire _10868_;
wire _10869_;
wire _10870_;
wire _10871_;
wire _10872_;
wire _10873_;
wire _10874_;
wire _10875_;
wire _10876_;
wire _10877_;
wire _10878_;
wire _10879_;
wire _10880_;
wire _10881_;
wire _10882_;
wire _10883_;
wire _10884_;
wire _10885_;
wire _10886_;
wire _10887_;
wire _10888_;
wire _10889_;
wire _10890_;
wire _10891_;
wire _10892_;
wire _10893_;
wire _10894_;
wire _10895_;
wire _10896_;
wire _10897_;
wire _10898_;
wire _10899_;
wire _10900_;
wire _10901_;
wire _10902_;
wire _10903_;
wire _10904_;
wire _10905_;
wire _10906_;
wire _10907_;
wire _10908_;
wire _10909_;
wire _10910_;
wire _10911_;
wire _10912_;
wire _10913_;
wire _10914_;
wire _10915_;
wire _10916_;
wire _10917_;
wire _10918_;
wire _10919_;
wire _10920_;
wire _10921_;
wire _10922_;
wire _10923_;
wire _10924_;
wire _10925_;
wire _10926_;
wire _10927_;
wire _10928_;
wire _10929_;
wire _10930_;
wire _10931_;
wire _10932_;
wire _10933_;
wire _10934_;
wire _10935_;
wire _10936_;
wire _10937_;
wire _10938_;
wire _10939_;
wire _10940_;
wire _10941_;
wire _10942_;
wire _10943_;
wire _10944_;
wire _10945_;
wire _10946_;
wire _10947_;
wire _10948_;
wire _10949_;
wire _10950_;
wire _10951_;
wire _10952_;
wire _10953_;
wire _10954_;
wire _10955_;
wire _10956_;
wire _10957_;
wire _10958_;
wire _10959_;
wire _10960_;
wire _10961_;
wire _10962_;
wire _10963_;
wire _10964_;
wire _10965_;
wire _10966_;
wire _10967_;
wire _10968_;
wire _10969_;
wire _10970_;
wire _10971_;
wire _10972_;
wire _10973_;
wire _10974_;
wire _10975_;
wire _10976_;
wire _10977_;
wire _10978_;
wire _10979_;
wire _10980_;
wire _10981_;
wire _10982_;
wire _10983_;
wire _10984_;
wire _10985_;
wire _10986_;
wire _10987_;
wire _10988_;
wire _10989_;
wire _10990_;
wire _10991_;
wire _10992_;
wire _10993_;
wire _10994_;
wire _10995_;
wire _10996_;
wire _10997_;
wire _10998_;
wire _10999_;
wire _11000_;
wire _11001_;
wire _11002_;
wire _11003_;
wire _11004_;
wire _11005_;
wire _11006_;
wire _11007_;
wire _11008_;
wire _11009_;
wire _11010_;
wire _11011_;
wire _11012_;
wire _11013_;
wire _11014_;
wire _11015_;
wire _11016_;
wire _11017_;
wire _11018_;
wire _11019_;
wire _11020_;
wire _11021_;
wire _11022_;
wire _11023_;
wire _11024_;
wire _11025_;
wire _11026_;
wire _11027_;
wire _11028_;
wire _11029_;
wire _11030_;
wire _11031_;
wire _11032_;
wire _11033_;
wire _11034_;
wire _11035_;
wire _11036_;
wire _11037_;
wire _11038_;
wire _11039_;
wire _11040_;
wire _11041_;
wire _11042_;
wire _11043_;
wire _11044_;
wire _11045_;
wire _11046_;
wire _11047_;
wire _11048_;
wire _11049_;
wire _11050_;
wire _11051_;
wire _11052_;
wire _11053_;
wire _11054_;
wire _11055_;
wire _11056_;
wire _11057_;
wire _11058_;
wire _11059_;
wire _11060_;
wire _11061_;
wire _11062_;
wire _11063_;
wire _11064_;
wire _11065_;
wire _11066_;
wire _11067_;
wire _11068_;
wire _11069_;
wire _11070_;
wire _11071_;
wire _11072_;
wire _11073_;
wire _11074_;
wire _11075_;
wire _11076_;
wire _11077_;
wire _11078_;
wire _11079_;
wire _11080_;
wire _11081_;
wire _11082_;
wire _11083_;
wire _11084_;
wire _11085_;
wire _11086_;
wire _11087_;
wire _11088_;
wire _11089_;
wire _11090_;
wire _11091_;
wire _11092_;
wire _11093_;
wire _11094_;
wire _11095_;
wire _11096_;
wire _11097_;
wire _11098_;
wire _11099_;
wire _11100_;
wire _11101_;
wire _11102_;
wire _11103_;
wire _11104_;
wire _11105_;
wire _11106_;
wire _11107_;
wire _11108_;
wire _11109_;
wire _11110_;
wire _11111_;
wire _11112_;
wire _11113_;
wire _11114_;
wire _11115_;
wire _11116_;
wire _11117_;
wire _11118_;
wire _11119_;
wire _11120_;
wire _11121_;
wire _11122_;
wire _11123_;
wire _11124_;
wire _11125_;
wire _11126_;
wire _11127_;
wire _11128_;
wire _11129_;
wire _11130_;
wire _11131_;
wire _11132_;
wire _11133_;
wire _11134_;
wire _11135_;
wire _11136_;
wire _11137_;
wire _11138_;
wire _11139_;
wire _11140_;
wire _11141_;
wire _11142_;
wire _11143_;
wire _11144_;
wire _11145_;
wire _11146_;
wire _11147_;
wire _11148_;
wire _11149_;
wire _11150_;
wire _11151_;
wire _11152_;
wire _11153_;
wire _11154_;
wire _11155_;
wire _11156_;
wire _11157_;
wire _11158_;
wire _11159_;
wire _11160_;
wire _11161_;
wire _11162_;
wire _11163_;
wire _11164_;
wire _11165_;
wire _11166_;
wire _11167_;
wire _11168_;
wire _11169_;
wire _11170_;
wire _11171_;
wire _11172_;
wire _11173_;
wire _11174_;
wire _11175_;
wire _11176_;
wire _11177_;
wire _11178_;
wire _11179_;
wire _11180_;
wire _11181_;
wire _11182_;
wire _11183_;
wire _11184_;
wire _11185_;
wire _11186_;
wire _11187_;
wire _11188_;
wire _11189_;
wire _11190_;
wire _11191_;
wire _11192_;
wire _11193_;
wire _11194_;
wire _11195_;
wire _11196_;
wire _11197_;
wire _11198_;
wire _11199_;
wire _11200_;
wire _11201_;
wire _11202_;
wire _11203_;
wire _11204_;
wire _11205_;
wire _11206_;
wire _11207_;
wire _11208_;
wire _11209_;
wire _11210_;
wire _11211_;
wire _11212_;
wire _11213_;
wire _11214_;
wire _11215_;
wire _11216_;
wire _11217_;
wire _11218_;
wire _11219_;
wire _11220_;
wire _11221_;
wire _11222_;
wire _11223_;
wire _11224_;
wire _11225_;
wire _11226_;
wire _11227_;
wire _11228_;
wire _11229_;
wire _11230_;
wire _11231_;
wire _11232_;
wire _11233_;
wire _11234_;
wire _11235_;
wire _11236_;
wire _11237_;
wire _11238_;
wire _11239_;
wire _11240_;
wire _11241_;
wire _11242_;
wire _11243_;
wire _11244_;
wire _11245_;
wire _11246_;
wire _11247_;
wire _11248_;
wire _11249_;
wire _11250_;
wire _11251_;
wire _11252_;
wire _11253_;
wire _11254_;
wire _11255_;
wire _11256_;
wire _11257_;
wire _11258_;
wire _11259_;
wire _11260_;
wire _11261_;
wire _11262_;
wire _11263_;
wire _11264_;
wire _11265_;
wire _11266_;
wire _11267_;
wire _11268_;
wire _11269_;
wire _11270_;
wire _11271_;
wire _11272_;
wire _11273_;
wire _11274_;
wire _11275_;
wire _11276_;
wire _11277_;
wire _11278_;
wire _11279_;
wire _11280_;
wire _11281_;
wire _11282_;
wire _11283_;
wire _11284_;
wire _11285_;
wire _11286_;
wire _11287_;
wire _11288_;
wire _11289_;
wire _11290_;
wire _11291_;
wire _11292_;
wire _11293_;
wire _11294_;
wire _11295_;
wire _11296_;
wire _11297_;
wire _11298_;
wire _11299_;
wire _11300_;
wire _11301_;
wire _11302_;
wire _11303_;
wire _11304_;
wire _11305_;
wire _11306_;
wire _11307_;
wire _11308_;
wire _11309_;
wire _11310_;
wire _11311_;
wire _11312_;
wire _11313_;
wire _11314_;
wire _11315_;
wire _11316_;
wire _11317_;
wire _11318_;
wire _11319_;
wire _11320_;
wire _11321_;
wire _11322_;
wire _11323_;
wire _11324_;
wire _11325_;
wire _11326_;
wire _11327_;
wire _11328_;
wire _11329_;
wire _11330_;
wire _11331_;
wire _11332_;
wire _11333_;
wire _11334_;
wire _11335_;
wire _11336_;
wire _11337_;
wire _11338_;
wire _11339_;
wire _11340_;
wire _11341_;
wire _11342_;
wire _11343_;
wire _11344_;
wire _11345_;
wire _11346_;
wire _11347_;
wire _11348_;
wire _11349_;
wire _11350_;
wire _11351_;
wire _11352_;
wire _11353_;
wire _11354_;
wire _11355_;
wire _11356_;
wire _11357_;
wire _11358_;
wire _11359_;
wire _11360_;
wire _11361_;
wire _11362_;
wire _11363_;
wire _11364_;
wire _11365_;
wire _11366_;
wire _11367_;
wire _11368_;
wire _11369_;
wire _11370_;
wire _11371_;
wire _11372_;
wire _11373_;
wire _11374_;
wire _11375_;
wire _11376_;
wire _11377_;
wire _11378_;
wire _11379_;
wire _11380_;
wire _11381_;
wire _11382_;
wire _11383_;
wire _11384_;
wire _11385_;
wire _11386_;
wire _11387_;
wire _11388_;
wire _11389_;
wire _11390_;
wire _11391_;
wire _11392_;
wire _11393_;
wire _11394_;
wire _11395_;
wire _11396_;
wire _11397_;
wire _11398_;
wire _11399_;
wire _11400_;
wire _11401_;
wire _11402_;
wire _11403_;
wire _11404_;
wire _11405_;
wire _11406_;
wire _11407_;
wire _11408_;
wire _11409_;
wire _11410_;
wire _11411_;
wire _11412_;
wire _11413_;
wire _11414_;
wire _11415_;
wire _11416_;
wire _11417_;
wire _11418_;
wire _11419_;
wire _11420_;
wire _11421_;
wire _11422_;
wire _11423_;
wire _11424_;
wire _11425_;
wire _11426_;
wire _11427_;
wire _11428_;
wire _11429_;
wire _11430_;
wire _11431_;
wire _11432_;
wire _11433_;
wire _11434_;
wire _11435_;
wire _11436_;
wire _11437_;
wire _11438_;
wire _11439_;
wire _11440_;
wire _11441_;
wire _11442_;
wire _11443_;
wire _11444_;
wire _11445_;
wire _11446_;
wire _11447_;
wire _11448_;
wire _11449_;
wire _11450_;
wire _11451_;
wire _11452_;
wire _11453_;
wire _11454_;
wire _11455_;
wire _11456_;
wire _11457_;
wire _11458_;
wire _11459_;
wire _11460_;
wire _11461_;
wire _11462_;
wire _11463_;
wire _11464_;
wire _11465_;
wire _11466_;
wire _11467_;
wire _11468_;
wire _11469_;
wire _11470_;
wire _11471_;
wire _11472_;
wire _11473_;
wire _11474_;
wire _11475_;
wire _11476_;
wire _11477_;
wire _11478_;
wire _11479_;
wire _11480_;
wire _11481_;
wire _11482_;
wire _11483_;
wire _11484_;
wire _11485_;
wire _11486_;
wire _11487_;
wire _11488_;
wire _11489_;
wire _11490_;
wire _11491_;
wire _11492_;
wire _11493_;
wire _11494_;
wire _11495_;
wire _11496_;
wire _11497_;
wire _11498_;
wire _11499_;
wire _11500_;
wire _11501_;
wire _11502_;
wire _11503_;
wire _11504_;
wire _11505_;
wire _11506_;
wire _11507_;
wire _11508_;
wire _11509_;
wire _11510_;
wire _11511_;
wire _11512_;
wire _11513_;
wire _11514_;
wire _11515_;
wire _11516_;
wire _11517_;
wire _11518_;
wire _11519_;
wire _11520_;
wire _11521_;
wire _11522_;
wire _11523_;
wire _11524_;
wire _11525_;
wire _11526_;
wire _11527_;
wire _11528_;
wire _11529_;
wire _11530_;
wire _11531_;
wire _11532_;
wire _11533_;
wire _11534_;
wire _11535_;
wire _11536_;
wire _11537_;
wire _11538_;
wire _11539_;
wire _11540_;
wire _11541_;
wire _11542_;
wire _11543_;
wire _11544_;
wire _11545_;
wire _11546_;
wire _11547_;
wire _11548_;
wire _11549_;
wire _11550_;
wire _11551_;
wire _11552_;
wire _11553_;
wire _11554_;
wire _11555_;
wire _11556_;
wire _11557_;
wire _11558_;
wire _11559_;
wire _11560_;
wire _11561_;
wire _11562_;
wire _11563_;
wire _11564_;
wire _11565_;
wire _11566_;
wire _11567_;
wire _11568_;
wire _11569_;
wire _11570_;
wire _11571_;
wire _11572_;
wire _11573_;
wire _11574_;
wire _11575_;
wire _11576_;
wire _11577_;
wire _11578_;
wire _11579_;
wire _11580_;
wire _11581_;
wire _11582_;
wire _11583_;
wire _11584_;
wire _11585_;
wire _11586_;
wire _11587_;
wire _11588_;
wire _11589_;
wire _11590_;
wire _11591_;
wire _11592_;
wire _11593_;
wire _11594_;
wire _11595_;
wire _11596_;
wire _11597_;
wire _11598_;
wire _11599_;
wire _11600_;
wire _11601_;
wire _11602_;
wire _11603_;
wire _11604_;
wire _11605_;
wire _11606_;
wire _11607_;
wire _11608_;
wire _11609_;
wire _11610_;
wire _11611_;
wire _11612_;
wire _11613_;
wire _11614_;
wire _11615_;
wire _11616_;
wire _11617_;
wire _11618_;
wire _11619_;
wire _11620_;
wire _11621_;
wire _11622_;
wire _11623_;
wire _11624_;
wire _11625_;
wire _11626_;
wire _11627_;
wire _11628_;
wire _11629_;
wire _11630_;
wire _11631_;
wire _11632_;
wire _11633_;
wire _11634_;
wire _11635_;
wire _11636_;
wire _11637_;
wire _11638_;
wire _11639_;
wire _11640_;
wire _11641_;
wire _11642_;
wire _11643_;
wire _11644_;
wire _11645_;
wire _11646_;
wire _11647_;
wire _11648_;
wire _11649_;
wire _11650_;
wire _11651_;
wire _11652_;
wire _11653_;
wire _11654_;
wire _11655_;
wire _11656_;
wire _11657_;
wire _11658_;
wire _11659_;
wire _11660_;
wire _11661_;
wire _11662_;
wire _11663_;
wire _11664_;
wire _11665_;
wire _11666_;
wire _11667_;
wire _11668_;
wire _11669_;
wire _11670_;
wire _11671_;
wire _11672_;
wire _11673_;
wire _11674_;
wire _11675_;
wire _11676_;
wire _11677_;
wire _11678_;
wire _11679_;
wire _11680_;
wire _11681_;
wire _11682_;
wire _11683_;
wire _11684_;
wire _11685_;
wire _11686_;
wire _11687_;
wire _11688_;
wire _11689_;
wire _11690_;
wire _11691_;
wire _11692_;
wire _11693_;
wire _11694_;
wire _11695_;
wire _11696_;
wire _11697_;
wire _11698_;
wire _11699_;
wire _11700_;
wire _11701_;
wire _11702_;
wire _11703_;
wire _11704_;
wire _11705_;
wire _11706_;
wire _11707_;
wire _11708_;
wire _11709_;
wire _11710_;
wire _11711_;
wire _11712_;
wire _11713_;
wire _11714_;
wire _11715_;
wire _11716_;
wire _11717_;
wire _11718_;
wire _11719_;
wire _11720_;
wire _11721_;
wire _11722_;
wire _11723_;
wire _11724_;
wire _11725_;
wire _11726_;
wire _11727_;
wire _11728_;
wire _11729_;
wire _11730_;
wire _11731_;
wire _11732_;
wire _11733_;
wire _11734_;
wire _11735_;
wire _11736_;
wire _11737_;
wire _11738_;
wire _11739_;
wire _11740_;
wire _11741_;
wire _11742_;
wire _11743_;
wire _11744_;
wire _11745_;
wire _11746_;
wire _11747_;
wire _11748_;
wire _11749_;
wire _11750_;
wire _11751_;
wire _11752_;
wire _11753_;
wire _11754_;
wire _11755_;
wire _11756_;
wire _11757_;
wire _11758_;
wire _11759_;
wire _11760_;
wire _11761_;
wire _11762_;
wire _11763_;
wire _11764_;
wire _11765_;
wire _11766_;
wire _11767_;
wire _11768_;
wire _11769_;
wire _11770_;
wire _11771_;
wire _11772_;
wire _11773_;
wire _11774_;
wire _11775_;
wire _11776_;
wire _11777_;
wire _11778_;
wire _11779_;
wire _11780_;
wire _11781_;
wire _11782_;
wire _11783_;
wire _11784_;
wire _11785_;
wire _11786_;
wire _11787_;
wire _11788_;
wire _11789_;
wire _11790_;
wire _11791_;
wire _11792_;
wire _11793_;
wire _11794_;
wire _11795_;
wire _11796_;
wire _11797_;
wire _11798_;
wire _11799_;
wire _11800_;
wire _11801_;
wire _11802_;
wire _11803_;
wire _11804_;
wire _11805_;
wire _11806_;
wire _11807_;
wire _11808_;
wire _11809_;
wire _11810_;
wire _11811_;
wire _11812_;
wire _11813_;
wire _11814_;
wire _11815_;
wire _11816_;
wire _11817_;
wire _11818_;
wire _11819_;
wire _11820_;
wire _11821_;
wire _11822_;
wire _11823_;
wire _11824_;
wire _11825_;
wire _11826_;
wire _11827_;
wire _11828_;
wire _11829_;
wire _11830_;
wire _11831_;
wire _11832_;
wire _11833_;
wire _11834_;
wire _11835_;
wire _11836_;
wire _11837_;
wire _11838_;
wire _11839_;
wire _11840_;
wire _11841_;
wire _11842_;
wire _11843_;
wire _11844_;
wire _11845_;
wire _11846_;
wire _11847_;
wire _11848_;
wire _11849_;
wire _11850_;
wire _11851_;
wire _11852_;
wire _11853_;
wire _11854_;
wire _11855_;
wire _11856_;
wire _11857_;
wire _11858_;
wire _11859_;
wire _11860_;
wire _11861_;
wire _11862_;
wire _11863_;
wire _11864_;
wire _11865_;
wire _11866_;
wire _11867_;
wire _11868_;
wire _11869_;
wire _11870_;
wire _11871_;
wire _11872_;
wire _11873_;
wire _11874_;
wire _11875_;
wire _11876_;
wire _11877_;
wire _11878_;
wire _11879_;
wire _11880_;
wire _11881_;
wire _11882_;
wire _11883_;
wire _11884_;
wire _11885_;
wire _11886_;
wire _11887_;
wire _11888_;
wire _11889_;
wire _11890_;
wire _11891_;
wire _11892_;
wire _11893_;
wire _11894_;
wire _11895_;
wire _11896_;
wire _11897_;
wire _11898_;
wire _11899_;
wire _11900_;
wire _11901_;
wire _11902_;
wire _11903_;
wire _11904_;
wire _11905_;
wire _11906_;
wire _11907_;
wire _11908_;
wire _11909_;
wire _11910_;
wire _11911_;
wire _11912_;
wire _11913_;
wire _11914_;
wire _11915_;
wire _11916_;
wire _11917_;
wire _11918_;
wire _11919_;
wire _11920_;
wire _11921_;
wire _11922_;
wire _11923_;
wire _11924_;
wire _11925_;
wire _11926_;
wire _11927_;
wire _11928_;
wire _11929_;
wire _11930_;
wire _11931_;
wire _11932_;
wire _11933_;
wire _11934_;
wire _11935_;
wire _11936_;
wire _11937_;
wire _11938_;
wire _11939_;
wire _11940_;
wire _11941_;
wire _11942_;
wire _11943_;
wire _11944_;
wire _11945_;
wire _11946_;
wire _11947_;
wire _11948_;
wire _11949_;
wire _11950_;
wire _11951_;
wire _11952_;
wire _11953_;
wire _11954_;
wire _11955_;
wire _11956_;
wire _11957_;
wire _11958_;
wire _11959_;
wire _11960_;
wire _11961_;
wire _11962_;
wire _11963_;
wire _11964_;
wire _11965_;
wire _11966_;
wire _11967_;
wire _11968_;
wire _11969_;
wire _11970_;
wire _11971_;
wire _11972_;
wire _11973_;
wire _11974_;
wire _11975_;
wire _11976_;
wire _11977_;
wire _11978_;
wire _11979_;
wire _11980_;
wire _11981_;
wire _11982_;
wire _11983_;
wire _11984_;
wire _11985_;
wire _11986_;
wire _11987_;
wire _11988_;
wire _11989_;
wire _11990_;
wire _11991_;
wire _11992_;
wire _11993_;
wire _11994_;
wire _11995_;
wire _11996_;
wire _11997_;
wire _11998_;
wire _11999_;
wire _12000_;
wire _12001_;
wire _12002_;
wire _12003_;
wire _12004_;
wire _12005_;
wire _12006_;
wire _12007_;
wire _12008_;
wire _12009_;
wire _12010_;
wire _12011_;
wire _12012_;
wire _12013_;
wire _12014_;
wire _12015_;
wire _12016_;
wire _12017_;
wire _12018_;
wire _12019_;
wire _12020_;
wire _12021_;
wire _12022_;
wire _12023_;
wire _12024_;
wire _12025_;
wire _12026_;
wire _12027_;
wire _12028_;
wire _12029_;
wire _12030_;
wire _12031_;
wire _12032_;
wire _12033_;
wire _12034_;
wire _12035_;
wire _12036_;
wire _12037_;
wire _12038_;
wire _12039_;
wire _12040_;
wire _12041_;
wire _12042_;
wire _12043_;
wire _12044_;
wire _12045_;
wire _12046_;
wire _12047_;
wire _12048_;
wire _12049_;
wire _12050_;
wire _12051_;
wire _12052_;
wire _12053_;
wire _12054_;
wire _12055_;
wire _12056_;
wire _12057_;
wire _12058_;
wire _12059_;
wire _12060_;
wire _12061_;
wire _12062_;
wire _12063_;
wire _12064_;
wire _12065_;
wire _12066_;
wire _12067_;
wire _12068_;
wire _12069_;
wire _12070_;
wire _12071_;
wire _12072_;
wire _12073_;
wire _12074_;
wire _12075_;
wire _12076_;
wire _12077_;
wire _12078_;
wire _12079_;
wire _12080_;
wire _12081_;
wire _12082_;
wire _12083_;
wire _12084_;
wire _12085_;
wire _12086_;
wire _12087_;
wire _12088_;
wire _12089_;
wire _12090_;
wire _12091_;
wire _12092_;
wire _12093_;
wire _12094_;
wire _12095_;
wire _12096_;
wire _12097_;
wire _12098_;
wire _12099_;
wire _12100_;
wire _12101_;
wire _12102_;
wire _12103_;
wire _12104_;
wire _12105_;
wire _12106_;
wire _12107_;
wire _12108_;
wire _12109_;
wire _12110_;
wire _12111_;
wire _12112_;
wire _12113_;
wire _12114_;
wire _12115_;
wire _12116_;
wire _12117_;
wire _12118_;
wire _12119_;
wire _12120_;
wire _12121_;
wire _12122_;
wire _12123_;
wire _12124_;
wire _12125_;
wire _12126_;
wire _12127_;
wire _12128_;
wire _12129_;
wire _12130_;
wire _12131_;
wire _12132_;
wire _12133_;
wire _12134_;
wire _12135_;
wire _12136_;
wire _12137_;
wire _12138_;
wire _12139_;
wire _12140_;
wire _12141_;
wire _12142_;
wire _12143_;
wire _12144_;
wire _12145_;
wire _12146_;
wire _12147_;
wire _12148_;
wire _12149_;
wire _12150_;
wire _12151_;
wire _12152_;
wire _12153_;
wire _12154_;
wire _12155_;
wire _12156_;
wire _12157_;
wire _12158_;
wire _12159_;
wire _12160_;
wire _12161_;
wire _12162_;
wire _12163_;
wire _12164_;
wire _12165_;
wire _12166_;
wire _12167_;
wire _12168_;
wire _12169_;
wire _12170_;
wire _12171_;
wire _12172_;
wire _12173_;
wire _12174_;
wire _12175_;
wire _12176_;
wire _12177_;
wire _12178_;
wire _12179_;
wire _12180_;
wire _12181_;
wire _12182_;
wire _12183_;
wire _12184_;
wire _12185_;
wire _12186_;
wire _12187_;
wire _12188_;
wire _12189_;
wire _12190_;
wire _12191_;
wire _12192_;
wire _12193_;
wire _12194_;
wire _12195_;
wire _12196_;
wire _12197_;
wire _12198_;
wire _12199_;
wire _12200_;
wire _12201_;
wire _12202_;
wire _12203_;
wire _12204_;
wire _12205_;
wire _12206_;
wire _12207_;
wire _12208_;
wire _12209_;
wire _12210_;
wire _12211_;
wire _12212_;
wire _12213_;
wire _12214_;
wire _12215_;
wire _12216_;
wire _12217_;
wire _12218_;
wire _12219_;
wire _12220_;
wire _12221_;
wire _12222_;
wire _12223_;
wire _12224_;
wire _12225_;
wire _12226_;
wire _12227_;
wire _12228_;
wire _12229_;
wire _12230_;
wire _12231_;
wire _12232_;
wire _12233_;
wire _12234_;
wire _12235_;
wire _12236_;
wire _12237_;
wire _12238_;
wire _12239_;
wire _12240_;
wire _12241_;
wire _12242_;
wire _12243_;
wire _12244_;
wire _12245_;
wire _12246_;
wire _12247_;
wire _12248_;
wire _12249_;
wire _12250_;
wire _12251_;
wire _12252_;
wire _12253_;
wire _12254_;
wire _12255_;
wire _12256_;
wire _12257_;
wire _12258_;
wire _12259_;
wire _12260_;
wire _12261_;
wire _12262_;
wire _12263_;
wire _12264_;
wire _12265_;
wire _12266_;
wire _12267_;
wire _12268_;
wire _12269_;
wire _12270_;
wire _12271_;
wire _12272_;
wire _12273_;
wire _12274_;
wire _12275_;
wire _12276_;
wire _12277_;
wire _12278_;
wire _12279_;
wire _12280_;
wire _12281_;
wire _12282_;
wire _12283_;
wire _12284_;
wire _12285_;
wire _12286_;
wire _12287_;
wire _12288_;
wire _12289_;
wire _12290_;
wire _12291_;
wire _12292_;
wire _12293_;
wire _12294_;
wire _12295_;
wire _12296_;
wire _12297_;
wire _12298_;
wire _12299_;
wire _12300_;
wire _12301_;
wire _12302_;
wire _12303_;
wire _12304_;
wire _12305_;
wire _12306_;
wire _12307_;
wire _12308_;
wire _12309_;
wire _12310_;
wire _12311_;
wire _12312_;
wire _12313_;
wire _12314_;
wire _12315_;
wire _12316_;
wire _12317_;
wire _12318_;
wire _12319_;
wire _12320_;
wire _12321_;
wire _12322_;
wire _12323_;
wire _12324_;
wire _12325_;
wire _12326_;
wire _12327_;
wire _12328_;
wire _12329_;
wire _12330_;
wire _12331_;
wire _12332_;
wire _12333_;
wire _12334_;
wire _12335_;
wire _12336_;
wire _12337_;
wire _12338_;
wire _12339_;
wire _12340_;
wire _12341_;
wire _12342_;
wire _12343_;
wire _12344_;
wire _12345_;
wire _12346_;
wire _12347_;
wire _12348_;
wire _12349_;
wire _12350_;
wire _12351_;
wire _12352_;
wire _12353_;
wire _12354_;
wire _12355_;
wire _12356_;
wire _12357_;
wire _12358_;
wire _12359_;
wire _12360_;
wire _12361_;
wire _12362_;
wire _12363_;
wire _12364_;
wire _12365_;
wire _12366_;
wire _12367_;
wire _12368_;
wire _12369_;
wire _12370_;
wire _12371_;
wire _12372_;
wire _12373_;
wire _12374_;
wire _12375_;
wire _12376_;
wire _12377_;
wire _12378_;
wire _12379_;
wire _12380_;
wire _12381_;
wire _12382_;
wire _12383_;
wire _12384_;
wire _12385_;
wire _12386_;
wire _12387_;
wire _12388_;
wire _12389_;
wire _12390_;
wire _12391_;
wire _12392_;
wire _12393_;
wire _12394_;
wire _12395_;
wire _12396_;
wire _12397_;
wire _12398_;
wire _12399_;
wire _12400_;
wire _12401_;
wire _12402_;
wire _12403_;
wire _12404_;
wire _12405_;
wire _12406_;
wire _12407_;
wire _12408_;
wire _12409_;
wire _12410_;
wire _12411_;
wire _12412_;
wire _12413_;
wire _12414_;
wire _12415_;
wire _12416_;
wire _12417_;
wire _12418_;
wire _12419_;
wire _12420_;
wire _12421_;
wire _12422_;
wire _12423_;
wire _12424_;
wire _12425_;
wire _12426_;
wire _12427_;
wire _12428_;
wire _12429_;
wire _12430_;
wire _12431_;
wire _12432_;
wire _12433_;
wire _12434_;
wire _12435_;
wire _12436_;
wire _12437_;
wire _12438_;
wire _12439_;
wire _12440_;
wire _12441_;
wire _12442_;
wire _12443_;
wire _12444_;
wire _12445_;
wire _12446_;
wire _12447_;
wire _12448_;
wire _12449_;
wire _12450_;
wire _12451_;
wire _12452_;
wire _12453_;
wire _12454_;
wire _12455_;
wire _12456_;
wire _12457_;
wire _12458_;
wire _12459_;
wire _12460_;
wire _12461_;
wire _12462_;
wire _12463_;
wire _12464_;
wire _12465_;
wire _12466_;
wire _12467_;
wire _12468_;
wire _12469_;
wire _12470_;
wire _12471_;
wire _12472_;
wire _12473_;
wire _12474_;
wire _12475_;
wire _12476_;
wire _12477_;
wire _12478_;
wire _12479_;
wire _12480_;
wire _12481_;
wire _12482_;
wire _12483_;
wire _12484_;
wire _12485_;
wire _12486_;
wire _12487_;
wire _12488_;
wire _12489_;
wire _12490_;
wire _12491_;
wire _12492_;
wire _12493_;
wire _12494_;
wire _12495_;
wire _12496_;
wire _12497_;
wire _12498_;
wire _12499_;
wire _12500_;
wire _12501_;
wire _12502_;
wire _12503_;
wire _12504_;
wire _12505_;
wire _12506_;
wire _12507_;
wire _12508_;
wire _12509_;
wire _12510_;
wire _12511_;
wire _12512_;
wire _12513_;
wire _12514_;
wire _12515_;
wire _12516_;
wire _12517_;
wire _12518_;
wire _12519_;
wire _12520_;
wire _12521_;
wire _12522_;
wire _12523_;
wire _12524_;
wire _12525_;
wire _12526_;
wire _12527_;
wire _12528_;
wire _12529_;
wire _12530_;
wire _12531_;
wire _12532_;
wire _12533_;
wire _12534_;
wire _12535_;
wire _12536_;
wire _12537_;
wire _12538_;
wire _12539_;
wire _12540_;
wire _12541_;
wire _12542_;
wire _12543_;
wire _12544_;
wire _12545_;
wire _12546_;
wire _12547_;
wire _12548_;
wire _12549_;
wire _12550_;
wire _12551_;
wire _12552_;
wire _12553_;
wire _12554_;
wire _12555_;
wire _12556_;
wire _12557_;
wire _12558_;
wire _12559_;
wire _12560_;
wire _12561_;
wire _12562_;
wire _12563_;
wire _12564_;
wire _12565_;
wire _12566_;
wire _12567_;
wire _12568_;
wire _12569_;
wire _12570_;
wire _12571_;
wire _12572_;
wire _12573_;
wire _12574_;
wire _12575_;
wire _12576_;
wire _12577_;
wire _12578_;
wire _12579_;
wire _12580_;
wire _12581_;
wire _12582_;
wire _12583_;
wire _12584_;
wire _12585_;
wire _12586_;
wire _12587_;
wire _12588_;
wire _12589_;
wire _12590_;
wire _12591_;
wire _12592_;
wire _12593_;
wire _12594_;
wire _12595_;
wire _12596_;
wire _12597_;
wire _12598_;
wire _12599_;
wire _12600_;
wire _12601_;
wire _12602_;
wire _12603_;
wire _12604_;
wire _12605_;
wire _12606_;
wire _12607_;
wire _12608_;
wire _12609_;
wire _12610_;
wire _12611_;
wire _12612_;
wire _12613_;
wire _12614_;
wire _12615_;
wire _12616_;
wire _12617_;
wire _12618_;
wire _12619_;
wire _12620_;
wire _12621_;
wire _12622_;
wire _12623_;
wire _12624_;
wire _12625_;
wire _12626_;
wire _12627_;
wire _12628_;
wire _12629_;
wire _12630_;
wire _12631_;
wire _12632_;
wire _12633_;
wire _12634_;
wire _12635_;
wire _12636_;
wire _12637_;
wire _12638_;
wire _12639_;
wire _12640_;
wire _12641_;
wire _12642_;
wire _12643_;
wire _12644_;
wire _12645_;
wire _12646_;
wire _12647_;
wire _12648_;
wire _12649_;
wire _12650_;
wire _12651_;
wire _12652_;
wire _12653_;
wire _12654_;
wire _12655_;
wire _12656_;
wire _12657_;
wire _12658_;
wire _12659_;
wire _12660_;
wire _12661_;
wire _12662_;
wire _12663_;
wire _12664_;
wire _12665_;
wire _12666_;
wire _12667_;
wire _12668_;
wire _12669_;
wire _12670_;
wire _12671_;
wire _12672_;
wire _12673_;
wire _12674_;
wire _12675_;
wire _12676_;
wire _12677_;
wire _12678_;
wire _12679_;
wire _12680_;
wire _12681_;
wire _12682_;
wire _12683_;
wire _12684_;
wire _12685_;
wire _12686_;
wire _12687_;
wire _12688_;
wire _12689_;
wire _12690_;
wire _12691_;
wire _12692_;
wire _12693_;
wire _12694_;
wire _12695_;
wire _12696_;
wire _12697_;
wire _12698_;
wire _12699_;
wire _12700_;
wire _12701_;
wire _12702_;
wire _12703_;
wire _12704_;
wire _12705_;
wire _12706_;
wire _12707_;
wire _12708_;
wire _12709_;
wire _12710_;
wire _12711_;
wire _12712_;
wire _12713_;
wire _12714_;
wire _12715_;
wire _12716_;
wire _12717_;
wire _12718_;
wire _12719_;
wire _12720_;
wire _12721_;
wire _12722_;
wire _12723_;
wire _12724_;
wire _12725_;
wire _12726_;
wire _12727_;
wire _12728_;
wire _12729_;
wire _12730_;
wire _12731_;
wire _12732_;
wire _12733_;
wire _12734_;
wire _12735_;
wire _12736_;
wire _12737_;
wire _12738_;
wire _12739_;
wire _12740_;
wire _12741_;
wire _12742_;
wire _12743_;
wire _12744_;
wire _12745_;
wire _12746_;
wire _12747_;
wire _12748_;
wire _12749_;
wire _12750_;
wire _12751_;
wire _12752_;
wire _12753_;
wire _12754_;
wire _12755_;
wire _12756_;
wire _12757_;
wire _12758_;
wire _12759_;
wire _12760_;
wire _12761_;
wire _12762_;
wire _12763_;
wire _12764_;
wire _12765_;
wire _12766_;
wire _12767_;
wire _12768_;
wire _12769_;
wire _12770_;
wire _12771_;
wire _12772_;
wire _12773_;
wire _12774_;
wire _12775_;
wire _12776_;
wire _12777_;
wire _12778_;
wire _12779_;
wire _12780_;
wire _12781_;
wire _12782_;
wire _12783_;
wire _12784_;
wire _12785_;
wire _12786_;
wire _12787_;
wire _12788_;
wire _12789_;
wire _12790_;
wire _12791_;
wire _12792_;
wire _12793_;
wire _12794_;
wire _12795_;
wire _12796_;
wire _12797_;
wire _12798_;
wire _12799_;
wire _12800_;
wire _12801_;
wire _12802_;
wire _12803_;
wire _12804_;
wire _12805_;
wire _12806_;
wire _12807_;
wire _12808_;
wire _12809_;
wire _12810_;
wire _12811_;
wire _12812_;
wire _12813_;
wire _12814_;
wire _12815_;
wire _12816_;
wire _12817_;
wire _12818_;
wire _12819_;
wire _12820_;
wire _12821_;
wire _12822_;
wire _12823_;
wire _12824_;
wire _12825_;
wire _12826_;
wire _12827_;
wire _12828_;
wire _12829_;
wire _12830_;
wire _12831_;
wire _12832_;
wire _12833_;
wire _12834_;
wire _12835_;
wire _12836_;
wire _12837_;
wire _12838_;
wire _12839_;
wire _12840_;
wire _12841_;
wire _12842_;
wire _12843_;
wire _12844_;
wire _12845_;
wire _12846_;
wire _12847_;
wire _12848_;
wire _12849_;
wire _12850_;
wire _12851_;
wire _12852_;
wire _12853_;
wire _12854_;
wire _12855_;
wire _12856_;
wire _12857_;
wire _12858_;
wire _12859_;
wire _12860_;
wire _12861_;
wire _12862_;
wire _12863_;
wire _12864_;
wire _12865_;
wire _12866_;
wire _12867_;
wire _12868_;
wire _12869_;
wire _12870_;
wire _12871_;
wire _12872_;
wire _12873_;
wire _12874_;
wire _12875_;
wire _12876_;
wire _12877_;
wire _12878_;
wire _12879_;
wire _12880_;
wire _12881_;
wire _12882_;
wire _12883_;
wire _12884_;
wire _12885_;
wire _12886_;
wire _12887_;
wire _12888_;
wire _12889_;
wire _12890_;
wire _12891_;
wire _12892_;
wire _12893_;
wire _12894_;
wire _12895_;
wire _12896_;
wire _12897_;
wire _12898_;
wire _12899_;
wire _12900_;
wire _12901_;
wire _12902_;
wire _12903_;
wire _12904_;
wire _12905_;
wire _12906_;
wire _12907_;
wire _12908_;
wire _12909_;
wire _12910_;
wire _12911_;
wire _12912_;
wire _12913_;
wire _12914_;
wire _12915_;
wire _12916_;
wire _12917_;
wire _12918_;
wire _12919_;
wire _12920_;
wire _12921_;
wire _12922_;
wire _12923_;
wire _12924_;
wire _12925_;
wire _12926_;
wire _12927_;
wire _12928_;
wire _12929_;
wire _12930_;
wire _12931_;
wire _12932_;
wire _12933_;
wire _12934_;
wire _12935_;
wire _12936_;
wire _12937_;
wire _12938_;
wire _12939_;
wire _12940_;
wire _12941_;
wire _12942_;
wire _12943_;
wire _12944_;
wire _12945_;
wire _12946_;
wire _12947_;
wire _12948_;
wire _12949_;
wire _12950_;
wire _12951_;
wire _12952_;
wire _12953_;
wire _12954_;
wire _12955_;
wire _12956_;
wire _12957_;
wire _12958_;
wire _12959_;
wire _12960_;
wire _12961_;
wire _12962_;
wire _12963_;
wire _12964_;
wire _12965_;
wire _12966_;
wire _12967_;
wire _12968_;
wire _12969_;
wire _12970_;
wire _12971_;
wire _12972_;
wire _12973_;
wire _12974_;
wire _12975_;
wire _12976_;
wire _12977_;
wire _12978_;
wire _12979_;
wire _12980_;
wire _12981_;
wire _12982_;
wire _12983_;
wire _12984_;
wire _12985_;
wire _12986_;
wire _12987_;
wire _12988_;
wire _12989_;
wire _12990_;
wire _12991_;
wire _12992_;
wire _12993_;
wire _12994_;
wire _12995_;
wire _12996_;
wire _12997_;
wire _12998_;
wire _12999_;
wire _13000_;
wire _13001_;
wire _13002_;
wire _13003_;
wire _13004_;
wire _13005_;
wire _13006_;
wire _13007_;
wire _13008_;
wire _13009_;
wire _13010_;
wire _13011_;
wire _13012_;
wire _13013_;
wire _13014_;
wire _13015_;
wire _13016_;
wire _13017_;
wire _13018_;
wire _13019_;
wire _13020_;
wire _13021_;
wire _13022_;
wire _13023_;
wire _13024_;
wire _13025_;
wire _13026_;
wire _13027_;
wire _13028_;
wire _13029_;
wire _13030_;
wire _13031_;
wire _13032_;
wire _13033_;
wire _13034_;
wire _13035_;
wire _13036_;
wire _13037_;
wire _13038_;
wire _13039_;
wire _13040_;
wire _13041_;
wire _13042_;
wire _13043_;
wire _13044_;
wire _13045_;
wire _13046_;
wire _13047_;
wire _13048_;
wire _13049_;
wire _13050_;
wire _13051_;
wire _13052_;
wire _13053_;
wire _13054_;
wire _13055_;
wire _13056_;
wire _13057_;
wire _13058_;
wire _13059_;
wire _13060_;
wire _13061_;
wire _13062_;
wire _13063_;
wire _13064_;
wire _13065_;
wire _13066_;
wire _13067_;
wire _13068_;
wire _13069_;
wire _13070_;
wire _13071_;
wire _13072_;
wire _13073_;
wire _13074_;
wire _13075_;
wire _13076_;
wire _13077_;
wire _13078_;
wire _13079_;
wire _13080_;
wire _13081_;
wire _13082_;
wire _13083_;
wire _13084_;
wire _13085_;
wire _13086_;
wire _13087_;
wire _13088_;
wire _13089_;
wire _13090_;
wire _13091_;
wire _13092_;
wire _13093_;
wire _13094_;
wire _13095_;
wire _13096_;
wire _13097_;
wire _13098_;
wire _13099_;
wire _13100_;
wire _13101_;
wire _13102_;
wire _13103_;
wire _13104_;
wire _13105_;
wire _13106_;
wire _13107_;
wire _13108_;
wire _13109_;
wire _13110_;
wire _13111_;
wire _13112_;
wire _13113_;
wire _13114_;
wire _13115_;
wire _13116_;
wire _13117_;
wire _13118_;
wire _13119_;
wire _13120_;
wire _13121_;
wire _13122_;
wire _13123_;
wire _13124_;
wire _13125_;
wire _13126_;
wire _13127_;
wire _13128_;
wire _13129_;
wire _13130_;
wire _13131_;
wire _13132_;
wire _13133_;
wire _13134_;
wire _13135_;
wire _13136_;
wire _13137_;
wire _13138_;
wire _13139_;
wire _13140_;
wire _13141_;
wire _13142_;
wire _13143_;
wire _13144_;
wire _13145_;
wire _13146_;
wire _13147_;
wire _13148_;
wire _13149_;
wire _13150_;
wire _13151_;
wire _13152_;
wire _13153_;
wire _13154_;
wire _13155_;
wire _13156_;
wire _13157_;
wire _13158_;
wire _13159_;
wire _13160_;
wire _13161_;
wire _13162_;
wire _13163_;
wire _13164_;
wire _13165_;
wire _13166_;
wire _13167_;
wire _13168_;
wire _13169_;
wire _13170_;
wire _13171_;
wire _13172_;
wire _13173_;
wire _13174_;
wire _13175_;
wire _13176_;
wire _13177_;
wire _13178_;
wire _13179_;
wire _13180_;
wire _13181_;
wire _13182_;
wire _13183_;
wire _13184_;
wire _13185_;
wire _13186_;
wire _13187_;
wire _13188_;
wire _13189_;
wire _13190_;
wire _13191_;
wire _13192_;
wire _13193_;
wire _13194_;
wire _13195_;
wire _13196_;
wire _13197_;
wire _13198_;
wire _13199_;
wire _13200_;
wire _13201_;
wire _13202_;
wire _13203_;
wire _13204_;
wire _13205_;
wire _13206_;
wire _13207_;
wire _13208_;
wire _13209_;
wire _13210_;
wire _13211_;
wire _13212_;
wire _13213_;
wire _13214_;
wire _13215_;
wire _13216_;
wire _13217_;
wire _13218_;
wire _13219_;
wire _13220_;
wire _13221_;
wire _13222_;
wire _13223_;
wire _13224_;
wire _13225_;
wire _13226_;
wire _13227_;
wire _13228_;
wire _13229_;
wire _13230_;
wire _13231_;
wire _13232_;
wire _13233_;
wire _13234_;
wire _13235_;
wire _13236_;
wire _13237_;
wire _13238_;
wire _13239_;
wire _13240_;
wire _13241_;
wire _13242_;
wire _13243_;
wire _13244_;
wire _13245_;
wire _13246_;
wire _13247_;
wire _13248_;
wire _13249_;
wire _13250_;
wire _13251_;
wire _13252_;
wire _13253_;
wire _13254_;
wire _13255_;
wire _13256_;
wire _13257_;
wire _13258_;
wire _13259_;
wire _13260_;
wire _13261_;
wire _13262_;
wire _13263_;
wire _13264_;
wire _13265_;
wire _13266_;
wire _13267_;
wire _13268_;
wire _13269_;
wire _13270_;
wire _13271_;
wire _13272_;
wire _13273_;
wire _13274_;
wire _13275_;
wire _13276_;
wire _13277_;
wire _13278_;
wire _13279_;
wire _13280_;
wire _13281_;
wire _13282_;
wire _13283_;
wire _13284_;
wire _13285_;
wire _13286_;
wire _13287_;
wire _13288_;
wire _13289_;
wire _13290_;
wire _13291_;
wire _13292_;
wire _13293_;
wire _13294_;
wire _13295_;
wire _13296_;
wire _13297_;
wire _13298_;
wire _13299_;
wire _13300_;
wire _13301_;
wire _13302_;
wire _13303_;
wire _13304_;
wire _13305_;
wire _13306_;
wire _13307_;
wire _13308_;
wire _13309_;
wire _13310_;
wire _13311_;
wire _13312_;
wire _13313_;
wire _13314_;
wire _13315_;
wire _13316_;
wire _13317_;
wire _13318_;
wire _13319_;
wire _13320_;
wire _13321_;
wire _13322_;
wire _13323_;
wire _13324_;
wire _13325_;
wire _13326_;
wire _13327_;
wire _13328_;
wire _13329_;
wire _13330_;
wire _13331_;
wire _13332_;
wire _13333_;
wire _13334_;
wire _13335_;
wire _13336_;
wire _13337_;
wire _13338_;
wire _13339_;
wire _13340_;
wire _13341_;
wire _13342_;
wire _13343_;
wire _13344_;
wire _13345_;
wire _13346_;
wire _13347_;
wire _13348_;
wire _13349_;
wire _13350_;
wire _13351_;
wire _13352_;
wire _13353_;
wire _13354_;
wire _13355_;
wire _13356_;
wire _13357_;
wire _13358_;
wire _13359_;
wire _13360_;
wire _13361_;
wire _13362_;
wire _13363_;
wire _13364_;
wire _13365_;
wire _13366_;
wire _13367_;
wire _13368_;
wire _13369_;
wire _13370_;
wire _13371_;
wire _13372_;
wire _13373_;
wire _13374_;
wire _13375_;
wire _13376_;
wire _13377_;
wire _13378_;
wire _13379_;
wire _13380_;
wire _13381_;
wire _13382_;
wire _13383_;
wire _13384_;
wire _13385_;
wire _13386_;
wire _13387_;
wire _13388_;
wire _13389_;
wire _13390_;
wire _13391_;
wire _13392_;
wire _13393_;
wire _13394_;
wire _13395_;
wire _13396_;
wire _13397_;
wire _13398_;
wire _13399_;
wire _13400_;
wire _13401_;
wire _13402_;
wire _13403_;
wire _13404_;
wire _13405_;
wire _13406_;
wire _13407_;
wire _13408_;
wire _13409_;
wire _13410_;
wire _13411_;
wire _13412_;
wire _13413_;
wire _13414_;
wire _13415_;
wire _13416_;
wire _13417_;
wire _13418_;
wire _13419_;
wire _13420_;
wire _13421_;
wire _13422_;
wire _13423_;
wire _13424_;
wire _13425_;
wire _13426_;
wire _13427_;
wire _13428_;
wire _13429_;
wire _13430_;
wire _13431_;
wire _13432_;
wire _13433_;
wire _13434_;
wire _13435_;
wire _13436_;
wire _13437_;
wire _13438_;
wire _13439_;
wire _13440_;
wire _13441_;
wire _13442_;
wire _13443_;
wire _13444_;
wire _13445_;
wire _13446_;
wire _13447_;
wire _13448_;
wire _13449_;
wire _13450_;
wire _13451_;
wire _13452_;
wire _13453_;
wire _13454_;
wire _13455_;
wire _13456_;
wire _13457_;
wire _13458_;
wire _13459_;
wire _13460_;
wire _13461_;
wire _13462_;
wire _13463_;
wire _13464_;
wire _13465_;
wire _13466_;
wire _13467_;
wire _13468_;
wire _13469_;
wire _13470_;
wire _13471_;
wire _13472_;
wire _13473_;
wire _13474_;
wire _13475_;
wire _13476_;
wire _13477_;
wire _13478_;
wire _13479_;
wire _13480_;
wire _13481_;
wire _13482_;
wire _13483_;
wire _13484_;
wire _13485_;
wire _13486_;
wire _13487_;
wire _13488_;
wire _13489_;
wire _13490_;
wire _13491_;
wire _13492_;
wire _13493_;
wire _13494_;
wire _13495_;
wire _13496_;
wire _13497_;
wire _13498_;
wire _13499_;
wire _13500_;
wire _13501_;
wire _13502_;
wire _13503_;
wire _13504_;
wire _13505_;
wire _13506_;
wire _13507_;
wire _13508_;
wire _13509_;
wire _13510_;
wire _13511_;
wire _13512_;
wire _13513_;
wire _13514_;
wire _13515_;
wire _13516_;
wire _13517_;
wire _13518_;
wire _13519_;
wire _13520_;
wire _13521_;
wire _13522_;
wire _13523_;
wire _13524_;
wire _13525_;
wire _13526_;
wire _13527_;
wire _13528_;
wire _13529_;
wire _13530_;
wire _13531_;
wire _13532_;
wire _13533_;
wire _13534_;
wire _13535_;
wire _13536_;
wire _13537_;
wire _13538_;
wire _13539_;
wire _13540_;
wire _13541_;
wire _13542_;
wire _13543_;
wire _13544_;
wire _13545_;
wire _13546_;
wire _13547_;
wire _13548_;
wire _13549_;
wire _13550_;
wire _13551_;
wire _13552_;
wire _13553_;
wire _13554_;
wire _13555_;
wire _13556_;
wire _13557_;
wire _13558_;
wire _13559_;
wire _13560_;
wire _13561_;
wire _13562_;
wire _13563_;
wire _13564_;
wire _13565_;
wire _13566_;
wire _13567_;
wire _13568_;
wire _13569_;
wire _13570_;
wire _13571_;
wire _13572_;
wire _13573_;
wire _13574_;
wire _13575_;
wire _13576_;
wire _13577_;
wire _13578_;
wire _13579_;
wire _13580_;
wire _13581_;
wire _13582_;
wire _13583_;
wire _13584_;
wire _13585_;
wire _13586_;
wire _13587_;
wire _13588_;
wire _13589_;
wire _13590_;
wire _13591_;
wire _13592_;
wire _13593_;
wire _13594_;
wire _13595_;
wire _13596_;
wire _13597_;
wire _13598_;
wire _13599_;
wire _13600_;
wire _13601_;
wire _13602_;
wire _13603_;
wire _13604_;
wire _13605_;
wire _13606_;
wire _13607_;
wire _13608_;
wire _13609_;
wire _13610_;
wire _13611_;
wire _13612_;
wire _13613_;
wire _13614_;
wire _13615_;
wire _13616_;
wire _13617_;
wire _13618_;
wire _13619_;
wire _13620_;
wire _13621_;
wire _13622_;
wire _13623_;
wire _13624_;
wire _13625_;
wire _13626_;
wire _13627_;
wire _13628_;
wire _13629_;
wire _13630_;
wire _13631_;
wire _13632_;
wire _13633_;
wire _13634_;
wire _13635_;
wire _13636_;
wire _13637_;
wire _13638_;
wire _13639_;
wire _13640_;
wire _13641_;
wire _13642_;
wire _13643_;
wire _13644_;
wire _13645_;
wire _13646_;
wire _13647_;
wire _13648_;
wire _13649_;
wire _13650_;
wire _13651_;
wire _13652_;
wire _13653_;
wire _13654_;
wire _13655_;
wire _13656_;
wire _13657_;
wire _13658_;
wire _13659_;
wire _13660_;
wire _13661_;
wire _13662_;
wire _13663_;
wire _13664_;
wire _13665_;
wire _13666_;
wire _13667_;
wire _13668_;
wire _13669_;
wire _13670_;
wire _13671_;
wire _13672_;
wire _13673_;
wire _13674_;
wire _13675_;
wire _13676_;
wire _13677_;
wire _13678_;
wire _13679_;
wire _13680_;
wire _13681_;
wire _13682_;
wire _13683_;
wire _13684_;
wire _13685_;
wire _13686_;
wire _13687_;
wire _13688_;
wire _13689_;
wire _13690_;
wire _13691_;
wire _13692_;
wire _13693_;
wire _13694_;
wire _13695_;
wire _13696_;
wire _13697_;
wire _13698_;
wire _13699_;
wire _13700_;
wire _13701_;
wire _13702_;
wire _13703_;
wire _13704_;
wire _13705_;
wire _13706_;
wire _13707_;
wire _13708_;
wire _13709_;
wire _13710_;
wire _13711_;
wire _13712_;
wire _13713_;
wire _13714_;
wire _13715_;
wire _13716_;
wire _13717_;
wire _13718_;
wire _13719_;
wire _13720_;
wire _13721_;
wire _13722_;
wire _13723_;
wire _13724_;
wire _13725_;
wire _13726_;
wire _13727_;
wire _13728_;
wire _13729_;
wire _13730_;
wire _13731_;
wire _13732_;
wire _13733_;
wire _13734_;
wire _13735_;
wire _13736_;
wire _13737_;
wire _13738_;
wire _13739_;
wire _13740_;
wire _13741_;
wire _13742_;
wire _13743_;
wire _13744_;
wire _13745_;
wire _13746_;
wire _13747_;
wire _13748_;
wire _13749_;
wire _13750_;
wire _13751_;
wire _13752_;
wire _13753_;
wire _13754_;
wire _13755_;
wire _13756_;
wire _13757_;
wire _13758_;
wire _13759_;
wire _13760_;
wire _13761_;
wire _13762_;
wire _13763_;
wire _13764_;
wire _13765_;
wire _13766_;
wire _13767_;
wire _13768_;
wire _13769_;
wire _13770_;
wire _13771_;
wire _13772_;
wire _13773_;
wire _13774_;
wire _13775_;
wire _13776_;
wire _13777_;
wire _13778_;
wire _13779_;
wire _13780_;
wire _13781_;
wire _13782_;
wire _13783_;
wire _13784_;
wire _13785_;
wire _13786_;
wire _13787_;
wire _13788_;
wire _13789_;
wire _13790_;
wire _13791_;
wire _13792_;
wire _13793_;
wire _13794_;
wire _13795_;
wire _13796_;
wire _13797_;
wire _13798_;
wire _13799_;
wire _13800_;
wire _13801_;
wire _13802_;
wire _13803_;
wire _13804_;
wire _13805_;
wire _13806_;
wire _13807_;
wire _13808_;
wire _13809_;
wire _13810_;
wire _13811_;
wire _13812_;
wire _13813_;
wire _13814_;
wire _13815_;
wire _13816_;
wire _13817_;
wire _13818_;
wire _13819_;
wire _13820_;
wire _13821_;
wire _13822_;
wire _13823_;
wire _13824_;
wire _13825_;
wire _13826_;
wire _13827_;
wire _13828_;
wire _13829_;
wire _13830_;
wire _13831_;
wire _13832_;
wire _13833_;
wire _13834_;
wire _13835_;
wire _13836_;
wire _13837_;
wire _13838_;
wire _13839_;
wire _13840_;
wire _13841_;
wire _13842_;
wire _13843_;
wire _13844_;
wire _13845_;
wire _13846_;
wire _13847_;
wire _13848_;
wire _13849_;
wire _13850_;
wire _13851_;
wire _13852_;
wire _13853_;
wire _13854_;
wire _13855_;
wire _13856_;
wire _13857_;
wire _13858_;
wire _13859_;
wire _13860_;
wire _13861_;
wire _13862_;
wire _13863_;
wire _13864_;
wire _13865_;
wire _13866_;
wire _13867_;
wire _13868_;
wire _13869_;
wire _13870_;
wire _13871_;
wire _13872_;
wire _13873_;
wire _13874_;
wire _13875_;
wire _13876_;
wire _13877_;
wire _13878_;
wire _13879_;
wire _13880_;
wire _13881_;
wire _13882_;
wire _13883_;
wire _13884_;
wire _13885_;
wire _13886_;
wire _13887_;
wire _13888_;
wire _13889_;
wire _13890_;
wire _13891_;
wire _13892_;
wire _13893_;
wire _13894_;
wire _13895_;
wire _13896_;
wire _13897_;
wire _13898_;
wire _13899_;
wire _13900_;
wire _13901_;
wire _13902_;
wire _13903_;
wire _13904_;
wire _13905_;
wire _13906_;
wire _13907_;
wire _13908_;
wire _13909_;
wire _13910_;
wire _13911_;
wire _13912_;
wire _13913_;
wire _13914_;
wire _13915_;
wire _13916_;
wire _13917_;
wire _13918_;
wire _13919_;
wire _13920_;
wire _13921_;
wire _13922_;
wire _13923_;
wire _13924_;
wire _13925_;
wire _13926_;
wire _13927_;
wire _13928_;
wire _13929_;
wire _13930_;
wire _13931_;
wire _13932_;
wire _13933_;
wire _13934_;
wire _13935_;
wire _13936_;
wire _13937_;
wire _13938_;
wire _13939_;
wire _13940_;
wire _13941_;
wire _13942_;
wire _13943_;
wire _13944_;
wire _13945_;
wire _13946_;
wire _13947_;
wire _13948_;
wire _13949_;
wire _13950_;
wire _13951_;
wire _13952_;
wire _13953_;
wire _13954_;
wire _13955_;
wire _13956_;
wire _13957_;
wire _13958_;
wire _13959_;
wire _13960_;
wire _13961_;
wire _13962_;
wire _13963_;
wire _13964_;
wire _13965_;
wire _13966_;
wire _13967_;
wire _13968_;
wire _13969_;
wire _13970_;
wire _13971_;
wire _13972_;
wire _13973_;
wire _13974_;
wire _13975_;
wire _13976_;
wire _13977_;
wire _13978_;
wire _13979_;
wire _13980_;
wire _13981_;
wire _13982_;
wire _13983_;
wire _13984_;
wire _13985_;
wire _13986_;
wire _13987_;
wire _13988_;
wire _13989_;
wire _13990_;
wire _13991_;
wire _13992_;
wire _13993_;
wire _13994_;
wire _13995_;
wire _13996_;
wire _13997_;
wire _13998_;
wire _13999_;
wire _14000_;
wire _14001_;
wire _14002_;
wire _14003_;
wire _14004_;
wire _14005_;
wire _14006_;
wire _14007_;
wire _14008_;
wire _14009_;
wire _14010_;
wire _14011_;
wire _14012_;
wire _14013_;
wire _14014_;
wire _14015_;
wire _14016_;
wire _14017_;
wire _14018_;
wire _14019_;
wire _14020_;
wire _14021_;
wire _14022_;
wire _14023_;
wire _14024_;
wire _14025_;
wire _14026_;
wire _14027_;
wire _14028_;
wire _14029_;
wire _14030_;
wire _14031_;
wire _14032_;
wire _14033_;
wire _14034_;
wire _14035_;
wire _14036_;
wire _14037_;
wire _14038_;
wire _14039_;
wire _14040_;
wire _14041_;
wire _14042_;
wire _14043_;
wire _14044_;
wire _14045_;
wire _14046_;
wire _14047_;
wire _14048_;
wire _14049_;
wire _14050_;
wire _14051_;
wire _14052_;
wire _14053_;
wire _14054_;
wire _14055_;
wire _14056_;
wire _14057_;
wire _14058_;
wire _14059_;
wire _14060_;
wire _14061_;
wire _14062_;
wire _14063_;
wire _14064_;
wire _14065_;
wire _14066_;
wire _14067_;
wire _14068_;
wire _14069_;
wire _14070_;
wire _14071_;
wire _14072_;
wire _14073_;
wire _14074_;
wire _14075_;
wire _14076_;
wire _14077_;
wire _14078_;
wire _14079_;
wire _14080_;
wire _14081_;
wire _14082_;
wire _14083_;
wire _14084_;
wire _14085_;
wire _14086_;
wire _14087_;
wire _14088_;
wire _14089_;
wire _14090_;
wire _14091_;
wire _14092_;
wire _14093_;
wire _14094_;
wire _14095_;
wire _14096_;
wire _14097_;
wire _14098_;
wire _14099_;
wire _14100_;
wire _14101_;
wire _14102_;
wire _14103_;
wire _14104_;
wire _14105_;
wire _14106_;
wire _14107_;
wire _14108_;
wire _14109_;
wire _14110_;
wire _14111_;
wire _14112_;
wire _14113_;
wire _14114_;
wire _14115_;
wire _14116_;
wire _14117_;
wire _14118_;
wire _14119_;
wire _14120_;
wire _14121_;
wire _14122_;
wire _14123_;
wire _14124_;
wire _14125_;
wire _14126_;
wire _14127_;
wire _14128_;
wire _14129_;
wire _14130_;
wire _14131_;
wire _14132_;
wire _14133_;
wire _14134_;
wire _14135_;
wire _14136_;
wire _14137_;
wire _14138_;
wire _14139_;
wire _14140_;
wire _14141_;
wire _14142_;
wire _14143_;
wire _14144_;
wire _14145_;
wire _14146_;
wire _14147_;
wire _14148_;
wire _14149_;
wire _14150_;
wire _14151_;
wire _14152_;
wire _14153_;
wire _14154_;
wire _14155_;
wire _14156_;
wire _14157_;
wire _14158_;
wire _14159_;
wire _14160_;
wire _14161_;
wire _14162_;
wire _14163_;
wire _14164_;
wire _14165_;
wire _14166_;
wire _14167_;
wire _14168_;
wire _14169_;
wire _14170_;
wire _14171_;
wire _14172_;
wire _14173_;
wire _14174_;
wire _14175_;
wire _14176_;
wire _14177_;
wire _14178_;
wire _14179_;
wire _14180_;
wire _14181_;
wire _14182_;
wire _14183_;
wire _14184_;
wire _14185_;
wire _14186_;
wire _14187_;
wire _14188_;
wire _14189_;
wire _14190_;
wire _14191_;
wire _14192_;
wire _14193_;
wire _14194_;
wire _14195_;
wire _14196_;
wire _14197_;
wire _14198_;
wire _14199_;
wire _14200_;
wire _14201_;
wire _14202_;
wire _14203_;
wire _14204_;
wire _14205_;
wire _14206_;
wire _14207_;
wire _14208_;
wire _14209_;
wire _14210_;
wire _14211_;
wire _14212_;
wire _14213_;
wire _14214_;
wire _14215_;
wire _14216_;
wire _14217_;
wire _14218_;
wire _14219_;
wire _14220_;
wire _14221_;
wire _14222_;
wire _14223_;
wire _14224_;
wire _14225_;
wire _14226_;
wire _14227_;
wire _14228_;
wire _14229_;
wire _14230_;
wire _14231_;
wire _14232_;
wire _14233_;
wire _14234_;
wire _14235_;
wire _14236_;
wire _14237_;
wire _14238_;
wire _14239_;
wire _14240_;
wire _14241_;
wire _14242_;
wire _14243_;
wire _14244_;
wire _14245_;
wire _14246_;
wire _14247_;
wire _14248_;
wire _14249_;
wire _14250_;
wire _14251_;
wire _14252_;
wire _14253_;
wire _14254_;
wire _14255_;
wire _14256_;
wire _14257_;
wire _14258_;
wire _14259_;
wire _14260_;
wire _14261_;
wire _14262_;
wire _14263_;
wire _14264_;
wire _14265_;
wire _14266_;
wire _14267_;
wire _14268_;
wire _14269_;
wire _14270_;
wire _14271_;
wire _14272_;
wire _14273_;
wire _14274_;
wire _14275_;
wire _14276_;
wire _14277_;
wire _14278_;
wire _14279_;
wire _14280_;
wire _14281_;
wire _14282_;
wire _14283_;
wire _14284_;
wire _14285_;
wire _14286_;
wire _14287_;
wire _14288_;
wire _14289_;
wire _14290_;
wire _14291_;
wire _14292_;
wire _14293_;
wire _14294_;
wire _14295_;
wire _14296_;
wire _14297_;
wire _14298_;
wire _14299_;
wire _14300_;
wire _14301_;
wire _14302_;
wire _14303_;
wire _14304_;
wire _14305_;
wire _14306_;
wire _14307_;
wire _14308_;
wire _14309_;
wire _14310_;
wire _14311_;
wire _14312_;
wire _14313_;
wire _14314_;
wire _14315_;
wire _14316_;
wire _14317_;
wire _14318_;
wire _14319_;
wire _14320_;
wire _14321_;
wire _14322_;
wire _14323_;
wire _14324_;
wire _14325_;
wire _14326_;
wire _14327_;
wire _14328_;
wire _14329_;
wire _14330_;
wire _14331_;
wire _14332_;
wire _14333_;
wire _14334_;
wire _14335_;
wire _14336_;
wire _14337_;
wire _14338_;
wire _14339_;
wire _14340_;
wire _14341_;
wire _14342_;
wire _14343_;
wire _14344_;
wire _14345_;
wire _14346_;
wire _14347_;
wire _14348_;
wire _14349_;
wire _14350_;
wire _14351_;
wire _14352_;
wire _14353_;
wire _14354_;
wire _14355_;
wire _14356_;
wire _14357_;
wire _14358_;
wire _14359_;
wire _14360_;
wire _14361_;
wire _14362_;
wire _14363_;
wire _14364_;
wire _14365_;
wire _14366_;
wire _14367_;
wire _14368_;
wire _14369_;
wire _14370_;
wire _14371_;
wire _14372_;
wire _14373_;
wire _14374_;
wire _14375_;
wire _14376_;
wire _14377_;
wire _14378_;
wire _14379_;
wire _14380_;
wire _14381_;
wire _14382_;
wire _14383_;
wire _14384_;
wire _14385_;
wire _14386_;
wire _14387_;
wire _14388_;
wire _14389_;
wire _14390_;
wire _14391_;
wire _14392_;
wire _14393_;
wire _14394_;
wire _14395_;
wire _14396_;
wire _14397_;
wire _14398_;
wire _14399_;
wire _14400_;
wire _14401_;
wire _14402_;
wire _14403_;
wire _14404_;
wire _14405_;
wire _14406_;
wire _14407_;
wire _14408_;
wire _14409_;
wire _14410_;
wire _14411_;
wire _14412_;
wire _14413_;
wire _14414_;
wire _14415_;
wire _14416_;
wire _14417_;
wire _14418_;
wire _14419_;
wire _14420_;
wire _14421_;
wire _14422_;
wire _14423_;
wire _14424_;
wire _14425_;
wire _14426_;
wire _14427_;
wire _14428_;
wire _14429_;
wire _14430_;
wire _14431_;
wire _14432_;
wire _14433_;
wire _14434_;
wire _14435_;
wire _14436_;
wire _14437_;
wire _14438_;
wire _14439_;
wire _14440_;
wire _14441_;
wire _14442_;
wire _14443_;
wire _14444_;
wire _14445_;
wire _14446_;
wire _14447_;
wire _14448_;
wire _14449_;
wire _14450_;
wire _14451_;
wire _14452_;
wire _14453_;
wire _14454_;
wire _14455_;
wire _14456_;
wire _14457_;
wire _14458_;
wire _14459_;
wire _14460_;
wire _14461_;
wire _14462_;
wire _14463_;
wire _14464_;
wire _14465_;
wire _14466_;
wire _14467_;
wire _14468_;
wire _14469_;
wire _14470_;
wire _14471_;
wire _14472_;
wire _14473_;
wire _14474_;
wire _14475_;
wire _14476_;
wire _14477_;
wire _14478_;
wire _14479_;
wire _14480_;
wire _14481_;
wire _14482_;
wire _14483_;
wire _14484_;
wire _14485_;
wire _14486_;
wire _14487_;
wire _14488_;
wire _14489_;
wire _14490_;
wire _14491_;
wire _14492_;
wire _14493_;
wire _14494_;
wire _14495_;
wire _14496_;
wire _14497_;
wire _14498_;
wire _14499_;
wire _14500_;
wire _14501_;
wire _14502_;
wire _14503_;
wire _14504_;
wire _14505_;
wire _14506_;
wire _14507_;
wire _14508_;
wire _14509_;
wire _14510_;
wire _14511_;
wire _14512_;
wire _14513_;
wire _14514_;
wire _14515_;
wire _14516_;
wire _14517_;
wire _14518_;
wire _14519_;
wire _14520_;
wire _14521_;
wire _14522_;
wire _14523_;
wire _14524_;
wire _14525_;
wire _14526_;
wire _14527_;
wire _14528_;
wire _14529_;
wire _14530_;
wire _14531_;
wire _14532_;
wire _14533_;
wire _14534_;
wire _14535_;
wire _14536_;
wire _14537_;
wire _14538_;
wire _14539_;
wire _14540_;
wire _14541_;
wire _14542_;
wire _14543_;
wire _14544_;
wire _14545_;
wire _14546_;
wire _14547_;
wire _14548_;
wire _14549_;
wire _14550_;
wire _14551_;
wire _14552_;
wire _14553_;
wire _14554_;
wire _14555_;
wire _14556_;
wire _14557_;
wire _14558_;
wire _14559_;
wire _14560_;
wire _14561_;
wire _14562_;
wire _14563_;
wire _14564_;
wire _14565_;
wire _14566_;
wire _14567_;
wire _14568_;
wire _14569_;
wire _14570_;
wire _14571_;
wire _14572_;
wire _14573_;
wire _14574_;
wire _14575_;
wire _14576_;
wire _14577_;
wire _14578_;
wire _14579_;
wire _14580_;
wire _14581_;
wire _14582_;
wire _14583_;
wire _14584_;
wire _14585_;
wire _14586_;
wire _14587_;
wire _14588_;
wire _14589_;
wire _14590_;
wire _14591_;
wire _14592_;
wire _14593_;
wire _14594_;
wire _14595_;
wire _14596_;
wire _14597_;
wire _14598_;
wire _14599_;
wire _14600_;
wire _14601_;
wire _14602_;
wire _14603_;
wire _14604_;
wire _14605_;
wire _14606_;
wire _14607_;
wire _14608_;
wire _14609_;
wire _14610_;
wire _14611_;
wire _14612_;
wire _14613_;
wire _14614_;
wire _14615_;
wire _14616_;
wire _14617_;
wire _14618_;
wire _14619_;
wire _14620_;
wire _14621_;
wire _14622_;
wire _14623_;
wire _14624_;
wire _14625_;
wire _14626_;
wire _14627_;
wire _14628_;
wire _14629_;
wire _14630_;
wire _14631_;
wire _14632_;
wire _14633_;
wire _14634_;
wire _14635_;
wire _14636_;
wire _14637_;
wire _14638_;
wire _14639_;
wire _14640_;
wire _14641_;
wire _14642_;
wire _14643_;
wire _14644_;
wire _14645_;
wire _14646_;
wire _14647_;
wire _14648_;
wire _14649_;
wire _14650_;
wire _14651_;
wire _14652_;
wire _14653_;
wire _14654_;
wire _14655_;
wire _14656_;
wire _14657_;
wire _14658_;
wire _14659_;
wire _14660_;
wire _14661_;
wire _14662_;
wire _14663_;
wire _14664_;
wire _14665_;
wire _14666_;
wire _14667_;
wire _14668_;
wire _14669_;
wire _14670_;
wire _14671_;
wire _14672_;
wire _14673_;
wire _14674_;
wire _14675_;
wire _14676_;
wire _14677_;
wire _14678_;
wire _14679_;
wire _14680_;
wire _14681_;
wire _14682_;
wire _14683_;
wire _14684_;
wire _14685_;
wire _14686_;
wire _14687_;
wire _14688_;
wire _14689_;
wire _14690_;
wire _14691_;
wire _14692_;
wire _14693_;
wire _14694_;
wire _14695_;
wire _14696_;
wire _14697_;
wire _14698_;
wire _14699_;
wire _14700_;
wire _14701_;
wire _14702_;
wire _14703_;
wire _14704_;
wire _14705_;
wire _14706_;
wire _14707_;
wire _14708_;
wire _14709_;
wire _14710_;
wire _14711_;
wire _14712_;
wire _14713_;
wire _14714_;
wire _14715_;
wire _14716_;
wire _14717_;
wire _14718_;
wire _14719_;
wire _14720_;
wire _14721_;
wire _14722_;
wire _14723_;
wire _14724_;
wire _14725_;
wire _14726_;
wire _14727_;
wire _14728_;
wire _14729_;
wire _14730_;
wire _14731_;
wire _14732_;
wire _14733_;
wire _14734_;
wire _14735_;
wire _14736_;
wire _14737_;
wire _14738_;
wire _14739_;
wire _14740_;
wire _14741_;
wire _14742_;
wire _14743_;
wire _14744_;
wire _14745_;
wire _14746_;
wire _14747_;
wire _14748_;
wire _14749_;
wire _14750_;
wire _14751_;
wire _14752_;
wire _14753_;
wire _14754_;
wire _14755_;
wire _14756_;
wire _14757_;
wire _14758_;
wire _14759_;
wire _14760_;
wire _14761_;
wire _14762_;
wire _14763_;
wire _14764_;
wire _14765_;
wire _14766_;
wire _14767_;
wire _14768_;
wire _14769_;
wire _14770_;
wire _14771_;
wire _14772_;
wire _14773_;
wire _14774_;
wire _14775_;
wire _14776_;
wire _14777_;
wire _14778_;
wire _14779_;
wire _14780_;
wire _14781_;
wire _14782_;
wire _14783_;
wire _14784_;
wire _14785_;
wire _14786_;
wire _14787_;
wire _14788_;
wire _14789_;
wire _14790_;
wire _14791_;
wire _14792_;
wire _14793_;
wire _14794_;
wire _14795_;
wire _14796_;
wire _14797_;
wire _14798_;
wire _14799_;
wire _14800_;
wire _14801_;
wire _14802_;
wire _14803_;
wire _14804_;
wire _14805_;
wire _14806_;
wire _14807_;
wire _14808_;
wire _14809_;
wire _14810_;
wire _14811_;
wire _14812_;
wire _14813_;
wire _14814_;
wire _14815_;
wire _14816_;
wire _14817_;
wire _14818_;
wire _14819_;
wire _14820_;
wire _14821_;
wire _14822_;
wire _14823_;
wire _14824_;
wire _14825_;
wire _14826_;
wire _14827_;
wire _14828_;
wire _14829_;
wire _14830_;
wire _14831_;
wire _14832_;
wire _14833_;
wire _14834_;
wire _14835_;
wire _14836_;
wire _14837_;
wire _14838_;
wire _14839_;
wire _14840_;
wire _14841_;
wire _14842_;
wire _14843_;
wire _14844_;
wire _14845_;
wire _14846_;
wire _14847_;
wire _14848_;
wire _14849_;
wire _14850_;
wire _14851_;
wire _14852_;
wire _14853_;
wire _14854_;
wire _14855_;
wire _14856_;
wire _14857_;
wire _14858_;
wire _14859_;
wire _14860_;
wire _14861_;
wire _14862_;
wire _14863_;
wire _14864_;
wire _14865_;
wire _14866_;
wire _14867_;
wire _14868_;
wire _14869_;
wire _14870_;
wire _14871_;
wire _14872_;
wire _14873_;
wire _14874_;
wire _14875_;
wire _14876_;
wire _14877_;
wire _14878_;
wire _14879_;
wire _14880_;
wire _14881_;
wire _14882_;
wire _14883_;
wire _14884_;
wire _14885_;
wire _14886_;
wire _14887_;
wire _14888_;
wire _14889_;
wire _14890_;
wire _14891_;
wire _14892_;
wire _14893_;
wire _14894_;
wire _14895_;
wire _14896_;
wire _14897_;
wire _14898_;
wire _14899_;
wire _14900_;
wire _14901_;
wire _14902_;
wire _14903_;
wire _14904_;
wire _14905_;
wire _14906_;
wire _14907_;
wire _14908_;
wire _14909_;
wire _14910_;
wire _14911_;
wire _14912_;
wire _14913_;
wire _14914_;
wire _14915_;
wire _14916_;
wire _14917_;
wire _14918_;
wire _14919_;
wire _14920_;
wire _14921_;
wire _14922_;
wire _14923_;
wire _14924_;
wire _14925_;
wire _14926_;
wire _14927_;
wire _14928_;
wire _14929_;
wire _14930_;
wire _14931_;
wire _14932_;
wire _14933_;
wire _14934_;
wire _14935_;
wire _14936_;
wire _14937_;
wire _14938_;
wire _14939_;
wire _14940_;
wire _14941_;
wire _14942_;
wire _14943_;
wire _14944_;
wire _14945_;
wire _14946_;
wire _14947_;
wire _14948_;
wire _14949_;
wire _14950_;
wire _14951_;
wire _14952_;
wire _14953_;
wire _14954_;
wire _14955_;
wire _14956_;
wire _14957_;
wire _14958_;
wire _14959_;
wire _14960_;
wire _14961_;
wire _14962_;
wire _14963_;
wire _14964_;
wire _14965_;
wire _14966_;
wire _14967_;
wire _14968_;
wire _14969_;
wire _14970_;
wire _14971_;
wire _14972_;
wire _14973_;
wire _14974_;
wire _14975_;
wire _14976_;
wire _14977_;
wire _14978_;
wire _14979_;
wire _14980_;
wire _14981_;
wire _14982_;
wire _14983_;
wire _14984_;
wire _14985_;
wire _14986_;
wire _14987_;
wire _14988_;
wire _14989_;
wire _14990_;
wire _14991_;
wire _14992_;
wire _14993_;
wire _14994_;
wire _14995_;
wire _14996_;
wire _14997_;
wire _14998_;
wire _14999_;
wire _15000_;
wire _15001_;
wire _15002_;
wire _15003_;
wire _15004_;
wire _15005_;
wire _15006_;
wire _15007_;
wire _15008_;
wire _15009_;
wire _15010_;
wire _15011_;
wire _15012_;
wire _15013_;
wire _15014_;
wire _15015_;
wire _15016_;
wire _15017_;
wire _15018_;
wire _15019_;
wire _15020_;
wire _15021_;
wire _15022_;
wire _15023_;
wire _15024_;
wire _15025_;
wire _15026_;
wire _15027_;
wire _15028_;
wire _15029_;
wire _15030_;
wire _15031_;
wire _15032_;
wire _15033_;
wire _15034_;
wire _15035_;
wire _15036_;
wire _15037_;
wire _15038_;
wire _15039_;
wire _15040_;
wire _15041_;
wire _15042_;
wire _15043_;
wire _15044_;
wire _15045_;
wire _15046_;
wire _15047_;
wire _15048_;
wire _15049_;
wire _15050_;
wire _15051_;
wire _15052_;
wire _15053_;
wire _15054_;
wire _15055_;
wire _15056_;
wire _15057_;
wire _15058_;
wire _15059_;
wire _15060_;
wire _15061_;
wire _15062_;
wire _15063_;
wire _15064_;
wire _15065_;
wire _15066_;
wire _15067_;
wire _15068_;
wire _15069_;
wire _15070_;
wire _15071_;
wire _15072_;
wire _15073_;
wire _15074_;
wire _15075_;
wire _15076_;
wire _15077_;
wire _15078_;
wire _15079_;
wire _15080_;
wire _15081_;
wire _15082_;
wire _15083_;
wire _15084_;
wire _15085_;
wire _15086_;
wire _15087_;
wire _15088_;
wire _15089_;
wire _15090_;
wire _15091_;
wire _15092_;
wire _15093_;
wire _15094_;
wire _15095_;
wire _15096_;
wire _15097_;
wire _15098_;
wire _15099_;
wire _15100_;
wire _15101_;
wire _15102_;
wire _15103_;
wire _15104_;
wire _15105_;
wire _15106_;
wire _15107_;
wire _15108_;
wire _15109_;
wire _15110_;
wire _15111_;
wire _15112_;
wire _15113_;
wire _15114_;
wire _15115_;
wire _15116_;
wire _15117_;
wire _15118_;
wire _15119_;
wire _15120_;
wire _15121_;
wire _15122_;
wire _15123_;
wire _15124_;
wire _15125_;
wire _15126_;
wire _15127_;
wire _15128_;
wire _15129_;
wire _15130_;
wire _15131_;
wire _15132_;
wire _15133_;
wire _15134_;
wire _15135_;
wire _15136_;
wire _15137_;
wire _15138_;
wire _15139_;
wire _15140_;
wire _15141_;
wire _15142_;
wire _15143_;
wire _15144_;
wire _15145_;
wire _15146_;
wire _15147_;
wire _15148_;
wire _15149_;
wire _15150_;
wire _15151_;
wire _15152_;
wire _15153_;
wire _15154_;
wire _15155_;
wire _15156_;
wire _15157_;
wire _15158_;
wire _15159_;
wire _15160_;
wire _15161_;
wire _15162_;
wire _15163_;
wire _15164_;
wire _15165_;
wire _15166_;
wire _15167_;
wire _15168_;
wire _15169_;
wire _15170_;
wire _15171_;
wire _15172_;
wire _15173_;
wire _15174_;
wire _15175_;
wire _15176_;
wire _15177_;
wire _15178_;
wire _15179_;
wire _15180_;
wire _15181_;
wire _15182_;
wire _15183_;
wire _15184_;
wire _15185_;
wire _15186_;
wire _15187_;
wire _15188_;
wire _15189_;
wire _15190_;
wire _15191_;
wire _15192_;
wire _15193_;
wire _15194_;
wire _15195_;
wire _15196_;
wire _15197_;
wire _15198_;
wire _15199_;
wire _15200_;
wire _15201_;
wire _15202_;
wire _15203_;
wire _15204_;
wire _15205_;
wire _15206_;
wire _15207_;
wire _15208_;
wire _15209_;
wire _15210_;
wire _15211_;
wire _15212_;
wire _15213_;
wire _15214_;
wire _15215_;
wire _15216_;
wire _15217_;
wire _15218_;
wire _15219_;
wire _15220_;
wire _15221_;
wire _15222_;
wire _15223_;
wire _15224_;
wire _15225_;
wire _15226_;
wire _15227_;
wire _15228_;
wire _15229_;
wire _15230_;
wire _15231_;
wire _15232_;
wire _15233_;
wire _15234_;
wire _15235_;
wire _15236_;
wire _15237_;
wire _15238_;
wire _15239_;
wire _15240_;
wire _15241_;
wire _15242_;
wire _15243_;
wire _15244_;
wire _15245_;
wire _15246_;
wire _15247_;
wire _15248_;
wire _15249_;
wire _15250_;
wire _15251_;
wire _15252_;
wire _15253_;
wire _15254_;
wire _15255_;
wire _15256_;
wire _15257_;
wire _15258_;
wire _15259_;
wire _15260_;
wire _15261_;
wire _15262_;
wire _15263_;
wire _15264_;
wire _15265_;
wire _15266_;
wire _15267_;
wire _15268_;
wire _15269_;
wire _15270_;
wire _15271_;
wire _15272_;
wire _15273_;
wire _15274_;
wire _15275_;
wire _15276_;
wire _15277_;
wire _15278_;
wire _15279_;
wire _15280_;
wire _15281_;
wire _15282_;
wire _15283_;
wire _15284_;
wire _15285_;
wire _15286_;
wire _15287_;
wire _15288_;
wire _15289_;
wire _15290_;
wire _15291_;
wire _15292_;
wire _15293_;
wire _15294_;
wire _15295_;
wire _15296_;
wire _15297_;
wire _15298_;
wire _15299_;
wire _15300_;
wire _15301_;
wire _15302_;
wire _15303_;
wire _15304_;
wire _15305_;
wire _15306_;
wire _15307_;
wire _15308_;
wire _15309_;
wire _15310_;
wire _15311_;
wire _15312_;
wire _15313_;
wire _15314_;
wire _15315_;
wire _15316_;
wire _15317_;
wire _15318_;
wire _15319_;
wire _15320_;
wire _15321_;
wire _15322_;
wire _15323_;
wire _15324_;
wire _15325_;
wire _15326_;
wire _15327_;
wire _15328_;
wire _15329_;
wire _15330_;
wire _15331_;
wire _15332_;
wire _15333_;
wire _15334_;
wire _15335_;
wire _15336_;
wire _15337_;
wire _15338_;
wire _15339_;
wire _15340_;
wire _15341_;
wire _15342_;
wire _15343_;
wire _15344_;
wire _15345_;
wire _15346_;
wire _15347_;
wire _15348_;
wire _15349_;
wire _15350_;
wire _15351_;
wire _15352_;
wire _15353_;
wire _15354_;
wire _15355_;
wire _15356_;
wire _15357_;
wire _15358_;
wire _15359_;
wire _15360_;
wire _15361_;
wire _15362_;
wire _15363_;
wire _15364_;
wire _15365_;
wire _15366_;
wire _15367_;
wire _15368_;
wire _15369_;
wire _15370_;
wire _15371_;
wire _15372_;
wire _15373_;
wire _15374_;
wire _15375_;
wire _15376_;
wire _15377_;
wire _15378_;
wire _15379_;
wire _15380_;
wire _15381_;
wire _15382_;
wire _15383_;
wire _15384_;
wire _15385_;
wire _15386_;
wire _15387_;
wire _15388_;
wire _15389_;
wire _15390_;
wire _15391_;
wire _15392_;
wire _15393_;
wire _15394_;
wire _15395_;
wire _15396_;
wire _15397_;
wire _15398_;
wire _15399_;
wire _15400_;
wire _15401_;
wire _15402_;
wire _15403_;
wire _15404_;
wire _15405_;
wire _15406_;
wire _15407_;
wire _15408_;
wire _15409_;
wire _15410_;
wire _15411_;
wire _15412_;
wire _15413_;
wire _15414_;
wire _15415_;
wire _15416_;
wire _15417_;
wire _15418_;
wire _15419_;
wire _15420_;
wire _15421_;
wire _15422_;
wire _15423_;
wire _15424_;
wire _15425_;
wire _15426_;
wire _15427_;
wire _15428_;
wire _15429_;
wire _15430_;
wire _15431_;
wire _15432_;
wire _15433_;
wire _15434_;
wire _15435_;
wire _15436_;
wire _15437_;
wire _15438_;
wire _15439_;
wire _15440_;
wire _15441_;
wire _15442_;
wire _15443_;
wire _15444_;
wire _15445_;
wire _15446_;
wire _15447_;
wire _15448_;
wire _15449_;
wire _15450_;
wire _15451_;
wire _15452_;
wire _15453_;
wire _15454_;
wire _15455_;
wire _15456_;
wire _15457_;
wire _15458_;
wire _15459_;
wire _15460_;
wire _15461_;
wire _15462_;
wire _15463_;
wire _15464_;
wire _15465_;
wire _15466_;
wire _15467_;
wire _15468_;
wire _15469_;
wire _15470_;
wire _15471_;
wire _15472_;
wire _15473_;
wire _15474_;
wire _15475_;
wire _15476_;
wire _15477_;
wire _15478_;
wire _15479_;
wire _15480_;
wire _15481_;
wire _15482_;
wire _15483_;
wire _15484_;
wire _15485_;
wire _15486_;
wire _15487_;
wire _15488_;
wire _15489_;
wire _15490_;
wire _15491_;
wire _15492_;
wire _15493_;
wire _15494_;
wire _15495_;
wire _15496_;
wire _15497_;
wire _15498_;
wire _15499_;
wire _15500_;
wire _15501_;
wire _15502_;
wire _15503_;
wire _15504_;
wire _15505_;
wire _15506_;
wire _15507_;
wire _15508_;
wire _15509_;
wire _15510_;
wire _15511_;
wire _15512_;
wire _15513_;
wire _15514_;
wire _15515_;
wire _15516_;
wire _15517_;
wire _15518_;
wire _15519_;
wire _15520_;
wire _15521_;
wire _15522_;
wire _15523_;
wire _15524_;
wire _15525_;
wire _15526_;
wire _15527_;
wire _15528_;
wire _15529_;
wire _15530_;
wire _15531_;
wire _15532_;
wire _15533_;
wire _15534_;
wire _15535_;
wire _15536_;
wire _15537_;
wire _15538_;
wire _15539_;
wire _15540_;
wire _15541_;
wire _15542_;
wire _15543_;
wire _15544_;
wire _15545_;
wire _15546_;
wire _15547_;
wire _15548_;
wire _15549_;
wire _15550_;
wire _15551_;
wire _15552_;
wire _15553_;
wire _15554_;
wire _15555_;
wire _15556_;
wire _15557_;
wire _15558_;
wire _15559_;
wire _15560_;
wire _15561_;
wire _15562_;
wire _15563_;
wire _15564_;
wire _15565_;
wire _15566_;
wire _15567_;
wire _15568_;
wire _15569_;
wire _15570_;
wire _15571_;
wire _15572_;
wire _15573_;
wire _15574_;
wire _15575_;
wire _15576_;
wire _15577_;
wire _15578_;
wire _15579_;
wire _15580_;
wire _15581_;
wire _15582_;
wire _15583_;
wire _15584_;
wire _15585_;
wire _15586_;
wire _15587_;
wire _15588_;
wire _15589_;
wire _15590_;
wire _15591_;
wire _15592_;
wire _15593_;
wire _15594_;
wire _15595_;
wire _15596_;
wire _15597_;
wire _15598_;
wire _15599_;
wire _15600_;
wire _15601_;
wire _15602_;
wire _15603_;
wire _15604_;
wire _15605_;
wire _15606_;
wire _15607_;
wire _15608_;
wire _15609_;
wire _15610_;
wire _15611_;
wire _15612_;
wire _15613_;
wire _15614_;
wire _15615_;
wire _15616_;
wire _15617_;
wire _15618_;
wire _15619_;
wire _15620_;
wire _15621_;
wire _15622_;
wire _15623_;
wire _15624_;
wire _15625_;
wire _15626_;
wire _15627_;
wire _15628_;
wire _15629_;
wire _15630_;
wire _15631_;
wire _15632_;
wire _15633_;
wire _15634_;
wire _15635_;
wire _15636_;
wire _15637_;
wire _15638_;
wire _15639_;
wire _15640_;
wire _15641_;
wire _15642_;
wire _15643_;
wire _15644_;
wire _15645_;
wire _15646_;
wire _15647_;
wire _15648_;
wire _15649_;
wire _15650_;
wire _15651_;
wire _15652_;
wire _15653_;
wire _15654_;
wire _15655_;
wire _15656_;
wire _15657_;
wire _15658_;
wire _15659_;
wire _15660_;
wire _15661_;
wire _15662_;
wire _15663_;
wire _15664_;
wire _15665_;
wire _15666_;
wire _15667_;
wire _15668_;
wire _15669_;
wire _15670_;
wire _15671_;
wire _15672_;
wire _15673_;
wire _15674_;
wire _15675_;
wire _15676_;
wire _15677_;
wire _15678_;
wire _15679_;
wire _15680_;
wire _15681_;
wire _15682_;
wire _15683_;
wire _15684_;
wire _15685_;
wire _15686_;
wire _15687_;
wire _15688_;
wire _15689_;
wire _15690_;
wire _15691_;
wire _15692_;
wire _15693_;
wire _15694_;
wire _15695_;
wire _15696_;
wire _15697_;
wire _15698_;
wire _15699_;
wire _15700_;
wire _15701_;
wire _15702_;
wire _15703_;
wire _15704_;
wire _15705_;
wire _15706_;
wire _15707_;
wire _15708_;
wire _15709_;
wire _15710_;
wire _15711_;
wire _15712_;
wire _15713_;
wire _15714_;
wire _15715_;
wire _15716_;
wire _15717_;
wire _15718_;
wire _15719_;
wire _15720_;
wire _15721_;
wire _15722_;
wire _15723_;
wire _15724_;
wire _15725_;
wire _15726_;
wire _15727_;
wire _15728_;
wire _15729_;
wire _15730_;
wire _15731_;
wire _15732_;
wire _15733_;
wire _15734_;
wire _15735_;
wire _15736_;
wire _15737_;
wire _15738_;
wire _15739_;
wire _15740_;
wire _15741_;
wire _15742_;
wire _15743_;
wire _15744_;
wire _15745_;
wire _15746_;
wire _15747_;
wire _15748_;
wire _15749_;
wire _15750_;
wire _15751_;
wire _15752_;
wire _15753_;
wire _15754_;
wire _15755_;
wire _15756_;
wire _15757_;
wire _15758_;
wire _15759_;
wire _15760_;
wire _15761_;
wire _15762_;
wire _15763_;
wire _15764_;
wire _15765_;
wire _15766_;
wire _15767_;
wire _15768_;
wire _15769_;
wire _15770_;
wire _15771_;
wire _15772_;
wire _15773_;
wire _15774_;
wire _15775_;
wire _15776_;
wire _15777_;
wire _15778_;
wire _15779_;
wire _15780_;
wire _15781_;
wire _15782_;
wire _15783_;
wire _15784_;
wire _15785_;
wire _15786_;
wire _15787_;
wire _15788_;
wire _15789_;
wire _15790_;
wire _15791_;
wire _15792_;
wire _15793_;
wire _15794_;
wire _15795_;
wire _15796_;
wire _15797_;
wire _15798_;
wire _15799_;
wire _15800_;
wire _15801_;
wire _15802_;
wire _15803_;
wire _15804_;
wire _15805_;
wire _15806_;
wire _15807_;
wire _15808_;
wire _15809_;
wire _15810_;
wire _15811_;
wire _15812_;
wire _15813_;
wire _15814_;
wire _15815_;
wire _15816_;
wire _15817_;
wire _15818_;
wire _15819_;
wire _15820_;
wire _15821_;
wire _15822_;
wire _15823_;
wire _15824_;
wire _15825_;
wire _15826_;
wire _15827_;
wire _15828_;
wire _15829_;
wire _15830_;
wire _15831_;
wire _15832_;
wire _15833_;
wire _15834_;
wire _15835_;
wire _15836_;
wire _15837_;
wire _15838_;
wire _15839_;
wire _15840_;
wire _15841_;
wire _15842_;
wire _15843_;
wire _15844_;
wire _15845_;
wire _15846_;
wire _15847_;
wire _15848_;
wire _15849_;
wire _15850_;
wire _15851_;
wire _15852_;
wire _15853_;
wire _15854_;
wire _15855_;
wire _15856_;
wire _15857_;
wire _15858_;
wire _15859_;
wire _15860_;
wire _15861_;
wire _15862_;
wire _15863_;
wire _15864_;
wire _15865_;
wire _15866_;
wire _15867_;
wire _15868_;
wire _15869_;
wire _15870_;
wire _15871_;
wire _15872_;
wire _15873_;
wire _15874_;
wire _15875_;
wire _15876_;
wire _15877_;
wire _15878_;
wire _15879_;
wire _15880_;
wire _15881_;
wire _15882_;
wire _15883_;
wire _15884_;
wire _15885_;
wire _15886_;
wire _15887_;
wire _15888_;
wire _15889_;
wire _15890_;
wire _15891_;
wire _15892_;
wire _15893_;
wire _15894_;
wire _15895_;
wire _15896_;
wire _15897_;
wire _15898_;
wire _15899_;
wire _15900_;
wire _15901_;
wire _15902_;
wire _15903_;
wire _15904_;
wire _15905_;
wire _15906_;
wire _15907_;
wire _15908_;
wire _15909_;
wire _15910_;
wire _15911_;
wire _15912_;
wire _15913_;
wire _15914_;
wire _15915_;
wire _15916_;
wire _15917_;
wire _15918_;
wire _15919_;
wire _15920_;
wire _15921_;
wire _15922_;
wire _15923_;
wire _15924_;
wire _15925_;
wire _15926_;
wire _15927_;
wire _15928_;
wire _15929_;
wire _15930_;
wire _15931_;
wire _15932_;
wire _15933_;
wire _15934_;
wire _15935_;
wire _15936_;
wire _15937_;
wire _15938_;
wire _15939_;
wire _15940_;
wire _15941_;
wire _15942_;
wire _15943_;
wire _15944_;
wire _15945_;
wire _15946_;
wire _15947_;
wire _15948_;
wire _15949_;
wire _15950_;
wire _15951_;
wire _15952_;
wire _15953_;
wire _15954_;
wire _15955_;
wire _15956_;
wire _15957_;
wire _15958_;
wire _15959_;
wire _15960_;
wire _15961_;
wire _15962_;
wire _15963_;
wire _15964_;
wire _15965_;
wire _15966_;
wire _15967_;
wire _15968_;
wire _15969_;
wire _15970_;
wire _15971_;
wire _15972_;
wire _15973_;
wire _15974_;
wire _15975_;
wire _15976_;
wire _15977_;
wire _15978_;
wire _15979_;
wire _15980_;
wire _15981_;
wire _15982_;
wire _15983_;
wire _15984_;
wire _15985_;
wire _15986_;
wire _15987_;
wire _15988_;
wire _15989_;
wire _15990_;
wire _15991_;
wire _15992_;
wire _15993_;
wire _15994_;
wire _15995_;
wire _15996_;
wire _15997_;
wire _15998_;
wire _15999_;
wire _16000_;
wire _16001_;
wire _16002_;
wire _16003_;
wire _16004_;
wire _16005_;
wire _16006_;
wire _16007_;
wire _16008_;
wire _16009_;
wire _16010_;
wire _16011_;
wire _16012_;
wire _16013_;
wire _16014_;
wire _16015_;
wire _16016_;
wire _16017_;
wire _16018_;
wire _16019_;
wire _16020_;
wire _16021_;
wire _16022_;
wire _16023_;
wire _16024_;
wire _16025_;
wire _16026_;
wire _16027_;
wire _16028_;
wire _16029_;
wire _16030_;
wire _16031_;
wire _16032_;
wire _16033_;
wire _16034_;
wire _16035_;
wire _16036_;
wire _16037_;
wire _16038_;
wire _16039_;
wire _16040_;
wire _16041_;
wire _16042_;
wire _16043_;
wire _16044_;
wire _16045_;
wire _16046_;
wire _16047_;
wire _16048_;
wire _16049_;
wire _16050_;
wire _16051_;
wire _16052_;
wire _16053_;
wire _16054_;
wire _16055_;
wire _16056_;
wire _16057_;
wire _16058_;
wire _16059_;
wire _16060_;
wire _16061_;
wire _16062_;
wire _16063_;
wire _16064_;
wire _16065_;
wire _16066_;
wire _16067_;
wire _16068_;
wire _16069_;
wire _16070_;
wire _16071_;
wire _16072_;
wire _16073_;
wire _16074_;
wire _16075_;
wire _16076_;
wire _16077_;
wire _16078_;
wire _16079_;
wire _16080_;
wire _16081_;
wire _16082_;
wire _16083_;
wire _16084_;
wire _16085_;
wire _16086_;
wire _16087_;
wire _16088_;
wire _16089_;
wire _16090_;
wire _16091_;
wire _16092_;
wire _16093_;
wire _16094_;
wire _16095_;
wire _16096_;
wire _16097_;
wire _16098_;
wire _16099_;
wire _16100_;
wire _16101_;
wire _16102_;
wire _16103_;
wire _16104_;
wire _16105_;
wire _16106_;
wire _16107_;
wire _16108_;
wire _16109_;
wire _16110_;
wire _16111_;
wire _16112_;
wire _16113_;
wire _16114_;
wire _16115_;
wire _16116_;
wire _16117_;
wire _16118_;
wire _16119_;
wire _16120_;
wire _16121_;
wire _16122_;
wire _16123_;
wire _16124_;
wire _16125_;
wire _16126_;
wire _16127_;
wire _16128_;
wire _16129_;
wire _16130_;
wire _16131_;
wire _16132_;
wire _16133_;
wire _16134_;
wire _16135_;
wire _16136_;
wire _16137_;
wire _16138_;
wire _16139_;
wire _16140_;
wire _16141_;
wire _16142_;
wire _16143_;
wire _16144_;
wire _16145_;
wire _16146_;
wire _16147_;
wire _16148_;
wire _16149_;
wire _16150_;
wire _16151_;
wire _16152_;
wire _16153_;
wire _16154_;
wire _16155_;
wire _16156_;
wire _16157_;
wire _16158_;
wire _16159_;
wire _16160_;
wire _16161_;
wire _16162_;
wire _16163_;
wire _16164_;
wire _16165_;
wire _16166_;
wire _16167_;
wire _16168_;
wire _16169_;
wire _16170_;
wire _16171_;
wire _16172_;
wire _16173_;
wire _16174_;
wire _16175_;
wire _16176_;
wire _16177_;
wire _16178_;
wire _16179_;
wire _16180_;
wire _16181_;
wire _16182_;
wire _16183_;
wire _16184_;
wire _16185_;
wire _16186_;
wire _16187_;
wire _16188_;
wire _16189_;
wire _16190_;
wire _16191_;
wire _16192_;
wire _16193_;
wire _16194_;
wire _16195_;
wire _16196_;
wire _16197_;
wire _16198_;
wire _16199_;
wire _16200_;
wire _16201_;
wire _16202_;
wire _16203_;
wire _16204_;
wire _16205_;
wire _16206_;
wire _16207_;
wire _16208_;
wire _16209_;
wire _16210_;
wire _16211_;
wire _16212_;
wire _16213_;
wire _16214_;
wire _16215_;
wire _16216_;
wire _16217_;
wire _16218_;
wire _16219_;
wire _16220_;
wire _16221_;
wire _16222_;
wire _16223_;
wire _16224_;
wire _16225_;
wire _16226_;
wire _16227_;
wire _16228_;
wire _16229_;
wire _16230_;
wire _16231_;
wire _16232_;
wire _16233_;
wire _16234_;
wire _16235_;
wire _16236_;
wire _16237_;
wire _16238_;
wire _16239_;
wire _16240_;
wire _16241_;
wire _16242_;
wire _16243_;
wire _16244_;
wire _16245_;
wire _16246_;
wire _16247_;
wire _16248_;
wire _16249_;
wire _16250_;
wire _16251_;
wire _16252_;
wire _16253_;
wire _16254_;
wire _16255_;
wire _16256_;
wire _16257_;
wire _16258_;
wire _16259_;
wire _16260_;
wire _16261_;
wire _16262_;
wire _16263_;
wire _16264_;
wire _16265_;
wire _16266_;
wire _16267_;
wire _16268_;
wire _16269_;
wire _16270_;
wire _16271_;
wire _16272_;
wire _16273_;
wire _16274_;
wire _16275_;
wire _16276_;
wire _16277_;
wire _16278_;
wire _16279_;
wire _16280_;
wire _16281_;
wire _16282_;
wire _16283_;
wire _16284_;
wire _16285_;
wire _16286_;
wire _16287_;
wire _16288_;
wire _16289_;
wire _16290_;
wire _16291_;
wire _16292_;
wire _16293_;
wire _16294_;
wire _16295_;
wire _16296_;
wire _16297_;
wire _16298_;
wire _16299_;
wire _16300_;
wire _16301_;
wire _16302_;
wire _16303_;
wire _16304_;
wire _16305_;
wire _16306_;
wire _16307_;
wire _16308_;
wire _16309_;
wire _16310_;
wire _16311_;
wire _16312_;
wire _16313_;
wire _16314_;
wire _16315_;
wire _16316_;
wire _16317_;
wire _16318_;
wire _16319_;
wire _16320_;
wire _16321_;
wire _16322_;
wire _16323_;
wire _16324_;
wire _16325_;
wire _16326_;
wire _16327_;
wire _16328_;
wire _16329_;
wire _16330_;
wire _16331_;
wire _16332_;
wire _16333_;
wire _16334_;
wire _16335_;
wire _16336_;
wire _16337_;
wire _16338_;
wire _16339_;
wire _16340_;
wire _16341_;
wire _16342_;
wire _16343_;
wire _16344_;
wire _16345_;
wire _16346_;
wire _16347_;
wire _16348_;
wire _16349_;
wire _16350_;
wire _16351_;
wire _16352_;
wire _16353_;
wire _16354_;
wire _16355_;
wire _16356_;
wire _16357_;
wire _16358_;
wire _16359_;
wire _16360_;
wire _16361_;
wire _16362_;
wire _16363_;
wire _16364_;
wire _16365_;
wire _16366_;
wire _16367_;
wire _16368_;
wire _16369_;
wire _16370_;
wire _16371_;
wire _16372_;
wire _16373_;
wire _16374_;
wire _16375_;
wire _16376_;
wire _16377_;
wire _16378_;
wire _16379_;
wire _16380_;
wire _16381_;
wire _16382_;
wire _16383_;
wire _16384_;
wire _16385_;
wire _16386_;
wire _16387_;
wire _16388_;
wire _16389_;
wire _16390_;
wire _16391_;
wire _16392_;
wire _16393_;
wire _16394_;
wire _16395_;
wire _16396_;
wire _16397_;
wire _16398_;
wire _16399_;
wire _16400_;
wire _16401_;
wire _16402_;
wire _16403_;
wire _16404_;
wire _16405_;
wire _16406_;
wire _16407_;
wire _16408_;
wire _16409_;
wire _16410_;
wire _16411_;
wire _16412_;
wire _16413_;
wire _16414_;
wire _16415_;
wire _16416_;
wire _16417_;
wire _16418_;
wire _16419_;
wire _16420_;
wire _16421_;
wire _16422_;
wire _16423_;
wire _16424_;
wire _16425_;
wire _16426_;
wire _16427_;
wire _16428_;
wire _16429_;
wire _16430_;
wire _16431_;
wire _16432_;
wire _16433_;
wire _16434_;
wire _16435_;
wire _16436_;
wire _16437_;
wire _16438_;
wire _16439_;
wire _16440_;
wire _16441_;
wire _16442_;
wire _16443_;
wire _16444_;
wire _16445_;
wire _16446_;
wire _16447_;
wire _16448_;
wire _16449_;
wire _16450_;
wire _16451_;
wire _16452_;
wire _16453_;
wire _16454_;
wire _16455_;
wire _16456_;
wire _16457_;
wire _16458_;
wire _16459_;
wire _16460_;
wire _16461_;
wire _16462_;
wire _16463_;
wire _16464_;
wire _16465_;
wire _16466_;
wire _16467_;
wire _16468_;
wire _16469_;
wire _16470_;
wire _16471_;
wire _16472_;
wire _16473_;
wire _16474_;
wire _16475_;
wire _16476_;
wire _16477_;
wire _16478_;
wire _16479_;
wire _16480_;
wire _16481_;
wire _16482_;
wire _16483_;
wire _16484_;
wire _16485_;
wire _16486_;
wire _16487_;
wire _16488_;
wire _16489_;
wire _16490_;
wire _16491_;
wire _16492_;
wire _16493_;
wire _16494_;
wire _16495_;
wire _16496_;
wire _16497_;
wire _16498_;
wire _16499_;
wire _16500_;
wire _16501_;
wire _16502_;
wire _16503_;
wire _16504_;
wire _16505_;
wire _16506_;
wire _16507_;
wire _16508_;
wire _16509_;
wire _16510_;
wire _16511_;
wire _16512_;
wire _16513_;
wire _16514_;
wire _16515_;
wire _16516_;
wire _16517_;
wire _16518_;
wire _16519_;
wire _16520_;
wire _16521_;
wire _16522_;
wire _16523_;
wire _16524_;
wire _16525_;
wire _16526_;
wire _16527_;
wire _16528_;
wire _16529_;
wire _16530_;
wire _16531_;
wire _16532_;
wire _16533_;
wire _16534_;
wire _16535_;
wire _16536_;
wire _16537_;
wire _16538_;
wire _16539_;
wire _16540_;
wire _16541_;
wire _16542_;
wire _16543_;
wire _16544_;
wire _16545_;
wire _16546_;
wire _16547_;
wire _16548_;
wire _16549_;
wire _16550_;
wire _16551_;
wire _16552_;
wire _16553_;
wire _16554_;
wire _16555_;
wire _16556_;
wire _16557_;
wire _16558_;
wire _16559_;
wire _16560_;
wire _16561_;
wire _16562_;
wire _16563_;
wire _16564_;
wire _16565_;
wire _16566_;
wire _16567_;
wire _16568_;
wire _16569_;
wire _16570_;
wire _16571_;
wire _16572_;
wire _16573_;
wire _16574_;
wire _16575_;
wire _16576_;
wire _16577_;
wire _16578_;
wire _16579_;
wire _16580_;
wire _16581_;
wire _16582_;
wire _16583_;
wire _16584_;
wire _16585_;
wire _16586_;
wire _16587_;
wire _16588_;
wire _16589_;
wire _16590_;
wire _16591_;
wire _16592_;
wire _16593_;
wire _16594_;
wire _16595_;
wire _16596_;
wire _16597_;
wire _16598_;
wire _16599_;
wire _16600_;
wire _16601_;
wire _16602_;
wire _16603_;
wire _16604_;
wire _16605_;
wire _16606_;
wire _16607_;
wire _16608_;
wire _16609_;
wire _16610_;
wire _16611_;
wire _16612_;
wire _16613_;
wire _16614_;
wire _16615_;
wire _16616_;
wire _16617_;
wire _16618_;
wire _16619_;
wire _16620_;
wire _16621_;
wire _16622_;
wire _16623_;
wire _16624_;
wire _16625_;
wire _16626_;
wire _16627_;
wire _16628_;
wire _16629_;
wire _16630_;
wire _16631_;
wire _16632_;
wire _16633_;
wire _16634_;
wire _16635_;
wire _16636_;
wire _16637_;
wire _16638_;
wire _16639_;
wire _16640_;
wire _16641_;
wire _16642_;
wire _16643_;
wire _16644_;
wire _16645_;
wire _16646_;
wire _16647_;
wire _16648_;
wire _16649_;
wire _16650_;
wire _16651_;
wire _16652_;
wire _16653_;
wire _16654_;
wire _16655_;
wire _16656_;
wire _16657_;
wire _16658_;
wire _16659_;
wire _16660_;
wire _16661_;
wire _16662_;
wire _16663_;
wire _16664_;
wire _16665_;
wire _16666_;
wire _16667_;
wire _16668_;
wire _16669_;
wire _16670_;
wire _16671_;
wire _16672_;
wire _16673_;
wire _16674_;
wire _16675_;
wire _16676_;
wire _16677_;
wire _16678_;
wire _16679_;
wire _16680_;
wire _16681_;
wire _16682_;
wire _16683_;
wire _16684_;
wire _16685_;
wire _16686_;
wire _16687_;
wire _16688_;
wire _16689_;
wire _16690_;
wire _16691_;
wire _16692_;
wire _16693_;
wire _16694_;
wire _16695_;
wire _16696_;
wire _16697_;
wire _16698_;
wire _16699_;
wire _16700_;
wire _16701_;
wire _16702_;
wire _16703_;
wire _16704_;
wire _16705_;
wire _16706_;
wire _16707_;
wire _16708_;
wire _16709_;
wire _16710_;
wire _16711_;
wire _16712_;
wire _16713_;
wire _16714_;
wire _16715_;
wire _16716_;
wire _16717_;
wire _16718_;
wire _16719_;
wire _16720_;
wire _16721_;
wire _16722_;
wire _16723_;
wire _16724_;
wire _16725_;
wire _16726_;
wire _16727_;
wire _16728_;
wire _16729_;
wire _16730_;
wire _16731_;
wire _16732_;
wire _16733_;
wire _16734_;
wire _16735_;
wire _16736_;
wire _16737_;
wire _16738_;
wire _16739_;
wire _16740_;
wire _16741_;
wire _16742_;
wire _16743_;
wire _16744_;
wire _16745_;
wire _16746_;
wire _16747_;
wire _16748_;
wire _16749_;
wire _16750_;
wire _16751_;
wire _16752_;
wire _16753_;
wire _16754_;
wire _16755_;
wire _16756_;
wire _16757_;
wire _16758_;
wire _16759_;
wire _16760_;
wire _16761_;
wire _16762_;
wire _16763_;
wire _16764_;
wire _16765_;
wire _16766_;
wire _16767_;
wire _16768_;
wire _16769_;
wire _16770_;
wire _16771_;
wire _16772_;
wire _16773_;
wire _16774_;
wire _16775_;
wire _16776_;
wire _16777_;
wire _16778_;
wire _16779_;
wire _16780_;
wire _16781_;
wire _16782_;
wire _16783_;
wire _16784_;
wire _16785_;
wire _16786_;
wire _16787_;
wire _16788_;
wire _16789_;
wire _16790_;
wire _16791_;
wire _16792_;
wire _16793_;
wire _16794_;
wire _16795_;
wire _16796_;
wire _16797_;
wire _16798_;
wire _16799_;
wire _16800_;
wire _16801_;
wire _16802_;
wire _16803_;
wire _16804_;
wire _16805_;
wire _16806_;
wire _16807_;
wire _16808_;
wire _16809_;
wire _16810_;
wire _16811_;
wire _16812_;
wire _16813_;
wire _16814_;
wire _16815_;
wire _16816_;
wire _16817_;
wire _16818_;
wire _16819_;
wire _16820_;
wire _16821_;
wire _16822_;
wire _16823_;
wire _16824_;
wire _16825_;
wire _16826_;
wire _16827_;
wire _16828_;
wire _16829_;
wire _16830_;
wire _16831_;
wire _16832_;
wire _16833_;
wire _16834_;
wire _16835_;
wire _16836_;
wire _16837_;
wire _16838_;
wire _16839_;
wire _16840_;
wire _16841_;
wire _16842_;
wire _16843_;
wire _16844_;
wire _16845_;
wire _16846_;
wire _16847_;
wire _16848_;
wire _16849_;
wire _16850_;
wire _16851_;
wire _16852_;
wire _16853_;
wire _16854_;
wire _16855_;
wire _16856_;
wire _16857_;
wire _16858_;
wire _16859_;
wire _16860_;
wire _16861_;
wire _16862_;
wire _16863_;
wire _16864_;
wire _16865_;
wire _16866_;
wire _16867_;
wire _16868_;
wire _16869_;
wire _16870_;
wire _16871_;
wire _16872_;
wire _16873_;
wire _16874_;
wire _16875_;
wire _16876_;
wire _16877_;
wire _16878_;
wire _16879_;
wire _16880_;
wire _16881_;
wire _16882_;
wire _16883_;
wire _16884_;
wire _16885_;
wire _16886_;
wire _16887_;
wire _16888_;
wire _16889_;
wire _16890_;
wire _16891_;
wire _16892_;
wire _16893_;
wire _16894_;
wire _16895_;
wire _16896_;
wire _16897_;
wire _16898_;
wire _16899_;
wire _16900_;
wire _16901_;
wire _16902_;
wire _16903_;
wire _16904_;
wire _16905_;
wire _16906_;
wire _16907_;
wire _16908_;
wire _16909_;
wire _16910_;
wire _16911_;
wire _16912_;
wire _16913_;
wire _16914_;
wire _16915_;
wire _16916_;
wire _16917_;
wire _16918_;
wire _16919_;
wire _16920_;
wire _16921_;
wire _16922_;
wire _16923_;
wire _16924_;
wire _16925_;
wire _16926_;
wire _16927_;
wire _16928_;
wire _16929_;
wire _16930_;
wire _16931_;
wire _16932_;
wire _16933_;
wire _16934_;
wire _16935_;
wire _16936_;
wire _16937_;
wire _16938_;
wire _16939_;
wire _16940_;
wire _16941_;
wire _16942_;
wire _16943_;
wire _16944_;
wire _16945_;
wire _16946_;
wire _16947_;
wire _16948_;
wire _16949_;
wire _16950_;
wire _16951_;
wire _16952_;
wire _16953_;
wire _16954_;
wire _16955_;
wire _16956_;
wire _16957_;
wire _16958_;
wire _16959_;
wire _16960_;
wire _16961_;
wire _16962_;
wire _16963_;
wire _16964_;
wire _16965_;
wire _16966_;
wire _16967_;
wire _16968_;
wire _16969_;
wire _16970_;
wire _16971_;
wire _16972_;
wire _16973_;
wire _16974_;
wire _16975_;
wire _16976_;
wire _16977_;
wire _16978_;
wire _16979_;
wire _16980_;
wire _16981_;
wire _16982_;
wire _16983_;
wire _16984_;
wire _16985_;
wire _16986_;
wire _16987_;
wire _16988_;
wire _16989_;
wire _16990_;
wire _16991_;
wire _16992_;
wire _16993_;
wire _16994_;
wire _16995_;
wire _16996_;
wire _16997_;
wire _16998_;
wire _16999_;
wire _17000_;
wire _17001_;
wire _17002_;
wire _17003_;
wire _17004_;
wire _17005_;
wire _17006_;
wire _17007_;
wire _17008_;
wire _17009_;
wire _17010_;
wire _17011_;
wire _17012_;
wire _17013_;
wire _17014_;
wire _17015_;
wire _17016_;
wire _17017_;
wire _17018_;
wire _17019_;
wire _17020_;
wire _17021_;
wire _17022_;
wire _17023_;
wire _17024_;
wire _17025_;
wire _17026_;
wire _17027_;
wire _17028_;
wire _17029_;
wire _17030_;
wire _17031_;
wire _17032_;
wire _17033_;
wire _17034_;
wire _17035_;
wire _17036_;
wire _17037_;
wire _17038_;
wire _17039_;
wire _17040_;
wire _17041_;
wire _17042_;
wire _17043_;
wire _17044_;
wire _17045_;
wire _17046_;
wire _17047_;
wire _17048_;
wire _17049_;
wire _17050_;
wire _17051_;
wire _17052_;
wire _17053_;
wire _17054_;
wire _17055_;
wire _17056_;
wire _17057_;
wire _17058_;
wire _17059_;
wire _17060_;
wire _17061_;
wire _17062_;
wire _17063_;
wire _17064_;
wire _17065_;
wire _17066_;
wire _17067_;
wire _17068_;
wire _17069_;
wire _17070_;
wire _17071_;
wire _17072_;
wire _17073_;
wire _17074_;
wire _17075_;
wire _17076_;
wire _17077_;
wire _17078_;
wire _17079_;
wire _17080_;
wire _17081_;
wire _17082_;
wire _17083_;
wire _17084_;
wire _17085_;
wire _17086_;
wire _17087_;
wire _17088_;
wire _17089_;
wire _17090_;
wire _17091_;
wire _17092_;
wire _17093_;
wire _17094_;
wire _17095_;
wire _17096_;
wire _17097_;
wire _17098_;
wire _17099_;
wire _17100_;
wire _17101_;
wire _17102_;
wire _17103_;
wire _17104_;
wire _17105_;
wire _17106_;
wire _17107_;
wire _17108_;
wire _17109_;
wire _17110_;
wire _17111_;
wire _17112_;
wire _17113_;
wire _17114_;
wire _17115_;
wire _17116_;
wire _17117_;
wire _17118_;
wire _17119_;
wire _17120_;
wire _17121_;
wire _17122_;
wire _17123_;
wire _17124_;
wire _17125_;
wire _17126_;
wire _17127_;
wire _17128_;
wire _17129_;
wire _17130_;
wire _17131_;
wire _17132_;
wire _17133_;
wire _17134_;
wire _17135_;
wire _17136_;
wire _17137_;
wire _17138_;
wire _17139_;
wire _17140_;
wire _17141_;
wire _17142_;
wire _17143_;
wire _17144_;
wire _17145_;
wire _17146_;
wire _17147_;
wire _17148_;
wire _17149_;
wire _17150_;
wire _17151_;
wire _17152_;
wire _17153_;
wire _17154_;
wire _17155_;
wire _17156_;
wire _17157_;
wire _17158_;
wire _17159_;
wire _17160_;
wire _17161_;
wire _17162_;
wire _17163_;
wire _17164_;
wire _17165_;
wire _17166_;
wire _17167_;
wire _17168_;
wire _17169_;
wire _17170_;
wire _17171_;
wire _17172_;
wire _17173_;
wire _17174_;
wire _17175_;
wire _17176_;
wire _17177_;
wire _17178_;
wire _17179_;
wire _17180_;
wire _17181_;
wire _17182_;
wire _17183_;
wire _17184_;
wire _17185_;
wire _17186_;
wire _17187_;
wire _17188_;
wire _17189_;
wire _17190_;
wire _17191_;
wire _17192_;
wire _17193_;
wire _17194_;
wire _17195_;
wire _17196_;
wire _17197_;
wire _17198_;
wire _17199_;
wire _17200_;
wire _17201_;
wire _17202_;
wire _17203_;
wire _17204_;
wire _17205_;
wire _17206_;
wire _17207_;
wire _17208_;
wire _17209_;
wire _17210_;
wire _17211_;
wire _17212_;
wire _17213_;
wire _17214_;
wire _17215_;
wire _17216_;
wire _17217_;
wire _17218_;
wire _17219_;
wire _17220_;
wire _17221_;
wire _17222_;
wire _17223_;
wire _17224_;
wire _17225_;
wire _17226_;
wire _17227_;
wire _17228_;
wire _17229_;
wire _17230_;
wire _17231_;
wire _17232_;
wire _17233_;
wire _17234_;
wire _17235_;
wire _17236_;
wire _17237_;
wire _17238_;
wire _17239_;
wire _17240_;
wire _17241_;
wire _17242_;
wire _17243_;
wire _17244_;
wire _17245_;
wire _17246_;
wire _17247_;
wire _17248_;
wire _17249_;
wire _17250_;
wire _17251_;
wire _17252_;
wire _17253_;
wire _17254_;
wire _17255_;
wire _17256_;
wire _17257_;
wire _17258_;
wire _17259_;
wire _17260_;
wire _17261_;
wire _17262_;
wire _17263_;
wire _17264_;
wire _17265_;
wire _17266_;
wire _17267_;
wire _17268_;
wire _17269_;
wire _17270_;
wire _17271_;
wire _17272_;
wire _17273_;
wire _17274_;
wire _17275_;
wire _17276_;
wire _17277_;
wire _17278_;
wire _17279_;
wire _17280_;
wire _17281_;
wire _17282_;
wire _17283_;
wire _17284_;
wire _17285_;
wire _17286_;
wire _17287_;
wire _17288_;
wire _17289_;
wire _17290_;
wire _17291_;
wire _17292_;
wire _17293_;
wire _17294_;
wire _17295_;
wire _17296_;
wire _17297_;
wire _17298_;
wire _17299_;
wire _17300_;
wire _17301_;
wire _17302_;
wire _17303_;
wire _17304_;
wire _17305_;
wire _17306_;
wire _17307_;
wire _17308_;
wire _17309_;
wire _17310_;
wire _17311_;
wire _17312_;
wire _17313_;
wire _17314_;
wire _17315_;
wire _17316_;
wire _17317_;
wire _17318_;
wire _17319_;
wire _17320_;
wire _17321_;
wire _17322_;
wire _17323_;
wire _17324_;
wire _17325_;
wire _17326_;
wire _17327_;
wire _17328_;
wire _17329_;
wire _17330_;
wire _17331_;
wire _17332_;
wire _17333_;
wire _17334_;
wire _17335_;
wire _17336_;
wire _17337_;
wire _17338_;
wire _17339_;
wire _17340_;
wire _17341_;
wire _17342_;
wire _17343_;
wire _17344_;
wire _17345_;
wire _17346_;
wire _17347_;
wire _17348_;
wire _17349_;
wire _17350_;
wire _17351_;
wire _17352_;
wire _17353_;
wire _17354_;
wire _17355_;
wire _17356_;
wire _17357_;
wire _17358_;
wire _17359_;
wire _17360_;
wire _17361_;
wire _17362_;
wire _17363_;
wire _17364_;
wire _17365_;
wire _17366_;
wire _17367_;
wire _17368_;
wire _17369_;
wire _17370_;
wire _17371_;
wire _17372_;
wire _17373_;
wire _17374_;
wire _17375_;
wire _17376_;
wire _17377_;
wire _17378_;
wire _17379_;
wire _17380_;
wire _17381_;
wire _17382_;
wire _17383_;
wire _17384_;
wire _17385_;
wire _17386_;
wire _17387_;
wire _17388_;
wire _17389_;
wire _17390_;
wire _17391_;
wire _17392_;
wire _17393_;
wire _17394_;
wire _17395_;
wire _17396_;
wire _17397_;
wire _17398_;
wire _17399_;
wire _17400_;
wire _17401_;
wire _17402_;
wire _17403_;
wire _17404_;
wire _17405_;
wire _17406_;
wire _17407_;
wire _17408_;
wire _17409_;
wire _17410_;
wire _17411_;
wire _17412_;
wire _17413_;
wire _17414_;
wire _17415_;
wire _17416_;
wire _17417_;
wire _17418_;
wire _17419_;
wire _17420_;
wire _17421_;
wire _17422_;
wire _17423_;
wire _17424_;
wire _17425_;
wire _17426_;
wire _17427_;
wire _17428_;
wire _17429_;
wire _17430_;
wire _17431_;
wire _17432_;
wire _17433_;
wire _17434_;
wire _17435_;
wire _17436_;
wire _17437_;
wire _17438_;
wire _17439_;
wire _17440_;
wire _17441_;
wire _17442_;
wire _17443_;
wire _17444_;
wire _17445_;
wire _17446_;
wire _17447_;
wire _17448_;
wire _17449_;
wire _17450_;
wire _17451_;
wire _17452_;
wire _17453_;
wire _17454_;
wire _17455_;
wire _17456_;
wire _17457_;
wire _17458_;
wire _17459_;
wire _17460_;
wire _17461_;
wire _17462_;
wire _17463_;
wire _17464_;
wire _17465_;
wire _17466_;
wire _17467_;
wire _17468_;
wire _17469_;
wire _17470_;
wire _17471_;
wire _17472_;
wire _17473_;
wire _17474_;
wire _17475_;
wire _17476_;
wire _17477_;
wire _17478_;
wire _17479_;
wire _17480_;
wire _17481_;
wire _17482_;
wire _17483_;
wire _17484_;
wire _17485_;
wire _17486_;
wire _17487_;
wire _17488_;
wire _17489_;
wire _17490_;
wire _17491_;
wire _17492_;
wire _17493_;
wire _17494_;
wire _17495_;
wire _17496_;
wire _17497_;
wire _17498_;
wire _17499_;
wire _17500_;
wire _17501_;
wire _17502_;
wire _17503_;
wire _17504_;
wire _17505_;
wire _17506_;
wire _17507_;
wire _17508_;
wire _17509_;
wire _17510_;
wire _17511_;
wire _17512_;
wire _17513_;
wire _17514_;
wire _17515_;
wire _17516_;
wire _17517_;
wire _17518_;
wire _17519_;
wire _17520_;
wire _17521_;
wire _17522_;
wire _17523_;
wire _17524_;
wire _17525_;
wire _17526_;
wire _17527_;
wire _17528_;
wire _17529_;
wire _17530_;
wire _17531_;
wire _17532_;
wire _17533_;
wire _17534_;
wire _17535_;
wire _17536_;
wire _17537_;
wire _17538_;
wire _17539_;
wire _17540_;
wire _17541_;
wire _17542_;
wire _17543_;
wire _17544_;
wire _17545_;
wire _17546_;
wire _17547_;
wire _17548_;
wire _17549_;
wire _17550_;
wire _17551_;
wire _17552_;
wire _17553_;
wire _17554_;
wire _17555_;
wire _17556_;
wire _17557_;
wire _17558_;
wire _17559_;
wire _17560_;
wire _17561_;
wire _17562_;
wire _17563_;
wire _17564_;
wire _17565_;
wire _17566_;
wire _17567_;
wire _17568_;
wire _17569_;
wire _17570_;
wire _17571_;
wire _17572_;
wire _17573_;
wire _17574_;
wire _17575_;
wire _17576_;
wire _17577_;
wire _17578_;
wire _17579_;
wire _17580_;
wire _17581_;
wire _17582_;
wire _17583_;
wire _17584_;
wire _17585_;
wire _17586_;
wire _17587_;
wire _17588_;
wire _17589_;
wire _17590_;
wire _17591_;
wire _17592_;
wire _17593_;
wire _17594_;
wire _17595_;
wire _17596_;
wire _17597_;
wire _17598_;
wire _17599_;
wire _17600_;
wire _17601_;
wire _17602_;
wire _17603_;
wire _17604_;
wire _17605_;
wire _17606_;
wire _17607_;
wire _17608_;
wire _17609_;
wire _17610_;
wire _17611_;
wire _17612_;
wire _17613_;
wire _17614_;
wire _17615_;
wire _17616_;
wire _17617_;
wire _17618_;
wire _17619_;
wire _17620_;
wire _17621_;
wire _17622_;
wire _17623_;
wire _17624_;
wire _17625_;
wire _17626_;
wire _17627_;
wire _17628_;
wire _17629_;
wire _17630_;
wire _17631_;
wire _17632_;
wire _17633_;
wire _17634_;
wire _17635_;
wire _17636_;
wire _17637_;
wire _17638_;
wire _17639_;
wire _17640_;
wire _17641_;
wire _17642_;
wire _17643_;
wire _17644_;
wire _17645_;
wire _17646_;
wire _17647_;
wire _17648_;
wire _17649_;
wire _17650_;
wire _17651_;
wire _17652_;
wire _17653_;
wire _17654_;
wire _17655_;
wire _17656_;
wire _17657_;
wire _17658_;
wire _17659_;
wire _17660_;
wire _17661_;
wire _17662_;
wire _17663_;
wire _17664_;
wire _17665_;
wire _17666_;
wire _17667_;
wire _17668_;
wire _17669_;
wire _17670_;
wire _17671_;
wire _17672_;
wire _17673_;
wire _17674_;
wire _17675_;
wire _17676_;
wire _17677_;
wire _17678_;
wire _17679_;
wire _17680_;
wire _17681_;
wire _17682_;
wire _17683_;
wire _17684_;
wire _17685_;
wire _17686_;
wire _17687_;
wire _17688_;
wire _17689_;
wire _17690_;
wire _17691_;
wire _17692_;
wire _17693_;
wire _17694_;
wire _17695_;
wire _17696_;
wire _17697_;
wire _17698_;
wire _17699_;
wire _17700_;
wire _17701_;
wire _17702_;
wire _17703_;
wire _17704_;
wire _17705_;
wire _17706_;
wire _17707_;
wire _17708_;
wire _17709_;
wire _17710_;
wire _17711_;
wire _17712_;
wire _17713_;
wire _17714_;
wire _17715_;
wire _17716_;
wire _17717_;
wire _17718_;
wire _17719_;
wire _17720_;
wire _17721_;
wire _17722_;
wire _17723_;
wire _17724_;
wire _17725_;
wire _17726_;
wire _17727_;
wire _17728_;
wire _17729_;
wire _17730_;
wire _17731_;
wire _17732_;
wire _17733_;
wire _17734_;
wire _17735_;
wire _17736_;
wire _17737_;
wire _17738_;
wire _17739_;
wire _17740_;
wire _17741_;
wire _17742_;
wire _17743_;
wire _17744_;
wire _17745_;
wire _17746_;
wire _17747_;
wire _17748_;
wire _17749_;
wire _17750_;
wire _17751_;
wire _17752_;
wire _17753_;
wire _17754_;
wire _17755_;
wire _17756_;
wire _17757_;
wire _17758_;
wire _17759_;
wire _17760_;
wire _17761_;
wire _17762_;
wire _17763_;
wire _17764_;
wire _17765_;
wire _17766_;
wire _17767_;
wire _17768_;
wire _17769_;
wire _17770_;
wire _17771_;
wire _17772_;
wire _17773_;
wire _17774_;
wire _17775_;
wire _17776_;
wire _17777_;
wire _17778_;
wire _17779_;
wire _17780_;
wire _17781_;
wire _17782_;
wire _17783_;
wire _17784_;
wire _17785_;
wire _17786_;
wire _17787_;
wire _17788_;
wire _17789_;
wire _17790_;
wire _17791_;
wire _17792_;
wire _17793_;
wire _17794_;
wire _17795_;
wire _17796_;
wire _17797_;
wire _17798_;
wire _17799_;
wire _17800_;
wire _17801_;
wire _17802_;
wire _17803_;
wire _17804_;
wire _17805_;
wire _17806_;
wire _17807_;
wire _17808_;
wire _17809_;
wire _17810_;
wire _17811_;
wire _17812_;
wire _17813_;
wire _17814_;
wire _17815_;
wire _17816_;
wire _17817_;
wire _17818_;
wire _17819_;
wire _17820_;
wire _17821_;
wire _17822_;
wire _17823_;
wire _17824_;
wire _17825_;
wire _17826_;
wire _17827_;
wire _17828_;
wire _17829_;
wire _17830_;
wire _17831_;
wire _17832_;
wire _17833_;
wire _17834_;
wire _17835_;
wire _17836_;
wire _17837_;
wire _17838_;
wire _17839_;
wire _17840_;
wire _17841_;
wire _17842_;
wire _17843_;
wire _17844_;
wire _17845_;
wire _17846_;
wire _17847_;
wire _17848_;
wire _17849_;
wire _17850_;
wire _17851_;
wire _17852_;
wire _17853_;
wire _17854_;
wire _17855_;
wire _17856_;
wire _17857_;
wire _17858_;
wire _17859_;
wire _17860_;
wire _17861_;
wire _17862_;
wire _17863_;
wire _17864_;
wire _17865_;
wire _17866_;
wire _17867_;
wire _17868_;
wire _17869_;
wire _17870_;
wire _17871_;
wire _17872_;
wire _17873_;
wire _17874_;
wire _17875_;
wire _17876_;
wire _17877_;
wire _17878_;
wire _17879_;
wire _17880_;
wire _17881_;
wire _17882_;
wire _17883_;
wire _17884_;
wire _17885_;
wire _17886_;
wire _17887_;
wire _17888_;
wire _17889_;
wire _17890_;
wire _17891_;
wire _17892_;
wire _17893_;
wire _17894_;
wire _17895_;
wire _17896_;
wire _17897_;
wire _17898_;
wire _17899_;
wire _17900_;
wire _17901_;
wire _17902_;
wire _17903_;
wire _17904_;
wire _17905_;
wire _17906_;
wire _17907_;
wire _17908_;
wire _17909_;
wire _17910_;
wire _17911_;
wire _17912_;
wire _17913_;
wire _17914_;
wire _17915_;
wire _17916_;
wire _17917_;
wire _17918_;
wire _17919_;
wire _17920_;
wire _17921_;
wire _17922_;
wire _17923_;
wire _17924_;
wire _17925_;
wire _17926_;
wire _17927_;
wire _17928_;
wire _17929_;
wire _17930_;
wire _17931_;
wire _17932_;
wire _17933_;
wire _17934_;
wire _17935_;
wire _17936_;
wire _17937_;
wire _17938_;
wire _17939_;
wire _17940_;
wire _17941_;
wire _17942_;
wire _17943_;
wire _17944_;
wire _17945_;
wire _17946_;
wire _17947_;
wire _17948_;
wire _17949_;
wire _17950_;
wire _17951_;
wire _17952_;
wire _17953_;
wire _17954_;
wire _17955_;
wire _17956_;
wire _17957_;
wire _17958_;
wire _17959_;
wire _17960_;
wire _17961_;
wire _17962_;
wire _17963_;
wire _17964_;
wire _17965_;
wire _17966_;
wire _17967_;
wire _17968_;
wire _17969_;
wire _17970_;
wire _17971_;
wire _17972_;
wire _17973_;
wire _17974_;
wire _17975_;
wire _17976_;
wire _17977_;
wire _17978_;
wire _17979_;
wire _17980_;
wire _17981_;
wire _17982_;
wire _17983_;
wire _17984_;
wire _17985_;
wire _17986_;
wire _17987_;
wire _17988_;
wire _17989_;
wire _17990_;
wire _17991_;
wire _17992_;
wire _17993_;
wire _17994_;
wire _17995_;
wire _17996_;
wire _17997_;
wire _17998_;
wire _17999_;
wire _18000_;
wire _18001_;
wire _18002_;
wire _18003_;
wire _18004_;
wire _18005_;
wire _18006_;
wire _18007_;
wire _18008_;
wire _18009_;
wire _18010_;
wire _18011_;
wire _18012_;
wire _18013_;
wire _18014_;
wire _18015_;
wire _18016_;
wire _18017_;
wire _18018_;
wire _18019_;
wire _18020_;
wire _18021_;
wire _18022_;
wire _18023_;
wire _18024_;
wire _18025_;
wire _18026_;
wire _18027_;
wire _18028_;
wire _18029_;
wire _18030_;
wire _18031_;
wire _18032_;
wire _18033_;
wire _18034_;
wire _18035_;
wire _18036_;
wire _18037_;
wire _18038_;
wire _18039_;
wire _18040_;
wire _18041_;
wire _18042_;
wire _18043_;
wire _18044_;
wire _18045_;
wire _18046_;
wire _18047_;
wire _18048_;
wire _18049_;
wire _18050_;
wire _18051_;
wire _18052_;
wire _18053_;
wire _18054_;
wire _18055_;
wire _18056_;
wire _18057_;
wire _18058_;
wire _18059_;
wire _18060_;
wire _18061_;
wire _18062_;
wire _18063_;
wire _18064_;
wire _18065_;
wire _18066_;
wire _18067_;
wire _18068_;
wire _18069_;
wire _18070_;
wire _18071_;
wire _18072_;
wire _18073_;
wire _18074_;
wire _18075_;
wire _18076_;
wire _18077_;
wire _18078_;
wire _18079_;
wire _18080_;
wire _18081_;
wire _18082_;
wire _18083_;
wire _18084_;
wire _18085_;
wire _18086_;
wire _18087_;
wire _18088_;
wire _18089_;
wire _18090_;
wire _18091_;
wire _18092_;
wire _18093_;
wire _18094_;
wire _18095_;
wire _18096_;
wire _18097_;
wire _18098_;
wire _18099_;
wire _18100_;
wire _18101_;
wire _18102_;
wire _18103_;
wire _18104_;
wire _18105_;
wire _18106_;
wire _18107_;
wire _18108_;
wire _18109_;
wire _18110_;
wire _18111_;
wire _18112_;
wire _18113_;
wire _18114_;
wire _18115_;
wire _18116_;
wire _18117_;
wire _18118_;
wire _18119_;
wire _18120_;
wire _18121_;
wire _18122_;
wire _18123_;
wire _18124_;
wire _18125_;
wire _18126_;
wire _18127_;
wire _18128_;
wire _18129_;
wire _18130_;
wire _18131_;
wire _18132_;
wire _18133_;
wire _18134_;
wire _18135_;
wire _18136_;
wire _18137_;
wire _18138_;
wire _18139_;
wire _18140_;
wire _18141_;
wire _18142_;
wire _18143_;
wire _18144_;
wire _18145_;
wire _18146_;
wire _18147_;
wire _18148_;
wire _18149_;
wire _18150_;
wire _18151_;
wire _18152_;
wire _18153_;
wire _18154_;
wire _18155_;
wire _18156_;
wire _18157_;
wire _18158_;
wire _18159_;
wire _18160_;
wire _18161_;
wire _18162_;
wire _18163_;
wire _18164_;
wire _18165_;
wire _18166_;
wire _18167_;
wire _18168_;
wire _18169_;
wire _18170_;
wire _18171_;
wire _18172_;
wire _18173_;
wire _18174_;
wire _18175_;
wire _18176_;
wire _18177_;
wire _18178_;
wire _18179_;
wire _18180_;
wire _18181_;
wire _18182_;
wire _18183_;
wire _18184_;
wire _18185_;
wire _18186_;
wire _18187_;
wire _18188_;
wire _18189_;
wire _18190_;
wire _18191_;
wire _18192_;
wire _18193_;
wire _18194_;
wire _18195_;
wire _18196_;
wire _18197_;
wire _18198_;
wire _18199_;
wire _18200_;
wire _18201_;
wire _18202_;
wire _18203_;
wire _18204_;
wire _18205_;
wire _18206_;
wire _18207_;
wire _18208_;
wire _18209_;
wire _18210_;
wire _18211_;
wire _18212_;
wire _18213_;
wire _18214_;
wire _18215_;
wire _18216_;
wire _18217_;
wire _18218_;
wire _18219_;
wire _18220_;
wire _18221_;
wire _18222_;
wire _18223_;
wire _18224_;
wire _18225_;
wire _18226_;
wire _18227_;
wire _18228_;
wire _18229_;
wire _18230_;
wire _18231_;
wire _18232_;
wire _18233_;
wire _18234_;
wire _18235_;
wire _18236_;
wire _18237_;
wire _18238_;
wire _18239_;
wire _18240_;
wire _18241_;
wire _18242_;
wire _18243_;
wire _18244_;
wire _18245_;
wire _18246_;
wire _18247_;
wire _18248_;
wire _18249_;
wire _18250_;
wire _18251_;
wire _18252_;
wire _18253_;
wire _18254_;
wire _18255_;
wire _18256_;
wire _18257_;
wire _18258_;
wire _18259_;
wire _18260_;
wire _18261_;
wire _18262_;
wire _18263_;
wire _18264_;
wire _18265_;
wire _18266_;
wire _18267_;
wire _18268_;
wire _18269_;
wire _18270_;
wire _18271_;
wire _18272_;
wire _18273_;
wire _18274_;
wire _18275_;
wire _18276_;
wire _18277_;
wire _18278_;
wire _18279_;
wire _18280_;
wire _18281_;
wire _18282_;
wire _18283_;
wire _18284_;
wire _18285_;
wire _18286_;
wire _18287_;
wire _18288_;
wire _18289_;
wire _18290_;
wire _18291_;
wire _18292_;
wire _18293_;
wire _18294_;
wire _18295_;
wire _18296_;
wire _18297_;
wire _18298_;
wire _18299_;
wire _18300_;
wire _18301_;
wire _18302_;
wire _18303_;
wire _18304_;
wire _18305_;
wire _18306_;
wire _18307_;
wire _18308_;
wire _18309_;
wire _18310_;
wire _18311_;
wire _18312_;
wire _18313_;
wire _18314_;
wire _18315_;
wire _18316_;
wire _18317_;
wire _18318_;
wire _18319_;
wire _18320_;
wire _18321_;
wire _18322_;
wire _18323_;
wire _18324_;
wire _18325_;
wire _18326_;
wire _18327_;
wire _18328_;
wire _18329_;
wire _18330_;
wire _18331_;
wire _18332_;
wire _18333_;
wire _18334_;
wire _18335_;
wire _18336_;
wire _18337_;
wire _18338_;
wire _18339_;
wire _18340_;
wire _18341_;
wire _18342_;
wire _18343_;
wire _18344_;
wire _18345_;
wire _18346_;
wire _18347_;
wire _18348_;
wire _18349_;
wire _18350_;
wire _18351_;
wire _18352_;
wire _18353_;
wire _18354_;
wire _18355_;
wire _18356_;
wire _18357_;
wire _18358_;
wire _18359_;
wire _18360_;
wire _18361_;
wire _18362_;
wire _18363_;
wire _18364_;
wire _18365_;
wire _18366_;
wire _18367_;
wire _18368_;
wire _18369_;
wire _18370_;
wire _18371_;
wire _18372_;
wire _18373_;
wire _18374_;
wire _18375_;
wire _18376_;
wire _18377_;
wire _18378_;
wire _18379_;
wire _18380_;
wire _18381_;
wire _18382_;
wire _18383_;
wire _18384_;
wire _18385_;
wire _18386_;
wire _18387_;
wire _18388_;
wire _18389_;
wire _18390_;
wire _18391_;
wire _18392_;
wire _18393_;
wire _18394_;
wire _18395_;
wire _18396_;
wire _18397_;
wire _18398_;
wire _18399_;
wire _18400_;
wire _18401_;
wire _18402_;
wire _18403_;
wire _18404_;
wire _18405_;
wire _18406_;
wire _18407_;
wire _18408_;
wire _18409_;
wire _18410_;
wire _18411_;
wire _18412_;
wire _18413_;
wire _18414_;
wire _18415_;
wire _18416_;
wire _18417_;
wire _18418_;
wire _18419_;
wire _18420_;
wire _18421_;
wire _18422_;
wire _18423_;
wire _18424_;
wire _18425_;
wire _18426_;
wire _18427_;
wire _18428_;
wire _18429_;
wire _18430_;
wire _18431_;
wire _18432_;
wire _18433_;
wire _18434_;
wire _18435_;
wire _18436_;
wire _18437_;
wire _18438_;
wire _18439_;
wire _18440_;
wire _18441_;
wire _18442_;
wire _18443_;
wire _18444_;
wire _18445_;
wire _18446_;
wire _18447_;
wire _18448_;
wire _18449_;
wire _18450_;
wire _18451_;
wire _18452_;
wire _18453_;
wire _18454_;
wire _18455_;
wire _18456_;
wire _18457_;
wire _18458_;
wire _18459_;
wire _18460_;
wire _18461_;
wire _18462_;
wire _18463_;
wire _18464_;
wire _18465_;
wire _18466_;
wire _18467_;
wire _18468_;
wire _18469_;
wire _18470_;
wire _18471_;
wire _18472_;
wire _18473_;
wire _18474_;
wire _18475_;
wire _18476_;
wire _18477_;
wire _18478_;
wire _18479_;
wire _18480_;
wire _18481_;
wire _18482_;
wire _18483_;
wire _18484_;
wire _18485_;
wire _18486_;
wire _18487_;
wire _18488_;
wire _18489_;
wire _18490_;
wire _18491_;
wire _18492_;
wire _18493_;
wire _18494_;
wire _18495_;
wire _18496_;
wire _18497_;
wire _18498_;
wire _18499_;
wire _18500_;
wire _18501_;
wire _18502_;
wire _18503_;
wire _18504_;
wire _18505_;
wire _18506_;
wire _18507_;
wire _18508_;
wire _18509_;
wire _18510_;
wire _18511_;
wire _18512_;
wire _18513_;
wire _18514_;
wire _18515_;
wire _18516_;
wire _18517_;
wire _18518_;
wire _18519_;
wire _18520_;
wire _18521_;
wire _18522_;
wire _18523_;
wire _18524_;
wire _18525_;
wire _18526_;
wire _18527_;
wire _18528_;
wire _18529_;
wire _18530_;
wire _18531_;
wire _18532_;
wire _18533_;
wire _18534_;
wire _18535_;
wire _18536_;
wire _18537_;
wire _18538_;
wire _18539_;
wire _18540_;
wire _18541_;
wire _18542_;
wire _18543_;
wire _18544_;
wire _18545_;
wire _18546_;
wire _18547_;
wire _18548_;
wire _18549_;
wire _18550_;
wire _18551_;
wire _18552_;
wire _18553_;
wire _18554_;
wire _18555_;
wire _18556_;
wire _18557_;
wire _18558_;
wire _18559_;
wire _18560_;
wire _18561_;
wire _18562_;
wire _18563_;
wire _18564_;
wire _18565_;
wire _18566_;
wire _18567_;
wire _18568_;
wire _18569_;
wire _18570_;
wire _18571_;
wire _18572_;
wire _18573_;
wire _18574_;
wire _18575_;
wire _18576_;
wire _18577_;
wire _18578_;
wire _18579_;
wire _18580_;
wire _18581_;
wire _18582_;
wire _18583_;
wire _18584_;
wire _18585_;
wire _18586_;
wire _18587_;
wire _18588_;
wire _18589_;
wire _18590_;
wire _18591_;
wire _18592_;
wire _18593_;
wire _18594_;
wire _18595_;
wire _18596_;
wire _18597_;
wire _18598_;
wire _18599_;
wire _18600_;
wire _18601_;
wire _18602_;
wire _18603_;
wire _18604_;
wire _18605_;
wire _18606_;
wire _18607_;
wire _18608_;
wire _18609_;
wire _18610_;
wire _18611_;
wire _18612_;
wire _18613_;
wire _18614_;
wire _18615_;
wire _18616_;
wire _18617_;
wire _18618_;
wire _18619_;
wire _18620_;
wire _18621_;
wire _18622_;
wire _18623_;
wire _18624_;
wire _18625_;
wire _18626_;
wire _18627_;
wire _18628_;
wire _18629_;
wire _18630_;
wire _18631_;
wire _18632_;
wire _18633_;
wire _18634_;
wire _18635_;
wire _18636_;
wire _18637_;
wire _18638_;
wire _18639_;
wire _18640_;
wire _18641_;
wire _18642_;
wire _18643_;
wire _18644_;
wire _18645_;
wire _18646_;
wire _18647_;
wire _18648_;
wire _18649_;
wire _18650_;
wire _18651_;
wire _18652_;
wire _18653_;
wire _18654_;
wire _18655_;
wire _18656_;
wire _18657_;
wire _18658_;
wire _18659_;
wire _18660_;
wire _18661_;
wire _18662_;
wire _18663_;
wire _18664_;
wire _18665_;
wire _18666_;
wire _18667_;
wire _18668_;
wire _18669_;
wire _18670_;
wire _18671_;
wire _18672_;
wire _18673_;
wire _18674_;
wire _18675_;
wire _18676_;
wire _18677_;
wire _18678_;
wire _18679_;
wire _18680_;
wire _18681_;
wire _18682_;
wire _18683_;
wire _18684_;
wire _18685_;
wire _18686_;
wire _18687_;
wire _18688_;
wire _18689_;
wire _18690_;
wire _18691_;
wire _18692_;
wire _18693_;
wire _18694_;
wire _18695_;
wire _18696_;
wire _18697_;
wire _18698_;
wire _18699_;
wire _18700_;
wire _18701_;
wire _18702_;
wire _18703_;
wire _18704_;
wire _18705_;
wire _18706_;
wire _18707_;
wire _18708_;
wire _18709_;
wire _18710_;
wire _18711_;
wire _18712_;
wire _18713_;
wire _18714_;
wire _18715_;
wire _18716_;
wire _18717_;
wire _18718_;
wire _18719_;
wire _18720_;
wire _18721_;
wire _18722_;
wire _18723_;
wire _18724_;
wire _18725_;
wire _18726_;
wire _18727_;
wire _18728_;
wire _18729_;
wire _18730_;
wire _18731_;
wire _18732_;
wire _18733_;
wire _18734_;
wire _18735_;
wire _18736_;
wire _18737_;
wire _18738_;
wire _18739_;
wire _18740_;
wire _18741_;
wire _18742_;
wire _18743_;
wire _18744_;
wire _18745_;
wire _18746_;
wire _18747_;
wire _18748_;
wire _18749_;
wire _18750_;
wire _18751_;
wire _18752_;
wire _18753_;
wire _18754_;
wire _18755_;
wire _18756_;
wire _18757_;
wire _18758_;
wire _18759_;
wire _18760_;
wire _18761_;
wire _18762_;
wire _18763_;
wire _18764_;
wire _18765_;
wire _18766_;
wire _18767_;
wire _18768_;
wire _18769_;
wire _18770_;
wire _18771_;
wire _18772_;
wire _18773_;
wire _18774_;
wire _18775_;
wire _18776_;
wire _18777_;
wire _18778_;
wire _18779_;
wire _18780_;
wire _18781_;
wire _18782_;
wire _18783_;
wire _18784_;
wire _18785_;
wire _18786_;
wire _18787_;
wire _18788_;
wire _18789_;
wire _18790_;
wire _18791_;
wire _18792_;
wire _18793_;
wire _18794_;
wire _18795_;
wire _18796_;
wire _18797_;
wire _18798_;
wire _18799_;
wire _18800_;
wire _18801_;
wire _18802_;
wire _18803_;
wire _18804_;
wire _18805_;
wire _18806_;
wire _18807_;
wire _18808_;
wire _18809_;
wire _18810_;
wire _18811_;
wire _18812_;
wire _18813_;
wire _18814_;
wire _18815_;
wire _18816_;
wire _18817_;
wire _18818_;
wire _18819_;
wire _18820_;
wire _18821_;
wire _18822_;
wire _18823_;
wire _18824_;
wire _18825_;
wire _18826_;
wire _18827_;
wire _18828_;
wire _18829_;
wire _18830_;
wire _18831_;
wire _18832_;
wire _18833_;
wire _18834_;
wire _18835_;
wire _18836_;
wire _18837_;
wire _18838_;
wire _18839_;
wire _18840_;
wire _18841_;
wire _18842_;
wire _18843_;
wire _18844_;
wire _18845_;
wire _18846_;
wire _18847_;
wire _18848_;
wire _18849_;
wire _18850_;
wire _18851_;
wire _18852_;
wire _18853_;
wire _18854_;
wire _18855_;
wire _18856_;
wire _18857_;
wire _18858_;
wire _18859_;
wire _18860_;
wire _18861_;
wire _18862_;
wire _18863_;
wire _18864_;
wire _18865_;
wire _18866_;
wire _18867_;
wire _18868_;
wire _18869_;
wire _18870_;
wire _18871_;
wire _18872_;
wire _18873_;
wire _18874_;
wire _18875_;
wire _18876_;
wire _18877_;
wire _18878_;
wire _18879_;
wire _18880_;
wire _18881_;
wire _18882_;
wire _18883_;
wire _18884_;
wire _18885_;
wire _18886_;
wire _18887_;
wire _18888_;
wire _18889_;
wire _18890_;
wire _18891_;
wire _18892_;
wire _18893_;
wire _18894_;
wire _18895_;
wire _18896_;
wire _18897_;
wire _18898_;
wire _18899_;
wire _18900_;
wire _18901_;
wire _18902_;
wire _18903_;
wire _18904_;
wire _18905_;
wire _18906_;
wire _18907_;
wire _18908_;
wire _18909_;
wire _18910_;
wire _18911_;
wire _18912_;
wire _18913_;
wire _18914_;
wire _18915_;
wire _18916_;
wire _18917_;
wire _18918_;
wire _18919_;
wire _18920_;
wire _18921_;
wire _18922_;
wire _18923_;
wire _18924_;
wire _18925_;
wire _18926_;
wire _18927_;
wire _18928_;
wire _18929_;
wire _18930_;
wire _18931_;
wire _18932_;
wire _18933_;
wire _18934_;
wire _18935_;
wire _18936_;
wire _18937_;
wire _18938_;
wire _18939_;
wire _18940_;
wire _18941_;
wire _18942_;
wire _18943_;
wire _18944_;
wire _18945_;
wire _18946_;
wire _18947_;
wire _18948_;
wire _18949_;
wire _18950_;
wire _18951_;
wire _18952_;
wire _18953_;
wire _18954_;
wire _18955_;
wire _18956_;
wire _18957_;
wire _18958_;
wire _18959_;
wire _18960_;
wire _18961_;
wire _18962_;
wire _18963_;
wire _18964_;
wire _18965_;
wire _18966_;
wire _18967_;
wire _18968_;
wire _18969_;
wire _18970_;
wire _18971_;
wire _18972_;
wire _18973_;
wire _18974_;
wire _18975_;
wire _18976_;
wire _18977_;
wire _18978_;
wire _18979_;
wire _18980_;
wire _18981_;
wire _18982_;
wire _18983_;
wire _18984_;
wire _18985_;
wire _18986_;
wire _18987_;
wire _18988_;
wire _18989_;
wire _18990_;
wire _18991_;
wire _18992_;
wire _18993_;
wire _18994_;
wire _18995_;
wire _18996_;
wire _18997_;
wire _18998_;
wire _18999_;
wire _19000_;
wire _19001_;
wire _19002_;
wire _19003_;
wire _19004_;
wire _19005_;
wire _19006_;
wire _19007_;
wire _19008_;
wire _19009_;
wire _19010_;
wire _19011_;
wire _19012_;
wire _19013_;
wire _19014_;
wire _19015_;
wire _19016_;
wire _19017_;
wire _19018_;
wire _19019_;
wire _19020_;
wire _19021_;
wire _19022_;
wire _19023_;
wire _19024_;
wire _19025_;
wire _19026_;
wire _19027_;
wire _19028_;
wire _19029_;
wire _19030_;
wire _19031_;
wire _19032_;
wire _19033_;
wire _19034_;
wire _19035_;
wire _19036_;
wire _19037_;
wire _19038_;
wire _19039_;
wire _19040_;
wire _19041_;
wire _19042_;
wire _19043_;
wire _19044_;
wire _19045_;
wire _19046_;
wire _19047_;
wire _19048_;
wire _19049_;
wire _19050_;
wire _19051_;
wire _19052_;
wire _19053_;
wire _19054_;
wire _19055_;
wire _19056_;
wire _19057_;
wire _19058_;
wire _19059_;
wire _19060_;
wire _19061_;
wire _19062_;
wire _19063_;
wire _19064_;
wire _19065_;
wire _19066_;
wire _19067_;
wire _19068_;
wire _19069_;
wire _19070_;
wire _19071_;
wire _19072_;
wire _19073_;
wire _19074_;
wire _19075_;
wire _19076_;
wire _19077_;
wire _19078_;
wire _19079_;
wire _19080_;
wire _19081_;
wire _19082_;
wire _19083_;
wire _19084_;
wire _19085_;
wire _19086_;
wire _19087_;
wire _19088_;
wire _19089_;
wire _19090_;
wire _19091_;
wire _19092_;
wire _19093_;
wire _19094_;
wire _19095_;
wire _19096_;
wire _19097_;
wire _19098_;
wire _19099_;
wire _19100_;
wire _19101_;
wire _19102_;
wire _19103_;
wire _19104_;
wire _19105_;
wire _19106_;
wire _19107_;
wire _19108_;
wire _19109_;
wire _19110_;
wire _19111_;
wire _19112_;
wire _19113_;
wire _19114_;
wire _19115_;
wire _19116_;
wire _19117_;
wire _19118_;
wire _19119_;
wire _19120_;
wire _19121_;
wire _19122_;
wire _19123_;
wire _19124_;
wire _19125_;
wire _19126_;
wire _19127_;
wire _19128_;
wire _19129_;
wire _19130_;
wire _19131_;
wire _19132_;
wire _19133_;
wire _19134_;
wire _19135_;
wire _19136_;
wire _19137_;
wire _19138_;
wire _19139_;
wire _19140_;
wire _19141_;
wire _19142_;
wire _19143_;
wire _19144_;
wire _19145_;
wire _19146_;
wire _19147_;
wire _19148_;
wire _19149_;
wire _19150_;
wire _19151_;
wire _19152_;
wire _19153_;
wire _19154_;
wire _19155_;
wire _19156_;
wire _19157_;
wire _19158_;
wire _19159_;
wire _19160_;
wire _19161_;
wire _19162_;
wire _19163_;
wire _19164_;
wire _19165_;
wire _19166_;
wire _19167_;
wire _19168_;
wire _19169_;
wire _19170_;
wire _19171_;
wire _19172_;
wire _19173_;
wire _19174_;
wire _19175_;
wire _19176_;
wire _19177_;
wire _19178_;
wire _19179_;
wire _19180_;
wire _19181_;
wire _19182_;
wire _19183_;
wire _19184_;
wire _19185_;
wire _19186_;
wire _19187_;
wire _19188_;
wire _19189_;
wire _19190_;
wire _19191_;
wire _19192_;
wire _19193_;
wire _19194_;
wire _19195_;
wire _19196_;
wire _19197_;
wire _19198_;
wire _19199_;
wire _19200_;
wire _19201_;
wire _19202_;
wire _19203_;
wire _19204_;
wire _19205_;
wire _19206_;
wire _19207_;
wire _19208_;
wire _19209_;
wire _19210_;
wire _19211_;
wire _19212_;
wire _19213_;
wire _19214_;
wire _19215_;
wire _19216_;
wire _19217_;
wire _19218_;
wire _19219_;
wire _19220_;
wire _19221_;
wire _19222_;
wire _19223_;
wire _19224_;
wire _19225_;
wire _19226_;
wire _19227_;
wire _19228_;
wire _19229_;
wire _19230_;
wire _19231_;
wire _19232_;
wire _19233_;
wire _19234_;
wire _19235_;
wire _19236_;
wire _19237_;
wire _19238_;
wire _19239_;
wire _19240_;
wire _19241_;
wire _19242_;
wire _19243_;
wire _19244_;
wire _19245_;
wire _19246_;
wire _19247_;
wire _19248_;
wire _19249_;
wire _19250_;
wire _19251_;
wire _19252_;
wire _19253_;
wire _19254_;
wire _19255_;
wire _19256_;
wire _19257_;
wire _19258_;
wire _19259_;
wire _19260_;
wire _19261_;
wire _19262_;
wire _19263_;
wire _19264_;
wire _19265_;
wire _19266_;
wire _19267_;
wire _19268_;
wire _19269_;
wire _19270_;
wire _19271_;
wire _19272_;
wire _19273_;
wire _19274_;
wire _19275_;
wire _19276_;
wire _19277_;
wire _19278_;
wire _19279_;
wire _19280_;
wire _19281_;
wire _19282_;
wire _19283_;
wire _19284_;
wire _19285_;
wire _19286_;
wire _19287_;
wire _19288_;
wire _19289_;
wire _19290_;
wire _19291_;
wire _19292_;
wire _19293_;
wire _19294_;
wire _19295_;
wire _19296_;
wire _19297_;
wire _19298_;
wire _19299_;
wire _19300_;
wire _19301_;
wire _19302_;
wire _19303_;
wire _19304_;
wire _19305_;
wire _19306_;
wire _19307_;
wire _19308_;
wire _19309_;
wire _19310_;
wire _19311_;
wire _19312_;
wire _19313_;
wire _19314_;
wire _19315_;
wire _19316_;
wire _19317_;
wire _19318_;
wire _19319_;
wire _19320_;
wire _19321_;
wire _19322_;
wire _19323_;
wire _19324_;
wire _19325_;
wire _19326_;
wire _19327_;
wire _19328_;
wire _19329_;
wire _19330_;
wire _19331_;
wire _19332_;
wire _19333_;
wire _19334_;
wire _19335_;
wire _19336_;
wire _19337_;
wire _19338_;
wire _19339_;
wire _19340_;
wire _19341_;
wire _19342_;
wire _19343_;
wire _19344_;
wire _19345_;
wire _19346_;
wire _19347_;
wire _19348_;
wire _19349_;
wire _19350_;
wire _19351_;
wire _19352_;
wire _19353_;
wire _19354_;
wire _19355_;
wire _19356_;
wire _19357_;
wire _19358_;
wire _19359_;
wire _19360_;
wire _19361_;
wire _19362_;
wire _19363_;
wire _19364_;
wire _19365_;
wire _19366_;
wire _19367_;
wire _19368_;
wire _19369_;
wire _19370_;
wire _19371_;
wire _19372_;
wire _19373_;
wire _19374_;
wire _19375_;
wire _19376_;
wire _19377_;
wire _19378_;
wire _19379_;
wire _19380_;
wire _19381_;
wire _19382_;
wire _19383_;
wire _19384_;
wire _19385_;
wire _19386_;
wire _19387_;
wire _19388_;
wire _19389_;
wire _19390_;
wire _19391_;
wire _19392_;
wire _19393_;
wire _19394_;
wire _19395_;
wire _19396_;
wire _19397_;
wire _19398_;
wire _19399_;
wire _19400_;
wire _19401_;
wire _19402_;
wire _19403_;
wire _19404_;
wire _19405_;
wire _19406_;
wire _19407_;
wire _19408_;
wire _19409_;
wire _19410_;
wire _19411_;
wire _19412_;
wire _19413_;
wire _19414_;
wire _19415_;
wire _19416_;
wire _19417_;
wire _19418_;
wire _19419_;
wire _19420_;
wire _19421_;
wire _19422_;
wire _19423_;
wire _19424_;
wire _19425_;
wire _19426_;
wire _19427_;
wire _19428_;
wire _19429_;
wire _19430_;
wire _19431_;
wire _19432_;
wire _19433_;
wire _19434_;
wire _19435_;
wire _19436_;
wire _19437_;
wire _19438_;
wire _19439_;
wire _19440_;
wire _19441_;
wire _19442_;
wire _19443_;
wire _19444_;
wire _19445_;
wire _19446_;
wire _19447_;
wire _19448_;
wire _19449_;
wire _19450_;
wire _19451_;
wire _19452_;
wire _19453_;
wire _19454_;
wire _19455_;
wire _19456_;
wire _19457_;
wire _19458_;
wire _19459_;
wire _19460_;
wire _19461_;
wire _19462_;
wire _19463_;
wire _19464_;
wire _19465_;
wire _19466_;
wire _19467_;
wire _19468_;
wire _19469_;
wire _19470_;
wire _19471_;
wire _19472_;
wire _19473_;
wire _19474_;
wire _19475_;
wire _19476_;
wire _19477_;
wire _19478_;
wire _19479_;
wire _19480_;
wire _19481_;
wire _19482_;
wire _19483_;
wire _19484_;
wire _19485_;
wire _19486_;
wire _19487_;
wire _19488_;
wire _19489_;
wire _19490_;
wire _19491_;
wire _19492_;
wire _19493_;
wire _19494_;
wire _19495_;
wire _19496_;
wire _19497_;
wire _19498_;
wire _19499_;
wire _19500_;
wire _19501_;
wire _19502_;
wire _19503_;
wire _19504_;
wire _19505_;
wire _19506_;
wire _19507_;
wire _19508_;
wire _19509_;
wire _19510_;
wire _19511_;
wire _19512_;
wire _19513_;
wire _19514_;
wire _19515_;
wire _19516_;
wire _19517_;
wire _19518_;
wire _19519_;
wire _19520_;
wire _19521_;
wire _19522_;
wire _19523_;
wire _19524_;
wire _19525_;
wire _19526_;
wire _19527_;
wire _19528_;
wire _19529_;
wire _19530_;
wire _19531_;
wire _19532_;
wire _19533_;
wire _19534_;
wire _19535_;
wire _19536_;
wire _19537_;
wire _19538_;
wire _19539_;
wire _19540_;
wire _19541_;
wire _19542_;
wire _19543_;
wire _19544_;
wire _19545_;
wire _19546_;
wire _19547_;
wire _19548_;
wire _19549_;
wire _19550_;
wire _19551_;
wire _19552_;
wire _19553_;
wire _19554_;
wire _19555_;
wire _19556_;
wire _19557_;
wire _19558_;
wire _19559_;
wire _19560_;
wire _19561_;
wire _19562_;
wire _19563_;
wire _19564_;
wire _19565_;
wire _19566_;
wire _19567_;
wire _19568_;
wire _19569_;
wire _19570_;
wire _19571_;
wire _19572_;
wire _19573_;
wire _19574_;
wire _19575_;
wire _19576_;
wire _19577_;
wire _19578_;
wire _19579_;
wire _19580_;
wire _19581_;
wire _19582_;
wire _19583_;
wire _19584_;
wire _19585_;
wire _19586_;
wire _19587_;
wire _19588_;
wire _19589_;
wire _19590_;
wire _19591_;
wire _19592_;
wire _19593_;
wire _19594_;
wire _19595_;
wire _19596_;
wire _19597_;
wire _19598_;
wire _19599_;
wire _19600_;
wire _19601_;
wire _19602_;
wire _19603_;
wire _19604_;
wire _19605_;
wire _19606_;
wire _19607_;
wire _19608_;
wire _19609_;
wire _19610_;
wire _19611_;
wire _19612_;
wire _19613_;
wire _19614_;
wire _19615_;
wire _19616_;
wire _19617_;
wire _19618_;
wire _19619_;
wire _19620_;
wire _19621_;
wire _19622_;
wire _19623_;
wire _19624_;
wire _19625_;
wire _19626_;
wire _19627_;
wire _19628_;
wire _19629_;
wire _19630_;
wire _19631_;
wire _19632_;
wire _19633_;
wire _19634_;
wire _19635_;
wire _19636_;
wire _19637_;
wire _19638_;
wire _19639_;
wire _19640_;
wire _19641_;
wire _19642_;
wire _19643_;
wire _19644_;
wire _19645_;
wire _19646_;
wire _19647_;
wire _19648_;
wire _19649_;
wire _19650_;
wire _19651_;
wire _19652_;
wire _19653_;
wire _19654_;
wire _19655_;
wire _19656_;
wire _19657_;
wire _19658_;
wire _19659_;
wire _19660_;
wire _19661_;
wire _19662_;
wire _19663_;
wire _19664_;
wire _19665_;
wire _19666_;
wire _19667_;
wire _19668_;
wire _19669_;
wire _19670_;
wire _19671_;
wire _19672_;
wire _19673_;
wire _19674_;
wire _19675_;
wire _19676_;
wire _19677_;
wire _19678_;
wire _19679_;
wire _19680_;
wire _19681_;
wire _19682_;
wire _19683_;
wire _19684_;
wire _19685_;
wire _19686_;
wire _19687_;
wire _19688_;
wire _19689_;
wire _19690_;
wire _19691_;
wire _19692_;
wire _19693_;
wire _19694_;
wire _19695_;
wire _19696_;
wire _19697_;
wire _19698_;
wire _19699_;
wire _19700_;
wire _19701_;
wire _19702_;
wire _19703_;
wire _19704_;
wire _19705_;
wire _19706_;
wire _19707_;
wire _19708_;
wire _19709_;
wire _19710_;
wire _19711_;
wire _19712_;
wire _19713_;
wire _19714_;
wire _19715_;
wire _19716_;
wire _19717_;
wire _19718_;
wire _19719_;
wire _19720_;
wire _19721_;
wire _19722_;
wire _19723_;
wire _19724_;
wire _19725_;
wire _19726_;
wire _19727_;
wire _19728_;
wire _19729_;
wire _19730_;
wire _19731_;
wire _19732_;
wire _19733_;
wire _19734_;
wire _19735_;
wire _19736_;
wire _19737_;
wire _19738_;
wire _19739_;
wire _19740_;
wire _19741_;
wire _19742_;
wire _19743_;
wire _19744_;
wire _19745_;
wire _19746_;
wire _19747_;
wire _19748_;
wire _19749_;
wire _19750_;
wire _19751_;
wire _19752_;
wire _19753_;
wire _19754_;
wire _19755_;
wire _19756_;
wire _19757_;
wire _19758_;
wire _19759_;
wire _19760_;
wire _19761_;
wire _19762_;
wire _19763_;
wire _19764_;
wire _19765_;
wire _19766_;
wire _19767_;
wire _19768_;
wire _19769_;
wire _19770_;
wire _19771_;
wire _19772_;
wire _19773_;
wire _19774_;
wire _19775_;
wire _19776_;
wire _19777_;
wire _19778_;
wire _19779_;
wire _19780_;
wire _19781_;
wire _19782_;
wire _19783_;
wire _19784_;
wire _19785_;
wire _19786_;
wire _19787_;
wire _19788_;
wire _19789_;
wire _19790_;
wire _19791_;
wire _19792_;
wire _19793_;
wire _19794_;
wire _19795_;
wire _19796_;
wire _19797_;
wire _19798_;
wire _19799_;
wire _19800_;
wire _19801_;
wire _19802_;
wire _19803_;
wire _19804_;
wire _19805_;
wire _19806_;
wire _19807_;
wire _19808_;
wire _19809_;
wire _19810_;
wire _19811_;
wire _19812_;
wire _19813_;
wire _19814_;
wire _19815_;
wire _19816_;
wire _19817_;
wire _19818_;
wire _19819_;
wire _19820_;
wire _19821_;
wire _19822_;
wire _19823_;
wire _19824_;
wire _19825_;
wire _19826_;
wire _19827_;
wire _19828_;
wire _19829_;
wire _19830_;
wire _19831_;
wire _19832_;
wire _19833_;
wire _19834_;
wire _19835_;
wire _19836_;
wire _19837_;
wire _19838_;
wire _19839_;
wire _19840_;
wire _19841_;
wire _19842_;
wire _19843_;
wire _19844_;
wire _19845_;
wire _19846_;
wire _19847_;
wire _19848_;
wire _19849_;
wire _19850_;
wire _19851_;
wire _19852_;
wire _19853_;
wire _19854_;
wire _19855_;
wire _19856_;
wire _19857_;
wire _19858_;
wire _19859_;
wire _19860_;
wire _19861_;
wire _19862_;
wire _19863_;
wire _19864_;
wire _19865_;
wire _19866_;
wire _19867_;
wire _19868_;
wire _19869_;
wire _19870_;
wire _19871_;
wire _19872_;
wire _19873_;
wire _19874_;
wire _19875_;
wire _19876_;
wire _19877_;
wire _19878_;
wire _19879_;
wire _19880_;
wire _19881_;
wire _19882_;
wire _19883_;
wire _19884_;
wire _19885_;
wire _19886_;
wire _19887_;
wire _19888_;
wire _19889_;
wire _19890_;
wire _19891_;
wire _19892_;
wire _19893_;
wire _19894_;
wire _19895_;
wire _19896_;
wire _19897_;
wire _19898_;
wire _19899_;
wire _19900_;
wire _19901_;
wire _19902_;
wire _19903_;
wire _19904_;
wire _19905_;
wire _19906_;
wire _19907_;
wire _19908_;
wire _19909_;
wire _19910_;
wire _19911_;
wire _19912_;
wire _19913_;
wire _19914_;
wire _19915_;
wire _19916_;
wire _19917_;
wire _19918_;
wire _19919_;
wire _19920_;
wire _19921_;
wire _19922_;
wire _19923_;
wire _19924_;
wire _19925_;
wire _19926_;
wire _19927_;
wire _19928_;
wire _19929_;
wire _19930_;
wire _19931_;
wire _19932_;
wire _19933_;
wire _19934_;
wire _19935_;
wire _19936_;
wire _19937_;
wire _19938_;
wire _19939_;
wire _19940_;
wire _19941_;
wire _19942_;
wire _19943_;
wire _19944_;
wire _19945_;
wire _19946_;
wire _19947_;
wire _19948_;
wire _19949_;
wire _19950_;
wire _19951_;
wire _19952_;
wire _19953_;
wire _19954_;
wire _19955_;
wire _19956_;
wire _19957_;
wire _19958_;
wire _19959_;
wire _19960_;
wire _19961_;
wire _19962_;
wire _19963_;
wire _19964_;
wire _19965_;
wire _19966_;
wire _19967_;
wire _19968_;
wire _19969_;
wire _19970_;
wire _19971_;
wire _19972_;
wire _19973_;
wire _19974_;
wire _19975_;
wire _19976_;
wire _19977_;
wire _19978_;
wire _19979_;
wire _19980_;
wire _19981_;
wire _19982_;
wire _19983_;
wire _19984_;
wire _19985_;
wire _19986_;
wire _19987_;
wire _19988_;
wire _19989_;
wire _19990_;
wire _19991_;
wire _19992_;
wire _19993_;
wire _19994_;
wire _19995_;
wire _19996_;
wire _19997_;
wire _19998_;
wire _19999_;
wire _20000_;
wire _20001_;
wire _20002_;
wire _20003_;
wire _20004_;
wire _20005_;
wire _20006_;
wire _20007_;
wire _20008_;
wire _20009_;
wire _20010_;
wire _20011_;
wire _20012_;
wire _20013_;
wire _20014_;
wire _20015_;
wire _20016_;
wire _20017_;
wire _20018_;
wire _20019_;
wire _20020_;
wire _20021_;
wire _20022_;
wire _20023_;
wire _20024_;
wire _20025_;
wire _20026_;
wire _20027_;
wire _20028_;
wire _20029_;
wire _20030_;
wire _20031_;
wire _20032_;
wire _20033_;
wire _20034_;
wire _20035_;
wire _20036_;
wire _20037_;
wire _20038_;
wire _20039_;
wire _20040_;
wire _20041_;
wire _20042_;
wire _20043_;
wire _20044_;
wire _20045_;
wire _20046_;
wire _20047_;
wire _20048_;
wire _20049_;
wire _20050_;
wire _20051_;
wire _20052_;
wire _20053_;
wire _20054_;
wire _20055_;
wire _20056_;
wire _20057_;
wire _20058_;
wire _20059_;
wire _20060_;
wire _20061_;
wire _20062_;
wire _20063_;
wire _20064_;
wire _20065_;
wire _20066_;
wire _20067_;
wire _20068_;
wire _20069_;
wire _20070_;
wire _20071_;
wire _20072_;
wire _20073_;
wire _20074_;
wire _20075_;
wire _20076_;
wire _20077_;
wire _20078_;
wire _20079_;
wire _20080_;
wire _20081_;
wire _20082_;
wire _20083_;
wire _20084_;
wire _20085_;
wire _20086_;
wire _20087_;
wire _20088_;
wire _20089_;
wire _20090_;
wire _20091_;
wire _20092_;
wire _20093_;
wire _20094_;
wire _20095_;
wire _20096_;
wire _20097_;
wire _20098_;
wire _20099_;
wire _20100_;
wire _20101_;
wire _20102_;
wire _20103_;
wire _20104_;
wire _20105_;
wire _20106_;
wire _20107_;
wire _20108_;
wire _20109_;
wire _20110_;
wire _20111_;
wire _20112_;
wire _20113_;
wire _20114_;
wire _20115_;
wire _20116_;
wire _20117_;
wire _20118_;
wire _20119_;
wire _20120_;
wire _20121_;
wire _20122_;
wire _20123_;
wire _20124_;
wire _20125_;
wire _20126_;
wire _20127_;
wire _20128_;
wire _20129_;
wire _20130_;
wire _20131_;
wire _20132_;
wire _20133_;
wire _20134_;
wire _20135_;
wire _20136_;
wire _20137_;
wire _20138_;
wire _20139_;
wire _20140_;
wire _20141_;
wire _20142_;
wire _20143_;
wire _20144_;
wire _20145_;
wire _20146_;
wire _20147_;
wire _20148_;
wire _20149_;
wire _20150_;
wire _20151_;
wire _20152_;
wire _20153_;
wire _20154_;
wire _20155_;
wire _20156_;
wire _20157_;
wire _20158_;
wire _20159_;
wire _20160_;
wire _20161_;
wire _20162_;
wire _20163_;
wire _20164_;
wire _20165_;
wire _20166_;
wire _20167_;
wire _20168_;
wire _20169_;
wire _20170_;
wire _20171_;
wire _20172_;
wire _20173_;
wire _20174_;
wire _20175_;
wire _20176_;
wire _20177_;
wire _20178_;
wire _20179_;
wire _20180_;
wire _20181_;
wire _20182_;
wire _20183_;
wire _20184_;
wire _20185_;
wire _20186_;
wire _20187_;
wire _20188_;
wire _20189_;
wire _20190_;
wire _20191_;
wire _20192_;
wire _20193_;
wire _20194_;
wire _20195_;
wire _20196_;
wire _20197_;
wire _20198_;
wire _20199_;
wire _20200_;
wire _20201_;
wire _20202_;
wire _20203_;
wire _20204_;
wire _20205_;
wire _20206_;
wire _20207_;
wire _20208_;
wire _20209_;
wire _20210_;
wire _20211_;
wire _20212_;
wire _20213_;
wire _20214_;
wire _20215_;
wire _20216_;
wire _20217_;
wire _20218_;
wire _20219_;
wire _20220_;
wire _20221_;
wire _20222_;
wire _20223_;
wire _20224_;
wire _20225_;
wire _20226_;
wire _20227_;
wire _20228_;
wire _20229_;
wire _20230_;
wire _20231_;
wire _20232_;
wire _20233_;
wire _20234_;
wire _20235_;
wire _20236_;
wire _20237_;
wire _20238_;
wire _20239_;
wire _20240_;
wire _20241_;
wire _20242_;
wire _20243_;
wire _20244_;
wire _20245_;
wire _20246_;
wire _20247_;
wire _20248_;
wire _20249_;
wire _20250_;
wire _20251_;
wire _20252_;
wire _20253_;
wire _20254_;
wire _20255_;
wire _20256_;
wire _20257_;
wire _20258_;
wire _20259_;
wire _20260_;
wire _20261_;
wire _20262_;
wire _20263_;
wire _20264_;
wire _20265_;
wire _20266_;
wire _20267_;
wire _20268_;
wire _20269_;
wire _20270_;
wire _20271_;
wire _20272_;
wire _20273_;
wire _20274_;
wire _20275_;
wire _20276_;
wire _20277_;
wire _20278_;
wire _20279_;
wire _20280_;
wire _20281_;
wire _20282_;
wire _20283_;
wire _20284_;
wire _20285_;
wire _20286_;
wire _20287_;
wire _20288_;
wire _20289_;
wire _20290_;
wire _20291_;
wire _20292_;
wire _20293_;
wire _20294_;
wire _20295_;
wire _20296_;
wire _20297_;
wire _20298_;
wire _20299_;
wire _20300_;
wire _20301_;
wire _20302_;
wire _20303_;
wire _20304_;
wire _20305_;
wire _20306_;
wire _20307_;
wire _20308_;
wire _20309_;
wire _20310_;
wire _20311_;
wire _20312_;
wire _20313_;
wire _20314_;
wire _20315_;
wire _20316_;
wire _20317_;
wire _20318_;
wire _20319_;
wire _20320_;
wire _20321_;
wire _20322_;
wire _20323_;
wire _20324_;
wire _20325_;
wire _20326_;
wire _20327_;
wire _20328_;
wire _20329_;
wire _20330_;
wire _20331_;
wire _20332_;
wire _20333_;
wire _20334_;
wire _20335_;
wire _20336_;
wire _20337_;
wire _20338_;
wire _20339_;
wire _20340_;
wire _20341_;
wire _20342_;
wire _20343_;
wire _20344_;
wire _20345_;
wire _20346_;
wire _20347_;
wire _20348_;
wire _20349_;
wire _20350_;
wire _20351_;
wire _20352_;
wire _20353_;
wire _20354_;
wire _20355_;
wire _20356_;
wire _20357_;
wire _20358_;
wire _20359_;
wire _20360_;
wire _20361_;
wire _20362_;
wire _20363_;
wire _20364_;
wire _20365_;
wire _20366_;
wire _20367_;
wire _20368_;
wire _20369_;
wire _20370_;
wire _20371_;
wire _20372_;
wire _20373_;
wire _20374_;
wire _20375_;
wire _20376_;
wire _20377_;
wire _20378_;
wire _20379_;
wire _20380_;
wire _20381_;
wire _20382_;
wire _20383_;
wire _20384_;
wire _20385_;
wire _20386_;
wire _20387_;
wire _20388_;
wire _20389_;
wire _20390_;
wire _20391_;
wire _20392_;
wire _20393_;
wire _20394_;
wire _20395_;
wire _20396_;
wire _20397_;
wire _20398_;
wire _20399_;
wire _20400_;
wire _20401_;
wire _20402_;
wire _20403_;
wire _20404_;
wire _20405_;
wire _20406_;
wire _20407_;
wire _20408_;
wire _20409_;
wire _20410_;
wire _20411_;
wire _20412_;
wire _20413_;
wire _20414_;
wire _20415_;
wire _20416_;
wire _20417_;
wire _20418_;
wire _20419_;
wire _20420_;
wire _20421_;
wire _20422_;
wire _20423_;
wire _20424_;
wire _20425_;
wire _20426_;
wire _20427_;
wire _20428_;
wire _20429_;
wire _20430_;
wire _20431_;
wire _20432_;
wire _20433_;
wire _20434_;
wire _20435_;
wire _20436_;
wire _20437_;
wire _20438_;
wire _20439_;
wire _20440_;
wire _20441_;
wire _20442_;
wire _20443_;
wire _20444_;
wire _20445_;
wire _20446_;
wire _20447_;
wire _20448_;
wire _20449_;
wire _20450_;
wire _20451_;
wire _20452_;
wire _20453_;
wire _20454_;
wire _20455_;
wire _20456_;
wire _20457_;
wire _20458_;
wire _20459_;
wire _20460_;
wire _20461_;
wire _20462_;
wire _20463_;
wire _20464_;
wire _20465_;
wire _20466_;
wire _20467_;
wire _20468_;
wire _20469_;
wire _20470_;
wire _20471_;
wire _20472_;
wire _20473_;
wire _20474_;
wire _20475_;
wire _20476_;
wire _20477_;
wire _20478_;
wire _20479_;
wire _20480_;
wire _20481_;
wire _20482_;
wire _20483_;
wire _20484_;
wire _20485_;
wire _20486_;
wire _20487_;
wire _20488_;
wire _20489_;
wire _20490_;
wire _20491_;
wire _20492_;
wire _20493_;
wire _20494_;
wire _20495_;
wire _20496_;
wire _20497_;
wire _20498_;
wire _20499_;
wire _20500_;
wire _20501_;
wire _20502_;
wire _20503_;
wire _20504_;
wire _20505_;
wire _20506_;
wire _20507_;
wire _20508_;
wire _20509_;
wire _20510_;
wire _20511_;
wire _20512_;
wire _20513_;
wire _20514_;
wire _20515_;
wire _20516_;
wire _20517_;
wire _20518_;
wire _20519_;
wire _20520_;
wire _20521_;
wire _20522_;
wire _20523_;
wire _20524_;
wire _20525_;
wire _20526_;
wire _20527_;
wire _20528_;
wire _20529_;
wire _20530_;
wire _20531_;
wire _20532_;
wire _20533_;
wire _20534_;
wire _20535_;
wire _20536_;
wire _20537_;
wire _20538_;
wire _20539_;
wire _20540_;
wire _20541_;
wire _20542_;
wire _20543_;
wire _20544_;
wire _20545_;
wire _20546_;
wire _20547_;
wire _20548_;
wire _20549_;
wire _20550_;
wire _20551_;
wire _20552_;
wire _20553_;
wire _20554_;
wire _20555_;
wire _20556_;
wire _20557_;
wire _20558_;
wire _20559_;
wire _20560_;
wire _20561_;
wire _20562_;
wire _20563_;
wire _20564_;
wire _20565_;
wire _20566_;
wire _20567_;
wire _20568_;
wire _20569_;
wire _20570_;
wire _20571_;
wire _20572_;
wire _20573_;
wire _20574_;
wire _20575_;
wire _20576_;
wire _20577_;
wire _20578_;
wire _20579_;
wire _20580_;
wire _20581_;
wire _20582_;
wire _20583_;
wire _20584_;
wire _20585_;
wire _20586_;
wire _20587_;
wire _20588_;
wire _20589_;
wire _20590_;
wire _20591_;
wire _20592_;
wire _20593_;
wire _20594_;
wire _20595_;
wire _20596_;
wire _20597_;
wire _20598_;
wire _20599_;
wire _20600_;
wire _20601_;
wire _20602_;
wire _20603_;
wire _20604_;
wire _20605_;
wire _20606_;
wire _20607_;
wire _20608_;
wire _20609_;
wire _20610_;
wire _20611_;
wire _20612_;
wire _20613_;
wire _20614_;
wire _20615_;
wire _20616_;
wire _20617_;
wire _20618_;
wire _20619_;
wire _20620_;
wire _20621_;
wire _20622_;
wire _20623_;
wire _20624_;
wire _20625_;
wire _20626_;
wire _20627_;
wire _20628_;
wire _20629_;
wire _20630_;
wire _20631_;
wire _20632_;
wire _20633_;
wire _20634_;
wire _20635_;
wire _20636_;
wire _20637_;
wire _20638_;
wire _20639_;
wire _20640_;
wire _20641_;
wire _20642_;
wire _20643_;
wire _20644_;
wire _20645_;
wire _20646_;
wire _20647_;
wire _20648_;
wire _20649_;
wire _20650_;
wire _20651_;
wire _20652_;
wire _20653_;
wire _20654_;
wire _20655_;
wire _20656_;
wire _20657_;
wire _20658_;
wire _20659_;
wire _20660_;
wire _20661_;
wire _20662_;
wire _20663_;
wire _20664_;
wire _20665_;
wire _20666_;
wire _20667_;
wire _20668_;
wire _20669_;
wire _20670_;
wire _20671_;
wire _20672_;
wire _20673_;
wire _20674_;
wire _20675_;
wire _20676_;
wire _20677_;
wire _20678_;
wire _20679_;
wire _20680_;
wire _20681_;
wire _20682_;
wire _20683_;
wire _20684_;
wire _20685_;
wire _20686_;
wire _20687_;
wire _20688_;
wire _20689_;
wire _20690_;
wire _20691_;
wire _20692_;
wire _20693_;
wire _20694_;
wire _20695_;
wire _20696_;
wire _20697_;
wire _20698_;
wire _20699_;
wire _20700_;
wire _20701_;
wire _20702_;
wire _20703_;
wire _20704_;
wire _20705_;
wire _20706_;
wire _20707_;
wire _20708_;
wire _20709_;
wire _20710_;
wire _20711_;
wire _20712_;
wire _20713_;
wire _20714_;
wire _20715_;
wire _20716_;
wire _20717_;
wire _20718_;
wire _20719_;
wire _20720_;
wire _20721_;
wire _20722_;
wire _20723_;
wire _20724_;
wire _20725_;
wire _20726_;
wire _20727_;
wire _20728_;
wire _20729_;
wire _20730_;
wire _20731_;
wire _20732_;
wire _20733_;
wire _20734_;
wire _20735_;
wire _20736_;
wire _20737_;
wire _20738_;
wire _20739_;
wire _20740_;
wire _20741_;
wire _20742_;
wire _20743_;
wire _20744_;
wire _20745_;
wire _20746_;
wire _20747_;
wire _20748_;
wire _20749_;
wire _20750_;
wire _20751_;
wire _20752_;
wire _20753_;
wire _20754_;
wire _20755_;
wire _20756_;
wire _20757_;
wire _20758_;
wire _20759_;
wire _20760_;
wire _20761_;
wire _20762_;
wire _20763_;
wire _20764_;
wire _20765_;
wire _20766_;
wire _20767_;
wire _20768_;
wire _20769_;
wire _20770_;
wire _20771_;
wire _20772_;
wire _20773_;
wire _20774_;
wire _20775_;
wire _20776_;
wire _20777_;
wire _20778_;
wire _20779_;
wire _20780_;
wire _20781_;
wire _20782_;
wire _20783_;
wire _20784_;
wire _20785_;
wire _20786_;
wire _20787_;
wire _20788_;
wire _20789_;
wire _20790_;
wire _20791_;
wire _20792_;
wire _20793_;
wire _20794_;
wire _20795_;
wire _20796_;
wire _20797_;
wire _20798_;
wire _20799_;
wire _20800_;
wire _20801_;
wire _20802_;
wire _20803_;
wire _20804_;
wire _20805_;
wire _20806_;
wire _20807_;
wire _20808_;
wire _20809_;
wire _20810_;
wire _20811_;
wire _20812_;
wire _20813_;
wire _20814_;
wire _20815_;
wire _20816_;
wire _20817_;
wire _20818_;
wire _20819_;
wire _20820_;
wire _20821_;
wire _20822_;
wire _20823_;
wire _20824_;
wire _20825_;
wire _20826_;
wire _20827_;
wire _20828_;
wire _20829_;
wire _20830_;
wire _20831_;
wire _20832_;
wire _20833_;
wire _20834_;
wire _20835_;
wire _20836_;
wire _20837_;
wire _20838_;
wire _20839_;
wire _20840_;
wire _20841_;
wire _20842_;
wire _20843_;
wire _20844_;
wire _20845_;
wire _20846_;
wire _20847_;
wire _20848_;
wire _20849_;
wire _20850_;
wire _20851_;
wire _20852_;
wire _20853_;
wire _20854_;
wire _20855_;
wire _20856_;
wire _20857_;
wire _20858_;
wire _20859_;
wire _20860_;
wire _20861_;
wire _20862_;
wire _20863_;
wire _20864_;
wire _20865_;
wire _20866_;
wire _20867_;
wire _20868_;
wire _20869_;
wire _20870_;
wire _20871_;
wire _20872_;
wire _20873_;
wire _20874_;
wire _20875_;
wire _20876_;
wire _20877_;
wire _20878_;
wire _20879_;
wire _20880_;
wire _20881_;
wire _20882_;
wire _20883_;
wire _20884_;
wire _20885_;
wire _20886_;
wire _20887_;
wire _20888_;
wire _20889_;
wire _20890_;
wire _20891_;
wire _20892_;
wire _20893_;
wire _20894_;
wire _20895_;
wire _20896_;
wire _20897_;
wire _20898_;
wire _20899_;
wire _20900_;
wire _20901_;
wire _20902_;
wire _20903_;
wire _20904_;
wire _20905_;
wire _20906_;
wire _20907_;
wire _20908_;
wire _20909_;
wire _20910_;
wire _20911_;
wire _20912_;
wire _20913_;
wire _20914_;
wire _20915_;
wire _20916_;
wire _20917_;
wire _20918_;
wire _20919_;
wire _20920_;
wire _20921_;
wire _20922_;
wire _20923_;
wire _20924_;
wire _20925_;
wire _20926_;
wire _20927_;
wire _20928_;
wire _20929_;
wire _20930_;
wire _20931_;
wire _20932_;
wire _20933_;
wire _20934_;
wire _20935_;
wire _20936_;
wire _20937_;
wire _20938_;
wire _20939_;
wire _20940_;
wire _20941_;
wire _20942_;
wire _20943_;
wire _20944_;
wire _20945_;
wire _20946_;
wire _20947_;
wire _20948_;
wire _20949_;
wire _20950_;
wire _20951_;
wire _20952_;
wire _20953_;
wire _20954_;
wire _20955_;
wire _20956_;
wire _20957_;
wire _20958_;
wire _20959_;
wire _20960_;
wire _20961_;
wire _20962_;
wire _20963_;
wire _20964_;
wire _20965_;
wire _20966_;
wire _20967_;
wire _20968_;
wire _20969_;
wire _20970_;
wire _20971_;
wire _20972_;
wire _20973_;
wire _20974_;
wire _20975_;
wire _20976_;
wire _20977_;
wire _20978_;
wire _20979_;
wire _20980_;
wire _20981_;
wire _20982_;
wire _20983_;
wire _20984_;
wire _20985_;
wire _20986_;
wire _20987_;
wire _20988_;
wire _20989_;
wire _20990_;
wire _20991_;
wire _20992_;
wire _20993_;
wire _20994_;
wire _20995_;
wire _20996_;
wire _20997_;
wire _20998_;
wire _20999_;
wire _21000_;
wire _21001_;
wire _21002_;
wire _21003_;
wire _21004_;
wire _21005_;
wire _21006_;
wire _21007_;
wire _21008_;
wire _21009_;
wire _21010_;
wire _21011_;
wire _21012_;
wire _21013_;
wire _21014_;
wire _21015_;
wire _21016_;
wire _21017_;
wire _21018_;
wire _21019_;
wire _21020_;
wire _21021_;
wire _21022_;
wire _21023_;
wire _21024_;
wire _21025_;
wire _21026_;
wire _21027_;
wire _21028_;
wire _21029_;
wire _21030_;
wire _21031_;
wire _21032_;
wire _21033_;
wire _21034_;
wire _21035_;
wire _21036_;
wire _21037_;
wire _21038_;
wire _21039_;
wire _21040_;
wire _21041_;
wire _21042_;
wire _21043_;
wire _21044_;
wire _21045_;
wire _21046_;
wire _21047_;
wire _21048_;
wire _21049_;
wire _21050_;
wire _21051_;
wire _21052_;
wire _21053_;
wire _21054_;
wire _21055_;
wire _21056_;
wire _21057_;
wire _21058_;
wire _21059_;
wire _21060_;
wire _21061_;
wire _21062_;
wire _21063_;
wire _21064_;
wire _21065_;
wire _21066_;
wire _21067_;
wire _21068_;
wire _21069_;
wire _21070_;
wire _21071_;
wire _21072_;
wire _21073_;
wire _21074_;
wire _21075_;
wire _21076_;
wire _21077_;
wire _21078_;
wire _21079_;
wire _21080_;
wire _21081_;
wire _21082_;
wire _21083_;
wire _21084_;
wire _21085_;
wire _21086_;
wire _21087_;
wire _21088_;
wire _21089_;
wire _21090_;
wire _21091_;
wire _21092_;
wire _21093_;
wire _21094_;
wire _21095_;
wire _21096_;
wire _21097_;
wire _21098_;
wire _21099_;
wire _21100_;
wire _21101_;
wire _21102_;
wire _21103_;
wire _21104_;
wire _21105_;
wire _21106_;
wire _21107_;
wire _21108_;
wire _21109_;
wire _21110_;
wire _21111_;
wire _21112_;
wire _21113_;
wire _21114_;
wire _21115_;
wire _21116_;
wire _21117_;
wire _21118_;
wire _21119_;
wire _21120_;
wire _21121_;
wire _21122_;
wire _21123_;
wire _21124_;
wire _21125_;
wire _21126_;
wire _21127_;
wire _21128_;
wire _21129_;
wire _21130_;
wire _21131_;
wire _21132_;
wire _21133_;
wire _21134_;
wire _21135_;
wire _21136_;
wire _21137_;
wire _21138_;
wire _21139_;
wire _21140_;
wire _21141_;
wire _21142_;
wire _21143_;
wire _21144_;
wire _21145_;
wire _21146_;
wire _21147_;
wire _21148_;
wire _21149_;
wire _21150_;
wire _21151_;
wire _21152_;
wire _21153_;
wire _21154_;
wire _21155_;
wire _21156_;
wire _21157_;
wire _21158_;
wire _21159_;
wire _21160_;
wire _21161_;
wire _21162_;
wire _21163_;
wire _21164_;
wire _21165_;
wire _21166_;
wire _21167_;
wire _21168_;
wire _21169_;
wire _21170_;
wire _21171_;
wire _21172_;
wire _21173_;
wire _21174_;
wire _21175_;
wire _21176_;
wire _21177_;
wire _21178_;
wire _21179_;
wire _21180_;
wire _21181_;
wire _21182_;
wire _21183_;
wire _21184_;
wire _21185_;
wire _21186_;
wire _21187_;
wire _21188_;
wire _21189_;
wire _21190_;
wire _21191_;
wire _21192_;
wire _21193_;
wire _21194_;
wire _21195_;
wire _21196_;
wire _21197_;
wire _21198_;
wire _21199_;
wire _21200_;
wire _21201_;
wire _21202_;
wire _21203_;
wire _21204_;
wire _21205_;
wire _21206_;
wire _21207_;
wire _21208_;
wire _21209_;
wire _21210_;
wire _21211_;
wire _21212_;
wire _21213_;
wire _21214_;
wire _21215_;
wire _21216_;
wire _21217_;
wire _21218_;
wire _21219_;
wire _21220_;
wire _21221_;
wire _21222_;
wire _21223_;
wire _21224_;
wire _21225_;
wire _21226_;
wire _21227_;
wire _21228_;
wire _21229_;
wire _21230_;
wire _21231_;
wire _21232_;
wire _21233_;
wire _21234_;
wire _21235_;
wire _21236_;
wire _21237_;
wire _21238_;
wire _21239_;
wire _21240_;
wire _21241_;
wire _21242_;
wire _21243_;
wire _21244_;
wire _21245_;
wire _21246_;
wire _21247_;
wire _21248_;
wire _21249_;
wire _21250_;
wire _21251_;
wire _21252_;
wire _21253_;
wire _21254_;
wire _21255_;
wire _21256_;
wire _21257_;
wire _21258_;
wire _21259_;
wire _21260_;
wire _21261_;
wire _21262_;
wire _21263_;
wire _21264_;
wire _21265_;
wire _21266_;
wire _21267_;
wire _21268_;
wire _21269_;
wire _21270_;
wire _21271_;
wire _21272_;
wire _21273_;
wire _21274_;
wire _21275_;
wire _21276_;
wire _21277_;
wire _21278_;
wire _21279_;
wire _21280_;
wire _21281_;
wire _21282_;
wire _21283_;
wire _21284_;
wire _21285_;
wire _21286_;
wire _21287_;
wire _21288_;
wire _21289_;
wire _21290_;
wire _21291_;
wire _21292_;
wire _21293_;
wire _21294_;
wire _21295_;
wire _21296_;
wire _21297_;
wire _21298_;
wire _21299_;
wire _21300_;
wire _21301_;
wire _21302_;
wire _21303_;
wire _21304_;
wire _21305_;
wire _21306_;
wire _21307_;
wire _21308_;
wire _21309_;
wire _21310_;
wire _21311_;
wire _21312_;
wire _21313_;
wire _21314_;
wire _21315_;
wire _21316_;
wire _21317_;
wire _21318_;
wire _21319_;
wire _21320_;
wire _21321_;
wire _21322_;
wire _21323_;
wire _21324_;
wire _21325_;
wire _21326_;
wire _21327_;
wire _21328_;
wire _21329_;
wire _21330_;
wire _21331_;
wire _21332_;
wire _21333_;
wire _21334_;
wire _21335_;
wire _21336_;
wire _21337_;
wire _21338_;
wire _21339_;
wire _21340_;
wire _21341_;
wire _21342_;
wire _21343_;
wire _21344_;
wire _21345_;
wire _21346_;
wire _21347_;
wire _21348_;
wire _21349_;
wire _21350_;
wire _21351_;
wire _21352_;
wire _21353_;
wire _21354_;
wire _21355_;
wire _21356_;
wire _21357_;
wire _21358_;
wire _21359_;
wire _21360_;
wire _21361_;
wire _21362_;
wire _21363_;
wire _21364_;
wire _21365_;
wire _21366_;
wire _21367_;
wire _21368_;
wire _21369_;
wire _21370_;
wire _21371_;
wire _21372_;
wire _21373_;
wire _21374_;
wire _21375_;
wire _21376_;
wire _21377_;
wire _21378_;
wire _21379_;
wire _21380_;
wire _21381_;
wire _21382_;
wire _21383_;
wire _21384_;
wire _21385_;
wire _21386_;
wire _21387_;
wire _21388_;
wire _21389_;
wire _21390_;
wire _21391_;
wire _21392_;
wire _21393_;
wire _21394_;
wire _21395_;
wire _21396_;
wire _21397_;
wire _21398_;
wire _21399_;
wire _21400_;
wire _21401_;
wire _21402_;
wire _21403_;
wire _21404_;
wire _21405_;
wire _21406_;
wire _21407_;
wire _21408_;
wire _21409_;
wire _21410_;
wire _21411_;
wire _21412_;
wire _21413_;
wire _21414_;
wire _21415_;
wire _21416_;
wire _21417_;
wire _21418_;
wire _21419_;
wire _21420_;
wire _21421_;
wire _21422_;
wire _21423_;
wire _21424_;
wire _21425_;
wire _21426_;
wire _21427_;
wire _21428_;
wire _21429_;
wire _21430_;
wire _21431_;
wire _21432_;
wire _21433_;
wire _21434_;
wire _21435_;
wire _21436_;
wire _21437_;
wire _21438_;
wire _21439_;
wire _21440_;
wire _21441_;
wire _21442_;
wire _21443_;
wire _21444_;
wire _21445_;
wire _21446_;
wire _21447_;
wire _21448_;
wire _21449_;
wire _21450_;
wire _21451_;
wire _21452_;
wire _21453_;
wire _21454_;
wire _21455_;
wire _21456_;
wire _21457_;
wire _21458_;
wire _21459_;
wire _21460_;
wire _21461_;
wire _21462_;
wire _21463_;
wire _21464_;
wire _21465_;
wire _21466_;
wire _21467_;
wire _21468_;
wire _21469_;
wire _21470_;
wire _21471_;
wire _21472_;
wire _21473_;
wire _21474_;
wire _21475_;
wire _21476_;
wire _21477_;
wire _21478_;
wire _21479_;
wire _21480_;
wire _21481_;
wire _21482_;
wire _21483_;
wire _21484_;
wire _21485_;
wire _21486_;
wire _21487_;
wire _21488_;
wire _21489_;
wire _21490_;
wire _21491_;
wire _21492_;
wire _21493_;
wire _21494_;
wire _21495_;
wire _21496_;
wire _21497_;
wire _21498_;
wire _21499_;
wire _21500_;
wire _21501_;
wire _21502_;
wire _21503_;
wire _21504_;
wire _21505_;
wire _21506_;
wire _21507_;
wire _21508_;
wire _21509_;
wire _21510_;
wire _21511_;
wire _21512_;
wire _21513_;
wire _21514_;
wire _21515_;
wire _21516_;
wire _21517_;
wire _21518_;
wire _21519_;
wire _21520_;
wire _21521_;
wire _21522_;
wire _21523_;
wire _21524_;
wire _21525_;
wire _21526_;
wire _21527_;
wire _21528_;
wire _21529_;
wire _21530_;
wire _21531_;
wire _21532_;
wire _21533_;
wire _21534_;
wire _21535_;
wire _21536_;
wire _21537_;
wire _21538_;
wire _21539_;
wire _21540_;
wire _21541_;
wire _21542_;
wire _21543_;
wire _21544_;
wire _21545_;
wire _21546_;
wire _21547_;
wire _21548_;
wire _21549_;
wire _21550_;
wire _21551_;
wire _21552_;
wire _21553_;
wire _21554_;
wire _21555_;
wire _21556_;
wire _21557_;
wire _21558_;
wire _21559_;
wire _21560_;
wire _21561_;
wire _21562_;
wire _21563_;
wire _21564_;
wire _21565_;
wire _21566_;
wire _21567_;
wire _21568_;
wire _21569_;
wire _21570_;
wire _21571_;
wire _21572_;
wire _21573_;
wire _21574_;
wire _21575_;
wire _21576_;
wire _21577_;
wire _21578_;
wire _21579_;
wire _21580_;
wire _21581_;
wire _21582_;
wire _21583_;
wire _21584_;
wire _21585_;
wire _21586_;
wire _21587_;
wire _21588_;
wire _21589_;
wire _21590_;
wire _21591_;
wire _21592_;
wire _21593_;
wire _21594_;
wire _21595_;
wire _21596_;
wire _21597_;
wire _21598_;
wire _21599_;
wire _21600_;
wire _21601_;
wire _21602_;
wire _21603_;
wire _21604_;
wire _21605_;
wire _21606_;
wire _21607_;
wire _21608_;
wire _21609_;
wire _21610_;
wire _21611_;
wire _21612_;
wire _21613_;
wire _21614_;
wire _21615_;
wire _21616_;
wire _21617_;
wire _21618_;
wire _21619_;
wire _21620_;
wire _21621_;
wire _21622_;
wire _21623_;
wire _21624_;
wire _21625_;
wire _21626_;
wire _21627_;
wire _21628_;
wire _21629_;
wire _21630_;
wire _21631_;
wire _21632_;
wire _21633_;
wire _21634_;
wire _21635_;
wire _21636_;
wire _21637_;
wire _21638_;
wire _21639_;
wire _21640_;
wire _21641_;
wire _21642_;
wire _21643_;
wire _21644_;
wire _21645_;
wire _21646_;
wire _21647_;
wire _21648_;
wire _21649_;
wire _21650_;
wire _21651_;
wire _21652_;
wire _21653_;
wire _21654_;
wire _21655_;
wire _21656_;
wire _21657_;
wire _21658_;
wire _21659_;
wire _21660_;
wire _21661_;
wire _21662_;
wire _21663_;
wire _21664_;
wire _21665_;
wire _21666_;
wire _21667_;
wire _21668_;
wire _21669_;
wire _21670_;
wire _21671_;
wire _21672_;
wire _21673_;
wire _21674_;
wire _21675_;
wire _21676_;
wire _21677_;
wire _21678_;
wire _21679_;
wire _21680_;
wire _21681_;
wire _21682_;
wire _21683_;
wire _21684_;
wire _21685_;
wire _21686_;
wire _21687_;
wire _21688_;
wire _21689_;
wire _21690_;
wire _21691_;
wire _21692_;
wire _21693_;
wire _21694_;
wire _21695_;
wire _21696_;
wire _21697_;
wire _21698_;
wire _21699_;
wire _21700_;
wire _21701_;
wire _21702_;
wire _21703_;
wire _21704_;
wire _21705_;
wire _21706_;
wire _21707_;
wire _21708_;
wire _21709_;
wire _21710_;
wire _21711_;
wire _21712_;
wire _21713_;
wire _21714_;
wire _21715_;
wire _21716_;
wire _21717_;
wire _21718_;
wire _21719_;
wire _21720_;
wire _21721_;
wire _21722_;
wire _21723_;
wire _21724_;
wire _21725_;
wire _21726_;
wire _21727_;
wire _21728_;
wire _21729_;
wire _21730_;
wire _21731_;
wire _21732_;
wire _21733_;
wire _21734_;
wire _21735_;
wire _21736_;
wire _21737_;
wire _21738_;
wire _21739_;
wire _21740_;
wire _21741_;
wire _21742_;
wire _21743_;
wire _21744_;
wire _21745_;
wire _21746_;
wire _21747_;
wire _21748_;
wire _21749_;
wire _21750_;
wire _21751_;
wire _21752_;
wire _21753_;
wire _21754_;
wire _21755_;
wire _21756_;
wire _21757_;
wire _21758_;
wire _21759_;
wire _21760_;
wire _21761_;
wire _21762_;
wire _21763_;
wire _21764_;
wire _21765_;
wire _21766_;
wire _21767_;
wire _21768_;
wire _21769_;
wire _21770_;
wire _21771_;
wire _21772_;
wire _21773_;
wire _21774_;
wire _21775_;
wire _21776_;
wire _21777_;
wire _21778_;
wire _21779_;
wire _21780_;
wire _21781_;
wire _21782_;
wire _21783_;
wire _21784_;
wire _21785_;
wire _21786_;
wire _21787_;
wire _21788_;
wire _21789_;
wire _21790_;
wire _21791_;
wire _21792_;
wire _21793_;
wire _21794_;
wire _21795_;
wire _21796_;
wire _21797_;
wire _21798_;
wire _21799_;
wire _21800_;
wire _21801_;
wire _21802_;
wire _21803_;
wire _21804_;
wire _21805_;
wire _21806_;
wire _21807_;
wire _21808_;
wire _21809_;
wire _21810_;
wire _21811_;
wire _21812_;
wire _21813_;
wire _21814_;
wire _21815_;
wire _21816_;
wire _21817_;
wire _21818_;
wire _21819_;
wire _21820_;
wire _21821_;
wire _21822_;
wire _21823_;
wire _21824_;
wire _21825_;
wire _21826_;
wire _21827_;
wire _21828_;
wire _21829_;
wire _21830_;
wire _21831_;
wire _21832_;
wire _21833_;
wire _21834_;
wire _21835_;
wire _21836_;
wire _21837_;
wire _21838_;
wire _21839_;
wire _21840_;
wire _21841_;
wire _21842_;
wire _21843_;
wire _21844_;
wire _21845_;
wire _21846_;
wire _21847_;
wire _21848_;
wire _21849_;
wire _21850_;
wire _21851_;
wire _21852_;
wire _21853_;
wire _21854_;
wire _21855_;
wire _21856_;
wire _21857_;
wire _21858_;
wire _21859_;
wire _21860_;
wire _21861_;
wire _21862_;
wire _21863_;
wire _21864_;
wire _21865_;
wire _21866_;
wire _21867_;
wire _21868_;
wire _21869_;
wire _21870_;
wire _21871_;
wire _21872_;
wire _21873_;
wire _21874_;
wire _21875_;
wire _21876_;
wire _21877_;
wire _21878_;
wire _21879_;
wire _21880_;
wire _21881_;
wire _21882_;
wire _21883_;
wire _21884_;
wire _21885_;
wire _21886_;
wire _21887_;
wire _21888_;
wire _21889_;
wire _21890_;
wire _21891_;
wire _21892_;
wire _21893_;
wire _21894_;
wire _21895_;
wire _21896_;
wire _21897_;
wire _21898_;
wire _21899_;
wire _21900_;
wire _21901_;
wire _21902_;
wire _21903_;
wire _21904_;
wire _21905_;
wire _21906_;
wire _21907_;
wire _21908_;
wire _21909_;
wire _21910_;
wire _21911_;
wire _21912_;
wire _21913_;
wire _21914_;
wire _21915_;
wire _21916_;
wire _21917_;
wire _21918_;
wire _21919_;
wire _21920_;
wire _21921_;
wire _21922_;
wire _21923_;
wire _21924_;
wire _21925_;
wire _21926_;
wire _21927_;
wire _21928_;
wire _21929_;
wire _21930_;
wire _21931_;
wire _21932_;
wire _21933_;
wire _21934_;
wire _21935_;
wire _21936_;
wire _21937_;
wire _21938_;
wire _21939_;
wire _21940_;
wire _21941_;
wire _21942_;
wire _21943_;
wire _21944_;
wire _21945_;
wire _21946_;
wire _21947_;
wire _21948_;
wire _21949_;
wire _21950_;
wire _21951_;
wire _21952_;
wire _21953_;
wire _21954_;
wire _21955_;
wire _21956_;
wire _21957_;
wire _21958_;
wire _21959_;
wire _21960_;
wire _21961_;
wire _21962_;
wire _21963_;
wire _21964_;
wire _21965_;
wire _21966_;
wire _21967_;
wire _21968_;
wire _21969_;
wire _21970_;
wire _21971_;
wire _21972_;
wire _21973_;
wire _21974_;
wire _21975_;
wire _21976_;
wire _21977_;
wire _21978_;
wire _21979_;
wire _21980_;
wire _21981_;
wire _21982_;
wire _21983_;
wire _21984_;
wire _21985_;
wire _21986_;
wire _21987_;
wire _21988_;
wire _21989_;
wire _21990_;
wire _21991_;
wire _21992_;
wire _21993_;
wire _21994_;
wire _21995_;
wire _21996_;
wire _21997_;
wire _21998_;
wire _21999_;
wire _22000_;
wire _22001_;
wire _22002_;
wire _22003_;
wire _22004_;
wire _22005_;
wire _22006_;
wire _22007_;
wire _22008_;
wire _22009_;
wire _22010_;
wire _22011_;
wire _22012_;
wire _22013_;
wire _22014_;
wire _22015_;
wire _22016_;
wire _22017_;
wire _22018_;
wire _22019_;
wire _22020_;
wire _22021_;
wire _22022_;
wire _22023_;
wire _22024_;
wire _22025_;
wire _22026_;
wire _22027_;
wire _22028_;
wire _22029_;
wire _22030_;
wire _22031_;
wire _22032_;
wire _22033_;
wire _22034_;
wire _22035_;
wire _22036_;
wire _22037_;
wire _22038_;
wire _22039_;
wire _22040_;
wire _22041_;
wire _22042_;
wire _22043_;
wire _22044_;
wire _22045_;
wire _22046_;
wire _22047_;
wire _22048_;
wire _22049_;
wire _22050_;
wire _22051_;
wire _22052_;
wire _22053_;
wire _22054_;
wire _22055_;
wire _22056_;
wire _22057_;
wire _22058_;
wire _22059_;
wire _22060_;
wire _22061_;
wire _22062_;
wire _22063_;
wire _22064_;
wire _22065_;
wire _22066_;
wire _22067_;
wire _22068_;
wire _22069_;
wire _22070_;
wire _22071_;
wire _22072_;
wire _22073_;
wire _22074_;
wire _22075_;
wire _22076_;
wire _22077_;
wire _22078_;
wire _22079_;
wire _22080_;
wire _22081_;
wire _22082_;
wire _22083_;
wire _22084_;
wire _22085_;
wire _22086_;
wire _22087_;
wire _22088_;
wire _22089_;
wire _22090_;
wire _22091_;
wire _22092_;
wire _22093_;
wire _22094_;
wire _22095_;
wire _22096_;
wire _22097_;
wire _22098_;
wire _22099_;
wire _22100_;
wire _22101_;
wire _22102_;
wire _22103_;
wire _22104_;
wire _22105_;
wire _22106_;
wire _22107_;
wire _22108_;
wire _22109_;
wire _22110_;
wire _22111_;
wire _22112_;
wire _22113_;
wire _22114_;
wire _22115_;
wire _22116_;
wire _22117_;
wire _22118_;
wire _22119_;
wire _22120_;
wire _22121_;
wire _22122_;
wire _22123_;
wire _22124_;
wire _22125_;
wire _22126_;
wire _22127_;
wire _22128_;
wire _22129_;
wire _22130_;
wire _22131_;
wire _22132_;
wire _22133_;
wire _22134_;
wire _22135_;
wire _22136_;
wire _22137_;
wire _22138_;
wire _22139_;
wire _22140_;
wire _22141_;
wire _22142_;
wire _22143_;
wire _22144_;
wire _22145_;
wire _22146_;
wire _22147_;
wire _22148_;
wire _22149_;
wire _22150_;
wire _22151_;
wire _22152_;
wire _22153_;
wire _22154_;
wire _22155_;
wire _22156_;
wire _22157_;
wire _22158_;
wire _22159_;
wire _22160_;
wire _22161_;
wire _22162_;
wire _22163_;
wire _22164_;
wire _22165_;
wire _22166_;
wire _22167_;
wire _22168_;
wire _22169_;
wire _22170_;
wire _22171_;
wire _22172_;
wire _22173_;
wire _22174_;
wire _22175_;
wire _22176_;
wire _22177_;
wire _22178_;
wire _22179_;
wire _22180_;
wire _22181_;
wire _22182_;
wire _22183_;
wire _22184_;
wire _22185_;
wire _22186_;
wire _22187_;
wire _22188_;
wire _22189_;
wire _22190_;
wire _22191_;
wire _22192_;
wire _22193_;
wire _22194_;
wire _22195_;
wire _22196_;
wire _22197_;
wire _22198_;
wire _22199_;
wire _22200_;
wire _22201_;
wire _22202_;
wire _22203_;
wire _22204_;
wire _22205_;
wire _22206_;
wire _22207_;
wire _22208_;
wire _22209_;
wire _22210_;
wire _22211_;
wire _22212_;
wire _22213_;
wire _22214_;
wire _22215_;
wire _22216_;
wire _22217_;
wire _22218_;
wire _22219_;
wire _22220_;
wire _22221_;
wire _22222_;
wire _22223_;
wire _22224_;
wire _22225_;
wire _22226_;
wire _22227_;
wire _22228_;
wire _22229_;
wire _22230_;
wire _22231_;
wire _22232_;
wire _22233_;
wire _22234_;
wire _22235_;
wire _22236_;
wire _22237_;
wire _22238_;
wire _22239_;
wire _22240_;
wire _22241_;
wire _22242_;
wire _22243_;
wire _22244_;
wire _22245_;
wire _22246_;
wire _22247_;
wire _22248_;
wire _22249_;
wire _22250_;
wire _22251_;
wire _22252_;
wire _22253_;
wire _22254_;
wire _22255_;
wire _22256_;
wire _22257_;
wire _22258_;
wire _22259_;
wire _22260_;
wire _22261_;
wire _22262_;
wire _22263_;
wire _22264_;
wire _22265_;
wire _22266_;
wire _22267_;
wire _22268_;
wire _22269_;
wire _22270_;
wire _22271_;
wire _22272_;
wire _22273_;
wire _22274_;
wire _22275_;
wire _22276_;
wire _22277_;
wire _22278_;
wire _22279_;
wire _22280_;
wire _22281_;
wire _22282_;
wire _22283_;
wire _22284_;
wire _22285_;
wire _22286_;
wire _22287_;
wire _22288_;
wire _22289_;
wire _22290_;
wire _22291_;
wire _22292_;
wire _22293_;
wire _22294_;
wire _22295_;
wire _22296_;
wire _22297_;
wire _22298_;
wire _22299_;
wire _22300_;
wire _22301_;
wire _22302_;
wire _22303_;
wire _22304_;
wire _22305_;
wire _22306_;
wire _22307_;
wire _22308_;
wire _22309_;
wire _22310_;
wire _22311_;
wire _22312_;
wire _22313_;
wire _22314_;
wire _22315_;
wire _22316_;
wire _22317_;
wire _22318_;
wire _22319_;
wire _22320_;
wire _22321_;
wire _22322_;
wire _22323_;
wire _22324_;
wire _22325_;
wire _22326_;
wire _22327_;
wire _22328_;
wire _22329_;
wire _22330_;
wire _22331_;
wire _22332_;
wire _22333_;
wire _22334_;
wire _22335_;
wire _22336_;
wire _22337_;
wire _22338_;
wire _22339_;
wire _22340_;
wire _22341_;
wire _22342_;
wire _22343_;
wire _22344_;
wire _22345_;
wire _22346_;
wire _22347_;
wire _22348_;
wire _22349_;
wire _22350_;
wire _22351_;
wire _22352_;
wire _22353_;
wire _22354_;
wire _22355_;
wire _22356_;
wire _22357_;
wire _22358_;
wire _22359_;
wire _22360_;
wire _22361_;
wire _22362_;
wire _22363_;
wire _22364_;
wire _22365_;
wire _22366_;
wire _22367_;
wire _22368_;
wire _22369_;
wire _22370_;
wire _22371_;
wire _22372_;
wire _22373_;
wire _22374_;
wire _22375_;
wire _22376_;
wire _22377_;
wire _22378_;
wire _22379_;
wire _22380_;
wire _22381_;
wire _22382_;
wire _22383_;
wire _22384_;
wire _22385_;
wire _22386_;
wire _22387_;
wire _22388_;
wire _22389_;
wire _22390_;
wire _22391_;
wire _22392_;
wire _22393_;
wire _22394_;
wire _22395_;
wire _22396_;
wire _22397_;
wire _22398_;
wire _22399_;
wire _22400_;
wire _22401_;
wire _22402_;
wire _22403_;
wire _22404_;
wire _22405_;
wire _22406_;
wire _22407_;
wire _22408_;
wire _22409_;
wire _22410_;
wire _22411_;
wire _22412_;
wire _22413_;
wire _22414_;
wire _22415_;
wire _22416_;
wire _22417_;
wire _22418_;
wire _22419_;
wire _22420_;
wire _22421_;
wire _22422_;
wire _22423_;
wire _22424_;
wire _22425_;
wire _22426_;
wire _22427_;
wire _22428_;
wire _22429_;
wire _22430_;
wire _22431_;
wire _22432_;
wire _22433_;
wire _22434_;
wire _22435_;
wire _22436_;
wire _22437_;
wire _22438_;
wire _22439_;
wire _22440_;
wire _22441_;
wire _22442_;
wire _22443_;
wire _22444_;
wire _22445_;
wire _22446_;
wire _22447_;
wire _22448_;
wire _22449_;
wire _22450_;
wire _22451_;
wire _22452_;
wire _22453_;
wire _22454_;
wire _22455_;
wire _22456_;
wire _22457_;
wire _22458_;
wire _22459_;
wire _22460_;
wire _22461_;
wire _22462_;
wire _22463_;
wire _22464_;
wire _22465_;
wire _22466_;
wire _22467_;
wire _22468_;
wire _22469_;
wire _22470_;
wire _22471_;
wire _22472_;
wire _22473_;
wire _22474_;
wire _22475_;
wire _22476_;
wire _22477_;
wire _22478_;
wire _22479_;
wire _22480_;
wire _22481_;
wire _22482_;
wire _22483_;
wire _22484_;
wire _22485_;
wire _22486_;
wire _22487_;
wire _22488_;
wire _22489_;
wire _22490_;
wire _22491_;
wire _22492_;
wire _22493_;
wire _22494_;
wire _22495_;
wire _22496_;
wire _22497_;
wire _22498_;
wire _22499_;
wire _22500_;
wire _22501_;
wire _22502_;
wire _22503_;
wire _22504_;
wire _22505_;
wire _22506_;
wire _22507_;
wire _22508_;
wire _22509_;
wire _22510_;
wire _22511_;
wire _22512_;
wire _22513_;
wire _22514_;
wire _22515_;
wire _22516_;
wire _22517_;
wire _22518_;
wire _22519_;
wire _22520_;
wire _22521_;
wire _22522_;
wire _22523_;
wire _22524_;
wire _22525_;
wire _22526_;
wire _22527_;
wire _22528_;
wire _22529_;
wire _22530_;
wire _22531_;
wire _22532_;
wire _22533_;
wire _22534_;
wire _22535_;
wire _22536_;
wire _22537_;
wire _22538_;
wire _22539_;
wire _22540_;
wire _22541_;
wire _22542_;
wire _22543_;
wire _22544_;
wire _22545_;
wire _22546_;
wire _22547_;
wire _22548_;
wire _22549_;
wire _22550_;
wire _22551_;
wire _22552_;
wire _22553_;
wire _22554_;
wire _22555_;
wire _22556_;
wire _22557_;
wire _22558_;
wire _22559_;
wire _22560_;
wire _22561_;
wire _22562_;
wire _22563_;
wire _22564_;
wire _22565_;
wire _22566_;
wire _22567_;
wire _22568_;
wire _22569_;
wire _22570_;
wire _22571_;
wire _22572_;
wire _22573_;
wire _22574_;
wire _22575_;
wire _22576_;
wire _22577_;
wire _22578_;
wire _22579_;
wire _22580_;
wire _22581_;
wire _22582_;
wire _22583_;
wire _22584_;
wire _22585_;
wire _22586_;
wire _22587_;
wire _22588_;
wire _22589_;
wire _22590_;
wire _22591_;
wire _22592_;
wire _22593_;
wire _22594_;
wire _22595_;
wire _22596_;
wire _22597_;
wire _22598_;
wire _22599_;
wire _22600_;
wire _22601_;
wire _22602_;
wire _22603_;
wire _22604_;
wire _22605_;
wire _22606_;
wire _22607_;
wire _22608_;
wire _22609_;
wire _22610_;
wire _22611_;
wire _22612_;
wire _22613_;
wire _22614_;
wire _22615_;
wire _22616_;
wire _22617_;
wire _22618_;
wire _22619_;
wire _22620_;
wire _22621_;
wire _22622_;
wire _22623_;
wire _22624_;
wire _22625_;
wire _22626_;
wire _22627_;
wire _22628_;
wire _22629_;
wire _22630_;
wire _22631_;
wire _22632_;
wire _22633_;
wire _22634_;
wire _22635_;
wire _22636_;
wire _22637_;
wire _22638_;
wire _22639_;
wire _22640_;
wire _22641_;
wire _22642_;
wire _22643_;
wire _22644_;
wire _22645_;
wire _22646_;
wire _22647_;
wire _22648_;
wire _22649_;
wire _22650_;
wire _22651_;
wire _22652_;
wire _22653_;
wire _22654_;
wire _22655_;
wire _22656_;
wire _22657_;
wire _22658_;
wire _22659_;
wire _22660_;
wire _22661_;
wire _22662_;
wire _22663_;
wire _22664_;
wire _22665_;
wire _22666_;
wire _22667_;
wire _22668_;
wire _22669_;
wire _22670_;
wire _22671_;
wire _22672_;
wire _22673_;
wire _22674_;
wire _22675_;
wire _22676_;
wire _22677_;
wire _22678_;
wire _22679_;
wire _22680_;
wire _22681_;
wire _22682_;
wire _22683_;
wire _22684_;
wire _22685_;
wire _22686_;
wire _22687_;
wire _22688_;
wire _22689_;
wire _22690_;
wire _22691_;
wire _22692_;
wire _22693_;
wire _22694_;
wire _22695_;
wire _22696_;
wire _22697_;
wire _22698_;
wire _22699_;
wire _22700_;
wire _22701_;
wire _22702_;
wire _22703_;
wire _22704_;
wire _22705_;
wire _22706_;
wire _22707_;
wire _22708_;
wire _22709_;
wire _22710_;
wire _22711_;
wire _22712_;
wire _22713_;
wire _22714_;
wire _22715_;
wire _22716_;
wire _22717_;
wire _22718_;
wire _22719_;
wire _22720_;
wire _22721_;
wire _22722_;
wire _22723_;
wire _22724_;
wire _22725_;
wire _22726_;
wire _22727_;
wire _22728_;
wire _22729_;
wire _22730_;
wire _22731_;
wire _22732_;
wire _22733_;
wire _22734_;
wire _22735_;
wire _22736_;
wire _22737_;
wire _22738_;
wire _22739_;
wire _22740_;
wire _22741_;
wire _22742_;
wire _22743_;
wire _22744_;
wire _22745_;
wire _22746_;
wire _22747_;
wire _22748_;
wire _22749_;
wire _22750_;
wire _22751_;
wire _22752_;
wire _22753_;
wire _22754_;
wire _22755_;
wire _22756_;
wire _22757_;
wire _22758_;
wire _22759_;
wire _22760_;
wire _22761_;
wire _22762_;
wire _22763_;
wire _22764_;
wire _22765_;
wire _22766_;
wire _22767_;
wire _22768_;
wire _22769_;
wire _22770_;
wire _22771_;
wire _22772_;
wire _22773_;
wire _22774_;
wire _22775_;
wire _22776_;
wire _22777_;
wire _22778_;
wire _22779_;
wire _22780_;
wire _22781_;
wire _22782_;
wire _22783_;
wire _22784_;
wire _22785_;
wire _22786_;
wire _22787_;
wire _22788_;
wire _22789_;
wire _22790_;
wire _22791_;
wire _22792_;
wire _22793_;
wire _22794_;
wire _22795_;
wire _22796_;
wire _22797_;
wire _22798_;
wire _22799_;
wire _22800_;
wire _22801_;
wire _22802_;
wire _22803_;
wire _22804_;
wire _22805_;
wire _22806_;
wire _22807_;
wire _22808_;
wire _22809_;
wire _22810_;
wire _22811_;
wire _22812_;
wire _22813_;
wire _22814_;
wire _22815_;
wire _22816_;
wire _22817_;
wire _22818_;
wire _22819_;
wire _22820_;
wire _22821_;
wire _22822_;
wire _22823_;
wire _22824_;
wire _22825_;
wire _22826_;
wire _22827_;
wire _22828_;
wire _22829_;
wire _22830_;
wire _22831_;
wire _22832_;
wire _22833_;
wire _22834_;
wire _22835_;
wire _22836_;
wire _22837_;
wire _22838_;
wire _22839_;
wire _22840_;
wire _22841_;
wire _22842_;
wire _22843_;
wire _22844_;
wire _22845_;
wire _22846_;
wire _22847_;
wire _22848_;
wire _22849_;
wire _22850_;
wire _22851_;
wire _22852_;
wire _22853_;
wire _22854_;
wire _22855_;
wire _22856_;
wire _22857_;
wire _22858_;
wire _22859_;
wire _22860_;
wire _22861_;
wire _22862_;
wire _22863_;
wire _22864_;
wire _22865_;
wire _22866_;
wire _22867_;
wire _22868_;
wire _22869_;
wire _22870_;
wire _22871_;
wire _22872_;
wire _22873_;
wire _22874_;
wire _22875_;
wire _22876_;
wire _22877_;
wire _22878_;
wire _22879_;
wire _22880_;
wire _22881_;
wire _22882_;
wire _22883_;
wire _22884_;
wire _22885_;
wire _22886_;
wire _22887_;
wire _22888_;
wire _22889_;
wire _22890_;
wire _22891_;
wire _22892_;
wire _22893_;
wire _22894_;
wire _22895_;
wire _22896_;
wire _22897_;
wire _22898_;
wire _22899_;
wire _22900_;
wire _22901_;
wire _22902_;
wire _22903_;
wire _22904_;
wire _22905_;
wire _22906_;
wire _22907_;
wire _22908_;
wire _22909_;
wire _22910_;
wire _22911_;
wire _22912_;
wire _22913_;
wire _22914_;
wire _22915_;
wire _22916_;
wire _22917_;
wire _22918_;
wire _22919_;
wire _22920_;
wire _22921_;
wire _22922_;
wire _22923_;
wire _22924_;
wire _22925_;
wire _22926_;
wire _22927_;
wire _22928_;
wire _22929_;
wire _22930_;
wire _22931_;
wire _22932_;
wire _22933_;
wire _22934_;
wire _22935_;
wire _22936_;
wire _22937_;
wire _22938_;
wire _22939_;
wire _22940_;
wire _22941_;
wire _22942_;
wire _22943_;
wire _22944_;
wire _22945_;
wire _22946_;
wire _22947_;
wire _22948_;
wire _22949_;
wire _22950_;
wire _22951_;
wire _22952_;
wire _22953_;
wire _22954_;
wire _22955_;
wire _22956_;
wire _22957_;
wire _22958_;
wire _22959_;
wire _22960_;
wire _22961_;
wire _22962_;
wire _22963_;
wire _22964_;
wire _22965_;
wire _22966_;
wire _22967_;
wire _22968_;
wire _22969_;
wire _22970_;
wire _22971_;
wire _22972_;
wire _22973_;
wire _22974_;
wire _22975_;
wire _22976_;
wire _22977_;
wire _22978_;
wire _22979_;
wire _22980_;
wire _22981_;
wire _22982_;
wire _22983_;
wire _22984_;
wire _22985_;
wire _22986_;
wire _22987_;
wire _22988_;
wire _22989_;
wire _22990_;
wire _22991_;
wire _22992_;
wire _22993_;
wire _22994_;
wire _22995_;
wire _22996_;
wire _22997_;
wire _22998_;
wire _22999_;
wire _23000_;
wire _23001_;
wire _23002_;
wire _23003_;
wire _23004_;
wire _23005_;
wire _23006_;
wire _23007_;
wire _23008_;
wire _23009_;
wire _23010_;
wire _23011_;
wire _23012_;
wire _23013_;
wire _23014_;
wire _23015_;
wire _23016_;
wire _23017_;
wire _23018_;
wire _23019_;
wire _23020_;
wire _23021_;
wire _23022_;
wire _23023_;
wire _23024_;
wire _23025_;
wire _23026_;
wire _23027_;
wire _23028_;
wire _23029_;
wire _23030_;
wire _23031_;
wire _23032_;
wire _23033_;
wire _23034_;
wire _23035_;
wire _23036_;
wire _23037_;
wire _23038_;
wire _23039_;
wire _23040_;
wire _23041_;
wire _23042_;
wire _23043_;
wire _23044_;
wire _23045_;
wire _23046_;
wire _23047_;
wire _23048_;
wire _23049_;
wire _23050_;
wire _23051_;
wire _23052_;
wire _23053_;
wire _23054_;
wire _23055_;
wire _23056_;
wire _23057_;
wire _23058_;
wire _23059_;
wire _23060_;
wire _23061_;
wire _23062_;
wire _23063_;
wire _23064_;
wire _23065_;
wire _23066_;
wire _23067_;
wire _23068_;
wire _23069_;
wire _23070_;
wire _23071_;
wire _23072_;
wire _23073_;
wire _23074_;
wire _23075_;
wire _23076_;
wire _23077_;
wire _23078_;
wire _23079_;
wire _23080_;
wire _23081_;
wire _23082_;
wire _23083_;
wire _23084_;
wire _23085_;
wire _23086_;
wire _23087_;
wire _23088_;
wire _23089_;
wire _23090_;
wire _23091_;
wire _23092_;
wire _23093_;
wire _23094_;
wire _23095_;
wire _23096_;
wire _23097_;
wire _23098_;
wire _23099_;
wire _23100_;
wire _23101_;
wire _23102_;
wire _23103_;
wire _23104_;
wire _23105_;
wire _23106_;
wire _23107_;
wire _23108_;
wire _23109_;
wire _23110_;
wire _23111_;
wire _23112_;
wire _23113_;
wire _23114_;
wire _23115_;
wire _23116_;
wire _23117_;
wire _23118_;
wire _23119_;
wire _23120_;
wire _23121_;
wire _23122_;
wire _23123_;
wire _23124_;
wire _23125_;
wire _23126_;
wire _23127_;
wire _23128_;
wire _23129_;
wire _23130_;
wire _23131_;
wire _23132_;
wire _23133_;
wire _23134_;
wire _23135_;
wire _23136_;
wire _23137_;
wire _23138_;
wire _23139_;
wire _23140_;
wire _23141_;
wire _23142_;
wire _23143_;
wire _23144_;
wire _23145_;
wire _23146_;
wire _23147_;
wire _23148_;
wire _23149_;
wire _23150_;
wire _23151_;
wire _23152_;
wire _23153_;
wire _23154_;
wire _23155_;
wire _23156_;
wire _23157_;
wire _23158_;
wire _23159_;
wire _23160_;
wire _23161_;
wire _23162_;
wire _23163_;
wire _23164_;
wire _23165_;
wire _23166_;
wire _23167_;
wire _23168_;
wire _23169_;
wire _23170_;
wire _23171_;
wire _23172_;
wire _23173_;
wire _23174_;
wire _23175_;
wire _23176_;
wire _23177_;
wire _23178_;
wire _23179_;
wire _23180_;
wire _23181_;
wire _23182_;
wire _23183_;
wire _23184_;
wire _23185_;
wire _23186_;
wire _23187_;
wire _23188_;
wire _23189_;
wire _23190_;
wire _23191_;
wire _23192_;
wire _23193_;
wire _23194_;
wire _23195_;
wire _23196_;
wire _23197_;
wire _23198_;
wire _23199_;
wire _23200_;
wire _23201_;
wire _23202_;
wire _23203_;
wire _23204_;
wire _23205_;
wire _23206_;
wire _23207_;
wire _23208_;
wire _23209_;
wire _23210_;
wire _23211_;
wire _23212_;
wire _23213_;
wire _23214_;
wire _23215_;
wire _23216_;
wire _23217_;
wire _23218_;
wire _23219_;
wire _23220_;
wire _23221_;
wire _23222_;
wire _23223_;
wire _23224_;
wire _23225_;
wire _23226_;
wire _23227_;
wire _23228_;
wire _23229_;
wire _23230_;
wire _23231_;
wire _23232_;
wire _23233_;
wire _23234_;
wire _23235_;
wire _23236_;
wire _23237_;
wire _23238_;
wire _23239_;
wire _23240_;
wire _23241_;
wire _23242_;
wire _23243_;
wire _23244_;
wire _23245_;
wire _23246_;
wire _23247_;
wire _23248_;
wire _23249_;
wire _23250_;
wire _23251_;
wire _23252_;
wire _23253_;
wire _23254_;
wire _23255_;
wire _23256_;
wire _23257_;
wire _23258_;
wire _23259_;
wire _23260_;
wire _23261_;
wire _23262_;
wire _23263_;
wire _23264_;
wire _23265_;
wire _23266_;
wire _23267_;
wire _23268_;
wire _23269_;
wire _23270_;
wire _23271_;
wire _23272_;
wire _23273_;
wire _23274_;
wire _23275_;
wire _23276_;
wire _23277_;
wire _23278_;
wire _23279_;
wire _23280_;
wire _23281_;
wire _23282_;
wire _23283_;
wire _23284_;
wire _23285_;
wire _23286_;
wire _23287_;
wire _23288_;
wire _23289_;
wire _23290_;
wire _23291_;
wire _23292_;
wire _23293_;
wire _23294_;
wire _23295_;
wire _23296_;
wire _23297_;
wire _23298_;
wire _23299_;
wire _23300_;
wire _23301_;
wire _23302_;
wire _23303_;
wire _23304_;
wire _23305_;
wire _23306_;
wire _23307_;
wire _23308_;
wire _23309_;
wire _23310_;
wire _23311_;
wire _23312_;
wire _23313_;
wire _23314_;
wire _23315_;
wire _23316_;
wire _23317_;
wire _23318_;
wire _23319_;
wire _23320_;
wire _23321_;
wire _23322_;
wire _23323_;
wire _23324_;
wire _23325_;
wire _23326_;
wire _23327_;
wire _23328_;
wire _23329_;
wire _23330_;
wire _23331_;
wire _23332_;
wire _23333_;
wire _23334_;
wire _23335_;
wire _23336_;
wire _23337_;
wire _23338_;
wire _23339_;
wire _23340_;
wire _23341_;
wire _23342_;
wire _23343_;
wire _23344_;
wire _23345_;
wire _23346_;
wire _23347_;
wire _23348_;
wire _23349_;
wire _23350_;
wire _23351_;
wire _23352_;
wire _23353_;
wire _23354_;
wire _23355_;
wire _23356_;
wire _23357_;
wire _23358_;
wire _23359_;
wire _23360_;
wire _23361_;
wire _23362_;
wire _23363_;
wire _23364_;
wire _23365_;
wire _23366_;
wire _23367_;
wire _23368_;
wire _23369_;
wire _23370_;
wire _23371_;
wire _23372_;
wire _23373_;
wire _23374_;
wire _23375_;
wire _23376_;
wire _23377_;
wire _23378_;
wire _23379_;
wire _23380_;
wire _23381_;
wire _23382_;
wire _23383_;
wire _23384_;
wire _23385_;
wire _23386_;
wire _23387_;
wire _23388_;
wire _23389_;
wire _23390_;
wire _23391_;
wire _23392_;
wire _23393_;
wire _23394_;
wire _23395_;
wire _23396_;
wire _23397_;
wire _23398_;
wire _23399_;
wire _23400_;
wire _23401_;
wire _23402_;
wire _23403_;
wire _23404_;
wire _23405_;
wire _23406_;
wire _23407_;
wire _23408_;
wire _23409_;
wire _23410_;
wire _23411_;
wire _23412_;
wire _23413_;
wire _23414_;
wire _23415_;
wire _23416_;
wire _23417_;
wire _23418_;
wire _23419_;
wire _23420_;
wire _23421_;
wire _23422_;
wire _23423_;
wire _23424_;
wire _23425_;
wire _23426_;
wire _23427_;
wire _23428_;
wire _23429_;
wire _23430_;
wire _23431_;
wire _23432_;
wire _23433_;
wire _23434_;
wire _23435_;
wire _23436_;
wire _23437_;
wire _23438_;
wire _23439_;
wire _23440_;
wire _23441_;
wire _23442_;
wire _23443_;
wire _23444_;
wire _23445_;
wire _23446_;
wire _23447_;
wire _23448_;
wire _23449_;
wire _23450_;
wire _23451_;
wire _23452_;
wire _23453_;
wire _23454_;
wire _23455_;
wire _23456_;
wire _23457_;
wire _23458_;
wire _23459_;
wire _23460_;
wire _23461_;
wire _23462_;
wire _23463_;
wire _23464_;
wire _23465_;
wire _23466_;
wire _23467_;
wire _23468_;
wire _23469_;
wire _23470_;
wire _23471_;
wire _23472_;
wire _23473_;
wire _23474_;
wire _23475_;
wire _23476_;
wire _23477_;
wire _23478_;
wire _23479_;
wire _23480_;
wire _23481_;
wire _23482_;
wire _23483_;
wire _23484_;
wire _23485_;
wire _23486_;
wire _23487_;
wire _23488_;
wire _23489_;
wire _23490_;
wire _23491_;
wire _23492_;
wire _23493_;
wire _23494_;
wire _23495_;
wire _23496_;
wire _23497_;
wire _23498_;
wire _23499_;
wire _23500_;
wire _23501_;
wire _23502_;
wire _23503_;
wire _23504_;
wire _23505_;
wire _23506_;
wire _23507_;
wire _23508_;
wire _23509_;
wire _23510_;
wire _23511_;
wire _23512_;
wire _23513_;
wire _23514_;
wire _23515_;
wire _23516_;
wire _23517_;
wire _23518_;
wire _23519_;
wire _23520_;
wire _23521_;
wire _23522_;
wire _23523_;
wire _23524_;
wire _23525_;
wire _23526_;
wire _23527_;
wire _23528_;
wire _23529_;
wire _23530_;
wire _23531_;
wire _23532_;
wire _23533_;
wire _23534_;
wire _23535_;
wire _23536_;
wire _23537_;
wire _23538_;
wire _23539_;
wire _23540_;
wire _23541_;
wire _23542_;
wire _23543_;
wire _23544_;
wire _23545_;
wire _23546_;
wire _23547_;
wire _23548_;
wire _23549_;
wire _23550_;
wire _23551_;
wire _23552_;
wire _23553_;
wire _23554_;
wire _23555_;
wire _23556_;
wire _23557_;
wire _23558_;
wire _23559_;
wire _23560_;
wire _23561_;
wire _23562_;
wire _23563_;
wire _23564_;
wire _23565_;
wire _23566_;
wire _23567_;
wire _23568_;
wire _23569_;
wire _23570_;
wire _23571_;
wire _23572_;
wire _23573_;
wire _23574_;
wire _23575_;
wire _23576_;
wire _23577_;
wire _23578_;
wire _23579_;
wire _23580_;
wire _23581_;
wire _23582_;
wire _23583_;
wire _23584_;
wire _23585_;
wire _23586_;
wire _23587_;
wire _23588_;
wire _23589_;
wire _23590_;
wire _23591_;
wire _23592_;
wire _23593_;
wire _23594_;
wire _23595_;
wire _23596_;
wire _23597_;
wire _23598_;
wire _23599_;
wire _23600_;
wire _23601_;
wire _23602_;
wire _23603_;
wire _23604_;
wire _23605_;
wire _23606_;
wire _23607_;
wire _23608_;
wire _23609_;
wire _23610_;
wire _23611_;
wire _23612_;
wire _23613_;
wire _23614_;
wire _23615_;
wire _23616_;
wire _23617_;
wire _23618_;
wire _23619_;
wire _23620_;
wire _23621_;
wire _23622_;
wire _23623_;
wire _23624_;
wire _23625_;
wire _23626_;
wire _23627_;
wire _23628_;
wire _23629_;
wire _23630_;
wire _23631_;
wire _23632_;
wire _23633_;
wire _23634_;
wire _23635_;
wire _23636_;
wire _23637_;
wire _23638_;
wire _23639_;
wire _23640_;
wire _23641_;
wire _23642_;
wire _23643_;
wire _23644_;
wire _23645_;
wire _23646_;
wire _23647_;
wire _23648_;
wire _23649_;
wire _23650_;
wire _23651_;
wire _23652_;
wire _23653_;
wire _23654_;
wire _23655_;
wire _23656_;
wire _23657_;
wire _23658_;
wire _23659_;
wire _23660_;
wire _23661_;
wire _23662_;
wire _23663_;
wire _23664_;
wire _23665_;
wire _23666_;
wire _23667_;
wire _23668_;
wire _23669_;
wire _23670_;
wire _23671_;
wire _23672_;
wire _23673_;
wire _23674_;
wire _23675_;
wire _23676_;
wire _23677_;
wire _23678_;
wire _23679_;
wire _23680_;
wire _23681_;
wire _23682_;
wire _23683_;
wire _23684_;
wire _23685_;
wire _23686_;
wire _23687_;
wire _23688_;
wire _23689_;
wire _23690_;
wire _23691_;
wire _23692_;
wire _23693_;
wire _23694_;
wire _23695_;
wire _23696_;
wire _23697_;
wire _23698_;
wire _23699_;
wire _23700_;
wire _23701_;
wire _23702_;
wire _23703_;
wire _23704_;
wire _23705_;
wire _23706_;
wire _23707_;
wire _23708_;
wire _23709_;
wire _23710_;
wire _23711_;
wire _23712_;
wire _23713_;
wire _23714_;
wire _23715_;
wire _23716_;
wire _23717_;
wire _23718_;
wire _23719_;
wire _23720_;
wire _23721_;
wire _23722_;
wire _23723_;
wire _23724_;
wire _23725_;
wire _23726_;
wire _23727_;
wire _23728_;
wire _23729_;
wire _23730_;
wire _23731_;
wire _23732_;
wire _23733_;
wire _23734_;
wire _23735_;
wire _23736_;
wire _23737_;
wire _23738_;
wire _23739_;
wire _23740_;
wire _23741_;
wire _23742_;
wire _23743_;
wire _23744_;
wire _23745_;
wire _23746_;
wire _23747_;
wire _23748_;
wire _23749_;
wire _23750_;
wire _23751_;
wire _23752_;
wire _23753_;
wire _23754_;
wire _23755_;
wire _23756_;
wire _23757_;
wire _23758_;
wire _23759_;
wire _23760_;
wire _23761_;
wire _23762_;
wire _23763_;
wire _23764_;
wire _23765_;
wire _23766_;
wire _23767_;
wire _23768_;
wire _23769_;
wire _23770_;
wire _23771_;
wire _23772_;
wire _23773_;
wire _23774_;
wire _23775_;
wire _23776_;
wire _23777_;
wire _23778_;
wire _23779_;
wire _23780_;
wire _23781_;
wire _23782_;
wire _23783_;
wire _23784_;
wire _23785_;
wire _23786_;
wire _23787_;
wire _23788_;
wire _23789_;
wire _23790_;
wire _23791_;
wire _23792_;
wire _23793_;
wire _23794_;
wire _23795_;
wire _23796_;
wire _23797_;
wire _23798_;
wire _23799_;
wire _23800_;
wire _23801_;
wire _23802_;
wire _23803_;
wire _23804_;
wire _23805_;
wire _23806_;
wire _23807_;
wire _23808_;
wire _23809_;
wire _23810_;
wire _23811_;
wire _23812_;
wire _23813_;
wire _23814_;
wire _23815_;
wire _23816_;
wire _23817_;
wire _23818_;
wire _23819_;
wire _23820_;
wire _23821_;
wire _23822_;
wire _23823_;
wire _23824_;
wire _23825_;
wire _23826_;
wire _23827_;
wire _23828_;
wire _23829_;
wire _23830_;
wire _23831_;
wire _23832_;
wire _23833_;
wire _23834_;
wire _23835_;
wire _23836_;
wire _23837_;
wire _23838_;
wire _23839_;
wire _23840_;
wire _23841_;
wire _23842_;
wire _23843_;
wire _23844_;
wire _23845_;
wire _23846_;
wire _23847_;
wire _23848_;
wire _23849_;
wire _23850_;
wire _23851_;
wire _23852_;
wire _23853_;
wire _23854_;
wire _23855_;
wire _23856_;
wire _23857_;
wire _23858_;
wire _23859_;
wire _23860_;
wire _23861_;
wire _23862_;
wire _23863_;
wire _23864_;
wire _23865_;
wire _23866_;
wire _23867_;
wire _23868_;
wire _23869_;
wire _23870_;
wire _23871_;
wire _23872_;
wire _23873_;
wire _23874_;
wire _23875_;
wire _23876_;
wire _23877_;
wire _23878_;
wire _23879_;
wire _23880_;
wire _23881_;
wire _23882_;
wire _23883_;
wire _23884_;
wire _23885_;
wire _23886_;
wire _23887_;
wire _23888_;
wire _23889_;
wire _23890_;
wire _23891_;
wire _23892_;
wire _23893_;
wire _23894_;
wire _23895_;
wire _23896_;
wire _23897_;
wire _23898_;
wire _23899_;
wire _23900_;
wire _23901_;
wire _23902_;
wire _23903_;
wire _23904_;
wire _23905_;
wire _23906_;
wire _23907_;
wire _23908_;
wire _23909_;
wire _23910_;
wire _23911_;
wire _23912_;
wire _23913_;
wire _23914_;
wire _23915_;
wire _23916_;
wire _23917_;
wire _23918_;
wire _23919_;
wire _23920_;
wire _23921_;
wire _23922_;
wire _23923_;
wire _23924_;
wire _23925_;
wire _23926_;
wire _23927_;
wire _23928_;
wire _23929_;
wire _23930_;
wire _23931_;
wire _23932_;
wire _23933_;
wire _23934_;
wire _23935_;
wire _23936_;
wire _23937_;
wire _23938_;
wire _23939_;
wire _23940_;
wire _23941_;
wire _23942_;
wire _23943_;
wire _23944_;
wire _23945_;
wire _23946_;
wire _23947_;
wire _23948_;
wire _23949_;
wire _23950_;
wire _23951_;
wire _23952_;
wire _23953_;
wire _23954_;
wire _23955_;
wire _23956_;
wire _23957_;
wire _23958_;
wire _23959_;
wire _23960_;
wire _23961_;
wire _23962_;
wire _23963_;
wire _23964_;
wire _23965_;
wire _23966_;
wire _23967_;
wire _23968_;
wire _23969_;
wire _23970_;
wire _23971_;
wire _23972_;
wire _23973_;
wire _23974_;
wire _23975_;
wire _23976_;
wire _23977_;
wire _23978_;
wire _23979_;
wire _23980_;
wire _23981_;
wire _23982_;
wire _23983_;
wire _23984_;
wire _23985_;
wire _23986_;
wire _23987_;
wire _23988_;
wire _23989_;
wire _23990_;
wire _23991_;
wire _23992_;
wire _23993_;
wire _23994_;
wire _23995_;
wire _23996_;
wire _23997_;
wire _23998_;
wire _23999_;
wire _24000_;
wire _24001_;
wire _24002_;
wire _24003_;
wire _24004_;
wire _24005_;
wire _24006_;
wire _24007_;
wire _24008_;
wire _24009_;
wire _24010_;
wire _24011_;
wire _24012_;
wire _24013_;
wire _24014_;
wire _24015_;
wire _24016_;
wire _24017_;
wire _24018_;
wire _24019_;
wire _24020_;
wire _24021_;
wire _24022_;
wire _24023_;
wire _24024_;
wire _24025_;
wire _24026_;
wire _24027_;
wire _24028_;
wire _24029_;
wire _24030_;
wire _24031_;
wire _24032_;
wire _24033_;
wire _24034_;
wire _24035_;
wire _24036_;
wire _24037_;
wire _24038_;
wire _24039_;
wire _24040_;
wire _24041_;
wire _24042_;
wire _24043_;
wire _24044_;
wire _24045_;
wire _24046_;
wire _24047_;
wire _24048_;
wire _24049_;
wire _24050_;
wire _24051_;
wire _24052_;
wire _24053_;
wire _24054_;
wire _24055_;
wire _24056_;
wire _24057_;
wire _24058_;
wire _24059_;
wire _24060_;
wire _24061_;
wire _24062_;
wire _24063_;
wire _24064_;
wire _24065_;
wire _24066_;
wire _24067_;
wire _24068_;
wire _24069_;
wire _24070_;
wire _24071_;
wire _24072_;
wire _24073_;
wire _24074_;
wire _24075_;
wire _24076_;
wire _24077_;
wire _24078_;
wire _24079_;
wire _24080_;
wire _24081_;
wire _24082_;
wire _24083_;
wire _24084_;
wire _24085_;
wire _24086_;
wire _24087_;
wire _24088_;
wire _24089_;
wire _24090_;
wire _24091_;
wire _24092_;
wire _24093_;
wire _24094_;
wire _24095_;
wire _24096_;
wire _24097_;
wire _24098_;
wire _24099_;
wire _24100_;
wire _24101_;
wire _24102_;
wire _24103_;
wire _24104_;
wire _24105_;
wire _24106_;
wire _24107_;
wire _24108_;
wire _24109_;
wire _24110_;
wire _24111_;
wire _24112_;
wire _24113_;
wire _24114_;
wire _24115_;
wire _24116_;
wire _24117_;
wire _24118_;
wire _24119_;
wire _24120_;
wire _24121_;
wire _24122_;
wire _24123_;
wire _24124_;
wire _24125_;
wire _24126_;
wire _24127_;
wire _24128_;
wire _24129_;
wire _24130_;
wire _24131_;
wire _24132_;
wire _24133_;
wire _24134_;
wire _24135_;
wire _24136_;
wire _24137_;
wire _24138_;
wire _24139_;
wire _24140_;
wire _24141_;
wire _24142_;
wire _24143_;
wire _24144_;
wire _24145_;
wire _24146_;
wire _24147_;
wire _24148_;
wire _24149_;
wire _24150_;
wire _24151_;
wire _24152_;
wire _24153_;
wire _24154_;
wire _24155_;
wire _24156_;
wire _24157_;
wire _24158_;
wire _24159_;
wire _24160_;
wire _24161_;
wire _24162_;
wire _24163_;
wire _24164_;
wire _24165_;
wire _24166_;
wire _24167_;
wire _24168_;
wire _24169_;
wire _24170_;
wire _24171_;
wire _24172_;
wire _24173_;
wire _24174_;
wire _24175_;
wire _24176_;
wire _24177_;
wire _24178_;
wire _24179_;
wire _24180_;
wire _24181_;
wire _24182_;
wire _24183_;
wire _24184_;
wire _24185_;
wire _24186_;
wire _24187_;
wire _24188_;
wire _24189_;
wire _24190_;
wire _24191_;
wire _24192_;
wire _24193_;
wire _24194_;
wire _24195_;
wire _24196_;
wire _24197_;
wire _24198_;
wire _24199_;
wire _24200_;
wire _24201_;
wire _24202_;
wire _24203_;
wire _24204_;
wire _24205_;
wire _24206_;
wire _24207_;
wire _24208_;
wire _24209_;
wire _24210_;
wire _24211_;
wire _24212_;
wire _24213_;
wire _24214_;
wire _24215_;
wire _24216_;
wire _24217_;
wire _24218_;
wire _24219_;
wire _24220_;
wire _24221_;
wire _24222_;
wire _24223_;
wire _24224_;
wire _24225_;
wire _24226_;
wire _24227_;
wire _24228_;
wire _24229_;
wire _24230_;
wire _24231_;
wire _24232_;
wire _24233_;
wire _24234_;
wire _24235_;
wire _24236_;
wire _24237_;
wire _24238_;
wire _24239_;
wire _24240_;
wire _24241_;
wire _24242_;
wire _24243_;
wire _24244_;
wire _24245_;
wire _24246_;
wire _24247_;
wire _24248_;
wire _24249_;
wire _24250_;
wire _24251_;
wire _24252_;
wire _24253_;
wire _24254_;
wire _24255_;
wire _24256_;
wire _24257_;
wire _24258_;
wire _24259_;
wire _24260_;
wire _24261_;
wire _24262_;
wire _24263_;
wire _24264_;
wire _24265_;
wire _24266_;
wire _24267_;
wire _24268_;
wire _24269_;
wire _24270_;
wire _24271_;
wire _24272_;
wire _24273_;
wire _24274_;
wire _24275_;
wire _24276_;
wire _24277_;
wire _24278_;
wire _24279_;
wire _24280_;
wire _24281_;
wire _24282_;
wire _24283_;
wire _24284_;
wire _24285_;
wire _24286_;
wire _24287_;
wire _24288_;
wire _24289_;
wire _24290_;
wire _24291_;
wire _24292_;
wire _24293_;
wire _24294_;
wire _24295_;
wire _24296_;
wire _24297_;
wire _24298_;
wire _24299_;
wire _24300_;
wire _24301_;
wire _24302_;
wire _24303_;
wire _24304_;
wire _24305_;
wire _24306_;
wire _24307_;
wire _24308_;
wire _24309_;
wire _24310_;
wire _24311_;
wire _24312_;
wire _24313_;
wire _24314_;
wire _24315_;
wire _24316_;
wire _24317_;
wire _24318_;
wire _24319_;
wire _24320_;
wire _24321_;
wire _24322_;
wire _24323_;
wire _24324_;
wire _24325_;
wire _24326_;
wire _24327_;
wire _24328_;
wire _24329_;
wire _24330_;
wire _24331_;
wire _24332_;
wire _24333_;
wire _24334_;
wire _24335_;
wire _24336_;
wire _24337_;
wire _24338_;
wire _24339_;
wire _24340_;
wire _24341_;
wire _24342_;
wire _24343_;
wire _24344_;
wire _24345_;
wire _24346_;
wire _24347_;
wire _24348_;
wire _24349_;
wire _24350_;
wire _24351_;
wire _24352_;
wire _24353_;
wire _24354_;
wire _24355_;
wire _24356_;
wire _24357_;
wire _24358_;
wire _24359_;
wire _24360_;
wire _24361_;
wire _24362_;
wire _24363_;
wire _24364_;
wire _24365_;
wire _24366_;
wire _24367_;
wire _24368_;
wire _24369_;
wire _24370_;
wire _24371_;
wire _24372_;
wire _24373_;
wire _24374_;
wire _24375_;
wire _24376_;
wire _24377_;
wire _24378_;
wire _24379_;
wire _24380_;
wire _24381_;
wire _24382_;
wire _24383_;
wire _24384_;
wire _24385_;
wire _24386_;
wire _24387_;
wire _24388_;
wire _24389_;
wire _24390_;
wire _24391_;
wire _24392_;
wire _24393_;
wire _24394_;
wire _24395_;
wire _24396_;
wire _24397_;
wire _24398_;
wire _24399_;
wire _24400_;
wire _24401_;
wire _24402_;
wire _24403_;
wire _24404_;
wire _24405_;
wire _24406_;
wire _24407_;
wire _24408_;
wire _24409_;
wire _24410_;
wire _24411_;
wire _24412_;
wire _24413_;
wire _24414_;
wire _24415_;
wire _24416_;
wire _24417_;
wire _24418_;
wire _24419_;
wire _24420_;
wire _24421_;
wire _24422_;
wire _24423_;
wire _24424_;
wire _24425_;
wire _24426_;
wire _24427_;
wire _24428_;
wire _24429_;
wire _24430_;
wire _24431_;
wire _24432_;
wire _24433_;
wire _24434_;
wire _24435_;
wire _24436_;
wire _24437_;
wire _24438_;
wire _24439_;
wire _24440_;
wire _24441_;
wire _24442_;
wire _24443_;
wire _24444_;
wire _24445_;
wire _24446_;
wire _24447_;
wire _24448_;
wire _24449_;
wire _24450_;
wire _24451_;
wire _24452_;
wire _24453_;
wire _24454_;
wire _24455_;
wire _24456_;
wire _24457_;
wire _24458_;
wire _24459_;
wire _24460_;
wire _24461_;
wire _24462_;
wire _24463_;
wire _24464_;
wire _24465_;
wire _24466_;
wire _24467_;
wire _24468_;
wire _24469_;
wire _24470_;
wire _24471_;
wire _24472_;
wire _24473_;
wire _24474_;
wire _24475_;
wire _24476_;
wire _24477_;
wire _24478_;
wire _24479_;
wire _24480_;
wire _24481_;
wire _24482_;
wire _24483_;
wire _24484_;
wire _24485_;
wire _24486_;
wire _24487_;
wire _24488_;
wire _24489_;
wire _24490_;
wire _24491_;
wire _24492_;
wire _24493_;
wire _24494_;
wire _24495_;
wire _24496_;
wire _24497_;
wire _24498_;
wire _24499_;
wire _24500_;
wire _24501_;
wire _24502_;
wire _24503_;
wire _24504_;
wire _24505_;
wire _24506_;
wire _24507_;
wire _24508_;
wire _24509_;
wire _24510_;
wire _24511_;
wire _24512_;
wire _24513_;
wire _24514_;
wire _24515_;
wire _24516_;
wire _24517_;
wire _24518_;
wire _24519_;
wire _24520_;
wire _24521_;
wire _24522_;
wire _24523_;
wire _24524_;
wire _24525_;
wire _24526_;
wire _24527_;
wire _24528_;
wire _24529_;
wire _24530_;
wire _24531_;
wire _24532_;
wire _24533_;
wire _24534_;
wire _24535_;
wire _24536_;
wire _24537_;
wire _24538_;
wire _24539_;
wire _24540_;
wire _24541_;
wire _24542_;
wire _24543_;
wire _24544_;
wire _24545_;
wire _24546_;
wire _24547_;
wire _24548_;
wire _24549_;
wire _24550_;
wire _24551_;
wire _24552_;
wire _24553_;
wire _24554_;
wire _24555_;
wire _24556_;
wire _24557_;
wire _24558_;
wire _24559_;
wire _24560_;
wire _24561_;
wire _24562_;
wire _24563_;
wire _24564_;
wire _24565_;
wire _24566_;
wire _24567_;
wire _24568_;
wire _24569_;
wire _24570_;
wire _24571_;
wire _24572_;
wire _24573_;
wire _24574_;
wire _24575_;
wire _24576_;
wire _24577_;
wire _24578_;
wire _24579_;
wire _24580_;
wire _24581_;
wire _24582_;
wire _24583_;
wire _24584_;
wire _24585_;
wire _24586_;
wire _24587_;
wire _24588_;
wire _24589_;
wire _24590_;
wire _24591_;
wire _24592_;
wire _24593_;
wire _24594_;
wire _24595_;
wire _24596_;
wire _24597_;
wire _24598_;
wire _24599_;
wire _24600_;
wire _24601_;
wire _24602_;
wire _24603_;
wire _24604_;
wire _24605_;
wire _24606_;
wire _24607_;
wire _24608_;
wire _24609_;
wire _24610_;
wire _24611_;
wire _24612_;
wire _24613_;
wire _24614_;
wire _24615_;
wire _24616_;
wire _24617_;
wire _24618_;
wire _24619_;
wire _24620_;
wire _24621_;
wire _24622_;
wire _24623_;
wire _24624_;
wire _24625_;
wire _24626_;
wire _24627_;
wire _24628_;
wire _24629_;
wire _24630_;
wire _24631_;
wire _24632_;
wire _24633_;
wire _24634_;
wire _24635_;
wire _24636_;
wire _24637_;
wire _24638_;
wire _24639_;
wire _24640_;
wire _24641_;
wire _24642_;
wire _24643_;
wire _24644_;
wire _24645_;
wire _24646_;
wire _24647_;
wire _24648_;
wire _24649_;
wire _24650_;
wire _24651_;
wire _24652_;
wire _24653_;
wire _24654_;
wire _24655_;
wire _24656_;
wire _24657_;
wire _24658_;
wire _24659_;
wire _24660_;
wire _24661_;
wire _24662_;
wire _24663_;
wire _24664_;
wire _24665_;
wire _24666_;
wire _24667_;
wire _24668_;
wire _24669_;
wire _24670_;
wire _24671_;
wire _24672_;
wire _24673_;
wire _24674_;
wire _24675_;
wire _24676_;
wire _24677_;
wire _24678_;
wire _24679_;
wire _24680_;
wire _24681_;
wire _24682_;
wire _24683_;
wire _24684_;
wire _24685_;
wire _24686_;
wire _24687_;
wire _24688_;
wire _24689_;
wire _24690_;
wire _24691_;
wire _24692_;
wire _24693_;
wire _24694_;
wire _24695_;
wire _24696_;
wire _24697_;
wire _24698_;
wire _24699_;
wire _24700_;
wire _24701_;
wire _24702_;
wire _24703_;
wire _24704_;
wire _24705_;
wire _24706_;
wire _24707_;
wire _24708_;
wire _24709_;
wire _24710_;
wire _24711_;
wire _24712_;
wire _24713_;
wire _24714_;
wire _24715_;
wire _24716_;
wire _24717_;
wire _24718_;
wire _24719_;
wire _24720_;
wire _24721_;
wire _24722_;
wire _24723_;
wire _24724_;
wire _24725_;
wire _24726_;
wire _24727_;
wire _24728_;
wire _24729_;
wire _24730_;
wire _24731_;
wire _24732_;
wire _24733_;
wire _24734_;
wire _24735_;
wire _24736_;
wire _24737_;
wire _24738_;
wire _24739_;
wire _24740_;
wire _24741_;
wire _24742_;
wire _24743_;
wire _24744_;
wire _24745_;
wire _24746_;
wire _24747_;
wire _24748_;
wire _24749_;
wire _24750_;
wire _24751_;
wire _24752_;
wire _24753_;
wire _24754_;
wire _24755_;
wire _24756_;
wire _24757_;
wire _24758_;
wire _24759_;
wire _24760_;
wire _24761_;
wire _24762_;
wire _24763_;
wire _24764_;
wire _24765_;
wire _24766_;
wire _24767_;
wire _24768_;
wire _24769_;
wire _24770_;
wire _24771_;
wire _24772_;
wire _24773_;
wire _24774_;
wire _24775_;
wire _24776_;
wire _24777_;
wire _24778_;
wire _24779_;
wire _24780_;
wire _24781_;
wire _24782_;
wire _24783_;
wire _24784_;
wire _24785_;
wire _24786_;
wire _24787_;
wire _24788_;
wire _24789_;
wire _24790_;
wire _24791_;
wire _24792_;
wire _24793_;
wire _24794_;
wire _24795_;
wire _24796_;
wire _24797_;
wire _24798_;
wire _24799_;
wire _24800_;
wire _24801_;
wire _24802_;
wire _24803_;
wire _24804_;
wire _24805_;
wire _24806_;
wire _24807_;
wire _24808_;
wire _24809_;
wire _24810_;
wire _24811_;
wire _24812_;
wire _24813_;
wire _24814_;
wire _24815_;
wire _24816_;
wire _24817_;
wire _24818_;
wire _24819_;
wire _24820_;
wire _24821_;
wire _24822_;
wire _24823_;
wire _24824_;
wire _24825_;
wire _24826_;
wire _24827_;
wire _24828_;
wire _24829_;
wire _24830_;
wire _24831_;
wire _24832_;
wire _24833_;
wire _24834_;
wire _24835_;
wire _24836_;
wire _24837_;
wire _24838_;
wire _24839_;
wire _24840_;
wire _24841_;
wire _24842_;
wire _24843_;
wire _24844_;
wire _24845_;
wire _24846_;
wire _24847_;
wire _24848_;
wire _24849_;
wire _24850_;
wire _24851_;
wire _24852_;
wire _24853_;
wire _24854_;
wire _24855_;
wire _24856_;
wire _24857_;
wire _24858_;
wire _24859_;
wire _24860_;
wire _24861_;
wire _24862_;
wire _24863_;
wire _24864_;
wire _24865_;
wire _24866_;
wire _24867_;
wire _24868_;
wire _24869_;
wire _24870_;
wire _24871_;
wire _24872_;
wire _24873_;
wire _24874_;
wire _24875_;
wire _24876_;
wire _24877_;
wire _24878_;
wire _24879_;
wire _24880_;
wire _24881_;
wire _24882_;
wire _24883_;
wire _24884_;
wire _24885_;
wire _24886_;
wire _24887_;
wire _24888_;
wire _24889_;
wire _24890_;
wire _24891_;
wire _24892_;
wire _24893_;
wire _24894_;
wire _24895_;
wire _24896_;
wire _24897_;
wire _24898_;
wire _24899_;
wire _24900_;
wire _24901_;
wire _24902_;
wire _24903_;
wire _24904_;
wire _24905_;
wire _24906_;
wire _24907_;
wire _24908_;
wire _24909_;
wire _24910_;
wire _24911_;
wire _24912_;
wire _24913_;
wire _24914_;
wire _24915_;
wire _24916_;
wire _24917_;
wire _24918_;
wire _24919_;
wire _24920_;
wire _24921_;
wire _24922_;
wire _24923_;
wire _24924_;
wire _24925_;
wire _24926_;
wire _24927_;
wire _24928_;
wire _24929_;
wire _24930_;
wire _24931_;
wire _24932_;
wire _24933_;
wire _24934_;
wire _24935_;
wire _24936_;
wire _24937_;
wire _24938_;
wire _24939_;
wire _24940_;
wire _24941_;
wire _24942_;
wire _24943_;
wire _24944_;
wire _24945_;
wire _24946_;
wire _24947_;
wire _24948_;
wire _24949_;
wire _24950_;
wire _24951_;
wire _24952_;
wire _24953_;
wire _24954_;
wire _24955_;
wire _24956_;
wire _24957_;
wire _24958_;
wire _24959_;
wire _24960_;
wire _24961_;
wire _24962_;
wire _24963_;
wire _24964_;
wire _24965_;
wire _24966_;
wire _24967_;
wire _24968_;
wire _24969_;
wire _24970_;
wire _24971_;
wire _24972_;
wire _24973_;
wire _24974_;
wire _24975_;
wire _24976_;
wire _24977_;
wire _24978_;
wire _24979_;
wire _24980_;
wire _24981_;
wire _24982_;
wire _24983_;
wire _24984_;
wire _24985_;
wire _24986_;
wire _24987_;
wire _24988_;
wire _24989_;
wire _24990_;
wire _24991_;
wire _24992_;
wire _24993_;
wire _24994_;
wire _24995_;
wire _24996_;
wire _24997_;
wire _24998_;
wire _24999_;
wire _25000_;
wire _25001_;
wire _25002_;
wire _25003_;
wire _25004_;
wire _25005_;
wire _25006_;
wire _25007_;
wire _25008_;
wire _25009_;
wire _25010_;
wire _25011_;
wire _25012_;
wire _25013_;
wire _25014_;
wire _25015_;
wire _25016_;
wire _25017_;
wire _25018_;
wire _25019_;
wire _25020_;
wire _25021_;
wire _25022_;
wire _25023_;
wire _25024_;
wire _25025_;
wire _25026_;
wire _25027_;
wire _25028_;
wire _25029_;
wire _25030_;
wire _25031_;
wire _25032_;
wire _25033_;
wire _25034_;
wire _25035_;
wire _25036_;
wire _25037_;
wire _25038_;
wire _25039_;
wire _25040_;
wire _25041_;
wire _25042_;
wire _25043_;
wire _25044_;
wire _25045_;
wire _25046_;
wire _25047_;
wire _25048_;
wire _25049_;
wire _25050_;
wire _25051_;
wire _25052_;
wire _25053_;
wire _25054_;
wire _25055_;
wire _25056_;
wire _25057_;
wire _25058_;
wire _25059_;
wire _25060_;
wire _25061_;
wire _25062_;
wire _25063_;
wire _25064_;
wire _25065_;
wire _25066_;
wire _25067_;
wire _25068_;
wire _25069_;
wire _25070_;
wire _25071_;
wire _25072_;
wire _25073_;
wire _25074_;
wire _25075_;
wire _25076_;
wire _25077_;
wire _25078_;
wire _25079_;
wire _25080_;
wire _25081_;
wire _25082_;
wire _25083_;
wire _25084_;
wire _25085_;
wire _25086_;
wire _25087_;
wire _25088_;
wire _25089_;
wire _25090_;
wire _25091_;
wire _25092_;
wire _25093_;
wire _25094_;
wire _25095_;
wire _25096_;
wire _25097_;
wire _25098_;
wire _25099_;
wire _25100_;
wire _25101_;
wire _25102_;
wire _25103_;
wire _25104_;
wire _25105_;
wire _25106_;
wire _25107_;
wire _25108_;
wire _25109_;
wire _25110_;
wire _25111_;
wire _25112_;
wire _25113_;
wire _25114_;
wire _25115_;
wire _25116_;
wire _25117_;
wire _25118_;
wire _25119_;
wire _25120_;
wire _25121_;
wire _25122_;
wire _25123_;
wire _25124_;
wire _25125_;
wire _25126_;
wire _25127_;
wire _25128_;
wire _25129_;
wire _25130_;
wire _25131_;
wire _25132_;
wire _25133_;
wire _25134_;
wire _25135_;
wire _25136_;
wire _25137_;
wire _25138_;
wire _25139_;
wire _25140_;
wire _25141_;
wire _25142_;
wire _25143_;
wire _25144_;
wire _25145_;
wire _25146_;
wire _25147_;
wire _25148_;
wire _25149_;
wire _25150_;
wire _25151_;
wire _25152_;
wire _25153_;
wire _25154_;
wire _25155_;
wire _25156_;
wire _25157_;
wire _25158_;
wire _25159_;
wire _25160_;
wire _25161_;
wire _25162_;
wire _25163_;
wire _25164_;
wire _25165_;
wire _25166_;
wire _25167_;
wire _25168_;
wire _25169_;
wire _25170_;
wire _25171_;
wire _25172_;
wire _25173_;
wire _25174_;
wire _25175_;
wire _25176_;
wire _25177_;
wire _25178_;
wire _25179_;
wire _25180_;
wire _25181_;
wire _25182_;
wire _25183_;
wire _25184_;
wire _25185_;
wire _25186_;
wire _25187_;
wire _25188_;
wire _25189_;
wire _25190_;
wire _25191_;
wire _25192_;
wire _25193_;
wire _25194_;
wire _25195_;
wire _25196_;
wire _25197_;
wire _25198_;
wire _25199_;
wire _25200_;
wire _25201_;
wire _25202_;
wire _25203_;
wire _25204_;
wire _25205_;
wire _25206_;
wire _25207_;
wire _25208_;
wire _25209_;
wire _25210_;
wire _25211_;
wire _25212_;
wire _25213_;
wire _25214_;
wire _25215_;
wire _25216_;
wire _25217_;
wire _25218_;
wire _25219_;
wire _25220_;
wire _25221_;
wire _25222_;
wire _25223_;
wire _25224_;
wire _25225_;
wire _25226_;
wire _25227_;
wire _25228_;
wire _25229_;
wire _25230_;
wire _25231_;
wire _25232_;
wire _25233_;
wire _25234_;
wire _25235_;
wire _25236_;
wire _25237_;
wire _25238_;
wire _25239_;
wire _25240_;
wire _25241_;
wire _25242_;
wire _25243_;
wire _25244_;
wire _25245_;
wire _25246_;
wire _25247_;
wire _25248_;
wire _25249_;
wire _25250_;
wire _25251_;
wire _25252_;
wire _25253_;
wire _25254_;
wire _25255_;
wire _25256_;
wire _25257_;
wire _25258_;
wire _25259_;
wire _25260_;
wire _25261_;
wire _25262_;
wire _25263_;
wire _25264_;
wire _25265_;
wire _25266_;
wire _25267_;
wire _25268_;
wire _25269_;
wire _25270_;
wire _25271_;
wire _25272_;
wire _25273_;
wire _25274_;
wire _25275_;
wire _25276_;
wire _25277_;
wire _25278_;
wire _25279_;
wire _25280_;
wire _25281_;
wire _25282_;
wire _25283_;
wire _25284_;
wire _25285_;
wire _25286_;
wire _25287_;
wire _25288_;
wire _25289_;
wire _25290_;
wire _25291_;
wire _25292_;
wire _25293_;
wire _25294_;
wire _25295_;
wire _25296_;
wire _25297_;
wire _25298_;
wire _25299_;
wire _25300_;
wire _25301_;
wire _25302_;
wire _25303_;
wire _25304_;
wire _25305_;
wire _25306_;
wire _25307_;
wire _25308_;
wire _25309_;
wire _25310_;
wire _25311_;
wire _25312_;
wire _25313_;
wire _25314_;
wire _25315_;
wire _25316_;
wire _25317_;
wire _25318_;
wire _25319_;
wire _25320_;
wire _25321_;
wire _25322_;
wire _25323_;
wire _25324_;
wire _25325_;
wire _25326_;
wire _25327_;
wire _25328_;
wire _25329_;
wire _25330_;
wire _25331_;
wire _25332_;
wire _25333_;
wire _25334_;
wire _25335_;
wire _25336_;
wire _25337_;
wire _25338_;
wire _25339_;
wire _25340_;
wire _25341_;
wire _25342_;
wire _25343_;
wire _25344_;
wire _25345_;
wire _25346_;
wire _25347_;
wire _25348_;
wire _25349_;
wire _25350_;
wire _25351_;
wire _25352_;
wire _25353_;
wire _25354_;
wire _25355_;
wire _25356_;
wire _25357_;
wire _25358_;
wire _25359_;
wire _25360_;
wire _25361_;
wire _25362_;
wire _25363_;
wire _25364_;
wire _25365_;
wire _25366_;
wire _25367_;
wire _25368_;
wire _25369_;
wire _25370_;
wire _25371_;
wire _25372_;
wire _25373_;
wire _25374_;
wire _25375_;
wire _25376_;
wire _25377_;
wire _25378_;
wire _25379_;
wire _25380_;
wire _25381_;
wire _25382_;
wire _25383_;
wire _25384_;
wire _25385_;
wire _25386_;
wire _25387_;
wire _25388_;
wire _25389_;
wire _25390_;
wire _25391_;
wire _25392_;
wire _25393_;
wire _25394_;
wire _25395_;
wire _25396_;
wire _25397_;
wire _25398_;
wire _25399_;
wire _25400_;
wire _25401_;
wire _25402_;
wire _25403_;
wire _25404_;
wire _25405_;
wire _25406_;
wire _25407_;
wire _25408_;
wire _25409_;
wire _25410_;
wire _25411_;
wire _25412_;
wire _25413_;
wire _25414_;
wire _25415_;
wire _25416_;
wire _25417_;
wire _25418_;
wire _25419_;
wire _25420_;
wire _25421_;
wire _25422_;
wire _25423_;
wire _25424_;
wire _25425_;
wire _25426_;
wire _25427_;
wire _25428_;
wire _25429_;
wire _25430_;
wire _25431_;
wire _25432_;
wire _25433_;
wire _25434_;
wire _25435_;
wire _25436_;
wire _25437_;
wire _25438_;
wire _25439_;
wire _25440_;
wire _25441_;
wire _25442_;
wire _25443_;
wire _25444_;
wire _25445_;
wire _25446_;
wire _25447_;
wire _25448_;
wire _25449_;
wire _25450_;
wire _25451_;
wire _25452_;
wire _25453_;
wire _25454_;
wire _25455_;
wire _25456_;
wire _25457_;
wire _25458_;
wire _25459_;
wire _25460_;
wire _25461_;
wire _25462_;
wire _25463_;
wire _25464_;
wire _25465_;
wire _25466_;
wire _25467_;
wire _25468_;
wire _25469_;
wire _25470_;
wire _25471_;
wire _25472_;
wire _25473_;
wire _25474_;
wire _25475_;
wire _25476_;
wire _25477_;
wire _25478_;
wire _25479_;
wire _25480_;
wire _25481_;
wire _25482_;
wire _25483_;
wire _25484_;
wire _25485_;
wire _25486_;
wire _25487_;
wire _25488_;
wire _25489_;
wire _25490_;
wire _25491_;
wire _25492_;
wire _25493_;
wire _25494_;
wire _25495_;
wire _25496_;
wire _25497_;
wire _25498_;
wire _25499_;
wire _25500_;
wire _25501_;
wire _25502_;
wire _25503_;
wire _25504_;
wire _25505_;
wire _25506_;
wire _25507_;
wire _25508_;
wire _25509_;
wire _25510_;
wire _25511_;
wire _25512_;
wire _25513_;
wire _25514_;
wire _25515_;
wire _25516_;
wire _25517_;
wire _25518_;
wire _25519_;
wire _25520_;
wire _25521_;
wire _25522_;
wire _25523_;
wire _25524_;
wire _25525_;
wire _25526_;
wire _25527_;
wire _25528_;
wire _25529_;
wire _25530_;
wire _25531_;
wire _25532_;
wire _25533_;
wire _25534_;
wire _25535_;
wire _25536_;
wire _25537_;
wire _25538_;
wire _25539_;
wire _25540_;
wire _25541_;
wire _25542_;
wire _25543_;
wire _25544_;
wire _25545_;
wire _25546_;
wire _25547_;
wire _25548_;
wire _25549_;
wire _25550_;
wire _25551_;
wire _25552_;
wire _25553_;
wire _25554_;
wire _25555_;
wire _25556_;
wire _25557_;
wire _25558_;
wire _25559_;
wire _25560_;
wire _25561_;
wire _25562_;
wire _25563_;
wire _25564_;
wire _25565_;
wire _25566_;
wire _25567_;
wire _25568_;
wire _25569_;
wire _25570_;
wire _25571_;
wire _25572_;
wire _25573_;
wire _25574_;
wire _25575_;
wire _25576_;
wire _25577_;
wire _25578_;
wire _25579_;
wire _25580_;
wire _25581_;
wire _25582_;
wire _25583_;
wire _25584_;
wire _25585_;
wire _25586_;
wire _25587_;
wire _25588_;
wire _25589_;
wire _25590_;
wire _25591_;
wire _25592_;
wire _25593_;
wire _25594_;
wire _25595_;
wire _25596_;
wire _25597_;
wire _25598_;
wire _25599_;
wire _25600_;
wire _25601_;
wire _25602_;
wire _25603_;
wire _25604_;
wire _25605_;
wire _25606_;
wire _25607_;
wire _25608_;
wire _25609_;
wire _25610_;
wire _25611_;
wire _25612_;
wire _25613_;
wire _25614_;
wire _25615_;
wire _25616_;
wire _25617_;
wire _25618_;
wire _25619_;
wire _25620_;
wire _25621_;
wire _25622_;
wire _25623_;
wire _25624_;
wire _25625_;
wire _25626_;
wire _25627_;
wire _25628_;
wire _25629_;
wire _25630_;
wire _25631_;
wire _25632_;
wire _25633_;
wire _25634_;
wire _25635_;
wire _25636_;
wire _25637_;
wire _25638_;
wire _25639_;
wire _25640_;
wire _25641_;
wire _25642_;
wire _25643_;
wire _25644_;
wire _25645_;
wire _25646_;
wire _25647_;
wire _25648_;
wire _25649_;
wire _25650_;
wire _25651_;
wire _25652_;
wire _25653_;
wire _25654_;
wire _25655_;
wire _25656_;
wire _25657_;
wire _25658_;
wire _25659_;
wire _25660_;
wire _25661_;
wire _25662_;
wire _25663_;
wire _25664_;
wire _25665_;
wire _25666_;
wire _25667_;
wire _25668_;
wire _25669_;
wire _25670_;
wire _25671_;
wire _25672_;
wire _25673_;
wire _25674_;
wire _25675_;
wire _25676_;
wire _25677_;
wire _25678_;
wire _25679_;
wire _25680_;
wire _25681_;
wire _25682_;
wire _25683_;
wire _25684_;
wire _25685_;
wire _25686_;
wire _25687_;
wire _25688_;
wire _25689_;
wire _25690_;
wire _25691_;
wire _25692_;
wire _25693_;
wire _25694_;
wire _25695_;
wire _25696_;
wire _25697_;
wire _25698_;
wire _25699_;
wire _25700_;
wire _25701_;
wire _25702_;
wire _25703_;
wire _25704_;
wire _25705_;
wire _25706_;
wire _25707_;
wire _25708_;
wire _25709_;
wire _25710_;
wire _25711_;
wire _25712_;
wire _25713_;
wire _25714_;
wire _25715_;
wire _25716_;
wire _25717_;
wire _25718_;
wire _25719_;
wire _25720_;
wire _25721_;
wire _25722_;
wire _25723_;
wire _25724_;
wire _25725_;
wire _25726_;
wire _25727_;
wire _25728_;
wire _25729_;
wire _25730_;
wire _25731_;
wire _25732_;
wire _25733_;
wire _25734_;
wire _25735_;
wire _25736_;
wire _25737_;
wire _25738_;
wire _25739_;
wire _25740_;
wire _25741_;
wire _25742_;
wire _25743_;
wire _25744_;
wire _25745_;
wire _25746_;
wire _25747_;
wire _25748_;
wire _25749_;
wire _25750_;
wire _25751_;
wire _25752_;
wire _25753_;
wire _25754_;
wire _25755_;
wire _25756_;
wire _25757_;
wire _25758_;
wire _25759_;
wire _25760_;
wire _25761_;
wire _25762_;
wire _25763_;
wire _25764_;
wire _25765_;
wire _25766_;
wire _25767_;
wire _25768_;
wire _25769_;
wire _25770_;
wire _25771_;
wire _25772_;
wire _25773_;
wire _25774_;
wire _25775_;
wire _25776_;
wire _25777_;
wire _25778_;
wire _25779_;
wire _25780_;
wire _25781_;
wire _25782_;
wire _25783_;
wire _25784_;
wire _25785_;
wire _25786_;
wire _25787_;
wire _25788_;
wire _25789_;
wire _25790_;
wire _25791_;
wire _25792_;
wire _25793_;
wire _25794_;
wire _25795_;
wire _25796_;
wire _25797_;
wire _25798_;
wire _25799_;
wire _25800_;
wire _25801_;
wire _25802_;
wire _25803_;
wire _25804_;
wire _25805_;
wire _25806_;
wire _25807_;
wire _25808_;
wire _25809_;
wire _25810_;
wire _25811_;
wire _25812_;
wire _25813_;
wire _25814_;
wire _25815_;
wire _25816_;
wire _25817_;
wire _25818_;
wire _25819_;
wire _25820_;
wire _25821_;
wire _25822_;
wire _25823_;
wire _25824_;
wire _25825_;
wire _25826_;
wire _25827_;
wire _25828_;
wire _25829_;
wire _25830_;
wire _25831_;
wire _25832_;
wire _25833_;
wire _25834_;
wire _25835_;
wire _25836_;
wire _25837_;
wire _25838_;
wire _25839_;
wire _25840_;
wire _25841_;
wire _25842_;
wire _25843_;
wire _25844_;
wire _25845_;
wire _25846_;
wire _25847_;
wire _25848_;
wire _25849_;
wire _25850_;
wire _25851_;
wire _25852_;
wire _25853_;
wire _25854_;
wire _25855_;
wire _25856_;
wire _25857_;
wire _25858_;
wire _25859_;
wire _25860_;
wire _25861_;
wire _25862_;
wire _25863_;
wire _25864_;
wire _25865_;
wire _25866_;
wire _25867_;
wire _25868_;
wire _25869_;
wire _25870_;
wire _25871_;
wire _25872_;
wire _25873_;
wire _25874_;
wire _25875_;
wire _25876_;
wire _25877_;
wire _25878_;
wire _25879_;
wire _25880_;
wire _25881_;
wire _25882_;
wire _25883_;
wire _25884_;
wire _25885_;
wire _25886_;
wire _25887_;
wire _25888_;
wire _25889_;
wire _25890_;
wire _25891_;
wire _25892_;
wire _25893_;
wire _25894_;
wire _25895_;
wire _25896_;
wire _25897_;
wire _25898_;
wire _25899_;
wire _25900_;
wire _25901_;
wire _25902_;
wire _25903_;
wire _25904_;
wire _25905_;
wire _25906_;
wire _25907_;
wire _25908_;
wire _25909_;
wire _25910_;
wire _25911_;
wire _25912_;
wire _25913_;
wire _25914_;
wire _25915_;
wire _25916_;
wire _25917_;
wire _25918_;
wire _25919_;
wire _25920_;
wire _25921_;
wire _25922_;
wire _25923_;
wire _25924_;
wire _25925_;
wire _25926_;
wire _25927_;
wire _25928_;
wire _25929_;
wire _25930_;
wire _25931_;
wire _25932_;
wire _25933_;
wire _25934_;
wire _25935_;
wire _25936_;
wire _25937_;
wire _25938_;
wire _25939_;
wire _25940_;
wire _25941_;
wire _25942_;
wire _25943_;
wire _25944_;
wire _25945_;
wire _25946_;
wire _25947_;
wire _25948_;
wire _25949_;
wire _25950_;
wire _25951_;
wire _25952_;
wire _25953_;
wire _25954_;
wire _25955_;
wire _25956_;
wire _25957_;
wire _25958_;
wire _25959_;
wire _25960_;
wire _25961_;
wire _25962_;
wire _25963_;
wire _25964_;
wire _25965_;
wire _25966_;
wire _25967_;
wire _25968_;
wire _25969_;
wire _25970_;
wire _25971_;
wire _25972_;
wire _25973_;
wire _25974_;
wire _25975_;
wire _25976_;
wire _25977_;
wire _25978_;
wire _25979_;
wire _25980_;
wire _25981_;
wire _25982_;
wire _25983_;
wire _25984_;
wire _25985_;
wire _25986_;
wire _25987_;
wire _25988_;
wire _25989_;
wire _25990_;
wire _25991_;
wire _25992_;
wire _25993_;
wire _25994_;
wire _25995_;
wire _25996_;
wire _25997_;
wire _25998_;
wire _25999_;
wire _26000_;
wire _26001_;
wire _26002_;
wire _26003_;
wire _26004_;
wire _26005_;
wire _26006_;
wire _26007_;
wire _26008_;
wire _26009_;
wire _26010_;
wire _26011_;
wire _26012_;
wire _26013_;
wire _26014_;
wire _26015_;
wire _26016_;
wire _26017_;
wire _26018_;
wire _26019_;
wire _26020_;
wire _26021_;
wire _26022_;
wire _26023_;
wire _26024_;
wire _26025_;
wire _26026_;
wire _26027_;
wire _26028_;
wire _26029_;
wire _26030_;
wire _26031_;
wire _26032_;
wire _26033_;
wire _26034_;
wire _26035_;
wire _26036_;
wire _26037_;
wire _26038_;
wire _26039_;
wire _26040_;
wire _26041_;
wire _26042_;
wire _26043_;
wire _26044_;
wire _26045_;
wire _26046_;
wire _26047_;
wire _26048_;
wire _26049_;
wire _26050_;
wire _26051_;
wire _26052_;
wire _26053_;
wire _26054_;
wire _26055_;
wire _26056_;
wire _26057_;
wire _26058_;
wire _26059_;
wire _26060_;
wire _26061_;
wire _26062_;
wire _26063_;
wire _26064_;
wire _26065_;
wire _26066_;
wire _26067_;
wire _26068_;
wire _26069_;
wire _26070_;
wire _26071_;
wire _26072_;
wire _26073_;
wire _26074_;
wire _26075_;
wire _26076_;
wire _26077_;
wire _26078_;
wire _26079_;
wire _26080_;
wire _26081_;
wire _26082_;
wire _26083_;
wire _26084_;
wire _26085_;
wire _26086_;
wire _26087_;
wire _26088_;
wire _26089_;
wire _26090_;
wire _26091_;
wire _26092_;
wire _26093_;
wire _26094_;
wire _26095_;
wire _26096_;
wire _26097_;
wire _26098_;
wire _26099_;
wire _26100_;
wire _26101_;
wire _26102_;
wire _26103_;
wire _26104_;
wire _26105_;
wire _26106_;
wire _26107_;
wire _26108_;
wire _26109_;
wire _26110_;
wire _26111_;
wire _26112_;
wire _26113_;
wire _26114_;
wire _26115_;
wire _26116_;
wire _26117_;
wire _26118_;
wire _26119_;
wire _26120_;
wire _26121_;
wire _26122_;
wire _26123_;
wire _26124_;
wire _26125_;
wire _26126_;
wire _26127_;
wire _26128_;
wire _26129_;
wire _26130_;
wire _26131_;
wire _26132_;
wire _26133_;
wire _26134_;
wire _26135_;
wire _26136_;
wire _26137_;
wire _26138_;
wire _26139_;
wire _26140_;
wire _26141_;
wire _26142_;
wire _26143_;
wire _26144_;
wire _26145_;
wire _26146_;
wire _26147_;
wire _26148_;
wire _26149_;
wire _26150_;
wire _26151_;
wire _26152_;
wire _26153_;
wire _26154_;
wire _26155_;
wire _26156_;
wire _26157_;
wire _26158_;
wire _26159_;
wire _26160_;
wire _26161_;
wire _26162_;
wire _26163_;
wire _26164_;
wire _26165_;
wire _26166_;
wire _26167_;
wire _26168_;
wire _26169_;
wire _26170_;
wire _26171_;
wire _26172_;
wire _26173_;
wire _26174_;
wire _26175_;
wire _26176_;
wire _26177_;
wire _26178_;
wire _26179_;
wire _26180_;
wire _26181_;
wire _26182_;
wire _26183_;
wire _26184_;
wire _26185_;
wire _26186_;
wire _26187_;
wire _26188_;
wire _26189_;
wire _26190_;
wire _26191_;
wire _26192_;
wire _26193_;
wire _26194_;
wire _26195_;
wire _26196_;
wire _26197_;
wire _26198_;
wire _26199_;
wire _26200_;
wire _26201_;
wire _26202_;
wire _26203_;
wire _26204_;
wire _26205_;
wire _26206_;
wire _26207_;
wire _26208_;
wire _26209_;
wire _26210_;
wire _26211_;
wire _26212_;
wire _26213_;
wire _26214_;
wire _26215_;
wire _26216_;
wire _26217_;
wire _26218_;
wire _26219_;
wire _26220_;
wire _26221_;
wire _26222_;
wire _26223_;
wire _26224_;
wire _26225_;
wire _26226_;
wire _26227_;
wire _26228_;
wire _26229_;
wire _26230_;
wire _26231_;
wire _26232_;
wire _26233_;
wire _26234_;
wire _26235_;
wire _26236_;
wire _26237_;
wire _26238_;
wire _26239_;
wire _26240_;
wire _26241_;
wire _26242_;
wire _26243_;
wire _26244_;
wire _26245_;
wire _26246_;
wire _26247_;
wire _26248_;
wire _26249_;
wire _26250_;
wire _26251_;
wire _26252_;
wire _26253_;
wire _26254_;
wire _26255_;
wire _26256_;
wire _26257_;
wire _26258_;
wire _26259_;
wire _26260_;
wire _26261_;
wire _26262_;
wire _26263_;
wire _26264_;
wire _26265_;
wire _26266_;
wire _26267_;
wire _26268_;
wire _26269_;
wire _26270_;
wire _26271_;
wire _26272_;
wire _26273_;
wire _26274_;
wire _26275_;
wire _26276_;
wire _26277_;
wire _26278_;
wire _26279_;
wire _26280_;
wire _26281_;
wire _26282_;
wire _26283_;
wire _26284_;
wire _26285_;
wire _26286_;
wire _26287_;
wire _26288_;
wire _26289_;
wire _26290_;
wire _26291_;
wire _26292_;
wire _26293_;
wire _26294_;
wire _26295_;
wire _26296_;
wire _26297_;
wire _26298_;
wire _26299_;
wire _26300_;
wire _26301_;
wire _26302_;
wire _26303_;
wire _26304_;
wire _26305_;
wire _26306_;
wire _26307_;
wire _26308_;
wire _26309_;
wire _26310_;
wire _26311_;
wire _26312_;
wire _26313_;
wire _26314_;
wire _26315_;
wire _26316_;
wire _26317_;
wire _26318_;
wire _26319_;
wire _26320_;
wire _26321_;
wire _26322_;
wire _26323_;
wire _26324_;
wire _26325_;
wire _26326_;
wire _26327_;
wire _26328_;
wire _26329_;
wire _26330_;
wire _26331_;
wire _26332_;
wire _26333_;
wire _26334_;
wire _26335_;
wire _26336_;
wire _26337_;
wire _26338_;
wire _26339_;
wire _26340_;
wire _26341_;
wire _26342_;
wire _26343_;
wire _26344_;
wire _26345_;
wire _26346_;
wire _26347_;
wire _26348_;
wire _26349_;
wire _26350_;
wire _26351_;
wire _26352_;
wire _26353_;
wire _26354_;
wire _26355_;
wire _26356_;
wire _26357_;
wire _26358_;
wire _26359_;
wire _26360_;
wire _26361_;
wire _26362_;
wire _26363_;
wire _26364_;
wire _26365_;
wire _26366_;
wire _26367_;
wire _26368_;
wire _26369_;
wire _26370_;
wire _26371_;
wire _26372_;
wire _26373_;
wire _26374_;
wire _26375_;
wire _26376_;
wire _26377_;
wire _26378_;
wire _26379_;
wire _26380_;
wire _26381_;
wire _26382_;
wire _26383_;
wire _26384_;
wire _26385_;
wire _26386_;
wire _26387_;
wire _26388_;
wire _26389_;
wire _26390_;
wire _26391_;
wire _26392_;
wire _26393_;
wire _26394_;
wire _26395_;
wire _26396_;
wire _26397_;
wire _26398_;
wire _26399_;
wire _26400_;
wire _26401_;
wire _26402_;
wire _26403_;
wire _26404_;
wire _26405_;
wire _26406_;
wire _26407_;
wire _26408_;
wire _26409_;
wire _26410_;
wire _26411_;
wire _26412_;
wire _26413_;
wire _26414_;
wire _26415_;
wire _26416_;
wire _26417_;
wire _26418_;
wire _26419_;
wire _26420_;
wire _26421_;
wire _26422_;
wire _26423_;
wire _26424_;
wire _26425_;
wire _26426_;
wire _26427_;
wire _26428_;
wire _26429_;
wire _26430_;
wire _26431_;
wire _26432_;
wire _26433_;
wire _26434_;
wire _26435_;
wire _26436_;
wire _26437_;
wire _26438_;
wire _26439_;
wire _26440_;
wire _26441_;
wire _26442_;
wire _26443_;
wire _26444_;
wire _26445_;
wire _26446_;
wire _26447_;
wire _26448_;
wire _26449_;
wire _26450_;
wire _26451_;
wire _26452_;
wire _26453_;
wire _26454_;
wire _26455_;
wire _26456_;
wire _26457_;
wire _26458_;
wire _26459_;
wire _26460_;
wire _26461_;
wire _26462_;
wire _26463_;
wire _26464_;
wire _26465_;
wire _26466_;
wire _26467_;
wire _26468_;
wire _26469_;
wire _26470_;
wire _26471_;
wire _26472_;
wire _26473_;
wire _26474_;
wire _26475_;
wire _26476_;
wire _26477_;
wire _26478_;
wire _26479_;
wire _26480_;
wire _26481_;
wire _26482_;
wire _26483_;
wire _26484_;
wire _26485_;
wire _26486_;
wire _26487_;
wire _26488_;
wire _26489_;
wire _26490_;
wire _26491_;
wire _26492_;
wire _26493_;
wire _26494_;
wire _26495_;
wire _26496_;
wire _26497_;
wire _26498_;
wire _26499_;
wire _26500_;
wire _26501_;
wire _26502_;
wire _26503_;
wire _26504_;
wire _26505_;
wire _26506_;
wire _26507_;
wire _26508_;
wire _26509_;
wire _26510_;
wire _26511_;
wire _26512_;
wire _26513_;
wire _26514_;
wire _26515_;
wire _26516_;
wire _26517_;
wire _26518_;
wire _26519_;
wire _26520_;
wire _26521_;
wire _26522_;
wire _26523_;
wire _26524_;
wire _26525_;
wire _26526_;
wire _26527_;
wire _26528_;
wire _26529_;
wire _26530_;
wire _26531_;
wire _26532_;
wire _26533_;
wire _26534_;
wire _26535_;
wire _26536_;
wire _26537_;
wire _26538_;
wire _26539_;
wire _26540_;
wire _26541_;
wire _26542_;
wire _26543_;
wire _26544_;
wire _26545_;
wire _26546_;
wire _26547_;
wire _26548_;
wire _26549_;
wire _26550_;
wire _26551_;
wire _26552_;
wire _26553_;
wire _26554_;
wire _26555_;
wire _26556_;
wire _26557_;
wire _26558_;
wire _26559_;
wire _26560_;
wire _26561_;
wire _26562_;
wire _26563_;
wire _26564_;
wire _26565_;
wire _26566_;
wire _26567_;
wire _26568_;
wire _26569_;
wire _26570_;
wire _26571_;
wire _26572_;
wire _26573_;
wire _26574_;
wire _26575_;
wire _26576_;
wire _26577_;
wire _26578_;
wire _26579_;
wire _26580_;
wire _26581_;
wire _26582_;
wire _26583_;
wire _26584_;
wire _26585_;
wire _26586_;
wire _26587_;
wire _26588_;
wire _26589_;
wire _26590_;
wire _26591_;
wire _26592_;
wire _26593_;
wire _26594_;
wire _26595_;
wire _26596_;
wire _26597_;
wire _26598_;
wire _26599_;
wire _26600_;
wire _26601_;
wire _26602_;
wire _26603_;
wire _26604_;
wire _26605_;
wire _26606_;
wire _26607_;
wire _26608_;
wire _26609_;
wire _26610_;
wire _26611_;
wire _26612_;
wire _26613_;
wire _26614_;
wire _26615_;
wire _26616_;
wire _26617_;
wire _26618_;
wire _26619_;
wire _26620_;
wire _26621_;
wire _26622_;
wire _26623_;
wire _26624_;
wire _26625_;
wire _26626_;
wire _26627_;
wire _26628_;
wire _26629_;
wire _26630_;
wire _26631_;
wire _26632_;
wire _26633_;
wire _26634_;
wire _26635_;
wire _26636_;
wire _26637_;
wire _26638_;
wire _26639_;
wire _26640_;
wire _26641_;
wire _26642_;
wire _26643_;
wire _26644_;
wire _26645_;
wire _26646_;
wire _26647_;
wire _26648_;
wire _26649_;
wire _26650_;
wire _26651_;
wire _26652_;
wire _26653_;
wire _26654_;
wire _26655_;
wire _26656_;
wire _26657_;
wire _26658_;
wire _26659_;
wire _26660_;
wire _26661_;
wire _26662_;
wire _26663_;
wire _26664_;
wire _26665_;
wire _26666_;
wire _26667_;
wire _26668_;
wire _26669_;
wire _26670_;
wire _26671_;
wire _26672_;
wire _26673_;
wire _26674_;
wire _26675_;
wire _26676_;
wire _26677_;
wire _26678_;
wire _26679_;
wire _26680_;
wire _26681_;
wire _26682_;
wire _26683_;
wire _26684_;
wire _26685_;
wire _26686_;
wire _26687_;
wire _26688_;
wire _26689_;
wire _26690_;
wire _26691_;
wire _26692_;
wire _26693_;
wire _26694_;
wire _26695_;
wire _26696_;
wire _26697_;
wire _26698_;
wire _26699_;
wire _26700_;
wire _26701_;
wire _26702_;
wire _26703_;
wire _26704_;
wire _26705_;
wire _26706_;
wire _26707_;
wire _26708_;
wire _26709_;
wire _26710_;
wire _26711_;
wire _26712_;
wire _26713_;
wire _26714_;
wire _26715_;
wire _26716_;
wire _26717_;
wire _26718_;
wire _26719_;
wire _26720_;
wire _26721_;
wire _26722_;
wire _26723_;
wire _26724_;
wire _26725_;
wire _26726_;
wire _26727_;
wire _26728_;
wire _26729_;
wire _26730_;
wire _26731_;
wire _26732_;
wire _26733_;
wire _26734_;
wire _26735_;
wire _26736_;
wire _26737_;
wire _26738_;
wire _26739_;
wire _26740_;
wire _26741_;
wire _26742_;
wire _26743_;
wire _26744_;
wire _26745_;
wire _26746_;
wire _26747_;
wire _26748_;
wire _26749_;
wire _26750_;
wire _26751_;
wire _26752_;
wire _26753_;
wire _26754_;
wire _26755_;
wire _26756_;
wire _26757_;
wire _26758_;
wire _26759_;
wire _26760_;
wire _26761_;
wire _26762_;
wire _26763_;
wire _26764_;
wire _26765_;
wire _26766_;
wire _26767_;
wire _26768_;
wire _26769_;
wire _26770_;
wire _26771_;
wire _26772_;
wire _26773_;
wire _26774_;
wire _26775_;
wire _26776_;
wire _26777_;
wire _26778_;
wire _26779_;
wire _26780_;
wire _26781_;
wire _26782_;
wire _26783_;
wire _26784_;
wire _26785_;
wire _26786_;
wire _26787_;
wire _26788_;
wire _26789_;
wire _26790_;
wire _26791_;
wire _26792_;
wire _26793_;
wire _26794_;
wire _26795_;
wire _26796_;
wire _26797_;
wire _26798_;
wire _26799_;
wire _26800_;
wire _26801_;
wire _26802_;
wire _26803_;
wire _26804_;
wire _26805_;
wire _26806_;
wire _26807_;
wire _26808_;
wire _26809_;
wire _26810_;
wire _26811_;
wire _26812_;
wire _26813_;
wire _26814_;
wire _26815_;
wire _26816_;
wire _26817_;
wire _26818_;
wire _26819_;
wire _26820_;
wire _26821_;
wire _26822_;
wire _26823_;
wire _26824_;
wire _26825_;
wire _26826_;
wire _26827_;
wire _26828_;
wire _26829_;
wire _26830_;
wire _26831_;
wire _26832_;
wire _26833_;
wire _26834_;
wire _26835_;
wire _26836_;
wire _26837_;
wire _26838_;
wire _26839_;
wire _26840_;
wire _26841_;
wire _26842_;
wire _26843_;
wire _26844_;
wire _26845_;
wire _26846_;
wire _26847_;
wire _26848_;
wire _26849_;
wire _26850_;
wire _26851_;
wire _26852_;
wire _26853_;
wire _26854_;
wire _26855_;
wire _26856_;
wire _26857_;
wire _26858_;
wire _26859_;
wire _26860_;
wire _26861_;
wire _26862_;
wire _26863_;
wire _26864_;
wire _26865_;
wire _26866_;
wire _26867_;
wire _26868_;
wire _26869_;
wire _26870_;
wire _26871_;
wire _26872_;
wire _26873_;
wire _26874_;
wire _26875_;
wire _26876_;
wire _26877_;
wire _26878_;
wire _26879_;
wire _26880_;
wire _26881_;
wire _26882_;
wire _26883_;
wire _26884_;
wire _26885_;
wire _26886_;
wire _26887_;
wire _26888_;
wire _26889_;
wire _26890_;
wire _26891_;
wire _26892_;
wire _26893_;
wire _26894_;
wire _26895_;
wire _26896_;
wire _26897_;
wire _26898_;
wire _26899_;
wire _26900_;
wire _26901_;
wire _26902_;
wire _26903_;
wire _26904_;
wire _26905_;
wire _26906_;
wire _26907_;
wire _26908_;
wire _26909_;
wire _26910_;
wire _26911_;
wire _26912_;
wire _26913_;
wire _26914_;
wire _26915_;
wire _26916_;
wire _26917_;
wire _26918_;
wire _26919_;
wire _26920_;
wire _26921_;
wire _26922_;
wire _26923_;
wire _26924_;
wire _26925_;
wire _26926_;
wire _26927_;
wire _26928_;
wire _26929_;
wire _26930_;
wire _26931_;
wire _26932_;
wire _26933_;
wire _26934_;
wire _26935_;
wire _26936_;
wire _26937_;
wire _26938_;
wire _26939_;
wire _26940_;
wire _26941_;
wire _26942_;
wire _26943_;
wire _26944_;
wire _26945_;
wire _26946_;
wire _26947_;
wire _26948_;
wire _26949_;
wire _26950_;
wire _26951_;
wire _26952_;
wire _26953_;
wire _26954_;
wire _26955_;
wire _26956_;
wire _26957_;
wire _26958_;
wire _26959_;
wire _26960_;
wire _26961_;
wire _26962_;
wire _26963_;
wire _26964_;
wire _26965_;
wire _26966_;
wire _26967_;
wire _26968_;
wire _26969_;
wire _26970_;
wire _26971_;
wire _26972_;
wire _26973_;
wire _26974_;
wire _26975_;
wire _26976_;
wire _26977_;
wire _26978_;
wire _26979_;
wire _26980_;
wire _26981_;
wire _26982_;
wire _26983_;
wire _26984_;
wire _26985_;
wire _26986_;
wire _26987_;
wire _26988_;
wire _26989_;
wire _26990_;
wire _26991_;
wire _26992_;
wire _26993_;
wire _26994_;
wire _26995_;
wire _26996_;
wire _26997_;
wire _26998_;
wire _26999_;
wire _27000_;
wire _27001_;
wire _27002_;
wire _27003_;
wire _27004_;
wire _27005_;
wire _27006_;
wire _27007_;
wire _27008_;
wire _27009_;
wire _27010_;
wire _27011_;
wire _27012_;
wire _27013_;
wire _27014_;
wire _27015_;
wire _27016_;
wire _27017_;
wire _27018_;
wire _27019_;
wire _27020_;
wire _27021_;
wire _27022_;
wire _27023_;
wire _27024_;
wire _27025_;
wire _27026_;
wire _27027_;
wire _27028_;
wire _27029_;
wire _27030_;
wire _27031_;
wire _27032_;
wire _27033_;
wire _27034_;
wire _27035_;
wire _27036_;
wire _27037_;
wire _27038_;
wire _27039_;
wire _27040_;
wire _27041_;
wire _27042_;
wire _27043_;
wire _27044_;
wire _27045_;
wire _27046_;
wire _27047_;
wire _27048_;
wire _27049_;
wire _27050_;
wire _27051_;
wire _27052_;
wire _27053_;
wire _27054_;
wire _27055_;
wire _27056_;
wire _27057_;
wire _27058_;
wire _27059_;
wire _27060_;
wire _27061_;
wire _27062_;
wire _27063_;
wire _27064_;
wire _27065_;
wire _27066_;
wire _27067_;
wire _27068_;
wire _27069_;
wire _27070_;
wire _27071_;
wire _27072_;
wire _27073_;
wire _27074_;
wire _27075_;
wire _27076_;
wire _27077_;
wire _27078_;
wire _27079_;
wire _27080_;
wire _27081_;
wire _27082_;
wire _27083_;
wire _27084_;
wire _27085_;
wire _27086_;
wire _27087_;
wire _27088_;
wire _27089_;
wire _27090_;
wire _27091_;
wire _27092_;
wire _27093_;
wire _27094_;
wire _27095_;
wire _27096_;
wire _27097_;
wire _27098_;
wire _27099_;
wire _27100_;
wire _27101_;
wire _27102_;
wire _27103_;
wire _27104_;
wire _27105_;
wire _27106_;
wire _27107_;
wire _27108_;
wire _27109_;
wire _27110_;
wire _27111_;
wire _27112_;
wire _27113_;
wire _27114_;
wire _27115_;
wire _27116_;
wire _27117_;
wire _27118_;
wire _27119_;
wire _27120_;
wire _27121_;
wire _27122_;
wire _27123_;
wire _27124_;
wire _27125_;
wire _27126_;
wire _27127_;
wire _27128_;
wire _27129_;
wire _27130_;
wire _27131_;
wire _27132_;
wire _27133_;
wire _27134_;
wire _27135_;
wire _27136_;
wire _27137_;
wire _27138_;
wire _27139_;
wire _27140_;
wire _27141_;
wire _27142_;
wire _27143_;
wire _27144_;
wire _27145_;
wire _27146_;
wire _27147_;
wire _27148_;
wire _27149_;
wire _27150_;
wire _27151_;
wire _27152_;
wire _27153_;
wire _27154_;
wire _27155_;
wire _27156_;
wire _27157_;
wire _27158_;
wire _27159_;
wire _27160_;
wire _27161_;
wire _27162_;
wire _27163_;
wire _27164_;
wire _27165_;
wire _27166_;
wire _27167_;
wire _27168_;
wire _27169_;
wire _27170_;
wire _27171_;
wire _27172_;
wire _27173_;
wire _27174_;
wire _27175_;
wire _27176_;
wire _27177_;
wire _27178_;
wire _27179_;
wire _27180_;
wire _27181_;
wire _27182_;
wire _27183_;
wire _27184_;
wire _27185_;
wire _27186_;
wire _27187_;
wire _27188_;
wire _27189_;
wire _27190_;
wire _27191_;
wire _27192_;
wire _27193_;
wire _27194_;
wire _27195_;
wire _27196_;
wire _27197_;
wire _27198_;
wire _27199_;
wire _27200_;
wire _27201_;
wire _27202_;
wire _27203_;
wire _27204_;
wire _27205_;
wire _27206_;
wire _27207_;
wire _27208_;
wire _27209_;
wire _27210_;
wire _27211_;
wire _27212_;
wire _27213_;
wire _27214_;
wire _27215_;
wire _27216_;
wire _27217_;
wire _27218_;
wire _27219_;
wire _27220_;
wire _27221_;
wire _27222_;
wire _27223_;
wire _27224_;
wire _27225_;
wire _27226_;
wire _27227_;
wire _27228_;
wire _27229_;
wire _27230_;
wire _27231_;
wire _27232_;
wire _27233_;
wire _27234_;
wire _27235_;
wire _27236_;
wire _27237_;
wire _27238_;
wire _27239_;
wire _27240_;
wire _27241_;
wire _27242_;
wire _27243_;
wire _27244_;
wire _27245_;
wire _27246_;
wire _27247_;
wire _27248_;
wire _27249_;
wire _27250_;
wire _27251_;
wire _27252_;
wire _27253_;
wire _27254_;
wire _27255_;
wire _27256_;
wire _27257_;
wire _27258_;
wire _27259_;
wire _27260_;
wire _27261_;
wire _27262_;
wire _27263_;
wire _27264_;
wire _27265_;
wire _27266_;
wire _27267_;
wire _27268_;
wire _27269_;
wire _27270_;
wire _27271_;
wire _27272_;
wire _27273_;
wire _27274_;
wire _27275_;
wire _27276_;
wire _27277_;
wire _27278_;
wire _27279_;
wire _27280_;
wire _27281_;
wire _27282_;
wire _27283_;
wire _27284_;
wire _27285_;
wire _27286_;
wire _27287_;
wire _27288_;
wire _27289_;
wire _27290_;
wire _27291_;
wire _27292_;
wire _27293_;
wire _27294_;
wire _27295_;
wire _27296_;
wire _27297_;
wire _27298_;
wire _27299_;
wire _27300_;
wire _27301_;
wire _27302_;
wire _27303_;
wire _27304_;
wire _27305_;
wire _27306_;
wire _27307_;
wire _27308_;
wire _27309_;
wire _27310_;
wire _27311_;
wire _27312_;
wire _27313_;
wire _27314_;
wire _27315_;
wire _27316_;
wire _27317_;
wire _27318_;
wire _27319_;
wire _27320_;
wire _27321_;
wire _27322_;
wire _27323_;
wire _27324_;
wire _27325_;
wire _27326_;
wire _27327_;
wire _27328_;
wire _27329_;
wire _27330_;
wire _27331_;
wire _27332_;
wire _27333_;
wire _27334_;
wire _27335_;
wire _27336_;
wire _27337_;
wire _27338_;
wire _27339_;
wire _27340_;
wire _27341_;
wire _27342_;
wire _27343_;
wire _27344_;
wire _27345_;
wire _27346_;
wire _27347_;
wire _27348_;
wire _27349_;
wire _27350_;
wire _27351_;
wire _27352_;
wire _27353_;
wire _27354_;
wire _27355_;
wire _27356_;
wire _27357_;
wire _27358_;
wire _27359_;
wire _27360_;
wire _27361_;
wire _27362_;
wire _27363_;
wire _27364_;
wire _27365_;
wire _27366_;
wire _27367_;
wire _27368_;
wire _27369_;
wire _27370_;
wire _27371_;
wire _27372_;
wire _27373_;
wire _27374_;
wire _27375_;
wire _27376_;
wire _27377_;
wire _27378_;
wire _27379_;
wire _27380_;
wire _27381_;
wire _27382_;
wire _27383_;
wire _27384_;
wire _27385_;
wire _27386_;
wire _27387_;
wire _27388_;
wire _27389_;
wire _27390_;
wire _27391_;
wire _27392_;
wire _27393_;
wire _27394_;
wire _27395_;
wire _27396_;
wire _27397_;
wire _27398_;
wire _27399_;
wire _27400_;
wire _27401_;
wire _27402_;
wire _27403_;
wire _27404_;
wire _27405_;
wire _27406_;
wire _27407_;
wire _27408_;
wire _27409_;
wire _27410_;
wire _27411_;
wire _27412_;
wire _27413_;
wire _27414_;
wire _27415_;
wire _27416_;
wire _27417_;
wire _27418_;
wire _27419_;
wire _27420_;
wire _27421_;
wire _27422_;
wire _27423_;
wire _27424_;
wire _27425_;
wire _27426_;
wire _27427_;
wire _27428_;
wire _27429_;
wire _27430_;
wire _27431_;
wire _27432_;
wire _27433_;
wire _27434_;
wire _27435_;
wire _27436_;
wire _27437_;
wire _27438_;
wire _27439_;
wire _27440_;
wire _27441_;
wire _27442_;
wire _27443_;
wire _27444_;
wire _27445_;
wire _27446_;
wire _27447_;
wire _27448_;
wire _27449_;
wire _27450_;
wire _27451_;
wire _27452_;
wire _27453_;
wire _27454_;
wire _27455_;
wire _27456_;
wire _27457_;
wire _27458_;
wire _27459_;
wire _27460_;
wire _27461_;
wire _27462_;
wire _27463_;
wire _27464_;
wire _27465_;
wire _27466_;
wire _27467_;
wire _27468_;
wire _27469_;
wire _27470_;
wire _27471_;
wire _27472_;
wire _27473_;
wire _27474_;
wire _27475_;
wire _27476_;
wire _27477_;
wire _27478_;
wire _27479_;
wire _27480_;
wire _27481_;
wire _27482_;
wire _27483_;
wire _27484_;
wire _27485_;
wire _27486_;
wire _27487_;
wire _27488_;
wire _27489_;
wire _27490_;
wire _27491_;
wire _27492_;
wire _27493_;
wire _27494_;
wire _27495_;
wire _27496_;
wire _27497_;
wire _27498_;
wire _27499_;
wire _27500_;
wire _27501_;
wire _27502_;
wire _27503_;
wire _27504_;
wire _27505_;
wire _27506_;
wire _27507_;
wire _27508_;
wire _27509_;
wire _27510_;
wire _27511_;
wire _27512_;
wire _27513_;
wire _27514_;
wire _27515_;
wire _27516_;
wire _27517_;
wire _27518_;
wire _27519_;
wire _27520_;
wire _27521_;
wire _27522_;
wire _27523_;
wire _27524_;
wire _27525_;
wire _27526_;
wire _27527_;
wire _27528_;
wire _27529_;
wire _27530_;
wire _27531_;
wire _27532_;
wire _27533_;
wire _27534_;
wire _27535_;
wire _27536_;
wire _27537_;
wire _27538_;
wire _27539_;
wire _27540_;
wire _27541_;
wire _27542_;
wire _27543_;
wire _27544_;
wire _27545_;
wire _27546_;
wire _27547_;
wire _27548_;
wire _27549_;
wire _27550_;
wire _27551_;
wire _27552_;
wire _27553_;
wire _27554_;
wire _27555_;
wire _27556_;
wire _27557_;
wire _27558_;
wire _27559_;
wire _27560_;
wire _27561_;
wire _27562_;
wire _27563_;
wire _27564_;
wire _27565_;
wire _27566_;
wire _27567_;
wire _27568_;
wire _27569_;
wire _27570_;
wire _27571_;
wire _27572_;
wire _27573_;
wire _27574_;
wire _27575_;
wire _27576_;
wire _27577_;
wire _27578_;
wire _27579_;
wire _27580_;
wire _27581_;
wire _27582_;
wire _27583_;
wire _27584_;
wire _27585_;
wire _27586_;
wire _27587_;
wire _27588_;
wire _27589_;
wire _27590_;
wire _27591_;
wire _27592_;
wire _27593_;
wire _27594_;
wire _27595_;
wire _27596_;
wire _27597_;
wire _27598_;
wire _27599_;
wire _27600_;
wire _27601_;
wire _27602_;
wire _27603_;
wire _27604_;
wire _27605_;
wire _27606_;
wire _27607_;
wire _27608_;
wire _27609_;
wire _27610_;
wire _27611_;
wire _27612_;
wire _27613_;
wire _27614_;
wire _27615_;
wire _27616_;
wire _27617_;
wire _27618_;
wire _27619_;
wire _27620_;
wire _27621_;
wire _27622_;
wire _27623_;
wire _27624_;
wire _27625_;
wire _27626_;
wire _27627_;
wire _27628_;
wire _27629_;
wire _27630_;
wire _27631_;
wire _27632_;
wire _27633_;
wire _27634_;
wire _27635_;
wire _27636_;
wire _27637_;
wire _27638_;
wire _27639_;
wire _27640_;
wire _27641_;
wire _27642_;
wire _27643_;
wire _27644_;
wire _27645_;
wire _27646_;
wire _27647_;
wire _27648_;
wire _27649_;
wire _27650_;
wire _27651_;
wire _27652_;
wire _27653_;
wire _27654_;
wire _27655_;
wire _27656_;
wire _27657_;
wire _27658_;
wire _27659_;
wire _27660_;
wire _27661_;
wire _27662_;
wire _27663_;
wire _27664_;
wire _27665_;
wire _27666_;
wire _27667_;
wire _27668_;
wire _27669_;
wire _27670_;
wire _27671_;
wire _27672_;
wire _27673_;
wire _27674_;
wire _27675_;
wire _27676_;
wire _27677_;
wire _27678_;
wire _27679_;
wire _27680_;
wire _27681_;
wire _27682_;
wire _27683_;
wire _27684_;
wire _27685_;
wire _27686_;
wire _27687_;
wire _27688_;
wire _27689_;
wire _27690_;
wire _27691_;
wire _27692_;
wire _27693_;
wire _27694_;
wire _27695_;
wire _27696_;
wire _27697_;
wire _27698_;
wire _27699_;
wire _27700_;
wire _27701_;
wire _27702_;
wire _27703_;
wire _27704_;
wire _27705_;
wire _27706_;
wire _27707_;
wire _27708_;
wire _27709_;
wire _27710_;
wire _27711_;
wire _27712_;
wire _27713_;
wire _27714_;
wire _27715_;
wire _27716_;
wire _27717_;
wire _27718_;
wire _27719_;
wire _27720_;
wire _27721_;
wire _27722_;
wire _27723_;
wire _27724_;
wire _27725_;
wire _27726_;
wire _27727_;
wire _27728_;
wire _27729_;
wire _27730_;
wire _27731_;
wire _27732_;
wire _27733_;
wire _27734_;
wire _27735_;
wire _27736_;
wire _27737_;
wire _27738_;
wire _27739_;
wire _27740_;
wire _27741_;
wire _27742_;
wire _27743_;
wire _27744_;
wire _27745_;
wire _27746_;
wire _27747_;
wire _27748_;
wire _27749_;
wire _27750_;
wire _27751_;
wire _27752_;
wire _27753_;
wire _27754_;
wire _27755_;
wire _27756_;
wire _27757_;
wire _27758_;
wire _27759_;
wire _27760_;
wire _27761_;
wire _27762_;
wire _27763_;
wire _27764_;
wire _27765_;
wire _27766_;
wire _27767_;
wire _27768_;
wire _27769_;
wire _27770_;
wire _27771_;
wire _27772_;
wire _27773_;
wire _27774_;
wire _27775_;
wire _27776_;
wire _27777_;
wire _27778_;
wire _27779_;
wire _27780_;
wire _27781_;
wire _27782_;
wire _27783_;
wire _27784_;
wire _27785_;
wire _27786_;
wire _27787_;
wire _27788_;
wire _27789_;
wire _27790_;
wire _27791_;
wire _27792_;
wire _27793_;
wire _27794_;
wire _27795_;
wire _27796_;
wire _27797_;
wire _27798_;
wire _27799_;
wire _27800_;
wire _27801_;
wire _27802_;
wire _27803_;
wire _27804_;
wire _27805_;
wire _27806_;
wire _27807_;
wire _27808_;
wire _27809_;
wire _27810_;
wire _27811_;
wire _27812_;
wire _27813_;
wire _27814_;
wire _27815_;
wire _27816_;
wire _27817_;
wire _27818_;
wire _27819_;
wire _27820_;
wire _27821_;
wire _27822_;
wire _27823_;
wire _27824_;
wire _27825_;
wire _27826_;
wire _27827_;
wire _27828_;
wire _27829_;
wire _27830_;
wire _27831_;
wire _27832_;
wire _27833_;
wire _27834_;
wire _27835_;
wire _27836_;
wire _27837_;
wire _27838_;
wire _27839_;
wire _27840_;
wire _27841_;
wire _27842_;
wire _27843_;
wire _27844_;
wire _27845_;
wire _27846_;
wire _27847_;
wire _27848_;
wire _27849_;
wire _27850_;
wire _27851_;
wire _27852_;
wire _27853_;
wire _27854_;
wire _27855_;
wire _27856_;
wire _27857_;
wire _27858_;
wire _27859_;
wire _27860_;
wire _27861_;
wire _27862_;
wire _27863_;
wire _27864_;
wire _27865_;
wire _27866_;
wire _27867_;
wire _27868_;
wire _27869_;
wire _27870_;
wire _27871_;
wire _27872_;
wire _27873_;
wire _27874_;
wire _27875_;
wire _27876_;
wire _27877_;
wire _27878_;
wire _27879_;
wire _27880_;
wire _27881_;
wire _27882_;
wire _27883_;
wire _27884_;
wire _27885_;
wire _27886_;
wire _27887_;
wire _27888_;
wire _27889_;
wire _27890_;
wire _27891_;
wire _27892_;
wire _27893_;
wire _27894_;
wire _27895_;
wire _27896_;
wire _27897_;
wire _27898_;
wire _27899_;
wire _27900_;
wire _27901_;
wire _27902_;
wire _27903_;
wire _27904_;
wire _27905_;
wire _27906_;
wire _27907_;
wire _27908_;
wire _27909_;
wire _27910_;
wire _27911_;
wire _27912_;
wire _27913_;
wire _27914_;
wire _27915_;
wire _27916_;
wire _27917_;
wire _27918_;
wire _27919_;
wire _27920_;
wire _27921_;
wire _27922_;
wire _27923_;
wire _27924_;
wire _27925_;
wire _27926_;
wire _27927_;
wire _27928_;
wire _27929_;
wire _27930_;
wire _27931_;
wire _27932_;
wire _27933_;
wire _27934_;
wire _27935_;
wire _27936_;
wire _27937_;
wire _27938_;
wire _27939_;
wire _27940_;
wire _27941_;
wire _27942_;
wire _27943_;
wire _27944_;
wire _27945_;
wire _27946_;
wire _27947_;
wire _27948_;
wire _27949_;
wire _27950_;
wire _27951_;
wire _27952_;
wire _27953_;
wire _27954_;
wire _27955_;
wire _27956_;
wire _27957_;
wire _27958_;
wire _27959_;
wire _27960_;
wire _27961_;
wire _27962_;
wire _27963_;
wire _27964_;
wire _27965_;
wire _27966_;
wire _27967_;
wire _27968_;
wire _27969_;
wire _27970_;
wire _27971_;
wire _27972_;
wire _27973_;
wire _27974_;
wire _27975_;
wire _27976_;
wire _27977_;
wire _27978_;
wire _27979_;
wire _27980_;
wire _27981_;
wire _27982_;
wire _27983_;
wire _27984_;
wire _27985_;
wire _27986_;
wire _27987_;
wire _27988_;
wire _27989_;
wire _27990_;
wire _27991_;
wire _27992_;
wire _27993_;
wire _27994_;
wire _27995_;
wire _27996_;
wire _27997_;
wire _27998_;
wire _27999_;
wire _28000_;
wire _28001_;
wire _28002_;
wire _28003_;
wire _28004_;
wire _28005_;
wire _28006_;
wire _28007_;
wire _28008_;
wire _28009_;
wire _28010_;
wire _28011_;
wire _28012_;
wire _28013_;
wire _28014_;
wire _28015_;
wire _28016_;
wire _28017_;
wire _28018_;
wire _28019_;
wire _28020_;
wire _28021_;
wire _28022_;
wire _28023_;
wire _28024_;
wire _28025_;
wire _28026_;
wire _28027_;
wire _28028_;
wire _28029_;
wire _28030_;
wire _28031_;
wire _28032_;
wire _28033_;
wire _28034_;
wire _28035_;
wire _28036_;
wire _28037_;
wire _28038_;
wire _28039_;
wire _28040_;
wire _28041_;
wire _28042_;
wire _28043_;
wire _28044_;
wire _28045_;
wire _28046_;
wire _28047_;
wire _28048_;
wire _28049_;
wire _28050_;
wire _28051_;
wire _28052_;
wire _28053_;
wire _28054_;
wire _28055_;
wire _28056_;
wire _28057_;
wire _28058_;
wire _28059_;
wire _28060_;
wire _28061_;
wire _28062_;
wire _28063_;
wire _28064_;
wire _28065_;
wire _28066_;
wire _28067_;
wire _28068_;
wire _28069_;
wire _28070_;
wire _28071_;
wire _28072_;
wire _28073_;
wire _28074_;
wire _28075_;
wire _28076_;
wire _28077_;
wire _28078_;
wire _28079_;
wire _28080_;
wire _28081_;
wire _28082_;
wire _28083_;
wire _28084_;
wire _28085_;
wire _28086_;
wire _28087_;
wire _28088_;
wire _28089_;
wire _28090_;
wire _28091_;
wire _28092_;
wire _28093_;
wire _28094_;
wire _28095_;
wire _28096_;
wire _28097_;
wire _28098_;
wire _28099_;
wire _28100_;
wire _28101_;
wire _28102_;
wire _28103_;
wire _28104_;
wire _28105_;
wire _28106_;
wire _28107_;
wire _28108_;
wire _28109_;
wire _28110_;
wire _28111_;
wire _28112_;
wire _28113_;
wire _28114_;
wire _28115_;
wire _28116_;
wire _28117_;
wire _28118_;
wire _28119_;
wire _28120_;
wire _28121_;
wire _28122_;
wire _28123_;
wire _28124_;
wire _28125_;
wire _28126_;
wire _28127_;
wire _28128_;
wire _28129_;
wire _28130_;
wire _28131_;
wire _28132_;
wire _28133_;
wire _28134_;
wire _28135_;
wire _28136_;
wire _28137_;
wire _28138_;
wire _28139_;
wire _28140_;
wire _28141_;
wire _28142_;
wire _28143_;
wire _28144_;
wire _28145_;
wire _28146_;
wire _28147_;
wire _28148_;
wire _28149_;
wire _28150_;
wire _28151_;
wire _28152_;
wire _28153_;
wire _28154_;
wire _28155_;
wire _28156_;
wire _28157_;
wire _28158_;
wire _28159_;
wire _28160_;
wire _28161_;
wire _28162_;
wire _28163_;
wire _28164_;
wire _28165_;
wire _28166_;
wire _28167_;
wire _28168_;
wire _28169_;
wire _28170_;
wire _28171_;
wire _28172_;
wire _28173_;
wire _28174_;
wire _28175_;
wire _28176_;
wire _28177_;
wire _28178_;
wire _28179_;
wire _28180_;
wire _28181_;
wire _28182_;
wire _28183_;
wire _28184_;
wire _28185_;
wire _28186_;
wire _28187_;
wire _28188_;
wire _28189_;
wire _28190_;
wire _28191_;
wire _28192_;
wire _28193_;
wire _28194_;
wire _28195_;
wire _28196_;
wire _28197_;
wire _28198_;
wire _28199_;
wire _28200_;
wire _28201_;
wire _28202_;
wire _28203_;
wire _28204_;
wire _28205_;
wire _28206_;
wire _28207_;
wire _28208_;
wire _28209_;
wire _28210_;
wire _28211_;
wire _28212_;
wire _28213_;
wire _28214_;
wire _28215_;
wire _28216_;
wire _28217_;
wire _28218_;
wire _28219_;
wire _28220_;
wire _28221_;
wire _28222_;
wire _28223_;
wire _28224_;
wire _28225_;
wire _28226_;
wire _28227_;
wire _28228_;
wire _28229_;
wire _28230_;
wire _28231_;
wire _28232_;
wire _28233_;
wire _28234_;
wire _28235_;
wire _28236_;
wire _28237_;
wire _28238_;
wire _28239_;
wire _28240_;
wire _28241_;
wire _28242_;
wire _28243_;
wire _28244_;
wire _28245_;
wire _28246_;
wire _28247_;
wire _28248_;
wire _28249_;
wire _28250_;
wire _28251_;
wire _28252_;
wire _28253_;
wire _28254_;
wire _28255_;
wire _28256_;
wire _28257_;
wire _28258_;
wire _28259_;
wire _28260_;
wire _28261_;
wire _28262_;
wire _28263_;
wire _28264_;
wire _28265_;
wire _28266_;
wire _28267_;
wire _28268_;
wire _28269_;
wire _28270_;
wire _28271_;
wire _28272_;
wire _28273_;
wire _28274_;
wire _28275_;
wire _28276_;
wire _28277_;
wire _28278_;
wire _28279_;
wire _28280_;
wire _28281_;
wire _28282_;
wire _28283_;
wire _28284_;
wire _28285_;
wire _28286_;
wire _28287_;
wire _28288_;
wire _28289_;
wire _28290_;
wire _28291_;
wire _28292_;
wire _28293_;
wire _28294_;
wire _28295_;
wire _28296_;
wire _28297_;
wire _28298_;
wire _28299_;
wire _28300_;
wire _28301_;
wire _28302_;
wire _28303_;
wire _28304_;
wire _28305_;
wire _28306_;
wire _28307_;
wire _28308_;
wire _28309_;
wire _28310_;
wire _28311_;
wire _28312_;
wire _28313_;
wire _28314_;
wire _28315_;
wire _28316_;
wire _28317_;
wire _28318_;
wire _28319_;
wire _28320_;
wire _28321_;
wire _28322_;
wire _28323_;
wire _28324_;
wire _28325_;
wire _28326_;
wire _28327_;
wire _28328_;
wire _28329_;
wire _28330_;
wire _28331_;
wire _28332_;
wire _28333_;
wire _28334_;
wire _28335_;
wire _28336_;
wire _28337_;
wire _28338_;
wire _28339_;
wire _28340_;
wire _28341_;
wire _28342_;
wire _28343_;
wire _28344_;
wire _28345_;
wire _28346_;
wire _28347_;
wire _28348_;
wire _28349_;
wire _28350_;
wire _28351_;
wire _28352_;
wire _28353_;
wire _28354_;
wire _28355_;
wire _28356_;
wire _28357_;
wire _28358_;
wire _28359_;
wire _28360_;
wire _28361_;
wire _28362_;
wire _28363_;
wire _28364_;
wire _28365_;
wire _28366_;
wire _28367_;
wire _28368_;
wire _28369_;
wire _28370_;
wire _28371_;
wire _28372_;
wire _28373_;
wire _28374_;
wire _28375_;
wire _28376_;
wire _28377_;
wire _28378_;
wire _28379_;
wire _28380_;
wire _28381_;
wire _28382_;
wire _28383_;
wire _28384_;
wire _28385_;
wire _28386_;
wire _28387_;
wire _28388_;
wire _28389_;
wire _28390_;
wire _28391_;
wire _28392_;
wire _28393_;
wire _28394_;
wire _28395_;
wire _28396_;
wire _28397_;
wire _28398_;
wire _28399_;
wire _28400_;
wire _28401_;
wire _28402_;
wire _28403_;
wire _28404_;
wire _28405_;
wire _28406_;
wire _28407_;
wire _28408_;
wire _28409_;
wire _28410_;
wire _28411_;
wire _28412_;
wire _28413_;
wire _28414_;
wire _28415_;
wire _28416_;
wire _28417_;
wire _28418_;
wire _28419_;
wire _28420_;
wire _28421_;
wire _28422_;
wire _28423_;
wire _28424_;
wire _28425_;
wire _28426_;
wire _28427_;
wire _28428_;
wire _28429_;
wire _28430_;
wire _28431_;
wire _28432_;
wire _28433_;
wire _28434_;
wire _28435_;
wire _28436_;
wire _28437_;
wire _28438_;
wire _28439_;
wire _28440_;
wire _28441_;
wire _28442_;
wire _28443_;
wire _28444_;
wire _28445_;
wire _28446_;
wire _28447_;
wire _28448_;
wire _28449_;
wire _28450_;
wire _28451_;
wire _28452_;
wire _28453_;
wire _28454_;
wire _28455_;
wire _28456_;
wire _28457_;
wire _28458_;
wire _28459_;
wire _28460_;
wire _28461_;
wire _28462_;
wire _28463_;
wire _28464_;
wire _28465_;
wire _28466_;
wire _28467_;
wire _28468_;
wire _28469_;
wire _28470_;
wire _28471_;
wire _28472_;
wire _28473_;
wire _28474_;
wire _28475_;
wire _28476_;
wire _28477_;
wire _28478_;
wire _28479_;
wire _28480_;
wire _28481_;
wire _28482_;
wire _28483_;
wire _28484_;
wire _28485_;
wire _28486_;
wire _28487_;
wire _28488_;
wire _28489_;
wire _28490_;
wire _28491_;
wire _28492_;
wire _28493_;
wire _28494_;
wire _28495_;
wire _28496_;
wire _28497_;
wire _28498_;
wire _28499_;
wire _28500_;
wire _28501_;
wire _28502_;
wire _28503_;
wire _28504_;
wire _28505_;
wire _28506_;
wire _28507_;
wire _28508_;
wire _28509_;
wire _28510_;
wire _28511_;
wire _28512_;
wire _28513_;
wire _28514_;
wire _28515_;
wire _28516_;
wire _28517_;
wire _28518_;
wire _28519_;
wire _28520_;
wire _28521_;
wire _28522_;
wire _28523_;
wire _28524_;
wire _28525_;
wire _28526_;
wire _28527_;
wire _28528_;
wire _28529_;
wire _28530_;
wire _28531_;
wire _28532_;
wire _28533_;
wire _28534_;
wire _28535_;
wire _28536_;
wire _28537_;
wire _28538_;
wire _28539_;
wire _28540_;
wire _28541_;
wire _28542_;
wire _28543_;
wire _28544_;
wire _28545_;
wire _28546_;
wire _28547_;
wire _28548_;
wire _28549_;
wire _28550_;
wire _28551_;
wire _28552_;
wire _28553_;
wire _28554_;
wire _28555_;
wire _28556_;
wire _28557_;
wire _28558_;
wire _28559_;
wire _28560_;
wire _28561_;
wire _28562_;
wire _28563_;
wire _28564_;
wire _28565_;
wire _28566_;
wire _28567_;
wire _28568_;
wire _28569_;
wire _28570_;
wire _28571_;
wire _28572_;
wire _28573_;
wire _28574_;
wire _28575_;
wire _28576_;
wire _28577_;
wire _28578_;
wire _28579_;
wire _28580_;
wire _28581_;
wire _28582_;
wire _28583_;
wire _28584_;
wire _28585_;
wire _28586_;
wire _28587_;
wire _28588_;
wire _28589_;
wire _28590_;
wire _28591_;
wire _28592_;
wire _28593_;
wire _28594_;
wire _28595_;
wire _28596_;
wire _28597_;
wire _28598_;
wire _28599_;
wire _28600_;
wire _28601_;
wire _28602_;
wire _28603_;
wire _28604_;
wire _28605_;
wire _28606_;
wire _28607_;
wire _28608_;
wire _28609_;
wire _28610_;
wire _28611_;
wire _28612_;
wire _28613_;
wire _28614_;
wire _28615_;
wire _28616_;
wire _28617_;
wire _28618_;
wire _28619_;
wire _28620_;
wire _28621_;
wire _28622_;
wire _28623_;
wire _28624_;
wire _28625_;
wire _28626_;
wire _28627_;
wire _28628_;
wire _28629_;
wire _28630_;
wire _28631_;
wire _28632_;
wire _28633_;
wire _28634_;
wire _28635_;
wire _28636_;
wire _28637_;
wire _28638_;
wire _28639_;
wire _28640_;
wire _28641_;
wire _28642_;
wire _28643_;
wire _28644_;
wire _28645_;
wire _28646_;
wire _28647_;
wire _28648_;
wire _28649_;
wire _28650_;
wire _28651_;
wire _28652_;
wire _28653_;
wire _28654_;
wire _28655_;
wire _28656_;
wire _28657_;
wire _28658_;
wire _28659_;
wire _28660_;
wire _28661_;
wire _28662_;
wire _28663_;
wire _28664_;
wire _28665_;
wire _28666_;
wire _28667_;
wire _28668_;
wire _28669_;
wire _28670_;
wire _28671_;
wire _28672_;
wire _28673_;
wire _28674_;
wire _28675_;
wire _28676_;
wire _28677_;
wire _28678_;
wire _28679_;
wire _28680_;
wire _28681_;
wire _28682_;
wire _28683_;
wire _28684_;
wire _28685_;
wire _28686_;
wire _28687_;
wire _28688_;
wire _28689_;
wire _28690_;
wire _28691_;
wire _28692_;
wire _28693_;
wire _28694_;
wire _28695_;
wire _28696_;
wire _28697_;
wire _28698_;
wire _28699_;
wire _28700_;
wire _28701_;
wire _28702_;
wire _28703_;
wire _28704_;
wire _28705_;
wire _28706_;
wire _28707_;
wire _28708_;
wire _28709_;
wire _28710_;
wire _28711_;
wire _28712_;
wire _28713_;
wire _28714_;
wire _28715_;
wire _28716_;
wire _28717_;
wire _28718_;
wire _28719_;
wire _28720_;
wire _28721_;
wire _28722_;
wire _28723_;
wire _28724_;
wire _28725_;
wire _28726_;
wire _28727_;
wire _28728_;
wire _28729_;
wire _28730_;
wire _28731_;
wire _28732_;
wire _28733_;
wire _28734_;
wire _28735_;
wire _28736_;
wire _28737_;
wire _28738_;
wire _28739_;
wire _28740_;
wire _28741_;
wire _28742_;
wire _28743_;
wire _28744_;
wire _28745_;
wire _28746_;
wire _28747_;
wire _28748_;
wire _28749_;
wire _28750_;
wire _28751_;
wire _28752_;
wire _28753_;
wire _28754_;
wire _28755_;
wire _28756_;
wire _28757_;
wire _28758_;
wire _28759_;
wire _28760_;
wire _28761_;
wire _28762_;
wire _28763_;
wire _28764_;
wire _28765_;
wire _28766_;
wire _28767_;
wire _28768_;
wire _28769_;
wire _28770_;
wire _28771_;
wire _28772_;
wire _28773_;
wire _28774_;
wire _28775_;
wire _28776_;
wire _28777_;
wire _28778_;
wire _28779_;
wire _28780_;
wire _28781_;
wire _28782_;
wire _28783_;
wire _28784_;
wire _28785_;
wire _28786_;
wire _28787_;
wire _28788_;
wire _28789_;
wire _28790_;
wire _28791_;
wire _28792_;
wire _28793_;
wire _28794_;
wire _28795_;
wire _28796_;
wire _28797_;
wire _28798_;
wire _28799_;
wire _28800_;
wire _28801_;
wire _28802_;
wire _28803_;
wire _28804_;
wire _28805_;
wire _28806_;
wire _28807_;
wire _28808_;
wire _28809_;
wire _28810_;
wire _28811_;
wire _28812_;
wire _28813_;
wire _28814_;
wire _28815_;
wire _28816_;
wire _28817_;
wire _28818_;
wire _28819_;
wire _28820_;
wire _28821_;
wire _28822_;
wire _28823_;
wire _28824_;
wire _28825_;
wire _28826_;
wire _28827_;
wire _28828_;
wire _28829_;
wire _28830_;
wire _28831_;
wire _28832_;
wire _28833_;
wire _28834_;
wire _28835_;
wire _28836_;
wire _28837_;
wire _28838_;
wire _28839_;
wire _28840_;
wire _28841_;
wire _28842_;
wire _28843_;
wire _28844_;
wire _28845_;
wire _28846_;
wire _28847_;
wire _28848_;
wire _28849_;
wire _28850_;
wire _28851_;
wire _28852_;
wire _28853_;
wire _28854_;
wire _28855_;
wire _28856_;
wire _28857_;
wire _28858_;
wire _28859_;
wire _28860_;
wire _28861_;
wire _28862_;
wire _28863_;
wire _28864_;
wire _28865_;
wire _28866_;
wire _28867_;
wire _28868_;
wire _28869_;
wire _28870_;
wire _28871_;
wire _28872_;
wire _28873_;
wire _28874_;
wire _28875_;
wire _28876_;
wire _28877_;
wire _28878_;
wire _28879_;
wire _28880_;
wire _28881_;
wire _28882_;
wire _28883_;
wire _28884_;
wire _28885_;
wire _28886_;
wire _28887_;
wire _28888_;
wire _28889_;
wire _28890_;
wire _28891_;
wire _28892_;
wire _28893_;
wire _28894_;
wire _28895_;
wire _28896_;
wire _28897_;
wire _28898_;
wire _28899_;
wire _28900_;
wire _28901_;
wire _28902_;
wire _28903_;
wire _28904_;
wire _28905_;
wire _28906_;
wire _28907_;
wire _28908_;
wire _28909_;
wire _28910_;
wire _28911_;
wire _28912_;
wire _28913_;
wire _28914_;
wire _28915_;
wire _28916_;
wire _28917_;
wire _28918_;
wire _28919_;
wire _28920_;
wire _28921_;
wire _28922_;
wire _28923_;
wire _28924_;
wire _28925_;
wire _28926_;
wire _28927_;
wire _28928_;
wire _28929_;
wire _28930_;
wire _28931_;
wire _28932_;
wire _28933_;
wire _28934_;
wire _28935_;
wire _28936_;
wire _28937_;
wire _28938_;
wire _28939_;
wire _28940_;
wire _28941_;
wire _28942_;
wire _28943_;
wire _28944_;
wire _28945_;
wire _28946_;
wire _28947_;
wire _28948_;
wire _28949_;
wire _28950_;
wire _28951_;
wire _28952_;
wire _28953_;
wire _28954_;
wire _28955_;
wire _28956_;
wire _28957_;
wire _28958_;
wire _28959_;
wire _28960_;
wire _28961_;
wire _28962_;
wire _28963_;
wire _28964_;
wire _28965_;
wire _28966_;
wire _28967_;
wire _28968_;
wire _28969_;
wire _28970_;
wire _28971_;
wire _28972_;
wire _28973_;
wire _28974_;
wire _28975_;
wire _28976_;
wire _28977_;
wire _28978_;
wire _28979_;
wire _28980_;
wire _28981_;
wire _28982_;
wire _28983_;
wire _28984_;
wire _28985_;
wire _28986_;
wire _28987_;
wire _28988_;
wire _28989_;
wire _28990_;
wire _28991_;
wire _28992_;
wire _28993_;
wire _28994_;
wire _28995_;
wire _28996_;
wire _28997_;
wire _28998_;
wire _28999_;
wire _29000_;
wire _29001_;
wire _29002_;
wire _29003_;
wire _29004_;
wire _29005_;
wire _29006_;
wire _29007_;
wire _29008_;
wire _29009_;
wire _29010_;
wire _29011_;
wire _29012_;
wire _29013_;
wire _29014_;
wire _29015_;
wire _29016_;
wire _29017_;
wire _29018_;
wire _29019_;
wire _29020_;
wire _29021_;
wire _29022_;
wire _29023_;
wire _29024_;
wire _29025_;
wire _29026_;
wire _29027_;
wire _29028_;
wire _29029_;
wire _29030_;
wire _29031_;
wire _29032_;
wire _29033_;
wire _29034_;
wire _29035_;
wire _29036_;
wire _29037_;
wire _29038_;
wire _29039_;
wire _29040_;
wire _29041_;
wire _29042_;
wire _29043_;
wire _29044_;
wire _29045_;
wire _29046_;
wire _29047_;
wire _29048_;
wire _29049_;
wire _29050_;
wire _29051_;
wire _29052_;
wire _29053_;
wire _29054_;
wire _29055_;
wire _29056_;
wire _29057_;
wire _29058_;
wire _29059_;
wire _29060_;
wire _29061_;
wire _29062_;
wire _29063_;
wire _29064_;
wire _29065_;
wire _29066_;
wire _29067_;
wire _29068_;
wire _29069_;
wire _29070_;
wire _29071_;
wire _29072_;
wire _29073_;
wire _29074_;
wire _29075_;
wire _29076_;
wire _29077_;
wire _29078_;
wire _29079_;
wire _29080_;
wire _29081_;
wire _29082_;
wire _29083_;
wire _29084_;
wire _29085_;
wire _29086_;
wire _29087_;
wire _29088_;
wire _29089_;
wire _29090_;
wire _29091_;
wire _29092_;
wire _29093_;
wire _29094_;
wire _29095_;
wire _29096_;
wire _29097_;
wire _29098_;
wire _29099_;
wire _29100_;
wire _29101_;
wire _29102_;
wire _29103_;
wire _29104_;
wire _29105_;
wire _29106_;
wire _29107_;
wire _29108_;
wire _29109_;
wire _29110_;
wire _29111_;
wire _29112_;
wire _29113_;
wire _29114_;
wire _29115_;
wire _29116_;
wire _29117_;
wire _29118_;
wire _29119_;
wire _29120_;
wire _29121_;
wire _29122_;
wire _29123_;
wire _29124_;
wire _29125_;
wire _29126_;
wire _29127_;
wire _29128_;
wire _29129_;
wire _29130_;
wire _29131_;
wire _29132_;
wire _29133_;
wire _29134_;
wire _29135_;
wire _29136_;
wire _29137_;
wire _29138_;
wire _29139_;
wire _29140_;
wire _29141_;
wire _29142_;
wire _29143_;
wire _29144_;
wire _29145_;
wire _29146_;
wire _29147_;
wire _29148_;
wire _29149_;
wire _29150_;
wire _29151_;
wire _29152_;
wire _29153_;
wire _29154_;
wire _29155_;
wire _29156_;
wire _29157_;
wire _29158_;
wire _29159_;
wire _29160_;
wire _29161_;
wire _29162_;
wire _29163_;
wire _29164_;
wire _29165_;
wire _29166_;
wire _29167_;
wire _29168_;
wire _29169_;
wire _29170_;
wire _29171_;
wire _29172_;
wire _29173_;
wire _29174_;
wire _29175_;
wire _29176_;
wire _29177_;
wire _29178_;
wire _29179_;
wire _29180_;
wire _29181_;
wire _29182_;
wire _29183_;
wire _29184_;
wire _29185_;
wire _29186_;
wire _29187_;
wire _29188_;
wire _29189_;
wire _29190_;
wire _29191_;
wire _29192_;
wire _29193_;
wire _29194_;
wire _29195_;
wire _29196_;
wire _29197_;
wire _29198_;
wire _29199_;
wire _29200_;
wire _29201_;
wire _29202_;
wire _29203_;
wire _29204_;
wire _29205_;
wire _29206_;
wire _29207_;
wire _29208_;
wire _29209_;
wire _29210_;
wire _29211_;
wire _29212_;
wire _29213_;
wire _29214_;
wire _29215_;
wire _29216_;
wire _29217_;
wire _29218_;
wire _29219_;
wire _29220_;
wire _29221_;
wire _29222_;
wire _29223_;
wire _29224_;
wire _29225_;
wire _29226_;
wire _29227_;
wire _29228_;
wire _29229_;
wire _29230_;
wire _29231_;
wire _29232_;
wire _29233_;
wire _29234_;
wire _29235_;
wire _29236_;
wire _29237_;
wire _29238_;
wire _29239_;
wire _29240_;
wire _29241_;
wire _29242_;
wire _29243_;
wire _29244_;
wire _29245_;
wire _29246_;
wire _29247_;
wire _29248_;
wire _29249_;
wire _29250_;
wire _29251_;
wire _29252_;
wire _29253_;
wire _29254_;
wire _29255_;
wire _29256_;
wire _29257_;
wire _29258_;
wire _29259_;
wire _29260_;
wire _29261_;
wire _29262_;
wire _29263_;
wire _29264_;
wire _29265_;
wire _29266_;
wire _29267_;
wire _29268_;
wire _29269_;
wire _29270_;
wire _29271_;
wire _29272_;
wire _29273_;
wire _29274_;
wire _29275_;
wire _29276_;
wire _29277_;
wire _29278_;
wire _29279_;
wire _29280_;
wire _29281_;
wire _29282_;
wire _29283_;
wire _29284_;
wire _29285_;
wire _29286_;
wire _29287_;
wire _29288_;
wire _29289_;
wire _29290_;
wire _29291_;
wire _29292_;
wire _29293_;
wire _29294_;
wire _29295_;
wire _29296_;
wire _29297_;
wire _29298_;
wire _29299_;
wire _29300_;
wire _29301_;
wire _29302_;
wire _29303_;
wire _29304_;
wire _29305_;
wire _29306_;
wire _29307_;
wire _29308_;
wire _29309_;
wire _29310_;
wire _29311_;
wire _29312_;
wire _29313_;
wire _29314_;
wire _29315_;
wire _29316_;
wire _29317_;
wire _29318_;
wire _29319_;
wire _29320_;
wire _29321_;
wire _29322_;
wire _29323_;
wire _29324_;
wire _29325_;
wire _29326_;
wire _29327_;
wire _29328_;
wire _29329_;
wire _29330_;
wire _29331_;
wire _29332_;
wire _29333_;
wire _29334_;
wire _29335_;
wire _29336_;
wire _29337_;
wire _29338_;
wire _29339_;
wire _29340_;
wire _29341_;
wire _29342_;
wire _29343_;
wire _29344_;
wire _29345_;
wire _29346_;
wire _29347_;
wire _29348_;
wire _29349_;
wire _29350_;
wire _29351_;
wire _29352_;
wire _29353_;
wire _29354_;
wire _29355_;
wire _29356_;
wire _29357_;
wire _29358_;
wire _29359_;
wire _29360_;
wire _29361_;
wire _29362_;
wire _29363_;
wire _29364_;
wire _29365_;
wire _29366_;
wire _29367_;
wire _29368_;
wire _29369_;
wire _29370_;
wire _29371_;
wire _29372_;
wire _29373_;
wire _29374_;
wire _29375_;
wire _29376_;
wire _29377_;
wire _29378_;
wire _29379_;
wire _29380_;
wire _29381_;
wire _29382_;
wire _29383_;
wire _29384_;
wire _29385_;
wire _29386_;
wire _29387_;
wire _29388_;
wire _29389_;
wire _29390_;
wire _29391_;
wire _29392_;
wire _29393_;
wire _29394_;
wire _29395_;
wire _29396_;
wire _29397_;
wire _29398_;
wire _29399_;
wire _29400_;
wire _29401_;
wire _29402_;
wire _29403_;
wire _29404_;
wire _29405_;
wire _29406_;
wire _29407_;
wire _29408_;
wire _29409_;
wire _29410_;
wire _29411_;
wire _29412_;
wire _29413_;
wire _29414_;
wire _29415_;
wire _29416_;
wire _29417_;
wire _29418_;
wire _29419_;
wire _29420_;
wire _29421_;
wire _29422_;
wire _29423_;
wire _29424_;
wire _29425_;
wire _29426_;
wire _29427_;
wire _29428_;
wire _29429_;
wire _29430_;
wire _29431_;
wire _29432_;
wire _29433_;
wire _29434_;
wire _29435_;
wire _29436_;
wire _29437_;
wire _29438_;
wire _29439_;
wire _29440_;
wire _29441_;
wire _29442_;
wire _29443_;
wire _29444_;
wire _29445_;
wire _29446_;
wire _29447_;
wire _29448_;
wire _29449_;
wire _29450_;
wire _29451_;
wire _29452_;
wire _29453_;
wire _29454_;
wire _29455_;
wire _29456_;
wire _29457_;
wire _29458_;
wire _29459_;
wire _29460_;
wire _29461_;
wire _29462_;
wire _29463_;
wire _29464_;
wire _29465_;
wire _29466_;
wire _29467_;
wire _29468_;
wire _29469_;
wire _29470_;
wire _29471_;
wire _29472_;
wire _29473_;
wire _29474_;
wire _29475_;
wire _29476_;
wire _29477_;
wire _29478_;
wire _29479_;
wire _29480_;
wire _29481_;
wire _29482_;
wire _29483_;
wire _29484_;
wire _29485_;
wire _29486_;
wire _29487_;
wire _29488_;
wire _29489_;
wire _29490_;
wire _29491_;
wire _29492_;
wire _29493_;
wire _29494_;
wire _29495_;
wire _29496_;
wire _29497_;
wire _29498_;
wire _29499_;
wire _29500_;
wire _29501_;
wire _29502_;
wire _29503_;
wire _29504_;
wire _29505_;
wire _29506_;
wire _29507_;
wire _29508_;
wire _29509_;
wire _29510_;
wire _29511_;
wire _29512_;
wire _29513_;
wire _29514_;
wire _29515_;
wire _29516_;
wire _29517_;
wire _29518_;
wire _29519_;
wire _29520_;
wire _29521_;
wire _29522_;
wire _29523_;
wire _29524_;
wire _29525_;
wire _29526_;
wire _29527_;
wire _29528_;
wire _29529_;
wire _29530_;
wire _29531_;
wire _29532_;
wire _29533_;
wire _29534_;
wire _29535_;
wire _29536_;
wire _29537_;
wire _29538_;
wire _29539_;
wire _29540_;
wire _29541_;
wire _29542_;
wire _29543_;
wire _29544_;
wire _29545_;
wire _29546_;
wire _29547_;
wire _29548_;
wire _29549_;
wire _29550_;
wire _29551_;
wire _29552_;
wire _29553_;
wire _29554_;
wire _29555_;
wire _29556_;
wire _29557_;
wire _29558_;
wire _29559_;
wire _29560_;
wire _29561_;
wire _29562_;
wire _29563_;
wire _29564_;
wire _29565_;
wire _29566_;
wire _29567_;
wire _29568_;
wire _29569_;
wire _29570_;
wire _29571_;
wire _29572_;
wire _29573_;
wire _29574_;
wire _29575_;
wire _29576_;
wire _29577_;
wire _29578_;
wire _29579_;
wire _29580_;
wire _29581_;
wire _29582_;
wire _29583_;
wire _29584_;
wire _29585_;
wire _29586_;
wire _29587_;
wire _29588_;
wire _29589_;
wire _29590_;
wire _29591_;
wire _29592_;
wire _29593_;
wire _29594_;
wire _29595_;
wire _29596_;
wire _29597_;
wire _29598_;
wire _29599_;
wire _29600_;
wire _29601_;
wire _29602_;
wire _29603_;
wire _29604_;
wire _29605_;
wire _29606_;
wire _29607_;
wire _29608_;
wire _29609_;
wire _29610_;
wire _29611_;
wire _29612_;
wire _29613_;
wire _29614_;
wire _29615_;
wire _29616_;
wire _29617_;
wire _29618_;
wire _29619_;
wire _29620_;
wire _29621_;
wire _29622_;
wire _29623_;
wire _29624_;
wire _29625_;
wire _29626_;
wire _29627_;
wire _29628_;
wire _29629_;
wire _29630_;
wire _29631_;
wire _29632_;
wire _29633_;
wire _29634_;
wire _29635_;
wire _29636_;
wire _29637_;
wire _29638_;
wire _29639_;
wire _29640_;
wire _29641_;
wire _29642_;
wire _29643_;
wire _29644_;
wire _29645_;
wire _29646_;
wire _29647_;
wire _29648_;
wire _29649_;
wire _29650_;
wire _29651_;
wire _29652_;
wire _29653_;
wire _29654_;
wire _29655_;
wire _29656_;
wire _29657_;
wire _29658_;
wire _29659_;
wire _29660_;
wire _29661_;
wire _29662_;
wire _29663_;
wire _29664_;
wire _29665_;
wire _29666_;
wire _29667_;
wire _29668_;
wire _29669_;
wire _29670_;
wire _29671_;
wire _29672_;
wire _29673_;
wire _29674_;
wire _29675_;
wire _29676_;
wire _29677_;
wire _29678_;
wire _29679_;
wire _29680_;
wire _29681_;
wire _29682_;
wire _29683_;
wire _29684_;
wire _29685_;
wire _29686_;
wire _29687_;
wire _29688_;
wire _29689_;
wire _29690_;
wire _29691_;
wire _29692_;
wire _29693_;
wire _29694_;
wire _29695_;
wire _29696_;
wire _29697_;
wire _29698_;
wire _29699_;
wire _29700_;
wire _29701_;
wire _29702_;
wire _29703_;
wire _29704_;
wire _29705_;
wire _29706_;
wire _29707_;
wire _29708_;
wire _29709_;
wire _29710_;
wire _29711_;
wire _29712_;
wire _29713_;
wire _29714_;
wire _29715_;
wire _29716_;
wire _29717_;
wire _29718_;
wire _29719_;
wire _29720_;
wire _29721_;
wire _29722_;
wire _29723_;
wire _29724_;
wire _29725_;
wire _29726_;
wire _29727_;
wire _29728_;
wire _29729_;
wire _29730_;
wire _29731_;
wire _29732_;
wire _29733_;
wire _29734_;
wire _29735_;
wire _29736_;
wire _29737_;
wire _29738_;
wire _29739_;
wire _29740_;
wire _29741_;
wire _29742_;
wire _29743_;
wire _29744_;
wire _29745_;
wire _29746_;
wire _29747_;
wire _29748_;
wire _29749_;
wire _29750_;
wire _29751_;
wire _29752_;
wire _29753_;
wire _29754_;
wire _29755_;
wire _29756_;
wire _29757_;
wire _29758_;
wire _29759_;
wire _29760_;
wire _29761_;
wire _29762_;
wire _29763_;
wire _29764_;
wire _29765_;
wire _29766_;
wire _29767_;
wire _29768_;
wire _29769_;
wire _29770_;
wire _29771_;
wire _29772_;
wire _29773_;
wire _29774_;
wire _29775_;
wire _29776_;
wire _29777_;
wire _29778_;
wire _29779_;
wire _29780_;
wire _29781_;
wire _29782_;
wire _29783_;
wire _29784_;
wire _29785_;
wire _29786_;
wire _29787_;
wire _29788_;
wire _29789_;
wire _29790_;
wire _29791_;
wire _29792_;
wire _29793_;
wire _29794_;
wire _29795_;
wire _29796_;
wire _29797_;
wire _29798_;
wire _29799_;
wire _29800_;
wire _29801_;
wire _29802_;
wire _29803_;
wire _29804_;
wire _29805_;
wire _29806_;
wire _29807_;
wire _29808_;
wire _29809_;
wire _29810_;
wire _29811_;
wire _29812_;
wire _29813_;
wire _29814_;
wire _29815_;
wire _29816_;
wire _29817_;
wire _29818_;
wire _29819_;
wire _29820_;
wire _29821_;
wire _29822_;
wire _29823_;
wire _29824_;
wire _29825_;
wire _29826_;
wire _29827_;
wire _29828_;
wire _29829_;
wire _29830_;
wire _29831_;
wire _29832_;
wire _29833_;
wire _29834_;
wire _29835_;
wire _29836_;
wire _29837_;
wire _29838_;
wire _29839_;
wire _29840_;
wire _29841_;
wire _29842_;
wire _29843_;
wire _29844_;
wire _29845_;
wire _29846_;
wire _29847_;
wire _29848_;
wire _29849_;
wire _29850_;
wire _29851_;
wire _29852_;
wire _29853_;
wire _29854_;
wire _29855_;
wire _29856_;
wire _29857_;
wire _29858_;
wire _29859_;
wire _29860_;
wire _29861_;
wire _29862_;
wire _29863_;
wire _29864_;
wire _29865_;
wire _29866_;
wire _29867_;
wire _29868_;
wire _29869_;
wire _29870_;
wire _29871_;
wire _29872_;
wire _29873_;
wire _29874_;
wire _29875_;
wire _29876_;
wire _29877_;
wire _29878_;
wire _29879_;
wire _29880_;
wire _29881_;
wire _29882_;
wire _29883_;
wire _29884_;
wire _29885_;
wire _29886_;
wire _29887_;
wire _29888_;
wire _29889_;
wire _29890_;
wire _29891_;
wire _29892_;
wire _29893_;
wire _29894_;
wire _29895_;
wire _29896_;
wire _29897_;
wire _29898_;
wire _29899_;
wire _29900_;
wire _29901_;
wire _29902_;
wire _29903_;
wire _29904_;
wire _29905_;
wire _29906_;
wire _29907_;
wire _29908_;
wire _29909_;
wire _29910_;
wire _29911_;
wire _29912_;
wire _29913_;
wire _29914_;
wire _29915_;
wire _29916_;
wire _29917_;
wire _29918_;
wire _29919_;
wire _29920_;
wire _29921_;
wire _29922_;
wire _29923_;
wire _29924_;
wire _29925_;
wire _29926_;
wire _29927_;
wire _29928_;
wire _29929_;
wire _29930_;
wire _29931_;
wire _29932_;
wire _29933_;
wire _29934_;
wire _29935_;
wire _29936_;
wire _29937_;
wire _29938_;
wire _29939_;
wire _29940_;
wire _29941_;
wire _29942_;
wire _29943_;
wire _29944_;
wire _29945_;
wire _29946_;
wire _29947_;
wire _29948_;
wire _29949_;
wire _29950_;
wire _29951_;
wire _29952_;
wire _29953_;
wire _29954_;
wire _29955_;
wire _29956_;
wire _29957_;
wire _29958_;
wire _29959_;
wire _29960_;
wire _29961_;
wire _29962_;
wire _29963_;
wire _29964_;
wire _29965_;
wire _29966_;
wire _29967_;
wire _29968_;
wire _29969_;
wire _29970_;
wire _29971_;
wire _29972_;
wire _29973_;
wire _29974_;
wire _29975_;
wire _29976_;
wire _29977_;
wire _29978_;
wire _29979_;
wire _29980_;
wire _29981_;
wire _29982_;
wire _29983_;
wire _29984_;
wire _29985_;
wire _29986_;
wire _29987_;
wire _29988_;
wire _29989_;
wire _29990_;
wire _29991_;
wire _29992_;
wire _29993_;
wire _29994_;
wire _29995_;
wire _29996_;
wire _29997_;
wire _29998_;
wire _29999_;
wire _30000_;
wire _30001_;
wire _30002_;
wire _30003_;
wire _30004_;
wire _30005_;
wire _30006_;
wire _30007_;
wire _30008_;
wire _30009_;
wire _30010_;
wire _30011_;
wire _30012_;
wire _30013_;
wire _30014_;
wire _30015_;
wire _30016_;
wire _30017_;
wire _30018_;
wire _30019_;
wire _30020_;
wire _30021_;
wire _30022_;
wire _30023_;
wire _30024_;
wire _30025_;
wire _30026_;
wire _30027_;
wire _30028_;
wire _30029_;
wire _30030_;
wire _30031_;
wire _30032_;
wire _30033_;
wire _30034_;
wire _30035_;
wire _30036_;
wire _30037_;
wire _30038_;
wire _30039_;
wire _30040_;
wire _30041_;
wire _30042_;
wire _30043_;
wire _30044_;
wire _30045_;
wire _30046_;
wire _30047_;
wire _30048_;
wire _30049_;
wire _30050_;
wire _30051_;
wire _30052_;
wire _30053_;
wire _30054_;
wire _30055_;
wire _30056_;
wire _30057_;
wire _30058_;
wire _30059_;
wire _30060_;
wire _30061_;
wire _30062_;
wire _30063_;
wire _30064_;
wire _30065_;
wire _30066_;
wire _30067_;
wire _30068_;
wire _30069_;
wire _30070_;
wire _30071_;
wire _30072_;
wire _30073_;
wire _30074_;
wire _30075_;
wire _30076_;
wire _30077_;
wire _30078_;
wire _30079_;
wire _30080_;
wire _30081_;
wire _30082_;
wire _30083_;
wire _30084_;
wire _30085_;
wire _30086_;
wire _30087_;
wire _30088_;
wire _30089_;
wire _30090_;
wire _30091_;
wire _30092_;
wire _30093_;
wire _30094_;
wire _30095_;
wire _30096_;
wire _30097_;
wire _30098_;
wire _30099_;
wire _30100_;
wire _30101_;
wire _30102_;
wire _30103_;
wire _30104_;
wire _30105_;
wire _30106_;
wire _30107_;
wire _30108_;
wire _30109_;
wire _30110_;
wire _30111_;
wire _30112_;
wire _30113_;
wire _30114_;
wire _30115_;
wire _30116_;
wire _30117_;
wire _30118_;
wire _30119_;
wire _30120_;
wire _30121_;
wire _30122_;
wire _30123_;
wire _30124_;
wire _30125_;
wire _30126_;
wire _30127_;
wire _30128_;
wire _30129_;
wire _30130_;
wire _30131_;
wire _30132_;
wire _30133_;
wire _30134_;
wire _30135_;
wire _30136_;
wire _30137_;
wire _30138_;
wire _30139_;
wire _30140_;
wire _30141_;
wire _30142_;
wire _30143_;
wire _30144_;
wire _30145_;
wire _30146_;
wire _30147_;
wire _30148_;
wire _30149_;
wire _30150_;
wire _30151_;
wire _30152_;
wire _30153_;
wire _30154_;
wire _30155_;
wire _30156_;
wire _30157_;
wire _30158_;
wire _30159_;
wire _30160_;
wire _30161_;
wire _30162_;
wire _30163_;
wire _30164_;
wire _30165_;
wire _30166_;
wire _30167_;
wire _30168_;
wire _30169_;
wire _30170_;
wire _30171_;
wire _30172_;
wire _30173_;
wire _30174_;
wire _30175_;
wire _30176_;
wire _30177_;
wire _30178_;
wire _30179_;
wire _30180_;
wire _30181_;
wire _30182_;
wire _30183_;
wire _30184_;
wire _30185_;
wire _30186_;
wire _30187_;
wire _30188_;
wire _30189_;
wire _30190_;
wire _30191_;
wire _30192_;
wire _30193_;
wire _30194_;
wire _30195_;
wire _30196_;
wire _30197_;
wire _30198_;
wire _30199_;
wire _30200_;
wire _30201_;
wire _30202_;
wire _30203_;
wire _30204_;
wire _30205_;
wire _30206_;
wire _30207_;
wire _30208_;
wire _30209_;
wire _30210_;
wire _30211_;
wire _30212_;
wire _30213_;
wire _30214_;
wire _30215_;
wire _30216_;
wire _30217_;
wire _30218_;
wire _30219_;
wire _30220_;
wire _30221_;
wire _30222_;
wire _30223_;
wire _30224_;
wire _30225_;
wire _30226_;
wire _30227_;
wire _30228_;
wire _30229_;
wire _30230_;
wire _30231_;
wire _30232_;
wire _30233_;
wire _30234_;
wire _30235_;
wire _30236_;
wire _30237_;
wire _30238_;
wire _30239_;
wire _30240_;
wire _30241_;
wire _30242_;
wire _30243_;
wire _30244_;
wire _30245_;
wire _30246_;
wire _30247_;
wire _30248_;
wire _30249_;
wire _30250_;
wire _30251_;
wire _30252_;
wire _30253_;
wire _30254_;
wire _30255_;
wire _30256_;
wire _30257_;
wire _30258_;
wire _30259_;
wire _30260_;
wire _30261_;
wire _30262_;
wire _30263_;
wire _30264_;
wire _30265_;
wire _30266_;
wire _30267_;
wire _30268_;
wire _30269_;
wire _30270_;
wire _30271_;
wire _30272_;
wire _30273_;
wire _30274_;
wire _30275_;
wire _30276_;
wire _30277_;
wire _30278_;
wire _30279_;
wire _30280_;
wire _30281_;
wire _30282_;
wire _30283_;
wire _30284_;
wire _30285_;
wire _30286_;
wire _30287_;
wire _30288_;
wire _30289_;
wire _30290_;
wire _30291_;
wire _30292_;
wire _30293_;
wire _30294_;
wire _30295_;
wire _30296_;
wire _30297_;
wire _30298_;
wire _30299_;
wire _30300_;
wire _30301_;
wire _30302_;
wire _30303_;
wire _30304_;
wire _30305_;
wire _30306_;
wire _30307_;
wire _30308_;
wire _30309_;
wire _30310_;
wire _30311_;
wire _30312_;
wire _30313_;
wire _30314_;
wire _30315_;
wire _30316_;
wire _30317_;
wire _30318_;
wire _30319_;
wire _30320_;
wire _30321_;
wire _30322_;
wire _30323_;
wire _30324_;
wire _30325_;
wire _30326_;
wire _30327_;
wire _30328_;
wire _30329_;
wire _30330_;
wire _30331_;
wire _30332_;
wire _30333_;
wire _30334_;
wire _30335_;
wire _30336_;
wire _30337_;
wire _30338_;
wire _30339_;
wire _30340_;
wire _30341_;
wire _30342_;
wire _30343_;
wire _30344_;
wire _30345_;
wire _30346_;
wire _30347_;
wire _30348_;
wire _30349_;
wire _30350_;
wire _30351_;
wire _30352_;
wire _30353_;
wire _30354_;
wire _30355_;
wire _30356_;
wire _30357_;
wire _30358_;
wire _30359_;
wire _30360_;
wire _30361_;
wire _30362_;
wire _30363_;
wire _30364_;
wire _30365_;
wire _30366_;
wire _30367_;
wire _30368_;
wire _30369_;
wire _30370_;
wire _30371_;
wire _30372_;
wire _30373_;
wire _30374_;
wire _30375_;
wire _30376_;
wire _30377_;
wire _30378_;
wire _30379_;
wire _30380_;
wire _30381_;
wire _30382_;
wire _30383_;
wire _30384_;
wire _30385_;
wire _30386_;
wire _30387_;
wire _30388_;
wire _30389_;
wire _30390_;
wire _30391_;
wire _30392_;
wire _30393_;
wire _30394_;
wire _30395_;
wire _30396_;
wire _30397_;
wire _30398_;
wire _30399_;
wire _30400_;
wire _30401_;
wire _30402_;
wire _30403_;
wire _30404_;
wire _30405_;
wire _30406_;
wire _30407_;
wire _30408_;
wire _30409_;
wire _30410_;
wire _30411_;
wire _30412_;
wire _30413_;
wire _30414_;
wire _30415_;
wire _30416_;
wire _30417_;
wire _30418_;
wire _30419_;
wire _30420_;
wire _30421_;
wire _30422_;
wire _30423_;
wire _30424_;
wire _30425_;
wire _30426_;
wire _30427_;
wire _30428_;
wire _30429_;
wire _30430_;
wire _30431_;
wire _30432_;
wire _30433_;
wire _30434_;
wire _30435_;
wire _30436_;
wire _30437_;
wire _30438_;
wire _30439_;
wire _30440_;
wire _30441_;
wire _30442_;
wire _30443_;
wire _30444_;
wire _30445_;
wire _30446_;
wire _30447_;
wire _30448_;
wire _30449_;
wire _30450_;
wire _30451_;
wire _30452_;
wire _30453_;
wire _30454_;
wire _30455_;
wire _30456_;
wire _30457_;
wire _30458_;
wire _30459_;
wire _30460_;
wire _30461_;
wire _30462_;
wire _30463_;
wire _30464_;
wire _30465_;
wire _30466_;
wire _30467_;
wire _30468_;
wire _30469_;
wire _30470_;
wire _30471_;
wire _30472_;
wire _30473_;
wire _30474_;
wire _30475_;
wire _30476_;
wire _30477_;
wire _30478_;
wire _30479_;
wire _30480_;
wire _30481_;
wire _30482_;
wire _30483_;
wire _30484_;
wire _30485_;
wire _30486_;
wire _30487_;
wire _30488_;
wire _30489_;
wire _30490_;
wire _30491_;
wire _30492_;
wire _30493_;
wire _30494_;
wire _30495_;
wire _30496_;
wire _30497_;
wire _30498_;
wire _30499_;
wire _30500_;
wire _30501_;
wire _30502_;
wire _30503_;
wire _30504_;
wire _30505_;
wire _30506_;
wire _30507_;
wire _30508_;
wire _30509_;
wire _30510_;
wire _30511_;
wire _30512_;
wire _30513_;
wire _30514_;
wire _30515_;
wire _30516_;
wire _30517_;
wire _30518_;
wire _30519_;
wire _30520_;
wire _30521_;
wire _30522_;
wire _30523_;
wire _30524_;
wire _30525_;
wire _30526_;
wire _30527_;
wire _30528_;
wire _30529_;
wire _30530_;
wire _30531_;
wire _30532_;
wire _30533_;
wire _30534_;
wire _30535_;
wire _30536_;
wire _30537_;
wire _30538_;
wire _30539_;
wire _30540_;
wire _30541_;
wire _30542_;
wire _30543_;
wire _30544_;
wire _30545_;
wire _30546_;
wire _30547_;
wire _30548_;
wire _30549_;
wire _30550_;
wire _30551_;
wire _30552_;
wire _30553_;
wire _30554_;
wire _30555_;
wire _30556_;
wire _30557_;
wire _30558_;
wire _30559_;
wire _30560_;
wire _30561_;
wire _30562_;
wire _30563_;
wire _30564_;
wire _30565_;
wire _30566_;
wire _30567_;
wire _30568_;
wire _30569_;
wire _30570_;
wire _30571_;
wire _30572_;
wire _30573_;
wire _30574_;
wire _30575_;
wire _30576_;
wire _30577_;
wire _30578_;
wire _30579_;
wire _30580_;
wire _30581_;
wire _30582_;
wire _30583_;
wire _30584_;
wire _30585_;
wire _30586_;
wire _30587_;
wire _30588_;
wire _30589_;
wire _30590_;
wire _30591_;
wire _30592_;
wire _30593_;
wire _30594_;
wire _30595_;
wire _30596_;
wire _30597_;
wire _30598_;
wire _30599_;
wire _30600_;
wire _30601_;
wire _30602_;
wire _30603_;
wire _30604_;
wire _30605_;
wire _30606_;
wire _30607_;
wire _30608_;
wire _30609_;
wire _30610_;
wire _30611_;
wire _30612_;
wire _30613_;
wire _30614_;
wire _30615_;
wire _30616_;
wire _30617_;
wire _30618_;
wire _30619_;
wire _30620_;
wire _30621_;
wire _30622_;
wire _30623_;
wire _30624_;
wire _30625_;
wire _30626_;
wire _30627_;
wire _30628_;
wire _30629_;
wire _30630_;
wire _30631_;
wire _30632_;
wire _30633_;
wire _30634_;
wire _30635_;
wire _30636_;
wire _30637_;
wire _30638_;
wire _30639_;
wire _30640_;
wire _30641_;
wire _30642_;
wire _30643_;
wire _30644_;
wire _30645_;
wire _30646_;
wire _30647_;
wire _30648_;
wire _30649_;
wire _30650_;
wire _30651_;
wire _30652_;
wire _30653_;
wire _30654_;
wire _30655_;
wire _30656_;
wire _30657_;
wire _30658_;
wire _30659_;
wire _30660_;
wire _30661_;
wire _30662_;
wire _30663_;
wire _30664_;
wire _30665_;
wire _30666_;
wire _30667_;
wire _30668_;
wire _30669_;
wire _30670_;
wire _30671_;
wire _30672_;
wire _30673_;
wire _30674_;
wire _30675_;
wire _30676_;
wire _30677_;
wire _30678_;
wire _30679_;
wire _30680_;
wire _30681_;
wire _30682_;
wire _30683_;
wire _30684_;
wire _30685_;
wire _30686_;
wire _30687_;
wire _30688_;
wire _30689_;
wire _30690_;
wire _30691_;
wire _30692_;
wire _30693_;
wire _30694_;
wire _30695_;
wire _30696_;
wire _30697_;
wire _30698_;
wire _30699_;
wire _30700_;
wire _30701_;
wire _30702_;
wire _30703_;
wire _30704_;
wire _30705_;
wire _30706_;
wire _30707_;
wire _30708_;
wire _30709_;
wire _30710_;
wire _30711_;
wire _30712_;
wire _30713_;
wire _30714_;
wire _30715_;
wire _30716_;
wire _30717_;
wire _30718_;
wire _30719_;
wire _30720_;
wire _30721_;
wire _30722_;
wire _30723_;
wire _30724_;
wire _30725_;
wire _30726_;
wire _30727_;
wire _30728_;
wire _30729_;
wire _30730_;
wire _30731_;
wire _30732_;
wire _30733_;
wire _30734_;
wire _30735_;
wire _30736_;
wire _30737_;
wire _30738_;
wire _30739_;
wire _30740_;
wire _30741_;
wire _30742_;
wire _30743_;
wire _30744_;
wire _30745_;
wire _30746_;
wire _30747_;
wire _30748_;
wire _30749_;
wire _30750_;
wire _30751_;
wire _30752_;
wire _30753_;
wire _30754_;
wire _30755_;
wire _30756_;
wire _30757_;
wire _30758_;
wire _30759_;
wire _30760_;
wire _30761_;
wire _30762_;
wire _30763_;
wire _30764_;
wire _30765_;
wire _30766_;
wire _30767_;
wire _30768_;
wire _30769_;
wire _30770_;
wire _30771_;
wire _30772_;
wire _30773_;
wire _30774_;
wire _30775_;
wire _30776_;
wire _30777_;
wire _30778_;
wire _30779_;
wire _30780_;
wire _30781_;
wire _30782_;
wire _30783_;
wire _30784_;
wire _30785_;
wire _30786_;
wire _30787_;
wire _30788_;
wire _30789_;
wire _30790_;
wire _30791_;
wire _30792_;
wire _30793_;
wire _30794_;
wire _30795_;
wire _30796_;
wire _30797_;
wire _30798_;
wire _30799_;
wire _30800_;
wire _30801_;
wire _30802_;
wire _30803_;
wire _30804_;
wire _30805_;
wire _30806_;
wire _30807_;
wire _30808_;
wire _30809_;
wire _30810_;
wire _30811_;
wire _30812_;
wire _30813_;
wire _30814_;
wire _30815_;
wire _30816_;
wire _30817_;
wire _30818_;
wire _30819_;
wire _30820_;
wire _30821_;
wire _30822_;
wire _30823_;
wire _30824_;
wire _30825_;
wire _30826_;
wire _30827_;
wire _30828_;
wire _30829_;
wire _30830_;
wire _30831_;
wire _30832_;
wire _30833_;
wire _30834_;
wire _30835_;
wire _30836_;
wire _30837_;
wire _30838_;
wire _30839_;
wire _30840_;
wire _30841_;
wire _30842_;
wire _30843_;
wire _30844_;
wire _30845_;
wire _30846_;
wire _30847_;
wire _30848_;
wire _30849_;
wire _30850_;
wire _30851_;
wire _30852_;
wire _30853_;
wire _30854_;
wire _30855_;
wire _30856_;
wire _30857_;
wire _30858_;
wire _30859_;
wire _30860_;
wire _30861_;
wire _30862_;
wire _30863_;
wire _30864_;
wire _30865_;
wire _30866_;
wire _30867_;
wire _30868_;
wire _30869_;
wire _30870_;
wire _30871_;
wire _30872_;
wire _30873_;
wire _30874_;
wire _30875_;
wire _30876_;
wire _30877_;
wire _30878_;
wire _30879_;
wire _30880_;
wire _30881_;
wire _30882_;
wire _30883_;
wire _30884_;
wire _30885_;
wire _30886_;
wire _30887_;
wire _30888_;
wire _30889_;
wire _30890_;
wire _30891_;
wire _30892_;
wire _30893_;
wire _30894_;
wire _30895_;
wire _30896_;
wire _30897_;
wire _30898_;
wire _30899_;
wire _30900_;
wire _30901_;
wire _30902_;
wire _30903_;
wire _30904_;
wire _30905_;
wire _30906_;
wire _30907_;
wire _30908_;
wire _30909_;
wire _30910_;
wire _30911_;
wire _30912_;
wire _30913_;
wire _30914_;
wire _30915_;
wire _30916_;
wire _30917_;
wire _30918_;
wire _30919_;
wire _30920_;
wire _30921_;
wire _30922_;
wire _30923_;
wire _30924_;
wire _30925_;
wire _30926_;
wire _30927_;
wire _30928_;
wire _30929_;
wire _30930_;
wire _30931_;
wire _30932_;
wire _30933_;
wire _30934_;
wire _30935_;
wire _30936_;
wire _30937_;
wire _30938_;
wire _30939_;
wire _30940_;
wire _30941_;
wire _30942_;
wire _30943_;
wire _30944_;
wire _30945_;
wire _30946_;
wire _30947_;
wire _30948_;
wire _30949_;
wire _30950_;
wire _30951_;
wire _30952_;
wire _30953_;
wire _30954_;
wire _30955_;
wire _30956_;
wire _30957_;
wire _30958_;
wire _30959_;
wire _30960_;
wire _30961_;
wire _30962_;
wire _30963_;
wire _30964_;
wire _30965_;
wire _30966_;
wire _30967_;
wire _30968_;
wire _30969_;
wire _30970_;
wire _30971_;
wire _30972_;
wire _30973_;
wire _30974_;
wire _30975_;
wire _30976_;
wire _30977_;
wire _30978_;
wire _30979_;
wire _30980_;
wire _30981_;
wire _30982_;
wire _30983_;
wire _30984_;
wire _30985_;
wire _30986_;
wire _30987_;
wire _30988_;
wire _30989_;
wire _30990_;
wire _30991_;
wire _30992_;
wire _30993_;
wire _30994_;
wire _30995_;
wire _30996_;
wire _30997_;
wire _30998_;
wire _30999_;
wire _31000_;
wire _31001_;
wire _31002_;
wire _31003_;
wire _31004_;
wire _31005_;
wire _31006_;
wire _31007_;
wire _31008_;
wire _31009_;
wire _31010_;
wire _31011_;
wire _31012_;
wire _31013_;
wire _31014_;
wire _31015_;
wire _31016_;
wire _31017_;
wire _31018_;
wire _31019_;
wire _31020_;
wire _31021_;
wire _31022_;
wire _31023_;
wire _31024_;
wire _31025_;
wire _31026_;
wire _31027_;
wire _31028_;
wire _31029_;
wire _31030_;
wire _31031_;
wire _31032_;
wire _31033_;
wire _31034_;
wire _31035_;
wire _31036_;
wire _31037_;
wire _31038_;
wire _31039_;
wire _31040_;
wire _31041_;
wire _31042_;
wire _31043_;
wire _31044_;
wire _31045_;
wire _31046_;
wire _31047_;
wire _31048_;
wire _31049_;
wire _31050_;
wire _31051_;
wire _31052_;
wire _31053_;
wire _31054_;
wire _31055_;
wire _31056_;
wire _31057_;
wire _31058_;
wire _31059_;
wire _31060_;
wire _31061_;
wire _31062_;
wire _31063_;
wire _31064_;
wire _31065_;
wire _31066_;
wire _31067_;
wire _31068_;
wire _31069_;
wire _31070_;
wire _31071_;
wire _31072_;
wire _31073_;
wire _31074_;
wire _31075_;
wire _31076_;
wire _31077_;
wire _31078_;
wire _31079_;
wire _31080_;
wire _31081_;
wire _31082_;
wire _31083_;
wire _31084_;
wire _31085_;
wire _31086_;
wire _31087_;
wire _31088_;
wire _31089_;
wire _31090_;
wire _31091_;
wire _31092_;
wire _31093_;
wire _31094_;
wire _31095_;
wire _31096_;
wire _31097_;
wire _31098_;
wire _31099_;
wire _31100_;
wire _31101_;
wire _31102_;
wire _31103_;
wire _31104_;
wire _31105_;
wire _31106_;
wire _31107_;
wire _31108_;
wire _31109_;
wire _31110_;
wire _31111_;
wire _31112_;
wire _31113_;
wire _31114_;
wire _31115_;
wire _31116_;
wire _31117_;
wire _31118_;
wire _31119_;
wire _31120_;
wire _31121_;
wire _31122_;
wire _31123_;
wire _31124_;
wire _31125_;
wire _31126_;
wire _31127_;
wire _31128_;
wire _31129_;
wire _31130_;
wire _31131_;
wire _31132_;
wire _31133_;
wire _31134_;
wire _31135_;
wire _31136_;
wire _31137_;
wire _31138_;
wire _31139_;
wire _31140_;
wire _31141_;
wire _31142_;
wire _31143_;
wire _31144_;
wire _31145_;
wire _31146_;
wire _31147_;
wire _31148_;
wire _31149_;
wire _31150_;
wire _31151_;
wire _31152_;
wire _31153_;
wire _31154_;
wire _31155_;
wire _31156_;
wire _31157_;
wire _31158_;
wire _31159_;
wire _31160_;
wire _31161_;
wire _31162_;
wire _31163_;
wire _31164_;
wire _31165_;
wire _31166_;
wire _31167_;
wire _31168_;
wire _31169_;
wire _31170_;
wire _31171_;
wire _31172_;
wire _31173_;
wire _31174_;
wire _31175_;
wire _31176_;
wire _31177_;
wire _31178_;
wire _31179_;
wire _31180_;
wire _31181_;
wire _31182_;
wire _31183_;
wire _31184_;
wire _31185_;
wire _31186_;
wire _31187_;
wire _31188_;
wire _31189_;
wire _31190_;
wire _31191_;
wire _31192_;
wire _31193_;
wire _31194_;
wire _31195_;
wire _31196_;
wire _31197_;
wire _31198_;
wire _31199_;
wire _31200_;
wire _31201_;
wire _31202_;
wire _31203_;
wire _31204_;
wire _31205_;
wire _31206_;
wire _31207_;
wire _31208_;
wire _31209_;
wire _31210_;
wire _31211_;
wire _31212_;
wire _31213_;
wire _31214_;
wire _31215_;
wire _31216_;
wire _31217_;
wire _31218_;
wire _31219_;
wire _31220_;
wire _31221_;
wire _31222_;
wire _31223_;
wire _31224_;
wire _31225_;
wire _31226_;
wire _31227_;
wire _31228_;
wire _31229_;
wire _31230_;
wire _31231_;
wire _31232_;
wire _31233_;
wire _31234_;
wire _31235_;
wire _31236_;
wire _31237_;
wire _31238_;
wire _31239_;
wire _31240_;
wire _31241_;
wire _31242_;
wire _31243_;
wire _31244_;
wire _31245_;
wire _31246_;
wire _31247_;
wire _31248_;
wire _31249_;
wire _31250_;
wire _31251_;
wire _31252_;
wire _31253_;
wire _31254_;
wire _31255_;
wire _31256_;
wire _31257_;
wire _31258_;
wire _31259_;
wire _31260_;
wire _31261_;
wire _31262_;
wire _31263_;
wire _31264_;
wire _31265_;
wire _31266_;
wire _31267_;
wire _31268_;
wire _31269_;
wire _31270_;
wire _31271_;
wire _31272_;
wire _31273_;
wire _31274_;
wire _31275_;
wire _31276_;
wire _31277_;
wire _31278_;
wire _31279_;
wire _31280_;
wire _31281_;
wire _31282_;
wire _31283_;
wire _31284_;
wire _31285_;
wire _31286_;
wire _31287_;
wire _31288_;
wire _31289_;
wire _31290_;
wire _31291_;
wire _31292_;
wire _31293_;
wire _31294_;
wire _31295_;
wire _31296_;
wire _31297_;
wire _31298_;
wire _31299_;
wire _31300_;
wire _31301_;
wire _31302_;
wire _31303_;
wire _31304_;
wire _31305_;
wire _31306_;
wire _31307_;
wire _31308_;
wire _31309_;
wire _31310_;
wire _31311_;
wire _31312_;
wire _31313_;
wire _31314_;
wire _31315_;
wire _31316_;
wire _31317_;
wire _31318_;
wire _31319_;
wire _31320_;
wire _31321_;
wire _31322_;
wire _31323_;
wire _31324_;
wire _31325_;
wire _31326_;
wire _31327_;
wire _31328_;
wire _31329_;
wire _31330_;
wire _31331_;
wire _31332_;
wire _31333_;
wire _31334_;
wire _31335_;
wire _31336_;
wire _31337_;
wire _31338_;
wire _31339_;
wire _31340_;
wire _31341_;
wire _31342_;
wire _31343_;
wire _31344_;
wire _31345_;
wire _31346_;
wire _31347_;
wire _31348_;
wire _31349_;
wire _31350_;
wire _31351_;
wire _31352_;
wire _31353_;
wire _31354_;
wire _31355_;
wire _31356_;
wire _31357_;
wire _31358_;
wire _31359_;
wire _31360_;
wire _31361_;
wire _31362_;
wire _31363_;
wire _31364_;
wire _31365_;
wire _31366_;
wire _31367_;
wire _31368_;
wire _31369_;
wire _31370_;
wire _31371_;
wire _31372_;
wire _31373_;
wire _31374_;
wire _31375_;
wire _31376_;
wire _31377_;
wire _31378_;
wire _31379_;
wire _31380_;
wire _31381_;
wire _31382_;
wire _31383_;
wire _31384_;
wire _31385_;
wire _31386_;
wire _31387_;
wire _31388_;
wire _31389_;
wire _31390_;
wire _31391_;
wire _31392_;
wire _31393_;
wire _31394_;
wire _31395_;
wire _31396_;
wire _31397_;
wire _31398_;
wire _31399_;
wire _31400_;
wire _31401_;
wire _31402_;
wire _31403_;
wire _31404_;
wire _31405_;
wire _31406_;
wire _31407_;
wire _31408_;
wire _31409_;
wire _31410_;
wire _31411_;
wire _31412_;
wire _31413_;
wire _31414_;
wire _31415_;
wire _31416_;
wire _31417_;
wire _31418_;
wire _31419_;
wire _31420_;
wire _31421_;
wire _31422_;
wire _31423_;
wire _31424_;
wire _31425_;
wire _31426_;
wire _31427_;
wire _31428_;
wire _31429_;
wire _31430_;
wire _31431_;
wire _31432_;
wire _31433_;
wire _31434_;
wire _31435_;
wire _31436_;
wire _31437_;
wire _31438_;
wire _31439_;
wire _31440_;
wire _31441_;
wire _31442_;
wire _31443_;
wire _31444_;
wire _31445_;
wire _31446_;
wire _31447_;
wire _31448_;
wire _31449_;
wire _31450_;
wire _31451_;
wire _31452_;
wire _31453_;
wire _31454_;
wire _31455_;
wire _31456_;
wire _31457_;
wire _31458_;
wire _31459_;
wire _31460_;
wire _31461_;
wire _31462_;
wire _31463_;
wire _31464_;
wire _31465_;
wire _31466_;
wire _31467_;
wire _31468_;
wire _31469_;
wire _31470_;
wire _31471_;
wire _31472_;
wire _31473_;
wire _31474_;
wire _31475_;
wire _31476_;
wire _31477_;
wire _31478_;
wire _31479_;
wire _31480_;
wire _31481_;
wire _31482_;
wire _31483_;
wire _31484_;
wire _31485_;
wire _31486_;
wire _31487_;
wire _31488_;
wire _31489_;
wire _31490_;
wire _31491_;
wire _31492_;
wire _31493_;
wire _31494_;
wire _31495_;
wire _31496_;
wire _31497_;
wire _31498_;
wire _31499_;
wire _31500_;
wire _31501_;
wire _31502_;
wire _31503_;
wire _31504_;
wire _31505_;
wire _31506_;
wire _31507_;
wire _31508_;
wire _31509_;
wire _31510_;
wire _31511_;
wire _31512_;
wire _31513_;
wire _31514_;
wire _31515_;
wire _31516_;
wire _31517_;
wire _31518_;
wire _31519_;
wire _31520_;
wire _31521_;
wire _31522_;
wire _31523_;
wire _31524_;
wire _31525_;
wire _31526_;
wire _31527_;
wire _31528_;
wire _31529_;
wire _31530_;
wire _31531_;
wire _31532_;
wire _31533_;
wire _31534_;
wire _31535_;
wire _31536_;
wire _31537_;
wire _31538_;
wire _31539_;
wire _31540_;
wire _31541_;
wire _31542_;
wire _31543_;
wire _31544_;
wire _31545_;
wire _31546_;
wire _31547_;
wire _31548_;
wire _31549_;
wire _31550_;
wire _31551_;
wire _31552_;
wire _31553_;
wire _31554_;
wire _31555_;
wire _31556_;
wire _31557_;
wire _31558_;
wire _31559_;
wire _31560_;
wire _31561_;
wire _31562_;
wire _31563_;
wire _31564_;
wire _31565_;
wire _31566_;
wire _31567_;
wire _31568_;
wire _31569_;
wire _31570_;
wire _31571_;
wire _31572_;
wire _31573_;
wire _31574_;
wire _31575_;
wire _31576_;
wire _31577_;
wire _31578_;
wire _31579_;
wire _31580_;
wire _31581_;
wire _31582_;
wire _31583_;
wire _31584_;
wire _31585_;
wire _31586_;
wire _31587_;
wire _31588_;
wire _31589_;
wire _31590_;
wire _31591_;
wire _31592_;
wire _31593_;
wire _31594_;
wire _31595_;
wire _31596_;
wire _31597_;
wire _31598_;
wire _31599_;
wire _31600_;
wire _31601_;
wire _31602_;
wire _31603_;
wire _31604_;
wire _31605_;
wire _31606_;
wire _31607_;
wire _31608_;
wire _31609_;
wire _31610_;
wire _31611_;
wire _31612_;
wire _31613_;
wire _31614_;
wire _31615_;
wire _31616_;
wire _31617_;
wire _31618_;
wire _31619_;
wire _31620_;
wire _31621_;
wire _31622_;
wire _31623_;
wire _31624_;
wire _31625_;
wire _31626_;
wire _31627_;
wire _31628_;
wire _31629_;
wire _31630_;
wire _31631_;
wire _31632_;
wire _31633_;
wire _31634_;
wire _31635_;
wire _31636_;
wire _31637_;
wire _31638_;
wire _31639_;
wire _31640_;
wire _31641_;
wire _31642_;
wire _31643_;
wire _31644_;
wire _31645_;
wire _31646_;
wire _31647_;
wire _31648_;
wire _31649_;
wire _31650_;
wire _31651_;
wire _31652_;
wire _31653_;
wire _31654_;
wire _31655_;
wire _31656_;
wire _31657_;
wire _31658_;
wire _31659_;
wire _31660_;
wire _31661_;
wire _31662_;
wire _31663_;
wire _31664_;
wire _31665_;
wire _31666_;
wire _31667_;
wire _31668_;
wire _31669_;
wire _31670_;
wire _31671_;
wire _31672_;
wire _31673_;
wire _31674_;
wire _31675_;
wire _31676_;
wire _31677_;
wire _31678_;
wire _31679_;
wire _31680_;
wire _31681_;
wire _31682_;
wire _31683_;
wire _31684_;
wire _31685_;
wire _31686_;
wire _31687_;
wire _31688_;
wire _31689_;
wire _31690_;
wire _31691_;
wire _31692_;
wire _31693_;
wire _31694_;
wire _31695_;
wire _31696_;
wire _31697_;
wire _31698_;
wire _31699_;
wire _31700_;
wire _31701_;
wire _31702_;
wire _31703_;
wire _31704_;
wire _31705_;
wire _31706_;
wire _31707_;
wire _31708_;
wire _31709_;
wire _31710_;
wire _31711_;
wire _31712_;
wire _31713_;
wire _31714_;
wire _31715_;
wire _31716_;
wire _31717_;
wire _31718_;
wire _31719_;
wire _31720_;
wire _31721_;
wire _31722_;
wire _31723_;
wire _31724_;
wire _31725_;
wire _31726_;
wire _31727_;
wire _31728_;
wire _31729_;
wire _31730_;
wire _31731_;
wire _31732_;
wire _31733_;
wire _31734_;
wire _31735_;
wire _31736_;
wire _31737_;
wire _31738_;
wire _31739_;
wire _31740_;
wire _31741_;
wire _31742_;
wire _31743_;
wire _31744_;
wire _31745_;
wire _31746_;
wire _31747_;
wire _31748_;
wire _31749_;
wire _31750_;
wire _31751_;
wire _31752_;
wire _31753_;
wire _31754_;
wire _31755_;
wire _31756_;
wire _31757_;
wire _31758_;
wire _31759_;
wire _31760_;
wire _31761_;
wire _31762_;
wire _31763_;
wire _31764_;
wire _31765_;
wire _31766_;
wire _31767_;
wire _31768_;
wire _31769_;
wire _31770_;
wire _31771_;
wire _31772_;
wire _31773_;
wire _31774_;
wire _31775_;
wire _31776_;
wire _31777_;
wire _31778_;
wire _31779_;
wire _31780_;
wire _31781_;
wire _31782_;
wire _31783_;
wire _31784_;
wire _31785_;
wire _31786_;
wire _31787_;
wire _31788_;
wire _31789_;
wire _31790_;
wire _31791_;
wire _31792_;
wire _31793_;
wire _31794_;
wire _31795_;
wire _31796_;
wire _31797_;
wire _31798_;
wire _31799_;
wire _31800_;
wire _31801_;
wire _31802_;
wire _31803_;
wire _31804_;
wire _31805_;
wire _31806_;
wire _31807_;
wire _31808_;
wire _31809_;
wire _31810_;
wire _31811_;
wire _31812_;
wire _31813_;
wire _31814_;
wire _31815_;
wire _31816_;
wire _31817_;
wire _31818_;
wire _31819_;
wire _31820_;
wire _31821_;
wire _31822_;
wire _31823_;
wire _31824_;
wire _31825_;
wire _31826_;
wire _31827_;
wire _31828_;
wire _31829_;
wire _31830_;
wire _31831_;
wire _31832_;
wire _31833_;
wire _31834_;
wire _31835_;
wire _31836_;
wire _31837_;
wire _31838_;
wire _31839_;
wire _31840_;
wire _31841_;
wire _31842_;
wire _31843_;
wire _31844_;
wire _31845_;
wire _31846_;
wire _31847_;
wire _31848_;
wire _31849_;
wire _31850_;
wire _31851_;
wire _31852_;
wire _31853_;
wire _31854_;
wire _31855_;
wire _31856_;
wire _31857_;
wire _31858_;
wire _31859_;
wire _31860_;
wire _31861_;
wire _31862_;
wire _31863_;
wire _31864_;
wire _31865_;
wire _31866_;
wire _31867_;
wire _31868_;
wire _31869_;
wire _31870_;
wire _31871_;
wire _31872_;
wire _31873_;
wire _31874_;
wire _31875_;
wire _31876_;
wire _31877_;
wire _31878_;
wire _31879_;
wire _31880_;
wire _31881_;
wire _31882_;
wire _31883_;
wire _31884_;
wire _31885_;
wire _31886_;
wire _31887_;
wire _31888_;
wire _31889_;
wire _31890_;
wire _31891_;
wire _31892_;
wire _31893_;
wire _31894_;
wire _31895_;
wire _31896_;
wire _31897_;
wire _31898_;
wire _31899_;
wire _31900_;
wire _31901_;
wire _31902_;
wire _31903_;
wire _31904_;
wire _31905_;
wire _31906_;
wire _31907_;
wire _31908_;
wire _31909_;
wire _31910_;
wire _31911_;
wire _31912_;
wire _31913_;
wire _31914_;
wire _31915_;
wire _31916_;
wire _31917_;
wire _31918_;
wire _31919_;
wire _31920_;
wire _31921_;
wire _31922_;
wire _31923_;
wire _31924_;
wire _31925_;
wire _31926_;
wire _31927_;
wire _31928_;
wire _31929_;
wire _31930_;
wire _31931_;
wire _31932_;
wire _31933_;
wire _31934_;
wire _31935_;
wire _31936_;
wire _31937_;
wire _31938_;
wire _31939_;
wire _31940_;
wire _31941_;
wire _31942_;
wire _31943_;
wire _31944_;
wire _31945_;
wire _31946_;
wire _31947_;
wire _31948_;
wire _31949_;
wire _31950_;
wire _31951_;
wire _31952_;
wire _31953_;
wire _31954_;
wire _31955_;
wire _31956_;
wire _31957_;
wire _31958_;
wire _31959_;
wire _31960_;
wire _31961_;
wire _31962_;
wire _31963_;
wire _31964_;
wire _31965_;
wire _31966_;
wire _31967_;
wire _31968_;
wire _31969_;
wire _31970_;
wire _31971_;
wire _31972_;
wire _31973_;
wire _31974_;
wire _31975_;
wire _31976_;
wire _31977_;
wire _31978_;
wire _31979_;
wire _31980_;
wire _31981_;
wire _31982_;
wire _31983_;
wire _31984_;
wire _31985_;
wire _31986_;
wire _31987_;
wire _31988_;
wire _31989_;
wire _31990_;
wire _31991_;
wire _31992_;
wire _31993_;
wire _31994_;
wire _31995_;
wire _31996_;
wire _31997_;
wire _31998_;
wire _31999_;
wire _32000_;
wire _32001_;
wire _32002_;
wire _32003_;
wire _32004_;
wire _32005_;
wire _32006_;
wire _32007_;
wire _32008_;
wire _32009_;
wire _32010_;
wire _32011_;
wire _32012_;
wire _32013_;
wire _32014_;
wire _32015_;
wire _32016_;
wire _32017_;
wire _32018_;
wire _32019_;
wire _32020_;
wire _32021_;
wire _32022_;
wire _32023_;
wire _32024_;
wire _32025_;
wire _32026_;
wire _32027_;
wire _32028_;
wire _32029_;
wire _32030_;
wire _32031_;
wire _32032_;
wire _32033_;
wire _32034_;
wire _32035_;
wire _32036_;
wire _32037_;
wire _32038_;
wire _32039_;
wire _32040_;
wire _32041_;
wire _32042_;
wire _32043_;
wire _32044_;
wire _32045_;
wire _32046_;
wire _32047_;
wire _32048_;
wire _32049_;
wire _32050_;
wire _32051_;
wire _32052_;
wire _32053_;
wire _32054_;
wire _32055_;
wire _32056_;
wire _32057_;
wire _32058_;
wire _32059_;
wire _32060_;
wire _32061_;
wire _32062_;
wire _32063_;
wire _32064_;
wire _32065_;
wire _32066_;
wire _32067_;
wire _32068_;
wire _32069_;
wire _32070_;
wire _32071_;
wire _32072_;
wire _32073_;
wire _32074_;
wire _32075_;
wire _32076_;
wire _32077_;
wire _32078_;
wire _32079_;
wire _32080_;
wire _32081_;
wire _32082_;
wire _32083_;
wire _32084_;
wire _32085_;
wire _32086_;
wire _32087_;
wire _32088_;
wire _32089_;
wire _32090_;
wire _32091_;
wire _32092_;
wire _32093_;
wire _32094_;
wire _32095_;
wire _32096_;
wire _32097_;
wire _32098_;
wire _32099_;
wire _32100_;
wire _32101_;
wire _32102_;
wire _32103_;
wire _32104_;
wire _32105_;
wire _32106_;
wire _32107_;
wire _32108_;
wire _32109_;
wire _32110_;
wire _32111_;
wire _32112_;
wire _32113_;
wire _32114_;
wire _32115_;
wire _32116_;
wire _32117_;
wire _32118_;
wire _32119_;
wire _32120_;
wire _32121_;
wire _32122_;
wire _32123_;
wire _32124_;
wire _32125_;
wire _32126_;
wire _32127_;
wire _32128_;
wire _32129_;
wire _32130_;
wire _32131_;
wire _32132_;
wire _32133_;
wire _32134_;
wire _32135_;
wire _32136_;
wire _32137_;
wire _32138_;
wire _32139_;
wire _32140_;
wire _32141_;
wire _32142_;
wire _32143_;
wire _32144_;
wire _32145_;
wire _32146_;
wire _32147_;
wire _32148_;
wire _32149_;
wire _32150_;
wire _32151_;
wire _32152_;
wire _32153_;
wire _32154_;
wire _32155_;
wire _32156_;
wire _32157_;
wire _32158_;
wire _32159_;
wire _32160_;
wire _32161_;
wire _32162_;
wire _32163_;
wire _32164_;
wire _32165_;
wire _32166_;
wire _32167_;
wire _32168_;
wire _32169_;
wire _32170_;
wire _32171_;
wire _32172_;
wire _32173_;
wire _32174_;
wire _32175_;
wire _32176_;
wire _32177_;
wire _32178_;
wire _32179_;
wire _32180_;
wire _32181_;
wire _32182_;
wire _32183_;
wire _32184_;
wire _32185_;
wire _32186_;
wire _32187_;
wire _32188_;
wire _32189_;
wire _32190_;
wire _32191_;
wire _32192_;
wire _32193_;
wire _32194_;
wire _32195_;
wire _32196_;
wire _32197_;
wire _32198_;
wire _32199_;
wire _32200_;
wire _32201_;
wire _32202_;
wire _32203_;
wire _32204_;
wire _32205_;
wire _32206_;
wire _32207_;
wire _32208_;
wire _32209_;
wire _32210_;
wire _32211_;
wire _32212_;
wire _32213_;
wire _32214_;
wire _32215_;
wire _32216_;
wire _32217_;
wire _32218_;
wire _32219_;
wire _32220_;
wire _32221_;
wire _32222_;
wire _32223_;
wire _32224_;
wire _32225_;
wire _32226_;
wire _32227_;
wire _32228_;
wire _32229_;
wire _32230_;
wire _32231_;
wire _32232_;
wire _32233_;
wire _32234_;
wire _32235_;
wire _32236_;
wire _32237_;
wire _32238_;
wire _32239_;
wire _32240_;
wire _32241_;
wire _32242_;
wire _32243_;
wire _32244_;
wire _32245_;
wire _32246_;
wire _32247_;
wire _32248_;
wire _32249_;
wire _32250_;
wire _32251_;
wire _32252_;
wire _32253_;
wire _32254_;
wire _32255_;
wire _32256_;
wire _32257_;
wire _32258_;
wire _32259_;
wire _32260_;
wire _32261_;
wire _32262_;
wire _32263_;
wire _32264_;
wire _32265_;
wire _32266_;
wire _32267_;
wire _32268_;
wire _32269_;
wire _32270_;
wire _32271_;
wire _32272_;
wire _32273_;
wire _32274_;
wire _32275_;
wire _32276_;
wire _32277_;
wire _32278_;
wire _32279_;
wire _32280_;
wire _32281_;
wire _32282_;
wire _32283_;
wire _32284_;
wire _32285_;
wire _32286_;
wire _32287_;
wire _32288_;
wire _32289_;
wire _32290_;
wire _32291_;
wire _32292_;
wire _32293_;
wire _32294_;
wire _32295_;
wire _32296_;
wire _32297_;
wire _32298_;
wire _32299_;
wire _32300_;
wire _32301_;
wire _32302_;
wire _32303_;
wire _32304_;
wire _32305_;
wire _32306_;
wire _32307_;
wire _32308_;
wire _32309_;
wire _32310_;
wire _32311_;
wire _32312_;
wire _32313_;
wire _32314_;
wire _32315_;
wire _32316_;
wire _32317_;
wire _32318_;
wire _32319_;
wire _32320_;
wire _32321_;
wire _32322_;
wire _32323_;
wire _32324_;
wire _32325_;
wire _32326_;
wire _32327_;
wire _32328_;
wire _32329_;
wire _32330_;
wire _32331_;
wire _32332_;
wire _32333_;
wire _32334_;
wire _32335_;
wire _32336_;
wire _32337_;
wire _32338_;
wire _32339_;
wire _32340_;
wire _32341_;
wire _32342_;
wire _32343_;
wire _32344_;
wire _32345_;
wire _32346_;
wire _32347_;
wire _32348_;
wire _32349_;
wire _32350_;
wire _32351_;
wire _32352_;
wire _32353_;
wire _32354_;
wire _32355_;
wire _32356_;
wire _32357_;
wire _32358_;
wire _32359_;
wire _32360_;
wire _32361_;
wire _32362_;
wire _32363_;
wire _32364_;
wire _32365_;
wire _32366_;
wire _32367_;
wire _32368_;
wire _32369_;
wire _32370_;
wire _32371_;
wire _32372_;
wire _32373_;
wire _32374_;
wire _32375_;
wire _32376_;
wire _32377_;
wire _32378_;
wire _32379_;
wire _32380_;
wire _32381_;
wire _32382_;
wire _32383_;
wire _32384_;
wire _32385_;
wire _32386_;
wire _32387_;
wire _32388_;
wire _32389_;
wire _32390_;
wire _32391_;
wire _32392_;
wire _32393_;
wire _32394_;
wire _32395_;
wire _32396_;
wire _32397_;
wire _32398_;
wire _32399_;
wire _32400_;
wire _32401_;
wire _32402_;
wire _32403_;
wire _32404_;
wire _32405_;
wire _32406_;
wire _32407_;
wire _32408_;
wire _32409_;
wire _32410_;
wire _32411_;
wire _32412_;
wire _32413_;
wire _32414_;
wire _32415_;
wire _32416_;
wire _32417_;
wire _32418_;
wire _32419_;
wire _32420_;
wire _32421_;
wire _32422_;
wire _32423_;
wire _32424_;
wire _32425_;
wire _32426_;
wire _32427_;
wire _32428_;
wire _32429_;
wire _32430_;
wire _32431_;
wire _32432_;
wire _32433_;
wire _32434_;
wire _32435_;
wire _32436_;
wire _32437_;
wire _32438_;
wire _32439_;
wire _32440_;
wire _32441_;
wire _32442_;
wire _32443_;
wire _32444_;
wire _32445_;
wire _32446_;
wire _32447_;
wire _32448_;
wire _32449_;
wire _32450_;
wire _32451_;
wire _32452_;
wire _32453_;
wire _32454_;
wire _32455_;
wire _32456_;
wire _32457_;
wire _32458_;
wire _32459_;
wire _32460_;
wire _32461_;
wire _32462_;
wire _32463_;
wire _32464_;
wire _32465_;
wire _32466_;
wire _32467_;
wire _32468_;
wire _32469_;
wire _32470_;
wire _32471_;
wire _32472_;
wire _32473_;
wire _32474_;
wire _32475_;
wire _32476_;
wire _32477_;
wire _32478_;
wire _32479_;
wire _32480_;
wire _32481_;
wire _32482_;
wire _32483_;
wire _32484_;
wire _32485_;
wire _32486_;
wire _32487_;
wire _32488_;
wire _32489_;
wire _32490_;
wire _32491_;
wire _32492_;
wire _32493_;
wire _32494_;
wire _32495_;
wire _32496_;
wire _32497_;
wire _32498_;
wire _32499_;
wire _32500_;
wire _32501_;
wire _32502_;
wire _32503_;
wire _32504_;
wire _32505_;
wire _32506_;
wire _32507_;
wire _32508_;
wire _32509_;
wire _32510_;
wire _32511_;
wire _32512_;
wire _32513_;
wire _32514_;
wire _32515_;
wire _32516_;
wire _32517_;
wire _32518_;
wire _32519_;
wire _32520_;
wire _32521_;
wire _32522_;
wire _32523_;
wire _32524_;
wire _32525_;
wire _32526_;
wire _32527_;
wire _32528_;
wire _32529_;
wire _32530_;
wire _32531_;
wire _32532_;
wire _32533_;
wire _32534_;
wire _32535_;
wire _32536_;
wire _32537_;
wire _32538_;
wire _32539_;
wire _32540_;
wire _32541_;
wire _32542_;
wire _32543_;
wire _32544_;
wire _32545_;
wire _32546_;
wire _32547_;
wire _32548_;
wire _32549_;
wire _32550_;
wire _32551_;
wire _32552_;
wire _32553_;
wire _32554_;
wire _32555_;
wire _32556_;
wire _32557_;
wire _32558_;
wire _32559_;
wire _32560_;
wire _32561_;
wire _32562_;
wire _32563_;
wire _32564_;
wire _32565_;
wire _32566_;
wire _32567_;
wire _32568_;
wire _32569_;
wire _32570_;
wire _32571_;
wire _32572_;
wire _32573_;
wire _32574_;
wire _32575_;
wire _32576_;
wire _32577_;
wire _32578_;
wire _32579_;
wire _32580_;
wire _32581_;
wire _32582_;
wire _32583_;
wire _32584_;
wire _32585_;
wire _32586_;
wire _32587_;
wire _32588_;
wire _32589_;
wire _32590_;
wire _32591_;
wire _32592_;
wire _32593_;
wire _32594_;
wire _32595_;
wire _32596_;
wire _32597_;
wire _32598_;
wire _32599_;
wire _32600_;
wire _32601_;
wire _32602_;
wire _32603_;
wire _32604_;
wire _32605_;
wire _32606_;
wire _32607_;
wire _32608_;
wire _32609_;
wire _32610_;
wire _32611_;
wire _32612_;
wire _32613_;
wire _32614_;
wire _32615_;
wire _32616_;
wire _32617_;
wire _32618_;
wire _32619_;
wire _32620_;
wire _32621_;
wire _32622_;
wire _32623_;
wire _32624_;
wire _32625_;
wire _32626_;
wire _32627_;
wire _32628_;
wire _32629_;
wire _32630_;
wire _32631_;
wire _32632_;
wire _32633_;
wire _32634_;
wire _32635_;
wire _32636_;
wire _32637_;
wire _32638_;
wire _32639_;
wire _32640_;
wire _32641_;
wire _32642_;
wire _32643_;
wire _32644_;
wire _32645_;
wire _32646_;
wire _32647_;
wire _32648_;
wire _32649_;
wire _32650_;
wire _32651_;
wire _32652_;
wire _32653_;
wire _32654_;
wire _32655_;
wire _32656_;
wire _32657_;
wire _32658_;
wire _32659_;
wire _32660_;
wire _32661_;
wire _32662_;
wire _32663_;
wire _32664_;
wire _32665_;
wire _32666_;
wire _32667_;
wire _32668_;
wire _32669_;
wire _32670_;
wire _32671_;
wire _32672_;
wire _32673_;
wire _32674_;
wire _32675_;
wire _32676_;
wire _32677_;
wire _32678_;
wire _32679_;
wire _32680_;
wire _32681_;
wire _32682_;
wire _32683_;
wire _32684_;
wire _32685_;
wire _32686_;
wire _32687_;
wire _32688_;
wire _32689_;
wire _32690_;
wire _32691_;
wire _32692_;
wire _32693_;
wire _32694_;
wire _32695_;
wire _32696_;
wire _32697_;
wire _32698_;
wire _32699_;
wire _32700_;
wire _32701_;
wire _32702_;
wire _32703_;
wire _32704_;
wire _32705_;
wire _32706_;
wire _32707_;
wire _32708_;
wire _32709_;
wire _32710_;
wire _32711_;
wire _32712_;
wire _32713_;
wire _32714_;
wire _32715_;
wire _32716_;
wire _32717_;
wire _32718_;
wire _32719_;
wire _32720_;
wire _32721_;
wire _32722_;
wire _32723_;
wire _32724_;
wire _32725_;
wire _32726_;
wire _32727_;
wire _32728_;
wire _32729_;
wire _32730_;
wire _32731_;
wire _32732_;
wire _32733_;
wire _32734_;
wire _32735_;
wire _32736_;
wire _32737_;
wire _32738_;
wire _32739_;
wire _32740_;
wire _32741_;
wire _32742_;
wire _32743_;
wire _32744_;
wire _32745_;
wire _32746_;
wire _32747_;
wire _32748_;
wire _32749_;
wire _32750_;
wire _32751_;
wire _32752_;
wire _32753_;
wire _32754_;
wire _32755_;
wire _32756_;
wire _32757_;
wire _32758_;
wire _32759_;
wire _32760_;
wire _32761_;
wire _32762_;
wire _32763_;
wire _32764_;
wire _32765_;
wire _32766_;
wire _32767_;
wire _32768_;
wire _32769_;
wire _32770_;
wire _32771_;
wire _32772_;
wire _32773_;
wire _32774_;
wire _32775_;
wire _32776_;
wire _32777_;
wire _32778_;
wire _32779_;
wire _32780_;
wire _32781_;
wire _32782_;
wire _32783_;
wire _32784_;
wire _32785_;
wire _32786_;
wire _32787_;
wire _32788_;
wire _32789_;
wire _32790_;
wire _32791_;
wire _32792_;
wire _32793_;
wire _32794_;
wire _32795_;
wire _32796_;
wire _32797_;
wire _32798_;
wire _32799_;
wire _32800_;
wire _32801_;
wire _32802_;
wire _32803_;
wire _32804_;
wire _32805_;
wire _32806_;
wire _32807_;
wire _32808_;
wire _32809_;
wire _32810_;
wire _32811_;
wire _32812_;
wire _32813_;
wire _32814_;
wire _32815_;
wire _32816_;
wire _32817_;
wire _32818_;
wire _32819_;
wire _32820_;
wire _32821_;
wire _32822_;
wire _32823_;
wire _32824_;
wire _32825_;
wire _32826_;
wire _32827_;
wire _32828_;
wire _32829_;
wire _32830_;
wire _32831_;
wire _32832_;
wire _32833_;
wire _32834_;
wire _32835_;
wire _32836_;
wire _32837_;
wire _32838_;
wire _32839_;
wire _32840_;
wire _32841_;
wire _32842_;
wire _32843_;
wire _32844_;
wire _32845_;
wire _32846_;
wire _32847_;
wire _32848_;
wire _32849_;
wire _32850_;
wire _32851_;
wire _32852_;
wire _32853_;
wire _32854_;
wire _32855_;
wire _32856_;
wire _32857_;
wire _32858_;
wire _32859_;
wire _32860_;
wire _32861_;
wire _32862_;
wire _32863_;
wire _32864_;
wire _32865_;
wire _32866_;
wire _32867_;
wire _32868_;
wire _32869_;
wire _32870_;
wire _32871_;
wire _32872_;
wire _32873_;
wire _32874_;
wire _32875_;
wire _32876_;
wire _32877_;
wire _32878_;
wire _32879_;
wire _32880_;
wire _32881_;
wire _32882_;
wire _32883_;
wire _32884_;
wire _32885_;
wire _32886_;
wire _32887_;
wire _32888_;
wire _32889_;
wire _32890_;
wire _32891_;
wire _32892_;
wire _32893_;
wire _32894_;
wire _32895_;
wire _32896_;
wire _32897_;
wire _32898_;
wire _32899_;
wire _32900_;
wire _32901_;
wire _32902_;
wire _32903_;
wire _32904_;
wire _32905_;
wire _32906_;
wire _32907_;
wire _32908_;
wire _32909_;
wire _32910_;
wire _32911_;
wire _32912_;
wire _32913_;
wire _32914_;
wire _32915_;
wire _32916_;
wire _32917_;
wire _32918_;
wire _32919_;
wire _32920_;
wire _32921_;
wire _32922_;
wire _32923_;
wire _32924_;
wire _32925_;
wire _32926_;
wire _32927_;
wire _32928_;
wire _32929_;
wire _32930_;
wire _32931_;
wire _32932_;
wire _32933_;
wire _32934_;
wire _32935_;
wire _32936_;
wire _32937_;
wire _32938_;
wire _32939_;
wire _32940_;
wire _32941_;
wire _32942_;
wire _32943_;
wire _32944_;
wire _32945_;
wire _32946_;
wire _32947_;
wire _32948_;
wire _32949_;
wire _32950_;
wire _32951_;
wire _32952_;
wire _32953_;
wire _32954_;
wire _32955_;
wire _32956_;
wire _32957_;
wire _32958_;
wire _32959_;
wire _32960_;
wire _32961_;
wire _32962_;
wire _32963_;
wire _32964_;
wire _32965_;
wire _32966_;
wire _32967_;
wire _32968_;
wire _32969_;
wire _32970_;
wire _32971_;
wire _32972_;
wire _32973_;
wire _32974_;
wire _32975_;
wire _32976_;
wire _32977_;
wire _32978_;
wire _32979_;
wire _32980_;
wire _32981_;
wire _32982_;
wire _32983_;
wire _32984_;
wire _32985_;
wire _32986_;
wire _32987_;
wire _32988_;
wire _32989_;
wire _32990_;
wire _32991_;
wire _32992_;
wire _32993_;
wire _32994_;
wire _32995_;
wire _32996_;
wire _32997_;
wire _32998_;
wire _32999_;
wire _33000_;
wire _33001_;
wire _33002_;
wire _33003_;
wire _33004_;
wire _33005_;
wire _33006_;
wire _33007_;
wire _33008_;
wire _33009_;
wire _33010_;
wire _33011_;
wire _33012_;
wire _33013_;
wire _33014_;
wire _33015_;
wire _33016_;
wire _33017_;
wire _33018_;
wire _33019_;
wire _33020_;
wire _33021_;
wire _33022_;
wire _33023_;
wire _33024_;
wire _33025_;
wire _33026_;
wire _33027_;
wire _33028_;
wire _33029_;
wire _33030_;
wire _33031_;
wire _33032_;
wire _33033_;
wire _33034_;
wire _33035_;
wire _33036_;
wire _33037_;
wire _33038_;
wire _33039_;
wire _33040_;
wire _33041_;
wire _33042_;
wire _33043_;
wire _33044_;
wire _33045_;
wire _33046_;
wire _33047_;
wire _33048_;
wire _33049_;
wire _33050_;
wire _33051_;
wire _33052_;
wire _33053_;
wire _33054_;
wire _33055_;
wire _33056_;
wire _33057_;
wire _33058_;
wire _33059_;
wire _33060_;
wire _33061_;
wire _33062_;
wire _33063_;
wire _33064_;
wire _33065_;
wire _33066_;
wire _33067_;
wire _33068_;
wire _33069_;
wire _33070_;
wire _33071_;
wire _33072_;
wire _33073_;
wire _33074_;
wire _33075_;
wire _33076_;
wire _33077_;
wire _33078_;
wire _33079_;
wire _33080_;
wire _33081_;
wire _33082_;
wire _33083_;
wire _33084_;
wire _33085_;
wire _33086_;
wire _33087_;
wire _33088_;
wire _33089_;
wire _33090_;
wire _33091_;
wire _33092_;
wire _33093_;
wire _33094_;
wire _33095_;
wire _33096_;
wire _33097_;
wire _33098_;
wire _33099_;
wire _33100_;
wire _33101_;
wire _33102_;
wire _33103_;
wire _33104_;
wire _33105_;
wire _33106_;
wire _33107_;
wire _33108_;
wire _33109_;
wire _33110_;
wire _33111_;
wire _33112_;
wire _33113_;
wire _33114_;
wire _33115_;
wire _33116_;
wire _33117_;
wire _33118_;
wire _33119_;
wire _33120_;
wire _33121_;
wire _33122_;
wire _33123_;
wire _33124_;
wire _33125_;
wire _33126_;
wire _33127_;
wire _33128_;
wire _33129_;
wire _33130_;
wire _33131_;
wire _33132_;
wire _33133_;
wire _33134_;
wire _33135_;
wire _33136_;
wire _33137_;
wire _33138_;
wire _33139_;
wire _33140_;
wire _33141_;
wire _33142_;
wire _33143_;
wire _33144_;
wire _33145_;
wire _33146_;
wire _33147_;
wire _33148_;
wire _33149_;
wire _33150_;
wire _33151_;
wire _33152_;
wire _33153_;
wire _33154_;
wire _33155_;
wire _33156_;
wire _33157_;
wire _33158_;
wire _33159_;
wire _33160_;
wire _33161_;
wire _33162_;
wire _33163_;
wire _33164_;
wire _33165_;
wire _33166_;
wire _33167_;
wire _33168_;
wire _33169_;
wire _33170_;
wire _33171_;
wire _33172_;
wire _33173_;
wire _33174_;
wire _33175_;
wire _33176_;
wire _33177_;
wire _33178_;
wire _33179_;
wire _33180_;
wire _33181_;
wire _33182_;
wire _33183_;
wire _33184_;
wire _33185_;
wire _33186_;
wire _33187_;
wire _33188_;
wire _33189_;
wire _33190_;
wire _33191_;
wire _33192_;
wire _33193_;
wire _33194_;
wire _33195_;
wire _33196_;
wire _33197_;
wire _33198_;
wire _33199_;
wire _33200_;
wire _33201_;
wire _33202_;
wire _33203_;
wire _33204_;
wire _33205_;
wire _33206_;
wire _33207_;
wire _33208_;
wire _33209_;
wire _33210_;
wire _33211_;
wire _33212_;
wire _33213_;
wire _33214_;
wire _33215_;
wire _33216_;
wire _33217_;
wire _33218_;
wire _33219_;
wire _33220_;
wire _33221_;
wire _33222_;
wire _33223_;
wire _33224_;
wire _33225_;
wire _33226_;
wire _33227_;
wire _33228_;
wire _33229_;
wire _33230_;
wire _33231_;
wire _33232_;
wire _33233_;
wire _33234_;
wire _33235_;
wire _33236_;
wire _33237_;
wire _33238_;
wire _33239_;
wire _33240_;
wire _33241_;
wire _33242_;
wire _33243_;
wire _33244_;
wire _33245_;
wire _33246_;
wire _33247_;
wire _33248_;
wire _33249_;
wire _33250_;
wire _33251_;
wire _33252_;
wire _33253_;
wire _33254_;
wire _33255_;
wire _33256_;
wire _33257_;
wire _33258_;
wire _33259_;
wire _33260_;
wire _33261_;
wire _33262_;
wire _33263_;
wire _33264_;
wire _33265_;
wire _33266_;
wire _33267_;
wire _33268_;
wire _33269_;
wire _33270_;
wire _33271_;
wire _33272_;
wire _33273_;
wire _33274_;
wire _33275_;
wire _33276_;
wire _33277_;
wire _33278_;
wire _33279_;
wire _33280_;
wire _33281_;
wire _33282_;
wire _33283_;
wire _33284_;
wire _33285_;
wire _33286_;
wire _33287_;
wire _33288_;
wire _33289_;
wire _33290_;
wire _33291_;
wire _33292_;
wire _33293_;
wire _33294_;
wire _33295_;
wire _33296_;
wire _33297_;
wire _33298_;
wire _33299_;
wire _33300_;
wire _33301_;
wire _33302_;
wire _33303_;
wire _33304_;
wire _33305_;
wire _33306_;
wire _33307_;
wire _33308_;
wire _33309_;
wire _33310_;
wire _33311_;
wire _33312_;
wire _33313_;
wire _33314_;
wire _33315_;
wire _33316_;
wire _33317_;
wire _33318_;
wire _33319_;
wire _33320_;
wire _33321_;
wire _33322_;
wire _33323_;
wire _33324_;
wire _33325_;
wire _33326_;
wire _33327_;
wire _33328_;
wire _33329_;
wire _33330_;
wire _33331_;
wire _33332_;
wire _33333_;
wire _33334_;
wire _33335_;
wire _33336_;
wire _33337_;
wire _33338_;
wire _33339_;
wire _33340_;
wire _33341_;
wire _33342_;
wire _33343_;
wire _33344_;
wire _33345_;
wire _33346_;
wire _33347_;
wire _33348_;
wire _33349_;
wire _33350_;
wire _33351_;
wire _33352_;
wire _33353_;
wire _33354_;
wire _33355_;
wire _33356_;
wire _33357_;
wire _33358_;
wire _33359_;
wire _33360_;
wire _33361_;
wire _33362_;
wire _33363_;
wire _33364_;
wire _33365_;
wire _33366_;
wire _33367_;
wire _33368_;
wire _33369_;
wire _33370_;
wire _33371_;
wire _33372_;
wire _33373_;
wire _33374_;
wire _33375_;
wire _33376_;
wire _33377_;
wire _33378_;
wire _33379_;
wire _33380_;
wire _33381_;
wire _33382_;
wire _33383_;
wire _33384_;
wire _33385_;
wire _33386_;
wire _33387_;
wire _33388_;
wire _33389_;
wire _33390_;
wire _33391_;
wire _33392_;
wire _33393_;
wire _33394_;
wire _33395_;
wire _33396_;
wire _33397_;
wire _33398_;
wire _33399_;
wire _33400_;
wire _33401_;
wire _33402_;
wire _33403_;
wire _33404_;
wire _33405_;
wire _33406_;
wire _33407_;
wire _33408_;
wire _33409_;
wire _33410_;
wire _33411_;
wire _33412_;
wire _33413_;
wire _33414_;
wire _33415_;
wire _33416_;
wire _33417_;
wire _33418_;
wire _33419_;
wire _33420_;
wire _33421_;
wire _33422_;
wire _33423_;
wire _33424_;
wire _33425_;
wire _33426_;
wire _33427_;
wire _33428_;
wire _33429_;
wire _33430_;
wire _33431_;
wire _33432_;
wire _33433_;
wire _33434_;
wire _33435_;
wire _33436_;
wire _33437_;
wire _33438_;
wire _33439_;
wire _33440_;
wire _33441_;
wire _33442_;
wire _33443_;
wire _33444_;
wire _33445_;
wire _33446_;
wire _33447_;
wire _33448_;
wire _33449_;
wire _33450_;
wire _33451_;
wire _33452_;
wire _33453_;
wire _33454_;
wire _33455_;
wire _33456_;
wire _33457_;
wire _33458_;
wire _33459_;
wire _33460_;
wire _33461_;
wire _33462_;
wire _33463_;
wire _33464_;
wire _33465_;
wire _33466_;
wire _33467_;
wire _33468_;
wire _33469_;
wire _33470_;
wire _33471_;
wire _33472_;
wire _33473_;
wire _33474_;
wire _33475_;
wire _33476_;
wire _33477_;
wire _33478_;
wire _33479_;
wire _33480_;
wire _33481_;
wire _33482_;
wire _33483_;
wire _33484_;
wire _33485_;
wire _33486_;
wire _33487_;
wire _33488_;
wire _33489_;
wire _33490_;
wire _33491_;
wire _33492_;
wire _33493_;
wire _33494_;
wire _33495_;
wire _33496_;
wire _33497_;
wire _33498_;
wire _33499_;
wire _33500_;
wire _33501_;
wire _33502_;
wire _33503_;
wire _33504_;
wire _33505_;
wire _33506_;
wire _33507_;
wire _33508_;
wire _33509_;
wire _33510_;
wire _33511_;
wire _33512_;
wire _33513_;
wire _33514_;
wire _33515_;
wire _33516_;
wire _33517_;
wire _33518_;
wire _33519_;
wire _33520_;
wire _33521_;
wire _33522_;
wire _33523_;
wire _33524_;
wire _33525_;
wire _33526_;
wire _33527_;
wire _33528_;
wire _33529_;
wire _33530_;
wire _33531_;
wire _33532_;
wire _33533_;
wire _33534_;
wire _33535_;
wire _33536_;
wire _33537_;
wire _33538_;
wire _33539_;
wire _33540_;
wire _33541_;
wire _33542_;
wire _33543_;
wire _33544_;
wire _33545_;
wire _33546_;
wire _33547_;
wire _33548_;
wire _33549_;
wire _33550_;
wire _33551_;
wire _33552_;
wire _33553_;
wire _33554_;
wire _33555_;
wire _33556_;
wire _33557_;
wire _33558_;
wire _33559_;
wire _33560_;
wire _33561_;
wire _33562_;
wire _33563_;
wire _33564_;
wire _33565_;
wire _33566_;
wire _33567_;
wire _33568_;
wire _33569_;
wire _33570_;
wire _33571_;
wire _33572_;
wire _33573_;
wire _33574_;
wire _33575_;
wire _33576_;
wire _33577_;
wire _33578_;
wire _33579_;
wire _33580_;
wire _33581_;
wire _33582_;
wire _33583_;
wire _33584_;
wire _33585_;
wire _33586_;
wire _33587_;
wire _33588_;
wire _33589_;
wire _33590_;
wire _33591_;
wire _33592_;
wire _33593_;
wire _33594_;
wire _33595_;
wire _33596_;
wire _33597_;
wire _33598_;
wire _33599_;
wire _33600_;
wire _33601_;
wire _33602_;
wire _33603_;
wire _33604_;
wire _33605_;
wire _33606_;
wire _33607_;
wire _33608_;
wire _33609_;
wire _33610_;
wire _33611_;
wire _33612_;
wire _33613_;
wire _33614_;
wire _33615_;
wire _33616_;
wire _33617_;
wire _33618_;
wire _33619_;
wire _33620_;
wire _33621_;
wire _33622_;
wire _33623_;
wire _33624_;
wire _33625_;
wire _33626_;
wire _33627_;
wire _33628_;
wire _33629_;
wire _33630_;
wire _33631_;
wire _33632_;
wire _33633_;
wire _33634_;
wire _33635_;
wire _33636_;
wire _33637_;
wire _33638_;
wire _33639_;
wire _33640_;
wire _33641_;
wire _33642_;
wire _33643_;
wire _33644_;
wire _33645_;
wire _33646_;
wire _33647_;
wire _33648_;
wire _33649_;
wire _33650_;
wire _33651_;
wire _33652_;
wire _33653_;
wire _33654_;
wire _33655_;
wire _33656_;
wire _33657_;
wire _33658_;
wire _33659_;
wire _33660_;
wire _33661_;
wire _33662_;
wire _33663_;
wire _33664_;
wire _33665_;
wire _33666_;
wire _33667_;
wire _33668_;
wire _33669_;
wire _33670_;
wire _33671_;
wire _33672_;
wire _33673_;
wire _33674_;
wire _33675_;
wire _33676_;
wire _33677_;
wire _33678_;
wire _33679_;
wire _33680_;
wire _33681_;
wire _33682_;
wire _33683_;
wire _33684_;
wire _33685_;
wire _33686_;
wire _33687_;
wire _33688_;
wire _33689_;
wire _33690_;
wire _33691_;
wire _33692_;
wire _33693_;
wire _33694_;
wire _33695_;
wire _33696_;
wire _33697_;
wire _33698_;
wire _33699_;
wire _33700_;
wire _33701_;
wire _33702_;
wire _33703_;
wire _33704_;
wire _33705_;
wire _33706_;
wire _33707_;
wire _33708_;
wire _33709_;
wire _33710_;
wire _33711_;
wire _33712_;
wire _33713_;
wire _33714_;
wire _33715_;
wire _33716_;
wire _33717_;
wire _33718_;
wire _33719_;
wire _33720_;
wire _33721_;
wire _33722_;
wire _33723_;
wire _33724_;
wire _33725_;
wire _33726_;
wire _33727_;
wire _33728_;
wire _33729_;
wire _33730_;
wire _33731_;
wire _33732_;
wire _33733_;
wire _33734_;
wire _33735_;
wire _33736_;
wire _33737_;
wire _33738_;
wire _33739_;
wire _33740_;
wire _33741_;
wire _33742_;
wire _33743_;
wire _33744_;
wire _33745_;
wire _33746_;
wire _33747_;
wire _33748_;
wire _33749_;
wire _33750_;
wire _33751_;
wire _33752_;
wire _33753_;
wire _33754_;
wire _33755_;
wire _33756_;
wire _33757_;
wire _33758_;
wire _33759_;
wire _33760_;
wire _33761_;
wire _33762_;
wire _33763_;
wire _33764_;
wire _33765_;
wire _33766_;
wire _33767_;
wire _33768_;
wire _33769_;
wire _33770_;
wire _33771_;
wire _33772_;
wire _33773_;
wire _33774_;
wire _33775_;
wire _33776_;
wire _33777_;
wire _33778_;
wire _33779_;
wire _33780_;
wire _33781_;
wire _33782_;
wire _33783_;
wire _33784_;
wire _33785_;
wire _33786_;
wire _33787_;
wire _33788_;
wire _33789_;
wire _33790_;
wire _33791_;
wire _33792_;
wire _33793_;
wire _33794_;
wire _33795_;
wire _33796_;
wire _33797_;
wire _33798_;
wire _33799_;
wire _33800_;
wire _33801_;
wire _33802_;
wire _33803_;
wire _33804_;
wire _33805_;
wire _33806_;
wire _33807_;
wire _33808_;
wire _33809_;
wire _33810_;
wire _33811_;
wire _33812_;
wire _33813_;
wire _33814_;
wire _33815_;
wire _33816_;
wire _33817_;
wire _33818_;
wire _33819_;
wire _33820_;
wire _33821_;
wire _33822_;
wire _33823_;
wire _33824_;
wire _33825_;
wire _33826_;
wire _33827_;
wire _33828_;
wire _33829_;
wire _33830_;
wire _33831_;
wire _33832_;
wire _33833_;
wire _33834_;
wire _33835_;
wire _33836_;
wire _33837_;
wire _33838_;
wire _33839_;
wire _33840_;
wire _33841_;
wire _33842_;
wire _33843_;
wire _33844_;
wire _33845_;
wire _33846_;
wire _33847_;
wire _33848_;
wire _33849_;
wire _33850_;
wire _33851_;
wire _33852_;
wire _33853_;
wire _33854_;
wire _33855_;
wire _33856_;
wire _33857_;
wire _33858_;
wire _33859_;
wire _33860_;
wire _33861_;
wire _33862_;
wire _33863_;
wire _33864_;
wire _33865_;
wire _33866_;
wire _33867_;
wire _33868_;
wire _33869_;
wire _33870_;
wire _33871_;
wire _33872_;
wire _33873_;
wire _33874_;
wire _33875_;
wire _33876_;
wire _33877_;
wire _33878_;
wire _33879_;
wire _33880_;
wire _33881_;
wire _33882_;
wire _33883_;
wire _33884_;
wire _33885_;
wire _33886_;
wire _33887_;
wire _33888_;
wire _33889_;
wire _33890_;
wire _33891_;
wire _33892_;
wire _33893_;
wire _33894_;
wire _33895_;
wire _33896_;
wire _33897_;
wire _33898_;
wire _33899_;
wire _33900_;
wire _33901_;
wire _33902_;
wire _33903_;
wire _33904_;
wire _33905_;
wire _33906_;
wire _33907_;
wire _33908_;
wire _33909_;
wire _33910_;
wire _33911_;
wire _33912_;
wire _33913_;
wire _33914_;
wire _33915_;
wire _33916_;
wire _33917_;
wire _33918_;
wire _33919_;
wire _33920_;
wire _33921_;
wire _33922_;
wire _33923_;
wire _33924_;
wire _33925_;
wire _33926_;
wire _33927_;
wire _33928_;
wire _33929_;
wire _33930_;
wire _33931_;
wire _33932_;
wire _33933_;
wire _33934_;
wire _33935_;
wire _33936_;
wire _33937_;
wire _33938_;
wire _33939_;
wire _33940_;
wire _33941_;
wire _33942_;
wire _33943_;
wire _33944_;
wire _33945_;
wire _33946_;
wire _33947_;
wire _33948_;
wire _33949_;
wire _33950_;
wire _33951_;
wire _33952_;
wire _33953_;
wire _33954_;
wire _33955_;
wire _33956_;
wire _33957_;
wire _33958_;
wire _33959_;
wire _33960_;
wire _33961_;
wire _33962_;
wire _33963_;
wire _33964_;
wire _33965_;
wire _33966_;
wire _33967_;
wire _33968_;
wire _33969_;
wire _33970_;
wire _33971_;
wire _33972_;
wire _33973_;
wire _33974_;
wire _33975_;
wire _33976_;
wire _33977_;
wire _33978_;
wire _33979_;
wire _33980_;
wire _33981_;
wire _33982_;
wire _33983_;
wire _33984_;
wire _33985_;
wire _33986_;
wire _33987_;
wire _33988_;
wire _33989_;
wire _33990_;
wire _33991_;
wire _33992_;
wire _33993_;
wire _33994_;
wire _33995_;
wire _33996_;
wire _33997_;
wire _33998_;
wire _33999_;
wire _34000_;
wire _34001_;
wire _34002_;
wire _34003_;
wire _34004_;
wire _34005_;
wire _34006_;
wire _34007_;
wire _34008_;
wire _34009_;
wire _34010_;
wire _34011_;
wire _34012_;
wire _34013_;
wire _34014_;
wire _34015_;
wire _34016_;
wire _34017_;
wire _34018_;
wire _34019_;
wire _34020_;
wire _34021_;
wire _34022_;
wire _34023_;
wire _34024_;
wire _34025_;
wire _34026_;
wire _34027_;
wire _34028_;
wire _34029_;
wire _34030_;
wire _34031_;
wire _34032_;
wire _34033_;
wire _34034_;
wire _34035_;
wire _34036_;
wire _34037_;
wire _34038_;
wire _34039_;
wire _34040_;
wire _34041_;
wire _34042_;
wire _34043_;
wire _34044_;
wire _34045_;
wire _34046_;
wire _34047_;
wire _34048_;
wire _34049_;
wire _34050_;
wire _34051_;
wire _34052_;
wire _34053_;
wire _34054_;
wire _34055_;
wire _34056_;
wire _34057_;
wire _34058_;
wire _34059_;
wire _34060_;
wire _34061_;
wire _34062_;
wire _34063_;
wire _34064_;
wire _34065_;
wire _34066_;
wire _34067_;
wire _34068_;
wire _34069_;
wire _34070_;
wire _34071_;
wire _34072_;
wire _34073_;
wire _34074_;
wire _34075_;
wire _34076_;
wire _34077_;
wire _34078_;
wire _34079_;
wire _34080_;
wire _34081_;
wire _34082_;
wire _34083_;
wire _34084_;
wire _34085_;
wire _34086_;
wire _34087_;
wire _34088_;
wire _34089_;
wire _34090_;
wire _34091_;
wire _34092_;
wire _34093_;
wire _34094_;
wire _34095_;
wire _34096_;
wire _34097_;
wire _34098_;
wire _34099_;
wire _34100_;
wire _34101_;
wire _34102_;
wire _34103_;
wire _34104_;
wire _34105_;
wire _34106_;
wire _34107_;
wire _34108_;
wire _34109_;
wire _34110_;
wire _34111_;
wire _34112_;
wire _34113_;
wire _34114_;
wire _34115_;
wire _34116_;
wire _34117_;
wire _34118_;
wire _34119_;
wire _34120_;
wire _34121_;
wire _34122_;
wire _34123_;
wire _34124_;
wire _34125_;
wire _34126_;
wire _34127_;
wire _34128_;
wire _34129_;
wire _34130_;
wire _34131_;
wire _34132_;
wire _34133_;
wire _34134_;
wire _34135_;
wire _34136_;
wire _34137_;
wire _34138_;
wire _34139_;
wire _34140_;
wire _34141_;
wire _34142_;
wire _34143_;
wire _34144_;
wire _34145_;
wire _34146_;
wire _34147_;
wire _34148_;
wire _34149_;
wire _34150_;
wire _34151_;
wire _34152_;
wire _34153_;
wire _34154_;
wire _34155_;
wire _34156_;
wire _34157_;
wire _34158_;
wire _34159_;
wire _34160_;
wire _34161_;
wire _34162_;
wire _34163_;
wire _34164_;
wire _34165_;
wire _34166_;
wire _34167_;
wire _34168_;
wire _34169_;
wire _34170_;
wire _34171_;
wire _34172_;
wire _34173_;
wire _34174_;
wire _34175_;
wire _34176_;
wire _34177_;
wire _34178_;
wire _34179_;
wire _34180_;
wire _34181_;
wire _34182_;
wire _34183_;
wire _34184_;
wire _34185_;
wire _34186_;
wire _34187_;
wire _34188_;
wire _34189_;
wire _34190_;
wire _34191_;
wire _34192_;
wire _34193_;
wire _34194_;
wire _34195_;
wire _34196_;
wire _34197_;
wire _34198_;
wire _34199_;
wire _34200_;
wire _34201_;
wire _34202_;
wire _34203_;
wire _34204_;
wire _34205_;
wire _34206_;
wire _34207_;
wire _34208_;
wire _34209_;
wire _34210_;
wire _34211_;
wire _34212_;
wire _34213_;
wire _34214_;
wire _34215_;
wire _34216_;
wire _34217_;
wire _34218_;
wire _34219_;
wire _34220_;
wire _34221_;
wire _34222_;
wire _34223_;
wire _34224_;
wire _34225_;
wire _34226_;
wire _34227_;
wire _34228_;
wire _34229_;
wire _34230_;
wire _34231_;
wire _34232_;
wire _34233_;
wire _34234_;
wire _34235_;
wire _34236_;
wire _34237_;
wire _34238_;
wire _34239_;
wire _34240_;
wire _34241_;
wire _34242_;
wire _34243_;
wire _34244_;
wire _34245_;
wire _34246_;
wire _34247_;
wire _34248_;
wire _34249_;
wire _34250_;
wire _34251_;
wire _34252_;
wire _34253_;
wire _34254_;
wire _34255_;
wire _34256_;
wire _34257_;
wire _34258_;
wire _34259_;
wire _34260_;
wire _34261_;
wire _34262_;
wire _34263_;
wire _34264_;
wire _34265_;
wire _34266_;
wire _34267_;
wire _34268_;
wire _34269_;
wire _34270_;
wire _34271_;
wire _34272_;
wire _34273_;
wire _34274_;
wire _34275_;
wire _34276_;
wire _34277_;
wire _34278_;
wire _34279_;
wire _34280_;
wire _34281_;
wire _34282_;
wire _34283_;
wire _34284_;
wire _34285_;
wire _34286_;
wire _34287_;
wire _34288_;
wire _34289_;
wire _34290_;
wire _34291_;
wire _34292_;
wire _34293_;
wire _34294_;
wire _34295_;
wire _34296_;
wire _34297_;
wire _34298_;
wire _34299_;
wire _34300_;
wire _34301_;
wire _34302_;
wire _34303_;
wire _34304_;
wire _34305_;
wire _34306_;
wire _34307_;
wire _34308_;
wire _34309_;
wire _34310_;
wire _34311_;
wire _34312_;
wire _34313_;
wire _34314_;
wire _34315_;
wire _34316_;
wire _34317_;
wire _34318_;
wire _34319_;
wire _34320_;
wire _34321_;
wire _34322_;
wire _34323_;
wire _34324_;
wire _34325_;
wire _34326_;
wire _34327_;
wire _34328_;
wire _34329_;
wire _34330_;
wire _34331_;
wire _34332_;
wire _34333_;
wire _34334_;
wire _34335_;
wire _34336_;
wire _34337_;
wire _34338_;
wire _34339_;
wire _34340_;
wire _34341_;
wire _34342_;
wire _34343_;
wire _34344_;
wire _34345_;
wire _34346_;
wire _34347_;
wire _34348_;
wire _34349_;
wire _34350_;
wire _34351_;
wire _34352_;
wire _34353_;
wire _34354_;
wire _34355_;
wire _34356_;
wire _34357_;
wire _34358_;
wire _34359_;
wire _34360_;
wire _34361_;
wire _34362_;
wire _34363_;
wire _34364_;
wire _34365_;
wire _34366_;
wire _34367_;
wire _34368_;
wire _34369_;
wire _34370_;
wire _34371_;
wire _34372_;
wire _34373_;
wire _34374_;
wire _34375_;
wire _34376_;
wire _34377_;
wire _34378_;
wire _34379_;
wire _34380_;
wire _34381_;
wire _34382_;
wire _34383_;
wire _34384_;
wire _34385_;
wire _34386_;
wire _34387_;
wire _34388_;
wire _34389_;
wire _34390_;
wire _34391_;
wire _34392_;
wire _34393_;
wire _34394_;
wire _34395_;
wire _34396_;
wire _34397_;
wire _34398_;
wire _34399_;
wire _34400_;
wire _34401_;
wire _34402_;
wire _34403_;
wire _34404_;
wire _34405_;
wire _34406_;
wire _34407_;
wire _34408_;
wire _34409_;
wire _34410_;
wire _34411_;
wire _34412_;
wire _34413_;
wire _34414_;
wire _34415_;
wire _34416_;
wire _34417_;
wire _34418_;
wire _34419_;
wire _34420_;
wire _34421_;
wire _34422_;
wire _34423_;
wire _34424_;
wire _34425_;
wire _34426_;
wire _34427_;
wire _34428_;
wire _34429_;
wire _34430_;
wire _34431_;
wire _34432_;
wire _34433_;
wire _34434_;
wire _34435_;
wire _34436_;
wire _34437_;
wire _34438_;
wire _34439_;
wire _34440_;
wire _34441_;
wire _34442_;
wire _34443_;
wire _34444_;
wire _34445_;
wire _34446_;
wire _34447_;
wire _34448_;
wire _34449_;
wire _34450_;
wire _34451_;
wire _34452_;
wire _34453_;
wire _34454_;
wire _34455_;
wire _34456_;
wire _34457_;
wire _34458_;
wire _34459_;
wire _34460_;
wire _34461_;
wire _34462_;
wire _34463_;
wire _34464_;
wire _34465_;
wire _34466_;
wire _34467_;
wire _34468_;
wire _34469_;
wire _34470_;
wire _34471_;
wire _34472_;
wire _34473_;
wire _34474_;
wire _34475_;
wire _34476_;
wire _34477_;
wire _34478_;
wire _34479_;
wire _34480_;
wire _34481_;
wire _34482_;
wire _34483_;
wire _34484_;
wire _34485_;
wire _34486_;
wire _34487_;
wire _34488_;
wire _34489_;
wire _34490_;
wire _34491_;
wire _34492_;
wire _34493_;
wire _34494_;
wire _34495_;
wire _34496_;
wire _34497_;
wire _34498_;
wire _34499_;
wire _34500_;
wire _34501_;
wire _34502_;
wire _34503_;
wire _34504_;
wire _34505_;
wire _34506_;
wire _34507_;
wire _34508_;
wire _34509_;
wire _34510_;
wire _34511_;
wire _34512_;
wire _34513_;
wire _34514_;
wire _34515_;
wire _34516_;
wire _34517_;
wire _34518_;
wire _34519_;
wire _34520_;
wire _34521_;
wire _34522_;
wire _34523_;
wire _34524_;
wire _34525_;
wire _34526_;
wire _34527_;
wire _34528_;
wire _34529_;
wire _34530_;
wire _34531_;
wire _34532_;
wire _34533_;
wire _34534_;
wire _34535_;
wire _34536_;
wire _34537_;
wire _34538_;
wire _34539_;
wire _34540_;
wire _34541_;
wire _34542_;
wire _34543_;
wire _34544_;
wire _34545_;
wire _34546_;
wire _34547_;
wire _34548_;
wire _34549_;
wire _34550_;
wire _34551_;
wire _34552_;
wire _34553_;
wire _34554_;
wire _34555_;
wire _34556_;
wire _34557_;
wire _34558_;
wire _34559_;
wire _34560_;
wire _34561_;
wire _34562_;
wire _34563_;
wire _34564_;
wire _34565_;
wire _34566_;
wire _34567_;
wire _34568_;
wire _34569_;
wire _34570_;
wire _34571_;
wire _34572_;
wire _34573_;
wire _34574_;
wire _34575_;
wire _34576_;
wire _34577_;
wire _34578_;
wire _34579_;
wire _34580_;
wire _34581_;
wire _34582_;
wire _34583_;
wire _34584_;
wire _34585_;
wire _34586_;
wire _34587_;
wire _34588_;
wire _34589_;
wire _34590_;
wire _34591_;
wire _34592_;
wire _34593_;
wire _34594_;
wire _34595_;
wire _34596_;
wire _34597_;
wire _34598_;
wire _34599_;
wire _34600_;
wire _34601_;
wire _34602_;
wire _34603_;
wire _34604_;
wire _34605_;
wire _34606_;
wire _34607_;
wire _34608_;
wire _34609_;
wire _34610_;
wire _34611_;
wire _34612_;
wire _34613_;
wire _34614_;
wire _34615_;
wire _34616_;
wire _34617_;
wire _34618_;
wire _34619_;
wire _34620_;
wire _34621_;
wire _34622_;
wire _34623_;
wire _34624_;
wire _34625_;
wire _34626_;
wire _34627_;
wire _34628_;
wire _34629_;
wire _34630_;
wire _34631_;
wire _34632_;
wire _34633_;
wire _34634_;
wire _34635_;
wire _34636_;
wire _34637_;
wire _34638_;
wire _34639_;
wire _34640_;
wire _34641_;
wire _34642_;
wire _34643_;
wire _34644_;
wire _34645_;
wire _34646_;
wire _34647_;
wire _34648_;
wire _34649_;
wire _34650_;
wire _34651_;
wire _34652_;
wire _34653_;
wire _34654_;
wire _34655_;
wire _34656_;
wire _34657_;
wire _34658_;
wire _34659_;
wire _34660_;
wire _34661_;
wire _34662_;
wire _34663_;
wire _34664_;
wire _34665_;
wire _34666_;
wire _34667_;
wire _34668_;
wire _34669_;
wire _34670_;
wire _34671_;
wire _34672_;
wire _34673_;
wire _34674_;
wire _34675_;
wire _34676_;
wire _34677_;
wire _34678_;
wire _34679_;
wire _34680_;
wire _34681_;
wire _34682_;
wire _34683_;
wire _34684_;
wire _34685_;
wire _34686_;
wire _34687_;
wire _34688_;
wire _34689_;
wire _34690_;
wire _34691_;
wire _34692_;
wire _34693_;
wire _34694_;
wire _34695_;
wire _34696_;
wire _34697_;
wire _34698_;
wire _34699_;
wire _34700_;
wire _34701_;
wire _34702_;
wire _34703_;
wire _34704_;
wire _34705_;
wire _34706_;
wire _34707_;
wire _34708_;
wire _34709_;
wire _34710_;
wire _34711_;
wire _34712_;
wire _34713_;
wire _34714_;
wire _34715_;
wire _34716_;
wire _34717_;
wire _34718_;
wire _34719_;
wire _34720_;
wire _34721_;
wire _34722_;
wire _34723_;
wire _34724_;
wire _34725_;
wire _34726_;
wire _34727_;
wire _34728_;
wire _34729_;
wire _34730_;
wire _34731_;
wire _34732_;
wire _34733_;
wire _34734_;
wire _34735_;
wire _34736_;
wire _34737_;
wire _34738_;
wire _34739_;
wire _34740_;
wire _34741_;
wire _34742_;
wire _34743_;
wire _34744_;
wire _34745_;
wire _34746_;
wire _34747_;
wire _34748_;
wire _34749_;
wire _34750_;
wire _34751_;
wire _34752_;
wire _34753_;
wire _34754_;
wire _34755_;
wire _34756_;
wire _34757_;
wire _34758_;
wire _34759_;
wire _34760_;
wire _34761_;
wire _34762_;
wire _34763_;
wire _34764_;
wire _34765_;
wire _34766_;
wire _34767_;
wire _34768_;
wire _34769_;
wire _34770_;
wire _34771_;
wire _34772_;
wire _34773_;
wire _34774_;
wire _34775_;
wire _34776_;
wire _34777_;
wire _34778_;
wire _34779_;
wire _34780_;
wire _34781_;
wire _34782_;
wire _34783_;
wire _34784_;
wire _34785_;
wire _34786_;
wire _34787_;
wire _34788_;
wire _34789_;
wire _34790_;
wire _34791_;
wire _34792_;
wire _34793_;
wire _34794_;
wire _34795_;
wire _34796_;
wire _34797_;
wire _34798_;
wire _34799_;
wire _34800_;
wire _34801_;
wire _34802_;
wire _34803_;
wire _34804_;
wire _34805_;
wire _34806_;
wire _34807_;
wire _34808_;
wire _34809_;
wire _34810_;
wire _34811_;
wire _34812_;
wire _34813_;
wire _34814_;
wire _34815_;
wire _34816_;
wire _34817_;
wire _34818_;
wire _34819_;
wire _34820_;
wire _34821_;
wire _34822_;
wire _34823_;
wire _34824_;
wire _34825_;
wire _34826_;
wire _34827_;
wire _34828_;
wire _34829_;
wire _34830_;
wire _34831_;
wire _34832_;
wire _34833_;
wire _34834_;
wire _34835_;
wire _34836_;
wire _34837_;
wire _34838_;
wire _34839_;
wire _34840_;
wire _34841_;
wire _34842_;
wire _34843_;
wire _34844_;
wire _34845_;
wire _34846_;
wire _34847_;
wire _34848_;
wire _34849_;
wire _34850_;
wire _34851_;
wire _34852_;
wire _34853_;
wire _34854_;
wire _34855_;
wire _34856_;
wire _34857_;
wire _34858_;
wire _34859_;
wire _34860_;
wire _34861_;
wire _34862_;
wire _34863_;
wire _34864_;
wire _34865_;
wire _34866_;
wire _34867_;
wire _34868_;
wire _34869_;
wire _34870_;
wire _34871_;
wire _34872_;
wire _34873_;
wire _34874_;
wire _34875_;
wire _34876_;
wire _34877_;
wire _34878_;
wire _34879_;
wire _34880_;
wire _34881_;
wire _34882_;
wire _34883_;
wire _34884_;
wire _34885_;
wire _34886_;
wire _34887_;
wire _34888_;
wire _34889_;
wire _34890_;
wire _34891_;
wire _34892_;
wire _34893_;
wire _34894_;
wire _34895_;
wire _34896_;
wire _34897_;
wire _34898_;
wire _34899_;
wire _34900_;
wire _34901_;
wire _34902_;
wire _34903_;
wire _34904_;
wire _34905_;
wire _34906_;
wire _34907_;
wire _34908_;
wire _34909_;
wire _34910_;
wire _34911_;
wire _34912_;
wire _34913_;
wire _34914_;
wire _34915_;
wire _34916_;
wire _34917_;
wire _34918_;
wire _34919_;
wire _34920_;
wire _34921_;
wire _34922_;
wire _34923_;
wire _34924_;
wire _34925_;
wire _34926_;
wire _34927_;
wire _34928_;
wire _34929_;
wire _34930_;
wire _34931_;
wire _34932_;
wire _34933_;
wire _34934_;
wire _34935_;
wire _34936_;
wire _34937_;
wire _34938_;
wire _34939_;
wire _34940_;
wire _34941_;
wire _34942_;
wire _34943_;
wire _34944_;
wire _34945_;
wire _34946_;
wire _34947_;
wire _34948_;
wire _34949_;
wire _34950_;
wire _34951_;
wire _34952_;
wire _34953_;
wire _34954_;
wire _34955_;
wire _34956_;
wire _34957_;
wire _34958_;
wire _34959_;
wire _34960_;
wire _34961_;
wire _34962_;
wire _34963_;
wire _34964_;
wire _34965_;
wire _34966_;
wire _34967_;
wire _34968_;
wire _34969_;
wire _34970_;
wire _34971_;
wire _34972_;
wire _34973_;
wire _34974_;
wire _34975_;
wire _34976_;
wire _34977_;
wire _34978_;
wire _34979_;
wire _34980_;
wire _34981_;
wire _34982_;
wire _34983_;
wire _34984_;
wire _34985_;
wire _34986_;
wire _34987_;
wire _34988_;
wire _34989_;
wire _34990_;
wire _34991_;
wire _34992_;
wire _34993_;
wire _34994_;
wire _34995_;
wire _34996_;
wire _34997_;
wire _34998_;
wire _34999_;
wire _35000_;
wire _35001_;
wire _35002_;
wire _35003_;
wire _35004_;
wire _35005_;
wire _35006_;
wire _35007_;
wire _35008_;
wire _35009_;
wire _35010_;
wire _35011_;
wire _35012_;
wire _35013_;
wire _35014_;
wire _35015_;
wire _35016_;
wire _35017_;
wire _35018_;
wire _35019_;
wire _35020_;
wire _35021_;
wire _35022_;
wire _35023_;
wire _35024_;
wire _35025_;
wire _35026_;
wire _35027_;
wire _35028_;
wire _35029_;
wire _35030_;
wire _35031_;
wire _35032_;
wire _35033_;
wire _35034_;
wire _35035_;
wire _35036_;
wire _35037_;
wire _35038_;
wire _35039_;
wire _35040_;
wire _35041_;
wire _35042_;
wire _35043_;
wire _35044_;
wire _35045_;
wire _35046_;
wire _35047_;
wire _35048_;
wire _35049_;
wire _35050_;
wire _35051_;
wire _35052_;
wire _35053_;
wire _35054_;
wire _35055_;
wire _35056_;
wire _35057_;
wire _35058_;
wire _35059_;
wire _35060_;
wire _35061_;
wire _35062_;
wire _35063_;
wire _35064_;
wire _35065_;
wire _35066_;
wire _35067_;
wire _35068_;
wire _35069_;
wire _35070_;
wire _35071_;
wire _35072_;
wire _35073_;
wire _35074_;
wire _35075_;
wire _35076_;
wire _35077_;
wire _35078_;
wire _35079_;
wire _35080_;
wire _35081_;
wire _35082_;
wire _35083_;
wire _35084_;
wire _35085_;
wire _35086_;
wire _35087_;
wire _35088_;
wire _35089_;
wire _35090_;
wire _35091_;
wire _35092_;
wire _35093_;
wire _35094_;
wire _35095_;
wire _35096_;
wire _35097_;
wire _35098_;
wire _35099_;
wire _35100_;
wire _35101_;
wire _35102_;
wire _35103_;
wire _35104_;
wire _35105_;
wire _35106_;
wire _35107_;
wire _35108_;
wire _35109_;
wire _35110_;
wire _35111_;
wire _35112_;
wire _35113_;
wire _35114_;
wire _35115_;
wire _35116_;
wire _35117_;
wire _35118_;
wire _35119_;
wire _35120_;
wire _35121_;
wire _35122_;
wire _35123_;
wire _35124_;
wire _35125_;
wire _35126_;
wire _35127_;
wire _35128_;
wire _35129_;
wire _35130_;
wire _35131_;
wire _35132_;
wire _35133_;
wire _35134_;
wire _35135_;
wire _35136_;
wire _35137_;
wire _35138_;
wire _35139_;
wire _35140_;
wire _35141_;
wire _35142_;
wire _35143_;
wire _35144_;
wire _35145_;
wire _35146_;
wire _35147_;
wire _35148_;
wire _35149_;
wire _35150_;
wire _35151_;
wire _35152_;
wire _35153_;
wire _35154_;
wire _35155_;
wire _35156_;
wire _35157_;
wire _35158_;
wire _35159_;
wire _35160_;
wire _35161_;
wire _35162_;
wire _35163_;
wire _35164_;
wire _35165_;
wire _35166_;
wire _35167_;
wire _35168_;
wire _35169_;
wire _35170_;
wire _35171_;
wire _35172_;
wire _35173_;
wire _35174_;
wire _35175_;
wire _35176_;
wire _35177_;
wire _35178_;
wire _35179_;
wire _35180_;
wire _35181_;
wire _35182_;
wire _35183_;
wire _35184_;
wire _35185_;
wire _35186_;
wire _35187_;
wire _35188_;
wire _35189_;
wire _35190_;
wire _35191_;
wire _35192_;
wire _35193_;
wire _35194_;
wire _35195_;
wire _35196_;
wire _35197_;
wire _35198_;
wire _35199_;
wire _35200_;
wire _35201_;
wire _35202_;
wire _35203_;
wire _35204_;
wire _35205_;
wire _35206_;
wire _35207_;
wire _35208_;
wire _35209_;
wire _35210_;
wire _35211_;
wire _35212_;
wire _35213_;
wire _35214_;
wire _35215_;
wire _35216_;
wire _35217_;
wire _35218_;
wire _35219_;
wire _35220_;
wire _35221_;
wire _35222_;
wire _35223_;
wire _35224_;
wire _35225_;
wire _35226_;
wire _35227_;
wire _35228_;
wire _35229_;
wire _35230_;
wire _35231_;
wire _35232_;
wire _35233_;
wire _35234_;
wire _35235_;
wire _35236_;
wire _35237_;
wire _35238_;
wire _35239_;
wire _35240_;
wire _35241_;
wire _35242_;
wire _35243_;
wire _35244_;
wire _35245_;
wire _35246_;
wire _35247_;
wire _35248_;
wire _35249_;
wire _35250_;
wire _35251_;
wire _35252_;
wire _35253_;
wire _35254_;
wire _35255_;
wire _35256_;
wire _35257_;
wire _35258_;
wire _35259_;
wire _35260_;
wire _35261_;
wire _35262_;
wire _35263_;
wire _35264_;
wire _35265_;
wire _35266_;
wire _35267_;
wire _35268_;
wire _35269_;
wire _35270_;
wire _35271_;
wire _35272_;
wire _35273_;
wire _35274_;
wire _35275_;
wire _35276_;
wire _35277_;
wire _35278_;
wire _35279_;
wire _35280_;
wire _35281_;
wire _35282_;
wire _35283_;
wire _35284_;
wire _35285_;
wire _35286_;
wire _35287_;
wire _35288_;
wire _35289_;
wire _35290_;
wire _35291_;
wire _35292_;
wire _35293_;
wire _35294_;
wire _35295_;
wire _35296_;
wire _35297_;
wire _35298_;
wire _35299_;
wire _35300_;
wire _35301_;
wire _35302_;
wire _35303_;
wire _35304_;
wire _35305_;
wire _35306_;
wire _35307_;
wire _35308_;
wire _35309_;
wire _35310_;
wire _35311_;
wire _35312_;
wire _35313_;
wire _35314_;
wire _35315_;
wire _35316_;
wire _35317_;
wire _35318_;
wire _35319_;
wire _35320_;
wire _35321_;
wire _35322_;
wire _35323_;
wire _35324_;
wire _35325_;
wire _35326_;
wire _35327_;
wire _35328_;
wire _35329_;
wire _35330_;
wire _35331_;
wire _35332_;
wire _35333_;
wire _35334_;
wire _35335_;
wire _35336_;
wire _35337_;
wire _35338_;
wire _35339_;
wire _35340_;
wire _35341_;
wire _35342_;
wire _35343_;
wire _35344_;
wire _35345_;
wire _35346_;
wire _35347_;
wire _35348_;
wire _35349_;
wire _35350_;
wire _35351_;
wire _35352_;
wire _35353_;
wire _35354_;
wire _35355_;
wire _35356_;
wire _35357_;
wire _35358_;
wire _35359_;
wire _35360_;
wire _35361_;
wire _35362_;
wire _35363_;
wire _35364_;
wire _35365_;
wire _35366_;
wire _35367_;
wire _35368_;
wire _35369_;
wire _35370_;
wire _35371_;
wire _35372_;
wire _35373_;
wire _35374_;
wire _35375_;
wire _35376_;
wire _35377_;
wire _35378_;
wire _35379_;
wire _35380_;
wire _35381_;
wire _35382_;
wire _35383_;
wire _35384_;
wire _35385_;
wire _35386_;
wire _35387_;
wire _35388_;
wire _35389_;
wire _35390_;
wire _35391_;
wire _35392_;
wire _35393_;
wire _35394_;
wire _35395_;
wire _35396_;
wire _35397_;
wire _35398_;
wire _35399_;
wire _35400_;
wire _35401_;
wire _35402_;
wire _35403_;
wire _35404_;
wire _35405_;
wire _35406_;
wire _35407_;
wire _35408_;
wire _35409_;
wire _35410_;
wire _35411_;
wire _35412_;
wire _35413_;
wire _35414_;
wire _35415_;
wire _35416_;
wire _35417_;
wire _35418_;
wire _35419_;
wire _35420_;
wire _35421_;
wire _35422_;
wire _35423_;
wire _35424_;
wire _35425_;
wire _35426_;
wire _35427_;
wire _35428_;
wire _35429_;
wire _35430_;
wire _35431_;
wire _35432_;
wire _35433_;
wire _35434_;
wire _35435_;
wire _35436_;
wire _35437_;
wire _35438_;
wire _35439_;
wire _35440_;
wire _35441_;
wire _35442_;
wire _35443_;
wire _35444_;
wire _35445_;
wire _35446_;
wire _35447_;
wire _35448_;
wire _35449_;
wire _35450_;
wire _35451_;
wire _35452_;
wire _35453_;
wire _35454_;
wire _35455_;
wire _35456_;
wire _35457_;
wire _35458_;
wire _35459_;
wire _35460_;
wire _35461_;
wire _35462_;
wire _35463_;
wire _35464_;
wire _35465_;
wire _35466_;
wire _35467_;
wire _35468_;
wire _35469_;
wire _35470_;
wire _35471_;
wire _35472_;
wire _35473_;
wire _35474_;
wire _35475_;
wire _35476_;
wire _35477_;
wire _35478_;
wire _35479_;
wire _35480_;
wire _35481_;
wire _35482_;
wire _35483_;
wire _35484_;
wire _35485_;
wire _35486_;
wire _35487_;
wire _35488_;
wire _35489_;
wire _35490_;
wire _35491_;
wire _35492_;
wire _35493_;
wire _35494_;
wire _35495_;
wire _35496_;
wire _35497_;
wire _35498_;
wire _35499_;
wire _35500_;
wire _35501_;
wire _35502_;
wire _35503_;
wire _35504_;
wire _35505_;
wire _35506_;
wire _35507_;
wire _35508_;
wire _35509_;
wire _35510_;
wire _35511_;
wire _35512_;
wire _35513_;
wire _35514_;
wire _35515_;
wire _35516_;
wire _35517_;
wire _35518_;
wire _35519_;
wire _35520_;
wire _35521_;
wire _35522_;
wire _35523_;
wire _35524_;
wire _35525_;
wire _35526_;
wire _35527_;
wire _35528_;
wire _35529_;
wire _35530_;
wire _35531_;
wire _35532_;
wire _35533_;
wire _35534_;
wire _35535_;
wire _35536_;
wire _35537_;
wire _35538_;
wire _35539_;
wire _35540_;
wire _35541_;
wire _35542_;
wire _35543_;
wire _35544_;
wire _35545_;
wire _35546_;
wire _35547_;
wire _35548_;
wire _35549_;
wire _35550_;
wire _35551_;
wire _35552_;
wire _35553_;
wire _35554_;
wire _35555_;
wire _35556_;
wire _35557_;
wire _35558_;
wire _35559_;
wire _35560_;
wire _35561_;
wire _35562_;
wire _35563_;
wire _35564_;
wire _35565_;
wire _35566_;
wire _35567_;
wire _35568_;
wire _35569_;
wire _35570_;
wire _35571_;
wire _35572_;
wire _35573_;
wire _35574_;
wire _35575_;
wire _35576_;
wire _35577_;
wire _35578_;
wire _35579_;
wire _35580_;
wire _35581_;
wire _35582_;
wire _35583_;
wire _35584_;
wire _35585_;
wire _35586_;
wire _35587_;
wire _35588_;
wire _35589_;
wire _35590_;
wire _35591_;
wire _35592_;
wire _35593_;
wire _35594_;
wire _35595_;
wire _35596_;
wire _35597_;
wire _35598_;
wire _35599_;
wire _35600_;
wire _35601_;
wire _35602_;
wire _35603_;
wire _35604_;
wire _35605_;
wire _35606_;
wire _35607_;
wire _35608_;
wire _35609_;
wire _35610_;
wire _35611_;
wire _35612_;
wire _35613_;
wire _35614_;
wire _35615_;
wire _35616_;
wire _35617_;
wire _35618_;
wire _35619_;
wire _35620_;
wire _35621_;
wire _35622_;
wire _35623_;
wire _35624_;
wire _35625_;
wire _35626_;
wire _35627_;
wire _35628_;
wire _35629_;
wire _35630_;
wire _35631_;
wire _35632_;
wire _35633_;
wire _35634_;
wire _35635_;
wire _35636_;
wire _35637_;
wire _35638_;
wire _35639_;
wire _35640_;
wire _35641_;
wire _35642_;
wire _35643_;
wire _35644_;
wire _35645_;
wire _35646_;
wire _35647_;
wire _35648_;
wire _35649_;
wire _35650_;
wire _35651_;
wire _35652_;
wire _35653_;
wire _35654_;
wire _35655_;
wire _35656_;
wire _35657_;
wire _35658_;
wire _35659_;
wire _35660_;
wire _35661_;
wire _35662_;
wire _35663_;
wire _35664_;
wire _35665_;
wire _35666_;
wire _35667_;
wire _35668_;
wire _35669_;
wire _35670_;
wire _35671_;
wire _35672_;
wire _35673_;
wire _35674_;
wire _35675_;
wire _35676_;
wire _35677_;
wire _35678_;
wire _35679_;
wire _35680_;
wire _35681_;
wire _35682_;
wire _35683_;
wire _35684_;
wire _35685_;
wire _35686_;
wire _35687_;
wire _35688_;
wire _35689_;
wire _35690_;
wire _35691_;
wire _35692_;
wire _35693_;
wire _35694_;
wire _35695_;
wire _35696_;
wire _35697_;
wire _35698_;
wire _35699_;
wire _35700_;
wire _35701_;
wire _35702_;
wire _35703_;
wire _35704_;
wire _35705_;
wire _35706_;
wire _35707_;
wire _35708_;
wire _35709_;
wire _35710_;
wire _35711_;
wire _35712_;
wire _35713_;
wire _35714_;
wire _35715_;
wire _35716_;
wire _35717_;
wire _35718_;
wire _35719_;
wire _35720_;
wire _35721_;
wire _35722_;
wire _35723_;
wire _35724_;
wire _35725_;
wire _35726_;
wire _35727_;
wire _35728_;
wire _35729_;
wire _35730_;
wire _35731_;
wire _35732_;
wire _35733_;
wire _35734_;
wire _35735_;
wire _35736_;
wire _35737_;
wire _35738_;
wire _35739_;
wire _35740_;
wire _35741_;
wire _35742_;
wire _35743_;
wire _35744_;
wire _35745_;
wire _35746_;
wire _35747_;
wire _35748_;
wire _35749_;
wire _35750_;
wire _35751_;
wire _35752_;
wire _35753_;
wire _35754_;
wire _35755_;
wire _35756_;
wire _35757_;
wire _35758_;
wire _35759_;
wire _35760_;
wire _35761_;
wire _35762_;
wire _35763_;
wire _35764_;
wire _35765_;
wire _35766_;
wire _35767_;
wire _35768_;
wire _35769_;
wire _35770_;
wire _35771_;
wire _35772_;
wire _35773_;
wire _35774_;
wire _35775_;
wire _35776_;
wire _35777_;
wire _35778_;
wire _35779_;
wire _35780_;
wire _35781_;
wire _35782_;
wire _35783_;
wire _35784_;
wire _35785_;
wire _35786_;
wire _35787_;
wire _35788_;
wire _35789_;
wire _35790_;
wire _35791_;
wire _35792_;
wire _35793_;
wire _35794_;
wire _35795_;
wire _35796_;
wire _35797_;
wire _35798_;
wire _35799_;
wire _35800_;
wire _35801_;
wire _35802_;
wire _35803_;
wire _35804_;
wire _35805_;
wire _35806_;
wire _35807_;
wire _35808_;
wire _35809_;
wire _35810_;
wire _35811_;
wire _35812_;
wire _35813_;
wire _35814_;
wire _35815_;
wire _35816_;
wire _35817_;
wire _35818_;
wire _35819_;
wire _35820_;
wire _35821_;
wire _35822_;
wire _35823_;
wire _35824_;
wire _35825_;
wire _35826_;
wire _35827_;
wire _35828_;
wire _35829_;
wire _35830_;
wire _35831_;
wire _35832_;
wire _35833_;
wire _35834_;
wire _35835_;
wire _35836_;
wire _35837_;
wire _35838_;
wire _35839_;
wire _35840_;
wire _35841_;
wire _35842_;
wire _35843_;
wire _35844_;
wire _35845_;
wire _35846_;
wire _35847_;
wire _35848_;
wire _35849_;
wire _35850_;
wire _35851_;
wire _35852_;
wire _35853_;
wire _35854_;
wire _35855_;
wire _35856_;
wire _35857_;
wire _35858_;
wire _35859_;
wire _35860_;
wire _35861_;
wire _35862_;
wire _35863_;
wire _35864_;
wire _35865_;
wire _35866_;
wire _35867_;
wire _35868_;
wire _35869_;
wire _35870_;
wire _35871_;
wire _35872_;
wire _35873_;
wire _35874_;
wire _35875_;
wire _35876_;
wire _35877_;
wire _35878_;
wire _35879_;
wire _35880_;
wire _35881_;
wire _35882_;
wire _35883_;
wire _35884_;
wire _35885_;
wire _35886_;
wire _35887_;
wire _35888_;
wire _35889_;
wire _35890_;
wire _35891_;
wire _35892_;
wire _35893_;
wire _35894_;
wire _35895_;
wire _35896_;
wire _35897_;
wire _35898_;
wire _35899_;
wire _35900_;
wire _35901_;
wire _35902_;
wire _35903_;
wire _35904_;
wire _35905_;
wire _35906_;
wire _35907_;
wire _35908_;
wire _35909_;
wire _35910_;
wire _35911_;
wire _35912_;
wire _35913_;
wire _35914_;
wire _35915_;
wire _35916_;
wire _35917_;
wire _35918_;
wire _35919_;
wire _35920_;
wire _35921_;
wire _35922_;
wire _35923_;
wire _35924_;
wire _35925_;
wire _35926_;
wire _35927_;
wire _35928_;
wire _35929_;
wire _35930_;
wire _35931_;
wire _35932_;
wire _35933_;
wire _35934_;
wire _35935_;
wire _35936_;
wire _35937_;
wire _35938_;
wire _35939_;
wire _35940_;
wire _35941_;
wire _35942_;
wire _35943_;
wire _35944_;
wire _35945_;
wire _35946_;
wire _35947_;
wire _35948_;
wire _35949_;
wire _35950_;
wire _35951_;
wire _35952_;
wire _35953_;
wire _35954_;
wire _35955_;
wire _35956_;
wire _35957_;
wire _35958_;
wire _35959_;
wire _35960_;
wire _35961_;
wire _35962_;
wire _35963_;
wire _35964_;
wire _35965_;
wire _35966_;
wire _35967_;
wire _35968_;
wire _35969_;
wire _35970_;
wire _35971_;
wire _35972_;
wire _35973_;
wire _35974_;
wire _35975_;
wire _35976_;
wire _35977_;
wire _35978_;
wire _35979_;
wire _35980_;
wire _35981_;
wire _35982_;
wire _35983_;
wire _35984_;
wire _35985_;
wire _35986_;
wire _35987_;
wire _35988_;
wire _35989_;
wire _35990_;
wire _35991_;
wire _35992_;
wire _35993_;
wire _35994_;
wire _35995_;
wire _35996_;
wire _35997_;
wire _35998_;
wire _35999_;
wire _36000_;
wire _36001_;
wire _36002_;
wire _36003_;
wire _36004_;
wire _36005_;
wire _36006_;
wire _36007_;
wire _36008_;
wire _36009_;
wire _36010_;
wire _36011_;
wire _36012_;
wire _36013_;
wire _36014_;
wire _36015_;
wire _36016_;
wire _36017_;
wire _36018_;
wire _36019_;
wire _36020_;
wire _36021_;
wire _36022_;
wire _36023_;
wire _36024_;
wire _36025_;
wire _36026_;
wire _36027_;
wire _36028_;
wire _36029_;
wire _36030_;
wire _36031_;
wire _36032_;
wire _36033_;
wire _36034_;
wire _36035_;
wire _36036_;
wire _36037_;
wire _36038_;
wire _36039_;
wire _36040_;
wire _36041_;
wire _36042_;
wire _36043_;
wire _36044_;
wire _36045_;
wire _36046_;
wire _36047_;
wire _36048_;
wire _36049_;
wire _36050_;
wire _36051_;
wire _36052_;
wire _36053_;
wire _36054_;
wire _36055_;
wire _36056_;
wire _36057_;
wire _36058_;
wire _36059_;
wire _36060_;
wire _36061_;
wire _36062_;
wire _36063_;
wire _36064_;
wire _36065_;
wire _36066_;
wire _36067_;
wire _36068_;
wire _36069_;
wire _36070_;
wire _36071_;
wire _36072_;
wire _36073_;
wire _36074_;
wire _36075_;
wire _36076_;
wire _36077_;
wire _36078_;
wire _36079_;
wire _36080_;
wire _36081_;
wire _36082_;
wire _36083_;
wire _36084_;
wire _36085_;
wire _36086_;
wire _36087_;
wire _36088_;
wire _36089_;
wire _36090_;
wire _36091_;
wire _36092_;
wire _36093_;
wire _36094_;
wire _36095_;
wire _36096_;
wire _36097_;
wire _36098_;
wire _36099_;
wire _36100_;
wire _36101_;
wire _36102_;
wire _36103_;
wire _36104_;
wire _36105_;
wire _36106_;
wire _36107_;
wire _36108_;
wire _36109_;
wire _36110_;
wire _36111_;
wire _36112_;
wire _36113_;
wire _36114_;
wire _36115_;
wire _36116_;
wire _36117_;
wire _36118_;
wire _36119_;
wire _36120_;
wire _36121_;
wire _36122_;
wire _36123_;
wire _36124_;
wire _36125_;
wire _36126_;
wire _36127_;
wire _36128_;
wire _36129_;
wire _36130_;
wire _36131_;
wire _36132_;
wire _36133_;
wire _36134_;
wire _36135_;
wire _36136_;
wire _36137_;
wire _36138_;
wire _36139_;
wire _36140_;
wire _36141_;
wire _36142_;
wire _36143_;
wire _36144_;
wire _36145_;
wire _36146_;
wire _36147_;
wire _36148_;
wire _36149_;
wire _36150_;
wire _36151_;
wire _36152_;
wire _36153_;
wire _36154_;
wire _36155_;
wire _36156_;
wire _36157_;
wire _36158_;
wire _36159_;
wire _36160_;
wire _36161_;
wire _36162_;
wire _36163_;
wire _36164_;
wire _36165_;
wire _36166_;
wire _36167_;
wire _36168_;
wire _36169_;
wire _36170_;
wire _36171_;
wire _36172_;
wire _36173_;
wire _36174_;
wire _36175_;
wire _36176_;
wire _36177_;
wire _36178_;
wire _36179_;
wire _36180_;
wire _36181_;
wire _36182_;
wire _36183_;
wire _36184_;
wire _36185_;
wire _36186_;
wire _36187_;
wire _36188_;
wire _36189_;
wire _36190_;
wire _36191_;
wire _36192_;
wire _36193_;
wire _36194_;
wire _36195_;
wire _36196_;
wire _36197_;
wire _36198_;
wire _36199_;
wire _36200_;
wire _36201_;
wire _36202_;
wire _36203_;
wire _36204_;
wire _36205_;
wire _36206_;
wire _36207_;
wire _36208_;
wire _36209_;
wire _36210_;
wire _36211_;
wire _36212_;
wire _36213_;
wire _36214_;
wire _36215_;
wire _36216_;
wire _36217_;
wire _36218_;
wire _36219_;
wire _36220_;
wire _36221_;
wire _36222_;
wire _36223_;
wire _36224_;
wire _36225_;
wire _36226_;
wire _36227_;
wire _36228_;
wire _36229_;
wire _36230_;
wire _36231_;
wire _36232_;
wire _36233_;
wire _36234_;
wire _36235_;
wire _36236_;
wire _36237_;
wire _36238_;
wire _36239_;
wire _36240_;
wire _36241_;
wire _36242_;
wire _36243_;
wire _36244_;
wire _36245_;
wire _36246_;
wire _36247_;
wire _36248_;
wire _36249_;
wire _36250_;
wire _36251_;
wire _36252_;
wire _36253_;
wire _36254_;
wire _36255_;
wire _36256_;
wire _36257_;
wire _36258_;
wire _36259_;
wire _36260_;
wire _36261_;
wire _36262_;
wire _36263_;
wire _36264_;
wire _36265_;
wire _36266_;
wire _36267_;
wire _36268_;
wire _36269_;
wire _36270_;
wire _36271_;
wire _36272_;
wire _36273_;
wire _36274_;
wire _36275_;
wire _36276_;
wire _36277_;
wire _36278_;
wire _36279_;
wire _36280_;
wire _36281_;
wire _36282_;
wire _36283_;
wire _36284_;
wire _36285_;
wire _36286_;
wire _36287_;
wire _36288_;
wire _36289_;
wire _36290_;
wire _36291_;
wire _36292_;
wire _36293_;
wire _36294_;
wire _36295_;
wire _36296_;
wire _36297_;
wire _36298_;
wire _36299_;
wire _36300_;
wire _36301_;
wire _36302_;
wire _36303_;
wire _36304_;
wire _36305_;
wire _36306_;
wire _36307_;
wire _36308_;
wire _36309_;
wire _36310_;
wire _36311_;
wire _36312_;
wire _36313_;
wire _36314_;
wire _36315_;
wire _36316_;
wire _36317_;
wire _36318_;
wire _36319_;
wire _36320_;
wire _36321_;
wire _36322_;
wire _36323_;
wire _36324_;
wire _36325_;
wire _36326_;
wire _36327_;
wire _36328_;
wire _36329_;
wire _36330_;
wire _36331_;
wire _36332_;
wire _36333_;
wire _36334_;
wire _36335_;
wire _36336_;
wire _36337_;
wire _36338_;
wire _36339_;
wire _36340_;
wire _36341_;
wire _36342_;
wire _36343_;
wire _36344_;
wire _36345_;
wire _36346_;
wire _36347_;
wire _36348_;
wire _36349_;
wire _36350_;
wire _36351_;
wire _36352_;
wire _36353_;
wire _36354_;
wire _36355_;
wire _36356_;
wire _36357_;
wire _36358_;
wire _36359_;
wire _36360_;
wire _36361_;
wire _36362_;
wire _36363_;
wire _36364_;
wire _36365_;
wire _36366_;
wire _36367_;
wire _36368_;
wire _36369_;
wire _36370_;
wire _36371_;
wire _36372_;
wire _36373_;
wire _36374_;
wire _36375_;
wire _36376_;
wire _36377_;
wire _36378_;
wire _36379_;
wire _36380_;
wire _36381_;
wire _36382_;
wire _36383_;
wire _36384_;
wire _36385_;
wire _36386_;
wire _36387_;
wire _36388_;
wire _36389_;
wire _36390_;
wire _36391_;
wire _36392_;
wire _36393_;
wire _36394_;
wire _36395_;
wire _36396_;
wire _36397_;
wire _36398_;
wire _36399_;
wire _36400_;
wire _36401_;
wire _36402_;
wire _36403_;
wire _36404_;
wire _36405_;
wire _36406_;
wire _36407_;
wire _36408_;
wire _36409_;
wire _36410_;
wire _36411_;
wire _36412_;
wire _36413_;
wire _36414_;
wire _36415_;
wire _36416_;
wire _36417_;
wire _36418_;
wire _36419_;
wire _36420_;
wire _36421_;
wire _36422_;
wire _36423_;
wire _36424_;
wire _36425_;
wire _36426_;
wire _36427_;
wire _36428_;
wire _36429_;
wire _36430_;
wire _36431_;
wire _36432_;
wire _36433_;
wire _36434_;
wire _36435_;
wire _36436_;
wire _36437_;
wire _36438_;
wire _36439_;
wire _36440_;
wire _36441_;
wire _36442_;
wire _36443_;
wire _36444_;
wire _36445_;
wire _36446_;
wire _36447_;
wire _36448_;
wire _36449_;
wire _36450_;
wire _36451_;
wire _36452_;
wire _36453_;
wire _36454_;
wire _36455_;
wire _36456_;
wire _36457_;
wire _36458_;
wire _36459_;
wire _36460_;
wire _36461_;
wire _36462_;
wire _36463_;
wire _36464_;
wire _36465_;
wire _36466_;
wire _36467_;
wire _36468_;
wire _36469_;
wire _36470_;
wire _36471_;
wire _36472_;
wire _36473_;
wire _36474_;
wire _36475_;
wire _36476_;
wire _36477_;
wire _36478_;
wire _36479_;
wire _36480_;
wire _36481_;
wire _36482_;
wire _36483_;
wire _36484_;
wire _36485_;
wire _36486_;
wire _36487_;
wire _36488_;
wire _36489_;
wire _36490_;
wire _36491_;
wire _36492_;
wire _36493_;
wire _36494_;
wire _36495_;
wire _36496_;
wire _36497_;
wire _36498_;
wire _36499_;
wire _36500_;
wire _36501_;
wire _36502_;
wire _36503_;
wire _36504_;
wire _36505_;
wire _36506_;
wire _36507_;
wire _36508_;
wire _36509_;
wire _36510_;
wire _36511_;
wire _36512_;
wire _36513_;
wire _36514_;
wire _36515_;
wire _36516_;
wire _36517_;
wire _36518_;
wire _36519_;
wire _36520_;
wire _36521_;
wire _36522_;
wire _36523_;
wire _36524_;
wire _36525_;
wire _36526_;
wire _36527_;
wire _36528_;
wire _36529_;
wire _36530_;
wire _36531_;
wire _36532_;
wire _36533_;
wire _36534_;
wire _36535_;
wire _36536_;
wire _36537_;
wire _36538_;
wire _36539_;
wire _36540_;
wire _36541_;
wire _36542_;
wire _36543_;
wire _36544_;
wire _36545_;
wire _36546_;
wire _36547_;
wire _36548_;
wire _36549_;
wire _36550_;
wire _36551_;
wire _36552_;
wire _36553_;
wire _36554_;
wire _36555_;
wire _36556_;
wire _36557_;
wire _36558_;
wire _36559_;
wire _36560_;
wire _36561_;
wire _36562_;
wire _36563_;
wire _36564_;
wire _36565_;
wire _36566_;
wire _36567_;
wire _36568_;
wire _36569_;
wire _36570_;
wire _36571_;
wire _36572_;
wire _36573_;
wire _36574_;
wire _36575_;
wire _36576_;
wire _36577_;
wire _36578_;
wire _36579_;
wire _36580_;
wire _36581_;
wire _36582_;
wire _36583_;
wire _36584_;
wire _36585_;
wire _36586_;
wire _36587_;
wire _36588_;
wire _36589_;
wire _36590_;
wire _36591_;
wire _36592_;
wire _36593_;
wire _36594_;
wire _36595_;
wire _36596_;
wire _36597_;
wire _36598_;
wire _36599_;
wire _36600_;
wire _36601_;
wire _36602_;
wire _36603_;
wire _36604_;
wire _36605_;
wire _36606_;
wire _36607_;
wire _36608_;
wire _36609_;
wire _36610_;
wire _36611_;
wire _36612_;
wire _36613_;
wire _36614_;
wire _36615_;
wire _36616_;
wire _36617_;
wire _36618_;
wire _36619_;
wire _36620_;
wire _36621_;
wire _36622_;
wire _36623_;
wire _36624_;
wire _36625_;
wire _36626_;
wire _36627_;
wire _36628_;
wire _36629_;
wire _36630_;
wire _36631_;
wire _36632_;
wire _36633_;
wire _36634_;
wire _36635_;
wire _36636_;
wire _36637_;
wire _36638_;
wire _36639_;
wire _36640_;
wire _36641_;
wire _36642_;
wire _36643_;
wire _36644_;
wire _36645_;
wire _36646_;
wire _36647_;
wire _36648_;
wire _36649_;
wire _36650_;
wire _36651_;
wire _36652_;
wire _36653_;
wire _36654_;
wire _36655_;
wire _36656_;
wire _36657_;
wire _36658_;
wire _36659_;
wire _36660_;
wire _36661_;
wire _36662_;
wire _36663_;
wire _36664_;
wire _36665_;
wire _36666_;
wire _36667_;
wire _36668_;
wire _36669_;
wire _36670_;
wire _36671_;
wire _36672_;
wire _36673_;
wire _36674_;
wire _36675_;
wire _36676_;
wire _36677_;
wire _36678_;
wire _36679_;
wire _36680_;
wire _36681_;
wire _36682_;
wire _36683_;
wire _36684_;
wire _36685_;
wire _36686_;
wire _36687_;
wire _36688_;
wire _36689_;
wire _36690_;
wire _36691_;
wire _36692_;
wire _36693_;
wire _36694_;
wire _36695_;
wire _36696_;
wire _36697_;
wire _36698_;
wire _36699_;
wire _36700_;
wire _36701_;
wire _36702_;
wire _36703_;
wire _36704_;
wire _36705_;
wire _36706_;
wire _36707_;
wire _36708_;
wire _36709_;
wire _36710_;
wire _36711_;
wire _36712_;
wire _36713_;
wire _36714_;
wire _36715_;
wire _36716_;
wire _36717_;
wire _36718_;
wire _36719_;
wire _36720_;
wire _36721_;
wire _36722_;
wire _36723_;
wire _36724_;
wire _36725_;
wire _36726_;
wire _36727_;
wire _36728_;
wire _36729_;
wire _36730_;
wire _36731_;
wire _36732_;
wire _36733_;
wire _36734_;
wire _36735_;
wire _36736_;
wire _36737_;
wire _36738_;
wire _36739_;
wire _36740_;
wire _36741_;
wire _36742_;
wire _36743_;
wire _36744_;
wire _36745_;
wire _36746_;
wire _36747_;
wire _36748_;
wire _36749_;
wire _36750_;
wire _36751_;
wire _36752_;
wire _36753_;
wire _36754_;
wire _36755_;
wire _36756_;
wire _36757_;
wire _36758_;
wire _36759_;
wire _36760_;
wire _36761_;
wire _36762_;
wire _36763_;
wire _36764_;
wire _36765_;
wire _36766_;
wire _36767_;
wire _36768_;
wire _36769_;
wire _36770_;
wire _36771_;
wire _36772_;
wire _36773_;
wire _36774_;
wire _36775_;
wire _36776_;
wire _36777_;
wire _36778_;
wire _36779_;
wire _36780_;
wire _36781_;
wire _36782_;
wire _36783_;
wire _36784_;
wire _36785_;
wire _36786_;
wire _36787_;
wire _36788_;
wire _36789_;
wire _36790_;
wire _36791_;
wire _36792_;
wire _36793_;
wire _36794_;
wire _36795_;
wire _36796_;
wire _36797_;
wire _36798_;
wire _36799_;
wire _36800_;
wire _36801_;
wire _36802_;
wire _36803_;
wire _36804_;
wire _36805_;
wire _36806_;
wire _36807_;
wire _36808_;
wire _36809_;
wire _36810_;
wire _36811_;
wire _36812_;
wire _36813_;
wire _36814_;
wire _36815_;
wire _36816_;
wire _36817_;
wire _36818_;
wire _36819_;
wire _36820_;
wire _36821_;
wire _36822_;
wire _36823_;
wire _36824_;
wire _36825_;
wire _36826_;
wire _36827_;
wire _36828_;
wire _36829_;
wire _36830_;
wire _36831_;
wire _36832_;
wire _36833_;
wire _36834_;
wire _36835_;
wire _36836_;
wire _36837_;
wire _36838_;
wire _36839_;
wire _36840_;
wire _36841_;
wire _36842_;
wire _36843_;
wire _36844_;
wire _36845_;
wire _36846_;
wire _36847_;
wire _36848_;
wire _36849_;
wire _36850_;
wire _36851_;
wire _36852_;
wire _36853_;
wire _36854_;
wire _36855_;
wire _36856_;
wire _36857_;
wire _36858_;
wire _36859_;
wire _36860_;
wire _36861_;
wire _36862_;
wire _36863_;
wire _36864_;
wire _36865_;
wire _36866_;
wire _36867_;
wire _36868_;
wire _36869_;
wire _36870_;
wire _36871_;
wire _36872_;
wire _36873_;
wire _36874_;
wire _36875_;
wire _36876_;
wire _36877_;
wire _36878_;
wire _36879_;
wire _36880_;
wire _36881_;
wire _36882_;
wire _36883_;
wire _36884_;
wire _36885_;
wire _36886_;
wire _36887_;
wire _36888_;
wire _36889_;
wire _36890_;
wire _36891_;
wire _36892_;
wire _36893_;
wire _36894_;
wire _36895_;
wire _36896_;
wire _36897_;
wire _36898_;
wire _36899_;
wire _36900_;
wire _36901_;
wire _36902_;
wire _36903_;
wire _36904_;
wire _36905_;
wire _36906_;
wire _36907_;
wire _36908_;
wire _36909_;
wire _36910_;
wire _36911_;
wire _36912_;
wire _36913_;
wire _36914_;
wire _36915_;
wire _36916_;
wire _36917_;
wire _36918_;
wire _36919_;
wire _36920_;
wire _36921_;
wire _36922_;
wire _36923_;
wire _36924_;
wire _36925_;
wire _36926_;
wire _36927_;
wire _36928_;
wire _36929_;
wire _36930_;
wire _36931_;
wire _36932_;
wire _36933_;
wire _36934_;
wire _36935_;
wire _36936_;
wire _36937_;
wire _36938_;
wire _36939_;
wire _36940_;
wire _36941_;
wire _36942_;
wire _36943_;
wire _36944_;
wire _36945_;
wire _36946_;
wire _36947_;
wire _36948_;
wire _36949_;
wire _36950_;
wire _36951_;
wire _36952_;
wire _36953_;
wire _36954_;
wire _36955_;
wire _36956_;
wire _36957_;
wire _36958_;
wire _36959_;
wire _36960_;
wire _36961_;
wire _36962_;
wire _36963_;
wire _36964_;
wire _36965_;
wire _36966_;
wire _36967_;
wire _36968_;
wire _36969_;
wire _36970_;
wire _36971_;
wire _36972_;
wire _36973_;
wire _36974_;
wire _36975_;
wire _36976_;
wire _36977_;
wire _36978_;
wire _36979_;
wire _36980_;
wire _36981_;
wire _36982_;
wire _36983_;
wire _36984_;
wire _36985_;
wire _36986_;
wire _36987_;
wire _36988_;
wire _36989_;
wire _36990_;
wire _36991_;
wire _36992_;
wire _36993_;
wire _36994_;
wire _36995_;
wire _36996_;
wire _36997_;
wire _36998_;
wire _36999_;
wire _37000_;
wire _37001_;
wire _37002_;
wire _37003_;
wire _37004_;
wire _37005_;
wire _37006_;
wire _37007_;
wire _37008_;
wire _37009_;
wire _37010_;
wire _37011_;
wire _37012_;
wire _37013_;
wire _37014_;
wire _37015_;
wire _37016_;
wire _37017_;
wire _37018_;
wire _37019_;
wire _37020_;
wire _37021_;
wire _37022_;
wire _37023_;
wire _37024_;
wire _37025_;
wire _37026_;
wire _37027_;
wire _37028_;
wire _37029_;
wire _37030_;
wire _37031_;
wire _37032_;
wire _37033_;
wire _37034_;
wire _37035_;
wire _37036_;
wire _37037_;
wire _37038_;
wire _37039_;
wire _37040_;
wire _37041_;
wire _37042_;
wire _37043_;
wire _37044_;
wire _37045_;
wire _37046_;
wire _37047_;
wire _37048_;
wire _37049_;
wire _37050_;
wire _37051_;
wire _37052_;
wire _37053_;
wire _37054_;
wire _37055_;
wire _37056_;
wire _37057_;
wire _37058_;
wire _37059_;
wire _37060_;
wire _37061_;
wire _37062_;
wire _37063_;
wire _37064_;
wire _37065_;
wire _37066_;
wire _37067_;
wire _37068_;
wire _37069_;
wire _37070_;
wire _37071_;
wire _37072_;
wire _37073_;
wire _37074_;
wire _37075_;
wire _37076_;
wire _37077_;
wire _37078_;
wire _37079_;
wire _37080_;
wire _37081_;
wire _37082_;
wire _37083_;
wire _37084_;
wire _37085_;
wire _37086_;
wire _37087_;
wire _37088_;
wire _37089_;
wire _37090_;
wire _37091_;
wire _37092_;
wire _37093_;
wire _37094_;
wire _37095_;
wire _37096_;
wire _37097_;
wire _37098_;
wire _37099_;
wire _37100_;
wire _37101_;
wire _37102_;
wire _37103_;
wire _37104_;
wire _37105_;
wire _37106_;
wire _37107_;
wire _37108_;
wire _37109_;
wire _37110_;
wire _37111_;
wire _37112_;
wire _37113_;
wire _37114_;
wire _37115_;
wire _37116_;
wire _37117_;
wire _37118_;
wire _37119_;
wire _37120_;
wire _37121_;
wire _37122_;
wire _37123_;
wire _37124_;
wire _37125_;
wire _37126_;
wire _37127_;
wire _37128_;
wire _37129_;
wire _37130_;
wire _37131_;
wire _37132_;
wire _37133_;
wire _37134_;
wire _37135_;
wire _37136_;
wire _37137_;
wire _37138_;
wire _37139_;
wire _37140_;
wire _37141_;
wire _37142_;
wire _37143_;
wire _37144_;
wire _37145_;
wire _37146_;
wire _37147_;
wire _37148_;
wire _37149_;
wire _37150_;
wire _37151_;
wire _37152_;
wire _37153_;
wire _37154_;
wire _37155_;
wire _37156_;
wire _37157_;
wire _37158_;
wire _37159_;
wire _37160_;
wire _37161_;
wire _37162_;
wire _37163_;
wire _37164_;
wire _37165_;
wire _37166_;
wire _37167_;
wire _37168_;
wire _37169_;
wire _37170_;
wire _37171_;
wire _37172_;
wire _37173_;
wire _37174_;
wire _37175_;
wire _37176_;
wire _37177_;
wire _37178_;
wire _37179_;
wire _37180_;
wire _37181_;
wire _37182_;
wire _37183_;
wire _37184_;
wire _37185_;
wire _37186_;
wire _37187_;
wire _37188_;
wire _37189_;
wire _37190_;
wire _37191_;
wire _37192_;
wire _37193_;
wire _37194_;
wire _37195_;
wire _37196_;
wire _37197_;
wire _37198_;
wire _37199_;
wire _37200_;
wire _37201_;
wire _37202_;
wire _37203_;
wire _37204_;
wire _37205_;
wire _37206_;
wire _37207_;
wire _37208_;
wire _37209_;
wire _37210_;
wire _37211_;
wire _37212_;
wire _37213_;
wire _37214_;
wire _37215_;
wire _37216_;
wire _37217_;
wire _37218_;
wire _37219_;
wire _37220_;
wire _37221_;
wire _37222_;
wire _37223_;
wire _37224_;
wire _37225_;
wire _37226_;
wire _37227_;
wire _37228_;
wire _37229_;
wire _37230_;
wire _37231_;
wire _37232_;
wire _37233_;
wire _37234_;
wire _37235_;
wire _37236_;
wire _37237_;
wire _37238_;
wire _37239_;
wire _37240_;
wire _37241_;
wire _37242_;
wire _37243_;
wire _37244_;
wire _37245_;
wire _37246_;
wire _37247_;
wire _37248_;
wire _37249_;
wire _37250_;
wire _37251_;
wire _37252_;
wire _37253_;
wire _37254_;
wire _37255_;
wire _37256_;
wire _37257_;
wire _37258_;
wire _37259_;
wire _37260_;
wire _37261_;
wire _37262_;
wire _37263_;
wire _37264_;
wire _37265_;
wire _37266_;
wire _37267_;
wire _37268_;
wire _37269_;
wire _37270_;
wire _37271_;
wire _37272_;
wire _37273_;
wire _37274_;
wire _37275_;
wire _37276_;
wire _37277_;
wire _37278_;
wire _37279_;
wire _37280_;
wire _37281_;
wire _37282_;
wire _37283_;
wire _37284_;
wire _37285_;
wire _37286_;
wire _37287_;
wire _37288_;
wire _37289_;
wire _37290_;
wire _37291_;
wire _37292_;
wire _37293_;
wire _37294_;
wire _37295_;
wire _37296_;
wire _37297_;
wire _37298_;
wire _37299_;
wire _37300_;
wire _37301_;
wire _37302_;
wire _37303_;
wire _37304_;
wire _37305_;
wire _37306_;
wire _37307_;
wire _37308_;
wire _37309_;
wire _37310_;
wire _37311_;
wire _37312_;
wire _37313_;
wire _37314_;
wire _37315_;
wire _37316_;
wire _37317_;
wire _37318_;
wire _37319_;
wire _37320_;
wire _37321_;
wire _37322_;
wire _37323_;
wire _37324_;
wire _37325_;
wire _37326_;
wire _37327_;
wire _37328_;
wire _37329_;
wire _37330_;
wire _37331_;
wire _37332_;
wire _37333_;
wire _37334_;
wire _37335_;
wire _37336_;
wire _37337_;
wire _37338_;
wire _37339_;
wire _37340_;
wire _37341_;
wire _37342_;
wire _37343_;
wire _37344_;
wire _37345_;
wire _37346_;
wire _37347_;
wire _37348_;
wire _37349_;
wire _37350_;
wire _37351_;
wire _37352_;
wire _37353_;
wire _37354_;
wire _37355_;
wire _37356_;
wire _37357_;
wire _37358_;
wire _37359_;
wire _37360_;
wire _37361_;
wire _37362_;
wire _37363_;
wire _37364_;
wire _37365_;
wire _37366_;
wire _37367_;
wire _37368_;
wire _37369_;
wire _37370_;
wire _37371_;
wire _37372_;
wire _37373_;
wire _37374_;
wire _37375_;
wire _37376_;
wire _37377_;
wire _37378_;
wire _37379_;
wire _37380_;
wire _37381_;
wire _37382_;
wire _37383_;
wire _37384_;
wire _37385_;
wire _37386_;
wire _37387_;
wire _37388_;
wire _37389_;
wire _37390_;
wire _37391_;
wire _37392_;
wire _37393_;
wire _37394_;
wire _37395_;
wire _37396_;
wire _37397_;
wire _37398_;
wire _37399_;
wire _37400_;
wire _37401_;
wire _37402_;
wire _37403_;
wire _37404_;
wire _37405_;
wire _37406_;
wire _37407_;
wire _37408_;
wire _37409_;
wire _37410_;
wire _37411_;
wire _37412_;
wire _37413_;
wire _37414_;
wire _37415_;
wire _37416_;
wire _37417_;
wire _37418_;
wire _37419_;
wire _37420_;
wire _37421_;
wire _37422_;
wire _37423_;
wire _37424_;
wire _37425_;
wire _37426_;
wire _37427_;
wire _37428_;
wire _37429_;
wire _37430_;
wire _37431_;
wire _37432_;
wire _37433_;
wire _37434_;
wire _37435_;
wire _37436_;
wire _37437_;
wire _37438_;
wire _37439_;
wire _37440_;
wire _37441_;
wire _37442_;
wire _37443_;
wire _37444_;
wire _37445_;
wire _37446_;
wire _37447_;
wire _37448_;
wire _37449_;
wire _37450_;
wire _37451_;
wire _37452_;
wire _37453_;
wire _37454_;
wire _37455_;
wire _37456_;
wire _37457_;
wire _37458_;
wire _37459_;
wire _37460_;
wire _37461_;
wire _37462_;
wire _37463_;
wire _37464_;
wire _37465_;
wire _37466_;
wire _37467_;
wire _37468_;
wire _37469_;
wire _37470_;
wire _37471_;
wire _37472_;
wire _37473_;
wire _37474_;
wire _37475_;
wire _37476_;
wire _37477_;
wire _37478_;
wire _37479_;
wire _37480_;
wire _37481_;
wire _37482_;
wire _37483_;
wire _37484_;
wire _37485_;
wire _37486_;
wire _37487_;
wire _37488_;
wire _37489_;
wire _37490_;
wire _37491_;
wire _37492_;
wire _37493_;
wire _37494_;
wire _37495_;
wire _37496_;
wire _37497_;
wire _37498_;
wire _37499_;
wire _37500_;
wire _37501_;
wire _37502_;
wire _37503_;
wire _37504_;
wire _37505_;
wire _37506_;
wire _37507_;
wire _37508_;
wire _37509_;
wire _37510_;
wire _37511_;
wire _37512_;
wire _37513_;
wire _37514_;
wire _37515_;
wire _37516_;
wire _37517_;
wire _37518_;
wire _37519_;
wire _37520_;
wire _37521_;
wire _37522_;
wire _37523_;
wire _37524_;
wire _37525_;
wire _37526_;
wire _37527_;
wire _37528_;
wire _37529_;
wire _37530_;
wire _37531_;
wire _37532_;
wire _37533_;
wire _37534_;
wire _37535_;
wire _37536_;
wire _37537_;
wire _37538_;
wire _37539_;
wire _37540_;
wire _37541_;
wire _37542_;
wire _37543_;
wire _37544_;
wire _37545_;
wire _37546_;
wire _37547_;
wire _37548_;
wire _37549_;
wire _37550_;
wire _37551_;
wire _37552_;
wire _37553_;
wire _37554_;
wire _37555_;
wire _37556_;
wire _37557_;
wire _37558_;
wire _37559_;
wire _37560_;
wire _37561_;
wire _37562_;
wire _37563_;
wire _37564_;
wire _37565_;
wire _37566_;
wire _37567_;
wire _37568_;
wire _37569_;
wire _37570_;
wire _37571_;
wire _37572_;
wire _37573_;
wire _37574_;
wire _37575_;
wire _37576_;
wire _37577_;
wire _37578_;
wire _37579_;
wire _37580_;
wire _37581_;
wire _37582_;
wire _37583_;
wire _37584_;
wire _37585_;
wire _37586_;
wire _37587_;
wire _37588_;
wire _37589_;
wire _37590_;
wire _37591_;
wire _37592_;
wire _37593_;
wire _37594_;
wire _37595_;
wire _37596_;
wire _37597_;
wire _37598_;
wire _37599_;
wire _37600_;
wire _37601_;
wire _37602_;
wire _37603_;
wire _37604_;
wire _37605_;
wire _37606_;
wire _37607_;
wire _37608_;
wire _37609_;
wire _37610_;
wire _37611_;
wire _37612_;
wire _37613_;
wire _37614_;
wire _37615_;
wire _37616_;
wire _37617_;
wire _37618_;
wire _37619_;
wire _37620_;
wire _37621_;
wire _37622_;
wire _37623_;
wire _37624_;
wire _37625_;
wire _37626_;
wire _37627_;
wire _37628_;
wire _37629_;
wire _37630_;
wire _37631_;
wire _37632_;
wire _37633_;
wire _37634_;
wire _37635_;
wire _37636_;
wire _37637_;
wire _37638_;
wire _37639_;
wire _37640_;
wire _37641_;
wire _37642_;
wire _37643_;
wire _37644_;
wire _37645_;
wire _37646_;
wire _37647_;
wire _37648_;
wire _37649_;
wire _37650_;
wire _37651_;
wire _37652_;
wire _37653_;
wire _37654_;
wire _37655_;
wire _37656_;
wire _37657_;
wire _37658_;
wire _37659_;
wire _37660_;
wire _37661_;
wire _37662_;
wire _37663_;
wire _37664_;
wire _37665_;
wire _37666_;
wire _37667_;
wire _37668_;
wire _37669_;
wire _37670_;
wire _37671_;
wire _37672_;
wire _37673_;
wire _37674_;
wire _37675_;
wire _37676_;
wire _37677_;
wire _37678_;
wire _37679_;
wire _37680_;
wire _37681_;
wire _37682_;
wire _37683_;
wire _37684_;
wire _37685_;
wire _37686_;
wire _37687_;
wire _37688_;
wire _37689_;
wire _37690_;
wire _37691_;
wire _37692_;
wire _37693_;
wire _37694_;
wire _37695_;
wire _37696_;
wire _37697_;
wire _37698_;
wire _37699_;
wire _37700_;
wire _37701_;
wire _37702_;
wire _37703_;
wire _37704_;
wire _37705_;
wire _37706_;
wire _37707_;
wire _37708_;
wire _37709_;
wire _37710_;
wire _37711_;
wire _37712_;
wire _37713_;
wire _37714_;
wire _37715_;
wire _37716_;
wire _37717_;
wire _37718_;
wire _37719_;
wire _37720_;
wire _37721_;
wire _37722_;
wire _37723_;
wire _37724_;
wire _37725_;
wire _37726_;
wire _37727_;
wire _37728_;
wire _37729_;
wire _37730_;
wire _37731_;
wire _37732_;
wire _37733_;
wire _37734_;
wire _37735_;
wire _37736_;
wire _37737_;
wire _37738_;
wire _37739_;
wire _37740_;
wire _37741_;
wire _37742_;
wire _37743_;
wire _37744_;
wire _37745_;
wire _37746_;
wire _37747_;
wire _37748_;
wire _37749_;
wire _37750_;
wire _37751_;
wire _37752_;
wire _37753_;
wire _37754_;
wire _37755_;
wire _37756_;
wire _37757_;
wire _37758_;
wire _37759_;
wire _37760_;
wire _37761_;
wire _37762_;
wire _37763_;
wire _37764_;
wire _37765_;
wire _37766_;
wire _37767_;
wire _37768_;
wire _37769_;
wire _37770_;
wire _37771_;
wire _37772_;
wire _37773_;
wire _37774_;
wire _37775_;
wire _37776_;
wire _37777_;
wire _37778_;
wire _37779_;
wire _37780_;
wire _37781_;
wire _37782_;
wire _37783_;
wire _37784_;
wire _37785_;
wire _37786_;
wire _37787_;
wire _37788_;
wire _37789_;
wire _37790_;
wire _37791_;
wire _37792_;
wire _37793_;
wire _37794_;
wire _37795_;
wire _37796_;
wire _37797_;
wire _37798_;
wire _37799_;
wire _37800_;
wire _37801_;
wire _37802_;
wire _37803_;
wire _37804_;
wire _37805_;
wire _37806_;
wire _37807_;
wire _37808_;
wire _37809_;
wire _37810_;
wire _37811_;
wire _37812_;
wire _37813_;
wire _37814_;
wire _37815_;
wire _37816_;
wire _37817_;
wire _37818_;
wire _37819_;
wire _37820_;
wire _37821_;
wire _37822_;
wire _37823_;
wire _37824_;
wire _37825_;
wire _37826_;
wire _37827_;
wire _37828_;
wire _37829_;
wire _37830_;
wire _37831_;
wire _37832_;
wire _37833_;
wire _37834_;
wire _37835_;
wire _37836_;
wire _37837_;
wire _37838_;
wire _37839_;
wire _37840_;
wire _37841_;
wire _37842_;
wire _37843_;
wire _37844_;
wire _37845_;
wire _37846_;
wire _37847_;
wire _37848_;
wire _37849_;
wire _37850_;
wire _37851_;
wire _37852_;
wire _37853_;
wire _37854_;
wire _37855_;
wire _37856_;
wire _37857_;
wire _37858_;
wire _37859_;
wire _37860_;
wire _37861_;
wire _37862_;
wire _37863_;
wire _37864_;
wire _37865_;
wire _37866_;
wire _37867_;
wire _37868_;
wire _37869_;
wire _37870_;
wire _37871_;
wire _37872_;
wire _37873_;
wire _37874_;
wire _37875_;
wire _37876_;
wire _37877_;
wire _37878_;
wire _37879_;
wire _37880_;
wire _37881_;
wire _37882_;
wire _37883_;
wire _37884_;
wire _37885_;
wire _37886_;
wire _37887_;
wire _37888_;
wire _37889_;
wire _37890_;
wire _37891_;
wire _37892_;
wire _37893_;
wire _37894_;
wire _37895_;
wire _37896_;
wire _37897_;
wire _37898_;
wire _37899_;
wire _37900_;
wire _37901_;
wire _37902_;
wire _37903_;
wire _37904_;
wire _37905_;
wire _37906_;
wire _37907_;
wire _37908_;
wire _37909_;
wire _37910_;
wire _37911_;
wire _37912_;
wire _37913_;
wire _37914_;
wire _37915_;
wire _37916_;
wire _37917_;
wire _37918_;
wire _37919_;
wire _37920_;
wire _37921_;
wire _37922_;
wire _37923_;
wire _37924_;
wire _37925_;
wire _37926_;
wire _37927_;
wire _37928_;
wire _37929_;
wire _37930_;
wire _37931_;
wire _37932_;
wire _37933_;
wire _37934_;
wire _37935_;
wire _37936_;
wire _37937_;
wire _37938_;
wire _37939_;
wire _37940_;
wire _37941_;
wire _37942_;
wire _37943_;
wire _37944_;
wire _37945_;
wire _37946_;
wire _37947_;
wire _37948_;
wire _37949_;
wire _37950_;
wire _37951_;
wire _37952_;
wire _37953_;
wire _37954_;
wire _37955_;
wire _37956_;
wire _37957_;
wire _37958_;
wire _37959_;
wire _37960_;
wire _37961_;
wire _37962_;
wire _37963_;
wire _37964_;
wire _37965_;
wire _37966_;
wire _37967_;
wire _37968_;
wire _37969_;
wire _37970_;
wire _37971_;
wire _37972_;
wire _37973_;
wire _37974_;
wire _37975_;
wire _37976_;
wire _37977_;
wire _37978_;
wire _37979_;
wire _37980_;
wire _37981_;
wire _37982_;
wire _37983_;
wire _37984_;
wire _37985_;
wire _37986_;
wire _37987_;
wire _37988_;
wire _37989_;
wire _37990_;
wire _37991_;
wire _37992_;
wire _37993_;
wire _37994_;
wire _37995_;
wire _37996_;
wire _37997_;
wire _37998_;
wire _37999_;
wire _38000_;
wire _38001_;
wire _38002_;
wire _38003_;
wire _38004_;
wire _38005_;
wire _38006_;
wire _38007_;
wire _38008_;
wire _38009_;
wire _38010_;
wire _38011_;
wire _38012_;
wire _38013_;
wire _38014_;
wire _38015_;
wire _38016_;
wire _38017_;
wire _38018_;
wire _38019_;
wire _38020_;
wire _38021_;
wire _38022_;
wire _38023_;
wire _38024_;
wire _38025_;
wire _38026_;
wire _38027_;
wire _38028_;
wire _38029_;
wire _38030_;
wire _38031_;
wire _38032_;
wire _38033_;
wire _38034_;
wire _38035_;
wire _38036_;
wire _38037_;
wire _38038_;
wire _38039_;
wire _38040_;
wire _38041_;
wire _38042_;
wire _38043_;
wire _38044_;
wire _38045_;
wire _38046_;
wire _38047_;
wire _38048_;
wire _38049_;
wire _38050_;
wire _38051_;
wire _38052_;
wire _38053_;
wire _38054_;
wire _38055_;
wire _38056_;
wire _38057_;
wire _38058_;
wire _38059_;
wire _38060_;
wire _38061_;
wire _38062_;
wire _38063_;
wire _38064_;
wire _38065_;
wire _38066_;
wire _38067_;
wire _38068_;
wire _38069_;
wire _38070_;
wire _38071_;
wire _38072_;
wire _38073_;
wire _38074_;
wire _38075_;
wire _38076_;
wire _38077_;
wire _38078_;
wire _38079_;
wire _38080_;
wire _38081_;
wire _38082_;
wire _38083_;
wire _38084_;
wire _38085_;
wire _38086_;
wire _38087_;
wire _38088_;
wire _38089_;
wire _38090_;
wire _38091_;
wire _38092_;
wire _38093_;
wire _38094_;
wire _38095_;
wire _38096_;
wire _38097_;
wire _38098_;
wire _38099_;
wire _38100_;
wire _38101_;
wire _38102_;
wire _38103_;
wire _38104_;
wire _38105_;
wire _38106_;
wire _38107_;
wire _38108_;
wire _38109_;
wire _38110_;
wire _38111_;
wire _38112_;
wire _38113_;
wire _38114_;
wire _38115_;
wire _38116_;
wire _38117_;
wire _38118_;
wire _38119_;
wire _38120_;
wire _38121_;
wire _38122_;
wire _38123_;
wire _38124_;
wire _38125_;
wire _38126_;
wire _38127_;
wire _38128_;
wire _38129_;
wire _38130_;
wire _38131_;
wire _38132_;
wire _38133_;
wire _38134_;
wire _38135_;
wire _38136_;
wire _38137_;
wire _38138_;
wire _38139_;
wire _38140_;
wire _38141_;
wire _38142_;
wire _38143_;
wire _38144_;
wire _38145_;
wire _38146_;
wire _38147_;
wire _38148_;
wire _38149_;
wire _38150_;
wire _38151_;
wire _38152_;
wire _38153_;
wire _38154_;
wire _38155_;
wire _38156_;
wire _38157_;
wire _38158_;
wire _38159_;
wire _38160_;
wire _38161_;
wire _38162_;
wire _38163_;
wire _38164_;
wire _38165_;
wire _38166_;
wire _38167_;
wire _38168_;
wire _38169_;
wire _38170_;
wire _38171_;
wire _38172_;
wire _38173_;
wire _38174_;
wire _38175_;
wire _38176_;
wire _38177_;
wire _38178_;
wire _38179_;
wire _38180_;
wire _38181_;
wire _38182_;
wire _38183_;
wire _38184_;
wire _38185_;
wire _38186_;
wire _38187_;
wire _38188_;
wire _38189_;
wire _38190_;
wire _38191_;
wire _38192_;
wire _38193_;
wire _38194_;
wire _38195_;
wire _38196_;
wire _38197_;
wire _38198_;
wire _38199_;
wire _38200_;
wire _38201_;
wire _38202_;
wire _38203_;
wire _38204_;
wire _38205_;
wire _38206_;
wire _38207_;
wire _38208_;
wire _38209_;
wire _38210_;
wire _38211_;
wire _38212_;
wire _38213_;
wire _38214_;
wire _38215_;
wire _38216_;
wire _38217_;
wire _38218_;
wire _38219_;
wire _38220_;
wire _38221_;
wire _38222_;
wire _38223_;
wire _38224_;
wire _38225_;
wire _38226_;
wire _38227_;
wire _38228_;
wire _38229_;
wire _38230_;
wire _38231_;
wire _38232_;
wire _38233_;
wire _38234_;
wire _38235_;
wire _38236_;
wire _38237_;
wire _38238_;
wire _38239_;
wire _38240_;
wire _38241_;
wire _38242_;
wire _38243_;
wire _38244_;
wire _38245_;
wire _38246_;
wire _38247_;
wire _38248_;
wire _38249_;
wire _38250_;
wire _38251_;
wire _38252_;
wire _38253_;
wire _38254_;
wire _38255_;
wire _38256_;
wire _38257_;
wire _38258_;
wire _38259_;
wire _38260_;
wire _38261_;
wire _38262_;
wire _38263_;
wire _38264_;
wire _38265_;
wire _38266_;
wire _38267_;
wire _38268_;
wire _38269_;
wire _38270_;
wire _38271_;
wire _38272_;
wire _38273_;
wire _38274_;
wire _38275_;
wire _38276_;
wire _38277_;
wire _38278_;
wire _38279_;
wire _38280_;
wire _38281_;
wire _38282_;
wire _38283_;
wire _38284_;
wire _38285_;
wire _38286_;
wire _38287_;
wire _38288_;
wire _38289_;
wire _38290_;
wire _38291_;
wire _38292_;
wire _38293_;
wire _38294_;
wire _38295_;
wire _38296_;
wire _38297_;
wire _38298_;
wire _38299_;
wire _38300_;
wire _38301_;
wire _38302_;
wire _38303_;
wire _38304_;
wire _38305_;
wire _38306_;
wire _38307_;
wire _38308_;
wire _38309_;
wire _38310_;
wire _38311_;
wire _38312_;
wire _38313_;
wire _38314_;
wire _38315_;
wire _38316_;
wire _38317_;
wire _38318_;
wire _38319_;
wire _38320_;
wire _38321_;
wire _38322_;
wire _38323_;
wire _38324_;
wire _38325_;
wire _38326_;
wire _38327_;
wire _38328_;
wire _38329_;
wire _38330_;
wire _38331_;
wire _38332_;
wire _38333_;
wire _38334_;
wire _38335_;
wire _38336_;
wire _38337_;
wire _38338_;
wire _38339_;
wire _38340_;
wire _38341_;
wire _38342_;
wire _38343_;
wire _38344_;
wire _38345_;
wire _38346_;
wire _38347_;
wire _38348_;
wire _38349_;
wire _38350_;
wire _38351_;
wire _38352_;
wire _38353_;
wire _38354_;
wire _38355_;
wire _38356_;
wire _38357_;
wire _38358_;
wire _38359_;
wire _38360_;
wire _38361_;
wire _38362_;
wire _38363_;
wire _38364_;
wire _38365_;
wire _38366_;
wire _38367_;
wire _38368_;
wire _38369_;
wire _38370_;
wire _38371_;
wire _38372_;
wire _38373_;
wire _38374_;
wire _38375_;
wire _38376_;
wire _38377_;
wire _38378_;
wire _38379_;
wire _38380_;
wire _38381_;
wire _38382_;
wire _38383_;
wire _38384_;
wire _38385_;
wire _38386_;
wire _38387_;
wire _38388_;
wire _38389_;
wire _38390_;
wire _38391_;
wire _38392_;
wire _38393_;
wire _38394_;
wire _38395_;
wire _38396_;
wire _38397_;
wire _38398_;
wire _38399_;
wire _38400_;
wire _38401_;
wire _38402_;
wire _38403_;
wire _38404_;
wire _38405_;
wire _38406_;
wire _38407_;
wire _38408_;
wire _38409_;
wire _38410_;
wire _38411_;
wire _38412_;
wire _38413_;
wire _38414_;
wire _38415_;
wire _38416_;
wire _38417_;
wire _38418_;
wire _38419_;
wire _38420_;
wire _38421_;
wire _38422_;
wire _38423_;
wire _38424_;
wire _38425_;
wire _38426_;
wire _38427_;
wire _38428_;
wire _38429_;
wire _38430_;
wire _38431_;
wire _38432_;
wire _38433_;
wire _38434_;
wire _38435_;
wire _38436_;
wire _38437_;
wire _38438_;
wire _38439_;
wire _38440_;
wire _38441_;
wire _38442_;
wire _38443_;
wire _38444_;
wire _38445_;
wire _38446_;
wire _38447_;
wire _38448_;
wire _38449_;
wire _38450_;
wire _38451_;
wire _38452_;
wire _38453_;
wire _38454_;
wire _38455_;
wire _38456_;
wire _38457_;
wire _38458_;
wire _38459_;
wire _38460_;
wire _38461_;
wire _38462_;
wire _38463_;
wire _38464_;
wire _38465_;
wire _38466_;
wire _38467_;
wire _38468_;
wire _38469_;
wire _38470_;
wire _38471_;
wire _38472_;
wire _38473_;
wire _38474_;
wire _38475_;
wire _38476_;
wire _38477_;
wire _38478_;
wire _38479_;
wire _38480_;
wire _38481_;
wire _38482_;
wire _38483_;
wire _38484_;
wire _38485_;
wire _38486_;
wire _38487_;
wire _38488_;
wire _38489_;
wire _38490_;
wire _38491_;
wire _38492_;
wire _38493_;
wire _38494_;
wire _38495_;
wire _38496_;
wire _38497_;
wire _38498_;
wire _38499_;
wire _38500_;
wire _38501_;
wire _38502_;
wire _38503_;
wire _38504_;
wire _38505_;
wire _38506_;
wire _38507_;
wire _38508_;
wire _38509_;
wire _38510_;
wire _38511_;
wire _38512_;
wire _38513_;
wire _38514_;
wire _38515_;
wire _38516_;
wire _38517_;
wire _38518_;
wire _38519_;
wire _38520_;
wire _38521_;
wire _38522_;
wire _38523_;
wire _38524_;
wire _38525_;
wire _38526_;
wire _38527_;
wire _38528_;
wire _38529_;
wire _38530_;
wire _38531_;
wire _38532_;
wire _38533_;
wire _38534_;
wire _38535_;
wire _38536_;
wire _38537_;
wire _38538_;
wire _38539_;
wire _38540_;
wire _38541_;
wire _38542_;
wire _38543_;
wire _38544_;
wire _38545_;
wire _38546_;
wire _38547_;
wire _38548_;
wire _38549_;
wire _38550_;
wire _38551_;
wire _38552_;
wire _38553_;
wire _38554_;
wire _38555_;
wire _38556_;
wire _38557_;
wire _38558_;
wire _38559_;
wire _38560_;
wire _38561_;
wire _38562_;
wire _38563_;
wire _38564_;
wire _38565_;
wire _38566_;
wire _38567_;
wire _38568_;
wire _38569_;
wire _38570_;
wire _38571_;
wire _38572_;
wire _38573_;
wire _38574_;
wire _38575_;
wire _38576_;
wire _38577_;
wire _38578_;
wire _38579_;
wire _38580_;
wire _38581_;
wire _38582_;
wire _38583_;
wire _38584_;
wire _38585_;
wire _38586_;
wire _38587_;
wire _38588_;
wire _38589_;
wire _38590_;
wire _38591_;
wire _38592_;
wire _38593_;
wire _38594_;
wire _38595_;
wire _38596_;
wire _38597_;
wire _38598_;
wire _38599_;
wire _38600_;
wire _38601_;
wire _38602_;
wire _38603_;
wire _38604_;
wire _38605_;
wire _38606_;
wire _38607_;
wire _38608_;
wire _38609_;
wire _38610_;
wire _38611_;
wire _38612_;
wire _38613_;
wire _38614_;
wire _38615_;
wire _38616_;
wire _38617_;
wire _38618_;
wire _38619_;
wire _38620_;
wire _38621_;
wire _38622_;
wire _38623_;
wire _38624_;
wire _38625_;
wire _38626_;
wire _38627_;
wire _38628_;
wire _38629_;
wire _38630_;
wire _38631_;
wire _38632_;
wire _38633_;
wire _38634_;
wire _38635_;
wire _38636_;
wire _38637_;
wire _38638_;
wire _38639_;
wire _38640_;
wire _38641_;
wire _38642_;
wire _38643_;
wire _38644_;
wire _38645_;
wire _38646_;
wire _38647_;
wire _38648_;
wire _38649_;
wire _38650_;
wire _38651_;
wire _38652_;
wire _38653_;
wire _38654_;
wire _38655_;
wire _38656_;
wire _38657_;
wire _38658_;
wire _38659_;
wire _38660_;
wire _38661_;
wire _38662_;
wire _38663_;
wire _38664_;
wire _38665_;
wire _38666_;
wire _38667_;
wire _38668_;
wire _38669_;
wire _38670_;
wire _38671_;
wire _38672_;
wire _38673_;
wire _38674_;
wire _38675_;
wire _38676_;
wire _38677_;
wire _38678_;
wire _38679_;
wire _38680_;
wire _38681_;
wire _38682_;
wire _38683_;
wire _38684_;
wire _38685_;
wire _38686_;
wire _38687_;
wire _38688_;
wire _38689_;
wire _38690_;
wire _38691_;
wire _38692_;
wire _38693_;
wire _38694_;
wire _38695_;
wire _38696_;
wire _38697_;
wire _38698_;
wire _38699_;
wire _38700_;
wire _38701_;
wire _38702_;
wire _38703_;
wire _38704_;
wire _38705_;
wire _38706_;
wire _38707_;
wire _38708_;
wire _38709_;
wire _38710_;
wire _38711_;
wire _38712_;
wire _38713_;
wire _38714_;
wire _38715_;
wire _38716_;
wire _38717_;
wire _38718_;
wire _38719_;
wire _38720_;
wire _38721_;
wire _38722_;
wire _38723_;
wire _38724_;
wire _38725_;
wire _38726_;
wire _38727_;
wire _38728_;
wire _38729_;
wire _38730_;
wire _38731_;
wire _38732_;
wire _38733_;
wire _38734_;
wire _38735_;
wire _38736_;
wire _38737_;
wire _38738_;
wire _38739_;
wire _38740_;
wire _38741_;
wire _38742_;
wire _38743_;
wire _38744_;
wire _38745_;
wire _38746_;
wire _38747_;
wire _38748_;
wire _38749_;
wire _38750_;
wire _38751_;
wire _38752_;
wire _38753_;
wire _38754_;
wire _38755_;
wire _38756_;
wire _38757_;
wire _38758_;
wire _38759_;
wire _38760_;
wire _38761_;
wire _38762_;
wire _38763_;
wire _38764_;
wire _38765_;
wire _38766_;
wire _38767_;
wire _38768_;
wire _38769_;
wire _38770_;
wire _38771_;
wire _38772_;
wire _38773_;
wire _38774_;
wire _38775_;
wire _38776_;
wire _38777_;
wire _38778_;
wire _38779_;
wire _38780_;
wire _38781_;
wire _38782_;
wire _38783_;
wire _38784_;
wire _38785_;
wire _38786_;
wire _38787_;
wire _38788_;
wire _38789_;
wire _38790_;
wire _38791_;
wire _38792_;
wire _38793_;
wire _38794_;
wire _38795_;
wire _38796_;
wire _38797_;
wire _38798_;
wire _38799_;
wire _38800_;
wire _38801_;
wire _38802_;
wire _38803_;
wire _38804_;
wire _38805_;
wire _38806_;
wire _38807_;
wire _38808_;
wire _38809_;
wire _38810_;
wire _38811_;
wire _38812_;
wire _38813_;
wire _38814_;
wire _38815_;
wire _38816_;
wire _38817_;
wire _38818_;
wire _38819_;
wire _38820_;
wire _38821_;
wire _38822_;
wire _38823_;
wire _38824_;
wire _38825_;
wire _38826_;
wire _38827_;
wire _38828_;
wire _38829_;
wire _38830_;
wire _38831_;
wire _38832_;
wire _38833_;
wire _38834_;
wire _38835_;
wire _38836_;
wire _38837_;
wire _38838_;
wire _38839_;
wire _38840_;
wire _38841_;
wire _38842_;
wire _38843_;
wire _38844_;
wire _38845_;
wire _38846_;
wire _38847_;
wire _38848_;
wire _38849_;
wire _38850_;
wire _38851_;
wire _38852_;
wire _38853_;
wire _38854_;
wire _38855_;
wire _38856_;
wire _38857_;
wire _38858_;
wire _38859_;
wire _38860_;
wire _38861_;
wire _38862_;
wire _38863_;
wire _38864_;
wire _38865_;
wire _38866_;
wire _38867_;
wire _38868_;
wire _38869_;
wire _38870_;
wire _38871_;
wire _38872_;
wire _38873_;
wire _38874_;
wire _38875_;
wire _38876_;
wire _38877_;
wire _38878_;
wire _38879_;
wire _38880_;
wire _38881_;
wire _38882_;
wire _38883_;
wire _38884_;
wire _38885_;
wire _38886_;
wire _38887_;
wire _38888_;
wire _38889_;
wire _38890_;
wire _38891_;
wire _38892_;
wire _38893_;
wire _38894_;
wire _38895_;
wire _38896_;
wire _38897_;
wire _38898_;
wire _38899_;
wire _38900_;
wire _38901_;
wire _38902_;
wire _38903_;
wire _38904_;
wire _38905_;
wire _38906_;
wire _38907_;
wire _38908_;
wire _38909_;
wire _38910_;
wire _38911_;
wire _38912_;
wire _38913_;
wire _38914_;
wire _38915_;
wire _38916_;
wire _38917_;
wire _38918_;
wire _38919_;
wire _38920_;
wire _38921_;
wire _38922_;
wire _38923_;
wire _38924_;
wire _38925_;
wire _38926_;
wire _38927_;
wire _38928_;
wire _38929_;
wire _38930_;
wire _38931_;
wire _38932_;
wire _38933_;
wire _38934_;
wire _38935_;
wire _38936_;
wire _38937_;
wire _38938_;
wire _38939_;
wire _38940_;
wire _38941_;
wire _38942_;
wire _38943_;
wire _38944_;
wire _38945_;
wire _38946_;
wire _38947_;
wire _38948_;
wire _38949_;
wire _38950_;
wire _38951_;
wire _38952_;
wire _38953_;
wire _38954_;
wire _38955_;
wire _38956_;
wire _38957_;
wire _38958_;
wire _38959_;
wire _38960_;
wire _38961_;
wire _38962_;
wire _38963_;
wire _38964_;
wire _38965_;
wire _38966_;
wire _38967_;
wire _38968_;
wire _38969_;
wire _38970_;
wire _38971_;
wire _38972_;
wire _38973_;
wire _38974_;
wire _38975_;
wire _38976_;
wire _38977_;
wire _38978_;
wire _38979_;
wire _38980_;
wire _38981_;
wire _38982_;
wire _38983_;
wire _38984_;
wire _38985_;
wire _38986_;
wire _38987_;
wire _38988_;
wire _38989_;
wire _38990_;
wire _38991_;
wire _38992_;
wire _38993_;
wire _38994_;
wire _38995_;
wire _38996_;
wire _38997_;
wire _38998_;
wire _38999_;
wire _39000_;
wire _39001_;
wire _39002_;
wire _39003_;
wire _39004_;
wire _39005_;
wire _39006_;
wire _39007_;
wire _39008_;
wire _39009_;
wire _39010_;
wire _39011_;
wire _39012_;
wire _39013_;
wire _39014_;
wire _39015_;
wire _39016_;
wire _39017_;
wire _39018_;
wire _39019_;
wire _39020_;
wire _39021_;
wire _39022_;
wire _39023_;
wire _39024_;
wire _39025_;
wire _39026_;
wire _39027_;
wire _39028_;
wire _39029_;
wire _39030_;
wire _39031_;
wire _39032_;
wire _39033_;
wire _39034_;
wire _39035_;
wire _39036_;
wire _39037_;
wire _39038_;
wire _39039_;
wire _39040_;
wire _39041_;
wire _39042_;
wire _39043_;
wire _39044_;
wire _39045_;
wire _39046_;
wire _39047_;
wire _39048_;
wire _39049_;
wire _39050_;
wire _39051_;
wire _39052_;
wire _39053_;
wire _39054_;
wire _39055_;
wire _39056_;
wire _39057_;
wire _39058_;
wire _39059_;
wire _39060_;
wire _39061_;
wire _39062_;
wire _39063_;
wire _39064_;
wire _39065_;
wire _39066_;
wire _39067_;
wire _39068_;
wire _39069_;
wire _39070_;
wire _39071_;
wire _39072_;
wire _39073_;
wire _39074_;
wire _39075_;
wire _39076_;
wire _39077_;
wire _39078_;
wire _39079_;
wire _39080_;
wire _39081_;
wire _39082_;
wire _39083_;
wire _39084_;
wire _39085_;
wire _39086_;
wire _39087_;
wire _39088_;
wire _39089_;
wire _39090_;
wire _39091_;
wire _39092_;
wire _39093_;
wire _39094_;
wire _39095_;
wire _39096_;
wire _39097_;
wire _39098_;
wire _39099_;
wire _39100_;
wire _39101_;
wire _39102_;
wire _39103_;
wire _39104_;
wire _39105_;
wire _39106_;
wire _39107_;
wire _39108_;
wire _39109_;
wire _39110_;
wire _39111_;
wire _39112_;
wire _39113_;
wire _39114_;
wire _39115_;
wire _39116_;
wire _39117_;
wire _39118_;
wire _39119_;
wire _39120_;
wire _39121_;
wire _39122_;
wire _39123_;
wire _39124_;
wire _39125_;
wire _39126_;
wire _39127_;
wire _39128_;
wire _39129_;
wire _39130_;
wire _39131_;
wire _39132_;
wire _39133_;
wire _39134_;
wire _39135_;
wire _39136_;
wire _39137_;
wire _39138_;
wire _39139_;
wire _39140_;
wire _39141_;
wire _39142_;
wire _39143_;
wire _39144_;
wire _39145_;
wire _39146_;
wire _39147_;
wire _39148_;
wire _39149_;
wire _39150_;
wire _39151_;
wire _39152_;
wire _39153_;
wire _39154_;
wire _39155_;
wire _39156_;
wire _39157_;
wire _39158_;
wire _39159_;
wire _39160_;
wire _39161_;
wire _39162_;
wire _39163_;
wire _39164_;
wire _39165_;
wire _39166_;
wire _39167_;
wire _39168_;
wire _39169_;
wire _39170_;
wire _39171_;
wire _39172_;
wire _39173_;
wire _39174_;
wire _39175_;
wire _39176_;
wire _39177_;
wire _39178_;
wire _39179_;
wire _39180_;
wire _39181_;
wire _39182_;
wire _39183_;
wire _39184_;
wire _39185_;
wire _39186_;
wire _39187_;
wire _39188_;
wire _39189_;
wire _39190_;
wire _39191_;
wire _39192_;
wire _39193_;
wire _39194_;
wire _39195_;
wire _39196_;
wire _39197_;
wire _39198_;
wire _39199_;
wire _39200_;
wire _39201_;
wire _39202_;
wire _39203_;
wire _39204_;
wire _39205_;
wire _39206_;
wire _39207_;
wire _39208_;
wire _39209_;
wire _39210_;
wire _39211_;
wire _39212_;
wire _39213_;
wire _39214_;
wire _39215_;
wire _39216_;
wire _39217_;
wire _39218_;
wire _39219_;
wire _39220_;
wire _39221_;
wire _39222_;
wire _39223_;
wire _39224_;
wire _39225_;
wire _39226_;
wire _39227_;
wire _39228_;
wire _39229_;
wire _39230_;
wire _39231_;
wire _39232_;
wire _39233_;
wire _39234_;
wire _39235_;
wire _39236_;
wire _39237_;
wire _39238_;
wire _39239_;
wire _39240_;
wire _39241_;
wire _39242_;
wire _39243_;
wire _39244_;
wire _39245_;
wire _39246_;
wire _39247_;
wire _39248_;
wire _39249_;
wire _39250_;
wire _39251_;
wire _39252_;
wire _39253_;
wire _39254_;
wire _39255_;
wire _39256_;
wire _39257_;
wire _39258_;
wire _39259_;
wire _39260_;
wire _39261_;
wire _39262_;
wire _39263_;
wire _39264_;
wire _39265_;
wire _39266_;
wire _39267_;
wire _39268_;
wire _39269_;
wire _39270_;
wire _39271_;
wire _39272_;
wire _39273_;
wire _39274_;
wire _39275_;
wire _39276_;
wire _39277_;
wire _39278_;
wire _39279_;
wire _39280_;
wire _39281_;
wire _39282_;
wire _39283_;
wire _39284_;
wire _39285_;
wire _39286_;
wire _39287_;
wire _39288_;
wire _39289_;
wire _39290_;
wire _39291_;
wire _39292_;
wire _39293_;
wire _39294_;
wire _39295_;
wire _39296_;
wire _39297_;
wire _39298_;
wire _39299_;
wire _39300_;
wire _39301_;
wire _39302_;
wire _39303_;
wire _39304_;
wire _39305_;
wire _39306_;
wire _39307_;
wire _39308_;
wire _39309_;
wire _39310_;
wire _39311_;
wire _39312_;
wire _39313_;
wire _39314_;
wire _39315_;
wire _39316_;
wire _39317_;
wire _39318_;
wire _39319_;
wire _39320_;
wire _39321_;
wire _39322_;
wire _39323_;
wire _39324_;
wire _39325_;
wire _39326_;
wire _39327_;
wire _39328_;
wire _39329_;
wire _39330_;
wire _39331_;
wire _39332_;
wire _39333_;
wire _39334_;
wire _39335_;
wire _39336_;
wire _39337_;
wire _39338_;
wire _39339_;
wire _39340_;
wire _39341_;
wire _39342_;
wire _39343_;
wire _39344_;
wire _39345_;
wire _39346_;
wire _39347_;
wire _39348_;
wire _39349_;
wire _39350_;
wire _39351_;
wire _39352_;
wire _39353_;
wire _39354_;
wire _39355_;
wire _39356_;
wire _39357_;
wire _39358_;
wire _39359_;
wire _39360_;
wire _39361_;
wire _39362_;
wire _39363_;
wire _39364_;
wire _39365_;
wire _39366_;
wire _39367_;
wire _39368_;
wire _39369_;
wire _39370_;
wire _39371_;
wire _39372_;
wire _39373_;
wire _39374_;
wire _39375_;
wire _39376_;
wire _39377_;
wire _39378_;
wire _39379_;
wire _39380_;
wire _39381_;
wire _39382_;
wire _39383_;
wire _39384_;
wire _39385_;
wire _39386_;
wire _39387_;
wire _39388_;
wire _39389_;
wire _39390_;
wire _39391_;
wire _39392_;
wire _39393_;
wire _39394_;
wire _39395_;
wire _39396_;
wire _39397_;
wire _39398_;
wire _39399_;
wire _39400_;
wire _39401_;
wire _39402_;
wire _39403_;
wire _39404_;
wire _39405_;
wire _39406_;
wire _39407_;
wire _39408_;
wire _39409_;
wire _39410_;
wire _39411_;
wire _39412_;
wire _39413_;
wire _39414_;
wire _39415_;
wire _39416_;
wire _39417_;
wire _39418_;
wire _39419_;
wire _39420_;
wire _39421_;
wire _39422_;
wire _39423_;
wire _39424_;
wire _39425_;
wire _39426_;
wire _39427_;
wire _39428_;
wire _39429_;
wire _39430_;
wire _39431_;
wire _39432_;
wire _39433_;
wire _39434_;
wire _39435_;
wire _39436_;
wire _39437_;
wire _39438_;
wire _39439_;
wire _39440_;
wire _39441_;
wire _39442_;
wire _39443_;
wire _39444_;
wire _39445_;
wire _39446_;
wire _39447_;
wire _39448_;
wire _39449_;
wire _39450_;
wire _39451_;
wire _39452_;
wire _39453_;
wire _39454_;
wire _39455_;
wire _39456_;
wire _39457_;
wire _39458_;
wire _39459_;
wire _39460_;
wire _39461_;
wire _39462_;
wire _39463_;
wire _39464_;
wire _39465_;
wire _39466_;
wire _39467_;
wire _39468_;
wire _39469_;
wire _39470_;
wire _39471_;
wire _39472_;
wire _39473_;
wire _39474_;
wire _39475_;
wire _39476_;
wire _39477_;
wire _39478_;
wire _39479_;
wire _39480_;
wire _39481_;
wire _39482_;
wire _39483_;
wire _39484_;
wire _39485_;
wire _39486_;
wire _39487_;
wire _39488_;
wire _39489_;
wire _39490_;
wire _39491_;
wire _39492_;
wire _39493_;
wire _39494_;
wire _39495_;
wire _39496_;
wire _39497_;
wire _39498_;
wire _39499_;
wire _39500_;
wire _39501_;
wire _39502_;
wire _39503_;
wire _39504_;
wire _39505_;
wire _39506_;
wire _39507_;
wire _39508_;
wire _39509_;
wire _39510_;
wire _39511_;
wire _39512_;
wire _39513_;
wire _39514_;
wire _39515_;
wire _39516_;
wire _39517_;
wire _39518_;
wire _39519_;
wire _39520_;
wire _39521_;
wire _39522_;
wire _39523_;
wire _39524_;
wire _39525_;
wire _39526_;
wire _39527_;
wire _39528_;
wire _39529_;
wire _39530_;
wire _39531_;
wire _39532_;
wire _39533_;
wire _39534_;
wire _39535_;
wire _39536_;
wire _39537_;
wire _39538_;
wire _39539_;
wire _39540_;
wire _39541_;
wire _39542_;
wire _39543_;
wire _39544_;
wire _39545_;
wire _39546_;
wire _39547_;
wire _39548_;
wire _39549_;
wire _39550_;
wire _39551_;
wire _39552_;
wire _39553_;
wire _39554_;
wire _39555_;
wire _39556_;
wire _39557_;
wire _39558_;
wire _39559_;
wire _39560_;
wire _39561_;
wire _39562_;
wire _39563_;
wire _39564_;
wire _39565_;
wire _39566_;
wire _39567_;
wire _39568_;
wire _39569_;
wire _39570_;
wire _39571_;
wire _39572_;
wire _39573_;
wire _39574_;
wire _39575_;
wire _39576_;
wire _39577_;
wire _39578_;
wire _39579_;
wire _39580_;
wire _39581_;
wire _39582_;
wire _39583_;
wire _39584_;
wire _39585_;
wire _39586_;
wire _39587_;
wire _39588_;
wire _39589_;
wire _39590_;
wire _39591_;
wire _39592_;
wire _39593_;
wire _39594_;
wire _39595_;
wire _39596_;
wire _39597_;
wire _39598_;
wire _39599_;
wire _39600_;
wire _39601_;
wire _39602_;
wire _39603_;
wire _39604_;
wire _39605_;
wire _39606_;
wire _39607_;
wire _39608_;
wire _39609_;
wire _39610_;
wire _39611_;
wire _39612_;
wire _39613_;
wire _39614_;
wire _39615_;
wire _39616_;
wire _39617_;
wire _39618_;
wire _39619_;
wire _39620_;
wire _39621_;
wire _39622_;
wire _39623_;
wire _39624_;
wire _39625_;
wire _39626_;
wire _39627_;
wire _39628_;
wire _39629_;
wire _39630_;
wire _39631_;
wire _39632_;
wire _39633_;
wire _39634_;
wire _39635_;
wire _39636_;
wire _39637_;
wire _39638_;
wire _39639_;
wire _39640_;
wire _39641_;
wire _39642_;
wire _39643_;
wire _39644_;
wire _39645_;
wire _39646_;
wire _39647_;
wire _39648_;
wire _39649_;
wire _39650_;
wire _39651_;
wire _39652_;
wire _39653_;
wire _39654_;
wire _39655_;
wire _39656_;
wire _39657_;
wire _39658_;
wire _39659_;
wire _39660_;
wire _39661_;
wire _39662_;
wire _39663_;
wire _39664_;
wire _39665_;
wire _39666_;
wire _39667_;
wire _39668_;
wire _39669_;
wire _39670_;
wire _39671_;
wire _39672_;
wire _39673_;
wire _39674_;
wire _39675_;
wire _39676_;
wire _39677_;
wire _39678_;
wire _39679_;
wire _39680_;
wire _39681_;
wire _39682_;
wire _39683_;
wire _39684_;
wire _39685_;
wire _39686_;
wire _39687_;
wire _39688_;
wire _39689_;
wire _39690_;
wire _39691_;
wire _39692_;
wire _39693_;
wire _39694_;
wire _39695_;
wire _39696_;
wire _39697_;
wire _39698_;
wire _39699_;
wire _39700_;
wire _39701_;
wire _39702_;
wire _39703_;
wire _39704_;
wire _39705_;
wire _39706_;
wire _39707_;
wire _39708_;
wire _39709_;
wire _39710_;
wire _39711_;
wire _39712_;
wire _39713_;
wire _39714_;
wire _39715_;
wire _39716_;
wire _39717_;
wire _39718_;
wire _39719_;
wire _39720_;
wire _39721_;
wire _39722_;
wire _39723_;
wire _39724_;
wire _39725_;
wire _39726_;
wire _39727_;
wire _39728_;
wire _39729_;
wire _39730_;
wire _39731_;
wire _39732_;
wire _39733_;
wire _39734_;
wire _39735_;
wire _39736_;
wire _39737_;
wire _39738_;
wire _39739_;
wire _39740_;
wire _39741_;
wire _39742_;
wire _39743_;
wire _39744_;
wire _39745_;
wire _39746_;
wire _39747_;
wire _39748_;
wire _39749_;
wire _39750_;
wire _39751_;
wire _39752_;
wire _39753_;
wire _39754_;
wire _39755_;
wire _39756_;
wire _39757_;
wire _39758_;
wire _39759_;
wire _39760_;
wire _39761_;
wire _39762_;
wire _39763_;
wire _39764_;
wire _39765_;
wire _39766_;
wire _39767_;
wire _39768_;
wire _39769_;
wire _39770_;
wire _39771_;
wire _39772_;
wire _39773_;
wire _39774_;
wire _39775_;
wire _39776_;
wire _39777_;
wire _39778_;
wire _39779_;
wire _39780_;
wire _39781_;
wire _39782_;
wire _39783_;
wire _39784_;
wire _39785_;
wire _39786_;
wire _39787_;
wire _39788_;
wire _39789_;
wire _39790_;
wire _39791_;
wire _39792_;
wire _39793_;
wire _39794_;
wire _39795_;
wire _39796_;
wire _39797_;
wire _39798_;
wire _39799_;
wire _39800_;
wire _39801_;
wire _39802_;
wire _39803_;
wire _39804_;
wire _39805_;
wire _39806_;
wire _39807_;
wire _39808_;
wire _39809_;
wire _39810_;
wire _39811_;
wire _39812_;
wire _39813_;
wire _39814_;
wire _39815_;
wire _39816_;
wire _39817_;
wire _39818_;
wire _39819_;
wire _39820_;
wire _39821_;
wire _39822_;
wire _39823_;
wire _39824_;
wire _39825_;
wire _39826_;
wire _39827_;
wire _39828_;
wire _39829_;
wire _39830_;
wire _39831_;
wire _39832_;
wire _39833_;
wire _39834_;
wire _39835_;
wire _39836_;
wire _39837_;
wire _39838_;
wire _39839_;
wire _39840_;
wire _39841_;
wire _39842_;
wire _39843_;
wire _39844_;
wire _39845_;
wire _39846_;
wire _39847_;
wire _39848_;
wire _39849_;
wire _39850_;
wire _39851_;
wire _39852_;
wire _39853_;
wire _39854_;
wire _39855_;
wire _39856_;
wire _39857_;
wire _39858_;
wire _39859_;
wire _39860_;
wire _39861_;
wire _39862_;
wire _39863_;
wire _39864_;
wire _39865_;
wire _39866_;
wire _39867_;
wire _39868_;
wire _39869_;
wire _39870_;
wire _39871_;
wire _39872_;
wire _39873_;
wire _39874_;
wire _39875_;
wire _39876_;
wire _39877_;
wire _39878_;
wire _39879_;
wire _39880_;
wire _39881_;
wire _39882_;
wire _39883_;
wire _39884_;
wire _39885_;
wire _39886_;
wire _39887_;
wire _39888_;
wire _39889_;
wire _39890_;
wire _39891_;
wire _39892_;
wire _39893_;
wire _39894_;
wire _39895_;
wire _39896_;
wire _39897_;
wire _39898_;
wire _39899_;
wire _39900_;
wire _39901_;
wire _39902_;
wire _39903_;
wire _39904_;
wire _39905_;
wire _39906_;
wire _39907_;
wire _39908_;
wire _39909_;
wire _39910_;
wire _39911_;
wire _39912_;
wire _39913_;
wire _39914_;
wire _39915_;
wire _39916_;
wire _39917_;
wire _39918_;
wire _39919_;
wire _39920_;
wire _39921_;
wire _39922_;
wire _39923_;
wire _39924_;
wire _39925_;
wire _39926_;
wire _39927_;
wire _39928_;
wire _39929_;
wire _39930_;
wire _39931_;
wire _39932_;
wire _39933_;
wire _39934_;
wire _39935_;
wire _39936_;
wire _39937_;
wire _39938_;
wire _39939_;
wire _39940_;
wire _39941_;
wire _39942_;
wire _39943_;
wire _39944_;
wire _39945_;
wire _39946_;
wire _39947_;
wire _39948_;
wire _39949_;
wire _39950_;
wire _39951_;
wire _39952_;
wire _39953_;
wire _39954_;
wire _39955_;
wire _39956_;
wire _39957_;
wire _39958_;
wire _39959_;
wire _39960_;
wire _39961_;
wire _39962_;
wire _39963_;
wire _39964_;
wire _39965_;
wire _39966_;
wire _39967_;
wire _39968_;
wire _39969_;
wire _39970_;
wire _39971_;
wire _39972_;
wire _39973_;
wire _39974_;
wire _39975_;
wire _39976_;
wire _39977_;
wire _39978_;
wire _39979_;
wire _39980_;
wire _39981_;
wire _39982_;
wire _39983_;
wire _39984_;
wire _39985_;
wire _39986_;
wire _39987_;
wire _39988_;
wire _39989_;
wire _39990_;
wire _39991_;
wire _39992_;
wire _39993_;
wire _39994_;
wire _39995_;
wire _39996_;
wire _39997_;
wire _39998_;
wire _39999_;
wire _40000_;
wire _40001_;
wire _40002_;
wire _40003_;
wire _40004_;
wire _40005_;
wire _40006_;
wire _40007_;
wire _40008_;
wire _40009_;
wire _40010_;
wire _40011_;
wire _40012_;
wire _40013_;
wire _40014_;
wire _40015_;
wire _40016_;
wire _40017_;
wire _40018_;
wire _40019_;
wire _40020_;
wire _40021_;
wire _40022_;
wire _40023_;
wire _40024_;
wire _40025_;
wire _40026_;
wire _40027_;
wire _40028_;
wire _40029_;
wire _40030_;
wire _40031_;
wire _40032_;
wire _40033_;
wire _40034_;
wire _40035_;
wire _40036_;
wire _40037_;
wire _40038_;
wire _40039_;
wire _40040_;
wire _40041_;
wire _40042_;
wire _40043_;
wire _40044_;
wire _40045_;
wire _40046_;
wire _40047_;
wire _40048_;
wire _40049_;
wire _40050_;
wire _40051_;
wire _40052_;
wire _40053_;
wire _40054_;
wire _40055_;
wire _40056_;
wire _40057_;
wire _40058_;
wire _40059_;
wire _40060_;
wire _40061_;
wire _40062_;
wire _40063_;
wire _40064_;
wire _40065_;
wire _40066_;
wire _40067_;
wire _40068_;
wire _40069_;
wire _40070_;
wire _40071_;
wire _40072_;
wire _40073_;
wire _40074_;
wire _40075_;
wire _40076_;
wire _40077_;
wire _40078_;
wire _40079_;
wire _40080_;
wire _40081_;
wire _40082_;
wire _40083_;
wire _40084_;
wire _40085_;
wire _40086_;
wire _40087_;
wire _40088_;
wire _40089_;
wire _40090_;
wire _40091_;
wire _40092_;
wire _40093_;
wire _40094_;
wire _40095_;
wire _40096_;
wire _40097_;
wire _40098_;
wire _40099_;
wire _40100_;
wire _40101_;
wire _40102_;
wire _40103_;
wire _40104_;
wire _40105_;
wire _40106_;
wire _40107_;
wire _40108_;
wire _40109_;
wire _40110_;
wire _40111_;
wire _40112_;
wire _40113_;
wire _40114_;
wire _40115_;
wire _40116_;
wire _40117_;
wire _40118_;
wire _40119_;
wire _40120_;
wire _40121_;
wire _40122_;
wire _40123_;
wire _40124_;
wire _40125_;
wire _40126_;
wire _40127_;
wire _40128_;
wire _40129_;
wire _40130_;
wire _40131_;
wire _40132_;
wire _40133_;
wire _40134_;
wire _40135_;
wire _40136_;
wire _40137_;
wire _40138_;
wire _40139_;
wire _40140_;
wire _40141_;
wire _40142_;
wire _40143_;
wire _40144_;
wire _40145_;
wire _40146_;
wire _40147_;
wire _40148_;
wire _40149_;
wire _40150_;
wire _40151_;
wire _40152_;
wire _40153_;
wire _40154_;
wire _40155_;
wire _40156_;
wire _40157_;
wire _40158_;
wire _40159_;
wire _40160_;
wire _40161_;
wire _40162_;
wire _40163_;
wire _40164_;
wire _40165_;
wire _40166_;
wire _40167_;
wire _40168_;
wire _40169_;
wire _40170_;
wire _40171_;
wire _40172_;
wire _40173_;
wire _40174_;
wire _40175_;
wire _40176_;
wire _40177_;
wire _40178_;
wire _40179_;
wire _40180_;
wire _40181_;
wire _40182_;
wire _40183_;
wire _40184_;
wire _40185_;
wire _40186_;
wire _40187_;
wire _40188_;
wire _40189_;
wire _40190_;
wire _40191_;
wire _40192_;
wire _40193_;
wire _40194_;
wire _40195_;
wire _40196_;
wire _40197_;
wire _40198_;
wire _40199_;
wire _40200_;
wire _40201_;
wire _40202_;
wire _40203_;
wire _40204_;
wire _40205_;
wire _40206_;
wire _40207_;
wire _40208_;
wire _40209_;
wire _40210_;
wire _40211_;
wire _40212_;
wire _40213_;
wire _40214_;
wire _40215_;
wire _40216_;
wire _40217_;
wire _40218_;
wire _40219_;
wire _40220_;
wire _40221_;
wire _40222_;
wire _40223_;
wire _40224_;
wire _40225_;
wire _40226_;
wire _40227_;
wire _40228_;
wire _40229_;
wire _40230_;
wire _40231_;
wire _40232_;
wire _40233_;
wire _40234_;
wire _40235_;
wire _40236_;
wire _40237_;
wire _40238_;
wire _40239_;
wire _40240_;
wire _40241_;
wire _40242_;
wire _40243_;
wire _40244_;
wire _40245_;
wire _40246_;
wire _40247_;
wire _40248_;
wire _40249_;
wire _40250_;
wire _40251_;
wire _40252_;
wire _40253_;
wire _40254_;
wire _40255_;
wire _40256_;
wire _40257_;
wire _40258_;
wire _40259_;
wire _40260_;
wire _40261_;
wire _40262_;
wire _40263_;
wire _40264_;
wire _40265_;
wire _40266_;
wire _40267_;
wire _40268_;
wire _40269_;
wire _40270_;
wire _40271_;
wire _40272_;
wire _40273_;
wire _40274_;
wire _40275_;
wire _40276_;
wire _40277_;
wire _40278_;
wire _40279_;
wire _40280_;
wire _40281_;
wire _40282_;
wire _40283_;
wire _40284_;
wire _40285_;
wire _40286_;
wire _40287_;
wire _40288_;
wire _40289_;
wire _40290_;
wire _40291_;
wire _40292_;
wire _40293_;
wire _40294_;
wire _40295_;
wire _40296_;
wire _40297_;
wire _40298_;
wire _40299_;
wire _40300_;
wire _40301_;
wire _40302_;
wire _40303_;
wire _40304_;
wire _40305_;
wire _40306_;
wire _40307_;
wire _40308_;
wire _40309_;
wire _40310_;
wire _40311_;
wire _40312_;
wire _40313_;
wire _40314_;
wire _40315_;
wire _40316_;
wire _40317_;
wire _40318_;
wire _40319_;
wire _40320_;
wire _40321_;
wire _40322_;
wire _40323_;
wire _40324_;
wire _40325_;
wire _40326_;
wire _40327_;
wire _40328_;
wire _40329_;
wire _40330_;
wire _40331_;
wire _40332_;
wire _40333_;
wire _40334_;
wire _40335_;
wire _40336_;
wire _40337_;
wire _40338_;
wire _40339_;
wire _40340_;
wire _40341_;
wire _40342_;
wire _40343_;
wire _40344_;
wire _40345_;
wire _40346_;
wire _40347_;
wire _40348_;
wire _40349_;
wire _40350_;
wire _40351_;
wire _40352_;
wire _40353_;
wire _40354_;
wire _40355_;
wire _40356_;
wire _40357_;
wire _40358_;
wire _40359_;
wire _40360_;
wire _40361_;
wire _40362_;
wire _40363_;
wire _40364_;
wire _40365_;
wire _40366_;
wire _40367_;
wire _40368_;
wire _40369_;
wire _40370_;
wire _40371_;
wire _40372_;
wire _40373_;
wire _40374_;
wire _40375_;
wire _40376_;
wire _40377_;
wire _40378_;
wire _40379_;
wire _40380_;
wire _40381_;
wire _40382_;
wire _40383_;
wire _40384_;
wire _40385_;
wire _40386_;
wire _40387_;
wire _40388_;
wire _40389_;
wire _40390_;
wire _40391_;
wire _40392_;
wire _40393_;
wire _40394_;
wire _40395_;
wire _40396_;
wire _40397_;
wire _40398_;
wire _40399_;
wire _40400_;
wire _40401_;
wire _40402_;
wire _40403_;
wire _40404_;
wire _40405_;
wire _40406_;
wire _40407_;
wire _40408_;
wire _40409_;
wire _40410_;
wire _40411_;
wire _40412_;
wire _40413_;
wire _40414_;
wire _40415_;
wire _40416_;
wire _40417_;
wire _40418_;
wire _40419_;
wire _40420_;
wire _40421_;
wire _40422_;
wire _40423_;
wire _40424_;
wire _40425_;
wire _40426_;
wire _40427_;
wire _40428_;
wire _40429_;
wire _40430_;
wire _40431_;
wire _40432_;
wire _40433_;
wire _40434_;
wire _40435_;
wire _40436_;
wire _40437_;
wire _40438_;
wire _40439_;
wire _40440_;
wire _40441_;
wire _40442_;
wire _40443_;
wire _40444_;
wire _40445_;
wire _40446_;
wire _40447_;
wire _40448_;
wire _40449_;
wire _40450_;
wire _40451_;
wire _40452_;
wire _40453_;
wire _40454_;
wire _40455_;
wire _40456_;
wire _40457_;
wire _40458_;
wire _40459_;
wire _40460_;
wire _40461_;
wire _40462_;
wire _40463_;
wire _40464_;
wire _40465_;
wire _40466_;
wire _40467_;
wire _40468_;
wire _40469_;
wire _40470_;
wire _40471_;
wire _40472_;
wire _40473_;
wire _40474_;
wire _40475_;
wire _40476_;
wire _40477_;
wire _40478_;
wire _40479_;
wire _40480_;
wire _40481_;
wire _40482_;
wire _40483_;
wire _40484_;
wire _40485_;
wire _40486_;
wire _40487_;
wire _40488_;
wire _40489_;
wire _40490_;
wire _40491_;
wire _40492_;
wire _40493_;
wire _40494_;
wire _40495_;
wire _40496_;
wire _40497_;
wire _40498_;
wire _40499_;
wire _40500_;
wire _40501_;
wire _40502_;
wire _40503_;
wire _40504_;
wire _40505_;
wire _40506_;
wire _40507_;
wire _40508_;
wire _40509_;
wire _40510_;
wire _40511_;
wire _40512_;
wire _40513_;
wire _40514_;
wire _40515_;
wire _40516_;
wire _40517_;
wire _40518_;
wire _40519_;
wire _40520_;
wire _40521_;
wire _40522_;
wire _40523_;
wire _40524_;
wire _40525_;
wire _40526_;
wire _40527_;
wire _40528_;
wire _40529_;
wire _40530_;
wire _40531_;
wire _40532_;
wire _40533_;
wire _40534_;
wire _40535_;
wire _40536_;
wire _40537_;
wire _40538_;
wire _40539_;
wire _40540_;
wire _40541_;
wire _40542_;
wire _40543_;
wire _40544_;
wire _40545_;
wire _40546_;
wire _40547_;
wire _40548_;
wire _40549_;
wire _40550_;
wire _40551_;
wire _40552_;
wire _40553_;
wire _40554_;
wire _40555_;
wire _40556_;
wire _40557_;
wire _40558_;
wire _40559_;
wire _40560_;
wire _40561_;
wire _40562_;
wire _40563_;
wire _40564_;
wire _40565_;
wire _40566_;
wire _40567_;
wire _40568_;
wire _40569_;
wire _40570_;
wire _40571_;
wire _40572_;
wire _40573_;
wire _40574_;
wire _40575_;
wire _40576_;
wire _40577_;
wire _40578_;
wire _40579_;
wire _40580_;
wire _40581_;
wire _40582_;
wire _40583_;
wire _40584_;
wire _40585_;
wire _40586_;
wire _40587_;
wire _40588_;
wire _40589_;
wire _40590_;
wire _40591_;
wire _40592_;
wire _40593_;
wire _40594_;
wire _40595_;
wire _40596_;
wire _40597_;
wire _40598_;
wire _40599_;
wire _40600_;
wire _40601_;
wire _40602_;
wire _40603_;
wire _40604_;
wire _40605_;
wire _40606_;
wire _40607_;
wire _40608_;
wire _40609_;
wire _40610_;
wire _40611_;
wire _40612_;
wire _40613_;
wire _40614_;
wire _40615_;
wire _40616_;
wire _40617_;
wire _40618_;
wire _40619_;
wire _40620_;
wire _40621_;
wire _40622_;
wire _40623_;
wire _40624_;
wire _40625_;
wire _40626_;
wire _40627_;
wire _40628_;
wire _40629_;
wire _40630_;
wire _40631_;
wire _40632_;
wire _40633_;
wire _40634_;
wire _40635_;
wire _40636_;
wire _40637_;
wire _40638_;
wire _40639_;
wire _40640_;
wire _40641_;
wire _40642_;
wire _40643_;
wire _40644_;
wire _40645_;
wire _40646_;
wire _40647_;
wire _40648_;
wire _40649_;
wire _40650_;
wire _40651_;
wire _40652_;
wire _40653_;
wire _40654_;
wire _40655_;
wire _40656_;
wire _40657_;
wire _40658_;
wire _40659_;
wire _40660_;
wire _40661_;
wire _40662_;
wire _40663_;
wire _40664_;
wire _40665_;
wire _40666_;
wire _40667_;
wire _40668_;
wire _40669_;
wire _40670_;
wire _40671_;
wire _40672_;
wire _40673_;
wire _40674_;
wire _40675_;
wire _40676_;
wire _40677_;
wire _40678_;
wire _40679_;
wire _40680_;
wire _40681_;
wire _40682_;
wire _40683_;
wire _40684_;
wire _40685_;
wire _40686_;
wire _40687_;
wire _40688_;
wire _40689_;
wire _40690_;
wire _40691_;
wire _40692_;
wire _40693_;
wire _40694_;
wire _40695_;
wire _40696_;
wire _40697_;
wire _40698_;
wire _40699_;
wire _40700_;
wire _40701_;
wire _40702_;
wire _40703_;
wire _40704_;
wire _40705_;
wire _40706_;
wire _40707_;
wire _40708_;
wire _40709_;
wire _40710_;
wire _40711_;
wire _40712_;
wire _40713_;
wire _40714_;
wire _40715_;
wire _40716_;
wire _40717_;
wire _40718_;
wire _40719_;
wire _40720_;
wire _40721_;
wire _40722_;
wire _40723_;
wire _40724_;
wire _40725_;
wire _40726_;
wire _40727_;
wire _40728_;
wire _40729_;
wire _40730_;
wire _40731_;
wire _40732_;
wire _40733_;
wire _40734_;
wire _40735_;
wire _40736_;
wire _40737_;
wire _40738_;
wire _40739_;
wire _40740_;
wire _40741_;
wire _40742_;
wire _40743_;
wire _40744_;
wire _40745_;
wire _40746_;
wire _40747_;
wire _40748_;
wire _40749_;
wire _40750_;
wire _40751_;
wire _40752_;
wire _40753_;
wire _40754_;
wire _40755_;
wire _40756_;
wire _40757_;
wire _40758_;
wire _40759_;
wire _40760_;
wire _40761_;
wire _40762_;
wire _40763_;
wire _40764_;
wire _40765_;
wire _40766_;
wire _40767_;
wire _40768_;
wire _40769_;
wire _40770_;
wire _40771_;
wire _40772_;
wire _40773_;
wire _40774_;
wire _40775_;
wire _40776_;
wire _40777_;
wire _40778_;
wire _40779_;
wire _40780_;
wire _40781_;
wire _40782_;
wire _40783_;
wire _40784_;
wire _40785_;
wire _40786_;
wire _40787_;
wire _40788_;
wire _40789_;
wire _40790_;
wire _40791_;
wire _40792_;
wire _40793_;
wire _40794_;
wire _40795_;
wire _40796_;
wire _40797_;
wire _40798_;
wire _40799_;
wire _40800_;
wire _40801_;
wire _40802_;
wire _40803_;
wire _40804_;
wire _40805_;
wire _40806_;
wire _40807_;
wire _40808_;
wire _40809_;
wire _40810_;
wire _40811_;
wire _40812_;
wire _40813_;
wire _40814_;
wire _40815_;
wire _40816_;
wire _40817_;
wire _40818_;
wire _40819_;
wire _40820_;
wire _40821_;
wire _40822_;
wire _40823_;
wire _40824_;
wire _40825_;
wire _40826_;
wire _40827_;
wire _40828_;
wire _40829_;
wire _40830_;
wire _40831_;
wire _40832_;
wire _40833_;
wire _40834_;
wire _40835_;
wire _40836_;
wire _40837_;
wire _40838_;
wire _40839_;
wire _40840_;
wire _40841_;
wire _40842_;
wire _40843_;
wire _40844_;
wire _40845_;
wire _40846_;
wire _40847_;
wire _40848_;
wire _40849_;
wire _40850_;
wire _40851_;
wire _40852_;
wire _40853_;
wire _40854_;
wire _40855_;
wire _40856_;
wire _40857_;
wire _40858_;
wire _40859_;
wire _40860_;
wire _40861_;
wire _40862_;
wire _40863_;
wire _40864_;
wire _40865_;
wire _40866_;
wire _40867_;
wire _40868_;
wire _40869_;
wire _40870_;
wire _40871_;
wire _40872_;
wire _40873_;
wire _40874_;
wire _40875_;
wire _40876_;
wire _40877_;
wire _40878_;
wire _40879_;
wire _40880_;
wire _40881_;
wire _40882_;
wire _40883_;
wire _40884_;
wire _40885_;
wire _40886_;
wire _40887_;
wire _40888_;
wire _40889_;
wire _40890_;
wire _40891_;
wire _40892_;
wire _40893_;
wire _40894_;
wire _40895_;
wire _40896_;
wire _40897_;
wire _40898_;
wire _40899_;
wire _40900_;
wire _40901_;
wire _40902_;
wire _40903_;
wire _40904_;
wire _40905_;
wire _40906_;
wire _40907_;
wire _40908_;
wire _40909_;
wire _40910_;
wire _40911_;
wire _40912_;
wire _40913_;
wire _40914_;
wire _40915_;
wire _40916_;
wire _40917_;
wire _40918_;
wire _40919_;
wire _40920_;
wire _40921_;
wire _40922_;
wire _40923_;
wire _40924_;
wire _40925_;
wire _40926_;
wire _40927_;
wire _40928_;
wire _40929_;
wire _40930_;
wire _40931_;
wire _40932_;
wire _40933_;
wire _40934_;
wire _40935_;
wire _40936_;
wire _40937_;
wire _40938_;
wire _40939_;
wire _40940_;
wire _40941_;
wire _40942_;
wire _40943_;
wire _40944_;
wire _40945_;
wire _40946_;
wire _40947_;
wire _40948_;
wire _40949_;
wire _40950_;
wire _40951_;
wire _40952_;
wire _40953_;
wire _40954_;
wire _40955_;
wire _40956_;
wire _40957_;
wire _40958_;
wire _40959_;
wire _40960_;
wire _40961_;
wire _40962_;
wire _40963_;
wire _40964_;
wire _40965_;
wire _40966_;
wire _40967_;
wire _40968_;
wire _40969_;
wire _40970_;
wire _40971_;
wire _40972_;
wire _40973_;
wire _40974_;
wire _40975_;
wire _40976_;
wire _40977_;
wire _40978_;
wire _40979_;
wire _40980_;
wire _40981_;
wire _40982_;
wire _40983_;
wire _40984_;
wire _40985_;
wire _40986_;
wire _40987_;
wire _40988_;
wire _40989_;
wire _40990_;
wire _40991_;
wire _40992_;
wire _40993_;
wire _40994_;
wire _40995_;
wire _40996_;
wire _40997_;
wire _40998_;
wire _40999_;
wire _41000_;
wire _41001_;
wire _41002_;
wire _41003_;
wire _41004_;
wire _41005_;
wire _41006_;
wire _41007_;
wire _41008_;
wire _41009_;
wire _41010_;
wire _41011_;
wire _41012_;
wire _41013_;
wire _41014_;
wire _41015_;
wire _41016_;
wire _41017_;
wire _41018_;
wire _41019_;
wire _41020_;
wire _41021_;
wire _41022_;
wire _41023_;
wire _41024_;
wire _41025_;
wire _41026_;
wire _41027_;
wire _41028_;
wire _41029_;
wire _41030_;
wire _41031_;
wire _41032_;
wire _41033_;
wire _41034_;
wire _41035_;
wire _41036_;
wire _41037_;
wire _41038_;
wire _41039_;
wire _41040_;
wire _41041_;
wire _41042_;
wire _41043_;
wire _41044_;
wire _41045_;
wire _41046_;
wire _41047_;
wire _41048_;
wire _41049_;
wire _41050_;
wire _41051_;
wire _41052_;
wire _41053_;
wire _41054_;
wire _41055_;
wire _41056_;
wire _41057_;
wire _41058_;
wire _41059_;
wire _41060_;
wire _41061_;
wire _41062_;
wire _41063_;
wire _41064_;
wire _41065_;
wire _41066_;
wire _41067_;
wire _41068_;
wire _41069_;
wire _41070_;
wire _41071_;
wire _41072_;
wire _41073_;
wire _41074_;
wire _41075_;
wire _41076_;
wire _41077_;
wire _41078_;
wire _41079_;
wire _41080_;
wire _41081_;
wire _41082_;
wire _41083_;
wire _41084_;
wire _41085_;
wire _41086_;
wire _41087_;
wire _41088_;
wire _41089_;
wire _41090_;
wire _41091_;
wire _41092_;
wire _41093_;
wire _41094_;
wire _41095_;
wire _41096_;
wire _41097_;
wire _41098_;
wire _41099_;
wire _41100_;
wire _41101_;
wire _41102_;
wire _41103_;
wire _41104_;
wire _41105_;
wire _41106_;
wire _41107_;
wire _41108_;
wire _41109_;
wire _41110_;
wire _41111_;
wire _41112_;
wire _41113_;
wire _41114_;
wire _41115_;
wire _41116_;
wire _41117_;
wire _41118_;
wire _41119_;
wire _41120_;
wire _41121_;
wire _41122_;
wire _41123_;
wire _41124_;
wire _41125_;
wire _41126_;
wire _41127_;
wire _41128_;
wire _41129_;
wire _41130_;
wire _41131_;
wire _41132_;
wire _41133_;
wire _41134_;
wire _41135_;
wire _41136_;
wire _41137_;
wire _41138_;
wire _41139_;
wire _41140_;
wire _41141_;
wire _41142_;
wire _41143_;
wire _41144_;
wire _41145_;
wire _41146_;
wire _41147_;
wire _41148_;
wire _41149_;
wire _41150_;
wire _41151_;
wire _41152_;
wire _41153_;
wire _41154_;
wire _41155_;
wire _41156_;
wire _41157_;
wire _41158_;
wire _41159_;
wire _41160_;
wire _41161_;
wire _41162_;
wire _41163_;
wire _41164_;
wire _41165_;
wire _41166_;
wire _41167_;
wire _41168_;
wire _41169_;
wire _41170_;
wire _41171_;
wire _41172_;
wire _41173_;
wire _41174_;
wire _41175_;
wire _41176_;
wire _41177_;
wire _41178_;
wire _41179_;
wire _41180_;
wire _41181_;
wire _41182_;
wire _41183_;
wire _41184_;
wire _41185_;
wire _41186_;
wire _41187_;
wire _41188_;
wire _41189_;
wire _41190_;
wire _41191_;
wire _41192_;
wire _41193_;
wire _41194_;
wire _41195_;
wire _41196_;
wire _41197_;
wire _41198_;
wire _41199_;
wire _41200_;
wire _41201_;
wire _41202_;
wire _41203_;
wire _41204_;
wire _41205_;
wire _41206_;
wire _41207_;
wire _41208_;
wire _41209_;
wire _41210_;
wire _41211_;
wire _41212_;
wire _41213_;
wire _41214_;
wire _41215_;
wire _41216_;
wire _41217_;
wire _41218_;
wire _41219_;
wire _41220_;
wire _41221_;
wire _41222_;
wire _41223_;
wire _41224_;
wire _41225_;
wire _41226_;
wire _41227_;
wire _41228_;
wire _41229_;
wire _41230_;
wire _41231_;
wire _41232_;
wire _41233_;
wire _41234_;
wire _41235_;
wire _41236_;
wire _41237_;
wire _41238_;
wire _41239_;
wire _41240_;
wire _41241_;
wire _41242_;
wire _41243_;
wire _41244_;
wire _41245_;
wire _41246_;
wire _41247_;
wire _41248_;
wire _41249_;
wire _41250_;
wire _41251_;
wire _41252_;
wire _41253_;
wire _41254_;
wire _41255_;
wire _41256_;
wire _41257_;
wire _41258_;
wire _41259_;
wire _41260_;
wire _41261_;
wire _41262_;
wire _41263_;
wire _41264_;
wire _41265_;
wire _41266_;
wire _41267_;
wire _41268_;
wire _41269_;
wire _41270_;
wire _41271_;
wire _41272_;
wire _41273_;
wire _41274_;
wire _41275_;
wire _41276_;
wire _41277_;
wire _41278_;
wire _41279_;
wire _41280_;
wire _41281_;
wire _41282_;
wire _41283_;
wire _41284_;
wire _41285_;
wire _41286_;
wire _41287_;
wire _41288_;
wire _41289_;
wire _41290_;
wire _41291_;
wire _41292_;
wire _41293_;
wire _41294_;
wire _41295_;
wire _41296_;
wire _41297_;
wire _41298_;
wire _41299_;
wire _41300_;
wire _41301_;
wire _41302_;
wire _41303_;
wire _41304_;
wire _41305_;
wire _41306_;
wire _41307_;
wire _41308_;
wire _41309_;
wire _41310_;
wire _41311_;
wire _41312_;
wire _41313_;
wire _41314_;
wire _41315_;
wire _41316_;
wire _41317_;
wire _41318_;
wire _41319_;
wire _41320_;
wire _41321_;
wire _41322_;
wire _41323_;
wire _41324_;
wire _41325_;
wire _41326_;
wire _41327_;
wire _41328_;
wire _41329_;
wire _41330_;
wire _41331_;
wire _41332_;
wire _41333_;
wire _41334_;
wire _41335_;
wire _41336_;
wire _41337_;
wire _41338_;
wire _41339_;
wire _41340_;
wire _41341_;
wire _41342_;
wire _41343_;
wire _41344_;
wire _41345_;
wire _41346_;
wire _41347_;
wire _41348_;
wire _41349_;
wire _41350_;
wire _41351_;
wire _41352_;
wire _41353_;
wire _41354_;
wire _41355_;
wire _41356_;
wire _41357_;
wire _41358_;
wire _41359_;
wire _41360_;
wire _41361_;
wire _41362_;
wire _41363_;
wire _41364_;
wire _41365_;
wire _41366_;
wire _41367_;
wire _41368_;
wire _41369_;
wire _41370_;
wire _41371_;
wire _41372_;
wire _41373_;
wire _41374_;
wire _41375_;
wire _41376_;
wire _41377_;
wire _41378_;
wire _41379_;
wire _41380_;
wire _41381_;
wire _41382_;
wire _41383_;
wire _41384_;
wire _41385_;
wire _41386_;
wire _41387_;
wire _41388_;
wire _41389_;
wire _41390_;
wire _41391_;
wire _41392_;
wire _41393_;
wire _41394_;
wire _41395_;
wire _41396_;
wire _41397_;
wire _41398_;
wire _41399_;
wire _41400_;
wire _41401_;
wire _41402_;
wire _41403_;
wire _41404_;
wire _41405_;
wire _41406_;
wire _41407_;
wire _41408_;
wire _41409_;
wire _41410_;
wire _41411_;
wire _41412_;
wire _41413_;
wire _41414_;
wire _41415_;
wire _41416_;
wire _41417_;
wire _41418_;
wire _41419_;
wire _41420_;
wire _41421_;
wire _41422_;
wire _41423_;
wire _41424_;
wire _41425_;
wire _41426_;
wire _41427_;
wire _41428_;
wire _41429_;
wire _41430_;
wire _41431_;
wire _41432_;
wire _41433_;
wire _41434_;
wire _41435_;
wire _41436_;
wire _41437_;
wire _41438_;
wire _41439_;
wire _41440_;
wire _41441_;
wire _41442_;
wire _41443_;
wire _41444_;
wire _41445_;
wire _41446_;
wire _41447_;
wire _41448_;
wire _41449_;
wire _41450_;
wire _41451_;
wire _41452_;
wire _41453_;
wire _41454_;
wire _41455_;
wire _41456_;
wire _41457_;
wire _41458_;
wire _41459_;
wire _41460_;
wire _41461_;
wire _41462_;
wire _41463_;
wire _41464_;
wire _41465_;
wire _41466_;
wire _41467_;
wire _41468_;
wire _41469_;
wire _41470_;
wire _41471_;
wire _41472_;
wire _41473_;
wire _41474_;
wire _41475_;
wire _41476_;
wire _41477_;
wire _41478_;
wire _41479_;
wire _41480_;
wire _41481_;
wire _41482_;
wire _41483_;
wire _41484_;
wire _41485_;
wire _41486_;
wire _41487_;
wire _41488_;
wire _41489_;
wire _41490_;
wire _41491_;
wire _41492_;
wire _41493_;
wire _41494_;
wire _41495_;
wire _41496_;
wire _41497_;
wire _41498_;
wire _41499_;
wire _41500_;
wire _41501_;
wire _41502_;
wire _41503_;
wire _41504_;
wire _41505_;
wire _41506_;
wire _41507_;
wire _41508_;
wire _41509_;
wire _41510_;
wire _41511_;
wire _41512_;
wire _41513_;
wire _41514_;
wire _41515_;
wire _41516_;
wire _41517_;
wire _41518_;
wire _41519_;
wire _41520_;
wire _41521_;
wire _41522_;
wire _41523_;
wire _41524_;
wire _41525_;
wire _41526_;
wire _41527_;
wire _41528_;
wire _41529_;
wire _41530_;
wire _41531_;
wire _41532_;
wire _41533_;
wire _41534_;
wire _41535_;
wire _41536_;
wire _41537_;
wire _41538_;
wire _41539_;
wire _41540_;
wire _41541_;
wire _41542_;
wire _41543_;
wire _41544_;
wire _41545_;
wire _41546_;
wire _41547_;
wire _41548_;
wire _41549_;
wire _41550_;
wire _41551_;
wire _41552_;
wire _41553_;
wire _41554_;
wire _41555_;
wire _41556_;
wire _41557_;
wire _41558_;
wire _41559_;
wire _41560_;
wire _41561_;
wire _41562_;
wire _41563_;
wire _41564_;
wire _41565_;
wire _41566_;
wire _41567_;
wire _41568_;
wire _41569_;
wire _41570_;
wire _41571_;
wire _41572_;
wire _41573_;
wire _41574_;
wire _41575_;
wire _41576_;
wire _41577_;
wire _41578_;
wire _41579_;
wire _41580_;
wire _41581_;
wire _41582_;
wire _41583_;
wire _41584_;
wire _41585_;
wire _41586_;
wire _41587_;
wire _41588_;
wire _41589_;
wire _41590_;
wire _41591_;
wire _41592_;
wire _41593_;
wire _41594_;
wire _41595_;
wire _41596_;
wire _41597_;
wire _41598_;
wire _41599_;
wire _41600_;
wire _41601_;
wire _41602_;
wire _41603_;
wire _41604_;
wire _41605_;
wire _41606_;
wire _41607_;
wire _41608_;
wire _41609_;
wire _41610_;
wire _41611_;
wire _41612_;
wire _41613_;
wire _41614_;
wire _41615_;
wire _41616_;
wire _41617_;
wire _41618_;
wire _41619_;
wire _41620_;
wire _41621_;
wire _41622_;
wire _41623_;
wire _41624_;
wire _41625_;
wire _41626_;
wire _41627_;
wire _41628_;
wire _41629_;
wire _41630_;
wire _41631_;
wire _41632_;
wire _41633_;
wire _41634_;
wire _41635_;
wire _41636_;
wire _41637_;
wire _41638_;
wire _41639_;
wire _41640_;
wire _41641_;
wire _41642_;
wire _41643_;
wire _41644_;
wire _41645_;
wire _41646_;
wire _41647_;
wire _41648_;
wire _41649_;
wire _41650_;
wire _41651_;
wire _41652_;
wire _41653_;
wire _41654_;
wire _41655_;
wire _41656_;
wire _41657_;
wire _41658_;
wire _41659_;
wire _41660_;
wire _41661_;
wire _41662_;
wire _41663_;
wire _41664_;
wire _41665_;
wire _41666_;
wire _41667_;
wire _41668_;
wire _41669_;
wire _41670_;
wire _41671_;
wire _41672_;
wire _41673_;
wire _41674_;
wire _41675_;
wire _41676_;
wire _41677_;
wire _41678_;
wire _41679_;
wire _41680_;
wire _41681_;
wire _41682_;
wire _41683_;
wire _41684_;
wire _41685_;
wire _41686_;
wire _41687_;
wire _41688_;
wire _41689_;
wire _41690_;
wire _41691_;
wire _41692_;
wire _41693_;
wire _41694_;
wire _41695_;
wire _41696_;
wire _41697_;
wire _41698_;
wire _41699_;
wire _41700_;
wire _41701_;
wire _41702_;
wire _41703_;
wire _41704_;
wire _41705_;
wire _41706_;
wire _41707_;
wire _41708_;
wire _41709_;
wire _41710_;
wire _41711_;
wire _41712_;
wire _41713_;
wire _41714_;
wire _41715_;
wire _41716_;
wire _41717_;
wire _41718_;
wire _41719_;
wire _41720_;
wire _41721_;
wire _41722_;
wire _41723_;
wire _41724_;
wire _41725_;
wire _41726_;
wire _41727_;
wire _41728_;
wire _41729_;
wire _41730_;
wire _41731_;
wire _41732_;
wire _41733_;
wire _41734_;
wire _41735_;
wire _41736_;
wire _41737_;
wire _41738_;
wire _41739_;
wire _41740_;
wire _41741_;
wire _41742_;
wire _41743_;
wire _41744_;
wire _41745_;
wire _41746_;
wire _41747_;
wire _41748_;
wire _41749_;
wire _41750_;
wire _41751_;
wire _41752_;
wire _41753_;
wire _41754_;
wire _41755_;
wire _41756_;
wire _41757_;
wire _41758_;
wire _41759_;
wire _41760_;
wire _41761_;
wire _41762_;
wire _41763_;
wire _41764_;
wire _41765_;
wire _41766_;
wire _41767_;
wire _41768_;
wire _41769_;
wire _41770_;
wire _41771_;
wire _41772_;
wire _41773_;
wire _41774_;
wire _41775_;
wire _41776_;
wire _41777_;
wire _41778_;
wire _41779_;
wire _41780_;
wire _41781_;
wire _41782_;
wire _41783_;
wire _41784_;
wire _41785_;
wire _41786_;
wire _41787_;
wire _41788_;
wire _41789_;
wire _41790_;
wire _41791_;
wire _41792_;
wire _41793_;
wire _41794_;
wire _41795_;
wire _41796_;
wire _41797_;
wire _41798_;
wire _41799_;
wire _41800_;
wire _41801_;
wire _41802_;
wire _41803_;
wire _41804_;
wire _41805_;
wire _41806_;
wire _41807_;
wire _41808_;
wire _41809_;
wire _41810_;
wire _41811_;
wire _41812_;
wire _41813_;
wire _41814_;
wire _41815_;
wire _41816_;
wire _41817_;
wire _41818_;
wire _41819_;
wire _41820_;
wire _41821_;
wire _41822_;
wire _41823_;
wire _41824_;
wire _41825_;
wire _41826_;
wire _41827_;
wire _41828_;
wire _41829_;
wire _41830_;
wire _41831_;
wire _41832_;
wire _41833_;
wire _41834_;
wire _41835_;
wire _41836_;
wire _41837_;
wire _41838_;
wire _41839_;
wire _41840_;
wire _41841_;
wire _41842_;
wire _41843_;
wire _41844_;
wire _41845_;
wire _41846_;
wire _41847_;
wire _41848_;
wire _41849_;
wire _41850_;
wire _41851_;
wire _41852_;
wire _41853_;
wire _41854_;
wire _41855_;
wire _41856_;
wire _41857_;
wire _41858_;
wire _41859_;
wire _41860_;
wire _41861_;
wire _41862_;
wire _41863_;
wire _41864_;
wire _41865_;
wire _41866_;
wire _41867_;
wire _41868_;
wire _41869_;
wire _41870_;
wire _41871_;
wire _41872_;
wire _41873_;
wire _41874_;
wire _41875_;
wire _41876_;
wire _41877_;
wire _41878_;
wire _41879_;
wire _41880_;
wire _41881_;
wire _41882_;
wire _41883_;
wire _41884_;
wire _41885_;
wire _41886_;
wire _41887_;
wire _41888_;
wire _41889_;
wire _41890_;
wire _41891_;
wire _41892_;
wire _41893_;
wire _41894_;
wire _41895_;
wire _41896_;
wire _41897_;
wire _41898_;
wire _41899_;
wire _41900_;
wire _41901_;
wire _41902_;
wire _41903_;
wire _41904_;
wire _41905_;
wire _41906_;
wire _41907_;
wire _41908_;
wire _41909_;
wire _41910_;
wire _41911_;
wire _41912_;
wire _41913_;
wire _41914_;
wire _41915_;
wire _41916_;
wire _41917_;
wire _41918_;
wire _41919_;
wire _41920_;
wire _41921_;
wire _41922_;
wire _41923_;
wire _41924_;
wire _41925_;
wire _41926_;
wire _41927_;
wire _41928_;
wire _41929_;
wire _41930_;
wire _41931_;
wire _41932_;
wire _41933_;
wire _41934_;
wire _41935_;
wire _41936_;
wire _41937_;
wire _41938_;
wire _41939_;
wire _41940_;
wire _41941_;
wire _41942_;
wire _41943_;
wire _41944_;
wire _41945_;
wire _41946_;
wire _41947_;
wire _41948_;
wire _41949_;
wire _41950_;
wire _41951_;
wire _41952_;
wire _41953_;
wire _41954_;
wire _41955_;
wire _41956_;
wire _41957_;
wire _41958_;
wire _41959_;
wire _41960_;
wire _41961_;
wire _41962_;
wire _41963_;
wire _41964_;
wire _41965_;
wire _41966_;
wire _41967_;
wire _41968_;
wire _41969_;
wire _41970_;
wire _41971_;
wire _41972_;
wire _41973_;
wire _41974_;
wire _41975_;
wire _41976_;
wire _41977_;
wire _41978_;
wire _41979_;
wire _41980_;
wire _41981_;
wire _41982_;
wire _41983_;
wire _41984_;
wire _41985_;
wire _41986_;
wire _41987_;
wire _41988_;
wire _41989_;
wire _41990_;
wire _41991_;
wire _41992_;
wire _41993_;
wire _41994_;
wire _41995_;
wire _41996_;
wire _41997_;
wire _41998_;
wire _41999_;
wire _42000_;
wire _42001_;
wire _42002_;
wire _42003_;
wire _42004_;
wire _42005_;
wire _42006_;
wire _42007_;
wire _42008_;
wire _42009_;
wire _42010_;
wire _42011_;
wire _42012_;
wire _42013_;
wire _42014_;
wire _42015_;
wire _42016_;
wire _42017_;
wire _42018_;
wire _42019_;
wire _42020_;
wire _42021_;
wire _42022_;
wire _42023_;
wire _42024_;
wire _42025_;
wire _42026_;
wire _42027_;
wire _42028_;
wire _42029_;
wire _42030_;
wire _42031_;
wire _42032_;
wire _42033_;
wire _42034_;
wire _42035_;
wire _42036_;
wire _42037_;
wire _42038_;
wire _42039_;
wire _42040_;
wire _42041_;
wire _42042_;
wire _42043_;
wire _42044_;
wire _42045_;
wire _42046_;
wire _42047_;
wire _42048_;
wire _42049_;
wire _42050_;
wire _42051_;
wire _42052_;
wire _42053_;
wire _42054_;
wire _42055_;
wire _42056_;
wire _42057_;
wire _42058_;
wire _42059_;
wire _42060_;
wire _42061_;
wire _42062_;
wire _42063_;
wire _42064_;
wire _42065_;
wire _42066_;
wire _42067_;
wire _42068_;
wire _42069_;
wire _42070_;
wire _42071_;
wire _42072_;
wire _42073_;
wire _42074_;
wire _42075_;
wire _42076_;
wire _42077_;
wire _42078_;
wire _42079_;
wire _42080_;
wire _42081_;
wire _42082_;
wire _42083_;
wire _42084_;
wire _42085_;
wire _42086_;
wire _42087_;
wire _42088_;
wire _42089_;
wire _42090_;
wire _42091_;
wire _42092_;
wire _42093_;
wire _42094_;
wire _42095_;
wire _42096_;
wire _42097_;
wire _42098_;
wire _42099_;
wire _42100_;
wire _42101_;
wire _42102_;
wire _42103_;
wire _42104_;
wire _42105_;
wire _42106_;
wire _42107_;
wire _42108_;
wire _42109_;
wire _42110_;
wire _42111_;
wire _42112_;
wire _42113_;
wire _42114_;
wire _42115_;
wire _42116_;
wire _42117_;
wire _42118_;
wire _42119_;
wire _42120_;
wire _42121_;
wire _42122_;
wire _42123_;
wire _42124_;
wire _42125_;
wire _42126_;
wire _42127_;
wire _42128_;
wire _42129_;
wire _42130_;
wire _42131_;
wire _42132_;
wire _42133_;
wire _42134_;
wire _42135_;
wire _42136_;
wire _42137_;
wire _42138_;
wire _42139_;
wire _42140_;
wire _42141_;
wire _42142_;
wire _42143_;
wire _42144_;
wire _42145_;
wire _42146_;
wire _42147_;
wire _42148_;
wire _42149_;
wire _42150_;
wire _42151_;
wire _42152_;
wire _42153_;
wire _42154_;
wire _42155_;
wire _42156_;
wire _42157_;
wire _42158_;
wire _42159_;
wire _42160_;
wire _42161_;
wire _42162_;
wire _42163_;
wire _42164_;
wire _42165_;
wire _42166_;
wire _42167_;
wire _42168_;
wire _42169_;
wire _42170_;
wire _42171_;
wire _42172_;
wire _42173_;
wire _42174_;
wire _42175_;
wire _42176_;
wire _42177_;
wire _42178_;
wire _42179_;
wire _42180_;
wire _42181_;
wire _42182_;
wire _42183_;
wire _42184_;
wire _42185_;
wire _42186_;
wire _42187_;
wire _42188_;
wire _42189_;
wire _42190_;
wire _42191_;
wire _42192_;
wire _42193_;
wire _42194_;
wire _42195_;
wire _42196_;
wire _42197_;
wire _42198_;
wire _42199_;
wire _42200_;
wire _42201_;
wire _42202_;
wire _42203_;
wire _42204_;
wire _42205_;
wire _42206_;
wire _42207_;
wire _42208_;
wire _42209_;
wire _42210_;
wire _42211_;
wire _42212_;
wire _42213_;
wire _42214_;
wire _42215_;
wire _42216_;
wire _42217_;
wire _42218_;
wire _42219_;
wire _42220_;
wire _42221_;
wire _42222_;
wire _42223_;
wire _42224_;
wire _42225_;
wire _42226_;
wire _42227_;
wire _42228_;
wire _42229_;
wire _42230_;
wire _42231_;
wire _42232_;
wire _42233_;
wire _42234_;
wire _42235_;
wire _42236_;
wire _42237_;
wire _42238_;
wire _42239_;
wire _42240_;
wire _42241_;
wire _42242_;
wire _42243_;
wire _42244_;
wire _42245_;
wire _42246_;
wire _42247_;
wire _42248_;
wire _42249_;
wire _42250_;
wire _42251_;
wire _42252_;
wire _42253_;
wire _42254_;
wire _42255_;
wire _42256_;
wire _42257_;
wire _42258_;
wire _42259_;
wire _42260_;
wire _42261_;
wire _42262_;
wire _42263_;
wire _42264_;
wire _42265_;
wire _42266_;
wire _42267_;
wire _42268_;
wire _42269_;
wire _42270_;
wire _42271_;
wire _42272_;
wire _42273_;
wire _42274_;
wire _42275_;
wire _42276_;
wire _42277_;
wire _42278_;
wire _42279_;
wire _42280_;
wire _42281_;
wire _42282_;
wire _42283_;
wire _42284_;
wire _42285_;
wire _42286_;
wire _42287_;
wire _42288_;
wire _42289_;
wire _42290_;
wire _42291_;
wire _42292_;
wire _42293_;
wire _42294_;
wire _42295_;
wire _42296_;
wire _42297_;
wire _42298_;
wire _42299_;
wire _42300_;
wire _42301_;
wire _42302_;
wire _42303_;
wire _42304_;
wire _42305_;
wire _42306_;
wire _42307_;
wire _42308_;
wire _42309_;
wire _42310_;
wire _42311_;
wire _42312_;
wire _42313_;
wire _42314_;
wire _42315_;
wire _42316_;
wire _42317_;
wire _42318_;
wire _42319_;
wire _42320_;
wire _42321_;
wire _42322_;
wire _42323_;
wire _42324_;
wire _42325_;
wire _42326_;
wire _42327_;
wire _42328_;
wire _42329_;
wire _42330_;
wire _42331_;
wire _42332_;
wire _42333_;
wire _42334_;
wire _42335_;
wire _42336_;
wire _42337_;
wire _42338_;
wire _42339_;
wire _42340_;
wire _42341_;
wire _42342_;
wire _42343_;
wire _42344_;
wire _42345_;
wire _42346_;
wire _42347_;
wire _42348_;
wire _42349_;
wire _42350_;
wire _42351_;
wire _42352_;
wire _42353_;
wire _42354_;
wire _42355_;
wire _42356_;
wire _42357_;
wire _42358_;
wire _42359_;
wire _42360_;
wire _42361_;
wire _42362_;
wire _42363_;
wire _42364_;
wire _42365_;
wire _42366_;
wire _42367_;
wire _42368_;
wire _42369_;
wire _42370_;
wire _42371_;
wire _42372_;
wire _42373_;
wire _42374_;
wire _42375_;
wire _42376_;
wire _42377_;
wire _42378_;
wire _42379_;
wire _42380_;
wire _42381_;
wire _42382_;
wire _42383_;
wire _42384_;
wire _42385_;
wire _42386_;
wire _42387_;
wire _42388_;
wire _42389_;
wire _42390_;
wire _42391_;
wire _42392_;
wire _42393_;
wire _42394_;
wire _42395_;
wire _42396_;
wire _42397_;
wire _42398_;
wire _42399_;
wire _42400_;
wire _42401_;
wire _42402_;
wire _42403_;
wire _42404_;
wire _42405_;
wire _42406_;
wire _42407_;
wire _42408_;
wire _42409_;
wire _42410_;
wire _42411_;
wire _42412_;
wire _42413_;
wire _42414_;
wire _42415_;
wire _42416_;
wire _42417_;
wire _42418_;
wire _42419_;
wire _42420_;
wire _42421_;
wire _42422_;
wire _42423_;
wire _42424_;
wire _42425_;
wire _42426_;
wire _42427_;
wire _42428_;
wire _42429_;
wire _42430_;
wire _42431_;
wire _42432_;
wire _42433_;
wire _42434_;
wire _42435_;
wire _42436_;
wire _42437_;
wire _42438_;
wire _42439_;
wire _42440_;
wire _42441_;
wire _42442_;
wire _42443_;
wire _42444_;
wire _42445_;
wire _42446_;
wire _42447_;
wire _42448_;
wire _42449_;
wire _42450_;
wire _42451_;
wire _42452_;
wire _42453_;
wire _42454_;
wire _42455_;
wire _42456_;
wire _42457_;
wire _42458_;
wire _42459_;
wire _42460_;
wire _42461_;
wire _42462_;
wire _42463_;
wire _42464_;
wire _42465_;
wire _42466_;
wire _42467_;
wire _42468_;
wire _42469_;
wire _42470_;
wire _42471_;
wire _42472_;
wire _42473_;
wire _42474_;
wire _42475_;
wire _42476_;
wire _42477_;
wire _42478_;
wire _42479_;
wire _42480_;
wire _42481_;
wire _42482_;
wire _42483_;
wire _42484_;
wire _42485_;
wire _42486_;
wire _42487_;
wire _42488_;
wire _42489_;
wire _42490_;
wire _42491_;
wire _42492_;
wire _42493_;
wire _42494_;
wire _42495_;
wire _42496_;
wire _42497_;
wire _42498_;
wire _42499_;
wire _42500_;
wire _42501_;
wire _42502_;
wire _42503_;
wire _42504_;
wire _42505_;
wire _42506_;
wire _42507_;
wire _42508_;
wire _42509_;
wire _42510_;
wire _42511_;
wire _42512_;
wire _42513_;
wire _42514_;
wire _42515_;
wire _42516_;
wire _42517_;
wire _42518_;
wire _42519_;
wire _42520_;
wire _42521_;
wire _42522_;
wire _42523_;
wire _42524_;
wire _42525_;
wire _42526_;
wire _42527_;
wire _42528_;
wire _42529_;
wire _42530_;
wire _42531_;
wire _42532_;
wire _42533_;
wire _42534_;
wire _42535_;
wire _42536_;
wire _42537_;
wire _42538_;
wire _42539_;
wire _42540_;
wire _42541_;
wire _42542_;
wire _42543_;
wire _42544_;
wire _42545_;
wire _42546_;
wire _42547_;
wire _42548_;
wire _42549_;
wire _42550_;
wire _42551_;
wire _42552_;
wire _42553_;
wire _42554_;
wire _42555_;
wire _42556_;
wire _42557_;
wire _42558_;
wire _42559_;
wire _42560_;
wire _42561_;
wire _42562_;
wire _42563_;
wire _42564_;
wire _42565_;
wire _42566_;
wire _42567_;
wire _42568_;
wire _42569_;
wire _42570_;
wire _42571_;
wire _42572_;
wire _42573_;
wire _42574_;
wire _42575_;
wire _42576_;
wire _42577_;
wire _42578_;
wire _42579_;
wire _42580_;
wire _42581_;
wire _42582_;
wire _42583_;
wire _42584_;
wire _42585_;
wire _42586_;
wire _42587_;
wire _42588_;
wire _42589_;
wire _42590_;
wire _42591_;
wire _42592_;
wire _42593_;
wire _42594_;
wire _42595_;
wire _42596_;
wire _42597_;
wire _42598_;
wire _42599_;
wire _42600_;
wire _42601_;
wire _42602_;
wire _42603_;
wire _42604_;
wire _42605_;
wire _42606_;
wire _42607_;
wire _42608_;
wire _42609_;
wire _42610_;
wire _42611_;
wire _42612_;
wire _42613_;
wire _42614_;
wire _42615_;
wire _42616_;
wire _42617_;
wire _42618_;
wire _42619_;
wire _42620_;
wire _42621_;
wire _42622_;
wire _42623_;
wire _42624_;
wire _42625_;
wire _42626_;
wire _42627_;
wire _42628_;
wire _42629_;
wire _42630_;
wire _42631_;
wire _42632_;
wire _42633_;
wire _42634_;
wire _42635_;
wire _42636_;
wire _42637_;
wire _42638_;
wire _42639_;
wire _42640_;
wire _42641_;
wire _42642_;
wire _42643_;
wire _42644_;
wire _42645_;
wire _42646_;
wire _42647_;
wire _42648_;
wire _42649_;
wire _42650_;
wire _42651_;
wire _42652_;
wire _42653_;
wire _42654_;
wire _42655_;
wire _42656_;
wire _42657_;
wire _42658_;
wire _42659_;
wire _42660_;
wire _42661_;
wire _42662_;
wire _42663_;
wire _42664_;
wire _42665_;
wire _42666_;
wire _42667_;
wire _42668_;
wire _42669_;
wire _42670_;
wire _42671_;
wire _42672_;
wire _42673_;
wire _42674_;
wire _42675_;
wire _42676_;
wire _42677_;
wire _42678_;
wire _42679_;
wire _42680_;
wire _42681_;
wire _42682_;
wire _42683_;
wire _42684_;
wire _42685_;
wire _42686_;
wire _42687_;
wire _42688_;
wire _42689_;
wire _42690_;
wire _42691_;
wire _42692_;
wire _42693_;
wire _42694_;
wire _42695_;
wire _42696_;
wire _42697_;
wire _42698_;
wire _42699_;
wire _42700_;
wire _42701_;
wire _42702_;
wire _42703_;
wire _42704_;
wire _42705_;
wire _42706_;
wire _42707_;
wire _42708_;
wire _42709_;
wire _42710_;
wire _42711_;
wire _42712_;
wire _42713_;
wire _42714_;
wire _42715_;
wire _42716_;
wire _42717_;
wire _42718_;
wire _42719_;
wire _42720_;
wire _42721_;
wire _42722_;
wire _42723_;
wire _42724_;
wire _42725_;
wire _42726_;
wire _42727_;
wire _42728_;
wire _42729_;
wire _42730_;
wire _42731_;
wire _42732_;
wire _42733_;
wire _42734_;
wire _42735_;
wire _42736_;
wire _42737_;
wire _42738_;
wire _42739_;
wire _42740_;
wire _42741_;
wire _42742_;
wire _42743_;
wire _42744_;
wire _42745_;
wire _42746_;
wire _42747_;
wire _42748_;
wire _42749_;
wire _42750_;
wire _42751_;
wire _42752_;
wire _42753_;
wire _42754_;
wire _42755_;
wire _42756_;
wire _42757_;
wire _42758_;
wire _42759_;
wire _42760_;
wire _42761_;
wire _42762_;
wire _42763_;
wire _42764_;
wire _42765_;
wire _42766_;
wire _42767_;
wire _42768_;
wire _42769_;
wire _42770_;
wire _42771_;
wire _42772_;
wire _42773_;
wire _42774_;
wire _42775_;
wire _42776_;
wire _42777_;
wire _42778_;
wire _42779_;
wire _42780_;
wire _42781_;
wire _42782_;
wire _42783_;
wire _42784_;
wire _42785_;
wire _42786_;
wire _42787_;
wire _42788_;
wire _42789_;
wire _42790_;
wire _42791_;
wire _42792_;
wire _42793_;
wire _42794_;
wire _42795_;
wire _42796_;
wire _42797_;
wire _42798_;
wire _42799_;
wire _42800_;
wire _42801_;
wire _42802_;
wire _42803_;
wire _42804_;
wire _42805_;
wire _42806_;
wire _42807_;
wire _42808_;
wire _42809_;
wire _42810_;
wire _42811_;
wire _42812_;
wire _42813_;
wire _42814_;
wire _42815_;
wire _42816_;
wire _42817_;
wire _42818_;
wire _42819_;
wire _42820_;
wire _42821_;
wire _42822_;
wire _42823_;
wire _42824_;
wire _42825_;
wire _42826_;
wire _42827_;
wire _42828_;
wire _42829_;
wire _42830_;
wire _42831_;
wire _42832_;
wire _42833_;
wire _42834_;
wire _42835_;
wire _42836_;
wire _42837_;
wire _42838_;
wire _42839_;
wire _42840_;
wire _42841_;
wire _42842_;
wire _42843_;
wire _42844_;
wire _42845_;
wire _42846_;
wire _42847_;
wire _42848_;
wire _42849_;
wire _42850_;
wire _42851_;
wire _42852_;
wire _42853_;
wire _42854_;
wire _42855_;
wire _42856_;
wire _42857_;
wire _42858_;
wire _42859_;
wire _42860_;
wire _42861_;
wire _42862_;
wire _42863_;
wire _42864_;
wire _42865_;
wire _42866_;
wire _42867_;
wire _42868_;
wire _42869_;
wire _42870_;
wire _42871_;
wire _42872_;
wire _42873_;
wire _42874_;
wire _42875_;
wire _42876_;
wire _42877_;
wire _42878_;
wire _42879_;
wire _42880_;
wire _42881_;
wire _42882_;
wire _42883_;
wire _42884_;
wire _42885_;
wire _42886_;
wire _42887_;
wire _42888_;
wire _42889_;
wire _42890_;
wire _42891_;
wire _42892_;
wire _42893_;
wire _42894_;
wire _42895_;
wire _42896_;
wire _42897_;
wire _42898_;
wire _42899_;
wire _42900_;
wire _42901_;
wire _42902_;
wire _42903_;
wire _42904_;
wire _42905_;
wire _42906_;
wire _42907_;
wire _42908_;
wire _42909_;
wire _42910_;
wire _42911_;
wire _42912_;
wire _42913_;
wire _42914_;
wire _42915_;
wire _42916_;
wire _42917_;
wire _42918_;
wire _42919_;
wire _42920_;
wire _42921_;
wire _42922_;
wire _42923_;
wire _42924_;
wire _42925_;
wire _42926_;
wire _42927_;
wire _42928_;
wire _42929_;
wire _42930_;
wire _42931_;
wire _42932_;
wire _42933_;
wire _42934_;
wire _42935_;
wire _42936_;
wire _42937_;
wire _42938_;
wire _42939_;
wire _42940_;
wire _42941_;
wire _42942_;
wire _42943_;
wire _42944_;
wire _42945_;
wire _42946_;
wire _42947_;
wire _42948_;
wire _42949_;
wire _42950_;
wire _42951_;
wire _42952_;
wire _42953_;
wire _42954_;
wire _42955_;
wire _42956_;
wire _42957_;
wire _42958_;
wire _42959_;
wire _42960_;
wire _42961_;
wire _42962_;
wire _42963_;
wire _42964_;
wire _42965_;
wire _42966_;
wire _42967_;
wire _42968_;
wire _42969_;
wire _42970_;
wire _42971_;
wire _42972_;
wire _42973_;
wire _42974_;
wire _42975_;
wire _42976_;
wire _42977_;
wire _42978_;
wire _42979_;
wire _42980_;
wire _42981_;
wire _42982_;
wire _42983_;
wire _42984_;
wire _42985_;
wire _42986_;
wire _42987_;
wire _42988_;
wire _42989_;
wire _42990_;
wire _42991_;
wire _42992_;
wire _42993_;
wire _42994_;
wire _42995_;
wire _42996_;
wire _42997_;
wire _42998_;
wire _42999_;
wire _43000_;
wire _43001_;
wire _43002_;
wire _43003_;
wire _43004_;
wire _43005_;
wire _43006_;
wire _43007_;
wire _43008_;
wire _43009_;
wire _43010_;
wire _43011_;
wire _43012_;
wire _43013_;
wire _43014_;
wire _43015_;
wire _43016_;
wire _43017_;
wire _43018_;
wire _43019_;
wire _43020_;
wire _43021_;
wire _43022_;
wire _43023_;
wire _43024_;
wire _43025_;
wire _43026_;
wire _43027_;
wire _43028_;
wire _43029_;
wire _43030_;
wire _43031_;
wire _43032_;
wire _43033_;
wire _43034_;
wire _43035_;
wire _43036_;
wire _43037_;
wire _43038_;
wire _43039_;
wire _43040_;
wire _43041_;
wire _43042_;
wire _43043_;
wire _43044_;
wire _43045_;
wire _43046_;
wire _43047_;
wire _43048_;
wire _43049_;
wire _43050_;
wire _43051_;
wire _43052_;
wire _43053_;
wire _43054_;
wire _43055_;
wire _43056_;
wire _43057_;
wire _43058_;
wire _43059_;
wire _43060_;
wire _43061_;
wire _43062_;
wire _43063_;
wire _43064_;
wire _43065_;
wire _43066_;
wire _43067_;
wire _43068_;
wire _43069_;
wire _43070_;
wire _43071_;
wire _43072_;
wire _43073_;
wire _43074_;
wire _43075_;
wire _43076_;
wire _43077_;
wire _43078_;
wire _43079_;
wire _43080_;
wire _43081_;
wire _43082_;
wire _43083_;
wire _43084_;
wire _43085_;
wire _43086_;
wire _43087_;
wire _43088_;
wire _43089_;
wire _43090_;
wire _43091_;
wire _43092_;
wire _43093_;
wire _43094_;
wire _43095_;
wire _43096_;
wire _43097_;
wire _43098_;
wire _43099_;
wire _43100_;
wire _43101_;
wire _43102_;
wire _43103_;
wire _43104_;
wire _43105_;
wire _43106_;
wire _43107_;
wire _43108_;
wire _43109_;
wire _43110_;
wire _43111_;
wire _43112_;
wire _43113_;
wire _43114_;
wire _43115_;
wire _43116_;
wire _43117_;
wire _43118_;
wire _43119_;
wire _43120_;
wire _43121_;
wire _43122_;
wire _43123_;
wire _43124_;
wire _43125_;
wire _43126_;
wire _43127_;
wire _43128_;
wire _43129_;
wire _43130_;
wire _43131_;
wire _43132_;
wire _43133_;
wire _43134_;
wire _43135_;
wire _43136_;
wire _43137_;
wire _43138_;
wire _43139_;
wire _43140_;
wire _43141_;
wire _43142_;
wire _43143_;
wire _43144_;
wire _43145_;
wire _43146_;
wire _43147_;
wire _43148_;
wire _43149_;
wire _43150_;
wire _43151_;
wire _43152_;
wire _43153_;
wire _43154_;
wire _43155_;
wire _43156_;
wire _43157_;
wire _43158_;
wire _43159_;
wire _43160_;
wire _43161_;
wire _43162_;
wire _43163_;
wire _43164_;
wire _43165_;
wire _43166_;
wire _43167_;
wire _43168_;
wire _43169_;
wire _43170_;
wire _43171_;
wire _43172_;
wire _43173_;
wire _43174_;
wire _43175_;
wire _43176_;
wire _43177_;
wire _43178_;
wire _43179_;
wire _43180_;
wire _43181_;
wire _43182_;
wire _43183_;
wire _43184_;
wire _43185_;
wire _43186_;
wire _43187_;
wire _43188_;
wire _43189_;
wire _43190_;
wire _43191_;
wire _43192_;
wire _43193_;
wire _43194_;
wire _43195_;
wire _43196_;
wire _43197_;
wire _43198_;
wire _43199_;
wire _43200_;
wire _43201_;
wire _43202_;
wire _43203_;
wire _43204_;
wire _43205_;
wire _43206_;
wire _43207_;
wire _43208_;
wire _43209_;
wire _43210_;
wire _43211_;
wire _43212_;
wire _43213_;
wire _43214_;
wire _43215_;
wire _43216_;
wire _43217_;
wire _43218_;
wire _43219_;
wire _43220_;
wire _43221_;
wire _43222_;
wire _43223_;
wire _43224_;
wire _43225_;
wire _43226_;
wire _43227_;
wire _43228_;
wire _43229_;
wire _43230_;
wire _43231_;
wire _43232_;
wire _43233_;
wire _43234_;
wire _43235_;
wire _43236_;
wire _43237_;
wire _43238_;
wire _43239_;
wire _43240_;
wire _43241_;
wire _43242_;
wire _43243_;
wire _43244_;
wire _43245_;
wire _43246_;
wire _43247_;
wire _43248_;
wire _43249_;
wire _43250_;
wire _43251_;
wire _43252_;
wire _43253_;
wire _43254_;
wire _43255_;
wire _43256_;
wire _43257_;
wire _43258_;
wire _43259_;
wire _43260_;
wire _43261_;
wire _43262_;
wire _43263_;
wire _43264_;
wire _43265_;
wire _43266_;
wire _43267_;
wire _43268_;
wire _43269_;
wire _43270_;
wire _43271_;
wire _43272_;
wire _43273_;
wire _43274_;
wire _43275_;
wire _43276_;
wire _43277_;
wire _43278_;
wire _43279_;
wire _43280_;
wire _43281_;
wire _43282_;
wire _43283_;
wire _43284_;
wire _43285_;
wire _43286_;
wire _43287_;
wire _43288_;
wire _43289_;
wire _43290_;
wire _43291_;
wire _43292_;
wire _43293_;
wire _43294_;
wire _43295_;
wire _43296_;
wire _43297_;
wire _43298_;
wire _43299_;
wire _43300_;
wire _43301_;
wire _43302_;
wire _43303_;
wire _43304_;
wire _43305_;
wire _43306_;
wire _43307_;
wire _43308_;
wire _43309_;
wire _43310_;
wire _43311_;
wire _43312_;
wire _43313_;
wire _43314_;
wire _43315_;
wire _43316_;
wire _43317_;
wire _43318_;
wire _43319_;
wire _43320_;
wire _43321_;
wire _43322_;
wire _43323_;
wire _43324_;
wire _43325_;
wire _43326_;
wire _43327_;
wire _43328_;
wire _43329_;
wire _43330_;
wire _43331_;
wire _43332_;
wire _43333_;
wire _43334_;
wire _43335_;
wire _43336_;
wire _43337_;
wire _43338_;
wire _43339_;
wire _43340_;
wire _43341_;
wire _43342_;
wire _43343_;
wire _43344_;
wire _43345_;
wire _43346_;
wire _43347_;
wire _43348_;
wire _43349_;
wire _43350_;
wire _43351_;
wire _43352_;
wire _43353_;
wire _43354_;
wire _43355_;
wire _43356_;
wire _43357_;
wire _43358_;
wire _43359_;
wire _43360_;
wire _43361_;
wire _43362_;
wire _43363_;
wire _43364_;
wire _43365_;
wire _43366_;
wire _43367_;
wire _43368_;
wire _43369_;
wire _43370_;
wire _43371_;
wire _43372_;
wire _43373_;
wire _43374_;
wire _43375_;
wire _43376_;
wire _43377_;
wire _43378_;
wire _43379_;
wire _43380_;
wire _43381_;
wire _43382_;
wire _43383_;
wire _43384_;
wire _43385_;
wire _43386_;
wire _43387_;
wire _43388_;
wire _43389_;
wire _43390_;
wire _43391_;
wire _43392_;
wire _43393_;
wire _43394_;
wire _43395_;
wire _43396_;
wire _43397_;
wire _43398_;
wire _43399_;
wire _43400_;
wire _43401_;
wire _43402_;
wire _43403_;
wire _43404_;
wire _43405_;
wire _43406_;
wire _43407_;
wire _43408_;
wire _43409_;
wire _43410_;
wire _43411_;
wire _43412_;
wire _43413_;
wire _43414_;
wire _43415_;
wire _43416_;
wire _43417_;
wire _43418_;
wire _43419_;
wire _43420_;
wire _43421_;
wire _43422_;
wire _43423_;
wire _43424_;
wire _43425_;
wire _43426_;
wire _43427_;
wire _43428_;
wire _43429_;
wire _43430_;
wire _43431_;
wire _43432_;
wire _43433_;
wire _43434_;
wire _43435_;
wire _43436_;
wire _43437_;
wire _43438_;
wire _43439_;
wire _43440_;
wire _43441_;
wire _43442_;
wire _43443_;
wire _43444_;
wire _43445_;
wire _43446_;
wire _43447_;
wire _43448_;
wire _43449_;
wire _43450_;
wire _43451_;
wire _43452_;
wire _43453_;
wire _43454_;
wire _43455_;
wire _43456_;
wire _43457_;
wire _43458_;
wire _43459_;
wire _43460_;
wire _43461_;
wire _43462_;
wire _43463_;
wire _43464_;
wire _43465_;
wire _43466_;
wire _43467_;
wire _43468_;
wire _43469_;
wire _43470_;
wire _43471_;
wire _43472_;
wire _43473_;
wire _43474_;
wire _43475_;
wire _43476_;
wire _43477_;
wire _43478_;
wire _43479_;
wire _43480_;
wire _43481_;
wire _43482_;
wire _43483_;
wire _43484_;
wire _43485_;
wire _43486_;
wire _43487_;
wire _43488_;
wire _43489_;
wire _43490_;
wire _43491_;
wire _43492_;
wire _43493_;
wire _43494_;
wire _43495_;
wire _43496_;
wire _43497_;
wire _43498_;
wire _43499_;
wire _43500_;
wire _43501_;
wire _43502_;
wire _43503_;
wire _43504_;
wire _43505_;
wire _43506_;
wire _43507_;
wire _43508_;
wire _43509_;
wire _43510_;
wire _43511_;
wire _43512_;
wire _43513_;
wire _43514_;
wire _43515_;
wire _43516_;
wire _43517_;
wire _43518_;
wire _43519_;
wire _43520_;
wire _43521_;
wire _43522_;
wire _43523_;
wire _43524_;
wire _43525_;
wire _43526_;
wire _43527_;
wire _43528_;
wire _43529_;
wire _43530_;
wire _43531_;
wire _43532_;
wire _43533_;
wire _43534_;
wire _43535_;
wire _43536_;
wire _43537_;
wire _43538_;
wire _43539_;
wire _43540_;
wire _43541_;
wire _43542_;
wire _43543_;
wire _43544_;
wire _43545_;
wire _43546_;
wire _43547_;
wire _43548_;
wire _43549_;
wire _43550_;
wire _43551_;
wire _43552_;
wire _43553_;
wire _43554_;
wire _43555_;
wire _43556_;
wire _43557_;
wire _43558_;
wire _43559_;
wire _43560_;
wire _43561_;
wire _43562_;
wire _43563_;
wire _43564_;
wire _43565_;
wire _43566_;
wire _43567_;
wire _43568_;
wire _43569_;
wire _43570_;
wire _43571_;
wire _43572_;
wire _43573_;
wire _43574_;
wire _43575_;
wire _43576_;
wire _43577_;
wire _43578_;
wire _43579_;
wire _43580_;
wire _43581_;
wire _43582_;
wire _43583_;
wire _43584_;
wire _43585_;
wire _43586_;
wire _43587_;
wire _43588_;
wire _43589_;
wire _43590_;
wire _43591_;
wire _43592_;
wire _43593_;
wire _43594_;
wire _43595_;
wire _43596_;
wire _43597_;
wire _43598_;
wire _43599_;
wire _43600_;
wire _43601_;
wire _43602_;
wire _43603_;
wire _43604_;
wire _43605_;
wire _43606_;
wire _43607_;
wire _43608_;
wire _43609_;
wire _43610_;
wire _43611_;
wire _43612_;
wire _43613_;
wire _43614_;
wire _43615_;
wire _43616_;
wire _43617_;
wire _43618_;
wire _43619_;
wire _43620_;
wire _43621_;
wire _43622_;
wire _43623_;
wire _43624_;
wire _43625_;
wire _43626_;
wire _43627_;
wire _43628_;
wire _43629_;
wire _43630_;
wire _43631_;
wire _43632_;
wire _43633_;
wire _43634_;
wire _43635_;
wire _43636_;
wire _43637_;
wire _43638_;
wire _43639_;
wire _43640_;
wire _43641_;
wire _43642_;
wire _43643_;
wire _43644_;
wire _43645_;
wire _43646_;
wire _43647_;
wire _43648_;
wire _43649_;
wire _43650_;
wire _43651_;
wire _43652_;
wire _43653_;
wire _43654_;
wire _43655_;
wire _43656_;
wire _43657_;
wire _43658_;
wire _43659_;
wire _43660_;
wire _43661_;
wire _43662_;
wire _43663_;
wire _43664_;
wire _43665_;
wire _43666_;
wire _43667_;
wire _43668_;
wire _43669_;
wire _43670_;
wire _43671_;
wire _43672_;
wire _43673_;
wire _43674_;
wire _43675_;
wire _43676_;
wire _43677_;
wire _43678_;
wire _43679_;
wire _43680_;
wire _43681_;
wire _43682_;
wire _43683_;
wire _43684_;
wire _43685_;
wire _43686_;
wire _43687_;
wire _43688_;
wire _43689_;
wire _43690_;
wire _43691_;
wire _43692_;
wire _43693_;
wire _43694_;
wire _43695_;
wire _43696_;
wire _43697_;
wire _43698_;
wire _43699_;
wire _43700_;
wire _43701_;
wire _43702_;
wire _43703_;
wire _43704_;
wire _43705_;
wire _43706_;
wire _43707_;
wire _43708_;
wire _43709_;
wire _43710_;
wire _43711_;
wire _43712_;
wire _43713_;
wire _43714_;
wire _43715_;
wire _43716_;
wire _43717_;
wire _43718_;
wire _43719_;
wire _43720_;
wire _43721_;
wire _43722_;
wire _43723_;
wire _43724_;
wire _43725_;
wire _43726_;
wire _43727_;
wire _43728_;
wire _43729_;
wire _43730_;
wire _43731_;
wire _43732_;
wire _43733_;
wire _43734_;
wire _43735_;
wire _43736_;
wire _43737_;
wire _43738_;
wire _43739_;
wire _43740_;
wire _43741_;
wire _43742_;
wire _43743_;
wire _43744_;
wire _43745_;
wire _43746_;
wire _43747_;
wire _43748_;
wire _43749_;
wire _43750_;
wire _43751_;
wire _43752_;
wire _43753_;
wire _43754_;
wire _43755_;
wire _43756_;
wire _43757_;
wire _43758_;
wire _43759_;
wire _43760_;
wire _43761_;
wire _43762_;
wire _43763_;
wire _43764_;
wire _43765_;
wire _43766_;
wire _43767_;
wire _43768_;
wire _43769_;
wire _43770_;
wire _43771_;
wire _43772_;
wire _43773_;
wire _43774_;
wire _43775_;
wire _43776_;
wire _43777_;
wire _43778_;
wire _43779_;
wire _43780_;
wire _43781_;
wire _43782_;
wire _43783_;
wire _43784_;
wire _43785_;
wire _43786_;
wire _43787_;
wire _43788_;
wire _43789_;
wire _43790_;
wire _43791_;
wire _43792_;
wire _43793_;
wire _43794_;
wire _43795_;
wire _43796_;
wire _43797_;
wire _43798_;
wire _43799_;
wire _43800_;
wire _43801_;
wire _43802_;
wire _43803_;
wire _43804_;
wire _43805_;
wire _43806_;
wire _43807_;
wire _43808_;
wire _43809_;
wire _43810_;
wire _43811_;
wire _43812_;
wire _43813_;
wire _43814_;
wire _43815_;
wire _43816_;
wire _43817_;
wire _43818_;
wire _43819_;
wire _43820_;
wire _43821_;
wire _43822_;
wire _43823_;
wire _43824_;
wire _43825_;
wire _43826_;
wire _43827_;
wire _43828_;
wire _43829_;
wire _43830_;
wire _43831_;
wire _43832_;
wire _43833_;
wire _43834_;
wire _43835_;
wire _43836_;
wire _43837_;
wire _43838_;
wire _43839_;
wire _43840_;
wire _43841_;
wire _43842_;
wire _43843_;
wire _43844_;
wire _43845_;
wire _43846_;
wire _43847_;
wire _43848_;
wire _43849_;
wire _43850_;
wire _43851_;
wire _43852_;
wire _43853_;
wire _43854_;
wire _43855_;
wire _43856_;
wire _43857_;
wire _43858_;
wire _43859_;
wire _43860_;
wire _43861_;
wire _43862_;
wire _43863_;
wire _43864_;
wire _43865_;
wire _43866_;
wire _43867_;
wire _43868_;
wire _43869_;
wire _43870_;
wire _43871_;
wire _43872_;
wire _43873_;
wire _43874_;
wire _43875_;
wire _43876_;
wire _43877_;
wire _43878_;
wire _43879_;
wire _43880_;
wire _43881_;
wire _43882_;
wire _43883_;
wire _43884_;
wire _43885_;
wire _43886_;
wire _43887_;
wire _43888_;
wire _43889_;
wire _43890_;
wire _43891_;
wire _43892_;
wire _43893_;
wire _43894_;
wire _43895_;
wire _43896_;
wire _43897_;
wire _43898_;
wire _43899_;
wire _43900_;
wire _43901_;
wire _43902_;
wire _43903_;
wire _43904_;
wire _43905_;
wire _43906_;
wire _43907_;
wire _43908_;
wire _43909_;
wire _43910_;
wire _43911_;
wire _43912_;
wire _43913_;
wire _43914_;
wire _43915_;
wire _43916_;
wire _43917_;
wire _43918_;
wire _43919_;
wire _43920_;
wire _43921_;
wire _43922_;
wire _43923_;
wire _43924_;
wire _43925_;
wire _43926_;
wire _43927_;
wire _43928_;
wire _43929_;
wire _43930_;
wire _43931_;
wire _43932_;
wire _43933_;
wire _43934_;
wire _43935_;
wire _43936_;
wire _43937_;
wire _43938_;
wire _43939_;
wire _43940_;
wire _43941_;
wire _43942_;
wire _43943_;
wire _43944_;
wire _43945_;
wire _43946_;
wire _43947_;
wire _43948_;
wire _43949_;
wire _43950_;
wire _43951_;
wire _43952_;
wire _43953_;
wire _43954_;
wire _43955_;
wire _43956_;
wire _43957_;
wire _43958_;
wire _43959_;
wire _43960_;
wire _43961_;
wire _43962_;
wire _43963_;
wire _43964_;
wire _43965_;
wire _43966_;
wire _43967_;
wire _43968_;
wire _43969_;
wire _43970_;
wire _43971_;
wire _43972_;
wire _43973_;
wire _43974_;
wire _43975_;
wire _43976_;
wire _43977_;
wire _43978_;
wire _43979_;
wire _43980_;
wire _43981_;
wire _43982_;
wire _43983_;
wire _43984_;
wire _43985_;
wire _43986_;
wire _43987_;
wire _43988_;
wire _43989_;
wire _43990_;
wire _43991_;
wire _43992_;
wire _43993_;
wire _43994_;
wire _43995_;
wire _43996_;
wire _43997_;
wire _43998_;
wire _43999_;
wire _44000_;
wire _44001_;
wire _44002_;
wire _44003_;
wire _44004_;
wire _44005_;
wire _44006_;
wire _44007_;
wire _44008_;
wire _44009_;
wire _44010_;
wire _44011_;
wire _44012_;
wire _44013_;
wire _44014_;
wire _44015_;
wire _44016_;
wire _44017_;
wire _44018_;
wire _44019_;
wire _44020_;
wire _44021_;
wire _44022_;
wire _44023_;
wire _44024_;
wire _44025_;
wire _44026_;
wire _44027_;
wire _44028_;
wire _44029_;
wire _44030_;
wire _44031_;
wire _44032_;
wire _44033_;
wire _44034_;
wire _44035_;
wire _44036_;
wire _44037_;
wire _44038_;
wire _44039_;
wire _44040_;
wire _44041_;
wire _44042_;
wire _44043_;
wire _44044_;
wire _44045_;
wire _44046_;
wire _44047_;
wire _44048_;
wire _44049_;
wire _44050_;
wire _44051_;
wire _44052_;
wire _44053_;
wire _44054_;
wire _44055_;
wire _44056_;
wire _44057_;
wire _44058_;
wire _44059_;
wire _44060_;
wire _44061_;
wire _44062_;
wire _44063_;
wire _44064_;
wire _44065_;
wire _44066_;
wire _44067_;
wire _44068_;
wire _44069_;
wire _44070_;
wire _44071_;
wire _44072_;
wire _44073_;
wire _44074_;
wire _44075_;
wire _44076_;
wire _44077_;
wire _44078_;
wire _44079_;
wire _44080_;
wire _44081_;
wire _44082_;
wire _44083_;
wire _44084_;
wire _44085_;
wire _44086_;
wire _44087_;
wire _44088_;
wire _44089_;
wire _44090_;
wire _44091_;
wire _44092_;
wire _44093_;
wire _44094_;
wire _44095_;
wire _44096_;
wire _44097_;
wire _44098_;
wire _44099_;
wire _44100_;
wire _44101_;
wire _44102_;
wire _44103_;
wire _44104_;
wire _44105_;
wire _44106_;
wire _44107_;
wire _44108_;
wire _44109_;
wire _44110_;
wire _44111_;
wire _44112_;
wire _44113_;
wire _44114_;
wire _44115_;
wire _44116_;
wire _44117_;
wire _44118_;
wire _44119_;
wire _44120_;
wire _44121_;
wire _44122_;
wire _44123_;
wire _44124_;
wire _44125_;
wire _44126_;
wire _44127_;
wire _44128_;
wire _44129_;
wire _44130_;
wire _44131_;
wire _44132_;
wire _44133_;
wire _44134_;
wire _44135_;
wire _44136_;
wire _44137_;
wire _44138_;
wire _44139_;
wire _44140_;
wire _44141_;
wire _44142_;
wire _44143_;
wire _44144_;
wire _44145_;
wire _44146_;
wire _44147_;
wire _44148_;
wire _44149_;
wire _44150_;
wire _44151_;
wire _44152_;
wire _44153_;
wire _44154_;
wire _44155_;
wire _44156_;
wire _44157_;
wire _44158_;
wire _44159_;
wire _44160_;
wire _44161_;
wire _44162_;
wire _44163_;
wire _44164_;
wire _44165_;
wire _44166_;
wire _44167_;
wire _44168_;
wire _44169_;
wire _44170_;
wire _44171_;
wire _44172_;
wire _44173_;
wire _44174_;
wire _44175_;
wire _44176_;
wire _44177_;
wire _44178_;
wire _44179_;
wire _44180_;
wire _44181_;
wire _44182_;
wire _44183_;
wire _44184_;
wire _44185_;
wire _44186_;
wire _44187_;
wire _44188_;
wire _44189_;
wire _44190_;
wire _44191_;
wire _44192_;
wire _44193_;
wire _44194_;
wire _44195_;
wire _44196_;
wire _44197_;
wire _44198_;
wire _44199_;
wire _44200_;
wire _44201_;
wire _44202_;
wire _44203_;
wire _44204_;
wire _44205_;
wire _44206_;
wire _44207_;
wire _44208_;
wire _44209_;
wire _44210_;
wire _44211_;
wire _44212_;
wire _44213_;
wire _44214_;
wire _44215_;
wire _44216_;
wire _44217_;
wire _44218_;
wire _44219_;
wire _44220_;
wire _44221_;
wire _44222_;
wire _44223_;
wire _44224_;
wire _44225_;
wire _44226_;
wire _44227_;
wire _44228_;
wire _44229_;
wire _44230_;
wire _44231_;
wire _44232_;
wire _44233_;
wire _44234_;
wire _44235_;
wire _44236_;
wire _44237_;
wire _44238_;
wire _44239_;
wire _44240_;
wire _44241_;
wire _44242_;
wire _44243_;
wire _44244_;
wire _44245_;
wire _44246_;
wire _44247_;
wire _44248_;
wire _44249_;
wire _44250_;
wire _44251_;
wire _44252_;
wire _44253_;
wire _44254_;
wire _44255_;
wire _44256_;
wire _44257_;
wire _44258_;
wire _44259_;
wire _44260_;
wire _44261_;
wire _44262_;
wire _44263_;
wire _44264_;
wire _44265_;
wire _44266_;
wire _44267_;
wire _44268_;
wire _44269_;
wire _44270_;
wire _44271_;
wire _44272_;
wire _44273_;
wire _44274_;
wire _44275_;
wire _44276_;
wire _44277_;
wire _44278_;
wire _44279_;
wire _44280_;
wire _44281_;
wire _44282_;
wire _44283_;
wire _44284_;
wire _44285_;
wire _44286_;
wire _44287_;
wire _44288_;
wire _44289_;
wire _44290_;
wire _44291_;
wire _44292_;
wire _44293_;
wire _44294_;
wire _44295_;
wire _44296_;
wire _44297_;
wire _44298_;
wire _44299_;
wire _44300_;
wire _44301_;
wire _44302_;
wire _44303_;
wire _44304_;
wire _44305_;
wire _44306_;
wire _44307_;
wire _44308_;
wire _44309_;
wire _44310_;
wire _44311_;
wire _44312_;
wire _44313_;
wire _44314_;
wire _44315_;
wire _44316_;
wire _44317_;
wire _44318_;
wire _44319_;
wire _44320_;
wire _44321_;
wire _44322_;
wire _44323_;
wire _44324_;
wire _44325_;
wire _44326_;
wire _44327_;
wire _44328_;
wire _44329_;
wire _44330_;
wire _44331_;
wire _44332_;
wire _44333_;
wire _44334_;
wire _44335_;
wire _44336_;
wire _44337_;
wire _44338_;
wire _44339_;
wire _44340_;
wire _44341_;
wire _44342_;
wire _44343_;
wire _44344_;
wire _44345_;
wire _44346_;
wire _44347_;
wire _44348_;
wire _44349_;
wire _44350_;
wire _44351_;
wire _44352_;
wire _44353_;
wire _44354_;
wire _44355_;
wire _44356_;
wire _44357_;
wire _44358_;
wire _44359_;
wire _44360_;
wire _44361_;
wire _44362_;
wire _44363_;
wire _44364_;
wire _44365_;
wire _44366_;
wire _44367_;
wire _44368_;
wire _44369_;
wire _44370_;
wire _44371_;
wire _44372_;
wire _44373_;
wire _44374_;
wire _44375_;
wire _44376_;
wire _44377_;
wire _44378_;
wire _44379_;
wire _44380_;
wire _44381_;
wire _44382_;
wire _44383_;
wire _44384_;
wire _44385_;
wire _44386_;
wire _44387_;
wire _44388_;
wire _44389_;
wire _44390_;
wire _44391_;
wire _44392_;
wire _44393_;
wire _44394_;
wire _44395_;
wire _44396_;
wire _44397_;
wire _44398_;
wire _44399_;
wire _44400_;
wire _44401_;
wire _44402_;
wire _44403_;
wire _44404_;
wire _44405_;
wire _44406_;
wire _44407_;
wire _44408_;
wire _44409_;
wire _44410_;
wire _44411_;
wire _44412_;
wire _44413_;
wire _44414_;
wire _44415_;
wire _44416_;
wire _44417_;
wire _44418_;
wire _44419_;
wire _44420_;
wire _44421_;
wire _44422_;
wire _44423_;
wire _44424_;
wire _44425_;
wire _44426_;
wire _44427_;
wire _44428_;
wire _44429_;
wire _44430_;
wire _44431_;
wire _44432_;
wire _44433_;
wire _44434_;
wire _44435_;
wire _44436_;
wire _44437_;
wire _44438_;
wire _44439_;
wire _44440_;
wire _44441_;
wire _44442_;
wire _44443_;
wire _44444_;
wire _44445_;
wire _44446_;
wire _44447_;
wire _44448_;
wire _44449_;
wire _44450_;
wire _44451_;
wire _44452_;
wire _44453_;
wire _44454_;
wire _44455_;
wire _44456_;
wire _44457_;
wire _44458_;
wire _44459_;
wire _44460_;
wire _44461_;
wire _44462_;
wire _44463_;
wire _44464_;
wire _44465_;
wire _44466_;
wire _44467_;
wire _44468_;
wire _44469_;
wire _44470_;
wire _44471_;
wire _44472_;
wire _44473_;
wire _44474_;
wire _44475_;
wire _44476_;
wire _44477_;
wire _44478_;
wire _44479_;
wire _44480_;
wire _44481_;
wire _44482_;
wire _44483_;
wire _44484_;
wire _44485_;
wire _44486_;
wire _44487_;
wire _44488_;
wire _44489_;
wire _44490_;
wire _44491_;
wire _44492_;
wire _44493_;
wire _44494_;
wire _44495_;
wire _44496_;
wire _44497_;
wire _44498_;
wire _44499_;
wire _44500_;
wire _44501_;
wire _44502_;
wire _44503_;
wire _44504_;
wire _44505_;
wire _44506_;
wire _44507_;
wire _44508_;
wire _44509_;
wire _44510_;
wire _44511_;
wire _44512_;
wire _44513_;
wire _44514_;
wire _44515_;
wire _44516_;
wire _44517_;
wire _44518_;
wire _44519_;
wire _44520_;
wire _44521_;
wire _44522_;
wire _44523_;
wire _44524_;
wire _44525_;
wire _44526_;
wire _44527_;
wire _44528_;
wire _44529_;
wire _44530_;
wire _44531_;
wire _44532_;
wire _44533_;
wire _44534_;
wire _44535_;
wire _44536_;
wire _44537_;
wire _44538_;
wire _44539_;
wire _44540_;
wire _44541_;
wire _44542_;
wire _44543_;
wire _44544_;
wire _44545_;
wire _44546_;
wire _44547_;
wire _44548_;
wire _44549_;
wire _44550_;
wire _44551_;
wire _44552_;
wire _44553_;
wire _44554_;
wire _44555_;
wire _44556_;
wire _44557_;
wire _44558_;
wire _44559_;
wire _44560_;
wire _44561_;
wire _44562_;
wire _44563_;
wire _44564_;
wire _44565_;
wire _44566_;
wire _44567_;
wire _44568_;
wire _44569_;
wire _44570_;
wire _44571_;
wire _44572_;
wire _44573_;
wire _44574_;
wire _44575_;
wire _44576_;
wire _44577_;
wire _44578_;
wire _44579_;
wire _44580_;
wire _44581_;
wire _44582_;
wire _44583_;
wire _44584_;
wire _44585_;
wire _44586_;
wire _44587_;
wire _44588_;
wire _44589_;
wire _44590_;
wire _44591_;
wire _44592_;
wire _44593_;
wire _44594_;
wire _44595_;
wire _44596_;
wire _44597_;
wire _44598_;
wire _44599_;
wire _44600_;
wire _44601_;
wire _44602_;
wire _44603_;
wire _44604_;
wire _44605_;
wire _44606_;
wire _44607_;
wire _44608_;
wire _44609_;
wire _44610_;
wire _44611_;
wire _44612_;
wire _44613_;
wire _44614_;
wire _44615_;
wire _44616_;
wire _44617_;
wire _44618_;
wire _44619_;
wire _44620_;
wire _44621_;
wire _44622_;
wire _44623_;
wire _44624_;
wire _44625_;
wire _44626_;
wire _44627_;
wire _44628_;
wire _44629_;
wire _44630_;
wire _44631_;
wire _44632_;
wire _44633_;
wire _44634_;
wire _44635_;
wire _44636_;
wire _44637_;
wire _44638_;
wire _44639_;
wire _44640_;
wire _44641_;
wire _44642_;
wire _44643_;
wire _44644_;
wire _44645_;
wire _44646_;
wire _44647_;
wire _44648_;
wire _44649_;
wire _44650_;
wire _44651_;
wire _44652_;
wire _44653_;
wire _44654_;
wire _44655_;
wire _44656_;
wire _44657_;
wire _44658_;
wire _44659_;
wire _44660_;
wire _44661_;
wire _44662_;
wire _44663_;
wire _44664_;
wire _44665_;
wire _44666_;
wire _44667_;
wire _44668_;
wire _44669_;
wire _44670_;
wire _44671_;
wire _44672_;
wire _44673_;
wire _44674_;
wire _44675_;
wire _44676_;
wire _44677_;
wire _44678_;
wire _44679_;
wire _44680_;
wire _44681_;
wire _44682_;
wire _44683_;
wire _44684_;
wire _44685_;
wire _44686_;
wire _44687_;
wire _44688_;
wire _44689_;
wire _44690_;
wire _44691_;
wire _44692_;
wire _44693_;
wire _44694_;
wire _44695_;
wire _44696_;
wire _44697_;
wire _44698_;
wire _44699_;
wire _44700_;
wire _44701_;
wire _44702_;
wire _44703_;
wire _44704_;
wire _44705_;
wire _44706_;
wire _44707_;
wire _44708_;
wire _44709_;
wire _44710_;
wire _44711_;
wire _44712_;
wire _44713_;
wire _44714_;
wire _44715_;
wire _44716_;
wire _44717_;
wire _44718_;
wire _44719_;
wire _44720_;
wire _44721_;
wire _44722_;
wire _44723_;
wire _44724_;
wire _44725_;
wire _44726_;
wire _44727_;
wire _44728_;
wire _44729_;
wire _44730_;
wire _44731_;
wire _44732_;
wire _44733_;
wire _44734_;
wire _44735_;
wire _44736_;
wire _44737_;
wire _44738_;
wire _44739_;
wire _44740_;
wire _44741_;
wire _44742_;
wire _44743_;
wire _44744_;
wire _44745_;
wire _44746_;
wire _44747_;
wire _44748_;
wire _44749_;
wire _44750_;
wire _44751_;
wire _44752_;
wire _44753_;
wire _44754_;
wire _44755_;
wire _44756_;
wire _44757_;
wire _44758_;
wire _44759_;
wire _44760_;
wire _44761_;
wire _44762_;
wire _44763_;
wire _44764_;
wire _44765_;
wire _44766_;
wire _44767_;
wire _44768_;
wire _44769_;
wire _44770_;
wire _44771_;
wire _44772_;
wire _44773_;
wire _44774_;
wire _44775_;
wire _44776_;
wire _44777_;
wire _44778_;
wire _44779_;
wire _44780_;
wire _44781_;
wire _44782_;
wire _44783_;
wire _44784_;
wire _44785_;
wire _44786_;
wire _44787_;
wire _44788_;
wire _44789_;
wire _44790_;
wire _44791_;
wire _44792_;
wire _44793_;
wire _44794_;
wire _44795_;
wire _44796_;
wire _44797_;
wire _44798_;
wire _44799_;
wire _44800_;
wire _44801_;
wire _44802_;
wire _44803_;
wire _44804_;
wire _44805_;
wire _44806_;
wire _44807_;
wire _44808_;
wire _44809_;
wire _44810_;
wire _44811_;
wire _44812_;
wire _44813_;
wire _44814_;
wire _44815_;
wire _44816_;
wire _44817_;
wire _44818_;
wire _44819_;
wire _44820_;
wire _44821_;
wire _44822_;
wire _44823_;
wire _44824_;
wire _44825_;
wire _44826_;
wire _44827_;
wire _44828_;
wire _44829_;
wire _44830_;
wire _44831_;
wire _44832_;
wire _44833_;
wire _44834_;
wire _44835_;
wire _44836_;
wire _44837_;
wire _44838_;
wire _44839_;
wire _44840_;
wire _44841_;
wire _44842_;
wire _44843_;
wire _44844_;
wire _44845_;
wire _44846_;
wire _44847_;
wire _44848_;
wire _44849_;
wire _44850_;
wire _44851_;
wire _44852_;
wire _44853_;
wire _44854_;
wire _44855_;
wire _44856_;
wire _44857_;
wire _44858_;
wire _44859_;
wire _44860_;
wire _44861_;
wire _44862_;
wire _44863_;
wire _44864_;
wire _44865_;
wire _44866_;
wire _44867_;
wire _44868_;
wire _44869_;
wire _44870_;
wire _44871_;
wire _44872_;
wire _44873_;
wire _44874_;
wire _44875_;
wire _44876_;
wire _44877_;
wire _44878_;
wire _44879_;
wire _44880_;
wire _44881_;
wire _44882_;
wire _44883_;
wire _44884_;
wire _44885_;
wire _44886_;
wire _44887_;
wire _44888_;
wire _44889_;
wire _44890_;
wire _44891_;
wire _44892_;
wire _44893_;
wire _44894_;
wire _44895_;
wire _44896_;
wire _44897_;
wire _44898_;
wire _44899_;
wire _44900_;
wire _44901_;
wire _44902_;
wire _44903_;
wire _44904_;
wire _44905_;
wire _44906_;
wire _44907_;
wire _44908_;
wire _44909_;
wire _44910_;
wire _44911_;
wire _44912_;
wire _44913_;
wire _44914_;
wire _44915_;
wire _44916_;
wire _44917_;
wire _44918_;
wire _44919_;
wire _44920_;
wire _44921_;
wire _44922_;
wire _44923_;
wire _44924_;
wire _44925_;
wire _44926_;
wire _44927_;
wire _44928_;
wire _44929_;
wire _44930_;
wire _44931_;
wire _44932_;
wire _44933_;
wire _44934_;
wire _44935_;
wire _44936_;
wire _44937_;
wire _44938_;
wire _44939_;
wire _44940_;
wire _44941_;
wire _44942_;
wire _44943_;
wire _44944_;
wire _44945_;
wire _44946_;
wire _44947_;
wire _44948_;
wire _44949_;
wire _44950_;
wire _44951_;
wire _44952_;
wire _44953_;
wire _44954_;
wire _44955_;
wire _44956_;
wire _44957_;
wire _44958_;
wire _44959_;
wire _44960_;
wire _44961_;
wire _44962_;
wire _44963_;
wire _44964_;
wire _44965_;
wire _44966_;
wire _44967_;
wire _44968_;
wire _44969_;
wire _44970_;
wire _44971_;
wire _44972_;
wire _44973_;
wire _44974_;
wire _44975_;
wire _44976_;
wire _44977_;
wire _44978_;
wire _44979_;
wire _44980_;
wire _44981_;
wire _44982_;
wire _44983_;
wire _44984_;
wire _44985_;
wire _44986_;
wire _44987_;
wire _44988_;
wire _44989_;
wire _44990_;
wire _44991_;
wire _44992_;
wire _44993_;
wire _44994_;
wire _44995_;
wire _44996_;
wire _44997_;
wire _44998_;
wire _44999_;
wire _45000_;
wire _45001_;
wire _45002_;
wire _45003_;
wire _45004_;
wire _45005_;
wire _45006_;
wire _45007_;
wire _45008_;
wire _45009_;
wire _45010_;
wire _45011_;
wire _45012_;
wire _45013_;
wire _45014_;
wire _45015_;
wire _45016_;
wire _45017_;
wire _45018_;
wire _45019_;
wire _45020_;
wire _45021_;
wire _45022_;
wire _45023_;
wire _45024_;
wire _45025_;
wire _45026_;
wire _45027_;
wire _45028_;
wire _45029_;
wire _45030_;
wire _45031_;
wire _45032_;
wire _45033_;
wire _45034_;
wire _45035_;
wire _45036_;
wire _45037_;
wire _45038_;
wire _45039_;
wire _45040_;
wire _45041_;
wire _45042_;
wire _45043_;
wire _45044_;
wire _45045_;
wire _45046_;
wire _45047_;
wire _45048_;
wire _45049_;
wire _45050_;
wire _45051_;
wire _45052_;
wire _45053_;
wire _45054_;
wire _45055_;
wire _45056_;
wire _45057_;
wire _45058_;
wire _45059_;
wire _45060_;
wire _45061_;
wire _45062_;
wire _45063_;
wire _45064_;
wire _45065_;
wire _45066_;
wire _45067_;
wire _45068_;
wire _45069_;
wire _45070_;
wire _45071_;
wire _45072_;
wire _45073_;
wire _45074_;
wire _45075_;
wire _45076_;
wire _45077_;
wire _45078_;
wire _45079_;
wire _45080_;
wire _45081_;
wire _45082_;
wire _45083_;
wire _45084_;
wire _45085_;
wire _45086_;
wire _45087_;
wire _45088_;
wire _45089_;
wire _45090_;
wire _45091_;
wire _45092_;
wire _45093_;
wire _45094_;
wire _45095_;
wire _45096_;
wire _45097_;
wire _45098_;
wire _45099_;
wire _45100_;
wire _45101_;
wire _45102_;
wire _45103_;
wire _45104_;
wire _45105_;
wire _45106_;
wire _45107_;
wire _45108_;
wire _45109_;
wire _45110_;
wire _45111_;
wire _45112_;
wire _45113_;
wire _45114_;
wire _45115_;
wire _45116_;
wire _45117_;
wire _45118_;
wire _45119_;
wire _45120_;
wire _45121_;
wire _45122_;
wire _45123_;
wire _45124_;
wire _45125_;
wire _45126_;
wire _45127_;
wire _45128_;
wire _45129_;
wire _45130_;
wire _45131_;
wire _45132_;
wire _45133_;
wire _45134_;
wire _45135_;
wire _45136_;
wire _45137_;
wire _45138_;
wire _45139_;
wire _45140_;
wire _45141_;
wire _45142_;
wire _45143_;
wire _45144_;
wire _45145_;
wire _45146_;
wire _45147_;
wire _45148_;
wire _45149_;
wire _45150_;
wire _45151_;
wire _45152_;
wire _45153_;
wire _45154_;
wire _45155_;
wire _45156_;
wire _45157_;
wire _45158_;
wire _45159_;
wire _45160_;
wire _45161_;
wire _45162_;
wire _45163_;
wire _45164_;
wire _45165_;
wire _45166_;
wire _45167_;
wire _45168_;
wire _45169_;
wire _45170_;
wire _45171_;
wire _45172_;
wire _45173_;
wire _45174_;
wire _45175_;
wire _45176_;
wire _45177_;
wire _45178_;
wire _45179_;
wire _45180_;
wire _45181_;
wire _45182_;
wire _45183_;
wire _45184_;
wire _45185_;
wire _45186_;
wire _45187_;
wire _45188_;
wire _45189_;
wire _45190_;
wire _45191_;
wire _45192_;
wire _45193_;
wire _45194_;
wire _45195_;
wire _45196_;
wire _45197_;
wire _45198_;
wire _45199_;
wire _45200_;
wire _45201_;
wire _45202_;
wire _45203_;
wire _45204_;
wire _45205_;
wire _45206_;
wire _45207_;
wire _45208_;
wire _45209_;
wire _45210_;
wire _45211_;
wire _45212_;
wire _45213_;
wire _45214_;
wire _45215_;
wire _45216_;
wire _45217_;
wire _45218_;
wire _45219_;
wire _45220_;
wire _45221_;
wire _45222_;
wire _45223_;
wire _45224_;
wire _45225_;
wire _45226_;
wire _45227_;
wire _45228_;
wire _45229_;
wire _45230_;
wire _45231_;
wire _45232_;
wire _45233_;
wire _45234_;
wire _45235_;
wire _45236_;
wire _45237_;
wire _45238_;
wire _45239_;
wire _45240_;
wire _45241_;
wire _45242_;
wire _45243_;
wire _45244_;
wire _45245_;
wire _45246_;
wire _45247_;
wire _45248_;
wire _45249_;
wire _45250_;
wire _45251_;
wire _45252_;
wire _45253_;
wire _45254_;
wire _45255_;
wire _45256_;
wire _45257_;
wire _45258_;
wire _45259_;
wire _45260_;
wire _45261_;
wire _45262_;
wire _45263_;
wire _45264_;
wire _45265_;
wire _45266_;
wire _45267_;
wire _45268_;
wire _45269_;
wire _45270_;
wire _45271_;
wire _45272_;
wire _45273_;
wire _45274_;
wire _45275_;
wire _45276_;
wire _45277_;
wire _45278_;
wire _45279_;
wire _45280_;
wire _45281_;
wire _45282_;
wire _45283_;
wire _45284_;
wire _45285_;
wire _45286_;
wire _45287_;
wire _45288_;
wire _45289_;
wire _45290_;
wire _45291_;
wire _45292_;
wire _45293_;
wire _45294_;
wire _45295_;
wire _45296_;
wire _45297_;
wire _45298_;
wire _45299_;
wire _45300_;
wire _45301_;
wire _45302_;
wire _45303_;
wire _45304_;
wire _45305_;
wire _45306_;
wire _45307_;
wire _45308_;
wire _45309_;
wire _45310_;
wire _45311_;
wire _45312_;
wire _45313_;
wire _45314_;
wire _45315_;
wire _45316_;
wire _45317_;
wire _45318_;
wire _45319_;
wire _45320_;
wire _45321_;
wire _45322_;
wire _45323_;
wire _45324_;
wire _45325_;
wire _45326_;
wire _45327_;
wire _45328_;
wire _45329_;
wire _45330_;
wire _45331_;
wire _45332_;
wire _45333_;
wire _45334_;
wire _45335_;
wire _45336_;
wire _45337_;
wire _45338_;
wire _45339_;
wire _45340_;
wire _45341_;
wire _45342_;
wire _45343_;
wire _45344_;
wire _45345_;
wire _45346_;
wire _45347_;
wire _45348_;
wire _45349_;
wire _45350_;
wire _45351_;
wire _45352_;
wire _45353_;
wire _45354_;
wire _45355_;
wire _45356_;
wire _45357_;
wire _45358_;
wire _45359_;
wire _45360_;
wire _45361_;
wire _45362_;
wire _45363_;
wire _45364_;
wire _45365_;
wire _45366_;
wire _45367_;
wire _45368_;
wire _45369_;
wire _45370_;
wire _45371_;
wire _45372_;
wire _45373_;
wire _45374_;
wire _45375_;
wire _45376_;
wire _45377_;
wire _45378_;
wire _45379_;
wire _45380_;
wire _45381_;
wire _45382_;
wire _45383_;
wire _45384_;
wire _45385_;
wire _45386_;
wire _45387_;
wire _45388_;
wire _45389_;
wire _45390_;
wire _45391_;
wire _45392_;
wire _45393_;
wire _45394_;
wire _45395_;
wire _45396_;
wire _45397_;
wire _45398_;
wire _45399_;
wire _45400_;
wire _45401_;
wire _45402_;
wire _45403_;
wire _45404_;
wire _45405_;
wire _45406_;
wire _45407_;
wire _45408_;
wire _45409_;
wire _45410_;
wire _45411_;
wire _45412_;
wire _45413_;
wire _45414_;
wire _45415_;
wire _45416_;
wire _45417_;
wire _45418_;
wire _45419_;
wire _45420_;
wire _45421_;
wire _45422_;
wire _45423_;
wire _45424_;
wire _45425_;
wire _45426_;
wire _45427_;
wire _45428_;
wire _45429_;
wire _45430_;
wire _45431_;
wire _45432_;
wire _45433_;
wire _45434_;
wire _45435_;
wire _45436_;
wire _45437_;
wire _45438_;
wire _45439_;
wire _45440_;
wire _45441_;
wire _45442_;
wire _45443_;
wire _45444_;
wire _45445_;
wire _45446_;
wire _45447_;
wire _45448_;
wire _45449_;
wire _45450_;
wire _45451_;
wire _45452_;
wire _45453_;
wire _45454_;
wire _45455_;
wire _45456_;
wire _45457_;
wire _45458_;
wire _45459_;
wire _45460_;
wire _45461_;
wire _45462_;
wire _45463_;
wire _45464_;
wire _45465_;
wire _45466_;
wire _45467_;
wire _45468_;
wire _45469_;
wire _45470_;
wire _45471_;
wire _45472_;
wire _45473_;
wire _45474_;
wire _45475_;
wire _45476_;
wire _45477_;
wire _45478_;
wire _45479_;
wire _45480_;
wire _45481_;
wire _45482_;
wire _45483_;
wire _45484_;
wire _45485_;
wire _45486_;
wire _45487_;
wire _45488_;
wire _45489_;
wire _45490_;
wire _45491_;
wire _45492_;
wire _45493_;
wire _45494_;
wire _45495_;
wire _45496_;
wire _45497_;
wire _45498_;
wire _45499_;
wire _45500_;
wire _45501_;
wire _45502_;
wire _45503_;
wire _45504_;
wire _45505_;
wire _45506_;
wire _45507_;
wire _45508_;
wire _45509_;
wire _45510_;
wire _45511_;
wire _45512_;
wire _45513_;
wire _45514_;
wire _45515_;
wire _45516_;
wire _45517_;
wire _45518_;
wire _45519_;
wire _45520_;
wire _45521_;
wire _45522_;
wire _45523_;
wire _45524_;
wire _45525_;
wire _45526_;
wire _45527_;
wire _45528_;
wire _45529_;
wire _45530_;
wire _45531_;
wire _45532_;
wire _45533_;
wire _45534_;
wire _45535_;
wire _45536_;
wire _45537_;
wire _45538_;
wire _45539_;
wire _45540_;
wire _45541_;
wire _45542_;
wire _45543_;
wire _45544_;
wire _45545_;
wire _45546_;
wire _45547_;
wire _45548_;
wire _45549_;
wire _45550_;
wire _45551_;
wire _45552_;
wire _45553_;
wire _45554_;
wire _45555_;
wire _45556_;
wire _45557_;
wire _45558_;
wire _45559_;
wire _45560_;
wire _45561_;
wire _45562_;
wire _45563_;
wire _45564_;
wire _45565_;
wire _45566_;
wire _45567_;
wire _45568_;
wire _45569_;
wire _45570_;
wire _45571_;
wire _45572_;
wire _45573_;
wire _45574_;
wire _45575_;
wire _45576_;
wire _45577_;
wire _45578_;
wire _45579_;
wire _45580_;
wire _45581_;
wire _45582_;
wire _45583_;
wire _45584_;
wire _45585_;
wire _45586_;
wire _45587_;
wire _45588_;
wire _45589_;
wire _45590_;
wire _45591_;
wire _45592_;
wire _45593_;
wire _45594_;
wire _45595_;
wire _45596_;
wire _45597_;
wire _45598_;
wire _45599_;
wire _45600_;
wire _45601_;
wire _45602_;
wire _45603_;
wire _45604_;
wire _45605_;
wire _45606_;
wire _45607_;
wire _45608_;
wire _45609_;
wire _45610_;
wire _45611_;
wire _45612_;
wire _45613_;
wire _45614_;
wire _45615_;
wire _45616_;
wire _45617_;
wire _45618_;
wire _45619_;
wire _45620_;
wire _45621_;
wire _45622_;
wire _45623_;
wire _45624_;
wire _45625_;
wire _45626_;
wire _45627_;
wire _45628_;
wire _45629_;
wire _45630_;
wire _45631_;
wire _45632_;
wire _45633_;
wire _45634_;
wire _45635_;
wire _45636_;
wire _45637_;
wire _45638_;
wire _45639_;
wire _45640_;
wire _45641_;
wire _45642_;
wire _45643_;
wire _45644_;
wire _45645_;
wire _45646_;
wire _45647_;
wire _45648_;
wire _45649_;
wire _45650_;
wire _45651_;
wire _45652_;
wire _45653_;
wire _45654_;
wire _45655_;
wire _45656_;
wire _45657_;
wire _45658_;
wire _45659_;
wire _45660_;
wire _45661_;
wire _45662_;
wire _45663_;
wire _45664_;
wire _45665_;
wire _45666_;
wire _45667_;
wire _45668_;
wire _45669_;
wire _45670_;
wire _45671_;
wire _45672_;
wire _45673_;
wire _45674_;
wire _45675_;
wire _45676_;
wire _45677_;
wire _45678_;
wire _45679_;
wire _45680_;
wire _45681_;
wire _45682_;
wire _45683_;
wire _45684_;
wire _45685_;
wire _45686_;
wire _45687_;
wire _45688_;
wire _45689_;
wire _45690_;
wire _45691_;
wire _45692_;
wire _45693_;
wire _45694_;
wire _45695_;
wire _45696_;
wire _45697_;
wire _45698_;
wire _45699_;
wire _45700_;
wire _45701_;
wire _45702_;
wire _45703_;
wire _45704_;
wire _45705_;
wire _45706_;
wire _45707_;
wire _45708_;
wire _45709_;
wire _45710_;
wire _45711_;
wire _45712_;
wire _45713_;
wire _45714_;
wire _45715_;
wire _45716_;
wire _45717_;
wire _45718_;
wire _45719_;
wire _45720_;
wire _45721_;
wire _45722_;
wire _45723_;
wire _45724_;
wire _45725_;
wire _45726_;
wire _45727_;
wire _45728_;
wire _45729_;
wire _45730_;
wire _45731_;
wire _45732_;
wire _45733_;
wire _45734_;
wire _45735_;
wire _45736_;
wire _45737_;
wire _45738_;
wire _45739_;
wire _45740_;
wire _45741_;
wire _45742_;
wire _45743_;
wire _45744_;
wire _45745_;
wire _45746_;
wire _45747_;
wire _45748_;
wire _45749_;
wire _45750_;
wire _45751_;
wire _45752_;
wire _45753_;
wire _45754_;
wire _45755_;
wire _45756_;
wire _45757_;
wire _45758_;
wire _45759_;
wire _45760_;
wire _45761_;
wire _45762_;
wire _45763_;
wire _45764_;
wire _45765_;
wire _45766_;
wire _45767_;
wire _45768_;
wire _45769_;
wire _45770_;
wire _45771_;
wire _45772_;
wire _45773_;
wire _45774_;
wire _45775_;
wire _45776_;
wire _45777_;
wire _45778_;
wire _45779_;
wire _45780_;
wire _45781_;
wire _45782_;
wire _45783_;
wire _45784_;
wire _45785_;
wire _45786_;
wire _45787_;
wire _45788_;
wire _45789_;
wire _45790_;
wire _45791_;
wire _45792_;
wire _45793_;
wire _45794_;
wire _45795_;
wire _45796_;
wire _45797_;
wire _45798_;
wire _45799_;
wire _45800_;
wire _45801_;
wire _45802_;
wire _45803_;
wire _45804_;
wire _45805_;
wire _45806_;
wire _45807_;
wire _45808_;
wire _45809_;
wire _45810_;
wire _45811_;
wire _45812_;
wire _45813_;
wire _45814_;
wire _45815_;
wire _45816_;
wire _45817_;
wire _45818_;
wire _45819_;
wire _45820_;
wire _45821_;
wire _45822_;
wire _45823_;
wire _45824_;
wire _45825_;
wire _45826_;
wire _45827_;
wire _45828_;
wire _45829_;
wire _45830_;
wire _45831_;
wire _45832_;
wire _45833_;
wire _45834_;
wire _45835_;
wire _45836_;
wire _45837_;
wire _45838_;
wire _45839_;
wire _45840_;
wire _45841_;
wire _45842_;
wire _45843_;
wire _45844_;
wire _45845_;
wire _45846_;
wire _45847_;
wire _45848_;
wire _45849_;
wire _45850_;
wire _45851_;
wire _45852_;
wire _45853_;
wire _45854_;
wire _45855_;
wire _45856_;
wire _45857_;
wire _45858_;
wire _45859_;
wire _45860_;
wire _45861_;
wire _45862_;
wire _45863_;
wire _45864_;
wire _45865_;
wire _45866_;
wire _45867_;
wire _45868_;
wire _45869_;
wire _45870_;
wire _45871_;
wire _45872_;
wire _45873_;
wire _45874_;
wire _45875_;
wire _45876_;
wire _45877_;
wire _45878_;
wire _45879_;
wire _45880_;
wire _45881_;
wire _45882_;
wire _45883_;
wire _45884_;
wire _45885_;
wire _45886_;
wire _45887_;
wire _45888_;
wire _45889_;
wire _45890_;
wire _45891_;
wire _45892_;
wire _45893_;
wire _45894_;
wire _45895_;
wire _45896_;
wire _45897_;
wire _45898_;
wire _45899_;
wire _45900_;
wire _45901_;
wire _45902_;
wire _45903_;
wire _45904_;
wire _45905_;
wire _45906_;
wire _45907_;
wire _45908_;
wire _45909_;
wire _45910_;
wire _45911_;
wire _45912_;
wire _45913_;
wire _45914_;
wire _45915_;
wire _45916_;
wire _45917_;
wire _45918_;
wire _45919_;
wire _45920_;
wire _45921_;
wire _45922_;
wire _45923_;
wire _45924_;
wire _45925_;
wire _45926_;
wire _45927_;
wire _45928_;
wire _45929_;
wire _45930_;
wire _45931_;
wire _45932_;
wire _45933_;
wire _45934_;
wire _45935_;
wire _45936_;
wire _45937_;
wire _45938_;
wire _45939_;
wire _45940_;
wire _45941_;
wire _45942_;
wire _45943_;
wire _45944_;
wire _45945_;
wire _45946_;
wire _45947_;
wire _45948_;
wire _45949_;
wire _45950_;
wire _45951_;
wire _45952_;
wire _45953_;
wire _45954_;
wire _45955_;
wire _45956_;
wire _45957_;
wire _45958_;
wire _45959_;
wire _45960_;
wire _45961_;
wire _45962_;
wire _45963_;
wire _45964_;
wire _45965_;
wire _45966_;
wire _45967_;
wire _45968_;
wire _45969_;
wire _45970_;
wire _45971_;
wire _45972_;
wire _45973_;
wire _45974_;
wire _45975_;
wire _45976_;
wire _45977_;
wire _45978_;
wire _45979_;
wire _45980_;
wire _45981_;
wire _45982_;
wire _45983_;
wire _45984_;
wire _45985_;
wire _45986_;
wire _45987_;
wire _45988_;
wire _45989_;
wire _45990_;
wire _45991_;
wire _45992_;
wire _45993_;
wire _45994_;
wire _45995_;
wire _45996_;
wire _45997_;
wire _45998_;
wire _45999_;
wire _46000_;
wire _46001_;
wire _46002_;
wire _46003_;
wire _46004_;
wire _46005_;
wire _46006_;
wire _46007_;
wire _46008_;
wire _46009_;
wire _46010_;
wire _46011_;
wire _46012_;
wire _46013_;
wire _46014_;
wire _46015_;
wire _46016_;
wire _46017_;
wire _46018_;
wire _46019_;
wire _46020_;
wire _46021_;
wire _46022_;
wire _46023_;
wire _46024_;
wire _46025_;
wire _46026_;
wire _46027_;
wire _46028_;
wire _46029_;
wire _46030_;
wire _46031_;
wire _46032_;
wire _46033_;
wire _46034_;
wire _46035_;
wire _46036_;
wire _46037_;
wire _46038_;
wire _46039_;
wire _46040_;
wire _46041_;
wire _46042_;
wire _46043_;
wire _46044_;
wire _46045_;
wire _46046_;
wire _46047_;
wire _46048_;
wire _46049_;
wire _46050_;
wire _46051_;
wire _46052_;
wire _46053_;
wire _46054_;
wire _46055_;
wire _46056_;
wire _46057_;
wire _46058_;
wire _46059_;
wire _46060_;
wire _46061_;
wire _46062_;
wire _46063_;
wire _46064_;
wire _46065_;
wire _46066_;
wire _46067_;
wire _46068_;
wire _46069_;
wire _46070_;
wire _46071_;
wire _46072_;
wire _46073_;
wire _46074_;
wire _46075_;
wire _46076_;
wire _46077_;
wire _46078_;
wire _46079_;
wire _46080_;
wire _46081_;
wire _46082_;
wire _46083_;
wire _46084_;
wire _46085_;
wire _46086_;
wire _46087_;
wire _46088_;
wire _46089_;
wire _46090_;
wire _46091_;
wire _46092_;
wire _46093_;
wire _46094_;
wire _46095_;
wire _46096_;
wire _46097_;
wire _46098_;
wire _46099_;
wire _46100_;
wire _46101_;
wire _46102_;
wire _46103_;
wire _46104_;
wire _46105_;
wire _46106_;
wire _46107_;
wire _46108_;
wire _46109_;
wire _46110_;
wire _46111_;
wire _46112_;
wire _46113_;
wire _46114_;
wire _46115_;
wire _46116_;
wire _46117_;
wire _46118_;
wire _46119_;
wire _46120_;
wire _46121_;
wire _46122_;
wire _46123_;
wire _46124_;
wire _46125_;
wire _46126_;
wire _46127_;
wire _46128_;
wire _46129_;
wire _46130_;
wire _46131_;
wire _46132_;
wire _46133_;
wire _46134_;
wire _46135_;
wire _46136_;
wire _46137_;
wire _46138_;
wire _46139_;
wire _46140_;
wire _46141_;
wire _46142_;
wire _46143_;
wire _46144_;
wire _46145_;
wire _46146_;
wire _46147_;
wire _46148_;
wire _46149_;
wire _46150_;
wire _46151_;
wire _46152_;
wire _46153_;
wire _46154_;
wire _46155_;
wire _46156_;
wire _46157_;
wire _46158_;
wire _46159_;
wire _46160_;
wire _46161_;
wire _46162_;
wire _46163_;
wire _46164_;
wire _46165_;
wire _46166_;
wire _46167_;
wire _46168_;
wire _46169_;
wire _46170_;
wire _46171_;
wire _46172_;
wire _46173_;
wire _46174_;
wire _46175_;
wire _46176_;
wire _46177_;
wire _46178_;
wire _46179_;
wire _46180_;
wire _46181_;
wire _46182_;
wire _46183_;
wire _46184_;
wire _46185_;
wire _46186_;
wire _46187_;
wire _46188_;
wire _46189_;
wire _46190_;
wire _46191_;
wire _46192_;
wire _46193_;
wire _46194_;
wire _46195_;
wire _46196_;
wire _46197_;
wire _46198_;
wire _46199_;
wire _46200_;
wire _46201_;
wire _46202_;
wire _46203_;
wire _46204_;
wire _46205_;
wire _46206_;
wire _46207_;
wire _46208_;
wire _46209_;
wire _46210_;
wire _46211_;
wire _46212_;
wire _46213_;
wire _46214_;
wire _46215_;
wire _46216_;
wire _46217_;
wire _46218_;
wire _46219_;
wire _46220_;
wire _46221_;
wire _46222_;
wire _46223_;
wire _46224_;
wire _46225_;
wire _46226_;
wire _46227_;
wire _46228_;
wire _46229_;
wire _46230_;
wire _46231_;
wire _46232_;
wire _46233_;
wire _46234_;
wire _46235_;
wire _46236_;
wire _46237_;
wire _46238_;
wire _46239_;
wire _46240_;
wire _46241_;
wire _46242_;
wire _46243_;
wire _46244_;
wire _46245_;
wire _46246_;
wire _46247_;
wire _46248_;
wire _46249_;
wire _46250_;
wire _46251_;
wire _46252_;
wire _46253_;
wire _46254_;
wire _46255_;
wire _46256_;
wire _46257_;
wire _46258_;
wire _46259_;
wire _46260_;
wire _46261_;
wire _46262_;
wire _46263_;
wire _46264_;
wire _46265_;
wire _46266_;
wire _46267_;
wire _46268_;
wire _46269_;
wire _46270_;
wire _46271_;
wire _46272_;
wire _46273_;
wire _46274_;
wire _46275_;
wire _46276_;
wire _46277_;
wire _46278_;
wire _46279_;
wire _46280_;
wire _46281_;
wire _46282_;
wire _46283_;
wire _46284_;
wire _46285_;
wire _46286_;
wire _46287_;
wire _46288_;
wire _46289_;
wire _46290_;
wire _46291_;
wire _46292_;
wire _46293_;
wire _46294_;
wire _46295_;
wire _46296_;
wire _46297_;
wire _46298_;
wire _46299_;
wire _46300_;
wire _46301_;
wire _46302_;
wire _46303_;
wire _46304_;
wire _46305_;
wire _46306_;
wire _46307_;
wire _46308_;
wire _46309_;
wire _46310_;
wire _46311_;
wire _46312_;
wire _46313_;
wire _46314_;
wire _46315_;
wire _46316_;
wire _46317_;
wire _46318_;
wire _46319_;
wire _46320_;
wire _46321_;
wire _46322_;
wire _46323_;
wire _46324_;
wire _46325_;
wire _46326_;
wire _46327_;
wire _46328_;
wire _46329_;
wire _46330_;
wire _46331_;
wire _46332_;
wire _46333_;
wire _46334_;
wire _46335_;
wire _46336_;
wire _46337_;
wire _46338_;
wire _46339_;
wire _46340_;
wire _46341_;
wire _46342_;
wire _46343_;
wire _46344_;
wire _46345_;
wire _46346_;
wire _46347_;
wire _46348_;
wire _46349_;
wire _46350_;
wire _46351_;
wire _46352_;
wire _46353_;
wire _46354_;
wire _46355_;
wire _46356_;
wire _46357_;
wire _46358_;
wire _46359_;
wire _46360_;
wire _46361_;
wire _46362_;
wire _46363_;
wire _46364_;
wire _46365_;
wire _46366_;
wire _46367_;
wire _46368_;
wire _46369_;
wire _46370_;
wire _46371_;
wire _46372_;
wire _46373_;
wire _46374_;
wire _46375_;
wire _46376_;
wire _46377_;
wire _46378_;
wire _46379_;
wire _46380_;
wire _46381_;
wire _46382_;
wire _46383_;
wire _46384_;
wire _46385_;
wire _46386_;
wire _46387_;
wire _46388_;
wire _46389_;
wire _46390_;
wire _46391_;
wire _46392_;
wire _46393_;
wire _46394_;
wire _46395_;
wire _46396_;
wire _46397_;
wire _46398_;
wire _46399_;
wire _46400_;
wire _46401_;
wire _46402_;
wire _46403_;
wire _46404_;
wire _46405_;
wire _46406_;
wire _46407_;
wire _46408_;
wire _46409_;
wire _46410_;
wire _46411_;
wire _46412_;
wire _46413_;
wire _46414_;
wire _46415_;
wire _46416_;
wire _46417_;
wire _46418_;
wire _46419_;
wire _46420_;
wire _46421_;
wire _46422_;
wire _46423_;
wire _46424_;
wire _46425_;
wire _46426_;
wire _46427_;
wire _46428_;
wire _46429_;
wire _46430_;
wire _46431_;
wire _46432_;
wire _46433_;
wire _46434_;
wire _46435_;
wire _46436_;
wire _46437_;
wire _46438_;
wire _46439_;
wire _46440_;
wire _46441_;
wire _46442_;
wire _46443_;
wire _46444_;
wire _46445_;
wire _46446_;
wire _46447_;
wire _46448_;
wire _46449_;
wire _46450_;
wire _46451_;
wire _46452_;
wire _46453_;
wire _46454_;
wire _46455_;
wire _46456_;
wire _46457_;
wire _46458_;
wire _46459_;
wire _46460_;
wire _46461_;
wire _46462_;
wire _46463_;
wire _46464_;
wire _46465_;
wire _46466_;
wire _46467_;
wire _46468_;
wire _46469_;
wire _46470_;
wire _46471_;
wire _46472_;
wire _46473_;
wire _46474_;
wire _46475_;
wire _46476_;
wire _46477_;
wire _46478_;
wire _46479_;
wire _46480_;
wire _46481_;
wire _46482_;
wire _46483_;
wire _46484_;
wire _46485_;
wire _46486_;
wire _46487_;
wire _46488_;
wire _46489_;
wire _46490_;
wire _46491_;
wire _46492_;
wire _46493_;
wire _46494_;
wire _46495_;
wire _46496_;
wire _46497_;
wire _46498_;
wire _46499_;
wire _46500_;
wire _46501_;
wire _46502_;
wire _46503_;
wire _46504_;
wire _46505_;
wire _46506_;
wire _46507_;
wire _46508_;
wire _46509_;
wire _46510_;
wire _46511_;
wire _46512_;
wire _46513_;
wire _46514_;
wire _46515_;
wire _46516_;
wire _46517_;
wire _46518_;
wire _46519_;
wire _46520_;
wire _46521_;
wire _46522_;
wire _46523_;
wire _46524_;
wire _46525_;
wire _46526_;
wire _46527_;
wire _46528_;
wire _46529_;
wire _46530_;
wire _46531_;
wire _46532_;
wire _46533_;
wire _46534_;
wire _46535_;
wire _46536_;
wire _46537_;
wire _46538_;
wire _46539_;
wire _46540_;
wire _46541_;
wire _46542_;
wire _46543_;
wire _46544_;
wire _46545_;
wire _46546_;
wire _46547_;
wire _46548_;
wire _46549_;
wire _46550_;
wire _46551_;
wire _46552_;
wire _46553_;
wire _46554_;
wire _46555_;
wire _46556_;
wire _46557_;
wire _46558_;
wire _46559_;
wire _46560_;
wire _46561_;
wire _46562_;
wire _46563_;
wire _46564_;
wire _46565_;
wire _46566_;
wire _46567_;
wire _46568_;
wire _46569_;
wire _46570_;
wire _46571_;
wire _46572_;
wire _46573_;
wire _46574_;
wire _46575_;
wire _46576_;
wire _46577_;
wire _46578_;
wire _46579_;
wire _46580_;
wire _46581_;
wire _46582_;
wire _46583_;
wire _46584_;
wire _46585_;
wire _46586_;
wire _46587_;
wire _46588_;
wire _46589_;
wire _46590_;
wire _46591_;
wire _46592_;
wire _46593_;
wire _46594_;
wire _46595_;
wire _46596_;
wire _46597_;
wire _46598_;
wire _46599_;
wire _46600_;
wire _46601_;
wire _46602_;
wire _46603_;
wire _46604_;
wire _46605_;
wire _46606_;
wire _46607_;
wire _46608_;
wire _46609_;
wire _46610_;
wire _46611_;
wire _46612_;
wire _46613_;
wire _46614_;
wire _46615_;
wire _46616_;
wire _46617_;
wire _46618_;
wire _46619_;
wire _46620_;
wire _46621_;
wire _46622_;
wire _46623_;
wire _46624_;
wire _46625_;
wire _46626_;
wire _46627_;
wire _46628_;
wire _46629_;
wire _46630_;
wire _46631_;
wire _46632_;
wire _46633_;
wire _46634_;
wire _46635_;
wire _46636_;
wire _46637_;
wire _46638_;
wire _46639_;
wire _46640_;
wire _46641_;
wire _46642_;
wire _46643_;
wire _46644_;
wire _46645_;
wire _46646_;
wire _46647_;
wire _46648_;
wire _46649_;
wire _46650_;
wire _46651_;
wire _46652_;
wire _46653_;
wire _46654_;
wire _46655_;
wire _46656_;
wire _46657_;
wire _46658_;
wire _46659_;
wire _46660_;
wire _46661_;
wire _46662_;
wire _46663_;
wire _46664_;
wire _46665_;
wire _46666_;
wire _46667_;
wire _46668_;
wire _46669_;
wire _46670_;
wire _46671_;
wire _46672_;
wire _46673_;
wire _46674_;
wire _46675_;
wire _46676_;
wire _46677_;
wire _46678_;
wire _46679_;
wire _46680_;
wire _46681_;
wire _46682_;
wire _46683_;
wire _46684_;
wire _46685_;
wire _46686_;
wire _46687_;
wire _46688_;
wire _46689_;
wire _46690_;
wire _46691_;
wire _46692_;
wire _46693_;
wire _46694_;
wire _46695_;
wire _46696_;
wire _46697_;
wire _46698_;
wire _46699_;
wire _46700_;
wire _46701_;
wire _46702_;
wire _46703_;
wire _46704_;
wire _46705_;
wire _46706_;
wire _46707_;
wire _46708_;
wire _46709_;
wire _46710_;
wire _46711_;
wire _46712_;
wire _46713_;
wire _46714_;
wire _46715_;
wire _46716_;
wire _46717_;
wire _46718_;
wire _46719_;
wire _46720_;
wire _46721_;
wire _46722_;
wire _46723_;
wire _46724_;
wire _46725_;
wire _46726_;
wire _46727_;
wire _46728_;
wire _46729_;
wire _46730_;
wire _46731_;
wire _46732_;
wire _46733_;
wire _46734_;
wire _46735_;
wire _46736_;
wire _46737_;
wire _46738_;
wire _46739_;
wire _46740_;
wire _46741_;
wire _46742_;
wire _46743_;
wire _46744_;
wire _46745_;
wire _46746_;
wire _46747_;
wire _46748_;
wire _46749_;
wire _46750_;
wire _46751_;
wire _46752_;
wire _46753_;
wire _46754_;
wire _46755_;
wire _46756_;
wire _46757_;
wire _46758_;
wire _46759_;
wire _46760_;
wire _46761_;
wire _46762_;
wire _46763_;
wire _46764_;
wire _46765_;
wire _46766_;
wire _46767_;
wire _46768_;
wire _46769_;
wire _46770_;
wire _46771_;
wire _46772_;
wire _46773_;
wire _46774_;
wire _46775_;
wire _46776_;
wire _46777_;
wire _46778_;
wire _46779_;
wire _46780_;
wire _46781_;
wire _46782_;
wire _46783_;
wire _46784_;
wire _46785_;
wire _46786_;
wire _46787_;
wire _46788_;
wire _46789_;
wire _46790_;
wire _46791_;
wire _46792_;
wire _46793_;
wire _46794_;
wire _46795_;
wire _46796_;
wire _46797_;
wire _46798_;
wire _46799_;
wire _46800_;
wire _46801_;
wire _46802_;
wire _46803_;
wire _46804_;
wire _46805_;
wire _46806_;
wire _46807_;
wire _46808_;
wire _46809_;
wire _46810_;
wire _46811_;
wire _46812_;
wire _46813_;
wire _46814_;
wire _46815_;
wire _46816_;
wire _46817_;
wire _46818_;
wire _46819_;
wire _46820_;
wire _46821_;
wire _46822_;
wire _46823_;
wire _46824_;
wire _46825_;
wire _46826_;
wire _46827_;
wire _46828_;
wire _46829_;
wire _46830_;
wire _46831_;
wire _46832_;
wire _46833_;
wire _46834_;
wire _46835_;
wire _46836_;
wire _46837_;
wire _46838_;
wire _46839_;
wire _46840_;
wire _46841_;
wire _46842_;
wire _46843_;
wire _46844_;
wire _46845_;
wire _46846_;
wire _46847_;
wire _46848_;
wire _46849_;
wire _46850_;
wire _46851_;
wire _46852_;
wire _46853_;
wire _46854_;
wire _46855_;
wire _46856_;
wire _46857_;
wire _46858_;
wire _46859_;
wire _46860_;
wire _46861_;
wire _46862_;
wire _46863_;
wire _46864_;
wire _46865_;
wire _46866_;
wire _46867_;
wire _46868_;
wire _46869_;
wire _46870_;
wire _46871_;
wire _46872_;
wire _46873_;
wire _46874_;
wire _46875_;
wire _46876_;
wire _46877_;
wire _46878_;
wire _46879_;
wire _46880_;
wire _46881_;
wire _46882_;
wire _46883_;
wire _46884_;
wire _46885_;
wire _46886_;
wire _46887_;
wire _46888_;
wire _46889_;
wire _46890_;
wire _46891_;
wire _46892_;
wire _46893_;
wire _46894_;
wire _46895_;
wire _46896_;
wire _46897_;
wire _46898_;
wire _46899_;
wire _46900_;
wire _46901_;
wire _46902_;
wire _46903_;
wire _46904_;
wire _46905_;
wire _46906_;
wire _46907_;
wire _46908_;
wire _46909_;
wire _46910_;
wire _46911_;
wire _46912_;
wire _46913_;
wire _46914_;
wire _46915_;
wire _46916_;
wire _46917_;
wire _46918_;
wire _46919_;
wire _46920_;
wire _46921_;
wire _46922_;
wire _46923_;
wire _46924_;
wire _46925_;
wire _46926_;
wire _46927_;
wire _46928_;
wire _46929_;
wire _46930_;
wire _46931_;
wire _46932_;
wire _46933_;
wire _46934_;
wire _46935_;
wire _46936_;
wire _46937_;
wire _46938_;
wire _46939_;
wire _46940_;
wire _46941_;
wire _46942_;
wire _46943_;
wire _46944_;
wire _46945_;
wire _46946_;
wire _46947_;
wire _46948_;
wire _46949_;
wire _46950_;
wire _46951_;
wire _46952_;
wire _46953_;
wire _46954_;
wire _46955_;
wire _46956_;
wire _46957_;
wire _46958_;
wire _46959_;
wire _46960_;
wire _46961_;
wire _46962_;
wire _46963_;
wire _46964_;
wire _46965_;
wire _46966_;
wire _46967_;
wire _46968_;
wire _46969_;
wire _46970_;
wire _46971_;
wire _46972_;
wire _46973_;
wire _46974_;
wire _46975_;
wire _46976_;
wire _46977_;
wire _46978_;
wire _46979_;
wire _46980_;
wire _46981_;
wire _46982_;
wire _46983_;
wire _46984_;
wire _46985_;
wire _46986_;
wire _46987_;
wire _46988_;
wire _46989_;
wire _46990_;
wire _46991_;
wire _46992_;
wire _46993_;
wire _46994_;
wire _46995_;
wire _46996_;
wire _46997_;
wire _46998_;
wire _46999_;
wire _47000_;
wire _47001_;
wire _47002_;
wire _47003_;
wire _47004_;
wire _47005_;
wire _47006_;
wire _47007_;
wire _47008_;
wire _47009_;
wire _47010_;
wire _47011_;
wire _47012_;
wire _47013_;
wire _47014_;
wire _47015_;
wire _47016_;
wire _47017_;
wire _47018_;
wire _47019_;
wire _47020_;
wire _47021_;
wire _47022_;
wire _47023_;
wire _47024_;
wire _47025_;
wire _47026_;
wire _47027_;
wire _47028_;
wire _47029_;
wire _47030_;
wire _47031_;
wire _47032_;
wire _47033_;
wire _47034_;
wire _47035_;
wire _47036_;
wire _47037_;
wire _47038_;
wire _47039_;
wire _47040_;
wire _47041_;
wire _47042_;
wire _47043_;
wire _47044_;
wire _47045_;
wire _47046_;
wire _47047_;
wire _47048_;
wire _47049_;
wire _47050_;
wire _47051_;
wire _47052_;
wire _47053_;
wire _47054_;
wire _47055_;
wire _47056_;
wire _47057_;
wire _47058_;
wire _47059_;
wire _47060_;
wire _47061_;
wire _47062_;
wire _47063_;
wire _47064_;
wire _47065_;
wire _47066_;
wire _47067_;
wire _47068_;
wire _47069_;
wire _47070_;
wire _47071_;
wire _47072_;
wire _47073_;
wire _47074_;
wire _47075_;
wire _47076_;
wire _47077_;
wire _47078_;
wire _47079_;
wire _47080_;
wire _47081_;
wire _47082_;
wire _47083_;
wire _47084_;
wire _47085_;
wire _47086_;
wire _47087_;
wire _47088_;
wire _47089_;
wire _47090_;
wire _47091_;
wire _47092_;
wire _47093_;
wire _47094_;
wire _47095_;
wire _47096_;
wire _47097_;
wire _47098_;
wire _47099_;
wire _47100_;
wire _47101_;
wire _47102_;
wire _47103_;
wire _47104_;
wire _47105_;
wire _47106_;
wire _47107_;
wire _47108_;
wire _47109_;
wire _47110_;
wire _47111_;
wire _47112_;
wire _47113_;
wire _47114_;
wire _47115_;
wire _47116_;
wire _47117_;
wire _47118_;
wire _47119_;
wire _47120_;
wire _47121_;
wire _47122_;
wire _47123_;
wire _47124_;
wire _47125_;
wire _47126_;
wire _47127_;
wire _47128_;
wire _47129_;
wire _47130_;
wire _47131_;
wire _47132_;
wire _47133_;
wire _47134_;
wire _47135_;
wire _47136_;
wire _47137_;
wire _47138_;
wire _47139_;
wire _47140_;
wire _47141_;
wire _47142_;
wire _47143_;
wire _47144_;
wire _47145_;
wire _47146_;
wire _47147_;
wire _47148_;
wire _47149_;
wire _47150_;
wire _47151_;
wire _47152_;
wire _47153_;
wire _47154_;
wire _47155_;
wire _47156_;
wire _47157_;
wire _47158_;
wire _47159_;
wire _47160_;
wire _47161_;
wire _47162_;
wire _47163_;
wire _47164_;
wire _47165_;
wire _47166_;
wire _47167_;
wire _47168_;
wire _47169_;
wire _47170_;
wire _47171_;
wire _47172_;
wire _47173_;
wire _47174_;
wire _47175_;
wire _47176_;
wire _47177_;
wire _47178_;
wire _47179_;
wire _47180_;
wire _47181_;
wire _47182_;
wire _47183_;
wire _47184_;
wire _47185_;
wire _47186_;
wire _47187_;
wire _47188_;
wire _47189_;
wire _47190_;
wire _47191_;
wire _47192_;
wire _47193_;
wire _47194_;
wire _47195_;
wire _47196_;
wire _47197_;
wire _47198_;
wire _47199_;
wire _47200_;
wire _47201_;
wire _47202_;
wire _47203_;
wire _47204_;
wire _47205_;
wire _47206_;
wire _47207_;
wire _47208_;
wire _47209_;
wire _47210_;
wire _47211_;
wire _47212_;
wire _47213_;
wire _47214_;
wire _47215_;
wire _47216_;
wire _47217_;
wire _47218_;
wire _47219_;
wire _47220_;
wire _47221_;
wire _47222_;
wire _47223_;
wire _47224_;
wire _47225_;
wire _47226_;
wire _47227_;
wire _47228_;
wire _47229_;
wire _47230_;
wire _47231_;
wire _47232_;
wire _47233_;
wire _47234_;
wire _47235_;
wire _47236_;
wire _47237_;
wire _47238_;
wire _47239_;
wire _47240_;
wire _47241_;
wire _47242_;
wire _47243_;
wire _47244_;
wire _47245_;
wire _47246_;
wire _47247_;
wire _47248_;
wire _47249_;
wire _47250_;
wire _47251_;
wire _47252_;
wire _47253_;
wire _47254_;
wire _47255_;
wire _47256_;
wire _47257_;
wire _47258_;
wire _47259_;
wire _47260_;
wire _47261_;
wire _47262_;
wire _47263_;
wire _47264_;
wire _47265_;
wire _47266_;
wire _47267_;
wire _47268_;
wire _47269_;
wire _47270_;
wire _47271_;
wire _47272_;
wire _47273_;
wire _47274_;
wire _47275_;
wire _47276_;
wire _47277_;
wire _47278_;
wire _47279_;
wire _47280_;
wire _47281_;
wire _47282_;
wire _47283_;
wire _47284_;
wire _47285_;
wire _47286_;
wire _47287_;
wire _47288_;
wire _47289_;
wire _47290_;
wire _47291_;
wire _47292_;
wire _47293_;
wire _47294_;
wire _47295_;
wire _47296_;
wire _47297_;
wire _47298_;
wire _47299_;
wire _47300_;
wire _47301_;
wire _47302_;
wire _47303_;
wire _47304_;
wire _47305_;
wire _47306_;
wire _47307_;
wire _47308_;
wire _47309_;
wire _47310_;
wire _47311_;
wire _47312_;
wire _47313_;
wire _47314_;
wire _47315_;
wire _47316_;
wire _47317_;
wire _47318_;
wire _47319_;
wire _47320_;
wire _47321_;
wire _47322_;
wire _47323_;
wire _47324_;
wire _47325_;
wire _47326_;
wire _47327_;
wire _47328_;
wire _47329_;
wire _47330_;
wire _47331_;
wire _47332_;
wire _47333_;
wire _47334_;
wire _47335_;
wire _47336_;
wire _47337_;
wire _47338_;
wire _47339_;
wire _47340_;
wire _47341_;
wire _47342_;
wire _47343_;
wire _47344_;
wire _47345_;
wire _47346_;
wire _47347_;
wire _47348_;
wire _47349_;
wire _47350_;
wire _47351_;
wire _47352_;
wire _47353_;
wire _47354_;
wire _47355_;
wire _47356_;
wire _47357_;
wire _47358_;
wire _47359_;
wire _47360_;
wire _47361_;
wire _47362_;
wire _47363_;
wire _47364_;
wire _47365_;
wire _47366_;
wire _47367_;
wire _47368_;
wire _47369_;
wire _47370_;
wire _47371_;
wire _47372_;
wire _47373_;
wire _47374_;
wire _47375_;
wire _47376_;
wire _47377_;
wire _47378_;
wire _47379_;
wire _47380_;
wire _47381_;
wire _47382_;
wire _47383_;
wire _47384_;
wire _47385_;
wire _47386_;
wire _47387_;
wire _47388_;
wire _47389_;
wire _47390_;
wire _47391_;
wire _47392_;
wire _47393_;
wire _47394_;
wire _47395_;
wire _47396_;
wire _47397_;
wire _47398_;
wire _47399_;
wire _47400_;
wire _47401_;
wire _47402_;
wire _47403_;
wire _47404_;
wire _47405_;
wire _47406_;
wire _47407_;
wire _47408_;
wire _47409_;
wire _47410_;
wire _47411_;
wire _47412_;
wire _47413_;
wire _47414_;
wire _47415_;
wire _47416_;
wire _47417_;
wire _47418_;
wire _47419_;
wire _47420_;
wire _47421_;
wire _47422_;
wire _47423_;
wire _47424_;
wire _47425_;
wire _47426_;
wire _47427_;
wire _47428_;
wire _47429_;
wire _47430_;
wire _47431_;
wire _47432_;
wire _47433_;
wire _47434_;
wire _47435_;
wire _47436_;
wire _47437_;
wire _47438_;
wire _47439_;
wire _47440_;
wire _47441_;
wire _47442_;
wire _47443_;
wire _47444_;
wire _47445_;
wire _47446_;
wire _47447_;
wire _47448_;
wire _47449_;
wire _47450_;
wire _47451_;
wire _47452_;
wire _47453_;
wire _47454_;
wire _47455_;
wire _47456_;
wire _47457_;
wire _47458_;
wire _47459_;
wire _47460_;
wire _47461_;
wire _47462_;
wire _47463_;
wire _47464_;
wire _47465_;
wire _47466_;
wire _47467_;
wire _47468_;
wire _47469_;
wire _47470_;
wire _47471_;
wire _47472_;
wire _47473_;
wire _47474_;
wire _47475_;
wire _47476_;
wire _47477_;
wire _47478_;
wire _47479_;
wire _47480_;
wire _47481_;
wire _47482_;
wire _47483_;
wire _47484_;
wire _47485_;
wire _47486_;
wire _47487_;
wire _47488_;
wire _47489_;
wire _47490_;
wire _47491_;
wire _47492_;
wire _47493_;
wire _47494_;
wire _47495_;
wire _47496_;
wire _47497_;
wire _47498_;
wire _47499_;
wire _47500_;
wire _47501_;
wire _47502_;
wire _47503_;
wire _47504_;
wire _47505_;
wire _47506_;
wire _47507_;
wire _47508_;
wire _47509_;
wire _47510_;
wire _47511_;
wire _47512_;
wire _47513_;
wire _47514_;
wire _47515_;
wire _47516_;
wire _47517_;
wire _47518_;
wire _47519_;
wire _47520_;
wire _47521_;
wire _47522_;
wire _47523_;
wire _47524_;
wire _47525_;
wire _47526_;
wire _47527_;
wire _47528_;
wire _47529_;
wire _47530_;
wire _47531_;
wire _47532_;
wire _47533_;
wire _47534_;
wire _47535_;
wire _47536_;
wire _47537_;
wire _47538_;
wire _47539_;
wire _47540_;
wire _47541_;
wire _47542_;
wire _47543_;
wire _47544_;
wire _47545_;
wire _47546_;
wire _47547_;
wire _47548_;
wire _47549_;
wire _47550_;
wire _47551_;
wire _47552_;
wire _47553_;
wire _47554_;
wire _47555_;
wire _47556_;
wire _47557_;
wire _47558_;
wire _47559_;
wire _47560_;
wire _47561_;
wire _47562_;
wire _47563_;
wire _47564_;
wire _47565_;
wire _47566_;
wire _47567_;
wire _47568_;
wire _47569_;
wire _47570_;
wire _47571_;
wire _47572_;
wire _47573_;
wire _47574_;
wire _47575_;
wire _47576_;
wire _47577_;
wire _47578_;
wire _47579_;
wire _47580_;
wire _47581_;
wire _47582_;
wire _47583_;
wire _47584_;
wire _47585_;
wire _47586_;
wire _47587_;
wire _47588_;
wire _47589_;
wire _47590_;
wire _47591_;
wire _47592_;
wire _47593_;
wire _47594_;
wire _47595_;
wire _47596_;
wire _47597_;
wire _47598_;
wire _47599_;
wire _47600_;
wire _47601_;
wire _47602_;
wire _47603_;
wire _47604_;
wire _47605_;
wire _47606_;
wire _47607_;
wire _47608_;
wire _47609_;
wire _47610_;
wire _47611_;
wire _47612_;
wire _47613_;
wire _47614_;
wire _47615_;
wire _47616_;
wire _47617_;
wire _47618_;
wire _47619_;
wire _47620_;
wire _47621_;
wire _47622_;
wire _47623_;
wire _47624_;
wire _47625_;
wire _47626_;
wire _47627_;
wire _47628_;
wire _47629_;
wire _47630_;
wire _47631_;
wire _47632_;
wire _47633_;
wire _47634_;
wire _47635_;
wire _47636_;
wire _47637_;
wire _47638_;
wire _47639_;
wire _47640_;
wire _47641_;
wire _47642_;
wire _47643_;
wire _47644_;
wire _47645_;
wire _47646_;
wire _47647_;
wire _47648_;
wire _47649_;
wire _47650_;
wire _47651_;
wire _47652_;
wire _47653_;
wire _47654_;
wire _47655_;
wire _47656_;
wire _47657_;
wire _47658_;
wire _47659_;
wire _47660_;
wire _47661_;
wire _47662_;
wire _47663_;
wire _47664_;
wire _47665_;
wire _47666_;
wire _47667_;
wire _47668_;
wire _47669_;
wire _47670_;
wire _47671_;
wire _47672_;
wire _47673_;
wire _47674_;
wire _47675_;
wire _47676_;
wire _47677_;
wire _47678_;
wire _47679_;
wire _47680_;
wire _47681_;
wire _47682_;
wire _47683_;
wire _47684_;
wire _47685_;
wire _47686_;
wire _47687_;
wire _47688_;
wire _47689_;
wire _47690_;
wire _47691_;
wire _47692_;
wire _47693_;
wire _47694_;
wire _47695_;
wire _47696_;
wire _47697_;
wire _47698_;
wire _47699_;
wire _47700_;
wire _47701_;
wire _47702_;
wire _47703_;
wire _47704_;
wire _47705_;
wire _47706_;
wire _47707_;
wire _47708_;
wire _47709_;
wire _47710_;
wire _47711_;
wire _47712_;
wire _47713_;
wire _47714_;
wire _47715_;
wire _47716_;
wire _47717_;
wire _47718_;
wire _47719_;
wire _47720_;
wire _47721_;
wire _47722_;
wire _47723_;
wire _47724_;
wire _47725_;
wire _47726_;
wire _47727_;
wire _47728_;
wire _47729_;
wire _47730_;
wire _47731_;
wire _47732_;
wire _47733_;
wire _47734_;
wire _47735_;
wire _47736_;
wire _47737_;
wire _47738_;
wire _47739_;
wire _47740_;
wire _47741_;
wire _47742_;
wire _47743_;
wire _47744_;
wire _47745_;
wire _47746_;
wire _47747_;
wire _47748_;
wire _47749_;
wire _47750_;
wire _47751_;
wire _47752_;
wire _47753_;
wire _47754_;
wire _47755_;
wire _47756_;
wire _47757_;
wire _47758_;
wire _47759_;
wire _47760_;
wire _47761_;
wire _47762_;
wire _47763_;
wire _47764_;
wire _47765_;
wire _47766_;
wire _47767_;
wire _47768_;
wire _47769_;
wire _47770_;
wire _47771_;
wire _47772_;
wire _47773_;
wire _47774_;
wire _47775_;
wire _47776_;
wire _47777_;
wire _47778_;
wire _47779_;
wire _47780_;
wire _47781_;
wire _47782_;
wire _47783_;
wire _47784_;
wire _47785_;
wire _47786_;
wire _47787_;
wire _47788_;
wire _47789_;
wire _47790_;
wire _47791_;
wire _47792_;
wire _47793_;
wire _47794_;
wire _47795_;
wire _47796_;
wire _47797_;
wire _47798_;
wire _47799_;
wire _47800_;
wire _47801_;
wire _47802_;
wire _47803_;
wire _47804_;
wire _47805_;
wire _47806_;
wire _47807_;
wire _47808_;
wire _47809_;
wire _47810_;
wire _47811_;
wire _47812_;
wire _47813_;
wire _47814_;
wire _47815_;
wire _47816_;
wire _47817_;
wire _47818_;
wire _47819_;
wire _47820_;
wire _47821_;
wire _47822_;
wire _47823_;
wire _47824_;
wire _47825_;
wire _47826_;
wire _47827_;
wire _47828_;
wire _47829_;
wire _47830_;
wire _47831_;
wire _47832_;
wire _47833_;
wire _47834_;
wire _47835_;
wire _47836_;
wire _47837_;
wire _47838_;
wire _47839_;
wire _47840_;
wire _47841_;
wire _47842_;
wire _47843_;
wire _47844_;
wire _47845_;
wire _47846_;
wire _47847_;
wire _47848_;
wire _47849_;
wire _47850_;
wire _47851_;
wire _47852_;
wire _47853_;
wire _47854_;
wire _47855_;
wire _47856_;
wire _47857_;
wire _47858_;
wire _47859_;
wire _47860_;
wire _47861_;
wire _47862_;
wire _47863_;
wire _47864_;
wire _47865_;
wire _47866_;
wire _47867_;
wire _47868_;
wire _47869_;
wire _47870_;
wire _47871_;
wire _47872_;
wire _47873_;
wire _47874_;
wire _47875_;
wire _47876_;
wire _47877_;
wire _47878_;
wire _47879_;
wire _47880_;
wire _47881_;
wire _47882_;
wire _47883_;
wire _47884_;
wire _47885_;
wire _47886_;
wire _47887_;
wire _47888_;
wire _47889_;
wire _47890_;
wire _47891_;
wire _47892_;
wire _47893_;
wire _47894_;
wire _47895_;
wire _47896_;
wire _47897_;
wire _47898_;
wire _47899_;
wire _47900_;
wire _47901_;
wire _47902_;
wire _47903_;
wire _47904_;
wire _47905_;
wire _47906_;
wire _47907_;
wire _47908_;
wire _47909_;
wire _47910_;
wire _47911_;
wire _47912_;
wire _47913_;
wire _47914_;
wire _47915_;
wire _47916_;
wire _47917_;
wire _47918_;
wire _47919_;
wire _47920_;
wire _47921_;
wire _47922_;
wire _47923_;
wire _47924_;
wire _47925_;
wire _47926_;
wire _47927_;
wire _47928_;
wire _47929_;
wire _47930_;
wire _47931_;
wire _47932_;
wire _47933_;
wire _47934_;
wire _47935_;
wire _47936_;
wire _47937_;
wire _47938_;
wire _47939_;
wire _47940_;
wire _47941_;
wire _47942_;
wire _47943_;
wire _47944_;
wire _47945_;
wire _47946_;
wire _47947_;
wire _47948_;
wire _47949_;
wire _47950_;
wire _47951_;
wire _47952_;
wire _47953_;
wire _47954_;
wire _47955_;
wire _47956_;
wire _47957_;
wire _47958_;
wire _47959_;
wire _47960_;
wire _47961_;
wire _47962_;
wire _47963_;
wire _47964_;
wire _47965_;
wire _47966_;
wire _47967_;
wire _47968_;
wire _47969_;
wire _47970_;
wire _47971_;
wire _47972_;
wire _47973_;
wire _47974_;
wire _47975_;
wire _47976_;
wire _47977_;
wire _47978_;
wire _47979_;
wire _47980_;
wire _47981_;
wire _47982_;
wire _47983_;
wire _47984_;
wire _47985_;
wire _47986_;
wire _47987_;
wire _47988_;
wire _47989_;
wire _47990_;
wire _47991_;
wire _47992_;
wire _47993_;
wire _47994_;
wire _47995_;
wire _47996_;
wire _47997_;
wire _47998_;
wire _47999_;
wire _48000_;
wire _48001_;
wire _48002_;
wire _48003_;
wire _48004_;
wire _48005_;
wire _48006_;
wire _48007_;
wire _48008_;
wire _48009_;
wire _48010_;
wire _48011_;
wire _48012_;
wire _48013_;
wire _48014_;
wire _48015_;
wire _48016_;
wire _48017_;
wire _48018_;
wire _48019_;
wire _48020_;
wire _48021_;
wire _48022_;
wire _48023_;
wire _48024_;
wire _48025_;
wire _48026_;
wire _48027_;
wire _48028_;
wire _48029_;
wire _48030_;
wire _48031_;
wire _48032_;
wire _48033_;
wire _48034_;
wire _48035_;
wire _48036_;
wire _48037_;
wire _48038_;
wire _48039_;
wire _48040_;
wire _48041_;
wire _48042_;
wire _48043_;
wire _48044_;
wire _48045_;
wire _48046_;
wire _48047_;
wire _48048_;
wire _48049_;
wire _48050_;
wire _48051_;
wire _48052_;
wire _48053_;
wire _48054_;
wire _48055_;
wire _48056_;
wire _48057_;
wire _48058_;
wire _48059_;
wire _48060_;
wire _48061_;
wire _48062_;
wire _48063_;
wire _48064_;
wire _48065_;
wire _48066_;
wire _48067_;
wire _48068_;
wire _48069_;
wire _48070_;
wire _48071_;
wire _48072_;
wire _48073_;
wire _48074_;
wire _48075_;
wire _48076_;
wire _48077_;
wire _48078_;
wire _48079_;
wire _48080_;
wire _48081_;
wire _48082_;
wire _48083_;
wire _48084_;
wire _48085_;
wire _48086_;
wire _48087_;
wire _48088_;
wire _48089_;
wire _48090_;
wire _48091_;
wire _48092_;
wire _48093_;
wire _48094_;
wire _48095_;
wire _48096_;
wire _48097_;
wire _48098_;
wire _48099_;
wire _48100_;
wire _48101_;
wire _48102_;
wire _48103_;
wire _48104_;
wire _48105_;
wire _48106_;
wire _48107_;
wire _48108_;
wire _48109_;
wire _48110_;
wire _48111_;
wire _48112_;
wire _48113_;
wire _48114_;
wire _48115_;
wire _48116_;
wire _48117_;
wire _48118_;
wire _48119_;
wire _48120_;
wire _48121_;
wire _48122_;
wire _48123_;
wire _48124_;
wire _48125_;
wire _48126_;
wire _48127_;
wire _48128_;
wire _48129_;
wire _48130_;
wire _48131_;
wire _48132_;
wire _48133_;
wire _48134_;
wire _48135_;
wire _48136_;
wire _48137_;
wire _48138_;
wire _48139_;
wire _48140_;
wire _48141_;
wire _48142_;
wire _48143_;
wire _48144_;
wire _48145_;
wire _48146_;
wire _48147_;
wire _48148_;
wire _48149_;
wire _48150_;
wire _48151_;
wire _48152_;
wire _48153_;
wire _48154_;
wire _48155_;
wire _48156_;
wire _48157_;
wire _48158_;
wire _48159_;
wire _48160_;
wire _48161_;
wire _48162_;
wire _48163_;
wire _48164_;
wire _48165_;
wire _48166_;
wire _48167_;
wire _48168_;
wire _48169_;
wire _48170_;
wire _48171_;
wire _48172_;
wire _48173_;
wire _48174_;
wire _48175_;
wire _48176_;
wire _48177_;
wire _48178_;
wire _48179_;
wire _48180_;
wire _48181_;
wire _48182_;
wire _48183_;
wire _48184_;
wire _48185_;
wire _48186_;
wire _48187_;
wire _48188_;
wire _48189_;
wire _48190_;
wire _48191_;
wire _48192_;
wire _48193_;
wire _48194_;
wire _48195_;
wire _48196_;
wire _48197_;
wire _48198_;
wire _48199_;
wire _48200_;
wire _48201_;
wire _48202_;
wire _48203_;
wire _48204_;
wire _48205_;
wire _48206_;
wire _48207_;
wire _48208_;
wire _48209_;
wire _48210_;
wire _48211_;
wire _48212_;
wire _48213_;
wire _48214_;
wire _48215_;
wire _48216_;
wire _48217_;
wire _48218_;
wire _48219_;
wire _48220_;
wire _48221_;
wire _48222_;
wire _48223_;
wire _48224_;
wire _48225_;
wire _48226_;
wire _48227_;
wire _48228_;
wire _48229_;
wire _48230_;
wire _48231_;
wire _48232_;
wire _48233_;
wire _48234_;
wire _48235_;
wire _48236_;
wire _48237_;
wire _48238_;
wire _48239_;
wire _48240_;
wire _48241_;
wire _48242_;
wire _48243_;
wire _48244_;
wire _48245_;
wire _48246_;
wire _48247_;
wire _48248_;
wire _48249_;
wire _48250_;
wire _48251_;
wire _48252_;
wire _48253_;
wire _48254_;
wire _48255_;
wire _48256_;
wire _48257_;
wire _48258_;
wire _48259_;
wire _48260_;
wire _48261_;
wire _48262_;
wire _48263_;
wire _48264_;
wire _48265_;
wire _48266_;
wire _48267_;
wire _48268_;
wire _48269_;
wire _48270_;
wire _48271_;
wire _48272_;
wire _48273_;
wire _48274_;
wire _48275_;
wire _48276_;
wire _48277_;
wire _48278_;
wire _48279_;
wire _48280_;
wire _48281_;
wire _48282_;
wire _48283_;
wire _48284_;
wire _48285_;
wire _48286_;
wire _48287_;
wire _48288_;
wire _48289_;
wire _48290_;
wire _48291_;
wire _48292_;
wire _48293_;
wire _48294_;
wire _48295_;
wire _48296_;
wire _48297_;
wire _48298_;
wire _48299_;
wire _48300_;
wire _48301_;
wire _48302_;
wire _48303_;
wire _48304_;
wire _48305_;
wire _48306_;
wire _48307_;
wire _48308_;
wire _48309_;
wire _48310_;
wire _48311_;
wire _48312_;
wire _48313_;
wire _48314_;
wire _48315_;
wire _48316_;
wire _48317_;
wire _48318_;
wire _48319_;
wire _48320_;
wire _48321_;
wire _48322_;
wire _48323_;
wire _48324_;
wire _48325_;
wire _48326_;
wire _48327_;
wire _48328_;
wire _48329_;
wire _48330_;
wire _48331_;
wire _48332_;
wire _48333_;
wire _48334_;
wire _48335_;
wire _48336_;
wire _48337_;
wire _48338_;
wire _48339_;
wire _48340_;
wire _48341_;
wire _48342_;
wire _48343_;
wire _48344_;
wire _48345_;
wire _48346_;
wire _48347_;
wire _48348_;
wire _48349_;
wire _48350_;
wire _48351_;
wire _48352_;
wire _48353_;
wire _48354_;
wire _48355_;
wire _48356_;
wire _48357_;
wire _48358_;
wire _48359_;
wire _48360_;
wire _48361_;
wire _48362_;
wire _48363_;
wire _48364_;
wire _48365_;
wire _48366_;
wire _48367_;
wire _48368_;
wire _48369_;
wire _48370_;
wire _48371_;
wire _48372_;
wire _48373_;
wire _48374_;
wire _48375_;
wire _48376_;
wire _48377_;
wire _48378_;
wire _48379_;
wire _48380_;
wire _48381_;
wire _48382_;
wire _48383_;
wire _48384_;
wire _48385_;
wire _48386_;
wire _48387_;
wire _48388_;
wire _48389_;
wire _48390_;
wire _48391_;
wire _48392_;
wire _48393_;
wire _48394_;
wire _48395_;
wire _48396_;
wire _48397_;
wire _48398_;
wire _48399_;
wire _48400_;
wire _48401_;
wire _48402_;
wire _48403_;
wire _48404_;
wire _48405_;
wire _48406_;
wire _48407_;
wire _48408_;
wire _48409_;
wire _48410_;
wire _48411_;
wire _48412_;
wire _48413_;
wire _48414_;
wire _48415_;
wire _48416_;
wire _48417_;
wire _48418_;
wire _48419_;
wire _48420_;
wire _48421_;
wire _48422_;
wire _48423_;
wire _48424_;
wire _48425_;
wire _48426_;
wire _48427_;
wire _48428_;
wire _48429_;
wire _48430_;
wire _48431_;
wire _48432_;
wire _48433_;
wire _48434_;
wire _48435_;
wire _48436_;
wire _48437_;
wire _48438_;
wire _48439_;
wire _48440_;
wire _48441_;
wire _48442_;
wire _48443_;
wire _48444_;
wire _48445_;
wire _48446_;
wire _48447_;
wire _48448_;
wire _48449_;
wire _48450_;
wire _48451_;
wire _48452_;
wire _48453_;
wire _48454_;
wire _48455_;
wire _48456_;
wire _48457_;
wire _48458_;
wire _48459_;
wire _48460_;
wire _48461_;
wire _48462_;
wire _48463_;
wire _48464_;
wire _48465_;
wire _48466_;
wire _48467_;
wire _48468_;
wire _48469_;
wire _48470_;
wire _48471_;
wire _48472_;
wire _48473_;
wire _48474_;
wire _48475_;
wire _48476_;
wire _48477_;
wire _48478_;
wire _48479_;
wire _48480_;
wire _48481_;
wire _48482_;
wire _48483_;
wire _48484_;
wire _48485_;
wire _48486_;
wire _48487_;
wire _48488_;
wire _48489_;
wire _48490_;
wire _48491_;
wire _48492_;
wire _48493_;
wire _48494_;
wire _48495_;
wire _48496_;
wire _48497_;
wire _48498_;
wire _48499_;
wire _48500_;
wire _48501_;
wire _48502_;
wire _48503_;
wire _48504_;
wire _48505_;
wire _48506_;
wire _48507_;
wire _48508_;
wire _48509_;
wire _48510_;
wire _48511_;
wire _48512_;
wire _48513_;
wire _48514_;
wire _48515_;
wire _48516_;
wire _48517_;
wire _48518_;
wire _48519_;
wire _48520_;
wire _48521_;
wire _48522_;
wire _48523_;
wire _48524_;
wire _48525_;
wire _48526_;
wire _48527_;
wire _48528_;
wire _48529_;
wire _48530_;
wire _48531_;
wire _48532_;
wire _48533_;
wire _48534_;
wire _48535_;
wire _48536_;
wire _48537_;
wire _48538_;
wire _48539_;
wire _48540_;
wire _48541_;
wire _48542_;
wire _48543_;
wire _48544_;
wire _48545_;
wire _48546_;
wire _48547_;
wire _48548_;
wire _48549_;
wire _48550_;
wire _48551_;
wire _48552_;
wire _48553_;
wire _48554_;
wire _48555_;
wire _48556_;
wire _48557_;
wire _48558_;
wire _48559_;
wire _48560_;
wire _48561_;
wire _48562_;
wire _48563_;
wire _48564_;
wire _48565_;
wire _48566_;
wire _48567_;
wire _48568_;
wire _48569_;
wire _48570_;
wire _48571_;
wire _48572_;
wire _48573_;
wire _48574_;
wire _48575_;
wire _48576_;
wire _48577_;
wire _48578_;
wire _48579_;
wire _48580_;
wire _48581_;
wire _48582_;
wire _48583_;
wire _48584_;
wire _48585_;
wire _48586_;
wire _48587_;
wire _48588_;
wire _48589_;
wire _48590_;
wire _48591_;
wire _48592_;
wire _48593_;
wire _48594_;
wire _48595_;
wire _48596_;
wire _48597_;
wire _48598_;
wire _48599_;
wire _48600_;
wire _48601_;
wire _48602_;
wire _48603_;
wire _48604_;
wire _48605_;
wire _48606_;
wire _48607_;
wire _48608_;
wire _48609_;
wire _48610_;
wire _48611_;
wire _48612_;
wire _48613_;
wire _48614_;
wire _48615_;
wire _48616_;
wire _48617_;
wire _48618_;
wire _48619_;
wire _48620_;
wire _48621_;
wire _48622_;
wire _48623_;
wire _48624_;
wire _48625_;
wire _48626_;
wire _48627_;
wire _48628_;
wire _48629_;
wire _48630_;
wire _48631_;
wire _48632_;
wire _48633_;
wire _48634_;
wire _48635_;
wire _48636_;
wire _48637_;
wire _48638_;
wire _48639_;
wire _48640_;
wire _48641_;
wire _48642_;
wire _48643_;
wire _48644_;
wire _48645_;
wire _48646_;
wire _48647_;
wire _48648_;
wire _48649_;
wire _48650_;
wire _48651_;
wire _48652_;
wire _48653_;
wire _48654_;
wire _48655_;
wire _48656_;
wire _48657_;
wire _48658_;
wire _48659_;
wire _48660_;
wire _48661_;
wire _48662_;
wire _48663_;
wire _48664_;
wire _48665_;
wire _48666_;
wire _48667_;
wire _48668_;
wire _48669_;
wire _48670_;
wire _48671_;
wire _48672_;
wire _48673_;
wire _48674_;
wire _48675_;
wire _48676_;
wire _48677_;
wire _48678_;
wire _48679_;
wire _48680_;
wire _48681_;
wire _48682_;
wire _48683_;
wire _48684_;
wire _48685_;
wire _48686_;
wire _48687_;
wire _48688_;
wire _48689_;
wire _48690_;
wire _48691_;
wire _48692_;
wire _48693_;
wire _48694_;
wire _48695_;
wire _48696_;
wire _48697_;
wire _48698_;
wire _48699_;
wire _48700_;
wire _48701_;
wire _48702_;
wire _48703_;
wire _48704_;
wire _48705_;
wire _48706_;
wire _48707_;
wire _48708_;
wire _48709_;
wire _48710_;
wire _48711_;
wire _48712_;
wire _48713_;
wire _48714_;
wire _48715_;
wire _48716_;
wire _48717_;
wire _48718_;
wire _48719_;
wire _48720_;
wire _48721_;
wire _48722_;
wire _48723_;
wire _48724_;
wire _48725_;
wire _48726_;
wire _48727_;
wire _48728_;
wire _48729_;
wire _48730_;
wire _48731_;
wire _48732_;
wire _48733_;
wire _48734_;
wire _48735_;
wire _48736_;
wire _48737_;
wire _48738_;
wire _48739_;
wire _48740_;
wire _48741_;
wire _48742_;
wire _48743_;
wire _48744_;
wire _48745_;
wire _48746_;
wire _48747_;
wire _48748_;
wire _48749_;
wire _48750_;
wire _48751_;
wire _48752_;
wire _48753_;
wire _48754_;
wire _48755_;
wire _48756_;
wire _48757_;
wire _48758_;
wire _48759_;
wire _48760_;
wire _48761_;
wire _48762_;
wire _48763_;
wire _48764_;
wire _48765_;
wire _48766_;
wire _48767_;
wire _48768_;
wire _48769_;
wire _48770_;
wire _48771_;
wire _48772_;
wire _48773_;
wire _48774_;
wire _48775_;
wire _48776_;
wire _48777_;
wire _48778_;
wire _48779_;
wire _48780_;
wire _48781_;
wire _48782_;
wire _48783_;
wire _48784_;
wire _48785_;
wire _48786_;
wire _48787_;
wire _48788_;
wire _48789_;
wire _48790_;
wire _48791_;
wire _48792_;
wire _48793_;
wire _48794_;
wire _48795_;
wire _48796_;
wire _48797_;
wire _48798_;
wire _48799_;
wire _48800_;
wire _48801_;
wire _48802_;
wire _48803_;
wire _48804_;
wire _48805_;
wire _48806_;
wire _48807_;
wire _48808_;
wire _48809_;
wire _48810_;
wire _48811_;
wire _48812_;
wire _48813_;
wire _48814_;
wire _48815_;
wire _48816_;
wire _48817_;
wire _48818_;
wire _48819_;
wire _48820_;
wire _48821_;
wire _48822_;
wire _48823_;
wire _48824_;
wire _48825_;
wire _48826_;
wire _48827_;
wire _48828_;
wire _48829_;
wire _48830_;
wire _48831_;
wire _48832_;
wire _48833_;
wire _48834_;
wire _48835_;
wire _48836_;
wire _48837_;
wire _48838_;
wire _48839_;
wire _48840_;
wire _48841_;
wire _48842_;
wire _48843_;
wire _48844_;
wire _48845_;
wire _48846_;
wire _48847_;
wire _48848_;
wire _48849_;
wire _48850_;
wire _48851_;
wire _48852_;
wire _48853_;
wire _48854_;
wire _48855_;
wire _48856_;
wire _48857_;
wire _48858_;
wire _48859_;
wire _48860_;
wire _48861_;
wire _48862_;
wire _48863_;
wire _48864_;
wire _48865_;
wire _48866_;
wire _48867_;
wire _48868_;
wire _48869_;
wire _48870_;
wire _48871_;
wire _48872_;
wire _48873_;
wire _48874_;
wire _48875_;
wire _48876_;
wire _48877_;
wire _48878_;
wire _48879_;
wire _48880_;
wire _48881_;
wire _48882_;
wire _48883_;
wire _48884_;
wire _48885_;
wire _48886_;
wire _48887_;
wire _48888_;
wire _48889_;
wire _48890_;
wire _48891_;
wire _48892_;
wire _48893_;
wire _48894_;
wire _48895_;
wire _48896_;
wire _48897_;
wire _48898_;
wire _48899_;
wire _48900_;
wire _48901_;
wire _48902_;
wire _48903_;
wire _48904_;
wire _48905_;
wire _48906_;
wire _48907_;
wire _48908_;
wire _48909_;
wire _48910_;
wire _48911_;
wire _48912_;
wire _48913_;
wire _48914_;
wire _48915_;
wire _48916_;
wire _48917_;
wire _48918_;
wire _48919_;
wire _48920_;
wire _48921_;
wire _48922_;
wire _48923_;
wire _48924_;
wire _48925_;
wire _48926_;
wire _48927_;
wire _48928_;
wire _48929_;
wire _48930_;
wire _48931_;
wire _48932_;
wire _48933_;
wire _48934_;
wire _48935_;
wire _48936_;
wire _48937_;
wire _48938_;
wire _48939_;
wire _48940_;
wire _48941_;
wire _48942_;
wire _48943_;
wire _48944_;
wire _48945_;
wire _48946_;
wire _48947_;
wire _48948_;
wire _48949_;
wire _48950_;
wire _48951_;
wire _48952_;
wire _48953_;
wire _48954_;
wire _48955_;
wire _48956_;
wire _48957_;
wire _48958_;
wire _48959_;
wire _48960_;
wire _48961_;
wire _48962_;
wire _48963_;
wire _48964_;
wire _48965_;
wire _48966_;
wire _48967_;
wire _48968_;
wire _48969_;
wire _48970_;
wire _48971_;
wire _48972_;
wire _48973_;
wire _48974_;
wire _48975_;
wire _48976_;
wire _48977_;
wire _48978_;
wire _48979_;
wire _48980_;
wire _48981_;
wire _48982_;
wire _48983_;
wire _48984_;
wire _48985_;
wire _48986_;
wire _48987_;
wire _48988_;
wire _48989_;
wire _48990_;
wire _48991_;
wire _48992_;
wire _48993_;
wire _48994_;
wire _48995_;
wire _48996_;
wire _48997_;
wire _48998_;
wire _48999_;
wire _49000_;
wire _49001_;
wire _49002_;
wire _49003_;
wire _49004_;
wire _49005_;
wire _49006_;
wire _49007_;
wire _49008_;
wire _49009_;
wire _49010_;
wire _49011_;
wire _49012_;
wire _49013_;
wire _49014_;
wire _49015_;
wire _49016_;
wire _49017_;
wire _49018_;
wire _49019_;
wire _49020_;
wire _49021_;
wire _49022_;
wire _49023_;
wire _49024_;
wire _49025_;
wire _49026_;
wire _49027_;
wire _49028_;
wire _49029_;
wire _49030_;
wire _49031_;
wire _49032_;
wire _49033_;
wire _49034_;
wire _49035_;
wire _49036_;
wire _49037_;
wire _49038_;
wire _49039_;
wire _49040_;
wire _49041_;
wire _49042_;
wire _49043_;
wire _49044_;
wire _49045_;
wire _49046_;
wire _49047_;
wire _49048_;
wire _49049_;
wire _49050_;
wire _49051_;
wire _49052_;
wire _49053_;
wire _49054_;
wire _49055_;
wire _49056_;
wire _49057_;
wire _49058_;
wire _49059_;
wire _49060_;
wire _49061_;
wire _49062_;
wire _49063_;
wire _49064_;
wire _49065_;
wire _49066_;
wire _49067_;
wire _49068_;
wire _49069_;
wire _49070_;
wire _49071_;
wire _49072_;
wire _49073_;
wire _49074_;
wire _49075_;
wire _49076_;
wire _49077_;
wire _49078_;
wire _49079_;
wire _49080_;
wire _49081_;
wire _49082_;
wire _49083_;
wire _49084_;
wire _49085_;
wire _49086_;
wire _49087_;
wire _49088_;
wire _49089_;
wire _49090_;
wire _49091_;
wire _49092_;
wire _49093_;
wire _49094_;
wire _49095_;
wire _49096_;
wire _49097_;
wire _49098_;
wire _49099_;
wire _49100_;
wire _49101_;
wire _49102_;
wire _49103_;
wire _49104_;
wire _49105_;
wire _49106_;
wire _49107_;
wire _49108_;
wire _49109_;
wire _49110_;
wire _49111_;
wire _49112_;
wire _49113_;
wire _49114_;
wire _49115_;
wire _49116_;
wire _49117_;
wire _49118_;
wire _49119_;
wire _49120_;
wire _49121_;
wire _49122_;
wire _49123_;
wire _49124_;
wire _49125_;
wire _49126_;
wire _49127_;
wire _49128_;
wire _49129_;
wire _49130_;
wire _49131_;
wire _49132_;
wire _49133_;
wire _49134_;
wire _49135_;
wire _49136_;
wire _49137_;
wire _49138_;
wire _49139_;
wire _49140_;
wire _49141_;
wire _49142_;
wire _49143_;
wire _49144_;
wire _49145_;
wire _49146_;
wire _49147_;
wire _49148_;
wire _49149_;
wire _49150_;
wire _49151_;
wire _49152_;
wire _49153_;
wire _49154_;
wire _49155_;
wire _49156_;
wire _49157_;
wire _49158_;
wire _49159_;
wire _49160_;
wire _49161_;
wire _49162_;
wire _49163_;
wire _49164_;
wire _49165_;
wire _49166_;
wire _49167_;
wire _49168_;
wire _49169_;
wire _49170_;
wire _49171_;
wire _49172_;
wire _49173_;
wire _49174_;
wire _49175_;
wire _49176_;
wire _49177_;
wire _49178_;
wire _49179_;
wire _49180_;
wire _49181_;
wire _49182_;
wire _49183_;
wire _49184_;
wire _49185_;
wire _49186_;
wire _49187_;
wire _49188_;
wire _49189_;
wire _49190_;
wire _49191_;
wire _49192_;
wire _49193_;
wire _49194_;
wire _49195_;
wire _49196_;
wire _49197_;
wire _49198_;
wire _49199_;
wire _49200_;
wire _49201_;
wire _49202_;
wire _49203_;
wire _49204_;
wire _49205_;
wire _49206_;
wire _49207_;
wire _49208_;
wire _49209_;
wire _49210_;
wire _49211_;
wire _49212_;
wire _49213_;
wire _49214_;
wire _49215_;
wire _49216_;
wire _49217_;
wire _49218_;
wire _49219_;
wire _49220_;
wire _49221_;
wire _49222_;
wire _49223_;
wire _49224_;
wire _49225_;
wire _49226_;
wire _49227_;
wire _49228_;
wire _49229_;
wire _49230_;
wire _49231_;
wire _49232_;
wire _49233_;
wire _49234_;
wire _49235_;
wire _49236_;
wire _49237_;
wire _49238_;
wire _49239_;
wire _49240_;
wire _49241_;
wire _49242_;
wire _49243_;
wire _49244_;
wire _49245_;
wire _49246_;
wire _49247_;
wire _49248_;
wire _49249_;
wire _49250_;
wire _49251_;
wire _49252_;
wire _49253_;
wire _49254_;
wire _49255_;
wire _49256_;
wire _49257_;
wire _49258_;
wire _49259_;
wire _49260_;
wire _49261_;
wire _49262_;
wire _49263_;
wire _49264_;
wire _49265_;
wire _49266_;
wire _49267_;
wire _49268_;
wire _49269_;
wire _49270_;
wire _49271_;
wire _49272_;
wire _49273_;
wire _49274_;
wire _49275_;
wire _49276_;
wire _49277_;
wire _49278_;
wire _49279_;
wire _49280_;
wire _49281_;
wire _49282_;
wire _49283_;
wire _49284_;
wire _49285_;
wire _49286_;
wire _49287_;
wire _49288_;
wire _49289_;
wire _49290_;
wire _49291_;
wire _49292_;
wire _49293_;
wire _49294_;
wire _49295_;
wire _49296_;
wire _49297_;
wire _49298_;
wire _49299_;
wire _49300_;
wire _49301_;
wire _49302_;
wire _49303_;
wire _49304_;
wire _49305_;
wire _49306_;
wire _49307_;
wire _49308_;
wire _49309_;
wire _49310_;
wire _49311_;
wire _49312_;
wire _49313_;
wire _49314_;
wire _49315_;
wire _49316_;
wire _49317_;
wire _49318_;
wire _49319_;
wire _49320_;
wire _49321_;
wire _49322_;
wire _49323_;
wire _49324_;
wire _49325_;
wire _49326_;
wire _49327_;
wire _49328_;
wire _49329_;
wire _49330_;
wire _49331_;
wire _49332_;
wire _49333_;
wire _49334_;
wire _49335_;
wire _49336_;
wire _49337_;
wire _49338_;
wire _49339_;
wire _49340_;
wire _49341_;
wire _49342_;
wire _49343_;
wire _49344_;
wire _49345_;
wire _49346_;
wire _49347_;
wire _49348_;
wire _49349_;
wire _49350_;
wire _49351_;
wire _49352_;
wire _49353_;
wire _49354_;
wire _49355_;
wire _49356_;
wire _49357_;
wire _49358_;
wire _49359_;
wire _49360_;
wire _49361_;
wire _49362_;
wire _49363_;
wire _49364_;
wire _49365_;
wire _49366_;
wire _49367_;
wire _49368_;
wire _49369_;
wire _49370_;
wire _49371_;
wire _49372_;
wire _49373_;
wire _49374_;
wire _49375_;
wire _49376_;
wire _49377_;
wire _49378_;
wire _49379_;
wire _49380_;
wire _49381_;
wire _49382_;
wire _49383_;
wire _49384_;
wire _49385_;
wire _49386_;
wire _49387_;
wire _49388_;
wire _49389_;
wire _49390_;
wire _49391_;
wire _49392_;
wire _49393_;
wire _49394_;
wire _49395_;
wire _49396_;
wire _49397_;
wire _49398_;
wire _49399_;
wire _49400_;
wire _49401_;
wire _49402_;
wire _49403_;
wire _49404_;
wire _49405_;
wire _49406_;
wire _49407_;
wire _49408_;
wire _49409_;
wire _49410_;
wire _49411_;
wire _49412_;
wire _49413_;
wire _49414_;
wire _49415_;
wire _49416_;
wire _49417_;
wire _49418_;
wire _49419_;
wire _49420_;
wire _49421_;
wire _49422_;
wire _49423_;
wire _49424_;
wire _49425_;
wire _49426_;
wire _49427_;
wire _49428_;
wire _49429_;
wire _49430_;
wire _49431_;
wire _49432_;
wire _49433_;
wire _49434_;
wire _49435_;
wire _49436_;
wire _49437_;
wire _49438_;
wire _49439_;
wire _49440_;
wire _49441_;
wire _49442_;
wire _49443_;
wire _49444_;
wire _49445_;
wire _49446_;
wire _49447_;
wire _49448_;
wire _49449_;
wire _49450_;
wire _49451_;
wire _49452_;
wire _49453_;
wire _49454_;
wire _49455_;
wire _49456_;
wire _49457_;
wire _49458_;
wire _49459_;
wire _49460_;
wire _49461_;
wire _49462_;
wire _49463_;
wire _49464_;
wire _49465_;
wire _49466_;
wire _49467_;
wire _49468_;
wire _49469_;
wire _49470_;
wire _49471_;
wire _49472_;
wire _49473_;
wire _49474_;
wire _49475_;
wire _49476_;
wire _49477_;
wire _49478_;
wire _49479_;
wire _49480_;
wire _49481_;
wire _49482_;
wire _49483_;
wire _49484_;
wire _49485_;
wire _49486_;
wire _49487_;
wire _49488_;
wire _49489_;
wire _49490_;
wire _49491_;
wire _49492_;
wire _49493_;
wire _49494_;
wire _49495_;
wire _49496_;
wire _49497_;
wire _49498_;
wire _49499_;
wire _49500_;
wire _49501_;
wire _49502_;
wire _49503_;
wire _49504_;
wire _49505_;
wire _49506_;
wire _49507_;
wire _49508_;
wire _49509_;
wire _49510_;
wire _49511_;
wire _49512_;
wire _49513_;
wire _49514_;
wire _49515_;
wire _49516_;
wire _49517_;
wire _49518_;
wire _49519_;
wire _49520_;
wire _49521_;
wire _49522_;
wire _49523_;
wire _49524_;
wire _49525_;
wire _49526_;
wire _49527_;
wire _49528_;
wire _49529_;
wire _49530_;
wire _49531_;
wire _49532_;
wire _49533_;
wire _49534_;
wire _49535_;
wire _49536_;
wire _49537_;
wire _49538_;
wire _49539_;
wire _49540_;
wire _49541_;
wire _49542_;
wire _49543_;
wire _49544_;
wire _49545_;
wire _49546_;
wire _49547_;
wire _49548_;
wire _49549_;
wire _49550_;
wire _49551_;
wire _49552_;
wire _49553_;
wire _49554_;
wire _49555_;
wire _49556_;
wire _49557_;
wire _49558_;
wire _49559_;
wire _49560_;
wire _49561_;
wire _49562_;
wire _49563_;
wire _49564_;
wire _49565_;
wire _49566_;
wire _49567_;
wire _49568_;
wire _49569_;
wire _49570_;
wire _49571_;
wire _49572_;
wire _49573_;
wire _49574_;
wire _49575_;
wire _49576_;
wire _49577_;
wire _49578_;
wire _49579_;
wire _49580_;
wire _49581_;
wire _49582_;
wire _49583_;
wire _49584_;
wire _49585_;
wire _49586_;
wire _49587_;
wire _49588_;
wire _49589_;
wire _49590_;
wire _49591_;
wire _49592_;
wire _49593_;
wire _49594_;
wire _49595_;
wire _49596_;
wire _49597_;
wire _49598_;
wire _49599_;
wire _49600_;
wire _49601_;
wire _49602_;
wire _49603_;
wire _49604_;
wire _49605_;
wire _49606_;
wire _49607_;
wire _49608_;
wire _49609_;
wire _49610_;
wire _49611_;
wire _49612_;
wire _49613_;
wire _49614_;
wire _49615_;
wire _49616_;
wire _49617_;
wire _49618_;
wire _49619_;
wire _49620_;
wire _49621_;
wire _49622_;
wire _49623_;
wire _49624_;
wire _49625_;
wire _49626_;
wire _49627_;
wire _49628_;
wire _49629_;
wire _49630_;
wire _49631_;
wire _49632_;
wire _49633_;
wire _49634_;
wire _49635_;
wire _49636_;
wire _49637_;
wire _49638_;
wire _49639_;
wire _49640_;
wire _49641_;
wire _49642_;
wire _49643_;
wire _49644_;
wire _49645_;
wire _49646_;
wire _49647_;
wire _49648_;
wire _49649_;
wire _49650_;
wire _49651_;
wire _49652_;
wire _49653_;
wire _49654_;
wire _49655_;
wire _49656_;
wire _49657_;
wire _49658_;
wire _49659_;
wire _49660_;
wire _49661_;
wire _49662_;
wire _49663_;
wire _49664_;
wire _49665_;
wire _49666_;
wire _49667_;
wire _49668_;
wire _49669_;
wire _49670_;
wire _49671_;
wire _49672_;
wire _49673_;
wire _49674_;
wire _49675_;
wire _49676_;
wire _49677_;
wire _49678_;
wire _49679_;
wire _49680_;
wire _49681_;
wire _49682_;
wire _49683_;
wire _49684_;
wire _49685_;
wire _49686_;
wire _49687_;
wire _49688_;
wire _49689_;
wire _49690_;
wire _49691_;
wire _49692_;
wire _49693_;
wire _49694_;
wire _49695_;
wire _49696_;
wire _49697_;
wire _49698_;
wire _49699_;
wire _49700_;
wire _49701_;
wire _49702_;
wire _49703_;
wire _49704_;
wire _49705_;
wire _49706_;
wire _49707_;
wire _49708_;
wire _49709_;
wire _49710_;
wire _49711_;
wire _49712_;
wire _49713_;
wire _49714_;
wire _49715_;
wire _49716_;
wire _49717_;
wire _49718_;
wire _49719_;
wire _49720_;
wire _49721_;
wire _49722_;
wire _49723_;
wire _49724_;
wire _49725_;
wire _49726_;
wire _49727_;
wire _49728_;
wire _49729_;
wire _49730_;
wire _49731_;
wire _49732_;
wire _49733_;
wire _49734_;
wire _49735_;
wire _49736_;
wire _49737_;
wire _49738_;
wire _49739_;
wire _49740_;
wire _49741_;
wire _49742_;
wire _49743_;
wire _49744_;
wire _49745_;
wire _49746_;
wire _49747_;
wire _49748_;
wire _49749_;
wire _49750_;
wire _49751_;
wire _49752_;
wire _49753_;
wire _49754_;
wire _49755_;
wire _49756_;
wire _49757_;
wire _49758_;
wire _49759_;
wire _49760_;
wire _49761_;
wire _49762_;
wire _49763_;
wire _49764_;
wire _49765_;
wire _49766_;
wire _49767_;
wire _49768_;
wire _49769_;
wire _49770_;
wire _49771_;
wire _49772_;
wire _49773_;
wire _49774_;
wire _49775_;
wire _49776_;
wire _49777_;
wire _49778_;
wire _49779_;
wire _49780_;
wire _49781_;
wire _49782_;
wire _49783_;
wire _49784_;
wire _49785_;
wire _49786_;
wire _49787_;
wire _49788_;
wire _49789_;
wire _49790_;
wire _49791_;
wire _49792_;
wire _49793_;
wire _49794_;
wire _49795_;
wire _49796_;
wire _49797_;
wire _49798_;
wire _49799_;
wire _49800_;
wire _49801_;
wire _49802_;
wire _49803_;
wire _49804_;
wire _49805_;
wire _49806_;
wire _49807_;
wire _49808_;
wire _49809_;
wire _49810_;
wire _49811_;
wire _49812_;
wire _49813_;
wire _49814_;
wire _49815_;
wire _49816_;
wire _49817_;
wire _49818_;
wire _49819_;
wire _49820_;
wire _49821_;
wire _49822_;
wire _49823_;
wire _49824_;
wire _49825_;
wire _49826_;
wire _49827_;
wire _49828_;
wire _49829_;
wire _49830_;
wire _49831_;
wire _49832_;
wire _49833_;
wire _49834_;
wire _49835_;
wire _49836_;
wire _49837_;
wire _49838_;
wire _49839_;
wire _49840_;
wire _49841_;
wire _49842_;
wire _49843_;
wire _49844_;
wire _49845_;
wire _49846_;
wire _49847_;
wire _49848_;
wire _49849_;
wire _49850_;
wire _49851_;
wire _49852_;
wire _49853_;
wire _49854_;
wire _49855_;
wire _49856_;
wire _49857_;
wire _49858_;
wire _49859_;
wire _49860_;
wire _49861_;
wire _49862_;
wire _49863_;
wire _49864_;
wire _49865_;
wire _49866_;
wire _49867_;
wire _49868_;
wire _49869_;
wire _49870_;
wire _49871_;
wire _49872_;
wire _49873_;
wire _49874_;
wire _49875_;
wire _49876_;
wire _49877_;
wire _49878_;
wire _49879_;
wire _49880_;
wire _49881_;
wire _49882_;
wire _49883_;
wire _49884_;
wire _49885_;
wire _49886_;
wire _49887_;
wire _49888_;
wire _49889_;
wire _49890_;
wire _49891_;
wire _49892_;
wire _49893_;
wire _49894_;
wire _49895_;
wire _49896_;
wire _49897_;
wire _49898_;
wire _49899_;
wire _49900_;
wire _49901_;
wire _49902_;
wire _49903_;
wire _49904_;
wire _49905_;
wire _49906_;
wire _49907_;
wire _49908_;
wire _49909_;
wire _49910_;
wire _49911_;
wire _49912_;
wire _49913_;
wire _49914_;
wire _49915_;
wire _49916_;
wire _49917_;
wire _49918_;
wire _49919_;
wire _49920_;
wire _49921_;
wire _49922_;
wire _49923_;
wire _49924_;
wire _49925_;
wire _49926_;
wire _49927_;
wire _49928_;
wire _49929_;
wire _49930_;
wire _49931_;
wire _49932_;
wire _49933_;
wire _49934_;
wire _49935_;
wire _49936_;
wire _49937_;
wire _49938_;
wire _49939_;
wire _49940_;
wire _49941_;
wire _49942_;
wire _49943_;
wire _49944_;
wire _49945_;
wire _49946_;
wire _49947_;
wire _49948_;
wire _49949_;
wire _49950_;
wire _49951_;
wire _49952_;
wire _49953_;
wire _49954_;
wire _49955_;
wire _49956_;
wire _49957_;
wire _49958_;
wire _49959_;
wire _49960_;
wire _49961_;
wire _49962_;
wire _49963_;
wire _49964_;
wire _49965_;
wire _49966_;
wire _49967_;
wire _49968_;
wire _49969_;
wire _49970_;
wire _49971_;
wire _49972_;
wire _49973_;
wire _49974_;
wire _49975_;
wire _49976_;
wire _49977_;
wire _49978_;
wire _49979_;
wire _49980_;
wire _49981_;
wire _49982_;
wire _49983_;
wire _49984_;
wire _49985_;
wire _49986_;
wire _49987_;
wire _49988_;
wire _49989_;
wire _49990_;
wire _49991_;
wire _49992_;
wire _49993_;
wire _49994_;
wire _49995_;
wire _49996_;
wire _49997_;
wire _49998_;
wire _49999_;
wire _50000_;
wire _50001_;
wire _50002_;
wire _50003_;
wire _50004_;
wire _50005_;
wire _50006_;
wire _50007_;
wire _50008_;
wire _50009_;
wire _50010_;
wire _50011_;
wire _50012_;
wire _50013_;
wire _50014_;
wire _50015_;
wire _50016_;
wire _50017_;
wire _50018_;
wire _50019_;
wire _50020_;
wire _50021_;
wire _50022_;
wire _50023_;
wire _50024_;
wire _50025_;
wire _50026_;
wire _50027_;
wire _50028_;
wire _50029_;
wire _50030_;
wire _50031_;
wire _50032_;
wire _50033_;
wire _50034_;
wire _50035_;
wire _50036_;
wire _50037_;
wire _50038_;
wire _50039_;
wire _50040_;
wire _50041_;
wire _50042_;
wire _50043_;
wire _50044_;
wire _50045_;
wire _50046_;
wire _50047_;
wire _50048_;
wire _50049_;
wire _50050_;
wire _50051_;
wire _50052_;
wire _50053_;
wire _50054_;
wire _50055_;
wire _50056_;
wire _50057_;
wire _50058_;
wire _50059_;
wire _50060_;
wire _50061_;
wire _50062_;
wire _50063_;
wire _50064_;
wire _50065_;
wire _50066_;
wire _50067_;
wire _50068_;
wire _50069_;
wire _50070_;
wire _50071_;
wire _50072_;
wire _50073_;
wire _50074_;
wire _50075_;
wire _50076_;
wire _50077_;
wire _50078_;
wire _50079_;
wire _50080_;
wire _50081_;
wire _50082_;
wire _50083_;
wire _50084_;
wire _50085_;
wire _50086_;
wire _50087_;
wire _50088_;
wire _50089_;
wire _50090_;
wire _50091_;
wire _50092_;
wire _50093_;
wire _50094_;
wire _50095_;
wire _50096_;
wire _50097_;
wire _50098_;
wire _50099_;
wire _50100_;
wire _50101_;
wire _50102_;
wire _50103_;
wire _50104_;
wire _50105_;
wire _50106_;
wire _50107_;
wire _50108_;
wire _50109_;
wire _50110_;
wire _50111_;
wire _50112_;
wire _50113_;
wire _50114_;
wire _50115_;
wire _50116_;
wire _50117_;
wire _50118_;
wire _50119_;
wire _50120_;
wire _50121_;
wire _50122_;
wire _50123_;
wire _50124_;
wire _50125_;
wire _50126_;
wire _50127_;
wire _50128_;
wire _50129_;
wire _50130_;
wire _50131_;
wire _50132_;
wire _50133_;
wire _50134_;
wire _50135_;
wire _50136_;
wire _50137_;
wire _50138_;
wire _50139_;
wire _50140_;
wire _50141_;
wire _50142_;
wire _50143_;
wire _50144_;
wire _50145_;
wire _50146_;
wire _50147_;
wire _50148_;
wire _50149_;
wire _50150_;
wire _50151_;
wire _50152_;
wire _50153_;
wire _50154_;
wire _50155_;
wire _50156_;
wire _50157_;
wire _50158_;
wire _50159_;
wire _50160_;
wire _50161_;
wire _50162_;
wire _50163_;
wire _50164_;
wire _50165_;
wire _50166_;
wire _50167_;
wire _50168_;
wire _50169_;
wire _50170_;
wire _50171_;
wire _50172_;
wire _50173_;
wire _50174_;
wire _50175_;
wire _50176_;
wire _50177_;
wire _50178_;
wire _50179_;
wire _50180_;
wire _50181_;
wire _50182_;
wire _50183_;
wire _50184_;
wire _50185_;
wire _50186_;
wire _50187_;
wire _50188_;
wire _50189_;
wire _50190_;
wire _50191_;
wire _50192_;
wire _50193_;
wire _50194_;
wire _50195_;
wire _50196_;
wire _50197_;
wire _50198_;
wire _50199_;
wire _50200_;
wire _50201_;
wire _50202_;
wire _50203_;
wire _50204_;
wire _50205_;
wire _50206_;
wire _50207_;
wire _50208_;
wire _50209_;
wire _50210_;
wire _50211_;
wire _50212_;
wire _50213_;
wire _50214_;
wire _50215_;
wire _50216_;
wire _50217_;
wire _50218_;
wire _50219_;
wire _50220_;
wire _50221_;
wire _50222_;
wire _50223_;
wire _50224_;
wire _50225_;
wire _50226_;
wire _50227_;
wire _50228_;
wire _50229_;
wire _50230_;
wire _50231_;
wire _50232_;
wire _50233_;
wire _50234_;
wire _50235_;
wire _50236_;
wire _50237_;
wire _50238_;
wire _50239_;
wire _50240_;
wire _50241_;
wire _50242_;
wire _50243_;
wire _50244_;
wire _50245_;
wire _50246_;
wire _50247_;
wire _50248_;
wire _50249_;
wire _50250_;
wire _50251_;
wire _50252_;
wire _50253_;
wire _50254_;
wire _50255_;
wire _50256_;
wire _50257_;
wire _50258_;
wire _50259_;
wire _50260_;
wire _50261_;
wire _50262_;
wire _50263_;
wire _50264_;
wire _50265_;
wire _50266_;
wire _50267_;
wire _50268_;
wire _50269_;
wire _50270_;
wire _50271_;
wire _50272_;
wire _50273_;
wire _50274_;
wire _50275_;
wire _50276_;
wire _50277_;
wire _50278_;
wire _50279_;
wire _50280_;
wire _50281_;
wire _50282_;
wire _50283_;
wire _50284_;
wire _50285_;
wire _50286_;
wire _50287_;
wire _50288_;
wire _50289_;
wire _50290_;
wire _50291_;
wire _50292_;
wire _50293_;
wire _50294_;
wire _50295_;
wire _50296_;
wire _50297_;
wire _50298_;
wire _50299_;
wire _50300_;
wire _50301_;
wire _50302_;
wire _50303_;
wire _50304_;
wire _50305_;
wire _50306_;
wire _50307_;
wire _50308_;
wire _50309_;
wire _50310_;
wire _50311_;
wire _50312_;
wire _50313_;
wire _50314_;
wire _50315_;
wire _50316_;
wire _50317_;
wire _50318_;
wire _50319_;
wire _50320_;
wire _50321_;
wire _50322_;
wire _50323_;
wire _50324_;
wire _50325_;
wire _50326_;
wire _50327_;
wire _50328_;
wire _50329_;
wire _50330_;
wire _50331_;
wire _50332_;
wire _50333_;
wire _50334_;
wire _50335_;
wire _50336_;
wire _50337_;
wire _50338_;
wire _50339_;
wire _50340_;
wire _50341_;
wire _50342_;
wire _50343_;
wire _50344_;
wire _50345_;
wire _50346_;
wire _50347_;
wire _50348_;
wire _50349_;
wire _50350_;
wire _50351_;
wire _50352_;
wire _50353_;
wire _50354_;
wire _50355_;
wire _50356_;
wire _50357_;
wire _50358_;
wire _50359_;
wire _50360_;
wire _50361_;
wire _50362_;
wire _50363_;
wire _50364_;
wire _50365_;
wire _50366_;
wire _50367_;
wire _50368_;
wire _50369_;
wire _50370_;
wire _50371_;
wire _50372_;
wire _50373_;
wire _50374_;
wire _50375_;
wire _50376_;
wire _50377_;
wire _50378_;
wire _50379_;
wire _50380_;
wire _50381_;
wire _50382_;
wire _50383_;
wire _50384_;
wire _50385_;
wire _50386_;
wire _50387_;
wire _50388_;
wire _50389_;
wire _50390_;
wire _50391_;
wire _50392_;
wire _50393_;
wire _50394_;
wire _50395_;
wire _50396_;
wire _50397_;
wire _50398_;
wire _50399_;
wire _50400_;
wire _50401_;
wire _50402_;
wire _50403_;
wire _50404_;
wire _50405_;
wire _50406_;
wire _50407_;
wire _50408_;
wire _50409_;
wire _50410_;
wire _50411_;
wire _50412_;
wire _50413_;
wire _50414_;
wire _50415_;
wire _50416_;
wire _50417_;
wire _50418_;
wire _50419_;
wire _50420_;
wire _50421_;
wire _50422_;
wire _50423_;
wire _50424_;
wire _50425_;
wire _50426_;
wire _50427_;
wire _50428_;
wire _50429_;
wire _50430_;
wire _50431_;
wire _50432_;
wire _50433_;
wire _50434_;
wire _50435_;
wire _50436_;
wire _50437_;
wire _50438_;
wire _50439_;
wire _50440_;
wire _50441_;
wire _50442_;
wire _50443_;
wire _50444_;
wire _50445_;
wire _50446_;
wire _50447_;
wire _50448_;
wire _50449_;
wire _50450_;
wire _50451_;
wire _50452_;
wire _50453_;
wire _50454_;
wire _50455_;
wire _50456_;
wire _50457_;
wire _50458_;
wire _50459_;
wire _50460_;
wire _50461_;
wire _50462_;
wire _50463_;
wire _50464_;
wire _50465_;
wire _50466_;
wire _50467_;
wire _50468_;
wire _50469_;
wire _50470_;
wire _50471_;
wire _50472_;
wire _50473_;
wire _50474_;
wire _50475_;
wire _50476_;
wire _50477_;
wire _50478_;
wire _50479_;
wire _50480_;
wire _50481_;
wire _50482_;
wire _50483_;
wire _50484_;
wire _50485_;
wire _50486_;
wire _50487_;
wire _50488_;
wire _50489_;
wire _50490_;
wire _50491_;
wire _50492_;
wire _50493_;
wire _50494_;
wire _50495_;
wire _50496_;
wire _50497_;
wire _50498_;
wire _50499_;
wire _50500_;
wire _50501_;
wire _50502_;
wire _50503_;
wire _50504_;
wire _50505_;
wire _50506_;
wire _50507_;
wire _50508_;
wire _50509_;
wire _50510_;
wire _50511_;
wire _50512_;
wire _50513_;
wire _50514_;
wire _50515_;
wire _50516_;
wire _50517_;
wire _50518_;
wire _50519_;
wire _50520_;
wire _50521_;
wire _50522_;
wire _50523_;
wire _50524_;
wire _50525_;
wire _50526_;
wire _50527_;
wire _50528_;
wire _50529_;
wire _50530_;
wire _50531_;
wire _50532_;
wire _50533_;
wire _50534_;
wire _50535_;
wire _50536_;
wire _50537_;
wire _50538_;
wire _50539_;
wire _50540_;
wire _50541_;
wire _50542_;
wire _50543_;
wire _50544_;
wire _50545_;
wire _50546_;
wire _50547_;
wire _50548_;
wire _50549_;
wire _50550_;
wire _50551_;
wire _50552_;
wire _50553_;
wire _50554_;
wire _50555_;
wire _50556_;
wire _50557_;
wire _50558_;
wire _50559_;
wire _50560_;
wire _50561_;
wire _50562_;
wire _50563_;
wire _50564_;
wire _50565_;
wire _50566_;
wire _50567_;
wire _50568_;
wire _50569_;
wire _50570_;
wire _50571_;
wire _50572_;
wire _50573_;
wire _50574_;
wire _50575_;
wire _50576_;
wire _50577_;
wire _50578_;
wire _50579_;
wire _50580_;
wire _50581_;
wire _50582_;
wire _50583_;
wire _50584_;
wire _50585_;
wire _50586_;
wire _50587_;
wire _50588_;
wire _50589_;
wire _50590_;
wire _50591_;
wire _50592_;
wire _50593_;
wire _50594_;
wire _50595_;
wire _50596_;
wire _50597_;
wire _50598_;
wire _50599_;
wire _50600_;
wire _50601_;
wire _50602_;
wire _50603_;
wire _50604_;
wire _50605_;
wire _50606_;
wire _50607_;
wire _50608_;
wire _50609_;
wire _50610_;
wire _50611_;
wire _50612_;
wire _50613_;
wire _50614_;
wire _50615_;
wire _50616_;
wire _50617_;
wire _50618_;
wire _50619_;
wire _50620_;
wire _50621_;
wire _50622_;
wire _50623_;
wire _50624_;
wire _50625_;
wire _50626_;
wire _50627_;
wire _50628_;
wire _50629_;
wire _50630_;
wire _50631_;
wire _50632_;
wire _50633_;
wire _50634_;
wire _50635_;
wire _50636_;
wire _50637_;
wire _50638_;
wire _50639_;
wire _50640_;
wire _50641_;
wire _50642_;
wire _50643_;
wire _50644_;
wire _50645_;
wire _50646_;
wire _50647_;
wire _50648_;
wire _50649_;
wire _50650_;
wire _50651_;
wire _50652_;
wire _50653_;
wire _50654_;
wire _50655_;
wire _50656_;
wire _50657_;
wire _50658_;
wire _50659_;
wire _50660_;
wire _50661_;
wire _50662_;
wire _50663_;
wire _50664_;
wire _50665_;
wire _50666_;
wire _50667_;
wire _50668_;
wire _50669_;
wire _50670_;
wire _50671_;
wire _50672_;
wire _50673_;
wire _50674_;
wire _50675_;
wire _50676_;
wire _50677_;
wire _50678_;
wire _50679_;
wire _50680_;
wire _50681_;
wire _50682_;
wire _50683_;
wire _50684_;
wire _50685_;
wire _50686_;
wire _50687_;
wire _50688_;
wire _50689_;
wire _50690_;
wire _50691_;
wire _50692_;
wire _50693_;
wire _50694_;
wire _50695_;
wire _50696_;
wire _50697_;
wire _50698_;
wire _50699_;
wire _50700_;
wire _50701_;
wire _50702_;
wire _50703_;
wire _50704_;
wire _50705_;
wire _50706_;
wire _50707_;
wire _50708_;
wire _50709_;
wire _50710_;
wire _50711_;
wire _50712_;
wire _50713_;
wire _50714_;
wire _50715_;
wire _50716_;
wire _50717_;
wire _50718_;
wire _50719_;
wire _50720_;
wire _50721_;
wire _50722_;
wire _50723_;
wire _50724_;
wire _50725_;
wire _50726_;
wire _50727_;
wire _50728_;
wire _50729_;
wire _50730_;
wire _50731_;
wire _50732_;
wire _50733_;
wire _50734_;
wire _50735_;
wire _50736_;
wire _50737_;
wire _50738_;
wire _50739_;
wire _50740_;
wire _50741_;
wire _50742_;
wire _50743_;
wire _50744_;
wire _50745_;
wire _50746_;
wire _50747_;
wire _50748_;
wire _50749_;
wire _50750_;
wire _50751_;
wire _50752_;
wire _50753_;
wire _50754_;
wire _50755_;
wire _50756_;
wire _50757_;
wire _50758_;
wire _50759_;
wire _50760_;
wire _50761_;
wire _50762_;
wire _50763_;
wire _50764_;
wire _50765_;
wire _50766_;
wire _50767_;
wire _50768_;
wire _50769_;
wire _50770_;
wire _50771_;
wire _50772_;
wire _50773_;
wire _50774_;
wire _50775_;
wire _50776_;
wire _50777_;
wire _50778_;
wire _50779_;
wire _50780_;
wire _50781_;
wire _50782_;
wire _50783_;
wire _50784_;
wire _50785_;
wire _50786_;
wire _50787_;
wire _50788_;
wire _50789_;
wire _50790_;
wire _50791_;
wire _50792_;
wire _50793_;
wire _50794_;
wire _50795_;
wire _50796_;
wire _50797_;
wire _50798_;
wire _50799_;
wire _50800_;
wire _50801_;
wire _50802_;
wire _50803_;
wire _50804_;
wire _50805_;
wire _50806_;
wire _50807_;
wire _50808_;
wire _50809_;
wire _50810_;
wire _50811_;
wire _50812_;
wire _50813_;
wire _50814_;
wire _50815_;
wire _50816_;
wire _50817_;
wire _50818_;
wire _50819_;
wire _50820_;
wire _50821_;
wire _50822_;
wire _50823_;
wire _50824_;
wire _50825_;
wire _50826_;
wire _50827_;
wire _50828_;
wire _50829_;
wire _50830_;
wire _50831_;
wire _50832_;
wire _50833_;
wire _50834_;
wire _50835_;
wire _50836_;
wire _50837_;
wire _50838_;
wire _50839_;
wire _50840_;
wire _50841_;
wire _50842_;
wire _50843_;
wire _50844_;
wire _50845_;
wire _50846_;
wire _50847_;
wire _50848_;
wire _50849_;
wire _50850_;
wire _50851_;
wire _50852_;
wire _50853_;
wire _50854_;
wire _50855_;
wire _50856_;
wire _50857_;
wire _50858_;
wire _50859_;
wire _50860_;
wire _50861_;
wire _50862_;
wire _50863_;
wire _50864_;
wire _50865_;
wire _50866_;
wire _50867_;
wire _50868_;
wire _50869_;
wire _50870_;
wire _50871_;
wire _50872_;
wire _50873_;
wire _50874_;
wire _50875_;
wire _50876_;
wire _50877_;
wire _50878_;
wire _50879_;
wire _50880_;
wire _50881_;
wire _50882_;
wire _50883_;
wire _50884_;
wire _50885_;
wire _50886_;
wire _50887_;
wire _50888_;
wire _50889_;
wire _50890_;
wire _50891_;
wire _50892_;
wire _50893_;
wire _50894_;
wire _50895_;
wire _50896_;
wire _50897_;
wire _50898_;
wire _50899_;
wire _50900_;
wire _50901_;
wire _50902_;
wire _50903_;
wire _50904_;
wire _50905_;
wire _50906_;
wire _50907_;
wire _50908_;
wire _50909_;
wire _50910_;
wire _50911_;
wire _50912_;
wire _50913_;
wire _50914_;
wire _50915_;
wire _50916_;
wire _50917_;
wire _50918_;
wire _50919_;
wire _50920_;
wire _50921_;
wire _50922_;
wire _50923_;
wire _50924_;
wire _50925_;
wire _50926_;
wire _50927_;
wire _50928_;
wire _50929_;
wire _50930_;
wire _50931_;
wire _50932_;
wire _50933_;
wire _50934_;
wire _50935_;
wire _50936_;
wire _50937_;
wire _50938_;
wire _50939_;
wire _50940_;
wire _50941_;
wire _50942_;
wire _50943_;
wire _50944_;
wire _50945_;
wire _50946_;
wire _50947_;
wire _50948_;
wire _50949_;
wire _50950_;
wire _50951_;
wire _50952_;
wire _50953_;
wire _50954_;
wire _50955_;
wire _50956_;
wire _50957_;
wire _50958_;
wire _50959_;
wire _50960_;
wire _50961_;
wire _50962_;
wire _50963_;
wire _50964_;
wire _50965_;
wire _50966_;
wire _50967_;
wire _50968_;
wire _50969_;
wire _50970_;
wire _50971_;
wire _50972_;
wire _50973_;
wire _50974_;
wire _50975_;
wire _50976_;
wire _50977_;
wire _50978_;
wire _50979_;
wire _50980_;
wire _50981_;
wire _50982_;
wire _50983_;
wire _50984_;
wire _50985_;
wire _50986_;
wire _50987_;
wire _50988_;
wire _50989_;
wire _50990_;
wire _50991_;
wire _50992_;
wire _50993_;
wire _50994_;
wire _50995_;
wire _50996_;
wire _50997_;
wire _50998_;
wire _50999_;
wire _51000_;
wire _51001_;
wire _51002_;
wire _51003_;
wire _51004_;
wire _51005_;
wire _51006_;
wire _51007_;
wire _51008_;
wire _51009_;
wire _51010_;
wire _51011_;
wire _51012_;
wire _51013_;
wire _51014_;
wire _51015_;
wire _51016_;
wire _51017_;
wire _51018_;
wire _51019_;
wire _51020_;
wire _51021_;
wire _51022_;
wire _51023_;
wire _51024_;
wire _51025_;
wire _51026_;
wire _51027_;
wire _51028_;
wire _51029_;
wire _51030_;
wire _51031_;
wire _51032_;
wire _51033_;
wire _51034_;
wire _51035_;
wire _51036_;
wire _51037_;
wire _51038_;
wire _51039_;
wire _51040_;
wire _51041_;
wire _51042_;
wire _51043_;
wire _51044_;
wire _51045_;
wire _51046_;
wire _51047_;
wire _51048_;
wire _51049_;
wire _51050_;
wire _51051_;
wire _51052_;
wire _51053_;
wire _51054_;
wire _51055_;
wire _51056_;
wire _51057_;
wire _51058_;
wire _51059_;
wire _51060_;
wire _51061_;
wire _51062_;
wire _51063_;
wire _51064_;
wire _51065_;
wire _51066_;
wire _51067_;
wire _51068_;
wire _51069_;
wire _51070_;
wire _51071_;
wire _51072_;
wire _51073_;
wire _51074_;
wire _51075_;
wire _51076_;
wire _51077_;
wire _51078_;
wire _51079_;
wire _51080_;
wire _51081_;
wire _51082_;
wire _51083_;
wire _51084_;
wire _51085_;
wire _51086_;
wire _51087_;
wire _51088_;
wire _51089_;
wire _51090_;
wire _51091_;
wire _51092_;
wire _51093_;
wire _51094_;
wire _51095_;
wire _51096_;
wire _51097_;
wire _51098_;
wire _51099_;
wire _51100_;
wire _51101_;
wire _51102_;
wire _51103_;
wire _51104_;
wire _51105_;
wire _51106_;
wire _51107_;
wire _51108_;
wire _51109_;
wire _51110_;
wire _51111_;
wire _51112_;
wire _51113_;
wire _51114_;
wire _51115_;
wire _51116_;
wire _51117_;
wire _51118_;
wire _51119_;
wire _51120_;
wire _51121_;
wire _51122_;
wire _51123_;
wire _51124_;
wire _51125_;
wire _51126_;
wire _51127_;
wire _51128_;
wire _51129_;
wire _51130_;
wire _51131_;
wire _51132_;
wire _51133_;
wire _51134_;
wire _51135_;
wire _51136_;
wire _51137_;
wire _51138_;
wire _51139_;
wire _51140_;
wire _51141_;
wire _51142_;
wire _51143_;
wire _51144_;
wire _51145_;
wire _51146_;
wire _51147_;
wire _51148_;
wire _51149_;
wire _51150_;
wire _51151_;
wire _51152_;
wire _51153_;
wire _51154_;
wire _51155_;
wire _51156_;
wire _51157_;
wire _51158_;
wire _51159_;
wire _51160_;
wire _51161_;
wire _51162_;
wire _51163_;
wire _51164_;
wire _51165_;
wire _51166_;
wire _51167_;
wire _51168_;
wire _51169_;
wire _51170_;
wire _51171_;
wire _51172_;
wire _51173_;
wire _51174_;
wire _51175_;
wire _51176_;
wire _51177_;
wire _51178_;
wire _51179_;
wire _51180_;
wire _51181_;
wire _51182_;
wire _51183_;
wire _51184_;
wire _51185_;
wire _51186_;
wire _51187_;
wire _51188_;
wire _51189_;
wire _51190_;
wire _51191_;
wire _51192_;
wire _51193_;
wire _51194_;
wire _51195_;
wire _51196_;
wire _51197_;
wire _51198_;
wire _51199_;
wire _51200_;
wire _51201_;
wire _51202_;
wire _51203_;
wire _51204_;
wire _51205_;
wire _51206_;
wire _51207_;
wire _51208_;
wire _51209_;
wire _51210_;
wire _51211_;
wire _51212_;
wire _51213_;
wire _51214_;
wire _51215_;
wire _51216_;
wire _51217_;
wire _51218_;
wire _51219_;
wire _51220_;
wire _51221_;
wire _51222_;
wire _51223_;
wire _51224_;
wire _51225_;
wire _51226_;
wire _51227_;
wire _51228_;
wire _51229_;
wire _51230_;
wire _51231_;
wire _51232_;
wire _51233_;
wire _51234_;
wire _51235_;
wire _51236_;
wire _51237_;
wire _51238_;
wire _51239_;
wire _51240_;
wire _51241_;
wire _51242_;
wire _51243_;
wire _51244_;
wire _51245_;
wire _51246_;
wire _51247_;
wire _51248_;
wire _51249_;
wire _51250_;
wire _51251_;
wire _51252_;
wire _51253_;
wire _51254_;
wire _51255_;
wire _51256_;
wire _51257_;
wire _51258_;
wire _51259_;
wire _51260_;
wire _51261_;
wire _51262_;
wire _51263_;
wire _51264_;
wire _51265_;
wire _51266_;
wire _51267_;
wire _51268_;
wire _51269_;
wire _51270_;
wire _51271_;
wire _51272_;
wire _51273_;
wire _51274_;
wire _51275_;
wire _51276_;
wire _51277_;
wire _51278_;
wire _51279_;
wire _51280_;
wire _51281_;
wire _51282_;
wire _51283_;
wire _51284_;
wire _51285_;
wire _51286_;
wire _51287_;
wire _51288_;
wire _51289_;
wire _51290_;
wire _51291_;
wire _51292_;
wire _51293_;
wire _51294_;
wire _51295_;
wire _51296_;
wire _51297_;
wire _51298_;
wire _51299_;
wire _51300_;
wire _51301_;
wire _51302_;
wire _51303_;
wire _51304_;
wire _51305_;
wire _51306_;
wire _51307_;
wire _51308_;
wire _51309_;
wire _51310_;
wire _51311_;
wire _51312_;
wire _51313_;
wire _51314_;
wire _51315_;
wire _51316_;
wire _51317_;
wire _51318_;
wire _51319_;
wire _51320_;
wire _51321_;
wire _51322_;
wire _51323_;
wire _51324_;
wire _51325_;
wire _51326_;
wire _51327_;
wire _51328_;
wire _51329_;
wire _51330_;
wire _51331_;
wire _51332_;
wire _51333_;
wire _51334_;
wire _51335_;
wire _51336_;
wire _51337_;
wire _51338_;
wire _51339_;
wire _51340_;
wire _51341_;
wire _51342_;
wire _51343_;
wire _51344_;
wire _51345_;
wire _51346_;
wire _51347_;
wire _51348_;
wire _51349_;
wire _51350_;
wire _51351_;
wire _51352_;
wire _51353_;
wire _51354_;
wire _51355_;
wire _51356_;
wire _51357_;
wire _51358_;
wire _51359_;
wire _51360_;
wire _51361_;
wire _51362_;
wire _51363_;
wire _51364_;
wire _51365_;
wire _51366_;
wire _51367_;
wire _51368_;
wire _51369_;
wire _51370_;
wire _51371_;
wire _51372_;
wire _51373_;
wire _51374_;
wire _51375_;
wire _51376_;
wire _51377_;
wire _51378_;
wire _51379_;
wire _51380_;
wire _51381_;
wire _51382_;
wire _51383_;
wire _51384_;
wire _51385_;
wire _51386_;
wire _51387_;
wire _51388_;
wire _51389_;
wire _51390_;
wire _51391_;
wire _51392_;
wire _51393_;
wire _51394_;
wire _51395_;
wire _51396_;
wire _51397_;
wire _51398_;
wire _51399_;
wire _51400_;
wire _51401_;
wire _51402_;
wire _51403_;
wire _51404_;
wire _51405_;
wire _51406_;
wire _51407_;
wire _51408_;
wire _51409_;
wire _51410_;
wire _51411_;
wire _51412_;
wire _51413_;
wire _51414_;
wire _51415_;
wire _51416_;
wire _51417_;
wire _51418_;
wire _51419_;
wire _51420_;
wire _51421_;
wire _51422_;
wire _51423_;
wire _51424_;
wire _51425_;
wire _51426_;
wire _51427_;
wire _51428_;
wire _51429_;
wire _51430_;
wire _51431_;
wire _51432_;
wire _51433_;
wire _51434_;
wire _51435_;
wire _51436_;
wire _51437_;
wire _51438_;
wire _51439_;
wire _51440_;
wire _51441_;
wire _51442_;
wire _51443_;
wire _51444_;
wire _51445_;
wire _51446_;
wire _51447_;
wire _51448_;
wire _51449_;
wire _51450_;
wire _51451_;
wire _51452_;
wire _51453_;
wire _51454_;
wire _51455_;
wire _51456_;
wire _51457_;
wire _51458_;
wire _51459_;
wire _51460_;
wire _51461_;
wire _51462_;
wire _51463_;
wire _51464_;
wire _51465_;
wire _51466_;
wire _51467_;
wire _51468_;
wire _51469_;
wire _51470_;
wire _51471_;
wire _51472_;
wire _51473_;
wire _51474_;
wire _51475_;
wire _51476_;
wire _51477_;
wire _51478_;
wire _51479_;
wire _51480_;
wire _51481_;
wire _51482_;
wire _51483_;
wire _51484_;
wire _51485_;
wire _51486_;
wire _51487_;
wire _51488_;
wire _51489_;
wire _51490_;
wire _51491_;
wire _51492_;
wire _51493_;
wire _51494_;
wire _51495_;
wire _51496_;
wire _51497_;
wire _51498_;
wire _51499_;
wire _51500_;
wire _51501_;
wire _51502_;
wire _51503_;
wire _51504_;
wire _51505_;
wire _51506_;
wire _51507_;
wire _51508_;
wire _51509_;
wire _51510_;
wire _51511_;
wire _51512_;
wire _51513_;
wire _51514_;
wire _51515_;
wire _51516_;
wire _51517_;
wire _51518_;
wire _51519_;
wire _51520_;
wire _51521_;
wire _51522_;
wire _51523_;
wire _51524_;
wire _51525_;
wire _51526_;
wire _51527_;
wire _51528_;
wire _51529_;
wire _51530_;
wire _51531_;
wire _51532_;
wire _51533_;
wire _51534_;
wire _51535_;
wire _51536_;
wire _51537_;
wire _51538_;
wire _51539_;
wire _51540_;
wire _51541_;
wire _51542_;
wire _51543_;
wire _51544_;
wire _51545_;
wire _51546_;
wire _51547_;
wire _51548_;
wire _51549_;
wire _51550_;
wire _51551_;
wire _51552_;
wire _51553_;
wire _51554_;
wire _51555_;
wire _51556_;
wire _51557_;
wire _51558_;
wire _51559_;
wire _51560_;
wire _51561_;
wire _51562_;
wire _51563_;
wire _51564_;
wire _51565_;
wire _51566_;
wire _51567_;
wire _51568_;
wire _51569_;
wire _51570_;
wire _51571_;
wire _51572_;
wire _51573_;
wire _51574_;
wire _51575_;
wire _51576_;
wire _51577_;
wire _51578_;
wire _51579_;
wire _51580_;
wire _51581_;
wire _51582_;
wire _51583_;
wire _51584_;
wire _51585_;
wire _51586_;
wire _51587_;
wire _51588_;
wire _51589_;
wire _51590_;
wire _51591_;
wire _51592_;
wire _51593_;
wire _51594_;
wire _51595_;
wire _51596_;
wire _51597_;
wire _51598_;
wire _51599_;
wire _51600_;
wire _51601_;
wire _51602_;
wire _51603_;
wire _51604_;
wire _51605_;
wire _51606_;
wire _51607_;
wire _51608_;
wire _51609_;
wire _51610_;
wire _51611_;
wire _51612_;
wire _51613_;
wire _51614_;
wire _51615_;
wire _51616_;
wire _51617_;
wire _51618_;
wire _51619_;
wire _51620_;
wire _51621_;
wire _51622_;
wire _51623_;
wire _51624_;
wire _51625_;
wire _51626_;
wire _51627_;
wire _51628_;
wire _51629_;
wire _51630_;
wire _51631_;
wire _51632_;
wire _51633_;
wire _51634_;
wire _51635_;
wire _51636_;
wire _51637_;
wire _51638_;
wire _51639_;
wire _51640_;
wire _51641_;
wire _51642_;
wire _51643_;
wire _51644_;
wire _51645_;
wire _51646_;
wire _51647_;
wire _51648_;
wire _51649_;
wire _51650_;
wire _51651_;
wire _51652_;
wire _51653_;
wire _51654_;
wire _51655_;
wire _51656_;
wire _51657_;
wire _51658_;
wire _51659_;
wire _51660_;
wire _51661_;
wire _51662_;
wire _51663_;
wire _51664_;
wire _51665_;
wire _51666_;
wire _51667_;
wire _51668_;
wire _51669_;
wire _51670_;
wire _51671_;
wire _51672_;
wire _51673_;
wire _51674_;
wire _51675_;
wire _51676_;
wire _51677_;
wire _51678_;
wire _51679_;
wire _51680_;
wire _51681_;
wire _51682_;
wire _51683_;
wire _51684_;
wire _51685_;
wire _51686_;
wire _51687_;
wire _51688_;
wire _51689_;
wire _51690_;
wire _51691_;
wire _51692_;
wire _51693_;
wire _51694_;
wire _51695_;
wire _51696_;
wire _51697_;
wire _51698_;
wire _51699_;
wire _51700_;
wire _51701_;
wire _51702_;
wire _51703_;
wire _51704_;
wire _51705_;
wire _51706_;
wire _51707_;
wire _51708_;
wire _51709_;
wire _51710_;
wire _51711_;
wire _51712_;
wire _51713_;
wire _51714_;
wire _51715_;
wire _51716_;
wire _51717_;
wire _51718_;
wire _51719_;
wire _51720_;
wire _51721_;
wire _51722_;
wire _51723_;
wire _51724_;
wire _51725_;
wire _51726_;
wire _51727_;
wire _51728_;
wire _51729_;
wire _51730_;
wire _51731_;
wire _51732_;
wire _51733_;
wire _51734_;
wire _51735_;
wire _51736_;
wire _51737_;
wire _51738_;
wire _51739_;
wire _51740_;
wire _51741_;
wire _51742_;
wire _51743_;
wire _51744_;
wire _51745_;
wire _51746_;
wire _51747_;
wire _51748_;
wire _51749_;
wire _51750_;
wire _51751_;
wire _51752_;
wire _51753_;
wire _51754_;
wire _51755_;
wire _51756_;
wire _51757_;
wire _51758_;
wire _51759_;
wire _51760_;
wire _51761_;
wire _51762_;
wire _51763_;
wire _51764_;
wire _51765_;
wire _51766_;
wire _51767_;
wire _51768_;
wire _51769_;
wire _51770_;
wire _51771_;
wire _51772_;
wire _51773_;
wire _51774_;
wire _51775_;
wire _51776_;
wire _51777_;
wire _51778_;
wire _51779_;
wire _51780_;
wire _51781_;
wire _51782_;
wire _51783_;
wire _51784_;
wire _51785_;
wire _51786_;
wire _51787_;
wire _51788_;
wire _51789_;
wire _51790_;
wire _51791_;
wire _51792_;
wire _51793_;
wire _51794_;
wire _51795_;
wire _51796_;
wire _51797_;
wire _51798_;
wire _51799_;
wire _51800_;
wire _51801_;
wire _51802_;
wire _51803_;
wire _51804_;
wire _51805_;
wire _51806_;
wire _51807_;
wire _51808_;
wire _51809_;
wire _51810_;
wire _51811_;
wire _51812_;
wire _51813_;
wire _51814_;
wire _51815_;
wire _51816_;
wire _51817_;
wire _51818_;
wire _51819_;
wire _51820_;
wire _51821_;
wire _51822_;
wire _51823_;
wire _51824_;
wire _51825_;
wire _51826_;
wire _51827_;
wire _51828_;
wire _51829_;
wire _51830_;
wire _51831_;
wire _51832_;
wire _51833_;
wire _51834_;
wire _51835_;
wire _51836_;
wire _51837_;
wire _51838_;
wire _51839_;
wire _51840_;
wire _51841_;
wire _51842_;
wire _51843_;
wire _51844_;
wire _51845_;
wire _51846_;
wire _51847_;
wire _51848_;
wire _51849_;
wire _51850_;
wire _51851_;
wire _51852_;
wire _51853_;
wire _51854_;
wire _51855_;
wire _51856_;
wire _51857_;
wire _51858_;
wire _51859_;
wire _51860_;
wire _51861_;
wire _51862_;
wire _51863_;
wire _51864_;
wire _51865_;
wire _51866_;
wire _51867_;
wire _51868_;
wire _51869_;
wire _51870_;
wire _51871_;
wire _51872_;
wire _51873_;
wire _51874_;
wire _51875_;
wire _51876_;
wire _51877_;
wire _51878_;
wire _51879_;
wire _51880_;
wire _51881_;
wire _51882_;
wire _51883_;
wire _51884_;
wire _51885_;
wire _51886_;
wire _51887_;
wire _51888_;
wire _51889_;
wire _51890_;
wire _51891_;
wire _51892_;
wire _51893_;
wire _51894_;
wire _51895_;
wire _51896_;
wire _51897_;
wire _51898_;
wire _51899_;
wire _51900_;
wire _51901_;
wire _51902_;
wire _51903_;
wire _51904_;
wire _51905_;
wire _51906_;
wire _51907_;
wire _51908_;
wire _51909_;
wire _51910_;
wire _51911_;
wire _51912_;
wire _51913_;
wire _51914_;
wire _51915_;
wire _51916_;
wire _51917_;
wire _51918_;
wire _51919_;
wire _51920_;
wire _51921_;
wire _51922_;
wire _51923_;
wire _51924_;
wire _51925_;
wire _51926_;
wire _51927_;
wire _51928_;
wire _51929_;
wire _51930_;
wire _51931_;
wire _51932_;
wire _51933_;
wire _51934_;
wire _51935_;
wire _51936_;
wire _51937_;
wire _51938_;
wire _51939_;
wire _51940_;
wire _51941_;
wire _51942_;
wire _51943_;
wire _51944_;
wire _51945_;
wire _51946_;
wire _51947_;
wire _51948_;
wire _51949_;
wire _51950_;
wire _51951_;
wire _51952_;
wire _51953_;
wire _51954_;
wire _51955_;
wire _51956_;
wire _51957_;
wire _51958_;
wire _51959_;
wire _51960_;
wire _51961_;
wire _51962_;
wire _51963_;
wire _51964_;
wire _51965_;
wire _51966_;
wire _51967_;
wire _51968_;
wire _51969_;
wire _51970_;
wire _51971_;
wire _51972_;
wire _51973_;
wire _51974_;
wire _51975_;
wire _51976_;
wire _51977_;
wire _51978_;
wire _51979_;
wire _51980_;
wire _51981_;
wire _51982_;
wire _51983_;
wire _51984_;
wire _51985_;
wire _51986_;
wire _51987_;
wire _51988_;
wire _51989_;
wire _51990_;
wire _51991_;
wire _51992_;
wire _51993_;
wire _51994_;
wire _51995_;
wire _51996_;
wire _51997_;
wire _51998_;
wire _51999_;
wire _52000_;
wire _52001_;
wire _52002_;
wire _52003_;
wire _52004_;
wire _52005_;
wire _52006_;
wire _52007_;
wire _52008_;
wire _52009_;
wire _52010_;
wire _52011_;
wire _52012_;
wire _52013_;
wire _52014_;
wire _52015_;
wire _52016_;
wire _52017_;
wire _52018_;
wire _52019_;
wire _52020_;
wire _52021_;
wire _52022_;
wire _52023_;
wire _52024_;
wire _52025_;
wire _52026_;
wire _52027_;
wire _52028_;
wire _52029_;
wire _52030_;
wire _52031_;
wire _52032_;
wire _52033_;
wire _52034_;
wire _52035_;
wire _52036_;
wire _52037_;
wire _52038_;
wire _52039_;
wire _52040_;
wire _52041_;
wire _52042_;
wire _52043_;
wire _52044_;
wire _52045_;
wire _52046_;
wire _52047_;
wire _52048_;
wire _52049_;
wire _52050_;
wire _52051_;
wire _52052_;
wire _52053_;
wire _52054_;
wire _52055_;
wire _52056_;
wire _52057_;
wire _52058_;
wire _52059_;
wire _52060_;
wire _52061_;
wire _52062_;
wire _52063_;
wire _52064_;
wire _52065_;
wire _52066_;
wire _52067_;
wire _52068_;
wire _52069_;
wire _52070_;
wire _52071_;
wire _52072_;
wire _52073_;
wire _52074_;
wire _52075_;
wire _52076_;
wire _52077_;
wire _52078_;
wire _52079_;
wire _52080_;
wire _52081_;
wire _52082_;
wire _52083_;
wire _52084_;
wire _52085_;
wire _52086_;
wire _52087_;
wire _52088_;
wire _52089_;
wire _52090_;
wire _52091_;
wire _52092_;
wire _52093_;
wire _52094_;
wire _52095_;
wire _52096_;
wire _52097_;
wire _52098_;
wire _52099_;
wire _52100_;
wire _52101_;
wire _52102_;
wire _52103_;
wire _52104_;
wire _52105_;
wire _52106_;
wire _52107_;
wire _52108_;
wire _52109_;
wire _52110_;
wire _52111_;
wire _52112_;
wire _52113_;
wire _52114_;
wire _52115_;
wire _52116_;
wire _52117_;
wire _52118_;
wire _52119_;
wire _52120_;
wire _52121_;
wire _52122_;
wire _52123_;
wire _52124_;
wire _52125_;
wire _52126_;
wire _52127_;
wire _52128_;
wire _52129_;
wire _52130_;
wire _52131_;
wire _52132_;
wire _52133_;
wire _52134_;
wire _52135_;
wire _52136_;
wire _52137_;
wire _52138_;
wire _52139_;
wire _52140_;
wire _52141_;
wire _52142_;
wire _52143_;
wire _52144_;
wire _52145_;
wire _52146_;
wire _52147_;
wire _52148_;
wire _52149_;
wire _52150_;
wire _52151_;
wire _52152_;
wire _52153_;
wire _52154_;
wire _52155_;
wire _52156_;
wire _52157_;
wire _52158_;
wire _52159_;
wire _52160_;
wire _52161_;
wire _52162_;
wire _52163_;
wire _52164_;
wire _52165_;
wire _52166_;
wire _52167_;
wire _52168_;
wire _52169_;
wire _52170_;
wire _52171_;
wire _52172_;
wire _52173_;
wire _52174_;
wire _52175_;
wire _52176_;
wire _52177_;
wire _52178_;
wire _52179_;
wire _52180_;
wire _52181_;
wire _52182_;
wire _52183_;
wire _52184_;
wire _52185_;
wire _52186_;
wire _52187_;
wire _52188_;
wire _52189_;
wire _52190_;
wire _52191_;
wire _52192_;
wire _52193_;
wire _52194_;
wire _52195_;
wire _52196_;
wire _52197_;
wire _52198_;
wire _52199_;
wire _52200_;
wire _52201_;
wire _52202_;
wire _52203_;
wire _52204_;
wire _52205_;
wire _52206_;
wire _52207_;
wire _52208_;
wire _52209_;
wire _52210_;
wire _52211_;
wire _52212_;
wire _52213_;
wire _52214_;
wire _52215_;
wire _52216_;
wire _52217_;
wire _52218_;
wire _52219_;
wire _52220_;
wire _52221_;
wire _52222_;
wire _52223_;
wire _52224_;
wire _52225_;
wire _52226_;
wire _52227_;
wire _52228_;
wire _52229_;
wire _52230_;
wire _52231_;
wire _52232_;
wire _52233_;
wire _52234_;
wire _52235_;
wire _52236_;
wire _52237_;
wire _52238_;
wire _52239_;
wire _52240_;
wire _52241_;
wire _52242_;
wire _52243_;
wire _52244_;
wire _52245_;
wire _52246_;
wire _52247_;
wire _52248_;
wire _52249_;
wire _52250_;
wire _52251_;
wire _52252_;
wire _52253_;
wire _52254_;
wire _52255_;
wire _52256_;
wire _52257_;
wire _52258_;
wire _52259_;
wire _52260_;
wire _52261_;
wire _52262_;
wire _52263_;
wire _52264_;
wire _52265_;
wire _52266_;
wire _52267_;
wire _52268_;
wire _52269_;
wire _52270_;
wire _52271_;
wire _52272_;
wire _52273_;
wire _52274_;
wire _52275_;
wire _52276_;
wire _52277_;
wire _52278_;
wire _52279_;
wire _52280_;
wire _52281_;
wire _52282_;
wire _52283_;
wire _52284_;
wire _52285_;
wire _52286_;
wire _52287_;
wire _52288_;
wire _52289_;
wire _52290_;
wire _52291_;
wire _52292_;
wire _52293_;
wire _52294_;
wire _52295_;
wire _52296_;
wire _52297_;
wire _52298_;
wire _52299_;
wire _52300_;
wire _52301_;
wire _52302_;
wire _52303_;
wire _52304_;
wire _52305_;
wire _52306_;
wire _52307_;
wire _52308_;
wire _52309_;
wire _52310_;
wire _52311_;
wire _52312_;
wire _52313_;
wire _52314_;
wire _52315_;
wire _52316_;
wire _52317_;
wire _52318_;
wire _52319_;
wire _52320_;
wire _52321_;
wire _52322_;
wire _52323_;
wire _52324_;
wire _52325_;
wire _52326_;
wire _52327_;
wire _52328_;
wire _52329_;
wire _52330_;
wire _52331_;
wire _52332_;
wire _52333_;
wire _52334_;
wire _52335_;
wire _52336_;
wire _52337_;
wire _52338_;
wire _52339_;
wire _52340_;
wire _52341_;
wire _52342_;
wire _52343_;
wire _52344_;
wire _52345_;
wire _52346_;
wire _52347_;
wire _52348_;
wire _52349_;
wire _52350_;
wire _52351_;
wire _52352_;
wire _52353_;
wire _52354_;
wire _52355_;
wire _52356_;
wire _52357_;
wire _52358_;
wire _52359_;
wire _52360_;
wire _52361_;
wire _52362_;
wire _52363_;
wire _52364_;
wire _52365_;
wire _52366_;
wire _52367_;
wire _52368_;
wire _52369_;
wire _52370_;
wire _52371_;
wire _52372_;
wire _52373_;
wire _52374_;
wire _52375_;
wire _52376_;
wire _52377_;
wire _52378_;
wire _52379_;
wire _52380_;
wire _52381_;
wire _52382_;
wire _52383_;
wire _52384_;
wire _52385_;
wire _52386_;
wire _52387_;
wire _52388_;
wire _52389_;
wire _52390_;
wire _52391_;
wire _52392_;
wire _52393_;
wire _52394_;
wire _52395_;
wire _52396_;
wire _52397_;
wire _52398_;
wire _52399_;
wire _52400_;
wire _52401_;
wire _52402_;
wire _52403_;
wire _52404_;
wire _52405_;
wire _52406_;
wire _52407_;
wire _52408_;
wire _52409_;
wire _52410_;
wire _52411_;
wire _52412_;
wire _52413_;
wire _52414_;
wire _52415_;
wire _52416_;
wire _52417_;
wire _52418_;
wire _52419_;
wire _52420_;
wire _52421_;
wire _52422_;
wire _52423_;
wire _52424_;
wire _52425_;
wire _52426_;
wire _52427_;
wire _52428_;
wire _52429_;
wire _52430_;
wire _52431_;
wire _52432_;
wire _52433_;
wire _52434_;
wire _52435_;
wire _52436_;
wire _52437_;
wire _52438_;
wire _52439_;
wire _52440_;
wire _52441_;
wire _52442_;
wire _52443_;
wire _52444_;
wire _52445_;
wire _52446_;
wire _52447_;
wire _52448_;
wire _52449_;
wire _52450_;
wire _52451_;
wire _52452_;
wire _52453_;
wire _52454_;
wire _52455_;
wire _52456_;
wire _52457_;
wire _52458_;
wire _52459_;
wire _52460_;
wire _52461_;
wire _52462_;
wire _52463_;
wire _52464_;
wire _52465_;
wire _52466_;
wire _52467_;
wire _52468_;
wire _52469_;
wire _52470_;
wire _52471_;
wire _52472_;
wire _52473_;
wire _52474_;
wire _52475_;
wire _52476_;
wire _52477_;
wire _52478_;
wire _52479_;
wire _52480_;
wire _52481_;
wire _52482_;
wire _52483_;
wire _52484_;
wire _52485_;
wire _52486_;
wire _52487_;
wire _52488_;
wire _52489_;
wire _52490_;
wire _52491_;
wire _52492_;
wire _52493_;
wire _52494_;
wire _52495_;
wire _52496_;
wire _52497_;
wire _52498_;
wire _52499_;
wire _52500_;
wire _52501_;
wire _52502_;
wire _52503_;
wire _52504_;
wire _52505_;
wire _52506_;
wire _52507_;
wire _52508_;
wire _52509_;
wire _52510_;
wire _52511_;
wire _52512_;
wire _52513_;
wire _52514_;
wire _52515_;
wire _52516_;
wire _52517_;
wire _52518_;
wire _52519_;
wire _52520_;
wire _52521_;
wire _52522_;
wire _52523_;
wire _52524_;
wire _52525_;
wire _52526_;
wire _52527_;
wire _52528_;
wire _52529_;
wire _52530_;
wire _52531_;
wire _52532_;
wire _52533_;
wire _52534_;
wire _52535_;
wire _52536_;
wire _52537_;
wire _52538_;
wire _52539_;
wire _52540_;
wire _52541_;
wire _52542_;
wire _52543_;
wire _52544_;
wire _52545_;
wire _52546_;
wire _52547_;
wire _52548_;
wire _52549_;
wire _52550_;
wire _52551_;
wire _52552_;
wire _52553_;
wire _52554_;
wire _52555_;
wire _52556_;
wire _52557_;
wire _52558_;
wire _52559_;
wire _52560_;
wire _52561_;
wire _52562_;
wire _52563_;
wire _52564_;
wire _52565_;
wire _52566_;
wire _52567_;
wire _52568_;
wire _52569_;
wire _52570_;
wire _52571_;
wire _52572_;
wire _52573_;
wire _52574_;
wire _52575_;
wire _52576_;
wire _52577_;
wire _52578_;
wire _52579_;
wire _52580_;
wire _52581_;
wire _52582_;
wire _52583_;
wire _52584_;
wire _52585_;
wire _52586_;
wire _52587_;
wire _52588_;
wire _52589_;
wire _52590_;
wire _52591_;
wire _52592_;
wire _52593_;
wire _52594_;
wire _52595_;
wire _52596_;
wire _52597_;
wire _52598_;
wire _52599_;
wire _52600_;
wire _52601_;
wire _52602_;
wire _52603_;
wire _52604_;
wire _52605_;
wire _52606_;
wire _52607_;
wire _52608_;
wire _52609_;
wire _52610_;
wire _52611_;
wire _52612_;
wire _52613_;
wire _52614_;
wire _52615_;
wire _52616_;
wire _52617_;
wire _52618_;
wire _52619_;
wire _52620_;
wire _52621_;
wire _52622_;
wire _52623_;
wire _52624_;
wire _52625_;
wire _52626_;
wire _52627_;
wire _52628_;
wire _52629_;
wire _52630_;
wire _52631_;
wire _52632_;
wire _52633_;
wire _52634_;
wire _52635_;
wire _52636_;
wire _52637_;
wire _52638_;
wire _52639_;
wire _52640_;
wire _52641_;
wire _52642_;
wire _52643_;
wire _52644_;
wire _52645_;
wire _52646_;
wire _52647_;
wire _52648_;
wire _52649_;
wire _52650_;
wire _52651_;
wire _52652_;
wire _52653_;
wire _52654_;
wire _52655_;
wire _52656_;
wire _52657_;
wire _52658_;
wire _52659_;
wire _52660_;
wire _52661_;
wire _52662_;
wire _52663_;
wire _52664_;
wire _52665_;
wire _52666_;
wire _52667_;
wire _52668_;
wire _52669_;
wire _52670_;
wire _52671_;
wire _52672_;
wire _52673_;
wire _52674_;
wire _52675_;
wire _52676_;
wire _52677_;
wire _52678_;
wire _52679_;
wire _52680_;
wire _52681_;
wire _52682_;
wire _52683_;
wire _52684_;
wire _52685_;
wire _52686_;
wire _52687_;
wire _52688_;
wire _52689_;
wire _52690_;
wire _52691_;
wire _52692_;
wire _52693_;
wire _52694_;
wire _52695_;
wire _52696_;
wire _52697_;
wire _52698_;
wire _52699_;
wire _52700_;
wire _52701_;
wire _52702_;
wire _52703_;
wire _52704_;
wire _52705_;
wire _52706_;
wire _52707_;
wire _52708_;
wire _52709_;
wire _52710_;
wire _52711_;
wire _52712_;
wire _52713_;
wire _52714_;
wire _52715_;
wire _52716_;
wire _52717_;
wire _52718_;
wire _52719_;
wire _52720_;
wire _52721_;
wire _52722_;
wire _52723_;
wire _52724_;
wire _52725_;
wire _52726_;
wire _52727_;
wire _52728_;
wire _52729_;
wire _52730_;
wire _52731_;
wire _52732_;
wire _52733_;
wire _52734_;
wire _52735_;
wire _52736_;
wire _52737_;
wire _52738_;
wire _52739_;
wire _52740_;
wire _52741_;
wire _52742_;
wire _52743_;
wire _52744_;
wire _52745_;
wire _52746_;
wire _52747_;
wire _52748_;
wire _52749_;
wire _52750_;
wire _52751_;
wire _52752_;
wire _52753_;
wire _52754_;
wire _52755_;
wire _52756_;
wire _52757_;
wire _52758_;
wire _52759_;
wire _52760_;
wire _52761_;
wire _52762_;
wire _52763_;
wire _52764_;
wire _52765_;
wire _52766_;
wire _52767_;
wire _52768_;
wire _52769_;
wire _52770_;
wire _52771_;
wire _52772_;
wire _52773_;
wire _52774_;
wire _52775_;
wire _52776_;
wire _52777_;
wire _52778_;
wire _52779_;
wire _52780_;
wire _52781_;
wire _52782_;
wire _52783_;
wire _52784_;
wire _52785_;
wire _52786_;
wire _52787_;
wire _52788_;
wire _52789_;
wire _52790_;
wire _52791_;
wire _52792_;
wire _52793_;
wire _52794_;
wire _52795_;
wire _52796_;
wire _52797_;
wire _52798_;
wire _52799_;
wire _52800_;
wire _52801_;
wire _52802_;
wire _52803_;
wire _52804_;
wire _52805_;
wire _52806_;
wire _52807_;
wire _52808_;
wire _52809_;
wire _52810_;
wire _52811_;
wire _52812_;
wire _52813_;
wire _52814_;
wire _52815_;
wire _52816_;
wire _52817_;
wire _52818_;
wire _52819_;
wire _52820_;
wire _52821_;
wire _52822_;
wire _52823_;
wire _52824_;
wire _52825_;
wire _52826_;
wire _52827_;
wire _52828_;
wire _52829_;
wire _52830_;
wire _52831_;
wire _52832_;
wire _52833_;
wire _52834_;
wire _52835_;
wire _52836_;
wire _52837_;
wire _52838_;
wire _52839_;
wire _52840_;
wire _52841_;
wire _52842_;
wire _52843_;
wire _52844_;
wire _52845_;
wire _52846_;
wire _52847_;
wire _52848_;
wire _52849_;
wire _52850_;
wire _52851_;
wire _52852_;
wire _52853_;
wire _52854_;
wire _52855_;
wire _52856_;
wire _52857_;
wire _52858_;
wire _52859_;
wire _52860_;
wire _52861_;
wire _52862_;
wire _52863_;
wire _52864_;
wire _52865_;
wire _52866_;
wire _52867_;
wire _52868_;
wire _52869_;
wire _52870_;
wire _52871_;
wire _52872_;
wire _52873_;
wire _52874_;
wire _52875_;
wire _52876_;
wire _52877_;
wire _52878_;
wire _52879_;
wire _52880_;
wire _52881_;
wire _52882_;
wire _52883_;
wire _52884_;
wire _52885_;
wire _52886_;
wire _52887_;
wire _52888_;
wire _52889_;
wire _52890_;
wire _52891_;
wire _52892_;
wire _52893_;
wire _52894_;
wire _52895_;
wire _52896_;
wire _52897_;
wire _52898_;
wire _52899_;
wire _52900_;
wire _52901_;
wire _52902_;
wire _52903_;
wire _52904_;
wire _52905_;
wire _52906_;
wire _52907_;
wire _52908_;
wire _52909_;
wire _52910_;
wire _52911_;
wire _52912_;
wire _52913_;
wire _52914_;
wire _52915_;
wire _52916_;
wire _52917_;
wire _52918_;
wire _52919_;
wire _52920_;
wire _52921_;
wire _52922_;
wire _52923_;
wire _52924_;
wire _52925_;
wire _52926_;
wire _52927_;
wire _52928_;
wire _52929_;
wire _52930_;
wire _52931_;
wire _52932_;
wire _52933_;
wire _52934_;
wire _52935_;
wire _52936_;
wire _52937_;
wire _52938_;
wire _52939_;
wire _52940_;
wire _52941_;
wire _52942_;
wire _52943_;
wire _52944_;
wire _52945_;
wire _52946_;
wire _52947_;
wire _52948_;
wire _52949_;
wire _52950_;
wire _52951_;
wire _52952_;
wire _52953_;
wire _52954_;
wire _52955_;
wire _52956_;
wire _52957_;
wire _52958_;
wire _52959_;
wire _52960_;
wire _52961_;
wire _52962_;
wire _52963_;
wire _52964_;
wire _52965_;
wire _52966_;
wire _52967_;
wire _52968_;
wire _52969_;
wire _52970_;
wire _52971_;
wire _52972_;
wire _52973_;
wire _52974_;
wire _52975_;
wire _52976_;
wire _52977_;
wire _52978_;
wire _52979_;
wire _52980_;
wire _52981_;
wire _52982_;
wire _52983_;
wire _52984_;
wire _52985_;
wire _52986_;
wire _52987_;
wire _52988_;
wire _52989_;
wire _52990_;
wire _52991_;
wire _52992_;
wire _52993_;
wire _52994_;
wire _52995_;
wire _52996_;
wire _52997_;
wire _52998_;
wire _52999_;
wire _53000_;
wire _53001_;
wire _53002_;
wire _53003_;
wire _53004_;
wire _53005_;
wire _53006_;
wire _53007_;
wire _53008_;
wire _53009_;
wire _53010_;
wire _53011_;
wire _53012_;
wire _53013_;
wire _53014_;
wire _53015_;
wire _53016_;
wire _53017_;
wire _53018_;
wire _53019_;
wire _53020_;
wire _53021_;
wire _53022_;
wire _53023_;
wire _53024_;
wire _53025_;
wire _53026_;
wire _53027_;
wire _53028_;
wire _53029_;
wire _53030_;
wire _53031_;
wire _53032_;
wire _53033_;
wire _53034_;
wire _53035_;
wire _53036_;
wire _53037_;
wire _53038_;
wire _53039_;
wire _53040_;
wire _53041_;
wire _53042_;
wire _53043_;
wire _53044_;
wire _53045_;
wire _53046_;
wire _53047_;
wire _53048_;
wire _53049_;
wire _53050_;
wire _53051_;
wire _53052_;
wire _53053_;
wire _53054_;
wire _53055_;
wire _53056_;
wire _53057_;
wire _53058_;
wire _53059_;
wire _53060_;
wire _53061_;
wire _53062_;
wire _53063_;
wire _53064_;
wire _53065_;
wire _53066_;
wire _53067_;
wire _53068_;
wire _53069_;
wire _53070_;
wire _53071_;
wire _53072_;
wire _53073_;
wire _53074_;
wire _53075_;
wire _53076_;
wire _53077_;
wire _53078_;
wire _53079_;
wire _53080_;
wire _53081_;
wire _53082_;
wire _53083_;
wire _53084_;
wire _53085_;
wire _53086_;
wire _53087_;
wire _53088_;
wire _53089_;
wire _53090_;
wire _53091_;
wire _53092_;
wire _53093_;
wire _53094_;
wire _53095_;
wire _53096_;
wire _53097_;
wire _53098_;
wire _53099_;
wire _53100_;
wire _53101_;
wire _53102_;
wire _53103_;
wire _53104_;
wire _53105_;
wire _53106_;
wire _53107_;
wire _53108_;
wire _53109_;
wire _53110_;
wire _53111_;
wire _53112_;
wire _53113_;
wire _53114_;
wire _53115_;
wire _53116_;
wire _53117_;
wire _53118_;
wire _53119_;
wire _53120_;
wire _53121_;
wire _53122_;
wire _53123_;
wire _53124_;
wire _53125_;
wire _53126_;
wire _53127_;
wire _53128_;
wire _53129_;
wire _53130_;
wire _53131_;
wire _53132_;
wire _53133_;
wire _53134_;
wire _53135_;
wire _53136_;
wire _53137_;
wire _53138_;
wire _53139_;
wire _53140_;
wire _53141_;
wire _53142_;
wire _53143_;
wire _53144_;
wire _53145_;
wire _53146_;
wire _53147_;
wire _53148_;
wire _53149_;
wire _53150_;
wire _53151_;
wire _53152_;
wire _53153_;
wire _53154_;
wire _53155_;
wire _53156_;
wire _53157_;
wire _53158_;
wire _53159_;
wire _53160_;
wire _53161_;
wire _53162_;
wire _53163_;
wire _53164_;
wire _53165_;
wire _53166_;
wire _53167_;
wire _53168_;
wire _53169_;
wire _53170_;
wire _53171_;
wire _53172_;
wire _53173_;
wire _53174_;
wire _53175_;
wire _53176_;
wire _53177_;
wire _53178_;
wire _53179_;
wire _53180_;
wire _53181_;
wire _53182_;
wire _53183_;
wire _53184_;
wire _53185_;
wire _53186_;
wire _53187_;
wire _53188_;
wire _53189_;
wire _53190_;
wire _53191_;
wire _53192_;
wire _53193_;
wire _53194_;
wire _53195_;
wire _53196_;
wire _53197_;
wire _53198_;
wire _53199_;
wire _53200_;
wire _53201_;
wire _53202_;
wire _53203_;
wire _53204_;
wire _53205_;
wire _53206_;
wire _53207_;
wire _53208_;
wire _53209_;
wire _53210_;
wire _53211_;
wire _53212_;
wire _53213_;
wire _53214_;
wire _53215_;
wire _53216_;
wire _53217_;
wire _53218_;
wire _53219_;
wire _53220_;
wire _53221_;
wire _53222_;
wire _53223_;
wire _53224_;
wire _53225_;
wire _53226_;
wire _53227_;
wire _53228_;
wire _53229_;
wire _53230_;
wire _53231_;
wire _53232_;
wire _53233_;
wire _53234_;
wire _53235_;
wire _53236_;
wire _53237_;
wire _53238_;
wire _53239_;
wire _53240_;
wire _53241_;
wire _53242_;
wire _53243_;
wire _53244_;
wire _53245_;
wire _53246_;
wire _53247_;
wire _53248_;
wire _53249_;
wire _53250_;
wire _53251_;
wire _53252_;
wire _53253_;
wire _53254_;
wire _53255_;
wire _53256_;
wire _53257_;
wire _53258_;
wire _53259_;
wire _53260_;
wire _53261_;
wire _53262_;
wire _53263_;
wire _53264_;
wire _53265_;
wire _53266_;
wire _53267_;
wire _53268_;
wire _53269_;
wire _53270_;
wire _53271_;
wire _53272_;
wire _53273_;
wire _53274_;
wire _53275_;
wire _53276_;
wire _53277_;
wire _53278_;
wire _53279_;
wire _53280_;
wire _53281_;
wire _53282_;
wire _53283_;
wire _53284_;
wire _53285_;
wire _53286_;
wire _53287_;
wire _53288_;
wire _53289_;
wire _53290_;
wire _53291_;
wire _53292_;
wire _53293_;
wire _53294_;
wire _53295_;
wire _53296_;
wire _53297_;
wire _53298_;
wire _53299_;
wire _53300_;
wire _53301_;
wire _53302_;
wire _53303_;
wire _53304_;
wire _53305_;
wire _53306_;
wire _53307_;
wire _53308_;
wire _53309_;
wire _53310_;
wire _53311_;
wire _53312_;
wire _53313_;
wire _53314_;
wire _53315_;
wire _53316_;
wire _53317_;
wire _53318_;
wire _53319_;
wire _53320_;
wire _53321_;
wire _53322_;
wire _53323_;
wire _53324_;
wire _53325_;
wire _53326_;
wire _53327_;
wire _53328_;
wire _53329_;
wire _53330_;
wire _53331_;
wire _53332_;
wire _53333_;
wire _53334_;
wire _53335_;
wire _53336_;
wire _53337_;
wire _53338_;
wire _53339_;
wire _53340_;
wire _53341_;
wire _53342_;
wire _53343_;
wire _53344_;
wire _53345_;
wire _53346_;
wire _53347_;
wire _53348_;
wire _53349_;
wire _53350_;
wire _53351_;
wire _53352_;
wire _53353_;
wire _53354_;
wire _53355_;
wire _53356_;
wire _53357_;
wire _53358_;
wire _53359_;
wire _53360_;
wire _53361_;
wire _53362_;
wire _53363_;
wire _53364_;
wire _53365_;
wire _53366_;
wire _53367_;
wire _53368_;
wire _53369_;
wire _53370_;
wire _53371_;
wire _53372_;
wire _53373_;
wire _53374_;
wire _53375_;
wire _53376_;
wire _53377_;
wire _53378_;
wire _53379_;
wire _53380_;
wire _53381_;
wire _53382_;
wire _53383_;
wire _53384_;
wire _53385_;
wire _53386_;
wire _53387_;
wire _53388_;
wire _53389_;
wire _53390_;
wire _53391_;
wire _53392_;
wire _53393_;
wire _53394_;
wire _53395_;
wire _53396_;
wire _53397_;
wire _53398_;
wire _53399_;
wire _53400_;
wire _53401_;
wire _53402_;
wire _53403_;
wire _53404_;
wire _53405_;
wire _53406_;
wire _53407_;
wire _53408_;
wire _53409_;
wire _53410_;
wire _53411_;
wire _53412_;
wire _53413_;
wire _53414_;
wire _53415_;
wire _53416_;
wire _53417_;
wire _53418_;
wire _53419_;
wire _53420_;
wire _53421_;
wire _53422_;
wire _53423_;
wire _53424_;
wire _53425_;
wire _53426_;
wire _53427_;
wire _53428_;
wire _53429_;
wire _53430_;
wire _53431_;
wire _53432_;
wire _53433_;
wire _53434_;
wire _53435_;
wire _53436_;
wire _53437_;
wire _53438_;
wire _53439_;
wire _53440_;
wire _53441_;
wire _53442_;
wire _53443_;
wire _53444_;
wire _53445_;
wire _53446_;
wire _53447_;
wire _53448_;
wire _53449_;
wire _53450_;
wire _53451_;
wire _53452_;
wire _53453_;
wire _53454_;
wire _53455_;
wire _53456_;
wire _53457_;
wire _53458_;
wire _53459_;
wire _53460_;
wire _53461_;
wire _53462_;
wire _53463_;
wire _53464_;
wire _53465_;
wire _53466_;
wire _53467_;
wire _53468_;
wire _53469_;
wire _53470_;
wire _53471_;
wire _53472_;
wire _53473_;
wire _53474_;
wire _53475_;
wire _53476_;
wire _53477_;
wire _53478_;
wire _53479_;
wire _53480_;
wire _53481_;
wire _53482_;
wire _53483_;
wire _53484_;
wire _53485_;
wire _53486_;
wire _53487_;
wire _53488_;
wire _53489_;
wire _53490_;
wire _53491_;
wire _53492_;
wire _53493_;
wire _53494_;
wire _53495_;
wire _53496_;
wire _53497_;
wire _53498_;
wire _53499_;
wire _53500_;
wire _53501_;
wire _53502_;
wire _53503_;
wire _53504_;
wire _53505_;
wire _53506_;
wire _53507_;
wire _53508_;
wire _53509_;
wire _53510_;
wire _53511_;
wire _53512_;
wire _53513_;
wire _53514_;
wire _53515_;
wire _53516_;
wire _53517_;
wire _53518_;
wire _53519_;
wire _53520_;
wire _53521_;
wire _53522_;
wire _53523_;
wire _53524_;
wire _53525_;
wire _53526_;
wire _53527_;
wire _53528_;
wire _53529_;
wire _53530_;
wire _53531_;
wire _53532_;
wire _53533_;
wire _53534_;
wire _53535_;
wire _53536_;
wire _53537_;
wire _53538_;
wire _53539_;
wire _53540_;
wire _53541_;
wire _53542_;
wire _53543_;
wire _53544_;
wire _53545_;
wire _53546_;
wire _53547_;
wire _53548_;
wire _53549_;
wire _53550_;
wire _53551_;
wire _53552_;
wire _53553_;
wire _53554_;
wire _53555_;
wire _53556_;
wire _53557_;
wire _53558_;
wire _53559_;
wire _53560_;
wire _53561_;
wire _53562_;
wire _53563_;
wire _53564_;
wire _53565_;
wire _53566_;
wire _53567_;
wire _53568_;
wire _53569_;
wire _53570_;
wire _53571_;
wire _53572_;
wire _53573_;
wire _53574_;
wire _53575_;
wire _53576_;
wire _53577_;
wire _53578_;
wire _53579_;
wire _53580_;
wire _53581_;
wire _53582_;
wire _53583_;
wire _53584_;
wire _53585_;
wire _53586_;
wire _53587_;
wire _53588_;
wire _53589_;
wire _53590_;
wire _53591_;
wire _53592_;
wire _53593_;
wire _53594_;
wire _53595_;
wire _53596_;
wire _53597_;
wire _53598_;
wire _53599_;
wire _53600_;
wire _53601_;
wire _53602_;
wire _53603_;
wire _53604_;
wire _53605_;
wire _53606_;
wire _53607_;
wire _53608_;
wire _53609_;
wire _53610_;
wire _53611_;
wire _53612_;
wire _53613_;
wire _53614_;
wire _53615_;
wire _53616_;
wire _53617_;
wire _53618_;
wire _53619_;
wire _53620_;
wire _53621_;
wire _53622_;
wire _53623_;
wire _53624_;
wire _53625_;
wire _53626_;
wire _53627_;
wire _53628_;
wire _53629_;
wire _53630_;
wire _53631_;
wire _53632_;
wire _53633_;
wire _53634_;
wire _53635_;
wire _53636_;
wire _53637_;
wire _53638_;
wire _53639_;
wire _53640_;
wire _53641_;
wire _53642_;
wire _53643_;
wire _53644_;
wire _53645_;
wire _53646_;
wire _53647_;
wire _53648_;
wire _53649_;
wire _53650_;
wire _53651_;
wire _53652_;
wire _53653_;
wire _53654_;
wire _53655_;
wire _53656_;
wire _53657_;
wire _53658_;
wire _53659_;
wire _53660_;
wire _53661_;
wire _53662_;
wire _53663_;
wire _53664_;
wire _53665_;
wire _53666_;
wire _53667_;
wire _53668_;
wire _53669_;
wire _53670_;
wire _53671_;
wire _53672_;
wire _53673_;
wire _53674_;
wire _53675_;
wire _53676_;
wire _53677_;
wire _53678_;
wire _53679_;
wire _53680_;
wire _53681_;
wire _53682_;
wire _53683_;
wire _53684_;
wire _53685_;
wire _53686_;
wire _53687_;
wire _53688_;
wire _53689_;
wire _53690_;
wire _53691_;
wire _53692_;
wire _53693_;
wire _53694_;
wire _53695_;
wire _53696_;
wire _53697_;
wire _53698_;
wire _53699_;
wire _53700_;
wire _53701_;
wire _53702_;
wire _53703_;
wire _53704_;
wire _53705_;
wire _53706_;
wire _53707_;
wire _53708_;
wire _53709_;
wire _53710_;
wire _53711_;
wire _53712_;
wire _53713_;
wire _53714_;
wire _53715_;
wire _53716_;
wire _53717_;
wire _53718_;
wire _53719_;
wire _53720_;
wire _53721_;
wire _53722_;
wire _53723_;
wire _53724_;
wire _53725_;
wire _53726_;
wire _53727_;
wire _53728_;
wire _53729_;
wire _53730_;
wire _53731_;
wire _53732_;
wire _53733_;
wire _53734_;
wire _53735_;
wire _53736_;
wire _53737_;
wire _53738_;
wire _53739_;
wire _53740_;
wire _53741_;
wire _53742_;
wire _53743_;
wire _53744_;
wire _53745_;
wire _53746_;
wire _53747_;
wire _53748_;
wire _53749_;
wire _53750_;
wire _53751_;
wire _53752_;
wire _53753_;
wire _53754_;
wire _53755_;
wire _53756_;
wire _53757_;
wire _53758_;
wire _53759_;
wire _53760_;
wire _53761_;
wire _53762_;
wire _53763_;
wire _53764_;
wire _53765_;
wire _53766_;
wire _53767_;
wire _53768_;
wire _53769_;
wire _53770_;
wire _53771_;
wire _53772_;
wire _53773_;
wire _53774_;
wire _53775_;
wire _53776_;
wire _53777_;
wire _53778_;
wire _53779_;
wire _53780_;
wire _53781_;
wire _53782_;
wire _53783_;
wire _53784_;
wire _53785_;
wire _53786_;
wire _53787_;
wire _53788_;
wire _53789_;
wire _53790_;
wire _53791_;
wire _53792_;
wire _53793_;
wire _53794_;
wire _53795_;
wire _53796_;
wire _53797_;
wire _53798_;
wire _53799_;
wire _53800_;
wire _53801_;
wire _53802_;
wire _53803_;
wire _53804_;
wire _53805_;
wire _53806_;
wire _53807_;
wire _53808_;
wire _53809_;
wire _53810_;
wire _53811_;
wire _53812_;
wire _53813_;
wire _53814_;
wire _53815_;
wire _53816_;
wire _53817_;
wire _53818_;
wire _53819_;
wire _53820_;
wire _53821_;
wire _53822_;
wire _53823_;
wire _53824_;
wire _53825_;
wire _53826_;
wire _53827_;
wire _53828_;
wire _53829_;
wire _53830_;
wire _53831_;
wire _53832_;
wire _53833_;
wire _53834_;
wire _53835_;
wire _53836_;
wire _53837_;
wire _53838_;
wire _53839_;
wire _53840_;
wire _53841_;
wire _53842_;
wire _53843_;
wire _53844_;
wire _53845_;
wire _53846_;
wire _53847_;
wire _53848_;
wire _53849_;
wire _53850_;
wire _53851_;
wire _53852_;
wire _53853_;
wire _53854_;
wire _53855_;
wire _53856_;
wire _53857_;
wire _53858_;
wire _53859_;
wire _53860_;
wire _53861_;
wire _53862_;
wire _53863_;
wire _53864_;
wire _53865_;
wire _53866_;
wire _53867_;
wire _53868_;
wire _53869_;
wire _53870_;
wire _53871_;
wire _53872_;
wire _53873_;
wire _53874_;
wire _53875_;
wire _53876_;
wire _53877_;
wire _53878_;
wire _53879_;
wire _53880_;
wire _53881_;
wire _53882_;
wire _53883_;
wire _53884_;
wire _53885_;
wire _53886_;
wire _53887_;
wire _53888_;
wire _53889_;
wire _53890_;
wire _53891_;
wire _53892_;
wire _53893_;
wire _53894_;
wire _53895_;
wire _53896_;
wire _53897_;
wire _53898_;
wire _53899_;
wire _53900_;
wire _53901_;
wire _53902_;
wire _53903_;
wire _53904_;
wire _53905_;
wire _53906_;
wire _53907_;
wire _53908_;
wire _53909_;
wire _53910_;
wire _53911_;
wire _53912_;
wire _53913_;
wire _53914_;
wire _53915_;
wire _53916_;
wire _53917_;
wire _53918_;
wire _53919_;
wire _53920_;
wire _53921_;
wire _53922_;
wire _53923_;
wire _53924_;
wire _53925_;
wire _53926_;
wire _53927_;
wire _53928_;
wire _53929_;
wire _53930_;
wire _53931_;
wire _53932_;
wire _53933_;
wire _53934_;
wire _53935_;
wire _53936_;
wire _53937_;
wire _53938_;
wire _53939_;
wire _53940_;
wire _53941_;
wire _53942_;
wire _53943_;
wire _53944_;
wire _53945_;
wire _53946_;
wire _53947_;
wire _53948_;
wire _53949_;
wire _53950_;
wire _53951_;
wire _53952_;
wire _53953_;
wire _53954_;
wire _53955_;
wire _53956_;
wire _53957_;
wire _53958_;
wire _53959_;
wire _53960_;
wire _53961_;
wire _53962_;
wire _53963_;
wire _53964_;
wire _53965_;
wire _53966_;
wire _53967_;
wire _53968_;
wire _53969_;
wire _53970_;
wire _53971_;
wire _53972_;
wire _53973_;
wire _53974_;
wire _53975_;
wire _53976_;
wire _53977_;
wire _53978_;
wire _53979_;
wire _53980_;
wire _53981_;
wire _53982_;
wire _53983_;
wire _53984_;
wire _53985_;
wire _53986_;
wire _53987_;
wire _53988_;
wire _53989_;
wire _53990_;
wire _53991_;
wire _53992_;
wire _53993_;
wire _53994_;
wire _53995_;
wire _53996_;
wire _53997_;
wire _53998_;
wire _53999_;
wire _54000_;
wire _54001_;
wire _54002_;
wire _54003_;
wire _54004_;
wire _54005_;
wire _54006_;
wire _54007_;
wire _54008_;
wire _54009_;
wire _54010_;
wire _54011_;
wire _54012_;
wire _54013_;
wire _54014_;
wire _54015_;
wire _54016_;
wire _54017_;
wire _54018_;
wire _54019_;
wire _54020_;
wire _54021_;
wire _54022_;
wire _54023_;
wire _54024_;
wire _54025_;
wire _54026_;
wire _54027_;
wire _54028_;
wire _54029_;
wire _54030_;
wire _54031_;
wire _54032_;
wire _54033_;
wire _54034_;
wire _54035_;
wire _54036_;
wire _54037_;
wire _54038_;
wire _54039_;
wire _54040_;
wire _54041_;
wire _54042_;
wire _54043_;
wire _54044_;
wire _54045_;
wire _54046_;
wire _54047_;
wire _54048_;
wire _54049_;
wire _54050_;
wire _54051_;
wire _54052_;
wire _54053_;
wire _54054_;
wire _54055_;
wire _54056_;
wire _54057_;
wire _54058_;
wire _54059_;
wire _54060_;
wire _54061_;
wire _54062_;
wire _54063_;
wire _54064_;
wire _54065_;
wire _54066_;
wire _54067_;
wire _54068_;
wire _54069_;
wire _54070_;
wire _54071_;
wire _54072_;
wire _54073_;
wire _54074_;
wire _54075_;
wire _54076_;
wire _54077_;
wire _54078_;
wire _54079_;
wire _54080_;
wire _54081_;
wire _54082_;
wire _54083_;
wire _54084_;
wire _54085_;
wire _54086_;
wire _54087_;
wire _54088_;
wire _54089_;
wire _54090_;
wire _54091_;
wire _54092_;
wire _54093_;
wire _54094_;
wire _54095_;
wire _54096_;
wire _54097_;
wire _54098_;
wire _54099_;
wire _54100_;
wire _54101_;
wire _54102_;
wire _54103_;
wire _54104_;
wire _54105_;
wire _54106_;
wire _54107_;
wire _54108_;
wire _54109_;
wire _54110_;
wire _54111_;
wire _54112_;
wire _54113_;
wire _54114_;
wire _54115_;
wire _54116_;
wire _54117_;
wire _54118_;
wire _54119_;
wire _54120_;
wire _54121_;
wire _54122_;
wire _54123_;
wire _54124_;
wire _54125_;
wire _54126_;
wire _54127_;
wire _54128_;
wire _54129_;
wire _54130_;
wire _54131_;
wire _54132_;
wire _54133_;
wire _54134_;
wire _54135_;
wire _54136_;
wire _54137_;
wire _54138_;
wire _54139_;
wire _54140_;
wire _54141_;
wire _54142_;
wire _54143_;
wire _54144_;
wire _54145_;
wire _54146_;
wire _54147_;
wire _54148_;
wire _54149_;
wire _54150_;
wire _54151_;
wire _54152_;
wire _54153_;
wire _54154_;
wire _54155_;
wire _54156_;
wire _54157_;
wire _54158_;
wire _54159_;
wire _54160_;
wire _54161_;
wire _54162_;
wire _54163_;
wire _54164_;
wire _54165_;
wire _54166_;
wire _54167_;
wire _54168_;
wire _54169_;
wire _54170_;
wire _54171_;
wire _54172_;
wire _54173_;
wire _54174_;
wire _54175_;
wire _54176_;
wire _54177_;
wire _54178_;
wire _54179_;
wire _54180_;
wire _54181_;
wire _54182_;
wire _54183_;
wire _54184_;
wire _54185_;
wire _54186_;
wire _54187_;
wire _54188_;
wire _54189_;
wire _54190_;
wire _54191_;
wire _54192_;
wire _54193_;
wire _54194_;
wire _54195_;
wire _54196_;
wire _54197_;
wire _54198_;
wire _54199_;
wire _54200_;
wire _54201_;
wire _54202_;
wire _54203_;
wire _54204_;
wire _54205_;
wire _54206_;
wire _54207_;
wire _54208_;
wire _54209_;
wire _54210_;
wire _54211_;
wire _54212_;
wire _54213_;
wire _54214_;
wire _54215_;
wire _54216_;
wire _54217_;
wire _54218_;
wire _54219_;
wire _54220_;
wire _54221_;
wire _54222_;
wire _54223_;
wire _54224_;
wire _54225_;
wire _54226_;
wire _54227_;
wire _54228_;
wire _54229_;
wire _54230_;
wire _54231_;
wire _54232_;
wire _54233_;
wire _54234_;
wire _54235_;
wire _54236_;
wire _54237_;
wire _54238_;
wire _54239_;
wire _54240_;
wire _54241_;
wire _54242_;
wire _54243_;
wire _54244_;
wire _54245_;
wire _54246_;
wire _54247_;
wire _54248_;
wire _54249_;
wire _54250_;
wire _54251_;
wire _54252_;
wire _54253_;
wire _54254_;
wire _54255_;
wire _54256_;
wire _54257_;
wire _54258_;
wire _54259_;
wire _54260_;
wire _54261_;
wire _54262_;
wire _54263_;
wire _54264_;
wire _54265_;
wire _54266_;
wire _54267_;
wire _54268_;
wire _54269_;
wire _54270_;
wire _54271_;
wire _54272_;
wire _54273_;
wire _54274_;
wire _54275_;
wire _54276_;
wire _54277_;
wire _54278_;
wire _54279_;
wire _54280_;
wire _54281_;
wire _54282_;
wire _54283_;
wire _54284_;
wire _54285_;
wire _54286_;
wire _54287_;
wire _54288_;
wire _54289_;
wire _54290_;
wire _54291_;
wire _54292_;
wire _54293_;
wire _54294_;
wire _54295_;
wire _54296_;
wire _54297_;
wire _54298_;
wire _54299_;
wire _54300_;
wire _54301_;
wire _54302_;
wire _54303_;
wire _54304_;
wire _54305_;
wire _54306_;
wire _54307_;
wire _54308_;
wire _54309_;
wire _54310_;
wire _54311_;
wire _54312_;
wire _54313_;
wire _54314_;
wire _54315_;
wire _54316_;
wire _54317_;
wire _54318_;
wire _54319_;
wire _54320_;
wire _54321_;
wire _54322_;
wire _54323_;
wire _54324_;
wire _54325_;
wire _54326_;
wire _54327_;
wire _54328_;
wire _54329_;
wire _54330_;
wire _54331_;
wire _54332_;
wire _54333_;
wire _54334_;
wire _54335_;
wire _54336_;
wire _54337_;
wire _54338_;
wire _54339_;
wire _54340_;
wire _54341_;
wire _54342_;
wire _54343_;
wire _54344_;
wire _54345_;
wire _54346_;
wire _54347_;
wire _54348_;
wire _54349_;
wire _54350_;
wire _54351_;
wire _54352_;
wire _54353_;
wire _54354_;
wire _54355_;
wire _54356_;
wire _54357_;
wire _54358_;
wire _54359_;
wire _54360_;
wire _54361_;
wire _54362_;
wire _54363_;
wire _54364_;
wire _54365_;
wire _54366_;
wire _54367_;
wire _54368_;
wire _54369_;
wire _54370_;
wire _54371_;
wire _54372_;
wire _54373_;
wire _54374_;
wire _54375_;
wire _54376_;
wire _54377_;
wire _54378_;
wire _54379_;
wire _54380_;
wire _54381_;
wire _54382_;
wire _54383_;
wire _54384_;
wire _54385_;
wire _54386_;
wire _54387_;
wire _54388_;
wire _54389_;
wire _54390_;
wire _54391_;
wire _54392_;
wire _54393_;
wire _54394_;
wire _54395_;
wire _54396_;
wire _54397_;
wire _54398_;
wire _54399_;
wire _54400_;
wire _54401_;
wire _54402_;
wire _54403_;
wire _54404_;
wire _54405_;
wire _54406_;
wire _54407_;
wire _54408_;
wire _54409_;
wire _54410_;
wire _54411_;
wire _54412_;
wire _54413_;
wire _54414_;
wire _54415_;
wire _54416_;
wire _54417_;
wire _54418_;
wire _54419_;
wire _54420_;
wire _54421_;
wire _54422_;
wire _54423_;
wire _54424_;
wire _54425_;
wire _54426_;
wire _54427_;
wire _54428_;
wire _54429_;
wire _54430_;
wire _54431_;
wire _54432_;
wire _54433_;
wire _54434_;
wire _54435_;
wire _54436_;
wire _54437_;
wire _54438_;
wire _54439_;
wire _54440_;
wire _54441_;
wire _54442_;
wire _54443_;
wire _54444_;
wire _54445_;
wire _54446_;
wire _54447_;
wire _54448_;
wire _54449_;
wire _54450_;
wire _54451_;
wire _54452_;
wire _54453_;
wire _54454_;
wire _54455_;
wire _54456_;
wire _54457_;
wire _54458_;
wire _54459_;
wire _54460_;
wire _54461_;
wire _54462_;
wire _54463_;
wire _54464_;
wire _54465_;
wire _54466_;
wire _54467_;
wire _54468_;
wire _54469_;
wire _54470_;
wire _54471_;
wire _54472_;
wire _54473_;
wire _54474_;
wire _54475_;
wire _54476_;
wire _54477_;
wire _54478_;
wire _54479_;
wire _54480_;
wire _54481_;
wire _54482_;
wire _54483_;
wire _54484_;
wire _54485_;
wire _54486_;
wire _54487_;
wire _54488_;
wire _54489_;
wire _54490_;
wire _54491_;
wire _54492_;
wire _54493_;
wire _54494_;
wire _54495_;
wire _54496_;
wire _54497_;
wire _54498_;
wire _54499_;
wire _54500_;
wire _54501_;
wire _54502_;
wire _54503_;
wire _54504_;
wire _54505_;
wire _54506_;
wire _54507_;
wire _54508_;
wire _54509_;
wire _54510_;
wire _54511_;
wire _54512_;
wire _54513_;
wire _54514_;
wire _54515_;
wire _54516_;
wire _54517_;
wire _54518_;
wire _54519_;
wire _54520_;
wire _54521_;
wire _54522_;
wire _54523_;
wire _54524_;
wire _54525_;
wire _54526_;
wire _54527_;
wire _54528_;
wire _54529_;
wire _54530_;
wire _54531_;
wire _54532_;
wire _54533_;
wire _54534_;
wire _54535_;
wire _54536_;
wire _54537_;
wire _54538_;
wire _54539_;
wire _54540_;
wire _54541_;
wire _54542_;
wire _54543_;
wire _54544_;
wire _54545_;
wire _54546_;
wire _54547_;
wire _54548_;
wire _54549_;
wire _54550_;
wire _54551_;
wire _54552_;
wire _54553_;
wire _54554_;
wire _54555_;
wire _54556_;
wire _54557_;
wire _54558_;
wire _54559_;
wire _54560_;
wire _54561_;
wire _54562_;
wire _54563_;
wire _54564_;
wire _54565_;
wire _54566_;
wire _54567_;
wire _54568_;
wire _54569_;
wire _54570_;
wire _54571_;
wire _54572_;
wire _54573_;
wire _54574_;
wire _54575_;
wire _54576_;
wire _54577_;
wire _54578_;
wire _54579_;
wire _54580_;
wire _54581_;
wire _54582_;
wire _54583_;
wire _54584_;
wire _54585_;
wire _54586_;
wire _54587_;
wire _54588_;
wire _54589_;
wire _54590_;
wire _54591_;
wire _54592_;
wire _54593_;
wire _54594_;
wire _54595_;
wire _54596_;
wire _54597_;
wire _54598_;
wire _54599_;
wire _54600_;
wire _54601_;
wire _54602_;
wire _54603_;
wire _54604_;
wire _54605_;
wire _54606_;
wire _54607_;
wire _54608_;
wire _54609_;
wire _54610_;
wire _54611_;
wire _54612_;
wire _54613_;
wire _54614_;
wire _54615_;
wire _54616_;
wire _54617_;
wire _54618_;
wire _54619_;
wire _54620_;
wire _54621_;
wire _54622_;
wire _54623_;
wire _54624_;
wire _54625_;
wire _54626_;
wire _54627_;
wire _54628_;
wire _54629_;
wire _54630_;
wire _54631_;
wire _54632_;
wire _54633_;
wire _54634_;
wire _54635_;
wire _54636_;
wire _54637_;
wire _54638_;
wire _54639_;
wire _54640_;
wire _54641_;
wire _54642_;
wire _54643_;
wire _54644_;
wire _54645_;
wire _54646_;
wire _54647_;
wire _54648_;
wire _54649_;
wire _54650_;
wire _54651_;
wire _54652_;
wire _54653_;
wire _54654_;
wire _54655_;
wire _54656_;
wire _54657_;
wire _54658_;
wire _54659_;
wire _54660_;
wire _54661_;
wire _54662_;
wire _54663_;
wire _54664_;
wire _54665_;
wire _54666_;
wire _54667_;
wire _54668_;
wire _54669_;
wire _54670_;
wire _54671_;
wire _54672_;
wire _54673_;
wire _54674_;
wire _54675_;
wire _54676_;
wire _54677_;
wire _54678_;
wire _54679_;
wire _54680_;
wire _54681_;
wire _54682_;
wire _54683_;
wire _54684_;
wire _54685_;
wire _54686_;
wire _54687_;
wire _54688_;
wire _54689_;
wire _54690_;
wire _54691_;
wire _54692_;
wire _54693_;
wire _54694_;
wire _54695_;
wire _54696_;
wire _54697_;
wire _54698_;
wire _54699_;
wire _54700_;
wire _54701_;
wire _54702_;
wire _54703_;
wire _54704_;
wire _54705_;
wire _54706_;
wire _54707_;
wire _54708_;
wire _54709_;
wire _54710_;
wire _54711_;
wire _54712_;
wire _54713_;
wire _54714_;
wire _54715_;
wire _54716_;
wire _54717_;
wire _54718_;
wire _54719_;
wire _54720_;
wire _54721_;
wire _54722_;
wire _54723_;
wire _54724_;
wire _54725_;
wire _54726_;
wire _54727_;
wire _54728_;
wire _54729_;
wire _54730_;
wire _54731_;
wire _54732_;
wire _54733_;
wire _54734_;
wire _54735_;
wire _54736_;
wire _54737_;
wire _54738_;
wire _54739_;
wire _54740_;
wire _54741_;
wire _54742_;
wire _54743_;
wire _54744_;
wire _54745_;
wire _54746_;
wire _54747_;
wire _54748_;
wire _54749_;
wire _54750_;
wire _54751_;
wire _54752_;
wire _54753_;
wire _54754_;
wire _54755_;
wire _54756_;
wire _54757_;
wire _54758_;
wire _54759_;
wire _54760_;
wire _54761_;
wire _54762_;
wire _54763_;
wire _54764_;
wire _54765_;
wire _54766_;
wire _54767_;
wire _54768_;
wire _54769_;
wire _54770_;
wire _54771_;
wire _54772_;
wire _54773_;
wire _54774_;
wire _54775_;
wire _54776_;
wire _54777_;
wire _54778_;
wire _54779_;
wire _54780_;
wire _54781_;
wire _54782_;
wire _54783_;
wire _54784_;
wire _54785_;
wire _54786_;
wire _54787_;
wire _54788_;
wire _54789_;
wire _54790_;
wire _54791_;
wire _54792_;
wire _54793_;
wire _54794_;
wire _54795_;
wire _54796_;
wire _54797_;
wire _54798_;
wire _54799_;
wire _54800_;
wire _54801_;
wire _54802_;
wire _54803_;
wire _54804_;
wire _54805_;
wire _54806_;
wire _54807_;
wire _54808_;
wire _54809_;
wire _54810_;
wire _54811_;
wire _54812_;
wire _54813_;
wire _54814_;
wire _54815_;
wire _54816_;
wire _54817_;
wire _54818_;
wire _54819_;
wire _54820_;
wire _54821_;
wire _54822_;
wire _54823_;
wire _54824_;
wire _54825_;
wire _54826_;
wire _54827_;
wire _54828_;
wire _54829_;
wire _54830_;
wire _54831_;
wire _54832_;
wire _54833_;
wire _54834_;
wire _54835_;
wire _54836_;
wire _54837_;
wire _54838_;
wire _54839_;
wire _54840_;
wire _54841_;
wire _54842_;
wire _54843_;
wire _54844_;
wire _54845_;
wire _54846_;
wire _54847_;
wire _54848_;
wire _54849_;
wire _54850_;
wire _54851_;
wire _54852_;
wire _54853_;
wire _54854_;
wire _54855_;
wire _54856_;
wire _54857_;
wire _54858_;
wire _54859_;
wire _54860_;
wire _54861_;
wire _54862_;
wire _54863_;
wire _54864_;
wire _54865_;
wire _54866_;
wire _54867_;
wire _54868_;
wire _54869_;
wire _54870_;
wire _54871_;
wire _54872_;
wire _54873_;
wire _54874_;
wire _54875_;
wire _54876_;
wire _54877_;
wire _54878_;
wire _54879_;
wire _54880_;
wire _54881_;
wire _54882_;
wire _54883_;
wire _54884_;
wire _54885_;
wire _54886_;
wire _54887_;
wire _54888_;
wire _54889_;
wire _54890_;
wire _54891_;
wire _54892_;
wire _54893_;
wire _54894_;
wire _54895_;
wire _54896_;
wire _54897_;
wire _54898_;
wire _54899_;
wire _54900_;
wire _54901_;
wire _54902_;
wire _54903_;
wire _54904_;
wire _54905_;
wire _54906_;
wire _54907_;
wire _54908_;
wire _54909_;
wire _54910_;
wire _54911_;
wire _54912_;
wire _54913_;
wire _54914_;
wire _54915_;
wire _54916_;
wire _54917_;
wire _54918_;
wire _54919_;
wire _54920_;
wire _54921_;
wire _54922_;
wire _54923_;
wire _54924_;
wire _54925_;
wire _54926_;
wire _54927_;
wire _54928_;
wire _54929_;
wire _54930_;
wire _54931_;
wire _54932_;
wire _54933_;
wire _54934_;
wire _54935_;
wire _54936_;
wire _54937_;
wire _54938_;
wire _54939_;
wire _54940_;
wire _54941_;
wire _54942_;
wire _54943_;
wire _54944_;
wire _54945_;
wire _54946_;
wire _54947_;
wire _54948_;
wire _54949_;
wire _54950_;
wire _54951_;
wire _54952_;
wire _54953_;
wire _54954_;
wire _54955_;
wire _54956_;
wire _54957_;
wire _54958_;
wire _54959_;
wire _54960_;
wire _54961_;
wire _54962_;
wire _54963_;
wire _54964_;
wire _54965_;
wire _54966_;
wire _54967_;
wire _54968_;
wire _54969_;
wire _54970_;
wire _54971_;
wire _54972_;
wire _54973_;
wire _54974_;
wire _54975_;
wire _54976_;
wire _54977_;
wire _54978_;
wire _54979_;
wire _54980_;
wire _54981_;
wire _54982_;
wire _54983_;
wire _54984_;
wire _54985_;
wire _54986_;
wire _54987_;
wire _54988_;
wire _54989_;
wire _54990_;
wire _54991_;
wire _54992_;
wire _54993_;
wire _54994_;
wire _54995_;
wire _54996_;
wire _54997_;
wire _54998_;
wire _54999_;
wire _55000_;
wire _55001_;
wire _55002_;
wire _55003_;
wire _55004_;
wire _55005_;
wire _55006_;
wire _55007_;
wire _55008_;
wire _55009_;
wire _55010_;
wire _55011_;
wire _55012_;
wire _55013_;
wire _55014_;
wire _55015_;
wire _55016_;
wire _55017_;
wire _55018_;
wire _55019_;
wire _55020_;
wire _55021_;
wire _55022_;
wire _55023_;
wire _55024_;
wire _55025_;
wire _55026_;
wire _55027_;
wire _55028_;
wire _55029_;
wire _55030_;
wire _55031_;
wire _55032_;
wire _55033_;
wire _55034_;
wire _55035_;
wire _55036_;
wire _55037_;
wire _55038_;
wire _55039_;
wire _55040_;
wire _55041_;
wire _55042_;
wire _55043_;
wire _55044_;
wire _55045_;
wire _55046_;
wire _55047_;
wire _55048_;
wire _55049_;
wire _55050_;
wire _55051_;
wire _55052_;
wire _55053_;
wire _55054_;
wire _55055_;
wire _55056_;
wire _55057_;
wire _55058_;
wire _55059_;
wire _55060_;
wire _55061_;
wire _55062_;
wire _55063_;
wire _55064_;
wire _55065_;
wire _55066_;
wire _55067_;
wire _55068_;
wire _55069_;
wire _55070_;
wire _55071_;
wire _55072_;
wire _55073_;
wire _55074_;
wire _55075_;
wire _55076_;
wire _55077_;
wire _55078_;
wire _55079_;
wire _55080_;
wire _55081_;
wire _55082_;
wire _55083_;
wire _55084_;
wire _55085_;
wire _55086_;
wire _55087_;
wire _55088_;
wire _55089_;
wire _55090_;
wire _55091_;
wire _55092_;
wire _55093_;
wire _55094_;
wire _55095_;
wire _55096_;
wire _55097_;
wire _55098_;
wire _55099_;
wire _55100_;
wire _55101_;
wire _55102_;
wire _55103_;
wire _55104_;
wire _55105_;
wire _55106_;
wire _55107_;
wire _55108_;
wire _55109_;
wire _55110_;
wire _55111_;
wire _55112_;
wire _55113_;
wire _55114_;
wire _55115_;
wire _55116_;
wire _55117_;
wire _55118_;
wire _55119_;
wire _55120_;
wire _55121_;
wire _55122_;
wire _55123_;
wire _55124_;
wire _55125_;
wire _55126_;
wire _55127_;
wire _55128_;
wire _55129_;
wire _55130_;
wire _55131_;
wire _55132_;
wire _55133_;
wire _55134_;
wire _55135_;
wire _55136_;
wire _55137_;
wire _55138_;
wire _55139_;
wire _55140_;
wire _55141_;
wire _55142_;
wire _55143_;
wire _55144_;
wire _55145_;
wire _55146_;
wire _55147_;
wire _55148_;
wire _55149_;
wire _55150_;
wire _55151_;
wire _55152_;
wire _55153_;
wire _55154_;
wire _55155_;
wire _55156_;
wire _55157_;
wire _55158_;
wire _55159_;
wire _55160_;
wire _55161_;
wire _55162_;
wire _55163_;
wire _55164_;
wire _55165_;
wire _55166_;
wire _55167_;
wire _55168_;
wire _55169_;
wire _55170_;
wire _55171_;
wire _55172_;
wire _55173_;
wire _55174_;
wire _55175_;
wire _55176_;
wire _55177_;
wire _55178_;
wire _55179_;
wire _55180_;
wire _55181_;
wire _55182_;
wire _55183_;
wire _55184_;
wire _55185_;
wire _55186_;
wire _55187_;
wire _55188_;
wire _55189_;
wire _55190_;
wire _55191_;
wire _55192_;
wire _55193_;
wire _55194_;
wire _55195_;
wire _55196_;
wire _55197_;
wire _55198_;
wire _55199_;
wire _55200_;
wire _55201_;
wire _55202_;
wire _55203_;
wire _55204_;
wire _55205_;
wire _55206_;
wire _55207_;
wire _55208_;
wire _55209_;
wire _55210_;
wire _55211_;
wire _55212_;
wire _55213_;
wire _55214_;
wire _55215_;
wire _55216_;
wire _55217_;
wire _55218_;
wire _55219_;
wire _55220_;
wire _55221_;
wire _55222_;
wire _55223_;
wire _55224_;
wire _55225_;
wire _55226_;
wire _55227_;
wire _55228_;
wire _55229_;
wire _55230_;
wire _55231_;
wire _55232_;
wire _55233_;
wire _55234_;
wire _55235_;
wire _55236_;
wire _55237_;
wire _55238_;
wire _55239_;
wire _55240_;
wire _55241_;
wire _55242_;
wire _55243_;
wire _55244_;
wire _55245_;
wire _55246_;
wire _55247_;
wire _55248_;
wire _55249_;
wire _55250_;
wire _55251_;
wire _55252_;
wire _55253_;
wire _55254_;
wire _55255_;
wire _55256_;
wire _55257_;
wire _55258_;
wire _55259_;
wire _55260_;
wire _55261_;
wire _55262_;
wire _55263_;
wire _55264_;
wire _55265_;
wire _55266_;
wire _55267_;
wire _55268_;
wire _55269_;
wire _55270_;
wire _55271_;
wire _55272_;
wire _55273_;
wire _55274_;
wire _55275_;
wire _55276_;
wire _55277_;
wire _55278_;
wire _55279_;
wire _55280_;
wire _55281_;
wire _55282_;
wire _55283_;
wire _55284_;
wire _55285_;
wire _55286_;
wire _55287_;
wire _55288_;
wire _55289_;
wire _55290_;
wire _55291_;
wire _55292_;
wire _55293_;
wire _55294_;
wire _55295_;
wire _55296_;
wire _55297_;
wire _55298_;
wire _55299_;
wire _55300_;
wire _55301_;
wire _55302_;
wire _55303_;
wire _55304_;
wire _55305_;
wire _55306_;
wire _55307_;
wire _55308_;
wire _55309_;
wire _55310_;
wire _55311_;
wire _55312_;
wire _55313_;
wire _55314_;
wire _55315_;
wire _55316_;
wire _55317_;
wire _55318_;
wire _55319_;
wire _55320_;
wire _55321_;
wire _55322_;
wire _55323_;
wire _55324_;
wire _55325_;
wire _55326_;
wire _55327_;
wire _55328_;
wire _55329_;
wire _55330_;
wire _55331_;
wire _55332_;
wire _55333_;
wire _55334_;
wire _55335_;
wire _55336_;
wire _55337_;
wire _55338_;
wire _55339_;
wire _55340_;
wire _55341_;
wire _55342_;
wire _55343_;
wire _55344_;
wire _55345_;
wire _55346_;
wire _55347_;
wire _55348_;
wire _55349_;
wire _55350_;
wire _55351_;
wire _55352_;
wire _55353_;
wire _55354_;
wire _55355_;
wire _55356_;
wire _55357_;
wire _55358_;
wire _55359_;
wire _55360_;
wire _55361_;
wire _55362_;
wire _55363_;
wire _55364_;
wire _55365_;
wire _55366_;
wire _55367_;
wire _55368_;
wire _55369_;
wire _55370_;
wire _55371_;
wire _55372_;
wire _55373_;
wire _55374_;
wire _55375_;
wire _55376_;
wire _55377_;
wire _55378_;
wire _55379_;
wire _55380_;
wire _55381_;
wire _55382_;
wire _55383_;
wire _55384_;
wire _55385_;
wire _55386_;
wire _55387_;
wire _55388_;
wire _55389_;
wire _55390_;
wire _55391_;
wire _55392_;
wire _55393_;
wire _55394_;
wire _55395_;
wire _55396_;
wire _55397_;
wire _55398_;
wire _55399_;
wire _55400_;
wire _55401_;
wire _55402_;
wire _55403_;
wire _55404_;
wire _55405_;
wire _55406_;
wire _55407_;
wire _55408_;
wire _55409_;
wire _55410_;
wire _55411_;
wire _55412_;
wire _55413_;
wire _55414_;
wire _55415_;
wire _55416_;
wire _55417_;
wire _55418_;
wire _55419_;
wire _55420_;
wire _55421_;
wire _55422_;
wire _55423_;
wire _55424_;
wire _55425_;
wire _55426_;
wire _55427_;
wire _55428_;
wire _55429_;
wire _55430_;
wire _55431_;
wire _55432_;
wire _55433_;
wire _55434_;
wire _55435_;
wire _55436_;
wire _55437_;
wire _55438_;
wire _55439_;
wire _55440_;
wire _55441_;
wire _55442_;
wire _55443_;
wire _55444_;
wire _55445_;
wire _55446_;
wire _55447_;
wire _55448_;
wire _55449_;
wire _55450_;
wire _55451_;
wire _55452_;
wire _55453_;
wire _55454_;
wire _55455_;
wire _55456_;
wire _55457_;
wire _55458_;
wire _55459_;
wire _55460_;
wire _55461_;
wire _55462_;
wire _55463_;
wire _55464_;
wire _55465_;
wire _55466_;
wire _55467_;
wire _55468_;
wire _55469_;
wire _55470_;
wire _55471_;
wire _55472_;
wire _55473_;
wire _55474_;
wire _55475_;
wire _55476_;
wire _55477_;
wire _55478_;
wire _55479_;
wire _55480_;
wire _55481_;
wire _55482_;
wire _55483_;
wire _55484_;
wire _55485_;
wire _55486_;
wire _55487_;
wire _55488_;
wire _55489_;
wire _55490_;
wire _55491_;
wire _55492_;
wire _55493_;
wire _55494_;
wire _55495_;
wire _55496_;
wire _55497_;
wire _55498_;
wire _55499_;
wire _55500_;
wire _55501_;
wire _55502_;
wire _55503_;
wire _55504_;
wire _55505_;
wire _55506_;
wire _55507_;
wire _55508_;
wire _55509_;
wire _55510_;
wire _55511_;
wire _55512_;
wire _55513_;
wire _55514_;
wire _55515_;
wire _55516_;
wire _55517_;
wire _55518_;
wire _55519_;
wire _55520_;
wire _55521_;
wire _55522_;
wire _55523_;
wire _55524_;
wire _55525_;
wire _55526_;
wire _55527_;
wire _55528_;
wire _55529_;
wire _55530_;
wire _55531_;
wire _55532_;
wire _55533_;
wire _55534_;
wire _55535_;
wire _55536_;
wire _55537_;
wire _55538_;
wire _55539_;
wire _55540_;
wire _55541_;
wire _55542_;
wire _55543_;
wire _55544_;
wire _55545_;
wire _55546_;
wire _55547_;
wire _55548_;
wire _55549_;
wire _55550_;
wire _55551_;
wire _55552_;
wire _55553_;
wire _55554_;
wire _55555_;
wire _55556_;
wire _55557_;
wire _55558_;
wire _55559_;
wire _55560_;
wire _55561_;
wire _55562_;
wire _55563_;
wire _55564_;
wire _55565_;
wire _55566_;
wire _55567_;
wire _55568_;
wire _55569_;
wire _55570_;
wire _55571_;
wire _55572_;
wire _55573_;
wire _55574_;
wire _55575_;
wire _55576_;
wire _55577_;
wire _55578_;
wire _55579_;
wire _55580_;
wire _55581_;
wire _55582_;
wire _55583_;
wire _55584_;
wire _55585_;
wire _55586_;
wire _55587_;
wire _55588_;
wire _55589_;
wire _55590_;
wire _55591_;
wire _55592_;
wire _55593_;
wire _55594_;
wire _55595_;
wire _55596_;
wire _55597_;
wire _55598_;
wire _55599_;
wire _55600_;
wire _55601_;
wire _55602_;
wire _55603_;
wire _55604_;
wire _55605_;
wire _55606_;
wire _55607_;
wire _55608_;
wire _55609_;
wire _55610_;
wire _55611_;
wire _55612_;
wire _55613_;
wire _55614_;
wire _55615_;
wire _55616_;
wire _55617_;
wire _55618_;
wire _55619_;
wire _55620_;
wire _55621_;
wire _55622_;
wire _55623_;
wire _55624_;
wire _55625_;
wire _55626_;
wire _55627_;
wire _55628_;
wire _55629_;
wire _55630_;
wire _55631_;
wire _55632_;
wire _55633_;
wire _55634_;
wire _55635_;
wire _55636_;
wire _55637_;
wire _55638_;
wire _55639_;
wire _55640_;
wire _55641_;
wire _55642_;
wire _55643_;
wire _55644_;
wire _55645_;
wire _55646_;
wire _55647_;
wire _55648_;
wire _55649_;
wire _55650_;
wire _55651_;
wire _55652_;
wire _55653_;
wire _55654_;
wire _55655_;
wire _55656_;
wire _55657_;
wire _55658_;
wire _55659_;
wire _55660_;
wire _55661_;
wire _55662_;
wire _55663_;
wire _55664_;
wire _55665_;
wire _55666_;
wire _55667_;
wire _55668_;
wire _55669_;
wire _55670_;
wire _55671_;
wire _55672_;
wire _55673_;
wire _55674_;
wire _55675_;
wire _55676_;
wire _55677_;
wire _55678_;
wire _55679_;
wire _55680_;
wire _55681_;
wire _55682_;
wire _55683_;
wire _55684_;
wire _55685_;
wire _55686_;
wire _55687_;
wire _55688_;
wire _55689_;
wire _55690_;
wire _55691_;
wire _55692_;
wire _55693_;
wire _55694_;
wire _55695_;
wire _55696_;
wire _55697_;
wire _55698_;
wire _55699_;
wire _55700_;
wire _55701_;
wire _55702_;
wire _55703_;
wire _55704_;
wire _55705_;
wire _55706_;
wire _55707_;
wire _55708_;
wire _55709_;
wire _55710_;
wire _55711_;
wire _55712_;
wire _55713_;
wire _55714_;
wire _55715_;
wire _55716_;
wire _55717_;
wire _55718_;
wire _55719_;
wire _55720_;
wire _55721_;
wire _55722_;
wire _55723_;
wire _55724_;
wire _55725_;
wire _55726_;
wire _55727_;
wire _55728_;
wire _55729_;
wire _55730_;
wire _55731_;
wire _55732_;
wire _55733_;
wire _55734_;
wire _55735_;
wire _55736_;
wire _55737_;
wire _55738_;
wire _55739_;
wire _55740_;
wire _55741_;
wire _55742_;
wire _55743_;
wire _55744_;
wire _55745_;
wire _55746_;
wire _55747_;
wire _55748_;
wire _55749_;
wire _55750_;
wire _55751_;
wire _55752_;
wire _55753_;
wire _55754_;
wire _55755_;
wire _55756_;
wire _55757_;
wire _55758_;
wire _55759_;
wire _55760_;
wire _55761_;
wire _55762_;
wire _55763_;
wire _55764_;
wire _55765_;
wire _55766_;
wire _55767_;
wire _55768_;
wire _55769_;
wire _55770_;
wire _55771_;
wire _55772_;
wire _55773_;
wire _55774_;
wire _55775_;
wire _55776_;
wire _55777_;
wire _55778_;
wire _55779_;
wire _55780_;
wire _55781_;
wire _55782_;
wire _55783_;
wire _55784_;
wire _55785_;
wire _55786_;
wire _55787_;
wire _55788_;
wire _55789_;
wire _55790_;
wire _55791_;
wire _55792_;
wire _55793_;
wire _55794_;
wire _55795_;
wire _55796_;
wire _55797_;
wire _55798_;
wire _55799_;
wire _55800_;
wire _55801_;
wire _55802_;
wire _55803_;
wire _55804_;
wire _55805_;
wire _55806_;
wire _55807_;
wire _55808_;
wire _55809_;
wire _55810_;
wire _55811_;
wire _55812_;
wire _55813_;
wire _55814_;
wire _55815_;
wire _55816_;
wire _55817_;
wire _55818_;
wire _55819_;
wire _55820_;
wire _55821_;
wire _55822_;
wire _55823_;
wire _55824_;
wire _55825_;
wire _55826_;
wire _55827_;
wire _55828_;
wire _55829_;
wire _55830_;
wire _55831_;
wire _55832_;
wire _55833_;
wire _55834_;
wire _55835_;
wire _55836_;
wire _55837_;
wire _55838_;
wire _55839_;
wire _55840_;
wire _55841_;
wire _55842_;
wire _55843_;
wire _55844_;
wire _55845_;
wire _55846_;
wire _55847_;
wire _55848_;
wire _55849_;
wire _55850_;
wire _55851_;
wire _55852_;
wire _55853_;
wire _55854_;
wire _55855_;
wire _55856_;
wire _55857_;
wire _55858_;
wire _55859_;
wire _55860_;
wire _55861_;
wire _55862_;
wire _55863_;
wire _55864_;
wire _55865_;
wire _55866_;
wire _55867_;
wire _55868_;
wire _55869_;
wire _55870_;
wire _55871_;
wire _55872_;
wire _55873_;
wire _55874_;
wire _55875_;
wire _55876_;
wire _55877_;
wire _55878_;
wire _55879_;
wire _55880_;
wire _55881_;
wire _55882_;
wire _55883_;
wire _55884_;
wire _55885_;
wire _55886_;
wire _55887_;
wire _55888_;
wire _55889_;
wire _55890_;
wire _55891_;
wire _55892_;
wire _55893_;
wire _55894_;
wire _55895_;
wire _55896_;
wire _55897_;
wire _55898_;
wire _55899_;
wire _55900_;
wire _55901_;
wire _55902_;
wire _55903_;
wire _55904_;
wire _55905_;
wire _55906_;
wire _55907_;
wire _55908_;
wire _55909_;
wire _55910_;
wire _55911_;
wire _55912_;
wire _55913_;
wire _55914_;
wire _55915_;
wire _55916_;
wire _55917_;
wire _55918_;
wire _55919_;
wire _55920_;
wire _55921_;
wire _55922_;
wire _55923_;
wire _55924_;
wire _55925_;
wire _55926_;
wire _55927_;
wire _55928_;
wire _55929_;
wire _55930_;
wire _55931_;
wire _55932_;
wire _55933_;
wire _55934_;
wire _55935_;
wire _55936_;
wire _55937_;
wire _55938_;
wire _55939_;
wire _55940_;
wire _55941_;
wire _55942_;
wire _55943_;
wire _55944_;
wire _55945_;
wire _55946_;
wire _55947_;
wire _55948_;
wire _55949_;
wire _55950_;
wire _55951_;
wire _55952_;
wire _55953_;
wire _55954_;
wire _55955_;
wire _55956_;
wire _55957_;
wire _55958_;
wire _55959_;
wire _55960_;
wire _55961_;
wire _55962_;
wire _55963_;
wire _55964_;
wire _55965_;
wire _55966_;
wire _55967_;
wire _55968_;
wire _55969_;
wire _55970_;
wire _55971_;
wire _55972_;
wire _55973_;
wire _55974_;
wire _55975_;
wire _55976_;
wire _55977_;
wire _55978_;
wire _55979_;
wire _55980_;
wire _55981_;
wire _55982_;
wire _55983_;
wire _55984_;
wire _55985_;
wire _55986_;
wire _55987_;
wire _55988_;
wire _55989_;
wire _55990_;
wire _55991_;
wire _55992_;
wire _55993_;
wire _55994_;
wire _55995_;
wire _55996_;
wire _55997_;
wire _55998_;
wire _55999_;
wire _56000_;
wire _56001_;
wire _56002_;
wire _56003_;
wire _56004_;
wire _56005_;
wire _56006_;
wire _56007_;
wire _56008_;
wire _56009_;
wire _56010_;
wire _56011_;
wire _56012_;
wire _56013_;
wire _56014_;
wire _56015_;
wire _56016_;
wire _56017_;
wire _56018_;
wire _56019_;
wire _56020_;
wire _56021_;
wire _56022_;
wire _56023_;
wire _56024_;
wire _56025_;
wire _56026_;
wire _56027_;
wire _56028_;
wire _56029_;
wire _56030_;
wire _56031_;
wire _56032_;
wire _56033_;
wire _56034_;
wire _56035_;
wire _56036_;
wire _56037_;
wire _56038_;
wire _56039_;
wire _56040_;
wire _56041_;
wire _56042_;
wire _56043_;
wire _56044_;
wire _56045_;
wire _56046_;
wire _56047_;
wire _56048_;
wire _56049_;
wire _56050_;
wire _56051_;
wire _56052_;
wire _56053_;
wire _56054_;
wire _56055_;
wire _56056_;
wire _56057_;
wire _56058_;
wire _56059_;
wire _56060_;
wire _56061_;
wire _56062_;
wire _56063_;
wire _56064_;
wire _56065_;
wire _56066_;
wire _56067_;
wire _56068_;
wire _56069_;
wire _56070_;
wire _56071_;
wire _56072_;
wire _56073_;
wire _56074_;
wire _56075_;
wire _56076_;
wire _56077_;
wire _56078_;
wire _56079_;
wire _56080_;
wire _56081_;
wire _56082_;
wire _56083_;
wire _56084_;
wire _56085_;
wire _56086_;
wire _56087_;
wire _56088_;
wire _56089_;
wire _56090_;
wire _56091_;
wire _56092_;
wire _56093_;
wire _56094_;
wire _56095_;
wire _56096_;
wire _56097_;
wire _56098_;
wire _56099_;
wire _56100_;
wire _56101_;
wire _56102_;
wire _56103_;
wire _56104_;
wire _56105_;
wire _56106_;
wire _56107_;
wire _56108_;
wire _56109_;
wire _56110_;
wire _56111_;
wire _56112_;
wire _56113_;
wire _56114_;
wire _56115_;
wire _56116_;
wire _56117_;
wire _56118_;
wire _56119_;
wire _56120_;
wire _56121_;
wire _56122_;
wire _56123_;
wire _56124_;
wire _56125_;
wire _56126_;
wire _56127_;
wire _56128_;
wire _56129_;
wire _56130_;
wire _56131_;
wire _56132_;
wire _56133_;
wire _56134_;
wire _56135_;
wire _56136_;
wire _56137_;
wire _56138_;
wire _56139_;
wire _56140_;
wire _56141_;
wire _56142_;
wire _56143_;
wire _56144_;
wire _56145_;
wire _56146_;
wire _56147_;
wire _56148_;
wire _56149_;
wire _56150_;
wire _56151_;
wire _56152_;
wire _56153_;
wire _56154_;
wire _56155_;
wire _56156_;
wire _56157_;
wire _56158_;
wire _56159_;
wire _56160_;
wire _56161_;
wire _56162_;
wire _56163_;
wire _56164_;
wire _56165_;
wire _56166_;
wire _56167_;
wire _56168_;
wire _56169_;
wire _56170_;
wire _56171_;
wire _56172_;
wire _56173_;
wire _56174_;
wire _56175_;
wire _56176_;
wire _56177_;
wire _56178_;
wire _56179_;
wire _56180_;
wire _56181_;
wire _56182_;
wire _56183_;
wire _56184_;
wire _56185_;
wire _56186_;
wire _56187_;
wire _56188_;
wire _56189_;
wire _56190_;
wire _56191_;
wire _56192_;
wire _56193_;
wire _56194_;
wire _56195_;
wire _56196_;
wire _56197_;
wire _56198_;
wire _56199_;
wire _56200_;
wire _56201_;
wire _56202_;
wire _56203_;
wire _56204_;
wire _56205_;
wire _56206_;
wire _56207_;
wire _56208_;
wire _56209_;
wire _56210_;
wire _56211_;
wire _56212_;
wire _56213_;
wire _56214_;
wire _56215_;
wire _56216_;
wire _56217_;
wire _56218_;
wire _56219_;
wire _56220_;
wire _56221_;
wire _56222_;
wire _56223_;
wire _56224_;
wire _56225_;
wire _56226_;
wire _56227_;
wire _56228_;
wire _56229_;
wire _56230_;
wire _56231_;
wire _56232_;
wire _56233_;
wire _56234_;
wire _56235_;
wire _56236_;
wire _56237_;
wire _56238_;
wire _56239_;
wire _56240_;
wire _56241_;
wire _56242_;
wire _56243_;
wire _56244_;
wire _56245_;
wire _56246_;
wire _56247_;
wire _56248_;
wire _56249_;
wire _56250_;
wire _56251_;
wire _56252_;
wire _56253_;
wire _56254_;
wire _56255_;
wire _56256_;
wire _56257_;
wire _56258_;
wire _56259_;
wire _56260_;
wire _56261_;
wire _56262_;
wire _56263_;
wire _56264_;
wire _56265_;
wire _56266_;
wire _56267_;
wire _56268_;
wire _56269_;
wire _56270_;
wire _56271_;
wire _56272_;
wire _56273_;
wire _56274_;
wire _56275_;
wire _56276_;
wire _56277_;
wire _56278_;
wire _56279_;
wire _56280_;
wire _56281_;
wire _56282_;
wire _56283_;
wire _56284_;
wire _56285_;
wire _56286_;
wire _56287_;
wire _56288_;
wire _56289_;
wire _56290_;
wire _56291_;
wire _56292_;
wire _56293_;
wire _56294_;
wire _56295_;
wire _56296_;
wire _56297_;
wire _56298_;
wire _56299_;
wire _56300_;
wire _56301_;
wire _56302_;
wire _56303_;
wire _56304_;
wire _56305_;
wire _56306_;
wire _56307_;
wire _56308_;
wire _56309_;
wire _56310_;
wire _56311_;
wire _56312_;
wire _56313_;
wire _56314_;
wire _56315_;
wire _56316_;
wire _56317_;
wire _56318_;
wire _56319_;
wire _56320_;
wire _56321_;
wire _56322_;
wire _56323_;
wire _56324_;
wire _56325_;
wire _56326_;
wire _56327_;
wire _56328_;
wire _56329_;
wire _56330_;
wire _56331_;
wire _56332_;
wire _56333_;
wire _56334_;
wire _56335_;
wire _56336_;
wire _56337_;
wire _56338_;
wire _56339_;
wire _56340_;
wire _56341_;
wire _56342_;
wire _56343_;
wire _56344_;
wire _56345_;
wire _56346_;
wire _56347_;
wire _56348_;
wire _56349_;
wire _56350_;
wire _56351_;
wire _56352_;
wire _56353_;
wire _56354_;
wire _56355_;
wire _56356_;
wire _56357_;
wire _56358_;
wire _56359_;
wire _56360_;
wire _56361_;
wire _56362_;
wire _56363_;
wire _56364_;
wire _56365_;
wire _56366_;
wire _56367_;
wire _56368_;
wire _56369_;
wire _56370_;
wire _56371_;
wire _56372_;
wire _56373_;
wire _56374_;
wire _56375_;
wire _56376_;
wire _56377_;
wire _56378_;
wire _56379_;
wire _56380_;
wire _56381_;
wire _56382_;
wire _56383_;
wire _56384_;
wire _56385_;
wire _56386_;
wire _56387_;
wire _56388_;
wire _56389_;
wire _56390_;
wire _56391_;
wire _56392_;
wire _56393_;
wire _56394_;
wire _56395_;
wire _56396_;
wire _56397_;
wire _56398_;
wire _56399_;
wire _56400_;
wire _56401_;
wire _56402_;
wire _56403_;
wire _56404_;
wire _56405_;
wire _56406_;
wire _56407_;
wire _56408_;
wire _56409_;
wire _56410_;
wire _56411_;
wire _56412_;
wire _56413_;
wire _56414_;
wire _56415_;
wire _56416_;
wire _56417_;
wire _56418_;
wire _56419_;
wire _56420_;
wire _56421_;
wire _56422_;
wire _56423_;
wire _56424_;
wire _56425_;
wire _56426_;
wire _56427_;
wire _56428_;
wire _56429_;
wire _56430_;
wire _56431_;
wire _56432_;
wire _56433_;
wire _56434_;
wire _56435_;
wire _56436_;
wire _56437_;
wire _56438_;
wire _56439_;
wire _56440_;
wire _56441_;
wire _56442_;
wire _56443_;
wire _56444_;
wire _56445_;
wire _56446_;
wire _56447_;
wire _56448_;
wire _56449_;
wire _56450_;
wire _56451_;
wire _56452_;
wire _56453_;
wire _56454_;
wire _56455_;
wire _56456_;
wire _56457_;
wire _56458_;
wire _56459_;
wire _56460_;
wire _56461_;
wire _56462_;
wire _56463_;
wire _56464_;
wire _56465_;
wire _56466_;
wire _56467_;
wire _56468_;
wire _56469_;
wire _56470_;
wire _56471_;
wire _56472_;
wire _56473_;
wire _56474_;
wire _56475_;
wire _56476_;
wire _56477_;
wire _56478_;
wire _56479_;
wire _56480_;
wire _56481_;
wire _56482_;
wire _56483_;
wire _56484_;
wire _56485_;
wire _56486_;
wire _56487_;
wire _56488_;
wire _56489_;
wire _56490_;
wire _56491_;
wire _56492_;
wire _56493_;
wire _56494_;
wire _56495_;
wire _56496_;
wire _56497_;
wire _56498_;
wire _56499_;
wire _56500_;
wire _56501_;
wire _56502_;
wire _56503_;
wire _56504_;
wire _56505_;
wire _56506_;
wire _56507_;
wire _56508_;
wire _56509_;
wire _56510_;
wire _56511_;
wire _56512_;
wire _56513_;
wire _56514_;
wire _56515_;
wire _56516_;
wire _56517_;
wire _56518_;
wire _56519_;
wire _56520_;
wire _56521_;
wire _56522_;
wire _56523_;
wire _56524_;
wire _56525_;
wire _56526_;
wire _56527_;
wire _56528_;
wire _56529_;
wire _56530_;
wire _56531_;
wire _56532_;
wire _56533_;
wire _56534_;
wire _56535_;
wire _56536_;
wire _56537_;
wire _56538_;
wire _56539_;
wire _56540_;
wire _56541_;
wire _56542_;
wire _56543_;
wire _56544_;
wire _56545_;
wire _56546_;
wire _56547_;
wire _56548_;
wire _56549_;
wire _56550_;
wire _56551_;
wire _56552_;
wire _56553_;
wire _56554_;
wire _56555_;
wire _56556_;
wire _56557_;
wire _56558_;
wire _56559_;
wire _56560_;
wire _56561_;
wire _56562_;
wire _56563_;
wire _56564_;
wire _56565_;
wire _56566_;
wire _56567_;
wire _56568_;
wire _56569_;
wire _56570_;
wire _56571_;
wire _56572_;
wire _56573_;
wire _56574_;
wire _56575_;
wire _56576_;
wire _56577_;
wire _56578_;
wire _56579_;
wire _56580_;
wire _56581_;
wire _56582_;
wire _56583_;
wire _56584_;
wire _56585_;
wire _56586_;
wire _56587_;
wire _56588_;
wire _56589_;
wire _56590_;
wire _56591_;
wire _56592_;
wire _56593_;
wire _56594_;
wire _56595_;
wire _56596_;
wire _56597_;
wire _56598_;
wire _56599_;
wire _56600_;
wire _56601_;
wire _56602_;
wire _56603_;
wire _56604_;
wire _56605_;
wire _56606_;
wire _56607_;
wire _56608_;
wire _56609_;
wire _56610_;
wire _56611_;
wire _56612_;
wire _56613_;
wire _56614_;
wire _56615_;
wire _56616_;
wire _56617_;
wire _56618_;
wire _56619_;
wire _56620_;
wire _56621_;
wire _56622_;
wire _56623_;
wire _56624_;
wire _56625_;
wire _56626_;
wire _56627_;
wire _56628_;
wire _56629_;
wire _56630_;
wire _56631_;
wire _56632_;
wire _56633_;
wire _56634_;
wire _56635_;
wire _56636_;
wire _56637_;
wire _56638_;
wire _56639_;
wire _56640_;
wire _56641_;
wire _56642_;
wire _56643_;
wire _56644_;
wire _56645_;
wire _56646_;
wire _56647_;
wire _56648_;
wire _56649_;
wire _56650_;
wire _56651_;
wire _56652_;
wire _56653_;
wire _56654_;
wire _56655_;
wire _56656_;
wire _56657_;
wire _56658_;
wire _56659_;
wire _56660_;
wire _56661_;
wire _56662_;
wire _56663_;
wire _56664_;
wire _56665_;
wire _56666_;
wire _56667_;
wire _56668_;
wire _56669_;
wire _56670_;
wire _56671_;
wire _56672_;
wire _56673_;
wire _56674_;
wire _56675_;
wire _56676_;
wire _56677_;
wire _56678_;
wire _56679_;
wire _56680_;
wire _56681_;
wire _56682_;
wire _56683_;
wire _56684_;
wire _56685_;
wire _56686_;
wire _56687_;
wire _56688_;
wire _56689_;
wire _56690_;
wire _56691_;
wire _56692_;
wire _56693_;
wire _56694_;
wire _56695_;
wire _56696_;
wire _56697_;
wire _56698_;
wire _56699_;
wire _56700_;
wire _56701_;
wire _56702_;
wire _56703_;
wire _56704_;
wire _56705_;
wire _56706_;
wire _56707_;
wire _56708_;
wire _56709_;
wire _56710_;
wire _56711_;
wire _56712_;
wire _56713_;
wire _56714_;
wire _56715_;
wire _56716_;
wire _56717_;
wire _56718_;
wire _56719_;
wire _56720_;
wire _56721_;
wire _56722_;
wire _56723_;
wire _56724_;
wire _56725_;
wire _56726_;
wire _56727_;
wire _56728_;
wire _56729_;
wire _56730_;
wire _56731_;
wire _56732_;
wire _56733_;
wire _56734_;
wire _56735_;
wire _56736_;
wire _56737_;
wire _56738_;
wire _56739_;
wire _56740_;
wire _56741_;
wire _56742_;
wire _56743_;
wire _56744_;
wire _56745_;
wire _56746_;
wire _56747_;
wire _56748_;
wire _56749_;
wire _56750_;
wire _56751_;
wire _56752_;
wire _56753_;
wire _56754_;
wire _56755_;
wire _56756_;
wire _56757_;
wire _56758_;
wire _56759_;
wire _56760_;
wire _56761_;
wire _56762_;
wire _56763_;
wire _56764_;
wire _56765_;
wire _56766_;
wire _56767_;
wire _56768_;
wire _56769_;
wire _56770_;
wire _56771_;
wire _56772_;
wire _56773_;
wire _56774_;
wire _56775_;
wire _56776_;
wire _56777_;
wire _56778_;
wire _56779_;
wire _56780_;
wire _56781_;
wire _56782_;
wire _56783_;
wire _56784_;
wire _56785_;
wire _56786_;
wire _56787_;
wire _56788_;
wire _56789_;
wire _56790_;
wire _56791_;
wire _56792_;
wire _56793_;
wire _56794_;
wire _56795_;
wire _56796_;
wire _56797_;
wire _56798_;
wire _56799_;
wire _56800_;
wire _56801_;
wire _56802_;
wire _56803_;
wire _56804_;
wire _56805_;
wire _56806_;
wire _56807_;
wire _56808_;
wire _56809_;
wire _56810_;
wire _56811_;
wire _56812_;
wire _56813_;
wire _56814_;
wire _56815_;
wire _56816_;
wire _56817_;
wire _56818_;
wire _56819_;
wire _56820_;
wire _56821_;
wire _56822_;
wire _56823_;
wire _56824_;
wire _56825_;
wire _56826_;
wire _56827_;
wire _56828_;
wire _56829_;
wire _56830_;
wire _56831_;
wire _56832_;
wire _56833_;
wire _56834_;
wire _56835_;
wire _56836_;
wire _56837_;
wire _56838_;
wire _56839_;
wire _56840_;
wire _56841_;
wire _56842_;
wire _56843_;
wire _56844_;
wire _56845_;
wire _56846_;
wire _56847_;
wire _56848_;
wire _56849_;
wire _56850_;
wire _56851_;
wire _56852_;
wire _56853_;
wire _56854_;
wire _56855_;
wire _56856_;
wire _56857_;
wire _56858_;
wire _56859_;
wire _56860_;
wire _56861_;
wire _56862_;
wire _56863_;
wire _56864_;
wire _56865_;
wire _56866_;
wire _56867_;
wire _56868_;
wire _56869_;
wire _56870_;
wire _56871_;
wire _56872_;
wire _56873_;
wire _56874_;
wire _56875_;
wire _56876_;
wire _56877_;
wire _56878_;
wire _56879_;
wire _56880_;
wire _56881_;
wire _56882_;
wire _56883_;
wire _56884_;
wire _56885_;
wire _56886_;
wire _56887_;
wire _56888_;
wire _56889_;
wire _56890_;
wire _56891_;
wire _56892_;
wire _56893_;
wire _56894_;
wire _56895_;
wire _56896_;
wire _56897_;
wire _56898_;
wire _56899_;
wire _56900_;
wire _56901_;
wire _56902_;
wire _56903_;
wire _56904_;
wire _56905_;
wire _56906_;
wire _56907_;
wire _56908_;
wire _56909_;
wire _56910_;
wire _56911_;
wire _56912_;
wire _56913_;
wire _56914_;
wire _56915_;
wire _56916_;
wire _56917_;
wire _56918_;
wire _56919_;
wire _56920_;
wire _56921_;
wire _56922_;
wire _56923_;
wire _56924_;
wire _56925_;
wire _56926_;
wire _56927_;
wire _56928_;
wire _56929_;
wire _56930_;
wire _56931_;
wire _56932_;
wire _56933_;
wire _56934_;
wire _56935_;
wire _56936_;
wire _56937_;
wire _56938_;
wire _56939_;
wire _56940_;
wire _56941_;
wire _56942_;
wire _56943_;
wire _56944_;
wire _56945_;
wire _56946_;
wire _56947_;
wire _56948_;
wire _56949_;
wire _56950_;
wire _56951_;
wire _56952_;
wire _56953_;
wire _56954_;
wire _56955_;
wire _56956_;
wire _56957_;
wire _56958_;
wire _56959_;
wire _56960_;
wire _56961_;
wire _56962_;
wire _56963_;
wire _56964_;
wire _56965_;
wire _56966_;
wire _56967_;
wire _56968_;
wire _56969_;
wire _56970_;
wire _56971_;
wire _56972_;
wire _56973_;
wire _56974_;
wire _56975_;
wire _56976_;
wire _56977_;
wire _56978_;
wire _56979_;
wire _56980_;
wire _56981_;
wire _56982_;
wire _56983_;
wire _56984_;
wire _56985_;
wire _56986_;
wire _56987_;
wire _56988_;
wire _56989_;
wire _56990_;
wire _56991_;
wire _56992_;
wire _56993_;
wire _56994_;
wire _56995_;
wire _56996_;
wire _56997_;
wire _56998_;
wire _56999_;
wire _57000_;
wire _57001_;
wire _57002_;
wire _57003_;
wire _57004_;
wire _57005_;
wire _57006_;
wire _57007_;
wire _57008_;
wire _57009_;
wire _57010_;
wire _57011_;
wire _57012_;
wire _57013_;
wire _57014_;
wire _57015_;
wire _57016_;
wire _57017_;
wire _57018_;
wire _57019_;
wire _57020_;
wire _57021_;
wire _57022_;
wire _57023_;
wire _57024_;
wire _57025_;
wire _57026_;
wire _57027_;
wire _57028_;
wire _57029_;
wire _57030_;
wire _57031_;
wire _57032_;
wire _57033_;
wire _57034_;
wire _57035_;
wire _57036_;
wire _57037_;
wire _57038_;
wire _57039_;
wire _57040_;
wire _57041_;
wire _57042_;
wire _57043_;
wire _57044_;
wire _57045_;
wire _57046_;
wire _57047_;
wire _57048_;
wire _57049_;
wire _57050_;
wire _57051_;
wire _57052_;
wire _57053_;
wire _57054_;
wire _57055_;
wire _57056_;
wire _57057_;
wire _57058_;
wire _57059_;
wire _57060_;
wire _57061_;
wire _57062_;
wire _57063_;
wire _57064_;
wire _57065_;
wire _57066_;
wire _57067_;
wire _57068_;
wire _57069_;
wire _57070_;
wire _57071_;
wire _57072_;
wire _57073_;
wire _57074_;
wire _57075_;
wire _57076_;
wire _57077_;
wire _57078_;
wire _57079_;
wire _57080_;
wire _57081_;
wire _57082_;
wire _57083_;
wire _57084_;
wire _57085_;
wire _57086_;
wire _57087_;
wire _57088_;
wire _57089_;
wire _57090_;
wire _57091_;
wire _57092_;
wire _57093_;
wire _57094_;
wire _57095_;
wire _57096_;
wire _57097_;
wire _57098_;
wire _57099_;
wire _57100_;
wire _57101_;
wire _57102_;
wire _57103_;
wire _57104_;
wire _57105_;
wire _57106_;
wire _57107_;
wire _57108_;
wire _57109_;
wire _57110_;
wire _57111_;
wire _57112_;
wire _57113_;
wire _57114_;
wire _57115_;
wire _57116_;
wire _57117_;
wire _57118_;
wire _57119_;
wire _57120_;
wire _57121_;
wire _57122_;
wire _57123_;
wire _57124_;
wire _57125_;
wire _57126_;
wire _57127_;
wire _57128_;
wire _57129_;
wire _57130_;
wire _57131_;
wire _57132_;
wire _57133_;
wire _57134_;
wire _57135_;
wire _57136_;
wire _57137_;
wire _57138_;
wire _57139_;
wire _57140_;
wire _57141_;
wire _57142_;
wire _57143_;
wire _57144_;
wire _57145_;
wire _57146_;
wire _57147_;
wire _57148_;
wire _57149_;
wire _57150_;
wire _57151_;
wire _57152_;
wire _57153_;
wire _57154_;
wire _57155_;
wire _57156_;
wire _57157_;
wire _57158_;
wire _57159_;
wire _57160_;
wire _57161_;
wire _57162_;
wire _57163_;
wire _57164_;
wire _57165_;
wire _57166_;
wire _57167_;
wire _57168_;
wire _57169_;
wire _57170_;
wire _57171_;
wire _57172_;
wire _57173_;
wire _57174_;
wire _57175_;
wire _57176_;
wire _57177_;
wire _57178_;
wire _57179_;
wire _57180_;
wire _57181_;
wire _57182_;
wire _57183_;
wire _57184_;
wire _57185_;
wire _57186_;
wire _57187_;
wire _57188_;
wire _57189_;
wire _57190_;
wire _57191_;
wire _57192_;
wire _57193_;
wire _57194_;
wire _57195_;
wire _57196_;
wire _57197_;
wire _57198_;
wire _57199_;
wire _57200_;
wire _57201_;
wire _57202_;
wire _57203_;
wire _57204_;
wire _57205_;
wire _57206_;
wire _57207_;
wire _57208_;
wire _57209_;
wire _57210_;
wire _57211_;
wire _57212_;
wire _57213_;
wire _57214_;
wire _57215_;
wire _57216_;
wire _57217_;
wire _57218_;
wire _57219_;
wire _57220_;
wire _57221_;
wire _57222_;
wire _57223_;
wire _57224_;
wire _57225_;
wire _57226_;
wire _57227_;
wire _57228_;
wire _57229_;
wire _57230_;
wire _57231_;
wire _57232_;
wire _57233_;
wire _57234_;
wire _57235_;
wire _57236_;
wire _57237_;
wire _57238_;
wire _57239_;
wire _57240_;
wire _57241_;
wire _57242_;
wire _57243_;
wire _57244_;
wire _57245_;
wire _57246_;
wire _57247_;
wire _57248_;
wire _57249_;
wire _57250_;
wire _57251_;
wire _57252_;
wire _57253_;
wire _57254_;
wire _57255_;
wire _57256_;
wire _57257_;
wire _57258_;
wire _57259_;
wire _57260_;
wire _57261_;
wire _57262_;
wire _57263_;
wire _57264_;
wire _57265_;
wire _57266_;
wire _57267_;
wire _57268_;
wire _57269_;
wire _57270_;
wire _57271_;
wire _57272_;
wire _57273_;
wire _57274_;
wire _57275_;
wire _57276_;
wire _57277_;
wire _57278_;
wire _57279_;
wire _57280_;
wire _57281_;
wire _57282_;
wire _57283_;
wire _57284_;
wire _57285_;
wire _57286_;
wire _57287_;
wire _57288_;
wire _57289_;
wire _57290_;
wire _57291_;
wire _57292_;
wire _57293_;
wire _57294_;
wire _57295_;
wire _57296_;
wire _57297_;
wire _57298_;
wire _57299_;
wire _57300_;
wire _57301_;
wire _57302_;
wire _57303_;
wire _57304_;
wire _57305_;
wire _57306_;
wire _57307_;
wire _57308_;
wire _57309_;
wire _57310_;
wire _57311_;
wire _57312_;
wire _57313_;
wire _57314_;
wire _57315_;
wire _57316_;
wire _57317_;
wire _57318_;
wire _57319_;
wire _57320_;
wire _57321_;
wire _57322_;
wire _57323_;
wire _57324_;
wire _57325_;
wire _57326_;
wire _57327_;
wire _57328_;
wire _57329_;
wire _57330_;
wire _57331_;
wire _57332_;
wire _57333_;
wire _57334_;
wire _57335_;
wire _57336_;
wire _57337_;
wire _57338_;
wire _57339_;
wire _57340_;
wire _57341_;
wire _57342_;
wire _57343_;
wire _57344_;
wire _57345_;
wire _57346_;
wire _57347_;
wire _57348_;
wire _57349_;
wire _57350_;
wire _57351_;
wire _57352_;
wire _57353_;
wire _57354_;
wire _57355_;
wire _57356_;
wire _57357_;
wire _57358_;
wire _57359_;
wire _57360_;
wire _57361_;
wire _57362_;
wire _57363_;
wire _57364_;
wire _57365_;
wire _57366_;
wire _57367_;
wire _57368_;
wire _57369_;
wire _57370_;
wire _57371_;
wire _57372_;
wire _57373_;
wire _57374_;
wire _57375_;
wire _57376_;
wire _57377_;
wire _57378_;
wire _57379_;
wire _57380_;
wire _57381_;
wire _57382_;
wire _57383_;
wire _57384_;
wire _57385_;
wire _57386_;
wire _57387_;
wire _57388_;
wire _57389_;
wire _57390_;
wire _57391_;
wire _57392_;
wire _57393_;
wire _57394_;
wire _57395_;
wire _57396_;
wire _57397_;
wire _57398_;
wire _57399_;
wire _57400_;
wire _57401_;
wire _57402_;
wire _57403_;
wire _57404_;
wire _57405_;
wire _57406_;
wire _57407_;
wire _57408_;
wire _57409_;
wire _57410_;
wire _57411_;
wire _57412_;
wire _57413_;
wire _57414_;
wire _57415_;
wire _57416_;
wire _57417_;
wire _57418_;
wire _57419_;
wire _57420_;
wire _57421_;
wire _57422_;
wire _57423_;
wire _57424_;
wire _57425_;
wire _57426_;
wire _57427_;
wire _57428_;
wire _57429_;
wire _57430_;
wire _57431_;
wire _57432_;
wire _57433_;
wire _57434_;
wire _57435_;
wire _57436_;
wire _57437_;
wire _57438_;
wire _57439_;
wire _57440_;
wire _57441_;
wire _57442_;
wire _57443_;
wire _57444_;
wire _57445_;
wire _57446_;
wire _57447_;
wire _57448_;
wire _57449_;
wire _57450_;
wire _57451_;
wire _57452_;
wire _57453_;
wire _57454_;
wire _57455_;
wire _57456_;
wire _57457_;
wire _57458_;
wire _57459_;
wire _57460_;
wire _57461_;
wire _57462_;
wire _57463_;
wire _57464_;
wire _57465_;
wire _57466_;
wire _57467_;
wire _57468_;
wire _57469_;
wire _57470_;
wire _57471_;
wire _57472_;
wire _57473_;
wire _57474_;
wire _57475_;
wire _57476_;
wire _57477_;
wire _57478_;
wire _57479_;
wire _57480_;
wire _57481_;
wire _57482_;
wire _57483_;
wire _57484_;
wire _57485_;
wire _57486_;
wire _57487_;
wire _57488_;
wire _57489_;
wire _57490_;
wire _57491_;
wire _57492_;
wire _57493_;
wire _57494_;
wire _57495_;
wire _57496_;
wire _57497_;
wire _57498_;
wire _57499_;
wire _57500_;
wire _57501_;
wire _57502_;
wire _57503_;
wire _57504_;
wire _57505_;
wire _57506_;
wire _57507_;
wire _57508_;
wire _57509_;
wire _57510_;
wire _57511_;
wire _57512_;
wire _57513_;
wire _57514_;
wire _57515_;
wire _57516_;
wire _57517_;
wire _57518_;
wire _57519_;
wire _57520_;
wire _57521_;
wire _57522_;
wire _57523_;
wire _57524_;
wire _57525_;
wire _57526_;
wire _57527_;
wire _57528_;
wire _57529_;
wire _57530_;
wire _57531_;
wire _57532_;
wire _57533_;
wire _57534_;
wire _57535_;
wire _57536_;
wire _57537_;
wire _57538_;
wire _57539_;
wire _57540_;
wire _57541_;
wire _57542_;
wire _57543_;
wire _57544_;
wire _57545_;
wire _57546_;
wire _57547_;
wire _57548_;
wire _57549_;
wire _57550_;
wire _57551_;
wire _57552_;
wire _57553_;
wire _57554_;
wire _57555_;
wire _57556_;
wire _57557_;
wire _57558_;
wire _57559_;
wire _57560_;
wire _57561_;
wire _57562_;
wire _57563_;
wire _57564_;
wire _57565_;
wire _57566_;
wire _57567_;
wire _57568_;
wire _57569_;
wire _57570_;
wire _57571_;
wire _57572_;
wire _57573_;
wire _57574_;
wire _57575_;
wire _57576_;
wire _57577_;
wire _57578_;
wire _57579_;
wire _57580_;
wire _57581_;
wire _57582_;
wire _57583_;
wire _57584_;
wire _57585_;
wire _57586_;
wire _57587_;
wire _57588_;
wire _57589_;
wire _57590_;
wire _57591_;
wire _57592_;
wire _57593_;
wire _57594_;
wire _57595_;
wire _57596_;
wire _57597_;
wire _57598_;
wire _57599_;
wire _57600_;
wire _57601_;
wire _57602_;
wire _57603_;
wire _57604_;
wire _57605_;
wire _57606_;
wire _57607_;
wire _57608_;
wire _57609_;
wire _57610_;
wire _57611_;
wire _57612_;
wire _57613_;
wire _57614_;
wire _57615_;
wire _57616_;
wire _57617_;
wire _57618_;
wire _57619_;
wire _57620_;
wire _57621_;
wire _57622_;
wire _57623_;
wire _57624_;
wire _57625_;
wire _57626_;
wire _57627_;
wire _57628_;
wire _57629_;
wire _57630_;
wire _57631_;
wire _57632_;
wire _57633_;
wire _57634_;
wire _57635_;
wire _57636_;
wire _57637_;
wire _57638_;
wire _57639_;
wire _57640_;
wire _57641_;
wire _57642_;
wire _57643_;
wire _57644_;
wire _57645_;
wire _57646_;
wire _57647_;
wire _57648_;
wire _57649_;
wire _57650_;
wire _57651_;
wire _57652_;
wire _57653_;
wire _57654_;
wire _57655_;
wire _57656_;
wire _57657_;
wire _57658_;
wire _57659_;
wire _57660_;
wire _57661_;
wire _57662_;
wire _57663_;
wire _57664_;
wire _57665_;
wire _57666_;
wire _57667_;
wire _57668_;
wire _57669_;
wire _57670_;
wire _57671_;
wire _57672_;
wire _57673_;
wire _57674_;
wire _57675_;
wire _57676_;
wire _57677_;
wire _57678_;
wire _57679_;
wire _57680_;
wire _57681_;
wire _57682_;
wire _57683_;
wire _57684_;
wire _57685_;
wire _57686_;
wire _57687_;
wire _57688_;
wire _57689_;
wire _57690_;
wire _57691_;
wire _57692_;
wire _57693_;
wire _57694_;
wire _57695_;
wire _57696_;
wire _57697_;
wire _57698_;
wire _57699_;
wire _57700_;
wire _57701_;
wire _57702_;
wire _57703_;
wire _57704_;
wire _57705_;
wire _57706_;
wire _57707_;
wire _57708_;
wire _57709_;
wire _57710_;
wire _57711_;
wire _57712_;
wire _57713_;
wire _57714_;
wire _57715_;
wire _57716_;
wire _57717_;
wire _57718_;
wire _57719_;
wire _57720_;
wire _57721_;
wire _57722_;
wire _57723_;
wire _57724_;
wire _57725_;
wire _57726_;
wire _57727_;
wire _57728_;
wire _57729_;
wire _57730_;
wire _57731_;
wire _57732_;
wire _57733_;
wire _57734_;
wire _57735_;
wire _57736_;
wire _57737_;
wire _57738_;
wire _57739_;
wire _57740_;
wire _57741_;
wire _57742_;
wire _57743_;
wire _57744_;
wire _57745_;
wire _57746_;
wire _57747_;
wire _57748_;
wire _57749_;
wire _57750_;
wire _57751_;
wire _57752_;
wire _57753_;
wire _57754_;
wire _57755_;
wire _57756_;
wire _57757_;
wire _57758_;
wire _57759_;
wire _57760_;
wire _57761_;
wire _57762_;
wire _57763_;
wire _57764_;
wire _57765_;
wire _57766_;
wire _57767_;
wire _57768_;
wire _57769_;
wire _57770_;
wire _57771_;
wire _57772_;
wire _57773_;
wire _57774_;
wire _57775_;
wire _57776_;
wire _57777_;
wire _57778_;
wire _57779_;
wire _57780_;
wire _57781_;
wire _57782_;
wire _57783_;
wire _57784_;
wire _57785_;
wire _57786_;
wire _57787_;
wire _57788_;
wire _57789_;
wire _57790_;
wire _57791_;
wire _57792_;
wire _57793_;
wire _57794_;
wire _57795_;
wire _57796_;
wire _57797_;
wire _57798_;
wire _57799_;
wire _57800_;
wire _57801_;
wire _57802_;
wire _57803_;
wire _57804_;
wire _57805_;
wire _57806_;
wire _57807_;
wire _57808_;
wire _57809_;
wire _57810_;
wire _57811_;
wire _57812_;
wire _57813_;
wire _57814_;
wire _57815_;
wire _57816_;
wire _57817_;
wire _57818_;
wire _57819_;
wire _57820_;
wire _57821_;
wire _57822_;
wire _57823_;
wire _57824_;
wire _57825_;
wire _57826_;
wire _57827_;
wire _57828_;
wire _57829_;
wire _57830_;
wire _57831_;
wire _57832_;
wire _57833_;
wire _57834_;
wire _57835_;
wire _57836_;
wire _57837_;
wire _57838_;
wire _57839_;
wire _57840_;
wire _57841_;
wire _57842_;
wire _57843_;
wire _57844_;
wire _57845_;
wire _57846_;
wire _57847_;
wire _57848_;
wire _57849_;
wire _57850_;
wire _57851_;
wire _57852_;
wire _57853_;
wire _57854_;
wire _57855_;
wire _57856_;
wire _57857_;
wire _57858_;
wire _57859_;
wire _57860_;
wire _57861_;
wire _57862_;
wire _57863_;
wire _57864_;
wire _57865_;
wire _57866_;
wire _57867_;
wire _57868_;
wire _57869_;
wire _57870_;
wire _57871_;
wire _57872_;
wire _57873_;
wire _57874_;
wire _57875_;
wire _57876_;
wire _57877_;
wire _57878_;
wire _57879_;
wire _57880_;
wire _57881_;
wire _57882_;
wire _57883_;
wire _57884_;
wire _57885_;
wire _57886_;
wire _57887_;
wire _57888_;
wire _57889_;
wire _57890_;
wire _57891_;
wire _57892_;
wire _57893_;
wire _57894_;
wire _57895_;
wire _57896_;
wire _57897_;
wire _57898_;
wire _57899_;
wire _57900_;
wire _57901_;
wire _57902_;
wire _57903_;
wire _57904_;
wire _57905_;
wire _57906_;
wire _57907_;
wire _57908_;
wire _57909_;
wire _57910_;
wire _57911_;
wire _57912_;
wire _57913_;
wire _57914_;
wire _57915_;
wire _57916_;
wire _57917_;
wire _57918_;
wire _57919_;
wire _57920_;
wire _57921_;
wire _57922_;
wire _57923_;
wire _57924_;
wire _57925_;
wire _57926_;
wire _57927_;
wire _57928_;
wire _57929_;
wire _57930_;
wire _57931_;
wire _57932_;
wire _57933_;
wire _57934_;
wire _57935_;
wire _57936_;
wire _57937_;
wire _57938_;
wire _57939_;
wire _57940_;
wire _57941_;
wire _57942_;
wire _57943_;
wire _57944_;
wire _57945_;
wire _57946_;
wire _57947_;
wire _57948_;
wire _57949_;
wire _57950_;
wire _57951_;
wire _57952_;
wire _57953_;
wire _57954_;
wire _57955_;
wire _57956_;
wire _57957_;
wire _57958_;
wire _57959_;
wire _57960_;
wire _57961_;
wire _57962_;
wire _57963_;
wire _57964_;
wire _57965_;
wire _57966_;
wire _57967_;
wire _57968_;
wire _57969_;
wire _57970_;
wire _57971_;
wire _57972_;
wire _57973_;
wire _57974_;
wire _57975_;
wire _57976_;
wire _57977_;
wire _57978_;
wire _57979_;
wire _57980_;
wire _57981_;
wire _57982_;
wire _57983_;
wire _57984_;
wire _57985_;
wire _57986_;
wire _57987_;
wire _57988_;
wire _57989_;
wire _57990_;
wire _57991_;
wire _57992_;
wire _57993_;
wire _57994_;
wire _57995_;
wire _57996_;
wire _57997_;
wire _57998_;
wire _57999_;
wire _58000_;
wire _58001_;
wire _58002_;
wire _58003_;
wire _58004_;
wire _58005_;
wire _58006_;
wire _58007_;
wire _58008_;
wire _58009_;
wire _58010_;
wire _58011_;
wire _58012_;
wire _58013_;
wire _58014_;
wire _58015_;
wire _58016_;
wire _58017_;
wire _58018_;
wire _58019_;
wire _58020_;
wire _58021_;
wire _58022_;
wire _58023_;
wire _58024_;
wire _58025_;
wire _58026_;
wire _58027_;
wire _58028_;
wire _58029_;
wire _58030_;
wire _58031_;
wire _58032_;
wire _58033_;
wire _58034_;
wire _58035_;
wire _58036_;
wire _58037_;
wire _58038_;
wire _58039_;
wire _58040_;
wire _58041_;
wire _58042_;
wire _58043_;
wire _58044_;
wire _58045_;
wire _58046_;
wire _58047_;
wire _58048_;
wire _58049_;
wire _58050_;
wire _58051_;
wire _58052_;
wire _58053_;
wire _58054_;
wire _58055_;
wire _58056_;
wire _58057_;
wire _58058_;
wire _58059_;
wire _58060_;
wire _58061_;
wire _58062_;
wire _58063_;
wire _58064_;
wire _58065_;
wire _58066_;
wire _58067_;
wire _58068_;
wire _58069_;
wire _58070_;
wire _58071_;
wire _58072_;
wire _58073_;
wire _58074_;
wire _58075_;
wire _58076_;
wire _58077_;
wire _58078_;
wire _58079_;
wire _58080_;
wire _58081_;
wire _58082_;
wire _58083_;
wire _58084_;
wire _58085_;
wire _58086_;
wire _58087_;
wire _58088_;
wire _58089_;
wire _58090_;
wire _58091_;
wire _58092_;
wire _58093_;
wire _58094_;
wire _58095_;
wire _58096_;
wire _58097_;
wire _58098_;
wire _58099_;
wire _58100_;
wire _58101_;
wire _58102_;
wire _58103_;
wire _58104_;
wire _58105_;
wire _58106_;
wire _58107_;
wire _58108_;
wire _58109_;
wire _58110_;
wire _58111_;
wire _58112_;
wire _58113_;
wire _58114_;
wire _58115_;
wire _58116_;
wire _58117_;
wire _58118_;
wire _58119_;
wire _58120_;
wire _58121_;
wire _58122_;
wire _58123_;
wire _58124_;
wire _58125_;
wire _58126_;
wire _58127_;
wire _58128_;
wire _58129_;
wire _58130_;
wire _58131_;
wire _58132_;
wire _58133_;
wire _58134_;
wire _58135_;
wire _58136_;
wire _58137_;
wire _58138_;
wire _58139_;
wire _58140_;
wire _58141_;
wire _58142_;
wire _58143_;
wire _58144_;
wire _58145_;
wire _58146_;
wire _58147_;
wire _58148_;
wire _58149_;
wire _58150_;
wire _58151_;
wire _58152_;
wire _58153_;
wire _58154_;
wire _58155_;
wire _58156_;
wire _58157_;
wire _58158_;
wire _58159_;
wire _58160_;
wire _58161_;
wire _58162_;
wire _58163_;
wire _58164_;
wire _58165_;
wire _58166_;
wire _58167_;
wire _58168_;
wire _58169_;
wire _58170_;
wire _58171_;
wire _58172_;
wire _58173_;
wire _58174_;
wire _58175_;
wire _58176_;
wire _58177_;
wire _58178_;
wire _58179_;
wire _58180_;
wire _58181_;
wire _58182_;
wire _58183_;
wire _58184_;
wire _58185_;
wire _58186_;
wire _58187_;
wire _58188_;
wire _58189_;
wire _58190_;
wire _58191_;
wire _58192_;
wire _58193_;
wire _58194_;
wire _58195_;
wire _58196_;
wire _58197_;
wire _58198_;
wire _58199_;
wire _58200_;
wire _58201_;
wire _58202_;
wire _58203_;
wire _58204_;
wire _58205_;
wire _58206_;
wire _58207_;
wire _58208_;
wire _58209_;
wire _58210_;
wire _58211_;
wire _58212_;
wire _58213_;
wire _58214_;
wire _58215_;
wire _58216_;
wire _58217_;
wire _58218_;
wire _58219_;
wire _58220_;
wire _58221_;
wire _58222_;
wire _58223_;
wire _58224_;
wire _58225_;
wire _58226_;
wire _58227_;
wire _58228_;
wire _58229_;
wire _58230_;
wire _58231_;
wire _58232_;
wire _58233_;
wire _58234_;
wire _58235_;
wire _58236_;
wire _58237_;
wire _58238_;
wire _58239_;
wire _58240_;
wire _58241_;
wire _58242_;
wire _58243_;
wire _58244_;
wire _58245_;
wire _58246_;
wire _58247_;
wire _58248_;
wire _58249_;
wire _58250_;
wire _58251_;
wire _58252_;
wire _58253_;
wire _58254_;
wire _58255_;
wire _58256_;
wire _58257_;
wire _58258_;
wire _58259_;
wire _58260_;
wire _58261_;
wire _58262_;
wire _58263_;
wire _58264_;
wire _58265_;
wire _58266_;
wire _58267_;
wire _58268_;
wire _58269_;
wire _58270_;
wire _58271_;
wire _58272_;
wire _58273_;
wire _58274_;
wire _58275_;
wire _58276_;
wire _58277_;
wire _58278_;
wire _58279_;
wire _58280_;
wire _58281_;
wire _58282_;
wire _58283_;
wire _58284_;
wire _58285_;
wire _58286_;
wire _58287_;
wire _58288_;
wire _58289_;
wire _58290_;
wire _58291_;
wire _58292_;
wire _58293_;
wire _58294_;
wire _58295_;
wire _58296_;
wire _58297_;
wire _58298_;
wire _58299_;
wire _58300_;
wire _58301_;
wire _58302_;
wire _58303_;
wire _58304_;
wire _58305_;
wire _58306_;
wire _58307_;
wire _58308_;
wire _58309_;
wire _58310_;
wire _58311_;
wire _58312_;
wire _58313_;
wire _58314_;
wire _58315_;
wire _58316_;
wire _58317_;
wire _58318_;
wire _58319_;
wire _58320_;
wire _58321_;
wire _58322_;
wire _58323_;
wire _58324_;
wire _58325_;
wire _58326_;
wire _58327_;
wire _58328_;
wire _58329_;
wire _58330_;
wire _58331_;
wire _58332_;
wire _58333_;
wire _58334_;
wire _58335_;
wire _58336_;
wire _58337_;
wire _58338_;
wire _58339_;
wire _58340_;
wire _58341_;
wire _58342_;
wire _58343_;
wire _58344_;
wire _58345_;
wire _58346_;
wire _58347_;
wire _58348_;
wire _58349_;
wire _58350_;
wire _58351_;
wire _58352_;
wire _58353_;
wire _58354_;
wire _58355_;
wire _58356_;
wire _58357_;
wire _58358_;
wire _58359_;
wire _58360_;
wire _58361_;
wire _58362_;
wire _58363_;
wire _58364_;
wire _58365_;
wire _58366_;
wire _58367_;
wire _58368_;
wire _58369_;
wire _58370_;
wire _58371_;
wire _58372_;
wire _58373_;
wire _58374_;
wire _58375_;
wire _58376_;
wire _58377_;
wire _58378_;
wire _58379_;
wire _58380_;
wire _58381_;
wire _58382_;
wire _58383_;
wire _58384_;
wire _58385_;
wire _58386_;
wire _58387_;
wire _58388_;
wire _58389_;
wire _58390_;
wire _58391_;
wire _58392_;
wire _58393_;
wire _58394_;
wire _58395_;
wire _58396_;
wire _58397_;
wire _58398_;
wire _58399_;
wire _58400_;
wire _58401_;
wire _58402_;
wire _58403_;
wire _58404_;
wire _58405_;
wire _58406_;
wire _58407_;
wire _58408_;
wire _58409_;
wire _58410_;
wire _58411_;
wire _58412_;
wire _58413_;
wire _58414_;
wire _58415_;
wire _58416_;
wire _58417_;
wire _58418_;
wire _58419_;
wire _58420_;
wire _58421_;
wire _58422_;
wire _58423_;
wire _58424_;
wire _58425_;
wire _58426_;
wire _58427_;
wire _58428_;
wire _58429_;
wire _58430_;
wire _58431_;
wire _58432_;
wire _58433_;
wire _58434_;
wire _58435_;
wire _58436_;
wire _58437_;
wire _58438_;
wire _58439_;
wire _58440_;
wire _58441_;
wire _58442_;
wire _58443_;
wire _58444_;
wire _58445_;
wire _58446_;
wire _58447_;
wire _58448_;
wire _58449_;
wire _58450_;
wire _58451_;
wire _58452_;
wire _58453_;
wire _58454_;
wire _58455_;
wire _58456_;
wire _58457_;
wire _58458_;
wire _58459_;
wire _58460_;
wire _58461_;
wire _58462_;
wire _58463_;
wire _58464_;
wire _58465_;
wire _58466_;
wire _58467_;
wire _58468_;
wire _58469_;
wire _58470_;
wire _58471_;
wire _58472_;
wire _58473_;
wire _58474_;
wire _58475_;
wire _58476_;
wire _58477_;
wire _58478_;
wire _58479_;
wire _58480_;
wire _58481_;
wire _58482_;
wire _58483_;
wire _58484_;
wire _58485_;
wire _58486_;
wire _58487_;
wire _58488_;
wire _58489_;
wire _58490_;
wire _58491_;
wire _58492_;
wire _58493_;
wire _58494_;
wire _58495_;
wire _58496_;
wire _58497_;
wire _58498_;
wire _58499_;
wire _58500_;
wire _58501_;
wire _58502_;
wire _58503_;
wire _58504_;
wire _58505_;
wire _58506_;
wire _58507_;
wire _58508_;
wire _58509_;
wire _58510_;
wire _58511_;
wire _58512_;
wire _58513_;
wire _58514_;
wire _58515_;
wire _58516_;
wire _58517_;
wire _58518_;
wire _58519_;
wire _58520_;
wire _58521_;
wire _58522_;
wire _58523_;
wire _58524_;
wire _58525_;
wire _58526_;
wire _58527_;
wire _58528_;
wire _58529_;
wire _58530_;
wire _58531_;
wire _58532_;
wire _58533_;
wire _58534_;
wire _58535_;
wire _58536_;
wire _58537_;
wire _58538_;
wire _58539_;
wire _58540_;
wire _58541_;
wire _58542_;
wire _58543_;
wire _58544_;
wire _58545_;
wire _58546_;
wire _58547_;
wire _58548_;
wire _58549_;
wire _58550_;
wire _58551_;
wire _58552_;
wire _58553_;
wire _58554_;
wire _58555_;
wire _58556_;
wire _58557_;
wire _58558_;
wire _58559_;
wire _58560_;
wire _58561_;
wire _58562_;
wire _58563_;
wire _58564_;
wire _58565_;
wire _58566_;
wire _58567_;
wire _58568_;
wire _58569_;
wire _58570_;
wire _58571_;
wire _58572_;
wire _58573_;
wire _58574_;
wire _58575_;
wire _58576_;
wire _58577_;
wire _58578_;
wire _58579_;
wire _58580_;
wire _58581_;
wire _58582_;
wire _58583_;
wire _58584_;
wire _58585_;
wire _58586_;
wire _58587_;
wire _58588_;
wire _58589_;
wire _58590_;
wire _58591_;
wire _58592_;
wire _58593_;
wire _58594_;
wire _58595_;
wire _58596_;
wire _58597_;
wire _58598_;
wire _58599_;
wire _58600_;
wire _58601_;
wire _58602_;
wire _58603_;
wire _58604_;
wire _58605_;
wire _58606_;
wire _58607_;
wire _58608_;
wire _58609_;
wire _58610_;
wire _58611_;
wire _58612_;
wire _58613_;
wire _58614_;
wire _58615_;
wire _58616_;
wire _58617_;
wire _58618_;
wire _58619_;
wire _58620_;
wire _58621_;
wire _58622_;
wire _58623_;
wire _58624_;
wire _58625_;
wire _58626_;
wire _58627_;
wire _58628_;
wire _58629_;
wire _58630_;
wire _58631_;
wire _58632_;
wire _58633_;
wire _58634_;
wire _58635_;
wire _58636_;
wire _58637_;
wire _58638_;
wire _58639_;
wire _58640_;
wire _58641_;
wire _58642_;
wire _58643_;
wire _58644_;
wire _58645_;
wire _58646_;
wire _58647_;
wire _58648_;
wire _58649_;
wire _58650_;
wire _58651_;
wire _58652_;
wire _58653_;
wire _58654_;
wire _58655_;
wire _58656_;
wire _58657_;
wire _58658_;
wire _58659_;
wire _58660_;
wire _58661_;
wire _58662_;
wire _58663_;
wire _58664_;
wire _58665_;
wire _58666_;
wire _58667_;
wire _58668_;
wire _58669_;
wire _58670_;
wire _58671_;
wire _58672_;
wire _58673_;
wire _58674_;
wire _58675_;
wire _58676_;
wire _58677_;
wire _58678_;
wire _58679_;
wire _58680_;
wire _58681_;
wire _58682_;
wire _58683_;
wire _58684_;
wire _58685_;
wire _58686_;
wire _58687_;
wire _58688_;
wire _58689_;
wire _58690_;
wire _58691_;
wire _58692_;
wire _58693_;
wire _58694_;
wire _58695_;
wire _58696_;
wire _58697_;
wire _58698_;
wire _58699_;
wire _58700_;
wire _58701_;
wire _58702_;
wire _58703_;
wire _58704_;
wire _58705_;
wire _58706_;
wire _58707_;
wire _58708_;
wire _58709_;
wire _58710_;
wire _58711_;
wire _58712_;
wire _58713_;
wire _58714_;
wire _58715_;
wire _58716_;
wire _58717_;
wire _58718_;
wire _58719_;
wire _58720_;
wire _58721_;
wire _58722_;
wire _58723_;
wire _58724_;
wire _58725_;
wire _58726_;
wire _58727_;
wire _58728_;
wire _58729_;
wire _58730_;
wire _58731_;
wire _58732_;
wire _58733_;
wire _58734_;
wire _58735_;
wire _58736_;
wire _58737_;
wire _58738_;
wire _58739_;
wire _58740_;
wire _58741_;
wire _58742_;
wire _58743_;
wire _58744_;
wire _58745_;
wire _58746_;
wire _58747_;
wire _58748_;
wire _58749_;
wire _58750_;
wire _58751_;
wire _58752_;
wire _58753_;
wire _58754_;
wire _58755_;
wire _58756_;
wire _58757_;
wire _58758_;
wire _58759_;
wire _58760_;
wire _58761_;
wire _58762_;
wire _58763_;
wire _58764_;
wire _58765_;
wire _58766_;
wire _58767_;
wire _58768_;
wire _58769_;
wire _58770_;
wire _58771_;
wire _58772_;
wire _58773_;
wire _58774_;
wire _58775_;
wire _58776_;
wire _58777_;
wire _58778_;
wire _58779_;
wire _58780_;
wire _58781_;
wire _58782_;
wire _58783_;
wire _58784_;
wire _58785_;
wire _58786_;
wire _58787_;
wire _58788_;
wire _58789_;
wire _58790_;
wire _58791_;
wire _58792_;
wire _58793_;
wire _58794_;
wire _58795_;
wire _58796_;
wire _58797_;
wire _58798_;
wire _58799_;
wire _58800_;
wire _58801_;
wire _58802_;
wire _58803_;
wire _58804_;
wire _58805_;
wire _58806_;
wire _58807_;
wire _58808_;
wire _58809_;
wire _58810_;
wire _58811_;
wire _58812_;
wire _58813_;
wire _58814_;
wire _58815_;
wire _58816_;
wire _58817_;
wire _58818_;
wire _58819_;
wire _58820_;
wire _58821_;
wire _58822_;
wire _58823_;
wire _58824_;
wire _58825_;
wire _58826_;
wire _58827_;
wire _58828_;
wire _58829_;
wire _58830_;
wire _58831_;
wire _58832_;
wire _58833_;
wire _58834_;
wire _58835_;
wire _58836_;
wire _58837_;
wire _58838_;
wire _58839_;
wire _58840_;
wire _58841_;
wire _58842_;
wire _58843_;
wire _58844_;
wire _58845_;
wire _58846_;
wire _58847_;
wire _58848_;
wire _58849_;
wire _58850_;
wire _58851_;
wire _58852_;
wire _58853_;
wire _58854_;
wire _58855_;
wire _58856_;
wire _58857_;
wire _58858_;
wire _58859_;
wire _58860_;
wire _58861_;
wire _58862_;
wire _58863_;
wire _58864_;
wire _58865_;
wire _58866_;
wire _58867_;
wire _58868_;
wire _58869_;
wire _58870_;
wire _58871_;
wire _58872_;
wire _58873_;
wire _58874_;
wire _58875_;
wire _58876_;
wire _58877_;
wire _58878_;
wire _58879_;
wire _58880_;
wire _58881_;
wire _58882_;
wire _58883_;
wire _58884_;
wire _58885_;
wire _58886_;
wire _58887_;
wire _58888_;
wire _58889_;
wire _58890_;
wire _58891_;
wire _58892_;
wire _58893_;
wire _58894_;
wire _58895_;
wire _58896_;
wire _58897_;
wire _58898_;
wire _58899_;
wire _58900_;
wire _58901_;
wire _58902_;
wire _58903_;
wire _58904_;
wire _58905_;
wire _58906_;
wire _58907_;
wire _58908_;
wire _58909_;
wire _58910_;
wire _58911_;
wire _58912_;
wire _58913_;
wire _58914_;
wire _58915_;
wire _58916_;
wire _58917_;
wire _58918_;
wire _58919_;
wire _58920_;
wire _58921_;
wire _58922_;
wire _58923_;
wire _58924_;
wire _58925_;
wire _58926_;
wire _58927_;
wire _58928_;
wire _58929_;
wire _58930_;
wire _58931_;
wire _58932_;
wire _58933_;
wire _58934_;
wire _58935_;
wire _58936_;
wire _58937_;
wire _58938_;
wire _58939_;
wire _58940_;
wire _58941_;
wire _58942_;
wire _58943_;
wire _58944_;
wire _58945_;
wire _58946_;
wire _58947_;
wire _58948_;
wire _58949_;
wire _58950_;
wire _58951_;
wire _58952_;
wire _58953_;
wire _58954_;
wire _58955_;
wire _58956_;
wire _58957_;
wire _58958_;
wire _58959_;
wire _58960_;
wire _58961_;
wire _58962_;
wire _58963_;
wire _58964_;
wire _58965_;
wire _58966_;
wire _58967_;
wire _58968_;
wire _58969_;
wire _58970_;
wire _58971_;
wire _58972_;
wire _58973_;
wire _58974_;
wire _58975_;
wire _58976_;
wire _58977_;
wire _58978_;
wire _58979_;
wire _58980_;
wire _58981_;
wire _58982_;
wire _58983_;
wire _58984_;
wire _58985_;
wire _58986_;
wire _58987_;
wire _58988_;
wire _58989_;
wire _58990_;
wire _58991_;
wire _58992_;
wire _58993_;
wire _58994_;
wire _58995_;
wire _58996_;
wire _58997_;
wire _58998_;
wire _58999_;
wire _59000_;
wire _59001_;
wire _59002_;
wire _59003_;
wire _59004_;
wire _59005_;
wire _59006_;
wire _59007_;
wire _59008_;
wire _59009_;
wire _59010_;
wire _59011_;
wire _59012_;
wire _59013_;
wire _59014_;
wire _59015_;
wire _59016_;
wire _59017_;
wire _59018_;
wire _59019_;
wire _59020_;
wire _59021_;
wire _59022_;
wire _59023_;
wire _59024_;
wire _59025_;
wire _59026_;
wire _59027_;
wire _59028_;
wire _59029_;
wire _59030_;
wire _59031_;
wire _59032_;
wire _59033_;
wire _59034_;
wire _59035_;
wire _59036_;
wire _59037_;
wire _59038_;
wire _59039_;
wire _59040_;
wire _59041_;
wire _59042_;
wire _59043_;
wire _59044_;
wire _59045_;
wire _59046_;
wire _59047_;
wire _59048_;
wire _59049_;
wire _59050_;
wire _59051_;
wire _59052_;
wire _59053_;
wire _59054_;
wire _59055_;
wire _59056_;
wire _59057_;
wire _59058_;
wire _59059_;
wire _59060_;
wire _59061_;
wire _59062_;
wire _59063_;
wire _59064_;
wire _59065_;
wire _59066_;
wire _59067_;
wire _59068_;
wire _59069_;
wire _59070_;
wire _59071_;
wire _59072_;
wire _59073_;
wire _59074_;
wire _59075_;
wire _59076_;
wire _59077_;
wire _59078_;
wire _59079_;
wire _59080_;
wire _59081_;
wire _59082_;
wire _59083_;
wire _59084_;
wire _59085_;
wire _59086_;
wire _59087_;
wire _59088_;
wire _59089_;
wire _59090_;
wire _59091_;
wire _59092_;
wire _59093_;
wire _59094_;
wire _59095_;
wire _59096_;
wire _59097_;
wire _59098_;
wire _59099_;
wire _59100_;
wire _59101_;
wire _59102_;
wire _59103_;
wire _59104_;
wire _59105_;
wire _59106_;
wire _59107_;
wire _59108_;
wire _59109_;
wire _59110_;
wire _59111_;
wire _59112_;
wire _59113_;
wire _59114_;
wire _59115_;
wire _59116_;
wire _59117_;
wire _59118_;
wire _59119_;
wire _59120_;
wire _59121_;
wire _59122_;
wire _59123_;
wire _59124_;
wire _59125_;
wire _59126_;
wire _59127_;
wire _59128_;
wire _59129_;
wire _59130_;
wire _59131_;
wire _59132_;
wire _59133_;
wire _59134_;
wire _59135_;
wire _59136_;
wire _59137_;
wire _59138_;
wire _59139_;
wire _59140_;
wire _59141_;
wire _59142_;
wire _59143_;
wire _59144_;
wire _59145_;
wire _59146_;
wire _59147_;
wire _59148_;
wire _59149_;
wire _59150_;
wire _59151_;
wire _59152_;
wire _59153_;
wire _59154_;
wire _59155_;
wire _59156_;
wire _59157_;
wire _59158_;
wire _59159_;
wire _59160_;
wire _59161_;
wire _59162_;
wire _59163_;
wire _59164_;
wire _59165_;
wire _59166_;
wire _59167_;
wire _59168_;
wire _59169_;
wire _59170_;
wire _59171_;
wire _59172_;
wire _59173_;
wire _59174_;
wire _59175_;
wire _59176_;
wire _59177_;
wire _59178_;
wire _59179_;
wire _59180_;
wire _59181_;
wire _59182_;
wire _59183_;
wire _59184_;
wire _59185_;
wire _59186_;
wire _59187_;
wire _59188_;
wire _59189_;
wire _59190_;
wire _59191_;
wire _59192_;
wire _59193_;
wire _59194_;
wire _59195_;
wire _59196_;
wire _59197_;
wire _59198_;
wire _59199_;
wire _59200_;
wire _59201_;
wire _59202_;
wire _59203_;
wire _59204_;
wire _59205_;
wire _59206_;
wire _59207_;
wire _59208_;
wire _59209_;
wire _59210_;
wire _59211_;
wire _59212_;
wire _59213_;
wire _59214_;
wire _59215_;
wire _59216_;
wire _59217_;
wire _59218_;
wire _59219_;
wire _59220_;
wire _59221_;
wire _59222_;
wire _59223_;
wire _59224_;
wire _59225_;
wire _59226_;
wire _59227_;
wire _59228_;
wire _59229_;
wire _59230_;
wire _59231_;
wire _59232_;
wire _59233_;
wire _59234_;
wire _59235_;
wire _59236_;
wire _59237_;
wire _59238_;
wire _59239_;
wire _59240_;
wire _59241_;
wire _59242_;
wire _59243_;
wire _59244_;
wire _59245_;
wire _59246_;
wire _59247_;
wire _59248_;
wire _59249_;
wire _59250_;
wire _59251_;
wire _59252_;
wire _59253_;
wire _59254_;
wire _59255_;
wire _59256_;
wire _59257_;
wire _59258_;
wire _59259_;
wire _59260_;
wire _59261_;
wire _59262_;
wire _59263_;
wire _59264_;
wire _59265_;
wire _59266_;
wire _59267_;
wire _59268_;
wire _59269_;
wire _59270_;
wire _59271_;
wire _59272_;
wire _59273_;
wire _59274_;
wire _59275_;
wire _59276_;
wire _59277_;
wire _59278_;
wire _59279_;
wire _59280_;
wire _59281_;
wire _59282_;
wire _59283_;
wire _59284_;
wire _59285_;
wire _59286_;
wire _59287_;
wire _59288_;
wire _59289_;
wire _59290_;
wire _59291_;
wire _59292_;
wire _59293_;
wire _59294_;
wire _59295_;
wire _59296_;
wire _59297_;
wire _59298_;
wire _59299_;
wire _59300_;
wire _59301_;
wire _59302_;
wire _59303_;
wire _59304_;
wire _59305_;
wire _59306_;
wire _59307_;
wire _59308_;
wire _59309_;
wire _59310_;
wire _59311_;
wire _59312_;
wire _59313_;
wire _59314_;
wire _59315_;
wire _59316_;
wire _59317_;
wire _59318_;
wire _59319_;
wire _59320_;
wire _59321_;
wire _59322_;
wire _59323_;
wire _59324_;
wire _59325_;
wire _59326_;
wire _59327_;
wire _59328_;
wire _59329_;
wire _59330_;
wire _59331_;
wire _59332_;
wire _59333_;
wire _59334_;
wire _59335_;
wire _59336_;
wire _59337_;
wire _59338_;
wire _59339_;
wire _59340_;
wire _59341_;
wire _59342_;
wire _59343_;
wire _59344_;
wire _59345_;
wire _59346_;
wire _59347_;
wire _59348_;
wire _59349_;
wire _59350_;
wire _59351_;
wire _59352_;
wire _59353_;
wire _59354_;
wire _59355_;
wire _59356_;
wire _59357_;
wire _59358_;
wire _59359_;
wire _59360_;
wire _59361_;
wire _59362_;
wire _59363_;
wire _59364_;
wire _59365_;
wire _59366_;
wire _59367_;
wire _59368_;
wire _59369_;
wire _59370_;
wire _59371_;
wire _59372_;
wire _59373_;
wire _59374_;
wire _59375_;
wire _59376_;
wire _59377_;
wire _59378_;
wire _59379_;
wire _59380_;
wire _59381_;
wire _59382_;
wire _59383_;
wire _59384_;
wire _59385_;
wire _59386_;
wire _59387_;
wire _59388_;
wire _59389_;
wire _59390_;
wire _59391_;
wire _59392_;
wire _59393_;
wire _59394_;
wire _59395_;
wire _59396_;
wire _59397_;
wire _59398_;
wire _59399_;
wire _59400_;
wire _59401_;
wire _59402_;
wire _59403_;
wire _59404_;
wire _59405_;
wire _59406_;
wire _59407_;
wire _59408_;
wire _59409_;
wire _59410_;
wire _59411_;
wire _59412_;
wire _59413_;
wire _59414_;
wire _59415_;
wire _59416_;
wire _59417_;
wire _59418_;
wire _59419_;
wire _59420_;
wire _59421_;
wire _59422_;
wire _59423_;
wire _59424_;
wire _59425_;
wire _59426_;
wire _59427_;
wire _59428_;
wire _59429_;
wire _59430_;
wire _59431_;
wire _59432_;
wire _59433_;
wire _59434_;
wire _59435_;
wire _59436_;
wire _59437_;
wire _59438_;
wire _59439_;
wire _59440_;
wire _59441_;
wire _59442_;
wire _59443_;
wire _59444_;
wire _59445_;
wire _59446_;
wire _59447_;
wire _59448_;
wire _59449_;
wire _59450_;
wire _59451_;
wire _59452_;
wire _59453_;
wire _59454_;
wire _59455_;
wire _59456_;
wire _59457_;
wire _59458_;
wire _59459_;
wire _59460_;
wire _59461_;
wire _59462_;
wire _59463_;
wire _59464_;
wire _59465_;
wire _59466_;
wire _59467_;
wire _59468_;
wire _59469_;
wire _59470_;
wire _59471_;
wire _59472_;
wire _59473_;
wire _59474_;
wire _59475_;
wire _59476_;
wire _59477_;
wire _59478_;
wire _59479_;
wire _59480_;
wire _59481_;
wire _59482_;
wire _59483_;
wire _59484_;
wire _59485_;
wire _59486_;
wire _59487_;
wire _59488_;
wire _59489_;
wire _59490_;
wire _59491_;
wire _59492_;
wire _59493_;
wire _59494_;
wire _59495_;
wire _59496_;
wire _59497_;
wire _59498_;
wire _59499_;
wire _59500_;
wire _59501_;
wire _59502_;
wire _59503_;
wire _59504_;
wire _59505_;
wire _59506_;
wire _59507_;
wire _59508_;
wire _59509_;
wire _59510_;
wire _59511_;
wire _59512_;
wire _59513_;
wire _59514_;
wire _59515_;
wire _59516_;
wire _59517_;
wire _59518_;
wire _59519_;
wire _59520_;
wire _59521_;
wire _59522_;
wire _59523_;
wire _59524_;
wire _59525_;
wire _59526_;
wire _59527_;
wire _59528_;
wire _59529_;
wire _59530_;
wire _59531_;
wire _59532_;
wire _59533_;
wire _59534_;
wire _59535_;
wire _59536_;
wire _59537_;
wire _59538_;
wire _59539_;
wire _59540_;
wire _59541_;
wire _59542_;
wire _59543_;
wire _59544_;
wire _59545_;
wire _59546_;
wire _59547_;
wire _59548_;
wire _59549_;
wire _59550_;
wire _59551_;
wire _59552_;
wire _59553_;
wire _59554_;
wire _59555_;
wire _59556_;
wire _59557_;
wire _59558_;
wire _59559_;
wire _59560_;
wire _59561_;
wire _59562_;
wire _59563_;
wire _59564_;
wire _59565_;
wire _59566_;
wire _59567_;
wire _59568_;
wire _59569_;
wire _59570_;
wire _59571_;
wire _59572_;
wire _59573_;
wire _59574_;
wire _59575_;
wire _59576_;
wire _59577_;
wire _59578_;
wire _59579_;
wire _59580_;
wire _59581_;
wire _59582_;
wire _59583_;
wire _59584_;
wire _59585_;
wire _59586_;
wire _59587_;
wire _59588_;
wire _59589_;
wire _59590_;
wire _59591_;
wire _59592_;
wire _59593_;
wire _59594_;
wire _59595_;
wire _59596_;
wire _59597_;
wire _59598_;
wire _59599_;
wire _59600_;
wire _59601_;
wire _59602_;
wire _59603_;
wire _59604_;
wire _59605_;
wire _59606_;
wire _59607_;
wire _59608_;
wire _59609_;
wire _59610_;
wire _59611_;
wire _59612_;
wire _59613_;
wire _59614_;
wire _59615_;
wire _59616_;
wire _59617_;
wire _59618_;
wire _59619_;
wire _59620_;
wire _59621_;
wire _59622_;
wire _59623_;
wire _59624_;
wire _59625_;
wire _59626_;
wire _59627_;
wire _59628_;
wire _59629_;
wire _59630_;
wire _59631_;
wire _59632_;
wire _59633_;
wire _59634_;
wire _59635_;
wire _59636_;
wire _59637_;
wire _59638_;
wire _59639_;
wire _59640_;
wire _59641_;
wire _59642_;
wire _59643_;
wire _59644_;
wire _59645_;
wire _59646_;
wire _59647_;
wire _59648_;
wire _59649_;
wire _59650_;
wire _59651_;
wire _59652_;
wire _59653_;
wire _59654_;
wire _59655_;
wire _59656_;
wire _59657_;
wire _59658_;
wire _59659_;
wire _59660_;
wire _59661_;
wire _59662_;
wire _59663_;
wire _59664_;
wire _59665_;
wire _59666_;
wire _59667_;
wire _59668_;
wire _59669_;
wire _59670_;
wire _59671_;
wire _59672_;
wire _59673_;
wire _59674_;
wire _59675_;
wire _59676_;
wire _59677_;
wire _59678_;
wire _59679_;
wire _59680_;
wire _59681_;
wire _59682_;
wire _59683_;
wire _59684_;
wire _59685_;
wire _59686_;
wire _59687_;
wire _59688_;
wire _59689_;
wire _59690_;
wire _59691_;
wire _59692_;
wire _59693_;
wire _59694_;
wire _59695_;
wire _59696_;
wire _59697_;
wire _59698_;
wire _59699_;
wire _59700_;
wire _59701_;
wire _59702_;
wire _59703_;
wire _59704_;
wire _59705_;
wire _59706_;
wire _59707_;
wire _59708_;
wire _59709_;
wire _59710_;
wire _59711_;
wire _59712_;
wire _59713_;
wire _59714_;
wire _59715_;
wire _59716_;
wire _59717_;
wire _59718_;
wire _59719_;
wire _59720_;
wire _59721_;
wire _59722_;
wire _59723_;
wire _59724_;
wire _59725_;
wire _59726_;
wire _59727_;
wire _59728_;
wire _59729_;
wire _59730_;
wire _59731_;
wire _59732_;
wire _59733_;
wire _59734_;
wire _59735_;
wire _59736_;
wire _59737_;
wire _59738_;
wire _59739_;
wire _59740_;
wire _59741_;
wire _59742_;
wire _59743_;
wire _59744_;
wire _59745_;
wire _59746_;
wire _59747_;
wire _59748_;
wire _59749_;
wire _59750_;
wire _59751_;
wire _59752_;
wire _59753_;
wire _59754_;
wire _59755_;
wire _59756_;
wire _59757_;
wire _59758_;
wire _59759_;
wire _59760_;
wire _59761_;
wire _59762_;
wire _59763_;
wire _59764_;
wire _59765_;
wire _59766_;
wire _59767_;
wire _59768_;
wire _59769_;
wire _59770_;
wire _59771_;
wire _59772_;
wire _59773_;
wire _59774_;
wire _59775_;
wire _59776_;
wire _59777_;
wire _59778_;
wire _59779_;
wire _59780_;
wire _59781_;
wire _59782_;
wire _59783_;
wire _59784_;
wire _59785_;
wire _59786_;
wire _59787_;
wire _59788_;
wire _59789_;
wire _59790_;
wire _59791_;
wire _59792_;
wire _59793_;
wire _59794_;
wire _59795_;
wire _59796_;
wire _59797_;
wire _59798_;
wire _59799_;
wire _59800_;
wire _59801_;
wire _59802_;
wire _59803_;
wire _59804_;
wire _59805_;
wire _59806_;
wire _59807_;
wire _59808_;
wire _59809_;
wire _59810_;
wire _59811_;
wire _59812_;
wire _59813_;
wire _59814_;
wire _59815_;
wire _59816_;
wire _59817_;
wire _59818_;
wire _59819_;
wire _59820_;
wire _59821_;
wire _59822_;
wire _59823_;
wire _59824_;
wire _59825_;
wire _59826_;
wire _59827_;
wire _59828_;
wire _59829_;
wire _59830_;
wire _59831_;
wire _59832_;
wire _59833_;
wire _59834_;
wire _59835_;
wire _59836_;
wire _59837_;
wire _59838_;
wire _59839_;
wire _59840_;
wire _59841_;
wire _59842_;
wire _59843_;
wire _59844_;
wire _59845_;
wire _59846_;
wire _59847_;
wire _59848_;
wire _59849_;
wire _59850_;
wire _59851_;
wire _59852_;
wire _59853_;
wire _59854_;
wire _59855_;
wire _59856_;
wire _59857_;
wire _59858_;
wire _59859_;
wire _59860_;
wire _59861_;
wire _59862_;
wire _59863_;
wire _59864_;
wire _59865_;
wire _59866_;
wire _59867_;
wire _59868_;
wire _59869_;
wire _59870_;
wire _59871_;
wire _59872_;
wire _59873_;
wire _59874_;
wire _59875_;
wire _59876_;
wire _59877_;
wire _59878_;
wire _59879_;
wire _59880_;
wire _59881_;
wire _59882_;
wire _59883_;
wire _59884_;
wire _59885_;
wire _59886_;
wire _59887_;
wire _59888_;
wire _59889_;
wire _59890_;
wire _59891_;
wire _59892_;
wire _59893_;
wire _59894_;
wire _59895_;
wire _59896_;
wire _59897_;
wire _59898_;
wire _59899_;
wire _59900_;
wire _59901_;
wire _59902_;
wire _59903_;
wire _59904_;
wire _59905_;
wire _59906_;
wire _59907_;
wire _59908_;
wire _59909_;
wire _59910_;
wire _59911_;
wire _59912_;
wire _59913_;
wire _59914_;
wire _59915_;
wire _59916_;
wire _59917_;
wire _59918_;
wire _59919_;
wire _59920_;
wire _59921_;
wire _59922_;
wire _59923_;
wire _59924_;
wire _59925_;
wire _59926_;
wire _59927_;
wire _59928_;
wire _59929_;
wire _59930_;
wire _59931_;
wire _59932_;
wire _59933_;
wire _59934_;
wire _59935_;
wire _59936_;
wire _59937_;
wire _59938_;
wire _59939_;
wire _59940_;
wire _59941_;
wire _59942_;
wire _59943_;
wire _59944_;
wire _59945_;
wire _59946_;
wire _59947_;
wire _59948_;
wire _59949_;
wire _59950_;
wire _59951_;
wire _59952_;
wire _59953_;
wire _59954_;
wire _59955_;
wire _59956_;
wire _59957_;
wire _59958_;
wire _59959_;
wire _59960_;
wire _59961_;
wire _59962_;
wire _59963_;
wire _59964_;
wire _59965_;
wire _59966_;
wire _59967_;
wire _59968_;
wire _59969_;
wire _59970_;
wire _59971_;
wire _59972_;
wire _59973_;
wire _59974_;
wire _59975_;
wire _59976_;
wire _59977_;
wire _59978_;
wire _59979_;
wire _59980_;
wire _59981_;
wire _59982_;
wire _59983_;
wire _59984_;
wire _59985_;
wire _59986_;
wire _59987_;
wire _59988_;
wire _59989_;
wire _59990_;
wire _59991_;
wire _59992_;
wire _59993_;
wire _59994_;
wire _59995_;
wire _59996_;
wire _59997_;
wire _59998_;
wire _59999_;
wire _60000_;
wire _60001_;
wire _60002_;
wire _60003_;
wire _60004_;
wire _60005_;
wire _60006_;
wire _60007_;
wire _60008_;
wire _60009_;
wire _60010_;
wire _60011_;
wire _60012_;
wire _60013_;
wire _60014_;
wire _60015_;
wire _60016_;
wire _60017_;
wire _60018_;
wire _60019_;
wire _60020_;
wire _60021_;
wire _60022_;
wire _60023_;
wire _60024_;
wire _60025_;
wire _60026_;
wire _60027_;
wire _60028_;
wire _60029_;
wire _60030_;
wire _60031_;
wire _60032_;
wire _60033_;
wire _60034_;
wire _60035_;
wire _60036_;
wire _60037_;
wire _60038_;
wire _60039_;
wire _60040_;
wire _60041_;
wire _60042_;
wire _60043_;
wire _60044_;
wire _60045_;
wire _60046_;
wire _60047_;
wire _60048_;
wire _60049_;
wire _60050_;
wire _60051_;
wire _60052_;
wire _60053_;
wire _60054_;
wire _60055_;
wire _60056_;
wire _60057_;
wire _60058_;
wire _60059_;
wire _60060_;
wire _60061_;
wire _60062_;
wire _60063_;
wire _60064_;
wire _60065_;
wire _60066_;
wire _60067_;
wire _60068_;
wire _60069_;
wire _60070_;
wire _60071_;
wire _60072_;
wire _60073_;
wire _60074_;
wire _60075_;
wire _60076_;
wire _60077_;
wire _60078_;
wire _60079_;
wire _60080_;
wire _60081_;
wire _60082_;
wire _60083_;
wire _60084_;
wire _60085_;
wire _60086_;
wire _60087_;
wire _60088_;
wire _60089_;
wire _60090_;
wire _60091_;
wire _60092_;
wire _60093_;
wire _60094_;
wire _60095_;
wire _60096_;
wire _60097_;
wire _60098_;
wire _60099_;
wire _60100_;
wire _60101_;
wire _60102_;
wire _60103_;
wire _60104_;
wire _60105_;
wire _60106_;
wire _60107_;
wire _60108_;
wire _60109_;
wire _60110_;
wire _60111_;
wire _60112_;
wire _60113_;
wire _60114_;
wire _60115_;
wire _60116_;
wire _60117_;
wire _60118_;
wire _60119_;
wire _60120_;
wire _60121_;
wire _60122_;
wire _60123_;
wire _60124_;
wire _60125_;
wire _60126_;
wire _60127_;
wire _60128_;
wire _60129_;
wire _60130_;
wire _60131_;
wire _60132_;
wire _60133_;
wire _60134_;
wire _60135_;
wire _60136_;
wire _60137_;
wire _60138_;
wire _60139_;
wire _60140_;
wire _60141_;
wire _60142_;
wire _60143_;
wire _60144_;
wire _60145_;
wire _60146_;
wire _60147_;
wire _60148_;
wire _60149_;
wire _60150_;
wire _60151_;
wire _60152_;
wire _60153_;
wire _60154_;
wire _60155_;
wire _60156_;
wire _60157_;
wire _60158_;
wire _60159_;
wire _60160_;
wire _60161_;
wire _60162_;
wire _60163_;
wire _60164_;
wire _60165_;
wire _60166_;
wire _60167_;
wire _60168_;
wire _60169_;
wire _60170_;
wire _60171_;
wire _60172_;
wire _60173_;
wire _60174_;
wire _60175_;
wire _60176_;
wire _60177_;
wire _60178_;
wire _60179_;
wire _60180_;
wire _60181_;
wire _60182_;
wire _60183_;
wire _60184_;
wire _60185_;
wire _60186_;
wire _60187_;
wire _60188_;
wire _60189_;
wire _60190_;
wire _60191_;
wire _60192_;
wire _60193_;
wire _60194_;
wire _60195_;
wire _60196_;
wire _60197_;
wire _60198_;
wire _60199_;
wire _60200_;
wire _60201_;
wire _60202_;
wire _60203_;
wire _60204_;
wire _60205_;
wire _60206_;
wire _60207_;
wire _60208_;
wire _60209_;
wire _60210_;
wire _60211_;
wire _60212_;
wire _60213_;
wire _60214_;
wire _60215_;
wire _60216_;
wire _60217_;
wire _60218_;
wire _60219_;
wire _60220_;
wire _60221_;
wire _60222_;
wire _60223_;
wire _60224_;
wire _60225_;
wire _60226_;
wire _60227_;
wire _60228_;
wire _60229_;
wire _60230_;
wire _60231_;
wire _60232_;
wire _60233_;
wire _60234_;
wire _60235_;
wire _60236_;
wire _60237_;
wire _60238_;
wire _60239_;
wire _60240_;
wire _60241_;
wire _60242_;
wire _60243_;
wire _60244_;
wire _60245_;
wire _60246_;
wire _60247_;
wire _60248_;
wire _60249_;
wire _60250_;
wire _60251_;
wire _60252_;
wire _60253_;
wire _60254_;
wire _60255_;
wire _60256_;
wire _60257_;
wire _60258_;
wire _60259_;
wire _60260_;
wire _60261_;
wire _60262_;
wire _60263_;
wire _60264_;
wire _60265_;
wire _60266_;
wire _60267_;
wire _60268_;
wire _60269_;
wire _60270_;
wire _60271_;
wire _60272_;
wire _60273_;
wire _60274_;
wire _60275_;
wire _60276_;
wire _60277_;
wire _60278_;
wire _60279_;
wire _60280_;
wire _60281_;
wire _60282_;
wire _60283_;
wire _60284_;
wire _60285_;
wire _60286_;
wire _60287_;
wire _60288_;
wire _60289_;
wire _60290_;
wire _60291_;
wire _60292_;
wire _60293_;
wire _60294_;
wire _60295_;
wire _60296_;
wire _60297_;
wire _60298_;
wire _60299_;
wire _60300_;
wire _60301_;
wire _60302_;
wire _60303_;
wire _60304_;
wire _60305_;
wire _60306_;
wire _60307_;
wire _60308_;
wire _60309_;
wire _60310_;
wire _60311_;
wire _60312_;
wire _60313_;
wire _60314_;
wire _60315_;
wire _60316_;
wire _60317_;
wire _60318_;
wire _60319_;
wire _60320_;
wire _60321_;
wire _60322_;
wire _60323_;
wire _60324_;
wire _60325_;
wire _60326_;
wire _60327_;
wire _60328_;
wire _60329_;
wire _60330_;
wire _60331_;
wire _60332_;
wire _60333_;
wire _60334_;
wire _60335_;
wire _60336_;
wire _60337_;
wire _60338_;
wire _60339_;
wire _60340_;
wire _60341_;
wire _60342_;
wire _60343_;
wire _60344_;
wire _60345_;
wire _60346_;
wire _60347_;
wire _60348_;
wire _60349_;
wire _60350_;
wire _60351_;
wire _60352_;
wire _60353_;
wire _60354_;
wire _60355_;
wire _60356_;
wire _60357_;
wire _60358_;
wire _60359_;
wire _60360_;
wire _60361_;
wire _60362_;
wire _60363_;
wire _60364_;
wire _60365_;
wire _60366_;
wire _60367_;
wire _60368_;
wire _60369_;
wire _60370_;
wire _60371_;
wire _60372_;
wire _60373_;
wire _60374_;
wire _60375_;
wire _60376_;
wire _60377_;
wire _60378_;
wire _60379_;
wire _60380_;
wire _60381_;
wire _60382_;
wire _60383_;
wire _60384_;
wire _60385_;
wire _60386_;
wire _60387_;
wire _60388_;
wire _60389_;
wire _60390_;
wire _60391_;
wire _60392_;
wire _60393_;
wire _60394_;
wire _60395_;
wire _60396_;
wire _60397_;
wire _60398_;
wire _60399_;
wire _60400_;
wire _60401_;
wire _60402_;
wire _60403_;
wire _60404_;
wire _60405_;
wire _60406_;
wire _60407_;
wire _60408_;
wire _60409_;
wire _60410_;
wire _60411_;
wire _60412_;
wire _60413_;
wire _60414_;
wire _60415_;
wire _60416_;
wire _60417_;
wire _60418_;
wire _60419_;
wire _60420_;
wire _60421_;
wire _60422_;
wire _60423_;
wire _60424_;
wire _60425_;
wire _60426_;
wire _60427_;
wire _60428_;
wire _60429_;
wire _60430_;
wire _60431_;
wire _60432_;
wire _60433_;
wire _60434_;
wire _60435_;
wire _60436_;
wire _60437_;
wire _60438_;
wire _60439_;
wire _60440_;
wire _60441_;
wire _60442_;
wire _60443_;
wire _60444_;
wire _60445_;
wire _60446_;
wire _60447_;
wire _60448_;
wire _60449_;
wire _60450_;
wire _60451_;
wire _60452_;
wire _60453_;
wire _60454_;
wire _60455_;
wire _60456_;
wire _60457_;
wire _60458_;
wire _60459_;
wire _60460_;
wire _60461_;
wire _60462_;
wire _60463_;
wire _60464_;
wire _60465_;
wire _60466_;
wire _60467_;
wire _60468_;
wire _60469_;
wire _60470_;
wire _60471_;
wire _60472_;
wire _60473_;
wire _60474_;
wire _60475_;
wire _60476_;
wire _60477_;
wire _60478_;
wire _60479_;
wire _60480_;
wire _60481_;
wire _60482_;
wire _60483_;
wire _60484_;
wire _60485_;
wire _60486_;
wire _60487_;
wire _60488_;
wire _60489_;
wire _60490_;
wire _60491_;
wire _60492_;
wire _60493_;
wire _60494_;
wire _60495_;
wire _60496_;
wire _60497_;
wire _60498_;
wire _60499_;
wire _60500_;
wire _60501_;
wire _60502_;
wire _60503_;
wire _60504_;
wire _60505_;
wire _60506_;
wire _60507_;
wire _60508_;
wire _60509_;
wire _60510_;
wire _60511_;
wire _60512_;
wire _60513_;
wire _60514_;
wire _60515_;
wire _60516_;
wire _60517_;
wire _60518_;
wire _60519_;
wire _60520_;
wire _60521_;
wire _60522_;
wire _60523_;
wire _60524_;
wire _60525_;
wire _60526_;
wire _60527_;
wire _60528_;
wire _60529_;
wire _60530_;
wire _60531_;
wire _60532_;
wire _60533_;
wire _60534_;
wire _60535_;
wire _60536_;
wire _60537_;
wire _60538_;
wire _60539_;
wire _60540_;
wire _60541_;
wire _60542_;
wire _60543_;
wire _60544_;
wire _60545_;
wire _60546_;
wire _60547_;
wire _60548_;
wire _60549_;
wire _60550_;
wire _60551_;
wire _60552_;
wire _60553_;
wire _60554_;
wire _60555_;
wire _60556_;
wire _60557_;
wire _60558_;
wire _60559_;
wire _60560_;
wire _60561_;
wire _60562_;
wire _60563_;
wire _60564_;
wire _60565_;
wire _60566_;
wire _60567_;
wire _60568_;
wire _60569_;
wire _60570_;
wire _60571_;
wire _60572_;
wire _60573_;
wire _60574_;
wire _60575_;
wire _60576_;
wire _60577_;
wire _60578_;
wire _60579_;
wire _60580_;
wire _60581_;
wire _60582_;
wire _60583_;
wire _60584_;
wire _60585_;
wire _60586_;
wire _60587_;
wire _60588_;
wire _60589_;
wire _60590_;
wire _60591_;
wire _60592_;
wire _60593_;
wire _60594_;
wire _60595_;
wire _60596_;
wire _60597_;
wire _60598_;
wire _60599_;
wire _60600_;
wire _60601_;
wire _60602_;
wire _60603_;
wire _60604_;
wire _60605_;
wire _60606_;
wire _60607_;
wire _60608_;
wire _60609_;
wire _60610_;
wire _60611_;
wire _60612_;
wire _60613_;
wire _60614_;
wire _60615_;
wire _60616_;
wire _60617_;
wire _60618_;
wire _60619_;
wire _60620_;
wire _60621_;
wire _60622_;
wire _60623_;
wire _60624_;
wire _60625_;
wire _60626_;
wire _60627_;
wire _60628_;
wire _60629_;
wire _60630_;
wire _60631_;
wire _60632_;
wire _60633_;
wire _60634_;
wire _60635_;
wire _60636_;
wire _60637_;
wire _60638_;
wire _60639_;
wire _60640_;
wire _60641_;
wire _60642_;
wire _60643_;
wire _60644_;
wire _60645_;
wire _60646_;
wire _60647_;
wire _60648_;
wire _60649_;
wire _60650_;
wire _60651_;
wire _60652_;
wire _60653_;
wire _60654_;
wire _60655_;
wire _60656_;
wire _60657_;
wire _60658_;
wire _60659_;
wire _60660_;
wire _60661_;
wire _60662_;
wire _60663_;
wire _60664_;
wire _60665_;
wire _60666_;
wire _60667_;
wire _60668_;
wire _60669_;
wire _60670_;
wire _60671_;
wire _60672_;
wire _60673_;
wire _60674_;
wire _60675_;
wire _60676_;
wire _60677_;
wire _60678_;
wire _60679_;
wire _60680_;
wire _60681_;
wire _60682_;
wire _60683_;
wire _60684_;
wire _60685_;
wire _60686_;
wire _60687_;
wire _60688_;
wire _60689_;
wire _60690_;
wire _60691_;
wire _60692_;
wire _60693_;
wire _60694_;
wire _60695_;
wire _60696_;
wire _60697_;
wire _60698_;
wire _60699_;
wire _60700_;
wire _60701_;
wire _60702_;
wire _60703_;
wire _60704_;
wire _60705_;
wire _60706_;
wire _60707_;
wire _60708_;
wire _60709_;
wire _60710_;
wire _60711_;
wire _60712_;
wire _60713_;
wire _60714_;
wire _60715_;
wire _60716_;
wire _60717_;
wire _60718_;
wire _60719_;
wire _60720_;
wire _60721_;
wire _60722_;
wire _60723_;
wire _60724_;
wire _60725_;
wire _60726_;
wire _60727_;
wire _60728_;
wire _60729_;
wire _60730_;
wire _60731_;
wire _60732_;
wire _60733_;
wire _60734_;
wire _60735_;
wire _60736_;
wire _60737_;
wire _60738_;
wire _60739_;
wire _60740_;
wire _60741_;
wire _60742_;
wire _60743_;
wire _60744_;
wire _60745_;
wire _60746_;
wire _60747_;
wire _60748_;
wire _60749_;
wire _60750_;
wire _60751_;
wire _60752_;
wire _60753_;
wire _60754_;
wire _60755_;
wire _60756_;
wire _60757_;
wire _60758_;
wire _60759_;
wire _60760_;
wire _60761_;
wire _60762_;
wire _60763_;
wire _60764_;
wire _60765_;
wire _60766_;
wire _60767_;
wire _60768_;
wire _60769_;
wire _60770_;
wire _60771_;
wire _60772_;
wire _60773_;
wire _60774_;
wire _60775_;
wire _60776_;
wire _60777_;
wire _60778_;
wire _60779_;
wire _60780_;
wire _60781_;
wire _60782_;
wire _60783_;
wire _60784_;
wire _60785_;
wire _60786_;
wire _60787_;
wire _60788_;
wire _60789_;
wire _60790_;
wire _60791_;
wire _60792_;
wire _60793_;
wire _60794_;
wire _60795_;
wire _60796_;
wire _60797_;
wire _60798_;
wire _60799_;
wire _60800_;
wire _60801_;
wire _60802_;
wire _60803_;
wire _60804_;
wire _60805_;
wire _60806_;
wire _60807_;
wire _60808_;
wire _60809_;
wire _60810_;
wire _60811_;
wire _60812_;
wire _60813_;
wire _60814_;
wire _60815_;
wire _60816_;
wire _60817_;
wire _60818_;
wire _60819_;
wire _60820_;
wire _60821_;
wire _60822_;
wire _60823_;
wire _60824_;
wire _60825_;
wire _60826_;
wire _60827_;
wire _60828_;
wire _60829_;
wire _60830_;
wire _60831_;
wire _60832_;
wire _60833_;
wire _60834_;
wire _60835_;
wire _60836_;
wire _60837_;
wire _60838_;
wire _60839_;
wire _60840_;
wire _60841_;
wire _60842_;
wire _60843_;
wire _60844_;
wire _60845_;
wire _60846_;
wire _60847_;
wire _60848_;
wire _60849_;
wire _60850_;
wire _60851_;
wire _60852_;
wire _60853_;
wire _60854_;
wire _60855_;
wire _60856_;
wire _60857_;
wire _60858_;
wire _60859_;
wire _60860_;
wire _60861_;
wire _60862_;
wire _60863_;
wire _60864_;
wire _60865_;
wire _60866_;
wire _60867_;
wire _60868_;
wire _60869_;
wire _60870_;
wire _60871_;
wire _60872_;
wire _60873_;
wire _60874_;
wire _60875_;
wire _60876_;
wire _60877_;
wire _60878_;
wire _60879_;
wire _60880_;
wire _60881_;
wire _60882_;
wire _60883_;
wire _60884_;
wire _60885_;
wire _60886_;
wire _60887_;
wire _60888_;
wire _60889_;
wire _60890_;
wire _60891_;
wire _60892_;
wire _60893_;
wire _60894_;
wire _60895_;
wire _60896_;
wire _60897_;
wire _60898_;
wire _60899_;
wire _60900_;
wire _60901_;
wire _60902_;
wire _60903_;
wire _60904_;
wire _60905_;
wire _60906_;
wire _60907_;
wire _60908_;
wire _60909_;
wire _60910_;
wire _60911_;
wire _60912_;
wire _60913_;
wire _60914_;
wire _60915_;
wire _60916_;
wire _60917_;
wire _60918_;
wire _60919_;
wire _60920_;
wire _60921_;
wire _60922_;
wire _60923_;
wire _60924_;
wire _60925_;
wire _60926_;
wire _60927_;
wire _60928_;
wire _60929_;
wire _60930_;
wire _60931_;
wire _60932_;
wire _60933_;
wire _60934_;
wire _60935_;
wire _60936_;
wire _60937_;
wire _60938_;
wire _60939_;
wire _60940_;
wire _60941_;
wire _60942_;
wire _60943_;
wire _60944_;
wire _60945_;
wire _60946_;
wire _60947_;
wire _60948_;
wire _60949_;
wire _60950_;
wire _60951_;
wire _60952_;
wire _60953_;
wire _60954_;
wire _60955_;
wire _60956_;
wire _60957_;
wire _60958_;
wire _60959_;
wire _60960_;
wire _60961_;
wire _60962_;
wire _60963_;
wire _60964_;
wire _60965_;
wire _60966_;
wire _60967_;
wire _60968_;
wire _60969_;
wire _60970_;
wire _60971_;
wire _60972_;
wire _60973_;
wire _60974_;
wire _60975_;
wire _60976_;
wire _60977_;
wire _60978_;
wire _60979_;
wire _60980_;
wire _60981_;
wire _60982_;
wire _60983_;
wire _60984_;
wire _60985_;
wire _60986_;
wire _60987_;
wire _60988_;
wire _60989_;
wire _60990_;
wire _60991_;
wire _60992_;
wire _60993_;
wire _60994_;
wire _60995_;
wire _60996_;
wire _60997_;
wire _60998_;
wire _60999_;
wire _61000_;
wire _61001_;
wire _61002_;
wire _61003_;
wire _61004_;
wire _61005_;
wire _61006_;
wire _61007_;
wire _61008_;
wire _61009_;
wire _61010_;
wire _61011_;
wire _61012_;
wire _61013_;
wire _61014_;
wire _61015_;
wire _61016_;
wire _61017_;
wire _61018_;
wire _61019_;
wire _61020_;
wire _61021_;
wire _61022_;
wire _61023_;
wire _61024_;
wire _61025_;
wire _61026_;
wire _61027_;
wire _61028_;
wire _61029_;
wire _61030_;
wire _61031_;
wire _61032_;
wire _61033_;
wire _61034_;
wire _61035_;
wire _61036_;
wire _61037_;
wire _61038_;
wire _61039_;
wire _61040_;
wire _61041_;
wire _61042_;
wire _61043_;
wire _61044_;
wire _61045_;
wire _61046_;
wire _61047_;
wire _61048_;
wire _61049_;
wire _61050_;
wire _61051_;
wire _61052_;
wire _61053_;
wire _61054_;
wire _61055_;
wire _61056_;
wire _61057_;
wire _61058_;
wire _61059_;
wire _61060_;
wire _61061_;
wire _61062_;
wire _61063_;
wire _61064_;
wire _61065_;
wire _61066_;
wire _61067_;
wire _61068_;
wire _61069_;
wire _61070_;
wire _61071_;
wire _61072_;
wire _61073_;
wire _61074_;
wire _61075_;
wire _61076_;
wire _61077_;
wire _61078_;
wire _61079_;
wire _61080_;
wire _61081_;
wire _61082_;
wire _61083_;
wire _61084_;
wire _61085_;
wire _61086_;
wire _61087_;
wire _61088_;
wire _61089_;
wire _61090_;
wire _61091_;
wire _61092_;
wire _61093_;
wire _61094_;
wire _61095_;
wire _61096_;
wire _61097_;
wire _61098_;
wire _61099_;
wire _61100_;
wire _61101_;
wire _61102_;
wire _61103_;
wire _61104_;
wire _61105_;
wire _61106_;
wire _61107_;
wire _61108_;
wire _61109_;
wire _61110_;
wire _61111_;
wire _61112_;
wire _61113_;
wire _61114_;
wire _61115_;
wire _61116_;
wire _61117_;
wire _61118_;
wire _61119_;
wire _61120_;
wire _61121_;
wire _61122_;
wire _61123_;
wire _61124_;
wire _61125_;
wire _61126_;
wire _61127_;
wire _61128_;
wire _61129_;
wire _61130_;
wire _61131_;
wire _61132_;
wire _61133_;
wire _61134_;
wire _61135_;
wire _61136_;
wire _61137_;
wire _61138_;
wire _61139_;
wire _61140_;
wire _61141_;
wire _61142_;
wire _61143_;
wire _61144_;
wire _61145_;
wire _61146_;
wire _61147_;
wire _61148_;
wire _61149_;
wire _61150_;
wire _61151_;
wire _61152_;
wire _61153_;
wire _61154_;
wire _61155_;
wire _61156_;
wire _61157_;
wire _61158_;
wire _61159_;
wire _61160_;
wire _61161_;
wire _61162_;
wire _61163_;
wire _61164_;
wire _61165_;
wire _61166_;
wire _61167_;
wire _61168_;
wire _61169_;
wire _61170_;
wire _61171_;
wire _61172_;
wire _61173_;
wire _61174_;
wire _61175_;
wire _61176_;
wire _61177_;
wire _61178_;
wire _61179_;
wire _61180_;
wire _61181_;
wire _61182_;
wire _61183_;
wire _61184_;
wire _61185_;
wire _61186_;
wire _61187_;
wire _61188_;
wire _61189_;
wire _61190_;
wire _61191_;
wire _61192_;
wire _61193_;
wire _61194_;
wire _61195_;
wire _61196_;
wire _61197_;
wire _61198_;
wire _61199_;
wire _61200_;
wire _61201_;
wire _61202_;
wire _61203_;
wire _61204_;
wire _61205_;
wire _61206_;
wire _61207_;
wire _61208_;
wire _61209_;
wire _61210_;
wire _61211_;
wire _61212_;
wire _61213_;
wire _61214_;
wire _61215_;
wire _61216_;
wire _61217_;
wire _61218_;
wire _61219_;
wire _61220_;
wire _61221_;
wire _61222_;
wire _61223_;
wire _61224_;
wire _61225_;
wire _61226_;
wire _61227_;
wire _61228_;
wire _61229_;
wire _61230_;
wire _61231_;
wire _61232_;
wire _61233_;
wire _61234_;
wire _61235_;
wire _61236_;
wire _61237_;
wire _61238_;
wire _61239_;
wire _61240_;
wire _61241_;
wire _61242_;
wire _61243_;
wire _61244_;
wire _61245_;
wire _61246_;
wire _61247_;
wire _61248_;
wire _61249_;
wire _61250_;
wire _61251_;
wire _61252_;
wire _61253_;
wire _61254_;
wire _61255_;
wire _61256_;
wire _61257_;
wire _61258_;
wire _61259_;
wire _61260_;
wire _61261_;
wire _61262_;
wire _61263_;
wire _61264_;
wire _61265_;
wire _61266_;
wire _61267_;
wire _61268_;
wire _61269_;
wire _61270_;
wire _61271_;
wire _61272_;
wire _61273_;
wire _61274_;
wire _61275_;
wire _61276_;
wire _61277_;
wire _61278_;
wire _61279_;
wire _61280_;
wire _61281_;
wire _61282_;
wire _61283_;
wire _61284_;
wire _61285_;
wire _61286_;
wire _61287_;
wire _61288_;
wire _61289_;
wire _61290_;
wire _61291_;
wire _61292_;
wire _61293_;
wire _61294_;
wire _61295_;
wire _61296_;
wire _61297_;
wire _61298_;
wire _61299_;
wire _61300_;
wire _61301_;
wire _61302_;
wire _61303_;
wire _61304_;
wire _61305_;
wire _61306_;
wire _61307_;
wire _61308_;
wire _61309_;
wire _61310_;
wire _61311_;
wire _61312_;
wire _61313_;
wire _61314_;
wire _61315_;
wire _61316_;
wire _61317_;
wire _61318_;
wire _61319_;
wire _61320_;
wire _61321_;
wire _61322_;
wire _61323_;
wire _61324_;
wire _61325_;
wire _61326_;
wire _61327_;
wire _61328_;
wire _61329_;
wire _61330_;
wire _61331_;
wire _61332_;
wire _61333_;
wire _61334_;
wire _61335_;
wire _61336_;
wire _61337_;
wire _61338_;
wire _61339_;
wire _61340_;
wire _61341_;
wire _61342_;
wire _61343_;
wire _61344_;
wire _61345_;
wire _61346_;
wire _61347_;
wire _61348_;
wire _61349_;
wire _61350_;
wire _61351_;
wire _61352_;
wire _61353_;
wire _61354_;
wire _61355_;
wire _61356_;
wire _61357_;
wire _61358_;
wire _61359_;
wire _61360_;
wire _61361_;
wire _61362_;
wire _61363_;
wire _61364_;
wire _61365_;
wire _61366_;
wire _61367_;
wire _61368_;
wire _61369_;
wire _61370_;
wire _61371_;
wire _61372_;
wire _61373_;
wire _61374_;
wire _61375_;
wire _61376_;
wire _61377_;
wire _61378_;
wire _61379_;
wire _61380_;
wire _61381_;
wire _61382_;
wire _61383_;
wire _61384_;
wire _61385_;
wire _61386_;
wire _61387_;
wire _61388_;
wire _61389_;
wire _61390_;
wire _61391_;
wire _61392_;
wire _61393_;
wire _61394_;
wire _61395_;
wire _61396_;
wire _61397_;
wire _61398_;
wire _61399_;
wire _61400_;
wire _61401_;
wire _61402_;
wire _61403_;
wire _61404_;
wire _61405_;
wire _61406_;
wire _61407_;
wire _61408_;
wire _61409_;
wire _61410_;
wire _61411_;
wire _61412_;
wire _61413_;
wire _61414_;
wire _61415_;
wire _61416_;
wire _61417_;
wire _61418_;
wire _61419_;
wire _61420_;
wire _61421_;
wire _61422_;
wire _61423_;
wire _61424_;
wire _61425_;
wire _61426_;
wire _61427_;
wire _61428_;
wire _61429_;
wire _61430_;
wire _61431_;
wire _61432_;
wire _61433_;
wire _61434_;
wire _61435_;
wire _61436_;
wire _61437_;
wire _61438_;
wire _61439_;
wire _61440_;
wire _61441_;
wire _61442_;
wire _61443_;
wire _61444_;
wire _61445_;
wire _61446_;
wire _61447_;
wire _61448_;
wire _61449_;
wire _61450_;
wire _61451_;
wire _61452_;
wire _61453_;
wire _61454_;
wire _61455_;
wire _61456_;
wire _61457_;
wire _61458_;
wire _61459_;
wire _61460_;
wire _61461_;
wire _61462_;
wire _61463_;
wire _61464_;
wire _61465_;
wire _61466_;
wire _61467_;
wire _61468_;
wire _61469_;
wire _61470_;
wire _61471_;
wire _61472_;
wire _61473_;
wire _61474_;
wire _61475_;
wire _61476_;
wire _61477_;
wire _61478_;
wire _61479_;
wire _61480_;
wire _61481_;
wire _61482_;
wire _61483_;
wire _61484_;
wire _61485_;
wire _61486_;
wire _61487_;
wire _61488_;
wire _61489_;
wire _61490_;
wire _61491_;
wire _61492_;
wire _61493_;
wire _61494_;
wire _61495_;
wire _61496_;
wire _61497_;
wire _61498_;
wire _61499_;
wire _61500_;
wire _61501_;
wire _61502_;
wire _61503_;
wire _61504_;
wire _61505_;
wire _61506_;
wire _61507_;
wire _61508_;
wire _61509_;
wire _61510_;
wire _61511_;
wire _61512_;
wire _61513_;
wire _61514_;
wire _61515_;
wire _61516_;
wire _61517_;
wire _61518_;
wire _61519_;
wire _61520_;
wire _61521_;
wire _61522_;
wire _61523_;
wire _61524_;
wire _61525_;
wire _61526_;
wire _61527_;
wire _61528_;
wire _61529_;
wire _61530_;
wire _61531_;
wire _61532_;
wire _61533_;
wire _61534_;
wire _61535_;
wire _61536_;
wire _61537_;
wire _61538_;
wire _61539_;
wire _61540_;
wire _61541_;
wire _61542_;
wire _61543_;
wire _61544_;
wire _61545_;
wire _61546_;
wire _61547_;
wire _61548_;
wire _61549_;
wire _61550_;
wire _61551_;
wire _61552_;
wire _61553_;
wire _61554_;
wire _61555_;
wire _61556_;
wire _61557_;
wire _61558_;
wire _61559_;
wire _61560_;
wire _61561_;
wire _61562_;
wire _61563_;
wire _61564_;
wire _61565_;
wire _61566_;
wire _61567_;
wire _61568_;
wire _61569_;
wire _61570_;
wire _61571_;
wire _61572_;
wire _61573_;
wire _61574_;
wire _61575_;
wire _61576_;
wire _61577_;
wire _61578_;
wire _61579_;
wire _61580_;
wire _61581_;
wire _61582_;
wire _61583_;
wire _61584_;
wire _61585_;
wire _61586_;
wire _61587_;
wire _61588_;
wire _61589_;
wire _61590_;
wire _61591_;
wire _61592_;
wire _61593_;
wire _61594_;
wire _61595_;
wire _61596_;
wire _61597_;
wire _61598_;
wire _61599_;
wire _61600_;
wire _61601_;
wire _61602_;
wire _61603_;
wire _61604_;
wire _61605_;
wire _61606_;
wire _61607_;
wire _61608_;
wire _61609_;
wire _61610_;
wire _61611_;
wire _61612_;
wire _61613_;
wire _61614_;
wire _61615_;
wire _61616_;
wire _61617_;
wire _61618_;
wire _61619_;
wire _61620_;
wire _61621_;
wire _61622_;
wire _61623_;
wire _61624_;
wire _61625_;
wire _61626_;
wire _61627_;
wire _61628_;
wire _61629_;
wire _61630_;
wire _61631_;
wire _61632_;
wire _61633_;
wire _61634_;
wire _61635_;
wire _61636_;
wire _61637_;
wire _61638_;
wire _61639_;
wire _61640_;
wire _61641_;
wire _61642_;
wire _61643_;
wire _61644_;
wire _61645_;
wire _61646_;
wire _61647_;
wire _61648_;
wire _61649_;
wire _61650_;
wire _61651_;
wire _61652_;
wire _61653_;
wire _61654_;
wire _61655_;
wire _61656_;
wire _61657_;
wire _61658_;
wire _61659_;
wire _61660_;
wire _61661_;
wire _61662_;
wire _61663_;
wire _61664_;
wire _61665_;
wire _61666_;
wire _61667_;
wire _61668_;
wire _61669_;
wire _61670_;
wire _61671_;
wire _61672_;
wire _61673_;
wire _61674_;
wire _61675_;
wire _61676_;
wire _61677_;
wire _61678_;
wire _61679_;
wire _61680_;
wire _61681_;
wire _61682_;
wire _61683_;
wire _61684_;
wire _61685_;
wire _61686_;
wire _61687_;
wire _61688_;
wire _61689_;
wire _61690_;
wire _61691_;
wire _61692_;
wire _61693_;
wire _61694_;
wire _61695_;
wire _61696_;
wire _61697_;
wire _61698_;
wire _61699_;
wire _61700_;
wire _61701_;
wire _61702_;
wire _61703_;
wire _61704_;
wire _61705_;
wire _61706_;
wire _61707_;
wire _61708_;
wire _61709_;
wire _61710_;
wire _61711_;
wire _61712_;
wire _61713_;
wire _61714_;
wire _61715_;
wire _61716_;
wire _61717_;
wire _61718_;
wire _61719_;
wire _61720_;
wire _61721_;
wire _61722_;
wire _61723_;
wire _61724_;
wire _61725_;
wire _61726_;
wire _61727_;
wire _61728_;
wire _61729_;
wire _61730_;
wire _61731_;
wire _61732_;
wire _61733_;
wire _61734_;
wire _61735_;
wire _61736_;
wire _61737_;
wire _61738_;
wire _61739_;
wire _61740_;
wire _61741_;
wire _61742_;
wire _61743_;
wire _61744_;
wire _61745_;
wire _61746_;
wire _61747_;
wire _61748_;
wire _61749_;
wire _61750_;
wire _61751_;
wire _61752_;
wire _61753_;
wire _61754_;
wire _61755_;
wire _61756_;
wire _61757_;
wire _61758_;
wire _61759_;
wire _61760_;
wire _61761_;
wire _61762_;
wire _61763_;
wire _61764_;
wire _61765_;
wire _61766_;
wire _61767_;
wire _61768_;
wire _61769_;
wire _61770_;
wire _61771_;
wire _61772_;
wire _61773_;
wire _61774_;
wire _61775_;
wire _61776_;
wire _61777_;
wire _61778_;
wire _61779_;
wire _61780_;
wire _61781_;
wire _61782_;
wire _61783_;
wire _61784_;
wire _61785_;
wire _61786_;
wire _61787_;
wire _61788_;
wire _61789_;
wire _61790_;
wire _61791_;
wire _61792_;
wire _61793_;
wire _61794_;
wire _61795_;
wire _61796_;
wire _61797_;
wire _61798_;
wire _61799_;
wire _61800_;
wire _61801_;
wire _61802_;
wire _61803_;
wire _61804_;
wire _61805_;
wire _61806_;
wire _61807_;
wire _61808_;
wire _61809_;
wire _61810_;
wire _61811_;
wire _61812_;
wire _61813_;
wire _61814_;
wire _61815_;
wire _61816_;
wire _61817_;
wire _61818_;
wire _61819_;
wire _61820_;
wire _61821_;
wire _61822_;
wire _61823_;
wire _61824_;
wire _61825_;
wire _61826_;
wire _61827_;
wire _61828_;
wire _61829_;
wire _61830_;
wire _61831_;
wire _61832_;
wire _61833_;
wire _61834_;
wire _61835_;
wire _61836_;
wire _61837_;
wire _61838_;
wire _61839_;
wire _61840_;
wire _61841_;
wire _61842_;
wire _61843_;
wire _61844_;
wire _61845_;
wire _61846_;
wire _61847_;
wire _61848_;
wire _61849_;
wire _61850_;
wire _61851_;
wire _61852_;
wire _61853_;
wire _61854_;
wire _61855_;
wire _61856_;
wire _61857_;
wire _61858_;
wire _61859_;
wire _61860_;
wire _61861_;
wire _61862_;
wire _61863_;
wire _61864_;
wire _61865_;
wire _61866_;
wire _61867_;
wire _61868_;
wire _61869_;
wire _61870_;
wire _61871_;
wire _61872_;
wire _61873_;
wire _61874_;
wire _61875_;
wire _61876_;
wire _61877_;
wire _61878_;
wire _61879_;
wire _61880_;
wire _61881_;
wire _61882_;
wire _61883_;
wire _61884_;
wire _61885_;
wire _61886_;
wire _61887_;
wire _61888_;
wire _61889_;
wire _61890_;
wire _61891_;
wire _61892_;
wire _61893_;
wire _61894_;
wire _61895_;
wire _61896_;
wire _61897_;
wire _61898_;
wire _61899_;
wire _61900_;
wire _61901_;
wire _61902_;
wire _61903_;
wire _61904_;
wire _61905_;
wire _61906_;
wire _61907_;
wire _61908_;
wire _61909_;
wire _61910_;
wire _61911_;
wire _61912_;
wire _61913_;
wire _61914_;
wire _61915_;
wire _61916_;
wire _61917_;
wire _61918_;
wire _61919_;
wire _61920_;
wire _61921_;
wire _61922_;
wire _61923_;
wire _61924_;
wire _61925_;
wire _61926_;
wire _61927_;
wire _61928_;
wire _61929_;
wire _61930_;
wire _61931_;
wire _61932_;
wire _61933_;
wire _61934_;
wire _61935_;
wire _61936_;
wire _61937_;
wire _61938_;
wire _61939_;
wire _61940_;
wire _61941_;
wire _61942_;
wire _61943_;
wire _61944_;
wire _61945_;
wire _61946_;
wire _61947_;
wire _61948_;
wire _61949_;
wire _61950_;
wire _61951_;
wire _61952_;
wire _61953_;
wire _61954_;
wire _61955_;
wire _61956_;
wire _61957_;
wire _61958_;
wire _61959_;
wire _61960_;
wire _61961_;
wire _61962_;
wire _61963_;
wire _61964_;
wire _61965_;
wire _61966_;
wire _61967_;
wire _61968_;
wire _61969_;
wire _61970_;
wire _61971_;
wire _61972_;
wire _61973_;
wire _61974_;
wire _61975_;
wire _61976_;
wire _61977_;
wire _61978_;
wire _61979_;
wire _61980_;
wire _61981_;
wire _61982_;
wire _61983_;
wire _61984_;
wire _61985_;
wire _61986_;
wire _61987_;
wire _61988_;
wire _61989_;
wire _61990_;
wire _61991_;
wire _61992_;
wire _61993_;
wire _61994_;
wire _61995_;
wire _61996_;
wire _61997_;
wire _61998_;
wire _61999_;
wire _62000_;
wire _62001_;
wire _62002_;
wire _62003_;
wire _62004_;
wire _62005_;
wire _62006_;
wire _62007_;
wire _62008_;
wire _62009_;
wire _62010_;
wire _62011_;
wire _62012_;
wire _62013_;
wire _62014_;
wire _62015_;
wire _62016_;
wire _62017_;
wire _62018_;
wire _62019_;
wire _62020_;
wire _62021_;
wire _62022_;
wire _62023_;
wire _62024_;
wire _62025_;
wire _62026_;
wire _62027_;
wire _62028_;
wire _62029_;
wire _62030_;
wire _62031_;
wire _62032_;
wire _62033_;
wire _62034_;
wire _62035_;
wire _62036_;
wire _62037_;
wire _62038_;
wire _62039_;
wire _62040_;
wire _62041_;
wire _62042_;
wire _62043_;
wire _62044_;
wire _62045_;
wire _62046_;
wire _62047_;
wire _62048_;
wire _62049_;
wire _62050_;
wire _62051_;
wire _62052_;
wire _62053_;
wire _62054_;
wire _62055_;
wire _62056_;
wire _62057_;
wire _62058_;
wire _62059_;
wire _62060_;
wire _62061_;
wire _62062_;
wire _62063_;
wire _62064_;
wire _62065_;
wire _62066_;
wire _62067_;
wire _62068_;
wire _62069_;
wire _62070_;
wire _62071_;
wire _62072_;
wire _62073_;
wire _62074_;
wire _62075_;
wire _62076_;
wire _62077_;
wire _62078_;
wire _62079_;
wire _62080_;
wire _62081_;
wire _62082_;
wire _62083_;
wire _62084_;
wire _62085_;
wire _62086_;
wire _62087_;
wire _62088_;
wire _62089_;
wire _62090_;
wire _62091_;
wire _62092_;
wire _62093_;
wire _62094_;
wire _62095_;
wire _62096_;
wire _62097_;
wire _62098_;
wire _62099_;
wire _62100_;
wire _62101_;
wire _62102_;
wire _62103_;
wire _62104_;
wire _62105_;
wire _62106_;
wire _62107_;
wire _62108_;
wire _62109_;
wire _62110_;
wire _62111_;
wire _62112_;
wire _62113_;
wire _62114_;
wire _62115_;
wire _62116_;
wire _62117_;
wire _62118_;
wire _62119_;
wire _62120_;
wire _62121_;
wire _62122_;
wire _62123_;
wire _62124_;
wire _62125_;
wire _62126_;
wire _62127_;
wire _62128_;
wire _62129_;
wire _62130_;
wire _62131_;
wire _62132_;
wire _62133_;
wire _62134_;
wire _62135_;
wire _62136_;
wire _62137_;
wire _62138_;
wire _62139_;
wire _62140_;
wire _62141_;
wire _62142_;
wire _62143_;
wire _62144_;
wire _62145_;
wire _62146_;
wire _62147_;
wire _62148_;
wire _62149_;
wire _62150_;
wire _62151_;
wire _62152_;
wire _62153_;
wire _62154_;
wire _62155_;
wire _62156_;
wire _62157_;
wire _62158_;
wire _62159_;
wire _62160_;
wire _62161_;
wire _62162_;
wire _62163_;
wire _62164_;
wire _62165_;
wire _62166_;
wire _62167_;
wire _62168_;
wire _62169_;
wire _62170_;
wire _62171_;
wire _62172_;
wire _62173_;
wire _62174_;
wire _62175_;
wire _62176_;
wire _62177_;
wire _62178_;
wire _62179_;
wire _62180_;
wire _62181_;
wire _62182_;
wire _62183_;
wire _62184_;
wire _62185_;
wire _62186_;
wire _62187_;
wire _62188_;
wire _62189_;
wire _62190_;
wire _62191_;
wire _62192_;
wire _62193_;
wire _62194_;
wire _62195_;
wire _62196_;
wire _62197_;
wire _62198_;
wire _62199_;
wire _62200_;
wire _62201_;
wire _62202_;
wire _62203_;
wire _62204_;
wire _62205_;
wire _62206_;
wire _62207_;
wire _62208_;
wire _62209_;
wire _62210_;
wire _62211_;
wire _62212_;
wire _62213_;
wire _62214_;
wire _62215_;
wire _62216_;
wire _62217_;
wire _62218_;
wire _62219_;
wire _62220_;
wire _62221_;
wire _62222_;
wire _62223_;
wire _62224_;
wire _62225_;
wire _62226_;
wire _62227_;
wire _62228_;
wire _62229_;
wire _62230_;
wire _62231_;
wire _62232_;
wire _62233_;
wire _62234_;
wire _62235_;
wire _62236_;
wire _62237_;
wire _62238_;
wire _62239_;
wire _62240_;
wire _62241_;
wire _62242_;
wire _62243_;
wire _62244_;
wire _62245_;
wire _62246_;
wire _62247_;
wire _62248_;
wire _62249_;
wire _62250_;
wire _62251_;
wire _62252_;
wire _62253_;
wire _62254_;
wire _62255_;
wire _62256_;
wire _62257_;
wire _62258_;
wire _62259_;
wire _62260_;
wire _62261_;
wire _62262_;
wire _62263_;
wire _62264_;
wire _62265_;
wire _62266_;
wire _62267_;
wire _62268_;
wire _62269_;
wire _62270_;
wire _62271_;
wire _62272_;
wire _62273_;
wire _62274_;
wire _62275_;
wire _62276_;
wire _62277_;
wire _62278_;
wire _62279_;
wire _62280_;
wire _62281_;
wire _62282_;
wire _62283_;
wire _62284_;
wire _62285_;
wire _62286_;
wire _62287_;
wire _62288_;
wire _62289_;
wire _62290_;
wire _62291_;
wire _62292_;
wire _62293_;
wire _62294_;
wire _62295_;
wire _62296_;
wire _62297_;
wire _62298_;
wire _62299_;
wire _62300_;
wire _62301_;
wire _62302_;
wire _62303_;
wire _62304_;
wire _62305_;
wire _62306_;
wire _62307_;
wire _62308_;
wire _62309_;
wire _62310_;
wire _62311_;
wire _62312_;
wire _62313_;
wire _62314_;
wire _62315_;
wire _62316_;
wire _62317_;
wire _62318_;
wire _62319_;
wire _62320_;
wire _62321_;
wire _62322_;
wire _62323_;
wire _62324_;
wire _62325_;
wire _62326_;
wire _62327_;
wire _62328_;
wire _62329_;
wire _62330_;
wire _62331_;
wire _62332_;
wire _62333_;
wire _62334_;
wire _62335_;
wire _62336_;
wire _62337_;
wire _62338_;
wire _62339_;
wire _62340_;
wire _62341_;
wire _62342_;
wire _62343_;
wire _62344_;
wire _62345_;
wire _62346_;
wire _62347_;
wire _62348_;
wire _62349_;
wire _62350_;
wire _62351_;
wire _62352_;
wire _62353_;
wire _62354_;
wire _62355_;
wire _62356_;
wire _62357_;
wire _62358_;
wire _62359_;
wire _62360_;
wire _62361_;
wire _62362_;
wire _62363_;
wire _62364_;
wire _62365_;
wire _62366_;
wire _62367_;
wire _62368_;
wire _62369_;
wire _62370_;
wire _62371_;
wire _62372_;
wire _62373_;
wire _62374_;
wire _62375_;
wire _62376_;
wire _62377_;
wire _62378_;
wire _62379_;
wire _62380_;
wire _62381_;
wire _62382_;
wire _62383_;
wire _62384_;
wire _62385_;
wire _62386_;
wire _62387_;
wire _62388_;
wire _62389_;
wire _62390_;
wire _62391_;
wire _62392_;
wire _62393_;
wire _62394_;
wire _62395_;
wire _62396_;
wire _62397_;
wire _62398_;
wire _62399_;
wire _62400_;
wire _62401_;
wire _62402_;
wire _62403_;
wire _62404_;
wire _62405_;
wire _62406_;
wire _62407_;
wire _62408_;
wire _62409_;
wire _62410_;
wire _62411_;
wire _62412_;
wire _62413_;
wire _62414_;
wire _62415_;
wire _62416_;
wire _62417_;
wire _62418_;
wire _62419_;
wire _62420_;
wire _62421_;
wire _62422_;
wire _62423_;
wire _62424_;
wire _62425_;
wire _62426_;
wire _62427_;
wire _62428_;
wire _62429_;
wire _62430_;
wire _62431_;
wire _62432_;
wire _62433_;
wire _62434_;
wire _62435_;
wire _62436_;
wire _62437_;
wire _62438_;
wire _62439_;
wire _62440_;
wire _62441_;
wire _62442_;
wire _62443_;
wire _62444_;
wire _62445_;
wire _62446_;
wire _62447_;
wire _62448_;
wire _62449_;
wire _62450_;
wire _62451_;
wire _62452_;
wire _62453_;
wire _62454_;
wire _62455_;
wire _62456_;
wire _62457_;
wire _62458_;
wire _62459_;
wire _62460_;
wire _62461_;
wire _62462_;
wire _62463_;
wire _62464_;
wire _62465_;
wire _62466_;
wire _62467_;
wire _62468_;
wire _62469_;
wire _62470_;
wire _62471_;
wire _62472_;
wire _62473_;
wire _62474_;
wire _62475_;
wire _62476_;
wire _62477_;
wire _62478_;
wire _62479_;
wire _62480_;
wire _62481_;
wire _62482_;
wire _62483_;
wire _62484_;
wire _62485_;
wire _62486_;
wire _62487_;
wire _62488_;
wire _62489_;
wire _62490_;
wire _62491_;
wire _62492_;
wire _62493_;
wire _62494_;
wire _62495_;
wire _62496_;
wire _62497_;
wire _62498_;
wire _62499_;
wire _62500_;
wire _62501_;
wire _62502_;
wire _62503_;
wire _62504_;
wire _62505_;
wire _62506_;
wire _62507_;
wire _62508_;
wire _62509_;
wire _62510_;
wire _62511_;
wire _62512_;
wire _62513_;
wire _62514_;
wire _62515_;
wire _62516_;
wire _62517_;
wire _62518_;
wire _62519_;
wire _62520_;
wire _62521_;
wire _62522_;
wire _62523_;
wire _62524_;
wire _62525_;
wire _62526_;
wire _62527_;
wire _62528_;
wire _62529_;
wire _62530_;
wire _62531_;
wire _62532_;
wire _62533_;
wire _62534_;
wire _62535_;
wire _62536_;
wire _62537_;
wire _62538_;
wire _62539_;
wire _62540_;
wire _62541_;
wire _62542_;
wire _62543_;
wire _62544_;
wire _62545_;
wire _62546_;
wire _62547_;
wire _62548_;
wire _62549_;
wire _62550_;
wire _62551_;
wire _62552_;
wire _62553_;
wire _62554_;
wire _62555_;
wire _62556_;
wire _62557_;
wire _62558_;
wire _62559_;
wire _62560_;
wire _62561_;
wire _62562_;
wire _62563_;
wire _62564_;
wire _62565_;
wire _62566_;
wire _62567_;
wire _62568_;
wire _62569_;
wire _62570_;
wire _62571_;
wire _62572_;
wire _62573_;
wire _62574_;
wire _62575_;
wire _62576_;
wire _62577_;
wire _62578_;
wire _62579_;
wire _62580_;
wire _62581_;
wire _62582_;
wire _62583_;
wire _62584_;
wire _62585_;
wire _62586_;
wire _62587_;
wire _62588_;
wire _62589_;
wire _62590_;
wire _62591_;
wire _62592_;
wire _62593_;
wire _62594_;
wire _62595_;
wire _62596_;
wire _62597_;
wire _62598_;
wire _62599_;
wire _62600_;
wire _62601_;
wire _62602_;
wire _62603_;
wire _62604_;
wire _62605_;
wire _62606_;
wire _62607_;
wire _62608_;
wire _62609_;
wire _62610_;
wire _62611_;
wire _62612_;
wire _62613_;
wire _62614_;
wire _62615_;
wire _62616_;
wire _62617_;
wire _62618_;
wire _62619_;
wire _62620_;
wire _62621_;
wire _62622_;
wire _62623_;
wire _62624_;
wire _62625_;
wire _62626_;
wire _62627_;
wire _62628_;
wire _62629_;
wire _62630_;
wire _62631_;
wire _62632_;
wire _62633_;
wire _62634_;
wire _62635_;
wire _62636_;
wire _62637_;
wire _62638_;
wire _62639_;
wire _62640_;
wire _62641_;
wire _62642_;
wire _62643_;
wire _62644_;
wire _62645_;
wire _62646_;
wire _62647_;
wire _62648_;
wire _62649_;
wire _62650_;
wire _62651_;
wire _62652_;
wire _62653_;
wire _62654_;
wire _62655_;
wire _62656_;
wire _62657_;
wire _62658_;
wire _62659_;
wire _62660_;
wire _62661_;
wire _62662_;
wire _62663_;
wire _62664_;
wire _62665_;
wire _62666_;
wire _62667_;
wire _62668_;
wire _62669_;
wire _62670_;
wire _62671_;
wire _62672_;
wire _62673_;
wire _62674_;
wire _62675_;
wire _62676_;
wire _62677_;
wire _62678_;
wire _62679_;
wire _62680_;
wire _62681_;
wire _62682_;
wire _62683_;
wire _62684_;
wire _62685_;
wire _62686_;
wire _62687_;
wire _62688_;
wire _62689_;
wire _62690_;
wire _62691_;
wire _62692_;
wire _62693_;
wire _62694_;
wire _62695_;
wire _62696_;
wire _62697_;
wire _62698_;
wire _62699_;
wire _62700_;
wire _62701_;
wire _62702_;
wire _62703_;
wire _62704_;
wire _62705_;
wire _62706_;
wire _62707_;
wire _62708_;
wire _62709_;
wire _62710_;
wire _62711_;
wire _62712_;
wire _62713_;
wire _62714_;
wire _62715_;
wire _62716_;
wire _62717_;
wire _62718_;
wire _62719_;
wire _62720_;
wire _62721_;
wire _62722_;
wire _62723_;
wire _62724_;
wire _62725_;
wire _62726_;
wire _62727_;
wire _62728_;
wire _62729_;
wire _62730_;
wire _62731_;
wire _62732_;
wire _62733_;
wire _62734_;
wire _62735_;
wire _62736_;
wire _62737_;
wire _62738_;
wire _62739_;
wire _62740_;
wire _62741_;
wire _62742_;
wire _62743_;
wire _62744_;
wire _62745_;
wire _62746_;
wire _62747_;
wire _62748_;
wire _62749_;
wire _62750_;
wire _62751_;
wire _62752_;
wire _62753_;
wire _62754_;
wire _62755_;
wire _62756_;
wire _62757_;
wire _62758_;
wire _62759_;
wire _62760_;
wire _62761_;
wire _62762_;
wire _62763_;
wire _62764_;
wire _62765_;
wire _62766_;
wire _62767_;
wire _62768_;
wire _62769_;
wire _62770_;
wire _62771_;
wire _62772_;
wire _62773_;
wire _62774_;
wire _62775_;
wire _62776_;
wire _62777_;
wire _62778_;
wire _62779_;
wire _62780_;
wire _62781_;
wire _62782_;
wire _62783_;
wire _62784_;
wire _62785_;
wire _62786_;
wire _62787_;
wire _62788_;
wire _62789_;
wire _62790_;
wire _62791_;
wire _62792_;
wire _62793_;
wire _62794_;
wire _62795_;
wire _62796_;
wire _62797_;
wire _62798_;
wire _62799_;
wire _62800_;
wire _62801_;
wire _62802_;
wire _62803_;
wire _62804_;
wire _62805_;
wire _62806_;
wire _62807_;
wire _62808_;
wire _62809_;
wire _62810_;
wire _62811_;
wire _62812_;
wire _62813_;
wire _62814_;
wire _62815_;
wire _62816_;
wire _62817_;
wire _62818_;
wire _62819_;
wire _62820_;
wire _62821_;
wire _62822_;
wire _62823_;
wire _62824_;
wire _62825_;
wire _62826_;
wire _62827_;
wire _62828_;
wire _62829_;
wire _62830_;
wire _62831_;
wire _62832_;
wire _62833_;
wire _62834_;
wire _62835_;
wire _62836_;
wire _62837_;
wire _62838_;
wire _62839_;
wire _62840_;
wire _62841_;
wire _62842_;
wire _62843_;
wire _62844_;
wire _62845_;
wire _62846_;
wire _62847_;
wire _62848_;
wire _62849_;
wire _62850_;
wire _62851_;
wire _62852_;
wire _62853_;
wire _62854_;
wire _62855_;
wire _62856_;
wire _62857_;
wire _62858_;
wire _62859_;
wire _62860_;
wire _62861_;
wire _62862_;
wire _62863_;
wire _62864_;
wire _62865_;
wire _62866_;
wire _62867_;
wire _62868_;
wire _62869_;
wire _62870_;
wire _62871_;
wire _62872_;
wire _62873_;
wire _62874_;
wire _62875_;
wire _62876_;
wire _62877_;
wire _62878_;
wire _62879_;
wire _62880_;
wire _62881_;
wire _62882_;
wire _62883_;
wire _62884_;
wire _62885_;
wire _62886_;
wire _62887_;
wire _62888_;
wire _62889_;
wire _62890_;
wire _62891_;
wire _62892_;
wire _62893_;
wire _62894_;
wire _62895_;
wire _62896_;
wire _62897_;
wire _62898_;
wire _62899_;
wire _62900_;
wire _62901_;
wire _62902_;
wire _62903_;
wire _62904_;
wire _62905_;
wire _62906_;
wire _62907_;
wire _62908_;
wire _62909_;
wire _62910_;
wire _62911_;
wire _62912_;
wire _62913_;
wire _62914_;
wire _62915_;
wire _62916_;
wire _62917_;
wire _62918_;
wire _62919_;
wire _62920_;
wire _62921_;
wire _62922_;
wire _62923_;
wire _62924_;
wire _62925_;
wire _62926_;
wire _62927_;
wire _62928_;
wire _62929_;
wire _62930_;
wire _62931_;
wire _62932_;
wire _62933_;
wire _62934_;
wire _62935_;
wire _62936_;
wire _62937_;
wire _62938_;
wire _62939_;
wire _62940_;
wire _62941_;
wire _62942_;
wire _62943_;
wire _62944_;
wire _62945_;
wire _62946_;
wire _62947_;
wire _62948_;
wire _62949_;
wire _62950_;
wire _62951_;
wire _62952_;
wire _62953_;
wire _62954_;
wire _62955_;
wire _62956_;
wire _62957_;
wire _62958_;
wire _62959_;
wire _62960_;
wire _62961_;
wire _62962_;
wire _62963_;
wire _62964_;
wire _62965_;
wire _62966_;
wire _62967_;
wire _62968_;
wire _62969_;
wire _62970_;
wire _62971_;
wire _62972_;
wire _62973_;
wire _62974_;
wire _62975_;
wire _62976_;
wire _62977_;
wire _62978_;
wire _62979_;
wire _62980_;
wire _62981_;
wire _62982_;
wire _62983_;
wire _62984_;
wire _62985_;
wire _62986_;
wire _62987_;
wire _62988_;
wire _62989_;
wire _62990_;
wire _62991_;
wire _62992_;
wire _62993_;
wire _62994_;
wire _62995_;
wire _62996_;
wire _62997_;
wire _62998_;
wire _62999_;
wire _63000_;
wire _63001_;
wire _63002_;
wire _63003_;
wire _63004_;
wire _63005_;
wire _63006_;
wire _63007_;
wire _63008_;
wire _63009_;
wire _63010_;
wire _63011_;
wire _63012_;
wire _63013_;
wire _63014_;
wire _63015_;
wire _63016_;
wire _63017_;
wire _63018_;
wire _63019_;
wire _63020_;
wire _63021_;
wire _63022_;
wire _63023_;
wire _63024_;
wire _63025_;
wire _63026_;
wire _63027_;
wire _63028_;
wire _63029_;
wire _63030_;
wire _63031_;
wire _63032_;
wire _63033_;
wire _63034_;
wire _63035_;
wire _63036_;
wire _63037_;
wire _63038_;
wire _63039_;
wire _63040_;
wire _63041_;
wire _63042_;
wire _63043_;
wire _63044_;
wire _63045_;
wire _63046_;
wire _63047_;
wire _63048_;
wire _63049_;
wire _63050_;
wire _63051_;
wire _63052_;
wire _63053_;
wire _63054_;
wire _63055_;
wire _63056_;
wire _63057_;
wire _63058_;
wire _63059_;
wire _63060_;
wire _63061_;
wire _63062_;
wire _63063_;
wire _63064_;
wire _63065_;
wire _63066_;
wire _63067_;
wire _63068_;
wire _63069_;
wire _63070_;
wire _63071_;
wire _63072_;
wire _63073_;
wire _63074_;
wire _63075_;
wire _63076_;
wire _63077_;
wire _63078_;
wire _63079_;
wire _63080_;
wire _63081_;
wire _63082_;
wire _63083_;
wire _63084_;
wire _63085_;
wire _63086_;
wire _63087_;
wire _63088_;
wire _63089_;
wire _63090_;
wire _63091_;
wire _63092_;
wire _63093_;
wire _63094_;
wire _63095_;
wire _63096_;
wire _63097_;
wire _63098_;
wire _63099_;
wire _63100_;
wire _63101_;
wire _63102_;
wire _63103_;
wire _63104_;
wire _63105_;
wire _63106_;
wire _63107_;
wire _63108_;
wire _63109_;
wire _63110_;
wire _63111_;
wire _63112_;
wire _63113_;
wire _63114_;
wire _63115_;
wire _63116_;
wire _63117_;
wire _63118_;
wire _63119_;
wire _63120_;
wire _63121_;
wire _63122_;
wire _63123_;
wire _63124_;
wire _63125_;
wire _63126_;
wire _63127_;
wire _63128_;
wire _63129_;
wire _63130_;
wire _63131_;
wire _63132_;
wire _63133_;
wire _63134_;
wire _63135_;
wire _63136_;
wire _63137_;
wire _63138_;
wire _63139_;
wire _63140_;
wire _63141_;
wire _63142_;
wire _63143_;
wire _63144_;
wire _63145_;
wire _63146_;
wire _63147_;
wire _63148_;
wire _63149_;
wire _63150_;
wire _63151_;
wire _63152_;
wire _63153_;
wire _63154_;
wire _63155_;
wire _63156_;
wire _63157_;
wire _63158_;
wire _63159_;
wire _63160_;
wire _63161_;
wire _63162_;
wire _63163_;
wire _63164_;
wire _63165_;
wire _63166_;
wire _63167_;
wire _63168_;
wire _63169_;
wire _63170_;
wire _63171_;
wire _63172_;
wire _63173_;
wire _63174_;
wire _63175_;
wire _63176_;
wire _63177_;
wire _63178_;
wire _63179_;
wire _63180_;
wire _63181_;
wire _63182_;
wire _63183_;
wire _63184_;
wire _63185_;
wire _63186_;
wire _63187_;
wire _63188_;
wire _63189_;
wire _63190_;
wire _63191_;
wire _63192_;
wire _63193_;
wire _63194_;
wire _63195_;
wire _63196_;
wire _63197_;
wire _63198_;
wire _63199_;
wire _63200_;
wire _63201_;
wire _63202_;
wire _63203_;
wire _63204_;
wire _63205_;
wire _63206_;
wire _63207_;
wire _63208_;
wire _63209_;
wire _63210_;
wire _63211_;
wire _63212_;
wire _63213_;
wire _63214_;
wire _63215_;
wire _63216_;
wire _63217_;
wire _63218_;
wire _63219_;
wire _63220_;
wire _63221_;
wire _63222_;
wire _63223_;
wire _63224_;
wire _63225_;
wire _63226_;
wire _63227_;
wire _63228_;
wire _63229_;
wire _63230_;
wire _63231_;
wire _63232_;
wire _63233_;
wire _63234_;
wire _63235_;
wire _63236_;
wire _63237_;
wire _63238_;
wire _63239_;
wire _63240_;
wire _63241_;
wire _63242_;
wire _63243_;
wire _63244_;
wire _63245_;
wire _63246_;
wire _63247_;
wire _63248_;
wire _63249_;
wire _63250_;
wire _63251_;
wire _63252_;
wire _63253_;
wire _63254_;
wire _63255_;
wire _63256_;
wire _63257_;
wire _63258_;
wire _63259_;
wire _63260_;
wire _63261_;
wire _63262_;
wire _63263_;
wire _63264_;
wire _63265_;
wire _63266_;
wire _63267_;
wire _63268_;
wire _63269_;
wire _63270_;
wire _63271_;
wire _63272_;
wire _63273_;
wire _63274_;
wire _63275_;
wire _63276_;
wire _63277_;
wire _63278_;
wire _63279_;
wire _63280_;
wire _63281_;
wire _63282_;
wire _63283_;
wire _63284_;
wire _63285_;
wire _63286_;
wire _63287_;
wire _63288_;
wire _63289_;
wire _63290_;
wire _63291_;
wire _63292_;
wire _63293_;
wire _63294_;
wire _63295_;
wire _63296_;
wire _63297_;
wire _63298_;
wire _63299_;
wire _63300_;
wire _63301_;
wire _63302_;
wire _63303_;
wire _63304_;
wire _63305_;
wire _63306_;
wire _63307_;
wire _63308_;
wire _63309_;
wire _63310_;
wire _63311_;
wire _63312_;
wire _63313_;
wire _63314_;
wire _63315_;
wire _63316_;
wire _63317_;
wire _63318_;
wire _63319_;
wire _63320_;
wire _63321_;
wire _63322_;
wire _63323_;
wire _63324_;
wire _63325_;
wire _63326_;
wire _63327_;
wire _63328_;
wire _63329_;
wire _63330_;
wire _63331_;
wire _63332_;
wire _63333_;
wire _63334_;
wire _63335_;
wire _63336_;
wire _63337_;
wire _63338_;
wire _63339_;
wire _63340_;
wire _63341_;
wire _63342_;
wire _63343_;
wire _63344_;
wire _63345_;
wire _63346_;
wire _63347_;
wire _63348_;
wire _63349_;
wire _63350_;
wire _63351_;
wire _63352_;
wire _63353_;
wire _63354_;
wire _63355_;
wire _63356_;
wire _63357_;
wire _63358_;
wire _63359_;
wire _63360_;
wire _63361_;
wire _63362_;
wire _63363_;
wire _63364_;
wire _63365_;
wire _63366_;
wire _63367_;
wire _63368_;
wire _63369_;
wire _63370_;
wire _63371_;
wire _63372_;
wire _63373_;
wire _63374_;
wire _63375_;
wire _63376_;
wire _63377_;
wire _63378_;
wire _63379_;
wire _63380_;
wire _63381_;
wire _63382_;
wire _63383_;
wire _63384_;
wire _63385_;
wire _63386_;
wire _63387_;
wire _63388_;
wire _63389_;
wire _63390_;
wire _63391_;
wire _63392_;
wire _63393_;
wire _63394_;
wire _63395_;
wire _63396_;
wire _63397_;
wire _63398_;
wire _63399_;
wire _63400_;
wire _63401_;
wire _63402_;
wire _63403_;
wire _63404_;
wire _63405_;
wire _63406_;
wire _63407_;
wire _63408_;
wire _63409_;
wire _63410_;
wire _63411_;
wire _63412_;
wire _63413_;
wire _63414_;
wire _63415_;
wire _63416_;
wire _63417_;
wire _63418_;
wire _63419_;
wire _63420_;
wire _63421_;
wire _63422_;
wire _63423_;
wire _63424_;
wire _63425_;
wire _63426_;
wire _63427_;
wire _63428_;
wire _63429_;
wire _63430_;
wire _63431_;
wire _63432_;
wire _63433_;
wire _63434_;
wire _63435_;
wire _63436_;
wire _63437_;
wire _63438_;
wire _63439_;
wire _63440_;
wire _63441_;
wire _63442_;
wire _63443_;
wire _63444_;
wire _63445_;
wire _63446_;
wire _63447_;
wire _63448_;
wire _63449_;
wire _63450_;
wire _63451_;
wire _63452_;
wire _63453_;
wire _63454_;
wire _63455_;
wire _63456_;
wire _63457_;
wire _63458_;
wire _63459_;
wire _63460_;
wire _63461_;
wire _63462_;
wire _63463_;
wire _63464_;
wire _63465_;
wire _63466_;
wire _63467_;
wire _63468_;
wire _63469_;
wire _63470_;
wire _63471_;
wire _63472_;
wire _63473_;
wire _63474_;
wire _63475_;
wire _63476_;
wire _63477_;
wire _63478_;
wire _63479_;
wire _63480_;
wire _63481_;
wire _63482_;
wire _63483_;
wire _63484_;
wire _63485_;
wire _63486_;
wire _63487_;
wire _63488_;
wire _63489_;
wire _63490_;
wire _63491_;
wire _63492_;
wire _63493_;
wire _63494_;
wire _63495_;
wire _63496_;
wire _63497_;
wire _63498_;
wire _63499_;
wire _63500_;
wire _63501_;
wire _63502_;
wire _63503_;
wire _63504_;
wire _63505_;
wire _63506_;
wire _63507_;
wire _63508_;
wire _63509_;
wire _63510_;
wire _63511_;
wire _63512_;
wire _63513_;
wire _63514_;
wire _63515_;
wire _63516_;
wire _63517_;
wire _63518_;
wire _63519_;
wire _63520_;
wire _63521_;
wire _63522_;
wire _63523_;
wire _63524_;
wire _63525_;
wire _63526_;
wire _63527_;
wire _63528_;
wire _63529_;
wire _63530_;
wire _63531_;
wire _63532_;
wire _63533_;
wire _63534_;
wire _63535_;
wire _63536_;
wire _63537_;
wire _63538_;
wire _63539_;
wire _63540_;
wire _63541_;
wire _63542_;
wire _63543_;
wire _63544_;
wire _63545_;
wire _63546_;
wire _63547_;
wire _63548_;
wire _63549_;
wire _63550_;
wire _63551_;
wire _63552_;
wire _63553_;
wire _63554_;
wire _63555_;
wire _63556_;
wire _63557_;
wire _63558_;
wire _63559_;
wire _63560_;
wire _63561_;
wire _63562_;
wire _63563_;
wire _63564_;
wire _63565_;
wire _63566_;
wire _63567_;
wire _63568_;
wire _63569_;
wire _63570_;
wire _63571_;
wire _63572_;
wire _63573_;
wire _63574_;
wire _63575_;
wire _63576_;
wire _63577_;
wire _63578_;
wire _63579_;
wire _63580_;
wire _63581_;
wire _63582_;
wire _63583_;
wire _63584_;
wire _63585_;
wire _63586_;
wire _63587_;
wire _63588_;
wire _63589_;
wire _63590_;
wire _63591_;
wire _63592_;
wire _63593_;
wire _63594_;
wire _63595_;
wire _63596_;
wire _63597_;
wire _63598_;
wire _63599_;
wire _63600_;
wire _63601_;
wire _63602_;
wire _63603_;
wire _63604_;
wire _63605_;
wire _63606_;
wire _63607_;
wire _63608_;
wire _63609_;
wire _63610_;
wire _63611_;
wire _63612_;
wire _63613_;
wire _63614_;
wire _63615_;
wire _63616_;
wire _63617_;
wire _63618_;
wire _63619_;
wire _63620_;
wire _63621_;
wire _63622_;
wire _63623_;
wire _63624_;
wire _63625_;
wire _63626_;
wire _63627_;
wire _63628_;
wire _63629_;
wire _63630_;
wire _63631_;
wire _63632_;
wire _63633_;
wire _63634_;
wire _63635_;
wire _63636_;
wire _63637_;
wire _63638_;
wire _63639_;
wire _63640_;
wire _63641_;
wire _63642_;
wire _63643_;
wire _63644_;
wire _63645_;
wire _63646_;
wire _63647_;
wire _63648_;
wire _63649_;
wire _63650_;
wire _63651_;
wire _63652_;
wire _63653_;
wire _63654_;
wire _63655_;
wire _63656_;
wire _63657_;
wire _63658_;
wire _63659_;
wire _63660_;
wire _63661_;
wire _63662_;
wire _63663_;
wire _63664_;
wire _63665_;
wire _63666_;
wire _63667_;
wire _63668_;
wire _63669_;
wire _63670_;
wire _63671_;
wire _63672_;
wire _63673_;
wire _63674_;
wire _63675_;
wire _63676_;
wire _63677_;
wire _63678_;
wire _63679_;
wire _63680_;
wire _63681_;
wire _63682_;
wire _63683_;
wire _63684_;
wire _63685_;
wire _63686_;
wire _63687_;
wire _63688_;
wire _63689_;
wire _63690_;
wire _63691_;
wire _63692_;
wire _63693_;
wire _63694_;
wire _63695_;
wire _63696_;
wire _63697_;
wire _63698_;
wire _63699_;
wire _63700_;
wire _63701_;
wire _63702_;
wire _63703_;
wire _63704_;
wire _63705_;
wire _63706_;
wire _63707_;
wire _63708_;
wire _63709_;
wire _63710_;
wire _63711_;
wire _63712_;
wire _63713_;
wire _63714_;
wire _63715_;
wire _63716_;
wire _63717_;
wire _63718_;
wire _63719_;
wire _63720_;
wire _63721_;
wire _63722_;
wire _63723_;
wire _63724_;
wire _63725_;
wire _63726_;
wire _63727_;
wire _63728_;
wire _63729_;
wire _63730_;
wire _63731_;
wire _63732_;
wire _63733_;
wire _63734_;
wire _63735_;
wire _63736_;
wire _63737_;
wire _63738_;
wire _63739_;
wire _63740_;
wire _63741_;
wire _63742_;
wire _63743_;
wire _63744_;
wire _63745_;
wire _63746_;
wire _63747_;
wire _63748_;
wire _63749_;
wire _63750_;
wire _63751_;
wire _63752_;
wire _63753_;
wire _63754_;
wire _63755_;
wire _63756_;
wire _63757_;
wire _63758_;
wire _63759_;
wire _63760_;
wire _63761_;
wire _63762_;
wire _63763_;
wire _63764_;
wire _63765_;
wire _63766_;
wire _63767_;
wire _63768_;
wire _63769_;
wire _63770_;
wire _63771_;
wire _63772_;
wire _63773_;
wire _63774_;
wire _63775_;
wire _63776_;
wire _63777_;
wire _63778_;
wire _63779_;
wire _63780_;
wire _63781_;
wire _63782_;
wire _63783_;
wire _63784_;
wire _63785_;
wire _63786_;
wire _63787_;
wire _63788_;
wire _63789_;
wire _63790_;
wire _63791_;
wire _63792_;
wire _63793_;
wire _63794_;
wire _63795_;
wire _63796_;
wire _63797_;
wire _63798_;
wire _63799_;
wire _63800_;
wire _63801_;
wire _63802_;
wire _63803_;
wire _63804_;
wire _63805_;
wire _63806_;
wire _63807_;
wire _63808_;
wire _63809_;
wire _63810_;
wire _63811_;
wire _63812_;
wire _63813_;
wire _63814_;
wire _63815_;
wire _63816_;
wire _63817_;
wire _63818_;
wire _63819_;
wire _63820_;
wire _63821_;
wire _63822_;
wire _63823_;
wire _63824_;
wire _63825_;
wire _63826_;
wire _63827_;
wire _63828_;
wire _63829_;
wire _63830_;
wire _63831_;
wire _63832_;
wire _63833_;
wire _63834_;
wire _63835_;
wire _63836_;
wire _63837_;
wire _63838_;
wire _63839_;
wire _63840_;
wire _63841_;
wire _63842_;
wire _63843_;
wire _63844_;
wire _63845_;
wire _63846_;
wire _63847_;
wire _63848_;
wire _63849_;
wire _63850_;
wire _63851_;
wire _63852_;
wire _63853_;
wire _63854_;
wire _63855_;
wire _63856_;
wire _63857_;
wire _63858_;
wire _63859_;
wire _63860_;
wire _63861_;
wire _63862_;
wire _63863_;
wire _63864_;
wire _63865_;
wire _63866_;
wire _63867_;
wire _63868_;
wire _63869_;
wire _63870_;
wire _63871_;
wire _63872_;
wire _63873_;
wire _63874_;
wire _63875_;
wire _63876_;
wire _63877_;
wire _63878_;
wire _63879_;
wire _63880_;
wire _63881_;
wire _63882_;
wire _63883_;
wire _63884_;
wire _63885_;
wire _63886_;
wire _63887_;
wire _63888_;
wire _63889_;
wire _63890_;
wire _63891_;
wire _63892_;
wire _63893_;
wire _63894_;
wire _63895_;
wire _63896_;
wire _63897_;
wire _63898_;
wire _63899_;
wire _63900_;
wire _63901_;
wire _63902_;
wire _63903_;
wire _63904_;
wire _63905_;
wire _63906_;
wire _63907_;
wire _63908_;
wire _63909_;
wire _63910_;
wire _63911_;
wire _63912_;
wire _63913_;
wire _63914_;
wire _63915_;
wire _63916_;
wire _63917_;
wire _63918_;
wire _63919_;
wire _63920_;
wire _63921_;
wire _63922_;
wire _63923_;
wire _63924_;
wire _63925_;
wire _63926_;
wire _63927_;
wire _63928_;
wire _63929_;
wire _63930_;
wire _63931_;
wire _63932_;
wire _63933_;
wire _63934_;
wire _63935_;
wire _63936_;
wire _63937_;
wire _63938_;
wire _63939_;
wire _63940_;
wire _63941_;
wire _63942_;
wire _63943_;
wire _63944_;
wire _63945_;
wire _63946_;
wire _63947_;
wire _63948_;
wire _63949_;
wire _63950_;
wire _63951_;
wire _63952_;
wire _63953_;
wire _63954_;
wire _63955_;
wire _63956_;
wire _63957_;
wire _63958_;
wire _63959_;
wire _63960_;
wire _63961_;
wire _63962_;
wire _63963_;
wire _63964_;
wire _63965_;
wire _63966_;
wire _63967_;
wire _63968_;
wire _63969_;
wire _63970_;
wire _63971_;
wire _63972_;
wire _63973_;
wire _63974_;
wire _63975_;
wire _63976_;
wire _63977_;
wire _63978_;
wire _63979_;
wire _63980_;
wire _63981_;
wire _63982_;
wire _63983_;
wire _63984_;
wire _63985_;
wire _63986_;
wire _63987_;
wire _63988_;
wire _63989_;
wire _63990_;
wire _63991_;
wire _63992_;
wire _63993_;
wire _63994_;
wire _63995_;
wire _63996_;
wire _63997_;
wire _63998_;
wire _63999_;
wire _64000_;
wire _64001_;
wire _64002_;
wire _64003_;
wire _64004_;
wire _64005_;
wire _64006_;
wire _64007_;
wire _64008_;
wire _64009_;
wire _64010_;
wire _64011_;
wire _64012_;
wire _64013_;
wire _64014_;
wire _64015_;
wire _64016_;
wire _64017_;
wire _64018_;
wire _64019_;
wire _64020_;
wire _64021_;
wire _64022_;
wire _64023_;
wire _64024_;
wire _64025_;
wire _64026_;
wire _64027_;
wire _64028_;
wire _64029_;
wire _64030_;
wire _64031_;
wire _64032_;
wire _64033_;
wire _64034_;
wire _64035_;
wire _64036_;
wire _64037_;
wire _64038_;
wire _64039_;
wire _64040_;
wire _64041_;
wire _64042_;
wire _64043_;
wire _64044_;
wire _64045_;
wire _64046_;
wire _64047_;
wire _64048_;
wire _64049_;
wire _64050_;
wire _64051_;
wire _64052_;
wire _64053_;
wire _64054_;
wire _64055_;
wire _64056_;
wire _64057_;
wire _64058_;
wire _64059_;
wire _64060_;
wire _64061_;
wire _64062_;
wire _64063_;
wire _64064_;
wire _64065_;
wire _64066_;
wire _64067_;
wire _64068_;
wire _64069_;
wire _64070_;
wire _64071_;
wire _64072_;
wire _64073_;
wire _64074_;
wire _64075_;
wire _64076_;
wire _64077_;
wire _64078_;
wire _64079_;
wire _64080_;
wire _64081_;
wire _64082_;
wire _64083_;
wire _64084_;
wire _64085_;
wire _64086_;
wire _64087_;
wire _64088_;
wire _64089_;
wire _64090_;
wire _64091_;
wire _64092_;
wire _64093_;
wire _64094_;
wire _64095_;
wire _64096_;
wire _64097_;
wire _64098_;
wire _64099_;
wire _64100_;
wire _64101_;
wire _64102_;
wire _64103_;
wire _64104_;
wire _64105_;
wire _64106_;
wire _64107_;
wire _64108_;
wire _64109_;
wire _64110_;
wire _64111_;
wire _64112_;
wire _64113_;
wire _64114_;
wire _64115_;
wire _64116_;
wire _64117_;
wire _64118_;
wire _64119_;
wire _64120_;
wire _64121_;
wire _64122_;
wire _64123_;
wire _64124_;
wire _64125_;
wire _64126_;
wire _64127_;
wire _64128_;
wire _64129_;
wire _64130_;
wire _64131_;
wire _64132_;
wire _64133_;
wire _64134_;
wire _64135_;
wire _64136_;
wire _64137_;
wire _64138_;
wire _64139_;
wire _64140_;
wire _64141_;
wire _64142_;
wire _64143_;
wire _64144_;
wire _64145_;
wire _64146_;
wire _64147_;
wire _64148_;
wire _64149_;
wire _64150_;
wire _64151_;
wire _64152_;
wire _64153_;
wire _64154_;
wire _64155_;
wire _64156_;
wire _64157_;
wire _64158_;
wire _64159_;
wire _64160_;
wire _64161_;
wire _64162_;
wire _64163_;
wire _64164_;
wire _64165_;
wire _64166_;
wire _64167_;
wire _64168_;
wire _64169_;
wire _64170_;
wire _64171_;
wire _64172_;
wire _64173_;
wire _64174_;
wire _64175_;
wire _64176_;
wire _64177_;
wire _64178_;
wire _64179_;
wire _64180_;
wire _64181_;
wire _64182_;
wire _64183_;
wire _64184_;
wire _64185_;
wire _64186_;
wire _64187_;
wire _64188_;
wire _64189_;
wire _64190_;
wire _64191_;
wire _64192_;
wire _64193_;
wire _64194_;
wire _64195_;
wire _64196_;
wire _64197_;
wire _64198_;
wire _64199_;
wire _64200_;
wire _64201_;
wire _64202_;
wire _64203_;
wire _64204_;
wire _64205_;
wire _64206_;
wire _64207_;
wire _64208_;
wire _64209_;
wire _64210_;
wire _64211_;
wire _64212_;
wire _64213_;
wire _64214_;
wire _64215_;
wire _64216_;
wire _64217_;
wire _64218_;
wire _64219_;
wire _64220_;
wire _64221_;
wire _64222_;
wire _64223_;
wire _64224_;
wire _64225_;
wire _64226_;
wire _64227_;
wire _64228_;
wire _64229_;
wire _64230_;
wire _64231_;
wire _64232_;
wire _64233_;
wire _64234_;
wire _64235_;
wire _64236_;
wire _64237_;
wire _64238_;
wire _64239_;
wire _64240_;
wire _64241_;
wire _64242_;
wire _64243_;
wire _64244_;
wire _64245_;
wire _64246_;
wire _64247_;
wire _64248_;
wire _64249_;
wire _64250_;
wire _64251_;
wire _64252_;
wire _64253_;
wire _64254_;
wire _64255_;
wire _64256_;
wire _64257_;
wire _64258_;
wire _64259_;
wire _64260_;
wire _64261_;
wire _64262_;
wire _64263_;
wire _64264_;
wire _64265_;
wire _64266_;
wire _64267_;
wire _64268_;
wire _64269_;
wire _64270_;
wire _64271_;
wire _64272_;
wire _64273_;
wire _64274_;
wire _64275_;
wire _64276_;
wire _64277_;
wire _64278_;
wire _64279_;
wire _64280_;
wire _64281_;
wire _64282_;
wire _64283_;
wire _64284_;
wire _64285_;
wire _64286_;
wire _64287_;
wire _64288_;
wire _64289_;
wire _64290_;
wire _64291_;
wire _64292_;
wire _64293_;
wire _64294_;
wire _64295_;
wire _64296_;
wire _64297_;
wire _64298_;
wire _64299_;
wire _64300_;
wire _64301_;
wire _64302_;
wire _64303_;
wire _64304_;
wire _64305_;
wire _64306_;
wire _64307_;
wire _64308_;
wire _64309_;
wire _64310_;
wire _64311_;
wire _64312_;
wire _64313_;
wire _64314_;
wire _64315_;
wire _64316_;
wire _64317_;
wire _64318_;
wire _64319_;
wire _64320_;
wire _64321_;
wire _64322_;
wire _64323_;
wire _64324_;
wire _64325_;
wire _64326_;
wire _64327_;
wire _64328_;
wire _64329_;
wire _64330_;
wire _64331_;
wire _64332_;
wire _64333_;
wire _64334_;
wire _64335_;
wire _64336_;
wire _64337_;
wire _64338_;
wire _64339_;
wire _64340_;
wire _64341_;
wire _64342_;
wire _64343_;
wire _64344_;
wire _64345_;
wire _64346_;
wire _64347_;
wire _64348_;
wire _64349_;
wire _64350_;
wire _64351_;
wire _64352_;
wire _64353_;
wire _64354_;
wire _64355_;
wire _64356_;
wire _64357_;
wire _64358_;
wire _64359_;
wire _64360_;
wire _64361_;
wire _64362_;
wire _64363_;
wire _64364_;
wire _64365_;
wire _64366_;
wire _64367_;
wire _64368_;
wire _64369_;
wire _64370_;
wire _64371_;
wire _64372_;
wire _64373_;
wire _64374_;
wire _64375_;
wire _64376_;
wire _64377_;
wire _64378_;
wire _64379_;
wire _64380_;
wire _64381_;
wire _64382_;
wire _64383_;
wire _64384_;
wire _64385_;
wire _64386_;
wire _64387_;
wire _64388_;
wire _64389_;
wire _64390_;
wire _64391_;
wire _64392_;
wire _64393_;
wire _64394_;
wire _64395_;
wire _64396_;
wire _64397_;
wire _64398_;
wire _64399_;
wire _64400_;
wire _64401_;
wire _64402_;
wire _64403_;
wire _64404_;
wire _64405_;
wire _64406_;
wire _64407_;
wire _64408_;
wire _64409_;
wire _64410_;
wire _64411_;
wire _64412_;
wire _64413_;
wire _64414_;
wire _64415_;
wire _64416_;
wire _64417_;
wire _64418_;
wire _64419_;
wire _64420_;
wire _64421_;
wire _64422_;
wire _64423_;
wire _64424_;
wire _64425_;
wire _64426_;
wire _64427_;
wire _64428_;
wire _64429_;
wire _64430_;
wire _64431_;
wire _64432_;
wire _64433_;
wire _64434_;
wire _64435_;
wire _64436_;
wire _64437_;
wire _64438_;
wire _64439_;
wire _64440_;
wire _64441_;
wire _64442_;
wire _64443_;
wire _64444_;
wire _64445_;
wire _64446_;
wire _64447_;
wire _64448_;
wire _64449_;
wire _64450_;
wire _64451_;
wire _64452_;
wire _64453_;
wire _64454_;
wire _64455_;
wire _64456_;
wire _64457_;
wire _64458_;
wire _64459_;
wire _64460_;
wire _64461_;
wire _64462_;
wire _64463_;
wire _64464_;
wire _64465_;
wire _64466_;
wire _64467_;
wire _64468_;
wire _64469_;
wire _64470_;
wire _64471_;
wire _64472_;
wire _64473_;
wire _64474_;
wire _64475_;
wire _64476_;
wire _64477_;
wire _64478_;
wire _64479_;
wire _64480_;
wire _64481_;
wire _64482_;
wire _64483_;
wire _64484_;
wire _64485_;
wire _64486_;
wire _64487_;
wire _64488_;
wire _64489_;
wire _64490_;
wire _64491_;
wire _64492_;
wire _64493_;
wire _64494_;
wire _64495_;
wire _64496_;
wire _64497_;
wire _64498_;
wire _64499_;
wire _64500_;
wire _64501_;
wire _64502_;
wire _64503_;
wire _64504_;
wire _64505_;
wire _64506_;
wire _64507_;
wire _64508_;
wire _64509_;
wire _64510_;
wire _64511_;
wire _64512_;
wire _64513_;
wire _64514_;
wire _64515_;
wire _64516_;
wire _64517_;
wire _64518_;
wire _64519_;
wire _64520_;
wire _64521_;
wire _64522_;
wire _64523_;
wire _64524_;
wire _64525_;
wire _64526_;
wire _64527_;
wire _64528_;
wire _64529_;
wire _64530_;
wire _64531_;
wire _64532_;
wire _64533_;
wire _64534_;
wire _64535_;
wire _64536_;
wire _64537_;
wire _64538_;
wire _64539_;
wire _64540_;
wire _64541_;
wire _64542_;
wire _64543_;
wire _64544_;
wire _64545_;
wire _64546_;
wire _64547_;
wire _64548_;
wire _64549_;
wire _64550_;
wire _64551_;
wire _64552_;
wire _64553_;
wire _64554_;
wire _64555_;
wire _64556_;
wire _64557_;
wire _64558_;
wire _64559_;
wire _64560_;
wire _64561_;
wire _64562_;
wire _64563_;
wire _64564_;
wire _64565_;
wire _64566_;
wire _64567_;
wire _64568_;
wire _64569_;
wire _64570_;
wire _64571_;
wire _64572_;
wire _64573_;
wire _64574_;
wire _64575_;
wire _64576_;
wire _64577_;
wire _64578_;
wire _64579_;
wire _64580_;
wire _64581_;
wire _64582_;
wire _64583_;
wire _64584_;
wire _64585_;
wire _64586_;
wire _64587_;
wire _64588_;
wire _64589_;
wire _64590_;
wire _64591_;
wire _64592_;
wire _64593_;
wire _64594_;
wire _64595_;
wire _64596_;
wire _64597_;
wire _64598_;
wire _64599_;
wire _64600_;
wire _64601_;
wire _64602_;
wire _64603_;
wire _64604_;
wire _64605_;
wire _64606_;
wire _64607_;
wire _64608_;
wire _64609_;
wire _64610_;
wire _64611_;
wire _64612_;
wire _64613_;
wire _64614_;
wire _64615_;
wire _64616_;
wire _64617_;
wire _64618_;
wire _64619_;
wire _64620_;
wire _64621_;
wire _64622_;
wire _64623_;
wire _64624_;
wire _64625_;
wire _64626_;
wire _64627_;
wire _64628_;
wire _64629_;
wire _64630_;
wire _64631_;
wire _64632_;
wire _64633_;
wire _64634_;
wire _64635_;
wire _64636_;
wire _64637_;
wire _64638_;
wire _64639_;
wire _64640_;
wire _64641_;
wire _64642_;
wire _64643_;
wire _64644_;
wire _64645_;
wire _64646_;
wire _64647_;
wire _64648_;
wire _64649_;
wire _64650_;
wire _64651_;
wire _64652_;
wire _64653_;
wire _64654_;
wire _64655_;
wire _64656_;
wire _64657_;
wire _64658_;
wire _64659_;
wire _64660_;
wire _64661_;
wire _64662_;
wire _64663_;
wire _64664_;
wire _64665_;
wire _64666_;
wire _64667_;
wire _64668_;
wire _64669_;
wire _64670_;
wire _64671_;
wire _64672_;
wire _64673_;
wire _64674_;
wire _64675_;
wire _64676_;
wire _64677_;
wire _64678_;
wire _64679_;
wire _64680_;
wire _64681_;
wire _64682_;
wire _64683_;
wire _64684_;
wire _64685_;
wire _64686_;
wire _64687_;
wire _64688_;
wire _64689_;
wire _64690_;
wire _64691_;
wire _64692_;
wire _64693_;
wire _64694_;
wire _64695_;
wire _64696_;
wire _64697_;
wire _64698_;
wire _64699_;
wire _64700_;
wire _64701_;
wire _64702_;
wire _64703_;
wire _64704_;
wire _64705_;
wire _64706_;
wire _64707_;
wire _64708_;
wire _64709_;
wire _64710_;
wire _64711_;
wire _64712_;
wire _64713_;
wire _64714_;
wire _64715_;
wire _64716_;
wire _64717_;
wire _64718_;
wire _64719_;
wire _64720_;
wire _64721_;
wire _64722_;
wire _64723_;
wire _64724_;
wire _64725_;
wire _64726_;
wire _64727_;
wire _64728_;
wire _64729_;
wire _64730_;
wire _64731_;
wire _64732_;
wire _64733_;
wire _64734_;
wire _64735_;
wire _64736_;
wire _64737_;
wire _64738_;
wire _64739_;
wire _64740_;
wire _64741_;
wire _64742_;
wire _64743_;
wire _64744_;
wire _64745_;
wire _64746_;
wire _64747_;
wire _64748_;
wire _64749_;
wire _64750_;
wire _64751_;
wire _64752_;
wire _64753_;
wire _64754_;
wire _64755_;
wire _64756_;
wire _64757_;
wire _64758_;
wire _64759_;
wire _64760_;
wire _64761_;
wire _64762_;
wire _64763_;
wire _64764_;
wire _64765_;
wire _64766_;
wire _64767_;
wire _64768_;
wire _64769_;
wire _64770_;
wire _64771_;
wire _64772_;
wire _64773_;
wire _64774_;
wire _64775_;
wire _64776_;
wire _64777_;
wire _64778_;
wire _64779_;
wire _64780_;
wire _64781_;
wire _64782_;
wire _64783_;
wire _64784_;
wire _64785_;
wire _64786_;
wire _64787_;
wire _64788_;
wire _64789_;
wire _64790_;
wire _64791_;
wire _64792_;
wire _64793_;
wire _64794_;
wire _64795_;
wire _64796_;
wire _64797_;
wire _64798_;
wire _64799_;
wire _64800_;
wire _64801_;
wire _64802_;
wire _64803_;
wire _64804_;
wire _64805_;
wire _64806_;
wire _64807_;
wire _64808_;
wire _64809_;
wire _64810_;
wire _64811_;
wire _64812_;
wire _64813_;
wire _64814_;
wire _64815_;
wire _64816_;
wire _64817_;
wire _64818_;
wire _64819_;
wire _64820_;
wire _64821_;
wire _64822_;
wire _64823_;
wire _64824_;
wire _64825_;
wire _64826_;
wire _64827_;
wire _64828_;
wire _64829_;
wire _64830_;
wire _64831_;
wire _64832_;
wire _64833_;
wire _64834_;
wire _64835_;
wire _64836_;
wire _64837_;
wire _64838_;
wire _64839_;
wire _64840_;
wire _64841_;
wire _64842_;
wire _64843_;
wire _64844_;
wire _64845_;
wire _64846_;
wire _64847_;
wire _64848_;
wire _64849_;
wire _64850_;
wire _64851_;
wire _64852_;
wire _64853_;
wire _64854_;
wire _64855_;
wire _64856_;
wire _64857_;
wire _64858_;
wire _64859_;
wire _64860_;
wire _64861_;
wire _64862_;
wire _64863_;
wire _64864_;
wire _64865_;
wire _64866_;
wire _64867_;
wire _64868_;
wire _64869_;
wire _64870_;
wire _64871_;
wire _64872_;
wire _64873_;
wire _64874_;
wire _64875_;
wire _64876_;
wire _64877_;
wire _64878_;
wire _64879_;
wire _64880_;
wire _64881_;
wire _64882_;
wire _64883_;
wire _64884_;
wire _64885_;
wire _64886_;
wire _64887_;
wire _64888_;
wire _64889_;
wire _64890_;
wire _64891_;
wire _64892_;
wire _64893_;
wire _64894_;
wire _64895_;
wire _64896_;
wire _64897_;
wire _64898_;
wire _64899_;
wire _64900_;
wire _64901_;
wire _64902_;
wire _64903_;
wire _64904_;
wire _64905_;
wire _64906_;
wire _64907_;
wire _64908_;
wire _64909_;
wire _64910_;
wire _64911_;
wire _64912_;
wire _64913_;
wire _64914_;
wire _64915_;
wire _64916_;
wire _64917_;
wire _64918_;
wire _64919_;
wire _64920_;
wire _64921_;
wire _64922_;
wire _64923_;
wire _64924_;
wire _64925_;
wire _64926_;
wire _64927_;
wire _64928_;
wire _64929_;
wire _64930_;
wire _64931_;
wire _64932_;
wire _64933_;
wire _64934_;
wire _64935_;
wire _64936_;
wire _64937_;
wire _64938_;
wire _64939_;
wire _64940_;
wire _64941_;
wire _64942_;
wire _64943_;
wire _64944_;
wire _64945_;
wire _64946_;
wire _64947_;
wire _64948_;
wire _64949_;
wire _64950_;
wire _64951_;
wire _64952_;
wire _64953_;
wire _64954_;
wire _64955_;
wire _64956_;
wire _64957_;
wire _64958_;
wire _64959_;
wire _64960_;
wire _64961_;
wire _64962_;
wire _64963_;
wire _64964_;
wire _64965_;
wire _64966_;
wire _64967_;
wire _64968_;
wire _64969_;
wire _64970_;
wire _64971_;
wire _64972_;
wire _64973_;
wire _64974_;
wire _64975_;
wire _64976_;
wire _64977_;
wire _64978_;
wire _64979_;
wire _64980_;
wire _64981_;
wire _64982_;
wire _64983_;
wire _64984_;
wire _64985_;
wire _64986_;
wire _64987_;
wire _64988_;
wire _64989_;
wire _64990_;
wire _64991_;
wire _64992_;
wire _64993_;
wire _64994_;
wire _64995_;
wire _64996_;
wire _64997_;
wire _64998_;
wire _64999_;
wire _65000_;
wire _65001_;
wire _65002_;
wire _65003_;
wire _65004_;
wire _65005_;
wire _65006_;
wire _65007_;
wire _65008_;
wire _65009_;
wire _65010_;
wire _65011_;
wire _65012_;
wire _65013_;
wire _65014_;
wire _65015_;
wire _65016_;
wire _65017_;
wire _65018_;
wire _65019_;
wire _65020_;
wire _65021_;
wire _65022_;
wire _65023_;
wire _65024_;
wire _65025_;
wire _65026_;
wire _65027_;
wire _65028_;
wire _65029_;
wire _65030_;
wire _65031_;
wire _65032_;
wire _65033_;
wire _65034_;
wire _65035_;
wire _65036_;
wire _65037_;
wire _65038_;
wire _65039_;
wire _65040_;
wire _65041_;
wire _65042_;
wire _65043_;
wire _65044_;
wire _65045_;
wire _65046_;
wire _65047_;
wire _65048_;
wire _65049_;
wire _65050_;
wire _65051_;
wire _65052_;
wire _65053_;
wire _65054_;
wire _65055_;
wire _65056_;
wire _65057_;
wire _65058_;
wire _65059_;
wire _65060_;
wire _65061_;
wire _65062_;
wire _65063_;
wire _65064_;
wire _65065_;
wire _65066_;
wire _65067_;
wire _65068_;
wire _65069_;
wire _65070_;
wire _65071_;
wire _65072_;
wire _65073_;
wire _65074_;
wire _65075_;
wire _65076_;
wire _65077_;
wire _65078_;
wire _65079_;
wire _65080_;
wire _65081_;
wire _65082_;
wire _65083_;
wire _65084_;
wire _65085_;
wire _65086_;
wire _65087_;
wire _65088_;
wire _65089_;
wire _65090_;
wire _65091_;
wire _65092_;
wire _65093_;
wire _65094_;
wire _65095_;
wire _65096_;
wire _65097_;
wire _65098_;
wire _65099_;
wire _65100_;
wire _65101_;
wire _65102_;
wire _65103_;
wire _65104_;
wire _65105_;
wire _65106_;
wire _65107_;
wire _65108_;
wire _65109_;
wire _65110_;
wire _65111_;
wire _65112_;
wire _65113_;
wire _65114_;
wire _65115_;
wire _65116_;
wire _65117_;
wire _65118_;
wire _65119_;
wire _65120_;
wire _65121_;
wire _65122_;
wire _65123_;
wire _65124_;
wire _65125_;
wire _65126_;
wire _65127_;
wire _65128_;
wire _65129_;
wire _65130_;
wire _65131_;
wire _65132_;
wire _65133_;
wire _65134_;
wire _65135_;
wire _65136_;
wire _65137_;
wire _65138_;
wire _65139_;
wire _65140_;
wire _65141_;
wire _65142_;
wire _65143_;
wire _65144_;
wire _65145_;
wire _65146_;
wire _65147_;
wire _65148_;
wire _65149_;
wire _65150_;
wire _65151_;
wire _65152_;
wire _65153_;
wire _65154_;
wire _65155_;
wire _65156_;
wire _65157_;
wire _65158_;
wire _65159_;
wire _65160_;
wire _65161_;
wire _65162_;
wire _65163_;
wire _65164_;
wire _65165_;
wire _65166_;
wire _65167_;
wire _65168_;
wire _65169_;
wire _65170_;
wire _65171_;
wire _65172_;
wire _65173_;
wire _65174_;
wire _65175_;
wire _65176_;
wire _65177_;
wire _65178_;
wire _65179_;
wire _65180_;
wire _65181_;
wire _65182_;
wire _65183_;
wire _65184_;
wire _65185_;
wire _65186_;
wire _65187_;
wire _65188_;
wire _65189_;
wire _65190_;
wire _65191_;
wire _65192_;
wire _65193_;
wire _65194_;
wire _65195_;
wire _65196_;
wire _65197_;
wire _65198_;
wire _65199_;
wire _65200_;
wire _65201_;
wire _65202_;
wire _65203_;
wire _65204_;
wire _65205_;
wire _65206_;
wire _65207_;
wire _65208_;
wire _65209_;
wire _65210_;
wire _65211_;
wire _65212_;
wire _65213_;
wire _65214_;
wire _65215_;
wire _65216_;
wire _65217_;
wire _65218_;
wire _65219_;
wire _65220_;
wire _65221_;
wire _65222_;
wire _65223_;
wire _65224_;
wire _65225_;
wire _65226_;
wire _65227_;
wire _65228_;
wire _65229_;
wire _65230_;
wire _65231_;
wire _65232_;
wire _65233_;
wire _65234_;
wire _65235_;
wire _65236_;
wire _65237_;
wire _65238_;
wire _65239_;
wire _65240_;
wire _65241_;
wire _65242_;
wire _65243_;
wire _65244_;
wire _65245_;
wire _65246_;
wire _65247_;
wire _65248_;
wire _65249_;
wire _65250_;
wire _65251_;
wire _65252_;
wire _65253_;
wire _65254_;
wire _65255_;
wire _65256_;
wire _65257_;
wire _65258_;
wire _65259_;
wire _65260_;
wire _65261_;
wire _65262_;
wire _65263_;
wire _65264_;
wire _65265_;
wire _65266_;
wire _65267_;
wire _65268_;
wire _65269_;
wire _65270_;
wire _65271_;
wire _65272_;
wire _65273_;
wire _65274_;
wire _65275_;
wire _65276_;
wire _65277_;
wire _65278_;
wire _65279_;
wire _65280_;
wire _65281_;
wire _65282_;
wire _65283_;
wire _65284_;
wire _65285_;
wire _65286_;
wire _65287_;
wire _65288_;
wire _65289_;
wire _65290_;
wire _65291_;
wire _65292_;
wire _65293_;
wire _65294_;
wire _65295_;
wire _65296_;
wire _65297_;
wire _65298_;
wire _65299_;
wire _65300_;
wire _65301_;
wire _65302_;
wire _65303_;
wire _65304_;
wire _65305_;
wire _65306_;
wire _65307_;
wire _65308_;
wire _65309_;
wire _65310_;
wire _65311_;
wire _65312_;
wire _65313_;
wire _65314_;
wire _65315_;
wire _65316_;
wire _65317_;
wire _65318_;
wire _65319_;
wire _65320_;
wire _65321_;
wire _65322_;
wire _65323_;
wire _65324_;
wire _65325_;
wire _65326_;
wire _65327_;
wire _65328_;
wire _65329_;
wire _65330_;
wire _65331_;
wire _65332_;
wire _65333_;
wire _65334_;
wire _65335_;
wire _65336_;
wire _65337_;
wire _65338_;
wire _65339_;
wire _65340_;
wire _65341_;
wire _65342_;
wire _65343_;
wire _65344_;
wire _65345_;
wire _65346_;
wire _65347_;
wire _65348_;
wire _65349_;
wire _65350_;
wire _65351_;
wire _65352_;
wire _65353_;
wire _65354_;
wire _65355_;
wire _65356_;
wire _65357_;
wire _65358_;
wire _65359_;
wire _65360_;
wire _65361_;
wire _65362_;
wire _65363_;
wire _65364_;
wire _65365_;
wire _65366_;
wire _65367_;
wire _65368_;
wire _65369_;
wire _65370_;
wire _65371_;
wire _65372_;
wire _65373_;
wire _65374_;
wire _65375_;
wire _65376_;
wire _65377_;
wire _65378_;
wire _65379_;
wire _65380_;
wire _65381_;
wire _65382_;
wire _65383_;
wire _65384_;
wire _65385_;
wire _65386_;
wire _65387_;
wire _65388_;
wire _65389_;
wire _65390_;
wire _65391_;
wire _65392_;
wire _65393_;
wire _65394_;
wire _65395_;
wire _65396_;
wire _65397_;
wire _65398_;
wire _65399_;
wire _65400_;
wire _65401_;
wire _65402_;
wire _65403_;
wire _65404_;
wire _65405_;
wire _65406_;
wire _65407_;
wire _65408_;
wire _65409_;
wire _65410_;
wire _65411_;
wire _65412_;
wire _65413_;
wire _65414_;
wire _65415_;
wire _65416_;
wire _65417_;
wire _65418_;
wire _65419_;
wire _65420_;
wire _65421_;
wire _65422_;
wire _65423_;
wire _65424_;
wire _65425_;
wire _65426_;
wire _65427_;
wire _65428_;
wire _65429_;
wire _65430_;
wire _65431_;
wire _65432_;
wire _65433_;
wire _65434_;
wire _65435_;
wire _65436_;
wire _65437_;
wire _65438_;
wire _65439_;
wire _65440_;
wire _65441_;
wire _65442_;
wire _65443_;
wire _65444_;
wire _65445_;
wire _65446_;
wire _65447_;
wire _65448_;
wire _65449_;
wire _65450_;
wire _65451_;
wire _65452_;
wire _65453_;
wire _65454_;
wire _65455_;
wire _65456_;
wire _65457_;
wire _65458_;
wire _65459_;
wire _65460_;
wire _65461_;
wire _65462_;
wire _65463_;
wire _65464_;
wire _65465_;
wire _65466_;
wire _65467_;
wire _65468_;
wire _65469_;
wire _65470_;
wire _65471_;
wire _65472_;
wire _65473_;
wire _65474_;
wire _65475_;
wire _65476_;
wire _65477_;
wire _65478_;
wire _65479_;
wire _65480_;
wire _65481_;
wire _65482_;
wire _65483_;
wire _65484_;
wire _65485_;
wire _65486_;
wire _65487_;
wire _65488_;
wire _65489_;
wire _65490_;
wire _65491_;
wire _65492_;
wire _65493_;
wire _65494_;
wire _65495_;
wire _65496_;
wire _65497_;
wire _65498_;
wire _65499_;
wire _65500_;
wire _65501_;
wire _65502_;
wire _65503_;
wire _65504_;
wire _65505_;
wire _65506_;
wire _65507_;
wire _65508_;
wire _65509_;
wire _65510_;
wire _65511_;
wire _65512_;
wire _65513_;
wire _65514_;
wire _65515_;
wire _65516_;
wire _65517_;
wire _65518_;
wire _65519_;
wire _65520_;
wire _65521_;
wire _65522_;
wire _65523_;
wire _65524_;
wire _65525_;
wire _65526_;
wire _65527_;
wire _65528_;
wire _65529_;
wire _65530_;
wire _65531_;
wire _65532_;
wire _65533_;
wire _65534_;
wire _65535_;
wire _65536_;
wire _65537_;
wire _65538_;
wire _65539_;
wire _65540_;
wire _65541_;
wire _65542_;
wire _65543_;
wire _65544_;
wire _65545_;
wire _65546_;
wire _65547_;
wire _65548_;
wire _65549_;
wire _65550_;
wire _65551_;
wire _65552_;
wire _65553_;
wire _65554_;
wire _65555_;
wire _65556_;
wire _65557_;
wire _65558_;
wire _65559_;
wire _65560_;
wire _65561_;
wire _65562_;
wire _65563_;
wire _65564_;
wire _65565_;
wire _65566_;
wire _65567_;
wire _65568_;
wire _65569_;
wire _65570_;
wire _65571_;
wire _65572_;
wire _65573_;
wire _65574_;
wire _65575_;
wire _65576_;
wire _65577_;
wire _65578_;
wire _65579_;
wire _65580_;
wire _65581_;
wire _65582_;
wire _65583_;
wire _65584_;
wire _65585_;
wire _65586_;
wire _65587_;
wire _65588_;
wire _65589_;
wire _65590_;
wire _65591_;
wire _65592_;
wire _65593_;
wire _65594_;
wire _65595_;
wire _65596_;
wire _65597_;
wire _65598_;
wire _65599_;
wire _65600_;
wire _65601_;
wire _65602_;
wire _65603_;
wire _65604_;
wire _65605_;
wire _65606_;
wire _65607_;
wire _65608_;
wire _65609_;
wire _65610_;
wire _65611_;
wire _65612_;
wire _65613_;
wire _65614_;
wire _65615_;
wire _65616_;
wire _65617_;
wire _65618_;
wire _65619_;
wire _65620_;
wire _65621_;
wire _65622_;
wire _65623_;
wire _65624_;
wire _65625_;
wire _65626_;
wire _65627_;
wire _65628_;
wire _65629_;
wire _65630_;
wire _65631_;
wire _65632_;
wire _65633_;
wire _65634_;
wire _65635_;
wire _65636_;
wire _65637_;
wire _65638_;
wire _65639_;
wire _65640_;
wire _65641_;
wire _65642_;
wire _65643_;
wire _65644_;
wire _65645_;
wire _65646_;
wire _65647_;
wire _65648_;
wire _65649_;
wire _65650_;
wire _65651_;
wire _65652_;
wire _65653_;
wire _65654_;
wire _65655_;
wire _65656_;
wire _65657_;
wire _65658_;
wire _65659_;
wire _65660_;
wire _65661_;
wire _65662_;
wire _65663_;
wire _65664_;
wire _65665_;
wire _65666_;
wire _65667_;
wire _65668_;
wire _65669_;
wire _65670_;
wire _65671_;
wire _65672_;
wire _65673_;
wire _65674_;
wire _65675_;
wire _65676_;
wire _65677_;
wire _65678_;
wire _65679_;
wire _65680_;
wire _65681_;
wire _65682_;
wire _65683_;
wire _65684_;
wire _65685_;
wire _65686_;
wire _65687_;
wire _65688_;
wire _65689_;
wire _65690_;
wire _65691_;
wire _65692_;
wire _65693_;
wire _65694_;
wire _65695_;
wire _65696_;
wire _65697_;
wire _65698_;
wire _65699_;
wire _65700_;
wire _65701_;
wire _65702_;
wire _65703_;
wire _65704_;
wire _65705_;
wire _65706_;
wire _65707_;
wire _65708_;
wire _65709_;
wire _65710_;
wire _65711_;
wire _65712_;
wire _65713_;
wire _65714_;
wire _65715_;
wire _65716_;
wire _65717_;
wire _65718_;
wire _65719_;
wire _65720_;
wire _65721_;
wire _65722_;
wire _65723_;
wire _65724_;
wire _65725_;
wire _65726_;
wire _65727_;
wire _65728_;
wire _65729_;
wire _65730_;
wire _65731_;
wire _65732_;
wire _65733_;
wire _65734_;
wire _65735_;
wire _65736_;
wire _65737_;
wire _65738_;
wire _65739_;
wire _65740_;
wire _65741_;
wire _65742_;
wire _65743_;
wire _65744_;
wire _65745_;
wire _65746_;
wire _65747_;
wire _65748_;
wire _65749_;
wire _65750_;
wire _65751_;
wire _65752_;
wire _65753_;
wire _65754_;
wire _65755_;
wire _65756_;
wire _65757_;
wire _65758_;
wire _65759_;
wire _65760_;
wire _65761_;
wire _65762_;
wire _65763_;
wire _65764_;
wire _65765_;
wire _65766_;
wire _65767_;
wire _65768_;
wire _65769_;
wire _65770_;
wire _65771_;
wire _65772_;
wire _65773_;
wire _65774_;
wire _65775_;
wire _65776_;
wire _65777_;
wire _65778_;
wire _65779_;
wire _65780_;
wire _65781_;
wire _65782_;
wire _65783_;
wire _65784_;
wire _65785_;
wire _65786_;
wire _65787_;
wire _65788_;
wire _65789_;
wire _65790_;
wire _65791_;
wire _65792_;
wire _65793_;
wire _65794_;
wire _65795_;
wire _65796_;
wire _65797_;
wire _65798_;
wire _65799_;
wire _65800_;
wire _65801_;
wire _65802_;
wire _65803_;
wire _65804_;
wire _65805_;
wire _65806_;
wire _65807_;
wire _65808_;
wire _65809_;
wire _65810_;
wire _65811_;
wire _65812_;
wire _65813_;
wire _65814_;
wire _65815_;
wire _65816_;
wire _65817_;
wire _65818_;
wire _65819_;
wire _65820_;
wire _65821_;
wire _65822_;
wire _65823_;
wire _65824_;
wire _65825_;
wire _65826_;
wire _65827_;
wire _65828_;
wire _65829_;
wire _65830_;
wire _65831_;
wire _65832_;
wire _65833_;
wire _65834_;
wire _65835_;
wire _65836_;
wire _65837_;
wire _65838_;
wire _65839_;
wire _65840_;
wire _65841_;
wire _65842_;
wire _65843_;
wire _65844_;
wire _65845_;
wire _65846_;
wire _65847_;
wire _65848_;
wire _65849_;
wire _65850_;
wire _65851_;
wire _65852_;
wire _65853_;
wire _65854_;
wire _65855_;
wire _65856_;
wire _65857_;
wire _65858_;
wire _65859_;
wire _65860_;
wire _65861_;
wire _65862_;
wire _65863_;
wire _65864_;
wire _65865_;
wire _65866_;
wire _65867_;
wire _65868_;
wire _65869_;
wire _65870_;
wire _65871_;
wire _65872_;
wire _65873_;
wire _65874_;
wire _65875_;
wire _65876_;
wire _65877_;
wire _65878_;
wire _65879_;
wire _65880_;
wire _65881_;
wire _65882_;
wire _65883_;
wire _65884_;
wire _65885_;
wire _65886_;
wire _65887_;
wire _65888_;
wire _65889_;
wire _65890_;
wire _65891_;
wire _65892_;
wire _65893_;
wire _65894_;
wire _65895_;
wire _65896_;
wire _65897_;
wire _65898_;
wire _65899_;
wire _65900_;
wire _65901_;
wire _65902_;
wire _65903_;
wire _65904_;
wire _65905_;
wire _65906_;
wire _65907_;
wire _65908_;
wire _65909_;
wire _65910_;
wire _65911_;
wire _65912_;
wire _65913_;
wire _65914_;
wire _65915_;
wire _65916_;
wire _65917_;
wire _65918_;
wire _65919_;
wire _65920_;
wire _65921_;
wire _65922_;
wire _65923_;
wire _65924_;
wire _65925_;
wire _65926_;
wire _65927_;
wire _65928_;
wire _65929_;
wire _65930_;
wire _65931_;
wire _65932_;
wire _65933_;
wire _65934_;
wire _65935_;
wire _65936_;
wire _65937_;
wire _65938_;
wire _65939_;
wire _65940_;
wire _65941_;
wire _65942_;
wire _65943_;
wire _65944_;
wire _65945_;
wire _65946_;
wire _65947_;
wire _65948_;
wire _65949_;
wire _65950_;
wire _65951_;
wire _65952_;
wire _65953_;
wire _65954_;
wire _65955_;
wire _65956_;
wire _65957_;
wire _65958_;
wire _65959_;
wire _65960_;
wire _65961_;
wire _65962_;
wire _65963_;
wire _65964_;
wire _65965_;
wire _65966_;
wire _65967_;
wire _65968_;
wire _65969_;
wire _65970_;
wire _65971_;
wire _65972_;
wire _65973_;
wire _65974_;
wire _65975_;
wire _65976_;
wire _65977_;
wire _65978_;
wire _65979_;
wire _65980_;
wire _65981_;
wire _65982_;
wire _65983_;
wire _65984_;
wire _65985_;
wire _65986_;
wire _65987_;
wire _65988_;
wire _65989_;
wire _65990_;
wire _65991_;
wire _65992_;
wire _65993_;
wire _65994_;
wire _65995_;
wire _65996_;
wire _65997_;
wire _65998_;
wire _65999_;
wire _66000_;
wire _66001_;
wire _66002_;
wire _66003_;
wire _66004_;
wire _66005_;
wire _66006_;
wire _66007_;
wire _66008_;
wire _66009_;
wire _66010_;
wire _66011_;
wire _66012_;
wire _66013_;
wire _66014_;
wire _66015_;
wire _66016_;
wire _66017_;
wire _66018_;
wire _66019_;
wire _66020_;
wire _66021_;
wire _66022_;
wire _66023_;
wire _66024_;
wire _66025_;
wire _66026_;
wire _66027_;
wire _66028_;
wire _66029_;
wire _66030_;
wire _66031_;
wire _66032_;
wire _66033_;
wire _66034_;
wire _66035_;
wire _66036_;
wire _66037_;
wire _66038_;
wire _66039_;
wire _66040_;
wire _66041_;
wire _66042_;
wire _66043_;
wire _66044_;
wire _66045_;
wire _66046_;
wire _66047_;
wire _66048_;
wire _66049_;
wire _66050_;
wire _66051_;
wire _66052_;
wire _66053_;
wire _66054_;
wire _66055_;
wire _66056_;
wire _66057_;
wire _66058_;
wire _66059_;
wire _66060_;
wire _66061_;
wire _66062_;
wire _66063_;
wire _66064_;
wire _66065_;
wire _66066_;
wire _66067_;
wire _66068_;
wire _66069_;
wire _66070_;
wire _66071_;
wire _66072_;
wire _66073_;
wire _66074_;
wire _66075_;
wire _66076_;
wire _66077_;
wire _66078_;
wire _66079_;
wire _66080_;
wire _66081_;
wire _66082_;
wire _66083_;
wire _66084_;
wire _66085_;
wire _66086_;
wire _66087_;
wire _66088_;
wire _66089_;
wire _66090_;
wire _66091_;
wire _66092_;
wire _66093_;
wire _66094_;
wire _66095_;
wire _66096_;
wire _66097_;
wire _66098_;
wire _66099_;
wire _66100_;
wire _66101_;
wire _66102_;
wire _66103_;
wire _66104_;
wire _66105_;
wire _66106_;
wire _66107_;
wire _66108_;
wire _66109_;
wire _66110_;
wire _66111_;
wire _66112_;
wire _66113_;
wire _66114_;
wire _66115_;
wire _66116_;
wire _66117_;
wire _66118_;
wire _66119_;
wire _66120_;
wire _66121_;
wire _66122_;
wire _66123_;
wire _66124_;
wire _66125_;
wire _66126_;
wire _66127_;
wire _66128_;
wire _66129_;
wire _66130_;
wire _66131_;
wire _66132_;
wire _66133_;
wire _66134_;
wire _66135_;
wire _66136_;
wire _66137_;
wire _66138_;
wire _66139_;
wire _66140_;
wire _66141_;
wire _66142_;
wire _66143_;
wire _66144_;
wire _66145_;
wire _66146_;
wire _66147_;
wire _66148_;
wire _66149_;
wire _66150_;
wire _66151_;
wire _66152_;
wire _66153_;
wire _66154_;
wire _66155_;
wire _66156_;
wire _66157_;
wire _66158_;
wire _66159_;
wire _66160_;
wire _66161_;
wire _66162_;
wire _66163_;
wire _66164_;
wire _66165_;
wire _66166_;
wire _66167_;
wire _66168_;
wire _66169_;
wire _66170_;
wire _66171_;
wire _66172_;
wire _66173_;
wire _66174_;
wire _66175_;
wire _66176_;
wire _66177_;
wire _66178_;
wire _66179_;
wire _66180_;
wire _66181_;
wire _66182_;
wire _66183_;
wire _66184_;
wire _66185_;
wire _66186_;
wire _66187_;
wire _66188_;
wire _66189_;
wire _66190_;
wire _66191_;
wire _66192_;
wire _66193_;
wire _66194_;
wire _66195_;
wire _66196_;
wire _66197_;
wire _66198_;
wire _66199_;
wire _66200_;
wire _66201_;
wire _66202_;
wire _66203_;
wire _66204_;
wire _66205_;
wire _66206_;
wire _66207_;
wire _66208_;
wire _66209_;
wire _66210_;
wire _66211_;
wire _66212_;
wire _66213_;
wire _66214_;
wire _66215_;
wire _66216_;
wire _66217_;
wire _66218_;
wire _66219_;
wire _66220_;
wire _66221_;
wire _66222_;
wire _66223_;
wire _66224_;
wire _66225_;
wire _66226_;
wire _66227_;
wire _66228_;
wire _66229_;
wire _66230_;
wire _66231_;
wire _66232_;
wire _66233_;
wire _66234_;
wire _66235_;
wire _66236_;
wire _66237_;
wire _66238_;
wire _66239_;
wire _66240_;
wire _66241_;
wire _66242_;
wire _66243_;
wire _66244_;
wire _66245_;
wire _66246_;
wire _66247_;
wire _66248_;
wire _66249_;
wire _66250_;
wire _66251_;
wire _66252_;
wire _66253_;
wire _66254_;
wire _66255_;
wire _66256_;
wire _66257_;
wire _66258_;
wire _66259_;
wire _66260_;
wire _66261_;
wire _66262_;
wire _66263_;
wire _66264_;
wire _66265_;
wire _66266_;
wire _66267_;
wire _66268_;
wire _66269_;
wire _66270_;
wire _66271_;
wire _66272_;
wire _66273_;
wire _66274_;
wire _66275_;
wire _66276_;
wire _66277_;
wire _66278_;
wire _66279_;
wire _66280_;
wire _66281_;
wire _66282_;
wire _66283_;
wire _66284_;
wire _66285_;
wire _66286_;
wire _66287_;
wire _66288_;
wire _66289_;
wire _66290_;
wire _66291_;
wire _66292_;
wire _66293_;
wire _66294_;
wire _66295_;
wire _66296_;
wire _66297_;
wire _66298_;
wire _66299_;
wire _66300_;
wire _66301_;
wire _66302_;
wire _66303_;
wire _66304_;
wire _66305_;
wire _66306_;
wire _66307_;
wire _66308_;
wire _66309_;
wire _66310_;
wire _66311_;
wire _66312_;
wire _66313_;
wire _66314_;
wire _66315_;
wire _66316_;
wire _66317_;
wire _66318_;
wire _66319_;
wire _66320_;
wire _66321_;
wire _66322_;
wire _66323_;
wire _66324_;
wire _66325_;
wire _66326_;
wire _66327_;
wire _66328_;
wire _66329_;
wire _66330_;
wire _66331_;
wire _66332_;
wire _66333_;
wire _66334_;
wire _66335_;
wire _66336_;
wire _66337_;
wire _66338_;
wire _66339_;
wire _66340_;
wire _66341_;
wire _66342_;
wire _66343_;
wire _66344_;
wire _66345_;
wire _66346_;
wire _66347_;
wire _66348_;
wire _66349_;
wire _66350_;
wire _66351_;
wire _66352_;
wire _66353_;
wire _66354_;
wire _66355_;
wire _66356_;
wire _66357_;
wire _66358_;
wire _66359_;
wire _66360_;
wire _66361_;
wire _66362_;
wire _66363_;
wire _66364_;
wire _66365_;
wire _66366_;
wire _66367_;
wire _66368_;
wire _66369_;
wire _66370_;
wire _66371_;
wire _66372_;
wire _66373_;
wire _66374_;
wire _66375_;
wire _66376_;
wire _66377_;
wire _66378_;
wire _66379_;
wire _66380_;
wire _66381_;
wire _66382_;
wire _66383_;
wire _66384_;
wire _66385_;
wire _66386_;
wire _66387_;
wire _66388_;
wire _66389_;
wire _66390_;
wire _66391_;
wire _66392_;
wire _66393_;
wire _66394_;
wire _66395_;
wire _66396_;
wire _66397_;
wire _66398_;
wire _66399_;
wire _66400_;
wire _66401_;
wire _66402_;
wire _66403_;
wire _66404_;
wire _66405_;
wire _66406_;
wire _66407_;
wire _66408_;
wire _66409_;
wire _66410_;
wire _66411_;
wire _66412_;
wire _66413_;
wire _66414_;
wire _66415_;
wire _66416_;
wire _66417_;
wire _66418_;
wire _66419_;
wire _66420_;
wire _66421_;
wire _66422_;
wire _66423_;
wire _66424_;
wire _66425_;
wire _66426_;
wire _66427_;
wire _66428_;
wire _66429_;
wire _66430_;
wire _66431_;
wire _66432_;
wire _66433_;
wire _66434_;
wire _66435_;
wire _66436_;
wire _66437_;
wire _66438_;
wire _66439_;
wire _66440_;
wire _66441_;
wire _66442_;
wire _66443_;
wire _66444_;
wire _66445_;
wire _66446_;
wire _66447_;
wire _66448_;
wire _66449_;
wire _66450_;
wire _66451_;
wire _66452_;
wire _66453_;
wire _66454_;
wire _66455_;
wire _66456_;
wire _66457_;
wire _66458_;
wire _66459_;
wire _66460_;
wire _66461_;
wire _66462_;
wire _66463_;
wire _66464_;
wire _66465_;
wire _66466_;
wire _66467_;
wire _66468_;
wire _66469_;
wire _66470_;
wire _66471_;
wire _66472_;
wire _66473_;
wire _66474_;
wire _66475_;
wire _66476_;
wire _66477_;
wire _66478_;
wire _66479_;
wire _66480_;
wire _66481_;
wire _66482_;
wire _66483_;
wire _66484_;
wire _66485_;
wire _66486_;
wire _66487_;
wire _66488_;
wire _66489_;
wire _66490_;
wire _66491_;
wire _66492_;
wire _66493_;
wire _66494_;
wire _66495_;
wire _66496_;
wire _66497_;
wire _66498_;
wire _66499_;
wire _66500_;
wire _66501_;
wire _66502_;
wire _66503_;
wire _66504_;
wire _66505_;
wire _66506_;
wire _66507_;
wire _66508_;
wire _66509_;
wire _66510_;
wire _66511_;
wire _66512_;
wire _66513_;
wire _66514_;
wire _66515_;
wire _66516_;
wire _66517_;
wire _66518_;
wire _66519_;
wire _66520_;
wire _66521_;
wire _66522_;
wire _66523_;
wire _66524_;
wire _66525_;
wire _66526_;
wire _66527_;
wire _66528_;
wire _66529_;
wire _66530_;
wire _66531_;
wire _66532_;
wire _66533_;
wire _66534_;
wire _66535_;
wire _66536_;
wire _66537_;
wire _66538_;
wire _66539_;
wire _66540_;
wire _66541_;
wire _66542_;
wire _66543_;
wire _66544_;
wire _66545_;
wire _66546_;
wire _66547_;
wire _66548_;
wire _66549_;
wire _66550_;
wire _66551_;
wire _66552_;
wire _66553_;
wire _66554_;
wire _66555_;
wire _66556_;
wire _66557_;
wire _66558_;
wire _66559_;
wire _66560_;
wire _66561_;
wire _66562_;
wire _66563_;
wire _66564_;
wire _66565_;
wire _66566_;
wire _66567_;
wire _66568_;
wire _66569_;
wire _66570_;
wire _66571_;
wire _66572_;
wire _66573_;
wire _66574_;
wire _66575_;
wire _66576_;
wire _66577_;
wire _66578_;
wire _66579_;
wire _66580_;
wire _66581_;
wire _66582_;
wire _66583_;
wire _66584_;
wire _66585_;
wire _66586_;
wire _66587_;
wire _66588_;
wire _66589_;
wire _66590_;
wire _66591_;
wire _66592_;
wire _66593_;
wire _66594_;
wire _66595_;
wire _66596_;
wire _66597_;
wire _66598_;
wire _66599_;
wire _66600_;
wire _66601_;
wire _66602_;
wire _66603_;
wire _66604_;
wire _66605_;
wire _66606_;
wire _66607_;
wire _66608_;
wire _66609_;
wire _66610_;
wire _66611_;
wire _66612_;
wire _66613_;
wire _66614_;
wire _66615_;
wire _66616_;
wire _66617_;
wire _66618_;
wire _66619_;
wire _66620_;
wire _66621_;
wire _66622_;
wire _66623_;
wire _66624_;
wire _66625_;
wire _66626_;
wire _66627_;
wire _66628_;
wire _66629_;
wire _66630_;
wire _66631_;
wire _66632_;
wire _66633_;
wire _66634_;
wire _66635_;
wire _66636_;
wire _66637_;
wire _66638_;
wire _66639_;
wire _66640_;
wire _66641_;
wire _66642_;
wire _66643_;
wire _66644_;
wire _66645_;
wire _66646_;
wire _66647_;
wire _66648_;
wire _66649_;
wire _66650_;
wire _66651_;
wire _66652_;
wire _66653_;
wire _66654_;
wire _66655_;
wire _66656_;
wire _66657_;
wire _66658_;
wire _66659_;
wire _66660_;
wire _66661_;
wire _66662_;
wire _66663_;
wire _66664_;
wire _66665_;
wire _66666_;
wire _66667_;
wire _66668_;
wire _66669_;
wire _66670_;
wire _66671_;
wire _66672_;
wire _66673_;
wire _66674_;
wire _66675_;
wire _66676_;
wire _66677_;
wire _66678_;
wire _66679_;
wire _66680_;
wire _66681_;
wire _66682_;
wire _66683_;
wire _66684_;
wire _66685_;
wire _66686_;
wire _66687_;
wire _66688_;
wire _66689_;
wire _66690_;
wire _66691_;
wire _66692_;
wire _66693_;
wire _66694_;
wire _66695_;
wire _66696_;
wire _66697_;
wire _66698_;
wire _66699_;
wire _66700_;
wire _66701_;
wire _66702_;
wire _66703_;
wire _66704_;
wire _66705_;
wire _66706_;
wire _66707_;
wire _66708_;
wire _66709_;
wire _66710_;
wire _66711_;
wire _66712_;
wire _66713_;
wire _66714_;
wire _66715_;
wire _66716_;
wire _66717_;
wire _66718_;
wire _66719_;
wire _66720_;
wire _66721_;
wire _66722_;
wire _66723_;
wire _66724_;
wire _66725_;
wire _66726_;
wire _66727_;
wire _66728_;
wire _66729_;
wire _66730_;
wire _66731_;
wire _66732_;
wire _66733_;
wire _66734_;
wire _66735_;
wire _66736_;
wire _66737_;
wire _66738_;
wire _66739_;
wire _66740_;
wire _66741_;
wire _66742_;
wire _66743_;
wire _66744_;
wire _66745_;
wire _66746_;
wire _66747_;
wire _66748_;
wire _66749_;
wire _66750_;
wire _66751_;
wire _66752_;
wire _66753_;
wire _66754_;
wire _66755_;
wire _66756_;
wire _66757_;
wire _66758_;
wire _66759_;
wire _66760_;
wire _66761_;
wire _66762_;
wire _66763_;
wire _66764_;
wire _66765_;
wire _66766_;
wire _66767_;
wire _66768_;
wire _66769_;
wire _66770_;
wire _66771_;
wire _66772_;
wire _66773_;
wire _66774_;
wire _66775_;
wire _66776_;
wire _66777_;
wire _66778_;
wire _66779_;
wire _66780_;
wire _66781_;
wire _66782_;
wire _66783_;
wire _66784_;
wire _66785_;
wire _66786_;
wire _66787_;
wire _66788_;
wire _66789_;
wire _66790_;
wire _66791_;
wire _66792_;
wire _66793_;
wire _66794_;
wire _66795_;
wire _66796_;
wire _66797_;
wire _66798_;
wire _66799_;
wire _66800_;
wire _66801_;
wire _66802_;
wire _66803_;
wire _66804_;
wire _66805_;
wire _66806_;
wire _66807_;
wire _66808_;
wire _66809_;
wire _66810_;
wire _66811_;
wire _66812_;
wire _66813_;
wire _66814_;
wire _66815_;
wire _66816_;
wire _66817_;
wire _66818_;
wire _66819_;
wire _66820_;
wire _66821_;
wire _66822_;
wire _66823_;
wire _66824_;
wire _66825_;
wire _66826_;
wire _66827_;
wire _66828_;
wire _66829_;
wire _66830_;
wire _66831_;
wire _66832_;
wire _66833_;
wire _66834_;
wire _66835_;
wire _66836_;
wire _66837_;
wire _66838_;
wire _66839_;
wire _66840_;
wire _66841_;
wire _66842_;
wire _66843_;
wire _66844_;
wire _66845_;
wire _66846_;
wire _66847_;
wire _66848_;
wire _66849_;
wire _66850_;
wire _66851_;
wire _66852_;
wire _66853_;
wire _66854_;
wire _66855_;
wire _66856_;
wire _66857_;
wire _66858_;
wire _66859_;
wire _66860_;
wire _66861_;
wire _66862_;
wire _66863_;
wire _66864_;
wire _66865_;
wire _66866_;
wire _66867_;
wire _66868_;
wire _66869_;
wire _66870_;
wire _66871_;
wire _66872_;
wire _66873_;
wire _66874_;
wire _66875_;
wire _66876_;
wire _66877_;
wire _66878_;
wire _66879_;
wire _66880_;
wire _66881_;
wire _66882_;
wire _66883_;
wire _66884_;
wire _66885_;
wire _66886_;
wire _66887_;
wire _66888_;
wire _66889_;
wire _66890_;
wire _66891_;
wire _66892_;
wire _66893_;
wire _66894_;
wire _66895_;
wire _66896_;
wire _66897_;
wire _66898_;
wire _66899_;
wire _66900_;
wire _66901_;
wire _66902_;
wire _66903_;
wire _66904_;
wire _66905_;
wire _66906_;
wire _66907_;
wire _66908_;
wire _66909_;
wire _66910_;
wire _66911_;
wire _66912_;
wire _66913_;
wire _66914_;
wire _66915_;
wire _66916_;
wire _66917_;
wire _66918_;
wire _66919_;
wire _66920_;
wire _66921_;
wire _66922_;
wire _66923_;
wire _66924_;
wire _66925_;
wire _66926_;
wire _66927_;
wire _66928_;
wire _66929_;
wire _66930_;
wire _66931_;
wire _66932_;
wire _66933_;
wire _66934_;
wire _66935_;
wire _66936_;
wire _66937_;
wire _66938_;
wire _66939_;
wire _66940_;
wire _66941_;
wire _66942_;
wire _66943_;
wire _66944_;
wire _66945_;
wire _66946_;
wire _66947_;
wire _66948_;
wire _66949_;
wire _66950_;
wire _66951_;
wire _66952_;
wire _66953_;
wire _66954_;
wire _66955_;
wire _66956_;
wire _66957_;
wire _66958_;
wire _66959_;
wire _66960_;
wire _66961_;
wire _66962_;
wire _66963_;
wire _66964_;
wire _66965_;
wire _66966_;
wire _66967_;
wire _66968_;
wire _66969_;
wire _66970_;
wire _66971_;
wire _66972_;
wire _66973_;
wire _66974_;
wire _66975_;
wire _66976_;
wire _66977_;
wire _66978_;
wire _66979_;
wire _66980_;
wire _66981_;
wire _66982_;
wire _66983_;
wire _66984_;
wire _66985_;
wire _66986_;
wire _66987_;
wire _66988_;
wire _66989_;
wire _66990_;
wire _66991_;
wire _66992_;
wire _66993_;
wire _66994_;
wire _66995_;
wire _66996_;
wire _66997_;
wire _66998_;
wire _66999_;
wire _67000_;
wire _67001_;
wire _67002_;
wire _67003_;
wire _67004_;
wire _67005_;
wire _67006_;
wire _67007_;
wire _67008_;
wire _67009_;
wire _67010_;
wire _67011_;
wire _67012_;
wire _67013_;
wire _67014_;
wire _67015_;
wire _67016_;
wire _67017_;
wire _67018_;
wire _67019_;
wire _67020_;
wire _67021_;
wire _67022_;
wire _67023_;
wire _67024_;
wire _67025_;
wire _67026_;
wire _67027_;
wire _67028_;
wire _67029_;
wire _67030_;
wire _67031_;
wire _67032_;
wire _67033_;
wire _67034_;
wire _67035_;
wire _67036_;
wire _67037_;
wire _67038_;
wire _67039_;
wire _67040_;
wire _67041_;
wire _67042_;
wire _67043_;
wire _67044_;
wire _67045_;
wire _67046_;
wire _67047_;
wire _67048_;
wire _67049_;
wire _67050_;
wire _67051_;
wire _67052_;
wire _67053_;
wire _67054_;
wire _67055_;
wire _67056_;
wire _67057_;
wire _67058_;
wire _67059_;
wire _67060_;
wire _67061_;
wire _67062_;
wire _67063_;
wire _67064_;
wire _67065_;
wire _67066_;
wire _67067_;
wire _67068_;
wire _67069_;
wire _67070_;
wire _67071_;
wire _67072_;
wire _67073_;
wire _67074_;
wire _67075_;
wire _67076_;
wire _67077_;
wire _67078_;
wire _67079_;
wire _67080_;
wire _67081_;
wire _67082_;
wire _67083_;
wire _67084_;
wire _67085_;
wire _67086_;
wire _67087_;
wire _67088_;
wire _67089_;
wire _67090_;
wire _67091_;
wire _67092_;
wire _67093_;
wire _67094_;
wire _67095_;
wire _67096_;
wire _67097_;
wire _67098_;
wire _67099_;
wire _67100_;
wire _67101_;
wire _67102_;
wire _67103_;
wire _67104_;
wire _67105_;
wire _67106_;
wire _67107_;
wire _67108_;
wire _67109_;
wire _67110_;
wire _67111_;
wire _67112_;
wire _67113_;
wire _67114_;
wire _67115_;
wire _67116_;
wire _67117_;
wire _67118_;
wire _67119_;
wire _67120_;
wire _67121_;
wire _67122_;
wire _67123_;
wire _67124_;
wire _67125_;
wire _67126_;
wire _67127_;
wire _67128_;
wire _67129_;
wire _67130_;
wire _67131_;
wire _67132_;
wire _67133_;
wire _67134_;
wire _67135_;
wire _67136_;
wire _67137_;
wire _67138_;
wire _67139_;
wire _67140_;
wire _67141_;
wire _67142_;
wire _67143_;
wire _67144_;
wire _67145_;
wire _67146_;
wire _67147_;
wire _67148_;
wire _67149_;
wire _67150_;
wire _67151_;
wire _67152_;
wire _67153_;
wire _67154_;
wire _67155_;
wire _67156_;
wire _67157_;
wire _67158_;
wire _67159_;
wire _67160_;
wire _67161_;
wire _67162_;
wire _67163_;
wire _67164_;
wire _67165_;
wire _67166_;
wire _67167_;
wire _67168_;
wire _67169_;
wire _67170_;
wire _67171_;
wire _67172_;
wire _67173_;
wire _67174_;
wire _67175_;
wire _67176_;
wire _67177_;
wire _67178_;
wire _67179_;
wire _67180_;
wire _67181_;
wire _67182_;
wire _67183_;
wire _67184_;
wire _67185_;
wire _67186_;
wire _67187_;
wire _67188_;
wire _67189_;
wire _67190_;
wire _67191_;
wire _67192_;
wire _67193_;
wire _67194_;
wire _67195_;
wire _67196_;
wire _67197_;
wire _67198_;
wire _67199_;
wire _67200_;
wire _67201_;
wire _67202_;
wire _67203_;
wire _67204_;
wire _67205_;
wire _67206_;
wire _67207_;
wire _67208_;
wire _67209_;
wire _67210_;
wire _67211_;
wire _67212_;
wire _67213_;
wire _67214_;
wire _67215_;
wire _67216_;
wire _67217_;
wire _67218_;
wire _67219_;
wire _67220_;
wire _67221_;
wire _67222_;
wire _67223_;
wire _67224_;
wire _67225_;
wire _67226_;
wire _67227_;
wire _67228_;
wire _67229_;
wire _67230_;
wire _67231_;
wire _67232_;
wire _67233_;
wire _67234_;
wire _67235_;
wire _67236_;
wire _67237_;
wire _67238_;
wire _67239_;
wire _67240_;
wire _67241_;
wire _67242_;
wire _67243_;
wire _67244_;
wire _67245_;
wire _67246_;
wire _67247_;
wire _67248_;
wire _67249_;
wire _67250_;
wire _67251_;
wire _67252_;
wire _67253_;
wire _67254_;
wire _67255_;
wire _67256_;
wire _67257_;
wire _67258_;
wire _67259_;
wire _67260_;
wire _67261_;
wire _67262_;
wire _67263_;
wire _67264_;
wire _67265_;
wire _67266_;
wire _67267_;
wire _67268_;
wire _67269_;
wire _67270_;
wire _67271_;
wire _67272_;
wire _67273_;
wire _67274_;
wire _67275_;
wire _67276_;
wire _67277_;
wire _67278_;
wire _67279_;
wire _67280_;
wire _67281_;
wire _67282_;
wire _67283_;
wire _67284_;
wire _67285_;
wire _67286_;
wire _67287_;
wire _67288_;
wire _67289_;
wire _67290_;
wire _67291_;
wire _67292_;
wire _67293_;
wire _67294_;
wire _67295_;
wire _67296_;
wire _67297_;
wire _67298_;
wire _67299_;
wire _67300_;
wire _67301_;
wire _67302_;
wire _67303_;
wire _67304_;
wire _67305_;
wire _67306_;
wire _67307_;
wire _67308_;
wire _67309_;
wire _67310_;
wire _67311_;
wire _67312_;
wire _67313_;
wire _67314_;
wire _67315_;
wire _67316_;
wire _67317_;
wire _67318_;
wire _67319_;
wire _67320_;
wire _67321_;
wire _67322_;
wire _67323_;
wire _67324_;
wire _67325_;
wire _67326_;
wire _67327_;
wire _67328_;
wire _67329_;
wire _67330_;
wire _67331_;
wire _67332_;
wire _67333_;
wire _67334_;
wire _67335_;
wire _67336_;
wire _67337_;
wire _67338_;
wire _67339_;
wire _67340_;
wire _67341_;
wire _67342_;
wire _67343_;
wire _67344_;
wire _67345_;
wire _67346_;
wire _67347_;
wire _67348_;
wire _67349_;
wire _67350_;
wire _67351_;
wire _67352_;
wire _67353_;
wire _67354_;
wire _67355_;
wire _67356_;
wire _67357_;
wire _67358_;
wire _67359_;
wire _67360_;
wire _67361_;
wire _67362_;
wire _67363_;
wire _67364_;
wire _67365_;
wire _67366_;
wire _67367_;
wire _67368_;
wire _67369_;
wire _67370_;
wire _67371_;
wire _67372_;
wire _67373_;
wire _67374_;
wire _67375_;
wire _67376_;
wire _67377_;
wire _67378_;
wire _67379_;
wire _67380_;
wire _67381_;
wire _67382_;
wire _67383_;
wire _67384_;
wire _67385_;
wire _67386_;
wire _67387_;
wire _67388_;
wire _67389_;
wire _67390_;
wire _67391_;
wire _67392_;
wire _67393_;
wire _67394_;
wire _67395_;
wire _67396_;
wire _67397_;
wire _67398_;
wire _67399_;
wire _67400_;
wire _67401_;
wire _67402_;
wire _67403_;
wire _67404_;
wire _67405_;
wire _67406_;
wire _67407_;
wire _67408_;
wire _67409_;
wire _67410_;
wire _67411_;
wire _67412_;
wire _67413_;
wire _67414_;
wire _67415_;
wire _67416_;
wire _67417_;
wire _67418_;
wire _67419_;
wire _67420_;
wire _67421_;
wire _67422_;
wire _67423_;
wire _67424_;
wire _67425_;
wire _67426_;
wire _67427_;
wire _67428_;
wire _67429_;
wire _67430_;
wire _67431_;
wire _67432_;
wire _67433_;
wire _67434_;
wire _67435_;
wire _67436_;
wire _67437_;
wire _67438_;
wire _67439_;
wire _67440_;
wire _67441_;
wire _67442_;
wire _67443_;
wire _67444_;
wire _67445_;
wire _67446_;
wire _67447_;
wire _67448_;
wire _67449_;
wire _67450_;
wire _67451_;
wire _67452_;
wire _67453_;
wire _67454_;
wire _67455_;
wire _67456_;
wire _67457_;
wire _67458_;
wire _67459_;
wire _67460_;
wire _67461_;
wire _67462_;
wire _67463_;
wire _67464_;
wire _67465_;
wire _67466_;
wire _67467_;
wire _67468_;
wire _67469_;
wire _67470_;
wire _67471_;
wire _67472_;
wire _67473_;
wire _67474_;
wire _67475_;
wire _67476_;
wire _67477_;
wire _67478_;
wire _67479_;
wire _67480_;
wire _67481_;
wire _67482_;
wire _67483_;
wire _67484_;
wire _67485_;
wire _67486_;
wire _67487_;
wire _67488_;
wire _67489_;
wire _67490_;
wire _67491_;
wire _67492_;
wire _67493_;
wire _67494_;
wire _67495_;
wire _67496_;
wire _67497_;
wire _67498_;
wire _67499_;
wire _67500_;
wire _67501_;
wire _67502_;
wire _67503_;
wire _67504_;
wire _67505_;
wire _67506_;
wire _67507_;
wire _67508_;
wire _67509_;
wire _67510_;
wire _67511_;
wire _67512_;
wire _67513_;
wire _67514_;
wire _67515_;
wire _67516_;
wire _67517_;
wire _67518_;
wire _67519_;
wire _67520_;
wire _67521_;
wire _67522_;
wire _67523_;
wire _67524_;
wire _67525_;
wire _67526_;
wire _67527_;
wire _67528_;
wire _67529_;
wire _67530_;
wire _67531_;
wire _67532_;
wire _67533_;
wire _67534_;
wire _67535_;
wire _67536_;
wire _67537_;
wire _67538_;
wire _67539_;
wire _67540_;
wire _67541_;
wire _67542_;
wire _67543_;
wire _67544_;
wire _67545_;
wire _67546_;
wire _67547_;
wire _67548_;
wire _67549_;
wire _67550_;
wire _67551_;
wire _67552_;
wire _67553_;
wire _67554_;
wire _67555_;
wire _67556_;
wire _67557_;
wire _67558_;
wire _67559_;
wire _67560_;
wire _67561_;
wire _67562_;
wire _67563_;
wire _67564_;
wire _67565_;
wire _67566_;
wire _67567_;
wire _67568_;
wire _67569_;
wire _67570_;
wire _67571_;
wire _67572_;
wire _67573_;
wire _67574_;
wire _67575_;
wire _67576_;
wire _67577_;
wire _67578_;
wire _67579_;
wire _67580_;
wire _67581_;
wire _67582_;
wire _67583_;
wire _67584_;
wire _67585_;
wire _67586_;
wire _67587_;
wire _67588_;
wire _67589_;
wire _67590_;
wire _67591_;
wire _67592_;
wire _67593_;
wire _67594_;
wire _67595_;
wire _67596_;
wire _67597_;
wire _67598_;
wire _67599_;
wire _67600_;
wire _67601_;
wire _67602_;
wire _67603_;
wire _67604_;
wire _67605_;
wire _67606_;
wire _67607_;
wire _67608_;
wire _67609_;
wire _67610_;
wire _67611_;
wire _67612_;
wire _67613_;
wire _67614_;
wire _67615_;
wire _67616_;
wire _67617_;
wire _67618_;
wire _67619_;
wire _67620_;
wire _67621_;
wire _67622_;
wire _67623_;
wire _67624_;
wire _67625_;
wire _67626_;
wire _67627_;
wire _67628_;
wire _67629_;
wire _67630_;
wire _67631_;
wire _67632_;
wire _67633_;
wire _67634_;
wire _67635_;
wire _67636_;
wire _67637_;
wire _67638_;
wire _67639_;
wire _67640_;
wire _67641_;
wire _67642_;
wire _67643_;
wire _67644_;
wire _67645_;
wire _67646_;
wire _67647_;
wire _67648_;
wire _67649_;
wire _67650_;
wire _67651_;
wire _67652_;
wire _67653_;
wire _67654_;
wire _67655_;
wire _67656_;
wire _67657_;
wire _67658_;
wire _67659_;
wire _67660_;
wire _67661_;
wire _67662_;
wire _67663_;
wire _67664_;
wire _67665_;
wire _67666_;
wire _67667_;
wire _67668_;
wire _67669_;
wire _67670_;
wire _67671_;
wire _67672_;
wire _67673_;
wire _67674_;
wire _67675_;
wire _67676_;
wire _67677_;
wire _67678_;
wire _67679_;
wire _67680_;
wire _67681_;
wire _67682_;
wire _67683_;
wire _67684_;
wire _67685_;
wire _67686_;
wire _67687_;
wire _67688_;
wire _67689_;
wire _67690_;
wire _67691_;
wire _67692_;
wire _67693_;
wire _67694_;
wire _67695_;
wire _67696_;
wire _67697_;
wire _67698_;
wire _67699_;
wire _67700_;
wire _67701_;
wire _67702_;
wire _67703_;
wire _67704_;
wire _67705_;
wire _67706_;
wire _67707_;
wire _67708_;
wire _67709_;
wire _67710_;
wire _67711_;
wire _67712_;
wire _67713_;
wire _67714_;
wire _67715_;
wire _67716_;
wire _67717_;
wire _67718_;
wire _67719_;
wire _67720_;
wire _67721_;
wire _67722_;
wire _67723_;
wire _67724_;
wire _67725_;
wire _67726_;
wire _67727_;
wire _67728_;
wire _67729_;
wire _67730_;
wire _67731_;
wire _67732_;
wire _67733_;
wire _67734_;
wire _67735_;
wire _67736_;
wire _67737_;
wire _67738_;
wire _67739_;
wire _67740_;
wire _67741_;
wire _67742_;
wire _67743_;
wire _67744_;
wire _67745_;
wire _67746_;
wire _67747_;
wire _67748_;
wire _67749_;
wire _67750_;
wire _67751_;
wire _67752_;
wire _67753_;
wire _67754_;
wire _67755_;
wire _67756_;
wire _67757_;
wire _67758_;
wire _67759_;
wire _67760_;
wire _67761_;
wire _67762_;
wire _67763_;
wire _67764_;
wire _67765_;
wire _67766_;
wire _67767_;
wire _67768_;
wire _67769_;
wire _67770_;
wire _67771_;
wire _67772_;
wire _67773_;
wire _67774_;
wire _67775_;
wire _67776_;
wire _67777_;
wire _67778_;
wire _67779_;
wire _67780_;
wire _67781_;
wire _67782_;
wire _67783_;
wire _67784_;
wire _67785_;
wire _67786_;
wire _67787_;
wire _67788_;
wire _67789_;
wire _67790_;
wire _67791_;
wire _67792_;
wire _67793_;
wire _67794_;
wire _67795_;
wire _67796_;
wire _67797_;
wire _67798_;
wire _67799_;
wire _67800_;
wire _67801_;
wire _67802_;
wire _67803_;
wire _67804_;
wire _67805_;
wire _67806_;
wire _67807_;
wire _67808_;
wire _67809_;
wire _67810_;
wire _67811_;
wire _67812_;
wire _67813_;
wire _67814_;
wire _67815_;
wire _67816_;
wire _67817_;
wire _67818_;
wire _67819_;
wire _67820_;
wire _67821_;
wire _67822_;
wire _67823_;
wire _67824_;
wire _67825_;
wire _67826_;
wire _67827_;
wire _67828_;
wire _67829_;
wire _67830_;
wire _67831_;
wire _67832_;
wire _67833_;
wire _67834_;
wire _67835_;
wire _67836_;
wire _67837_;
wire _67838_;
wire _67839_;
wire _67840_;
wire _67841_;
wire _67842_;
wire _67843_;
wire _67844_;
wire _67845_;
wire _67846_;
wire _67847_;
wire _67848_;
wire _67849_;
wire _67850_;
wire _67851_;
wire _67852_;
wire _67853_;
wire _67854_;
wire _67855_;
wire _67856_;
wire _67857_;
wire _67858_;
wire _67859_;
wire _67860_;
wire _67861_;
wire _67862_;
wire _67863_;
wire _67864_;
wire _67865_;
wire _67866_;
wire _67867_;
wire _67868_;
wire _67869_;
wire _67870_;
wire _67871_;
wire _67872_;
wire _67873_;
wire _67874_;
wire _67875_;
wire _67876_;
wire _67877_;
wire _67878_;
wire _67879_;
wire _67880_;
wire _67881_;
wire _67882_;
wire _67883_;
wire _67884_;
wire _67885_;
wire _67886_;
wire _67887_;
wire _67888_;
wire _67889_;
wire _67890_;
wire _67891_;
wire _67892_;
wire _67893_;
wire _67894_;
wire _67895_;
wire _67896_;
wire _67897_;
wire _67898_;
wire _67899_;
wire _67900_;
wire _67901_;
wire _67902_;
wire _67903_;
wire _67904_;
wire _67905_;
wire _67906_;
wire _67907_;
wire _67908_;
wire _67909_;
wire _67910_;
wire _67911_;
wire _67912_;
wire _67913_;
wire _67914_;
wire _67915_;
wire _67916_;
wire _67917_;
wire _67918_;
wire _67919_;
wire _67920_;
wire _67921_;
wire _67922_;
wire _67923_;
wire _67924_;
wire _67925_;
wire _67926_;
wire _67927_;
wire _67928_;
wire _67929_;
wire _67930_;
wire _67931_;
wire _67932_;
wire _67933_;
wire _67934_;
wire _67935_;
wire _67936_;
wire _67937_;
wire _67938_;
wire _67939_;
wire _67940_;
wire _67941_;
wire _67942_;
wire _67943_;
wire _67944_;
wire _67945_;
wire _67946_;
wire _67947_;
wire _67948_;
wire _67949_;
wire _67950_;
wire _67951_;
wire _67952_;
wire _67953_;
wire _67954_;
wire _67955_;
wire _67956_;
wire _67957_;
wire _67958_;
wire _67959_;
wire _67960_;
wire _67961_;
wire _67962_;
wire _67963_;
wire _67964_;
wire _67965_;
wire _67966_;
wire _67967_;
wire _67968_;
wire _67969_;
wire _67970_;
wire _67971_;
wire _67972_;
wire _67973_;
wire _67974_;
wire _67975_;
wire _67976_;
wire _67977_;
wire _67978_;
wire _67979_;
wire _67980_;
wire _67981_;
wire _67982_;
wire _67983_;
wire _67984_;
wire _67985_;
wire _67986_;
wire _67987_;
wire _67988_;
wire _67989_;
wire _67990_;
wire _67991_;
wire _67992_;
wire _67993_;
wire _67994_;
wire _67995_;
wire _67996_;
wire _67997_;
wire _67998_;
wire _67999_;
wire _68000_;
wire _68001_;
wire _68002_;
wire _68003_;
wire _68004_;
wire _68005_;
wire _68006_;
wire _68007_;
wire _68008_;
wire _68009_;
wire _68010_;
wire _68011_;
wire _68012_;
wire _68013_;
wire _68014_;
wire _68015_;
wire _68016_;
wire _68017_;
wire _68018_;
wire _68019_;
wire _68020_;
wire _68021_;
wire _68022_;
wire _68023_;
wire _68024_;
wire _68025_;
wire _68026_;
wire _68027_;
wire _68028_;
wire _68029_;
wire _68030_;
wire _68031_;
wire _68032_;
wire _68033_;
wire _68034_;
wire _68035_;
wire _68036_;
wire _68037_;
wire _68038_;
wire _68039_;
wire _68040_;
wire _68041_;
wire _68042_;
wire _68043_;
wire _68044_;
wire _68045_;
wire _68046_;
wire _68047_;
wire _68048_;
wire _68049_;
wire _68050_;
wire _68051_;
wire _68052_;
wire _68053_;
wire _68054_;
wire _68055_;
wire _68056_;
wire _68057_;
wire _68058_;
wire _68059_;
wire _68060_;
wire _68061_;
wire _68062_;
wire _68063_;
wire _68064_;
wire _68065_;
wire _68066_;
wire _68067_;
wire _68068_;
wire _68069_;
wire _68070_;
wire _68071_;
wire _68072_;
wire _68073_;
wire _68074_;
wire _68075_;
wire _68076_;
wire _68077_;
wire _68078_;
wire _68079_;
wire _68080_;
wire _68081_;
wire _68082_;
wire _68083_;
wire _68084_;
wire _68085_;
wire _68086_;
wire _68087_;
wire _68088_;
wire _68089_;
wire _68090_;
wire _68091_;
wire _68092_;
wire _68093_;
wire _68094_;
wire _68095_;
wire _68096_;
wire _68097_;
wire _68098_;
wire _68099_;
wire _68100_;
wire _68101_;
wire _68102_;
wire _68103_;
wire _68104_;
wire _68105_;
wire _68106_;
wire _68107_;
wire _68108_;
wire _68109_;
wire _68110_;
wire _68111_;
wire _68112_;
wire _68113_;
wire _68114_;
wire _68115_;
wire _68116_;
wire _68117_;
wire _68118_;
wire _68119_;
wire _68120_;
wire _68121_;
wire _68122_;
wire _68123_;
wire _68124_;
wire _68125_;
wire _68126_;
wire _68127_;
wire _68128_;
wire _68129_;
wire _68130_;
wire _68131_;
wire _68132_;
wire _68133_;
wire _68134_;
wire _68135_;
wire _68136_;
wire _68137_;
wire _68138_;
wire _68139_;
wire _68140_;
wire _68141_;
wire _68142_;
wire _68143_;
wire _68144_;
wire _68145_;
wire _68146_;
wire _68147_;
wire _68148_;
wire _68149_;
wire _68150_;
wire _68151_;
wire _68152_;
wire _68153_;
wire _68154_;
wire _68155_;
wire _68156_;
wire _68157_;
wire _68158_;
wire _68159_;
wire _68160_;
wire _68161_;
wire _68162_;
wire _68163_;
wire _68164_;
wire _68165_;
wire _68166_;
wire _68167_;
wire _68168_;
wire _68169_;
wire _68170_;
wire _68171_;
wire _68172_;
wire _68173_;
wire _68174_;
wire _68175_;
wire _68176_;
wire _68177_;
wire _68178_;
wire _68179_;
wire _68180_;
wire _68181_;
wire _68182_;
wire _68183_;
wire _68184_;
wire _68185_;
wire _68186_;
wire _68187_;
wire _68188_;
wire _68189_;
wire _68190_;
wire _68191_;
wire _68192_;
wire _68193_;
wire _68194_;
wire _68195_;
wire _68196_;
wire _68197_;
wire _68198_;
wire _68199_;
wire _68200_;
wire _68201_;
wire _68202_;
wire _68203_;
wire _68204_;
wire _68205_;
wire _68206_;
wire _68207_;
wire _68208_;
wire _68209_;
wire _68210_;
wire _68211_;
wire _68212_;
wire _68213_;
wire _68214_;
wire _68215_;
wire _68216_;
wire _68217_;
wire _68218_;
wire _68219_;
wire _68220_;
wire _68221_;
wire _68222_;
wire _68223_;
wire _68224_;
wire _68225_;
wire _68226_;
wire _68227_;
wire _68228_;
wire _68229_;
wire _68230_;
wire _68231_;
wire _68232_;
wire _68233_;
wire _68234_;
wire _68235_;
wire _68236_;
wire _68237_;
wire _68238_;
wire _68239_;
wire _68240_;
wire _68241_;
wire _68242_;
wire _68243_;
wire _68244_;
wire _68245_;
wire _68246_;
wire _68247_;
wire _68248_;
wire _68249_;
wire _68250_;
wire _68251_;
wire _68252_;
wire _68253_;
wire _68254_;
wire _68255_;
wire _68256_;
wire _68257_;
wire _68258_;
wire _68259_;
wire _68260_;
wire _68261_;
wire _68262_;
wire _68263_;
wire _68264_;
wire _68265_;
wire _68266_;
wire _68267_;
wire _68268_;
wire _68269_;
wire _68270_;
wire _68271_;
wire _68272_;
wire _68273_;
wire _68274_;
wire _68275_;
wire _68276_;
wire _68277_;
wire _68278_;
wire _68279_;
wire _68280_;
wire _68281_;
wire _68282_;
wire _68283_;
wire _68284_;
wire _68285_;
wire _68286_;
wire _68287_;
wire _68288_;
wire _68289_;
wire _68290_;
wire _68291_;
wire _68292_;
wire _68293_;
wire _68294_;
wire _68295_;
wire _68296_;
wire _68297_;
wire _68298_;
wire _68299_;
wire _68300_;
wire _68301_;
wire _68302_;
wire _68303_;
wire _68304_;
wire _68305_;
wire _68306_;
wire _68307_;
wire _68308_;
wire _68309_;
wire _68310_;
wire _68311_;
wire _68312_;
wire _68313_;
wire _68314_;
wire _68315_;
wire _68316_;
wire _68317_;
wire _68318_;
wire _68319_;
wire _68320_;
wire _68321_;
wire _68322_;
wire _68323_;
wire _68324_;
wire _68325_;
wire _68326_;
wire _68327_;
wire _68328_;
wire _68329_;
wire _68330_;
wire _68331_;
wire _68332_;
wire _68333_;
wire _68334_;
wire _68335_;
wire _68336_;
wire _68337_;
wire _68338_;
wire _68339_;
wire _68340_;
wire _68341_;
wire _68342_;
wire _68343_;
wire _68344_;
wire _68345_;
wire _68346_;
wire _68347_;
wire _68348_;
wire _68349_;
wire _68350_;
wire _68351_;
wire _68352_;
wire _68353_;
wire _68354_;
wire _68355_;
wire _68356_;
wire _68357_;
wire _68358_;
wire _68359_;
wire _68360_;
wire _68361_;
wire _68362_;
wire _68363_;
wire _68364_;
wire _68365_;
wire _68366_;
wire _68367_;
wire _68368_;
wire _68369_;
wire _68370_;
wire _68371_;
wire _68372_;
wire _68373_;
wire _68374_;
wire _68375_;
wire _68376_;
wire _68377_;
wire _68378_;
wire _68379_;
wire _68380_;
wire _68381_;
wire _68382_;
wire _68383_;
wire _68384_;
wire _68385_;
wire _68386_;
wire _68387_;
wire _68388_;
wire _68389_;
wire _68390_;
wire _68391_;
wire _68392_;
wire _68393_;
wire _68394_;
wire _68395_;
wire _68396_;
wire _68397_;
wire _68398_;
wire _68399_;
wire _68400_;
wire _68401_;
wire _68402_;
wire _68403_;
wire _68404_;
wire _68405_;
wire _68406_;
wire _68407_;
wire _68408_;
wire _68409_;
wire _68410_;
wire _68411_;
wire _68412_;
wire _68413_;
wire _68414_;
wire _68415_;
wire _68416_;
wire _68417_;
wire _68418_;
wire _68419_;
wire _68420_;
wire _68421_;
wire _68422_;
wire _68423_;
wire _68424_;
wire _68425_;
wire _68426_;
wire _68427_;
wire _68428_;
wire _68429_;
wire _68430_;
wire _68431_;
wire _68432_;
wire _68433_;
wire _68434_;
wire _68435_;
wire _68436_;
wire _68437_;
wire _68438_;
wire _68439_;
wire _68440_;
wire _68441_;
wire _68442_;
wire _68443_;
wire _68444_;
wire _68445_;
wire _68446_;
wire _68447_;
wire _68448_;
wire _68449_;
wire _68450_;
wire _68451_;
wire _68452_;
wire _68453_;
wire _68454_;
wire _68455_;
wire _68456_;
wire _68457_;
wire _68458_;
wire _68459_;
wire _68460_;
wire _68461_;
wire _68462_;
wire _68463_;
wire _68464_;
wire _68465_;
wire _68466_;
wire _68467_;
wire _68468_;
wire _68469_;
wire _68470_;
wire _68471_;
wire _68472_;
wire _68473_;
wire _68474_;
wire _68475_;
wire _68476_;
wire _68477_;
wire _68478_;
wire _68479_;
wire _68480_;
wire _68481_;
wire _68482_;
wire _68483_;
wire _68484_;
wire _68485_;
wire _68486_;
wire _68487_;
wire _68488_;
wire _68489_;
wire _68490_;
wire _68491_;
wire _68492_;
wire _68493_;
wire _68494_;
wire _68495_;
wire _68496_;
wire _68497_;
wire _68498_;
wire _68499_;
wire _68500_;
wire _68501_;
wire _68502_;
wire _68503_;
wire _68504_;
wire _68505_;
wire _68506_;
wire _68507_;
wire _68508_;
wire _68509_;
wire _68510_;
wire _68511_;
wire _68512_;
wire _68513_;
wire _68514_;
wire _68515_;
wire _68516_;
wire _68517_;
wire _68518_;
wire _68519_;
wire _68520_;
wire _68521_;
wire _68522_;
wire _68523_;
wire _68524_;
wire _68525_;
wire _68526_;
wire _68527_;
wire _68528_;
wire _68529_;
wire _68530_;
wire _68531_;
wire _68532_;
wire _68533_;
wire _68534_;
wire _68535_;
wire _68536_;
wire _68537_;
wire _68538_;
wire _68539_;
wire _68540_;
wire _68541_;
wire _68542_;
wire _68543_;
wire _68544_;
wire _68545_;
wire _68546_;
wire _68547_;
wire _68548_;
wire _68549_;
wire _68550_;
wire _68551_;
wire _68552_;
wire _68553_;
wire _68554_;
wire _68555_;
wire _68556_;
wire _68557_;
wire _68558_;
wire _68559_;
wire _68560_;
wire _68561_;
wire _68562_;
wire _68563_;
wire _68564_;
wire _68565_;
wire _68566_;
wire _68567_;
wire _68568_;
wire _68569_;
wire _68570_;
wire _68571_;
wire _68572_;
wire _68573_;
wire _68574_;
wire _68575_;
wire _68576_;
wire _68577_;
wire _68578_;
wire _68579_;
wire _68580_;
wire _68581_;
wire _68582_;
wire _68583_;
wire _68584_;
wire _68585_;
wire _68586_;
wire _68587_;
wire _68588_;
wire _68589_;
wire _68590_;
wire _68591_;
wire _68592_;
wire _68593_;
wire _68594_;
wire _68595_;
wire _68596_;
wire _68597_;
wire _68598_;
wire _68599_;
wire _68600_;
wire _68601_;
wire _68602_;
wire _68603_;
wire _68604_;
wire _68605_;
wire _68606_;
wire _68607_;
wire _68608_;
wire _68609_;
wire _68610_;
wire _68611_;
wire _68612_;
wire _68613_;
wire _68614_;
wire _68615_;
wire _68616_;
wire _68617_;
wire _68618_;
wire _68619_;
wire _68620_;
wire _68621_;
wire _68622_;
wire _68623_;
wire _68624_;
wire _68625_;
wire _68626_;
wire _68627_;
wire _68628_;
wire _68629_;
wire _68630_;
wire _68631_;
wire _68632_;
wire _68633_;
wire _68634_;
wire _68635_;
wire _68636_;
wire _68637_;
wire _68638_;
wire _68639_;
wire _68640_;
wire _68641_;
wire _68642_;
wire _68643_;
wire _68644_;
wire _68645_;
wire _68646_;
wire _68647_;
wire _68648_;
wire _68649_;
wire _68650_;
wire _68651_;
wire _68652_;
wire _68653_;
wire _68654_;
wire _68655_;
wire _68656_;
wire _68657_;
wire _68658_;
wire _68659_;
wire _68660_;
wire _68661_;
wire _68662_;
wire _68663_;
wire _68664_;
wire _68665_;
wire _68666_;
wire _68667_;
wire _68668_;
wire _68669_;
wire _68670_;
wire _68671_;
wire _68672_;
wire _68673_;
wire _68674_;
wire _68675_;
wire _68676_;
wire _68677_;
wire _68678_;
wire _68679_;
wire _68680_;
wire _68681_;
wire _68682_;
wire _68683_;
wire _68684_;
wire _68685_;
wire _68686_;
wire _68687_;
wire _68688_;
wire _68689_;
wire _68690_;
wire _68691_;
wire _68692_;
wire _68693_;
wire _68694_;
wire _68695_;
wire _68696_;
wire _68697_;
wire _68698_;
wire _68699_;
wire _68700_;
wire _68701_;
wire _68702_;
wire _68703_;
wire _68704_;
wire _68705_;
wire _68706_;
wire _68707_;
wire _68708_;
wire _68709_;
wire _68710_;
wire _68711_;
wire _68712_;
wire _68713_;
wire _68714_;
wire _68715_;
wire _68716_;
wire _68717_;
wire _68718_;
wire _68719_;
wire _68720_;
wire _68721_;
wire _68722_;
wire _68723_;
wire _68724_;
wire _68725_;
wire _68726_;
wire _68727_;
wire _68728_;
wire _68729_;
wire _68730_;
wire _68731_;
wire _68732_;
wire _68733_;
wire _68734_;
wire _68735_;
wire _68736_;
wire _68737_;
wire _68738_;
wire _68739_;
wire _68740_;
wire _68741_;
wire _68742_;
wire _68743_;
wire _68744_;
wire _68745_;
wire _68746_;
wire _68747_;
wire _68748_;
wire _68749_;
wire _68750_;
wire _68751_;
wire _68752_;
wire _68753_;
wire _68754_;
wire _68755_;
wire _68756_;
wire _68757_;
wire _68758_;
wire _68759_;
wire _68760_;
wire _68761_;
wire _68762_;
wire _68763_;
wire _68764_;
wire _68765_;
wire _68766_;
wire _68767_;
wire _68768_;
wire _68769_;
wire _68770_;
wire _68771_;
wire _68772_;
wire _68773_;
wire _68774_;
wire _68775_;
wire _68776_;
wire _68777_;
wire _68778_;
wire _68779_;
wire _68780_;
wire _68781_;
wire _68782_;
wire _68783_;
wire _68784_;
wire _68785_;
wire _68786_;
wire _68787_;
wire _68788_;
wire _68789_;
wire _68790_;
wire _68791_;
wire _68792_;
wire _68793_;
wire _68794_;
wire _68795_;
wire _68796_;
wire _68797_;
wire _68798_;
wire _68799_;
wire _68800_;
wire _68801_;
wire _68802_;
wire _68803_;
wire _68804_;
wire _68805_;
wire _68806_;
wire _68807_;
wire _68808_;
wire _68809_;
wire _68810_;
wire _68811_;
wire _68812_;
wire _68813_;
wire _68814_;
wire _68815_;
wire _68816_;
wire _68817_;
wire _68818_;
wire _68819_;
wire _68820_;
wire _68821_;
wire _68822_;
wire _68823_;
wire _68824_;
wire _68825_;
wire _68826_;
wire _68827_;
wire _68828_;
wire _68829_;
wire _68830_;
wire _68831_;
wire _68832_;
wire _68833_;
wire _68834_;
wire _68835_;
wire _68836_;
wire _68837_;
wire _68838_;
wire _68839_;
wire _68840_;
wire _68841_;
wire _68842_;
wire _68843_;
wire _68844_;
wire _68845_;
wire _68846_;
wire _68847_;
wire _68848_;
wire _68849_;
wire _68850_;
wire _68851_;
wire _68852_;
wire _68853_;
wire _68854_;
wire _68855_;
wire _68856_;
wire _68857_;
wire _68858_;
wire _68859_;
wire _68860_;
wire _68861_;
wire _68862_;
wire _68863_;
wire _68864_;
wire _68865_;
wire _68866_;
wire _68867_;
wire _68868_;
wire _68869_;
wire _68870_;
wire _68871_;
wire _68872_;
wire _68873_;
wire _68874_;
wire _68875_;
wire _68876_;
wire _68877_;
wire _68878_;
wire _68879_;
wire _68880_;
wire _68881_;
wire _68882_;
wire _68883_;
wire _68884_;
wire _68885_;
wire _68886_;
wire _68887_;
wire _68888_;
wire _68889_;
wire _68890_;
wire _68891_;
wire _68892_;
wire _68893_;
wire _68894_;
wire _68895_;
wire _68896_;
wire _68897_;
wire _68898_;
wire _68899_;
wire _68900_;
wire _68901_;
wire _68902_;
wire _68903_;
wire _68904_;
wire _68905_;
wire _68906_;
wire _68907_;
wire _68908_;
wire _68909_;
wire _68910_;
wire _68911_;
wire _68912_;
wire _68913_;
wire _68914_;
wire _68915_;
wire _68916_;
wire _68917_;
wire _68918_;
wire _68919_;
wire _68920_;
wire _68921_;
wire _68922_;
wire _68923_;
wire _68924_;
wire _68925_;
wire _68926_;
wire _68927_;
wire _68928_;
wire _68929_;
wire _68930_;
wire _68931_;
wire _68932_;
wire _68933_;
wire _68934_;
wire _68935_;
wire _68936_;
wire _68937_;
wire _68938_;
wire _68939_;
wire _68940_;
wire _68941_;
wire _68942_;
wire _68943_;
wire _68944_;
wire _68945_;
wire _68946_;
wire _68947_;
wire _68948_;
wire _68949_;
wire _68950_;
wire _68951_;
wire _68952_;
wire _68953_;
wire _68954_;
wire _68955_;
wire _68956_;
wire _68957_;
wire _68958_;
wire _68959_;
wire _68960_;
wire _68961_;
wire _68962_;
wire _68963_;
wire _68964_;
wire _68965_;
wire _68966_;
wire _68967_;
wire _68968_;
wire _68969_;
wire _68970_;
wire _68971_;
wire _68972_;
wire _68973_;
wire _68974_;
wire _68975_;
wire _68976_;
wire _68977_;
wire _68978_;
wire _68979_;
wire _68980_;
wire _68981_;
wire _68982_;
wire _68983_;
wire _68984_;
wire _68985_;
wire _68986_;
wire _68987_;
wire _68988_;
wire _68989_;
wire _68990_;
wire _68991_;
wire _68992_;
wire _68993_;
wire _68994_;
wire _68995_;
wire _68996_;
wire _68997_;
wire _68998_;
wire _68999_;
wire _69000_;
wire _69001_;
wire _69002_;
wire _69003_;
wire _69004_;
wire _69005_;
wire _69006_;
wire _69007_;
wire _69008_;
wire _69009_;
wire _69010_;
wire _69011_;
wire _69012_;
wire _69013_;
wire _69014_;
wire _69015_;
wire _69016_;
wire _69017_;
wire _69018_;
wire _69019_;
wire _69020_;
wire _69021_;
wire _69022_;
wire _69023_;
wire _69024_;
wire _69025_;
wire _69026_;
wire _69027_;
wire _69028_;
wire _69029_;
wire _69030_;
wire _69031_;
wire _69032_;
wire _69033_;
wire _69034_;
wire _69035_;
wire _69036_;
wire _69037_;
wire _69038_;
wire _69039_;
wire _69040_;
wire _69041_;
wire _69042_;
wire _69043_;
wire _69044_;
wire _69045_;
wire _69046_;
wire _69047_;
wire _69048_;
wire _69049_;
wire _69050_;
wire _69051_;
wire _69052_;
wire _69053_;
wire _69054_;
wire _69055_;
wire _69056_;
wire _69057_;
wire _69058_;
wire _69059_;
wire _69060_;
wire _69061_;
wire _69062_;
wire _69063_;
wire _69064_;
wire _69065_;
wire _69066_;
wire _69067_;
wire _69068_;
wire _69069_;
wire _69070_;
wire _69071_;
wire _69072_;
wire _69073_;
wire _69074_;
wire _69075_;
wire _69076_;
wire _69077_;
wire _69078_;
wire _69079_;
wire _69080_;
wire _69081_;
wire _69082_;
wire _69083_;
wire _69084_;
wire _69085_;
wire _69086_;
wire _69087_;
wire _69088_;
wire _69089_;
wire _69090_;
wire _69091_;
wire _69092_;
wire _69093_;
wire _69094_;
wire _69095_;
wire _69096_;
wire _69097_;
wire _69098_;
wire _69099_;
wire _69100_;
wire _69101_;
wire _69102_;
wire _69103_;
wire _69104_;
wire _69105_;
wire _69106_;
wire _69107_;
wire _69108_;
wire _69109_;
wire _69110_;
wire _69111_;
wire _69112_;
wire _69113_;
wire _69114_;
wire _69115_;
wire _69116_;
wire _69117_;
wire _69118_;
wire _69119_;
wire _69120_;
wire _69121_;
wire _69122_;
wire _69123_;
wire _69124_;
wire _69125_;
wire _69126_;
wire _69127_;
wire _69128_;
wire _69129_;
wire _69130_;
wire _69131_;
wire _69132_;
wire _69133_;
wire _69134_;
wire _69135_;
wire _69136_;
wire _69137_;
wire _69138_;
wire _69139_;
wire _69140_;
wire _69141_;
wire _69142_;
wire _69143_;
wire _69144_;
wire _69145_;
wire _69146_;
wire _69147_;
wire _69148_;
wire _69149_;
wire _69150_;
wire _69151_;
wire _69152_;
wire _69153_;
wire _69154_;
wire _69155_;
wire _69156_;
wire _69157_;
wire _69158_;
wire _69159_;
wire _69160_;
wire _69161_;
wire _69162_;
wire _69163_;
wire _69164_;
wire _69165_;
wire _69166_;
wire _69167_;
wire _69168_;
wire _69169_;
wire _69170_;
wire _69171_;
wire _69172_;
wire _69173_;
wire _69174_;
wire _69175_;
wire _69176_;
wire _69177_;
wire _69178_;
wire _69179_;
wire _69180_;
wire _69181_;
wire _69182_;
wire _69183_;
wire _69184_;
wire _69185_;
wire _69186_;
wire _69187_;
wire _69188_;
wire _69189_;
wire _69190_;
wire _69191_;
wire _69192_;
wire _69193_;
wire _69194_;
wire _69195_;
wire _69196_;
wire _69197_;
wire _69198_;
wire _69199_;
wire _69200_;
wire _69201_;
wire _69202_;
wire _69203_;
wire _69204_;
wire _69205_;
wire _69206_;
wire _69207_;
wire _69208_;
wire _69209_;
wire _69210_;
wire _69211_;
wire _69212_;
wire _69213_;
wire _69214_;
wire _69215_;
wire _69216_;
wire _69217_;
wire _69218_;
wire _69219_;
wire _69220_;
wire _69221_;
wire _69222_;
wire _69223_;
wire _69224_;
wire _69225_;
wire _69226_;
wire _69227_;
wire _69228_;
wire _69229_;
wire _69230_;
wire _69231_;
wire _69232_;
wire _69233_;
wire _69234_;
wire _69235_;
wire _69236_;
wire _69237_;
wire _69238_;
wire _69239_;
wire _69240_;
wire _69241_;
wire _69242_;
wire _69243_;
wire _69244_;
wire _69245_;
wire _69246_;
wire _69247_;
wire _69248_;
wire _69249_;
wire _69250_;
wire _69251_;
wire _69252_;
wire _69253_;
wire _69254_;
wire _69255_;
wire _69256_;
wire _69257_;
wire _69258_;
wire _69259_;
wire _69260_;
wire _69261_;
wire _69262_;
wire _69263_;
wire _69264_;
wire _69265_;
wire _69266_;
wire _69267_;
wire _69268_;
wire _69269_;
wire _69270_;
wire _69271_;
wire _69272_;
wire _69273_;
wire _69274_;
wire _69275_;
wire _69276_;
wire _69277_;
wire _69278_;
wire _69279_;
wire _69280_;
wire _69281_;
wire _69282_;
wire _69283_;
wire _69284_;
wire _69285_;
wire _69286_;
wire _69287_;
wire _69288_;
wire _69289_;
wire _69290_;
wire _69291_;
wire _69292_;
wire _69293_;
wire _69294_;
wire _69295_;
wire _69296_;
wire _69297_;
wire _69298_;
wire _69299_;
wire _69300_;
wire _69301_;
wire _69302_;
wire _69303_;
wire _69304_;
wire _69305_;
wire _69306_;
wire _69307_;
wire _69308_;
wire _69309_;
wire _69310_;
wire _69311_;
wire _69312_;
wire _69313_;
wire _69314_;
wire _69315_;
wire _69316_;
wire _69317_;
wire _69318_;
wire _69319_;
wire _69320_;
wire _69321_;
wire _69322_;
wire _69323_;
wire _69324_;
wire _69325_;
wire _69326_;
wire _69327_;
wire _69328_;
wire _69329_;
wire _69330_;
wire _69331_;
wire _69332_;
wire _69333_;
wire _69334_;
wire _69335_;
wire _69336_;
wire _69337_;
wire _69338_;
wire _69339_;
wire _69340_;
wire _69341_;
wire _69342_;
wire _69343_;
wire _69344_;
wire _69345_;
wire _69346_;
wire _69347_;
wire _69348_;
wire _69349_;
wire _69350_;
wire _69351_;
wire _69352_;
wire _69353_;
wire _69354_;
wire _69355_;
wire _69356_;
wire _69357_;
wire _69358_;
wire _69359_;
wire _69360_;
wire _69361_;
wire _69362_;
wire _69363_;
wire _69364_;
wire _69365_;
wire _69366_;
wire _69367_;
wire _69368_;
wire _69369_;
wire _69370_;
wire _69371_;
wire _69372_;
wire _69373_;
wire _69374_;
wire _69375_;
wire _69376_;
wire _69377_;
wire _69378_;
wire _69379_;
wire _69380_;
wire _69381_;
wire _69382_;
wire _69383_;
wire _69384_;
wire _69385_;
wire _69386_;
wire _69387_;
wire _69388_;
wire _69389_;
wire _69390_;
wire _69391_;
wire _69392_;
wire _69393_;
wire _69394_;
wire _69395_;
wire _69396_;
wire _69397_;
wire _69398_;
wire _69399_;
wire _69400_;
wire _69401_;
wire _69402_;
wire _69403_;
wire _69404_;
wire _69405_;
wire _69406_;
wire _69407_;
wire _69408_;
wire _69409_;
wire _69410_;
wire _69411_;
wire _69412_;
wire _69413_;
wire _69414_;
wire _69415_;
wire _69416_;
wire _69417_;
wire _69418_;
wire _69419_;
wire _69420_;
wire _69421_;
wire _69422_;
wire _69423_;
wire _69424_;
wire _69425_;
wire _69426_;
wire _69427_;
wire _69428_;
wire _69429_;
wire _69430_;
wire _69431_;
wire _69432_;
wire _69433_;
wire _69434_;
wire _69435_;
wire _69436_;
wire _69437_;
wire _69438_;
wire _69439_;
wire _69440_;
wire _69441_;
wire _69442_;
wire _69443_;
wire _69444_;
wire _69445_;
wire _69446_;
wire _69447_;
wire _69448_;
wire _69449_;
wire _69450_;
wire _69451_;
wire _69452_;
wire _69453_;
wire _69454_;
wire _69455_;
wire _69456_;
wire _69457_;
wire _69458_;
wire _69459_;
wire _69460_;
wire _69461_;
wire _69462_;
wire _69463_;
wire _69464_;
wire _69465_;
wire _69466_;
wire _69467_;
wire _69468_;
wire _69469_;
wire _69470_;
wire _69471_;
wire _69472_;
wire _69473_;
wire _69474_;
wire _69475_;
wire _69476_;
wire _69477_;
wire _69478_;
wire _69479_;
wire _69480_;
wire _69481_;
wire _69482_;
wire _69483_;
wire _69484_;
wire _69485_;
wire _69486_;
wire _69487_;
wire _69488_;
wire _69489_;
wire _69490_;
wire _69491_;
wire _69492_;
wire _69493_;
wire _69494_;
wire _69495_;
wire _69496_;
wire _69497_;
wire _69498_;
wire _69499_;
wire _69500_;
wire _69501_;
wire _69502_;
wire _69503_;
wire _69504_;
wire _69505_;
wire _69506_;
wire _69507_;
wire _69508_;
wire _69509_;
wire _69510_;
wire _69511_;
wire _69512_;
wire _69513_;
wire _69514_;
wire _69515_;
wire _69516_;
wire _69517_;
wire _69518_;
wire _69519_;
wire _69520_;
wire _69521_;
wire _69522_;
wire _69523_;
wire _69524_;
wire _69525_;
wire _69526_;
wire _69527_;
wire _69528_;
wire _69529_;
wire _69530_;
wire _69531_;
wire _69532_;
wire _69533_;
wire _69534_;
wire _69535_;
wire _69536_;
wire _69537_;
wire _69538_;
wire _69539_;
wire _69540_;
wire _69541_;
wire _69542_;
wire _69543_;
wire _69544_;
wire _69545_;
wire _69546_;
wire _69547_;
wire _69548_;
wire _69549_;
wire _69550_;
wire _69551_;
wire _69552_;
wire _69553_;
wire _69554_;
wire _69555_;
wire _69556_;
wire _69557_;
wire _69558_;
wire _69559_;
wire _69560_;
wire _69561_;
wire _69562_;
wire _69563_;
wire _69564_;
wire _69565_;
wire _69566_;
wire _69567_;
wire _69568_;
wire _69569_;
wire _69570_;
wire _69571_;
wire _69572_;
wire _69573_;
wire _69574_;
wire _69575_;
wire _69576_;
wire _69577_;
wire _69578_;
wire _69579_;
wire _69580_;
wire _69581_;
wire _69582_;
wire _69583_;
wire _69584_;
wire _69585_;
wire _69586_;
wire _69587_;
wire _69588_;
wire _69589_;
wire _69590_;
wire _69591_;
wire _69592_;
wire _69593_;
wire _69594_;
wire _69595_;
wire _69596_;
wire _69597_;
wire _69598_;
wire _69599_;
wire _69600_;
wire _69601_;
wire _69602_;
wire _69603_;
wire _69604_;
wire _69605_;
wire _69606_;
wire _69607_;
wire _69608_;
wire _69609_;
wire _69610_;
wire _69611_;
wire _69612_;
wire _69613_;
wire _69614_;
wire _69615_;
wire _69616_;
wire _69617_;
wire _69618_;
wire _69619_;
wire _69620_;
wire _69621_;
wire _69622_;
wire _69623_;
wire _69624_;
wire _69625_;
wire _69626_;
wire _69627_;
wire _69628_;
wire _69629_;
wire _69630_;
wire _69631_;
wire _69632_;
wire _69633_;
wire _69634_;
wire _69635_;
wire _69636_;
wire _69637_;
wire _69638_;
wire _69639_;
wire _69640_;
wire _69641_;
wire _69642_;
wire _69643_;
wire _69644_;
wire _69645_;
wire _69646_;
wire _69647_;
wire _69648_;
wire _69649_;
wire _69650_;
wire _69651_;
wire _69652_;
wire _69653_;
wire _69654_;
wire _69655_;
wire _69656_;
wire _69657_;
wire _69658_;
wire _69659_;
wire _69660_;
wire _69661_;
wire _69662_;
wire _69663_;
wire _69664_;
wire _69665_;
wire _69666_;
wire _69667_;
wire _69668_;
wire _69669_;
wire _69670_;
wire _69671_;
wire _69672_;
wire _69673_;
wire _69674_;
wire _69675_;
wire _69676_;
wire _69677_;
wire _69678_;
wire _69679_;
wire _69680_;
wire _69681_;
wire _69682_;
wire _69683_;
wire _69684_;
wire _69685_;
wire _69686_;
wire _69687_;
wire _69688_;
wire _69689_;
wire _69690_;
wire _69691_;
wire _69692_;
wire _69693_;
wire _69694_;
wire _69695_;
wire _69696_;
wire _69697_;
wire _69698_;
wire _69699_;
wire _69700_;
wire _69701_;
wire _69702_;
wire _69703_;
wire _69704_;
wire _69705_;
wire _69706_;
wire _69707_;
wire _69708_;
wire _69709_;
wire _69710_;
wire _69711_;
wire _69712_;
wire _69713_;
wire _69714_;
wire _69715_;
wire _69716_;
wire _69717_;
wire _69718_;
wire _69719_;
wire _69720_;
wire _69721_;
wire _69722_;
wire _69723_;
wire _69724_;
wire _69725_;
wire _69726_;
wire _69727_;
wire _69728_;
wire _69729_;
wire _69730_;
wire _69731_;
wire _69732_;
wire _69733_;
wire _69734_;
wire _69735_;
wire _69736_;
wire _69737_;
wire _69738_;
wire _69739_;
wire _69740_;
wire _69741_;
wire _69742_;
wire _69743_;
wire _69744_;
wire _69745_;
wire _69746_;
wire _69747_;
wire _69748_;
wire _69749_;
wire _69750_;
wire _69751_;
wire _69752_;
wire _69753_;
wire _69754_;
wire _69755_;
wire _69756_;
wire _69757_;
wire _69758_;
wire _69759_;
wire _69760_;
wire _69761_;
wire _69762_;
wire _69763_;
wire _69764_;
wire _69765_;
wire _69766_;
wire _69767_;
wire _69768_;
wire _69769_;
wire _69770_;
wire _69771_;
wire _69772_;
wire _69773_;
wire _69774_;
wire _69775_;
wire _69776_;
wire _69777_;
wire _69778_;
wire _69779_;
wire _69780_;
wire _69781_;
wire _69782_;
wire _69783_;
wire _69784_;
wire _69785_;
wire _69786_;
wire _69787_;
wire _69788_;
wire _69789_;
wire _69790_;
wire _69791_;
wire _69792_;
wire _69793_;
wire _69794_;
wire _69795_;
wire _69796_;
wire _69797_;
wire _69798_;
wire _69799_;
wire _69800_;
wire _69801_;
wire _69802_;
wire _69803_;
wire _69804_;
wire _69805_;
wire _69806_;
wire _69807_;
wire _69808_;
wire _69809_;
wire _69810_;
wire _69811_;
wire _69812_;
wire _69813_;
wire _69814_;
wire _69815_;
wire _69816_;
wire _69817_;
wire _69818_;
wire _69819_;
wire _69820_;
wire _69821_;
wire _69822_;
wire _69823_;
wire _69824_;
wire _69825_;
wire _69826_;
wire _69827_;
wire _69828_;
wire _69829_;
wire _69830_;
wire _69831_;
wire _69832_;
wire _69833_;
wire _69834_;
wire _69835_;
wire _69836_;
wire _69837_;
wire _69838_;
wire _69839_;
wire _69840_;
wire _69841_;
wire _69842_;
wire _69843_;
wire _69844_;
wire _69845_;
wire _69846_;
wire _69847_;
wire _69848_;
wire _69849_;
wire _69850_;
wire _69851_;
wire _69852_;
wire _69853_;
wire _69854_;
wire _69855_;
wire _69856_;
wire _69857_;
wire _69858_;
wire _69859_;
wire _69860_;
wire _69861_;
wire _69862_;
wire _69863_;
wire _69864_;
wire _69865_;
wire _69866_;
wire _69867_;
wire _69868_;
wire _69869_;
wire _69870_;
wire _69871_;
wire _69872_;
wire _69873_;
wire _69874_;
wire _69875_;
wire _69876_;
wire _69877_;
wire _69878_;
wire _69879_;
wire _69880_;
wire _69881_;
wire _69882_;
wire _69883_;
wire _69884_;
wire _69885_;
wire _69886_;
wire _69887_;
wire _69888_;
wire _69889_;
wire _69890_;
wire _69891_;
wire _69892_;
wire _69893_;
wire _69894_;
wire _69895_;
wire _69896_;
wire _69897_;
wire _69898_;
wire _69899_;
wire _69900_;
wire _69901_;
wire _69902_;
wire _69903_;
wire _69904_;
wire _69905_;
wire _69906_;
wire _69907_;
wire _69908_;
wire _69909_;
wire _69910_;
wire _69911_;
wire _69912_;
wire _69913_;
wire _69914_;
wire _69915_;
wire _69916_;
wire _69917_;
wire _69918_;
wire _69919_;
wire _69920_;
wire _69921_;
wire _69922_;
wire _69923_;
wire _69924_;
wire _69925_;
wire _69926_;
wire _69927_;
wire _69928_;
wire _69929_;
wire _69930_;
wire _69931_;
wire _69932_;
wire _69933_;
wire _69934_;
wire _69935_;
wire _69936_;
wire _69937_;
wire _69938_;
wire _69939_;
wire _69940_;
wire _69941_;
wire _69942_;
wire _69943_;
wire _69944_;
wire _69945_;
wire _69946_;
wire _69947_;
wire _69948_;
wire _69949_;
wire _69950_;
wire _69951_;
wire _69952_;
wire _69953_;
wire _69954_;
wire _69955_;
wire _69956_;
wire _69957_;
wire _69958_;
wire _69959_;
wire _69960_;
wire _69961_;
wire _69962_;
wire _69963_;
wire _69964_;
wire _69965_;
wire _69966_;
wire _69967_;
wire _69968_;
wire _69969_;
wire _69970_;
wire _69971_;
wire _69972_;
wire _69973_;
wire _69974_;
wire _69975_;
wire _69976_;
wire _69977_;
wire _69978_;
wire _69979_;
wire _69980_;
wire _69981_;
wire _69982_;
wire _69983_;
wire _69984_;
wire _69985_;
wire _69986_;
wire _69987_;
wire _69988_;
wire _69989_;
wire _69990_;
wire _69991_;
wire _69992_;
wire _69993_;
wire _69994_;
wire _69995_;
wire _69996_;
wire _69997_;
wire _69998_;
wire _69999_;
wire _70000_;
wire _70001_;
wire _70002_;
wire _70003_;
wire _70004_;
wire _70005_;
wire _70006_;
wire _70007_;
wire _70008_;
wire _70009_;
wire _70010_;
wire _70011_;
wire _70012_;
wire _70013_;
wire _70014_;
wire _70015_;
wire _70016_;
wire _70017_;
wire _70018_;
wire _70019_;
wire _70020_;
wire _70021_;
wire _70022_;
wire _70023_;
wire _70024_;
wire _70025_;
wire _70026_;
wire _70027_;
wire _70028_;
wire _70029_;
wire _70030_;
wire _70031_;
wire _70032_;
wire _70033_;
wire _70034_;
wire _70035_;
wire _70036_;
wire _70037_;
wire _70038_;
wire _70039_;
wire _70040_;
wire _70041_;
wire _70042_;
wire _70043_;
wire _70044_;
wire _70045_;
wire _70046_;
wire _70047_;
wire _70048_;
wire _70049_;
wire _70050_;
wire _70051_;
wire _70052_;
wire _70053_;
wire _70054_;
wire _70055_;
wire _70056_;
wire _70057_;
wire _70058_;
wire _70059_;
wire _70060_;
wire _70061_;
wire _70062_;
wire _70063_;
wire _70064_;
wire _70065_;
wire _70066_;
wire _70067_;
wire _70068_;
wire _70069_;
wire _70070_;
wire _70071_;
wire _70072_;
wire _70073_;
wire _70074_;
wire _70075_;
wire _70076_;
wire _70077_;
wire _70078_;
wire _70079_;
wire _70080_;
wire _70081_;
wire _70082_;
wire _70083_;
wire _70084_;
wire _70085_;
wire _70086_;
wire _70087_;
wire _70088_;
wire _70089_;
wire _70090_;
wire _70091_;
wire _70092_;
wire _70093_;
wire _70094_;
wire _70095_;
wire _70096_;
wire _70097_;
wire _70098_;
wire _70099_;
wire _70100_;
wire _70101_;
wire _70102_;
wire _70103_;
wire _70104_;
wire _70105_;
wire _70106_;
wire _70107_;
wire _70108_;
wire _70109_;
wire _70110_;
wire _70111_;
wire _70112_;
wire _70113_;
wire _70114_;
wire _70115_;
wire _70116_;
wire _70117_;
wire _70118_;
wire _70119_;
wire _70120_;
wire _70121_;
wire _70122_;
wire _70123_;
wire _70124_;
wire _70125_;
wire _70126_;
wire _70127_;
wire _70128_;
wire _70129_;
wire _70130_;
wire _70131_;
wire _70132_;
wire _70133_;
wire _70134_;
wire _70135_;
wire _70136_;
wire _70137_;
wire _70138_;
wire _70139_;
wire _70140_;
wire _70141_;
wire _70142_;
wire _70143_;
wire _70144_;
wire _70145_;
wire _70146_;
wire _70147_;
wire _70148_;
wire _70149_;
wire _70150_;
wire _70151_;
wire _70152_;
wire _70153_;
wire _70154_;
wire _70155_;
wire _70156_;
wire _70157_;
wire _70158_;
wire _70159_;
wire _70160_;
wire _70161_;
wire _70162_;
wire _70163_;
wire _70164_;
wire _70165_;
wire _70166_;
wire _70167_;
wire _70168_;
wire _70169_;
wire _70170_;
wire _70171_;
wire _70172_;
wire _70173_;
wire _70174_;
wire _70175_;
wire _70176_;
wire _70177_;
wire _70178_;
wire _70179_;
wire _70180_;
wire _70181_;
wire _70182_;
wire _70183_;
wire _70184_;
wire _70185_;
wire _70186_;
wire _70187_;
wire _70188_;
wire _70189_;
wire _70190_;
wire _70191_;
wire _70192_;
wire _70193_;
wire _70194_;
wire _70195_;
wire _70196_;
wire _70197_;
wire _70198_;
wire _70199_;
wire _70200_;
wire _70201_;
wire _70202_;
wire _70203_;
wire _70204_;
wire _70205_;
wire _70206_;
wire _70207_;
wire _70208_;
wire _70209_;
wire _70210_;
wire _70211_;
wire _70212_;
wire _70213_;
wire _70214_;
wire _70215_;
wire _70216_;
wire _70217_;
wire _70218_;
wire _70219_;
wire _70220_;
wire _70221_;
wire _70222_;
wire _70223_;
wire _70224_;
wire _70225_;
wire _70226_;
wire _70227_;
wire _70228_;
wire _70229_;
wire _70230_;
wire _70231_;
wire _70232_;
wire _70233_;
wire _70234_;
wire _70235_;
wire _70236_;
wire _70237_;
wire _70238_;
wire _70239_;
wire _70240_;
wire _70241_;
wire _70242_;
wire _70243_;
wire _70244_;
wire _70245_;
wire _70246_;
wire _70247_;
wire _70248_;
wire _70249_;
wire _70250_;
wire _70251_;
wire _70252_;
wire _70253_;
wire _70254_;
wire _70255_;
wire _70256_;
wire _70257_;
wire _70258_;
wire _70259_;
wire _70260_;
wire _70261_;
wire _70262_;
wire _70263_;
wire _70264_;
wire _70265_;
wire _70266_;
wire _70267_;
wire _70268_;
wire _70269_;
wire _70270_;
wire _70271_;
wire _70272_;
wire _70273_;
wire _70274_;
wire _70275_;
wire _70276_;
wire _70277_;
wire _70278_;
wire _70279_;
wire _70280_;
wire _70281_;
wire _70282_;
wire _70283_;
wire _70284_;
wire _70285_;
wire _70286_;
wire _70287_;
wire _70288_;
wire _70289_;
wire _70290_;
wire _70291_;
wire _70292_;
wire _70293_;
wire _70294_;
wire _70295_;
wire _70296_;
wire _70297_;
wire _70298_;
wire _70299_;
wire _70300_;
wire _70301_;
wire _70302_;
wire _70303_;
wire _70304_;
wire _70305_;
wire _70306_;
wire _70307_;
wire _70308_;
wire _70309_;
wire _70310_;
wire _70311_;
wire _70312_;
wire _70313_;
wire _70314_;
wire _70315_;
wire _70316_;
wire _70317_;
wire _70318_;
wire _70319_;
wire _70320_;
wire _70321_;
wire _70322_;
wire _70323_;
wire _70324_;
wire _70325_;
wire _70326_;
wire _70327_;
wire _70328_;
wire _70329_;
wire _70330_;
wire _70331_;
wire _70332_;
wire _70333_;
wire _70334_;
wire _70335_;
wire _70336_;
wire _70337_;
wire _70338_;
wire _70339_;
wire _70340_;
wire _70341_;
wire _70342_;
wire _70343_;
wire _70344_;
wire _70345_;
wire _70346_;
wire _70347_;
wire _70348_;
wire _70349_;
wire _70350_;
wire _70351_;
wire _70352_;
wire _70353_;
wire _70354_;
wire _70355_;
wire _70356_;
wire _70357_;
wire _70358_;
wire _70359_;
wire _70360_;
wire _70361_;
wire _70362_;
wire _70363_;
wire _70364_;
wire _70365_;
wire _70366_;
wire _70367_;
wire _70368_;
wire _70369_;
wire _70370_;
wire _70371_;
wire _70372_;
wire _70373_;
wire _70374_;
wire _70375_;
wire _70376_;
wire _70377_;
wire _70378_;
wire _70379_;
wire _70380_;
wire _70381_;
wire _70382_;
wire _70383_;
wire _70384_;
wire _70385_;
wire _70386_;
wire _70387_;
wire _70388_;
wire _70389_;
wire _70390_;
wire _70391_;
wire _70392_;
wire _70393_;
wire _70394_;
wire _70395_;
wire _70396_;
wire _70397_;
wire _70398_;
wire _70399_;
wire _70400_;
wire _70401_;
wire _70402_;
wire _70403_;
wire _70404_;
wire _70405_;
wire _70406_;
wire _70407_;
wire _70408_;
wire _70409_;
wire _70410_;
wire _70411_;
wire _70412_;
wire _70413_;
wire _70414_;
wire _70415_;
wire _70416_;
wire _70417_;
wire _70418_;
wire _70419_;
wire _70420_;
wire _70421_;
wire _70422_;
wire _70423_;
wire _70424_;
wire _70425_;
wire _70426_;
wire _70427_;
wire _70428_;
wire _70429_;
wire _70430_;
wire _70431_;
wire _70432_;
wire _70433_;
wire _70434_;
wire _70435_;
wire _70436_;
wire _70437_;
wire _70438_;
wire _70439_;
wire _70440_;
wire _70441_;
wire _70442_;
wire _70443_;
wire _70444_;
wire _70445_;
wire _70446_;
wire _70447_;
wire _70448_;
wire _70449_;
wire _70450_;
wire _70451_;
wire _70452_;
wire _70453_;
wire _70454_;
wire _70455_;
wire _70456_;
wire _70457_;
wire _70458_;
wire _70459_;
wire _70460_;
wire _70461_;
wire _70462_;
wire _70463_;
wire _70464_;
wire _70465_;
wire _70466_;
wire _70467_;
wire _70468_;
wire _70469_;
wire _70470_;
wire _70471_;
wire _70472_;
wire _70473_;
wire _70474_;
wire _70475_;
wire _70476_;
wire _70477_;
wire _70478_;
wire _70479_;
wire _70480_;
wire _70481_;
wire _70482_;
wire _70483_;
wire _70484_;
wire _70485_;
wire _70486_;
wire _70487_;
wire _70488_;
wire _70489_;
wire _70490_;
wire _70491_;
wire _70492_;
wire _70493_;
wire _70494_;
wire _70495_;
wire _70496_;
wire _70497_;
wire _70498_;
wire _70499_;
wire _70500_;
wire _70501_;
wire _70502_;
wire _70503_;
wire _70504_;
wire _70505_;
wire _70506_;
wire _70507_;
wire _70508_;
wire _70509_;
wire _70510_;
wire _70511_;
wire _70512_;
wire _70513_;
wire _70514_;
wire _70515_;
wire _70516_;
wire _70517_;
wire _70518_;
wire _70519_;
wire _70520_;
wire _70521_;
wire _70522_;
wire _70523_;
wire _70524_;
wire _70525_;
wire _70526_;
wire _70527_;
wire _70528_;
wire _70529_;
wire _70530_;
wire _70531_;
wire _70532_;
wire _70533_;
wire _70534_;
wire _70535_;
wire _70536_;
wire _70537_;
wire _70538_;
wire _70539_;
wire _70540_;
wire _70541_;
wire _70542_;
wire _70543_;
wire _70544_;
wire _70545_;
wire _70546_;
wire _70547_;
wire _70548_;
wire _70549_;
wire _70550_;
wire _70551_;
wire _70552_;
wire _70553_;
wire _70554_;
wire _70555_;
wire _70556_;
wire _70557_;
wire _70558_;
wire _70559_;
wire _70560_;
wire _70561_;
wire _70562_;
wire _70563_;
wire _70564_;
wire _70565_;
wire _70566_;
wire _70567_;
wire _70568_;
wire _70569_;
wire _70570_;
wire _70571_;
wire _70572_;
wire _70573_;
wire _70574_;
wire _70575_;
wire _70576_;
wire _70577_;
wire _70578_;
wire _70579_;
wire _70580_;
wire _70581_;
wire _70582_;
wire _70583_;
wire _70584_;
wire _70585_;
wire _70586_;
wire _70587_;
wire _70588_;
wire _70589_;
wire _70590_;
wire _70591_;
wire _70592_;
wire _70593_;
wire _70594_;
wire _70595_;
wire _70596_;
wire _70597_;
wire _70598_;
wire _70599_;
wire _70600_;
wire _70601_;
wire _70602_;
wire _70603_;
wire _70604_;
wire _70605_;
wire _70606_;
wire _70607_;
wire _70608_;
wire _70609_;
wire _70610_;
wire _70611_;
wire _70612_;
wire _70613_;
wire _70614_;
wire _70615_;
wire _70616_;
wire _70617_;
wire _70618_;
wire _70619_;
wire _70620_;
wire _70621_;
wire _70622_;
wire _70623_;
wire _70624_;
wire _70625_;
wire _70626_;
wire _70627_;
wire _70628_;
wire _70629_;
wire _70630_;
wire _70631_;
wire _70632_;
wire _70633_;
wire _70634_;
wire _70635_;
wire _70636_;
wire _70637_;
wire _70638_;
wire _70639_;
wire _70640_;
wire _70641_;
wire _70642_;
wire _70643_;
wire _70644_;
wire _70645_;
wire _70646_;
wire _70647_;
wire _70648_;
wire _70649_;
wire _70650_;
wire _70651_;
wire _70652_;
wire _70653_;
wire _70654_;
wire _70655_;
wire _70656_;
wire _70657_;
wire _70658_;
wire _70659_;
wire _70660_;
wire _70661_;
wire _70662_;
wire _70663_;
wire _70664_;
wire _70665_;
wire _70666_;
wire _70667_;
wire _70668_;
wire _70669_;
wire _70670_;
wire _70671_;
wire _70672_;
wire _70673_;
wire _70674_;
wire _70675_;
wire _70676_;
wire _70677_;
wire _70678_;
wire _70679_;
wire _70680_;
wire _70681_;
wire _70682_;
wire _70683_;
wire _70684_;
wire _70685_;
wire _70686_;
wire _70687_;
wire _70688_;
wire _70689_;
wire _70690_;
wire _70691_;
wire _70692_;
wire _70693_;
wire _70694_;
wire _70695_;
wire _70696_;
wire _70697_;
wire _70698_;
wire _70699_;
wire _70700_;
wire _70701_;
wire _70702_;
wire _70703_;
wire _70704_;
wire _70705_;
wire _70706_;
wire _70707_;
wire _70708_;
wire _70709_;
wire _70710_;
wire _70711_;
wire _70712_;
wire _70713_;
wire _70714_;
wire _70715_;
wire _70716_;
wire _70717_;
wire _70718_;
wire _70719_;
wire _70720_;
wire _70721_;
wire _70722_;
wire _70723_;
wire _70724_;
wire _70725_;
wire _70726_;
wire _70727_;
wire _70728_;
wire _70729_;
wire _70730_;
wire _70731_;
wire _70732_;
wire _70733_;
wire _70734_;
wire _70735_;
wire _70736_;
wire _70737_;
wire _70738_;
wire _70739_;
wire _70740_;
wire _70741_;
wire _70742_;
wire _70743_;
wire _70744_;
wire _70745_;
wire _70746_;
wire _70747_;
wire _70748_;
wire _70749_;
wire _70750_;
wire _70751_;
wire _70752_;
wire _70753_;
wire _70754_;
wire _70755_;
wire _70756_;
wire _70757_;
wire _70758_;
wire _70759_;
wire _70760_;
wire _70761_;
wire _70762_;
wire _70763_;
wire _70764_;
wire _70765_;
wire _70766_;
wire _70767_;
wire _70768_;
wire _70769_;
wire _70770_;
wire _70771_;
wire _70772_;
wire _70773_;
wire _70774_;
wire _70775_;
wire _70776_;
wire _70777_;
wire _70778_;
wire _70779_;
wire _70780_;
wire _70781_;
wire _70782_;
wire _70783_;
wire _70784_;
wire _70785_;
wire _70786_;
wire _70787_;
wire _70788_;
wire _70789_;
wire _70790_;
wire _70791_;
wire _70792_;
wire _70793_;
wire _70794_;
wire _70795_;
wire _70796_;
wire _70797_;
wire _70798_;
wire _70799_;
wire _70800_;
wire _70801_;
wire _70802_;
wire _70803_;
wire _70804_;
wire _70805_;
wire _70806_;
wire _70807_;
wire _70808_;
wire _70809_;
wire _70810_;
wire _70811_;
wire _70812_;
wire _70813_;
wire _70814_;
wire _70815_;
wire _70816_;
wire _70817_;
wire _70818_;
wire _70819_;
wire _70820_;
wire _70821_;
wire _70822_;
wire _70823_;
wire _70824_;
wire _70825_;
wire _70826_;
wire _70827_;
wire _70828_;
wire _70829_;
wire _70830_;
wire _70831_;
wire _70832_;
wire _70833_;
wire _70834_;
wire _70835_;
wire _70836_;
wire _70837_;
wire _70838_;
wire _70839_;
wire _70840_;
wire _70841_;
wire _70842_;
wire _70843_;
wire _70844_;
wire _70845_;
wire _70846_;
wire _70847_;
wire _70848_;
wire _70849_;
wire _70850_;
wire _70851_;
wire _70852_;
wire _70853_;
wire _70854_;
wire _70855_;
wire _70856_;
wire _70857_;
wire _70858_;
wire _70859_;
wire _70860_;
wire _70861_;
wire _70862_;
wire _70863_;
wire _70864_;
wire _70865_;
wire _70866_;
wire _70867_;
wire _70868_;
wire _70869_;
wire _70870_;
wire _70871_;
wire _70872_;
wire _70873_;
wire _70874_;
wire _70875_;
wire _70876_;
wire _70877_;
wire _70878_;
wire _70879_;
wire _70880_;
wire _70881_;
wire _70882_;
wire _70883_;
wire _70884_;
wire _70885_;
wire _70886_;
wire _70887_;
wire _70888_;
wire _70889_;
wire _70890_;
wire _70891_;
wire _70892_;
wire _70893_;
wire _70894_;
wire _70895_;
wire _70896_;
wire _70897_;
wire _70898_;
wire _70899_;
wire _70900_;
wire _70901_;
wire _70902_;
wire _70903_;
wire _70904_;
wire _70905_;
wire _70906_;
wire _70907_;
wire _70908_;
wire _70909_;
wire _70910_;
wire _70911_;
wire _70912_;
wire _70913_;
wire _70914_;
wire _70915_;
wire _70916_;
wire _70917_;
wire _70918_;
wire _70919_;
wire _70920_;
wire _70921_;
wire _70922_;
wire _70923_;
wire _70924_;
wire _70925_;
wire _70926_;
wire _70927_;
wire _70928_;
wire _70929_;
wire _70930_;
wire _70931_;
wire _70932_;
wire _70933_;
wire _70934_;
wire _70935_;
wire _70936_;
wire _70937_;
wire _70938_;
wire _70939_;
wire _70940_;
wire _70941_;
wire _70942_;
wire _70943_;
wire _70944_;
wire _70945_;
wire _70946_;
wire _70947_;
wire _70948_;
wire _70949_;
wire _70950_;
wire _70951_;
wire _70952_;
wire _70953_;
wire _70954_;
wire _70955_;
wire _70956_;
wire _70957_;
wire _70958_;
wire _70959_;
wire _70960_;
wire _70961_;
wire _70962_;
wire _70963_;
wire _70964_;
wire _70965_;
wire _70966_;
wire _70967_;
wire _70968_;
wire _70969_;
wire _70970_;
wire _70971_;
wire _70972_;
wire _70973_;
wire _70974_;
wire _70975_;
wire _70976_;
wire _70977_;
wire _70978_;
wire _70979_;
wire _70980_;
wire _70981_;
wire _70982_;
wire _70983_;
wire _70984_;
wire _70985_;
wire _70986_;
wire _70987_;
wire _70988_;
wire _70989_;
wire _70990_;
wire _70991_;
wire _70992_;
wire _70993_;
wire _70994_;
wire _70995_;
wire _70996_;
wire _70997_;
wire _70998_;
wire _70999_;
wire _71000_;
wire _71001_;
wire _71002_;
wire _71003_;
wire _71004_;
wire _71005_;
wire _71006_;
wire _71007_;
wire _71008_;
wire _71009_;
wire _71010_;
wire _71011_;
wire _71012_;
wire _71013_;
wire _71014_;
wire _71015_;
wire _71016_;
wire _71017_;
wire _71018_;
wire _71019_;
wire _71020_;
wire _71021_;
wire _71022_;
wire _71023_;
wire _71024_;
wire _71025_;
wire _71026_;
wire _71027_;
wire _71028_;
wire _71029_;
wire _71030_;
wire _71031_;
wire _71032_;
wire _71033_;
wire _71034_;
wire _71035_;
wire _71036_;
wire _71037_;
wire _71038_;
wire _71039_;
wire _71040_;
wire _71041_;
wire _71042_;
wire _71043_;
wire _71044_;
wire _71045_;
wire _71046_;
wire _71047_;
wire _71048_;
wire _71049_;
wire _71050_;
wire _71051_;
wire _71052_;
wire _71053_;
wire _71054_;
wire _71055_;
wire _71056_;
wire _71057_;
wire _71058_;
wire _71059_;
wire _71060_;
wire _71061_;
wire _71062_;
wire _71063_;
wire _71064_;
wire _71065_;
wire _71066_;
wire _71067_;
wire _71068_;
wire _71069_;
wire _71070_;
wire _71071_;
wire _71072_;
wire _71073_;
wire _71074_;
wire _71075_;
wire _71076_;
wire _71077_;
wire _71078_;
wire _71079_;
wire _71080_;
wire _71081_;
wire _71082_;
wire _71083_;
wire _71084_;
wire _71085_;
wire _71086_;
wire _71087_;
wire _71088_;
wire _71089_;
wire _71090_;
wire _71091_;
wire _71092_;
wire _71093_;
wire _71094_;
wire _71095_;
wire _71096_;
wire _71097_;
wire _71098_;
wire _71099_;
wire _71100_;
wire _71101_;
wire _71102_;
wire _71103_;
wire _71104_;
wire _71105_;
wire _71106_;
wire _71107_;
wire _71108_;
wire _71109_;
wire _71110_;
wire _71111_;
wire _71112_;
wire _71113_;
wire _71114_;
wire _71115_;
wire _71116_;
wire _71117_;
wire _71118_;
wire _71119_;
wire _71120_;
wire _71121_;
wire _71122_;
wire _71123_;
wire _71124_;
wire _71125_;
wire _71126_;
wire _71127_;
wire _71128_;
wire _71129_;
wire _71130_;
wire _71131_;
wire _71132_;
wire _71133_;
wire _71134_;
wire _71135_;
wire _71136_;
wire _71137_;
wire _71138_;
wire _71139_;
wire _71140_;
wire _71141_;
wire _71142_;
wire _71143_;
wire _71144_;
wire _71145_;
wire _71146_;
wire _71147_;
wire _71148_;
wire _71149_;
wire _71150_;
wire _71151_;
wire _71152_;
wire _71153_;
wire _71154_;
wire _71155_;
wire _71156_;
wire _71157_;
wire _71158_;
wire _71159_;
wire _71160_;
wire _71161_;
wire _71162_;
wire _71163_;
wire _71164_;
wire _71165_;
wire _71166_;
wire _71167_;
wire _71168_;
wire _71169_;
wire _71170_;
wire _71171_;
wire _71172_;
wire _71173_;
wire _71174_;
wire _71175_;
wire _71176_;
wire _71177_;
wire _71178_;
wire _71179_;
wire _71180_;
wire _71181_;
wire _71182_;
wire _71183_;
wire _71184_;
wire _71185_;
wire _71186_;
wire _71187_;
wire _71188_;
wire _71189_;
wire _71190_;
wire _71191_;
wire _71192_;
wire _71193_;
wire _71194_;
wire _71195_;
wire _71196_;
wire _71197_;
wire _71198_;
wire _71199_;
wire _71200_;
wire _71201_;
wire _71202_;
wire _71203_;
wire _71204_;
wire _71205_;
wire _71206_;
wire _71207_;
wire _71208_;
wire _71209_;
wire _71210_;
wire _71211_;
wire _71212_;
wire _71213_;
wire _71214_;
wire _71215_;
wire _71216_;
wire _71217_;
wire _71218_;
wire _71219_;
wire _71220_;
wire _71221_;
wire _71222_;
wire _71223_;
wire _71224_;
wire _71225_;
wire _71226_;
wire _71227_;
wire _71228_;
wire _71229_;
wire _71230_;
wire _71231_;
wire _71232_;
wire _71233_;
wire _71234_;
wire _71235_;
wire _71236_;
wire _71237_;
wire _71238_;
wire _71239_;
wire _71240_;
wire _71241_;
wire _71242_;
wire _71243_;
wire _71244_;
wire _71245_;
wire _71246_;
wire _71247_;
wire _71248_;
wire _71249_;
wire _71250_;
wire _71251_;
wire _71252_;
wire _71253_;
wire _71254_;
wire _71255_;
wire _71256_;
wire _71257_;
wire _71258_;
wire _71259_;
wire _71260_;
wire _71261_;
wire _71262_;
wire _71263_;
wire _71264_;
wire _71265_;
wire _71266_;
wire _71267_;
wire _71268_;
wire _71269_;
wire _71270_;
wire _71271_;
wire _71272_;
wire _71273_;
wire _71274_;
wire _71275_;
wire _71276_;
wire _71277_;
wire _71278_;
wire _71279_;
wire _71280_;
wire _71281_;
wire _71282_;
wire _71283_;
wire _71284_;
wire _71285_;
wire _71286_;
wire _71287_;
wire _71288_;
wire _71289_;
wire _71290_;
wire _71291_;
wire _71292_;
wire _71293_;
wire _71294_;
wire _71295_;
wire _71296_;
wire _71297_;
wire _71298_;
wire _71299_;
wire _71300_;
wire _71301_;
wire _71302_;
wire _71303_;
wire _71304_;
wire _71305_;
wire _71306_;
wire _71307_;
wire _71308_;
wire _71309_;
wire _71310_;
wire _71311_;
wire _71312_;
wire _71313_;
wire _71314_;
wire _71315_;
wire _71316_;
wire _71317_;
wire _71318_;
wire _71319_;
wire _71320_;
wire _71321_;
wire _71322_;
wire _71323_;
wire _71324_;
wire _71325_;
wire _71326_;
wire _71327_;
wire _71328_;
wire _71329_;
wire _71330_;
wire _71331_;
wire _71332_;
wire _71333_;
wire _71334_;
wire _71335_;
wire _71336_;
wire _71337_;
wire _71338_;
wire _71339_;
wire _71340_;
wire _71341_;
wire _71342_;
wire _71343_;
wire _71344_;
wire _71345_;
wire _71346_;
wire _71347_;
wire _71348_;
wire _71349_;
wire _71350_;
wire _71351_;
wire _71352_;
wire _71353_;
wire _71354_;
wire _71355_;
wire _71356_;
wire _71357_;
wire _71358_;
wire _71359_;
wire _71360_;
wire _71361_;
wire _71362_;
wire _71363_;
wire _71364_;
wire _71365_;
wire _71366_;
wire _71367_;
wire _71368_;
wire _71369_;
wire _71370_;
wire _71371_;
wire _71372_;
wire _71373_;
wire _71374_;
wire _71375_;
wire _71376_;
wire _71377_;
wire _71378_;
wire _71379_;
wire _71380_;
wire _71381_;
wire _71382_;
wire _71383_;
wire _71384_;
wire _71385_;
wire _71386_;
wire _71387_;
wire _71388_;
wire _71389_;
wire _71390_;
wire _71391_;
wire _71392_;
wire _71393_;
wire _71394_;
wire _71395_;
wire _71396_;
wire _71397_;
wire _71398_;
wire _71399_;
wire _71400_;
wire _71401_;
wire _71402_;
wire _71403_;
wire _71404_;
wire _71405_;
wire _71406_;
wire _71407_;
wire _71408_;
wire _71409_;
wire _71410_;
wire _71411_;
wire _71412_;
wire _71413_;
wire _71414_;
wire _71415_;
wire _71416_;
wire _71417_;
wire _71418_;
wire _71419_;
wire _71420_;
wire _71421_;
wire _71422_;
wire _71423_;
wire _71424_;
wire _71425_;
wire _71426_;
wire _71427_;
wire _71428_;
wire _71429_;
wire _71430_;
wire _71431_;
wire _71432_;
wire _71433_;
wire _71434_;
wire _71435_;
wire _71436_;
wire _71437_;
wire _71438_;
wire _71439_;
wire _71440_;
wire _71441_;
wire _71442_;
wire _71443_;
wire _71444_;
wire _71445_;
wire _71446_;
wire _71447_;
wire _71448_;
wire _71449_;
wire _71450_;
wire _71451_;
wire _71452_;
wire _71453_;
wire _71454_;
wire _71455_;
wire _71456_;
wire _71457_;
wire _71458_;
wire _71459_;
wire _71460_;
wire _71461_;
wire _71462_;
wire _71463_;
wire _71464_;
wire _71465_;
wire _71466_;
wire _71467_;
wire _71468_;
wire _71469_;
wire _71470_;
wire _71471_;
wire _71472_;
wire _71473_;
wire _71474_;
wire _71475_;
wire _71476_;
wire _71477_;
wire _71478_;
wire _71479_;
wire _71480_;
wire _71481_;
wire _71482_;
wire _71483_;
wire _71484_;
wire _71485_;
wire _71486_;
wire _71487_;
wire _71488_;
wire _71489_;
wire _71490_;
wire _71491_;
wire _71492_;
wire _71493_;
wire _71494_;
wire _71495_;
wire _71496_;
wire _71497_;
wire _71498_;
wire _71499_;
wire _71500_;
wire _71501_;
wire _71502_;
wire _71503_;
wire _71504_;
wire _71505_;
wire _71506_;
wire _71507_;
wire _71508_;
wire _71509_;
wire _71510_;
wire _71511_;
wire _71512_;
wire _71513_;
wire _71514_;
wire _71515_;
wire _71516_;
wire _71517_;
wire _71518_;
wire _71519_;
wire _71520_;
wire _71521_;
wire _71522_;
wire _71523_;
wire _71524_;
wire _71525_;
wire _71526_;
wire _71527_;
wire _71528_;
wire _71529_;
wire _71530_;
wire _71531_;
wire _71532_;
wire _71533_;
wire _71534_;
wire _71535_;
wire _71536_;
wire _71537_;
wire _71538_;
wire _71539_;
wire _71540_;
wire _71541_;
wire _71542_;
wire _71543_;
wire _71544_;
wire _71545_;
wire _71546_;
wire _71547_;
wire _71548_;
wire _71549_;
wire _71550_;
wire _71551_;
wire _71552_;
wire _71553_;
wire _71554_;
wire _71555_;
wire _71556_;
wire _71557_;
wire _71558_;
wire _71559_;
wire _71560_;
wire _71561_;
wire _71562_;
wire _71563_;
wire _71564_;
wire _71565_;
wire _71566_;
wire _71567_;
wire _71568_;
wire _71569_;
wire _71570_;
wire _71571_;
wire _71572_;
wire _71573_;
wire _71574_;
wire _71575_;
wire _71576_;
wire _71577_;
wire _71578_;
wire _71579_;
wire _71580_;
wire _71581_;
wire _71582_;
wire _71583_;
wire _71584_;
wire _71585_;
wire _71586_;
wire _71587_;
wire _71588_;
wire _71589_;
wire _71590_;
wire _71591_;
wire _71592_;
wire _71593_;
wire _71594_;
wire _71595_;
wire _71596_;
wire _71597_;
wire _71598_;
wire _71599_;
wire _71600_;
wire _71601_;
wire _71602_;
wire _71603_;
wire _71604_;
wire _71605_;
wire _71606_;
wire _71607_;
wire _71608_;
wire _71609_;
wire _71610_;
wire _71611_;
wire _71612_;
wire _71613_;
wire _71614_;
wire _71615_;
wire _71616_;
wire _71617_;
wire _71618_;
wire _71619_;
wire _71620_;
wire _71621_;
wire _71622_;
wire _71623_;
wire _71624_;
wire _71625_;
wire _71626_;
wire _71627_;
wire _71628_;
wire _71629_;
wire _71630_;
wire _71631_;
wire _71632_;
wire _71633_;
wire _71634_;
wire _71635_;
wire _71636_;
wire _71637_;
wire _71638_;
wire _71639_;
wire _71640_;
wire _71641_;
wire _71642_;
wire _71643_;
wire _71644_;
wire _71645_;
wire _71646_;
wire _71647_;
wire _71648_;
wire _71649_;
wire _71650_;
wire _71651_;
wire _71652_;
wire _71653_;
wire _71654_;
wire _71655_;
wire _71656_;
wire _71657_;
wire _71658_;
wire _71659_;
wire _71660_;
wire _71661_;
wire _71662_;
wire _71663_;
wire _71664_;
wire _71665_;
wire _71666_;
wire _71667_;
wire _71668_;
wire _71669_;
wire _71670_;
wire _71671_;
wire _71672_;
wire _71673_;
wire _71674_;
wire _71675_;
wire _71676_;
wire _71677_;
wire _71678_;
wire _71679_;
wire _71680_;
wire _71681_;
wire _71682_;
wire _71683_;
wire _71684_;
wire _71685_;
wire _71686_;
wire _71687_;
wire _71688_;
wire _71689_;
wire _71690_;
wire _71691_;
wire _71692_;
wire _71693_;
wire _71694_;
wire _71695_;
wire _71696_;
wire _71697_;
wire _71698_;
wire _71699_;
wire _71700_;
wire _71701_;
wire _71702_;
wire _71703_;
wire _71704_;
wire _71705_;
wire _71706_;
wire _71707_;
wire _71708_;
wire _71709_;
wire _71710_;
wire _71711_;
wire _71712_;
wire _71713_;
wire _71714_;
wire _71715_;
wire _71716_;
wire _71717_;
wire _71718_;
wire _71719_;
wire _71720_;
wire _71721_;
wire _71722_;
wire _71723_;
wire _71724_;
wire _71725_;
wire _71726_;
wire _71727_;
wire _71728_;
wire _71729_;
wire _71730_;
wire _71731_;
wire _71732_;
wire _71733_;
wire _71734_;
wire _71735_;
wire _71736_;
wire _71737_;
wire _71738_;
wire _71739_;
wire _71740_;
wire _71741_;
wire _71742_;
wire _71743_;
wire _71744_;
wire _71745_;
wire _71746_;
wire _71747_;
wire _71748_;
wire _71749_;
wire _71750_;
wire _71751_;
wire _71752_;
wire _71753_;
wire _71754_;
wire _71755_;
wire _71756_;
wire _71757_;
wire _71758_;
wire _71759_;
wire _71760_;
wire _71761_;
wire _71762_;
wire _71763_;
wire _71764_;
wire _71765_;
wire _71766_;
wire _71767_;
wire _71768_;
wire _71769_;
wire _71770_;
wire _71771_;
wire _71772_;
wire _71773_;
wire _71774_;
wire _71775_;
wire _71776_;
wire _71777_;
wire _71778_;
wire _71779_;
wire _71780_;
wire _71781_;
wire _71782_;
wire _71783_;
wire _71784_;
wire _71785_;
wire _71786_;
wire _71787_;
wire _71788_;
wire _71789_;
wire _71790_;
wire _71791_;
wire _71792_;
wire _71793_;
wire _71794_;
wire _71795_;
wire _71796_;
wire _71797_;
wire _71798_;
wire _71799_;
wire _71800_;
wire _71801_;
wire _71802_;
wire _71803_;
wire _71804_;
wire _71805_;
wire _71806_;
wire _71807_;
wire _71808_;
wire _71809_;
wire _71810_;
wire _71811_;
wire _71812_;
wire _71813_;
wire _71814_;
wire _71815_;
wire _71816_;
wire _71817_;
wire _71818_;
wire _71819_;
wire _71820_;
wire _71821_;
wire _71822_;
wire _71823_;
wire _71824_;
wire _71825_;
wire _71826_;
wire _71827_;
wire _71828_;
wire _71829_;
wire _71830_;
wire _71831_;
wire _71832_;
wire _71833_;
wire _71834_;
wire _71835_;
wire _71836_;
wire _71837_;
wire _71838_;
wire _71839_;
wire _71840_;
wire _71841_;
wire _71842_;
wire _71843_;
wire _71844_;
wire _71845_;
wire _71846_;
wire _71847_;
wire _71848_;
wire _71849_;
wire _71850_;
wire _71851_;
wire _71852_;
wire _71853_;
wire _71854_;
wire _71855_;
wire _71856_;
wire _71857_;
wire _71858_;
wire _71859_;
wire _71860_;
wire _71861_;
wire _71862_;
wire _71863_;
wire _71864_;
wire _71865_;
wire _71866_;
wire _71867_;
wire _71868_;
wire _71869_;
wire _71870_;
wire _71871_;
wire _71872_;
wire _71873_;
wire _71874_;
wire _71875_;
wire _71876_;
wire _71877_;
wire _71878_;
wire _71879_;
wire _71880_;
wire _71881_;
wire _71882_;
wire _71883_;
wire _71884_;
wire _71885_;
wire _71886_;
wire _71887_;
wire _71888_;
wire _71889_;
wire _71890_;
wire _71891_;
wire _71892_;
wire _71893_;
wire _71894_;
wire _71895_;
wire _71896_;
wire _71897_;
wire _71898_;
wire _71899_;
wire _71900_;
wire _71901_;
wire _71902_;
wire _71903_;
wire _71904_;
wire _71905_;
wire _71906_;
wire _71907_;
wire _71908_;
wire _71909_;
wire _71910_;
wire _71911_;
wire _71912_;
wire _71913_;
wire _71914_;
wire _71915_;
wire _71916_;
wire _71917_;
wire _71918_;
wire _71919_;
wire _71920_;
wire _71921_;
wire _71922_;
wire _71923_;
wire _71924_;
wire _71925_;
wire _71926_;
wire _71927_;
wire _71928_;
wire _71929_;
wire _71930_;
wire _71931_;
wire _71932_;
wire _71933_;
wire _71934_;
wire _71935_;
wire _71936_;
wire _71937_;
wire _71938_;
wire _71939_;
wire _71940_;
wire _71941_;
wire _71942_;
wire _71943_;
wire _71944_;
wire _71945_;
wire _71946_;
wire _71947_;
wire _71948_;
wire _71949_;
wire _71950_;
wire _71951_;
wire _71952_;
wire _71953_;
wire _71954_;
wire _71955_;
wire _71956_;
wire _71957_;
wire _71958_;
wire _71959_;
wire _71960_;
wire _71961_;
wire _71962_;
wire _71963_;
wire _71964_;
wire _71965_;
wire _71966_;
wire _71967_;
wire _71968_;
wire _71969_;
wire _71970_;
wire _71971_;
wire _71972_;
wire _71973_;
wire _71974_;
wire _71975_;
wire _71976_;
wire _71977_;
wire _71978_;
wire _71979_;
wire _71980_;
wire _71981_;
wire _71982_;
wire _71983_;
wire _71984_;
wire _71985_;
wire _71986_;
wire _71987_;
wire _71988_;
wire _71989_;
wire _71990_;
wire _71991_;
wire _71992_;
wire _71993_;
wire _71994_;
wire _71995_;
wire _71996_;
wire _71997_;
wire _71998_;
wire _71999_;
wire _72000_;
wire _72001_;
wire _72002_;
wire _72003_;
wire _72004_;
wire _72005_;
wire _72006_;
wire _72007_;
wire _72008_;
wire _72009_;
wire _72010_;
wire _72011_;
wire _72012_;
wire _72013_;
wire _72014_;
wire _72015_;
wire _72016_;
wire _72017_;
wire _72018_;
wire _72019_;
wire _72020_;
wire _72021_;
wire _72022_;
wire _72023_;
wire _72024_;
wire _72025_;
wire _72026_;
wire _72027_;
wire _72028_;
wire _72029_;
wire _72030_;
wire _72031_;
wire _72032_;
wire _72033_;
wire _72034_;
wire _72035_;
wire _72036_;
wire _72037_;
wire _72038_;
wire _72039_;
wire _72040_;
wire _72041_;
wire _72042_;
wire _72043_;
wire _72044_;
wire _72045_;
wire _72046_;
wire _72047_;
wire _72048_;
wire _72049_;
wire _72050_;
wire _72051_;
wire _72052_;
wire _72053_;
wire _72054_;
wire _72055_;
wire _72056_;
wire _72057_;
wire _72058_;
wire _72059_;
wire _72060_;
wire _72061_;
wire _72062_;
wire _72063_;
wire _72064_;
wire _72065_;
wire _72066_;
wire _72067_;
wire _72068_;
wire _72069_;
wire _72070_;
wire _72071_;
wire _72072_;
wire _72073_;
wire _72074_;
wire _72075_;
wire _72076_;
wire _72077_;
wire _72078_;
wire _72079_;
wire _72080_;
wire _72081_;
wire _72082_;
wire _72083_;
wire _72084_;
wire _72085_;
wire _72086_;
wire _72087_;
wire _72088_;
wire _72089_;
wire _72090_;
wire _72091_;
wire _72092_;
wire _72093_;
wire _72094_;
wire _72095_;
wire _72096_;
wire _72097_;
wire _72098_;
wire _72099_;
wire _72100_;
wire _72101_;
wire _72102_;
wire _72103_;
wire _72104_;
wire _72105_;
wire _72106_;
wire _72107_;
wire _72108_;
wire _72109_;
wire _72110_;
wire _72111_;
wire _72112_;
wire _72113_;
wire _72114_;
wire _72115_;
wire _72116_;
wire _72117_;
wire _72118_;
wire _72119_;
wire _72120_;
wire _72121_;
wire _72122_;
wire _72123_;
wire _72124_;
wire _72125_;
wire _72126_;
wire _72127_;
wire _72128_;
wire _72129_;
wire _72130_;
wire _72131_;
wire _72132_;
wire _72133_;
wire _72134_;
wire _72135_;
wire _72136_;
wire _72137_;
wire _72138_;
wire _72139_;
wire _72140_;
wire _72141_;
wire _72142_;
wire _72143_;
wire _72144_;
wire _72145_;
wire _72146_;
wire _72147_;
wire _72148_;
wire _72149_;
wire _72150_;
wire _72151_;
wire _72152_;
wire _72153_;
wire _72154_;
wire _72155_;
wire _72156_;
wire _72157_;
wire _72158_;
wire _72159_;
wire _72160_;
wire _72161_;
wire _72162_;
wire _72163_;
wire _72164_;
wire _72165_;
wire _72166_;
wire _72167_;
wire _72168_;
wire _72169_;
wire _72170_;
wire _72171_;
wire _72172_;
wire _72173_;
wire _72174_;
wire _72175_;
wire _72176_;
wire _72177_;
wire _72178_;
wire _72179_;
wire _72180_;
wire _72181_;
wire _72182_;
wire _72183_;
wire _72184_;
wire _72185_;
wire _72186_;
wire _72187_;
wire _72188_;
wire _72189_;
wire _72190_;
wire _72191_;
wire _72192_;
wire _72193_;
wire _72194_;
wire _72195_;
wire _72196_;
wire _72197_;
wire _72198_;
wire _72199_;
wire _72200_;
wire _72201_;
wire _72202_;
wire _72203_;
wire _72204_;
wire _72205_;
wire _72206_;
wire _72207_;
wire _72208_;
wire _72209_;
wire _72210_;
wire _72211_;
wire _72212_;
wire _72213_;
wire _72214_;
wire _72215_;
wire _72216_;
wire _72217_;
wire _72218_;
wire _72219_;
wire _72220_;
wire _72221_;
wire _72222_;
wire _72223_;
wire _72224_;
wire _72225_;
wire _72226_;
wire _72227_;
wire _72228_;
wire _72229_;
wire _72230_;
wire _72231_;
wire _72232_;
wire _72233_;
wire _72234_;
wire _72235_;
wire _72236_;
wire _72237_;
wire _72238_;
wire _72239_;
wire _72240_;
wire _72241_;
wire _72242_;
wire _72243_;
wire _72244_;
wire _72245_;
wire _72246_;
wire _72247_;
wire _72248_;
wire _72249_;
wire _72250_;
wire _72251_;
wire _72252_;
wire _72253_;
wire _72254_;
wire _72255_;
wire _72256_;
wire _72257_;
wire _72258_;
wire _72259_;
wire _72260_;
wire _72261_;
wire _72262_;
wire _72263_;
wire _72264_;
wire _72265_;
wire _72266_;
wire _72267_;
wire _72268_;
wire _72269_;
wire _72270_;
wire _72271_;
wire _72272_;
wire _72273_;
wire _72274_;
wire _72275_;
wire _72276_;
wire _72277_;
wire _72278_;
wire _72279_;
wire _72280_;
wire _72281_;
wire _72282_;
wire _72283_;
wire _72284_;
wire _72285_;
wire _72286_;
wire _72287_;
wire _72288_;
wire _72289_;
wire _72290_;
wire _72291_;
wire _72292_;
wire _72293_;
wire _72294_;
wire _72295_;
wire _72296_;
wire _72297_;
wire _72298_;
wire _72299_;
wire _72300_;
wire _72301_;
wire _72302_;
wire _72303_;
wire _72304_;
wire _72305_;
wire _72306_;
wire _72307_;
wire _72308_;
wire _72309_;
wire _72310_;
wire _72311_;
wire _72312_;
wire _72313_;
wire _72314_;
wire _72315_;
wire _72316_;
wire _72317_;
wire _72318_;
wire _72319_;
wire _72320_;
wire _72321_;
wire _72322_;
wire _72323_;
wire _72324_;
wire _72325_;
wire _72326_;
wire _72327_;
wire _72328_;
wire _72329_;
wire _72330_;
wire _72331_;
wire _72332_;
wire _72333_;
wire _72334_;
wire _72335_;
wire _72336_;
wire _72337_;
wire _72338_;
wire _72339_;
wire _72340_;
wire _72341_;
wire _72342_;
wire _72343_;
wire _72344_;
wire _72345_;
wire _72346_;
wire _72347_;
wire _72348_;
wire _72349_;
wire _72350_;
wire _72351_;
wire _72352_;
wire _72353_;
wire _72354_;
wire _72355_;
wire _72356_;
wire _72357_;
wire _72358_;
wire _72359_;
wire _72360_;
wire _72361_;
wire _72362_;
wire _72363_;
wire _72364_;
wire _72365_;
wire _72366_;
wire _72367_;
wire _72368_;
wire _72369_;
wire _72370_;
wire _72371_;
wire _72372_;
wire _72373_;
wire _72374_;
wire _72375_;
wire _72376_;
wire _72377_;
wire _72378_;
wire _72379_;
wire _72380_;
wire _72381_;
wire _72382_;
wire _72383_;
wire _72384_;
wire _72385_;
wire _72386_;
wire _72387_;
wire _72388_;
wire _72389_;
wire _72390_;
wire _72391_;
wire _72392_;
wire _72393_;
wire _72394_;
wire _72395_;
wire _72396_;
wire _72397_;
wire _72398_;
wire _72399_;
wire _72400_;
wire _72401_;
wire _72402_;
wire _72403_;
wire _72404_;
wire _72405_;
wire _72406_;
wire _72407_;
wire _72408_;
wire _72409_;
wire _72410_;
wire _72411_;
wire _72412_;
wire _72413_;
wire _72414_;
wire _72415_;
wire _72416_;
wire _72417_;
wire _72418_;
wire _72419_;
wire _72420_;
wire _72421_;
wire _72422_;
wire _72423_;
wire _72424_;
wire _72425_;
wire _72426_;
wire _72427_;
wire _72428_;
wire _72429_;
wire _72430_;
wire _72431_;
wire _72432_;
wire _72433_;
wire _72434_;
wire _72435_;
wire _72436_;
wire _72437_;
wire _72438_;
wire _72439_;
wire _72440_;
wire _72441_;
wire _72442_;
wire _72443_;
wire _72444_;
wire _72445_;
wire _72446_;
wire _72447_;
wire _72448_;
wire _72449_;
wire _72450_;
wire _72451_;
wire _72452_;
wire _72453_;
wire _72454_;
wire _72455_;
wire _72456_;
wire _72457_;
wire _72458_;
wire _72459_;
wire _72460_;
wire _72461_;
wire _72462_;
wire _72463_;
wire _72464_;
wire _72465_;
wire _72466_;
wire _72467_;
wire _72468_;
wire _72469_;
wire _72470_;
wire _72471_;
wire _72472_;
wire _72473_;
wire _72474_;
wire _72475_;
wire _72476_;
wire _72477_;
wire _72478_;
wire _72479_;
wire _72480_;
wire _72481_;
wire _72482_;
wire _72483_;
wire _72484_;
wire _72485_;
wire _72486_;
wire _72487_;
wire _72488_;
wire _72489_;
wire _72490_;
wire _72491_;
wire _72492_;
wire _72493_;
wire _72494_;
wire _72495_;
wire _72496_;
wire _72497_;
wire _72498_;
wire _72499_;
wire _72500_;
wire _72501_;
wire _72502_;
wire _72503_;
wire _72504_;
wire _72505_;
wire _72506_;
wire _72507_;
wire _72508_;
wire _72509_;
wire _72510_;
wire _72511_;
wire _72512_;
wire _72513_;
wire _72514_;
wire _72515_;
wire _72516_;
wire _72517_;
wire _72518_;
wire _72519_;
wire _72520_;
wire _72521_;
wire _72522_;
wire _72523_;
wire _72524_;
wire _72525_;
wire _72526_;
wire _72527_;
wire _72528_;
wire _72529_;
wire _72530_;
wire _72531_;
wire _72532_;
wire _72533_;
wire _72534_;
wire _72535_;
wire _72536_;
wire _72537_;
wire _72538_;
wire _72539_;
wire _72540_;
wire _72541_;
wire _72542_;
wire _72543_;
wire _72544_;
wire _72545_;
wire _72546_;
wire _72547_;
wire _72548_;
wire _72549_;
wire _72550_;
wire _72551_;
wire _72552_;
wire _72553_;
wire _72554_;
wire _72555_;
wire _72556_;
wire _72557_;
wire _72558_;
wire _72559_;
wire _72560_;
wire _72561_;
wire _72562_;
wire _72563_;
wire _72564_;
wire _72565_;
wire _72566_;
wire _72567_;
wire _72568_;
wire _72569_;
wire _72570_;
wire _72571_;
wire _72572_;
wire _72573_;
wire _72574_;
wire _72575_;
wire _72576_;
wire _72577_;
wire _72578_;
wire _72579_;
wire _72580_;
wire _72581_;
wire _72582_;
wire _72583_;
wire _72584_;
wire _72585_;
wire _72586_;
wire _72587_;
wire _72588_;
wire _72589_;
wire _72590_;
wire _72591_;
wire _72592_;
wire _72593_;
wire _72594_;
wire _72595_;
wire _72596_;
wire _72597_;
wire _72598_;
wire _72599_;
wire _72600_;
wire _72601_;
wire _72602_;
wire _72603_;
wire _72604_;
wire _72605_;
wire _72606_;
wire _72607_;
wire _72608_;
wire _72609_;
wire _72610_;
wire _72611_;
wire _72612_;
wire _72613_;
wire _72614_;
wire _72615_;
wire _72616_;
wire _72617_;
wire _72618_;
wire _72619_;
wire _72620_;
wire _72621_;
wire _72622_;
wire _72623_;
wire _72624_;
wire _72625_;
wire _72626_;
wire _72627_;
wire _72628_;
wire _72629_;
wire _72630_;
wire _72631_;
wire _72632_;
wire _72633_;
wire _72634_;
wire _72635_;
wire _72636_;
wire _72637_;
wire _72638_;
wire _72639_;
wire _72640_;
wire _72641_;
wire _72642_;
wire _72643_;
wire _72644_;
wire _72645_;
wire _72646_;
wire _72647_;
wire _72648_;
wire _72649_;
wire _72650_;
wire _72651_;
wire _72652_;
wire _72653_;
wire _72654_;
wire _72655_;
wire _72656_;
wire _72657_;
wire _72658_;
wire _72659_;
wire _72660_;
wire _72661_;
wire _72662_;
wire _72663_;
wire _72664_;
wire _72665_;
wire _72666_;
wire _72667_;
wire _72668_;
wire _72669_;
wire _72670_;
wire _72671_;
wire _72672_;
wire _72673_;
wire _72674_;
wire _72675_;
wire _72676_;
wire _72677_;
wire _72678_;
wire _72679_;
wire _72680_;
wire _72681_;
wire _72682_;
wire _72683_;
wire _72684_;
wire _72685_;
wire _72686_;
wire _72687_;
wire _72688_;
wire _72689_;
wire _72690_;
wire _72691_;
wire _72692_;
wire _72693_;
wire _72694_;
wire _72695_;
wire _72696_;
wire _72697_;
wire _72698_;
wire _72699_;
wire _72700_;
wire _72701_;
wire _72702_;
wire _72703_;
wire _72704_;
wire _72705_;
wire _72706_;
wire _72707_;
wire _72708_;
wire _72709_;
wire _72710_;
wire _72711_;
wire _72712_;
wire _72713_;
wire _72714_;
wire _72715_;
wire _72716_;
wire _72717_;
wire _72718_;
wire _72719_;
wire _72720_;
wire _72721_;
wire _72722_;
wire _72723_;
wire _72724_;
wire _72725_;
wire _72726_;
wire _72727_;
wire _72728_;
wire _72729_;
wire _72730_;
wire _72731_;
wire _72732_;
wire _72733_;
wire _72734_;
wire _72735_;
wire _72736_;
wire _72737_;
wire _72738_;
wire _72739_;
wire _72740_;
wire _72741_;
wire _72742_;
wire _72743_;
wire _72744_;
wire _72745_;
wire _72746_;
wire _72747_;
wire _72748_;
wire _72749_;
wire _72750_;
wire _72751_;
wire _72752_;
wire _72753_;
wire _72754_;
wire _72755_;
wire _72756_;
wire _72757_;
wire _72758_;
wire _72759_;
wire _72760_;
wire _72761_;
wire _72762_;
wire _72763_;
wire _72764_;
wire _72765_;
wire _72766_;
wire _72767_;
wire _72768_;
wire _72769_;
wire _72770_;
wire _72771_;
wire _72772_;
wire _72773_;
wire _72774_;
wire _72775_;
wire _72776_;
wire _72777_;
wire _72778_;
wire _72779_;
wire _72780_;
wire _72781_;
wire _72782_;
wire _72783_;
wire _72784_;
wire _72785_;
wire _72786_;
wire _72787_;
wire _72788_;
wire _72789_;
wire _72790_;
wire _72791_;
wire _72792_;
wire _72793_;
wire _72794_;
wire _72795_;
wire _72796_;
wire _72797_;
wire _72798_;
wire _72799_;
wire _72800_;
wire _72801_;
wire _72802_;
wire _72803_;
wire _72804_;
wire _72805_;
wire _72806_;
wire _72807_;
wire _72808_;
wire _72809_;
wire _72810_;
wire _72811_;
wire _72812_;
wire _72813_;
wire _72814_;
wire _72815_;
wire _72816_;
wire _72817_;
wire _72818_;
wire _72819_;
wire _72820_;
wire _72821_;
wire _72822_;
wire _72823_;
wire _72824_;
wire _72825_;
wire _72826_;
wire _72827_;
wire _72828_;
wire _72829_;
wire _72830_;
wire _72831_;
wire _72832_;
wire _72833_;
wire _72834_;
wire _72835_;
wire _72836_;
wire _72837_;
wire _72838_;
wire _72839_;
wire _72840_;
wire _72841_;
wire _72842_;
wire _72843_;
wire _72844_;
wire _72845_;
wire _72846_;
wire _72847_;
wire _72848_;
wire _72849_;
wire _72850_;
wire _72851_;
wire _72852_;
wire _72853_;
wire _72854_;
wire _72855_;
wire _72856_;
wire _72857_;
wire _72858_;
wire _72859_;
wire _72860_;
wire _72861_;
wire _72862_;
wire _72863_;
wire _72864_;
wire _72865_;
wire _72866_;
wire _72867_;
wire _72868_;
wire _72869_;
wire _72870_;
wire _72871_;
wire _72872_;
wire _72873_;
wire _72874_;
wire _72875_;
wire _72876_;
wire _72877_;
wire _72878_;
wire _72879_;
wire _72880_;
wire _72881_;
wire _72882_;
wire _72883_;
wire _72884_;
wire _72885_;
wire _72886_;
wire _72887_;
wire _72888_;
wire _72889_;
wire _72890_;
wire _72891_;
wire _72892_;
wire _72893_;
wire _72894_;
wire _72895_;
wire _72896_;
wire _72897_;
wire _72898_;
wire _72899_;
wire _72900_;
wire _72901_;
wire _72902_;
wire _72903_;
wire _72904_;
wire _72905_;
wire _72906_;
wire _72907_;
wire _72908_;
wire _72909_;
wire _72910_;
wire _72911_;
wire _72912_;
wire _72913_;
wire _72914_;
wire _72915_;
wire _72916_;
wire _72917_;
wire _72918_;
wire _72919_;
wire _72920_;
wire _72921_;
wire _72922_;
wire _72923_;
wire _72924_;
wire _72925_;
wire _72926_;
wire _72927_;
wire _72928_;
wire _72929_;
wire _72930_;
wire _72931_;
wire _72932_;
wire _72933_;
wire _72934_;
wire _72935_;
wire _72936_;
wire _72937_;
wire _72938_;
wire _72939_;
wire _72940_;
wire _72941_;
wire _72942_;
wire _72943_;
wire _72944_;
wire _72945_;
wire _72946_;
wire _72947_;
wire _72948_;
wire _72949_;
wire _72950_;
wire _72951_;
wire _72952_;
wire _72953_;
wire _72954_;
wire _72955_;
wire _72956_;
wire _72957_;
wire _72958_;
wire _72959_;
wire _72960_;
wire _72961_;
wire _72962_;
wire _72963_;
wire _72964_;
wire _72965_;
wire _72966_;
wire _72967_;
wire _72968_;
wire _72969_;
wire _72970_;
wire _72971_;
wire _72972_;
wire _72973_;
wire _72974_;
wire _72975_;
wire _72976_;
wire _72977_;
wire _72978_;
wire _72979_;
wire _72980_;
wire _72981_;
wire _72982_;
wire _72983_;
wire _72984_;
wire _72985_;
wire _72986_;
wire _72987_;
wire _72988_;
wire _72989_;
wire _72990_;
wire _72991_;
wire _72992_;
wire _72993_;
wire _72994_;
wire _72995_;
wire _72996_;
wire _72997_;
wire _72998_;
wire _72999_;
wire _73000_;
wire _73001_;
wire _73002_;
wire _73003_;
wire _73004_;
wire _73005_;
wire _73006_;
wire _73007_;
wire _73008_;
wire _73009_;
wire _73010_;
wire _73011_;
wire _73012_;
wire _73013_;
wire _73014_;
wire _73015_;
wire _73016_;
wire _73017_;
wire _73018_;
wire _73019_;
wire _73020_;
wire _73021_;
wire _73022_;
wire _73023_;
wire _73024_;
wire _73025_;
wire _73026_;
wire _73027_;
wire _73028_;
wire _73029_;
wire _73030_;
wire _73031_;
wire _73032_;
wire _73033_;
wire _73034_;
wire _73035_;
wire _73036_;
wire _73037_;
wire _73038_;
wire _73039_;
wire _73040_;
wire _73041_;
wire _73042_;
wire _73043_;
wire _73044_;
wire _73045_;
wire _73046_;
wire _73047_;
wire _73048_;
wire _73049_;
wire _73050_;
wire _73051_;
wire _73052_;
wire _73053_;
wire _73054_;
wire _73055_;
wire _73056_;
wire _73057_;
wire _73058_;
wire _73059_;
wire _73060_;
wire _73061_;
wire _73062_;
wire _73063_;
wire _73064_;
wire _73065_;
wire _73066_;
wire _73067_;
wire _73068_;
wire _73069_;
wire _73070_;
wire _73071_;
wire _73072_;
wire _73073_;
wire _73074_;
wire _73075_;
wire _73076_;
wire _73077_;
wire _73078_;
wire _73079_;
wire _73080_;
wire _73081_;
wire _73082_;
wire _73083_;
wire _73084_;
wire _73085_;
wire _73086_;
wire _73087_;
wire _73088_;
wire _73089_;
wire _73090_;
wire _73091_;
wire _73092_;
wire _73093_;
wire _73094_;
wire _73095_;
wire _73096_;
wire _73097_;
wire _73098_;
wire _73099_;
wire _73100_;
wire _73101_;
wire _73102_;
wire _73103_;
wire _73104_;
wire _73105_;
wire _73106_;
wire _73107_;
wire _73108_;
wire _73109_;
wire _73110_;
wire _73111_;
wire _73112_;
wire _73113_;
wire _73114_;
wire _73115_;
wire _73116_;
wire _73117_;
wire _73118_;
wire _73119_;
wire _73120_;
wire _73121_;
wire _73122_;
wire _73123_;
wire _73124_;
wire _73125_;
wire _73126_;
wire _73127_;
wire _73128_;
wire _73129_;
wire _73130_;
wire _73131_;
wire _73132_;
wire _73133_;
wire _73134_;
wire _73135_;
wire _73136_;
wire _73137_;
wire _73138_;
wire _73139_;
wire _73140_;
wire _73141_;
wire _73142_;
wire _73143_;
wire _73144_;
wire _73145_;
wire _73146_;
wire _73147_;
wire _73148_;
wire _73149_;
wire _73150_;
wire _73151_;
wire _73152_;
wire _73153_;
wire _73154_;
wire _73155_;
wire _73156_;
wire _73157_;
wire _73158_;
wire _73159_;
wire _73160_;
wire _73161_;
wire _73162_;
wire _73163_;
wire _73164_;
wire _73165_;
wire _73166_;
wire _73167_;
wire _73168_;
wire _73169_;
wire _73170_;
wire _73171_;
wire _73172_;
wire _73173_;
wire _73174_;
wire _73175_;
wire _73176_;
wire _73177_;
wire _73178_;
wire _73179_;
wire _73180_;
wire _73181_;
wire _73182_;
wire _73183_;
wire _73184_;
wire _73185_;
wire _73186_;
wire _73187_;
wire _73188_;
wire _73189_;
wire _73190_;
wire _73191_;
wire _73192_;
wire _73193_;
wire _73194_;
wire _73195_;
wire _73196_;
wire _73197_;
wire _73198_;
wire _73199_;
wire _73200_;
wire _73201_;
wire _73202_;
wire _73203_;
wire _73204_;
wire _73205_;
wire _73206_;
wire _73207_;
wire _73208_;
wire _73209_;
wire _73210_;
wire _73211_;
wire _73212_;
wire _73213_;
wire _73214_;
wire _73215_;
wire _73216_;
wire _73217_;
wire _73218_;
wire _73219_;
wire _73220_;
wire _73221_;
wire _73222_;
wire _73223_;
wire _73224_;
wire _73225_;
wire _73226_;
wire _73227_;
wire _73228_;
wire _73229_;
wire _73230_;
wire _73231_;
wire _73232_;
wire _73233_;
wire _73234_;
wire _73235_;
wire _73236_;
wire _73237_;
wire _73238_;
wire _73239_;
wire _73240_;
wire _73241_;
wire _73242_;
wire _73243_;
wire _73244_;
wire _73245_;
wire _73246_;
wire _73247_;
wire _73248_;
wire _73249_;
wire _73250_;
wire _73251_;
wire _73252_;
wire _73253_;
wire _73254_;
wire _73255_;
wire _73256_;
wire _73257_;
wire _73258_;
wire _73259_;
wire _73260_;
wire _73261_;
wire _73262_;
wire _73263_;
wire _73264_;
wire _73265_;
wire _73266_;
wire _73267_;
wire _73268_;
wire _73269_;
wire _73270_;
wire _73271_;
wire _73272_;
wire _73273_;
wire _73274_;
wire _73275_;
wire _73276_;
wire _73277_;
wire _73278_;
wire _73279_;
wire _73280_;
wire _73281_;
wire _73282_;
wire _73283_;
wire _73284_;
wire _73285_;
wire _73286_;
wire _73287_;
wire _73288_;
wire _73289_;
wire _73290_;
wire _73291_;
wire _73292_;
wire _73293_;
wire _73294_;
wire _73295_;
wire _73296_;
wire _73297_;
wire _73298_;
wire _73299_;
wire _73300_;
wire _73301_;
wire _73302_;
wire _73303_;
wire _73304_;
wire _73305_;
wire _73306_;
wire _73307_;
wire _73308_;
wire _73309_;
wire _73310_;
wire _73311_;
wire _73312_;
wire _73313_;
wire _73314_;
wire _73315_;
wire _73316_;
wire _73317_;
wire _73318_;
wire _73319_;
wire _73320_;
wire _73321_;
wire _73322_;
wire _73323_;
wire _73324_;
wire _73325_;
wire _73326_;
wire _73327_;
wire _73328_;
wire _73329_;
wire _73330_;
wire _73331_;
wire _73332_;
wire _73333_;
wire _73334_;
wire _73335_;
wire _73336_;
wire _73337_;
wire _73338_;
wire _73339_;
wire _73340_;
wire _73341_;
wire _73342_;
wire _73343_;
wire _73344_;
wire _73345_;
wire _73346_;
wire _73347_;
wire _73348_;
wire _73349_;
wire _73350_;
wire _73351_;
wire _73352_;
wire _73353_;
wire _73354_;
wire _73355_;
wire _73356_;
wire _73357_;
wire _73358_;
wire _73359_;
wire _73360_;
wire _73361_;
wire _73362_;
wire _73363_;
wire _73364_;
wire _73365_;
wire _73366_;
wire _73367_;
wire _73368_;
wire _73369_;
wire _73370_;
wire _73371_;
wire _73372_;
wire _73373_;
wire _73374_;
wire _73375_;
wire _73376_;
wire _73377_;
wire _73378_;
wire _73379_;
wire _73380_;
wire _73381_;
wire _73382_;
wire _73383_;
wire _73384_;
wire _73385_;
wire _73386_;
wire _73387_;
wire _73388_;
wire _73389_;
wire _73390_;
wire _73391_;
wire _73392_;
wire _73393_;
wire _73394_;
wire _73395_;
wire _73396_;
wire _73397_;
wire _73398_;
wire _73399_;
wire _73400_;
wire _73401_;
wire _73402_;
wire _73403_;
wire _73404_;
wire _73405_;
wire _73406_;
wire _73407_;
wire _73408_;
wire _73409_;
wire _73410_;
wire _73411_;
wire _73412_;
wire _73413_;
wire _73414_;
wire _73415_;
wire _73416_;
wire _73417_;
wire _73418_;
wire _73419_;
wire _73420_;
wire _73421_;
wire _73422_;
wire _73423_;
wire _73424_;
wire _73425_;
wire _73426_;
wire _73427_;
wire _73428_;
wire _73429_;
wire _73430_;
wire _73431_;
wire _73432_;
wire _73433_;
wire _73434_;
wire _73435_;
wire _73436_;
wire _73437_;
wire _73438_;
wire _73439_;
wire _73440_;
wire _73441_;
wire _73442_;
wire _73443_;
wire _73444_;
wire _73445_;
wire _73446_;
wire _73447_;
wire _73448_;
wire _73449_;
wire _73450_;
wire _73451_;
wire _73452_;
wire _73453_;
wire _73454_;
wire _73455_;
wire _73456_;
wire _73457_;
wire _73458_;
wire _73459_;
wire _73460_;
wire _73461_;
wire _73462_;
wire _73463_;
wire _73464_;
wire _73465_;
wire _73466_;
wire _73467_;
wire _73468_;
wire _73469_;
wire _73470_;
wire _73471_;
wire _73472_;
wire _73473_;
wire _73474_;
wire _73475_;
wire _73476_;
wire _73477_;
wire _73478_;
wire _73479_;
wire _73480_;
wire _73481_;
wire _73482_;
wire _73483_;
wire _73484_;
wire _73485_;
wire _73486_;
wire _73487_;
wire _73488_;
wire _73489_;
wire _73490_;
wire _73491_;
wire _73492_;
wire _73493_;
wire _73494_;
wire _73495_;
wire _73496_;
wire _73497_;
wire _73498_;
wire _73499_;
wire _73500_;
wire _73501_;
wire _73502_;
wire _73503_;
wire _73504_;
wire _73505_;
wire _73506_;
wire _73507_;
wire _73508_;
wire _73509_;
wire _73510_;
wire _73511_;
wire _73512_;
wire _73513_;
wire _73514_;
wire _73515_;
wire _73516_;
wire _73517_;
wire _73518_;
wire _73519_;
wire _73520_;
wire _73521_;
wire _73522_;
wire _73523_;
wire _73524_;
wire _73525_;
wire _73526_;
wire _73527_;
wire _73528_;
wire _73529_;
wire _73530_;
wire _73531_;
wire _73532_;
wire _73533_;
wire _73534_;
wire _73535_;
wire _73536_;
wire _73537_;
wire _73538_;
wire _73539_;
wire _73540_;
wire _73541_;
wire _73542_;
wire _73543_;
wire _73544_;
wire _73545_;
wire _73546_;
wire _73547_;
wire _73548_;
wire _73549_;
wire _73550_;
wire _73551_;
wire _73552_;
wire _73553_;
wire _73554_;
wire _73555_;
wire _73556_;
wire _73557_;
wire _73558_;
wire _73559_;
wire _73560_;
wire _73561_;
wire _73562_;
wire _73563_;
wire _73564_;
wire _73565_;
wire _73566_;
wire _73567_;
wire _73568_;
wire _73569_;
wire _73570_;
wire _73571_;
wire _73572_;
wire _73573_;
wire _73574_;
wire _73575_;
wire _73576_;
wire _73577_;
wire _73578_;
wire _73579_;
wire _73580_;
wire _73581_;
wire _73582_;
wire _73583_;
wire _73584_;
wire _73585_;
wire _73586_;
wire _73587_;
wire _73588_;
wire _73589_;
wire _73590_;
wire _73591_;
wire _73592_;
wire _73593_;
wire _73594_;
wire _73595_;
wire _73596_;
wire _73597_;
wire _73598_;
wire _73599_;
wire _73600_;
wire _73601_;
wire _73602_;
wire _73603_;
wire _73604_;
wire _73605_;
wire _73606_;
wire _73607_;
wire _73608_;
wire _73609_;
wire _73610_;
wire _73611_;
wire _73612_;
wire _73613_;
wire _73614_;
wire _73615_;
wire _73616_;
wire _73617_;
wire _73618_;
wire _73619_;
wire _73620_;
wire _73621_;
wire _73622_;
wire _73623_;
wire _73624_;
wire _73625_;
wire _73626_;
wire _73627_;
wire _73628_;
wire _73629_;
wire _73630_;
wire _73631_;
wire _73632_;
wire _73633_;
wire _73634_;
wire _73635_;
wire _73636_;
wire _73637_;
wire _73638_;
wire _73639_;
wire _73640_;
wire _73641_;
wire _73642_;
wire _73643_;
wire _73644_;
wire _73645_;
wire _73646_;
wire _73647_;
wire _73648_;
wire _73649_;
wire _73650_;
wire _73651_;
wire _73652_;
wire _73653_;
wire _73654_;
wire _73655_;
wire _73656_;
wire _73657_;
wire _73658_;
wire _73659_;
wire _73660_;
wire _73661_;
wire _73662_;
wire _73663_;
wire _73664_;
wire _73665_;
wire _73666_;
wire _73667_;
wire _73668_;
wire _73669_;
wire _73670_;
wire _73671_;
wire _73672_;
wire _73673_;
wire _73674_;
wire _73675_;
wire _73676_;
wire _73677_;
wire _73678_;
wire _73679_;
wire _73680_;
wire _73681_;
wire _73682_;
wire _73683_;
wire _73684_;
wire _73685_;
wire _73686_;
wire _73687_;
wire _73688_;
wire _73689_;
wire _73690_;
wire _73691_;
wire _73692_;
wire _73693_;
wire _73694_;
wire _73695_;
wire _73696_;
wire _73697_;
wire _73698_;
wire _73699_;
wire _73700_;
wire _73701_;
wire _73702_;
wire _73703_;
wire _73704_;
wire _73705_;
wire _73706_;
wire _73707_;
wire _73708_;
wire _73709_;
wire _73710_;
wire _73711_;
wire _73712_;
wire _73713_;
wire _73714_;
wire _73715_;
wire _73716_;
wire _73717_;
wire _73718_;
wire _73719_;
wire _73720_;
wire _73721_;
wire _73722_;
wire _73723_;
wire _73724_;
wire _73725_;
wire _73726_;
wire _73727_;
wire _73728_;
wire _73729_;
wire _73730_;
wire _73731_;
wire _73732_;
wire _73733_;
wire _73734_;
wire _73735_;
wire _73736_;
wire _73737_;
wire _73738_;
wire _73739_;
wire _73740_;
wire _73741_;
wire _73742_;
wire _73743_;
wire _73744_;
wire _73745_;
wire _73746_;
wire _73747_;
wire _73748_;
wire _73749_;
wire _73750_;
wire _73751_;
wire _73752_;
wire _73753_;
wire _73754_;
wire _73755_;
wire _73756_;
wire _73757_;
wire _73758_;
wire _73759_;
wire _73760_;
wire _73761_;
wire _73762_;
wire _73763_;
wire _73764_;
wire _73765_;
wire _73766_;
wire _73767_;
wire _73768_;
wire _73769_;
wire _73770_;
wire _73771_;
wire _73772_;
wire _73773_;
wire _73774_;
wire _73775_;
wire _73776_;
wire _73777_;
wire _73778_;
wire _73779_;
wire _73780_;
wire _73781_;
wire _73782_;
wire _73783_;
wire _73784_;
wire _73785_;
wire _73786_;
wire _73787_;
wire _73788_;
wire _73789_;
wire _73790_;
wire _73791_;
wire _73792_;
wire _73793_;
wire _73794_;
wire _73795_;
wire _73796_;
wire _73797_;
wire _73798_;
wire _73799_;
wire _73800_;
wire _73801_;
wire _73802_;
wire _73803_;
wire _73804_;
wire _73805_;
wire _73806_;
wire _73807_;
wire _73808_;
wire _73809_;
wire _73810_;
wire _73811_;
wire _73812_;
wire _73813_;
wire _73814_;
wire _73815_;
wire _73816_;
wire _73817_;
wire _73818_;
wire _73819_;
wire _73820_;
wire _73821_;
wire _73822_;
wire _73823_;
wire _73824_;
wire _73825_;
wire _73826_;
wire _73827_;
wire _73828_;
wire _73829_;
wire _73830_;
wire _73831_;
wire _73832_;
wire _73833_;
wire _73834_;
wire _73835_;
wire _73836_;
wire _73837_;
wire _73838_;
wire _73839_;
wire _73840_;
wire _73841_;
wire _73842_;
wire _73843_;
wire _73844_;
wire _73845_;
wire _73846_;
wire _73847_;
wire _73848_;
wire _73849_;
wire _73850_;
wire _73851_;
wire _73852_;
wire _73853_;
wire _73854_;
wire _73855_;
wire _73856_;
wire _73857_;
wire _73858_;
wire _73859_;
wire _73860_;
wire _73861_;
wire _73862_;
wire _73863_;
wire _73864_;
wire _73865_;
wire _73866_;
wire _73867_;
wire _73868_;
wire _73869_;
wire _73870_;
wire _73871_;
wire _73872_;
wire _73873_;
wire _73874_;
wire _73875_;
wire _73876_;
wire _73877_;
wire _73878_;
wire _73879_;
wire _73880_;
wire _73881_;
wire _73882_;
wire _73883_;
wire _73884_;
wire _73885_;
wire _73886_;
wire _73887_;
wire _73888_;
wire _73889_;
wire _73890_;
wire _73891_;
wire _73892_;
wire _73893_;
wire _73894_;
wire _73895_;
wire _73896_;
wire _73897_;
wire _73898_;
wire _73899_;
wire _73900_;
wire _73901_;
wire _73902_;
wire _73903_;
wire _73904_;
wire _73905_;
wire _73906_;
wire _73907_;
wire _73908_;
wire _73909_;
wire _73910_;
wire _73911_;
wire _73912_;
wire _73913_;
wire _73914_;
wire _73915_;
wire _73916_;
wire _73917_;
wire _73918_;
wire _73919_;
wire _73920_;
wire _73921_;
wire _73922_;
wire _73923_;
wire _73924_;
wire _73925_;
wire _73926_;
wire _73927_;
wire _73928_;
wire _73929_;
wire _73930_;
wire _73931_;
wire _73932_;
wire _73933_;
wire _73934_;
wire _73935_;
wire _73936_;
wire _73937_;
wire _73938_;
wire _73939_;
wire _73940_;
wire _73941_;
wire _73942_;
wire _73943_;
wire _73944_;
wire _73945_;
wire _73946_;
wire _73947_;
wire _73948_;
wire _73949_;
wire _73950_;
wire _73951_;
wire _73952_;
wire _73953_;
wire _73954_;
wire _73955_;
wire _73956_;
wire _73957_;
wire _73958_;
wire _73959_;
wire _73960_;
wire _73961_;
wire _73962_;
wire _73963_;
wire _73964_;
wire _73965_;
wire _73966_;
wire _73967_;
wire _73968_;
wire _73969_;
wire _73970_;
wire _73971_;
wire _73972_;
wire _73973_;
wire _73974_;
wire _73975_;
wire _73976_;
wire _73977_;
wire _73978_;
wire _73979_;
wire _73980_;
wire _73981_;
wire _73982_;
wire _73983_;
wire _73984_;
wire _73985_;
wire _73986_;
wire _73987_;
wire _73988_;
wire _73989_;
wire _73990_;
wire _73991_;
wire _73992_;
wire _73993_;
wire _73994_;
wire _73995_;
wire _73996_;
wire _73997_;
wire _73998_;
wire _73999_;
wire _74000_;
wire _74001_;
wire _74002_;
wire _74003_;
wire _74004_;
wire _74005_;
wire _74006_;
wire _74007_;
wire _74008_;
wire _74009_;
wire _74010_;
wire _74011_;
wire _74012_;
wire _74013_;
wire _74014_;
wire _74015_;
wire _74016_;
wire _74017_;
wire _74018_;
wire _74019_;
wire _74020_;
wire _74021_;
wire _74022_;
wire _74023_;
wire _74024_;
wire _74025_;
wire _74026_;
wire _74027_;
wire _74028_;
wire _74029_;
wire _74030_;
wire _74031_;
wire _74032_;
wire _74033_;
wire _74034_;
wire _74035_;
wire _74036_;
wire _74037_;
wire _74038_;
wire _74039_;
wire _74040_;
wire _74041_;
wire _74042_;
wire _74043_;
wire _74044_;
wire _74045_;
wire _74046_;
wire _74047_;
wire _74048_;
wire _74049_;
wire _74050_;
wire _74051_;
wire _74052_;
wire _74053_;
wire _74054_;
wire _74055_;
wire _74056_;
wire _74057_;
wire _74058_;
wire _74059_;
wire _74060_;
wire _74061_;
wire _74062_;
wire _74063_;
wire _74064_;
wire _74065_;
wire _74066_;
wire _74067_;
wire _74068_;
wire _74069_;
wire _74070_;
wire _74071_;
wire _74072_;
wire _74073_;
wire _74074_;
wire _74075_;
wire _74076_;
wire _74077_;
wire _74078_;
wire _74079_;
wire _74080_;
wire _74081_;
wire _74082_;
wire _74083_;
wire _74084_;
wire _74085_;
wire _74086_;
wire _74087_;
wire _74088_;
wire _74089_;
wire _74090_;
wire _74091_;
wire _74092_;
wire _74093_;
wire _74094_;
wire _74095_;
wire _74096_;
wire _74097_;
wire _74098_;
wire _74099_;
wire _74100_;
wire _74101_;
wire _74102_;
wire _74103_;
wire _74104_;
wire _74105_;
wire _74106_;
wire _74107_;
wire _74108_;
wire _74109_;
wire _74110_;
wire _74111_;
wire _74112_;
wire _74113_;
wire _74114_;
wire _74115_;
wire _74116_;
wire _74117_;
wire _74118_;
wire _74119_;
wire _74120_;
wire _74121_;
wire _74122_;
wire _74123_;
wire _74124_;
wire _74125_;
wire _74126_;
wire _74127_;
wire _74128_;
wire _74129_;
wire _74130_;
wire _74131_;
wire _74132_;
wire _74133_;
wire _74134_;
wire _74135_;
wire _74136_;
wire _74137_;
wire _74138_;
wire _74139_;
wire _74140_;
wire _74141_;
wire _74142_;
wire _74143_;
wire _74144_;
wire _74145_;
wire _74146_;
wire _74147_;
wire _74148_;
wire _74149_;
wire _74150_;
wire _74151_;
wire _74152_;
wire _74153_;
wire _74154_;
wire _74155_;
wire _74156_;
wire _74157_;
wire _74158_;
wire _74159_;
wire _74160_;
wire _74161_;
wire _74162_;
wire _74163_;
wire _74164_;
wire _74165_;
wire _74166_;
wire _74167_;
wire _74168_;
wire _74169_;
wire _74170_;
wire _74171_;
wire _74172_;
wire _74173_;
wire _74174_;
wire _74175_;
wire _74176_;
wire _74177_;
wire _74178_;
wire _74179_;
wire _74180_;
wire _74181_;
wire _74182_;
wire _74183_;
wire _74184_;
wire _74185_;
wire _74186_;
wire _74187_;
wire _74188_;
wire _74189_;
wire _74190_;
wire _74191_;
wire _74192_;
wire _74193_;
wire _74194_;
wire _74195_;
wire _74196_;
wire _74197_;
wire _74198_;
wire _74199_;
wire _74200_;
wire _74201_;
wire _74202_;
wire _74203_;
wire _74204_;
wire _74205_;
wire _74206_;
wire _74207_;
wire _74208_;
wire _74209_;
wire _74210_;
wire _74211_;
wire _74212_;
wire _74213_;
wire _74214_;
wire _74215_;
wire _74216_;
wire _74217_;
wire _74218_;
wire _74219_;
wire _74220_;
wire _74221_;
wire _74222_;
wire _74223_;
wire _74224_;
wire _74225_;
wire _74226_;
wire _74227_;
wire _74228_;
wire _74229_;
wire _74230_;
wire _74231_;
wire _74232_;
wire _74233_;
wire _74234_;
wire _74235_;
wire _74236_;
wire _74237_;
wire _74238_;
wire _74239_;
wire _74240_;
wire _74241_;
wire _74242_;
wire _74243_;
wire _74244_;
wire _74245_;
wire _74246_;
wire _74247_;
wire _74248_;
wire _74249_;
wire _74250_;
wire _74251_;
wire _74252_;
wire _74253_;
wire _74254_;
wire _74255_;
wire _74256_;
wire _74257_;
wire _74258_;
wire _74259_;
wire _74260_;
wire _74261_;
wire _74262_;
wire _74263_;
wire _74264_;
wire _74265_;
wire _74266_;
wire _74267_;
wire _74268_;
wire _74269_;
wire _74270_;
wire _74271_;
wire _74272_;
wire _74273_;
wire _74274_;
wire _74275_;
wire _74276_;
wire _74277_;
wire _74278_;
wire _74279_;
wire _74280_;
wire _74281_;
wire _74282_;
wire _74283_;
wire _74284_;
wire _74285_;
wire _74286_;
wire _74287_;
wire _74288_;
wire _74289_;
wire _74290_;
wire _74291_;
wire _74292_;
wire _74293_;
wire _74294_;
wire _74295_;
wire _74296_;
wire _74297_;
wire _74298_;
wire _74299_;
wire _74300_;
wire _74301_;
wire _74302_;
wire _74303_;
wire _74304_;
wire _74305_;
wire _74306_;
wire _74307_;
wire _74308_;
wire _74309_;
wire _74310_;
wire _74311_;
wire _74312_;
wire _74313_;
wire _74314_;
wire _74315_;
wire _74316_;
wire _74317_;
wire _74318_;
wire _74319_;
wire _74320_;
wire _74321_;
wire _74322_;
wire _74323_;
wire _74324_;
wire _74325_;
wire _74326_;
wire _74327_;
wire _74328_;
wire _74329_;
wire _74330_;
wire _74331_;
wire _74332_;
wire _74333_;
wire _74334_;
wire _74335_;
wire _74336_;
wire _74337_;
wire _74338_;
wire _74339_;
wire _74340_;
wire _74341_;
wire _74342_;
wire _74343_;
wire _74344_;
wire _74345_;
wire _74346_;
wire _74347_;
wire _74348_;
wire _74349_;
wire _74350_;
wire _74351_;
wire _74352_;
wire _74353_;
wire _74354_;
wire _74355_;
wire _74356_;
wire _74357_;
wire _74358_;
wire _74359_;
wire _74360_;
wire _74361_;
wire _74362_;
wire _74363_;
wire _74364_;
wire _74365_;
wire _74366_;
wire _74367_;
wire _74368_;
wire _74369_;
wire _74370_;
wire _74371_;
wire _74372_;
wire _74373_;
wire _74374_;
wire _74375_;
wire _74376_;
wire _74377_;
wire _74378_;
wire _74379_;
wire _74380_;
wire _74381_;
wire _74382_;
wire _74383_;
wire _74384_;
wire _74385_;
wire _74386_;
wire _74387_;
wire _74388_;
wire _74389_;
wire _74390_;
wire _74391_;
wire _74392_;
wire _74393_;
wire _74394_;
wire _74395_;
wire _74396_;
wire _74397_;
wire _74398_;
wire _74399_;
wire _74400_;
wire _74401_;
wire _74402_;
wire _74403_;
wire _74404_;
wire _74405_;
wire _74406_;
wire _74407_;
wire _74408_;
wire _74409_;
wire _74410_;
wire _74411_;
wire _74412_;
wire _74413_;
wire _74414_;
wire _74415_;
wire _74416_;
wire _74417_;
wire _74418_;
wire _74419_;
wire _74420_;
wire _74421_;
wire _74422_;
wire _74423_;
wire _74424_;
wire _74425_;
wire _74426_;
wire _74427_;
wire _74428_;
wire _74429_;
wire _74430_;
wire _74431_;
wire _74432_;
wire _74433_;
wire _74434_;
wire _74435_;
wire _74436_;
wire _74437_;
wire _74438_;
wire _74439_;
wire _74440_;
wire _74441_;
wire _74442_;
wire _74443_;
wire _74444_;
wire _74445_;
wire _74446_;
wire _74447_;
wire _74448_;
wire _74449_;
wire _74450_;
wire _74451_;
wire _74452_;
wire _74453_;
wire _74454_;
wire _74455_;
wire _74456_;
wire _74457_;
wire _74458_;
wire _74459_;
wire _74460_;
wire _74461_;
wire _74462_;
wire _74463_;
wire _74464_;
wire _74465_;
wire _74466_;
wire _74467_;
wire _74468_;
wire _74469_;
wire _74470_;
wire _74471_;
wire _74472_;
wire _74473_;
wire _74474_;
wire _74475_;
wire _74476_;
wire _74477_;
wire _74478_;
wire _74479_;
wire _74480_;
wire _74481_;
wire _74482_;
wire _74483_;
wire _74484_;
wire _74485_;
wire _74486_;
wire _74487_;
wire _74488_;
wire _74489_;
wire _74490_;
wire _74491_;
wire _74492_;
wire _74493_;
wire _74494_;
wire _74495_;
wire _74496_;
wire _74497_;
wire _74498_;
wire _74499_;
wire _74500_;
wire _74501_;
wire _74502_;
wire _74503_;
wire _74504_;
wire _74505_;
wire _74506_;
wire _74507_;
wire _74508_;
wire _74509_;
wire _74510_;
wire _74511_;
wire _74512_;
wire _74513_;
wire _74514_;
wire _74515_;
wire _74516_;
wire _74517_;
wire _74518_;
wire _74519_;
wire _74520_;
wire _74521_;
wire _74522_;
wire _74523_;
wire _74524_;
wire _74525_;
wire _74526_;
wire _74527_;
wire _74528_;
wire _74529_;
wire _74530_;
wire _74531_;
wire _74532_;
wire _74533_;
wire _74534_;
wire _74535_;
wire _74536_;
wire _74537_;
wire _74538_;
wire _74539_;
wire _74540_;
wire _74541_;
wire _74542_;
wire _74543_;
wire _74544_;
wire _74545_;
wire _74546_;
wire _74547_;
wire _74548_;
wire _74549_;
wire _74550_;
wire _74551_;
wire _74552_;
wire _74553_;
wire _74554_;
wire _74555_;
wire _74556_;
wire _74557_;
wire _74558_;
wire _74559_;
wire _74560_;
wire _74561_;
wire _74562_;
wire _74563_;
wire _74564_;
wire _74565_;
wire _74566_;
wire _74567_;
wire _74568_;
wire _74569_;
wire _74570_;
wire _74571_;
wire _74572_;
wire _74573_;
wire _74574_;
wire _74575_;
wire _74576_;
wire _74577_;
wire _74578_;
wire _74579_;
wire _74580_;
wire _74581_;
wire _74582_;
wire _74583_;
wire _74584_;
wire _74585_;
wire _74586_;
wire _74587_;
wire _74588_;
wire _74589_;
wire _74590_;
wire _74591_;
wire _74592_;
wire _74593_;
wire _74594_;
wire _74595_;
wire _74596_;
wire _74597_;
wire _74598_;
wire _74599_;
wire _74600_;
wire _74601_;
wire _74602_;
wire _74603_;
wire _74604_;
wire _74605_;
wire _74606_;
wire _74607_;
wire _74608_;
wire _74609_;
wire _74610_;
wire _74611_;
wire _74612_;
wire _74613_;
wire _74614_;
wire _74615_;
wire _74616_;
wire _74617_;
wire _74618_;
wire _74619_;
wire _74620_;
wire _74621_;
wire _74622_;
wire _74623_;
wire _74624_;
wire _74625_;
wire _74626_;
wire _74627_;
wire _74628_;
wire _74629_;
wire _74630_;
wire _74631_;
wire _74632_;
wire _74633_;
wire _74634_;
wire _74635_;
wire _74636_;
wire _74637_;
wire _74638_;
wire _74639_;
wire _74640_;
wire _74641_;
wire _74642_;
wire _74643_;
wire _74644_;
wire _74645_;
wire _74646_;
wire _74647_;
wire _74648_;
wire _74649_;
wire _74650_;
wire _74651_;
wire _74652_;
wire _74653_;
wire _74654_;
wire _74655_;
wire _74656_;
wire _74657_;
wire _74658_;
wire _74659_;
wire _74660_;
wire _74661_;
wire _74662_;
wire _74663_;
wire _74664_;
wire _74665_;
wire _74666_;
wire _74667_;
wire _74668_;
wire _74669_;
wire _74670_;
wire _74671_;
wire _74672_;
wire _74673_;
wire _74674_;
wire _74675_;
wire _74676_;
wire _74677_;
wire _74678_;
wire _74679_;
wire _74680_;
wire _74681_;
wire _74682_;
wire _74683_;
wire _74684_;
wire _74685_;
wire _74686_;
wire _74687_;
wire _74688_;
wire _74689_;
wire _74690_;
wire _74691_;
wire _74692_;
wire _74693_;
wire _74694_;
wire _74695_;
wire _74696_;
wire _74697_;
wire _74698_;
wire _74699_;
wire _74700_;
wire _74701_;
wire _74702_;
wire _74703_;
wire _74704_;
wire _74705_;
wire _74706_;
wire _74707_;
wire _74708_;
wire _74709_;
wire _74710_;
wire _74711_;
wire _74712_;
wire _74713_;
wire _74714_;
wire _74715_;
wire _74716_;
wire _74717_;
wire _74718_;
wire _74719_;
wire _74720_;
wire _74721_;
wire _74722_;
wire _74723_;
wire _74724_;
wire _74725_;
wire _74726_;
wire _74727_;
wire _74728_;
wire _74729_;
wire _74730_;
wire _74731_;
wire _74732_;
wire _74733_;
wire _74734_;
wire _74735_;
wire _74736_;
wire _74737_;
wire _74738_;
wire _74739_;
wire _74740_;
wire _74741_;
wire _74742_;
wire _74743_;
wire _74744_;
wire _74745_;
wire _74746_;
wire _74747_;
wire _74748_;
wire _74749_;
wire _74750_;
wire _74751_;
wire _74752_;
wire _74753_;
wire _74754_;
wire _74755_;
wire _74756_;
wire _74757_;
wire _74758_;
wire _74759_;
wire _74760_;
wire _74761_;
wire _74762_;
wire _74763_;
wire _74764_;
wire _74765_;
wire _74766_;
wire _74767_;
wire _74768_;
wire _74769_;
wire _74770_;
wire _74771_;
wire _74772_;
wire _74773_;
wire _74774_;
wire _74775_;
wire _74776_;
wire _74777_;
wire _74778_;
wire _74779_;
wire _74780_;
wire _74781_;
wire _74782_;
wire _74783_;
wire _74784_;
wire _74785_;
wire _74786_;
wire _74787_;
wire _74788_;
wire _74789_;
wire _74790_;
wire _74791_;
wire _74792_;
wire _74793_;
wire _74794_;
wire _74795_;
wire _74796_;
wire _74797_;
wire _74798_;
wire _74799_;
wire _74800_;
wire _74801_;
wire _74802_;
wire _74803_;
wire _74804_;
wire _74805_;
wire _74806_;
wire _74807_;
wire _74808_;
wire _74809_;
wire _74810_;
wire _74811_;
wire _74812_;
wire _74813_;
wire _74814_;
wire _74815_;
wire _74816_;
wire _74817_;
wire _74818_;
wire _74819_;
wire _74820_;
wire _74821_;
wire _74822_;
wire _74823_;
wire _74824_;
wire _74825_;
wire _74826_;
wire _74827_;
wire _74828_;
wire _74829_;
wire _74830_;
wire _74831_;
wire _74832_;
wire _74833_;
wire _74834_;
wire _74835_;
wire _74836_;
wire _74837_;
wire _74838_;
wire _74839_;
wire _74840_;
wire _74841_;
wire _74842_;
wire _74843_;
wire _74844_;
wire _74845_;
wire _74846_;
wire _74847_;
wire _74848_;
wire _74849_;
wire _74850_;
wire _74851_;
wire _74852_;
wire _74853_;
wire _74854_;
wire _74855_;
wire _74856_;
wire _74857_;
wire _74858_;
wire _74859_;
wire _74860_;
wire _74861_;
wire _74862_;
wire _74863_;
wire _74864_;
wire _74865_;
wire _74866_;
wire _74867_;
wire _74868_;
wire _74869_;
wire _74870_;
wire _74871_;
wire _74872_;
wire _74873_;
wire _74874_;
wire _74875_;
wire _74876_;
wire _74877_;
wire _74878_;
wire _74879_;
wire _74880_;
wire _74881_;
wire _74882_;
wire _74883_;
wire _74884_;
wire _74885_;
wire _74886_;
wire _74887_;
wire _74888_;
wire _74889_;
wire _74890_;
wire _74891_;
wire _74892_;
wire _74893_;
wire _74894_;
wire _74895_;
wire _74896_;
wire _74897_;
wire _74898_;
wire _74899_;
wire _74900_;
wire _74901_;
wire _74902_;
wire _74903_;
wire _74904_;
wire _74905_;
wire _74906_;
wire _74907_;
wire _74908_;
wire _74909_;
wire _74910_;
wire _74911_;
wire _74912_;
wire _74913_;
wire _74914_;
wire _74915_;
wire _74916_;
wire _74917_;
wire _74918_;
wire _74919_;
wire _74920_;
wire _74921_;
wire _74922_;
wire _74923_;
wire _74924_;
wire _74925_;
wire _74926_;
wire _74927_;
wire _74928_;
wire _74929_;
wire _74930_;
wire _74931_;
wire _74932_;
wire _74933_;
wire _74934_;
wire _74935_;
wire _74936_;
wire _74937_;
wire _74938_;
wire _74939_;
wire _74940_;
wire _74941_;
wire _74942_;
wire _74943_;
wire _74944_;
wire _74945_;
wire _74946_;
wire _74947_;
wire _74948_;
wire _74949_;
wire _74950_;
wire _74951_;
wire _74952_;
wire _74953_;
wire _74954_;
wire _74955_;
wire _74956_;
wire _74957_;
wire _74958_;
wire _74959_;
wire _74960_;
wire _74961_;
wire _74962_;
wire _74963_;
wire _74964_;
wire _74965_;
wire _74966_;
wire _74967_;
wire _74968_;
wire _74969_;
wire _74970_;
wire _74971_;
wire _74972_;
wire _74973_;
wire _74974_;
wire _74975_;
wire _74976_;
wire _74977_;
wire _74978_;
wire _74979_;
wire _74980_;
wire _74981_;
wire _74982_;
wire _74983_;
wire _74984_;
wire _74985_;
wire _74986_;
wire _74987_;
wire _74988_;
wire _74989_;
wire _74990_;
wire _74991_;
wire _74992_;
wire _74993_;
wire _74994_;
wire _74995_;
wire _74996_;
wire _74997_;
wire _74998_;
wire _74999_;
wire _75000_;
wire _75001_;
wire _75002_;
wire _75003_;
wire _75004_;
wire _75005_;
wire _75006_;
wire _75007_;
wire _75008_;
wire _75009_;
wire _75010_;
wire _75011_;
wire _75012_;
wire _75013_;
wire _75014_;
wire _75015_;
wire _75016_;
wire _75017_;
wire _75018_;
wire _75019_;
wire _75020_;
wire _75021_;
wire _75022_;
wire _75023_;
wire _75024_;
wire _75025_;
wire _75026_;
wire _75027_;
wire _75028_;
wire _75029_;
wire _75030_;
wire _75031_;
wire _75032_;
wire _75033_;
wire _75034_;
wire _75035_;
wire _75036_;
wire _75037_;
wire _75038_;
wire _75039_;
wire _75040_;
wire _75041_;
wire _75042_;
wire _75043_;
wire _75044_;
wire _75045_;
wire _75046_;
wire _75047_;
wire _75048_;
wire _75049_;
wire _75050_;
wire _75051_;
wire _75052_;
wire _75053_;
wire _75054_;
wire _75055_;
wire _75056_;
wire _75057_;
wire _75058_;
wire _75059_;
wire _75060_;
wire _75061_;
wire _75062_;
wire _75063_;
wire _75064_;
wire _75065_;
wire _75066_;
wire _75067_;
wire _75068_;
wire _75069_;
wire _75070_;
wire _75071_;
wire _75072_;
wire _75073_;
wire _75074_;
wire _75075_;
wire _75076_;
wire _75077_;
wire _75078_;
wire _75079_;
wire _75080_;
wire _75081_;
wire _75082_;
wire _75083_;
wire _75084_;
wire _75085_;
wire _75086_;
wire _75087_;
wire _75088_;
wire _75089_;
wire _75090_;
wire _75091_;
wire _75092_;
wire _75093_;
wire _75094_;
wire _75095_;
wire _75096_;
wire _75097_;
wire _75098_;
wire _75099_;
wire _75100_;
wire _75101_;
wire _75102_;
wire _75103_;
wire _75104_;
wire _75105_;
wire _75106_;
wire _75107_;
wire _75108_;
wire _75109_;
wire _75110_;
wire _75111_;
wire _75112_;
wire _75113_;
wire _75114_;
wire _75115_;
wire _75116_;
wire _75117_;
wire _75118_;
wire _75119_;
wire _75120_;
wire _75121_;
wire _75122_;
wire _75123_;
wire _75124_;
wire _75125_;
wire _75126_;
wire _75127_;
wire _75128_;
wire _75129_;
wire _75130_;
wire _75131_;
wire _75132_;
wire _75133_;
wire _75134_;
wire _75135_;
wire _75136_;
wire _75137_;
wire _75138_;
wire _75139_;
wire _75140_;
wire _75141_;
wire _75142_;
wire _75143_;
wire _75144_;
wire _75145_;
wire _75146_;
wire _75147_;
wire _75148_;
wire _75149_;
wire _75150_;
wire _75151_;
wire _75152_;
wire _75153_;
wire _75154_;
wire _75155_;
wire _75156_;
wire _75157_;
wire _75158_;
wire _75159_;
wire _75160_;
wire _75161_;
wire _75162_;
wire _75163_;
wire _75164_;
wire _75165_;
wire _75166_;
wire _75167_;
wire _75168_;
wire _75169_;
wire _75170_;
wire _75171_;
wire _75172_;
wire _75173_;
wire _75174_;
wire _75175_;
wire _75176_;
wire _75177_;
wire _75178_;
wire _75179_;
wire _75180_;
wire _75181_;
wire _75182_;
wire _75183_;
wire _75184_;
wire _75185_;
wire _75186_;
wire _75187_;
wire _75188_;
wire _75189_;
wire _75190_;
wire _75191_;
wire _75192_;
wire _75193_;
wire _75194_;
wire _75195_;
wire _75196_;
wire _75197_;
wire _75198_;
wire _75199_;
wire _75200_;
wire _75201_;
wire _75202_;
wire _75203_;
wire _75204_;
wire _75205_;
wire _75206_;
wire _75207_;
wire _75208_;
wire _75209_;
wire _75210_;
wire _75211_;
wire _75212_;
wire _75213_;
wire _75214_;
wire _75215_;
wire _75216_;
wire _75217_;
wire _75218_;
wire _75219_;
wire _75220_;
wire _75221_;
wire _75222_;
wire _75223_;
wire _75224_;
wire _75225_;
wire _75226_;
wire _75227_;
wire _75228_;
wire _75229_;
wire _75230_;
wire _75231_;
wire _75232_;
wire _75233_;
wire _75234_;
wire _75235_;
wire _75236_;
wire _75237_;
wire _75238_;
wire _75239_;
wire _75240_;
wire _75241_;
wire _75242_;
wire _75243_;
wire _75244_;
wire _75245_;
wire _75246_;
wire _75247_;
wire _75248_;
wire _75249_;
wire _75250_;
wire _75251_;
wire _75252_;
wire _75253_;
wire _75254_;
wire _75255_;
wire _75256_;
wire _75257_;
wire _75258_;
wire _75259_;
wire _75260_;
wire _75261_;
wire _75262_;
wire _75263_;
wire _75264_;
wire _75265_;
wire _75266_;
wire _75267_;
wire _75268_;
wire _75269_;
wire _75270_;
wire _75271_;
wire _75272_;
wire _75273_;
wire _75274_;
wire _75275_;
wire _75276_;
wire _75277_;
wire _75278_;
wire _75279_;
wire _75280_;
wire _75281_;
wire _75282_;
wire _75283_;
wire _75284_;
wire _75285_;
wire _75286_;
wire _75287_;
wire _75288_;
wire _75289_;
wire _75290_;
wire _75291_;
wire _75292_;
wire _75293_;
wire _75294_;
wire _75295_;
wire _75296_;
wire _75297_;
wire _75298_;
wire _75299_;
wire _75300_;
wire _75301_;
wire _75302_;
wire _75303_;
wire _75304_;
wire _75305_;
wire _75306_;
wire _75307_;
wire _75308_;
wire _75309_;
wire _75310_;
wire _75311_;
wire _75312_;
wire _75313_;
wire _75314_;
wire _75315_;
wire _75316_;
wire _75317_;
wire _75318_;
wire _75319_;
wire _75320_;
wire _75321_;
wire _75322_;
wire _75323_;
wire _75324_;
wire _75325_;
wire _75326_;
wire _75327_;
wire _75328_;
wire _75329_;
wire _75330_;
wire _75331_;
wire _75332_;
wire _75333_;
wire _75334_;
wire _75335_;
wire _75336_;
wire _75337_;
wire _75338_;
wire _75339_;
wire _75340_;
wire _75341_;
wire _75342_;
wire _75343_;
wire _75344_;
wire _75345_;
wire _75346_;
wire _75347_;
wire _75348_;
wire _75349_;
wire _75350_;
wire _75351_;
wire _75352_;
wire _75353_;
wire _75354_;
wire _75355_;
wire _75356_;
wire _75357_;
wire _75358_;
wire _75359_;
wire _75360_;
wire _75361_;
wire _75362_;
wire _75363_;
wire _75364_;
wire _75365_;
wire _75366_;
wire _75367_;
wire _75368_;
wire _75369_;
wire _75370_;
wire _75371_;
wire _75372_;
wire _75373_;
wire _75374_;
wire _75375_;
wire _75376_;
wire _75377_;
wire _75378_;
wire _75379_;
wire _75380_;
wire _75381_;
wire _75382_;
wire _75383_;
wire _75384_;
wire _75385_;
wire _75386_;
wire _75387_;
wire _75388_;
wire _75389_;
wire _75390_;
wire _75391_;
wire _75392_;
wire _75393_;
wire _75394_;
wire _75395_;
wire _75396_;
wire _75397_;
wire _75398_;
wire _75399_;
wire _75400_;
wire _75401_;
wire _75402_;
wire _75403_;
wire _75404_;
wire _75405_;
wire _75406_;
wire _75407_;
wire _75408_;
wire _75409_;
wire _75410_;
wire _75411_;
wire _75412_;
wire _75413_;
wire _75414_;
wire _75415_;
wire _75416_;
wire _75417_;
wire _75418_;
wire _75419_;
wire _75420_;
wire _75421_;
wire _75422_;
wire _75423_;
wire _75424_;
wire _75425_;
wire _75426_;
wire _75427_;
wire _75428_;
wire _75429_;
wire _75430_;
wire _75431_;
wire _75432_;
wire _75433_;
wire _75434_;
wire _75435_;
wire _75436_;
wire _75437_;
wire _75438_;
wire _75439_;
wire _75440_;
wire _75441_;
wire _75442_;
wire _75443_;
wire _75444_;
wire _75445_;
wire _75446_;
wire _75447_;
wire _75448_;
wire _75449_;
wire _75450_;
wire _75451_;
wire _75452_;
wire _75453_;
wire _75454_;
wire _75455_;
wire _75456_;
wire _75457_;
wire _75458_;
wire _75459_;
wire _75460_;
wire _75461_;
wire _75462_;
wire _75463_;
wire _75464_;
wire _75465_;
wire _75466_;
wire _75467_;
wire _75468_;
wire _75469_;
wire _75470_;
wire _75471_;
wire _75472_;
wire _75473_;
wire _75474_;
wire _75475_;
wire _75476_;
wire _75477_;
wire _75478_;
wire _75479_;
wire _75480_;
wire _75481_;
wire _75482_;
wire _75483_;
wire _75484_;
wire _75485_;
wire _75486_;
wire _75487_;
wire _75488_;
wire _75489_;
wire _75490_;
wire _75491_;
wire _75492_;
wire _75493_;
wire _75494_;
wire _75495_;
wire _75496_;
wire _75497_;
wire _75498_;
wire _75499_;
wire _75500_;
wire _75501_;
wire _75502_;
wire _75503_;
wire _75504_;
wire _75505_;
wire _75506_;
wire _75507_;
wire _75508_;
wire _75509_;
wire _75510_;
wire _75511_;
wire _75512_;
wire _75513_;
wire _75514_;
wire _75515_;
wire _75516_;
wire _75517_;
wire _75518_;
wire _75519_;
wire _75520_;
wire _75521_;
wire _75522_;
wire _75523_;
wire _75524_;
wire _75525_;
wire _75526_;
wire _75527_;
wire _75528_;
wire _75529_;
wire _75530_;
wire _75531_;
wire _75532_;
wire _75533_;
wire _75534_;
wire _75535_;
wire _75536_;
wire _75537_;
wire _75538_;
wire _75539_;
wire _75540_;
wire _75541_;
wire _75542_;
wire _75543_;
wire _75544_;
wire _75545_;
wire _75546_;
wire _75547_;
wire _75548_;
wire _75549_;
wire _75550_;
wire _75551_;
wire _75552_;
wire _75553_;
wire _75554_;
wire _75555_;
wire _75556_;
wire _75557_;
wire _75558_;
wire _75559_;
wire _75560_;
wire _75561_;
wire _75562_;
wire _75563_;
wire _75564_;
wire _75565_;
wire _75566_;
wire _75567_;
wire _75568_;
wire _75569_;
wire _75570_;
wire _75571_;
wire _75572_;
wire _75573_;
wire _75574_;
wire _75575_;
wire _75576_;
wire _75577_;
wire _75578_;
wire _75579_;
wire _75580_;
wire _75581_;
wire _75582_;
wire _75583_;
wire _75584_;
wire _75585_;
wire _75586_;
wire _75587_;
wire _75588_;
wire _75589_;
wire _75590_;
wire _75591_;
wire _75592_;
wire _75593_;
wire _75594_;
wire _75595_;
wire _75596_;
wire _75597_;
wire _75598_;
wire _75599_;
wire _75600_;
wire _75601_;
wire _75602_;
wire _75603_;
wire _75604_;
wire _75605_;
wire _75606_;
wire _75607_;
wire _75608_;
wire _75609_;
wire _75610_;
wire _75611_;
wire _75612_;
wire _75613_;
wire _75614_;
wire _75615_;
wire _75616_;
wire _75617_;
wire _75618_;
wire _75619_;
wire _75620_;
wire _75621_;
wire _75622_;
wire _75623_;
wire _75624_;
wire _75625_;
wire _75626_;
wire _75627_;
wire _75628_;
wire _75629_;
wire _75630_;
wire _75631_;
wire _75632_;
wire _75633_;
wire _75634_;
wire _75635_;
wire _75636_;
wire _75637_;
wire _75638_;
wire _75639_;
wire _75640_;
wire _75641_;
wire _75642_;
wire _75643_;
wire _75644_;
wire _75645_;
wire _75646_;
wire _75647_;
wire _75648_;
wire _75649_;
wire _75650_;
wire _75651_;
wire _75652_;
wire _75653_;
wire _75654_;
wire _75655_;
wire _75656_;
wire _75657_;
wire _75658_;
wire _75659_;
wire _75660_;
wire _75661_;
wire _75662_;
wire _75663_;
wire _75664_;
wire _75665_;
wire _75666_;
wire _75667_;
wire _75668_;
wire _75669_;
wire _75670_;
wire _75671_;
wire _75672_;
wire _75673_;
wire _75674_;
wire _75675_;
wire _75676_;
wire _75677_;
wire _75678_;
wire _75679_;
wire _75680_;
wire _75681_;
wire _75682_;
wire _75683_;
wire _75684_;
wire _75685_;
wire _75686_;
wire _75687_;
wire _75688_;
wire _75689_;
wire _75690_;
wire _75691_;
wire _75692_;
wire _75693_;
wire _75694_;
wire _75695_;
wire _75696_;
wire _75697_;
wire _75698_;
wire _75699_;
wire _75700_;
wire _75701_;
wire _75702_;
wire _75703_;
wire _75704_;
wire _75705_;
wire _75706_;
wire _75707_;
wire _75708_;
wire _75709_;
wire _75710_;
wire _75711_;
wire _75712_;
wire _75713_;
wire _75714_;
wire _75715_;
wire _75716_;
wire _75717_;
wire _75718_;
wire _75719_;
wire _75720_;
wire _75721_;
wire _75722_;
wire _75723_;
wire _75724_;
wire _75725_;
wire _75726_;
wire _75727_;
wire _75728_;
wire _75729_;
wire _75730_;
wire _75731_;
wire _75732_;
wire _75733_;
wire _75734_;
wire _75735_;
wire _75736_;
wire _75737_;
wire _75738_;
wire _75739_;
wire _75740_;
wire _75741_;
wire _75742_;
wire _75743_;
wire _75744_;
wire _75745_;
wire _75746_;
wire _75747_;
wire _75748_;
wire _75749_;
wire _75750_;
wire _75751_;
wire _75752_;
wire _75753_;
wire _75754_;
wire _75755_;
wire _75756_;
wire _75757_;
wire _75758_;
wire _75759_;
wire _75760_;
wire _75761_;
wire _75762_;
wire _75763_;
wire _75764_;
wire _75765_;
wire _75766_;
wire _75767_;
wire _75768_;
wire _75769_;
wire _75770_;
wire _75771_;
wire _75772_;
wire _75773_;
wire _75774_;
wire _75775_;
wire _75776_;
wire _75777_;
wire _75778_;
wire _75779_;
wire _75780_;
wire _75781_;
wire _75782_;
wire _75783_;
wire _75784_;
wire _75785_;
wire _75786_;
wire _75787_;
wire _75788_;
wire _75789_;
wire _75790_;
wire _75791_;
wire _75792_;
wire _75793_;
wire _75794_;
wire _75795_;
wire _75796_;
wire _75797_;
wire _75798_;
wire _75799_;
wire _75800_;
wire _75801_;
wire _75802_;
wire _75803_;
wire _75804_;
wire _75805_;
wire _75806_;
wire _75807_;
wire _75808_;
wire _75809_;
wire _75810_;
wire _75811_;
wire _75812_;
wire _75813_;
wire _75814_;
wire _75815_;
wire _75816_;
wire _75817_;
wire _75818_;
wire _75819_;
wire _75820_;
wire _75821_;
wire _75822_;
wire _75823_;
wire _75824_;
wire _75825_;
wire _75826_;
wire _75827_;
wire _75828_;
wire _75829_;
wire _75830_;
wire _75831_;
wire _75832_;
wire _75833_;
wire _75834_;
wire _75835_;
wire _75836_;
wire _75837_;
wire _75838_;
wire _75839_;
wire _75840_;
wire _75841_;
wire _75842_;
wire _75843_;
wire _75844_;
wire _75845_;
wire _75846_;
wire _75847_;
wire _75848_;
wire _75849_;
wire _75850_;
wire _75851_;
wire _75852_;
wire _75853_;
wire _75854_;
wire _75855_;
wire _75856_;
wire _75857_;
wire _75858_;
wire _75859_;
wire _75860_;
wire _75861_;
wire _75862_;
wire _75863_;
wire _75864_;
wire _75865_;
wire _75866_;
wire _75867_;
wire _75868_;
wire _75869_;
wire _75870_;
wire _75871_;
wire _75872_;
wire _75873_;
wire _75874_;
wire _75875_;
wire _75876_;
wire _75877_;
wire _75878_;
wire _75879_;
wire _75880_;
wire _75881_;
wire _75882_;
wire _75883_;
wire _75884_;
wire _75885_;
wire _75886_;
wire _75887_;
wire _75888_;
wire _75889_;
wire _75890_;
wire _75891_;
wire _75892_;
wire _75893_;
wire _75894_;
wire _75895_;
wire _75896_;
wire _75897_;
wire _75898_;
wire _75899_;
wire _75900_;
wire _75901_;
wire _75902_;
wire _75903_;
wire _75904_;
wire _75905_;
wire _75906_;
wire _75907_;
wire _75908_;
wire _75909_;
wire _75910_;
wire _75911_;
wire _75912_;
wire _75913_;
wire _75914_;
wire _75915_;
wire _75916_;
wire _75917_;
wire _75918_;
wire _75919_;
wire _75920_;
wire _75921_;
wire _75922_;
wire _75923_;
wire _75924_;
wire _75925_;
wire _75926_;
wire _75927_;
wire _75928_;
wire _75929_;
wire _75930_;
wire _75931_;
wire _75932_;
wire _75933_;
wire _75934_;
wire _75935_;
wire _75936_;
wire _75937_;
wire _75938_;
wire _75939_;
wire _75940_;
wire _75941_;
wire _75942_;
wire _75943_;
wire _75944_;
wire _75945_;
wire _75946_;
wire _75947_;
wire _75948_;
wire _75949_;
wire _75950_;
wire _75951_;
wire _75952_;
wire _75953_;
wire _75954_;
wire _75955_;
wire _75956_;
wire _75957_;
wire _75958_;
wire _75959_;
wire _75960_;
wire _75961_;
wire _75962_;
wire _75963_;
wire _75964_;
wire _75965_;
wire _75966_;
wire _75967_;
wire _75968_;
wire _75969_;
wire _75970_;
wire _75971_;
wire _75972_;
wire _75973_;
wire _75974_;
wire _75975_;
wire _75976_;
wire _75977_;
wire _75978_;
wire _75979_;
wire _75980_;
wire _75981_;
wire _75982_;
wire _75983_;
wire _75984_;
wire _75985_;
wire _75986_;
wire _75987_;
wire _75988_;
wire _75989_;
wire _75990_;
wire _75991_;
wire _75992_;
wire _75993_;
wire _75994_;
wire _75995_;
wire _75996_;
wire _75997_;
wire _75998_;
wire _75999_;
wire _76000_;
wire _76001_;
wire _76002_;
wire _76003_;
wire _76004_;
wire _76005_;
wire _76006_;
wire _76007_;
wire _76008_;
wire _76009_;
wire _76010_;
wire _76011_;
wire _76012_;
wire _76013_;
wire _76014_;
wire _76015_;
wire _76016_;
wire _76017_;
wire _76018_;
wire _76019_;
wire _76020_;
wire _76021_;
wire _76022_;
wire _76023_;
wire _76024_;
wire _76025_;
wire _76026_;
wire _76027_;
wire _76028_;
wire _76029_;
wire _76030_;
wire _76031_;
wire _76032_;
wire _76033_;
wire _76034_;
wire _76035_;
wire _76036_;
wire _76037_;
wire _76038_;
wire _76039_;
wire _76040_;
wire _76041_;
wire _76042_;
wire _76043_;
wire _76044_;
wire _76045_;
wire _76046_;
wire _76047_;
wire _76048_;
wire _76049_;
wire _76050_;
wire _76051_;
wire _76052_;
wire _76053_;
wire _76054_;
wire _76055_;
wire _76056_;
wire _76057_;
wire _76058_;
wire _76059_;
wire _76060_;
wire _76061_;
wire _76062_;
wire _76063_;
wire _76064_;
wire _76065_;
wire _76066_;
wire _76067_;
wire _76068_;
wire _76069_;
wire _76070_;
wire _76071_;
wire _76072_;
wire _76073_;
wire _76074_;
wire _76075_;
wire _76076_;
wire _76077_;
wire _76078_;
wire _76079_;
wire _76080_;
wire _76081_;
wire _76082_;
wire _76083_;
wire _76084_;
wire _76085_;
wire _76086_;
wire _76087_;
wire _76088_;
wire _76089_;
wire _76090_;
wire _76091_;
wire _76092_;
wire _76093_;
wire _76094_;
wire _76095_;
wire _76096_;
wire _76097_;
wire _76098_;
wire _76099_;
wire _76100_;
wire _76101_;
wire _76102_;
wire _76103_;
wire _76104_;
wire _76105_;
wire _76106_;
wire _76107_;
wire _76108_;
wire _76109_;
wire _76110_;
wire _76111_;
wire _76112_;
wire _76113_;
wire _76114_;
wire _76115_;
wire _76116_;
wire _76117_;
wire _76118_;
wire _76119_;
wire _76120_;
wire _76121_;
wire _76122_;
wire _76123_;
wire _76124_;
wire _76125_;
wire _76126_;
wire _76127_;
wire _76128_;
wire _76129_;
wire _76130_;
wire _76131_;
wire _76132_;
wire _76133_;
wire _76134_;
wire _76135_;
wire _76136_;
wire _76137_;
wire _76138_;
wire _76139_;
wire _76140_;
wire _76141_;
wire _76142_;
wire _76143_;
wire _76144_;
wire _76145_;
wire _76146_;
wire _76147_;
wire _76148_;
wire _76149_;
wire _76150_;
wire _76151_;
wire _76152_;
wire _76153_;
wire _76154_;
wire _76155_;
wire _76156_;
wire _76157_;
wire _76158_;
wire _76159_;
wire _76160_;
wire _76161_;
wire _76162_;
wire _76163_;
wire _76164_;
wire _76165_;
wire _76166_;
wire _76167_;
wire _76168_;
wire _76169_;
wire _76170_;
wire _76171_;
wire _76172_;
wire _76173_;
wire _76174_;
wire _76175_;
wire _76176_;
wire _76177_;
wire _76178_;
wire _76179_;
wire _76180_;
wire _76181_;
wire _76182_;
wire _76183_;
wire _76184_;
wire _76185_;
wire _76186_;
wire _76187_;
wire _76188_;
wire _76189_;
wire _76190_;
wire _76191_;
wire _76192_;
wire _76193_;
wire _76194_;
wire _76195_;
wire _76196_;
wire _76197_;
wire _76198_;
wire _76199_;
wire _76200_;
wire _76201_;
wire _76202_;
wire _76203_;
wire _76204_;
wire _76205_;
wire _76206_;
wire _76207_;
wire _76208_;
wire _76209_;
wire _76210_;
wire _76211_;
wire _76212_;
wire _76213_;
wire _76214_;
wire _76215_;
wire _76216_;
wire _76217_;
wire _76218_;
wire _76219_;
wire _76220_;
wire _76221_;
wire _76222_;
wire _76223_;
wire _76224_;
wire _76225_;
wire _76226_;
wire _76227_;
wire _76228_;
wire _76229_;
wire _76230_;
wire _76231_;
wire _76232_;
wire _76233_;
wire _76234_;
wire _76235_;
wire _76236_;
wire _76237_;
wire _76238_;
wire _76239_;
wire _76240_;
wire _76241_;
wire _76242_;
wire _76243_;
wire _76244_;
wire _76245_;
wire _76246_;
wire _76247_;
wire _76248_;
wire _76249_;
wire _76250_;
wire _76251_;
wire _76252_;
wire _76253_;
wire _76254_;
wire _76255_;
wire _76256_;
wire _76257_;
wire _76258_;
wire _76259_;
wire _76260_;
wire _76261_;
wire _76262_;
wire _76263_;
wire _76264_;
wire _76265_;
wire _76266_;
wire _76267_;
wire _76268_;
wire _76269_;
wire _76270_;
wire _76271_;
wire _76272_;
wire _76273_;
wire _76274_;
wire _76275_;
wire _76276_;
wire _76277_;
wire _76278_;
wire _76279_;
wire _76280_;
wire _76281_;
wire _76282_;
wire _76283_;
wire _76284_;
wire _76285_;
wire _76286_;
wire _76287_;
wire _76288_;
wire _76289_;
wire _76290_;
wire _76291_;
wire _76292_;
wire _76293_;
wire _76294_;
wire _76295_;
wire _76296_;
wire _76297_;
wire _76298_;
wire _76299_;
wire _76300_;
wire _76301_;
wire _76302_;
wire _76303_;
wire _76304_;
wire _76305_;
wire _76306_;
wire _76307_;
wire _76308_;
wire _76309_;
wire _76310_;
wire _76311_;
wire _76312_;
wire _76313_;
wire _76314_;
wire _76315_;
wire _76316_;
wire _76317_;
wire _76318_;
wire _76319_;
wire _76320_;
wire _76321_;
wire _76322_;
wire _76323_;
wire _76324_;
wire _76325_;
wire _76326_;
wire _76327_;
wire _76328_;
wire _76329_;
wire _76330_;
wire _76331_;
wire _76332_;
wire _76333_;
wire _76334_;
wire _76335_;
wire _76336_;
wire _76337_;
wire _76338_;
wire _76339_;
wire _76340_;
wire _76341_;
wire _76342_;
wire _76343_;
wire _76344_;
wire _76345_;
wire _76346_;
wire _76347_;
wire _76348_;
wire _76349_;
wire _76350_;
wire _76351_;
wire _76352_;
wire _76353_;
wire _76354_;
wire _76355_;
wire _76356_;
wire _76357_;
wire _76358_;
wire _76359_;
wire _76360_;
wire _76361_;
wire _76362_;
wire _76363_;
wire _76364_;
wire _76365_;
wire _76366_;
wire _76367_;
wire _76368_;
wire _76369_;
wire _76370_;
wire _76371_;
wire _76372_;
wire _76373_;
wire _76374_;
wire _76375_;
wire _76376_;
wire _76377_;
wire _76378_;
wire _76379_;
wire _76380_;
wire _76381_;
wire _76382_;
wire _76383_;
wire _76384_;
wire _76385_;
wire _76386_;
wire _76387_;
wire _76388_;
wire _76389_;
wire _76390_;
wire _76391_;
wire _76392_;
wire _76393_;
wire _76394_;
wire _76395_;
wire _76396_;
wire _76397_;
wire _76398_;
wire _76399_;
wire _76400_;
wire _76401_;
wire _76402_;
wire _76403_;
wire _76404_;
wire _76405_;
wire _76406_;
wire _76407_;
wire _76408_;
wire _76409_;
wire _76410_;
wire _76411_;
wire _76412_;
wire _76413_;
wire _76414_;
wire _76415_;
wire _76416_;
wire _76417_;
wire _76418_;
wire _76419_;
wire _76420_;
wire _76421_;
wire _76422_;
wire _76423_;
wire _76424_;
wire _76425_;
wire _76426_;
wire _76427_;
wire _76428_;
wire _76429_;
wire _76430_;
wire _76431_;
wire _76432_;
wire _76433_;
wire _76434_;
wire _76435_;
wire _76436_;
wire _76437_;
wire _76438_;
wire _76439_;
wire _76440_;
wire _76441_;
wire _76442_;
wire _76443_;
wire _76444_;
wire _76445_;
wire _76446_;
wire _76447_;
wire _76448_;
wire _76449_;
wire _76450_;
wire _76451_;
wire _76452_;
wire _76453_;
wire _76454_;
wire _76455_;
wire _76456_;
wire _76457_;
wire _76458_;
wire _76459_;
wire _76460_;
wire _76461_;
wire _76462_;
wire _76463_;
wire _76464_;
wire _76465_;
wire _76466_;
wire _76467_;
wire _76468_;
wire _76469_;
wire _76470_;
wire _76471_;
wire _76472_;
wire _76473_;
wire _76474_;
wire _76475_;
wire _76476_;
wire _76477_;
wire _76478_;
wire _76479_;
wire _76480_;
wire _76481_;
wire _76482_;
wire _76483_;
wire _76484_;
wire _76485_;
wire _76486_;
wire _76487_;
wire _76488_;
wire _76489_;
wire _76490_;
wire _76491_;
wire _76492_;
wire _76493_;
wire _76494_;
wire _76495_;
wire _76496_;
wire _76497_;
wire _76498_;
wire _76499_;
wire _76500_;
wire _76501_;
wire _76502_;
wire _76503_;
wire _76504_;
wire _76505_;
wire _76506_;
wire _76507_;
wire _76508_;
wire _76509_;
wire _76510_;
wire _76511_;
wire _76512_;
wire _76513_;
wire _76514_;
wire _76515_;
wire _76516_;
wire _76517_;
wire _76518_;
wire _76519_;
wire _76520_;
wire _76521_;
wire _76522_;
wire _76523_;
wire _76524_;
wire _76525_;
wire _76526_;
wire _76527_;
wire _76528_;
wire _76529_;
wire _76530_;
wire _76531_;
wire _76532_;
wire _76533_;
wire _76534_;
wire _76535_;
wire _76536_;
wire _76537_;
wire _76538_;
wire _76539_;
wire _76540_;
wire _76541_;
wire _76542_;
wire _76543_;
wire _76544_;
wire _76545_;
wire _76546_;
wire _76547_;
wire _76548_;
wire _76549_;
wire _76550_;
wire _76551_;
wire _76552_;
wire _76553_;
wire _76554_;
wire _76555_;
wire _76556_;
wire _76557_;
wire _76558_;
wire _76559_;
wire _76560_;
wire _76561_;
wire _76562_;
wire _76563_;
wire _76564_;
wire _76565_;
wire _76566_;
wire _76567_;
wire _76568_;
wire _76569_;
wire _76570_;
wire _76571_;
wire _76572_;
wire _76573_;
wire _76574_;
wire _76575_;
wire _76576_;
wire _76577_;
wire _76578_;
wire _76579_;
wire _76580_;
wire _76581_;
wire _76582_;
wire _76583_;
wire _76584_;
wire _76585_;
wire _76586_;
wire _76587_;
wire _76588_;
wire _76589_;
wire _76590_;
wire _76591_;
wire _76592_;
wire _76593_;
wire _76594_;
wire _76595_;
wire _76596_;
wire _76597_;
wire _76598_;
wire _76599_;
wire _76600_;
wire _76601_;
wire _76602_;
wire _76603_;
wire _76604_;
wire _76605_;
wire _76606_;
wire _76607_;
wire _76608_;
wire _76609_;
wire _76610_;
wire _76611_;
wire _76612_;
wire _76613_;
wire _76614_;
wire _76615_;
wire _76616_;
wire _76617_;
wire _76618_;
wire _76619_;
wire _76620_;
wire _76621_;
wire _76622_;
wire _76623_;
wire _76624_;
wire _76625_;
wire _76626_;
wire _76627_;
wire _76628_;
wire _76629_;
wire _76630_;
wire _76631_;
wire _76632_;
wire _76633_;
wire _76634_;
wire _76635_;
wire _76636_;
wire _76637_;
wire _76638_;
wire _76639_;
wire _76640_;
wire _76641_;
wire _76642_;
wire _76643_;
wire _76644_;
wire _76645_;
wire _76646_;
wire _76647_;
wire _76648_;
wire _76649_;
wire _76650_;
wire _76651_;
wire _76652_;
wire _76653_;
wire _76654_;
wire _76655_;
wire _76656_;
wire _76657_;
wire _76658_;
wire _76659_;
wire _76660_;
wire _76661_;
wire _76662_;
wire _76663_;
wire _76664_;
wire _76665_;
wire _76666_;
wire _76667_;
wire _76668_;
wire _76669_;
wire _76670_;
wire _76671_;
wire _76672_;
wire _76673_;
wire _76674_;
wire _76675_;
wire _76676_;
wire _76677_;
wire _76678_;
wire _76679_;
wire _76680_;
wire _76681_;
wire _76682_;
wire _76683_;
wire _76684_;
wire _76685_;
wire _76686_;
wire _76687_;
wire _76688_;
wire _76689_;
wire _76690_;
wire _76691_;
wire _76692_;
wire _76693_;
wire _76694_;
wire _76695_;
wire _76696_;
wire _76697_;
wire _76698_;
wire _76699_;
wire _76700_;
wire _76701_;
wire _76702_;
wire _76703_;
wire _76704_;
wire _76705_;
wire _76706_;
wire _76707_;
wire _76708_;
wire _76709_;
wire _76710_;
wire _76711_;
wire _76712_;
wire _76713_;
wire _76714_;
wire _76715_;
wire _76716_;
wire _76717_;
wire _76718_;
wire _76719_;
wire _76720_;
wire _76721_;
wire _76722_;
wire _76723_;
wire _76724_;
wire _76725_;
wire _76726_;
wire _76727_;
wire _76728_;
wire _76729_;
wire _76730_;
wire _76731_;
wire _76732_;
wire _76733_;
wire _76734_;
wire _76735_;
wire _76736_;
wire _76737_;
wire _76738_;
wire _76739_;
wire _76740_;
wire _76741_;
wire _76742_;
wire _76743_;
wire _76744_;
wire _76745_;
wire _76746_;
wire _76747_;
wire _76748_;
wire _76749_;
wire _76750_;
wire _76751_;
wire _76752_;
wire _76753_;
wire _76754_;
wire _76755_;
wire _76756_;
wire _76757_;
wire _76758_;
wire _76759_;
wire _76760_;
wire _76761_;
wire _76762_;
wire _76763_;
wire _76764_;
wire _76765_;
wire _76766_;
wire _76767_;
wire _76768_;
wire _76769_;
wire _76770_;
wire _76771_;
wire _76772_;
wire _76773_;
wire _76774_;
wire _76775_;
wire _76776_;
wire _76777_;
wire _76778_;
wire _76779_;
wire _76780_;
wire _76781_;
wire _76782_;
wire _76783_;
wire _76784_;
wire _76785_;
wire _76786_;
wire _76787_;
wire _76788_;
wire _76789_;
wire _76790_;
wire _76791_;
wire _76792_;
wire _76793_;
wire _76794_;
wire _76795_;
wire _76796_;
wire _76797_;
wire _76798_;
wire _76799_;
wire _76800_;
wire _76801_;
wire _76802_;
wire _76803_;
wire _76804_;
wire _76805_;
wire _76806_;
wire _76807_;
wire _76808_;
wire _76809_;
wire _76810_;
wire _76811_;
wire _76812_;
wire _76813_;
wire _76814_;
wire _76815_;
wire _76816_;
wire _76817_;
wire _76818_;
wire _76819_;
wire _76820_;
wire _76821_;
wire _76822_;
wire _76823_;
wire _76824_;
wire _76825_;
wire _76826_;
wire _76827_;
wire _76828_;
wire _76829_;
wire _76830_;
wire _76831_;
wire _76832_;
wire _76833_;
wire _76834_;
wire _76835_;
wire _76836_;
wire _76837_;
wire _76838_;
wire _76839_;
wire _76840_;
wire _76841_;
wire _76842_;
wire _76843_;
wire _76844_;
wire _76845_;
wire _76846_;
wire _76847_;
wire _76848_;
wire _76849_;
wire _76850_;
wire _76851_;
wire _76852_;
wire _76853_;
wire _76854_;
wire _76855_;
wire _76856_;
wire _76857_;
wire _76858_;
wire _76859_;
wire _76860_;
wire _76861_;
wire _76862_;
wire _76863_;
wire _76864_;
wire _76865_;
wire _76866_;
wire _76867_;
wire _76868_;
wire _76869_;
wire _76870_;
wire _76871_;
wire _76872_;
wire _76873_;
wire _76874_;
wire _76875_;
wire _76876_;
wire _76877_;
wire _76878_;
wire _76879_;
wire _76880_;
wire _76881_;
wire _76882_;
wire _76883_;
wire _76884_;
wire _76885_;
wire _76886_;
wire _76887_;
wire _76888_;
wire _76889_;
wire _76890_;
wire _76891_;
wire _76892_;
wire _76893_;
wire _76894_;
wire _76895_;
wire _76896_;
wire _76897_;
wire _76898_;
wire _76899_;
wire _76900_;
wire _76901_;
wire _76902_;
wire _76903_;
wire _76904_;
wire _76905_;
wire _76906_;
wire _76907_;
wire _76908_;
wire _76909_;
wire _76910_;
wire _76911_;
wire _76912_;
wire _76913_;
wire _76914_;
wire _76915_;
wire _76916_;
wire _76917_;
wire _76918_;
wire _76919_;
wire _76920_;
wire _76921_;
wire _76922_;
wire _76923_;
wire _76924_;
wire _76925_;
wire _76926_;
wire _76927_;
wire _76928_;
wire _76929_;
wire _76930_;
wire _76931_;
wire _76932_;
wire _76933_;
wire _76934_;
wire _76935_;
wire _76936_;
wire _76937_;
wire _76938_;
wire _76939_;
wire _76940_;
wire _76941_;
wire _76942_;
wire _76943_;
wire _76944_;
wire _76945_;
wire _76946_;
wire _76947_;
wire _76948_;
wire _76949_;
wire _76950_;
wire _76951_;
wire _76952_;
wire _76953_;
wire _76954_;
wire _76955_;
wire _76956_;
wire _76957_;
wire _76958_;
wire _76959_;
wire _76960_;
wire _76961_;
wire _76962_;
wire _76963_;
wire _76964_;
wire _76965_;
wire _76966_;
wire _76967_;
wire _76968_;
wire _76969_;
wire _76970_;
wire _76971_;
wire _76972_;
wire _76973_;
wire _76974_;
wire _76975_;
wire _76976_;
wire _76977_;
wire _76978_;
wire _76979_;
wire _76980_;
wire _76981_;
wire _76982_;
wire _76983_;
wire _76984_;
wire _76985_;
wire _76986_;
wire _76987_;
wire _76988_;
wire _76989_;
wire _76990_;
wire _76991_;
wire _76992_;
wire _76993_;
wire _76994_;
wire _76995_;
wire _76996_;
wire _76997_;
wire _76998_;
wire _76999_;
wire _77000_;
wire _77001_;
wire _77002_;
wire _77003_;
wire _77004_;
wire _77005_;
wire _77006_;
wire _77007_;
wire _77008_;
wire _77009_;
wire _77010_;
wire _77011_;
wire _77012_;
wire _77013_;
wire _77014_;
wire _77015_;
wire _77016_;
wire _77017_;
wire _77018_;
wire _77019_;
wire _77020_;
wire _77021_;
wire _77022_;
wire _77023_;
wire _77024_;
wire _77025_;
wire _77026_;
wire _77027_;
wire _77028_;
wire _77029_;
wire _77030_;
wire _77031_;
wire _77032_;
wire _77033_;
wire _77034_;
wire _77035_;
wire _77036_;
wire _77037_;
wire _77038_;
wire _77039_;
wire _77040_;
wire _77041_;
wire _77042_;
wire _77043_;
wire _77044_;
wire _77045_;
wire _77046_;
wire _77047_;
wire _77048_;
wire _77049_;
wire _77050_;
wire _77051_;
wire _77052_;
wire _77053_;
wire _77054_;
wire _77055_;
wire _77056_;
wire _77057_;
wire _77058_;
wire _77059_;
wire _77060_;
wire _77061_;
wire _77062_;
wire _77063_;
wire _77064_;
wire _77065_;
wire _77066_;
wire _77067_;
wire _77068_;
wire _77069_;
wire _77070_;
wire _77071_;
wire _77072_;
wire _77073_;
wire _77074_;
wire _77075_;
wire _77076_;
wire _77077_;
wire _77078_;
wire _77079_;
wire _77080_;
wire _77081_;
wire _77082_;
wire _77083_;
wire _77084_;
wire _77085_;
wire _77086_;
wire _77087_;
wire _77088_;
wire _77089_;
wire _77090_;
wire _77091_;
wire _77092_;
wire _77093_;
wire _77094_;
wire _77095_;
wire _77096_;
wire _77097_;
wire _77098_;
wire _77099_;
wire _77100_;
wire _77101_;
wire _77102_;
wire _77103_;
wire _77104_;
wire _77105_;
wire _77106_;
wire _77107_;
wire _77108_;
wire _77109_;
wire _77110_;
wire _77111_;
wire _77112_;
wire _77113_;
wire _77114_;
wire _77115_;
wire _77116_;
wire _77117_;
wire _77118_;
wire _77119_;
wire _77120_;
wire _77121_;
wire _77122_;
wire _77123_;
wire _77124_;
wire _77125_;
wire _77126_;
wire _77127_;
wire _77128_;
wire _77129_;
wire _77130_;
wire _77131_;
wire _77132_;
wire _77133_;
wire _77134_;
wire _77135_;
wire _77136_;
wire _77137_;
wire _77138_;
wire _77139_;
wire _77140_;
wire _77141_;
wire _77142_;
wire _77143_;
wire _77144_;
wire _77145_;
wire _77146_;
wire _77147_;
wire _77148_;
wire _77149_;
wire _77150_;
wire _77151_;
wire _77152_;
wire _77153_;
wire _77154_;
wire _77155_;
wire _77156_;
wire _77157_;
wire _77158_;
wire _77159_;
wire _77160_;
wire _77161_;
wire _77162_;
wire _77163_;
wire _77164_;
wire _77165_;
wire _77166_;
wire _77167_;
wire _77168_;
wire _77169_;
wire _77170_;
wire _77171_;
wire _77172_;
wire _77173_;
wire _77174_;
wire _77175_;
wire _77176_;
wire _77177_;
wire _77178_;
wire _77179_;
wire _77180_;
wire _77181_;
wire _77182_;
wire _77183_;
wire _77184_;
wire _77185_;
wire _77186_;
wire _77187_;
wire _77188_;
wire _77189_;
wire _77190_;
wire _77191_;
wire _77192_;
wire _77193_;
wire _77194_;
wire _77195_;
wire _77196_;
wire _77197_;
wire _77198_;
wire _77199_;
wire _77200_;
wire _77201_;
wire _77202_;
wire _77203_;
wire _77204_;
wire _77205_;
wire _77206_;
wire _77207_;
wire _77208_;
wire _77209_;
wire _77210_;
wire _77211_;
wire _77212_;
wire _77213_;
wire _77214_;
wire _77215_;
wire _77216_;
wire _77217_;
wire _77218_;
wire _77219_;
wire _77220_;
wire _77221_;
wire _77222_;
wire _77223_;
wire _77224_;
wire _77225_;
wire _77226_;
wire _77227_;
wire _77228_;
wire _77229_;
wire _77230_;
wire _77231_;
wire _77232_;
wire _77233_;
wire _77234_;
wire _77235_;
wire _77236_;
wire _77237_;
wire _77238_;
wire _77239_;
wire _77240_;
wire _77241_;
wire _77242_;
wire _77243_;
wire _77244_;
wire _77245_;
wire _77246_;
wire _77247_;
wire _77248_;
wire _77249_;
wire _77250_;
wire _77251_;
wire _77252_;
wire _77253_;
wire _77254_;
wire _77255_;
wire _77256_;
wire _77257_;
wire _77258_;
wire _77259_;
wire _77260_;
wire _77261_;
wire _77262_;
wire _77263_;
wire _77264_;
wire _77265_;
wire _77266_;
wire _77267_;
wire _77268_;
wire _77269_;
wire _77270_;
wire _77271_;
wire _77272_;
wire _77273_;
wire _77274_;
wire _77275_;
wire _77276_;
wire _77277_;
wire _77278_;
wire _77279_;
wire _77280_;
wire _77281_;
wire _77282_;
wire _77283_;
wire _77284_;
wire _77285_;
wire _77286_;
wire _77287_;
wire _77288_;
wire _77289_;
wire _77290_;
wire _77291_;
wire _77292_;
wire _77293_;
wire _77294_;
wire _77295_;
wire _77296_;
wire _77297_;
wire _77298_;
wire _77299_;
wire _77300_;
wire _77301_;
wire _77302_;
wire _77303_;
wire _77304_;
wire _77305_;
wire _77306_;
wire _77307_;
wire _77308_;
wire _77309_;
wire _77310_;
wire _77311_;
wire _77312_;
wire _77313_;
wire _77314_;
wire _77315_;
wire _77316_;
wire _77317_;
wire _77318_;
wire _77319_;
wire _77320_;
wire _77321_;
wire _77322_;
wire _77323_;
wire _77324_;
wire _77325_;
wire _77326_;
wire _77327_;
wire _77328_;
wire _77329_;
wire _77330_;
wire _77331_;
wire _77332_;
wire _77333_;
wire _77334_;
wire _77335_;
wire _77336_;
wire _77337_;
wire _77338_;
wire _77339_;
wire _77340_;
wire _77341_;
wire _77342_;
wire _77343_;
wire _77344_;
wire _77345_;
wire _77346_;
wire _77347_;
wire _77348_;
wire _77349_;
wire _77350_;
wire _77351_;
wire _77352_;
wire _77353_;
wire _77354_;
wire _77355_;
wire _77356_;
wire _77357_;
wire _77358_;
wire _77359_;
wire _77360_;
wire _77361_;
wire _77362_;
wire _77363_;
wire _77364_;
wire _77365_;
wire _77366_;
wire _77367_;
wire _77368_;
wire _77369_;
wire _77370_;
wire _77371_;
wire _77372_;
wire _77373_;
wire _77374_;
wire _77375_;
wire _77376_;
wire _77377_;
wire _77378_;
wire _77379_;
wire _77380_;
wire _77381_;
wire _77382_;
wire _77383_;
wire _77384_;
wire _77385_;
wire _77386_;
wire _77387_;
wire _77388_;
wire _77389_;
wire _77390_;
wire _77391_;
wire _77392_;
wire _77393_;
wire _77394_;
wire _77395_;
wire _77396_;
wire _77397_;
wire _77398_;
wire _77399_;
wire _77400_;
wire _77401_;
wire _77402_;
wire _77403_;
wire _77404_;
wire _77405_;
wire _77406_;
wire _77407_;
wire _77408_;
wire _77409_;
wire _77410_;
wire _77411_;
wire _77412_;
wire _77413_;
wire _77414_;
wire _77415_;
wire _77416_;
wire _77417_;
wire _77418_;
wire _77419_;
wire _77420_;
wire _77421_;
wire _77422_;
wire _77423_;
wire _77424_;
wire _77425_;
wire _77426_;
wire _77427_;
wire _77428_;
wire _77429_;
wire _77430_;
wire _77431_;
wire _77432_;
wire _77433_;
wire _77434_;
wire _77435_;
wire _77436_;
wire _77437_;
wire _77438_;
wire _77439_;
wire _77440_;
wire _77441_;
wire _77442_;
wire _77443_;
wire _77444_;
wire _77445_;
wire _77446_;
wire _77447_;
wire _77448_;
wire _77449_;
wire _77450_;
wire _77451_;
wire _77452_;
wire _77453_;
wire _77454_;
wire _77455_;
wire _77456_;
wire _77457_;
wire _77458_;
wire _77459_;
wire _77460_;
wire _77461_;
wire _77462_;
wire _77463_;
wire _77464_;
wire _77465_;
wire _77466_;
wire _77467_;
wire _77468_;
wire _77469_;
wire _77470_;
wire _77471_;
wire _77472_;
wire _77473_;
wire _77474_;
wire _77475_;
wire _77476_;
wire _77477_;
wire _77478_;
wire _77479_;
wire _77480_;
wire _77481_;
wire _77482_;
wire _77483_;
wire _77484_;
wire _77485_;
wire _77486_;
wire _77487_;
wire _77488_;
wire _77489_;
wire _77490_;
wire _77491_;
wire _77492_;
wire _77493_;
wire _77494_;
wire _77495_;
wire _77496_;
wire _77497_;
wire _77498_;
wire _77499_;
wire _77500_;
wire _77501_;
wire _77502_;
wire _77503_;
wire _77504_;
wire _77505_;
wire _77506_;
wire _77507_;
wire _77508_;
wire _77509_;
wire _77510_;
wire _77511_;
wire _77512_;
wire _77513_;
wire _77514_;
wire _77515_;
wire _77516_;
wire _77517_;
wire _77518_;
wire _77519_;
wire _77520_;
wire _77521_;
wire _77522_;
wire _77523_;
wire _77524_;
wire _77525_;
wire _77526_;
wire _77527_;
wire _77528_;
wire _77529_;
wire _77530_;
wire _77531_;
wire _77532_;
wire _77533_;
wire _77534_;
wire _77535_;
wire _77536_;
wire _77537_;
wire _77538_;
wire _77539_;
wire _77540_;
wire _77541_;
wire _77542_;
wire _77543_;
wire _77544_;
wire _77545_;
wire _77546_;
wire _77547_;
wire _77548_;
wire _77549_;
wire _77550_;
wire _77551_;
wire _77552_;
wire _77553_;
wire _77554_;
wire _77555_;
wire _77556_;
wire _77557_;
wire _77558_;
wire _77559_;
wire _77560_;
wire _77561_;
wire _77562_;
wire _77563_;
wire _77564_;
wire _77565_;
wire _77566_;
wire _77567_;
wire _77568_;
wire _77569_;
wire _77570_;
wire _77571_;
wire _77572_;
wire _77573_;
wire _77574_;
wire _77575_;
wire _77576_;
wire _77577_;
wire _77578_;
wire _77579_;
wire _77580_;
wire _77581_;
wire _77582_;
wire _77583_;
wire _77584_;
wire _77585_;
wire _77586_;
wire _77587_;
wire _77588_;
wire _77589_;
wire _77590_;
wire _77591_;
wire _77592_;
wire _77593_;
wire _77594_;
wire _77595_;
wire _77596_;
wire _77597_;
wire _77598_;
wire _77599_;
wire _77600_;
wire _77601_;
wire _77602_;
wire _77603_;
wire _77604_;
wire _77605_;
wire _77606_;
wire _77607_;
wire _77608_;
wire _77609_;
wire _77610_;
wire _77611_;
wire _77612_;
wire _77613_;
wire _77614_;
wire _77615_;
wire _77616_;
wire _77617_;
wire _77618_;
wire _77619_;
wire _77620_;
wire _77621_;
wire _77622_;
wire _77623_;
wire _77624_;
wire _77625_;
wire _77626_;
wire _77627_;
wire _77628_;
wire _77629_;
wire _77630_;
wire _77631_;
wire _77632_;
wire _77633_;
wire _77634_;
wire _77635_;
wire _77636_;
wire _77637_;
wire _77638_;
wire _77639_;
wire _77640_;
wire _77641_;
wire _77642_;
wire _77643_;
wire _77644_;
wire _77645_;
wire _77646_;
wire _77647_;
wire _77648_;
wire _77649_;
wire _77650_;
wire _77651_;
wire _77652_;
wire _77653_;
wire _77654_;
wire _77655_;
wire _77656_;
wire _77657_;
wire _77658_;
wire _77659_;
wire _77660_;
wire _77661_;
wire _77662_;
wire _77663_;
wire _77664_;
wire _77665_;
wire _77666_;
wire _77667_;
wire _77668_;
wire _77669_;
wire _77670_;
wire _77671_;
wire _77672_;
wire _77673_;
wire _77674_;
wire _77675_;
wire _77676_;
wire _77677_;
wire _77678_;
wire _77679_;
wire _77680_;
wire _77681_;
wire _77682_;
wire _77683_;
wire _77684_;
wire _77685_;
wire _77686_;
wire _77687_;
wire _77688_;
wire _77689_;
wire _77690_;
wire _77691_;
wire _77692_;
wire _77693_;
wire _77694_;
wire _77695_;
wire _77696_;
wire _77697_;
wire _77698_;
wire _77699_;
wire _77700_;
wire _77701_;
wire _77702_;
wire _77703_;
wire _77704_;
wire _77705_;
wire _77706_;
wire _77707_;
wire _77708_;
wire _77709_;
wire _77710_;
wire _77711_;
wire _77712_;
wire _77713_;
wire _77714_;
wire _77715_;
wire _77716_;
wire _77717_;
wire _77718_;
wire _77719_;
wire _77720_;
wire _77721_;
wire _77722_;
wire _77723_;
wire _77724_;
wire _77725_;
wire _77726_;
wire _77727_;
wire _77728_;
wire _77729_;
wire _77730_;
wire _77731_;
wire _77732_;
wire _77733_;
wire _77734_;
wire _77735_;
wire _77736_;
wire _77737_;
wire _77738_;
wire _77739_;
wire _77740_;
wire _77741_;
wire _77742_;
wire _77743_;
wire _77744_;
wire _77745_;
wire _77746_;
wire _77747_;
wire _77748_;
wire _77749_;
wire _77750_;
wire _77751_;
wire _77752_;
wire _77753_;
wire _77754_;
wire _77755_;
wire _77756_;
wire _77757_;
wire _77758_;
wire _77759_;
wire _77760_;
wire _77761_;
wire _77762_;
wire _77763_;
wire _77764_;
wire _77765_;
wire _77766_;
wire _77767_;
wire _77768_;
wire _77769_;
wire _77770_;
wire _77771_;
wire _77772_;
wire _77773_;
wire _77774_;
wire _77775_;
wire _77776_;
wire _77777_;
wire _77778_;
wire _77779_;
wire _77780_;
wire _77781_;
wire _77782_;
wire _77783_;
wire _77784_;
wire _77785_;
wire _77786_;
wire _77787_;
wire _77788_;
wire _77789_;
wire _77790_;
wire _77791_;
wire _77792_;
wire _77793_;
wire _77794_;
wire _77795_;
wire _77796_;
wire _77797_;
wire _77798_;
wire _77799_;
wire _77800_;
wire _77801_;
wire _77802_;
wire _77803_;
wire _77804_;
wire _77805_;
wire _77806_;
wire _77807_;
wire _77808_;
wire _77809_;
wire _77810_;
wire _77811_;
wire _77812_;
wire _77813_;
wire _77814_;
wire _77815_;
wire _77816_;
wire _77817_;
wire _77818_;
wire _77819_;
wire _77820_;
wire _77821_;
wire _77822_;
wire _77823_;
wire _77824_;
wire _77825_;
wire _77826_;
wire _77827_;
wire _77828_;
wire _77829_;
wire _77830_;
wire _77831_;
wire _77832_;
wire _77833_;
wire _77834_;
wire _77835_;
wire _77836_;
wire _77837_;
wire _77838_;
wire _77839_;
wire _77840_;
wire _77841_;
wire _77842_;
wire _77843_;
wire _77844_;
wire _77845_;
wire _77846_;
wire _77847_;
wire _77848_;
wire _77849_;
wire _77850_;
wire _77851_;
wire _77852_;
wire _77853_;
wire _77854_;
wire _77855_;
wire _77856_;
wire _77857_;
wire _77858_;
wire _77859_;
wire _77860_;
wire _77861_;
wire _77862_;
wire _77863_;
wire _77864_;
wire _77865_;
wire _77866_;
wire _77867_;
wire _77868_;
wire _77869_;
wire _77870_;
wire _77871_;
wire _77872_;
wire _77873_;
wire _77874_;
wire _77875_;
wire _77876_;
wire _77877_;
wire _77878_;
wire _77879_;
wire _77880_;
wire _77881_;
wire _77882_;
wire _77883_;
wire _77884_;
wire _77885_;
wire _77886_;
wire _77887_;
wire _77888_;
wire _77889_;
wire _77890_;
wire _77891_;
wire _77892_;
wire _77893_;
wire _77894_;
wire _77895_;
wire _77896_;
wire _77897_;
wire _77898_;
wire _77899_;
wire _77900_;
wire _77901_;
wire _77902_;
wire _77903_;
wire _77904_;
wire _77905_;
wire _77906_;
wire _77907_;
wire _77908_;
wire _77909_;
wire _77910_;
wire _77911_;
wire _77912_;
wire _77913_;
wire _77914_;
wire _77915_;
wire _77916_;
wire _77917_;
wire _77918_;
wire _77919_;
wire _77920_;
wire _77921_;
wire _77922_;
wire _77923_;
wire _77924_;
wire _77925_;
wire _77926_;
wire _77927_;
wire _77928_;
wire _77929_;
wire _77930_;
wire _77931_;
wire _77932_;
wire _77933_;
wire _77934_;
wire _77935_;
wire _77936_;
wire _77937_;
wire _77938_;
wire _77939_;
wire _77940_;
wire _77941_;
wire _77942_;
wire _77943_;
wire _77944_;
wire _77945_;
wire _77946_;
wire _77947_;
wire _77948_;
wire _77949_;
wire _77950_;
wire _77951_;
wire _77952_;
wire _77953_;
wire _77954_;
wire _77955_;
wire _77956_;
wire _77957_;
wire _77958_;
wire _77959_;
wire _77960_;
wire _77961_;
wire _77962_;
wire _77963_;
wire _77964_;
wire _77965_;
wire _77966_;
wire _77967_;
wire _77968_;
wire _77969_;
wire _77970_;
wire _77971_;
wire _77972_;
wire _77973_;
wire _77974_;
wire _77975_;
wire _77976_;
wire _77977_;
wire _77978_;
wire _77979_;
wire _77980_;
wire _77981_;
wire _77982_;
wire _77983_;
wire _77984_;
wire _77985_;
wire _77986_;
wire _77987_;
wire _77988_;
wire _77989_;
wire _77990_;
wire _77991_;
wire _77992_;
wire _77993_;
wire _77994_;
wire _77995_;
wire _77996_;
wire _77997_;
wire _77998_;
wire _77999_;
wire _78000_;
wire _78001_;
wire _78002_;
wire _78003_;
wire _78004_;
wire _78005_;
wire _78006_;
wire _78007_;
wire _78008_;
wire _78009_;
wire _78010_;
wire _78011_;
wire _78012_;
wire _78013_;
wire _78014_;
wire _78015_;
wire _78016_;
wire _78017_;
wire _78018_;
wire _78019_;
wire _78020_;
wire _78021_;
wire _78022_;
wire _78023_;
wire _78024_;
wire _78025_;
wire _78026_;
wire _78027_;
wire _78028_;
wire _78029_;
wire _78030_;
wire _78031_;
wire _78032_;
wire _78033_;
wire _78034_;
wire _78035_;
wire _78036_;
wire _78037_;
wire _78038_;
wire _78039_;
wire _78040_;
wire _78041_;
wire _78042_;
wire _78043_;
wire _78044_;
wire _78045_;
wire _78046_;
wire _78047_;
wire _78048_;
wire _78049_;
wire _78050_;
wire _78051_;
wire _78052_;
wire _78053_;
wire _78054_;
wire _78055_;
wire _78056_;
wire _78057_;
wire _78058_;
wire _78059_;
wire _78060_;
wire _78061_;
wire _78062_;
wire _78063_;
wire _78064_;
wire _78065_;
wire _78066_;
wire _78067_;
wire _78068_;
wire _78069_;
wire _78070_;
wire _78071_;
wire _78072_;
wire _78073_;
wire _78074_;
wire _78075_;
wire _78076_;
wire _78077_;
wire _78078_;
wire _78079_;
wire _78080_;
wire _78081_;
wire _78082_;
wire _78083_;
wire _78084_;
wire _78085_;
wire _78086_;
wire _78087_;
wire _78088_;
wire _78089_;
wire _78090_;
wire _78091_;
wire _78092_;
wire _78093_;
wire _78094_;
wire _78095_;
wire _78096_;
wire _78097_;
wire _78098_;
wire _78099_;
wire _78100_;
wire _78101_;
wire _78102_;
wire _78103_;
wire _78104_;
wire _78105_;
wire _78106_;
wire _78107_;
wire _78108_;
wire _78109_;
wire _78110_;
wire _78111_;
wire _78112_;
wire _78113_;
wire _78114_;
wire _78115_;
wire _78116_;
wire _78117_;
wire _78118_;
wire _78119_;
wire _78120_;
wire _78121_;
wire _78122_;
wire _78123_;
wire _78124_;
wire _78125_;
wire _78126_;
wire _78127_;
wire _78128_;
wire _78129_;
wire _78130_;
wire _78131_;
wire _78132_;
wire _78133_;
wire _78134_;
wire _78135_;
wire _78136_;
wire _78137_;
wire _78138_;
wire _78139_;
wire _78140_;
wire _78141_;
wire _78142_;
wire _78143_;
wire _78144_;
wire _78145_;
wire _78146_;
wire _78147_;
wire _78148_;
wire _78149_;
wire _78150_;
wire _78151_;
wire _78152_;
wire _78153_;
wire _78154_;
wire _78155_;
wire _78156_;
wire _78157_;
wire _78158_;
wire _78159_;
wire _78160_;
wire _78161_;
wire _78162_;
wire _78163_;
wire _78164_;
wire _78165_;
wire _78166_;
wire _78167_;
wire _78168_;
wire _78169_;
wire _78170_;
wire _78171_;
wire _78172_;
wire _78173_;
wire _78174_;
wire _78175_;
wire _78176_;
wire _78177_;
wire _78178_;
wire _78179_;
wire _78180_;
wire _78181_;
wire _78182_;
wire _78183_;
wire _78184_;
wire _78185_;
wire _78186_;
wire _78187_;
wire _78188_;
wire _78189_;
wire _78190_;
wire _78191_;
wire _78192_;
wire _78193_;
wire _78194_;
wire _78195_;
wire _78196_;
wire _78197_;
wire _78198_;
wire _78199_;
wire _78200_;
wire _78201_;
wire _78202_;
wire _78203_;
wire _78204_;
wire _78205_;
wire _78206_;
wire _78207_;
wire _78208_;
wire _78209_;
wire _78210_;
wire _78211_;
wire _78212_;
wire _78213_;
wire _78214_;
wire _78215_;
wire _78216_;
wire _78217_;
wire _78218_;
wire _78219_;
wire _78220_;
wire _78221_;
wire _78222_;
wire _78223_;
wire _78224_;
wire _78225_;
wire _78226_;
wire _78227_;
wire _78228_;
wire _78229_;
wire _78230_;
wire _78231_;
wire _78232_;
wire _78233_;
wire _78234_;
wire _78235_;
wire _78236_;
wire _78237_;
wire _78238_;
wire _78239_;
wire _78240_;
wire _78241_;
wire _78242_;
wire _78243_;
wire _78244_;
wire _78245_;
wire _78246_;
wire _78247_;
wire _78248_;
wire _78249_;
wire _78250_;
wire _78251_;
wire _78252_;
wire _78253_;
wire _78254_;
wire _78255_;
wire _78256_;
wire _78257_;
wire _78258_;
wire _78259_;
wire _78260_;
wire _78261_;
wire _78262_;
wire _78263_;
wire _78264_;
wire _78265_;
wire _78266_;
wire _78267_;
wire _78268_;
wire _78269_;
wire _78270_;
wire _78271_;
wire _78272_;
wire _78273_;
wire _78274_;
wire _78275_;
wire _78276_;
wire _78277_;
wire _78278_;
wire _78279_;
wire _78280_;
wire _78281_;
wire _78282_;
wire _78283_;
wire _78284_;
wire _78285_;
wire _78286_;
wire _78287_;
wire _78288_;
wire _78289_;
wire _78290_;
wire _78291_;
wire _78292_;
wire _78293_;
wire _78294_;
wire _78295_;
wire _78296_;
wire _78297_;
wire _78298_;
wire _78299_;
wire _78300_;
wire _78301_;
wire _78302_;
wire _78303_;
wire _78304_;
wire _78305_;
wire _78306_;
wire _78307_;
wire _78308_;
wire _78309_;
wire _78310_;
wire _78311_;
wire _78312_;
wire _78313_;
wire _78314_;
wire _78315_;
wire _78316_;
wire _78317_;
wire _78318_;
wire _78319_;
wire _78320_;
wire _78321_;
wire _78322_;
wire _78323_;
wire _78324_;
wire _78325_;
wire _78326_;
wire _78327_;
wire _78328_;
wire _78329_;
wire _78330_;
wire _78331_;
wire _78332_;
wire _78333_;
wire _78334_;
wire _78335_;
wire _78336_;
wire _78337_;
wire _78338_;
wire _78339_;
wire _78340_;
wire _78341_;
wire _78342_;
wire _78343_;
wire _78344_;
wire _78345_;
wire _78346_;
wire _78347_;
wire _78348_;
wire _78349_;
wire _78350_;
wire _78351_;
wire _78352_;
wire _78353_;
wire _78354_;
wire _78355_;
wire _78356_;
wire _78357_;
wire _78358_;
wire _78359_;
wire _78360_;
wire _78361_;
wire _78362_;
wire _78363_;
wire _78364_;
wire _78365_;
wire _78366_;
wire _78367_;
wire _78368_;
wire _78369_;
wire _78370_;
wire _78371_;
wire _78372_;
wire _78373_;
wire _78374_;
wire _78375_;
wire _78376_;
wire _78377_;
wire _78378_;
wire _78379_;
wire _78380_;
wire _78381_;
wire _78382_;
wire _78383_;
wire _78384_;
wire _78385_;
wire _78386_;
wire _78387_;
wire _78388_;
wire _78389_;
wire _78390_;
wire _78391_;
wire _78392_;
wire _78393_;
wire _78394_;
wire _78395_;
wire _78396_;
wire _78397_;
wire _78398_;
wire _78399_;
wire _78400_;
wire _78401_;
wire _78402_;
wire _78403_;
wire _78404_;
wire _78405_;
wire _78406_;
wire _78407_;
wire _78408_;
wire _78409_;
wire _78410_;
wire _78411_;
wire _78412_;
wire _78413_;
wire _78414_;
wire _78415_;
wire _78416_;
wire _78417_;
wire _78418_;
wire _78419_;
wire _78420_;
wire _78421_;
wire _78422_;
wire _78423_;
wire _78424_;
wire _78425_;
wire _78426_;
wire _78427_;
wire _78428_;
wire _78429_;
wire _78430_;
wire _78431_;
wire _78432_;
wire _78433_;
wire _78434_;
wire _78435_;
wire _78436_;
wire _78437_;
wire _78438_;
wire _78439_;
wire _78440_;
wire _78441_;
wire _78442_;
wire _78443_;
wire _78444_;
wire _78445_;
wire _78446_;
wire _78447_;
wire _78448_;
wire _78449_;
wire _78450_;
wire _78451_;
wire _78452_;
wire _78453_;
wire _78454_;
wire _78455_;
wire _78456_;
wire _78457_;
wire _78458_;
wire _78459_;
wire _78460_;
wire _78461_;
wire _78462_;
wire _78463_;
wire _78464_;
wire _78465_;
wire _78466_;
wire _78467_;
wire _78468_;
wire _78469_;
wire _78470_;
wire _78471_;
wire _78472_;
wire _78473_;
wire _78474_;
wire _78475_;
wire _78476_;
wire _78477_;
wire _78478_;
wire _78479_;
wire _78480_;
wire _78481_;
wire _78482_;
wire _78483_;
wire _78484_;
wire _78485_;
wire _78486_;
wire _78487_;
wire _78488_;
wire _78489_;
wire _78490_;
wire _78491_;
wire _78492_;
wire _78493_;
wire _78494_;
wire _78495_;
wire _78496_;
wire _78497_;
wire _78498_;
wire _78499_;
wire _78500_;
wire _78501_;
wire _78502_;
wire _78503_;
wire _78504_;
wire _78505_;
wire _78506_;
wire _78507_;
wire _78508_;
wire _78509_;
wire _78510_;
wire _78511_;
wire _78512_;
wire _78513_;
wire _78514_;
wire _78515_;
wire _78516_;
wire _78517_;
wire _78518_;
wire _78519_;
wire _78520_;
wire _78521_;
wire _78522_;
wire _78523_;
wire _78524_;
wire _78525_;
wire _78526_;
wire _78527_;
wire _78528_;
wire _78529_;
wire _78530_;
wire _78531_;
wire _78532_;
wire _78533_;
wire _78534_;
wire _78535_;
wire _78536_;
wire _78537_;
wire _78538_;
wire _78539_;
wire _78540_;
wire _78541_;
wire _78542_;
wire _78543_;
wire _78544_;
wire _78545_;
wire _78546_;
wire _78547_;
wire _78548_;
wire _78549_;
wire _78550_;
wire _78551_;
wire _78552_;
wire _78553_;
wire _78554_;
wire _78555_;
wire _78556_;
wire _78557_;
wire _78558_;
wire _78559_;
wire _78560_;
wire _78561_;
wire _78562_;
wire _78563_;
wire _78564_;
wire _78565_;
wire _78566_;
wire _78567_;
wire _78568_;
wire _78569_;
wire _78570_;
wire _78571_;
wire _78572_;
wire _78573_;
wire _78574_;
wire _78575_;
wire _78576_;
wire _78577_;
wire _78578_;
wire _78579_;
wire _78580_;
wire _78581_;
wire _78582_;
wire _78583_;
wire _78584_;
wire _78585_;
wire _78586_;
wire _78587_;
wire _78588_;
wire _78589_;
wire _78590_;
wire _78591_;
wire _78592_;
wire _78593_;
wire _78594_;
wire _78595_;
wire _78596_;
wire _78597_;
wire _78598_;
wire _78599_;
wire _78600_;
wire _78601_;
wire _78602_;
wire _78603_;
wire _78604_;
wire _78605_;
wire _78606_;
wire _78607_;
wire _78608_;
wire _78609_;
wire _78610_;
wire _78611_;
wire _78612_;
wire _78613_;
wire _78614_;
wire _78615_;
wire _78616_;
wire _78617_;
wire _78618_;
wire _78619_;
wire _78620_;
wire _78621_;
wire _78622_;
wire _78623_;
wire _78624_;
wire _78625_;
wire _78626_;
wire _78627_;
wire _78628_;
wire _78629_;
wire _78630_;
wire _78631_;
wire _78632_;
wire _78633_;
wire _78634_;
wire _78635_;
wire _78636_;
wire _78637_;
wire _78638_;
wire _78639_;
wire _78640_;
wire _78641_;
wire _78642_;
wire _78643_;
wire _78644_;
wire _78645_;
wire _78646_;
wire _78647_;
wire _78648_;
wire _78649_;
wire _78650_;
wire _78651_;
wire _78652_;
wire _78653_;
wire _78654_;
wire _78655_;
wire _78656_;
wire _78657_;
wire _78658_;
wire _78659_;
wire _78660_;
wire _78661_;
wire _78662_;
wire _78663_;
wire _78664_;
wire _78665_;
wire _78666_;
wire _78667_;
wire _78668_;
wire _78669_;
wire _78670_;
wire _78671_;
wire _78672_;
wire _78673_;
wire _78674_;
wire _78675_;
wire _78676_;
wire _78677_;
wire _78678_;
wire _78679_;
wire _78680_;
wire _78681_;
wire _78682_;
wire _78683_;
wire _78684_;
wire _78685_;
wire _78686_;
wire _78687_;
wire _78688_;
wire _78689_;
wire _78690_;
wire _78691_;
wire _78692_;
wire _78693_;
wire _78694_;
wire _78695_;
wire _78696_;
wire _78697_;
wire _78698_;
wire _78699_;
wire _78700_;
wire _78701_;
wire _78702_;
wire _78703_;
wire _78704_;
wire _78705_;
wire _78706_;
wire _78707_;
wire _78708_;
wire _78709_;
wire _78710_;
wire _78711_;
wire _78712_;
wire _78713_;
wire _78714_;
wire _78715_;
wire _78716_;
wire _78717_;
wire _78718_;
wire _78719_;
wire _78720_;
wire _78721_;
wire _78722_;
wire _78723_;
wire _78724_;
wire _78725_;
wire _78726_;
wire _78727_;
wire _78728_;
wire _78729_;
wire _78730_;
wire _78731_;
wire _78732_;
wire _78733_;
wire _78734_;
wire _78735_;
wire _78736_;
wire _78737_;
wire _78738_;
wire _78739_;
wire _78740_;
wire _78741_;
wire _78742_;
wire _78743_;
wire _78744_;
wire _78745_;
wire _78746_;
wire _78747_;
wire _78748_;
wire _78749_;
wire _78750_;
wire _78751_;
wire _78752_;
wire _78753_;
wire _78754_;
wire _78755_;
wire _78756_;
wire _78757_;
wire _78758_;
wire _78759_;
wire _78760_;
wire _78761_;
wire _78762_;
wire _78763_;
wire _78764_;
wire _78765_;
wire _78766_;
wire _78767_;
wire _78768_;
wire _78769_;
wire _78770_;
wire _78771_;
wire _78772_;
wire _78773_;
wire _78774_;
wire _78775_;
wire _78776_;
wire _78777_;
wire _78778_;
wire _78779_;
wire _78780_;
wire _78781_;
wire _78782_;
wire _78783_;
wire _78784_;
wire _78785_;
wire _78786_;
wire _78787_;
wire _78788_;
wire _78789_;
wire _78790_;
wire _78791_;
wire _78792_;
wire _78793_;
wire _78794_;
wire _78795_;
wire _78796_;
wire _78797_;
wire _78798_;
wire _78799_;
wire _78800_;
wire _78801_;
wire _78802_;
wire _78803_;
wire _78804_;
wire _78805_;
wire _78806_;
wire _78807_;
wire _78808_;
wire _78809_;
wire _78810_;
wire _78811_;
wire _78812_;
wire _78813_;
wire _78814_;
wire _78815_;
wire _78816_;
wire _78817_;
wire _78818_;
wire _78819_;
wire _78820_;
wire _78821_;
wire _78822_;
wire _78823_;
wire _78824_;
wire _78825_;
wire _78826_;
wire _78827_;
wire _78828_;
wire _78829_;
wire _78830_;
wire _78831_;
wire _78832_;
wire _78833_;
wire _78834_;
wire _78835_;
wire _78836_;
wire _78837_;
wire _78838_;
wire _78839_;
wire _78840_;
wire _78841_;
wire _78842_;
wire _78843_;
wire _78844_;
wire _78845_;
wire _78846_;
wire _78847_;
wire _78848_;
wire _78849_;
wire _78850_;
wire _78851_;
wire _78852_;
wire _78853_;
wire _78854_;
wire _78855_;
wire _78856_;
wire _78857_;
wire _78858_;
wire _78859_;
wire _78860_;
wire _78861_;
wire _78862_;
wire _78863_;
wire _78864_;
wire _78865_;
wire _78866_;
wire _78867_;
wire _78868_;
wire _78869_;
wire _78870_;
wire _78871_;
wire _78872_;
wire _78873_;
wire _78874_;
wire _78875_;
wire _78876_;
wire _78877_;
wire _78878_;
wire _78879_;
wire _78880_;
wire _78881_;
wire _78882_;
wire _78883_;
wire _78884_;
wire _78885_;
wire _78886_;
wire _78887_;
wire _78888_;
wire _78889_;
wire _78890_;
wire _78891_;
wire _78892_;
wire _78893_;
wire _78894_;
wire _78895_;
wire _78896_;
wire _78897_;
wire _78898_;
wire _78899_;
wire _78900_;
wire _78901_;
wire _78902_;
wire _78903_;
wire _78904_;
wire _78905_;
wire _78906_;
wire _78907_;
wire _78908_;
wire _78909_;
wire _78910_;
wire _78911_;
wire _78912_;
wire _78913_;
wire _78914_;
wire _78915_;
wire _78916_;
wire _78917_;
wire _78918_;
wire _78919_;
wire _78920_;
wire _78921_;
wire _78922_;
wire _78923_;
wire _78924_;
wire _78925_;
wire _78926_;
wire _78927_;
wire _78928_;
wire _78929_;
wire _78930_;
wire _78931_;
wire _78932_;
wire _78933_;
wire _78934_;
wire _78935_;
wire _78936_;
wire _78937_;
wire _78938_;
wire _78939_;
wire _78940_;
wire _78941_;
wire _78942_;
wire _78943_;
wire _78944_;
wire _78945_;
wire _78946_;
wire _78947_;
wire _78948_;
wire _78949_;
wire _78950_;
wire _78951_;
wire _78952_;
wire _78953_;
wire _78954_;
wire _78955_;
wire _78956_;
wire _78957_;
wire _78958_;
wire _78959_;
wire _78960_;
wire _78961_;
wire _78962_;
wire _78963_;
wire _78964_;
wire _78965_;
wire _78966_;
wire _78967_;
wire _78968_;
wire _78969_;
wire _78970_;
wire _78971_;
wire _78972_;
wire _78973_;
wire _78974_;
wire _78975_;
wire _78976_;
wire _78977_;
wire _78978_;
wire _78979_;
wire _78980_;
wire _78981_;
wire _78982_;
wire _78983_;
wire _78984_;
wire _78985_;
wire _78986_;
wire _78987_;
wire _78988_;
wire _78989_;
wire _78990_;
wire _78991_;
wire _78992_;
wire _78993_;
wire _78994_;
wire _78995_;
wire _78996_;
wire _78997_;
wire _78998_;
wire _78999_;
wire _79000_;
wire _79001_;
wire _79002_;
wire _79003_;
wire _79004_;
wire _79005_;
wire _79006_;
wire _79007_;
wire _79008_;
wire _79009_;
wire _79010_;
wire _79011_;
wire _79012_;
wire _79013_;
wire _79014_;
wire _79015_;
wire _79016_;
wire _79017_;
wire _79018_;
wire _79019_;
wire _79020_;
wire _79021_;
wire _79022_;
wire _79023_;
wire _79024_;
wire _79025_;
wire _79026_;
wire _79027_;
wire _79028_;
wire _79029_;
wire _79030_;
wire _79031_;
wire _79032_;
wire _79033_;
wire _79034_;
wire _79035_;
wire _79036_;
wire _79037_;
wire _79038_;
wire _79039_;
wire _79040_;
wire _79041_;
wire _79042_;
wire _79043_;
wire _79044_;
wire _79045_;
wire _79046_;
wire _79047_;
wire _79048_;
wire _79049_;
wire _79050_;
wire _79051_;
wire _79052_;
wire _79053_;
wire _79054_;
wire _79055_;
wire _79056_;
wire _79057_;
wire _79058_;
wire _79059_;
wire _79060_;
wire _79061_;
wire _79062_;
wire _79063_;
wire _79064_;
wire _79065_;
wire _79066_;
wire _79067_;
wire _79068_;
wire _79069_;
wire _79070_;
wire _79071_;
wire _79072_;
wire _79073_;
wire _79074_;
wire _79075_;
wire _79076_;
wire _79077_;
wire _79078_;
wire _79079_;
wire _79080_;
wire _79081_;
wire _79082_;
wire _79083_;
wire _79084_;
wire _79085_;
wire _79086_;
wire _79087_;
wire _79088_;
wire _79089_;
wire _79090_;
wire _79091_;
wire _79092_;
wire _79093_;
wire _79094_;
wire _79095_;
wire _79096_;
wire _79097_;
wire _79098_;
wire _79099_;
wire _79100_;
wire _79101_;
wire _79102_;
wire _79103_;
wire _79104_;
wire _79105_;
wire _79106_;
wire _79107_;
wire _79108_;
wire _79109_;
wire _79110_;
wire _79111_;
wire _79112_;
wire _79113_;
wire _79114_;
wire _79115_;
wire _79116_;
wire _79117_;
wire _79118_;
wire _79119_;
wire _79120_;
wire _79121_;
wire _79122_;
wire _79123_;
wire _79124_;
wire _79125_;
wire _79126_;
wire _79127_;
wire _79128_;
wire _79129_;
wire _79130_;
wire _79131_;
wire _79132_;
wire _79133_;
wire _79134_;
wire _79135_;
wire _79136_;
wire _79137_;
wire _79138_;
wire _79139_;
wire _79140_;
wire _79141_;
wire _79142_;
wire _79143_;
wire _79144_;
wire _79145_;
wire _79146_;
wire _79147_;
wire _79148_;
wire _79149_;
wire _79150_;
wire _79151_;
wire _79152_;
wire _79153_;
wire _79154_;
wire _79155_;
wire _79156_;
wire _79157_;
wire _79158_;
wire _79159_;
wire _79160_;
wire _79161_;
wire _79162_;
wire _79163_;
wire _79164_;
wire _79165_;
wire _79166_;
wire _79167_;
wire _79168_;
wire _79169_;
wire _79170_;
wire _79171_;
wire _79172_;
wire _79173_;
wire _79174_;
wire _79175_;
wire _79176_;
wire _79177_;
wire _79178_;
wire _79179_;
wire _79180_;
wire _79181_;
wire _79182_;
wire _79183_;
wire _79184_;
wire _79185_;
wire _79186_;
wire _79187_;
wire _79188_;
wire _79189_;
wire _79190_;
wire _79191_;
wire _79192_;
wire _79193_;
wire _79194_;
wire _79195_;
wire _79196_;
wire _79197_;
wire _79198_;
wire _79199_;
wire _79200_;
wire _79201_;
wire _79202_;
wire _79203_;
wire _79204_;
wire _79205_;
wire _79206_;
wire _79207_;
wire _79208_;
wire _79209_;
wire _79210_;
wire _79211_;
wire _79212_;
wire _79213_;
wire _79214_;
wire _79215_;
wire _79216_;
wire _79217_;
wire _79218_;
wire _79219_;
wire _79220_;
wire _79221_;
wire _79222_;
wire _79223_;
wire _79224_;
wire _79225_;
wire _79226_;
wire _79227_;
wire _79228_;
wire _79229_;
wire _79230_;
wire _79231_;
wire _79232_;
wire _79233_;
wire _79234_;
wire _79235_;
wire _79236_;
wire _79237_;
wire _79238_;
wire _79239_;
wire _79240_;
wire _79241_;
wire _79242_;
wire _79243_;
wire _79244_;
wire _79245_;
wire _79246_;
wire _79247_;
wire _79248_;
wire _79249_;
wire _79250_;
wire _79251_;
wire _79252_;
wire _79253_;
wire _79254_;
wire _79255_;
wire _79256_;
wire _79257_;
wire _79258_;
wire _79259_;
wire _79260_;
wire _79261_;
wire _79262_;
wire _79263_;
wire _79264_;
wire _79265_;
wire _79266_;
wire _79267_;
wire _79268_;
wire _79269_;
wire _79270_;
wire _79271_;
wire _79272_;
wire _79273_;
wire _79274_;
wire _79275_;
wire _79276_;
wire _79277_;
wire _79278_;
wire _79279_;
wire _79280_;
wire _79281_;
wire _79282_;
wire _79283_;
wire _79284_;
wire _79285_;
wire _79286_;
wire _79287_;
wire _79288_;
wire _79289_;
wire _79290_;
wire _79291_;
wire _79292_;
wire _79293_;
wire _79294_;
wire _79295_;
wire _79296_;
wire _79297_;
wire _79298_;
wire _79299_;
wire _79300_;
wire _79301_;
wire _79302_;
wire _79303_;
wire _79304_;
wire _79305_;
wire _79306_;
wire _79307_;
wire _79308_;
wire _79309_;
wire _79310_;
wire _79311_;
wire _79312_;
wire _79313_;
wire _79314_;
wire _79315_;
wire _79316_;
wire _79317_;
wire _79318_;
wire _79319_;
wire _79320_;
wire _79321_;
wire _79322_;
wire _79323_;
wire _79324_;
wire _79325_;
wire _79326_;
wire _79327_;
wire _79328_;
wire _79329_;
wire _79330_;
wire _79331_;
wire _79332_;
wire _79333_;
wire _79334_;
wire _79335_;
wire _79336_;
wire _79337_;
wire _79338_;
wire _79339_;
wire _79340_;
wire _79341_;
wire _79342_;
wire _79343_;
wire _79344_;
wire _79345_;
wire _79346_;
wire _79347_;
wire _79348_;
wire _79349_;
wire _79350_;
wire _79351_;
wire _79352_;
wire _79353_;
wire _79354_;
wire _79355_;
wire _79356_;
wire _79357_;
wire _79358_;
wire _79359_;
wire _79360_;
wire _79361_;
wire _79362_;
wire _79363_;
wire _79364_;
wire _79365_;
wire _79366_;
wire _79367_;
wire _79368_;
wire _79369_;
wire _79370_;
wire _79371_;
wire _79372_;
wire _79373_;
wire _79374_;
wire _79375_;
wire _79376_;
wire _79377_;
wire _79378_;
wire _79379_;
wire _79380_;
wire _79381_;
wire _79382_;
wire _79383_;
wire _79384_;
wire _79385_;
wire _79386_;
wire _79387_;
wire _79388_;
wire _79389_;
wire _79390_;
wire _79391_;
wire _79392_;
wire _79393_;
wire _79394_;
wire _79395_;
wire _79396_;
wire _79397_;
wire _79398_;
wire _79399_;
wire _79400_;
wire _79401_;
wire _79402_;
wire _79403_;
wire _79404_;
wire _79405_;
wire _79406_;
wire _79407_;
wire _79408_;
wire _79409_;
wire _79410_;
wire _79411_;
wire _79412_;
wire _79413_;
wire _79414_;
wire _79415_;
wire _79416_;
wire _79417_;
wire _79418_;
wire _79419_;
wire _79420_;
wire _79421_;
wire _79422_;
wire _79423_;
wire _79424_;
wire _79425_;
wire _79426_;
wire _79427_;
wire _79428_;
wire _79429_;
wire _79430_;
wire _79431_;
wire _79432_;
wire _79433_;
wire _79434_;
wire _79435_;
wire _79436_;
wire _79437_;
wire _79438_;
wire _79439_;
wire _79440_;
wire _79441_;
wire _79442_;
wire _79443_;
wire _79444_;
wire _79445_;
wire _79446_;
wire _79447_;
wire _79448_;
wire _79449_;
wire _79450_;
wire _79451_;
wire _79452_;
wire _79453_;
wire _79454_;
wire _79455_;
wire _79456_;
wire _79457_;
wire _79458_;
wire _79459_;
wire _79460_;
wire _79461_;
wire _79462_;
wire _79463_;
wire _79464_;
wire _79465_;
wire _79466_;
wire _79467_;
wire _79468_;
wire _79469_;
wire _79470_;
wire _79471_;
wire _79472_;
wire _79473_;
wire _79474_;
wire _79475_;
wire _79476_;
wire _79477_;
wire _79478_;
wire _79479_;
wire _79480_;
wire _79481_;
wire _79482_;
wire _79483_;
wire _79484_;
wire _79485_;
wire _79486_;
wire _79487_;
wire _79488_;
wire _79489_;
wire _79490_;
wire _79491_;
wire _79492_;
wire _79493_;
wire _79494_;
wire _79495_;
wire _79496_;
wire _79497_;
wire _79498_;
wire _79499_;
wire _79500_;
wire _79501_;
wire _79502_;
wire _79503_;
wire _79504_;
wire _79505_;
wire _79506_;
wire _79507_;
wire _79508_;
wire _79509_;
wire _79510_;
wire _79511_;
wire _79512_;
wire _79513_;
wire _79514_;
wire _79515_;
wire _79516_;
wire _79517_;
wire _79518_;
wire _79519_;
wire _79520_;
wire _79521_;
wire _79522_;
wire _79523_;
wire _79524_;
wire _79525_;
wire _79526_;
wire _79527_;
wire _79528_;
wire _79529_;
wire _79530_;
wire _79531_;
wire _79532_;
wire _79533_;
wire _79534_;
wire _79535_;
wire _79536_;
wire _79537_;
wire _79538_;
wire _79539_;
wire _79540_;
wire _79541_;
wire _79542_;
wire _79543_;
wire _79544_;
wire _79545_;
wire _79546_;
wire _79547_;
wire _79548_;
wire _79549_;
wire _79550_;
wire _79551_;
wire _79552_;
wire _79553_;
wire _79554_;
wire _79555_;
wire _79556_;
wire _79557_;
wire _79558_;
wire _79559_;
wire _79560_;
wire _79561_;
wire _79562_;
wire _79563_;
wire _79564_;
wire _79565_;
wire _79566_;
wire _79567_;
wire _79568_;
wire _79569_;
wire _79570_;
wire _79571_;
wire _79572_;
wire _79573_;
wire _79574_;
wire _79575_;
wire _79576_;
wire _79577_;
wire _79578_;
wire _79579_;
wire _79580_;
wire _79581_;
wire _79582_;
wire _79583_;
wire _79584_;
wire _79585_;
wire _79586_;
wire _79587_;
wire _79588_;
wire _79589_;
wire _79590_;
wire _79591_;
wire _79592_;
wire _79593_;
wire _79594_;
wire _79595_;
wire _79596_;
wire _79597_;
wire _79598_;
wire _79599_;
wire _79600_;
wire _79601_;
wire _79602_;
wire _79603_;
wire _79604_;
wire _79605_;
wire _79606_;
wire _79607_;
wire _79608_;
wire _79609_;
wire _79610_;
wire _79611_;
wire _79612_;
wire _79613_;
wire _79614_;
wire _79615_;
wire _79616_;
wire _79617_;
wire _79618_;
wire _79619_;
wire _79620_;
wire _79621_;
wire _79622_;
wire _79623_;
wire _79624_;
wire _79625_;
wire _79626_;
wire _79627_;
wire _79628_;
wire _79629_;
wire _79630_;
wire _79631_;
wire _79632_;
wire _79633_;
wire _79634_;
wire _79635_;
wire _79636_;
wire _79637_;
wire _79638_;
wire _79639_;
wire _79640_;
wire _79641_;
wire _79642_;
wire _79643_;
wire _79644_;
wire _79645_;
wire _79646_;
wire _79647_;
wire _79648_;
wire _79649_;
wire _79650_;
wire _79651_;
wire _79652_;
wire _79653_;
wire _79654_;
wire _79655_;
wire _79656_;
wire _79657_;
wire _79658_;
wire _79659_;
wire _79660_;
wire _79661_;
wire _79662_;
wire _79663_;
wire _79664_;
wire _79665_;
wire _79666_;
wire _79667_;
wire _79668_;
wire _79669_;
wire _79670_;
wire _79671_;
wire _79672_;
wire _79673_;
wire _79674_;
wire _79675_;
wire _79676_;
wire _79677_;
wire _79678_;
wire _79679_;
wire _79680_;
wire _79681_;
wire _79682_;
wire _79683_;
wire _79684_;
wire _79685_;
wire _79686_;
wire _79687_;
wire _79688_;
wire _79689_;
wire _79690_;
wire _79691_;
wire _79692_;
wire _79693_;
wire _79694_;
wire _79695_;
wire _79696_;
wire _79697_;
wire _79698_;
wire _79699_;
wire _79700_;
wire _79701_;
wire _79702_;
wire _79703_;
wire _79704_;
wire _79705_;
wire _79706_;
wire _79707_;
wire _79708_;
wire _79709_;
wire _79710_;
wire _79711_;
wire _79712_;
wire _79713_;
wire _79714_;
wire _79715_;
wire _79716_;
wire _79717_;
wire _79718_;
wire _79719_;
wire _79720_;
wire _79721_;
wire _79722_;
wire _79723_;
wire _79724_;
wire _79725_;
wire _79726_;
wire _79727_;
wire _79728_;
wire _79729_;
wire _79730_;
wire _79731_;
wire _79732_;
wire _79733_;
wire _79734_;
wire _79735_;
wire _79736_;
wire _79737_;
wire _79738_;
wire _79739_;
wire _79740_;
wire _79741_;
wire _79742_;
wire _79743_;
wire _79744_;
wire _79745_;
wire _79746_;
wire _79747_;
wire _79748_;
wire _79749_;
wire _79750_;
wire _79751_;
wire _79752_;
wire _79753_;
wire _79754_;
wire _79755_;
wire _79756_;
wire _79757_;
wire _79758_;
wire _79759_;
wire _79760_;
wire _79761_;
wire _79762_;
wire _79763_;
wire _79764_;
wire _79765_;
wire _79766_;
wire _79767_;
wire _79768_;
wire _79769_;
wire _79770_;
wire _79771_;
wire _79772_;
wire _79773_;
wire _79774_;
wire _79775_;
wire _79776_;
wire _79777_;
wire _79778_;
wire _79779_;
wire _79780_;
wire _79781_;
wire _79782_;
wire _79783_;
wire _79784_;
wire _79785_;
wire _79786_;
wire _79787_;
wire _79788_;
wire _79789_;
wire _79790_;
wire _79791_;
wire _79792_;
wire _79793_;
wire _79794_;
wire _79795_;
wire _79796_;
wire _79797_;
wire _79798_;
wire _79799_;
wire _79800_;
wire _79801_;
wire _79802_;
wire _79803_;
wire _79804_;
wire _79805_;
wire _79806_;
wire _79807_;
wire _79808_;
wire _79809_;
wire _79810_;
wire _79811_;
wire _79812_;
wire _79813_;
wire _79814_;
wire _79815_;
wire _79816_;
wire _79817_;
wire _79818_;
wire _79819_;
wire _79820_;
wire _79821_;
wire _79822_;
wire _79823_;
wire _79824_;
wire _79825_;
wire _79826_;
wire _79827_;
wire _79828_;
wire _79829_;
wire _79830_;
wire _79831_;
wire _79832_;
wire _79833_;
wire _79834_;
wire _79835_;
wire _79836_;
wire _79837_;
wire _79838_;
wire _79839_;
wire _79840_;
wire _79841_;
wire _79842_;
wire _79843_;
wire _79844_;
wire _79845_;
wire _79846_;
wire _79847_;
wire _79848_;
wire _79849_;
wire _79850_;
wire _79851_;
wire _79852_;
wire _79853_;
wire _79854_;
wire _79855_;
wire _79856_;
wire _79857_;
wire _79858_;
wire _79859_;
wire _79860_;
wire _79861_;
wire _79862_;
wire _79863_;
wire _79864_;
wire _79865_;
wire _79866_;
wire _79867_;
wire _79868_;
wire _79869_;
wire _79870_;
wire _79871_;
wire _79872_;
wire _79873_;
wire _79874_;
wire _79875_;
wire _79876_;
wire _79877_;
wire _79878_;
wire _79879_;
wire _79880_;
wire _79881_;
wire _79882_;
wire _79883_;
wire _79884_;
wire _79885_;
wire _79886_;
wire _79887_;
wire _79888_;
wire _79889_;
wire _79890_;
wire _79891_;
wire _79892_;
wire _79893_;
wire _79894_;
wire _79895_;
wire _79896_;
wire _79897_;
wire _79898_;
wire _79899_;
wire _79900_;
wire _79901_;
wire _79902_;
wire _79903_;
wire _79904_;
wire _79905_;
wire _79906_;
wire _79907_;
wire _79908_;
wire _79909_;
wire _79910_;
wire _79911_;
wire _79912_;
wire _79913_;
wire _79914_;
wire _79915_;
wire _79916_;
wire _79917_;
wire _79918_;
wire _79919_;
wire _79920_;
wire _79921_;
wire _79922_;
wire _79923_;
wire _79924_;
wire _79925_;
wire _79926_;
wire _79927_;
wire _79928_;
wire _79929_;
wire _79930_;
wire _79931_;
wire _79932_;
wire _79933_;
wire _79934_;
wire _79935_;
wire _79936_;
wire _79937_;
wire _79938_;
wire _79939_;
wire _79940_;
wire _79941_;
wire _79942_;
wire _79943_;
wire _79944_;
wire _79945_;
wire _79946_;
wire _79947_;
wire _79948_;
wire _79949_;
wire _79950_;
wire _79951_;
wire _79952_;
wire _79953_;
wire _79954_;
wire _79955_;
wire _79956_;
wire _79957_;
wire _79958_;
wire _79959_;
wire _79960_;
wire _79961_;
wire _79962_;
wire _79963_;
wire _79964_;
wire _79965_;
wire _79966_;
wire _79967_;
wire _79968_;
wire _79969_;
wire _79970_;
wire _79971_;
wire _79972_;
wire _79973_;
wire _79974_;
wire _79975_;
wire _79976_;
wire _79977_;
wire _79978_;
wire _79979_;
wire _79980_;
wire _79981_;
wire _79982_;
wire _79983_;
wire _79984_;
wire _79985_;
wire _79986_;
wire _79987_;
wire _79988_;
wire _79989_;
wire _79990_;
wire _79991_;
wire _79992_;
wire _79993_;
wire _79994_;
wire _79995_;
wire _79996_;
wire _79997_;
wire _79998_;
wire _79999_;
wire _80000_;
wire _80001_;
wire _80002_;
wire _80003_;
wire _80004_;
wire _80005_;
wire _80006_;
wire _80007_;
wire _80008_;
wire _80009_;
wire _80010_;
wire _80011_;
wire _80012_;
wire _80013_;
wire _80014_;
wire _80015_;
wire _80016_;
wire _80017_;
wire _80018_;
wire _80019_;
wire _80020_;
wire _80021_;
wire _80022_;
wire _80023_;
wire _80024_;
wire _80025_;
wire _80026_;
wire _80027_;
wire _80028_;
wire _80029_;
wire _80030_;
wire _80031_;
wire _80032_;
wire _80033_;
wire _80034_;
wire _80035_;
wire _80036_;
wire _80037_;
wire _80038_;
wire _80039_;
wire _80040_;
wire _80041_;
wire _80042_;
wire _80043_;
wire _80044_;
wire _80045_;
wire _80046_;
wire _80047_;
wire _80048_;
wire _80049_;
wire _80050_;
wire _80051_;
wire _80052_;
wire _80053_;
wire _80054_;
wire _80055_;
wire _80056_;
wire _80057_;
wire _80058_;
wire _80059_;
wire _80060_;
wire _80061_;
wire _80062_;
wire _80063_;
wire _80064_;
wire _80065_;
wire _80066_;
wire _80067_;
wire _80068_;
wire _80069_;
wire _80070_;
wire _80071_;
wire _80072_;
wire _80073_;
wire _80074_;
wire _80075_;
wire _80076_;
wire _80077_;
wire _80078_;
wire _80079_;
wire _80080_;
wire _80081_;
wire _80082_;
wire _80083_;
wire _80084_;
wire _80085_;
wire _80086_;
wire _80087_;
wire _80088_;
wire _80089_;
wire _80090_;
wire _80091_;
wire _80092_;
wire _80093_;
wire _80094_;
wire _80095_;
wire _80096_;
wire _80097_;
wire _80098_;
wire _80099_;
wire _80100_;
wire _80101_;
wire _80102_;
wire _80103_;
wire _80104_;
wire _80105_;
wire _80106_;
wire _80107_;
wire _80108_;
wire _80109_;
wire _80110_;
wire _80111_;
wire _80112_;
wire _80113_;
wire _80114_;
wire _80115_;
wire _80116_;
wire _80117_;
wire _80118_;
wire _80119_;
wire _80120_;
wire _80121_;
wire _80122_;
wire _80123_;
wire _80124_;
wire _80125_;
wire _80126_;
wire _80127_;
wire _80128_;
wire _80129_;
wire _80130_;
wire _80131_;
wire _80132_;
wire _80133_;
wire _80134_;
wire _80135_;
wire _80136_;
wire _80137_;
wire _80138_;
wire _80139_;
wire _80140_;
wire _80141_;
wire _80142_;
wire _80143_;
wire _80144_;
wire _80145_;
wire _80146_;
wire _80147_;
wire _80148_;
wire _80149_;
wire _80150_;
wire _80151_;
wire _80152_;
wire _80153_;
wire _80154_;
wire _80155_;
wire _80156_;
wire _80157_;
wire _80158_;
wire _80159_;
wire _80160_;
wire _80161_;
wire _80162_;
wire _80163_;
wire _80164_;
wire _80165_;
wire _80166_;
wire _80167_;
wire _80168_;
wire _80169_;
wire _80170_;
wire _80171_;
wire _80172_;
wire _80173_;
wire _80174_;
wire _80175_;
wire _80176_;
wire _80177_;
wire _80178_;
wire _80179_;
wire _80180_;
wire _80181_;
wire _80182_;
wire _80183_;
wire _80184_;
wire _80185_;
wire _80186_;
wire _80187_;
wire _80188_;
wire _80189_;
wire _80190_;
wire _80191_;
wire _80192_;
wire _80193_;
wire _80194_;
wire _80195_;
wire _80196_;
wire _80197_;
wire _80198_;
wire _80199_;
wire _80200_;
wire _80201_;
wire _80202_;
wire _80203_;
wire _80204_;
wire _80205_;
wire _80206_;
wire _80207_;
wire _80208_;
wire _80209_;
wire _80210_;
wire _80211_;
wire _80212_;
wire _80213_;
wire _80214_;
wire _80215_;
wire _80216_;
wire _80217_;
wire _80218_;
wire _80219_;
wire _80220_;
wire _80221_;
wire _80222_;
wire _80223_;
wire _80224_;
wire _80225_;
wire _80226_;
wire _80227_;
wire _80228_;
wire _80229_;
wire _80230_;
wire _80231_;
wire _80232_;
wire _80233_;
wire _80234_;
wire _80235_;
wire _80236_;
wire _80237_;
wire _80238_;
wire _80239_;
wire _80240_;
wire _80241_;
wire _80242_;
wire _80243_;
wire _80244_;
wire _80245_;
wire _80246_;
wire _80247_;
wire _80248_;
wire _80249_;
wire _80250_;
wire _80251_;
wire _80252_;
wire _80253_;
wire _80254_;
wire _80255_;
wire _80256_;
wire _80257_;
wire _80258_;
wire _80259_;
wire _80260_;
wire _80261_;
wire _80262_;
wire _80263_;
wire _80264_;
wire _80265_;
wire _80266_;
wire _80267_;
wire _80268_;
wire _80269_;
wire _80270_;
wire _80271_;
wire _80272_;
wire _80273_;
wire _80274_;
wire _80275_;
wire _80276_;
wire _80277_;
wire _80278_;
wire _80279_;
wire _80280_;
wire _80281_;
wire _80282_;
wire _80283_;
wire _80284_;
wire _80285_;
wire _80286_;
wire _80287_;
wire _80288_;
wire _80289_;
wire _80290_;
wire _80291_;
wire _80292_;
wire _80293_;
wire _80294_;
wire _80295_;
wire _80296_;
wire _80297_;
wire _80298_;
wire _80299_;
wire _80300_;
wire _80301_;
wire _80302_;
wire _80303_;
wire _80304_;
wire _80305_;
wire _80306_;
wire _80307_;
wire _80308_;
wire _80309_;
wire _80310_;
wire _80311_;
wire _80312_;
wire _80313_;
wire _80314_;
wire _80315_;
wire _80316_;
wire _80317_;
wire _80318_;
wire _80319_;
wire _80320_;
wire _80321_;
wire _80322_;
wire _80323_;
wire _80324_;
wire _80325_;
wire _80326_;
wire _80327_;
wire _80328_;
wire _80329_;
wire _80330_;
wire _80331_;
wire _80332_;
wire _80333_;
wire _80334_;
wire _80335_;
wire _80336_;
wire _80337_;
wire _80338_;
wire _80339_;
wire _80340_;
wire _80341_;
wire _80342_;
wire _80343_;
wire _80344_;
wire _80345_;
wire _80346_;
wire _80347_;
wire _80348_;
wire _80349_;
wire _80350_;
wire _80351_;
wire _80352_;
wire _80353_;
wire _80354_;
wire _80355_;
wire _80356_;
wire _80357_;
wire _80358_;
wire _80359_;
wire _80360_;
wire _80361_;
wire _80362_;
wire _80363_;
wire _80364_;
wire _80365_;
wire _80366_;
wire _80367_;
wire _80368_;
wire _80369_;
wire _80370_;
wire _80371_;
wire _80372_;
wire _80373_;
wire _80374_;
wire _80375_;
wire _80376_;
wire _80377_;
wire _80378_;
wire _80379_;
wire _80380_;
wire _80381_;
wire _80382_;
wire _80383_;
wire _80384_;
wire _80385_;
wire _80386_;
wire _80387_;
wire _80388_;
wire _80389_;
wire _80390_;
wire _80391_;
wire _80392_;
wire _80393_;
wire _80394_;
wire _80395_;
wire _80396_;
wire _80397_;
wire _80398_;
wire _80399_;
wire _80400_;
wire _80401_;
wire _80402_;
wire _80403_;
wire _80404_;
wire _80405_;
wire _80406_;
wire _80407_;
wire _80408_;
wire _80409_;
wire _80410_;
wire _80411_;
wire _80412_;
wire _80413_;
wire _80414_;
wire _80415_;
wire _80416_;
wire _80417_;
wire _80418_;
wire _80419_;
wire _80420_;
wire _80421_;
wire _80422_;
wire _80423_;
wire _80424_;
wire _80425_;
wire _80426_;
wire _80427_;
wire _80428_;
wire _80429_;
wire _80430_;
wire _80431_;
wire _80432_;
wire _80433_;
wire _80434_;
wire _80435_;
wire _80436_;
wire _80437_;
wire _80438_;
wire _80439_;
wire _80440_;
wire _80441_;
wire _80442_;
wire _80443_;
wire _80444_;
wire _80445_;
wire _80446_;
wire _80447_;
wire _80448_;
wire _80449_;
wire _80450_;
wire _80451_;
wire _80452_;
wire _80453_;
wire _80454_;
wire _80455_;
wire _80456_;
wire _80457_;
wire _80458_;
wire _80459_;
wire _80460_;
wire _80461_;
wire _80462_;
wire _80463_;
wire _80464_;
wire _80465_;
wire _80466_;
wire _80467_;
wire _80468_;
wire _80469_;
wire _80470_;
wire _80471_;
wire _80472_;
wire _80473_;
wire _80474_;
wire _80475_;
wire _80476_;
wire _80477_;
wire _80478_;
wire _80479_;
wire _80480_;
wire _80481_;
wire _80482_;
wire _80483_;
wire _80484_;
wire _80485_;
wire _80486_;
wire _80487_;
wire _80488_;
wire _80489_;
wire _80490_;
wire _80491_;
wire _80492_;
wire _80493_;
wire _80494_;
wire _80495_;
wire _80496_;
wire _80497_;
wire _80498_;
wire _80499_;
wire _80500_;
wire _80501_;
wire _80502_;
wire _80503_;
wire _80504_;
wire _80505_;
wire _80506_;
wire _80507_;
wire _80508_;
wire _80509_;
wire _80510_;
wire _80511_;
wire _80512_;
wire _80513_;
wire _80514_;
wire _80515_;
wire _80516_;
wire _80517_;
wire _80518_;
wire _80519_;
wire _80520_;
wire _80521_;
wire _80522_;
wire _80523_;
wire _80524_;
wire _80525_;
wire _80526_;
wire _80527_;
wire _80528_;
wire _80529_;
wire _80530_;
wire _80531_;
wire _80532_;
wire _80533_;
wire _80534_;
wire _80535_;
wire _80536_;
wire _80537_;
wire _80538_;
wire _80539_;
wire _80540_;
wire _80541_;
wire _80542_;
wire _80543_;
wire _80544_;
wire _80545_;
wire _80546_;
wire _80547_;
wire _80548_;
wire _80549_;
wire _80550_;
wire _80551_;
wire _80552_;
wire _80553_;
wire _80554_;
wire _80555_;
wire _80556_;
wire _80557_;
wire _80558_;
wire _80559_;
wire _80560_;
wire _80561_;
wire _80562_;
wire _80563_;
wire _80564_;
wire _80565_;
wire _80566_;
wire _80567_;
wire _80568_;
wire _80569_;
wire _80570_;
wire _80571_;
wire _80572_;
wire _80573_;
wire _80574_;
wire _80575_;
wire _80576_;
wire _80577_;
wire _80578_;
wire _80579_;
wire _80580_;
wire _80581_;
wire _80582_;
wire _80583_;
wire _80584_;
wire _80585_;
wire _80586_;
wire _80587_;
wire _80588_;
wire _80589_;
wire _80590_;
wire _80591_;
wire _80592_;
wire _80593_;
wire _80594_;
wire _80595_;
wire _80596_;
wire _80597_;
wire _80598_;
wire _80599_;
wire _80600_;
wire _80601_;
wire _80602_;
wire _80603_;
wire _80604_;
wire _80605_;
wire _80606_;
wire _80607_;
wire _80608_;
wire _80609_;
wire _80610_;
wire _80611_;
wire _80612_;
wire _80613_;
wire _80614_;
wire _80615_;
wire _80616_;
wire _80617_;
wire _80618_;
wire _80619_;
wire _80620_;
wire _80621_;
wire _80622_;
wire _80623_;
wire _80624_;
wire _80625_;
wire _80626_;
wire _80627_;
wire _80628_;
wire _80629_;
wire _80630_;
wire _80631_;
wire _80632_;
wire _80633_;
wire _80634_;
wire _80635_;
wire _80636_;
wire _80637_;
wire _80638_;
wire _80639_;
wire _80640_;
wire _80641_;
wire _80642_;
wire _80643_;
wire _80644_;
wire _80645_;
wire _80646_;
wire _80647_;
wire _80648_;
wire _80649_;
wire _80650_;
wire _80651_;
wire _80652_;
wire _80653_;
wire _80654_;
wire _80655_;
wire _80656_;
wire _80657_;
wire _80658_;
wire _80659_;
wire _80660_;
wire _80661_;
wire _80662_;
wire _80663_;
wire _80664_;
wire _80665_;
wire _80666_;
wire _80667_;
wire _80668_;
wire _80669_;
wire _80670_;
wire _80671_;
wire _80672_;
wire _80673_;
wire _80674_;
wire _80675_;
wire _80676_;
wire _80677_;
wire _80678_;
wire _80679_;
wire _80680_;
wire _80681_;
wire _80682_;
wire _80683_;
wire _80684_;
wire _80685_;
wire _80686_;
wire _80687_;
wire _80688_;
wire _80689_;
wire _80690_;
wire _80691_;
wire _80692_;
wire _80693_;
wire _80694_;
wire _80695_;
wire _80696_;
wire _80697_;
wire _80698_;
wire _80699_;
wire _80700_;
wire _80701_;
wire _80702_;
wire _80703_;
wire _80704_;
wire _80705_;
wire _80706_;
wire _80707_;
wire _80708_;
wire _80709_;
wire _80710_;
wire _80711_;
wire _80712_;
wire _80713_;
wire _80714_;
wire _80715_;
wire _80716_;
wire _80717_;
wire _80718_;
wire _80719_;
wire _80720_;
wire _80721_;
wire _80722_;
wire _80723_;
wire _80724_;
wire _80725_;
wire _80726_;
wire _80727_;
wire _80728_;
wire _80729_;
wire _80730_;
wire _80731_;
wire _80732_;
wire _80733_;
wire _80734_;
wire _80735_;
wire _80736_;
wire _80737_;
wire _80738_;
wire _80739_;
wire _80740_;
wire _80741_;
wire _80742_;
wire _80743_;
wire _80744_;
wire _80745_;
wire _80746_;
wire _80747_;
wire _80748_;
wire _80749_;
wire _80750_;
wire _80751_;
wire _80752_;
wire _80753_;
wire _80754_;
wire _80755_;
wire _80756_;
wire _80757_;
wire _80758_;
wire _80759_;
wire _80760_;
wire _80761_;
wire _80762_;
wire _80763_;
wire _80764_;
wire _80765_;
wire _80766_;
wire _80767_;
wire _80768_;
wire _80769_;
wire _80770_;
wire _80771_;
wire _80772_;
wire _80773_;
wire _80774_;
wire _80775_;
wire _80776_;
wire _80777_;
wire _80778_;
wire _80779_;
wire _80780_;
wire _80781_;
wire _80782_;
wire _80783_;
wire _80784_;
wire _80785_;
wire _80786_;
wire _80787_;
wire _80788_;
wire _80789_;
wire _80790_;
wire _80791_;
wire _80792_;
wire _80793_;
wire _80794_;
wire _80795_;
wire _80796_;
wire _80797_;
wire _80798_;
wire _80799_;
wire _80800_;
wire _80801_;
wire _80802_;
wire _80803_;
wire _80804_;
wire _80805_;
wire _80806_;
wire _80807_;
wire _80808_;
wire _80809_;
wire _80810_;
wire _80811_;
wire _80812_;
wire _80813_;
wire _80814_;
wire _80815_;
wire _80816_;
wire _80817_;
wire _80818_;
wire _80819_;
wire _80820_;
wire _80821_;
wire _80822_;
wire _80823_;
wire _80824_;
wire _80825_;
wire _80826_;
wire _80827_;
wire _80828_;
wire _80829_;
wire _80830_;
wire _80831_;
wire _80832_;
wire _80833_;
wire _80834_;
wire _80835_;
wire _80836_;
wire _80837_;
wire _80838_;
wire _80839_;
wire _80840_;
wire _80841_;
wire _80842_;
wire _80843_;
wire _80844_;
wire _80845_;
wire _80846_;
wire _80847_;
wire _80848_;
wire _80849_;
wire _80850_;
wire _80851_;
wire _80852_;
wire _80853_;
wire _80854_;
wire _80855_;
wire _80856_;
wire _80857_;
wire _80858_;
wire _80859_;
wire _80860_;
wire _80861_;
wire _80862_;
wire _80863_;
wire _80864_;
wire _80865_;
wire _80866_;
wire _80867_;
wire _80868_;
wire _80869_;
wire _80870_;
wire _80871_;
wire _80872_;
wire _80873_;
wire _80874_;
wire _80875_;
wire _80876_;
wire _80877_;
wire _80878_;
wire _80879_;
wire _80880_;
wire _80881_;
wire _80882_;
wire _80883_;
wire _80884_;
wire _80885_;
wire _80886_;
wire _80887_;
wire _80888_;
wire _80889_;
wire _80890_;
wire _80891_;
wire _80892_;
wire _80893_;
wire _80894_;
wire _80895_;
wire _80896_;
wire _80897_;
wire _80898_;
wire _80899_;
wire _80900_;
wire _80901_;
wire _80902_;
wire _80903_;
wire _80904_;
wire _80905_;
wire _80906_;
wire _80907_;
wire _80908_;
wire _80909_;
wire _80910_;
wire _80911_;
wire _80912_;
wire _80913_;
wire _80914_;
wire _80915_;
wire _80916_;
wire _80917_;
wire _80918_;
wire _80919_;
wire _80920_;
wire _80921_;
wire _80922_;
wire _80923_;
wire _80924_;
wire _80925_;
wire _80926_;
wire _80927_;
wire _80928_;
wire _80929_;
wire _80930_;
wire _80931_;
wire _80932_;
wire _80933_;
wire _80934_;
wire _80935_;
wire _80936_;
wire _80937_;
wire _80938_;
wire _80939_;
wire _80940_;
wire _80941_;
wire _80942_;
wire _80943_;
wire _80944_;
wire _80945_;
wire _80946_;
wire _80947_;
wire _80948_;
wire _80949_;
wire _80950_;
wire _80951_;
wire _80952_;
wire _80953_;
wire _80954_;
wire _80955_;
wire _80956_;
wire _80957_;
wire _80958_;
wire _80959_;
wire _80960_;
wire _80961_;
wire _80962_;
wire _80963_;
wire _80964_;
wire _80965_;
wire _80966_;
wire _80967_;
wire _80968_;
wire _80969_;
wire _80970_;
wire _80971_;
wire _80972_;
wire _80973_;
wire _80974_;
wire _80975_;
wire _80976_;
wire _80977_;
wire _80978_;
wire _80979_;
wire _80980_;
wire _80981_;
wire _80982_;
wire _80983_;
wire _80984_;
wire _80985_;
wire _80986_;
wire _80987_;
wire _80988_;
wire _80989_;
wire _80990_;
wire _80991_;
wire _80992_;
wire _80993_;
wire _80994_;
wire _80995_;
wire _80996_;
wire _80997_;
wire _80998_;
wire _80999_;
wire _81000_;
wire _81001_;
wire _81002_;
wire _81003_;
wire _81004_;
wire _81005_;
wire _81006_;
wire _81007_;
wire _81008_;
wire _81009_;
wire _81010_;
wire _81011_;
wire _81012_;
wire _81013_;
wire _81014_;
wire _81015_;
wire _81016_;
wire _81017_;
wire _81018_;
wire _81019_;
wire _81020_;
wire _81021_;
wire _81022_;
wire _81023_;
wire _81024_;
wire _81025_;
wire _81026_;
wire _81027_;
wire _81028_;
wire _81029_;
wire _81030_;
wire _81031_;
wire _81032_;
wire _81033_;
wire _81034_;
wire _81035_;
wire _81036_;
wire _81037_;
wire _81038_;
wire _81039_;
wire _81040_;
wire _81041_;
wire _81042_;
wire _81043_;
wire _81044_;
wire _81045_;
wire _81046_;
wire _81047_;
wire _81048_;
wire _81049_;
wire _81050_;
wire _81051_;
wire _81052_;
wire _81053_;
wire _81054_;
wire _81055_;
wire _81056_;
wire _81057_;
wire _81058_;
wire _81059_;
wire _81060_;
wire _81061_;
wire _81062_;
wire _81063_;
wire _81064_;
wire _81065_;
wire _81066_;
wire _81067_;
wire _81068_;
wire _81069_;
wire _81070_;
wire _81071_;
wire _81072_;
wire _81073_;
wire _81074_;
wire _81075_;
wire _81076_;
wire _81077_;
wire _81078_;
wire _81079_;
wire _81080_;
wire _81081_;
wire _81082_;
wire _81083_;
wire _81084_;
wire _81085_;
wire _81086_;
wire _81087_;
wire _81088_;
wire _81089_;
wire _81090_;
wire _81091_;
wire _81092_;
wire _81093_;
wire _81094_;
wire _81095_;
wire _81096_;
wire _81097_;
wire _81098_;
wire _81099_;
wire _81100_;
wire _81101_;
wire _81102_;
wire _81103_;
wire _81104_;
wire _81105_;
wire _81106_;
wire _81107_;
wire _81108_;
wire _81109_;
wire _81110_;
wire _81111_;
wire _81112_;
wire _81113_;
wire _81114_;
wire _81115_;
wire _81116_;
wire _81117_;
wire _81118_;
wire _81119_;
wire _81120_;
wire _81121_;
wire _81122_;
wire _81123_;
wire _81124_;
wire _81125_;
wire _81126_;
wire _81127_;
wire _81128_;
wire _81129_;
wire _81130_;
wire _81131_;
wire _81132_;
wire _81133_;
wire _81134_;
wire _81135_;
wire _81136_;
wire _81137_;
wire _81138_;
wire _81139_;
wire _81140_;
wire _81141_;
wire _81142_;
wire _81143_;
wire _81144_;
wire _81145_;
wire _81146_;
wire _81147_;
wire _81148_;
wire _81149_;
wire _81150_;
wire _81151_;
wire _81152_;
wire _81153_;
wire _81154_;
wire _81155_;
wire _81156_;
wire _81157_;
wire _81158_;
wire _81159_;
wire _81160_;
wire _81161_;
wire _81162_;
wire _81163_;
wire _81164_;
wire _81165_;
wire _81166_;
wire _81167_;
wire _81168_;
wire _81169_;
wire _81170_;
wire _81171_;
wire _81172_;
wire _81173_;
wire _81174_;
wire _81175_;
wire _81176_;
wire _81177_;
wire _81178_;
wire _81179_;
wire _81180_;
wire _81181_;
wire _81182_;
wire _81183_;
wire _81184_;
wire _81185_;
wire _81186_;
wire _81187_;
wire _81188_;
wire _81189_;
wire _81190_;
wire _81191_;
wire _81192_;
wire _81193_;
wire _81194_;
wire _81195_;
wire _81196_;
wire _81197_;
wire _81198_;
wire _81199_;
wire _81200_;
wire _81201_;
wire _81202_;
wire _81203_;
wire _81204_;
wire _81205_;
wire _81206_;
wire _81207_;
wire _81208_;
wire _81209_;
wire _81210_;
wire _81211_;
wire _81212_;
wire _81213_;
wire _81214_;
wire _81215_;
wire _81216_;
wire _81217_;
wire _81218_;
wire _81219_;
wire _81220_;
wire _81221_;
wire _81222_;
wire _81223_;
wire _81224_;
wire _81225_;
wire _81226_;
wire _81227_;
wire _81228_;
wire _81229_;
wire _81230_;
wire _81231_;
wire _81232_;
wire _81233_;
wire _81234_;
wire _81235_;
wire _81236_;
wire _81237_;
wire _81238_;
wire _81239_;
wire _81240_;
wire _81241_;
wire _81242_;
wire _81243_;
wire _81244_;
wire _81245_;
wire _81246_;
wire _81247_;
wire _81248_;
wire _81249_;
wire _81250_;
wire _81251_;
wire _81252_;
wire _81253_;
wire _81254_;
wire _81255_;
wire _81256_;
wire _81257_;
wire _81258_;
wire _81259_;
wire _81260_;
wire _81261_;
wire _81262_;
wire _81263_;
wire _81264_;
wire _81265_;
wire _81266_;
wire _81267_;
wire _81268_;
wire _81269_;
wire _81270_;
wire _81271_;
wire _81272_;
wire _81273_;
wire _81274_;
wire _81275_;
wire _81276_;
wire _81277_;
wire _81278_;
wire _81279_;
wire _81280_;
wire _81281_;
wire _81282_;
wire _81283_;
wire _81284_;
wire _81285_;
wire _81286_;
wire _81287_;
wire _81288_;
wire _81289_;
wire _81290_;
wire _81291_;
wire _81292_;
wire _81293_;
wire _81294_;
wire _81295_;
wire _81296_;
wire _81297_;
wire _81298_;
wire _81299_;
wire _81300_;
wire _81301_;
wire _81302_;
wire _81303_;
wire _81304_;
wire _81305_;
wire _81306_;
wire _81307_;
wire _81308_;
wire _81309_;
wire _81310_;
wire _81311_;
wire _81312_;
wire _81313_;
wire _81314_;
wire _81315_;
wire _81316_;
wire _81317_;
wire _81318_;
wire _81319_;
wire _81320_;
wire _81321_;
wire _81322_;
wire _81323_;
wire _81324_;
wire _81325_;
wire _81326_;
wire _81327_;
wire _81328_;
wire _81329_;
wire _81330_;
wire _81331_;
wire _81332_;
wire _81333_;
wire _81334_;
wire _81335_;
wire _81336_;
wire _81337_;
wire _81338_;
wire _81339_;
wire _81340_;
wire _81341_;
wire _81342_;
wire _81343_;
wire _81344_;
wire _81345_;
wire _81346_;
wire _81347_;
wire _81348_;
wire _81349_;
wire _81350_;
wire _81351_;
wire _81352_;
wire _81353_;
wire _81354_;
wire _81355_;
wire _81356_;
wire _81357_;
wire _81358_;
wire _81359_;
wire _81360_;
wire _81361_;
wire _81362_;
wire _81363_;
wire _81364_;
wire _81365_;
wire _81366_;
wire _81367_;
wire _81368_;
wire _81369_;
wire _81370_;
wire _81371_;
wire _81372_;
wire _81373_;
wire _81374_;
wire _81375_;
wire _81376_;
wire _81377_;
wire _81378_;
wire _81379_;
wire _81380_;
wire _81381_;
wire _81382_;
wire _81383_;
wire _81384_;
wire _81385_;
wire _81386_;
wire _81387_;
wire _81388_;
wire _81389_;
wire _81390_;
wire _81391_;
wire _81392_;
wire _81393_;
wire _81394_;
wire _81395_;
wire _81396_;
wire _81397_;
wire _81398_;
wire _81399_;
wire _81400_;
wire _81401_;
wire _81402_;
wire _81403_;
wire _81404_;
wire _81405_;
wire _81406_;
wire _81407_;
wire _81408_;
wire _81409_;
wire _81410_;
wire _81411_;
wire _81412_;
wire _81413_;
wire _81414_;
wire _81415_;
wire _81416_;
wire _81417_;
wire _81418_;
wire _81419_;
wire _81420_;
wire _81421_;
wire _81422_;
wire _81423_;
wire _81424_;
wire _81425_;
wire _81426_;
wire _81427_;
wire _81428_;
wire _81429_;
wire _81430_;
wire _81431_;
wire _81432_;
wire _81433_;
wire _81434_;
wire _81435_;
wire _81436_;
wire _81437_;
wire _81438_;
wire _81439_;
wire _81440_;
wire _81441_;
wire _81442_;
wire _81443_;
wire _81444_;
wire _81445_;
wire _81446_;
wire _81447_;
wire _81448_;
wire _81449_;
wire _81450_;
wire _81451_;
wire _81452_;
wire _81453_;
wire _81454_;
wire _81455_;
wire _81456_;
wire _81457_;
wire _81458_;
wire _81459_;
wire _81460_;
wire _81461_;
wire _81462_;
wire _81463_;
wire _81464_;
wire _81465_;
wire _81466_;
wire _81467_;
wire _81468_;
wire _81469_;
wire _81470_;
wire _81471_;
wire _81472_;
wire _81473_;
wire _81474_;
wire _81475_;
wire _81476_;
wire _81477_;
wire _81478_;
wire _81479_;
wire _81480_;
wire _81481_;
wire _81482_;
wire _81483_;
wire _81484_;
wire _81485_;
wire _81486_;
wire _81487_;
wire _81488_;
wire _81489_;
wire _81490_;
wire _81491_;
wire _81492_;
wire _81493_;
wire _81494_;
wire _81495_;
wire _81496_;
wire _81497_;
wire _81498_;
wire _81499_;
wire _81500_;
wire _81501_;
wire _81502_;
wire _81503_;
wire _81504_;
wire _81505_;
wire _81506_;
wire _81507_;
wire _81508_;
wire _81509_;
wire _81510_;
wire _81511_;
wire _81512_;
wire _81513_;
wire _81514_;
wire _81515_;
wire _81516_;
wire _81517_;
wire _81518_;
wire _81519_;
wire _81520_;
wire _81521_;
wire _81522_;
wire _81523_;
wire _81524_;
wire _81525_;
wire _81526_;
wire _81527_;
wire _81528_;
wire _81529_;
wire _81530_;
wire _81531_;
wire _81532_;
wire _81533_;
wire _81534_;
wire _81535_;
wire _81536_;
wire _81537_;
wire _81538_;
wire _81539_;
wire _81540_;
wire _81541_;
wire _81542_;
wire _81543_;
wire _81544_;
wire _81545_;
wire _81546_;
wire _81547_;
wire _81548_;
wire _81549_;
wire _81550_;
wire _81551_;
wire _81552_;
wire _81553_;
wire _81554_;
wire _81555_;
wire _81556_;
wire _81557_;
wire _81558_;
wire _81559_;
wire _81560_;
wire _81561_;
wire _81562_;
wire _81563_;
wire _81564_;
wire _81565_;
wire _81566_;
wire _81567_;
wire _81568_;
wire _81569_;
wire _81570_;
wire _81571_;
wire _81572_;
wire _81573_;
wire _81574_;
wire _81575_;
wire _81576_;
wire _81577_;
wire _81578_;
wire _81579_;
wire _81580_;
wire _81581_;
wire _81582_;
wire _81583_;
wire _81584_;
wire _81585_;
wire _81586_;
wire _81587_;
wire _81588_;
wire _81589_;
wire _81590_;
wire _81591_;
wire _81592_;
wire _81593_;
wire _81594_;
wire _81595_;
wire _81596_;
wire _81597_;
wire _81598_;
wire _81599_;
wire _81600_;
wire _81601_;
wire _81602_;
wire _81603_;
wire _81604_;
wire _81605_;
wire _81606_;
wire _81607_;
wire _81608_;
wire _81609_;
wire _81610_;
wire _81611_;
wire _81612_;
wire _81613_;
wire _81614_;
wire _81615_;
wire _81616_;
wire _81617_;
wire _81618_;
wire _81619_;
wire _81620_;
wire _81621_;
wire _81622_;
wire _81623_;
wire _81624_;
wire _81625_;
wire _81626_;
wire _81627_;
wire _81628_;
wire _81629_;
wire _81630_;
wire _81631_;
wire _81632_;
wire _81633_;
wire _81634_;
wire _81635_;
wire _81636_;
wire _81637_;
wire _81638_;
wire _81639_;
wire _81640_;
wire _81641_;
wire _81642_;
wire _81643_;
wire _81644_;
wire _81645_;
wire _81646_;
wire _81647_;
wire _81648_;
wire _81649_;
wire _81650_;
wire _81651_;
wire _81652_;
wire _81653_;
wire _81654_;
wire _81655_;
wire _81656_;
wire _81657_;
wire _81658_;
wire _81659_;
wire _81660_;
wire _81661_;
wire _81662_;
wire _81663_;
wire _81664_;
wire _81665_;
wire _81666_;
wire _81667_;
wire _81668_;
wire _81669_;
wire _81670_;
wire _81671_;
wire _81672_;
wire _81673_;
wire _81674_;
wire _81675_;
wire _81676_;
wire _81677_;
wire _81678_;
wire _81679_;
wire _81680_;
wire _81681_;
wire _81682_;
wire _81683_;
wire _81684_;
wire _81685_;
wire _81686_;
wire _81687_;
wire _81688_;
wire _81689_;
wire _81690_;
wire _81691_;
wire _81692_;
wire _81693_;
wire _81694_;
wire _81695_;
wire _81696_;
wire _81697_;
wire _81698_;
wire _81699_;
wire _81700_;
wire _81701_;
wire _81702_;
wire _81703_;
wire _81704_;
wire _81705_;
wire _81706_;
wire _81707_;
wire _81708_;
wire _81709_;
wire _81710_;
wire _81711_;
wire _81712_;
wire _81713_;
wire _81714_;
wire _81715_;
wire _81716_;
wire _81717_;
wire _81718_;
wire _81719_;
wire _81720_;
wire _81721_;
wire _81722_;
wire _81723_;
wire _81724_;
wire _81725_;
wire _81726_;
wire _81727_;
wire _81728_;
wire _81729_;
wire _81730_;
wire _81731_;
wire _81732_;
wire _81733_;
wire _81734_;
wire _81735_;
wire _81736_;
wire _81737_;
wire _81738_;
wire _81739_;
wire _81740_;
wire _81741_;
wire _81742_;
wire _81743_;
wire _81744_;
wire _81745_;
wire _81746_;
wire _81747_;
wire _81748_;
wire _81749_;
wire _81750_;
wire _81751_;
wire _81752_;
wire _81753_;
wire _81754_;
wire _81755_;
wire _81756_;
wire _81757_;
wire _81758_;
wire _81759_;
wire _81760_;
wire _81761_;
wire _81762_;
wire _81763_;
wire _81764_;
wire _81765_;
wire _81766_;
wire _81767_;
wire _81768_;
wire _81769_;
wire _81770_;
wire _81771_;
wire _81772_;
wire _81773_;
wire _81774_;
wire _81775_;
wire _81776_;
wire _81777_;
wire _81778_;
wire _81779_;
wire _81780_;
wire _81781_;
wire _81782_;
wire _81783_;
wire _81784_;
wire _81785_;
wire _81786_;
wire _81787_;
wire _81788_;
wire _81789_;
wire _81790_;
wire _81791_;
wire _81792_;
wire _81793_;
wire _81794_;
wire _81795_;
wire _81796_;
wire _81797_;
wire _81798_;
wire _81799_;
wire _81800_;
wire _81801_;
wire _81802_;
wire _81803_;
wire _81804_;
wire _81805_;
wire _81806_;
wire _81807_;
wire _81808_;
wire _81809_;
wire _81810_;
wire _81811_;
wire _81812_;
wire _81813_;
wire _81814_;
wire _81815_;
wire _81816_;
wire _81817_;
wire _81818_;
wire _81819_;
wire _81820_;
wire _81821_;
wire _81822_;
wire _81823_;
wire _81824_;
wire _81825_;
wire _81826_;
wire _81827_;
wire _81828_;
wire _81829_;
wire _81830_;
wire _81831_;
wire _81832_;
wire _81833_;
wire _81834_;
wire _81835_;
wire _81836_;
wire _81837_;
wire _81838_;
wire _81839_;
wire _81840_;
wire _81841_;
wire _81842_;
wire _81843_;
wire _81844_;
wire _81845_;
wire _81846_;
wire _81847_;
wire _81848_;
wire _81849_;
wire _81850_;
wire _81851_;
wire _81852_;
wire _81853_;
wire _81854_;
wire _81855_;
wire _81856_;
wire _81857_;
wire _81858_;
wire _81859_;
wire _81860_;
wire _81861_;
wire _81862_;
wire _81863_;
wire _81864_;
wire _81865_;
wire _81866_;
wire _81867_;
wire _81868_;
wire _81869_;
wire _81870_;
wire _81871_;
wire _81872_;
wire _81873_;
wire _81874_;
wire _81875_;
wire _81876_;
wire _81877_;
wire _81878_;
wire _81879_;
wire _81880_;
wire _81881_;
wire _81882_;
wire _81883_;
wire _81884_;
wire _81885_;
wire _81886_;
wire _81887_;
wire _81888_;
wire _81889_;
wire _81890_;
wire _81891_;
wire _81892_;
wire _81893_;
wire _81894_;
wire _81895_;
wire _81896_;
wire _81897_;
wire _81898_;
wire _81899_;
wire _81900_;
wire _81901_;
wire _81902_;
wire _81903_;
wire _81904_;
wire _81905_;
wire _81906_;
wire _81907_;
wire _81908_;
wire _81909_;
wire _81910_;
wire _81911_;
wire _81912_;
wire _81913_;
wire _81914_;
wire _81915_;
wire _81916_;
wire _81917_;
wire _81918_;
wire _81919_;
wire _81920_;
wire _81921_;
wire _81922_;
wire _81923_;
wire _81924_;
wire _81925_;
wire _81926_;
wire _81927_;
wire _81928_;
wire _81929_;
wire _81930_;
wire _81931_;
wire _81932_;
wire _81933_;
wire _81934_;
wire _81935_;
wire _81936_;
wire _81937_;
wire _81938_;
wire _81939_;
wire _81940_;
wire _81941_;
wire _81942_;
wire _81943_;
wire _81944_;
wire _81945_;
wire _81946_;
wire _81947_;
wire _81948_;
wire _81949_;
wire _81950_;
wire _81951_;
wire _81952_;
wire _81953_;
wire _81954_;
wire _81955_;
wire _81956_;
wire _81957_;
wire _81958_;
wire _81959_;
wire _81960_;
wire _81961_;
wire _81962_;
wire _81963_;
wire _81964_;
wire _81965_;
wire _81966_;
wire _81967_;
wire _81968_;
wire _81969_;
wire _81970_;
wire _81971_;
wire _81972_;
wire _81973_;
wire _81974_;
wire _81975_;
wire _81976_;
wire _81977_;
wire _81978_;
wire _81979_;
wire _81980_;
wire _81981_;
wire _81982_;
wire _81983_;
wire _81984_;
wire _81985_;
wire _81986_;
wire _81987_;
wire _81988_;
wire _81989_;
wire _81990_;
wire _81991_;
wire _81992_;
wire _81993_;
wire _81994_;
wire _81995_;
wire _81996_;
wire _81997_;
wire _81998_;
wire _81999_;
wire _82000_;
wire _82001_;
wire _82002_;
wire _82003_;
wire _82004_;
wire _82005_;
wire _82006_;
wire _82007_;
wire _82008_;
wire _82009_;
wire _82010_;
wire _82011_;
wire _82012_;
wire _82013_;
wire _82014_;
wire _82015_;
wire _82016_;
wire _82017_;
wire _82018_;
wire _82019_;
wire _82020_;
wire _82021_;
wire _82022_;
wire _82023_;
wire _82024_;
wire _82025_;
wire _82026_;
wire _82027_;
wire _82028_;
wire _82029_;
wire _82030_;
wire _82031_;
wire _82032_;
wire _82033_;
wire _82034_;
wire _82035_;
wire _82036_;
wire _82037_;
wire _82038_;
wire _82039_;
wire _82040_;
wire _82041_;
wire _82042_;
wire _82043_;
wire _82044_;
wire _82045_;
wire _82046_;
wire _82047_;
wire _82048_;
wire _82049_;
wire _82050_;
wire _82051_;
wire _82052_;
wire _82053_;
wire _82054_;
wire _82055_;
wire _82056_;
wire _82057_;
wire _82058_;
wire _82059_;
wire _82060_;
wire _82061_;
wire _82062_;
wire _82063_;
wire _82064_;
wire _82065_;
wire _82066_;
wire _82067_;
wire _82068_;
wire _82069_;
wire _82070_;
wire _82071_;
wire _82072_;
wire _82073_;
wire _82074_;
wire _82075_;
wire _82076_;
wire _82077_;
wire _82078_;
wire _82079_;
wire _82080_;
wire _82081_;
wire _82082_;
wire _82083_;
wire _82084_;
wire _82085_;
wire _82086_;
wire _82087_;
wire _82088_;
wire _82089_;
wire _82090_;
wire _82091_;
wire _82092_;
wire _82093_;
wire _82094_;
wire _82095_;
wire _82096_;
wire _82097_;
wire _82098_;
wire _82099_;
wire _82100_;
wire _82101_;
wire _82102_;
wire _82103_;
wire _82104_;
wire _82105_;
wire _82106_;
wire _82107_;
wire _82108_;
wire _82109_;
wire _82110_;
wire _82111_;
wire _82112_;
wire _82113_;
wire _82114_;
wire _82115_;
wire _82116_;
wire _82117_;
wire _82118_;
wire _82119_;
wire _82120_;
wire _82121_;
wire _82122_;
wire _82123_;
wire _82124_;
wire _82125_;
wire _82126_;
wire _82127_;
wire _82128_;
wire _82129_;
wire _82130_;
wire _82131_;
wire _82132_;
wire _82133_;
wire _82134_;
wire _82135_;
wire _82136_;
wire _82137_;
wire _82138_;
wire _82139_;
wire _82140_;
wire _82141_;
wire _82142_;
wire _82143_;
wire _82144_;
wire _82145_;
wire _82146_;
wire _82147_;
wire _82148_;
wire _82149_;
wire _82150_;
wire _82151_;
wire _82152_;
wire _82153_;
wire _82154_;
wire _82155_;
wire _82156_;
wire _82157_;
wire _82158_;
wire _82159_;
wire _82160_;
wire _82161_;
wire _82162_;
wire _82163_;
wire _82164_;
wire _82165_;
wire _82166_;
wire _82167_;
wire _82168_;
wire _82169_;
wire _82170_;
wire _82171_;
wire _82172_;
wire _82173_;
wire _82174_;
wire _82175_;
wire _82176_;
wire _82177_;
wire _82178_;
wire _82179_;
wire _82180_;
wire _82181_;
wire _82182_;
wire _82183_;
wire _82184_;
wire _82185_;
wire _82186_;
wire _82187_;
wire _82188_;
wire _82189_;
wire _82190_;
wire _82191_;
wire _82192_;
wire _82193_;
wire _82194_;
wire _82195_;
wire _82196_;
wire _82197_;
wire _82198_;
wire _82199_;
wire _82200_;
wire _82201_;
wire _82202_;
wire _82203_;
wire _82204_;
wire _82205_;
wire _82206_;
wire _82207_;
wire _82208_;
wire _82209_;
wire _82210_;
wire _82211_;
wire _82212_;
wire _82213_;
wire _82214_;
wire _82215_;
wire _82216_;
wire _82217_;
wire _82218_;
wire _82219_;
wire _82220_;
wire _82221_;
wire _82222_;
wire _82223_;
wire _82224_;
wire _82225_;
wire _82226_;
wire _82227_;
wire _82228_;
wire _82229_;
wire _82230_;
wire _82231_;
wire _82232_;
wire _82233_;
wire _82234_;
wire _82235_;
wire _82236_;
wire _82237_;
wire _82238_;
wire _82239_;
wire _82240_;
wire _82241_;
wire _82242_;
wire _82243_;
wire _82244_;
wire _82245_;
wire _82246_;
wire _82247_;
wire _82248_;
wire _82249_;
wire _82250_;
wire _82251_;
wire _82252_;
wire _82253_;
wire _82254_;
wire _82255_;
wire _82256_;
wire _82257_;
wire _82258_;
wire _82259_;
wire _82260_;
wire _82261_;
wire _82262_;
wire _82263_;
wire _82264_;
wire _82265_;
wire _82266_;
wire _82267_;
wire _82268_;
wire _82269_;
wire _82270_;
wire _82271_;
wire _82272_;
wire _82273_;
wire _82274_;
wire _82275_;
wire _82276_;
wire _82277_;
wire _82278_;
wire _82279_;
wire _82280_;
wire _82281_;
wire _82282_;
wire _82283_;
wire _82284_;
wire _82285_;
wire _82286_;
wire _82287_;
wire _82288_;
wire _82289_;
wire _82290_;
wire _82291_;
wire _82292_;
wire _82293_;
wire _82294_;
wire _82295_;
wire _82296_;
wire _82297_;
wire _82298_;
wire _82299_;
wire _82300_;
wire _82301_;
wire _82302_;
wire _82303_;
wire _82304_;
wire _82305_;
wire _82306_;
wire _82307_;
wire _82308_;
wire _82309_;
wire _82310_;
wire _82311_;
wire _82312_;
wire _82313_;
wire _82314_;
wire _82315_;
wire _82316_;
wire _82317_;
wire _82318_;
wire _82319_;
wire _82320_;
wire _82321_;
wire _82322_;
wire _82323_;
wire _82324_;
wire _82325_;
wire _82326_;
wire _82327_;
wire _82328_;
wire _82329_;
wire _82330_;
wire _82331_;
wire _82332_;
wire _82333_;
wire _82334_;
wire _82335_;
wire _82336_;
wire _82337_;
wire _82338_;
wire _82339_;
wire _82340_;
wire _82341_;
wire _82342_;
wire _82343_;
wire _82344_;
wire _82345_;
wire _82346_;
wire _82347_;
wire _82348_;
wire _82349_;
wire _82350_;
wire _82351_;
wire _82352_;
wire _82353_;
wire _82354_;
wire _82355_;
wire _82356_;
wire _82357_;
wire _82358_;
wire _82359_;
wire _82360_;
wire _82361_;
wire _82362_;
wire _82363_;
wire _82364_;
wire _82365_;
wire _82366_;
wire _82367_;
wire _82368_;
wire _82369_;
wire _82370_;
wire _82371_;
wire _82372_;
wire _82373_;
wire _82374_;
wire _82375_;
wire _82376_;
wire _82377_;
wire _82378_;
wire _82379_;
wire _82380_;
wire _82381_;
wire _82382_;
wire _82383_;
wire _82384_;
wire _82385_;
wire _82386_;
wire _82387_;
wire _82388_;
wire _82389_;
wire _82390_;
wire _82391_;
wire _82392_;
wire _82393_;
wire _82394_;
wire _82395_;
wire _82396_;
wire _82397_;
wire _82398_;
wire _82399_;
wire _82400_;
wire _82401_;
wire _82402_;
wire _82403_;
wire _82404_;
wire _82405_;
wire _82406_;
wire _82407_;
wire _82408_;
wire _82409_;
wire _82410_;
wire _82411_;
wire _82412_;
wire _82413_;
wire _82414_;
wire _82415_;
wire _82416_;
wire _82417_;
wire _82418_;
wire _82419_;
wire _82420_;
wire _82421_;
wire _82422_;
wire _82423_;
wire _82424_;
wire _82425_;
wire _82426_;
wire _82427_;
wire _82428_;
wire _82429_;
wire _82430_;
wire _82431_;
wire _82432_;
wire _82433_;
wire _82434_;
wire _82435_;
wire _82436_;
wire _82437_;
wire _82438_;
wire _82439_;
wire _82440_;
wire _82441_;
wire _82442_;
wire _82443_;
wire _82444_;
wire _82445_;
wire _82446_;
wire _82447_;
wire _82448_;
wire _82449_;
wire _82450_;
wire _82451_;
wire _82452_;
wire _82453_;
wire _82454_;
wire _82455_;
wire _82456_;
wire _82457_;
wire _82458_;
wire _82459_;
wire _82460_;
wire _82461_;
wire _82462_;
wire _82463_;
wire _82464_;
wire _82465_;
wire _82466_;
wire _82467_;
wire _82468_;
wire _82469_;
wire _82470_;
wire _82471_;
wire _82472_;
wire _82473_;
wire _82474_;
wire _82475_;
wire _82476_;
wire _82477_;
wire _82478_;
wire _82479_;
wire _82480_;
wire _82481_;
wire _82482_;
wire _82483_;
wire _82484_;
wire _82485_;
wire _82486_;
wire _82487_;
wire _82488_;
wire _82489_;
wire _82490_;
wire _82491_;
wire _82492_;
wire _82493_;
wire _82494_;
wire _82495_;
wire _82496_;
wire _82497_;
wire _82498_;
wire _82499_;
wire _82500_;
wire _82501_;
wire _82502_;
wire _82503_;
wire _82504_;
wire _82505_;
wire _82506_;
wire _82507_;
wire _82508_;
wire _82509_;
wire _82510_;
wire _82511_;
wire _82512_;
wire _82513_;
wire _82514_;
wire _82515_;
wire _82516_;
wire _82517_;
wire _82518_;
wire _82519_;
wire _82520_;
wire _82521_;
wire _82522_;
wire _82523_;
wire _82524_;
wire _82525_;
wire _82526_;
wire _82527_;
wire _82528_;
wire _82529_;
wire _82530_;
wire _82531_;
wire _82532_;
wire _82533_;
wire _82534_;
wire _82535_;
wire _82536_;
wire _82537_;
wire _82538_;
wire _82539_;
wire _82540_;
wire _82541_;
wire _82542_;
wire _82543_;
wire _82544_;
wire _82545_;
wire _82546_;
wire _82547_;
wire _82548_;
wire _82549_;
wire _82550_;
wire _82551_;
wire _82552_;
wire _82553_;
wire _82554_;
wire _82555_;
wire _82556_;
wire _82557_;
wire _82558_;
wire _82559_;
wire _82560_;
wire _82561_;
wire _82562_;
wire _82563_;
wire _82564_;
wire _82565_;
wire _82566_;
wire _82567_;
wire _82568_;
wire _82569_;
wire _82570_;
wire _82571_;
wire _82572_;
wire _82573_;
wire _82574_;
wire _82575_;
wire _82576_;
wire _82577_;
wire _82578_;
wire _82579_;
wire _82580_;
wire _82581_;
wire _82582_;
wire _82583_;
wire _82584_;
wire _82585_;
wire _82586_;
wire _82587_;
wire _82588_;
wire _82589_;
wire _82590_;
wire _82591_;
wire _82592_;
wire _82593_;
wire _82594_;
wire _82595_;
wire _82596_;
wire _82597_;
wire _82598_;
wire _82599_;
wire _82600_;
wire _82601_;
wire _82602_;
wire _82603_;
wire _82604_;
wire _82605_;
wire _82606_;
wire _82607_;
wire _82608_;
wire _82609_;
wire _82610_;
wire _82611_;
wire _82612_;
wire _82613_;
wire _82614_;
wire _82615_;
wire _82616_;
wire _82617_;
wire _82618_;
wire _82619_;
wire _82620_;
wire _82621_;
wire _82622_;
wire _82623_;
wire _82624_;
wire _82625_;
wire _82626_;
wire _82627_;
wire _82628_;
wire _82629_;
wire _82630_;
wire _82631_;
wire _82632_;
wire _82633_;
wire _82634_;
wire _82635_;
wire _82636_;
wire _82637_;
wire _82638_;
wire _82639_;
wire _82640_;
wire _82641_;
wire _82642_;
wire _82643_;
wire _82644_;
wire _82645_;
wire _82646_;
wire _82647_;
wire _82648_;
wire _82649_;
wire _82650_;
wire _82651_;
wire _82652_;
wire _82653_;
wire _82654_;
wire _82655_;
wire _82656_;
wire _82657_;
wire _82658_;
wire _82659_;
wire _82660_;
wire _82661_;
wire _82662_;
wire _82663_;
wire _82664_;
wire _82665_;
wire _82666_;
wire _82667_;
wire _82668_;
wire _82669_;
wire _82670_;
wire _82671_;
wire _82672_;
wire _82673_;
wire _82674_;
wire _82675_;
wire _82676_;
wire _82677_;
wire _82678_;
wire _82679_;
wire _82680_;
wire _82681_;
wire _82682_;
wire _82683_;
wire _82684_;
wire _82685_;
wire _82686_;
wire _82687_;
wire _82688_;
wire _82689_;
wire _82690_;
wire _82691_;
wire _82692_;
wire _82693_;
wire _82694_;
wire _82695_;
wire _82696_;
wire _82697_;
wire _82698_;
wire _82699_;
wire _82700_;
wire _82701_;
wire _82702_;
wire _82703_;
wire _82704_;
wire _82705_;
wire _82706_;
wire _82707_;
wire _82708_;
wire _82709_;
wire _82710_;
wire _82711_;
wire _82712_;
wire _82713_;
wire _82714_;
wire _82715_;
wire _82716_;
wire _82717_;
wire _82718_;
wire _82719_;
wire _82720_;
wire _82721_;
wire _82722_;
wire _82723_;
wire _82724_;
wire _82725_;
wire _82726_;
wire _82727_;
wire _82728_;
wire _82729_;
wire _82730_;
wire _82731_;
wire _82732_;
wire _82733_;
wire _82734_;
wire _82735_;
wire _82736_;
wire _82737_;
wire _82738_;
wire _82739_;
wire _82740_;
wire _82741_;
wire _82742_;
wire _82743_;
wire _82744_;
wire _82745_;
wire _82746_;
wire _82747_;
wire _82748_;
wire _82749_;
wire _82750_;
wire _82751_;
wire _82752_;
wire _82753_;
wire _82754_;
wire _82755_;
wire _82756_;
wire _82757_;
wire _82758_;
wire _82759_;
wire _82760_;
wire _82761_;
wire _82762_;
wire _82763_;
wire _82764_;
wire _82765_;
wire _82766_;
wire _82767_;
wire _82768_;
wire _82769_;
wire _82770_;
wire _82771_;
wire _82772_;
wire _82773_;
wire _82774_;
wire _82775_;
wire _82776_;
wire _82777_;
wire _82778_;
wire _82779_;
wire _82780_;
wire _82781_;
wire _82782_;
wire _82783_;
wire _82784_;
wire _82785_;
wire _82786_;
wire _82787_;
wire _82788_;
wire _82789_;
wire _82790_;
wire _82791_;
wire _82792_;
wire _82793_;
wire _82794_;
wire _82795_;
wire _82796_;
wire _82797_;
wire _82798_;
wire _82799_;
wire _82800_;
wire _82801_;
wire _82802_;
wire _82803_;
wire _82804_;
wire _82805_;
wire _82806_;
wire _82807_;
wire _82808_;
wire _82809_;
wire _82810_;
wire _82811_;
wire _82812_;
wire _82813_;
wire _82814_;
wire _82815_;
wire _82816_;
wire _82817_;
wire _82818_;
wire _82819_;
wire _82820_;
wire _82821_;
wire _82822_;
wire _82823_;
wire _82824_;
wire _82825_;
wire _82826_;
wire _82827_;
wire _82828_;
wire _82829_;
wire _82830_;
wire _82831_;
wire _82832_;
wire _82833_;
wire _82834_;
wire _82835_;
wire _82836_;
wire _82837_;
wire _82838_;
wire _82839_;
wire _82840_;
wire _82841_;
wire _82842_;
wire _82843_;
wire _82844_;
wire _82845_;
wire _82846_;
wire _82847_;
wire _82848_;
wire _82849_;
wire _82850_;
wire _82851_;
wire _82852_;
wire _82853_;
wire _82854_;
wire _82855_;
wire _82856_;
wire _82857_;
wire _82858_;
wire _82859_;
wire _82860_;
wire _82861_;
wire _82862_;
wire _82863_;
wire _82864_;
wire _82865_;
wire _82866_;
wire _82867_;
wire _82868_;
wire _82869_;
wire _82870_;
wire _82871_;
wire _82872_;
wire _82873_;
wire _82874_;
wire _82875_;
wire _82876_;
wire _82877_;
wire _82878_;
wire _82879_;
wire _82880_;
wire _82881_;
wire _82882_;
wire _82883_;
wire _82884_;
wire _82885_;
wire _82886_;
wire _82887_;
wire _82888_;
wire _82889_;
wire _82890_;
wire _82891_;
wire _82892_;
wire _82893_;
wire _82894_;
wire _82895_;
wire _82896_;
wire _82897_;
wire _82898_;
wire _82899_;
wire _82900_;
wire _82901_;
wire _82902_;
wire _82903_;
wire _82904_;
wire _82905_;
wire _82906_;
wire _82907_;
wire _82908_;
wire _82909_;
wire _82910_;
wire _82911_;
wire _82912_;
wire _82913_;
wire _82914_;
wire _82915_;
wire _82916_;
wire _82917_;
wire _82918_;
wire _82919_;
wire _82920_;
wire _82921_;
wire _82922_;
wire _82923_;
wire _82924_;
wire _82925_;
wire _82926_;
wire _82927_;
wire _82928_;
wire _82929_;
wire _82930_;
wire _82931_;
wire _82932_;
wire _82933_;
wire _82934_;
wire _82935_;
wire _82936_;
wire _82937_;
wire _82938_;
wire _82939_;
wire _82940_;
wire _82941_;
wire _82942_;
wire _82943_;
wire _82944_;
wire _82945_;
wire _82946_;
wire _82947_;
wire _82948_;
wire _82949_;
wire _82950_;
wire _82951_;
wire _82952_;
wire _82953_;
wire _82954_;
wire _82955_;
wire _82956_;
wire _82957_;
wire _82958_;
wire _82959_;
wire _82960_;
wire _82961_;
wire _82962_;
wire _82963_;
wire _82964_;
wire _82965_;
wire _82966_;
wire _82967_;
wire _82968_;
wire _82969_;
wire _82970_;
wire _82971_;
wire _82972_;
wire _82973_;
wire _82974_;
wire _82975_;
wire _82976_;
wire _82977_;
wire _82978_;
wire _82979_;
wire _82980_;
wire _82981_;
wire _82982_;
wire _82983_;
wire _82984_;
wire _82985_;
wire _82986_;
wire _82987_;
wire _82988_;
wire _82989_;
wire _82990_;
wire _82991_;
wire _82992_;
wire _82993_;
wire _82994_;
wire _82995_;
wire _82996_;
wire _82997_;
wire _82998_;
wire _82999_;
wire _83000_;
wire _83001_;
wire _83002_;
wire _83003_;
wire _83004_;
wire _83005_;
wire _83006_;
wire _83007_;
wire _83008_;
wire _83009_;
wire _83010_;
wire _83011_;
wire _83012_;
wire _83013_;
wire _83014_;
wire _83015_;
wire _83016_;
wire _83017_;
wire _83018_;
wire _83019_;
wire _83020_;
wire _83021_;
wire _83022_;
wire _83023_;
wire _83024_;
wire _83025_;
wire _83026_;
wire _83027_;
wire _83028_;
wire _83029_;
wire _83030_;
wire _83031_;
wire _83032_;
wire _83033_;
wire _83034_;
wire _83035_;
wire _83036_;
wire _83037_;
wire _83038_;
wire _83039_;
wire _83040_;
wire _83041_;
wire _83042_;
wire _83043_;
wire _83044_;
wire _83045_;
wire _83046_;
wire _83047_;
wire _83048_;
wire _83049_;
wire _83050_;
wire _83051_;
wire _83052_;
wire _83053_;
wire _83054_;
wire _83055_;
wire _83056_;
wire _83057_;
wire _83058_;
wire _83059_;
wire _83060_;
wire _83061_;
wire _83062_;
wire _83063_;
wire _83064_;
wire _83065_;
wire _83066_;
wire _83067_;
wire _83068_;
wire _83069_;
wire _83070_;
wire _83071_;
wire _83072_;
wire _83073_;
wire _83074_;
wire _83075_;
wire _83076_;
wire _83077_;
wire _83078_;
wire _83079_;
wire _83080_;
wire _83081_;
wire _83082_;
wire _83083_;
wire _83084_;
wire _83085_;
wire _83086_;
wire _83087_;
wire _83088_;
wire _83089_;
wire _83090_;
wire _83091_;
wire _83092_;
wire _83093_;
wire _83094_;
wire _83095_;
wire _83096_;
wire _83097_;
wire _83098_;
wire _83099_;
wire _83100_;
wire _83101_;
wire _83102_;
wire _83103_;
wire _83104_;
wire _83105_;
wire _83106_;
wire _83107_;
wire _83108_;
wire _83109_;
wire _83110_;
wire _83111_;
wire _83112_;
wire _83113_;
wire _83114_;
wire _83115_;
wire _83116_;
wire _83117_;
wire _83118_;
wire _83119_;
wire _83120_;
wire _83121_;
wire zeroWire;
wire oneWire;
assign zeroWire = 1'b0 /*99506*/;
assign oneWire = 1'b1 /*99506*/;
assign _69_ = ~D[0] /*99120*/;
assign _66_ = R_0[63] & _69_ /*99116*/;
assign _67_ = R_0[63] ^ _69_ /*99119*/;
assign _68_ = oneWire & _67_ /*99117*/;
assign _0_ = oneWire ^ _67_ /*99118*/;
assign _65_ = _66_ | _68_ /*99115*/;
assign _74_ = ~D[1] /*99114*/;
assign _71_ = R_0[64] & _74_ /*99110*/;
assign _72_ = R_0[64] ^ _74_ /*99113*/;
assign _73_ = _65_ & _72_ /*99111*/;
assign _1_ = _65_ ^ _72_ /*99112*/;
assign _70_ = _71_ | _73_ /*99109*/;
assign _79_ = ~D[2] /*99108*/;
assign _76_ = R_0[65] & _79_ /*99104*/;
assign _77_ = R_0[65] ^ _79_ /*99107*/;
assign _78_ = _70_ & _77_ /*99105*/;
assign _2_ = _70_ ^ _77_ /*99106*/;
assign _75_ = _76_ | _78_ /*99103*/;
assign _84_ = ~D[3] /*99102*/;
assign _81_ = R_0[66] & _84_ /*99098*/;
assign _82_ = R_0[66] ^ _84_ /*99101*/;
assign _83_ = _75_ & _82_ /*99099*/;
assign _3_ = _75_ ^ _82_ /*99100*/;
assign _80_ = _81_ | _83_ /*99097*/;
assign _89_ = ~D[4] /*99096*/;
assign _86_ = R_0[67] & _89_ /*99092*/;
assign _87_ = R_0[67] ^ _89_ /*99095*/;
assign _88_ = _80_ & _87_ /*99093*/;
assign _4_ = _80_ ^ _87_ /*99094*/;
assign _85_ = _86_ | _88_ /*99091*/;
assign _94_ = ~D[5] /*99090*/;
assign _91_ = R_0[68] & _94_ /*99086*/;
assign _92_ = R_0[68] ^ _94_ /*99089*/;
assign _93_ = _85_ & _92_ /*99087*/;
assign _5_ = _85_ ^ _92_ /*99088*/;
assign _90_ = _91_ | _93_ /*99085*/;
assign _99_ = ~D[6] /*99084*/;
assign _96_ = R_0[69] & _99_ /*99080*/;
assign _97_ = R_0[69] ^ _99_ /*99083*/;
assign _98_ = _90_ & _97_ /*99081*/;
assign _6_ = _90_ ^ _97_ /*99082*/;
assign _95_ = _96_ | _98_ /*99079*/;
assign _104_ = ~D[7] /*99078*/;
assign _101_ = R_0[70] & _104_ /*99074*/;
assign _102_ = R_0[70] ^ _104_ /*99077*/;
assign _103_ = _95_ & _102_ /*99075*/;
assign _7_ = _95_ ^ _102_ /*99076*/;
assign _100_ = _101_ | _103_ /*99073*/;
assign _109_ = ~D[8] /*99072*/;
assign _106_ = R_0[71] & _109_ /*99068*/;
assign _107_ = R_0[71] ^ _109_ /*99071*/;
assign _108_ = _100_ & _107_ /*99069*/;
assign _8_ = _100_ ^ _107_ /*99070*/;
assign _105_ = _106_ | _108_ /*99067*/;
assign _114_ = ~D[9] /*99066*/;
assign _111_ = R_0[72] & _114_ /*99062*/;
assign _112_ = R_0[72] ^ _114_ /*99065*/;
assign _113_ = _105_ & _112_ /*99063*/;
assign _9_ = _105_ ^ _112_ /*99064*/;
assign _110_ = _111_ | _113_ /*99061*/;
assign _119_ = ~D[10] /*99060*/;
assign _116_ = R_0[73] & _119_ /*99056*/;
assign _117_ = R_0[73] ^ _119_ /*99059*/;
assign _118_ = _110_ & _117_ /*99057*/;
assign _10_ = _110_ ^ _117_ /*99058*/;
assign _115_ = _116_ | _118_ /*99055*/;
assign _124_ = ~D[11] /*99054*/;
assign _121_ = R_0[74] & _124_ /*99050*/;
assign _122_ = R_0[74] ^ _124_ /*99053*/;
assign _123_ = _115_ & _122_ /*99051*/;
assign _11_ = _115_ ^ _122_ /*99052*/;
assign _120_ = _121_ | _123_ /*99049*/;
assign _129_ = ~D[12] /*99048*/;
assign _126_ = R_0[75] & _129_ /*99044*/;
assign _127_ = R_0[75] ^ _129_ /*99047*/;
assign _128_ = _120_ & _127_ /*99045*/;
assign _12_ = _120_ ^ _127_ /*99046*/;
assign _125_ = _126_ | _128_ /*99043*/;
assign _134_ = ~D[13] /*99042*/;
assign _131_ = R_0[76] & _134_ /*99038*/;
assign _132_ = R_0[76] ^ _134_ /*99041*/;
assign _133_ = _125_ & _132_ /*99039*/;
assign _13_ = _125_ ^ _132_ /*99040*/;
assign _130_ = _131_ | _133_ /*99037*/;
assign _139_ = ~D[14] /*99036*/;
assign _136_ = R_0[77] & _139_ /*99032*/;
assign _137_ = R_0[77] ^ _139_ /*99035*/;
assign _138_ = _130_ & _137_ /*99033*/;
assign _14_ = _130_ ^ _137_ /*99034*/;
assign _135_ = _136_ | _138_ /*99031*/;
assign _144_ = ~D[15] /*99030*/;
assign _141_ = R_0[78] & _144_ /*99026*/;
assign _142_ = R_0[78] ^ _144_ /*99029*/;
assign _143_ = _135_ & _142_ /*99027*/;
assign _15_ = _135_ ^ _142_ /*99028*/;
assign _140_ = _141_ | _143_ /*99025*/;
assign _149_ = ~D[16] /*99024*/;
assign _146_ = R_0[79] & _149_ /*99020*/;
assign _147_ = R_0[79] ^ _149_ /*99023*/;
assign _148_ = _140_ & _147_ /*99021*/;
assign _16_ = _140_ ^ _147_ /*99022*/;
assign _145_ = _146_ | _148_ /*99019*/;
assign _154_ = ~D[17] /*99018*/;
assign _151_ = R_0[80] & _154_ /*99014*/;
assign _152_ = R_0[80] ^ _154_ /*99017*/;
assign _153_ = _145_ & _152_ /*99015*/;
assign _17_ = _145_ ^ _152_ /*99016*/;
assign _150_ = _151_ | _153_ /*99013*/;
assign _159_ = ~D[18] /*99012*/;
assign _156_ = R_0[81] & _159_ /*99008*/;
assign _157_ = R_0[81] ^ _159_ /*99011*/;
assign _158_ = _150_ & _157_ /*99009*/;
assign _18_ = _150_ ^ _157_ /*99010*/;
assign _155_ = _156_ | _158_ /*99007*/;
assign _164_ = ~D[19] /*99006*/;
assign _161_ = R_0[82] & _164_ /*99002*/;
assign _162_ = R_0[82] ^ _164_ /*99005*/;
assign _163_ = _155_ & _162_ /*99003*/;
assign _19_ = _155_ ^ _162_ /*99004*/;
assign _160_ = _161_ | _163_ /*99001*/;
assign _169_ = ~D[20] /*99000*/;
assign _166_ = R_0[83] & _169_ /*98996*/;
assign _167_ = R_0[83] ^ _169_ /*98999*/;
assign _168_ = _160_ & _167_ /*98997*/;
assign _20_ = _160_ ^ _167_ /*98998*/;
assign _165_ = _166_ | _168_ /*98995*/;
assign _174_ = ~D[21] /*98994*/;
assign _171_ = R_0[84] & _174_ /*98990*/;
assign _172_ = R_0[84] ^ _174_ /*98993*/;
assign _173_ = _165_ & _172_ /*98991*/;
assign _21_ = _165_ ^ _172_ /*98992*/;
assign _170_ = _171_ | _173_ /*98989*/;
assign _179_ = ~D[22] /*98988*/;
assign _176_ = R_0[85] & _179_ /*98984*/;
assign _177_ = R_0[85] ^ _179_ /*98987*/;
assign _178_ = _170_ & _177_ /*98985*/;
assign _22_ = _170_ ^ _177_ /*98986*/;
assign _175_ = _176_ | _178_ /*98983*/;
assign _184_ = ~D[23] /*98982*/;
assign _181_ = R_0[86] & _184_ /*98978*/;
assign _182_ = R_0[86] ^ _184_ /*98981*/;
assign _183_ = _175_ & _182_ /*98979*/;
assign _23_ = _175_ ^ _182_ /*98980*/;
assign _180_ = _181_ | _183_ /*98977*/;
assign _189_ = ~D[24] /*98976*/;
assign _186_ = R_0[87] & _189_ /*98972*/;
assign _187_ = R_0[87] ^ _189_ /*98975*/;
assign _188_ = _180_ & _187_ /*98973*/;
assign _24_ = _180_ ^ _187_ /*98974*/;
assign _185_ = _186_ | _188_ /*98971*/;
assign _194_ = ~D[25] /*98970*/;
assign _191_ = R_0[88] & _194_ /*98966*/;
assign _192_ = R_0[88] ^ _194_ /*98969*/;
assign _193_ = _185_ & _192_ /*98967*/;
assign _25_ = _185_ ^ _192_ /*98968*/;
assign _190_ = _191_ | _193_ /*98965*/;
assign _199_ = ~D[26] /*98964*/;
assign _196_ = R_0[89] & _199_ /*98960*/;
assign _197_ = R_0[89] ^ _199_ /*98963*/;
assign _198_ = _190_ & _197_ /*98961*/;
assign _26_ = _190_ ^ _197_ /*98962*/;
assign _195_ = _196_ | _198_ /*98959*/;
assign _204_ = ~D[27] /*98958*/;
assign _201_ = R_0[90] & _204_ /*98954*/;
assign _202_ = R_0[90] ^ _204_ /*98957*/;
assign _203_ = _195_ & _202_ /*98955*/;
assign _27_ = _195_ ^ _202_ /*98956*/;
assign _200_ = _201_ | _203_ /*98953*/;
assign _209_ = ~D[28] /*98952*/;
assign _206_ = R_0[91] & _209_ /*98948*/;
assign _207_ = R_0[91] ^ _209_ /*98951*/;
assign _208_ = _200_ & _207_ /*98949*/;
assign _28_ = _200_ ^ _207_ /*98950*/;
assign _205_ = _206_ | _208_ /*98947*/;
assign _214_ = ~D[29] /*98946*/;
assign _211_ = R_0[92] & _214_ /*98942*/;
assign _212_ = R_0[92] ^ _214_ /*98945*/;
assign _213_ = _205_ & _212_ /*98943*/;
assign _29_ = _205_ ^ _212_ /*98944*/;
assign _210_ = _211_ | _213_ /*98941*/;
assign _219_ = ~D[30] /*98940*/;
assign _216_ = R_0[93] & _219_ /*98936*/;
assign _217_ = R_0[93] ^ _219_ /*98939*/;
assign _218_ = _210_ & _217_ /*98937*/;
assign _30_ = _210_ ^ _217_ /*98938*/;
assign _215_ = _216_ | _218_ /*98935*/;
assign _224_ = ~D[31] /*98934*/;
assign _221_ = R_0[94] & _224_ /*98930*/;
assign _222_ = R_0[94] ^ _224_ /*98933*/;
assign _223_ = _215_ & _222_ /*98931*/;
assign _31_ = _215_ ^ _222_ /*98932*/;
assign _220_ = _221_ | _223_ /*98929*/;
assign _229_ = ~D[32] /*98928*/;
assign _226_ = R_0[95] & _229_ /*98924*/;
assign _227_ = R_0[95] ^ _229_ /*98927*/;
assign _228_ = _220_ & _227_ /*98925*/;
assign _32_ = _220_ ^ _227_ /*98926*/;
assign _225_ = _226_ | _228_ /*98923*/;
assign _234_ = ~D[33] /*98922*/;
assign _231_ = R_0[96] & _234_ /*98918*/;
assign _232_ = R_0[96] ^ _234_ /*98921*/;
assign _233_ = _225_ & _232_ /*98919*/;
assign _33_ = _225_ ^ _232_ /*98920*/;
assign _230_ = _231_ | _233_ /*98917*/;
assign _239_ = ~D[34] /*98916*/;
assign _236_ = R_0[97] & _239_ /*98912*/;
assign _237_ = R_0[97] ^ _239_ /*98915*/;
assign _238_ = _230_ & _237_ /*98913*/;
assign _34_ = _230_ ^ _237_ /*98914*/;
assign _235_ = _236_ | _238_ /*98911*/;
assign _244_ = ~D[35] /*98910*/;
assign _241_ = R_0[98] & _244_ /*98906*/;
assign _242_ = R_0[98] ^ _244_ /*98909*/;
assign _243_ = _235_ & _242_ /*98907*/;
assign _35_ = _235_ ^ _242_ /*98908*/;
assign _240_ = _241_ | _243_ /*98905*/;
assign _249_ = ~D[36] /*98904*/;
assign _246_ = R_0[99] & _249_ /*98900*/;
assign _247_ = R_0[99] ^ _249_ /*98903*/;
assign _248_ = _240_ & _247_ /*98901*/;
assign _36_ = _240_ ^ _247_ /*98902*/;
assign _245_ = _246_ | _248_ /*98899*/;
assign _254_ = ~D[37] /*98898*/;
assign _251_ = R_0[100] & _254_ /*98894*/;
assign _252_ = R_0[100] ^ _254_ /*98897*/;
assign _253_ = _245_ & _252_ /*98895*/;
assign _37_ = _245_ ^ _252_ /*98896*/;
assign _250_ = _251_ | _253_ /*98893*/;
assign _259_ = ~D[38] /*98892*/;
assign _256_ = R_0[101] & _259_ /*98888*/;
assign _257_ = R_0[101] ^ _259_ /*98891*/;
assign _258_ = _250_ & _257_ /*98889*/;
assign _38_ = _250_ ^ _257_ /*98890*/;
assign _255_ = _256_ | _258_ /*98887*/;
assign _264_ = ~D[39] /*98886*/;
assign _261_ = R_0[102] & _264_ /*98882*/;
assign _262_ = R_0[102] ^ _264_ /*98885*/;
assign _263_ = _255_ & _262_ /*98883*/;
assign _39_ = _255_ ^ _262_ /*98884*/;
assign _260_ = _261_ | _263_ /*98881*/;
assign _269_ = ~D[40] /*98880*/;
assign _266_ = R_0[103] & _269_ /*98876*/;
assign _267_ = R_0[103] ^ _269_ /*98879*/;
assign _268_ = _260_ & _267_ /*98877*/;
assign _40_ = _260_ ^ _267_ /*98878*/;
assign _265_ = _266_ | _268_ /*98875*/;
assign _274_ = ~D[41] /*98874*/;
assign _271_ = R_0[104] & _274_ /*98870*/;
assign _272_ = R_0[104] ^ _274_ /*98873*/;
assign _273_ = _265_ & _272_ /*98871*/;
assign _41_ = _265_ ^ _272_ /*98872*/;
assign _270_ = _271_ | _273_ /*98869*/;
assign _279_ = ~D[42] /*98868*/;
assign _276_ = R_0[105] & _279_ /*98864*/;
assign _277_ = R_0[105] ^ _279_ /*98867*/;
assign _278_ = _270_ & _277_ /*98865*/;
assign _42_ = _270_ ^ _277_ /*98866*/;
assign _275_ = _276_ | _278_ /*98863*/;
assign _284_ = ~D[43] /*98862*/;
assign _281_ = R_0[106] & _284_ /*98858*/;
assign _282_ = R_0[106] ^ _284_ /*98861*/;
assign _283_ = _275_ & _282_ /*98859*/;
assign _43_ = _275_ ^ _282_ /*98860*/;
assign _280_ = _281_ | _283_ /*98857*/;
assign _289_ = ~D[44] /*98856*/;
assign _286_ = R_0[107] & _289_ /*98852*/;
assign _287_ = R_0[107] ^ _289_ /*98855*/;
assign _288_ = _280_ & _287_ /*98853*/;
assign _44_ = _280_ ^ _287_ /*98854*/;
assign _285_ = _286_ | _288_ /*98851*/;
assign _294_ = ~D[45] /*98850*/;
assign _291_ = R_0[108] & _294_ /*98846*/;
assign _292_ = R_0[108] ^ _294_ /*98849*/;
assign _293_ = _285_ & _292_ /*98847*/;
assign _45_ = _285_ ^ _292_ /*98848*/;
assign _290_ = _291_ | _293_ /*98845*/;
assign _299_ = ~D[46] /*98844*/;
assign _296_ = R_0[109] & _299_ /*98840*/;
assign _297_ = R_0[109] ^ _299_ /*98843*/;
assign _298_ = _290_ & _297_ /*98841*/;
assign _46_ = _290_ ^ _297_ /*98842*/;
assign _295_ = _296_ | _298_ /*98839*/;
assign _304_ = ~D[47] /*98838*/;
assign _301_ = R_0[110] & _304_ /*98834*/;
assign _302_ = R_0[110] ^ _304_ /*98837*/;
assign _303_ = _295_ & _302_ /*98835*/;
assign _47_ = _295_ ^ _302_ /*98836*/;
assign _300_ = _301_ | _303_ /*98833*/;
assign _309_ = ~D[48] /*98832*/;
assign _306_ = R_0[111] & _309_ /*98828*/;
assign _307_ = R_0[111] ^ _309_ /*98831*/;
assign _308_ = _300_ & _307_ /*98829*/;
assign _48_ = _300_ ^ _307_ /*98830*/;
assign _305_ = _306_ | _308_ /*98827*/;
assign _314_ = ~D[49] /*98826*/;
assign _311_ = R_0[112] & _314_ /*98822*/;
assign _312_ = R_0[112] ^ _314_ /*98825*/;
assign _313_ = _305_ & _312_ /*98823*/;
assign _49_ = _305_ ^ _312_ /*98824*/;
assign _310_ = _311_ | _313_ /*98821*/;
assign _319_ = ~D[50] /*98820*/;
assign _316_ = R_0[113] & _319_ /*98816*/;
assign _317_ = R_0[113] ^ _319_ /*98819*/;
assign _318_ = _310_ & _317_ /*98817*/;
assign _50_ = _310_ ^ _317_ /*98818*/;
assign _315_ = _316_ | _318_ /*98815*/;
assign _324_ = ~D[51] /*98814*/;
assign _321_ = R_0[114] & _324_ /*98810*/;
assign _322_ = R_0[114] ^ _324_ /*98813*/;
assign _323_ = _315_ & _322_ /*98811*/;
assign _51_ = _315_ ^ _322_ /*98812*/;
assign _320_ = _321_ | _323_ /*98809*/;
assign _329_ = ~D[52] /*98808*/;
assign _326_ = R_0[115] & _329_ /*98804*/;
assign _327_ = R_0[115] ^ _329_ /*98807*/;
assign _328_ = _320_ & _327_ /*98805*/;
assign _52_ = _320_ ^ _327_ /*98806*/;
assign _325_ = _326_ | _328_ /*98803*/;
assign _334_ = ~D[53] /*98802*/;
assign _331_ = R_0[116] & _334_ /*98798*/;
assign _332_ = R_0[116] ^ _334_ /*98801*/;
assign _333_ = _325_ & _332_ /*98799*/;
assign _53_ = _325_ ^ _332_ /*98800*/;
assign _330_ = _331_ | _333_ /*98797*/;
assign _339_ = ~D[54] /*98796*/;
assign _336_ = R_0[117] & _339_ /*98792*/;
assign _337_ = R_0[117] ^ _339_ /*98795*/;
assign _338_ = _330_ & _337_ /*98793*/;
assign _54_ = _330_ ^ _337_ /*98794*/;
assign _335_ = _336_ | _338_ /*98791*/;
assign _344_ = ~D[55] /*98790*/;
assign _341_ = R_0[118] & _344_ /*98786*/;
assign _342_ = R_0[118] ^ _344_ /*98789*/;
assign _343_ = _335_ & _342_ /*98787*/;
assign _55_ = _335_ ^ _342_ /*98788*/;
assign _340_ = _341_ | _343_ /*98785*/;
assign _349_ = ~D[56] /*98784*/;
assign _346_ = R_0[119] & _349_ /*98780*/;
assign _347_ = R_0[119] ^ _349_ /*98783*/;
assign _348_ = _340_ & _347_ /*98781*/;
assign _56_ = _340_ ^ _347_ /*98782*/;
assign _345_ = _346_ | _348_ /*98779*/;
assign _354_ = ~D[57] /*98778*/;
assign _351_ = R_0[120] & _354_ /*98774*/;
assign _352_ = R_0[120] ^ _354_ /*98777*/;
assign _353_ = _345_ & _352_ /*98775*/;
assign _57_ = _345_ ^ _352_ /*98776*/;
assign _350_ = _351_ | _353_ /*98773*/;
assign _359_ = ~D[58] /*98772*/;
assign _356_ = R_0[121] & _359_ /*98768*/;
assign _357_ = R_0[121] ^ _359_ /*98771*/;
assign _358_ = _350_ & _357_ /*98769*/;
assign _58_ = _350_ ^ _357_ /*98770*/;
assign _355_ = _356_ | _358_ /*98767*/;
assign _364_ = ~D[59] /*98766*/;
assign _361_ = R_0[122] & _364_ /*98762*/;
assign _362_ = R_0[122] ^ _364_ /*98765*/;
assign _363_ = _355_ & _362_ /*98763*/;
assign _59_ = _355_ ^ _362_ /*98764*/;
assign _360_ = _361_ | _363_ /*98761*/;
assign _369_ = ~D[60] /*98760*/;
assign _366_ = R_0[123] & _369_ /*98756*/;
assign _367_ = R_0[123] ^ _369_ /*98759*/;
assign _368_ = _360_ & _367_ /*98757*/;
assign _60_ = _360_ ^ _367_ /*98758*/;
assign _365_ = _366_ | _368_ /*98755*/;
assign _374_ = ~D[61] /*98754*/;
assign _371_ = R_0[124] & _374_ /*98750*/;
assign _372_ = R_0[124] ^ _374_ /*98753*/;
assign _373_ = _365_ & _372_ /*98751*/;
assign _61_ = _365_ ^ _372_ /*98752*/;
assign _370_ = _371_ | _373_ /*98749*/;
assign _379_ = ~D[62] /*98748*/;
assign _376_ = R_0[125] & _379_ /*98744*/;
assign _377_ = R_0[125] ^ _379_ /*98747*/;
assign _378_ = _370_ & _377_ /*98745*/;
assign _62_ = _370_ ^ _377_ /*98746*/;
assign _375_ = _376_ | _378_ /*98743*/;
assign _380_ = zeroWire & oneWire /*98738*/;
assign _381_ = zeroWire ^ oneWire /*98741*/;
assign _382_ = _375_ & _381_ /*98739*/;
assign _63_ = _375_ ^ _381_ /*98740*/;
assign Q[63] = _380_ | _382_ /*98737*/;
assign _451_ = ~Q[63] /*98353*/;
assign _450_ = _451_ & D[0] /*98352*/;
assign _453_ = _0_ & _450_ /*98347*/;
assign _454_ = _0_ ^ _450_ /*98350*/;
assign _455_ = zeroWire & _454_ /*98348*/;
assign _385_ = zeroWire ^ _454_ /*98349*/;
assign _452_ = _453_ | _455_ /*98346*/;
assign _457_ = ~Q[63] /*98345*/;
assign _456_ = _457_ & D[1] /*98344*/;
assign _459_ = _1_ & _456_ /*98339*/;
assign _460_ = _1_ ^ _456_ /*98342*/;
assign _461_ = _452_ & _460_ /*98340*/;
assign _386_ = _452_ ^ _460_ /*98341*/;
assign _458_ = _459_ | _461_ /*98338*/;
assign _463_ = ~Q[63] /*98337*/;
assign _462_ = _463_ & D[2] /*98336*/;
assign _465_ = _2_ & _462_ /*98331*/;
assign _466_ = _2_ ^ _462_ /*98334*/;
assign _467_ = _458_ & _466_ /*98332*/;
assign _387_ = _458_ ^ _466_ /*98333*/;
assign _464_ = _465_ | _467_ /*98330*/;
assign _469_ = ~Q[63] /*98329*/;
assign _468_ = _469_ & D[3] /*98328*/;
assign _471_ = _3_ & _468_ /*98323*/;
assign _472_ = _3_ ^ _468_ /*98326*/;
assign _473_ = _464_ & _472_ /*98324*/;
assign _388_ = _464_ ^ _472_ /*98325*/;
assign _470_ = _471_ | _473_ /*98322*/;
assign _475_ = ~Q[63] /*98321*/;
assign _474_ = _475_ & D[4] /*98320*/;
assign _477_ = _4_ & _474_ /*98315*/;
assign _478_ = _4_ ^ _474_ /*98318*/;
assign _479_ = _470_ & _478_ /*98316*/;
assign _389_ = _470_ ^ _478_ /*98317*/;
assign _476_ = _477_ | _479_ /*98314*/;
assign _481_ = ~Q[63] /*98313*/;
assign _480_ = _481_ & D[5] /*98312*/;
assign _483_ = _5_ & _480_ /*98307*/;
assign _484_ = _5_ ^ _480_ /*98310*/;
assign _485_ = _476_ & _484_ /*98308*/;
assign _390_ = _476_ ^ _484_ /*98309*/;
assign _482_ = _483_ | _485_ /*98306*/;
assign _487_ = ~Q[63] /*98305*/;
assign _486_ = _487_ & D[6] /*98304*/;
assign _489_ = _6_ & _486_ /*98299*/;
assign _490_ = _6_ ^ _486_ /*98302*/;
assign _491_ = _482_ & _490_ /*98300*/;
assign _391_ = _482_ ^ _490_ /*98301*/;
assign _488_ = _489_ | _491_ /*98298*/;
assign _493_ = ~Q[63] /*98297*/;
assign _492_ = _493_ & D[7] /*98296*/;
assign _495_ = _7_ & _492_ /*98291*/;
assign _496_ = _7_ ^ _492_ /*98294*/;
assign _497_ = _488_ & _496_ /*98292*/;
assign _392_ = _488_ ^ _496_ /*98293*/;
assign _494_ = _495_ | _497_ /*98290*/;
assign _499_ = ~Q[63] /*98289*/;
assign _498_ = _499_ & D[8] /*98288*/;
assign _501_ = _8_ & _498_ /*98283*/;
assign _502_ = _8_ ^ _498_ /*98286*/;
assign _503_ = _494_ & _502_ /*98284*/;
assign _393_ = _494_ ^ _502_ /*98285*/;
assign _500_ = _501_ | _503_ /*98282*/;
assign _505_ = ~Q[63] /*98281*/;
assign _504_ = _505_ & D[9] /*98280*/;
assign _507_ = _9_ & _504_ /*98275*/;
assign _508_ = _9_ ^ _504_ /*98278*/;
assign _509_ = _500_ & _508_ /*98276*/;
assign _394_ = _500_ ^ _508_ /*98277*/;
assign _506_ = _507_ | _509_ /*98274*/;
assign _511_ = ~Q[63] /*98273*/;
assign _510_ = _511_ & D[10] /*98272*/;
assign _513_ = _10_ & _510_ /*98267*/;
assign _514_ = _10_ ^ _510_ /*98270*/;
assign _515_ = _506_ & _514_ /*98268*/;
assign _395_ = _506_ ^ _514_ /*98269*/;
assign _512_ = _513_ | _515_ /*98266*/;
assign _517_ = ~Q[63] /*98265*/;
assign _516_ = _517_ & D[11] /*98264*/;
assign _519_ = _11_ & _516_ /*98259*/;
assign _520_ = _11_ ^ _516_ /*98262*/;
assign _521_ = _512_ & _520_ /*98260*/;
assign _396_ = _512_ ^ _520_ /*98261*/;
assign _518_ = _519_ | _521_ /*98258*/;
assign _523_ = ~Q[63] /*98257*/;
assign _522_ = _523_ & D[12] /*98256*/;
assign _525_ = _12_ & _522_ /*98251*/;
assign _526_ = _12_ ^ _522_ /*98254*/;
assign _527_ = _518_ & _526_ /*98252*/;
assign _397_ = _518_ ^ _526_ /*98253*/;
assign _524_ = _525_ | _527_ /*98250*/;
assign _529_ = ~Q[63] /*98249*/;
assign _528_ = _529_ & D[13] /*98248*/;
assign _531_ = _13_ & _528_ /*98243*/;
assign _532_ = _13_ ^ _528_ /*98246*/;
assign _533_ = _524_ & _532_ /*98244*/;
assign _398_ = _524_ ^ _532_ /*98245*/;
assign _530_ = _531_ | _533_ /*98242*/;
assign _535_ = ~Q[63] /*98241*/;
assign _534_ = _535_ & D[14] /*98240*/;
assign _537_ = _14_ & _534_ /*98235*/;
assign _538_ = _14_ ^ _534_ /*98238*/;
assign _539_ = _530_ & _538_ /*98236*/;
assign _399_ = _530_ ^ _538_ /*98237*/;
assign _536_ = _537_ | _539_ /*98234*/;
assign _541_ = ~Q[63] /*98233*/;
assign _540_ = _541_ & D[15] /*98232*/;
assign _543_ = _15_ & _540_ /*98227*/;
assign _544_ = _15_ ^ _540_ /*98230*/;
assign _545_ = _536_ & _544_ /*98228*/;
assign _400_ = _536_ ^ _544_ /*98229*/;
assign _542_ = _543_ | _545_ /*98226*/;
assign _547_ = ~Q[63] /*98225*/;
assign _546_ = _547_ & D[16] /*98224*/;
assign _549_ = _16_ & _546_ /*98219*/;
assign _550_ = _16_ ^ _546_ /*98222*/;
assign _551_ = _542_ & _550_ /*98220*/;
assign _401_ = _542_ ^ _550_ /*98221*/;
assign _548_ = _549_ | _551_ /*98218*/;
assign _553_ = ~Q[63] /*98217*/;
assign _552_ = _553_ & D[17] /*98216*/;
assign _555_ = _17_ & _552_ /*98211*/;
assign _556_ = _17_ ^ _552_ /*98214*/;
assign _557_ = _548_ & _556_ /*98212*/;
assign _402_ = _548_ ^ _556_ /*98213*/;
assign _554_ = _555_ | _557_ /*98210*/;
assign _559_ = ~Q[63] /*98209*/;
assign _558_ = _559_ & D[18] /*98208*/;
assign _561_ = _18_ & _558_ /*98203*/;
assign _562_ = _18_ ^ _558_ /*98206*/;
assign _563_ = _554_ & _562_ /*98204*/;
assign _403_ = _554_ ^ _562_ /*98205*/;
assign _560_ = _561_ | _563_ /*98202*/;
assign _565_ = ~Q[63] /*98201*/;
assign _564_ = _565_ & D[19] /*98200*/;
assign _567_ = _19_ & _564_ /*98195*/;
assign _568_ = _19_ ^ _564_ /*98198*/;
assign _569_ = _560_ & _568_ /*98196*/;
assign _404_ = _560_ ^ _568_ /*98197*/;
assign _566_ = _567_ | _569_ /*98194*/;
assign _571_ = ~Q[63] /*98193*/;
assign _570_ = _571_ & D[20] /*98192*/;
assign _573_ = _20_ & _570_ /*98187*/;
assign _574_ = _20_ ^ _570_ /*98190*/;
assign _575_ = _566_ & _574_ /*98188*/;
assign _405_ = _566_ ^ _574_ /*98189*/;
assign _572_ = _573_ | _575_ /*98186*/;
assign _577_ = ~Q[63] /*98185*/;
assign _576_ = _577_ & D[21] /*98184*/;
assign _579_ = _21_ & _576_ /*98179*/;
assign _580_ = _21_ ^ _576_ /*98182*/;
assign _581_ = _572_ & _580_ /*98180*/;
assign _406_ = _572_ ^ _580_ /*98181*/;
assign _578_ = _579_ | _581_ /*98178*/;
assign _583_ = ~Q[63] /*98177*/;
assign _582_ = _583_ & D[22] /*98176*/;
assign _585_ = _22_ & _582_ /*98171*/;
assign _586_ = _22_ ^ _582_ /*98174*/;
assign _587_ = _578_ & _586_ /*98172*/;
assign _407_ = _578_ ^ _586_ /*98173*/;
assign _584_ = _585_ | _587_ /*98170*/;
assign _589_ = ~Q[63] /*98169*/;
assign _588_ = _589_ & D[23] /*98168*/;
assign _591_ = _23_ & _588_ /*98163*/;
assign _592_ = _23_ ^ _588_ /*98166*/;
assign _593_ = _584_ & _592_ /*98164*/;
assign _408_ = _584_ ^ _592_ /*98165*/;
assign _590_ = _591_ | _593_ /*98162*/;
assign _595_ = ~Q[63] /*98161*/;
assign _594_ = _595_ & D[24] /*98160*/;
assign _597_ = _24_ & _594_ /*98155*/;
assign _598_ = _24_ ^ _594_ /*98158*/;
assign _599_ = _590_ & _598_ /*98156*/;
assign _409_ = _590_ ^ _598_ /*98157*/;
assign _596_ = _597_ | _599_ /*98154*/;
assign _601_ = ~Q[63] /*98153*/;
assign _600_ = _601_ & D[25] /*98152*/;
assign _603_ = _25_ & _600_ /*98147*/;
assign _604_ = _25_ ^ _600_ /*98150*/;
assign _605_ = _596_ & _604_ /*98148*/;
assign _410_ = _596_ ^ _604_ /*98149*/;
assign _602_ = _603_ | _605_ /*98146*/;
assign _607_ = ~Q[63] /*98145*/;
assign _606_ = _607_ & D[26] /*98144*/;
assign _609_ = _26_ & _606_ /*98139*/;
assign _610_ = _26_ ^ _606_ /*98142*/;
assign _611_ = _602_ & _610_ /*98140*/;
assign _411_ = _602_ ^ _610_ /*98141*/;
assign _608_ = _609_ | _611_ /*98138*/;
assign _613_ = ~Q[63] /*98137*/;
assign _612_ = _613_ & D[27] /*98136*/;
assign _615_ = _27_ & _612_ /*98131*/;
assign _616_ = _27_ ^ _612_ /*98134*/;
assign _617_ = _608_ & _616_ /*98132*/;
assign _412_ = _608_ ^ _616_ /*98133*/;
assign _614_ = _615_ | _617_ /*98130*/;
assign _619_ = ~Q[63] /*98129*/;
assign _618_ = _619_ & D[28] /*98128*/;
assign _621_ = _28_ & _618_ /*98123*/;
assign _622_ = _28_ ^ _618_ /*98126*/;
assign _623_ = _614_ & _622_ /*98124*/;
assign _413_ = _614_ ^ _622_ /*98125*/;
assign _620_ = _621_ | _623_ /*98122*/;
assign _625_ = ~Q[63] /*98121*/;
assign _624_ = _625_ & D[29] /*98120*/;
assign _627_ = _29_ & _624_ /*98115*/;
assign _628_ = _29_ ^ _624_ /*98118*/;
assign _629_ = _620_ & _628_ /*98116*/;
assign _414_ = _620_ ^ _628_ /*98117*/;
assign _626_ = _627_ | _629_ /*98114*/;
assign _631_ = ~Q[63] /*98113*/;
assign _630_ = _631_ & D[30] /*98112*/;
assign _633_ = _30_ & _630_ /*98107*/;
assign _634_ = _30_ ^ _630_ /*98110*/;
assign _635_ = _626_ & _634_ /*98108*/;
assign _415_ = _626_ ^ _634_ /*98109*/;
assign _632_ = _633_ | _635_ /*98106*/;
assign _637_ = ~Q[63] /*98105*/;
assign _636_ = _637_ & D[31] /*98104*/;
assign _639_ = _31_ & _636_ /*98099*/;
assign _640_ = _31_ ^ _636_ /*98102*/;
assign _641_ = _632_ & _640_ /*98100*/;
assign _416_ = _632_ ^ _640_ /*98101*/;
assign _638_ = _639_ | _641_ /*98098*/;
assign _643_ = ~Q[63] /*98097*/;
assign _642_ = _643_ & D[32] /*98096*/;
assign _645_ = _32_ & _642_ /*98091*/;
assign _646_ = _32_ ^ _642_ /*98094*/;
assign _647_ = _638_ & _646_ /*98092*/;
assign _417_ = _638_ ^ _646_ /*98093*/;
assign _644_ = _645_ | _647_ /*98090*/;
assign _649_ = ~Q[63] /*98089*/;
assign _648_ = _649_ & D[33] /*98088*/;
assign _651_ = _33_ & _648_ /*98083*/;
assign _652_ = _33_ ^ _648_ /*98086*/;
assign _653_ = _644_ & _652_ /*98084*/;
assign _418_ = _644_ ^ _652_ /*98085*/;
assign _650_ = _651_ | _653_ /*98082*/;
assign _655_ = ~Q[63] /*98081*/;
assign _654_ = _655_ & D[34] /*98080*/;
assign _657_ = _34_ & _654_ /*98075*/;
assign _658_ = _34_ ^ _654_ /*98078*/;
assign _659_ = _650_ & _658_ /*98076*/;
assign _419_ = _650_ ^ _658_ /*98077*/;
assign _656_ = _657_ | _659_ /*98074*/;
assign _661_ = ~Q[63] /*98073*/;
assign _660_ = _661_ & D[35] /*98072*/;
assign _663_ = _35_ & _660_ /*98067*/;
assign _664_ = _35_ ^ _660_ /*98070*/;
assign _665_ = _656_ & _664_ /*98068*/;
assign _420_ = _656_ ^ _664_ /*98069*/;
assign _662_ = _663_ | _665_ /*98066*/;
assign _667_ = ~Q[63] /*98065*/;
assign _666_ = _667_ & D[36] /*98064*/;
assign _669_ = _36_ & _666_ /*98059*/;
assign _670_ = _36_ ^ _666_ /*98062*/;
assign _671_ = _662_ & _670_ /*98060*/;
assign _421_ = _662_ ^ _670_ /*98061*/;
assign _668_ = _669_ | _671_ /*98058*/;
assign _673_ = ~Q[63] /*98057*/;
assign _672_ = _673_ & D[37] /*98056*/;
assign _675_ = _37_ & _672_ /*98051*/;
assign _676_ = _37_ ^ _672_ /*98054*/;
assign _677_ = _668_ & _676_ /*98052*/;
assign _422_ = _668_ ^ _676_ /*98053*/;
assign _674_ = _675_ | _677_ /*98050*/;
assign _679_ = ~Q[63] /*98049*/;
assign _678_ = _679_ & D[38] /*98048*/;
assign _681_ = _38_ & _678_ /*98043*/;
assign _682_ = _38_ ^ _678_ /*98046*/;
assign _683_ = _674_ & _682_ /*98044*/;
assign _423_ = _674_ ^ _682_ /*98045*/;
assign _680_ = _681_ | _683_ /*98042*/;
assign _685_ = ~Q[63] /*98041*/;
assign _684_ = _685_ & D[39] /*98040*/;
assign _687_ = _39_ & _684_ /*98035*/;
assign _688_ = _39_ ^ _684_ /*98038*/;
assign _689_ = _680_ & _688_ /*98036*/;
assign _424_ = _680_ ^ _688_ /*98037*/;
assign _686_ = _687_ | _689_ /*98034*/;
assign _691_ = ~Q[63] /*98033*/;
assign _690_ = _691_ & D[40] /*98032*/;
assign _693_ = _40_ & _690_ /*98027*/;
assign _694_ = _40_ ^ _690_ /*98030*/;
assign _695_ = _686_ & _694_ /*98028*/;
assign _425_ = _686_ ^ _694_ /*98029*/;
assign _692_ = _693_ | _695_ /*98026*/;
assign _697_ = ~Q[63] /*98025*/;
assign _696_ = _697_ & D[41] /*98024*/;
assign _699_ = _41_ & _696_ /*98019*/;
assign _700_ = _41_ ^ _696_ /*98022*/;
assign _701_ = _692_ & _700_ /*98020*/;
assign _426_ = _692_ ^ _700_ /*98021*/;
assign _698_ = _699_ | _701_ /*98018*/;
assign _703_ = ~Q[63] /*98017*/;
assign _702_ = _703_ & D[42] /*98016*/;
assign _705_ = _42_ & _702_ /*98011*/;
assign _706_ = _42_ ^ _702_ /*98014*/;
assign _707_ = _698_ & _706_ /*98012*/;
assign _427_ = _698_ ^ _706_ /*98013*/;
assign _704_ = _705_ | _707_ /*98010*/;
assign _709_ = ~Q[63] /*98009*/;
assign _708_ = _709_ & D[43] /*98008*/;
assign _711_ = _43_ & _708_ /*98003*/;
assign _712_ = _43_ ^ _708_ /*98006*/;
assign _713_ = _704_ & _712_ /*98004*/;
assign _428_ = _704_ ^ _712_ /*98005*/;
assign _710_ = _711_ | _713_ /*98002*/;
assign _715_ = ~Q[63] /*98001*/;
assign _714_ = _715_ & D[44] /*98000*/;
assign _717_ = _44_ & _714_ /*97995*/;
assign _718_ = _44_ ^ _714_ /*97998*/;
assign _719_ = _710_ & _718_ /*97996*/;
assign _429_ = _710_ ^ _718_ /*97997*/;
assign _716_ = _717_ | _719_ /*97994*/;
assign _721_ = ~Q[63] /*97993*/;
assign _720_ = _721_ & D[45] /*97992*/;
assign _723_ = _45_ & _720_ /*97987*/;
assign _724_ = _45_ ^ _720_ /*97990*/;
assign _725_ = _716_ & _724_ /*97988*/;
assign _430_ = _716_ ^ _724_ /*97989*/;
assign _722_ = _723_ | _725_ /*97986*/;
assign _727_ = ~Q[63] /*97985*/;
assign _726_ = _727_ & D[46] /*97984*/;
assign _729_ = _46_ & _726_ /*97979*/;
assign _730_ = _46_ ^ _726_ /*97982*/;
assign _731_ = _722_ & _730_ /*97980*/;
assign _431_ = _722_ ^ _730_ /*97981*/;
assign _728_ = _729_ | _731_ /*97978*/;
assign _733_ = ~Q[63] /*97977*/;
assign _732_ = _733_ & D[47] /*97976*/;
assign _735_ = _47_ & _732_ /*97971*/;
assign _736_ = _47_ ^ _732_ /*97974*/;
assign _737_ = _728_ & _736_ /*97972*/;
assign _432_ = _728_ ^ _736_ /*97973*/;
assign _734_ = _735_ | _737_ /*97970*/;
assign _739_ = ~Q[63] /*97969*/;
assign _738_ = _739_ & D[48] /*97968*/;
assign _741_ = _48_ & _738_ /*97963*/;
assign _742_ = _48_ ^ _738_ /*97966*/;
assign _743_ = _734_ & _742_ /*97964*/;
assign _433_ = _734_ ^ _742_ /*97965*/;
assign _740_ = _741_ | _743_ /*97962*/;
assign _745_ = ~Q[63] /*97961*/;
assign _744_ = _745_ & D[49] /*97960*/;
assign _747_ = _49_ & _744_ /*97955*/;
assign _748_ = _49_ ^ _744_ /*97958*/;
assign _749_ = _740_ & _748_ /*97956*/;
assign _434_ = _740_ ^ _748_ /*97957*/;
assign _746_ = _747_ | _749_ /*97954*/;
assign _751_ = ~Q[63] /*97953*/;
assign _750_ = _751_ & D[50] /*97952*/;
assign _753_ = _50_ & _750_ /*97947*/;
assign _754_ = _50_ ^ _750_ /*97950*/;
assign _755_ = _746_ & _754_ /*97948*/;
assign _435_ = _746_ ^ _754_ /*97949*/;
assign _752_ = _753_ | _755_ /*97946*/;
assign _757_ = ~Q[63] /*97945*/;
assign _756_ = _757_ & D[51] /*97944*/;
assign _759_ = _51_ & _756_ /*97939*/;
assign _760_ = _51_ ^ _756_ /*97942*/;
assign _761_ = _752_ & _760_ /*97940*/;
assign _436_ = _752_ ^ _760_ /*97941*/;
assign _758_ = _759_ | _761_ /*97938*/;
assign _763_ = ~Q[63] /*97937*/;
assign _762_ = _763_ & D[52] /*97936*/;
assign _765_ = _52_ & _762_ /*97931*/;
assign _766_ = _52_ ^ _762_ /*97934*/;
assign _767_ = _758_ & _766_ /*97932*/;
assign _437_ = _758_ ^ _766_ /*97933*/;
assign _764_ = _765_ | _767_ /*97930*/;
assign _769_ = ~Q[63] /*97929*/;
assign _768_ = _769_ & D[53] /*97928*/;
assign _771_ = _53_ & _768_ /*97923*/;
assign _772_ = _53_ ^ _768_ /*97926*/;
assign _773_ = _764_ & _772_ /*97924*/;
assign _438_ = _764_ ^ _772_ /*97925*/;
assign _770_ = _771_ | _773_ /*97922*/;
assign _775_ = ~Q[63] /*97921*/;
assign _774_ = _775_ & D[54] /*97920*/;
assign _777_ = _54_ & _774_ /*97915*/;
assign _778_ = _54_ ^ _774_ /*97918*/;
assign _779_ = _770_ & _778_ /*97916*/;
assign _439_ = _770_ ^ _778_ /*97917*/;
assign _776_ = _777_ | _779_ /*97914*/;
assign _781_ = ~Q[63] /*97913*/;
assign _780_ = _781_ & D[55] /*97912*/;
assign _783_ = _55_ & _780_ /*97907*/;
assign _784_ = _55_ ^ _780_ /*97910*/;
assign _785_ = _776_ & _784_ /*97908*/;
assign _440_ = _776_ ^ _784_ /*97909*/;
assign _782_ = _783_ | _785_ /*97906*/;
assign _787_ = ~Q[63] /*97905*/;
assign _786_ = _787_ & D[56] /*97904*/;
assign _789_ = _56_ & _786_ /*97899*/;
assign _790_ = _56_ ^ _786_ /*97902*/;
assign _791_ = _782_ & _790_ /*97900*/;
assign _441_ = _782_ ^ _790_ /*97901*/;
assign _788_ = _789_ | _791_ /*97898*/;
assign _793_ = ~Q[63] /*97897*/;
assign _792_ = _793_ & D[57] /*97896*/;
assign _795_ = _57_ & _792_ /*97891*/;
assign _796_ = _57_ ^ _792_ /*97894*/;
assign _797_ = _788_ & _796_ /*97892*/;
assign _442_ = _788_ ^ _796_ /*97893*/;
assign _794_ = _795_ | _797_ /*97890*/;
assign _799_ = ~Q[63] /*97889*/;
assign _798_ = _799_ & D[58] /*97888*/;
assign _801_ = _58_ & _798_ /*97883*/;
assign _802_ = _58_ ^ _798_ /*97886*/;
assign _803_ = _794_ & _802_ /*97884*/;
assign _443_ = _794_ ^ _802_ /*97885*/;
assign _800_ = _801_ | _803_ /*97882*/;
assign _805_ = ~Q[63] /*97881*/;
assign _804_ = _805_ & D[59] /*97880*/;
assign _807_ = _59_ & _804_ /*97875*/;
assign _808_ = _59_ ^ _804_ /*97878*/;
assign _809_ = _800_ & _808_ /*97876*/;
assign _444_ = _800_ ^ _808_ /*97877*/;
assign _806_ = _807_ | _809_ /*97874*/;
assign _811_ = ~Q[63] /*97873*/;
assign _810_ = _811_ & D[60] /*97872*/;
assign _813_ = _60_ & _810_ /*97867*/;
assign _814_ = _60_ ^ _810_ /*97870*/;
assign _815_ = _806_ & _814_ /*97868*/;
assign _445_ = _806_ ^ _814_ /*97869*/;
assign _812_ = _813_ | _815_ /*97866*/;
assign _817_ = ~Q[63] /*97865*/;
assign _816_ = _817_ & D[61] /*97864*/;
assign _819_ = _61_ & _816_ /*97859*/;
assign _820_ = _61_ ^ _816_ /*97862*/;
assign _821_ = _812_ & _820_ /*97860*/;
assign _446_ = _812_ ^ _820_ /*97861*/;
assign _818_ = _819_ | _821_ /*97858*/;
assign _823_ = ~Q[63] /*97857*/;
assign _822_ = _823_ & D[62] /*97856*/;
assign _825_ = _62_ & _822_ /*97851*/;
assign _826_ = _62_ ^ _822_ /*97854*/;
assign _827_ = _818_ & _826_ /*97852*/;
assign _447_ = _818_ ^ _826_ /*97853*/;
assign _824_ = _825_ | _827_ /*97850*/;
assign _829_ = ~Q[63] /*97849*/;
assign _828_ = _829_ & zeroWire /*97848*/;
assign _830_ = _63_ ^ _828_ /*97846*/;
assign _448_ = _830_ ^ _824_ /*97845*/;
assign _901_ = ~D[0] /*97591*/;
assign _898_ = R_0[62] & _901_ /*97587*/;
assign _899_ = R_0[62] ^ _901_ /*97590*/;
assign _900_ = oneWire & _899_ /*97588*/;
assign _833_ = oneWire ^ _899_ /*97589*/;
assign _897_ = _898_ | _900_ /*97586*/;
assign _906_ = ~D[1] /*97585*/;
assign _903_ = _385_ & _906_ /*97581*/;
assign _904_ = _385_ ^ _906_ /*97584*/;
assign _905_ = _897_ & _904_ /*97582*/;
assign _834_ = _897_ ^ _904_ /*97583*/;
assign _902_ = _903_ | _905_ /*97580*/;
assign _911_ = ~D[2] /*97579*/;
assign _908_ = _386_ & _911_ /*97575*/;
assign _909_ = _386_ ^ _911_ /*97578*/;
assign _910_ = _902_ & _909_ /*97576*/;
assign _835_ = _902_ ^ _909_ /*97577*/;
assign _907_ = _908_ | _910_ /*97574*/;
assign _916_ = ~D[3] /*97573*/;
assign _913_ = _387_ & _916_ /*97569*/;
assign _914_ = _387_ ^ _916_ /*97572*/;
assign _915_ = _907_ & _914_ /*97570*/;
assign _836_ = _907_ ^ _914_ /*97571*/;
assign _912_ = _913_ | _915_ /*97568*/;
assign _921_ = ~D[4] /*97567*/;
assign _918_ = _388_ & _921_ /*97563*/;
assign _919_ = _388_ ^ _921_ /*97566*/;
assign _920_ = _912_ & _919_ /*97564*/;
assign _837_ = _912_ ^ _919_ /*97565*/;
assign _917_ = _918_ | _920_ /*97562*/;
assign _926_ = ~D[5] /*97561*/;
assign _923_ = _389_ & _926_ /*97557*/;
assign _924_ = _389_ ^ _926_ /*97560*/;
assign _925_ = _917_ & _924_ /*97558*/;
assign _838_ = _917_ ^ _924_ /*97559*/;
assign _922_ = _923_ | _925_ /*97556*/;
assign _931_ = ~D[6] /*97555*/;
assign _928_ = _390_ & _931_ /*97551*/;
assign _929_ = _390_ ^ _931_ /*97554*/;
assign _930_ = _922_ & _929_ /*97552*/;
assign _839_ = _922_ ^ _929_ /*97553*/;
assign _927_ = _928_ | _930_ /*97550*/;
assign _936_ = ~D[7] /*97549*/;
assign _933_ = _391_ & _936_ /*97545*/;
assign _934_ = _391_ ^ _936_ /*97548*/;
assign _935_ = _927_ & _934_ /*97546*/;
assign _840_ = _927_ ^ _934_ /*97547*/;
assign _932_ = _933_ | _935_ /*97544*/;
assign _941_ = ~D[8] /*97543*/;
assign _938_ = _392_ & _941_ /*97539*/;
assign _939_ = _392_ ^ _941_ /*97542*/;
assign _940_ = _932_ & _939_ /*97540*/;
assign _841_ = _932_ ^ _939_ /*97541*/;
assign _937_ = _938_ | _940_ /*97538*/;
assign _946_ = ~D[9] /*97537*/;
assign _943_ = _393_ & _946_ /*97533*/;
assign _944_ = _393_ ^ _946_ /*97536*/;
assign _945_ = _937_ & _944_ /*97534*/;
assign _842_ = _937_ ^ _944_ /*97535*/;
assign _942_ = _943_ | _945_ /*97532*/;
assign _951_ = ~D[10] /*97531*/;
assign _948_ = _394_ & _951_ /*97527*/;
assign _949_ = _394_ ^ _951_ /*97530*/;
assign _950_ = _942_ & _949_ /*97528*/;
assign _843_ = _942_ ^ _949_ /*97529*/;
assign _947_ = _948_ | _950_ /*97526*/;
assign _956_ = ~D[11] /*97525*/;
assign _953_ = _395_ & _956_ /*97521*/;
assign _954_ = _395_ ^ _956_ /*97524*/;
assign _955_ = _947_ & _954_ /*97522*/;
assign _844_ = _947_ ^ _954_ /*97523*/;
assign _952_ = _953_ | _955_ /*97520*/;
assign _961_ = ~D[12] /*97519*/;
assign _958_ = _396_ & _961_ /*97515*/;
assign _959_ = _396_ ^ _961_ /*97518*/;
assign _960_ = _952_ & _959_ /*97516*/;
assign _845_ = _952_ ^ _959_ /*97517*/;
assign _957_ = _958_ | _960_ /*97514*/;
assign _966_ = ~D[13] /*97513*/;
assign _963_ = _397_ & _966_ /*97509*/;
assign _964_ = _397_ ^ _966_ /*97512*/;
assign _965_ = _957_ & _964_ /*97510*/;
assign _846_ = _957_ ^ _964_ /*97511*/;
assign _962_ = _963_ | _965_ /*97508*/;
assign _971_ = ~D[14] /*97507*/;
assign _968_ = _398_ & _971_ /*97503*/;
assign _969_ = _398_ ^ _971_ /*97506*/;
assign _970_ = _962_ & _969_ /*97504*/;
assign _847_ = _962_ ^ _969_ /*97505*/;
assign _967_ = _968_ | _970_ /*97502*/;
assign _976_ = ~D[15] /*97501*/;
assign _973_ = _399_ & _976_ /*97497*/;
assign _974_ = _399_ ^ _976_ /*97500*/;
assign _975_ = _967_ & _974_ /*97498*/;
assign _848_ = _967_ ^ _974_ /*97499*/;
assign _972_ = _973_ | _975_ /*97496*/;
assign _981_ = ~D[16] /*97495*/;
assign _978_ = _400_ & _981_ /*97491*/;
assign _979_ = _400_ ^ _981_ /*97494*/;
assign _980_ = _972_ & _979_ /*97492*/;
assign _849_ = _972_ ^ _979_ /*97493*/;
assign _977_ = _978_ | _980_ /*97490*/;
assign _986_ = ~D[17] /*97489*/;
assign _983_ = _401_ & _986_ /*97485*/;
assign _984_ = _401_ ^ _986_ /*97488*/;
assign _985_ = _977_ & _984_ /*97486*/;
assign _850_ = _977_ ^ _984_ /*97487*/;
assign _982_ = _983_ | _985_ /*97484*/;
assign _991_ = ~D[18] /*97483*/;
assign _988_ = _402_ & _991_ /*97479*/;
assign _989_ = _402_ ^ _991_ /*97482*/;
assign _990_ = _982_ & _989_ /*97480*/;
assign _851_ = _982_ ^ _989_ /*97481*/;
assign _987_ = _988_ | _990_ /*97478*/;
assign _996_ = ~D[19] /*97477*/;
assign _993_ = _403_ & _996_ /*97473*/;
assign _994_ = _403_ ^ _996_ /*97476*/;
assign _995_ = _987_ & _994_ /*97474*/;
assign _852_ = _987_ ^ _994_ /*97475*/;
assign _992_ = _993_ | _995_ /*97472*/;
assign _1001_ = ~D[20] /*97471*/;
assign _998_ = _404_ & _1001_ /*97467*/;
assign _999_ = _404_ ^ _1001_ /*97470*/;
assign _1000_ = _992_ & _999_ /*97468*/;
assign _853_ = _992_ ^ _999_ /*97469*/;
assign _997_ = _998_ | _1000_ /*97466*/;
assign _1006_ = ~D[21] /*97465*/;
assign _1003_ = _405_ & _1006_ /*97461*/;
assign _1004_ = _405_ ^ _1006_ /*97464*/;
assign _1005_ = _997_ & _1004_ /*97462*/;
assign _854_ = _997_ ^ _1004_ /*97463*/;
assign _1002_ = _1003_ | _1005_ /*97460*/;
assign _1011_ = ~D[22] /*97459*/;
assign _1008_ = _406_ & _1011_ /*97455*/;
assign _1009_ = _406_ ^ _1011_ /*97458*/;
assign _1010_ = _1002_ & _1009_ /*97456*/;
assign _855_ = _1002_ ^ _1009_ /*97457*/;
assign _1007_ = _1008_ | _1010_ /*97454*/;
assign _1016_ = ~D[23] /*97453*/;
assign _1013_ = _407_ & _1016_ /*97449*/;
assign _1014_ = _407_ ^ _1016_ /*97452*/;
assign _1015_ = _1007_ & _1014_ /*97450*/;
assign _856_ = _1007_ ^ _1014_ /*97451*/;
assign _1012_ = _1013_ | _1015_ /*97448*/;
assign _1021_ = ~D[24] /*97447*/;
assign _1018_ = _408_ & _1021_ /*97443*/;
assign _1019_ = _408_ ^ _1021_ /*97446*/;
assign _1020_ = _1012_ & _1019_ /*97444*/;
assign _857_ = _1012_ ^ _1019_ /*97445*/;
assign _1017_ = _1018_ | _1020_ /*97442*/;
assign _1026_ = ~D[25] /*97441*/;
assign _1023_ = _409_ & _1026_ /*97437*/;
assign _1024_ = _409_ ^ _1026_ /*97440*/;
assign _1025_ = _1017_ & _1024_ /*97438*/;
assign _858_ = _1017_ ^ _1024_ /*97439*/;
assign _1022_ = _1023_ | _1025_ /*97436*/;
assign _1031_ = ~D[26] /*97435*/;
assign _1028_ = _410_ & _1031_ /*97431*/;
assign _1029_ = _410_ ^ _1031_ /*97434*/;
assign _1030_ = _1022_ & _1029_ /*97432*/;
assign _859_ = _1022_ ^ _1029_ /*97433*/;
assign _1027_ = _1028_ | _1030_ /*97430*/;
assign _1036_ = ~D[27] /*97429*/;
assign _1033_ = _411_ & _1036_ /*97425*/;
assign _1034_ = _411_ ^ _1036_ /*97428*/;
assign _1035_ = _1027_ & _1034_ /*97426*/;
assign _860_ = _1027_ ^ _1034_ /*97427*/;
assign _1032_ = _1033_ | _1035_ /*97424*/;
assign _1041_ = ~D[28] /*97423*/;
assign _1038_ = _412_ & _1041_ /*97419*/;
assign _1039_ = _412_ ^ _1041_ /*97422*/;
assign _1040_ = _1032_ & _1039_ /*97420*/;
assign _861_ = _1032_ ^ _1039_ /*97421*/;
assign _1037_ = _1038_ | _1040_ /*97418*/;
assign _1046_ = ~D[29] /*97417*/;
assign _1043_ = _413_ & _1046_ /*97413*/;
assign _1044_ = _413_ ^ _1046_ /*97416*/;
assign _1045_ = _1037_ & _1044_ /*97414*/;
assign _862_ = _1037_ ^ _1044_ /*97415*/;
assign _1042_ = _1043_ | _1045_ /*97412*/;
assign _1051_ = ~D[30] /*97411*/;
assign _1048_ = _414_ & _1051_ /*97407*/;
assign _1049_ = _414_ ^ _1051_ /*97410*/;
assign _1050_ = _1042_ & _1049_ /*97408*/;
assign _863_ = _1042_ ^ _1049_ /*97409*/;
assign _1047_ = _1048_ | _1050_ /*97406*/;
assign _1056_ = ~D[31] /*97405*/;
assign _1053_ = _415_ & _1056_ /*97401*/;
assign _1054_ = _415_ ^ _1056_ /*97404*/;
assign _1055_ = _1047_ & _1054_ /*97402*/;
assign _864_ = _1047_ ^ _1054_ /*97403*/;
assign _1052_ = _1053_ | _1055_ /*97400*/;
assign _1061_ = ~D[32] /*97399*/;
assign _1058_ = _416_ & _1061_ /*97395*/;
assign _1059_ = _416_ ^ _1061_ /*97398*/;
assign _1060_ = _1052_ & _1059_ /*97396*/;
assign _865_ = _1052_ ^ _1059_ /*97397*/;
assign _1057_ = _1058_ | _1060_ /*97394*/;
assign _1066_ = ~D[33] /*97393*/;
assign _1063_ = _417_ & _1066_ /*97389*/;
assign _1064_ = _417_ ^ _1066_ /*97392*/;
assign _1065_ = _1057_ & _1064_ /*97390*/;
assign _866_ = _1057_ ^ _1064_ /*97391*/;
assign _1062_ = _1063_ | _1065_ /*97388*/;
assign _1071_ = ~D[34] /*97387*/;
assign _1068_ = _418_ & _1071_ /*97383*/;
assign _1069_ = _418_ ^ _1071_ /*97386*/;
assign _1070_ = _1062_ & _1069_ /*97384*/;
assign _867_ = _1062_ ^ _1069_ /*97385*/;
assign _1067_ = _1068_ | _1070_ /*97382*/;
assign _1076_ = ~D[35] /*97381*/;
assign _1073_ = _419_ & _1076_ /*97377*/;
assign _1074_ = _419_ ^ _1076_ /*97380*/;
assign _1075_ = _1067_ & _1074_ /*97378*/;
assign _868_ = _1067_ ^ _1074_ /*97379*/;
assign _1072_ = _1073_ | _1075_ /*97376*/;
assign _1081_ = ~D[36] /*97375*/;
assign _1078_ = _420_ & _1081_ /*97371*/;
assign _1079_ = _420_ ^ _1081_ /*97374*/;
assign _1080_ = _1072_ & _1079_ /*97372*/;
assign _869_ = _1072_ ^ _1079_ /*97373*/;
assign _1077_ = _1078_ | _1080_ /*97370*/;
assign _1086_ = ~D[37] /*97369*/;
assign _1083_ = _421_ & _1086_ /*97365*/;
assign _1084_ = _421_ ^ _1086_ /*97368*/;
assign _1085_ = _1077_ & _1084_ /*97366*/;
assign _870_ = _1077_ ^ _1084_ /*97367*/;
assign _1082_ = _1083_ | _1085_ /*97364*/;
assign _1091_ = ~D[38] /*97363*/;
assign _1088_ = _422_ & _1091_ /*97359*/;
assign _1089_ = _422_ ^ _1091_ /*97362*/;
assign _1090_ = _1082_ & _1089_ /*97360*/;
assign _871_ = _1082_ ^ _1089_ /*97361*/;
assign _1087_ = _1088_ | _1090_ /*97358*/;
assign _1096_ = ~D[39] /*97357*/;
assign _1093_ = _423_ & _1096_ /*97353*/;
assign _1094_ = _423_ ^ _1096_ /*97356*/;
assign _1095_ = _1087_ & _1094_ /*97354*/;
assign _872_ = _1087_ ^ _1094_ /*97355*/;
assign _1092_ = _1093_ | _1095_ /*97352*/;
assign _1101_ = ~D[40] /*97351*/;
assign _1098_ = _424_ & _1101_ /*97347*/;
assign _1099_ = _424_ ^ _1101_ /*97350*/;
assign _1100_ = _1092_ & _1099_ /*97348*/;
assign _873_ = _1092_ ^ _1099_ /*97349*/;
assign _1097_ = _1098_ | _1100_ /*97346*/;
assign _1106_ = ~D[41] /*97345*/;
assign _1103_ = _425_ & _1106_ /*97341*/;
assign _1104_ = _425_ ^ _1106_ /*97344*/;
assign _1105_ = _1097_ & _1104_ /*97342*/;
assign _874_ = _1097_ ^ _1104_ /*97343*/;
assign _1102_ = _1103_ | _1105_ /*97340*/;
assign _1111_ = ~D[42] /*97339*/;
assign _1108_ = _426_ & _1111_ /*97335*/;
assign _1109_ = _426_ ^ _1111_ /*97338*/;
assign _1110_ = _1102_ & _1109_ /*97336*/;
assign _875_ = _1102_ ^ _1109_ /*97337*/;
assign _1107_ = _1108_ | _1110_ /*97334*/;
assign _1116_ = ~D[43] /*97333*/;
assign _1113_ = _427_ & _1116_ /*97329*/;
assign _1114_ = _427_ ^ _1116_ /*97332*/;
assign _1115_ = _1107_ & _1114_ /*97330*/;
assign _876_ = _1107_ ^ _1114_ /*97331*/;
assign _1112_ = _1113_ | _1115_ /*97328*/;
assign _1121_ = ~D[44] /*97327*/;
assign _1118_ = _428_ & _1121_ /*97323*/;
assign _1119_ = _428_ ^ _1121_ /*97326*/;
assign _1120_ = _1112_ & _1119_ /*97324*/;
assign _877_ = _1112_ ^ _1119_ /*97325*/;
assign _1117_ = _1118_ | _1120_ /*97322*/;
assign _1126_ = ~D[45] /*97321*/;
assign _1123_ = _429_ & _1126_ /*97317*/;
assign _1124_ = _429_ ^ _1126_ /*97320*/;
assign _1125_ = _1117_ & _1124_ /*97318*/;
assign _878_ = _1117_ ^ _1124_ /*97319*/;
assign _1122_ = _1123_ | _1125_ /*97316*/;
assign _1131_ = ~D[46] /*97315*/;
assign _1128_ = _430_ & _1131_ /*97311*/;
assign _1129_ = _430_ ^ _1131_ /*97314*/;
assign _1130_ = _1122_ & _1129_ /*97312*/;
assign _879_ = _1122_ ^ _1129_ /*97313*/;
assign _1127_ = _1128_ | _1130_ /*97310*/;
assign _1136_ = ~D[47] /*97309*/;
assign _1133_ = _431_ & _1136_ /*97305*/;
assign _1134_ = _431_ ^ _1136_ /*97308*/;
assign _1135_ = _1127_ & _1134_ /*97306*/;
assign _880_ = _1127_ ^ _1134_ /*97307*/;
assign _1132_ = _1133_ | _1135_ /*97304*/;
assign _1141_ = ~D[48] /*97303*/;
assign _1138_ = _432_ & _1141_ /*97299*/;
assign _1139_ = _432_ ^ _1141_ /*97302*/;
assign _1140_ = _1132_ & _1139_ /*97300*/;
assign _881_ = _1132_ ^ _1139_ /*97301*/;
assign _1137_ = _1138_ | _1140_ /*97298*/;
assign _1146_ = ~D[49] /*97297*/;
assign _1143_ = _433_ & _1146_ /*97293*/;
assign _1144_ = _433_ ^ _1146_ /*97296*/;
assign _1145_ = _1137_ & _1144_ /*97294*/;
assign _882_ = _1137_ ^ _1144_ /*97295*/;
assign _1142_ = _1143_ | _1145_ /*97292*/;
assign _1151_ = ~D[50] /*97291*/;
assign _1148_ = _434_ & _1151_ /*97287*/;
assign _1149_ = _434_ ^ _1151_ /*97290*/;
assign _1150_ = _1142_ & _1149_ /*97288*/;
assign _883_ = _1142_ ^ _1149_ /*97289*/;
assign _1147_ = _1148_ | _1150_ /*97286*/;
assign _1156_ = ~D[51] /*97285*/;
assign _1153_ = _435_ & _1156_ /*97281*/;
assign _1154_ = _435_ ^ _1156_ /*97284*/;
assign _1155_ = _1147_ & _1154_ /*97282*/;
assign _884_ = _1147_ ^ _1154_ /*97283*/;
assign _1152_ = _1153_ | _1155_ /*97280*/;
assign _1161_ = ~D[52] /*97279*/;
assign _1158_ = _436_ & _1161_ /*97275*/;
assign _1159_ = _436_ ^ _1161_ /*97278*/;
assign _1160_ = _1152_ & _1159_ /*97276*/;
assign _885_ = _1152_ ^ _1159_ /*97277*/;
assign _1157_ = _1158_ | _1160_ /*97274*/;
assign _1166_ = ~D[53] /*97273*/;
assign _1163_ = _437_ & _1166_ /*97269*/;
assign _1164_ = _437_ ^ _1166_ /*97272*/;
assign _1165_ = _1157_ & _1164_ /*97270*/;
assign _886_ = _1157_ ^ _1164_ /*97271*/;
assign _1162_ = _1163_ | _1165_ /*97268*/;
assign _1171_ = ~D[54] /*97267*/;
assign _1168_ = _438_ & _1171_ /*97263*/;
assign _1169_ = _438_ ^ _1171_ /*97266*/;
assign _1170_ = _1162_ & _1169_ /*97264*/;
assign _887_ = _1162_ ^ _1169_ /*97265*/;
assign _1167_ = _1168_ | _1170_ /*97262*/;
assign _1176_ = ~D[55] /*97261*/;
assign _1173_ = _439_ & _1176_ /*97257*/;
assign _1174_ = _439_ ^ _1176_ /*97260*/;
assign _1175_ = _1167_ & _1174_ /*97258*/;
assign _888_ = _1167_ ^ _1174_ /*97259*/;
assign _1172_ = _1173_ | _1175_ /*97256*/;
assign _1181_ = ~D[56] /*97255*/;
assign _1178_ = _440_ & _1181_ /*97251*/;
assign _1179_ = _440_ ^ _1181_ /*97254*/;
assign _1180_ = _1172_ & _1179_ /*97252*/;
assign _889_ = _1172_ ^ _1179_ /*97253*/;
assign _1177_ = _1178_ | _1180_ /*97250*/;
assign _1186_ = ~D[57] /*97249*/;
assign _1183_ = _441_ & _1186_ /*97245*/;
assign _1184_ = _441_ ^ _1186_ /*97248*/;
assign _1185_ = _1177_ & _1184_ /*97246*/;
assign _890_ = _1177_ ^ _1184_ /*97247*/;
assign _1182_ = _1183_ | _1185_ /*97244*/;
assign _1191_ = ~D[58] /*97243*/;
assign _1188_ = _442_ & _1191_ /*97239*/;
assign _1189_ = _442_ ^ _1191_ /*97242*/;
assign _1190_ = _1182_ & _1189_ /*97240*/;
assign _891_ = _1182_ ^ _1189_ /*97241*/;
assign _1187_ = _1188_ | _1190_ /*97238*/;
assign _1196_ = ~D[59] /*97237*/;
assign _1193_ = _443_ & _1196_ /*97233*/;
assign _1194_ = _443_ ^ _1196_ /*97236*/;
assign _1195_ = _1187_ & _1194_ /*97234*/;
assign _892_ = _1187_ ^ _1194_ /*97235*/;
assign _1192_ = _1193_ | _1195_ /*97232*/;
assign _1201_ = ~D[60] /*97231*/;
assign _1198_ = _444_ & _1201_ /*97227*/;
assign _1199_ = _444_ ^ _1201_ /*97230*/;
assign _1200_ = _1192_ & _1199_ /*97228*/;
assign _893_ = _1192_ ^ _1199_ /*97229*/;
assign _1197_ = _1198_ | _1200_ /*97226*/;
assign _1206_ = ~D[61] /*97225*/;
assign _1203_ = _445_ & _1206_ /*97221*/;
assign _1204_ = _445_ ^ _1206_ /*97224*/;
assign _1205_ = _1197_ & _1204_ /*97222*/;
assign _894_ = _1197_ ^ _1204_ /*97223*/;
assign _1202_ = _1203_ | _1205_ /*97220*/;
assign _1211_ = ~D[62] /*97219*/;
assign _1208_ = _446_ & _1211_ /*97215*/;
assign _1209_ = _446_ ^ _1211_ /*97218*/;
assign _1210_ = _1202_ & _1209_ /*97216*/;
assign _895_ = _1202_ ^ _1209_ /*97217*/;
assign _1207_ = _1208_ | _1210_ /*97214*/;
assign _1212_ = _447_ & oneWire /*97209*/;
assign _1213_ = _447_ ^ oneWire /*97212*/;
assign _1214_ = _1207_ & _1213_ /*97210*/;
assign _896_ = _1207_ ^ _1213_ /*97211*/;
assign Q[62] = _1212_ | _1214_ /*97208*/;
assign _1347_ = ~Q[62] /*96823*/;
assign _1346_ = _1347_ & D[0] /*96822*/;
assign _1349_ = _833_ & _1346_ /*96817*/;
assign _1350_ = _833_ ^ _1346_ /*96820*/;
assign _1351_ = zeroWire & _1350_ /*96818*/;
assign _1281_ = zeroWire ^ _1350_ /*96819*/;
assign _1348_ = _1349_ | _1351_ /*96816*/;
assign _1353_ = ~Q[62] /*96815*/;
assign _1352_ = _1353_ & D[1] /*96814*/;
assign _1355_ = _834_ & _1352_ /*96809*/;
assign _1356_ = _834_ ^ _1352_ /*96812*/;
assign _1357_ = _1348_ & _1356_ /*96810*/;
assign _1282_ = _1348_ ^ _1356_ /*96811*/;
assign _1354_ = _1355_ | _1357_ /*96808*/;
assign _1359_ = ~Q[62] /*96807*/;
assign _1358_ = _1359_ & D[2] /*96806*/;
assign _1361_ = _835_ & _1358_ /*96801*/;
assign _1362_ = _835_ ^ _1358_ /*96804*/;
assign _1363_ = _1354_ & _1362_ /*96802*/;
assign _1283_ = _1354_ ^ _1362_ /*96803*/;
assign _1360_ = _1361_ | _1363_ /*96800*/;
assign _1365_ = ~Q[62] /*96799*/;
assign _1364_ = _1365_ & D[3] /*96798*/;
assign _1367_ = _836_ & _1364_ /*96793*/;
assign _1368_ = _836_ ^ _1364_ /*96796*/;
assign _1369_ = _1360_ & _1368_ /*96794*/;
assign _1284_ = _1360_ ^ _1368_ /*96795*/;
assign _1366_ = _1367_ | _1369_ /*96792*/;
assign _1371_ = ~Q[62] /*96791*/;
assign _1370_ = _1371_ & D[4] /*96790*/;
assign _1373_ = _837_ & _1370_ /*96785*/;
assign _1374_ = _837_ ^ _1370_ /*96788*/;
assign _1375_ = _1366_ & _1374_ /*96786*/;
assign _1285_ = _1366_ ^ _1374_ /*96787*/;
assign _1372_ = _1373_ | _1375_ /*96784*/;
assign _1377_ = ~Q[62] /*96783*/;
assign _1376_ = _1377_ & D[5] /*96782*/;
assign _1379_ = _838_ & _1376_ /*96777*/;
assign _1380_ = _838_ ^ _1376_ /*96780*/;
assign _1381_ = _1372_ & _1380_ /*96778*/;
assign _1286_ = _1372_ ^ _1380_ /*96779*/;
assign _1378_ = _1379_ | _1381_ /*96776*/;
assign _1383_ = ~Q[62] /*96775*/;
assign _1382_ = _1383_ & D[6] /*96774*/;
assign _1385_ = _839_ & _1382_ /*96769*/;
assign _1386_ = _839_ ^ _1382_ /*96772*/;
assign _1387_ = _1378_ & _1386_ /*96770*/;
assign _1287_ = _1378_ ^ _1386_ /*96771*/;
assign _1384_ = _1385_ | _1387_ /*96768*/;
assign _1389_ = ~Q[62] /*96767*/;
assign _1388_ = _1389_ & D[7] /*96766*/;
assign _1391_ = _840_ & _1388_ /*96761*/;
assign _1392_ = _840_ ^ _1388_ /*96764*/;
assign _1393_ = _1384_ & _1392_ /*96762*/;
assign _1288_ = _1384_ ^ _1392_ /*96763*/;
assign _1390_ = _1391_ | _1393_ /*96760*/;
assign _1395_ = ~Q[62] /*96759*/;
assign _1394_ = _1395_ & D[8] /*96758*/;
assign _1397_ = _841_ & _1394_ /*96753*/;
assign _1398_ = _841_ ^ _1394_ /*96756*/;
assign _1399_ = _1390_ & _1398_ /*96754*/;
assign _1289_ = _1390_ ^ _1398_ /*96755*/;
assign _1396_ = _1397_ | _1399_ /*96752*/;
assign _1401_ = ~Q[62] /*96751*/;
assign _1400_ = _1401_ & D[9] /*96750*/;
assign _1403_ = _842_ & _1400_ /*96745*/;
assign _1404_ = _842_ ^ _1400_ /*96748*/;
assign _1405_ = _1396_ & _1404_ /*96746*/;
assign _1290_ = _1396_ ^ _1404_ /*96747*/;
assign _1402_ = _1403_ | _1405_ /*96744*/;
assign _1407_ = ~Q[62] /*96743*/;
assign _1406_ = _1407_ & D[10] /*96742*/;
assign _1409_ = _843_ & _1406_ /*96737*/;
assign _1410_ = _843_ ^ _1406_ /*96740*/;
assign _1411_ = _1402_ & _1410_ /*96738*/;
assign _1291_ = _1402_ ^ _1410_ /*96739*/;
assign _1408_ = _1409_ | _1411_ /*96736*/;
assign _1413_ = ~Q[62] /*96735*/;
assign _1412_ = _1413_ & D[11] /*96734*/;
assign _1415_ = _844_ & _1412_ /*96729*/;
assign _1416_ = _844_ ^ _1412_ /*96732*/;
assign _1417_ = _1408_ & _1416_ /*96730*/;
assign _1292_ = _1408_ ^ _1416_ /*96731*/;
assign _1414_ = _1415_ | _1417_ /*96728*/;
assign _1419_ = ~Q[62] /*96727*/;
assign _1418_ = _1419_ & D[12] /*96726*/;
assign _1421_ = _845_ & _1418_ /*96721*/;
assign _1422_ = _845_ ^ _1418_ /*96724*/;
assign _1423_ = _1414_ & _1422_ /*96722*/;
assign _1293_ = _1414_ ^ _1422_ /*96723*/;
assign _1420_ = _1421_ | _1423_ /*96720*/;
assign _1425_ = ~Q[62] /*96719*/;
assign _1424_ = _1425_ & D[13] /*96718*/;
assign _1427_ = _846_ & _1424_ /*96713*/;
assign _1428_ = _846_ ^ _1424_ /*96716*/;
assign _1429_ = _1420_ & _1428_ /*96714*/;
assign _1294_ = _1420_ ^ _1428_ /*96715*/;
assign _1426_ = _1427_ | _1429_ /*96712*/;
assign _1431_ = ~Q[62] /*96711*/;
assign _1430_ = _1431_ & D[14] /*96710*/;
assign _1433_ = _847_ & _1430_ /*96705*/;
assign _1434_ = _847_ ^ _1430_ /*96708*/;
assign _1435_ = _1426_ & _1434_ /*96706*/;
assign _1295_ = _1426_ ^ _1434_ /*96707*/;
assign _1432_ = _1433_ | _1435_ /*96704*/;
assign _1437_ = ~Q[62] /*96703*/;
assign _1436_ = _1437_ & D[15] /*96702*/;
assign _1439_ = _848_ & _1436_ /*96697*/;
assign _1440_ = _848_ ^ _1436_ /*96700*/;
assign _1441_ = _1432_ & _1440_ /*96698*/;
assign _1296_ = _1432_ ^ _1440_ /*96699*/;
assign _1438_ = _1439_ | _1441_ /*96696*/;
assign _1443_ = ~Q[62] /*96695*/;
assign _1442_ = _1443_ & D[16] /*96694*/;
assign _1445_ = _849_ & _1442_ /*96689*/;
assign _1446_ = _849_ ^ _1442_ /*96692*/;
assign _1447_ = _1438_ & _1446_ /*96690*/;
assign _1297_ = _1438_ ^ _1446_ /*96691*/;
assign _1444_ = _1445_ | _1447_ /*96688*/;
assign _1449_ = ~Q[62] /*96687*/;
assign _1448_ = _1449_ & D[17] /*96686*/;
assign _1451_ = _850_ & _1448_ /*96681*/;
assign _1452_ = _850_ ^ _1448_ /*96684*/;
assign _1453_ = _1444_ & _1452_ /*96682*/;
assign _1298_ = _1444_ ^ _1452_ /*96683*/;
assign _1450_ = _1451_ | _1453_ /*96680*/;
assign _1455_ = ~Q[62] /*96679*/;
assign _1454_ = _1455_ & D[18] /*96678*/;
assign _1457_ = _851_ & _1454_ /*96673*/;
assign _1458_ = _851_ ^ _1454_ /*96676*/;
assign _1459_ = _1450_ & _1458_ /*96674*/;
assign _1299_ = _1450_ ^ _1458_ /*96675*/;
assign _1456_ = _1457_ | _1459_ /*96672*/;
assign _1461_ = ~Q[62] /*96671*/;
assign _1460_ = _1461_ & D[19] /*96670*/;
assign _1463_ = _852_ & _1460_ /*96665*/;
assign _1464_ = _852_ ^ _1460_ /*96668*/;
assign _1465_ = _1456_ & _1464_ /*96666*/;
assign _1300_ = _1456_ ^ _1464_ /*96667*/;
assign _1462_ = _1463_ | _1465_ /*96664*/;
assign _1467_ = ~Q[62] /*96663*/;
assign _1466_ = _1467_ & D[20] /*96662*/;
assign _1469_ = _853_ & _1466_ /*96657*/;
assign _1470_ = _853_ ^ _1466_ /*96660*/;
assign _1471_ = _1462_ & _1470_ /*96658*/;
assign _1301_ = _1462_ ^ _1470_ /*96659*/;
assign _1468_ = _1469_ | _1471_ /*96656*/;
assign _1473_ = ~Q[62] /*96655*/;
assign _1472_ = _1473_ & D[21] /*96654*/;
assign _1475_ = _854_ & _1472_ /*96649*/;
assign _1476_ = _854_ ^ _1472_ /*96652*/;
assign _1477_ = _1468_ & _1476_ /*96650*/;
assign _1302_ = _1468_ ^ _1476_ /*96651*/;
assign _1474_ = _1475_ | _1477_ /*96648*/;
assign _1479_ = ~Q[62] /*96647*/;
assign _1478_ = _1479_ & D[22] /*96646*/;
assign _1481_ = _855_ & _1478_ /*96641*/;
assign _1482_ = _855_ ^ _1478_ /*96644*/;
assign _1483_ = _1474_ & _1482_ /*96642*/;
assign _1303_ = _1474_ ^ _1482_ /*96643*/;
assign _1480_ = _1481_ | _1483_ /*96640*/;
assign _1485_ = ~Q[62] /*96639*/;
assign _1484_ = _1485_ & D[23] /*96638*/;
assign _1487_ = _856_ & _1484_ /*96633*/;
assign _1488_ = _856_ ^ _1484_ /*96636*/;
assign _1489_ = _1480_ & _1488_ /*96634*/;
assign _1304_ = _1480_ ^ _1488_ /*96635*/;
assign _1486_ = _1487_ | _1489_ /*96632*/;
assign _1491_ = ~Q[62] /*96631*/;
assign _1490_ = _1491_ & D[24] /*96630*/;
assign _1493_ = _857_ & _1490_ /*96625*/;
assign _1494_ = _857_ ^ _1490_ /*96628*/;
assign _1495_ = _1486_ & _1494_ /*96626*/;
assign _1305_ = _1486_ ^ _1494_ /*96627*/;
assign _1492_ = _1493_ | _1495_ /*96624*/;
assign _1497_ = ~Q[62] /*96623*/;
assign _1496_ = _1497_ & D[25] /*96622*/;
assign _1499_ = _858_ & _1496_ /*96617*/;
assign _1500_ = _858_ ^ _1496_ /*96620*/;
assign _1501_ = _1492_ & _1500_ /*96618*/;
assign _1306_ = _1492_ ^ _1500_ /*96619*/;
assign _1498_ = _1499_ | _1501_ /*96616*/;
assign _1503_ = ~Q[62] /*96615*/;
assign _1502_ = _1503_ & D[26] /*96614*/;
assign _1505_ = _859_ & _1502_ /*96609*/;
assign _1506_ = _859_ ^ _1502_ /*96612*/;
assign _1507_ = _1498_ & _1506_ /*96610*/;
assign _1307_ = _1498_ ^ _1506_ /*96611*/;
assign _1504_ = _1505_ | _1507_ /*96608*/;
assign _1509_ = ~Q[62] /*96607*/;
assign _1508_ = _1509_ & D[27] /*96606*/;
assign _1511_ = _860_ & _1508_ /*96601*/;
assign _1512_ = _860_ ^ _1508_ /*96604*/;
assign _1513_ = _1504_ & _1512_ /*96602*/;
assign _1308_ = _1504_ ^ _1512_ /*96603*/;
assign _1510_ = _1511_ | _1513_ /*96600*/;
assign _1515_ = ~Q[62] /*96599*/;
assign _1514_ = _1515_ & D[28] /*96598*/;
assign _1517_ = _861_ & _1514_ /*96593*/;
assign _1518_ = _861_ ^ _1514_ /*96596*/;
assign _1519_ = _1510_ & _1518_ /*96594*/;
assign _1309_ = _1510_ ^ _1518_ /*96595*/;
assign _1516_ = _1517_ | _1519_ /*96592*/;
assign _1521_ = ~Q[62] /*96591*/;
assign _1520_ = _1521_ & D[29] /*96590*/;
assign _1523_ = _862_ & _1520_ /*96585*/;
assign _1524_ = _862_ ^ _1520_ /*96588*/;
assign _1525_ = _1516_ & _1524_ /*96586*/;
assign _1310_ = _1516_ ^ _1524_ /*96587*/;
assign _1522_ = _1523_ | _1525_ /*96584*/;
assign _1527_ = ~Q[62] /*96583*/;
assign _1526_ = _1527_ & D[30] /*96582*/;
assign _1529_ = _863_ & _1526_ /*96577*/;
assign _1530_ = _863_ ^ _1526_ /*96580*/;
assign _1531_ = _1522_ & _1530_ /*96578*/;
assign _1311_ = _1522_ ^ _1530_ /*96579*/;
assign _1528_ = _1529_ | _1531_ /*96576*/;
assign _1533_ = ~Q[62] /*96575*/;
assign _1532_ = _1533_ & D[31] /*96574*/;
assign _1535_ = _864_ & _1532_ /*96569*/;
assign _1536_ = _864_ ^ _1532_ /*96572*/;
assign _1537_ = _1528_ & _1536_ /*96570*/;
assign _1312_ = _1528_ ^ _1536_ /*96571*/;
assign _1534_ = _1535_ | _1537_ /*96568*/;
assign _1539_ = ~Q[62] /*96567*/;
assign _1538_ = _1539_ & D[32] /*96566*/;
assign _1541_ = _865_ & _1538_ /*96561*/;
assign _1542_ = _865_ ^ _1538_ /*96564*/;
assign _1543_ = _1534_ & _1542_ /*96562*/;
assign _1313_ = _1534_ ^ _1542_ /*96563*/;
assign _1540_ = _1541_ | _1543_ /*96560*/;
assign _1545_ = ~Q[62] /*96559*/;
assign _1544_ = _1545_ & D[33] /*96558*/;
assign _1547_ = _866_ & _1544_ /*96553*/;
assign _1548_ = _866_ ^ _1544_ /*96556*/;
assign _1549_ = _1540_ & _1548_ /*96554*/;
assign _1314_ = _1540_ ^ _1548_ /*96555*/;
assign _1546_ = _1547_ | _1549_ /*96552*/;
assign _1551_ = ~Q[62] /*96551*/;
assign _1550_ = _1551_ & D[34] /*96550*/;
assign _1553_ = _867_ & _1550_ /*96545*/;
assign _1554_ = _867_ ^ _1550_ /*96548*/;
assign _1555_ = _1546_ & _1554_ /*96546*/;
assign _1315_ = _1546_ ^ _1554_ /*96547*/;
assign _1552_ = _1553_ | _1555_ /*96544*/;
assign _1557_ = ~Q[62] /*96543*/;
assign _1556_ = _1557_ & D[35] /*96542*/;
assign _1559_ = _868_ & _1556_ /*96537*/;
assign _1560_ = _868_ ^ _1556_ /*96540*/;
assign _1561_ = _1552_ & _1560_ /*96538*/;
assign _1316_ = _1552_ ^ _1560_ /*96539*/;
assign _1558_ = _1559_ | _1561_ /*96536*/;
assign _1563_ = ~Q[62] /*96535*/;
assign _1562_ = _1563_ & D[36] /*96534*/;
assign _1565_ = _869_ & _1562_ /*96529*/;
assign _1566_ = _869_ ^ _1562_ /*96532*/;
assign _1567_ = _1558_ & _1566_ /*96530*/;
assign _1317_ = _1558_ ^ _1566_ /*96531*/;
assign _1564_ = _1565_ | _1567_ /*96528*/;
assign _1569_ = ~Q[62] /*96527*/;
assign _1568_ = _1569_ & D[37] /*96526*/;
assign _1571_ = _870_ & _1568_ /*96521*/;
assign _1572_ = _870_ ^ _1568_ /*96524*/;
assign _1573_ = _1564_ & _1572_ /*96522*/;
assign _1318_ = _1564_ ^ _1572_ /*96523*/;
assign _1570_ = _1571_ | _1573_ /*96520*/;
assign _1575_ = ~Q[62] /*96519*/;
assign _1574_ = _1575_ & D[38] /*96518*/;
assign _1577_ = _871_ & _1574_ /*96513*/;
assign _1578_ = _871_ ^ _1574_ /*96516*/;
assign _1579_ = _1570_ & _1578_ /*96514*/;
assign _1319_ = _1570_ ^ _1578_ /*96515*/;
assign _1576_ = _1577_ | _1579_ /*96512*/;
assign _1581_ = ~Q[62] /*96511*/;
assign _1580_ = _1581_ & D[39] /*96510*/;
assign _1583_ = _872_ & _1580_ /*96505*/;
assign _1584_ = _872_ ^ _1580_ /*96508*/;
assign _1585_ = _1576_ & _1584_ /*96506*/;
assign _1320_ = _1576_ ^ _1584_ /*96507*/;
assign _1582_ = _1583_ | _1585_ /*96504*/;
assign _1587_ = ~Q[62] /*96503*/;
assign _1586_ = _1587_ & D[40] /*96502*/;
assign _1589_ = _873_ & _1586_ /*96497*/;
assign _1590_ = _873_ ^ _1586_ /*96500*/;
assign _1591_ = _1582_ & _1590_ /*96498*/;
assign _1321_ = _1582_ ^ _1590_ /*96499*/;
assign _1588_ = _1589_ | _1591_ /*96496*/;
assign _1593_ = ~Q[62] /*96495*/;
assign _1592_ = _1593_ & D[41] /*96494*/;
assign _1595_ = _874_ & _1592_ /*96489*/;
assign _1596_ = _874_ ^ _1592_ /*96492*/;
assign _1597_ = _1588_ & _1596_ /*96490*/;
assign _1322_ = _1588_ ^ _1596_ /*96491*/;
assign _1594_ = _1595_ | _1597_ /*96488*/;
assign _1599_ = ~Q[62] /*96487*/;
assign _1598_ = _1599_ & D[42] /*96486*/;
assign _1601_ = _875_ & _1598_ /*96481*/;
assign _1602_ = _875_ ^ _1598_ /*96484*/;
assign _1603_ = _1594_ & _1602_ /*96482*/;
assign _1323_ = _1594_ ^ _1602_ /*96483*/;
assign _1600_ = _1601_ | _1603_ /*96480*/;
assign _1605_ = ~Q[62] /*96479*/;
assign _1604_ = _1605_ & D[43] /*96478*/;
assign _1607_ = _876_ & _1604_ /*96473*/;
assign _1608_ = _876_ ^ _1604_ /*96476*/;
assign _1609_ = _1600_ & _1608_ /*96474*/;
assign _1324_ = _1600_ ^ _1608_ /*96475*/;
assign _1606_ = _1607_ | _1609_ /*96472*/;
assign _1611_ = ~Q[62] /*96471*/;
assign _1610_ = _1611_ & D[44] /*96470*/;
assign _1613_ = _877_ & _1610_ /*96465*/;
assign _1614_ = _877_ ^ _1610_ /*96468*/;
assign _1615_ = _1606_ & _1614_ /*96466*/;
assign _1325_ = _1606_ ^ _1614_ /*96467*/;
assign _1612_ = _1613_ | _1615_ /*96464*/;
assign _1617_ = ~Q[62] /*96463*/;
assign _1616_ = _1617_ & D[45] /*96462*/;
assign _1619_ = _878_ & _1616_ /*96457*/;
assign _1620_ = _878_ ^ _1616_ /*96460*/;
assign _1621_ = _1612_ & _1620_ /*96458*/;
assign _1326_ = _1612_ ^ _1620_ /*96459*/;
assign _1618_ = _1619_ | _1621_ /*96456*/;
assign _1623_ = ~Q[62] /*96455*/;
assign _1622_ = _1623_ & D[46] /*96454*/;
assign _1625_ = _879_ & _1622_ /*96449*/;
assign _1626_ = _879_ ^ _1622_ /*96452*/;
assign _1627_ = _1618_ & _1626_ /*96450*/;
assign _1327_ = _1618_ ^ _1626_ /*96451*/;
assign _1624_ = _1625_ | _1627_ /*96448*/;
assign _1629_ = ~Q[62] /*96447*/;
assign _1628_ = _1629_ & D[47] /*96446*/;
assign _1631_ = _880_ & _1628_ /*96441*/;
assign _1632_ = _880_ ^ _1628_ /*96444*/;
assign _1633_ = _1624_ & _1632_ /*96442*/;
assign _1328_ = _1624_ ^ _1632_ /*96443*/;
assign _1630_ = _1631_ | _1633_ /*96440*/;
assign _1635_ = ~Q[62] /*96439*/;
assign _1634_ = _1635_ & D[48] /*96438*/;
assign _1637_ = _881_ & _1634_ /*96433*/;
assign _1638_ = _881_ ^ _1634_ /*96436*/;
assign _1639_ = _1630_ & _1638_ /*96434*/;
assign _1329_ = _1630_ ^ _1638_ /*96435*/;
assign _1636_ = _1637_ | _1639_ /*96432*/;
assign _1641_ = ~Q[62] /*96431*/;
assign _1640_ = _1641_ & D[49] /*96430*/;
assign _1643_ = _882_ & _1640_ /*96425*/;
assign _1644_ = _882_ ^ _1640_ /*96428*/;
assign _1645_ = _1636_ & _1644_ /*96426*/;
assign _1330_ = _1636_ ^ _1644_ /*96427*/;
assign _1642_ = _1643_ | _1645_ /*96424*/;
assign _1647_ = ~Q[62] /*96423*/;
assign _1646_ = _1647_ & D[50] /*96422*/;
assign _1649_ = _883_ & _1646_ /*96417*/;
assign _1650_ = _883_ ^ _1646_ /*96420*/;
assign _1651_ = _1642_ & _1650_ /*96418*/;
assign _1331_ = _1642_ ^ _1650_ /*96419*/;
assign _1648_ = _1649_ | _1651_ /*96416*/;
assign _1653_ = ~Q[62] /*96415*/;
assign _1652_ = _1653_ & D[51] /*96414*/;
assign _1655_ = _884_ & _1652_ /*96409*/;
assign _1656_ = _884_ ^ _1652_ /*96412*/;
assign _1657_ = _1648_ & _1656_ /*96410*/;
assign _1332_ = _1648_ ^ _1656_ /*96411*/;
assign _1654_ = _1655_ | _1657_ /*96408*/;
assign _1659_ = ~Q[62] /*96407*/;
assign _1658_ = _1659_ & D[52] /*96406*/;
assign _1661_ = _885_ & _1658_ /*96401*/;
assign _1662_ = _885_ ^ _1658_ /*96404*/;
assign _1663_ = _1654_ & _1662_ /*96402*/;
assign _1333_ = _1654_ ^ _1662_ /*96403*/;
assign _1660_ = _1661_ | _1663_ /*96400*/;
assign _1665_ = ~Q[62] /*96399*/;
assign _1664_ = _1665_ & D[53] /*96398*/;
assign _1667_ = _886_ & _1664_ /*96393*/;
assign _1668_ = _886_ ^ _1664_ /*96396*/;
assign _1669_ = _1660_ & _1668_ /*96394*/;
assign _1334_ = _1660_ ^ _1668_ /*96395*/;
assign _1666_ = _1667_ | _1669_ /*96392*/;
assign _1671_ = ~Q[62] /*96391*/;
assign _1670_ = _1671_ & D[54] /*96390*/;
assign _1673_ = _887_ & _1670_ /*96385*/;
assign _1674_ = _887_ ^ _1670_ /*96388*/;
assign _1675_ = _1666_ & _1674_ /*96386*/;
assign _1335_ = _1666_ ^ _1674_ /*96387*/;
assign _1672_ = _1673_ | _1675_ /*96384*/;
assign _1677_ = ~Q[62] /*96383*/;
assign _1676_ = _1677_ & D[55] /*96382*/;
assign _1679_ = _888_ & _1676_ /*96377*/;
assign _1680_ = _888_ ^ _1676_ /*96380*/;
assign _1681_ = _1672_ & _1680_ /*96378*/;
assign _1336_ = _1672_ ^ _1680_ /*96379*/;
assign _1678_ = _1679_ | _1681_ /*96376*/;
assign _1683_ = ~Q[62] /*96375*/;
assign _1682_ = _1683_ & D[56] /*96374*/;
assign _1685_ = _889_ & _1682_ /*96369*/;
assign _1686_ = _889_ ^ _1682_ /*96372*/;
assign _1687_ = _1678_ & _1686_ /*96370*/;
assign _1337_ = _1678_ ^ _1686_ /*96371*/;
assign _1684_ = _1685_ | _1687_ /*96368*/;
assign _1689_ = ~Q[62] /*96367*/;
assign _1688_ = _1689_ & D[57] /*96366*/;
assign _1691_ = _890_ & _1688_ /*96361*/;
assign _1692_ = _890_ ^ _1688_ /*96364*/;
assign _1693_ = _1684_ & _1692_ /*96362*/;
assign _1338_ = _1684_ ^ _1692_ /*96363*/;
assign _1690_ = _1691_ | _1693_ /*96360*/;
assign _1695_ = ~Q[62] /*96359*/;
assign _1694_ = _1695_ & D[58] /*96358*/;
assign _1697_ = _891_ & _1694_ /*96353*/;
assign _1698_ = _891_ ^ _1694_ /*96356*/;
assign _1699_ = _1690_ & _1698_ /*96354*/;
assign _1339_ = _1690_ ^ _1698_ /*96355*/;
assign _1696_ = _1697_ | _1699_ /*96352*/;
assign _1701_ = ~Q[62] /*96351*/;
assign _1700_ = _1701_ & D[59] /*96350*/;
assign _1703_ = _892_ & _1700_ /*96345*/;
assign _1704_ = _892_ ^ _1700_ /*96348*/;
assign _1705_ = _1696_ & _1704_ /*96346*/;
assign _1340_ = _1696_ ^ _1704_ /*96347*/;
assign _1702_ = _1703_ | _1705_ /*96344*/;
assign _1707_ = ~Q[62] /*96343*/;
assign _1706_ = _1707_ & D[60] /*96342*/;
assign _1709_ = _893_ & _1706_ /*96337*/;
assign _1710_ = _893_ ^ _1706_ /*96340*/;
assign _1711_ = _1702_ & _1710_ /*96338*/;
assign _1341_ = _1702_ ^ _1710_ /*96339*/;
assign _1708_ = _1709_ | _1711_ /*96336*/;
assign _1713_ = ~Q[62] /*96335*/;
assign _1712_ = _1713_ & D[61] /*96334*/;
assign _1715_ = _894_ & _1712_ /*96329*/;
assign _1716_ = _894_ ^ _1712_ /*96332*/;
assign _1717_ = _1708_ & _1716_ /*96330*/;
assign _1342_ = _1708_ ^ _1716_ /*96331*/;
assign _1714_ = _1715_ | _1717_ /*96328*/;
assign _1719_ = ~Q[62] /*96327*/;
assign _1718_ = _1719_ & D[62] /*96326*/;
assign _1721_ = _895_ & _1718_ /*96321*/;
assign _1722_ = _895_ ^ _1718_ /*96324*/;
assign _1723_ = _1714_ & _1722_ /*96322*/;
assign _1343_ = _1714_ ^ _1722_ /*96323*/;
assign _1720_ = _1721_ | _1723_ /*96320*/;
assign _1725_ = ~Q[62] /*96319*/;
assign _1724_ = _1725_ & zeroWire /*96318*/;
assign _1726_ = _896_ ^ _1724_ /*96316*/;
assign _1344_ = _1726_ ^ _1720_ /*96315*/;
assign _1797_ = ~D[0] /*96061*/;
assign _1794_ = R_0[61] & _1797_ /*96057*/;
assign _1795_ = R_0[61] ^ _1797_ /*96060*/;
assign _1796_ = oneWire & _1795_ /*96058*/;
assign _1729_ = oneWire ^ _1795_ /*96059*/;
assign _1793_ = _1794_ | _1796_ /*96056*/;
assign _1802_ = ~D[1] /*96055*/;
assign _1799_ = _1281_ & _1802_ /*96051*/;
assign _1800_ = _1281_ ^ _1802_ /*96054*/;
assign _1801_ = _1793_ & _1800_ /*96052*/;
assign _1730_ = _1793_ ^ _1800_ /*96053*/;
assign _1798_ = _1799_ | _1801_ /*96050*/;
assign _1807_ = ~D[2] /*96049*/;
assign _1804_ = _1282_ & _1807_ /*96045*/;
assign _1805_ = _1282_ ^ _1807_ /*96048*/;
assign _1806_ = _1798_ & _1805_ /*96046*/;
assign _1731_ = _1798_ ^ _1805_ /*96047*/;
assign _1803_ = _1804_ | _1806_ /*96044*/;
assign _1812_ = ~D[3] /*96043*/;
assign _1809_ = _1283_ & _1812_ /*96039*/;
assign _1810_ = _1283_ ^ _1812_ /*96042*/;
assign _1811_ = _1803_ & _1810_ /*96040*/;
assign _1732_ = _1803_ ^ _1810_ /*96041*/;
assign _1808_ = _1809_ | _1811_ /*96038*/;
assign _1817_ = ~D[4] /*96037*/;
assign _1814_ = _1284_ & _1817_ /*96033*/;
assign _1815_ = _1284_ ^ _1817_ /*96036*/;
assign _1816_ = _1808_ & _1815_ /*96034*/;
assign _1733_ = _1808_ ^ _1815_ /*96035*/;
assign _1813_ = _1814_ | _1816_ /*96032*/;
assign _1822_ = ~D[5] /*96031*/;
assign _1819_ = _1285_ & _1822_ /*96027*/;
assign _1820_ = _1285_ ^ _1822_ /*96030*/;
assign _1821_ = _1813_ & _1820_ /*96028*/;
assign _1734_ = _1813_ ^ _1820_ /*96029*/;
assign _1818_ = _1819_ | _1821_ /*96026*/;
assign _1827_ = ~D[6] /*96025*/;
assign _1824_ = _1286_ & _1827_ /*96021*/;
assign _1825_ = _1286_ ^ _1827_ /*96024*/;
assign _1826_ = _1818_ & _1825_ /*96022*/;
assign _1735_ = _1818_ ^ _1825_ /*96023*/;
assign _1823_ = _1824_ | _1826_ /*96020*/;
assign _1832_ = ~D[7] /*96019*/;
assign _1829_ = _1287_ & _1832_ /*96015*/;
assign _1830_ = _1287_ ^ _1832_ /*96018*/;
assign _1831_ = _1823_ & _1830_ /*96016*/;
assign _1736_ = _1823_ ^ _1830_ /*96017*/;
assign _1828_ = _1829_ | _1831_ /*96014*/;
assign _1837_ = ~D[8] /*96013*/;
assign _1834_ = _1288_ & _1837_ /*96009*/;
assign _1835_ = _1288_ ^ _1837_ /*96012*/;
assign _1836_ = _1828_ & _1835_ /*96010*/;
assign _1737_ = _1828_ ^ _1835_ /*96011*/;
assign _1833_ = _1834_ | _1836_ /*96008*/;
assign _1842_ = ~D[9] /*96007*/;
assign _1839_ = _1289_ & _1842_ /*96003*/;
assign _1840_ = _1289_ ^ _1842_ /*96006*/;
assign _1841_ = _1833_ & _1840_ /*96004*/;
assign _1738_ = _1833_ ^ _1840_ /*96005*/;
assign _1838_ = _1839_ | _1841_ /*96002*/;
assign _1847_ = ~D[10] /*96001*/;
assign _1844_ = _1290_ & _1847_ /*95997*/;
assign _1845_ = _1290_ ^ _1847_ /*96000*/;
assign _1846_ = _1838_ & _1845_ /*95998*/;
assign _1739_ = _1838_ ^ _1845_ /*95999*/;
assign _1843_ = _1844_ | _1846_ /*95996*/;
assign _1852_ = ~D[11] /*95995*/;
assign _1849_ = _1291_ & _1852_ /*95991*/;
assign _1850_ = _1291_ ^ _1852_ /*95994*/;
assign _1851_ = _1843_ & _1850_ /*95992*/;
assign _1740_ = _1843_ ^ _1850_ /*95993*/;
assign _1848_ = _1849_ | _1851_ /*95990*/;
assign _1857_ = ~D[12] /*95989*/;
assign _1854_ = _1292_ & _1857_ /*95985*/;
assign _1855_ = _1292_ ^ _1857_ /*95988*/;
assign _1856_ = _1848_ & _1855_ /*95986*/;
assign _1741_ = _1848_ ^ _1855_ /*95987*/;
assign _1853_ = _1854_ | _1856_ /*95984*/;
assign _1862_ = ~D[13] /*95983*/;
assign _1859_ = _1293_ & _1862_ /*95979*/;
assign _1860_ = _1293_ ^ _1862_ /*95982*/;
assign _1861_ = _1853_ & _1860_ /*95980*/;
assign _1742_ = _1853_ ^ _1860_ /*95981*/;
assign _1858_ = _1859_ | _1861_ /*95978*/;
assign _1867_ = ~D[14] /*95977*/;
assign _1864_ = _1294_ & _1867_ /*95973*/;
assign _1865_ = _1294_ ^ _1867_ /*95976*/;
assign _1866_ = _1858_ & _1865_ /*95974*/;
assign _1743_ = _1858_ ^ _1865_ /*95975*/;
assign _1863_ = _1864_ | _1866_ /*95972*/;
assign _1872_ = ~D[15] /*95971*/;
assign _1869_ = _1295_ & _1872_ /*95967*/;
assign _1870_ = _1295_ ^ _1872_ /*95970*/;
assign _1871_ = _1863_ & _1870_ /*95968*/;
assign _1744_ = _1863_ ^ _1870_ /*95969*/;
assign _1868_ = _1869_ | _1871_ /*95966*/;
assign _1877_ = ~D[16] /*95965*/;
assign _1874_ = _1296_ & _1877_ /*95961*/;
assign _1875_ = _1296_ ^ _1877_ /*95964*/;
assign _1876_ = _1868_ & _1875_ /*95962*/;
assign _1745_ = _1868_ ^ _1875_ /*95963*/;
assign _1873_ = _1874_ | _1876_ /*95960*/;
assign _1882_ = ~D[17] /*95959*/;
assign _1879_ = _1297_ & _1882_ /*95955*/;
assign _1880_ = _1297_ ^ _1882_ /*95958*/;
assign _1881_ = _1873_ & _1880_ /*95956*/;
assign _1746_ = _1873_ ^ _1880_ /*95957*/;
assign _1878_ = _1879_ | _1881_ /*95954*/;
assign _1887_ = ~D[18] /*95953*/;
assign _1884_ = _1298_ & _1887_ /*95949*/;
assign _1885_ = _1298_ ^ _1887_ /*95952*/;
assign _1886_ = _1878_ & _1885_ /*95950*/;
assign _1747_ = _1878_ ^ _1885_ /*95951*/;
assign _1883_ = _1884_ | _1886_ /*95948*/;
assign _1892_ = ~D[19] /*95947*/;
assign _1889_ = _1299_ & _1892_ /*95943*/;
assign _1890_ = _1299_ ^ _1892_ /*95946*/;
assign _1891_ = _1883_ & _1890_ /*95944*/;
assign _1748_ = _1883_ ^ _1890_ /*95945*/;
assign _1888_ = _1889_ | _1891_ /*95942*/;
assign _1897_ = ~D[20] /*95941*/;
assign _1894_ = _1300_ & _1897_ /*95937*/;
assign _1895_ = _1300_ ^ _1897_ /*95940*/;
assign _1896_ = _1888_ & _1895_ /*95938*/;
assign _1749_ = _1888_ ^ _1895_ /*95939*/;
assign _1893_ = _1894_ | _1896_ /*95936*/;
assign _1902_ = ~D[21] /*95935*/;
assign _1899_ = _1301_ & _1902_ /*95931*/;
assign _1900_ = _1301_ ^ _1902_ /*95934*/;
assign _1901_ = _1893_ & _1900_ /*95932*/;
assign _1750_ = _1893_ ^ _1900_ /*95933*/;
assign _1898_ = _1899_ | _1901_ /*95930*/;
assign _1907_ = ~D[22] /*95929*/;
assign _1904_ = _1302_ & _1907_ /*95925*/;
assign _1905_ = _1302_ ^ _1907_ /*95928*/;
assign _1906_ = _1898_ & _1905_ /*95926*/;
assign _1751_ = _1898_ ^ _1905_ /*95927*/;
assign _1903_ = _1904_ | _1906_ /*95924*/;
assign _1912_ = ~D[23] /*95923*/;
assign _1909_ = _1303_ & _1912_ /*95919*/;
assign _1910_ = _1303_ ^ _1912_ /*95922*/;
assign _1911_ = _1903_ & _1910_ /*95920*/;
assign _1752_ = _1903_ ^ _1910_ /*95921*/;
assign _1908_ = _1909_ | _1911_ /*95918*/;
assign _1917_ = ~D[24] /*95917*/;
assign _1914_ = _1304_ & _1917_ /*95913*/;
assign _1915_ = _1304_ ^ _1917_ /*95916*/;
assign _1916_ = _1908_ & _1915_ /*95914*/;
assign _1753_ = _1908_ ^ _1915_ /*95915*/;
assign _1913_ = _1914_ | _1916_ /*95912*/;
assign _1922_ = ~D[25] /*95911*/;
assign _1919_ = _1305_ & _1922_ /*95907*/;
assign _1920_ = _1305_ ^ _1922_ /*95910*/;
assign _1921_ = _1913_ & _1920_ /*95908*/;
assign _1754_ = _1913_ ^ _1920_ /*95909*/;
assign _1918_ = _1919_ | _1921_ /*95906*/;
assign _1927_ = ~D[26] /*95905*/;
assign _1924_ = _1306_ & _1927_ /*95901*/;
assign _1925_ = _1306_ ^ _1927_ /*95904*/;
assign _1926_ = _1918_ & _1925_ /*95902*/;
assign _1755_ = _1918_ ^ _1925_ /*95903*/;
assign _1923_ = _1924_ | _1926_ /*95900*/;
assign _1932_ = ~D[27] /*95899*/;
assign _1929_ = _1307_ & _1932_ /*95895*/;
assign _1930_ = _1307_ ^ _1932_ /*95898*/;
assign _1931_ = _1923_ & _1930_ /*95896*/;
assign _1756_ = _1923_ ^ _1930_ /*95897*/;
assign _1928_ = _1929_ | _1931_ /*95894*/;
assign _1937_ = ~D[28] /*95893*/;
assign _1934_ = _1308_ & _1937_ /*95889*/;
assign _1935_ = _1308_ ^ _1937_ /*95892*/;
assign _1936_ = _1928_ & _1935_ /*95890*/;
assign _1757_ = _1928_ ^ _1935_ /*95891*/;
assign _1933_ = _1934_ | _1936_ /*95888*/;
assign _1942_ = ~D[29] /*95887*/;
assign _1939_ = _1309_ & _1942_ /*95883*/;
assign _1940_ = _1309_ ^ _1942_ /*95886*/;
assign _1941_ = _1933_ & _1940_ /*95884*/;
assign _1758_ = _1933_ ^ _1940_ /*95885*/;
assign _1938_ = _1939_ | _1941_ /*95882*/;
assign _1947_ = ~D[30] /*95881*/;
assign _1944_ = _1310_ & _1947_ /*95877*/;
assign _1945_ = _1310_ ^ _1947_ /*95880*/;
assign _1946_ = _1938_ & _1945_ /*95878*/;
assign _1759_ = _1938_ ^ _1945_ /*95879*/;
assign _1943_ = _1944_ | _1946_ /*95876*/;
assign _1952_ = ~D[31] /*95875*/;
assign _1949_ = _1311_ & _1952_ /*95871*/;
assign _1950_ = _1311_ ^ _1952_ /*95874*/;
assign _1951_ = _1943_ & _1950_ /*95872*/;
assign _1760_ = _1943_ ^ _1950_ /*95873*/;
assign _1948_ = _1949_ | _1951_ /*95870*/;
assign _1957_ = ~D[32] /*95869*/;
assign _1954_ = _1312_ & _1957_ /*95865*/;
assign _1955_ = _1312_ ^ _1957_ /*95868*/;
assign _1956_ = _1948_ & _1955_ /*95866*/;
assign _1761_ = _1948_ ^ _1955_ /*95867*/;
assign _1953_ = _1954_ | _1956_ /*95864*/;
assign _1962_ = ~D[33] /*95863*/;
assign _1959_ = _1313_ & _1962_ /*95859*/;
assign _1960_ = _1313_ ^ _1962_ /*95862*/;
assign _1961_ = _1953_ & _1960_ /*95860*/;
assign _1762_ = _1953_ ^ _1960_ /*95861*/;
assign _1958_ = _1959_ | _1961_ /*95858*/;
assign _1967_ = ~D[34] /*95857*/;
assign _1964_ = _1314_ & _1967_ /*95853*/;
assign _1965_ = _1314_ ^ _1967_ /*95856*/;
assign _1966_ = _1958_ & _1965_ /*95854*/;
assign _1763_ = _1958_ ^ _1965_ /*95855*/;
assign _1963_ = _1964_ | _1966_ /*95852*/;
assign _1972_ = ~D[35] /*95851*/;
assign _1969_ = _1315_ & _1972_ /*95847*/;
assign _1970_ = _1315_ ^ _1972_ /*95850*/;
assign _1971_ = _1963_ & _1970_ /*95848*/;
assign _1764_ = _1963_ ^ _1970_ /*95849*/;
assign _1968_ = _1969_ | _1971_ /*95846*/;
assign _1977_ = ~D[36] /*95845*/;
assign _1974_ = _1316_ & _1977_ /*95841*/;
assign _1975_ = _1316_ ^ _1977_ /*95844*/;
assign _1976_ = _1968_ & _1975_ /*95842*/;
assign _1765_ = _1968_ ^ _1975_ /*95843*/;
assign _1973_ = _1974_ | _1976_ /*95840*/;
assign _1982_ = ~D[37] /*95839*/;
assign _1979_ = _1317_ & _1982_ /*95835*/;
assign _1980_ = _1317_ ^ _1982_ /*95838*/;
assign _1981_ = _1973_ & _1980_ /*95836*/;
assign _1766_ = _1973_ ^ _1980_ /*95837*/;
assign _1978_ = _1979_ | _1981_ /*95834*/;
assign _1987_ = ~D[38] /*95833*/;
assign _1984_ = _1318_ & _1987_ /*95829*/;
assign _1985_ = _1318_ ^ _1987_ /*95832*/;
assign _1986_ = _1978_ & _1985_ /*95830*/;
assign _1767_ = _1978_ ^ _1985_ /*95831*/;
assign _1983_ = _1984_ | _1986_ /*95828*/;
assign _1992_ = ~D[39] /*95827*/;
assign _1989_ = _1319_ & _1992_ /*95823*/;
assign _1990_ = _1319_ ^ _1992_ /*95826*/;
assign _1991_ = _1983_ & _1990_ /*95824*/;
assign _1768_ = _1983_ ^ _1990_ /*95825*/;
assign _1988_ = _1989_ | _1991_ /*95822*/;
assign _1997_ = ~D[40] /*95821*/;
assign _1994_ = _1320_ & _1997_ /*95817*/;
assign _1995_ = _1320_ ^ _1997_ /*95820*/;
assign _1996_ = _1988_ & _1995_ /*95818*/;
assign _1769_ = _1988_ ^ _1995_ /*95819*/;
assign _1993_ = _1994_ | _1996_ /*95816*/;
assign _2002_ = ~D[41] /*95815*/;
assign _1999_ = _1321_ & _2002_ /*95811*/;
assign _2000_ = _1321_ ^ _2002_ /*95814*/;
assign _2001_ = _1993_ & _2000_ /*95812*/;
assign _1770_ = _1993_ ^ _2000_ /*95813*/;
assign _1998_ = _1999_ | _2001_ /*95810*/;
assign _2007_ = ~D[42] /*95809*/;
assign _2004_ = _1322_ & _2007_ /*95805*/;
assign _2005_ = _1322_ ^ _2007_ /*95808*/;
assign _2006_ = _1998_ & _2005_ /*95806*/;
assign _1771_ = _1998_ ^ _2005_ /*95807*/;
assign _2003_ = _2004_ | _2006_ /*95804*/;
assign _2012_ = ~D[43] /*95803*/;
assign _2009_ = _1323_ & _2012_ /*95799*/;
assign _2010_ = _1323_ ^ _2012_ /*95802*/;
assign _2011_ = _2003_ & _2010_ /*95800*/;
assign _1772_ = _2003_ ^ _2010_ /*95801*/;
assign _2008_ = _2009_ | _2011_ /*95798*/;
assign _2017_ = ~D[44] /*95797*/;
assign _2014_ = _1324_ & _2017_ /*95793*/;
assign _2015_ = _1324_ ^ _2017_ /*95796*/;
assign _2016_ = _2008_ & _2015_ /*95794*/;
assign _1773_ = _2008_ ^ _2015_ /*95795*/;
assign _2013_ = _2014_ | _2016_ /*95792*/;
assign _2022_ = ~D[45] /*95791*/;
assign _2019_ = _1325_ & _2022_ /*95787*/;
assign _2020_ = _1325_ ^ _2022_ /*95790*/;
assign _2021_ = _2013_ & _2020_ /*95788*/;
assign _1774_ = _2013_ ^ _2020_ /*95789*/;
assign _2018_ = _2019_ | _2021_ /*95786*/;
assign _2027_ = ~D[46] /*95785*/;
assign _2024_ = _1326_ & _2027_ /*95781*/;
assign _2025_ = _1326_ ^ _2027_ /*95784*/;
assign _2026_ = _2018_ & _2025_ /*95782*/;
assign _1775_ = _2018_ ^ _2025_ /*95783*/;
assign _2023_ = _2024_ | _2026_ /*95780*/;
assign _2032_ = ~D[47] /*95779*/;
assign _2029_ = _1327_ & _2032_ /*95775*/;
assign _2030_ = _1327_ ^ _2032_ /*95778*/;
assign _2031_ = _2023_ & _2030_ /*95776*/;
assign _1776_ = _2023_ ^ _2030_ /*95777*/;
assign _2028_ = _2029_ | _2031_ /*95774*/;
assign _2037_ = ~D[48] /*95773*/;
assign _2034_ = _1328_ & _2037_ /*95769*/;
assign _2035_ = _1328_ ^ _2037_ /*95772*/;
assign _2036_ = _2028_ & _2035_ /*95770*/;
assign _1777_ = _2028_ ^ _2035_ /*95771*/;
assign _2033_ = _2034_ | _2036_ /*95768*/;
assign _2042_ = ~D[49] /*95767*/;
assign _2039_ = _1329_ & _2042_ /*95763*/;
assign _2040_ = _1329_ ^ _2042_ /*95766*/;
assign _2041_ = _2033_ & _2040_ /*95764*/;
assign _1778_ = _2033_ ^ _2040_ /*95765*/;
assign _2038_ = _2039_ | _2041_ /*95762*/;
assign _2047_ = ~D[50] /*95761*/;
assign _2044_ = _1330_ & _2047_ /*95757*/;
assign _2045_ = _1330_ ^ _2047_ /*95760*/;
assign _2046_ = _2038_ & _2045_ /*95758*/;
assign _1779_ = _2038_ ^ _2045_ /*95759*/;
assign _2043_ = _2044_ | _2046_ /*95756*/;
assign _2052_ = ~D[51] /*95755*/;
assign _2049_ = _1331_ & _2052_ /*95751*/;
assign _2050_ = _1331_ ^ _2052_ /*95754*/;
assign _2051_ = _2043_ & _2050_ /*95752*/;
assign _1780_ = _2043_ ^ _2050_ /*95753*/;
assign _2048_ = _2049_ | _2051_ /*95750*/;
assign _2057_ = ~D[52] /*95749*/;
assign _2054_ = _1332_ & _2057_ /*95745*/;
assign _2055_ = _1332_ ^ _2057_ /*95748*/;
assign _2056_ = _2048_ & _2055_ /*95746*/;
assign _1781_ = _2048_ ^ _2055_ /*95747*/;
assign _2053_ = _2054_ | _2056_ /*95744*/;
assign _2062_ = ~D[53] /*95743*/;
assign _2059_ = _1333_ & _2062_ /*95739*/;
assign _2060_ = _1333_ ^ _2062_ /*95742*/;
assign _2061_ = _2053_ & _2060_ /*95740*/;
assign _1782_ = _2053_ ^ _2060_ /*95741*/;
assign _2058_ = _2059_ | _2061_ /*95738*/;
assign _2067_ = ~D[54] /*95737*/;
assign _2064_ = _1334_ & _2067_ /*95733*/;
assign _2065_ = _1334_ ^ _2067_ /*95736*/;
assign _2066_ = _2058_ & _2065_ /*95734*/;
assign _1783_ = _2058_ ^ _2065_ /*95735*/;
assign _2063_ = _2064_ | _2066_ /*95732*/;
assign _2072_ = ~D[55] /*95731*/;
assign _2069_ = _1335_ & _2072_ /*95727*/;
assign _2070_ = _1335_ ^ _2072_ /*95730*/;
assign _2071_ = _2063_ & _2070_ /*95728*/;
assign _1784_ = _2063_ ^ _2070_ /*95729*/;
assign _2068_ = _2069_ | _2071_ /*95726*/;
assign _2077_ = ~D[56] /*95725*/;
assign _2074_ = _1336_ & _2077_ /*95721*/;
assign _2075_ = _1336_ ^ _2077_ /*95724*/;
assign _2076_ = _2068_ & _2075_ /*95722*/;
assign _1785_ = _2068_ ^ _2075_ /*95723*/;
assign _2073_ = _2074_ | _2076_ /*95720*/;
assign _2082_ = ~D[57] /*95719*/;
assign _2079_ = _1337_ & _2082_ /*95715*/;
assign _2080_ = _1337_ ^ _2082_ /*95718*/;
assign _2081_ = _2073_ & _2080_ /*95716*/;
assign _1786_ = _2073_ ^ _2080_ /*95717*/;
assign _2078_ = _2079_ | _2081_ /*95714*/;
assign _2087_ = ~D[58] /*95713*/;
assign _2084_ = _1338_ & _2087_ /*95709*/;
assign _2085_ = _1338_ ^ _2087_ /*95712*/;
assign _2086_ = _2078_ & _2085_ /*95710*/;
assign _1787_ = _2078_ ^ _2085_ /*95711*/;
assign _2083_ = _2084_ | _2086_ /*95708*/;
assign _2092_ = ~D[59] /*95707*/;
assign _2089_ = _1339_ & _2092_ /*95703*/;
assign _2090_ = _1339_ ^ _2092_ /*95706*/;
assign _2091_ = _2083_ & _2090_ /*95704*/;
assign _1788_ = _2083_ ^ _2090_ /*95705*/;
assign _2088_ = _2089_ | _2091_ /*95702*/;
assign _2097_ = ~D[60] /*95701*/;
assign _2094_ = _1340_ & _2097_ /*95697*/;
assign _2095_ = _1340_ ^ _2097_ /*95700*/;
assign _2096_ = _2088_ & _2095_ /*95698*/;
assign _1789_ = _2088_ ^ _2095_ /*95699*/;
assign _2093_ = _2094_ | _2096_ /*95696*/;
assign _2102_ = ~D[61] /*95695*/;
assign _2099_ = _1341_ & _2102_ /*95691*/;
assign _2100_ = _1341_ ^ _2102_ /*95694*/;
assign _2101_ = _2093_ & _2100_ /*95692*/;
assign _1790_ = _2093_ ^ _2100_ /*95693*/;
assign _2098_ = _2099_ | _2101_ /*95690*/;
assign _2107_ = ~D[62] /*95689*/;
assign _2104_ = _1342_ & _2107_ /*95685*/;
assign _2105_ = _1342_ ^ _2107_ /*95688*/;
assign _2106_ = _2098_ & _2105_ /*95686*/;
assign _1791_ = _2098_ ^ _2105_ /*95687*/;
assign _2103_ = _2104_ | _2106_ /*95684*/;
assign _2108_ = _1343_ & oneWire /*95679*/;
assign _2109_ = _1343_ ^ oneWire /*95682*/;
assign _2110_ = _2103_ & _2109_ /*95680*/;
assign _1792_ = _2103_ ^ _2109_ /*95681*/;
assign Q[61] = _2108_ | _2110_ /*95678*/;
assign _2243_ = ~Q[61] /*95293*/;
assign _2242_ = _2243_ & D[0] /*95292*/;
assign _2245_ = _1729_ & _2242_ /*95287*/;
assign _2246_ = _1729_ ^ _2242_ /*95290*/;
assign _2247_ = zeroWire & _2246_ /*95288*/;
assign _2177_ = zeroWire ^ _2246_ /*95289*/;
assign _2244_ = _2245_ | _2247_ /*95286*/;
assign _2249_ = ~Q[61] /*95285*/;
assign _2248_ = _2249_ & D[1] /*95284*/;
assign _2251_ = _1730_ & _2248_ /*95279*/;
assign _2252_ = _1730_ ^ _2248_ /*95282*/;
assign _2253_ = _2244_ & _2252_ /*95280*/;
assign _2178_ = _2244_ ^ _2252_ /*95281*/;
assign _2250_ = _2251_ | _2253_ /*95278*/;
assign _2255_ = ~Q[61] /*95277*/;
assign _2254_ = _2255_ & D[2] /*95276*/;
assign _2257_ = _1731_ & _2254_ /*95271*/;
assign _2258_ = _1731_ ^ _2254_ /*95274*/;
assign _2259_ = _2250_ & _2258_ /*95272*/;
assign _2179_ = _2250_ ^ _2258_ /*95273*/;
assign _2256_ = _2257_ | _2259_ /*95270*/;
assign _2261_ = ~Q[61] /*95269*/;
assign _2260_ = _2261_ & D[3] /*95268*/;
assign _2263_ = _1732_ & _2260_ /*95263*/;
assign _2264_ = _1732_ ^ _2260_ /*95266*/;
assign _2265_ = _2256_ & _2264_ /*95264*/;
assign _2180_ = _2256_ ^ _2264_ /*95265*/;
assign _2262_ = _2263_ | _2265_ /*95262*/;
assign _2267_ = ~Q[61] /*95261*/;
assign _2266_ = _2267_ & D[4] /*95260*/;
assign _2269_ = _1733_ & _2266_ /*95255*/;
assign _2270_ = _1733_ ^ _2266_ /*95258*/;
assign _2271_ = _2262_ & _2270_ /*95256*/;
assign _2181_ = _2262_ ^ _2270_ /*95257*/;
assign _2268_ = _2269_ | _2271_ /*95254*/;
assign _2273_ = ~Q[61] /*95253*/;
assign _2272_ = _2273_ & D[5] /*95252*/;
assign _2275_ = _1734_ & _2272_ /*95247*/;
assign _2276_ = _1734_ ^ _2272_ /*95250*/;
assign _2277_ = _2268_ & _2276_ /*95248*/;
assign _2182_ = _2268_ ^ _2276_ /*95249*/;
assign _2274_ = _2275_ | _2277_ /*95246*/;
assign _2279_ = ~Q[61] /*95245*/;
assign _2278_ = _2279_ & D[6] /*95244*/;
assign _2281_ = _1735_ & _2278_ /*95239*/;
assign _2282_ = _1735_ ^ _2278_ /*95242*/;
assign _2283_ = _2274_ & _2282_ /*95240*/;
assign _2183_ = _2274_ ^ _2282_ /*95241*/;
assign _2280_ = _2281_ | _2283_ /*95238*/;
assign _2285_ = ~Q[61] /*95237*/;
assign _2284_ = _2285_ & D[7] /*95236*/;
assign _2287_ = _1736_ & _2284_ /*95231*/;
assign _2288_ = _1736_ ^ _2284_ /*95234*/;
assign _2289_ = _2280_ & _2288_ /*95232*/;
assign _2184_ = _2280_ ^ _2288_ /*95233*/;
assign _2286_ = _2287_ | _2289_ /*95230*/;
assign _2291_ = ~Q[61] /*95229*/;
assign _2290_ = _2291_ & D[8] /*95228*/;
assign _2293_ = _1737_ & _2290_ /*95223*/;
assign _2294_ = _1737_ ^ _2290_ /*95226*/;
assign _2295_ = _2286_ & _2294_ /*95224*/;
assign _2185_ = _2286_ ^ _2294_ /*95225*/;
assign _2292_ = _2293_ | _2295_ /*95222*/;
assign _2297_ = ~Q[61] /*95221*/;
assign _2296_ = _2297_ & D[9] /*95220*/;
assign _2299_ = _1738_ & _2296_ /*95215*/;
assign _2300_ = _1738_ ^ _2296_ /*95218*/;
assign _2301_ = _2292_ & _2300_ /*95216*/;
assign _2186_ = _2292_ ^ _2300_ /*95217*/;
assign _2298_ = _2299_ | _2301_ /*95214*/;
assign _2303_ = ~Q[61] /*95213*/;
assign _2302_ = _2303_ & D[10] /*95212*/;
assign _2305_ = _1739_ & _2302_ /*95207*/;
assign _2306_ = _1739_ ^ _2302_ /*95210*/;
assign _2307_ = _2298_ & _2306_ /*95208*/;
assign _2187_ = _2298_ ^ _2306_ /*95209*/;
assign _2304_ = _2305_ | _2307_ /*95206*/;
assign _2309_ = ~Q[61] /*95205*/;
assign _2308_ = _2309_ & D[11] /*95204*/;
assign _2311_ = _1740_ & _2308_ /*95199*/;
assign _2312_ = _1740_ ^ _2308_ /*95202*/;
assign _2313_ = _2304_ & _2312_ /*95200*/;
assign _2188_ = _2304_ ^ _2312_ /*95201*/;
assign _2310_ = _2311_ | _2313_ /*95198*/;
assign _2315_ = ~Q[61] /*95197*/;
assign _2314_ = _2315_ & D[12] /*95196*/;
assign _2317_ = _1741_ & _2314_ /*95191*/;
assign _2318_ = _1741_ ^ _2314_ /*95194*/;
assign _2319_ = _2310_ & _2318_ /*95192*/;
assign _2189_ = _2310_ ^ _2318_ /*95193*/;
assign _2316_ = _2317_ | _2319_ /*95190*/;
assign _2321_ = ~Q[61] /*95189*/;
assign _2320_ = _2321_ & D[13] /*95188*/;
assign _2323_ = _1742_ & _2320_ /*95183*/;
assign _2324_ = _1742_ ^ _2320_ /*95186*/;
assign _2325_ = _2316_ & _2324_ /*95184*/;
assign _2190_ = _2316_ ^ _2324_ /*95185*/;
assign _2322_ = _2323_ | _2325_ /*95182*/;
assign _2327_ = ~Q[61] /*95181*/;
assign _2326_ = _2327_ & D[14] /*95180*/;
assign _2329_ = _1743_ & _2326_ /*95175*/;
assign _2330_ = _1743_ ^ _2326_ /*95178*/;
assign _2331_ = _2322_ & _2330_ /*95176*/;
assign _2191_ = _2322_ ^ _2330_ /*95177*/;
assign _2328_ = _2329_ | _2331_ /*95174*/;
assign _2333_ = ~Q[61] /*95173*/;
assign _2332_ = _2333_ & D[15] /*95172*/;
assign _2335_ = _1744_ & _2332_ /*95167*/;
assign _2336_ = _1744_ ^ _2332_ /*95170*/;
assign _2337_ = _2328_ & _2336_ /*95168*/;
assign _2192_ = _2328_ ^ _2336_ /*95169*/;
assign _2334_ = _2335_ | _2337_ /*95166*/;
assign _2339_ = ~Q[61] /*95165*/;
assign _2338_ = _2339_ & D[16] /*95164*/;
assign _2341_ = _1745_ & _2338_ /*95159*/;
assign _2342_ = _1745_ ^ _2338_ /*95162*/;
assign _2343_ = _2334_ & _2342_ /*95160*/;
assign _2193_ = _2334_ ^ _2342_ /*95161*/;
assign _2340_ = _2341_ | _2343_ /*95158*/;
assign _2345_ = ~Q[61] /*95157*/;
assign _2344_ = _2345_ & D[17] /*95156*/;
assign _2347_ = _1746_ & _2344_ /*95151*/;
assign _2348_ = _1746_ ^ _2344_ /*95154*/;
assign _2349_ = _2340_ & _2348_ /*95152*/;
assign _2194_ = _2340_ ^ _2348_ /*95153*/;
assign _2346_ = _2347_ | _2349_ /*95150*/;
assign _2351_ = ~Q[61] /*95149*/;
assign _2350_ = _2351_ & D[18] /*95148*/;
assign _2353_ = _1747_ & _2350_ /*95143*/;
assign _2354_ = _1747_ ^ _2350_ /*95146*/;
assign _2355_ = _2346_ & _2354_ /*95144*/;
assign _2195_ = _2346_ ^ _2354_ /*95145*/;
assign _2352_ = _2353_ | _2355_ /*95142*/;
assign _2357_ = ~Q[61] /*95141*/;
assign _2356_ = _2357_ & D[19] /*95140*/;
assign _2359_ = _1748_ & _2356_ /*95135*/;
assign _2360_ = _1748_ ^ _2356_ /*95138*/;
assign _2361_ = _2352_ & _2360_ /*95136*/;
assign _2196_ = _2352_ ^ _2360_ /*95137*/;
assign _2358_ = _2359_ | _2361_ /*95134*/;
assign _2363_ = ~Q[61] /*95133*/;
assign _2362_ = _2363_ & D[20] /*95132*/;
assign _2365_ = _1749_ & _2362_ /*95127*/;
assign _2366_ = _1749_ ^ _2362_ /*95130*/;
assign _2367_ = _2358_ & _2366_ /*95128*/;
assign _2197_ = _2358_ ^ _2366_ /*95129*/;
assign _2364_ = _2365_ | _2367_ /*95126*/;
assign _2369_ = ~Q[61] /*95125*/;
assign _2368_ = _2369_ & D[21] /*95124*/;
assign _2371_ = _1750_ & _2368_ /*95119*/;
assign _2372_ = _1750_ ^ _2368_ /*95122*/;
assign _2373_ = _2364_ & _2372_ /*95120*/;
assign _2198_ = _2364_ ^ _2372_ /*95121*/;
assign _2370_ = _2371_ | _2373_ /*95118*/;
assign _2375_ = ~Q[61] /*95117*/;
assign _2374_ = _2375_ & D[22] /*95116*/;
assign _2377_ = _1751_ & _2374_ /*95111*/;
assign _2378_ = _1751_ ^ _2374_ /*95114*/;
assign _2379_ = _2370_ & _2378_ /*95112*/;
assign _2199_ = _2370_ ^ _2378_ /*95113*/;
assign _2376_ = _2377_ | _2379_ /*95110*/;
assign _2381_ = ~Q[61] /*95109*/;
assign _2380_ = _2381_ & D[23] /*95108*/;
assign _2383_ = _1752_ & _2380_ /*95103*/;
assign _2384_ = _1752_ ^ _2380_ /*95106*/;
assign _2385_ = _2376_ & _2384_ /*95104*/;
assign _2200_ = _2376_ ^ _2384_ /*95105*/;
assign _2382_ = _2383_ | _2385_ /*95102*/;
assign _2387_ = ~Q[61] /*95101*/;
assign _2386_ = _2387_ & D[24] /*95100*/;
assign _2389_ = _1753_ & _2386_ /*95095*/;
assign _2390_ = _1753_ ^ _2386_ /*95098*/;
assign _2391_ = _2382_ & _2390_ /*95096*/;
assign _2201_ = _2382_ ^ _2390_ /*95097*/;
assign _2388_ = _2389_ | _2391_ /*95094*/;
assign _2393_ = ~Q[61] /*95093*/;
assign _2392_ = _2393_ & D[25] /*95092*/;
assign _2395_ = _1754_ & _2392_ /*95087*/;
assign _2396_ = _1754_ ^ _2392_ /*95090*/;
assign _2397_ = _2388_ & _2396_ /*95088*/;
assign _2202_ = _2388_ ^ _2396_ /*95089*/;
assign _2394_ = _2395_ | _2397_ /*95086*/;
assign _2399_ = ~Q[61] /*95085*/;
assign _2398_ = _2399_ & D[26] /*95084*/;
assign _2401_ = _1755_ & _2398_ /*95079*/;
assign _2402_ = _1755_ ^ _2398_ /*95082*/;
assign _2403_ = _2394_ & _2402_ /*95080*/;
assign _2203_ = _2394_ ^ _2402_ /*95081*/;
assign _2400_ = _2401_ | _2403_ /*95078*/;
assign _2405_ = ~Q[61] /*95077*/;
assign _2404_ = _2405_ & D[27] /*95076*/;
assign _2407_ = _1756_ & _2404_ /*95071*/;
assign _2408_ = _1756_ ^ _2404_ /*95074*/;
assign _2409_ = _2400_ & _2408_ /*95072*/;
assign _2204_ = _2400_ ^ _2408_ /*95073*/;
assign _2406_ = _2407_ | _2409_ /*95070*/;
assign _2411_ = ~Q[61] /*95069*/;
assign _2410_ = _2411_ & D[28] /*95068*/;
assign _2413_ = _1757_ & _2410_ /*95063*/;
assign _2414_ = _1757_ ^ _2410_ /*95066*/;
assign _2415_ = _2406_ & _2414_ /*95064*/;
assign _2205_ = _2406_ ^ _2414_ /*95065*/;
assign _2412_ = _2413_ | _2415_ /*95062*/;
assign _2417_ = ~Q[61] /*95061*/;
assign _2416_ = _2417_ & D[29] /*95060*/;
assign _2419_ = _1758_ & _2416_ /*95055*/;
assign _2420_ = _1758_ ^ _2416_ /*95058*/;
assign _2421_ = _2412_ & _2420_ /*95056*/;
assign _2206_ = _2412_ ^ _2420_ /*95057*/;
assign _2418_ = _2419_ | _2421_ /*95054*/;
assign _2423_ = ~Q[61] /*95053*/;
assign _2422_ = _2423_ & D[30] /*95052*/;
assign _2425_ = _1759_ & _2422_ /*95047*/;
assign _2426_ = _1759_ ^ _2422_ /*95050*/;
assign _2427_ = _2418_ & _2426_ /*95048*/;
assign _2207_ = _2418_ ^ _2426_ /*95049*/;
assign _2424_ = _2425_ | _2427_ /*95046*/;
assign _2429_ = ~Q[61] /*95045*/;
assign _2428_ = _2429_ & D[31] /*95044*/;
assign _2431_ = _1760_ & _2428_ /*95039*/;
assign _2432_ = _1760_ ^ _2428_ /*95042*/;
assign _2433_ = _2424_ & _2432_ /*95040*/;
assign _2208_ = _2424_ ^ _2432_ /*95041*/;
assign _2430_ = _2431_ | _2433_ /*95038*/;
assign _2435_ = ~Q[61] /*95037*/;
assign _2434_ = _2435_ & D[32] /*95036*/;
assign _2437_ = _1761_ & _2434_ /*95031*/;
assign _2438_ = _1761_ ^ _2434_ /*95034*/;
assign _2439_ = _2430_ & _2438_ /*95032*/;
assign _2209_ = _2430_ ^ _2438_ /*95033*/;
assign _2436_ = _2437_ | _2439_ /*95030*/;
assign _2441_ = ~Q[61] /*95029*/;
assign _2440_ = _2441_ & D[33] /*95028*/;
assign _2443_ = _1762_ & _2440_ /*95023*/;
assign _2444_ = _1762_ ^ _2440_ /*95026*/;
assign _2445_ = _2436_ & _2444_ /*95024*/;
assign _2210_ = _2436_ ^ _2444_ /*95025*/;
assign _2442_ = _2443_ | _2445_ /*95022*/;
assign _2447_ = ~Q[61] /*95021*/;
assign _2446_ = _2447_ & D[34] /*95020*/;
assign _2449_ = _1763_ & _2446_ /*95015*/;
assign _2450_ = _1763_ ^ _2446_ /*95018*/;
assign _2451_ = _2442_ & _2450_ /*95016*/;
assign _2211_ = _2442_ ^ _2450_ /*95017*/;
assign _2448_ = _2449_ | _2451_ /*95014*/;
assign _2453_ = ~Q[61] /*95013*/;
assign _2452_ = _2453_ & D[35] /*95012*/;
assign _2455_ = _1764_ & _2452_ /*95007*/;
assign _2456_ = _1764_ ^ _2452_ /*95010*/;
assign _2457_ = _2448_ & _2456_ /*95008*/;
assign _2212_ = _2448_ ^ _2456_ /*95009*/;
assign _2454_ = _2455_ | _2457_ /*95006*/;
assign _2459_ = ~Q[61] /*95005*/;
assign _2458_ = _2459_ & D[36] /*95004*/;
assign _2461_ = _1765_ & _2458_ /*94999*/;
assign _2462_ = _1765_ ^ _2458_ /*95002*/;
assign _2463_ = _2454_ & _2462_ /*95000*/;
assign _2213_ = _2454_ ^ _2462_ /*95001*/;
assign _2460_ = _2461_ | _2463_ /*94998*/;
assign _2465_ = ~Q[61] /*94997*/;
assign _2464_ = _2465_ & D[37] /*94996*/;
assign _2467_ = _1766_ & _2464_ /*94991*/;
assign _2468_ = _1766_ ^ _2464_ /*94994*/;
assign _2469_ = _2460_ & _2468_ /*94992*/;
assign _2214_ = _2460_ ^ _2468_ /*94993*/;
assign _2466_ = _2467_ | _2469_ /*94990*/;
assign _2471_ = ~Q[61] /*94989*/;
assign _2470_ = _2471_ & D[38] /*94988*/;
assign _2473_ = _1767_ & _2470_ /*94983*/;
assign _2474_ = _1767_ ^ _2470_ /*94986*/;
assign _2475_ = _2466_ & _2474_ /*94984*/;
assign _2215_ = _2466_ ^ _2474_ /*94985*/;
assign _2472_ = _2473_ | _2475_ /*94982*/;
assign _2477_ = ~Q[61] /*94981*/;
assign _2476_ = _2477_ & D[39] /*94980*/;
assign _2479_ = _1768_ & _2476_ /*94975*/;
assign _2480_ = _1768_ ^ _2476_ /*94978*/;
assign _2481_ = _2472_ & _2480_ /*94976*/;
assign _2216_ = _2472_ ^ _2480_ /*94977*/;
assign _2478_ = _2479_ | _2481_ /*94974*/;
assign _2483_ = ~Q[61] /*94973*/;
assign _2482_ = _2483_ & D[40] /*94972*/;
assign _2485_ = _1769_ & _2482_ /*94967*/;
assign _2486_ = _1769_ ^ _2482_ /*94970*/;
assign _2487_ = _2478_ & _2486_ /*94968*/;
assign _2217_ = _2478_ ^ _2486_ /*94969*/;
assign _2484_ = _2485_ | _2487_ /*94966*/;
assign _2489_ = ~Q[61] /*94965*/;
assign _2488_ = _2489_ & D[41] /*94964*/;
assign _2491_ = _1770_ & _2488_ /*94959*/;
assign _2492_ = _1770_ ^ _2488_ /*94962*/;
assign _2493_ = _2484_ & _2492_ /*94960*/;
assign _2218_ = _2484_ ^ _2492_ /*94961*/;
assign _2490_ = _2491_ | _2493_ /*94958*/;
assign _2495_ = ~Q[61] /*94957*/;
assign _2494_ = _2495_ & D[42] /*94956*/;
assign _2497_ = _1771_ & _2494_ /*94951*/;
assign _2498_ = _1771_ ^ _2494_ /*94954*/;
assign _2499_ = _2490_ & _2498_ /*94952*/;
assign _2219_ = _2490_ ^ _2498_ /*94953*/;
assign _2496_ = _2497_ | _2499_ /*94950*/;
assign _2501_ = ~Q[61] /*94949*/;
assign _2500_ = _2501_ & D[43] /*94948*/;
assign _2503_ = _1772_ & _2500_ /*94943*/;
assign _2504_ = _1772_ ^ _2500_ /*94946*/;
assign _2505_ = _2496_ & _2504_ /*94944*/;
assign _2220_ = _2496_ ^ _2504_ /*94945*/;
assign _2502_ = _2503_ | _2505_ /*94942*/;
assign _2507_ = ~Q[61] /*94941*/;
assign _2506_ = _2507_ & D[44] /*94940*/;
assign _2509_ = _1773_ & _2506_ /*94935*/;
assign _2510_ = _1773_ ^ _2506_ /*94938*/;
assign _2511_ = _2502_ & _2510_ /*94936*/;
assign _2221_ = _2502_ ^ _2510_ /*94937*/;
assign _2508_ = _2509_ | _2511_ /*94934*/;
assign _2513_ = ~Q[61] /*94933*/;
assign _2512_ = _2513_ & D[45] /*94932*/;
assign _2515_ = _1774_ & _2512_ /*94927*/;
assign _2516_ = _1774_ ^ _2512_ /*94930*/;
assign _2517_ = _2508_ & _2516_ /*94928*/;
assign _2222_ = _2508_ ^ _2516_ /*94929*/;
assign _2514_ = _2515_ | _2517_ /*94926*/;
assign _2519_ = ~Q[61] /*94925*/;
assign _2518_ = _2519_ & D[46] /*94924*/;
assign _2521_ = _1775_ & _2518_ /*94919*/;
assign _2522_ = _1775_ ^ _2518_ /*94922*/;
assign _2523_ = _2514_ & _2522_ /*94920*/;
assign _2223_ = _2514_ ^ _2522_ /*94921*/;
assign _2520_ = _2521_ | _2523_ /*94918*/;
assign _2525_ = ~Q[61] /*94917*/;
assign _2524_ = _2525_ & D[47] /*94916*/;
assign _2527_ = _1776_ & _2524_ /*94911*/;
assign _2528_ = _1776_ ^ _2524_ /*94914*/;
assign _2529_ = _2520_ & _2528_ /*94912*/;
assign _2224_ = _2520_ ^ _2528_ /*94913*/;
assign _2526_ = _2527_ | _2529_ /*94910*/;
assign _2531_ = ~Q[61] /*94909*/;
assign _2530_ = _2531_ & D[48] /*94908*/;
assign _2533_ = _1777_ & _2530_ /*94903*/;
assign _2534_ = _1777_ ^ _2530_ /*94906*/;
assign _2535_ = _2526_ & _2534_ /*94904*/;
assign _2225_ = _2526_ ^ _2534_ /*94905*/;
assign _2532_ = _2533_ | _2535_ /*94902*/;
assign _2537_ = ~Q[61] /*94901*/;
assign _2536_ = _2537_ & D[49] /*94900*/;
assign _2539_ = _1778_ & _2536_ /*94895*/;
assign _2540_ = _1778_ ^ _2536_ /*94898*/;
assign _2541_ = _2532_ & _2540_ /*94896*/;
assign _2226_ = _2532_ ^ _2540_ /*94897*/;
assign _2538_ = _2539_ | _2541_ /*94894*/;
assign _2543_ = ~Q[61] /*94893*/;
assign _2542_ = _2543_ & D[50] /*94892*/;
assign _2545_ = _1779_ & _2542_ /*94887*/;
assign _2546_ = _1779_ ^ _2542_ /*94890*/;
assign _2547_ = _2538_ & _2546_ /*94888*/;
assign _2227_ = _2538_ ^ _2546_ /*94889*/;
assign _2544_ = _2545_ | _2547_ /*94886*/;
assign _2549_ = ~Q[61] /*94885*/;
assign _2548_ = _2549_ & D[51] /*94884*/;
assign _2551_ = _1780_ & _2548_ /*94879*/;
assign _2552_ = _1780_ ^ _2548_ /*94882*/;
assign _2553_ = _2544_ & _2552_ /*94880*/;
assign _2228_ = _2544_ ^ _2552_ /*94881*/;
assign _2550_ = _2551_ | _2553_ /*94878*/;
assign _2555_ = ~Q[61] /*94877*/;
assign _2554_ = _2555_ & D[52] /*94876*/;
assign _2557_ = _1781_ & _2554_ /*94871*/;
assign _2558_ = _1781_ ^ _2554_ /*94874*/;
assign _2559_ = _2550_ & _2558_ /*94872*/;
assign _2229_ = _2550_ ^ _2558_ /*94873*/;
assign _2556_ = _2557_ | _2559_ /*94870*/;
assign _2561_ = ~Q[61] /*94869*/;
assign _2560_ = _2561_ & D[53] /*94868*/;
assign _2563_ = _1782_ & _2560_ /*94863*/;
assign _2564_ = _1782_ ^ _2560_ /*94866*/;
assign _2565_ = _2556_ & _2564_ /*94864*/;
assign _2230_ = _2556_ ^ _2564_ /*94865*/;
assign _2562_ = _2563_ | _2565_ /*94862*/;
assign _2567_ = ~Q[61] /*94861*/;
assign _2566_ = _2567_ & D[54] /*94860*/;
assign _2569_ = _1783_ & _2566_ /*94855*/;
assign _2570_ = _1783_ ^ _2566_ /*94858*/;
assign _2571_ = _2562_ & _2570_ /*94856*/;
assign _2231_ = _2562_ ^ _2570_ /*94857*/;
assign _2568_ = _2569_ | _2571_ /*94854*/;
assign _2573_ = ~Q[61] /*94853*/;
assign _2572_ = _2573_ & D[55] /*94852*/;
assign _2575_ = _1784_ & _2572_ /*94847*/;
assign _2576_ = _1784_ ^ _2572_ /*94850*/;
assign _2577_ = _2568_ & _2576_ /*94848*/;
assign _2232_ = _2568_ ^ _2576_ /*94849*/;
assign _2574_ = _2575_ | _2577_ /*94846*/;
assign _2579_ = ~Q[61] /*94845*/;
assign _2578_ = _2579_ & D[56] /*94844*/;
assign _2581_ = _1785_ & _2578_ /*94839*/;
assign _2582_ = _1785_ ^ _2578_ /*94842*/;
assign _2583_ = _2574_ & _2582_ /*94840*/;
assign _2233_ = _2574_ ^ _2582_ /*94841*/;
assign _2580_ = _2581_ | _2583_ /*94838*/;
assign _2585_ = ~Q[61] /*94837*/;
assign _2584_ = _2585_ & D[57] /*94836*/;
assign _2587_ = _1786_ & _2584_ /*94831*/;
assign _2588_ = _1786_ ^ _2584_ /*94834*/;
assign _2589_ = _2580_ & _2588_ /*94832*/;
assign _2234_ = _2580_ ^ _2588_ /*94833*/;
assign _2586_ = _2587_ | _2589_ /*94830*/;
assign _2591_ = ~Q[61] /*94829*/;
assign _2590_ = _2591_ & D[58] /*94828*/;
assign _2593_ = _1787_ & _2590_ /*94823*/;
assign _2594_ = _1787_ ^ _2590_ /*94826*/;
assign _2595_ = _2586_ & _2594_ /*94824*/;
assign _2235_ = _2586_ ^ _2594_ /*94825*/;
assign _2592_ = _2593_ | _2595_ /*94822*/;
assign _2597_ = ~Q[61] /*94821*/;
assign _2596_ = _2597_ & D[59] /*94820*/;
assign _2599_ = _1788_ & _2596_ /*94815*/;
assign _2600_ = _1788_ ^ _2596_ /*94818*/;
assign _2601_ = _2592_ & _2600_ /*94816*/;
assign _2236_ = _2592_ ^ _2600_ /*94817*/;
assign _2598_ = _2599_ | _2601_ /*94814*/;
assign _2603_ = ~Q[61] /*94813*/;
assign _2602_ = _2603_ & D[60] /*94812*/;
assign _2605_ = _1789_ & _2602_ /*94807*/;
assign _2606_ = _1789_ ^ _2602_ /*94810*/;
assign _2607_ = _2598_ & _2606_ /*94808*/;
assign _2237_ = _2598_ ^ _2606_ /*94809*/;
assign _2604_ = _2605_ | _2607_ /*94806*/;
assign _2609_ = ~Q[61] /*94805*/;
assign _2608_ = _2609_ & D[61] /*94804*/;
assign _2611_ = _1790_ & _2608_ /*94799*/;
assign _2612_ = _1790_ ^ _2608_ /*94802*/;
assign _2613_ = _2604_ & _2612_ /*94800*/;
assign _2238_ = _2604_ ^ _2612_ /*94801*/;
assign _2610_ = _2611_ | _2613_ /*94798*/;
assign _2615_ = ~Q[61] /*94797*/;
assign _2614_ = _2615_ & D[62] /*94796*/;
assign _2617_ = _1791_ & _2614_ /*94791*/;
assign _2618_ = _1791_ ^ _2614_ /*94794*/;
assign _2619_ = _2610_ & _2618_ /*94792*/;
assign _2239_ = _2610_ ^ _2618_ /*94793*/;
assign _2616_ = _2617_ | _2619_ /*94790*/;
assign _2621_ = ~Q[61] /*94789*/;
assign _2620_ = _2621_ & zeroWire /*94788*/;
assign _2622_ = _1792_ ^ _2620_ /*94786*/;
assign _2240_ = _2622_ ^ _2616_ /*94785*/;
assign _2693_ = ~D[0] /*94531*/;
assign _2690_ = R_0[60] & _2693_ /*94527*/;
assign _2691_ = R_0[60] ^ _2693_ /*94530*/;
assign _2692_ = oneWire & _2691_ /*94528*/;
assign _2625_ = oneWire ^ _2691_ /*94529*/;
assign _2689_ = _2690_ | _2692_ /*94526*/;
assign _2698_ = ~D[1] /*94525*/;
assign _2695_ = _2177_ & _2698_ /*94521*/;
assign _2696_ = _2177_ ^ _2698_ /*94524*/;
assign _2697_ = _2689_ & _2696_ /*94522*/;
assign _2626_ = _2689_ ^ _2696_ /*94523*/;
assign _2694_ = _2695_ | _2697_ /*94520*/;
assign _2703_ = ~D[2] /*94519*/;
assign _2700_ = _2178_ & _2703_ /*94515*/;
assign _2701_ = _2178_ ^ _2703_ /*94518*/;
assign _2702_ = _2694_ & _2701_ /*94516*/;
assign _2627_ = _2694_ ^ _2701_ /*94517*/;
assign _2699_ = _2700_ | _2702_ /*94514*/;
assign _2708_ = ~D[3] /*94513*/;
assign _2705_ = _2179_ & _2708_ /*94509*/;
assign _2706_ = _2179_ ^ _2708_ /*94512*/;
assign _2707_ = _2699_ & _2706_ /*94510*/;
assign _2628_ = _2699_ ^ _2706_ /*94511*/;
assign _2704_ = _2705_ | _2707_ /*94508*/;
assign _2713_ = ~D[4] /*94507*/;
assign _2710_ = _2180_ & _2713_ /*94503*/;
assign _2711_ = _2180_ ^ _2713_ /*94506*/;
assign _2712_ = _2704_ & _2711_ /*94504*/;
assign _2629_ = _2704_ ^ _2711_ /*94505*/;
assign _2709_ = _2710_ | _2712_ /*94502*/;
assign _2718_ = ~D[5] /*94501*/;
assign _2715_ = _2181_ & _2718_ /*94497*/;
assign _2716_ = _2181_ ^ _2718_ /*94500*/;
assign _2717_ = _2709_ & _2716_ /*94498*/;
assign _2630_ = _2709_ ^ _2716_ /*94499*/;
assign _2714_ = _2715_ | _2717_ /*94496*/;
assign _2723_ = ~D[6] /*94495*/;
assign _2720_ = _2182_ & _2723_ /*94491*/;
assign _2721_ = _2182_ ^ _2723_ /*94494*/;
assign _2722_ = _2714_ & _2721_ /*94492*/;
assign _2631_ = _2714_ ^ _2721_ /*94493*/;
assign _2719_ = _2720_ | _2722_ /*94490*/;
assign _2728_ = ~D[7] /*94489*/;
assign _2725_ = _2183_ & _2728_ /*94485*/;
assign _2726_ = _2183_ ^ _2728_ /*94488*/;
assign _2727_ = _2719_ & _2726_ /*94486*/;
assign _2632_ = _2719_ ^ _2726_ /*94487*/;
assign _2724_ = _2725_ | _2727_ /*94484*/;
assign _2733_ = ~D[8] /*94483*/;
assign _2730_ = _2184_ & _2733_ /*94479*/;
assign _2731_ = _2184_ ^ _2733_ /*94482*/;
assign _2732_ = _2724_ & _2731_ /*94480*/;
assign _2633_ = _2724_ ^ _2731_ /*94481*/;
assign _2729_ = _2730_ | _2732_ /*94478*/;
assign _2738_ = ~D[9] /*94477*/;
assign _2735_ = _2185_ & _2738_ /*94473*/;
assign _2736_ = _2185_ ^ _2738_ /*94476*/;
assign _2737_ = _2729_ & _2736_ /*94474*/;
assign _2634_ = _2729_ ^ _2736_ /*94475*/;
assign _2734_ = _2735_ | _2737_ /*94472*/;
assign _2743_ = ~D[10] /*94471*/;
assign _2740_ = _2186_ & _2743_ /*94467*/;
assign _2741_ = _2186_ ^ _2743_ /*94470*/;
assign _2742_ = _2734_ & _2741_ /*94468*/;
assign _2635_ = _2734_ ^ _2741_ /*94469*/;
assign _2739_ = _2740_ | _2742_ /*94466*/;
assign _2748_ = ~D[11] /*94465*/;
assign _2745_ = _2187_ & _2748_ /*94461*/;
assign _2746_ = _2187_ ^ _2748_ /*94464*/;
assign _2747_ = _2739_ & _2746_ /*94462*/;
assign _2636_ = _2739_ ^ _2746_ /*94463*/;
assign _2744_ = _2745_ | _2747_ /*94460*/;
assign _2753_ = ~D[12] /*94459*/;
assign _2750_ = _2188_ & _2753_ /*94455*/;
assign _2751_ = _2188_ ^ _2753_ /*94458*/;
assign _2752_ = _2744_ & _2751_ /*94456*/;
assign _2637_ = _2744_ ^ _2751_ /*94457*/;
assign _2749_ = _2750_ | _2752_ /*94454*/;
assign _2758_ = ~D[13] /*94453*/;
assign _2755_ = _2189_ & _2758_ /*94449*/;
assign _2756_ = _2189_ ^ _2758_ /*94452*/;
assign _2757_ = _2749_ & _2756_ /*94450*/;
assign _2638_ = _2749_ ^ _2756_ /*94451*/;
assign _2754_ = _2755_ | _2757_ /*94448*/;
assign _2763_ = ~D[14] /*94447*/;
assign _2760_ = _2190_ & _2763_ /*94443*/;
assign _2761_ = _2190_ ^ _2763_ /*94446*/;
assign _2762_ = _2754_ & _2761_ /*94444*/;
assign _2639_ = _2754_ ^ _2761_ /*94445*/;
assign _2759_ = _2760_ | _2762_ /*94442*/;
assign _2768_ = ~D[15] /*94441*/;
assign _2765_ = _2191_ & _2768_ /*94437*/;
assign _2766_ = _2191_ ^ _2768_ /*94440*/;
assign _2767_ = _2759_ & _2766_ /*94438*/;
assign _2640_ = _2759_ ^ _2766_ /*94439*/;
assign _2764_ = _2765_ | _2767_ /*94436*/;
assign _2773_ = ~D[16] /*94435*/;
assign _2770_ = _2192_ & _2773_ /*94431*/;
assign _2771_ = _2192_ ^ _2773_ /*94434*/;
assign _2772_ = _2764_ & _2771_ /*94432*/;
assign _2641_ = _2764_ ^ _2771_ /*94433*/;
assign _2769_ = _2770_ | _2772_ /*94430*/;
assign _2778_ = ~D[17] /*94429*/;
assign _2775_ = _2193_ & _2778_ /*94425*/;
assign _2776_ = _2193_ ^ _2778_ /*94428*/;
assign _2777_ = _2769_ & _2776_ /*94426*/;
assign _2642_ = _2769_ ^ _2776_ /*94427*/;
assign _2774_ = _2775_ | _2777_ /*94424*/;
assign _2783_ = ~D[18] /*94423*/;
assign _2780_ = _2194_ & _2783_ /*94419*/;
assign _2781_ = _2194_ ^ _2783_ /*94422*/;
assign _2782_ = _2774_ & _2781_ /*94420*/;
assign _2643_ = _2774_ ^ _2781_ /*94421*/;
assign _2779_ = _2780_ | _2782_ /*94418*/;
assign _2788_ = ~D[19] /*94417*/;
assign _2785_ = _2195_ & _2788_ /*94413*/;
assign _2786_ = _2195_ ^ _2788_ /*94416*/;
assign _2787_ = _2779_ & _2786_ /*94414*/;
assign _2644_ = _2779_ ^ _2786_ /*94415*/;
assign _2784_ = _2785_ | _2787_ /*94412*/;
assign _2793_ = ~D[20] /*94411*/;
assign _2790_ = _2196_ & _2793_ /*94407*/;
assign _2791_ = _2196_ ^ _2793_ /*94410*/;
assign _2792_ = _2784_ & _2791_ /*94408*/;
assign _2645_ = _2784_ ^ _2791_ /*94409*/;
assign _2789_ = _2790_ | _2792_ /*94406*/;
assign _2798_ = ~D[21] /*94405*/;
assign _2795_ = _2197_ & _2798_ /*94401*/;
assign _2796_ = _2197_ ^ _2798_ /*94404*/;
assign _2797_ = _2789_ & _2796_ /*94402*/;
assign _2646_ = _2789_ ^ _2796_ /*94403*/;
assign _2794_ = _2795_ | _2797_ /*94400*/;
assign _2803_ = ~D[22] /*94399*/;
assign _2800_ = _2198_ & _2803_ /*94395*/;
assign _2801_ = _2198_ ^ _2803_ /*94398*/;
assign _2802_ = _2794_ & _2801_ /*94396*/;
assign _2647_ = _2794_ ^ _2801_ /*94397*/;
assign _2799_ = _2800_ | _2802_ /*94394*/;
assign _2808_ = ~D[23] /*94393*/;
assign _2805_ = _2199_ & _2808_ /*94389*/;
assign _2806_ = _2199_ ^ _2808_ /*94392*/;
assign _2807_ = _2799_ & _2806_ /*94390*/;
assign _2648_ = _2799_ ^ _2806_ /*94391*/;
assign _2804_ = _2805_ | _2807_ /*94388*/;
assign _2813_ = ~D[24] /*94387*/;
assign _2810_ = _2200_ & _2813_ /*94383*/;
assign _2811_ = _2200_ ^ _2813_ /*94386*/;
assign _2812_ = _2804_ & _2811_ /*94384*/;
assign _2649_ = _2804_ ^ _2811_ /*94385*/;
assign _2809_ = _2810_ | _2812_ /*94382*/;
assign _2818_ = ~D[25] /*94381*/;
assign _2815_ = _2201_ & _2818_ /*94377*/;
assign _2816_ = _2201_ ^ _2818_ /*94380*/;
assign _2817_ = _2809_ & _2816_ /*94378*/;
assign _2650_ = _2809_ ^ _2816_ /*94379*/;
assign _2814_ = _2815_ | _2817_ /*94376*/;
assign _2823_ = ~D[26] /*94375*/;
assign _2820_ = _2202_ & _2823_ /*94371*/;
assign _2821_ = _2202_ ^ _2823_ /*94374*/;
assign _2822_ = _2814_ & _2821_ /*94372*/;
assign _2651_ = _2814_ ^ _2821_ /*94373*/;
assign _2819_ = _2820_ | _2822_ /*94370*/;
assign _2828_ = ~D[27] /*94369*/;
assign _2825_ = _2203_ & _2828_ /*94365*/;
assign _2826_ = _2203_ ^ _2828_ /*94368*/;
assign _2827_ = _2819_ & _2826_ /*94366*/;
assign _2652_ = _2819_ ^ _2826_ /*94367*/;
assign _2824_ = _2825_ | _2827_ /*94364*/;
assign _2833_ = ~D[28] /*94363*/;
assign _2830_ = _2204_ & _2833_ /*94359*/;
assign _2831_ = _2204_ ^ _2833_ /*94362*/;
assign _2832_ = _2824_ & _2831_ /*94360*/;
assign _2653_ = _2824_ ^ _2831_ /*94361*/;
assign _2829_ = _2830_ | _2832_ /*94358*/;
assign _2838_ = ~D[29] /*94357*/;
assign _2835_ = _2205_ & _2838_ /*94353*/;
assign _2836_ = _2205_ ^ _2838_ /*94356*/;
assign _2837_ = _2829_ & _2836_ /*94354*/;
assign _2654_ = _2829_ ^ _2836_ /*94355*/;
assign _2834_ = _2835_ | _2837_ /*94352*/;
assign _2843_ = ~D[30] /*94351*/;
assign _2840_ = _2206_ & _2843_ /*94347*/;
assign _2841_ = _2206_ ^ _2843_ /*94350*/;
assign _2842_ = _2834_ & _2841_ /*94348*/;
assign _2655_ = _2834_ ^ _2841_ /*94349*/;
assign _2839_ = _2840_ | _2842_ /*94346*/;
assign _2848_ = ~D[31] /*94345*/;
assign _2845_ = _2207_ & _2848_ /*94341*/;
assign _2846_ = _2207_ ^ _2848_ /*94344*/;
assign _2847_ = _2839_ & _2846_ /*94342*/;
assign _2656_ = _2839_ ^ _2846_ /*94343*/;
assign _2844_ = _2845_ | _2847_ /*94340*/;
assign _2853_ = ~D[32] /*94339*/;
assign _2850_ = _2208_ & _2853_ /*94335*/;
assign _2851_ = _2208_ ^ _2853_ /*94338*/;
assign _2852_ = _2844_ & _2851_ /*94336*/;
assign _2657_ = _2844_ ^ _2851_ /*94337*/;
assign _2849_ = _2850_ | _2852_ /*94334*/;
assign _2858_ = ~D[33] /*94333*/;
assign _2855_ = _2209_ & _2858_ /*94329*/;
assign _2856_ = _2209_ ^ _2858_ /*94332*/;
assign _2857_ = _2849_ & _2856_ /*94330*/;
assign _2658_ = _2849_ ^ _2856_ /*94331*/;
assign _2854_ = _2855_ | _2857_ /*94328*/;
assign _2863_ = ~D[34] /*94327*/;
assign _2860_ = _2210_ & _2863_ /*94323*/;
assign _2861_ = _2210_ ^ _2863_ /*94326*/;
assign _2862_ = _2854_ & _2861_ /*94324*/;
assign _2659_ = _2854_ ^ _2861_ /*94325*/;
assign _2859_ = _2860_ | _2862_ /*94322*/;
assign _2868_ = ~D[35] /*94321*/;
assign _2865_ = _2211_ & _2868_ /*94317*/;
assign _2866_ = _2211_ ^ _2868_ /*94320*/;
assign _2867_ = _2859_ & _2866_ /*94318*/;
assign _2660_ = _2859_ ^ _2866_ /*94319*/;
assign _2864_ = _2865_ | _2867_ /*94316*/;
assign _2873_ = ~D[36] /*94315*/;
assign _2870_ = _2212_ & _2873_ /*94311*/;
assign _2871_ = _2212_ ^ _2873_ /*94314*/;
assign _2872_ = _2864_ & _2871_ /*94312*/;
assign _2661_ = _2864_ ^ _2871_ /*94313*/;
assign _2869_ = _2870_ | _2872_ /*94310*/;
assign _2878_ = ~D[37] /*94309*/;
assign _2875_ = _2213_ & _2878_ /*94305*/;
assign _2876_ = _2213_ ^ _2878_ /*94308*/;
assign _2877_ = _2869_ & _2876_ /*94306*/;
assign _2662_ = _2869_ ^ _2876_ /*94307*/;
assign _2874_ = _2875_ | _2877_ /*94304*/;
assign _2883_ = ~D[38] /*94303*/;
assign _2880_ = _2214_ & _2883_ /*94299*/;
assign _2881_ = _2214_ ^ _2883_ /*94302*/;
assign _2882_ = _2874_ & _2881_ /*94300*/;
assign _2663_ = _2874_ ^ _2881_ /*94301*/;
assign _2879_ = _2880_ | _2882_ /*94298*/;
assign _2888_ = ~D[39] /*94297*/;
assign _2885_ = _2215_ & _2888_ /*94293*/;
assign _2886_ = _2215_ ^ _2888_ /*94296*/;
assign _2887_ = _2879_ & _2886_ /*94294*/;
assign _2664_ = _2879_ ^ _2886_ /*94295*/;
assign _2884_ = _2885_ | _2887_ /*94292*/;
assign _2893_ = ~D[40] /*94291*/;
assign _2890_ = _2216_ & _2893_ /*94287*/;
assign _2891_ = _2216_ ^ _2893_ /*94290*/;
assign _2892_ = _2884_ & _2891_ /*94288*/;
assign _2665_ = _2884_ ^ _2891_ /*94289*/;
assign _2889_ = _2890_ | _2892_ /*94286*/;
assign _2898_ = ~D[41] /*94285*/;
assign _2895_ = _2217_ & _2898_ /*94281*/;
assign _2896_ = _2217_ ^ _2898_ /*94284*/;
assign _2897_ = _2889_ & _2896_ /*94282*/;
assign _2666_ = _2889_ ^ _2896_ /*94283*/;
assign _2894_ = _2895_ | _2897_ /*94280*/;
assign _2903_ = ~D[42] /*94279*/;
assign _2900_ = _2218_ & _2903_ /*94275*/;
assign _2901_ = _2218_ ^ _2903_ /*94278*/;
assign _2902_ = _2894_ & _2901_ /*94276*/;
assign _2667_ = _2894_ ^ _2901_ /*94277*/;
assign _2899_ = _2900_ | _2902_ /*94274*/;
assign _2908_ = ~D[43] /*94273*/;
assign _2905_ = _2219_ & _2908_ /*94269*/;
assign _2906_ = _2219_ ^ _2908_ /*94272*/;
assign _2907_ = _2899_ & _2906_ /*94270*/;
assign _2668_ = _2899_ ^ _2906_ /*94271*/;
assign _2904_ = _2905_ | _2907_ /*94268*/;
assign _2913_ = ~D[44] /*94267*/;
assign _2910_ = _2220_ & _2913_ /*94263*/;
assign _2911_ = _2220_ ^ _2913_ /*94266*/;
assign _2912_ = _2904_ & _2911_ /*94264*/;
assign _2669_ = _2904_ ^ _2911_ /*94265*/;
assign _2909_ = _2910_ | _2912_ /*94262*/;
assign _2918_ = ~D[45] /*94261*/;
assign _2915_ = _2221_ & _2918_ /*94257*/;
assign _2916_ = _2221_ ^ _2918_ /*94260*/;
assign _2917_ = _2909_ & _2916_ /*94258*/;
assign _2670_ = _2909_ ^ _2916_ /*94259*/;
assign _2914_ = _2915_ | _2917_ /*94256*/;
assign _2923_ = ~D[46] /*94255*/;
assign _2920_ = _2222_ & _2923_ /*94251*/;
assign _2921_ = _2222_ ^ _2923_ /*94254*/;
assign _2922_ = _2914_ & _2921_ /*94252*/;
assign _2671_ = _2914_ ^ _2921_ /*94253*/;
assign _2919_ = _2920_ | _2922_ /*94250*/;
assign _2928_ = ~D[47] /*94249*/;
assign _2925_ = _2223_ & _2928_ /*94245*/;
assign _2926_ = _2223_ ^ _2928_ /*94248*/;
assign _2927_ = _2919_ & _2926_ /*94246*/;
assign _2672_ = _2919_ ^ _2926_ /*94247*/;
assign _2924_ = _2925_ | _2927_ /*94244*/;
assign _2933_ = ~D[48] /*94243*/;
assign _2930_ = _2224_ & _2933_ /*94239*/;
assign _2931_ = _2224_ ^ _2933_ /*94242*/;
assign _2932_ = _2924_ & _2931_ /*94240*/;
assign _2673_ = _2924_ ^ _2931_ /*94241*/;
assign _2929_ = _2930_ | _2932_ /*94238*/;
assign _2938_ = ~D[49] /*94237*/;
assign _2935_ = _2225_ & _2938_ /*94233*/;
assign _2936_ = _2225_ ^ _2938_ /*94236*/;
assign _2937_ = _2929_ & _2936_ /*94234*/;
assign _2674_ = _2929_ ^ _2936_ /*94235*/;
assign _2934_ = _2935_ | _2937_ /*94232*/;
assign _2943_ = ~D[50] /*94231*/;
assign _2940_ = _2226_ & _2943_ /*94227*/;
assign _2941_ = _2226_ ^ _2943_ /*94230*/;
assign _2942_ = _2934_ & _2941_ /*94228*/;
assign _2675_ = _2934_ ^ _2941_ /*94229*/;
assign _2939_ = _2940_ | _2942_ /*94226*/;
assign _2948_ = ~D[51] /*94225*/;
assign _2945_ = _2227_ & _2948_ /*94221*/;
assign _2946_ = _2227_ ^ _2948_ /*94224*/;
assign _2947_ = _2939_ & _2946_ /*94222*/;
assign _2676_ = _2939_ ^ _2946_ /*94223*/;
assign _2944_ = _2945_ | _2947_ /*94220*/;
assign _2953_ = ~D[52] /*94219*/;
assign _2950_ = _2228_ & _2953_ /*94215*/;
assign _2951_ = _2228_ ^ _2953_ /*94218*/;
assign _2952_ = _2944_ & _2951_ /*94216*/;
assign _2677_ = _2944_ ^ _2951_ /*94217*/;
assign _2949_ = _2950_ | _2952_ /*94214*/;
assign _2958_ = ~D[53] /*94213*/;
assign _2955_ = _2229_ & _2958_ /*94209*/;
assign _2956_ = _2229_ ^ _2958_ /*94212*/;
assign _2957_ = _2949_ & _2956_ /*94210*/;
assign _2678_ = _2949_ ^ _2956_ /*94211*/;
assign _2954_ = _2955_ | _2957_ /*94208*/;
assign _2963_ = ~D[54] /*94207*/;
assign _2960_ = _2230_ & _2963_ /*94203*/;
assign _2961_ = _2230_ ^ _2963_ /*94206*/;
assign _2962_ = _2954_ & _2961_ /*94204*/;
assign _2679_ = _2954_ ^ _2961_ /*94205*/;
assign _2959_ = _2960_ | _2962_ /*94202*/;
assign _2968_ = ~D[55] /*94201*/;
assign _2965_ = _2231_ & _2968_ /*94197*/;
assign _2966_ = _2231_ ^ _2968_ /*94200*/;
assign _2967_ = _2959_ & _2966_ /*94198*/;
assign _2680_ = _2959_ ^ _2966_ /*94199*/;
assign _2964_ = _2965_ | _2967_ /*94196*/;
assign _2973_ = ~D[56] /*94195*/;
assign _2970_ = _2232_ & _2973_ /*94191*/;
assign _2971_ = _2232_ ^ _2973_ /*94194*/;
assign _2972_ = _2964_ & _2971_ /*94192*/;
assign _2681_ = _2964_ ^ _2971_ /*94193*/;
assign _2969_ = _2970_ | _2972_ /*94190*/;
assign _2978_ = ~D[57] /*94189*/;
assign _2975_ = _2233_ & _2978_ /*94185*/;
assign _2976_ = _2233_ ^ _2978_ /*94188*/;
assign _2977_ = _2969_ & _2976_ /*94186*/;
assign _2682_ = _2969_ ^ _2976_ /*94187*/;
assign _2974_ = _2975_ | _2977_ /*94184*/;
assign _2983_ = ~D[58] /*94183*/;
assign _2980_ = _2234_ & _2983_ /*94179*/;
assign _2981_ = _2234_ ^ _2983_ /*94182*/;
assign _2982_ = _2974_ & _2981_ /*94180*/;
assign _2683_ = _2974_ ^ _2981_ /*94181*/;
assign _2979_ = _2980_ | _2982_ /*94178*/;
assign _2988_ = ~D[59] /*94177*/;
assign _2985_ = _2235_ & _2988_ /*94173*/;
assign _2986_ = _2235_ ^ _2988_ /*94176*/;
assign _2987_ = _2979_ & _2986_ /*94174*/;
assign _2684_ = _2979_ ^ _2986_ /*94175*/;
assign _2984_ = _2985_ | _2987_ /*94172*/;
assign _2993_ = ~D[60] /*94171*/;
assign _2990_ = _2236_ & _2993_ /*94167*/;
assign _2991_ = _2236_ ^ _2993_ /*94170*/;
assign _2992_ = _2984_ & _2991_ /*94168*/;
assign _2685_ = _2984_ ^ _2991_ /*94169*/;
assign _2989_ = _2990_ | _2992_ /*94166*/;
assign _2998_ = ~D[61] /*94165*/;
assign _2995_ = _2237_ & _2998_ /*94161*/;
assign _2996_ = _2237_ ^ _2998_ /*94164*/;
assign _2997_ = _2989_ & _2996_ /*94162*/;
assign _2686_ = _2989_ ^ _2996_ /*94163*/;
assign _2994_ = _2995_ | _2997_ /*94160*/;
assign _3003_ = ~D[62] /*94159*/;
assign _3000_ = _2238_ & _3003_ /*94155*/;
assign _3001_ = _2238_ ^ _3003_ /*94158*/;
assign _3002_ = _2994_ & _3001_ /*94156*/;
assign _2687_ = _2994_ ^ _3001_ /*94157*/;
assign _2999_ = _3000_ | _3002_ /*94154*/;
assign _3004_ = _2239_ & oneWire /*94149*/;
assign _3005_ = _2239_ ^ oneWire /*94152*/;
assign _3006_ = _2999_ & _3005_ /*94150*/;
assign _2688_ = _2999_ ^ _3005_ /*94151*/;
assign Q[60] = _3004_ | _3006_ /*94148*/;
assign _3139_ = ~Q[60] /*93763*/;
assign _3138_ = _3139_ & D[0] /*93762*/;
assign _3141_ = _2625_ & _3138_ /*93757*/;
assign _3142_ = _2625_ ^ _3138_ /*93760*/;
assign _3143_ = zeroWire & _3142_ /*93758*/;
assign _3073_ = zeroWire ^ _3142_ /*93759*/;
assign _3140_ = _3141_ | _3143_ /*93756*/;
assign _3145_ = ~Q[60] /*93755*/;
assign _3144_ = _3145_ & D[1] /*93754*/;
assign _3147_ = _2626_ & _3144_ /*93749*/;
assign _3148_ = _2626_ ^ _3144_ /*93752*/;
assign _3149_ = _3140_ & _3148_ /*93750*/;
assign _3074_ = _3140_ ^ _3148_ /*93751*/;
assign _3146_ = _3147_ | _3149_ /*93748*/;
assign _3151_ = ~Q[60] /*93747*/;
assign _3150_ = _3151_ & D[2] /*93746*/;
assign _3153_ = _2627_ & _3150_ /*93741*/;
assign _3154_ = _2627_ ^ _3150_ /*93744*/;
assign _3155_ = _3146_ & _3154_ /*93742*/;
assign _3075_ = _3146_ ^ _3154_ /*93743*/;
assign _3152_ = _3153_ | _3155_ /*93740*/;
assign _3157_ = ~Q[60] /*93739*/;
assign _3156_ = _3157_ & D[3] /*93738*/;
assign _3159_ = _2628_ & _3156_ /*93733*/;
assign _3160_ = _2628_ ^ _3156_ /*93736*/;
assign _3161_ = _3152_ & _3160_ /*93734*/;
assign _3076_ = _3152_ ^ _3160_ /*93735*/;
assign _3158_ = _3159_ | _3161_ /*93732*/;
assign _3163_ = ~Q[60] /*93731*/;
assign _3162_ = _3163_ & D[4] /*93730*/;
assign _3165_ = _2629_ & _3162_ /*93725*/;
assign _3166_ = _2629_ ^ _3162_ /*93728*/;
assign _3167_ = _3158_ & _3166_ /*93726*/;
assign _3077_ = _3158_ ^ _3166_ /*93727*/;
assign _3164_ = _3165_ | _3167_ /*93724*/;
assign _3169_ = ~Q[60] /*93723*/;
assign _3168_ = _3169_ & D[5] /*93722*/;
assign _3171_ = _2630_ & _3168_ /*93717*/;
assign _3172_ = _2630_ ^ _3168_ /*93720*/;
assign _3173_ = _3164_ & _3172_ /*93718*/;
assign _3078_ = _3164_ ^ _3172_ /*93719*/;
assign _3170_ = _3171_ | _3173_ /*93716*/;
assign _3175_ = ~Q[60] /*93715*/;
assign _3174_ = _3175_ & D[6] /*93714*/;
assign _3177_ = _2631_ & _3174_ /*93709*/;
assign _3178_ = _2631_ ^ _3174_ /*93712*/;
assign _3179_ = _3170_ & _3178_ /*93710*/;
assign _3079_ = _3170_ ^ _3178_ /*93711*/;
assign _3176_ = _3177_ | _3179_ /*93708*/;
assign _3181_ = ~Q[60] /*93707*/;
assign _3180_ = _3181_ & D[7] /*93706*/;
assign _3183_ = _2632_ & _3180_ /*93701*/;
assign _3184_ = _2632_ ^ _3180_ /*93704*/;
assign _3185_ = _3176_ & _3184_ /*93702*/;
assign _3080_ = _3176_ ^ _3184_ /*93703*/;
assign _3182_ = _3183_ | _3185_ /*93700*/;
assign _3187_ = ~Q[60] /*93699*/;
assign _3186_ = _3187_ & D[8] /*93698*/;
assign _3189_ = _2633_ & _3186_ /*93693*/;
assign _3190_ = _2633_ ^ _3186_ /*93696*/;
assign _3191_ = _3182_ & _3190_ /*93694*/;
assign _3081_ = _3182_ ^ _3190_ /*93695*/;
assign _3188_ = _3189_ | _3191_ /*93692*/;
assign _3193_ = ~Q[60] /*93691*/;
assign _3192_ = _3193_ & D[9] /*93690*/;
assign _3195_ = _2634_ & _3192_ /*93685*/;
assign _3196_ = _2634_ ^ _3192_ /*93688*/;
assign _3197_ = _3188_ & _3196_ /*93686*/;
assign _3082_ = _3188_ ^ _3196_ /*93687*/;
assign _3194_ = _3195_ | _3197_ /*93684*/;
assign _3199_ = ~Q[60] /*93683*/;
assign _3198_ = _3199_ & D[10] /*93682*/;
assign _3201_ = _2635_ & _3198_ /*93677*/;
assign _3202_ = _2635_ ^ _3198_ /*93680*/;
assign _3203_ = _3194_ & _3202_ /*93678*/;
assign _3083_ = _3194_ ^ _3202_ /*93679*/;
assign _3200_ = _3201_ | _3203_ /*93676*/;
assign _3205_ = ~Q[60] /*93675*/;
assign _3204_ = _3205_ & D[11] /*93674*/;
assign _3207_ = _2636_ & _3204_ /*93669*/;
assign _3208_ = _2636_ ^ _3204_ /*93672*/;
assign _3209_ = _3200_ & _3208_ /*93670*/;
assign _3084_ = _3200_ ^ _3208_ /*93671*/;
assign _3206_ = _3207_ | _3209_ /*93668*/;
assign _3211_ = ~Q[60] /*93667*/;
assign _3210_ = _3211_ & D[12] /*93666*/;
assign _3213_ = _2637_ & _3210_ /*93661*/;
assign _3214_ = _2637_ ^ _3210_ /*93664*/;
assign _3215_ = _3206_ & _3214_ /*93662*/;
assign _3085_ = _3206_ ^ _3214_ /*93663*/;
assign _3212_ = _3213_ | _3215_ /*93660*/;
assign _3217_ = ~Q[60] /*93659*/;
assign _3216_ = _3217_ & D[13] /*93658*/;
assign _3219_ = _2638_ & _3216_ /*93653*/;
assign _3220_ = _2638_ ^ _3216_ /*93656*/;
assign _3221_ = _3212_ & _3220_ /*93654*/;
assign _3086_ = _3212_ ^ _3220_ /*93655*/;
assign _3218_ = _3219_ | _3221_ /*93652*/;
assign _3223_ = ~Q[60] /*93651*/;
assign _3222_ = _3223_ & D[14] /*93650*/;
assign _3225_ = _2639_ & _3222_ /*93645*/;
assign _3226_ = _2639_ ^ _3222_ /*93648*/;
assign _3227_ = _3218_ & _3226_ /*93646*/;
assign _3087_ = _3218_ ^ _3226_ /*93647*/;
assign _3224_ = _3225_ | _3227_ /*93644*/;
assign _3229_ = ~Q[60] /*93643*/;
assign _3228_ = _3229_ & D[15] /*93642*/;
assign _3231_ = _2640_ & _3228_ /*93637*/;
assign _3232_ = _2640_ ^ _3228_ /*93640*/;
assign _3233_ = _3224_ & _3232_ /*93638*/;
assign _3088_ = _3224_ ^ _3232_ /*93639*/;
assign _3230_ = _3231_ | _3233_ /*93636*/;
assign _3235_ = ~Q[60] /*93635*/;
assign _3234_ = _3235_ & D[16] /*93634*/;
assign _3237_ = _2641_ & _3234_ /*93629*/;
assign _3238_ = _2641_ ^ _3234_ /*93632*/;
assign _3239_ = _3230_ & _3238_ /*93630*/;
assign _3089_ = _3230_ ^ _3238_ /*93631*/;
assign _3236_ = _3237_ | _3239_ /*93628*/;
assign _3241_ = ~Q[60] /*93627*/;
assign _3240_ = _3241_ & D[17] /*93626*/;
assign _3243_ = _2642_ & _3240_ /*93621*/;
assign _3244_ = _2642_ ^ _3240_ /*93624*/;
assign _3245_ = _3236_ & _3244_ /*93622*/;
assign _3090_ = _3236_ ^ _3244_ /*93623*/;
assign _3242_ = _3243_ | _3245_ /*93620*/;
assign _3247_ = ~Q[60] /*93619*/;
assign _3246_ = _3247_ & D[18] /*93618*/;
assign _3249_ = _2643_ & _3246_ /*93613*/;
assign _3250_ = _2643_ ^ _3246_ /*93616*/;
assign _3251_ = _3242_ & _3250_ /*93614*/;
assign _3091_ = _3242_ ^ _3250_ /*93615*/;
assign _3248_ = _3249_ | _3251_ /*93612*/;
assign _3253_ = ~Q[60] /*93611*/;
assign _3252_ = _3253_ & D[19] /*93610*/;
assign _3255_ = _2644_ & _3252_ /*93605*/;
assign _3256_ = _2644_ ^ _3252_ /*93608*/;
assign _3257_ = _3248_ & _3256_ /*93606*/;
assign _3092_ = _3248_ ^ _3256_ /*93607*/;
assign _3254_ = _3255_ | _3257_ /*93604*/;
assign _3259_ = ~Q[60] /*93603*/;
assign _3258_ = _3259_ & D[20] /*93602*/;
assign _3261_ = _2645_ & _3258_ /*93597*/;
assign _3262_ = _2645_ ^ _3258_ /*93600*/;
assign _3263_ = _3254_ & _3262_ /*93598*/;
assign _3093_ = _3254_ ^ _3262_ /*93599*/;
assign _3260_ = _3261_ | _3263_ /*93596*/;
assign _3265_ = ~Q[60] /*93595*/;
assign _3264_ = _3265_ & D[21] /*93594*/;
assign _3267_ = _2646_ & _3264_ /*93589*/;
assign _3268_ = _2646_ ^ _3264_ /*93592*/;
assign _3269_ = _3260_ & _3268_ /*93590*/;
assign _3094_ = _3260_ ^ _3268_ /*93591*/;
assign _3266_ = _3267_ | _3269_ /*93588*/;
assign _3271_ = ~Q[60] /*93587*/;
assign _3270_ = _3271_ & D[22] /*93586*/;
assign _3273_ = _2647_ & _3270_ /*93581*/;
assign _3274_ = _2647_ ^ _3270_ /*93584*/;
assign _3275_ = _3266_ & _3274_ /*93582*/;
assign _3095_ = _3266_ ^ _3274_ /*93583*/;
assign _3272_ = _3273_ | _3275_ /*93580*/;
assign _3277_ = ~Q[60] /*93579*/;
assign _3276_ = _3277_ & D[23] /*93578*/;
assign _3279_ = _2648_ & _3276_ /*93573*/;
assign _3280_ = _2648_ ^ _3276_ /*93576*/;
assign _3281_ = _3272_ & _3280_ /*93574*/;
assign _3096_ = _3272_ ^ _3280_ /*93575*/;
assign _3278_ = _3279_ | _3281_ /*93572*/;
assign _3283_ = ~Q[60] /*93571*/;
assign _3282_ = _3283_ & D[24] /*93570*/;
assign _3285_ = _2649_ & _3282_ /*93565*/;
assign _3286_ = _2649_ ^ _3282_ /*93568*/;
assign _3287_ = _3278_ & _3286_ /*93566*/;
assign _3097_ = _3278_ ^ _3286_ /*93567*/;
assign _3284_ = _3285_ | _3287_ /*93564*/;
assign _3289_ = ~Q[60] /*93563*/;
assign _3288_ = _3289_ & D[25] /*93562*/;
assign _3291_ = _2650_ & _3288_ /*93557*/;
assign _3292_ = _2650_ ^ _3288_ /*93560*/;
assign _3293_ = _3284_ & _3292_ /*93558*/;
assign _3098_ = _3284_ ^ _3292_ /*93559*/;
assign _3290_ = _3291_ | _3293_ /*93556*/;
assign _3295_ = ~Q[60] /*93555*/;
assign _3294_ = _3295_ & D[26] /*93554*/;
assign _3297_ = _2651_ & _3294_ /*93549*/;
assign _3298_ = _2651_ ^ _3294_ /*93552*/;
assign _3299_ = _3290_ & _3298_ /*93550*/;
assign _3099_ = _3290_ ^ _3298_ /*93551*/;
assign _3296_ = _3297_ | _3299_ /*93548*/;
assign _3301_ = ~Q[60] /*93547*/;
assign _3300_ = _3301_ & D[27] /*93546*/;
assign _3303_ = _2652_ & _3300_ /*93541*/;
assign _3304_ = _2652_ ^ _3300_ /*93544*/;
assign _3305_ = _3296_ & _3304_ /*93542*/;
assign _3100_ = _3296_ ^ _3304_ /*93543*/;
assign _3302_ = _3303_ | _3305_ /*93540*/;
assign _3307_ = ~Q[60] /*93539*/;
assign _3306_ = _3307_ & D[28] /*93538*/;
assign _3309_ = _2653_ & _3306_ /*93533*/;
assign _3310_ = _2653_ ^ _3306_ /*93536*/;
assign _3311_ = _3302_ & _3310_ /*93534*/;
assign _3101_ = _3302_ ^ _3310_ /*93535*/;
assign _3308_ = _3309_ | _3311_ /*93532*/;
assign _3313_ = ~Q[60] /*93531*/;
assign _3312_ = _3313_ & D[29] /*93530*/;
assign _3315_ = _2654_ & _3312_ /*93525*/;
assign _3316_ = _2654_ ^ _3312_ /*93528*/;
assign _3317_ = _3308_ & _3316_ /*93526*/;
assign _3102_ = _3308_ ^ _3316_ /*93527*/;
assign _3314_ = _3315_ | _3317_ /*93524*/;
assign _3319_ = ~Q[60] /*93523*/;
assign _3318_ = _3319_ & D[30] /*93522*/;
assign _3321_ = _2655_ & _3318_ /*93517*/;
assign _3322_ = _2655_ ^ _3318_ /*93520*/;
assign _3323_ = _3314_ & _3322_ /*93518*/;
assign _3103_ = _3314_ ^ _3322_ /*93519*/;
assign _3320_ = _3321_ | _3323_ /*93516*/;
assign _3325_ = ~Q[60] /*93515*/;
assign _3324_ = _3325_ & D[31] /*93514*/;
assign _3327_ = _2656_ & _3324_ /*93509*/;
assign _3328_ = _2656_ ^ _3324_ /*93512*/;
assign _3329_ = _3320_ & _3328_ /*93510*/;
assign _3104_ = _3320_ ^ _3328_ /*93511*/;
assign _3326_ = _3327_ | _3329_ /*93508*/;
assign _3331_ = ~Q[60] /*93507*/;
assign _3330_ = _3331_ & D[32] /*93506*/;
assign _3333_ = _2657_ & _3330_ /*93501*/;
assign _3334_ = _2657_ ^ _3330_ /*93504*/;
assign _3335_ = _3326_ & _3334_ /*93502*/;
assign _3105_ = _3326_ ^ _3334_ /*93503*/;
assign _3332_ = _3333_ | _3335_ /*93500*/;
assign _3337_ = ~Q[60] /*93499*/;
assign _3336_ = _3337_ & D[33] /*93498*/;
assign _3339_ = _2658_ & _3336_ /*93493*/;
assign _3340_ = _2658_ ^ _3336_ /*93496*/;
assign _3341_ = _3332_ & _3340_ /*93494*/;
assign _3106_ = _3332_ ^ _3340_ /*93495*/;
assign _3338_ = _3339_ | _3341_ /*93492*/;
assign _3343_ = ~Q[60] /*93491*/;
assign _3342_ = _3343_ & D[34] /*93490*/;
assign _3345_ = _2659_ & _3342_ /*93485*/;
assign _3346_ = _2659_ ^ _3342_ /*93488*/;
assign _3347_ = _3338_ & _3346_ /*93486*/;
assign _3107_ = _3338_ ^ _3346_ /*93487*/;
assign _3344_ = _3345_ | _3347_ /*93484*/;
assign _3349_ = ~Q[60] /*93483*/;
assign _3348_ = _3349_ & D[35] /*93482*/;
assign _3351_ = _2660_ & _3348_ /*93477*/;
assign _3352_ = _2660_ ^ _3348_ /*93480*/;
assign _3353_ = _3344_ & _3352_ /*93478*/;
assign _3108_ = _3344_ ^ _3352_ /*93479*/;
assign _3350_ = _3351_ | _3353_ /*93476*/;
assign _3355_ = ~Q[60] /*93475*/;
assign _3354_ = _3355_ & D[36] /*93474*/;
assign _3357_ = _2661_ & _3354_ /*93469*/;
assign _3358_ = _2661_ ^ _3354_ /*93472*/;
assign _3359_ = _3350_ & _3358_ /*93470*/;
assign _3109_ = _3350_ ^ _3358_ /*93471*/;
assign _3356_ = _3357_ | _3359_ /*93468*/;
assign _3361_ = ~Q[60] /*93467*/;
assign _3360_ = _3361_ & D[37] /*93466*/;
assign _3363_ = _2662_ & _3360_ /*93461*/;
assign _3364_ = _2662_ ^ _3360_ /*93464*/;
assign _3365_ = _3356_ & _3364_ /*93462*/;
assign _3110_ = _3356_ ^ _3364_ /*93463*/;
assign _3362_ = _3363_ | _3365_ /*93460*/;
assign _3367_ = ~Q[60] /*93459*/;
assign _3366_ = _3367_ & D[38] /*93458*/;
assign _3369_ = _2663_ & _3366_ /*93453*/;
assign _3370_ = _2663_ ^ _3366_ /*93456*/;
assign _3371_ = _3362_ & _3370_ /*93454*/;
assign _3111_ = _3362_ ^ _3370_ /*93455*/;
assign _3368_ = _3369_ | _3371_ /*93452*/;
assign _3373_ = ~Q[60] /*93451*/;
assign _3372_ = _3373_ & D[39] /*93450*/;
assign _3375_ = _2664_ & _3372_ /*93445*/;
assign _3376_ = _2664_ ^ _3372_ /*93448*/;
assign _3377_ = _3368_ & _3376_ /*93446*/;
assign _3112_ = _3368_ ^ _3376_ /*93447*/;
assign _3374_ = _3375_ | _3377_ /*93444*/;
assign _3379_ = ~Q[60] /*93443*/;
assign _3378_ = _3379_ & D[40] /*93442*/;
assign _3381_ = _2665_ & _3378_ /*93437*/;
assign _3382_ = _2665_ ^ _3378_ /*93440*/;
assign _3383_ = _3374_ & _3382_ /*93438*/;
assign _3113_ = _3374_ ^ _3382_ /*93439*/;
assign _3380_ = _3381_ | _3383_ /*93436*/;
assign _3385_ = ~Q[60] /*93435*/;
assign _3384_ = _3385_ & D[41] /*93434*/;
assign _3387_ = _2666_ & _3384_ /*93429*/;
assign _3388_ = _2666_ ^ _3384_ /*93432*/;
assign _3389_ = _3380_ & _3388_ /*93430*/;
assign _3114_ = _3380_ ^ _3388_ /*93431*/;
assign _3386_ = _3387_ | _3389_ /*93428*/;
assign _3391_ = ~Q[60] /*93427*/;
assign _3390_ = _3391_ & D[42] /*93426*/;
assign _3393_ = _2667_ & _3390_ /*93421*/;
assign _3394_ = _2667_ ^ _3390_ /*93424*/;
assign _3395_ = _3386_ & _3394_ /*93422*/;
assign _3115_ = _3386_ ^ _3394_ /*93423*/;
assign _3392_ = _3393_ | _3395_ /*93420*/;
assign _3397_ = ~Q[60] /*93419*/;
assign _3396_ = _3397_ & D[43] /*93418*/;
assign _3399_ = _2668_ & _3396_ /*93413*/;
assign _3400_ = _2668_ ^ _3396_ /*93416*/;
assign _3401_ = _3392_ & _3400_ /*93414*/;
assign _3116_ = _3392_ ^ _3400_ /*93415*/;
assign _3398_ = _3399_ | _3401_ /*93412*/;
assign _3403_ = ~Q[60] /*93411*/;
assign _3402_ = _3403_ & D[44] /*93410*/;
assign _3405_ = _2669_ & _3402_ /*93405*/;
assign _3406_ = _2669_ ^ _3402_ /*93408*/;
assign _3407_ = _3398_ & _3406_ /*93406*/;
assign _3117_ = _3398_ ^ _3406_ /*93407*/;
assign _3404_ = _3405_ | _3407_ /*93404*/;
assign _3409_ = ~Q[60] /*93403*/;
assign _3408_ = _3409_ & D[45] /*93402*/;
assign _3411_ = _2670_ & _3408_ /*93397*/;
assign _3412_ = _2670_ ^ _3408_ /*93400*/;
assign _3413_ = _3404_ & _3412_ /*93398*/;
assign _3118_ = _3404_ ^ _3412_ /*93399*/;
assign _3410_ = _3411_ | _3413_ /*93396*/;
assign _3415_ = ~Q[60] /*93395*/;
assign _3414_ = _3415_ & D[46] /*93394*/;
assign _3417_ = _2671_ & _3414_ /*93389*/;
assign _3418_ = _2671_ ^ _3414_ /*93392*/;
assign _3419_ = _3410_ & _3418_ /*93390*/;
assign _3119_ = _3410_ ^ _3418_ /*93391*/;
assign _3416_ = _3417_ | _3419_ /*93388*/;
assign _3421_ = ~Q[60] /*93387*/;
assign _3420_ = _3421_ & D[47] /*93386*/;
assign _3423_ = _2672_ & _3420_ /*93381*/;
assign _3424_ = _2672_ ^ _3420_ /*93384*/;
assign _3425_ = _3416_ & _3424_ /*93382*/;
assign _3120_ = _3416_ ^ _3424_ /*93383*/;
assign _3422_ = _3423_ | _3425_ /*93380*/;
assign _3427_ = ~Q[60] /*93379*/;
assign _3426_ = _3427_ & D[48] /*93378*/;
assign _3429_ = _2673_ & _3426_ /*93373*/;
assign _3430_ = _2673_ ^ _3426_ /*93376*/;
assign _3431_ = _3422_ & _3430_ /*93374*/;
assign _3121_ = _3422_ ^ _3430_ /*93375*/;
assign _3428_ = _3429_ | _3431_ /*93372*/;
assign _3433_ = ~Q[60] /*93371*/;
assign _3432_ = _3433_ & D[49] /*93370*/;
assign _3435_ = _2674_ & _3432_ /*93365*/;
assign _3436_ = _2674_ ^ _3432_ /*93368*/;
assign _3437_ = _3428_ & _3436_ /*93366*/;
assign _3122_ = _3428_ ^ _3436_ /*93367*/;
assign _3434_ = _3435_ | _3437_ /*93364*/;
assign _3439_ = ~Q[60] /*93363*/;
assign _3438_ = _3439_ & D[50] /*93362*/;
assign _3441_ = _2675_ & _3438_ /*93357*/;
assign _3442_ = _2675_ ^ _3438_ /*93360*/;
assign _3443_ = _3434_ & _3442_ /*93358*/;
assign _3123_ = _3434_ ^ _3442_ /*93359*/;
assign _3440_ = _3441_ | _3443_ /*93356*/;
assign _3445_ = ~Q[60] /*93355*/;
assign _3444_ = _3445_ & D[51] /*93354*/;
assign _3447_ = _2676_ & _3444_ /*93349*/;
assign _3448_ = _2676_ ^ _3444_ /*93352*/;
assign _3449_ = _3440_ & _3448_ /*93350*/;
assign _3124_ = _3440_ ^ _3448_ /*93351*/;
assign _3446_ = _3447_ | _3449_ /*93348*/;
assign _3451_ = ~Q[60] /*93347*/;
assign _3450_ = _3451_ & D[52] /*93346*/;
assign _3453_ = _2677_ & _3450_ /*93341*/;
assign _3454_ = _2677_ ^ _3450_ /*93344*/;
assign _3455_ = _3446_ & _3454_ /*93342*/;
assign _3125_ = _3446_ ^ _3454_ /*93343*/;
assign _3452_ = _3453_ | _3455_ /*93340*/;
assign _3457_ = ~Q[60] /*93339*/;
assign _3456_ = _3457_ & D[53] /*93338*/;
assign _3459_ = _2678_ & _3456_ /*93333*/;
assign _3460_ = _2678_ ^ _3456_ /*93336*/;
assign _3461_ = _3452_ & _3460_ /*93334*/;
assign _3126_ = _3452_ ^ _3460_ /*93335*/;
assign _3458_ = _3459_ | _3461_ /*93332*/;
assign _3463_ = ~Q[60] /*93331*/;
assign _3462_ = _3463_ & D[54] /*93330*/;
assign _3465_ = _2679_ & _3462_ /*93325*/;
assign _3466_ = _2679_ ^ _3462_ /*93328*/;
assign _3467_ = _3458_ & _3466_ /*93326*/;
assign _3127_ = _3458_ ^ _3466_ /*93327*/;
assign _3464_ = _3465_ | _3467_ /*93324*/;
assign _3469_ = ~Q[60] /*93323*/;
assign _3468_ = _3469_ & D[55] /*93322*/;
assign _3471_ = _2680_ & _3468_ /*93317*/;
assign _3472_ = _2680_ ^ _3468_ /*93320*/;
assign _3473_ = _3464_ & _3472_ /*93318*/;
assign _3128_ = _3464_ ^ _3472_ /*93319*/;
assign _3470_ = _3471_ | _3473_ /*93316*/;
assign _3475_ = ~Q[60] /*93315*/;
assign _3474_ = _3475_ & D[56] /*93314*/;
assign _3477_ = _2681_ & _3474_ /*93309*/;
assign _3478_ = _2681_ ^ _3474_ /*93312*/;
assign _3479_ = _3470_ & _3478_ /*93310*/;
assign _3129_ = _3470_ ^ _3478_ /*93311*/;
assign _3476_ = _3477_ | _3479_ /*93308*/;
assign _3481_ = ~Q[60] /*93307*/;
assign _3480_ = _3481_ & D[57] /*93306*/;
assign _3483_ = _2682_ & _3480_ /*93301*/;
assign _3484_ = _2682_ ^ _3480_ /*93304*/;
assign _3485_ = _3476_ & _3484_ /*93302*/;
assign _3130_ = _3476_ ^ _3484_ /*93303*/;
assign _3482_ = _3483_ | _3485_ /*93300*/;
assign _3487_ = ~Q[60] /*93299*/;
assign _3486_ = _3487_ & D[58] /*93298*/;
assign _3489_ = _2683_ & _3486_ /*93293*/;
assign _3490_ = _2683_ ^ _3486_ /*93296*/;
assign _3491_ = _3482_ & _3490_ /*93294*/;
assign _3131_ = _3482_ ^ _3490_ /*93295*/;
assign _3488_ = _3489_ | _3491_ /*93292*/;
assign _3493_ = ~Q[60] /*93291*/;
assign _3492_ = _3493_ & D[59] /*93290*/;
assign _3495_ = _2684_ & _3492_ /*93285*/;
assign _3496_ = _2684_ ^ _3492_ /*93288*/;
assign _3497_ = _3488_ & _3496_ /*93286*/;
assign _3132_ = _3488_ ^ _3496_ /*93287*/;
assign _3494_ = _3495_ | _3497_ /*93284*/;
assign _3499_ = ~Q[60] /*93283*/;
assign _3498_ = _3499_ & D[60] /*93282*/;
assign _3501_ = _2685_ & _3498_ /*93277*/;
assign _3502_ = _2685_ ^ _3498_ /*93280*/;
assign _3503_ = _3494_ & _3502_ /*93278*/;
assign _3133_ = _3494_ ^ _3502_ /*93279*/;
assign _3500_ = _3501_ | _3503_ /*93276*/;
assign _3505_ = ~Q[60] /*93275*/;
assign _3504_ = _3505_ & D[61] /*93274*/;
assign _3507_ = _2686_ & _3504_ /*93269*/;
assign _3508_ = _2686_ ^ _3504_ /*93272*/;
assign _3509_ = _3500_ & _3508_ /*93270*/;
assign _3134_ = _3500_ ^ _3508_ /*93271*/;
assign _3506_ = _3507_ | _3509_ /*93268*/;
assign _3511_ = ~Q[60] /*93267*/;
assign _3510_ = _3511_ & D[62] /*93266*/;
assign _3513_ = _2687_ & _3510_ /*93261*/;
assign _3514_ = _2687_ ^ _3510_ /*93264*/;
assign _3515_ = _3506_ & _3514_ /*93262*/;
assign _3135_ = _3506_ ^ _3514_ /*93263*/;
assign _3512_ = _3513_ | _3515_ /*93260*/;
assign _3517_ = ~Q[60] /*93259*/;
assign _3516_ = _3517_ & zeroWire /*93258*/;
assign _3518_ = _2688_ ^ _3516_ /*93256*/;
assign _3136_ = _3518_ ^ _3512_ /*93255*/;
assign _3589_ = ~D[0] /*93001*/;
assign _3586_ = R_0[59] & _3589_ /*92997*/;
assign _3587_ = R_0[59] ^ _3589_ /*93000*/;
assign _3588_ = oneWire & _3587_ /*92998*/;
assign _3521_ = oneWire ^ _3587_ /*92999*/;
assign _3585_ = _3586_ | _3588_ /*92996*/;
assign _3594_ = ~D[1] /*92995*/;
assign _3591_ = _3073_ & _3594_ /*92991*/;
assign _3592_ = _3073_ ^ _3594_ /*92994*/;
assign _3593_ = _3585_ & _3592_ /*92992*/;
assign _3522_ = _3585_ ^ _3592_ /*92993*/;
assign _3590_ = _3591_ | _3593_ /*92990*/;
assign _3599_ = ~D[2] /*92989*/;
assign _3596_ = _3074_ & _3599_ /*92985*/;
assign _3597_ = _3074_ ^ _3599_ /*92988*/;
assign _3598_ = _3590_ & _3597_ /*92986*/;
assign _3523_ = _3590_ ^ _3597_ /*92987*/;
assign _3595_ = _3596_ | _3598_ /*92984*/;
assign _3604_ = ~D[3] /*92983*/;
assign _3601_ = _3075_ & _3604_ /*92979*/;
assign _3602_ = _3075_ ^ _3604_ /*92982*/;
assign _3603_ = _3595_ & _3602_ /*92980*/;
assign _3524_ = _3595_ ^ _3602_ /*92981*/;
assign _3600_ = _3601_ | _3603_ /*92978*/;
assign _3609_ = ~D[4] /*92977*/;
assign _3606_ = _3076_ & _3609_ /*92973*/;
assign _3607_ = _3076_ ^ _3609_ /*92976*/;
assign _3608_ = _3600_ & _3607_ /*92974*/;
assign _3525_ = _3600_ ^ _3607_ /*92975*/;
assign _3605_ = _3606_ | _3608_ /*92972*/;
assign _3614_ = ~D[5] /*92971*/;
assign _3611_ = _3077_ & _3614_ /*92967*/;
assign _3612_ = _3077_ ^ _3614_ /*92970*/;
assign _3613_ = _3605_ & _3612_ /*92968*/;
assign _3526_ = _3605_ ^ _3612_ /*92969*/;
assign _3610_ = _3611_ | _3613_ /*92966*/;
assign _3619_ = ~D[6] /*92965*/;
assign _3616_ = _3078_ & _3619_ /*92961*/;
assign _3617_ = _3078_ ^ _3619_ /*92964*/;
assign _3618_ = _3610_ & _3617_ /*92962*/;
assign _3527_ = _3610_ ^ _3617_ /*92963*/;
assign _3615_ = _3616_ | _3618_ /*92960*/;
assign _3624_ = ~D[7] /*92959*/;
assign _3621_ = _3079_ & _3624_ /*92955*/;
assign _3622_ = _3079_ ^ _3624_ /*92958*/;
assign _3623_ = _3615_ & _3622_ /*92956*/;
assign _3528_ = _3615_ ^ _3622_ /*92957*/;
assign _3620_ = _3621_ | _3623_ /*92954*/;
assign _3629_ = ~D[8] /*92953*/;
assign _3626_ = _3080_ & _3629_ /*92949*/;
assign _3627_ = _3080_ ^ _3629_ /*92952*/;
assign _3628_ = _3620_ & _3627_ /*92950*/;
assign _3529_ = _3620_ ^ _3627_ /*92951*/;
assign _3625_ = _3626_ | _3628_ /*92948*/;
assign _3634_ = ~D[9] /*92947*/;
assign _3631_ = _3081_ & _3634_ /*92943*/;
assign _3632_ = _3081_ ^ _3634_ /*92946*/;
assign _3633_ = _3625_ & _3632_ /*92944*/;
assign _3530_ = _3625_ ^ _3632_ /*92945*/;
assign _3630_ = _3631_ | _3633_ /*92942*/;
assign _3639_ = ~D[10] /*92941*/;
assign _3636_ = _3082_ & _3639_ /*92937*/;
assign _3637_ = _3082_ ^ _3639_ /*92940*/;
assign _3638_ = _3630_ & _3637_ /*92938*/;
assign _3531_ = _3630_ ^ _3637_ /*92939*/;
assign _3635_ = _3636_ | _3638_ /*92936*/;
assign _3644_ = ~D[11] /*92935*/;
assign _3641_ = _3083_ & _3644_ /*92931*/;
assign _3642_ = _3083_ ^ _3644_ /*92934*/;
assign _3643_ = _3635_ & _3642_ /*92932*/;
assign _3532_ = _3635_ ^ _3642_ /*92933*/;
assign _3640_ = _3641_ | _3643_ /*92930*/;
assign _3649_ = ~D[12] /*92929*/;
assign _3646_ = _3084_ & _3649_ /*92925*/;
assign _3647_ = _3084_ ^ _3649_ /*92928*/;
assign _3648_ = _3640_ & _3647_ /*92926*/;
assign _3533_ = _3640_ ^ _3647_ /*92927*/;
assign _3645_ = _3646_ | _3648_ /*92924*/;
assign _3654_ = ~D[13] /*92923*/;
assign _3651_ = _3085_ & _3654_ /*92919*/;
assign _3652_ = _3085_ ^ _3654_ /*92922*/;
assign _3653_ = _3645_ & _3652_ /*92920*/;
assign _3534_ = _3645_ ^ _3652_ /*92921*/;
assign _3650_ = _3651_ | _3653_ /*92918*/;
assign _3659_ = ~D[14] /*92917*/;
assign _3656_ = _3086_ & _3659_ /*92913*/;
assign _3657_ = _3086_ ^ _3659_ /*92916*/;
assign _3658_ = _3650_ & _3657_ /*92914*/;
assign _3535_ = _3650_ ^ _3657_ /*92915*/;
assign _3655_ = _3656_ | _3658_ /*92912*/;
assign _3664_ = ~D[15] /*92911*/;
assign _3661_ = _3087_ & _3664_ /*92907*/;
assign _3662_ = _3087_ ^ _3664_ /*92910*/;
assign _3663_ = _3655_ & _3662_ /*92908*/;
assign _3536_ = _3655_ ^ _3662_ /*92909*/;
assign _3660_ = _3661_ | _3663_ /*92906*/;
assign _3669_ = ~D[16] /*92905*/;
assign _3666_ = _3088_ & _3669_ /*92901*/;
assign _3667_ = _3088_ ^ _3669_ /*92904*/;
assign _3668_ = _3660_ & _3667_ /*92902*/;
assign _3537_ = _3660_ ^ _3667_ /*92903*/;
assign _3665_ = _3666_ | _3668_ /*92900*/;
assign _3674_ = ~D[17] /*92899*/;
assign _3671_ = _3089_ & _3674_ /*92895*/;
assign _3672_ = _3089_ ^ _3674_ /*92898*/;
assign _3673_ = _3665_ & _3672_ /*92896*/;
assign _3538_ = _3665_ ^ _3672_ /*92897*/;
assign _3670_ = _3671_ | _3673_ /*92894*/;
assign _3679_ = ~D[18] /*92893*/;
assign _3676_ = _3090_ & _3679_ /*92889*/;
assign _3677_ = _3090_ ^ _3679_ /*92892*/;
assign _3678_ = _3670_ & _3677_ /*92890*/;
assign _3539_ = _3670_ ^ _3677_ /*92891*/;
assign _3675_ = _3676_ | _3678_ /*92888*/;
assign _3684_ = ~D[19] /*92887*/;
assign _3681_ = _3091_ & _3684_ /*92883*/;
assign _3682_ = _3091_ ^ _3684_ /*92886*/;
assign _3683_ = _3675_ & _3682_ /*92884*/;
assign _3540_ = _3675_ ^ _3682_ /*92885*/;
assign _3680_ = _3681_ | _3683_ /*92882*/;
assign _3689_ = ~D[20] /*92881*/;
assign _3686_ = _3092_ & _3689_ /*92877*/;
assign _3687_ = _3092_ ^ _3689_ /*92880*/;
assign _3688_ = _3680_ & _3687_ /*92878*/;
assign _3541_ = _3680_ ^ _3687_ /*92879*/;
assign _3685_ = _3686_ | _3688_ /*92876*/;
assign _3694_ = ~D[21] /*92875*/;
assign _3691_ = _3093_ & _3694_ /*92871*/;
assign _3692_ = _3093_ ^ _3694_ /*92874*/;
assign _3693_ = _3685_ & _3692_ /*92872*/;
assign _3542_ = _3685_ ^ _3692_ /*92873*/;
assign _3690_ = _3691_ | _3693_ /*92870*/;
assign _3699_ = ~D[22] /*92869*/;
assign _3696_ = _3094_ & _3699_ /*92865*/;
assign _3697_ = _3094_ ^ _3699_ /*92868*/;
assign _3698_ = _3690_ & _3697_ /*92866*/;
assign _3543_ = _3690_ ^ _3697_ /*92867*/;
assign _3695_ = _3696_ | _3698_ /*92864*/;
assign _3704_ = ~D[23] /*92863*/;
assign _3701_ = _3095_ & _3704_ /*92859*/;
assign _3702_ = _3095_ ^ _3704_ /*92862*/;
assign _3703_ = _3695_ & _3702_ /*92860*/;
assign _3544_ = _3695_ ^ _3702_ /*92861*/;
assign _3700_ = _3701_ | _3703_ /*92858*/;
assign _3709_ = ~D[24] /*92857*/;
assign _3706_ = _3096_ & _3709_ /*92853*/;
assign _3707_ = _3096_ ^ _3709_ /*92856*/;
assign _3708_ = _3700_ & _3707_ /*92854*/;
assign _3545_ = _3700_ ^ _3707_ /*92855*/;
assign _3705_ = _3706_ | _3708_ /*92852*/;
assign _3714_ = ~D[25] /*92851*/;
assign _3711_ = _3097_ & _3714_ /*92847*/;
assign _3712_ = _3097_ ^ _3714_ /*92850*/;
assign _3713_ = _3705_ & _3712_ /*92848*/;
assign _3546_ = _3705_ ^ _3712_ /*92849*/;
assign _3710_ = _3711_ | _3713_ /*92846*/;
assign _3719_ = ~D[26] /*92845*/;
assign _3716_ = _3098_ & _3719_ /*92841*/;
assign _3717_ = _3098_ ^ _3719_ /*92844*/;
assign _3718_ = _3710_ & _3717_ /*92842*/;
assign _3547_ = _3710_ ^ _3717_ /*92843*/;
assign _3715_ = _3716_ | _3718_ /*92840*/;
assign _3724_ = ~D[27] /*92839*/;
assign _3721_ = _3099_ & _3724_ /*92835*/;
assign _3722_ = _3099_ ^ _3724_ /*92838*/;
assign _3723_ = _3715_ & _3722_ /*92836*/;
assign _3548_ = _3715_ ^ _3722_ /*92837*/;
assign _3720_ = _3721_ | _3723_ /*92834*/;
assign _3729_ = ~D[28] /*92833*/;
assign _3726_ = _3100_ & _3729_ /*92829*/;
assign _3727_ = _3100_ ^ _3729_ /*92832*/;
assign _3728_ = _3720_ & _3727_ /*92830*/;
assign _3549_ = _3720_ ^ _3727_ /*92831*/;
assign _3725_ = _3726_ | _3728_ /*92828*/;
assign _3734_ = ~D[29] /*92827*/;
assign _3731_ = _3101_ & _3734_ /*92823*/;
assign _3732_ = _3101_ ^ _3734_ /*92826*/;
assign _3733_ = _3725_ & _3732_ /*92824*/;
assign _3550_ = _3725_ ^ _3732_ /*92825*/;
assign _3730_ = _3731_ | _3733_ /*92822*/;
assign _3739_ = ~D[30] /*92821*/;
assign _3736_ = _3102_ & _3739_ /*92817*/;
assign _3737_ = _3102_ ^ _3739_ /*92820*/;
assign _3738_ = _3730_ & _3737_ /*92818*/;
assign _3551_ = _3730_ ^ _3737_ /*92819*/;
assign _3735_ = _3736_ | _3738_ /*92816*/;
assign _3744_ = ~D[31] /*92815*/;
assign _3741_ = _3103_ & _3744_ /*92811*/;
assign _3742_ = _3103_ ^ _3744_ /*92814*/;
assign _3743_ = _3735_ & _3742_ /*92812*/;
assign _3552_ = _3735_ ^ _3742_ /*92813*/;
assign _3740_ = _3741_ | _3743_ /*92810*/;
assign _3749_ = ~D[32] /*92809*/;
assign _3746_ = _3104_ & _3749_ /*92805*/;
assign _3747_ = _3104_ ^ _3749_ /*92808*/;
assign _3748_ = _3740_ & _3747_ /*92806*/;
assign _3553_ = _3740_ ^ _3747_ /*92807*/;
assign _3745_ = _3746_ | _3748_ /*92804*/;
assign _3754_ = ~D[33] /*92803*/;
assign _3751_ = _3105_ & _3754_ /*92799*/;
assign _3752_ = _3105_ ^ _3754_ /*92802*/;
assign _3753_ = _3745_ & _3752_ /*92800*/;
assign _3554_ = _3745_ ^ _3752_ /*92801*/;
assign _3750_ = _3751_ | _3753_ /*92798*/;
assign _3759_ = ~D[34] /*92797*/;
assign _3756_ = _3106_ & _3759_ /*92793*/;
assign _3757_ = _3106_ ^ _3759_ /*92796*/;
assign _3758_ = _3750_ & _3757_ /*92794*/;
assign _3555_ = _3750_ ^ _3757_ /*92795*/;
assign _3755_ = _3756_ | _3758_ /*92792*/;
assign _3764_ = ~D[35] /*92791*/;
assign _3761_ = _3107_ & _3764_ /*92787*/;
assign _3762_ = _3107_ ^ _3764_ /*92790*/;
assign _3763_ = _3755_ & _3762_ /*92788*/;
assign _3556_ = _3755_ ^ _3762_ /*92789*/;
assign _3760_ = _3761_ | _3763_ /*92786*/;
assign _3769_ = ~D[36] /*92785*/;
assign _3766_ = _3108_ & _3769_ /*92781*/;
assign _3767_ = _3108_ ^ _3769_ /*92784*/;
assign _3768_ = _3760_ & _3767_ /*92782*/;
assign _3557_ = _3760_ ^ _3767_ /*92783*/;
assign _3765_ = _3766_ | _3768_ /*92780*/;
assign _3774_ = ~D[37] /*92779*/;
assign _3771_ = _3109_ & _3774_ /*92775*/;
assign _3772_ = _3109_ ^ _3774_ /*92778*/;
assign _3773_ = _3765_ & _3772_ /*92776*/;
assign _3558_ = _3765_ ^ _3772_ /*92777*/;
assign _3770_ = _3771_ | _3773_ /*92774*/;
assign _3779_ = ~D[38] /*92773*/;
assign _3776_ = _3110_ & _3779_ /*92769*/;
assign _3777_ = _3110_ ^ _3779_ /*92772*/;
assign _3778_ = _3770_ & _3777_ /*92770*/;
assign _3559_ = _3770_ ^ _3777_ /*92771*/;
assign _3775_ = _3776_ | _3778_ /*92768*/;
assign _3784_ = ~D[39] /*92767*/;
assign _3781_ = _3111_ & _3784_ /*92763*/;
assign _3782_ = _3111_ ^ _3784_ /*92766*/;
assign _3783_ = _3775_ & _3782_ /*92764*/;
assign _3560_ = _3775_ ^ _3782_ /*92765*/;
assign _3780_ = _3781_ | _3783_ /*92762*/;
assign _3789_ = ~D[40] /*92761*/;
assign _3786_ = _3112_ & _3789_ /*92757*/;
assign _3787_ = _3112_ ^ _3789_ /*92760*/;
assign _3788_ = _3780_ & _3787_ /*92758*/;
assign _3561_ = _3780_ ^ _3787_ /*92759*/;
assign _3785_ = _3786_ | _3788_ /*92756*/;
assign _3794_ = ~D[41] /*92755*/;
assign _3791_ = _3113_ & _3794_ /*92751*/;
assign _3792_ = _3113_ ^ _3794_ /*92754*/;
assign _3793_ = _3785_ & _3792_ /*92752*/;
assign _3562_ = _3785_ ^ _3792_ /*92753*/;
assign _3790_ = _3791_ | _3793_ /*92750*/;
assign _3799_ = ~D[42] /*92749*/;
assign _3796_ = _3114_ & _3799_ /*92745*/;
assign _3797_ = _3114_ ^ _3799_ /*92748*/;
assign _3798_ = _3790_ & _3797_ /*92746*/;
assign _3563_ = _3790_ ^ _3797_ /*92747*/;
assign _3795_ = _3796_ | _3798_ /*92744*/;
assign _3804_ = ~D[43] /*92743*/;
assign _3801_ = _3115_ & _3804_ /*92739*/;
assign _3802_ = _3115_ ^ _3804_ /*92742*/;
assign _3803_ = _3795_ & _3802_ /*92740*/;
assign _3564_ = _3795_ ^ _3802_ /*92741*/;
assign _3800_ = _3801_ | _3803_ /*92738*/;
assign _3809_ = ~D[44] /*92737*/;
assign _3806_ = _3116_ & _3809_ /*92733*/;
assign _3807_ = _3116_ ^ _3809_ /*92736*/;
assign _3808_ = _3800_ & _3807_ /*92734*/;
assign _3565_ = _3800_ ^ _3807_ /*92735*/;
assign _3805_ = _3806_ | _3808_ /*92732*/;
assign _3814_ = ~D[45] /*92731*/;
assign _3811_ = _3117_ & _3814_ /*92727*/;
assign _3812_ = _3117_ ^ _3814_ /*92730*/;
assign _3813_ = _3805_ & _3812_ /*92728*/;
assign _3566_ = _3805_ ^ _3812_ /*92729*/;
assign _3810_ = _3811_ | _3813_ /*92726*/;
assign _3819_ = ~D[46] /*92725*/;
assign _3816_ = _3118_ & _3819_ /*92721*/;
assign _3817_ = _3118_ ^ _3819_ /*92724*/;
assign _3818_ = _3810_ & _3817_ /*92722*/;
assign _3567_ = _3810_ ^ _3817_ /*92723*/;
assign _3815_ = _3816_ | _3818_ /*92720*/;
assign _3824_ = ~D[47] /*92719*/;
assign _3821_ = _3119_ & _3824_ /*92715*/;
assign _3822_ = _3119_ ^ _3824_ /*92718*/;
assign _3823_ = _3815_ & _3822_ /*92716*/;
assign _3568_ = _3815_ ^ _3822_ /*92717*/;
assign _3820_ = _3821_ | _3823_ /*92714*/;
assign _3829_ = ~D[48] /*92713*/;
assign _3826_ = _3120_ & _3829_ /*92709*/;
assign _3827_ = _3120_ ^ _3829_ /*92712*/;
assign _3828_ = _3820_ & _3827_ /*92710*/;
assign _3569_ = _3820_ ^ _3827_ /*92711*/;
assign _3825_ = _3826_ | _3828_ /*92708*/;
assign _3834_ = ~D[49] /*92707*/;
assign _3831_ = _3121_ & _3834_ /*92703*/;
assign _3832_ = _3121_ ^ _3834_ /*92706*/;
assign _3833_ = _3825_ & _3832_ /*92704*/;
assign _3570_ = _3825_ ^ _3832_ /*92705*/;
assign _3830_ = _3831_ | _3833_ /*92702*/;
assign _3839_ = ~D[50] /*92701*/;
assign _3836_ = _3122_ & _3839_ /*92697*/;
assign _3837_ = _3122_ ^ _3839_ /*92700*/;
assign _3838_ = _3830_ & _3837_ /*92698*/;
assign _3571_ = _3830_ ^ _3837_ /*92699*/;
assign _3835_ = _3836_ | _3838_ /*92696*/;
assign _3844_ = ~D[51] /*92695*/;
assign _3841_ = _3123_ & _3844_ /*92691*/;
assign _3842_ = _3123_ ^ _3844_ /*92694*/;
assign _3843_ = _3835_ & _3842_ /*92692*/;
assign _3572_ = _3835_ ^ _3842_ /*92693*/;
assign _3840_ = _3841_ | _3843_ /*92690*/;
assign _3849_ = ~D[52] /*92689*/;
assign _3846_ = _3124_ & _3849_ /*92685*/;
assign _3847_ = _3124_ ^ _3849_ /*92688*/;
assign _3848_ = _3840_ & _3847_ /*92686*/;
assign _3573_ = _3840_ ^ _3847_ /*92687*/;
assign _3845_ = _3846_ | _3848_ /*92684*/;
assign _3854_ = ~D[53] /*92683*/;
assign _3851_ = _3125_ & _3854_ /*92679*/;
assign _3852_ = _3125_ ^ _3854_ /*92682*/;
assign _3853_ = _3845_ & _3852_ /*92680*/;
assign _3574_ = _3845_ ^ _3852_ /*92681*/;
assign _3850_ = _3851_ | _3853_ /*92678*/;
assign _3859_ = ~D[54] /*92677*/;
assign _3856_ = _3126_ & _3859_ /*92673*/;
assign _3857_ = _3126_ ^ _3859_ /*92676*/;
assign _3858_ = _3850_ & _3857_ /*92674*/;
assign _3575_ = _3850_ ^ _3857_ /*92675*/;
assign _3855_ = _3856_ | _3858_ /*92672*/;
assign _3864_ = ~D[55] /*92671*/;
assign _3861_ = _3127_ & _3864_ /*92667*/;
assign _3862_ = _3127_ ^ _3864_ /*92670*/;
assign _3863_ = _3855_ & _3862_ /*92668*/;
assign _3576_ = _3855_ ^ _3862_ /*92669*/;
assign _3860_ = _3861_ | _3863_ /*92666*/;
assign _3869_ = ~D[56] /*92665*/;
assign _3866_ = _3128_ & _3869_ /*92661*/;
assign _3867_ = _3128_ ^ _3869_ /*92664*/;
assign _3868_ = _3860_ & _3867_ /*92662*/;
assign _3577_ = _3860_ ^ _3867_ /*92663*/;
assign _3865_ = _3866_ | _3868_ /*92660*/;
assign _3874_ = ~D[57] /*92659*/;
assign _3871_ = _3129_ & _3874_ /*92655*/;
assign _3872_ = _3129_ ^ _3874_ /*92658*/;
assign _3873_ = _3865_ & _3872_ /*92656*/;
assign _3578_ = _3865_ ^ _3872_ /*92657*/;
assign _3870_ = _3871_ | _3873_ /*92654*/;
assign _3879_ = ~D[58] /*92653*/;
assign _3876_ = _3130_ & _3879_ /*92649*/;
assign _3877_ = _3130_ ^ _3879_ /*92652*/;
assign _3878_ = _3870_ & _3877_ /*92650*/;
assign _3579_ = _3870_ ^ _3877_ /*92651*/;
assign _3875_ = _3876_ | _3878_ /*92648*/;
assign _3884_ = ~D[59] /*92647*/;
assign _3881_ = _3131_ & _3884_ /*92643*/;
assign _3882_ = _3131_ ^ _3884_ /*92646*/;
assign _3883_ = _3875_ & _3882_ /*92644*/;
assign _3580_ = _3875_ ^ _3882_ /*92645*/;
assign _3880_ = _3881_ | _3883_ /*92642*/;
assign _3889_ = ~D[60] /*92641*/;
assign _3886_ = _3132_ & _3889_ /*92637*/;
assign _3887_ = _3132_ ^ _3889_ /*92640*/;
assign _3888_ = _3880_ & _3887_ /*92638*/;
assign _3581_ = _3880_ ^ _3887_ /*92639*/;
assign _3885_ = _3886_ | _3888_ /*92636*/;
assign _3894_ = ~D[61] /*92635*/;
assign _3891_ = _3133_ & _3894_ /*92631*/;
assign _3892_ = _3133_ ^ _3894_ /*92634*/;
assign _3893_ = _3885_ & _3892_ /*92632*/;
assign _3582_ = _3885_ ^ _3892_ /*92633*/;
assign _3890_ = _3891_ | _3893_ /*92630*/;
assign _3899_ = ~D[62] /*92629*/;
assign _3896_ = _3134_ & _3899_ /*92625*/;
assign _3897_ = _3134_ ^ _3899_ /*92628*/;
assign _3898_ = _3890_ & _3897_ /*92626*/;
assign _3583_ = _3890_ ^ _3897_ /*92627*/;
assign _3895_ = _3896_ | _3898_ /*92624*/;
assign _3900_ = _3135_ & oneWire /*92619*/;
assign _3901_ = _3135_ ^ oneWire /*92622*/;
assign _3902_ = _3895_ & _3901_ /*92620*/;
assign _3584_ = _3895_ ^ _3901_ /*92621*/;
assign Q[59] = _3900_ | _3902_ /*92618*/;
assign _4035_ = ~Q[59] /*92233*/;
assign _4034_ = _4035_ & D[0] /*92232*/;
assign _4037_ = _3521_ & _4034_ /*92227*/;
assign _4038_ = _3521_ ^ _4034_ /*92230*/;
assign _4039_ = zeroWire & _4038_ /*92228*/;
assign _3969_ = zeroWire ^ _4038_ /*92229*/;
assign _4036_ = _4037_ | _4039_ /*92226*/;
assign _4041_ = ~Q[59] /*92225*/;
assign _4040_ = _4041_ & D[1] /*92224*/;
assign _4043_ = _3522_ & _4040_ /*92219*/;
assign _4044_ = _3522_ ^ _4040_ /*92222*/;
assign _4045_ = _4036_ & _4044_ /*92220*/;
assign _3970_ = _4036_ ^ _4044_ /*92221*/;
assign _4042_ = _4043_ | _4045_ /*92218*/;
assign _4047_ = ~Q[59] /*92217*/;
assign _4046_ = _4047_ & D[2] /*92216*/;
assign _4049_ = _3523_ & _4046_ /*92211*/;
assign _4050_ = _3523_ ^ _4046_ /*92214*/;
assign _4051_ = _4042_ & _4050_ /*92212*/;
assign _3971_ = _4042_ ^ _4050_ /*92213*/;
assign _4048_ = _4049_ | _4051_ /*92210*/;
assign _4053_ = ~Q[59] /*92209*/;
assign _4052_ = _4053_ & D[3] /*92208*/;
assign _4055_ = _3524_ & _4052_ /*92203*/;
assign _4056_ = _3524_ ^ _4052_ /*92206*/;
assign _4057_ = _4048_ & _4056_ /*92204*/;
assign _3972_ = _4048_ ^ _4056_ /*92205*/;
assign _4054_ = _4055_ | _4057_ /*92202*/;
assign _4059_ = ~Q[59] /*92201*/;
assign _4058_ = _4059_ & D[4] /*92200*/;
assign _4061_ = _3525_ & _4058_ /*92195*/;
assign _4062_ = _3525_ ^ _4058_ /*92198*/;
assign _4063_ = _4054_ & _4062_ /*92196*/;
assign _3973_ = _4054_ ^ _4062_ /*92197*/;
assign _4060_ = _4061_ | _4063_ /*92194*/;
assign _4065_ = ~Q[59] /*92193*/;
assign _4064_ = _4065_ & D[5] /*92192*/;
assign _4067_ = _3526_ & _4064_ /*92187*/;
assign _4068_ = _3526_ ^ _4064_ /*92190*/;
assign _4069_ = _4060_ & _4068_ /*92188*/;
assign _3974_ = _4060_ ^ _4068_ /*92189*/;
assign _4066_ = _4067_ | _4069_ /*92186*/;
assign _4071_ = ~Q[59] /*92185*/;
assign _4070_ = _4071_ & D[6] /*92184*/;
assign _4073_ = _3527_ & _4070_ /*92179*/;
assign _4074_ = _3527_ ^ _4070_ /*92182*/;
assign _4075_ = _4066_ & _4074_ /*92180*/;
assign _3975_ = _4066_ ^ _4074_ /*92181*/;
assign _4072_ = _4073_ | _4075_ /*92178*/;
assign _4077_ = ~Q[59] /*92177*/;
assign _4076_ = _4077_ & D[7] /*92176*/;
assign _4079_ = _3528_ & _4076_ /*92171*/;
assign _4080_ = _3528_ ^ _4076_ /*92174*/;
assign _4081_ = _4072_ & _4080_ /*92172*/;
assign _3976_ = _4072_ ^ _4080_ /*92173*/;
assign _4078_ = _4079_ | _4081_ /*92170*/;
assign _4083_ = ~Q[59] /*92169*/;
assign _4082_ = _4083_ & D[8] /*92168*/;
assign _4085_ = _3529_ & _4082_ /*92163*/;
assign _4086_ = _3529_ ^ _4082_ /*92166*/;
assign _4087_ = _4078_ & _4086_ /*92164*/;
assign _3977_ = _4078_ ^ _4086_ /*92165*/;
assign _4084_ = _4085_ | _4087_ /*92162*/;
assign _4089_ = ~Q[59] /*92161*/;
assign _4088_ = _4089_ & D[9] /*92160*/;
assign _4091_ = _3530_ & _4088_ /*92155*/;
assign _4092_ = _3530_ ^ _4088_ /*92158*/;
assign _4093_ = _4084_ & _4092_ /*92156*/;
assign _3978_ = _4084_ ^ _4092_ /*92157*/;
assign _4090_ = _4091_ | _4093_ /*92154*/;
assign _4095_ = ~Q[59] /*92153*/;
assign _4094_ = _4095_ & D[10] /*92152*/;
assign _4097_ = _3531_ & _4094_ /*92147*/;
assign _4098_ = _3531_ ^ _4094_ /*92150*/;
assign _4099_ = _4090_ & _4098_ /*92148*/;
assign _3979_ = _4090_ ^ _4098_ /*92149*/;
assign _4096_ = _4097_ | _4099_ /*92146*/;
assign _4101_ = ~Q[59] /*92145*/;
assign _4100_ = _4101_ & D[11] /*92144*/;
assign _4103_ = _3532_ & _4100_ /*92139*/;
assign _4104_ = _3532_ ^ _4100_ /*92142*/;
assign _4105_ = _4096_ & _4104_ /*92140*/;
assign _3980_ = _4096_ ^ _4104_ /*92141*/;
assign _4102_ = _4103_ | _4105_ /*92138*/;
assign _4107_ = ~Q[59] /*92137*/;
assign _4106_ = _4107_ & D[12] /*92136*/;
assign _4109_ = _3533_ & _4106_ /*92131*/;
assign _4110_ = _3533_ ^ _4106_ /*92134*/;
assign _4111_ = _4102_ & _4110_ /*92132*/;
assign _3981_ = _4102_ ^ _4110_ /*92133*/;
assign _4108_ = _4109_ | _4111_ /*92130*/;
assign _4113_ = ~Q[59] /*92129*/;
assign _4112_ = _4113_ & D[13] /*92128*/;
assign _4115_ = _3534_ & _4112_ /*92123*/;
assign _4116_ = _3534_ ^ _4112_ /*92126*/;
assign _4117_ = _4108_ & _4116_ /*92124*/;
assign _3982_ = _4108_ ^ _4116_ /*92125*/;
assign _4114_ = _4115_ | _4117_ /*92122*/;
assign _4119_ = ~Q[59] /*92121*/;
assign _4118_ = _4119_ & D[14] /*92120*/;
assign _4121_ = _3535_ & _4118_ /*92115*/;
assign _4122_ = _3535_ ^ _4118_ /*92118*/;
assign _4123_ = _4114_ & _4122_ /*92116*/;
assign _3983_ = _4114_ ^ _4122_ /*92117*/;
assign _4120_ = _4121_ | _4123_ /*92114*/;
assign _4125_ = ~Q[59] /*92113*/;
assign _4124_ = _4125_ & D[15] /*92112*/;
assign _4127_ = _3536_ & _4124_ /*92107*/;
assign _4128_ = _3536_ ^ _4124_ /*92110*/;
assign _4129_ = _4120_ & _4128_ /*92108*/;
assign _3984_ = _4120_ ^ _4128_ /*92109*/;
assign _4126_ = _4127_ | _4129_ /*92106*/;
assign _4131_ = ~Q[59] /*92105*/;
assign _4130_ = _4131_ & D[16] /*92104*/;
assign _4133_ = _3537_ & _4130_ /*92099*/;
assign _4134_ = _3537_ ^ _4130_ /*92102*/;
assign _4135_ = _4126_ & _4134_ /*92100*/;
assign _3985_ = _4126_ ^ _4134_ /*92101*/;
assign _4132_ = _4133_ | _4135_ /*92098*/;
assign _4137_ = ~Q[59] /*92097*/;
assign _4136_ = _4137_ & D[17] /*92096*/;
assign _4139_ = _3538_ & _4136_ /*92091*/;
assign _4140_ = _3538_ ^ _4136_ /*92094*/;
assign _4141_ = _4132_ & _4140_ /*92092*/;
assign _3986_ = _4132_ ^ _4140_ /*92093*/;
assign _4138_ = _4139_ | _4141_ /*92090*/;
assign _4143_ = ~Q[59] /*92089*/;
assign _4142_ = _4143_ & D[18] /*92088*/;
assign _4145_ = _3539_ & _4142_ /*92083*/;
assign _4146_ = _3539_ ^ _4142_ /*92086*/;
assign _4147_ = _4138_ & _4146_ /*92084*/;
assign _3987_ = _4138_ ^ _4146_ /*92085*/;
assign _4144_ = _4145_ | _4147_ /*92082*/;
assign _4149_ = ~Q[59] /*92081*/;
assign _4148_ = _4149_ & D[19] /*92080*/;
assign _4151_ = _3540_ & _4148_ /*92075*/;
assign _4152_ = _3540_ ^ _4148_ /*92078*/;
assign _4153_ = _4144_ & _4152_ /*92076*/;
assign _3988_ = _4144_ ^ _4152_ /*92077*/;
assign _4150_ = _4151_ | _4153_ /*92074*/;
assign _4155_ = ~Q[59] /*92073*/;
assign _4154_ = _4155_ & D[20] /*92072*/;
assign _4157_ = _3541_ & _4154_ /*92067*/;
assign _4158_ = _3541_ ^ _4154_ /*92070*/;
assign _4159_ = _4150_ & _4158_ /*92068*/;
assign _3989_ = _4150_ ^ _4158_ /*92069*/;
assign _4156_ = _4157_ | _4159_ /*92066*/;
assign _4161_ = ~Q[59] /*92065*/;
assign _4160_ = _4161_ & D[21] /*92064*/;
assign _4163_ = _3542_ & _4160_ /*92059*/;
assign _4164_ = _3542_ ^ _4160_ /*92062*/;
assign _4165_ = _4156_ & _4164_ /*92060*/;
assign _3990_ = _4156_ ^ _4164_ /*92061*/;
assign _4162_ = _4163_ | _4165_ /*92058*/;
assign _4167_ = ~Q[59] /*92057*/;
assign _4166_ = _4167_ & D[22] /*92056*/;
assign _4169_ = _3543_ & _4166_ /*92051*/;
assign _4170_ = _3543_ ^ _4166_ /*92054*/;
assign _4171_ = _4162_ & _4170_ /*92052*/;
assign _3991_ = _4162_ ^ _4170_ /*92053*/;
assign _4168_ = _4169_ | _4171_ /*92050*/;
assign _4173_ = ~Q[59] /*92049*/;
assign _4172_ = _4173_ & D[23] /*92048*/;
assign _4175_ = _3544_ & _4172_ /*92043*/;
assign _4176_ = _3544_ ^ _4172_ /*92046*/;
assign _4177_ = _4168_ & _4176_ /*92044*/;
assign _3992_ = _4168_ ^ _4176_ /*92045*/;
assign _4174_ = _4175_ | _4177_ /*92042*/;
assign _4179_ = ~Q[59] /*92041*/;
assign _4178_ = _4179_ & D[24] /*92040*/;
assign _4181_ = _3545_ & _4178_ /*92035*/;
assign _4182_ = _3545_ ^ _4178_ /*92038*/;
assign _4183_ = _4174_ & _4182_ /*92036*/;
assign _3993_ = _4174_ ^ _4182_ /*92037*/;
assign _4180_ = _4181_ | _4183_ /*92034*/;
assign _4185_ = ~Q[59] /*92033*/;
assign _4184_ = _4185_ & D[25] /*92032*/;
assign _4187_ = _3546_ & _4184_ /*92027*/;
assign _4188_ = _3546_ ^ _4184_ /*92030*/;
assign _4189_ = _4180_ & _4188_ /*92028*/;
assign _3994_ = _4180_ ^ _4188_ /*92029*/;
assign _4186_ = _4187_ | _4189_ /*92026*/;
assign _4191_ = ~Q[59] /*92025*/;
assign _4190_ = _4191_ & D[26] /*92024*/;
assign _4193_ = _3547_ & _4190_ /*92019*/;
assign _4194_ = _3547_ ^ _4190_ /*92022*/;
assign _4195_ = _4186_ & _4194_ /*92020*/;
assign _3995_ = _4186_ ^ _4194_ /*92021*/;
assign _4192_ = _4193_ | _4195_ /*92018*/;
assign _4197_ = ~Q[59] /*92017*/;
assign _4196_ = _4197_ & D[27] /*92016*/;
assign _4199_ = _3548_ & _4196_ /*92011*/;
assign _4200_ = _3548_ ^ _4196_ /*92014*/;
assign _4201_ = _4192_ & _4200_ /*92012*/;
assign _3996_ = _4192_ ^ _4200_ /*92013*/;
assign _4198_ = _4199_ | _4201_ /*92010*/;
assign _4203_ = ~Q[59] /*92009*/;
assign _4202_ = _4203_ & D[28] /*92008*/;
assign _4205_ = _3549_ & _4202_ /*92003*/;
assign _4206_ = _3549_ ^ _4202_ /*92006*/;
assign _4207_ = _4198_ & _4206_ /*92004*/;
assign _3997_ = _4198_ ^ _4206_ /*92005*/;
assign _4204_ = _4205_ | _4207_ /*92002*/;
assign _4209_ = ~Q[59] /*92001*/;
assign _4208_ = _4209_ & D[29] /*92000*/;
assign _4211_ = _3550_ & _4208_ /*91995*/;
assign _4212_ = _3550_ ^ _4208_ /*91998*/;
assign _4213_ = _4204_ & _4212_ /*91996*/;
assign _3998_ = _4204_ ^ _4212_ /*91997*/;
assign _4210_ = _4211_ | _4213_ /*91994*/;
assign _4215_ = ~Q[59] /*91993*/;
assign _4214_ = _4215_ & D[30] /*91992*/;
assign _4217_ = _3551_ & _4214_ /*91987*/;
assign _4218_ = _3551_ ^ _4214_ /*91990*/;
assign _4219_ = _4210_ & _4218_ /*91988*/;
assign _3999_ = _4210_ ^ _4218_ /*91989*/;
assign _4216_ = _4217_ | _4219_ /*91986*/;
assign _4221_ = ~Q[59] /*91985*/;
assign _4220_ = _4221_ & D[31] /*91984*/;
assign _4223_ = _3552_ & _4220_ /*91979*/;
assign _4224_ = _3552_ ^ _4220_ /*91982*/;
assign _4225_ = _4216_ & _4224_ /*91980*/;
assign _4000_ = _4216_ ^ _4224_ /*91981*/;
assign _4222_ = _4223_ | _4225_ /*91978*/;
assign _4227_ = ~Q[59] /*91977*/;
assign _4226_ = _4227_ & D[32] /*91976*/;
assign _4229_ = _3553_ & _4226_ /*91971*/;
assign _4230_ = _3553_ ^ _4226_ /*91974*/;
assign _4231_ = _4222_ & _4230_ /*91972*/;
assign _4001_ = _4222_ ^ _4230_ /*91973*/;
assign _4228_ = _4229_ | _4231_ /*91970*/;
assign _4233_ = ~Q[59] /*91969*/;
assign _4232_ = _4233_ & D[33] /*91968*/;
assign _4235_ = _3554_ & _4232_ /*91963*/;
assign _4236_ = _3554_ ^ _4232_ /*91966*/;
assign _4237_ = _4228_ & _4236_ /*91964*/;
assign _4002_ = _4228_ ^ _4236_ /*91965*/;
assign _4234_ = _4235_ | _4237_ /*91962*/;
assign _4239_ = ~Q[59] /*91961*/;
assign _4238_ = _4239_ & D[34] /*91960*/;
assign _4241_ = _3555_ & _4238_ /*91955*/;
assign _4242_ = _3555_ ^ _4238_ /*91958*/;
assign _4243_ = _4234_ & _4242_ /*91956*/;
assign _4003_ = _4234_ ^ _4242_ /*91957*/;
assign _4240_ = _4241_ | _4243_ /*91954*/;
assign _4245_ = ~Q[59] /*91953*/;
assign _4244_ = _4245_ & D[35] /*91952*/;
assign _4247_ = _3556_ & _4244_ /*91947*/;
assign _4248_ = _3556_ ^ _4244_ /*91950*/;
assign _4249_ = _4240_ & _4248_ /*91948*/;
assign _4004_ = _4240_ ^ _4248_ /*91949*/;
assign _4246_ = _4247_ | _4249_ /*91946*/;
assign _4251_ = ~Q[59] /*91945*/;
assign _4250_ = _4251_ & D[36] /*91944*/;
assign _4253_ = _3557_ & _4250_ /*91939*/;
assign _4254_ = _3557_ ^ _4250_ /*91942*/;
assign _4255_ = _4246_ & _4254_ /*91940*/;
assign _4005_ = _4246_ ^ _4254_ /*91941*/;
assign _4252_ = _4253_ | _4255_ /*91938*/;
assign _4257_ = ~Q[59] /*91937*/;
assign _4256_ = _4257_ & D[37] /*91936*/;
assign _4259_ = _3558_ & _4256_ /*91931*/;
assign _4260_ = _3558_ ^ _4256_ /*91934*/;
assign _4261_ = _4252_ & _4260_ /*91932*/;
assign _4006_ = _4252_ ^ _4260_ /*91933*/;
assign _4258_ = _4259_ | _4261_ /*91930*/;
assign _4263_ = ~Q[59] /*91929*/;
assign _4262_ = _4263_ & D[38] /*91928*/;
assign _4265_ = _3559_ & _4262_ /*91923*/;
assign _4266_ = _3559_ ^ _4262_ /*91926*/;
assign _4267_ = _4258_ & _4266_ /*91924*/;
assign _4007_ = _4258_ ^ _4266_ /*91925*/;
assign _4264_ = _4265_ | _4267_ /*91922*/;
assign _4269_ = ~Q[59] /*91921*/;
assign _4268_ = _4269_ & D[39] /*91920*/;
assign _4271_ = _3560_ & _4268_ /*91915*/;
assign _4272_ = _3560_ ^ _4268_ /*91918*/;
assign _4273_ = _4264_ & _4272_ /*91916*/;
assign _4008_ = _4264_ ^ _4272_ /*91917*/;
assign _4270_ = _4271_ | _4273_ /*91914*/;
assign _4275_ = ~Q[59] /*91913*/;
assign _4274_ = _4275_ & D[40] /*91912*/;
assign _4277_ = _3561_ & _4274_ /*91907*/;
assign _4278_ = _3561_ ^ _4274_ /*91910*/;
assign _4279_ = _4270_ & _4278_ /*91908*/;
assign _4009_ = _4270_ ^ _4278_ /*91909*/;
assign _4276_ = _4277_ | _4279_ /*91906*/;
assign _4281_ = ~Q[59] /*91905*/;
assign _4280_ = _4281_ & D[41] /*91904*/;
assign _4283_ = _3562_ & _4280_ /*91899*/;
assign _4284_ = _3562_ ^ _4280_ /*91902*/;
assign _4285_ = _4276_ & _4284_ /*91900*/;
assign _4010_ = _4276_ ^ _4284_ /*91901*/;
assign _4282_ = _4283_ | _4285_ /*91898*/;
assign _4287_ = ~Q[59] /*91897*/;
assign _4286_ = _4287_ & D[42] /*91896*/;
assign _4289_ = _3563_ & _4286_ /*91891*/;
assign _4290_ = _3563_ ^ _4286_ /*91894*/;
assign _4291_ = _4282_ & _4290_ /*91892*/;
assign _4011_ = _4282_ ^ _4290_ /*91893*/;
assign _4288_ = _4289_ | _4291_ /*91890*/;
assign _4293_ = ~Q[59] /*91889*/;
assign _4292_ = _4293_ & D[43] /*91888*/;
assign _4295_ = _3564_ & _4292_ /*91883*/;
assign _4296_ = _3564_ ^ _4292_ /*91886*/;
assign _4297_ = _4288_ & _4296_ /*91884*/;
assign _4012_ = _4288_ ^ _4296_ /*91885*/;
assign _4294_ = _4295_ | _4297_ /*91882*/;
assign _4299_ = ~Q[59] /*91881*/;
assign _4298_ = _4299_ & D[44] /*91880*/;
assign _4301_ = _3565_ & _4298_ /*91875*/;
assign _4302_ = _3565_ ^ _4298_ /*91878*/;
assign _4303_ = _4294_ & _4302_ /*91876*/;
assign _4013_ = _4294_ ^ _4302_ /*91877*/;
assign _4300_ = _4301_ | _4303_ /*91874*/;
assign _4305_ = ~Q[59] /*91873*/;
assign _4304_ = _4305_ & D[45] /*91872*/;
assign _4307_ = _3566_ & _4304_ /*91867*/;
assign _4308_ = _3566_ ^ _4304_ /*91870*/;
assign _4309_ = _4300_ & _4308_ /*91868*/;
assign _4014_ = _4300_ ^ _4308_ /*91869*/;
assign _4306_ = _4307_ | _4309_ /*91866*/;
assign _4311_ = ~Q[59] /*91865*/;
assign _4310_ = _4311_ & D[46] /*91864*/;
assign _4313_ = _3567_ & _4310_ /*91859*/;
assign _4314_ = _3567_ ^ _4310_ /*91862*/;
assign _4315_ = _4306_ & _4314_ /*91860*/;
assign _4015_ = _4306_ ^ _4314_ /*91861*/;
assign _4312_ = _4313_ | _4315_ /*91858*/;
assign _4317_ = ~Q[59] /*91857*/;
assign _4316_ = _4317_ & D[47] /*91856*/;
assign _4319_ = _3568_ & _4316_ /*91851*/;
assign _4320_ = _3568_ ^ _4316_ /*91854*/;
assign _4321_ = _4312_ & _4320_ /*91852*/;
assign _4016_ = _4312_ ^ _4320_ /*91853*/;
assign _4318_ = _4319_ | _4321_ /*91850*/;
assign _4323_ = ~Q[59] /*91849*/;
assign _4322_ = _4323_ & D[48] /*91848*/;
assign _4325_ = _3569_ & _4322_ /*91843*/;
assign _4326_ = _3569_ ^ _4322_ /*91846*/;
assign _4327_ = _4318_ & _4326_ /*91844*/;
assign _4017_ = _4318_ ^ _4326_ /*91845*/;
assign _4324_ = _4325_ | _4327_ /*91842*/;
assign _4329_ = ~Q[59] /*91841*/;
assign _4328_ = _4329_ & D[49] /*91840*/;
assign _4331_ = _3570_ & _4328_ /*91835*/;
assign _4332_ = _3570_ ^ _4328_ /*91838*/;
assign _4333_ = _4324_ & _4332_ /*91836*/;
assign _4018_ = _4324_ ^ _4332_ /*91837*/;
assign _4330_ = _4331_ | _4333_ /*91834*/;
assign _4335_ = ~Q[59] /*91833*/;
assign _4334_ = _4335_ & D[50] /*91832*/;
assign _4337_ = _3571_ & _4334_ /*91827*/;
assign _4338_ = _3571_ ^ _4334_ /*91830*/;
assign _4339_ = _4330_ & _4338_ /*91828*/;
assign _4019_ = _4330_ ^ _4338_ /*91829*/;
assign _4336_ = _4337_ | _4339_ /*91826*/;
assign _4341_ = ~Q[59] /*91825*/;
assign _4340_ = _4341_ & D[51] /*91824*/;
assign _4343_ = _3572_ & _4340_ /*91819*/;
assign _4344_ = _3572_ ^ _4340_ /*91822*/;
assign _4345_ = _4336_ & _4344_ /*91820*/;
assign _4020_ = _4336_ ^ _4344_ /*91821*/;
assign _4342_ = _4343_ | _4345_ /*91818*/;
assign _4347_ = ~Q[59] /*91817*/;
assign _4346_ = _4347_ & D[52] /*91816*/;
assign _4349_ = _3573_ & _4346_ /*91811*/;
assign _4350_ = _3573_ ^ _4346_ /*91814*/;
assign _4351_ = _4342_ & _4350_ /*91812*/;
assign _4021_ = _4342_ ^ _4350_ /*91813*/;
assign _4348_ = _4349_ | _4351_ /*91810*/;
assign _4353_ = ~Q[59] /*91809*/;
assign _4352_ = _4353_ & D[53] /*91808*/;
assign _4355_ = _3574_ & _4352_ /*91803*/;
assign _4356_ = _3574_ ^ _4352_ /*91806*/;
assign _4357_ = _4348_ & _4356_ /*91804*/;
assign _4022_ = _4348_ ^ _4356_ /*91805*/;
assign _4354_ = _4355_ | _4357_ /*91802*/;
assign _4359_ = ~Q[59] /*91801*/;
assign _4358_ = _4359_ & D[54] /*91800*/;
assign _4361_ = _3575_ & _4358_ /*91795*/;
assign _4362_ = _3575_ ^ _4358_ /*91798*/;
assign _4363_ = _4354_ & _4362_ /*91796*/;
assign _4023_ = _4354_ ^ _4362_ /*91797*/;
assign _4360_ = _4361_ | _4363_ /*91794*/;
assign _4365_ = ~Q[59] /*91793*/;
assign _4364_ = _4365_ & D[55] /*91792*/;
assign _4367_ = _3576_ & _4364_ /*91787*/;
assign _4368_ = _3576_ ^ _4364_ /*91790*/;
assign _4369_ = _4360_ & _4368_ /*91788*/;
assign _4024_ = _4360_ ^ _4368_ /*91789*/;
assign _4366_ = _4367_ | _4369_ /*91786*/;
assign _4371_ = ~Q[59] /*91785*/;
assign _4370_ = _4371_ & D[56] /*91784*/;
assign _4373_ = _3577_ & _4370_ /*91779*/;
assign _4374_ = _3577_ ^ _4370_ /*91782*/;
assign _4375_ = _4366_ & _4374_ /*91780*/;
assign _4025_ = _4366_ ^ _4374_ /*91781*/;
assign _4372_ = _4373_ | _4375_ /*91778*/;
assign _4377_ = ~Q[59] /*91777*/;
assign _4376_ = _4377_ & D[57] /*91776*/;
assign _4379_ = _3578_ & _4376_ /*91771*/;
assign _4380_ = _3578_ ^ _4376_ /*91774*/;
assign _4381_ = _4372_ & _4380_ /*91772*/;
assign _4026_ = _4372_ ^ _4380_ /*91773*/;
assign _4378_ = _4379_ | _4381_ /*91770*/;
assign _4383_ = ~Q[59] /*91769*/;
assign _4382_ = _4383_ & D[58] /*91768*/;
assign _4385_ = _3579_ & _4382_ /*91763*/;
assign _4386_ = _3579_ ^ _4382_ /*91766*/;
assign _4387_ = _4378_ & _4386_ /*91764*/;
assign _4027_ = _4378_ ^ _4386_ /*91765*/;
assign _4384_ = _4385_ | _4387_ /*91762*/;
assign _4389_ = ~Q[59] /*91761*/;
assign _4388_ = _4389_ & D[59] /*91760*/;
assign _4391_ = _3580_ & _4388_ /*91755*/;
assign _4392_ = _3580_ ^ _4388_ /*91758*/;
assign _4393_ = _4384_ & _4392_ /*91756*/;
assign _4028_ = _4384_ ^ _4392_ /*91757*/;
assign _4390_ = _4391_ | _4393_ /*91754*/;
assign _4395_ = ~Q[59] /*91753*/;
assign _4394_ = _4395_ & D[60] /*91752*/;
assign _4397_ = _3581_ & _4394_ /*91747*/;
assign _4398_ = _3581_ ^ _4394_ /*91750*/;
assign _4399_ = _4390_ & _4398_ /*91748*/;
assign _4029_ = _4390_ ^ _4398_ /*91749*/;
assign _4396_ = _4397_ | _4399_ /*91746*/;
assign _4401_ = ~Q[59] /*91745*/;
assign _4400_ = _4401_ & D[61] /*91744*/;
assign _4403_ = _3582_ & _4400_ /*91739*/;
assign _4404_ = _3582_ ^ _4400_ /*91742*/;
assign _4405_ = _4396_ & _4404_ /*91740*/;
assign _4030_ = _4396_ ^ _4404_ /*91741*/;
assign _4402_ = _4403_ | _4405_ /*91738*/;
assign _4407_ = ~Q[59] /*91737*/;
assign _4406_ = _4407_ & D[62] /*91736*/;
assign _4409_ = _3583_ & _4406_ /*91731*/;
assign _4410_ = _3583_ ^ _4406_ /*91734*/;
assign _4411_ = _4402_ & _4410_ /*91732*/;
assign _4031_ = _4402_ ^ _4410_ /*91733*/;
assign _4408_ = _4409_ | _4411_ /*91730*/;
assign _4413_ = ~Q[59] /*91729*/;
assign _4412_ = _4413_ & zeroWire /*91728*/;
assign _4414_ = _3584_ ^ _4412_ /*91726*/;
assign _4032_ = _4414_ ^ _4408_ /*91725*/;
assign _4485_ = ~D[0] /*91471*/;
assign _4482_ = R_0[58] & _4485_ /*91467*/;
assign _4483_ = R_0[58] ^ _4485_ /*91470*/;
assign _4484_ = oneWire & _4483_ /*91468*/;
assign _4417_ = oneWire ^ _4483_ /*91469*/;
assign _4481_ = _4482_ | _4484_ /*91466*/;
assign _4490_ = ~D[1] /*91465*/;
assign _4487_ = _3969_ & _4490_ /*91461*/;
assign _4488_ = _3969_ ^ _4490_ /*91464*/;
assign _4489_ = _4481_ & _4488_ /*91462*/;
assign _4418_ = _4481_ ^ _4488_ /*91463*/;
assign _4486_ = _4487_ | _4489_ /*91460*/;
assign _4495_ = ~D[2] /*91459*/;
assign _4492_ = _3970_ & _4495_ /*91455*/;
assign _4493_ = _3970_ ^ _4495_ /*91458*/;
assign _4494_ = _4486_ & _4493_ /*91456*/;
assign _4419_ = _4486_ ^ _4493_ /*91457*/;
assign _4491_ = _4492_ | _4494_ /*91454*/;
assign _4500_ = ~D[3] /*91453*/;
assign _4497_ = _3971_ & _4500_ /*91449*/;
assign _4498_ = _3971_ ^ _4500_ /*91452*/;
assign _4499_ = _4491_ & _4498_ /*91450*/;
assign _4420_ = _4491_ ^ _4498_ /*91451*/;
assign _4496_ = _4497_ | _4499_ /*91448*/;
assign _4505_ = ~D[4] /*91447*/;
assign _4502_ = _3972_ & _4505_ /*91443*/;
assign _4503_ = _3972_ ^ _4505_ /*91446*/;
assign _4504_ = _4496_ & _4503_ /*91444*/;
assign _4421_ = _4496_ ^ _4503_ /*91445*/;
assign _4501_ = _4502_ | _4504_ /*91442*/;
assign _4510_ = ~D[5] /*91441*/;
assign _4507_ = _3973_ & _4510_ /*91437*/;
assign _4508_ = _3973_ ^ _4510_ /*91440*/;
assign _4509_ = _4501_ & _4508_ /*91438*/;
assign _4422_ = _4501_ ^ _4508_ /*91439*/;
assign _4506_ = _4507_ | _4509_ /*91436*/;
assign _4515_ = ~D[6] /*91435*/;
assign _4512_ = _3974_ & _4515_ /*91431*/;
assign _4513_ = _3974_ ^ _4515_ /*91434*/;
assign _4514_ = _4506_ & _4513_ /*91432*/;
assign _4423_ = _4506_ ^ _4513_ /*91433*/;
assign _4511_ = _4512_ | _4514_ /*91430*/;
assign _4520_ = ~D[7] /*91429*/;
assign _4517_ = _3975_ & _4520_ /*91425*/;
assign _4518_ = _3975_ ^ _4520_ /*91428*/;
assign _4519_ = _4511_ & _4518_ /*91426*/;
assign _4424_ = _4511_ ^ _4518_ /*91427*/;
assign _4516_ = _4517_ | _4519_ /*91424*/;
assign _4525_ = ~D[8] /*91423*/;
assign _4522_ = _3976_ & _4525_ /*91419*/;
assign _4523_ = _3976_ ^ _4525_ /*91422*/;
assign _4524_ = _4516_ & _4523_ /*91420*/;
assign _4425_ = _4516_ ^ _4523_ /*91421*/;
assign _4521_ = _4522_ | _4524_ /*91418*/;
assign _4530_ = ~D[9] /*91417*/;
assign _4527_ = _3977_ & _4530_ /*91413*/;
assign _4528_ = _3977_ ^ _4530_ /*91416*/;
assign _4529_ = _4521_ & _4528_ /*91414*/;
assign _4426_ = _4521_ ^ _4528_ /*91415*/;
assign _4526_ = _4527_ | _4529_ /*91412*/;
assign _4535_ = ~D[10] /*91411*/;
assign _4532_ = _3978_ & _4535_ /*91407*/;
assign _4533_ = _3978_ ^ _4535_ /*91410*/;
assign _4534_ = _4526_ & _4533_ /*91408*/;
assign _4427_ = _4526_ ^ _4533_ /*91409*/;
assign _4531_ = _4532_ | _4534_ /*91406*/;
assign _4540_ = ~D[11] /*91405*/;
assign _4537_ = _3979_ & _4540_ /*91401*/;
assign _4538_ = _3979_ ^ _4540_ /*91404*/;
assign _4539_ = _4531_ & _4538_ /*91402*/;
assign _4428_ = _4531_ ^ _4538_ /*91403*/;
assign _4536_ = _4537_ | _4539_ /*91400*/;
assign _4545_ = ~D[12] /*91399*/;
assign _4542_ = _3980_ & _4545_ /*91395*/;
assign _4543_ = _3980_ ^ _4545_ /*91398*/;
assign _4544_ = _4536_ & _4543_ /*91396*/;
assign _4429_ = _4536_ ^ _4543_ /*91397*/;
assign _4541_ = _4542_ | _4544_ /*91394*/;
assign _4550_ = ~D[13] /*91393*/;
assign _4547_ = _3981_ & _4550_ /*91389*/;
assign _4548_ = _3981_ ^ _4550_ /*91392*/;
assign _4549_ = _4541_ & _4548_ /*91390*/;
assign _4430_ = _4541_ ^ _4548_ /*91391*/;
assign _4546_ = _4547_ | _4549_ /*91388*/;
assign _4555_ = ~D[14] /*91387*/;
assign _4552_ = _3982_ & _4555_ /*91383*/;
assign _4553_ = _3982_ ^ _4555_ /*91386*/;
assign _4554_ = _4546_ & _4553_ /*91384*/;
assign _4431_ = _4546_ ^ _4553_ /*91385*/;
assign _4551_ = _4552_ | _4554_ /*91382*/;
assign _4560_ = ~D[15] /*91381*/;
assign _4557_ = _3983_ & _4560_ /*91377*/;
assign _4558_ = _3983_ ^ _4560_ /*91380*/;
assign _4559_ = _4551_ & _4558_ /*91378*/;
assign _4432_ = _4551_ ^ _4558_ /*91379*/;
assign _4556_ = _4557_ | _4559_ /*91376*/;
assign _4565_ = ~D[16] /*91375*/;
assign _4562_ = _3984_ & _4565_ /*91371*/;
assign _4563_ = _3984_ ^ _4565_ /*91374*/;
assign _4564_ = _4556_ & _4563_ /*91372*/;
assign _4433_ = _4556_ ^ _4563_ /*91373*/;
assign _4561_ = _4562_ | _4564_ /*91370*/;
assign _4570_ = ~D[17] /*91369*/;
assign _4567_ = _3985_ & _4570_ /*91365*/;
assign _4568_ = _3985_ ^ _4570_ /*91368*/;
assign _4569_ = _4561_ & _4568_ /*91366*/;
assign _4434_ = _4561_ ^ _4568_ /*91367*/;
assign _4566_ = _4567_ | _4569_ /*91364*/;
assign _4575_ = ~D[18] /*91363*/;
assign _4572_ = _3986_ & _4575_ /*91359*/;
assign _4573_ = _3986_ ^ _4575_ /*91362*/;
assign _4574_ = _4566_ & _4573_ /*91360*/;
assign _4435_ = _4566_ ^ _4573_ /*91361*/;
assign _4571_ = _4572_ | _4574_ /*91358*/;
assign _4580_ = ~D[19] /*91357*/;
assign _4577_ = _3987_ & _4580_ /*91353*/;
assign _4578_ = _3987_ ^ _4580_ /*91356*/;
assign _4579_ = _4571_ & _4578_ /*91354*/;
assign _4436_ = _4571_ ^ _4578_ /*91355*/;
assign _4576_ = _4577_ | _4579_ /*91352*/;
assign _4585_ = ~D[20] /*91351*/;
assign _4582_ = _3988_ & _4585_ /*91347*/;
assign _4583_ = _3988_ ^ _4585_ /*91350*/;
assign _4584_ = _4576_ & _4583_ /*91348*/;
assign _4437_ = _4576_ ^ _4583_ /*91349*/;
assign _4581_ = _4582_ | _4584_ /*91346*/;
assign _4590_ = ~D[21] /*91345*/;
assign _4587_ = _3989_ & _4590_ /*91341*/;
assign _4588_ = _3989_ ^ _4590_ /*91344*/;
assign _4589_ = _4581_ & _4588_ /*91342*/;
assign _4438_ = _4581_ ^ _4588_ /*91343*/;
assign _4586_ = _4587_ | _4589_ /*91340*/;
assign _4595_ = ~D[22] /*91339*/;
assign _4592_ = _3990_ & _4595_ /*91335*/;
assign _4593_ = _3990_ ^ _4595_ /*91338*/;
assign _4594_ = _4586_ & _4593_ /*91336*/;
assign _4439_ = _4586_ ^ _4593_ /*91337*/;
assign _4591_ = _4592_ | _4594_ /*91334*/;
assign _4600_ = ~D[23] /*91333*/;
assign _4597_ = _3991_ & _4600_ /*91329*/;
assign _4598_ = _3991_ ^ _4600_ /*91332*/;
assign _4599_ = _4591_ & _4598_ /*91330*/;
assign _4440_ = _4591_ ^ _4598_ /*91331*/;
assign _4596_ = _4597_ | _4599_ /*91328*/;
assign _4605_ = ~D[24] /*91327*/;
assign _4602_ = _3992_ & _4605_ /*91323*/;
assign _4603_ = _3992_ ^ _4605_ /*91326*/;
assign _4604_ = _4596_ & _4603_ /*91324*/;
assign _4441_ = _4596_ ^ _4603_ /*91325*/;
assign _4601_ = _4602_ | _4604_ /*91322*/;
assign _4610_ = ~D[25] /*91321*/;
assign _4607_ = _3993_ & _4610_ /*91317*/;
assign _4608_ = _3993_ ^ _4610_ /*91320*/;
assign _4609_ = _4601_ & _4608_ /*91318*/;
assign _4442_ = _4601_ ^ _4608_ /*91319*/;
assign _4606_ = _4607_ | _4609_ /*91316*/;
assign _4615_ = ~D[26] /*91315*/;
assign _4612_ = _3994_ & _4615_ /*91311*/;
assign _4613_ = _3994_ ^ _4615_ /*91314*/;
assign _4614_ = _4606_ & _4613_ /*91312*/;
assign _4443_ = _4606_ ^ _4613_ /*91313*/;
assign _4611_ = _4612_ | _4614_ /*91310*/;
assign _4620_ = ~D[27] /*91309*/;
assign _4617_ = _3995_ & _4620_ /*91305*/;
assign _4618_ = _3995_ ^ _4620_ /*91308*/;
assign _4619_ = _4611_ & _4618_ /*91306*/;
assign _4444_ = _4611_ ^ _4618_ /*91307*/;
assign _4616_ = _4617_ | _4619_ /*91304*/;
assign _4625_ = ~D[28] /*91303*/;
assign _4622_ = _3996_ & _4625_ /*91299*/;
assign _4623_ = _3996_ ^ _4625_ /*91302*/;
assign _4624_ = _4616_ & _4623_ /*91300*/;
assign _4445_ = _4616_ ^ _4623_ /*91301*/;
assign _4621_ = _4622_ | _4624_ /*91298*/;
assign _4630_ = ~D[29] /*91297*/;
assign _4627_ = _3997_ & _4630_ /*91293*/;
assign _4628_ = _3997_ ^ _4630_ /*91296*/;
assign _4629_ = _4621_ & _4628_ /*91294*/;
assign _4446_ = _4621_ ^ _4628_ /*91295*/;
assign _4626_ = _4627_ | _4629_ /*91292*/;
assign _4635_ = ~D[30] /*91291*/;
assign _4632_ = _3998_ & _4635_ /*91287*/;
assign _4633_ = _3998_ ^ _4635_ /*91290*/;
assign _4634_ = _4626_ & _4633_ /*91288*/;
assign _4447_ = _4626_ ^ _4633_ /*91289*/;
assign _4631_ = _4632_ | _4634_ /*91286*/;
assign _4640_ = ~D[31] /*91285*/;
assign _4637_ = _3999_ & _4640_ /*91281*/;
assign _4638_ = _3999_ ^ _4640_ /*91284*/;
assign _4639_ = _4631_ & _4638_ /*91282*/;
assign _4448_ = _4631_ ^ _4638_ /*91283*/;
assign _4636_ = _4637_ | _4639_ /*91280*/;
assign _4645_ = ~D[32] /*91279*/;
assign _4642_ = _4000_ & _4645_ /*91275*/;
assign _4643_ = _4000_ ^ _4645_ /*91278*/;
assign _4644_ = _4636_ & _4643_ /*91276*/;
assign _4449_ = _4636_ ^ _4643_ /*91277*/;
assign _4641_ = _4642_ | _4644_ /*91274*/;
assign _4650_ = ~D[33] /*91273*/;
assign _4647_ = _4001_ & _4650_ /*91269*/;
assign _4648_ = _4001_ ^ _4650_ /*91272*/;
assign _4649_ = _4641_ & _4648_ /*91270*/;
assign _4450_ = _4641_ ^ _4648_ /*91271*/;
assign _4646_ = _4647_ | _4649_ /*91268*/;
assign _4655_ = ~D[34] /*91267*/;
assign _4652_ = _4002_ & _4655_ /*91263*/;
assign _4653_ = _4002_ ^ _4655_ /*91266*/;
assign _4654_ = _4646_ & _4653_ /*91264*/;
assign _4451_ = _4646_ ^ _4653_ /*91265*/;
assign _4651_ = _4652_ | _4654_ /*91262*/;
assign _4660_ = ~D[35] /*91261*/;
assign _4657_ = _4003_ & _4660_ /*91257*/;
assign _4658_ = _4003_ ^ _4660_ /*91260*/;
assign _4659_ = _4651_ & _4658_ /*91258*/;
assign _4452_ = _4651_ ^ _4658_ /*91259*/;
assign _4656_ = _4657_ | _4659_ /*91256*/;
assign _4665_ = ~D[36] /*91255*/;
assign _4662_ = _4004_ & _4665_ /*91251*/;
assign _4663_ = _4004_ ^ _4665_ /*91254*/;
assign _4664_ = _4656_ & _4663_ /*91252*/;
assign _4453_ = _4656_ ^ _4663_ /*91253*/;
assign _4661_ = _4662_ | _4664_ /*91250*/;
assign _4670_ = ~D[37] /*91249*/;
assign _4667_ = _4005_ & _4670_ /*91245*/;
assign _4668_ = _4005_ ^ _4670_ /*91248*/;
assign _4669_ = _4661_ & _4668_ /*91246*/;
assign _4454_ = _4661_ ^ _4668_ /*91247*/;
assign _4666_ = _4667_ | _4669_ /*91244*/;
assign _4675_ = ~D[38] /*91243*/;
assign _4672_ = _4006_ & _4675_ /*91239*/;
assign _4673_ = _4006_ ^ _4675_ /*91242*/;
assign _4674_ = _4666_ & _4673_ /*91240*/;
assign _4455_ = _4666_ ^ _4673_ /*91241*/;
assign _4671_ = _4672_ | _4674_ /*91238*/;
assign _4680_ = ~D[39] /*91237*/;
assign _4677_ = _4007_ & _4680_ /*91233*/;
assign _4678_ = _4007_ ^ _4680_ /*91236*/;
assign _4679_ = _4671_ & _4678_ /*91234*/;
assign _4456_ = _4671_ ^ _4678_ /*91235*/;
assign _4676_ = _4677_ | _4679_ /*91232*/;
assign _4685_ = ~D[40] /*91231*/;
assign _4682_ = _4008_ & _4685_ /*91227*/;
assign _4683_ = _4008_ ^ _4685_ /*91230*/;
assign _4684_ = _4676_ & _4683_ /*91228*/;
assign _4457_ = _4676_ ^ _4683_ /*91229*/;
assign _4681_ = _4682_ | _4684_ /*91226*/;
assign _4690_ = ~D[41] /*91225*/;
assign _4687_ = _4009_ & _4690_ /*91221*/;
assign _4688_ = _4009_ ^ _4690_ /*91224*/;
assign _4689_ = _4681_ & _4688_ /*91222*/;
assign _4458_ = _4681_ ^ _4688_ /*91223*/;
assign _4686_ = _4687_ | _4689_ /*91220*/;
assign _4695_ = ~D[42] /*91219*/;
assign _4692_ = _4010_ & _4695_ /*91215*/;
assign _4693_ = _4010_ ^ _4695_ /*91218*/;
assign _4694_ = _4686_ & _4693_ /*91216*/;
assign _4459_ = _4686_ ^ _4693_ /*91217*/;
assign _4691_ = _4692_ | _4694_ /*91214*/;
assign _4700_ = ~D[43] /*91213*/;
assign _4697_ = _4011_ & _4700_ /*91209*/;
assign _4698_ = _4011_ ^ _4700_ /*91212*/;
assign _4699_ = _4691_ & _4698_ /*91210*/;
assign _4460_ = _4691_ ^ _4698_ /*91211*/;
assign _4696_ = _4697_ | _4699_ /*91208*/;
assign _4705_ = ~D[44] /*91207*/;
assign _4702_ = _4012_ & _4705_ /*91203*/;
assign _4703_ = _4012_ ^ _4705_ /*91206*/;
assign _4704_ = _4696_ & _4703_ /*91204*/;
assign _4461_ = _4696_ ^ _4703_ /*91205*/;
assign _4701_ = _4702_ | _4704_ /*91202*/;
assign _4710_ = ~D[45] /*91201*/;
assign _4707_ = _4013_ & _4710_ /*91197*/;
assign _4708_ = _4013_ ^ _4710_ /*91200*/;
assign _4709_ = _4701_ & _4708_ /*91198*/;
assign _4462_ = _4701_ ^ _4708_ /*91199*/;
assign _4706_ = _4707_ | _4709_ /*91196*/;
assign _4715_ = ~D[46] /*91195*/;
assign _4712_ = _4014_ & _4715_ /*91191*/;
assign _4713_ = _4014_ ^ _4715_ /*91194*/;
assign _4714_ = _4706_ & _4713_ /*91192*/;
assign _4463_ = _4706_ ^ _4713_ /*91193*/;
assign _4711_ = _4712_ | _4714_ /*91190*/;
assign _4720_ = ~D[47] /*91189*/;
assign _4717_ = _4015_ & _4720_ /*91185*/;
assign _4718_ = _4015_ ^ _4720_ /*91188*/;
assign _4719_ = _4711_ & _4718_ /*91186*/;
assign _4464_ = _4711_ ^ _4718_ /*91187*/;
assign _4716_ = _4717_ | _4719_ /*91184*/;
assign _4725_ = ~D[48] /*91183*/;
assign _4722_ = _4016_ & _4725_ /*91179*/;
assign _4723_ = _4016_ ^ _4725_ /*91182*/;
assign _4724_ = _4716_ & _4723_ /*91180*/;
assign _4465_ = _4716_ ^ _4723_ /*91181*/;
assign _4721_ = _4722_ | _4724_ /*91178*/;
assign _4730_ = ~D[49] /*91177*/;
assign _4727_ = _4017_ & _4730_ /*91173*/;
assign _4728_ = _4017_ ^ _4730_ /*91176*/;
assign _4729_ = _4721_ & _4728_ /*91174*/;
assign _4466_ = _4721_ ^ _4728_ /*91175*/;
assign _4726_ = _4727_ | _4729_ /*91172*/;
assign _4735_ = ~D[50] /*91171*/;
assign _4732_ = _4018_ & _4735_ /*91167*/;
assign _4733_ = _4018_ ^ _4735_ /*91170*/;
assign _4734_ = _4726_ & _4733_ /*91168*/;
assign _4467_ = _4726_ ^ _4733_ /*91169*/;
assign _4731_ = _4732_ | _4734_ /*91166*/;
assign _4740_ = ~D[51] /*91165*/;
assign _4737_ = _4019_ & _4740_ /*91161*/;
assign _4738_ = _4019_ ^ _4740_ /*91164*/;
assign _4739_ = _4731_ & _4738_ /*91162*/;
assign _4468_ = _4731_ ^ _4738_ /*91163*/;
assign _4736_ = _4737_ | _4739_ /*91160*/;
assign _4745_ = ~D[52] /*91159*/;
assign _4742_ = _4020_ & _4745_ /*91155*/;
assign _4743_ = _4020_ ^ _4745_ /*91158*/;
assign _4744_ = _4736_ & _4743_ /*91156*/;
assign _4469_ = _4736_ ^ _4743_ /*91157*/;
assign _4741_ = _4742_ | _4744_ /*91154*/;
assign _4750_ = ~D[53] /*91153*/;
assign _4747_ = _4021_ & _4750_ /*91149*/;
assign _4748_ = _4021_ ^ _4750_ /*91152*/;
assign _4749_ = _4741_ & _4748_ /*91150*/;
assign _4470_ = _4741_ ^ _4748_ /*91151*/;
assign _4746_ = _4747_ | _4749_ /*91148*/;
assign _4755_ = ~D[54] /*91147*/;
assign _4752_ = _4022_ & _4755_ /*91143*/;
assign _4753_ = _4022_ ^ _4755_ /*91146*/;
assign _4754_ = _4746_ & _4753_ /*91144*/;
assign _4471_ = _4746_ ^ _4753_ /*91145*/;
assign _4751_ = _4752_ | _4754_ /*91142*/;
assign _4760_ = ~D[55] /*91141*/;
assign _4757_ = _4023_ & _4760_ /*91137*/;
assign _4758_ = _4023_ ^ _4760_ /*91140*/;
assign _4759_ = _4751_ & _4758_ /*91138*/;
assign _4472_ = _4751_ ^ _4758_ /*91139*/;
assign _4756_ = _4757_ | _4759_ /*91136*/;
assign _4765_ = ~D[56] /*91135*/;
assign _4762_ = _4024_ & _4765_ /*91131*/;
assign _4763_ = _4024_ ^ _4765_ /*91134*/;
assign _4764_ = _4756_ & _4763_ /*91132*/;
assign _4473_ = _4756_ ^ _4763_ /*91133*/;
assign _4761_ = _4762_ | _4764_ /*91130*/;
assign _4770_ = ~D[57] /*91129*/;
assign _4767_ = _4025_ & _4770_ /*91125*/;
assign _4768_ = _4025_ ^ _4770_ /*91128*/;
assign _4769_ = _4761_ & _4768_ /*91126*/;
assign _4474_ = _4761_ ^ _4768_ /*91127*/;
assign _4766_ = _4767_ | _4769_ /*91124*/;
assign _4775_ = ~D[58] /*91123*/;
assign _4772_ = _4026_ & _4775_ /*91119*/;
assign _4773_ = _4026_ ^ _4775_ /*91122*/;
assign _4774_ = _4766_ & _4773_ /*91120*/;
assign _4475_ = _4766_ ^ _4773_ /*91121*/;
assign _4771_ = _4772_ | _4774_ /*91118*/;
assign _4780_ = ~D[59] /*91117*/;
assign _4777_ = _4027_ & _4780_ /*91113*/;
assign _4778_ = _4027_ ^ _4780_ /*91116*/;
assign _4779_ = _4771_ & _4778_ /*91114*/;
assign _4476_ = _4771_ ^ _4778_ /*91115*/;
assign _4776_ = _4777_ | _4779_ /*91112*/;
assign _4785_ = ~D[60] /*91111*/;
assign _4782_ = _4028_ & _4785_ /*91107*/;
assign _4783_ = _4028_ ^ _4785_ /*91110*/;
assign _4784_ = _4776_ & _4783_ /*91108*/;
assign _4477_ = _4776_ ^ _4783_ /*91109*/;
assign _4781_ = _4782_ | _4784_ /*91106*/;
assign _4790_ = ~D[61] /*91105*/;
assign _4787_ = _4029_ & _4790_ /*91101*/;
assign _4788_ = _4029_ ^ _4790_ /*91104*/;
assign _4789_ = _4781_ & _4788_ /*91102*/;
assign _4478_ = _4781_ ^ _4788_ /*91103*/;
assign _4786_ = _4787_ | _4789_ /*91100*/;
assign _4795_ = ~D[62] /*91099*/;
assign _4792_ = _4030_ & _4795_ /*91095*/;
assign _4793_ = _4030_ ^ _4795_ /*91098*/;
assign _4794_ = _4786_ & _4793_ /*91096*/;
assign _4479_ = _4786_ ^ _4793_ /*91097*/;
assign _4791_ = _4792_ | _4794_ /*91094*/;
assign _4796_ = _4031_ & oneWire /*91089*/;
assign _4797_ = _4031_ ^ oneWire /*91092*/;
assign _4798_ = _4791_ & _4797_ /*91090*/;
assign _4480_ = _4791_ ^ _4797_ /*91091*/;
assign Q[58] = _4796_ | _4798_ /*91088*/;
assign _4931_ = ~Q[58] /*90703*/;
assign _4930_ = _4931_ & D[0] /*90702*/;
assign _4933_ = _4417_ & _4930_ /*90697*/;
assign _4934_ = _4417_ ^ _4930_ /*90700*/;
assign _4935_ = zeroWire & _4934_ /*90698*/;
assign _4865_ = zeroWire ^ _4934_ /*90699*/;
assign _4932_ = _4933_ | _4935_ /*90696*/;
assign _4937_ = ~Q[58] /*90695*/;
assign _4936_ = _4937_ & D[1] /*90694*/;
assign _4939_ = _4418_ & _4936_ /*90689*/;
assign _4940_ = _4418_ ^ _4936_ /*90692*/;
assign _4941_ = _4932_ & _4940_ /*90690*/;
assign _4866_ = _4932_ ^ _4940_ /*90691*/;
assign _4938_ = _4939_ | _4941_ /*90688*/;
assign _4943_ = ~Q[58] /*90687*/;
assign _4942_ = _4943_ & D[2] /*90686*/;
assign _4945_ = _4419_ & _4942_ /*90681*/;
assign _4946_ = _4419_ ^ _4942_ /*90684*/;
assign _4947_ = _4938_ & _4946_ /*90682*/;
assign _4867_ = _4938_ ^ _4946_ /*90683*/;
assign _4944_ = _4945_ | _4947_ /*90680*/;
assign _4949_ = ~Q[58] /*90679*/;
assign _4948_ = _4949_ & D[3] /*90678*/;
assign _4951_ = _4420_ & _4948_ /*90673*/;
assign _4952_ = _4420_ ^ _4948_ /*90676*/;
assign _4953_ = _4944_ & _4952_ /*90674*/;
assign _4868_ = _4944_ ^ _4952_ /*90675*/;
assign _4950_ = _4951_ | _4953_ /*90672*/;
assign _4955_ = ~Q[58] /*90671*/;
assign _4954_ = _4955_ & D[4] /*90670*/;
assign _4957_ = _4421_ & _4954_ /*90665*/;
assign _4958_ = _4421_ ^ _4954_ /*90668*/;
assign _4959_ = _4950_ & _4958_ /*90666*/;
assign _4869_ = _4950_ ^ _4958_ /*90667*/;
assign _4956_ = _4957_ | _4959_ /*90664*/;
assign _4961_ = ~Q[58] /*90663*/;
assign _4960_ = _4961_ & D[5] /*90662*/;
assign _4963_ = _4422_ & _4960_ /*90657*/;
assign _4964_ = _4422_ ^ _4960_ /*90660*/;
assign _4965_ = _4956_ & _4964_ /*90658*/;
assign _4870_ = _4956_ ^ _4964_ /*90659*/;
assign _4962_ = _4963_ | _4965_ /*90656*/;
assign _4967_ = ~Q[58] /*90655*/;
assign _4966_ = _4967_ & D[6] /*90654*/;
assign _4969_ = _4423_ & _4966_ /*90649*/;
assign _4970_ = _4423_ ^ _4966_ /*90652*/;
assign _4971_ = _4962_ & _4970_ /*90650*/;
assign _4871_ = _4962_ ^ _4970_ /*90651*/;
assign _4968_ = _4969_ | _4971_ /*90648*/;
assign _4973_ = ~Q[58] /*90647*/;
assign _4972_ = _4973_ & D[7] /*90646*/;
assign _4975_ = _4424_ & _4972_ /*90641*/;
assign _4976_ = _4424_ ^ _4972_ /*90644*/;
assign _4977_ = _4968_ & _4976_ /*90642*/;
assign _4872_ = _4968_ ^ _4976_ /*90643*/;
assign _4974_ = _4975_ | _4977_ /*90640*/;
assign _4979_ = ~Q[58] /*90639*/;
assign _4978_ = _4979_ & D[8] /*90638*/;
assign _4981_ = _4425_ & _4978_ /*90633*/;
assign _4982_ = _4425_ ^ _4978_ /*90636*/;
assign _4983_ = _4974_ & _4982_ /*90634*/;
assign _4873_ = _4974_ ^ _4982_ /*90635*/;
assign _4980_ = _4981_ | _4983_ /*90632*/;
assign _4985_ = ~Q[58] /*90631*/;
assign _4984_ = _4985_ & D[9] /*90630*/;
assign _4987_ = _4426_ & _4984_ /*90625*/;
assign _4988_ = _4426_ ^ _4984_ /*90628*/;
assign _4989_ = _4980_ & _4988_ /*90626*/;
assign _4874_ = _4980_ ^ _4988_ /*90627*/;
assign _4986_ = _4987_ | _4989_ /*90624*/;
assign _4991_ = ~Q[58] /*90623*/;
assign _4990_ = _4991_ & D[10] /*90622*/;
assign _4993_ = _4427_ & _4990_ /*90617*/;
assign _4994_ = _4427_ ^ _4990_ /*90620*/;
assign _4995_ = _4986_ & _4994_ /*90618*/;
assign _4875_ = _4986_ ^ _4994_ /*90619*/;
assign _4992_ = _4993_ | _4995_ /*90616*/;
assign _4997_ = ~Q[58] /*90615*/;
assign _4996_ = _4997_ & D[11] /*90614*/;
assign _4999_ = _4428_ & _4996_ /*90609*/;
assign _5000_ = _4428_ ^ _4996_ /*90612*/;
assign _5001_ = _4992_ & _5000_ /*90610*/;
assign _4876_ = _4992_ ^ _5000_ /*90611*/;
assign _4998_ = _4999_ | _5001_ /*90608*/;
assign _5003_ = ~Q[58] /*90607*/;
assign _5002_ = _5003_ & D[12] /*90606*/;
assign _5005_ = _4429_ & _5002_ /*90601*/;
assign _5006_ = _4429_ ^ _5002_ /*90604*/;
assign _5007_ = _4998_ & _5006_ /*90602*/;
assign _4877_ = _4998_ ^ _5006_ /*90603*/;
assign _5004_ = _5005_ | _5007_ /*90600*/;
assign _5009_ = ~Q[58] /*90599*/;
assign _5008_ = _5009_ & D[13] /*90598*/;
assign _5011_ = _4430_ & _5008_ /*90593*/;
assign _5012_ = _4430_ ^ _5008_ /*90596*/;
assign _5013_ = _5004_ & _5012_ /*90594*/;
assign _4878_ = _5004_ ^ _5012_ /*90595*/;
assign _5010_ = _5011_ | _5013_ /*90592*/;
assign _5015_ = ~Q[58] /*90591*/;
assign _5014_ = _5015_ & D[14] /*90590*/;
assign _5017_ = _4431_ & _5014_ /*90585*/;
assign _5018_ = _4431_ ^ _5014_ /*90588*/;
assign _5019_ = _5010_ & _5018_ /*90586*/;
assign _4879_ = _5010_ ^ _5018_ /*90587*/;
assign _5016_ = _5017_ | _5019_ /*90584*/;
assign _5021_ = ~Q[58] /*90583*/;
assign _5020_ = _5021_ & D[15] /*90582*/;
assign _5023_ = _4432_ & _5020_ /*90577*/;
assign _5024_ = _4432_ ^ _5020_ /*90580*/;
assign _5025_ = _5016_ & _5024_ /*90578*/;
assign _4880_ = _5016_ ^ _5024_ /*90579*/;
assign _5022_ = _5023_ | _5025_ /*90576*/;
assign _5027_ = ~Q[58] /*90575*/;
assign _5026_ = _5027_ & D[16] /*90574*/;
assign _5029_ = _4433_ & _5026_ /*90569*/;
assign _5030_ = _4433_ ^ _5026_ /*90572*/;
assign _5031_ = _5022_ & _5030_ /*90570*/;
assign _4881_ = _5022_ ^ _5030_ /*90571*/;
assign _5028_ = _5029_ | _5031_ /*90568*/;
assign _5033_ = ~Q[58] /*90567*/;
assign _5032_ = _5033_ & D[17] /*90566*/;
assign _5035_ = _4434_ & _5032_ /*90561*/;
assign _5036_ = _4434_ ^ _5032_ /*90564*/;
assign _5037_ = _5028_ & _5036_ /*90562*/;
assign _4882_ = _5028_ ^ _5036_ /*90563*/;
assign _5034_ = _5035_ | _5037_ /*90560*/;
assign _5039_ = ~Q[58] /*90559*/;
assign _5038_ = _5039_ & D[18] /*90558*/;
assign _5041_ = _4435_ & _5038_ /*90553*/;
assign _5042_ = _4435_ ^ _5038_ /*90556*/;
assign _5043_ = _5034_ & _5042_ /*90554*/;
assign _4883_ = _5034_ ^ _5042_ /*90555*/;
assign _5040_ = _5041_ | _5043_ /*90552*/;
assign _5045_ = ~Q[58] /*90551*/;
assign _5044_ = _5045_ & D[19] /*90550*/;
assign _5047_ = _4436_ & _5044_ /*90545*/;
assign _5048_ = _4436_ ^ _5044_ /*90548*/;
assign _5049_ = _5040_ & _5048_ /*90546*/;
assign _4884_ = _5040_ ^ _5048_ /*90547*/;
assign _5046_ = _5047_ | _5049_ /*90544*/;
assign _5051_ = ~Q[58] /*90543*/;
assign _5050_ = _5051_ & D[20] /*90542*/;
assign _5053_ = _4437_ & _5050_ /*90537*/;
assign _5054_ = _4437_ ^ _5050_ /*90540*/;
assign _5055_ = _5046_ & _5054_ /*90538*/;
assign _4885_ = _5046_ ^ _5054_ /*90539*/;
assign _5052_ = _5053_ | _5055_ /*90536*/;
assign _5057_ = ~Q[58] /*90535*/;
assign _5056_ = _5057_ & D[21] /*90534*/;
assign _5059_ = _4438_ & _5056_ /*90529*/;
assign _5060_ = _4438_ ^ _5056_ /*90532*/;
assign _5061_ = _5052_ & _5060_ /*90530*/;
assign _4886_ = _5052_ ^ _5060_ /*90531*/;
assign _5058_ = _5059_ | _5061_ /*90528*/;
assign _5063_ = ~Q[58] /*90527*/;
assign _5062_ = _5063_ & D[22] /*90526*/;
assign _5065_ = _4439_ & _5062_ /*90521*/;
assign _5066_ = _4439_ ^ _5062_ /*90524*/;
assign _5067_ = _5058_ & _5066_ /*90522*/;
assign _4887_ = _5058_ ^ _5066_ /*90523*/;
assign _5064_ = _5065_ | _5067_ /*90520*/;
assign _5069_ = ~Q[58] /*90519*/;
assign _5068_ = _5069_ & D[23] /*90518*/;
assign _5071_ = _4440_ & _5068_ /*90513*/;
assign _5072_ = _4440_ ^ _5068_ /*90516*/;
assign _5073_ = _5064_ & _5072_ /*90514*/;
assign _4888_ = _5064_ ^ _5072_ /*90515*/;
assign _5070_ = _5071_ | _5073_ /*90512*/;
assign _5075_ = ~Q[58] /*90511*/;
assign _5074_ = _5075_ & D[24] /*90510*/;
assign _5077_ = _4441_ & _5074_ /*90505*/;
assign _5078_ = _4441_ ^ _5074_ /*90508*/;
assign _5079_ = _5070_ & _5078_ /*90506*/;
assign _4889_ = _5070_ ^ _5078_ /*90507*/;
assign _5076_ = _5077_ | _5079_ /*90504*/;
assign _5081_ = ~Q[58] /*90503*/;
assign _5080_ = _5081_ & D[25] /*90502*/;
assign _5083_ = _4442_ & _5080_ /*90497*/;
assign _5084_ = _4442_ ^ _5080_ /*90500*/;
assign _5085_ = _5076_ & _5084_ /*90498*/;
assign _4890_ = _5076_ ^ _5084_ /*90499*/;
assign _5082_ = _5083_ | _5085_ /*90496*/;
assign _5087_ = ~Q[58] /*90495*/;
assign _5086_ = _5087_ & D[26] /*90494*/;
assign _5089_ = _4443_ & _5086_ /*90489*/;
assign _5090_ = _4443_ ^ _5086_ /*90492*/;
assign _5091_ = _5082_ & _5090_ /*90490*/;
assign _4891_ = _5082_ ^ _5090_ /*90491*/;
assign _5088_ = _5089_ | _5091_ /*90488*/;
assign _5093_ = ~Q[58] /*90487*/;
assign _5092_ = _5093_ & D[27] /*90486*/;
assign _5095_ = _4444_ & _5092_ /*90481*/;
assign _5096_ = _4444_ ^ _5092_ /*90484*/;
assign _5097_ = _5088_ & _5096_ /*90482*/;
assign _4892_ = _5088_ ^ _5096_ /*90483*/;
assign _5094_ = _5095_ | _5097_ /*90480*/;
assign _5099_ = ~Q[58] /*90479*/;
assign _5098_ = _5099_ & D[28] /*90478*/;
assign _5101_ = _4445_ & _5098_ /*90473*/;
assign _5102_ = _4445_ ^ _5098_ /*90476*/;
assign _5103_ = _5094_ & _5102_ /*90474*/;
assign _4893_ = _5094_ ^ _5102_ /*90475*/;
assign _5100_ = _5101_ | _5103_ /*90472*/;
assign _5105_ = ~Q[58] /*90471*/;
assign _5104_ = _5105_ & D[29] /*90470*/;
assign _5107_ = _4446_ & _5104_ /*90465*/;
assign _5108_ = _4446_ ^ _5104_ /*90468*/;
assign _5109_ = _5100_ & _5108_ /*90466*/;
assign _4894_ = _5100_ ^ _5108_ /*90467*/;
assign _5106_ = _5107_ | _5109_ /*90464*/;
assign _5111_ = ~Q[58] /*90463*/;
assign _5110_ = _5111_ & D[30] /*90462*/;
assign _5113_ = _4447_ & _5110_ /*90457*/;
assign _5114_ = _4447_ ^ _5110_ /*90460*/;
assign _5115_ = _5106_ & _5114_ /*90458*/;
assign _4895_ = _5106_ ^ _5114_ /*90459*/;
assign _5112_ = _5113_ | _5115_ /*90456*/;
assign _5117_ = ~Q[58] /*90455*/;
assign _5116_ = _5117_ & D[31] /*90454*/;
assign _5119_ = _4448_ & _5116_ /*90449*/;
assign _5120_ = _4448_ ^ _5116_ /*90452*/;
assign _5121_ = _5112_ & _5120_ /*90450*/;
assign _4896_ = _5112_ ^ _5120_ /*90451*/;
assign _5118_ = _5119_ | _5121_ /*90448*/;
assign _5123_ = ~Q[58] /*90447*/;
assign _5122_ = _5123_ & D[32] /*90446*/;
assign _5125_ = _4449_ & _5122_ /*90441*/;
assign _5126_ = _4449_ ^ _5122_ /*90444*/;
assign _5127_ = _5118_ & _5126_ /*90442*/;
assign _4897_ = _5118_ ^ _5126_ /*90443*/;
assign _5124_ = _5125_ | _5127_ /*90440*/;
assign _5129_ = ~Q[58] /*90439*/;
assign _5128_ = _5129_ & D[33] /*90438*/;
assign _5131_ = _4450_ & _5128_ /*90433*/;
assign _5132_ = _4450_ ^ _5128_ /*90436*/;
assign _5133_ = _5124_ & _5132_ /*90434*/;
assign _4898_ = _5124_ ^ _5132_ /*90435*/;
assign _5130_ = _5131_ | _5133_ /*90432*/;
assign _5135_ = ~Q[58] /*90431*/;
assign _5134_ = _5135_ & D[34] /*90430*/;
assign _5137_ = _4451_ & _5134_ /*90425*/;
assign _5138_ = _4451_ ^ _5134_ /*90428*/;
assign _5139_ = _5130_ & _5138_ /*90426*/;
assign _4899_ = _5130_ ^ _5138_ /*90427*/;
assign _5136_ = _5137_ | _5139_ /*90424*/;
assign _5141_ = ~Q[58] /*90423*/;
assign _5140_ = _5141_ & D[35] /*90422*/;
assign _5143_ = _4452_ & _5140_ /*90417*/;
assign _5144_ = _4452_ ^ _5140_ /*90420*/;
assign _5145_ = _5136_ & _5144_ /*90418*/;
assign _4900_ = _5136_ ^ _5144_ /*90419*/;
assign _5142_ = _5143_ | _5145_ /*90416*/;
assign _5147_ = ~Q[58] /*90415*/;
assign _5146_ = _5147_ & D[36] /*90414*/;
assign _5149_ = _4453_ & _5146_ /*90409*/;
assign _5150_ = _4453_ ^ _5146_ /*90412*/;
assign _5151_ = _5142_ & _5150_ /*90410*/;
assign _4901_ = _5142_ ^ _5150_ /*90411*/;
assign _5148_ = _5149_ | _5151_ /*90408*/;
assign _5153_ = ~Q[58] /*90407*/;
assign _5152_ = _5153_ & D[37] /*90406*/;
assign _5155_ = _4454_ & _5152_ /*90401*/;
assign _5156_ = _4454_ ^ _5152_ /*90404*/;
assign _5157_ = _5148_ & _5156_ /*90402*/;
assign _4902_ = _5148_ ^ _5156_ /*90403*/;
assign _5154_ = _5155_ | _5157_ /*90400*/;
assign _5159_ = ~Q[58] /*90399*/;
assign _5158_ = _5159_ & D[38] /*90398*/;
assign _5161_ = _4455_ & _5158_ /*90393*/;
assign _5162_ = _4455_ ^ _5158_ /*90396*/;
assign _5163_ = _5154_ & _5162_ /*90394*/;
assign _4903_ = _5154_ ^ _5162_ /*90395*/;
assign _5160_ = _5161_ | _5163_ /*90392*/;
assign _5165_ = ~Q[58] /*90391*/;
assign _5164_ = _5165_ & D[39] /*90390*/;
assign _5167_ = _4456_ & _5164_ /*90385*/;
assign _5168_ = _4456_ ^ _5164_ /*90388*/;
assign _5169_ = _5160_ & _5168_ /*90386*/;
assign _4904_ = _5160_ ^ _5168_ /*90387*/;
assign _5166_ = _5167_ | _5169_ /*90384*/;
assign _5171_ = ~Q[58] /*90383*/;
assign _5170_ = _5171_ & D[40] /*90382*/;
assign _5173_ = _4457_ & _5170_ /*90377*/;
assign _5174_ = _4457_ ^ _5170_ /*90380*/;
assign _5175_ = _5166_ & _5174_ /*90378*/;
assign _4905_ = _5166_ ^ _5174_ /*90379*/;
assign _5172_ = _5173_ | _5175_ /*90376*/;
assign _5177_ = ~Q[58] /*90375*/;
assign _5176_ = _5177_ & D[41] /*90374*/;
assign _5179_ = _4458_ & _5176_ /*90369*/;
assign _5180_ = _4458_ ^ _5176_ /*90372*/;
assign _5181_ = _5172_ & _5180_ /*90370*/;
assign _4906_ = _5172_ ^ _5180_ /*90371*/;
assign _5178_ = _5179_ | _5181_ /*90368*/;
assign _5183_ = ~Q[58] /*90367*/;
assign _5182_ = _5183_ & D[42] /*90366*/;
assign _5185_ = _4459_ & _5182_ /*90361*/;
assign _5186_ = _4459_ ^ _5182_ /*90364*/;
assign _5187_ = _5178_ & _5186_ /*90362*/;
assign _4907_ = _5178_ ^ _5186_ /*90363*/;
assign _5184_ = _5185_ | _5187_ /*90360*/;
assign _5189_ = ~Q[58] /*90359*/;
assign _5188_ = _5189_ & D[43] /*90358*/;
assign _5191_ = _4460_ & _5188_ /*90353*/;
assign _5192_ = _4460_ ^ _5188_ /*90356*/;
assign _5193_ = _5184_ & _5192_ /*90354*/;
assign _4908_ = _5184_ ^ _5192_ /*90355*/;
assign _5190_ = _5191_ | _5193_ /*90352*/;
assign _5195_ = ~Q[58] /*90351*/;
assign _5194_ = _5195_ & D[44] /*90350*/;
assign _5197_ = _4461_ & _5194_ /*90345*/;
assign _5198_ = _4461_ ^ _5194_ /*90348*/;
assign _5199_ = _5190_ & _5198_ /*90346*/;
assign _4909_ = _5190_ ^ _5198_ /*90347*/;
assign _5196_ = _5197_ | _5199_ /*90344*/;
assign _5201_ = ~Q[58] /*90343*/;
assign _5200_ = _5201_ & D[45] /*90342*/;
assign _5203_ = _4462_ & _5200_ /*90337*/;
assign _5204_ = _4462_ ^ _5200_ /*90340*/;
assign _5205_ = _5196_ & _5204_ /*90338*/;
assign _4910_ = _5196_ ^ _5204_ /*90339*/;
assign _5202_ = _5203_ | _5205_ /*90336*/;
assign _5207_ = ~Q[58] /*90335*/;
assign _5206_ = _5207_ & D[46] /*90334*/;
assign _5209_ = _4463_ & _5206_ /*90329*/;
assign _5210_ = _4463_ ^ _5206_ /*90332*/;
assign _5211_ = _5202_ & _5210_ /*90330*/;
assign _4911_ = _5202_ ^ _5210_ /*90331*/;
assign _5208_ = _5209_ | _5211_ /*90328*/;
assign _5213_ = ~Q[58] /*90327*/;
assign _5212_ = _5213_ & D[47] /*90326*/;
assign _5215_ = _4464_ & _5212_ /*90321*/;
assign _5216_ = _4464_ ^ _5212_ /*90324*/;
assign _5217_ = _5208_ & _5216_ /*90322*/;
assign _4912_ = _5208_ ^ _5216_ /*90323*/;
assign _5214_ = _5215_ | _5217_ /*90320*/;
assign _5219_ = ~Q[58] /*90319*/;
assign _5218_ = _5219_ & D[48] /*90318*/;
assign _5221_ = _4465_ & _5218_ /*90313*/;
assign _5222_ = _4465_ ^ _5218_ /*90316*/;
assign _5223_ = _5214_ & _5222_ /*90314*/;
assign _4913_ = _5214_ ^ _5222_ /*90315*/;
assign _5220_ = _5221_ | _5223_ /*90312*/;
assign _5225_ = ~Q[58] /*90311*/;
assign _5224_ = _5225_ & D[49] /*90310*/;
assign _5227_ = _4466_ & _5224_ /*90305*/;
assign _5228_ = _4466_ ^ _5224_ /*90308*/;
assign _5229_ = _5220_ & _5228_ /*90306*/;
assign _4914_ = _5220_ ^ _5228_ /*90307*/;
assign _5226_ = _5227_ | _5229_ /*90304*/;
assign _5231_ = ~Q[58] /*90303*/;
assign _5230_ = _5231_ & D[50] /*90302*/;
assign _5233_ = _4467_ & _5230_ /*90297*/;
assign _5234_ = _4467_ ^ _5230_ /*90300*/;
assign _5235_ = _5226_ & _5234_ /*90298*/;
assign _4915_ = _5226_ ^ _5234_ /*90299*/;
assign _5232_ = _5233_ | _5235_ /*90296*/;
assign _5237_ = ~Q[58] /*90295*/;
assign _5236_ = _5237_ & D[51] /*90294*/;
assign _5239_ = _4468_ & _5236_ /*90289*/;
assign _5240_ = _4468_ ^ _5236_ /*90292*/;
assign _5241_ = _5232_ & _5240_ /*90290*/;
assign _4916_ = _5232_ ^ _5240_ /*90291*/;
assign _5238_ = _5239_ | _5241_ /*90288*/;
assign _5243_ = ~Q[58] /*90287*/;
assign _5242_ = _5243_ & D[52] /*90286*/;
assign _5245_ = _4469_ & _5242_ /*90281*/;
assign _5246_ = _4469_ ^ _5242_ /*90284*/;
assign _5247_ = _5238_ & _5246_ /*90282*/;
assign _4917_ = _5238_ ^ _5246_ /*90283*/;
assign _5244_ = _5245_ | _5247_ /*90280*/;
assign _5249_ = ~Q[58] /*90279*/;
assign _5248_ = _5249_ & D[53] /*90278*/;
assign _5251_ = _4470_ & _5248_ /*90273*/;
assign _5252_ = _4470_ ^ _5248_ /*90276*/;
assign _5253_ = _5244_ & _5252_ /*90274*/;
assign _4918_ = _5244_ ^ _5252_ /*90275*/;
assign _5250_ = _5251_ | _5253_ /*90272*/;
assign _5255_ = ~Q[58] /*90271*/;
assign _5254_ = _5255_ & D[54] /*90270*/;
assign _5257_ = _4471_ & _5254_ /*90265*/;
assign _5258_ = _4471_ ^ _5254_ /*90268*/;
assign _5259_ = _5250_ & _5258_ /*90266*/;
assign _4919_ = _5250_ ^ _5258_ /*90267*/;
assign _5256_ = _5257_ | _5259_ /*90264*/;
assign _5261_ = ~Q[58] /*90263*/;
assign _5260_ = _5261_ & D[55] /*90262*/;
assign _5263_ = _4472_ & _5260_ /*90257*/;
assign _5264_ = _4472_ ^ _5260_ /*90260*/;
assign _5265_ = _5256_ & _5264_ /*90258*/;
assign _4920_ = _5256_ ^ _5264_ /*90259*/;
assign _5262_ = _5263_ | _5265_ /*90256*/;
assign _5267_ = ~Q[58] /*90255*/;
assign _5266_ = _5267_ & D[56] /*90254*/;
assign _5269_ = _4473_ & _5266_ /*90249*/;
assign _5270_ = _4473_ ^ _5266_ /*90252*/;
assign _5271_ = _5262_ & _5270_ /*90250*/;
assign _4921_ = _5262_ ^ _5270_ /*90251*/;
assign _5268_ = _5269_ | _5271_ /*90248*/;
assign _5273_ = ~Q[58] /*90247*/;
assign _5272_ = _5273_ & D[57] /*90246*/;
assign _5275_ = _4474_ & _5272_ /*90241*/;
assign _5276_ = _4474_ ^ _5272_ /*90244*/;
assign _5277_ = _5268_ & _5276_ /*90242*/;
assign _4922_ = _5268_ ^ _5276_ /*90243*/;
assign _5274_ = _5275_ | _5277_ /*90240*/;
assign _5279_ = ~Q[58] /*90239*/;
assign _5278_ = _5279_ & D[58] /*90238*/;
assign _5281_ = _4475_ & _5278_ /*90233*/;
assign _5282_ = _4475_ ^ _5278_ /*90236*/;
assign _5283_ = _5274_ & _5282_ /*90234*/;
assign _4923_ = _5274_ ^ _5282_ /*90235*/;
assign _5280_ = _5281_ | _5283_ /*90232*/;
assign _5285_ = ~Q[58] /*90231*/;
assign _5284_ = _5285_ & D[59] /*90230*/;
assign _5287_ = _4476_ & _5284_ /*90225*/;
assign _5288_ = _4476_ ^ _5284_ /*90228*/;
assign _5289_ = _5280_ & _5288_ /*90226*/;
assign _4924_ = _5280_ ^ _5288_ /*90227*/;
assign _5286_ = _5287_ | _5289_ /*90224*/;
assign _5291_ = ~Q[58] /*90223*/;
assign _5290_ = _5291_ & D[60] /*90222*/;
assign _5293_ = _4477_ & _5290_ /*90217*/;
assign _5294_ = _4477_ ^ _5290_ /*90220*/;
assign _5295_ = _5286_ & _5294_ /*90218*/;
assign _4925_ = _5286_ ^ _5294_ /*90219*/;
assign _5292_ = _5293_ | _5295_ /*90216*/;
assign _5297_ = ~Q[58] /*90215*/;
assign _5296_ = _5297_ & D[61] /*90214*/;
assign _5299_ = _4478_ & _5296_ /*90209*/;
assign _5300_ = _4478_ ^ _5296_ /*90212*/;
assign _5301_ = _5292_ & _5300_ /*90210*/;
assign _4926_ = _5292_ ^ _5300_ /*90211*/;
assign _5298_ = _5299_ | _5301_ /*90208*/;
assign _5303_ = ~Q[58] /*90207*/;
assign _5302_ = _5303_ & D[62] /*90206*/;
assign _5305_ = _4479_ & _5302_ /*90201*/;
assign _5306_ = _4479_ ^ _5302_ /*90204*/;
assign _5307_ = _5298_ & _5306_ /*90202*/;
assign _4927_ = _5298_ ^ _5306_ /*90203*/;
assign _5304_ = _5305_ | _5307_ /*90200*/;
assign _5309_ = ~Q[58] /*90199*/;
assign _5308_ = _5309_ & zeroWire /*90198*/;
assign _5310_ = _4480_ ^ _5308_ /*90196*/;
assign _4928_ = _5310_ ^ _5304_ /*90195*/;
assign _5381_ = ~D[0] /*89941*/;
assign _5378_ = R_0[57] & _5381_ /*89937*/;
assign _5379_ = R_0[57] ^ _5381_ /*89940*/;
assign _5380_ = oneWire & _5379_ /*89938*/;
assign _5313_ = oneWire ^ _5379_ /*89939*/;
assign _5377_ = _5378_ | _5380_ /*89936*/;
assign _5386_ = ~D[1] /*89935*/;
assign _5383_ = _4865_ & _5386_ /*89931*/;
assign _5384_ = _4865_ ^ _5386_ /*89934*/;
assign _5385_ = _5377_ & _5384_ /*89932*/;
assign _5314_ = _5377_ ^ _5384_ /*89933*/;
assign _5382_ = _5383_ | _5385_ /*89930*/;
assign _5391_ = ~D[2] /*89929*/;
assign _5388_ = _4866_ & _5391_ /*89925*/;
assign _5389_ = _4866_ ^ _5391_ /*89928*/;
assign _5390_ = _5382_ & _5389_ /*89926*/;
assign _5315_ = _5382_ ^ _5389_ /*89927*/;
assign _5387_ = _5388_ | _5390_ /*89924*/;
assign _5396_ = ~D[3] /*89923*/;
assign _5393_ = _4867_ & _5396_ /*89919*/;
assign _5394_ = _4867_ ^ _5396_ /*89922*/;
assign _5395_ = _5387_ & _5394_ /*89920*/;
assign _5316_ = _5387_ ^ _5394_ /*89921*/;
assign _5392_ = _5393_ | _5395_ /*89918*/;
assign _5401_ = ~D[4] /*89917*/;
assign _5398_ = _4868_ & _5401_ /*89913*/;
assign _5399_ = _4868_ ^ _5401_ /*89916*/;
assign _5400_ = _5392_ & _5399_ /*89914*/;
assign _5317_ = _5392_ ^ _5399_ /*89915*/;
assign _5397_ = _5398_ | _5400_ /*89912*/;
assign _5406_ = ~D[5] /*89911*/;
assign _5403_ = _4869_ & _5406_ /*89907*/;
assign _5404_ = _4869_ ^ _5406_ /*89910*/;
assign _5405_ = _5397_ & _5404_ /*89908*/;
assign _5318_ = _5397_ ^ _5404_ /*89909*/;
assign _5402_ = _5403_ | _5405_ /*89906*/;
assign _5411_ = ~D[6] /*89905*/;
assign _5408_ = _4870_ & _5411_ /*89901*/;
assign _5409_ = _4870_ ^ _5411_ /*89904*/;
assign _5410_ = _5402_ & _5409_ /*89902*/;
assign _5319_ = _5402_ ^ _5409_ /*89903*/;
assign _5407_ = _5408_ | _5410_ /*89900*/;
assign _5416_ = ~D[7] /*89899*/;
assign _5413_ = _4871_ & _5416_ /*89895*/;
assign _5414_ = _4871_ ^ _5416_ /*89898*/;
assign _5415_ = _5407_ & _5414_ /*89896*/;
assign _5320_ = _5407_ ^ _5414_ /*89897*/;
assign _5412_ = _5413_ | _5415_ /*89894*/;
assign _5421_ = ~D[8] /*89893*/;
assign _5418_ = _4872_ & _5421_ /*89889*/;
assign _5419_ = _4872_ ^ _5421_ /*89892*/;
assign _5420_ = _5412_ & _5419_ /*89890*/;
assign _5321_ = _5412_ ^ _5419_ /*89891*/;
assign _5417_ = _5418_ | _5420_ /*89888*/;
assign _5426_ = ~D[9] /*89887*/;
assign _5423_ = _4873_ & _5426_ /*89883*/;
assign _5424_ = _4873_ ^ _5426_ /*89886*/;
assign _5425_ = _5417_ & _5424_ /*89884*/;
assign _5322_ = _5417_ ^ _5424_ /*89885*/;
assign _5422_ = _5423_ | _5425_ /*89882*/;
assign _5431_ = ~D[10] /*89881*/;
assign _5428_ = _4874_ & _5431_ /*89877*/;
assign _5429_ = _4874_ ^ _5431_ /*89880*/;
assign _5430_ = _5422_ & _5429_ /*89878*/;
assign _5323_ = _5422_ ^ _5429_ /*89879*/;
assign _5427_ = _5428_ | _5430_ /*89876*/;
assign _5436_ = ~D[11] /*89875*/;
assign _5433_ = _4875_ & _5436_ /*89871*/;
assign _5434_ = _4875_ ^ _5436_ /*89874*/;
assign _5435_ = _5427_ & _5434_ /*89872*/;
assign _5324_ = _5427_ ^ _5434_ /*89873*/;
assign _5432_ = _5433_ | _5435_ /*89870*/;
assign _5441_ = ~D[12] /*89869*/;
assign _5438_ = _4876_ & _5441_ /*89865*/;
assign _5439_ = _4876_ ^ _5441_ /*89868*/;
assign _5440_ = _5432_ & _5439_ /*89866*/;
assign _5325_ = _5432_ ^ _5439_ /*89867*/;
assign _5437_ = _5438_ | _5440_ /*89864*/;
assign _5446_ = ~D[13] /*89863*/;
assign _5443_ = _4877_ & _5446_ /*89859*/;
assign _5444_ = _4877_ ^ _5446_ /*89862*/;
assign _5445_ = _5437_ & _5444_ /*89860*/;
assign _5326_ = _5437_ ^ _5444_ /*89861*/;
assign _5442_ = _5443_ | _5445_ /*89858*/;
assign _5451_ = ~D[14] /*89857*/;
assign _5448_ = _4878_ & _5451_ /*89853*/;
assign _5449_ = _4878_ ^ _5451_ /*89856*/;
assign _5450_ = _5442_ & _5449_ /*89854*/;
assign _5327_ = _5442_ ^ _5449_ /*89855*/;
assign _5447_ = _5448_ | _5450_ /*89852*/;
assign _5456_ = ~D[15] /*89851*/;
assign _5453_ = _4879_ & _5456_ /*89847*/;
assign _5454_ = _4879_ ^ _5456_ /*89850*/;
assign _5455_ = _5447_ & _5454_ /*89848*/;
assign _5328_ = _5447_ ^ _5454_ /*89849*/;
assign _5452_ = _5453_ | _5455_ /*89846*/;
assign _5461_ = ~D[16] /*89845*/;
assign _5458_ = _4880_ & _5461_ /*89841*/;
assign _5459_ = _4880_ ^ _5461_ /*89844*/;
assign _5460_ = _5452_ & _5459_ /*89842*/;
assign _5329_ = _5452_ ^ _5459_ /*89843*/;
assign _5457_ = _5458_ | _5460_ /*89840*/;
assign _5466_ = ~D[17] /*89839*/;
assign _5463_ = _4881_ & _5466_ /*89835*/;
assign _5464_ = _4881_ ^ _5466_ /*89838*/;
assign _5465_ = _5457_ & _5464_ /*89836*/;
assign _5330_ = _5457_ ^ _5464_ /*89837*/;
assign _5462_ = _5463_ | _5465_ /*89834*/;
assign _5471_ = ~D[18] /*89833*/;
assign _5468_ = _4882_ & _5471_ /*89829*/;
assign _5469_ = _4882_ ^ _5471_ /*89832*/;
assign _5470_ = _5462_ & _5469_ /*89830*/;
assign _5331_ = _5462_ ^ _5469_ /*89831*/;
assign _5467_ = _5468_ | _5470_ /*89828*/;
assign _5476_ = ~D[19] /*89827*/;
assign _5473_ = _4883_ & _5476_ /*89823*/;
assign _5474_ = _4883_ ^ _5476_ /*89826*/;
assign _5475_ = _5467_ & _5474_ /*89824*/;
assign _5332_ = _5467_ ^ _5474_ /*89825*/;
assign _5472_ = _5473_ | _5475_ /*89822*/;
assign _5481_ = ~D[20] /*89821*/;
assign _5478_ = _4884_ & _5481_ /*89817*/;
assign _5479_ = _4884_ ^ _5481_ /*89820*/;
assign _5480_ = _5472_ & _5479_ /*89818*/;
assign _5333_ = _5472_ ^ _5479_ /*89819*/;
assign _5477_ = _5478_ | _5480_ /*89816*/;
assign _5486_ = ~D[21] /*89815*/;
assign _5483_ = _4885_ & _5486_ /*89811*/;
assign _5484_ = _4885_ ^ _5486_ /*89814*/;
assign _5485_ = _5477_ & _5484_ /*89812*/;
assign _5334_ = _5477_ ^ _5484_ /*89813*/;
assign _5482_ = _5483_ | _5485_ /*89810*/;
assign _5491_ = ~D[22] /*89809*/;
assign _5488_ = _4886_ & _5491_ /*89805*/;
assign _5489_ = _4886_ ^ _5491_ /*89808*/;
assign _5490_ = _5482_ & _5489_ /*89806*/;
assign _5335_ = _5482_ ^ _5489_ /*89807*/;
assign _5487_ = _5488_ | _5490_ /*89804*/;
assign _5496_ = ~D[23] /*89803*/;
assign _5493_ = _4887_ & _5496_ /*89799*/;
assign _5494_ = _4887_ ^ _5496_ /*89802*/;
assign _5495_ = _5487_ & _5494_ /*89800*/;
assign _5336_ = _5487_ ^ _5494_ /*89801*/;
assign _5492_ = _5493_ | _5495_ /*89798*/;
assign _5501_ = ~D[24] /*89797*/;
assign _5498_ = _4888_ & _5501_ /*89793*/;
assign _5499_ = _4888_ ^ _5501_ /*89796*/;
assign _5500_ = _5492_ & _5499_ /*89794*/;
assign _5337_ = _5492_ ^ _5499_ /*89795*/;
assign _5497_ = _5498_ | _5500_ /*89792*/;
assign _5506_ = ~D[25] /*89791*/;
assign _5503_ = _4889_ & _5506_ /*89787*/;
assign _5504_ = _4889_ ^ _5506_ /*89790*/;
assign _5505_ = _5497_ & _5504_ /*89788*/;
assign _5338_ = _5497_ ^ _5504_ /*89789*/;
assign _5502_ = _5503_ | _5505_ /*89786*/;
assign _5511_ = ~D[26] /*89785*/;
assign _5508_ = _4890_ & _5511_ /*89781*/;
assign _5509_ = _4890_ ^ _5511_ /*89784*/;
assign _5510_ = _5502_ & _5509_ /*89782*/;
assign _5339_ = _5502_ ^ _5509_ /*89783*/;
assign _5507_ = _5508_ | _5510_ /*89780*/;
assign _5516_ = ~D[27] /*89779*/;
assign _5513_ = _4891_ & _5516_ /*89775*/;
assign _5514_ = _4891_ ^ _5516_ /*89778*/;
assign _5515_ = _5507_ & _5514_ /*89776*/;
assign _5340_ = _5507_ ^ _5514_ /*89777*/;
assign _5512_ = _5513_ | _5515_ /*89774*/;
assign _5521_ = ~D[28] /*89773*/;
assign _5518_ = _4892_ & _5521_ /*89769*/;
assign _5519_ = _4892_ ^ _5521_ /*89772*/;
assign _5520_ = _5512_ & _5519_ /*89770*/;
assign _5341_ = _5512_ ^ _5519_ /*89771*/;
assign _5517_ = _5518_ | _5520_ /*89768*/;
assign _5526_ = ~D[29] /*89767*/;
assign _5523_ = _4893_ & _5526_ /*89763*/;
assign _5524_ = _4893_ ^ _5526_ /*89766*/;
assign _5525_ = _5517_ & _5524_ /*89764*/;
assign _5342_ = _5517_ ^ _5524_ /*89765*/;
assign _5522_ = _5523_ | _5525_ /*89762*/;
assign _5531_ = ~D[30] /*89761*/;
assign _5528_ = _4894_ & _5531_ /*89757*/;
assign _5529_ = _4894_ ^ _5531_ /*89760*/;
assign _5530_ = _5522_ & _5529_ /*89758*/;
assign _5343_ = _5522_ ^ _5529_ /*89759*/;
assign _5527_ = _5528_ | _5530_ /*89756*/;
assign _5536_ = ~D[31] /*89755*/;
assign _5533_ = _4895_ & _5536_ /*89751*/;
assign _5534_ = _4895_ ^ _5536_ /*89754*/;
assign _5535_ = _5527_ & _5534_ /*89752*/;
assign _5344_ = _5527_ ^ _5534_ /*89753*/;
assign _5532_ = _5533_ | _5535_ /*89750*/;
assign _5541_ = ~D[32] /*89749*/;
assign _5538_ = _4896_ & _5541_ /*89745*/;
assign _5539_ = _4896_ ^ _5541_ /*89748*/;
assign _5540_ = _5532_ & _5539_ /*89746*/;
assign _5345_ = _5532_ ^ _5539_ /*89747*/;
assign _5537_ = _5538_ | _5540_ /*89744*/;
assign _5546_ = ~D[33] /*89743*/;
assign _5543_ = _4897_ & _5546_ /*89739*/;
assign _5544_ = _4897_ ^ _5546_ /*89742*/;
assign _5545_ = _5537_ & _5544_ /*89740*/;
assign _5346_ = _5537_ ^ _5544_ /*89741*/;
assign _5542_ = _5543_ | _5545_ /*89738*/;
assign _5551_ = ~D[34] /*89737*/;
assign _5548_ = _4898_ & _5551_ /*89733*/;
assign _5549_ = _4898_ ^ _5551_ /*89736*/;
assign _5550_ = _5542_ & _5549_ /*89734*/;
assign _5347_ = _5542_ ^ _5549_ /*89735*/;
assign _5547_ = _5548_ | _5550_ /*89732*/;
assign _5556_ = ~D[35] /*89731*/;
assign _5553_ = _4899_ & _5556_ /*89727*/;
assign _5554_ = _4899_ ^ _5556_ /*89730*/;
assign _5555_ = _5547_ & _5554_ /*89728*/;
assign _5348_ = _5547_ ^ _5554_ /*89729*/;
assign _5552_ = _5553_ | _5555_ /*89726*/;
assign _5561_ = ~D[36] /*89725*/;
assign _5558_ = _4900_ & _5561_ /*89721*/;
assign _5559_ = _4900_ ^ _5561_ /*89724*/;
assign _5560_ = _5552_ & _5559_ /*89722*/;
assign _5349_ = _5552_ ^ _5559_ /*89723*/;
assign _5557_ = _5558_ | _5560_ /*89720*/;
assign _5566_ = ~D[37] /*89719*/;
assign _5563_ = _4901_ & _5566_ /*89715*/;
assign _5564_ = _4901_ ^ _5566_ /*89718*/;
assign _5565_ = _5557_ & _5564_ /*89716*/;
assign _5350_ = _5557_ ^ _5564_ /*89717*/;
assign _5562_ = _5563_ | _5565_ /*89714*/;
assign _5571_ = ~D[38] /*89713*/;
assign _5568_ = _4902_ & _5571_ /*89709*/;
assign _5569_ = _4902_ ^ _5571_ /*89712*/;
assign _5570_ = _5562_ & _5569_ /*89710*/;
assign _5351_ = _5562_ ^ _5569_ /*89711*/;
assign _5567_ = _5568_ | _5570_ /*89708*/;
assign _5576_ = ~D[39] /*89707*/;
assign _5573_ = _4903_ & _5576_ /*89703*/;
assign _5574_ = _4903_ ^ _5576_ /*89706*/;
assign _5575_ = _5567_ & _5574_ /*89704*/;
assign _5352_ = _5567_ ^ _5574_ /*89705*/;
assign _5572_ = _5573_ | _5575_ /*89702*/;
assign _5581_ = ~D[40] /*89701*/;
assign _5578_ = _4904_ & _5581_ /*89697*/;
assign _5579_ = _4904_ ^ _5581_ /*89700*/;
assign _5580_ = _5572_ & _5579_ /*89698*/;
assign _5353_ = _5572_ ^ _5579_ /*89699*/;
assign _5577_ = _5578_ | _5580_ /*89696*/;
assign _5586_ = ~D[41] /*89695*/;
assign _5583_ = _4905_ & _5586_ /*89691*/;
assign _5584_ = _4905_ ^ _5586_ /*89694*/;
assign _5585_ = _5577_ & _5584_ /*89692*/;
assign _5354_ = _5577_ ^ _5584_ /*89693*/;
assign _5582_ = _5583_ | _5585_ /*89690*/;
assign _5591_ = ~D[42] /*89689*/;
assign _5588_ = _4906_ & _5591_ /*89685*/;
assign _5589_ = _4906_ ^ _5591_ /*89688*/;
assign _5590_ = _5582_ & _5589_ /*89686*/;
assign _5355_ = _5582_ ^ _5589_ /*89687*/;
assign _5587_ = _5588_ | _5590_ /*89684*/;
assign _5596_ = ~D[43] /*89683*/;
assign _5593_ = _4907_ & _5596_ /*89679*/;
assign _5594_ = _4907_ ^ _5596_ /*89682*/;
assign _5595_ = _5587_ & _5594_ /*89680*/;
assign _5356_ = _5587_ ^ _5594_ /*89681*/;
assign _5592_ = _5593_ | _5595_ /*89678*/;
assign _5601_ = ~D[44] /*89677*/;
assign _5598_ = _4908_ & _5601_ /*89673*/;
assign _5599_ = _4908_ ^ _5601_ /*89676*/;
assign _5600_ = _5592_ & _5599_ /*89674*/;
assign _5357_ = _5592_ ^ _5599_ /*89675*/;
assign _5597_ = _5598_ | _5600_ /*89672*/;
assign _5606_ = ~D[45] /*89671*/;
assign _5603_ = _4909_ & _5606_ /*89667*/;
assign _5604_ = _4909_ ^ _5606_ /*89670*/;
assign _5605_ = _5597_ & _5604_ /*89668*/;
assign _5358_ = _5597_ ^ _5604_ /*89669*/;
assign _5602_ = _5603_ | _5605_ /*89666*/;
assign _5611_ = ~D[46] /*89665*/;
assign _5608_ = _4910_ & _5611_ /*89661*/;
assign _5609_ = _4910_ ^ _5611_ /*89664*/;
assign _5610_ = _5602_ & _5609_ /*89662*/;
assign _5359_ = _5602_ ^ _5609_ /*89663*/;
assign _5607_ = _5608_ | _5610_ /*89660*/;
assign _5616_ = ~D[47] /*89659*/;
assign _5613_ = _4911_ & _5616_ /*89655*/;
assign _5614_ = _4911_ ^ _5616_ /*89658*/;
assign _5615_ = _5607_ & _5614_ /*89656*/;
assign _5360_ = _5607_ ^ _5614_ /*89657*/;
assign _5612_ = _5613_ | _5615_ /*89654*/;
assign _5621_ = ~D[48] /*89653*/;
assign _5618_ = _4912_ & _5621_ /*89649*/;
assign _5619_ = _4912_ ^ _5621_ /*89652*/;
assign _5620_ = _5612_ & _5619_ /*89650*/;
assign _5361_ = _5612_ ^ _5619_ /*89651*/;
assign _5617_ = _5618_ | _5620_ /*89648*/;
assign _5626_ = ~D[49] /*89647*/;
assign _5623_ = _4913_ & _5626_ /*89643*/;
assign _5624_ = _4913_ ^ _5626_ /*89646*/;
assign _5625_ = _5617_ & _5624_ /*89644*/;
assign _5362_ = _5617_ ^ _5624_ /*89645*/;
assign _5622_ = _5623_ | _5625_ /*89642*/;
assign _5631_ = ~D[50] /*89641*/;
assign _5628_ = _4914_ & _5631_ /*89637*/;
assign _5629_ = _4914_ ^ _5631_ /*89640*/;
assign _5630_ = _5622_ & _5629_ /*89638*/;
assign _5363_ = _5622_ ^ _5629_ /*89639*/;
assign _5627_ = _5628_ | _5630_ /*89636*/;
assign _5636_ = ~D[51] /*89635*/;
assign _5633_ = _4915_ & _5636_ /*89631*/;
assign _5634_ = _4915_ ^ _5636_ /*89634*/;
assign _5635_ = _5627_ & _5634_ /*89632*/;
assign _5364_ = _5627_ ^ _5634_ /*89633*/;
assign _5632_ = _5633_ | _5635_ /*89630*/;
assign _5641_ = ~D[52] /*89629*/;
assign _5638_ = _4916_ & _5641_ /*89625*/;
assign _5639_ = _4916_ ^ _5641_ /*89628*/;
assign _5640_ = _5632_ & _5639_ /*89626*/;
assign _5365_ = _5632_ ^ _5639_ /*89627*/;
assign _5637_ = _5638_ | _5640_ /*89624*/;
assign _5646_ = ~D[53] /*89623*/;
assign _5643_ = _4917_ & _5646_ /*89619*/;
assign _5644_ = _4917_ ^ _5646_ /*89622*/;
assign _5645_ = _5637_ & _5644_ /*89620*/;
assign _5366_ = _5637_ ^ _5644_ /*89621*/;
assign _5642_ = _5643_ | _5645_ /*89618*/;
assign _5651_ = ~D[54] /*89617*/;
assign _5648_ = _4918_ & _5651_ /*89613*/;
assign _5649_ = _4918_ ^ _5651_ /*89616*/;
assign _5650_ = _5642_ & _5649_ /*89614*/;
assign _5367_ = _5642_ ^ _5649_ /*89615*/;
assign _5647_ = _5648_ | _5650_ /*89612*/;
assign _5656_ = ~D[55] /*89611*/;
assign _5653_ = _4919_ & _5656_ /*89607*/;
assign _5654_ = _4919_ ^ _5656_ /*89610*/;
assign _5655_ = _5647_ & _5654_ /*89608*/;
assign _5368_ = _5647_ ^ _5654_ /*89609*/;
assign _5652_ = _5653_ | _5655_ /*89606*/;
assign _5661_ = ~D[56] /*89605*/;
assign _5658_ = _4920_ & _5661_ /*89601*/;
assign _5659_ = _4920_ ^ _5661_ /*89604*/;
assign _5660_ = _5652_ & _5659_ /*89602*/;
assign _5369_ = _5652_ ^ _5659_ /*89603*/;
assign _5657_ = _5658_ | _5660_ /*89600*/;
assign _5666_ = ~D[57] /*89599*/;
assign _5663_ = _4921_ & _5666_ /*89595*/;
assign _5664_ = _4921_ ^ _5666_ /*89598*/;
assign _5665_ = _5657_ & _5664_ /*89596*/;
assign _5370_ = _5657_ ^ _5664_ /*89597*/;
assign _5662_ = _5663_ | _5665_ /*89594*/;
assign _5671_ = ~D[58] /*89593*/;
assign _5668_ = _4922_ & _5671_ /*89589*/;
assign _5669_ = _4922_ ^ _5671_ /*89592*/;
assign _5670_ = _5662_ & _5669_ /*89590*/;
assign _5371_ = _5662_ ^ _5669_ /*89591*/;
assign _5667_ = _5668_ | _5670_ /*89588*/;
assign _5676_ = ~D[59] /*89587*/;
assign _5673_ = _4923_ & _5676_ /*89583*/;
assign _5674_ = _4923_ ^ _5676_ /*89586*/;
assign _5675_ = _5667_ & _5674_ /*89584*/;
assign _5372_ = _5667_ ^ _5674_ /*89585*/;
assign _5672_ = _5673_ | _5675_ /*89582*/;
assign _5681_ = ~D[60] /*89581*/;
assign _5678_ = _4924_ & _5681_ /*89577*/;
assign _5679_ = _4924_ ^ _5681_ /*89580*/;
assign _5680_ = _5672_ & _5679_ /*89578*/;
assign _5373_ = _5672_ ^ _5679_ /*89579*/;
assign _5677_ = _5678_ | _5680_ /*89576*/;
assign _5686_ = ~D[61] /*89575*/;
assign _5683_ = _4925_ & _5686_ /*89571*/;
assign _5684_ = _4925_ ^ _5686_ /*89574*/;
assign _5685_ = _5677_ & _5684_ /*89572*/;
assign _5374_ = _5677_ ^ _5684_ /*89573*/;
assign _5682_ = _5683_ | _5685_ /*89570*/;
assign _5691_ = ~D[62] /*89569*/;
assign _5688_ = _4926_ & _5691_ /*89565*/;
assign _5689_ = _4926_ ^ _5691_ /*89568*/;
assign _5690_ = _5682_ & _5689_ /*89566*/;
assign _5375_ = _5682_ ^ _5689_ /*89567*/;
assign _5687_ = _5688_ | _5690_ /*89564*/;
assign _5692_ = _4927_ & oneWire /*89559*/;
assign _5693_ = _4927_ ^ oneWire /*89562*/;
assign _5694_ = _5687_ & _5693_ /*89560*/;
assign _5376_ = _5687_ ^ _5693_ /*89561*/;
assign Q[57] = _5692_ | _5694_ /*89558*/;
assign _5827_ = ~Q[57] /*89173*/;
assign _5826_ = _5827_ & D[0] /*89172*/;
assign _5829_ = _5313_ & _5826_ /*89167*/;
assign _5830_ = _5313_ ^ _5826_ /*89170*/;
assign _5831_ = zeroWire & _5830_ /*89168*/;
assign _5761_ = zeroWire ^ _5830_ /*89169*/;
assign _5828_ = _5829_ | _5831_ /*89166*/;
assign _5833_ = ~Q[57] /*89165*/;
assign _5832_ = _5833_ & D[1] /*89164*/;
assign _5835_ = _5314_ & _5832_ /*89159*/;
assign _5836_ = _5314_ ^ _5832_ /*89162*/;
assign _5837_ = _5828_ & _5836_ /*89160*/;
assign _5762_ = _5828_ ^ _5836_ /*89161*/;
assign _5834_ = _5835_ | _5837_ /*89158*/;
assign _5839_ = ~Q[57] /*89157*/;
assign _5838_ = _5839_ & D[2] /*89156*/;
assign _5841_ = _5315_ & _5838_ /*89151*/;
assign _5842_ = _5315_ ^ _5838_ /*89154*/;
assign _5843_ = _5834_ & _5842_ /*89152*/;
assign _5763_ = _5834_ ^ _5842_ /*89153*/;
assign _5840_ = _5841_ | _5843_ /*89150*/;
assign _5845_ = ~Q[57] /*89149*/;
assign _5844_ = _5845_ & D[3] /*89148*/;
assign _5847_ = _5316_ & _5844_ /*89143*/;
assign _5848_ = _5316_ ^ _5844_ /*89146*/;
assign _5849_ = _5840_ & _5848_ /*89144*/;
assign _5764_ = _5840_ ^ _5848_ /*89145*/;
assign _5846_ = _5847_ | _5849_ /*89142*/;
assign _5851_ = ~Q[57] /*89141*/;
assign _5850_ = _5851_ & D[4] /*89140*/;
assign _5853_ = _5317_ & _5850_ /*89135*/;
assign _5854_ = _5317_ ^ _5850_ /*89138*/;
assign _5855_ = _5846_ & _5854_ /*89136*/;
assign _5765_ = _5846_ ^ _5854_ /*89137*/;
assign _5852_ = _5853_ | _5855_ /*89134*/;
assign _5857_ = ~Q[57] /*89133*/;
assign _5856_ = _5857_ & D[5] /*89132*/;
assign _5859_ = _5318_ & _5856_ /*89127*/;
assign _5860_ = _5318_ ^ _5856_ /*89130*/;
assign _5861_ = _5852_ & _5860_ /*89128*/;
assign _5766_ = _5852_ ^ _5860_ /*89129*/;
assign _5858_ = _5859_ | _5861_ /*89126*/;
assign _5863_ = ~Q[57] /*89125*/;
assign _5862_ = _5863_ & D[6] /*89124*/;
assign _5865_ = _5319_ & _5862_ /*89119*/;
assign _5866_ = _5319_ ^ _5862_ /*89122*/;
assign _5867_ = _5858_ & _5866_ /*89120*/;
assign _5767_ = _5858_ ^ _5866_ /*89121*/;
assign _5864_ = _5865_ | _5867_ /*89118*/;
assign _5869_ = ~Q[57] /*89117*/;
assign _5868_ = _5869_ & D[7] /*89116*/;
assign _5871_ = _5320_ & _5868_ /*89111*/;
assign _5872_ = _5320_ ^ _5868_ /*89114*/;
assign _5873_ = _5864_ & _5872_ /*89112*/;
assign _5768_ = _5864_ ^ _5872_ /*89113*/;
assign _5870_ = _5871_ | _5873_ /*89110*/;
assign _5875_ = ~Q[57] /*89109*/;
assign _5874_ = _5875_ & D[8] /*89108*/;
assign _5877_ = _5321_ & _5874_ /*89103*/;
assign _5878_ = _5321_ ^ _5874_ /*89106*/;
assign _5879_ = _5870_ & _5878_ /*89104*/;
assign _5769_ = _5870_ ^ _5878_ /*89105*/;
assign _5876_ = _5877_ | _5879_ /*89102*/;
assign _5881_ = ~Q[57] /*89101*/;
assign _5880_ = _5881_ & D[9] /*89100*/;
assign _5883_ = _5322_ & _5880_ /*89095*/;
assign _5884_ = _5322_ ^ _5880_ /*89098*/;
assign _5885_ = _5876_ & _5884_ /*89096*/;
assign _5770_ = _5876_ ^ _5884_ /*89097*/;
assign _5882_ = _5883_ | _5885_ /*89094*/;
assign _5887_ = ~Q[57] /*89093*/;
assign _5886_ = _5887_ & D[10] /*89092*/;
assign _5889_ = _5323_ & _5886_ /*89087*/;
assign _5890_ = _5323_ ^ _5886_ /*89090*/;
assign _5891_ = _5882_ & _5890_ /*89088*/;
assign _5771_ = _5882_ ^ _5890_ /*89089*/;
assign _5888_ = _5889_ | _5891_ /*89086*/;
assign _5893_ = ~Q[57] /*89085*/;
assign _5892_ = _5893_ & D[11] /*89084*/;
assign _5895_ = _5324_ & _5892_ /*89079*/;
assign _5896_ = _5324_ ^ _5892_ /*89082*/;
assign _5897_ = _5888_ & _5896_ /*89080*/;
assign _5772_ = _5888_ ^ _5896_ /*89081*/;
assign _5894_ = _5895_ | _5897_ /*89078*/;
assign _5899_ = ~Q[57] /*89077*/;
assign _5898_ = _5899_ & D[12] /*89076*/;
assign _5901_ = _5325_ & _5898_ /*89071*/;
assign _5902_ = _5325_ ^ _5898_ /*89074*/;
assign _5903_ = _5894_ & _5902_ /*89072*/;
assign _5773_ = _5894_ ^ _5902_ /*89073*/;
assign _5900_ = _5901_ | _5903_ /*89070*/;
assign _5905_ = ~Q[57] /*89069*/;
assign _5904_ = _5905_ & D[13] /*89068*/;
assign _5907_ = _5326_ & _5904_ /*89063*/;
assign _5908_ = _5326_ ^ _5904_ /*89066*/;
assign _5909_ = _5900_ & _5908_ /*89064*/;
assign _5774_ = _5900_ ^ _5908_ /*89065*/;
assign _5906_ = _5907_ | _5909_ /*89062*/;
assign _5911_ = ~Q[57] /*89061*/;
assign _5910_ = _5911_ & D[14] /*89060*/;
assign _5913_ = _5327_ & _5910_ /*89055*/;
assign _5914_ = _5327_ ^ _5910_ /*89058*/;
assign _5915_ = _5906_ & _5914_ /*89056*/;
assign _5775_ = _5906_ ^ _5914_ /*89057*/;
assign _5912_ = _5913_ | _5915_ /*89054*/;
assign _5917_ = ~Q[57] /*89053*/;
assign _5916_ = _5917_ & D[15] /*89052*/;
assign _5919_ = _5328_ & _5916_ /*89047*/;
assign _5920_ = _5328_ ^ _5916_ /*89050*/;
assign _5921_ = _5912_ & _5920_ /*89048*/;
assign _5776_ = _5912_ ^ _5920_ /*89049*/;
assign _5918_ = _5919_ | _5921_ /*89046*/;
assign _5923_ = ~Q[57] /*89045*/;
assign _5922_ = _5923_ & D[16] /*89044*/;
assign _5925_ = _5329_ & _5922_ /*89039*/;
assign _5926_ = _5329_ ^ _5922_ /*89042*/;
assign _5927_ = _5918_ & _5926_ /*89040*/;
assign _5777_ = _5918_ ^ _5926_ /*89041*/;
assign _5924_ = _5925_ | _5927_ /*89038*/;
assign _5929_ = ~Q[57] /*89037*/;
assign _5928_ = _5929_ & D[17] /*89036*/;
assign _5931_ = _5330_ & _5928_ /*89031*/;
assign _5932_ = _5330_ ^ _5928_ /*89034*/;
assign _5933_ = _5924_ & _5932_ /*89032*/;
assign _5778_ = _5924_ ^ _5932_ /*89033*/;
assign _5930_ = _5931_ | _5933_ /*89030*/;
assign _5935_ = ~Q[57] /*89029*/;
assign _5934_ = _5935_ & D[18] /*89028*/;
assign _5937_ = _5331_ & _5934_ /*89023*/;
assign _5938_ = _5331_ ^ _5934_ /*89026*/;
assign _5939_ = _5930_ & _5938_ /*89024*/;
assign _5779_ = _5930_ ^ _5938_ /*89025*/;
assign _5936_ = _5937_ | _5939_ /*89022*/;
assign _5941_ = ~Q[57] /*89021*/;
assign _5940_ = _5941_ & D[19] /*89020*/;
assign _5943_ = _5332_ & _5940_ /*89015*/;
assign _5944_ = _5332_ ^ _5940_ /*89018*/;
assign _5945_ = _5936_ & _5944_ /*89016*/;
assign _5780_ = _5936_ ^ _5944_ /*89017*/;
assign _5942_ = _5943_ | _5945_ /*89014*/;
assign _5947_ = ~Q[57] /*89013*/;
assign _5946_ = _5947_ & D[20] /*89012*/;
assign _5949_ = _5333_ & _5946_ /*89007*/;
assign _5950_ = _5333_ ^ _5946_ /*89010*/;
assign _5951_ = _5942_ & _5950_ /*89008*/;
assign _5781_ = _5942_ ^ _5950_ /*89009*/;
assign _5948_ = _5949_ | _5951_ /*89006*/;
assign _5953_ = ~Q[57] /*89005*/;
assign _5952_ = _5953_ & D[21] /*89004*/;
assign _5955_ = _5334_ & _5952_ /*88999*/;
assign _5956_ = _5334_ ^ _5952_ /*89002*/;
assign _5957_ = _5948_ & _5956_ /*89000*/;
assign _5782_ = _5948_ ^ _5956_ /*89001*/;
assign _5954_ = _5955_ | _5957_ /*88998*/;
assign _5959_ = ~Q[57] /*88997*/;
assign _5958_ = _5959_ & D[22] /*88996*/;
assign _5961_ = _5335_ & _5958_ /*88991*/;
assign _5962_ = _5335_ ^ _5958_ /*88994*/;
assign _5963_ = _5954_ & _5962_ /*88992*/;
assign _5783_ = _5954_ ^ _5962_ /*88993*/;
assign _5960_ = _5961_ | _5963_ /*88990*/;
assign _5965_ = ~Q[57] /*88989*/;
assign _5964_ = _5965_ & D[23] /*88988*/;
assign _5967_ = _5336_ & _5964_ /*88983*/;
assign _5968_ = _5336_ ^ _5964_ /*88986*/;
assign _5969_ = _5960_ & _5968_ /*88984*/;
assign _5784_ = _5960_ ^ _5968_ /*88985*/;
assign _5966_ = _5967_ | _5969_ /*88982*/;
assign _5971_ = ~Q[57] /*88981*/;
assign _5970_ = _5971_ & D[24] /*88980*/;
assign _5973_ = _5337_ & _5970_ /*88975*/;
assign _5974_ = _5337_ ^ _5970_ /*88978*/;
assign _5975_ = _5966_ & _5974_ /*88976*/;
assign _5785_ = _5966_ ^ _5974_ /*88977*/;
assign _5972_ = _5973_ | _5975_ /*88974*/;
assign _5977_ = ~Q[57] /*88973*/;
assign _5976_ = _5977_ & D[25] /*88972*/;
assign _5979_ = _5338_ & _5976_ /*88967*/;
assign _5980_ = _5338_ ^ _5976_ /*88970*/;
assign _5981_ = _5972_ & _5980_ /*88968*/;
assign _5786_ = _5972_ ^ _5980_ /*88969*/;
assign _5978_ = _5979_ | _5981_ /*88966*/;
assign _5983_ = ~Q[57] /*88965*/;
assign _5982_ = _5983_ & D[26] /*88964*/;
assign _5985_ = _5339_ & _5982_ /*88959*/;
assign _5986_ = _5339_ ^ _5982_ /*88962*/;
assign _5987_ = _5978_ & _5986_ /*88960*/;
assign _5787_ = _5978_ ^ _5986_ /*88961*/;
assign _5984_ = _5985_ | _5987_ /*88958*/;
assign _5989_ = ~Q[57] /*88957*/;
assign _5988_ = _5989_ & D[27] /*88956*/;
assign _5991_ = _5340_ & _5988_ /*88951*/;
assign _5992_ = _5340_ ^ _5988_ /*88954*/;
assign _5993_ = _5984_ & _5992_ /*88952*/;
assign _5788_ = _5984_ ^ _5992_ /*88953*/;
assign _5990_ = _5991_ | _5993_ /*88950*/;
assign _5995_ = ~Q[57] /*88949*/;
assign _5994_ = _5995_ & D[28] /*88948*/;
assign _5997_ = _5341_ & _5994_ /*88943*/;
assign _5998_ = _5341_ ^ _5994_ /*88946*/;
assign _5999_ = _5990_ & _5998_ /*88944*/;
assign _5789_ = _5990_ ^ _5998_ /*88945*/;
assign _5996_ = _5997_ | _5999_ /*88942*/;
assign _6001_ = ~Q[57] /*88941*/;
assign _6000_ = _6001_ & D[29] /*88940*/;
assign _6003_ = _5342_ & _6000_ /*88935*/;
assign _6004_ = _5342_ ^ _6000_ /*88938*/;
assign _6005_ = _5996_ & _6004_ /*88936*/;
assign _5790_ = _5996_ ^ _6004_ /*88937*/;
assign _6002_ = _6003_ | _6005_ /*88934*/;
assign _6007_ = ~Q[57] /*88933*/;
assign _6006_ = _6007_ & D[30] /*88932*/;
assign _6009_ = _5343_ & _6006_ /*88927*/;
assign _6010_ = _5343_ ^ _6006_ /*88930*/;
assign _6011_ = _6002_ & _6010_ /*88928*/;
assign _5791_ = _6002_ ^ _6010_ /*88929*/;
assign _6008_ = _6009_ | _6011_ /*88926*/;
assign _6013_ = ~Q[57] /*88925*/;
assign _6012_ = _6013_ & D[31] /*88924*/;
assign _6015_ = _5344_ & _6012_ /*88919*/;
assign _6016_ = _5344_ ^ _6012_ /*88922*/;
assign _6017_ = _6008_ & _6016_ /*88920*/;
assign _5792_ = _6008_ ^ _6016_ /*88921*/;
assign _6014_ = _6015_ | _6017_ /*88918*/;
assign _6019_ = ~Q[57] /*88917*/;
assign _6018_ = _6019_ & D[32] /*88916*/;
assign _6021_ = _5345_ & _6018_ /*88911*/;
assign _6022_ = _5345_ ^ _6018_ /*88914*/;
assign _6023_ = _6014_ & _6022_ /*88912*/;
assign _5793_ = _6014_ ^ _6022_ /*88913*/;
assign _6020_ = _6021_ | _6023_ /*88910*/;
assign _6025_ = ~Q[57] /*88909*/;
assign _6024_ = _6025_ & D[33] /*88908*/;
assign _6027_ = _5346_ & _6024_ /*88903*/;
assign _6028_ = _5346_ ^ _6024_ /*88906*/;
assign _6029_ = _6020_ & _6028_ /*88904*/;
assign _5794_ = _6020_ ^ _6028_ /*88905*/;
assign _6026_ = _6027_ | _6029_ /*88902*/;
assign _6031_ = ~Q[57] /*88901*/;
assign _6030_ = _6031_ & D[34] /*88900*/;
assign _6033_ = _5347_ & _6030_ /*88895*/;
assign _6034_ = _5347_ ^ _6030_ /*88898*/;
assign _6035_ = _6026_ & _6034_ /*88896*/;
assign _5795_ = _6026_ ^ _6034_ /*88897*/;
assign _6032_ = _6033_ | _6035_ /*88894*/;
assign _6037_ = ~Q[57] /*88893*/;
assign _6036_ = _6037_ & D[35] /*88892*/;
assign _6039_ = _5348_ & _6036_ /*88887*/;
assign _6040_ = _5348_ ^ _6036_ /*88890*/;
assign _6041_ = _6032_ & _6040_ /*88888*/;
assign _5796_ = _6032_ ^ _6040_ /*88889*/;
assign _6038_ = _6039_ | _6041_ /*88886*/;
assign _6043_ = ~Q[57] /*88885*/;
assign _6042_ = _6043_ & D[36] /*88884*/;
assign _6045_ = _5349_ & _6042_ /*88879*/;
assign _6046_ = _5349_ ^ _6042_ /*88882*/;
assign _6047_ = _6038_ & _6046_ /*88880*/;
assign _5797_ = _6038_ ^ _6046_ /*88881*/;
assign _6044_ = _6045_ | _6047_ /*88878*/;
assign _6049_ = ~Q[57] /*88877*/;
assign _6048_ = _6049_ & D[37] /*88876*/;
assign _6051_ = _5350_ & _6048_ /*88871*/;
assign _6052_ = _5350_ ^ _6048_ /*88874*/;
assign _6053_ = _6044_ & _6052_ /*88872*/;
assign _5798_ = _6044_ ^ _6052_ /*88873*/;
assign _6050_ = _6051_ | _6053_ /*88870*/;
assign _6055_ = ~Q[57] /*88869*/;
assign _6054_ = _6055_ & D[38] /*88868*/;
assign _6057_ = _5351_ & _6054_ /*88863*/;
assign _6058_ = _5351_ ^ _6054_ /*88866*/;
assign _6059_ = _6050_ & _6058_ /*88864*/;
assign _5799_ = _6050_ ^ _6058_ /*88865*/;
assign _6056_ = _6057_ | _6059_ /*88862*/;
assign _6061_ = ~Q[57] /*88861*/;
assign _6060_ = _6061_ & D[39] /*88860*/;
assign _6063_ = _5352_ & _6060_ /*88855*/;
assign _6064_ = _5352_ ^ _6060_ /*88858*/;
assign _6065_ = _6056_ & _6064_ /*88856*/;
assign _5800_ = _6056_ ^ _6064_ /*88857*/;
assign _6062_ = _6063_ | _6065_ /*88854*/;
assign _6067_ = ~Q[57] /*88853*/;
assign _6066_ = _6067_ & D[40] /*88852*/;
assign _6069_ = _5353_ & _6066_ /*88847*/;
assign _6070_ = _5353_ ^ _6066_ /*88850*/;
assign _6071_ = _6062_ & _6070_ /*88848*/;
assign _5801_ = _6062_ ^ _6070_ /*88849*/;
assign _6068_ = _6069_ | _6071_ /*88846*/;
assign _6073_ = ~Q[57] /*88845*/;
assign _6072_ = _6073_ & D[41] /*88844*/;
assign _6075_ = _5354_ & _6072_ /*88839*/;
assign _6076_ = _5354_ ^ _6072_ /*88842*/;
assign _6077_ = _6068_ & _6076_ /*88840*/;
assign _5802_ = _6068_ ^ _6076_ /*88841*/;
assign _6074_ = _6075_ | _6077_ /*88838*/;
assign _6079_ = ~Q[57] /*88837*/;
assign _6078_ = _6079_ & D[42] /*88836*/;
assign _6081_ = _5355_ & _6078_ /*88831*/;
assign _6082_ = _5355_ ^ _6078_ /*88834*/;
assign _6083_ = _6074_ & _6082_ /*88832*/;
assign _5803_ = _6074_ ^ _6082_ /*88833*/;
assign _6080_ = _6081_ | _6083_ /*88830*/;
assign _6085_ = ~Q[57] /*88829*/;
assign _6084_ = _6085_ & D[43] /*88828*/;
assign _6087_ = _5356_ & _6084_ /*88823*/;
assign _6088_ = _5356_ ^ _6084_ /*88826*/;
assign _6089_ = _6080_ & _6088_ /*88824*/;
assign _5804_ = _6080_ ^ _6088_ /*88825*/;
assign _6086_ = _6087_ | _6089_ /*88822*/;
assign _6091_ = ~Q[57] /*88821*/;
assign _6090_ = _6091_ & D[44] /*88820*/;
assign _6093_ = _5357_ & _6090_ /*88815*/;
assign _6094_ = _5357_ ^ _6090_ /*88818*/;
assign _6095_ = _6086_ & _6094_ /*88816*/;
assign _5805_ = _6086_ ^ _6094_ /*88817*/;
assign _6092_ = _6093_ | _6095_ /*88814*/;
assign _6097_ = ~Q[57] /*88813*/;
assign _6096_ = _6097_ & D[45] /*88812*/;
assign _6099_ = _5358_ & _6096_ /*88807*/;
assign _6100_ = _5358_ ^ _6096_ /*88810*/;
assign _6101_ = _6092_ & _6100_ /*88808*/;
assign _5806_ = _6092_ ^ _6100_ /*88809*/;
assign _6098_ = _6099_ | _6101_ /*88806*/;
assign _6103_ = ~Q[57] /*88805*/;
assign _6102_ = _6103_ & D[46] /*88804*/;
assign _6105_ = _5359_ & _6102_ /*88799*/;
assign _6106_ = _5359_ ^ _6102_ /*88802*/;
assign _6107_ = _6098_ & _6106_ /*88800*/;
assign _5807_ = _6098_ ^ _6106_ /*88801*/;
assign _6104_ = _6105_ | _6107_ /*88798*/;
assign _6109_ = ~Q[57] /*88797*/;
assign _6108_ = _6109_ & D[47] /*88796*/;
assign _6111_ = _5360_ & _6108_ /*88791*/;
assign _6112_ = _5360_ ^ _6108_ /*88794*/;
assign _6113_ = _6104_ & _6112_ /*88792*/;
assign _5808_ = _6104_ ^ _6112_ /*88793*/;
assign _6110_ = _6111_ | _6113_ /*88790*/;
assign _6115_ = ~Q[57] /*88789*/;
assign _6114_ = _6115_ & D[48] /*88788*/;
assign _6117_ = _5361_ & _6114_ /*88783*/;
assign _6118_ = _5361_ ^ _6114_ /*88786*/;
assign _6119_ = _6110_ & _6118_ /*88784*/;
assign _5809_ = _6110_ ^ _6118_ /*88785*/;
assign _6116_ = _6117_ | _6119_ /*88782*/;
assign _6121_ = ~Q[57] /*88781*/;
assign _6120_ = _6121_ & D[49] /*88780*/;
assign _6123_ = _5362_ & _6120_ /*88775*/;
assign _6124_ = _5362_ ^ _6120_ /*88778*/;
assign _6125_ = _6116_ & _6124_ /*88776*/;
assign _5810_ = _6116_ ^ _6124_ /*88777*/;
assign _6122_ = _6123_ | _6125_ /*88774*/;
assign _6127_ = ~Q[57] /*88773*/;
assign _6126_ = _6127_ & D[50] /*88772*/;
assign _6129_ = _5363_ & _6126_ /*88767*/;
assign _6130_ = _5363_ ^ _6126_ /*88770*/;
assign _6131_ = _6122_ & _6130_ /*88768*/;
assign _5811_ = _6122_ ^ _6130_ /*88769*/;
assign _6128_ = _6129_ | _6131_ /*88766*/;
assign _6133_ = ~Q[57] /*88765*/;
assign _6132_ = _6133_ & D[51] /*88764*/;
assign _6135_ = _5364_ & _6132_ /*88759*/;
assign _6136_ = _5364_ ^ _6132_ /*88762*/;
assign _6137_ = _6128_ & _6136_ /*88760*/;
assign _5812_ = _6128_ ^ _6136_ /*88761*/;
assign _6134_ = _6135_ | _6137_ /*88758*/;
assign _6139_ = ~Q[57] /*88757*/;
assign _6138_ = _6139_ & D[52] /*88756*/;
assign _6141_ = _5365_ & _6138_ /*88751*/;
assign _6142_ = _5365_ ^ _6138_ /*88754*/;
assign _6143_ = _6134_ & _6142_ /*88752*/;
assign _5813_ = _6134_ ^ _6142_ /*88753*/;
assign _6140_ = _6141_ | _6143_ /*88750*/;
assign _6145_ = ~Q[57] /*88749*/;
assign _6144_ = _6145_ & D[53] /*88748*/;
assign _6147_ = _5366_ & _6144_ /*88743*/;
assign _6148_ = _5366_ ^ _6144_ /*88746*/;
assign _6149_ = _6140_ & _6148_ /*88744*/;
assign _5814_ = _6140_ ^ _6148_ /*88745*/;
assign _6146_ = _6147_ | _6149_ /*88742*/;
assign _6151_ = ~Q[57] /*88741*/;
assign _6150_ = _6151_ & D[54] /*88740*/;
assign _6153_ = _5367_ & _6150_ /*88735*/;
assign _6154_ = _5367_ ^ _6150_ /*88738*/;
assign _6155_ = _6146_ & _6154_ /*88736*/;
assign _5815_ = _6146_ ^ _6154_ /*88737*/;
assign _6152_ = _6153_ | _6155_ /*88734*/;
assign _6157_ = ~Q[57] /*88733*/;
assign _6156_ = _6157_ & D[55] /*88732*/;
assign _6159_ = _5368_ & _6156_ /*88727*/;
assign _6160_ = _5368_ ^ _6156_ /*88730*/;
assign _6161_ = _6152_ & _6160_ /*88728*/;
assign _5816_ = _6152_ ^ _6160_ /*88729*/;
assign _6158_ = _6159_ | _6161_ /*88726*/;
assign _6163_ = ~Q[57] /*88725*/;
assign _6162_ = _6163_ & D[56] /*88724*/;
assign _6165_ = _5369_ & _6162_ /*88719*/;
assign _6166_ = _5369_ ^ _6162_ /*88722*/;
assign _6167_ = _6158_ & _6166_ /*88720*/;
assign _5817_ = _6158_ ^ _6166_ /*88721*/;
assign _6164_ = _6165_ | _6167_ /*88718*/;
assign _6169_ = ~Q[57] /*88717*/;
assign _6168_ = _6169_ & D[57] /*88716*/;
assign _6171_ = _5370_ & _6168_ /*88711*/;
assign _6172_ = _5370_ ^ _6168_ /*88714*/;
assign _6173_ = _6164_ & _6172_ /*88712*/;
assign _5818_ = _6164_ ^ _6172_ /*88713*/;
assign _6170_ = _6171_ | _6173_ /*88710*/;
assign _6175_ = ~Q[57] /*88709*/;
assign _6174_ = _6175_ & D[58] /*88708*/;
assign _6177_ = _5371_ & _6174_ /*88703*/;
assign _6178_ = _5371_ ^ _6174_ /*88706*/;
assign _6179_ = _6170_ & _6178_ /*88704*/;
assign _5819_ = _6170_ ^ _6178_ /*88705*/;
assign _6176_ = _6177_ | _6179_ /*88702*/;
assign _6181_ = ~Q[57] /*88701*/;
assign _6180_ = _6181_ & D[59] /*88700*/;
assign _6183_ = _5372_ & _6180_ /*88695*/;
assign _6184_ = _5372_ ^ _6180_ /*88698*/;
assign _6185_ = _6176_ & _6184_ /*88696*/;
assign _5820_ = _6176_ ^ _6184_ /*88697*/;
assign _6182_ = _6183_ | _6185_ /*88694*/;
assign _6187_ = ~Q[57] /*88693*/;
assign _6186_ = _6187_ & D[60] /*88692*/;
assign _6189_ = _5373_ & _6186_ /*88687*/;
assign _6190_ = _5373_ ^ _6186_ /*88690*/;
assign _6191_ = _6182_ & _6190_ /*88688*/;
assign _5821_ = _6182_ ^ _6190_ /*88689*/;
assign _6188_ = _6189_ | _6191_ /*88686*/;
assign _6193_ = ~Q[57] /*88685*/;
assign _6192_ = _6193_ & D[61] /*88684*/;
assign _6195_ = _5374_ & _6192_ /*88679*/;
assign _6196_ = _5374_ ^ _6192_ /*88682*/;
assign _6197_ = _6188_ & _6196_ /*88680*/;
assign _5822_ = _6188_ ^ _6196_ /*88681*/;
assign _6194_ = _6195_ | _6197_ /*88678*/;
assign _6199_ = ~Q[57] /*88677*/;
assign _6198_ = _6199_ & D[62] /*88676*/;
assign _6201_ = _5375_ & _6198_ /*88671*/;
assign _6202_ = _5375_ ^ _6198_ /*88674*/;
assign _6203_ = _6194_ & _6202_ /*88672*/;
assign _5823_ = _6194_ ^ _6202_ /*88673*/;
assign _6200_ = _6201_ | _6203_ /*88670*/;
assign _6205_ = ~Q[57] /*88669*/;
assign _6204_ = _6205_ & zeroWire /*88668*/;
assign _6206_ = _5376_ ^ _6204_ /*88666*/;
assign _5824_ = _6206_ ^ _6200_ /*88665*/;
assign _6277_ = ~D[0] /*88411*/;
assign _6274_ = R_0[56] & _6277_ /*88407*/;
assign _6275_ = R_0[56] ^ _6277_ /*88410*/;
assign _6276_ = oneWire & _6275_ /*88408*/;
assign _6209_ = oneWire ^ _6275_ /*88409*/;
assign _6273_ = _6274_ | _6276_ /*88406*/;
assign _6282_ = ~D[1] /*88405*/;
assign _6279_ = _5761_ & _6282_ /*88401*/;
assign _6280_ = _5761_ ^ _6282_ /*88404*/;
assign _6281_ = _6273_ & _6280_ /*88402*/;
assign _6210_ = _6273_ ^ _6280_ /*88403*/;
assign _6278_ = _6279_ | _6281_ /*88400*/;
assign _6287_ = ~D[2] /*88399*/;
assign _6284_ = _5762_ & _6287_ /*88395*/;
assign _6285_ = _5762_ ^ _6287_ /*88398*/;
assign _6286_ = _6278_ & _6285_ /*88396*/;
assign _6211_ = _6278_ ^ _6285_ /*88397*/;
assign _6283_ = _6284_ | _6286_ /*88394*/;
assign _6292_ = ~D[3] /*88393*/;
assign _6289_ = _5763_ & _6292_ /*88389*/;
assign _6290_ = _5763_ ^ _6292_ /*88392*/;
assign _6291_ = _6283_ & _6290_ /*88390*/;
assign _6212_ = _6283_ ^ _6290_ /*88391*/;
assign _6288_ = _6289_ | _6291_ /*88388*/;
assign _6297_ = ~D[4] /*88387*/;
assign _6294_ = _5764_ & _6297_ /*88383*/;
assign _6295_ = _5764_ ^ _6297_ /*88386*/;
assign _6296_ = _6288_ & _6295_ /*88384*/;
assign _6213_ = _6288_ ^ _6295_ /*88385*/;
assign _6293_ = _6294_ | _6296_ /*88382*/;
assign _6302_ = ~D[5] /*88381*/;
assign _6299_ = _5765_ & _6302_ /*88377*/;
assign _6300_ = _5765_ ^ _6302_ /*88380*/;
assign _6301_ = _6293_ & _6300_ /*88378*/;
assign _6214_ = _6293_ ^ _6300_ /*88379*/;
assign _6298_ = _6299_ | _6301_ /*88376*/;
assign _6307_ = ~D[6] /*88375*/;
assign _6304_ = _5766_ & _6307_ /*88371*/;
assign _6305_ = _5766_ ^ _6307_ /*88374*/;
assign _6306_ = _6298_ & _6305_ /*88372*/;
assign _6215_ = _6298_ ^ _6305_ /*88373*/;
assign _6303_ = _6304_ | _6306_ /*88370*/;
assign _6312_ = ~D[7] /*88369*/;
assign _6309_ = _5767_ & _6312_ /*88365*/;
assign _6310_ = _5767_ ^ _6312_ /*88368*/;
assign _6311_ = _6303_ & _6310_ /*88366*/;
assign _6216_ = _6303_ ^ _6310_ /*88367*/;
assign _6308_ = _6309_ | _6311_ /*88364*/;
assign _6317_ = ~D[8] /*88363*/;
assign _6314_ = _5768_ & _6317_ /*88359*/;
assign _6315_ = _5768_ ^ _6317_ /*88362*/;
assign _6316_ = _6308_ & _6315_ /*88360*/;
assign _6217_ = _6308_ ^ _6315_ /*88361*/;
assign _6313_ = _6314_ | _6316_ /*88358*/;
assign _6322_ = ~D[9] /*88357*/;
assign _6319_ = _5769_ & _6322_ /*88353*/;
assign _6320_ = _5769_ ^ _6322_ /*88356*/;
assign _6321_ = _6313_ & _6320_ /*88354*/;
assign _6218_ = _6313_ ^ _6320_ /*88355*/;
assign _6318_ = _6319_ | _6321_ /*88352*/;
assign _6327_ = ~D[10] /*88351*/;
assign _6324_ = _5770_ & _6327_ /*88347*/;
assign _6325_ = _5770_ ^ _6327_ /*88350*/;
assign _6326_ = _6318_ & _6325_ /*88348*/;
assign _6219_ = _6318_ ^ _6325_ /*88349*/;
assign _6323_ = _6324_ | _6326_ /*88346*/;
assign _6332_ = ~D[11] /*88345*/;
assign _6329_ = _5771_ & _6332_ /*88341*/;
assign _6330_ = _5771_ ^ _6332_ /*88344*/;
assign _6331_ = _6323_ & _6330_ /*88342*/;
assign _6220_ = _6323_ ^ _6330_ /*88343*/;
assign _6328_ = _6329_ | _6331_ /*88340*/;
assign _6337_ = ~D[12] /*88339*/;
assign _6334_ = _5772_ & _6337_ /*88335*/;
assign _6335_ = _5772_ ^ _6337_ /*88338*/;
assign _6336_ = _6328_ & _6335_ /*88336*/;
assign _6221_ = _6328_ ^ _6335_ /*88337*/;
assign _6333_ = _6334_ | _6336_ /*88334*/;
assign _6342_ = ~D[13] /*88333*/;
assign _6339_ = _5773_ & _6342_ /*88329*/;
assign _6340_ = _5773_ ^ _6342_ /*88332*/;
assign _6341_ = _6333_ & _6340_ /*88330*/;
assign _6222_ = _6333_ ^ _6340_ /*88331*/;
assign _6338_ = _6339_ | _6341_ /*88328*/;
assign _6347_ = ~D[14] /*88327*/;
assign _6344_ = _5774_ & _6347_ /*88323*/;
assign _6345_ = _5774_ ^ _6347_ /*88326*/;
assign _6346_ = _6338_ & _6345_ /*88324*/;
assign _6223_ = _6338_ ^ _6345_ /*88325*/;
assign _6343_ = _6344_ | _6346_ /*88322*/;
assign _6352_ = ~D[15] /*88321*/;
assign _6349_ = _5775_ & _6352_ /*88317*/;
assign _6350_ = _5775_ ^ _6352_ /*88320*/;
assign _6351_ = _6343_ & _6350_ /*88318*/;
assign _6224_ = _6343_ ^ _6350_ /*88319*/;
assign _6348_ = _6349_ | _6351_ /*88316*/;
assign _6357_ = ~D[16] /*88315*/;
assign _6354_ = _5776_ & _6357_ /*88311*/;
assign _6355_ = _5776_ ^ _6357_ /*88314*/;
assign _6356_ = _6348_ & _6355_ /*88312*/;
assign _6225_ = _6348_ ^ _6355_ /*88313*/;
assign _6353_ = _6354_ | _6356_ /*88310*/;
assign _6362_ = ~D[17] /*88309*/;
assign _6359_ = _5777_ & _6362_ /*88305*/;
assign _6360_ = _5777_ ^ _6362_ /*88308*/;
assign _6361_ = _6353_ & _6360_ /*88306*/;
assign _6226_ = _6353_ ^ _6360_ /*88307*/;
assign _6358_ = _6359_ | _6361_ /*88304*/;
assign _6367_ = ~D[18] /*88303*/;
assign _6364_ = _5778_ & _6367_ /*88299*/;
assign _6365_ = _5778_ ^ _6367_ /*88302*/;
assign _6366_ = _6358_ & _6365_ /*88300*/;
assign _6227_ = _6358_ ^ _6365_ /*88301*/;
assign _6363_ = _6364_ | _6366_ /*88298*/;
assign _6372_ = ~D[19] /*88297*/;
assign _6369_ = _5779_ & _6372_ /*88293*/;
assign _6370_ = _5779_ ^ _6372_ /*88296*/;
assign _6371_ = _6363_ & _6370_ /*88294*/;
assign _6228_ = _6363_ ^ _6370_ /*88295*/;
assign _6368_ = _6369_ | _6371_ /*88292*/;
assign _6377_ = ~D[20] /*88291*/;
assign _6374_ = _5780_ & _6377_ /*88287*/;
assign _6375_ = _5780_ ^ _6377_ /*88290*/;
assign _6376_ = _6368_ & _6375_ /*88288*/;
assign _6229_ = _6368_ ^ _6375_ /*88289*/;
assign _6373_ = _6374_ | _6376_ /*88286*/;
assign _6382_ = ~D[21] /*88285*/;
assign _6379_ = _5781_ & _6382_ /*88281*/;
assign _6380_ = _5781_ ^ _6382_ /*88284*/;
assign _6381_ = _6373_ & _6380_ /*88282*/;
assign _6230_ = _6373_ ^ _6380_ /*88283*/;
assign _6378_ = _6379_ | _6381_ /*88280*/;
assign _6387_ = ~D[22] /*88279*/;
assign _6384_ = _5782_ & _6387_ /*88275*/;
assign _6385_ = _5782_ ^ _6387_ /*88278*/;
assign _6386_ = _6378_ & _6385_ /*88276*/;
assign _6231_ = _6378_ ^ _6385_ /*88277*/;
assign _6383_ = _6384_ | _6386_ /*88274*/;
assign _6392_ = ~D[23] /*88273*/;
assign _6389_ = _5783_ & _6392_ /*88269*/;
assign _6390_ = _5783_ ^ _6392_ /*88272*/;
assign _6391_ = _6383_ & _6390_ /*88270*/;
assign _6232_ = _6383_ ^ _6390_ /*88271*/;
assign _6388_ = _6389_ | _6391_ /*88268*/;
assign _6397_ = ~D[24] /*88267*/;
assign _6394_ = _5784_ & _6397_ /*88263*/;
assign _6395_ = _5784_ ^ _6397_ /*88266*/;
assign _6396_ = _6388_ & _6395_ /*88264*/;
assign _6233_ = _6388_ ^ _6395_ /*88265*/;
assign _6393_ = _6394_ | _6396_ /*88262*/;
assign _6402_ = ~D[25] /*88261*/;
assign _6399_ = _5785_ & _6402_ /*88257*/;
assign _6400_ = _5785_ ^ _6402_ /*88260*/;
assign _6401_ = _6393_ & _6400_ /*88258*/;
assign _6234_ = _6393_ ^ _6400_ /*88259*/;
assign _6398_ = _6399_ | _6401_ /*88256*/;
assign _6407_ = ~D[26] /*88255*/;
assign _6404_ = _5786_ & _6407_ /*88251*/;
assign _6405_ = _5786_ ^ _6407_ /*88254*/;
assign _6406_ = _6398_ & _6405_ /*88252*/;
assign _6235_ = _6398_ ^ _6405_ /*88253*/;
assign _6403_ = _6404_ | _6406_ /*88250*/;
assign _6412_ = ~D[27] /*88249*/;
assign _6409_ = _5787_ & _6412_ /*88245*/;
assign _6410_ = _5787_ ^ _6412_ /*88248*/;
assign _6411_ = _6403_ & _6410_ /*88246*/;
assign _6236_ = _6403_ ^ _6410_ /*88247*/;
assign _6408_ = _6409_ | _6411_ /*88244*/;
assign _6417_ = ~D[28] /*88243*/;
assign _6414_ = _5788_ & _6417_ /*88239*/;
assign _6415_ = _5788_ ^ _6417_ /*88242*/;
assign _6416_ = _6408_ & _6415_ /*88240*/;
assign _6237_ = _6408_ ^ _6415_ /*88241*/;
assign _6413_ = _6414_ | _6416_ /*88238*/;
assign _6422_ = ~D[29] /*88237*/;
assign _6419_ = _5789_ & _6422_ /*88233*/;
assign _6420_ = _5789_ ^ _6422_ /*88236*/;
assign _6421_ = _6413_ & _6420_ /*88234*/;
assign _6238_ = _6413_ ^ _6420_ /*88235*/;
assign _6418_ = _6419_ | _6421_ /*88232*/;
assign _6427_ = ~D[30] /*88231*/;
assign _6424_ = _5790_ & _6427_ /*88227*/;
assign _6425_ = _5790_ ^ _6427_ /*88230*/;
assign _6426_ = _6418_ & _6425_ /*88228*/;
assign _6239_ = _6418_ ^ _6425_ /*88229*/;
assign _6423_ = _6424_ | _6426_ /*88226*/;
assign _6432_ = ~D[31] /*88225*/;
assign _6429_ = _5791_ & _6432_ /*88221*/;
assign _6430_ = _5791_ ^ _6432_ /*88224*/;
assign _6431_ = _6423_ & _6430_ /*88222*/;
assign _6240_ = _6423_ ^ _6430_ /*88223*/;
assign _6428_ = _6429_ | _6431_ /*88220*/;
assign _6437_ = ~D[32] /*88219*/;
assign _6434_ = _5792_ & _6437_ /*88215*/;
assign _6435_ = _5792_ ^ _6437_ /*88218*/;
assign _6436_ = _6428_ & _6435_ /*88216*/;
assign _6241_ = _6428_ ^ _6435_ /*88217*/;
assign _6433_ = _6434_ | _6436_ /*88214*/;
assign _6442_ = ~D[33] /*88213*/;
assign _6439_ = _5793_ & _6442_ /*88209*/;
assign _6440_ = _5793_ ^ _6442_ /*88212*/;
assign _6441_ = _6433_ & _6440_ /*88210*/;
assign _6242_ = _6433_ ^ _6440_ /*88211*/;
assign _6438_ = _6439_ | _6441_ /*88208*/;
assign _6447_ = ~D[34] /*88207*/;
assign _6444_ = _5794_ & _6447_ /*88203*/;
assign _6445_ = _5794_ ^ _6447_ /*88206*/;
assign _6446_ = _6438_ & _6445_ /*88204*/;
assign _6243_ = _6438_ ^ _6445_ /*88205*/;
assign _6443_ = _6444_ | _6446_ /*88202*/;
assign _6452_ = ~D[35] /*88201*/;
assign _6449_ = _5795_ & _6452_ /*88197*/;
assign _6450_ = _5795_ ^ _6452_ /*88200*/;
assign _6451_ = _6443_ & _6450_ /*88198*/;
assign _6244_ = _6443_ ^ _6450_ /*88199*/;
assign _6448_ = _6449_ | _6451_ /*88196*/;
assign _6457_ = ~D[36] /*88195*/;
assign _6454_ = _5796_ & _6457_ /*88191*/;
assign _6455_ = _5796_ ^ _6457_ /*88194*/;
assign _6456_ = _6448_ & _6455_ /*88192*/;
assign _6245_ = _6448_ ^ _6455_ /*88193*/;
assign _6453_ = _6454_ | _6456_ /*88190*/;
assign _6462_ = ~D[37] /*88189*/;
assign _6459_ = _5797_ & _6462_ /*88185*/;
assign _6460_ = _5797_ ^ _6462_ /*88188*/;
assign _6461_ = _6453_ & _6460_ /*88186*/;
assign _6246_ = _6453_ ^ _6460_ /*88187*/;
assign _6458_ = _6459_ | _6461_ /*88184*/;
assign _6467_ = ~D[38] /*88183*/;
assign _6464_ = _5798_ & _6467_ /*88179*/;
assign _6465_ = _5798_ ^ _6467_ /*88182*/;
assign _6466_ = _6458_ & _6465_ /*88180*/;
assign _6247_ = _6458_ ^ _6465_ /*88181*/;
assign _6463_ = _6464_ | _6466_ /*88178*/;
assign _6472_ = ~D[39] /*88177*/;
assign _6469_ = _5799_ & _6472_ /*88173*/;
assign _6470_ = _5799_ ^ _6472_ /*88176*/;
assign _6471_ = _6463_ & _6470_ /*88174*/;
assign _6248_ = _6463_ ^ _6470_ /*88175*/;
assign _6468_ = _6469_ | _6471_ /*88172*/;
assign _6477_ = ~D[40] /*88171*/;
assign _6474_ = _5800_ & _6477_ /*88167*/;
assign _6475_ = _5800_ ^ _6477_ /*88170*/;
assign _6476_ = _6468_ & _6475_ /*88168*/;
assign _6249_ = _6468_ ^ _6475_ /*88169*/;
assign _6473_ = _6474_ | _6476_ /*88166*/;
assign _6482_ = ~D[41] /*88165*/;
assign _6479_ = _5801_ & _6482_ /*88161*/;
assign _6480_ = _5801_ ^ _6482_ /*88164*/;
assign _6481_ = _6473_ & _6480_ /*88162*/;
assign _6250_ = _6473_ ^ _6480_ /*88163*/;
assign _6478_ = _6479_ | _6481_ /*88160*/;
assign _6487_ = ~D[42] /*88159*/;
assign _6484_ = _5802_ & _6487_ /*88155*/;
assign _6485_ = _5802_ ^ _6487_ /*88158*/;
assign _6486_ = _6478_ & _6485_ /*88156*/;
assign _6251_ = _6478_ ^ _6485_ /*88157*/;
assign _6483_ = _6484_ | _6486_ /*88154*/;
assign _6492_ = ~D[43] /*88153*/;
assign _6489_ = _5803_ & _6492_ /*88149*/;
assign _6490_ = _5803_ ^ _6492_ /*88152*/;
assign _6491_ = _6483_ & _6490_ /*88150*/;
assign _6252_ = _6483_ ^ _6490_ /*88151*/;
assign _6488_ = _6489_ | _6491_ /*88148*/;
assign _6497_ = ~D[44] /*88147*/;
assign _6494_ = _5804_ & _6497_ /*88143*/;
assign _6495_ = _5804_ ^ _6497_ /*88146*/;
assign _6496_ = _6488_ & _6495_ /*88144*/;
assign _6253_ = _6488_ ^ _6495_ /*88145*/;
assign _6493_ = _6494_ | _6496_ /*88142*/;
assign _6502_ = ~D[45] /*88141*/;
assign _6499_ = _5805_ & _6502_ /*88137*/;
assign _6500_ = _5805_ ^ _6502_ /*88140*/;
assign _6501_ = _6493_ & _6500_ /*88138*/;
assign _6254_ = _6493_ ^ _6500_ /*88139*/;
assign _6498_ = _6499_ | _6501_ /*88136*/;
assign _6507_ = ~D[46] /*88135*/;
assign _6504_ = _5806_ & _6507_ /*88131*/;
assign _6505_ = _5806_ ^ _6507_ /*88134*/;
assign _6506_ = _6498_ & _6505_ /*88132*/;
assign _6255_ = _6498_ ^ _6505_ /*88133*/;
assign _6503_ = _6504_ | _6506_ /*88130*/;
assign _6512_ = ~D[47] /*88129*/;
assign _6509_ = _5807_ & _6512_ /*88125*/;
assign _6510_ = _5807_ ^ _6512_ /*88128*/;
assign _6511_ = _6503_ & _6510_ /*88126*/;
assign _6256_ = _6503_ ^ _6510_ /*88127*/;
assign _6508_ = _6509_ | _6511_ /*88124*/;
assign _6517_ = ~D[48] /*88123*/;
assign _6514_ = _5808_ & _6517_ /*88119*/;
assign _6515_ = _5808_ ^ _6517_ /*88122*/;
assign _6516_ = _6508_ & _6515_ /*88120*/;
assign _6257_ = _6508_ ^ _6515_ /*88121*/;
assign _6513_ = _6514_ | _6516_ /*88118*/;
assign _6522_ = ~D[49] /*88117*/;
assign _6519_ = _5809_ & _6522_ /*88113*/;
assign _6520_ = _5809_ ^ _6522_ /*88116*/;
assign _6521_ = _6513_ & _6520_ /*88114*/;
assign _6258_ = _6513_ ^ _6520_ /*88115*/;
assign _6518_ = _6519_ | _6521_ /*88112*/;
assign _6527_ = ~D[50] /*88111*/;
assign _6524_ = _5810_ & _6527_ /*88107*/;
assign _6525_ = _5810_ ^ _6527_ /*88110*/;
assign _6526_ = _6518_ & _6525_ /*88108*/;
assign _6259_ = _6518_ ^ _6525_ /*88109*/;
assign _6523_ = _6524_ | _6526_ /*88106*/;
assign _6532_ = ~D[51] /*88105*/;
assign _6529_ = _5811_ & _6532_ /*88101*/;
assign _6530_ = _5811_ ^ _6532_ /*88104*/;
assign _6531_ = _6523_ & _6530_ /*88102*/;
assign _6260_ = _6523_ ^ _6530_ /*88103*/;
assign _6528_ = _6529_ | _6531_ /*88100*/;
assign _6537_ = ~D[52] /*88099*/;
assign _6534_ = _5812_ & _6537_ /*88095*/;
assign _6535_ = _5812_ ^ _6537_ /*88098*/;
assign _6536_ = _6528_ & _6535_ /*88096*/;
assign _6261_ = _6528_ ^ _6535_ /*88097*/;
assign _6533_ = _6534_ | _6536_ /*88094*/;
assign _6542_ = ~D[53] /*88093*/;
assign _6539_ = _5813_ & _6542_ /*88089*/;
assign _6540_ = _5813_ ^ _6542_ /*88092*/;
assign _6541_ = _6533_ & _6540_ /*88090*/;
assign _6262_ = _6533_ ^ _6540_ /*88091*/;
assign _6538_ = _6539_ | _6541_ /*88088*/;
assign _6547_ = ~D[54] /*88087*/;
assign _6544_ = _5814_ & _6547_ /*88083*/;
assign _6545_ = _5814_ ^ _6547_ /*88086*/;
assign _6546_ = _6538_ & _6545_ /*88084*/;
assign _6263_ = _6538_ ^ _6545_ /*88085*/;
assign _6543_ = _6544_ | _6546_ /*88082*/;
assign _6552_ = ~D[55] /*88081*/;
assign _6549_ = _5815_ & _6552_ /*88077*/;
assign _6550_ = _5815_ ^ _6552_ /*88080*/;
assign _6551_ = _6543_ & _6550_ /*88078*/;
assign _6264_ = _6543_ ^ _6550_ /*88079*/;
assign _6548_ = _6549_ | _6551_ /*88076*/;
assign _6557_ = ~D[56] /*88075*/;
assign _6554_ = _5816_ & _6557_ /*88071*/;
assign _6555_ = _5816_ ^ _6557_ /*88074*/;
assign _6556_ = _6548_ & _6555_ /*88072*/;
assign _6265_ = _6548_ ^ _6555_ /*88073*/;
assign _6553_ = _6554_ | _6556_ /*88070*/;
assign _6562_ = ~D[57] /*88069*/;
assign _6559_ = _5817_ & _6562_ /*88065*/;
assign _6560_ = _5817_ ^ _6562_ /*88068*/;
assign _6561_ = _6553_ & _6560_ /*88066*/;
assign _6266_ = _6553_ ^ _6560_ /*88067*/;
assign _6558_ = _6559_ | _6561_ /*88064*/;
assign _6567_ = ~D[58] /*88063*/;
assign _6564_ = _5818_ & _6567_ /*88059*/;
assign _6565_ = _5818_ ^ _6567_ /*88062*/;
assign _6566_ = _6558_ & _6565_ /*88060*/;
assign _6267_ = _6558_ ^ _6565_ /*88061*/;
assign _6563_ = _6564_ | _6566_ /*88058*/;
assign _6572_ = ~D[59] /*88057*/;
assign _6569_ = _5819_ & _6572_ /*88053*/;
assign _6570_ = _5819_ ^ _6572_ /*88056*/;
assign _6571_ = _6563_ & _6570_ /*88054*/;
assign _6268_ = _6563_ ^ _6570_ /*88055*/;
assign _6568_ = _6569_ | _6571_ /*88052*/;
assign _6577_ = ~D[60] /*88051*/;
assign _6574_ = _5820_ & _6577_ /*88047*/;
assign _6575_ = _5820_ ^ _6577_ /*88050*/;
assign _6576_ = _6568_ & _6575_ /*88048*/;
assign _6269_ = _6568_ ^ _6575_ /*88049*/;
assign _6573_ = _6574_ | _6576_ /*88046*/;
assign _6582_ = ~D[61] /*88045*/;
assign _6579_ = _5821_ & _6582_ /*88041*/;
assign _6580_ = _5821_ ^ _6582_ /*88044*/;
assign _6581_ = _6573_ & _6580_ /*88042*/;
assign _6270_ = _6573_ ^ _6580_ /*88043*/;
assign _6578_ = _6579_ | _6581_ /*88040*/;
assign _6587_ = ~D[62] /*88039*/;
assign _6584_ = _5822_ & _6587_ /*88035*/;
assign _6585_ = _5822_ ^ _6587_ /*88038*/;
assign _6586_ = _6578_ & _6585_ /*88036*/;
assign _6271_ = _6578_ ^ _6585_ /*88037*/;
assign _6583_ = _6584_ | _6586_ /*88034*/;
assign _6588_ = _5823_ & oneWire /*88029*/;
assign _6589_ = _5823_ ^ oneWire /*88032*/;
assign _6590_ = _6583_ & _6589_ /*88030*/;
assign _6272_ = _6583_ ^ _6589_ /*88031*/;
assign Q[56] = _6588_ | _6590_ /*88028*/;
assign _6723_ = ~Q[56] /*87643*/;
assign _6722_ = _6723_ & D[0] /*87642*/;
assign _6725_ = _6209_ & _6722_ /*87637*/;
assign _6726_ = _6209_ ^ _6722_ /*87640*/;
assign _6727_ = zeroWire & _6726_ /*87638*/;
assign _6657_ = zeroWire ^ _6726_ /*87639*/;
assign _6724_ = _6725_ | _6727_ /*87636*/;
assign _6729_ = ~Q[56] /*87635*/;
assign _6728_ = _6729_ & D[1] /*87634*/;
assign _6731_ = _6210_ & _6728_ /*87629*/;
assign _6732_ = _6210_ ^ _6728_ /*87632*/;
assign _6733_ = _6724_ & _6732_ /*87630*/;
assign _6658_ = _6724_ ^ _6732_ /*87631*/;
assign _6730_ = _6731_ | _6733_ /*87628*/;
assign _6735_ = ~Q[56] /*87627*/;
assign _6734_ = _6735_ & D[2] /*87626*/;
assign _6737_ = _6211_ & _6734_ /*87621*/;
assign _6738_ = _6211_ ^ _6734_ /*87624*/;
assign _6739_ = _6730_ & _6738_ /*87622*/;
assign _6659_ = _6730_ ^ _6738_ /*87623*/;
assign _6736_ = _6737_ | _6739_ /*87620*/;
assign _6741_ = ~Q[56] /*87619*/;
assign _6740_ = _6741_ & D[3] /*87618*/;
assign _6743_ = _6212_ & _6740_ /*87613*/;
assign _6744_ = _6212_ ^ _6740_ /*87616*/;
assign _6745_ = _6736_ & _6744_ /*87614*/;
assign _6660_ = _6736_ ^ _6744_ /*87615*/;
assign _6742_ = _6743_ | _6745_ /*87612*/;
assign _6747_ = ~Q[56] /*87611*/;
assign _6746_ = _6747_ & D[4] /*87610*/;
assign _6749_ = _6213_ & _6746_ /*87605*/;
assign _6750_ = _6213_ ^ _6746_ /*87608*/;
assign _6751_ = _6742_ & _6750_ /*87606*/;
assign _6661_ = _6742_ ^ _6750_ /*87607*/;
assign _6748_ = _6749_ | _6751_ /*87604*/;
assign _6753_ = ~Q[56] /*87603*/;
assign _6752_ = _6753_ & D[5] /*87602*/;
assign _6755_ = _6214_ & _6752_ /*87597*/;
assign _6756_ = _6214_ ^ _6752_ /*87600*/;
assign _6757_ = _6748_ & _6756_ /*87598*/;
assign _6662_ = _6748_ ^ _6756_ /*87599*/;
assign _6754_ = _6755_ | _6757_ /*87596*/;
assign _6759_ = ~Q[56] /*87595*/;
assign _6758_ = _6759_ & D[6] /*87594*/;
assign _6761_ = _6215_ & _6758_ /*87589*/;
assign _6762_ = _6215_ ^ _6758_ /*87592*/;
assign _6763_ = _6754_ & _6762_ /*87590*/;
assign _6663_ = _6754_ ^ _6762_ /*87591*/;
assign _6760_ = _6761_ | _6763_ /*87588*/;
assign _6765_ = ~Q[56] /*87587*/;
assign _6764_ = _6765_ & D[7] /*87586*/;
assign _6767_ = _6216_ & _6764_ /*87581*/;
assign _6768_ = _6216_ ^ _6764_ /*87584*/;
assign _6769_ = _6760_ & _6768_ /*87582*/;
assign _6664_ = _6760_ ^ _6768_ /*87583*/;
assign _6766_ = _6767_ | _6769_ /*87580*/;
assign _6771_ = ~Q[56] /*87579*/;
assign _6770_ = _6771_ & D[8] /*87578*/;
assign _6773_ = _6217_ & _6770_ /*87573*/;
assign _6774_ = _6217_ ^ _6770_ /*87576*/;
assign _6775_ = _6766_ & _6774_ /*87574*/;
assign _6665_ = _6766_ ^ _6774_ /*87575*/;
assign _6772_ = _6773_ | _6775_ /*87572*/;
assign _6777_ = ~Q[56] /*87571*/;
assign _6776_ = _6777_ & D[9] /*87570*/;
assign _6779_ = _6218_ & _6776_ /*87565*/;
assign _6780_ = _6218_ ^ _6776_ /*87568*/;
assign _6781_ = _6772_ & _6780_ /*87566*/;
assign _6666_ = _6772_ ^ _6780_ /*87567*/;
assign _6778_ = _6779_ | _6781_ /*87564*/;
assign _6783_ = ~Q[56] /*87563*/;
assign _6782_ = _6783_ & D[10] /*87562*/;
assign _6785_ = _6219_ & _6782_ /*87557*/;
assign _6786_ = _6219_ ^ _6782_ /*87560*/;
assign _6787_ = _6778_ & _6786_ /*87558*/;
assign _6667_ = _6778_ ^ _6786_ /*87559*/;
assign _6784_ = _6785_ | _6787_ /*87556*/;
assign _6789_ = ~Q[56] /*87555*/;
assign _6788_ = _6789_ & D[11] /*87554*/;
assign _6791_ = _6220_ & _6788_ /*87549*/;
assign _6792_ = _6220_ ^ _6788_ /*87552*/;
assign _6793_ = _6784_ & _6792_ /*87550*/;
assign _6668_ = _6784_ ^ _6792_ /*87551*/;
assign _6790_ = _6791_ | _6793_ /*87548*/;
assign _6795_ = ~Q[56] /*87547*/;
assign _6794_ = _6795_ & D[12] /*87546*/;
assign _6797_ = _6221_ & _6794_ /*87541*/;
assign _6798_ = _6221_ ^ _6794_ /*87544*/;
assign _6799_ = _6790_ & _6798_ /*87542*/;
assign _6669_ = _6790_ ^ _6798_ /*87543*/;
assign _6796_ = _6797_ | _6799_ /*87540*/;
assign _6801_ = ~Q[56] /*87539*/;
assign _6800_ = _6801_ & D[13] /*87538*/;
assign _6803_ = _6222_ & _6800_ /*87533*/;
assign _6804_ = _6222_ ^ _6800_ /*87536*/;
assign _6805_ = _6796_ & _6804_ /*87534*/;
assign _6670_ = _6796_ ^ _6804_ /*87535*/;
assign _6802_ = _6803_ | _6805_ /*87532*/;
assign _6807_ = ~Q[56] /*87531*/;
assign _6806_ = _6807_ & D[14] /*87530*/;
assign _6809_ = _6223_ & _6806_ /*87525*/;
assign _6810_ = _6223_ ^ _6806_ /*87528*/;
assign _6811_ = _6802_ & _6810_ /*87526*/;
assign _6671_ = _6802_ ^ _6810_ /*87527*/;
assign _6808_ = _6809_ | _6811_ /*87524*/;
assign _6813_ = ~Q[56] /*87523*/;
assign _6812_ = _6813_ & D[15] /*87522*/;
assign _6815_ = _6224_ & _6812_ /*87517*/;
assign _6816_ = _6224_ ^ _6812_ /*87520*/;
assign _6817_ = _6808_ & _6816_ /*87518*/;
assign _6672_ = _6808_ ^ _6816_ /*87519*/;
assign _6814_ = _6815_ | _6817_ /*87516*/;
assign _6819_ = ~Q[56] /*87515*/;
assign _6818_ = _6819_ & D[16] /*87514*/;
assign _6821_ = _6225_ & _6818_ /*87509*/;
assign _6822_ = _6225_ ^ _6818_ /*87512*/;
assign _6823_ = _6814_ & _6822_ /*87510*/;
assign _6673_ = _6814_ ^ _6822_ /*87511*/;
assign _6820_ = _6821_ | _6823_ /*87508*/;
assign _6825_ = ~Q[56] /*87507*/;
assign _6824_ = _6825_ & D[17] /*87506*/;
assign _6827_ = _6226_ & _6824_ /*87501*/;
assign _6828_ = _6226_ ^ _6824_ /*87504*/;
assign _6829_ = _6820_ & _6828_ /*87502*/;
assign _6674_ = _6820_ ^ _6828_ /*87503*/;
assign _6826_ = _6827_ | _6829_ /*87500*/;
assign _6831_ = ~Q[56] /*87499*/;
assign _6830_ = _6831_ & D[18] /*87498*/;
assign _6833_ = _6227_ & _6830_ /*87493*/;
assign _6834_ = _6227_ ^ _6830_ /*87496*/;
assign _6835_ = _6826_ & _6834_ /*87494*/;
assign _6675_ = _6826_ ^ _6834_ /*87495*/;
assign _6832_ = _6833_ | _6835_ /*87492*/;
assign _6837_ = ~Q[56] /*87491*/;
assign _6836_ = _6837_ & D[19] /*87490*/;
assign _6839_ = _6228_ & _6836_ /*87485*/;
assign _6840_ = _6228_ ^ _6836_ /*87488*/;
assign _6841_ = _6832_ & _6840_ /*87486*/;
assign _6676_ = _6832_ ^ _6840_ /*87487*/;
assign _6838_ = _6839_ | _6841_ /*87484*/;
assign _6843_ = ~Q[56] /*87483*/;
assign _6842_ = _6843_ & D[20] /*87482*/;
assign _6845_ = _6229_ & _6842_ /*87477*/;
assign _6846_ = _6229_ ^ _6842_ /*87480*/;
assign _6847_ = _6838_ & _6846_ /*87478*/;
assign _6677_ = _6838_ ^ _6846_ /*87479*/;
assign _6844_ = _6845_ | _6847_ /*87476*/;
assign _6849_ = ~Q[56] /*87475*/;
assign _6848_ = _6849_ & D[21] /*87474*/;
assign _6851_ = _6230_ & _6848_ /*87469*/;
assign _6852_ = _6230_ ^ _6848_ /*87472*/;
assign _6853_ = _6844_ & _6852_ /*87470*/;
assign _6678_ = _6844_ ^ _6852_ /*87471*/;
assign _6850_ = _6851_ | _6853_ /*87468*/;
assign _6855_ = ~Q[56] /*87467*/;
assign _6854_ = _6855_ & D[22] /*87466*/;
assign _6857_ = _6231_ & _6854_ /*87461*/;
assign _6858_ = _6231_ ^ _6854_ /*87464*/;
assign _6859_ = _6850_ & _6858_ /*87462*/;
assign _6679_ = _6850_ ^ _6858_ /*87463*/;
assign _6856_ = _6857_ | _6859_ /*87460*/;
assign _6861_ = ~Q[56] /*87459*/;
assign _6860_ = _6861_ & D[23] /*87458*/;
assign _6863_ = _6232_ & _6860_ /*87453*/;
assign _6864_ = _6232_ ^ _6860_ /*87456*/;
assign _6865_ = _6856_ & _6864_ /*87454*/;
assign _6680_ = _6856_ ^ _6864_ /*87455*/;
assign _6862_ = _6863_ | _6865_ /*87452*/;
assign _6867_ = ~Q[56] /*87451*/;
assign _6866_ = _6867_ & D[24] /*87450*/;
assign _6869_ = _6233_ & _6866_ /*87445*/;
assign _6870_ = _6233_ ^ _6866_ /*87448*/;
assign _6871_ = _6862_ & _6870_ /*87446*/;
assign _6681_ = _6862_ ^ _6870_ /*87447*/;
assign _6868_ = _6869_ | _6871_ /*87444*/;
assign _6873_ = ~Q[56] /*87443*/;
assign _6872_ = _6873_ & D[25] /*87442*/;
assign _6875_ = _6234_ & _6872_ /*87437*/;
assign _6876_ = _6234_ ^ _6872_ /*87440*/;
assign _6877_ = _6868_ & _6876_ /*87438*/;
assign _6682_ = _6868_ ^ _6876_ /*87439*/;
assign _6874_ = _6875_ | _6877_ /*87436*/;
assign _6879_ = ~Q[56] /*87435*/;
assign _6878_ = _6879_ & D[26] /*87434*/;
assign _6881_ = _6235_ & _6878_ /*87429*/;
assign _6882_ = _6235_ ^ _6878_ /*87432*/;
assign _6883_ = _6874_ & _6882_ /*87430*/;
assign _6683_ = _6874_ ^ _6882_ /*87431*/;
assign _6880_ = _6881_ | _6883_ /*87428*/;
assign _6885_ = ~Q[56] /*87427*/;
assign _6884_ = _6885_ & D[27] /*87426*/;
assign _6887_ = _6236_ & _6884_ /*87421*/;
assign _6888_ = _6236_ ^ _6884_ /*87424*/;
assign _6889_ = _6880_ & _6888_ /*87422*/;
assign _6684_ = _6880_ ^ _6888_ /*87423*/;
assign _6886_ = _6887_ | _6889_ /*87420*/;
assign _6891_ = ~Q[56] /*87419*/;
assign _6890_ = _6891_ & D[28] /*87418*/;
assign _6893_ = _6237_ & _6890_ /*87413*/;
assign _6894_ = _6237_ ^ _6890_ /*87416*/;
assign _6895_ = _6886_ & _6894_ /*87414*/;
assign _6685_ = _6886_ ^ _6894_ /*87415*/;
assign _6892_ = _6893_ | _6895_ /*87412*/;
assign _6897_ = ~Q[56] /*87411*/;
assign _6896_ = _6897_ & D[29] /*87410*/;
assign _6899_ = _6238_ & _6896_ /*87405*/;
assign _6900_ = _6238_ ^ _6896_ /*87408*/;
assign _6901_ = _6892_ & _6900_ /*87406*/;
assign _6686_ = _6892_ ^ _6900_ /*87407*/;
assign _6898_ = _6899_ | _6901_ /*87404*/;
assign _6903_ = ~Q[56] /*87403*/;
assign _6902_ = _6903_ & D[30] /*87402*/;
assign _6905_ = _6239_ & _6902_ /*87397*/;
assign _6906_ = _6239_ ^ _6902_ /*87400*/;
assign _6907_ = _6898_ & _6906_ /*87398*/;
assign _6687_ = _6898_ ^ _6906_ /*87399*/;
assign _6904_ = _6905_ | _6907_ /*87396*/;
assign _6909_ = ~Q[56] /*87395*/;
assign _6908_ = _6909_ & D[31] /*87394*/;
assign _6911_ = _6240_ & _6908_ /*87389*/;
assign _6912_ = _6240_ ^ _6908_ /*87392*/;
assign _6913_ = _6904_ & _6912_ /*87390*/;
assign _6688_ = _6904_ ^ _6912_ /*87391*/;
assign _6910_ = _6911_ | _6913_ /*87388*/;
assign _6915_ = ~Q[56] /*87387*/;
assign _6914_ = _6915_ & D[32] /*87386*/;
assign _6917_ = _6241_ & _6914_ /*87381*/;
assign _6918_ = _6241_ ^ _6914_ /*87384*/;
assign _6919_ = _6910_ & _6918_ /*87382*/;
assign _6689_ = _6910_ ^ _6918_ /*87383*/;
assign _6916_ = _6917_ | _6919_ /*87380*/;
assign _6921_ = ~Q[56] /*87379*/;
assign _6920_ = _6921_ & D[33] /*87378*/;
assign _6923_ = _6242_ & _6920_ /*87373*/;
assign _6924_ = _6242_ ^ _6920_ /*87376*/;
assign _6925_ = _6916_ & _6924_ /*87374*/;
assign _6690_ = _6916_ ^ _6924_ /*87375*/;
assign _6922_ = _6923_ | _6925_ /*87372*/;
assign _6927_ = ~Q[56] /*87371*/;
assign _6926_ = _6927_ & D[34] /*87370*/;
assign _6929_ = _6243_ & _6926_ /*87365*/;
assign _6930_ = _6243_ ^ _6926_ /*87368*/;
assign _6931_ = _6922_ & _6930_ /*87366*/;
assign _6691_ = _6922_ ^ _6930_ /*87367*/;
assign _6928_ = _6929_ | _6931_ /*87364*/;
assign _6933_ = ~Q[56] /*87363*/;
assign _6932_ = _6933_ & D[35] /*87362*/;
assign _6935_ = _6244_ & _6932_ /*87357*/;
assign _6936_ = _6244_ ^ _6932_ /*87360*/;
assign _6937_ = _6928_ & _6936_ /*87358*/;
assign _6692_ = _6928_ ^ _6936_ /*87359*/;
assign _6934_ = _6935_ | _6937_ /*87356*/;
assign _6939_ = ~Q[56] /*87355*/;
assign _6938_ = _6939_ & D[36] /*87354*/;
assign _6941_ = _6245_ & _6938_ /*87349*/;
assign _6942_ = _6245_ ^ _6938_ /*87352*/;
assign _6943_ = _6934_ & _6942_ /*87350*/;
assign _6693_ = _6934_ ^ _6942_ /*87351*/;
assign _6940_ = _6941_ | _6943_ /*87348*/;
assign _6945_ = ~Q[56] /*87347*/;
assign _6944_ = _6945_ & D[37] /*87346*/;
assign _6947_ = _6246_ & _6944_ /*87341*/;
assign _6948_ = _6246_ ^ _6944_ /*87344*/;
assign _6949_ = _6940_ & _6948_ /*87342*/;
assign _6694_ = _6940_ ^ _6948_ /*87343*/;
assign _6946_ = _6947_ | _6949_ /*87340*/;
assign _6951_ = ~Q[56] /*87339*/;
assign _6950_ = _6951_ & D[38] /*87338*/;
assign _6953_ = _6247_ & _6950_ /*87333*/;
assign _6954_ = _6247_ ^ _6950_ /*87336*/;
assign _6955_ = _6946_ & _6954_ /*87334*/;
assign _6695_ = _6946_ ^ _6954_ /*87335*/;
assign _6952_ = _6953_ | _6955_ /*87332*/;
assign _6957_ = ~Q[56] /*87331*/;
assign _6956_ = _6957_ & D[39] /*87330*/;
assign _6959_ = _6248_ & _6956_ /*87325*/;
assign _6960_ = _6248_ ^ _6956_ /*87328*/;
assign _6961_ = _6952_ & _6960_ /*87326*/;
assign _6696_ = _6952_ ^ _6960_ /*87327*/;
assign _6958_ = _6959_ | _6961_ /*87324*/;
assign _6963_ = ~Q[56] /*87323*/;
assign _6962_ = _6963_ & D[40] /*87322*/;
assign _6965_ = _6249_ & _6962_ /*87317*/;
assign _6966_ = _6249_ ^ _6962_ /*87320*/;
assign _6967_ = _6958_ & _6966_ /*87318*/;
assign _6697_ = _6958_ ^ _6966_ /*87319*/;
assign _6964_ = _6965_ | _6967_ /*87316*/;
assign _6969_ = ~Q[56] /*87315*/;
assign _6968_ = _6969_ & D[41] /*87314*/;
assign _6971_ = _6250_ & _6968_ /*87309*/;
assign _6972_ = _6250_ ^ _6968_ /*87312*/;
assign _6973_ = _6964_ & _6972_ /*87310*/;
assign _6698_ = _6964_ ^ _6972_ /*87311*/;
assign _6970_ = _6971_ | _6973_ /*87308*/;
assign _6975_ = ~Q[56] /*87307*/;
assign _6974_ = _6975_ & D[42] /*87306*/;
assign _6977_ = _6251_ & _6974_ /*87301*/;
assign _6978_ = _6251_ ^ _6974_ /*87304*/;
assign _6979_ = _6970_ & _6978_ /*87302*/;
assign _6699_ = _6970_ ^ _6978_ /*87303*/;
assign _6976_ = _6977_ | _6979_ /*87300*/;
assign _6981_ = ~Q[56] /*87299*/;
assign _6980_ = _6981_ & D[43] /*87298*/;
assign _6983_ = _6252_ & _6980_ /*87293*/;
assign _6984_ = _6252_ ^ _6980_ /*87296*/;
assign _6985_ = _6976_ & _6984_ /*87294*/;
assign _6700_ = _6976_ ^ _6984_ /*87295*/;
assign _6982_ = _6983_ | _6985_ /*87292*/;
assign _6987_ = ~Q[56] /*87291*/;
assign _6986_ = _6987_ & D[44] /*87290*/;
assign _6989_ = _6253_ & _6986_ /*87285*/;
assign _6990_ = _6253_ ^ _6986_ /*87288*/;
assign _6991_ = _6982_ & _6990_ /*87286*/;
assign _6701_ = _6982_ ^ _6990_ /*87287*/;
assign _6988_ = _6989_ | _6991_ /*87284*/;
assign _6993_ = ~Q[56] /*87283*/;
assign _6992_ = _6993_ & D[45] /*87282*/;
assign _6995_ = _6254_ & _6992_ /*87277*/;
assign _6996_ = _6254_ ^ _6992_ /*87280*/;
assign _6997_ = _6988_ & _6996_ /*87278*/;
assign _6702_ = _6988_ ^ _6996_ /*87279*/;
assign _6994_ = _6995_ | _6997_ /*87276*/;
assign _6999_ = ~Q[56] /*87275*/;
assign _6998_ = _6999_ & D[46] /*87274*/;
assign _7001_ = _6255_ & _6998_ /*87269*/;
assign _7002_ = _6255_ ^ _6998_ /*87272*/;
assign _7003_ = _6994_ & _7002_ /*87270*/;
assign _6703_ = _6994_ ^ _7002_ /*87271*/;
assign _7000_ = _7001_ | _7003_ /*87268*/;
assign _7005_ = ~Q[56] /*87267*/;
assign _7004_ = _7005_ & D[47] /*87266*/;
assign _7007_ = _6256_ & _7004_ /*87261*/;
assign _7008_ = _6256_ ^ _7004_ /*87264*/;
assign _7009_ = _7000_ & _7008_ /*87262*/;
assign _6704_ = _7000_ ^ _7008_ /*87263*/;
assign _7006_ = _7007_ | _7009_ /*87260*/;
assign _7011_ = ~Q[56] /*87259*/;
assign _7010_ = _7011_ & D[48] /*87258*/;
assign _7013_ = _6257_ & _7010_ /*87253*/;
assign _7014_ = _6257_ ^ _7010_ /*87256*/;
assign _7015_ = _7006_ & _7014_ /*87254*/;
assign _6705_ = _7006_ ^ _7014_ /*87255*/;
assign _7012_ = _7013_ | _7015_ /*87252*/;
assign _7017_ = ~Q[56] /*87251*/;
assign _7016_ = _7017_ & D[49] /*87250*/;
assign _7019_ = _6258_ & _7016_ /*87245*/;
assign _7020_ = _6258_ ^ _7016_ /*87248*/;
assign _7021_ = _7012_ & _7020_ /*87246*/;
assign _6706_ = _7012_ ^ _7020_ /*87247*/;
assign _7018_ = _7019_ | _7021_ /*87244*/;
assign _7023_ = ~Q[56] /*87243*/;
assign _7022_ = _7023_ & D[50] /*87242*/;
assign _7025_ = _6259_ & _7022_ /*87237*/;
assign _7026_ = _6259_ ^ _7022_ /*87240*/;
assign _7027_ = _7018_ & _7026_ /*87238*/;
assign _6707_ = _7018_ ^ _7026_ /*87239*/;
assign _7024_ = _7025_ | _7027_ /*87236*/;
assign _7029_ = ~Q[56] /*87235*/;
assign _7028_ = _7029_ & D[51] /*87234*/;
assign _7031_ = _6260_ & _7028_ /*87229*/;
assign _7032_ = _6260_ ^ _7028_ /*87232*/;
assign _7033_ = _7024_ & _7032_ /*87230*/;
assign _6708_ = _7024_ ^ _7032_ /*87231*/;
assign _7030_ = _7031_ | _7033_ /*87228*/;
assign _7035_ = ~Q[56] /*87227*/;
assign _7034_ = _7035_ & D[52] /*87226*/;
assign _7037_ = _6261_ & _7034_ /*87221*/;
assign _7038_ = _6261_ ^ _7034_ /*87224*/;
assign _7039_ = _7030_ & _7038_ /*87222*/;
assign _6709_ = _7030_ ^ _7038_ /*87223*/;
assign _7036_ = _7037_ | _7039_ /*87220*/;
assign _7041_ = ~Q[56] /*87219*/;
assign _7040_ = _7041_ & D[53] /*87218*/;
assign _7043_ = _6262_ & _7040_ /*87213*/;
assign _7044_ = _6262_ ^ _7040_ /*87216*/;
assign _7045_ = _7036_ & _7044_ /*87214*/;
assign _6710_ = _7036_ ^ _7044_ /*87215*/;
assign _7042_ = _7043_ | _7045_ /*87212*/;
assign _7047_ = ~Q[56] /*87211*/;
assign _7046_ = _7047_ & D[54] /*87210*/;
assign _7049_ = _6263_ & _7046_ /*87205*/;
assign _7050_ = _6263_ ^ _7046_ /*87208*/;
assign _7051_ = _7042_ & _7050_ /*87206*/;
assign _6711_ = _7042_ ^ _7050_ /*87207*/;
assign _7048_ = _7049_ | _7051_ /*87204*/;
assign _7053_ = ~Q[56] /*87203*/;
assign _7052_ = _7053_ & D[55] /*87202*/;
assign _7055_ = _6264_ & _7052_ /*87197*/;
assign _7056_ = _6264_ ^ _7052_ /*87200*/;
assign _7057_ = _7048_ & _7056_ /*87198*/;
assign _6712_ = _7048_ ^ _7056_ /*87199*/;
assign _7054_ = _7055_ | _7057_ /*87196*/;
assign _7059_ = ~Q[56] /*87195*/;
assign _7058_ = _7059_ & D[56] /*87194*/;
assign _7061_ = _6265_ & _7058_ /*87189*/;
assign _7062_ = _6265_ ^ _7058_ /*87192*/;
assign _7063_ = _7054_ & _7062_ /*87190*/;
assign _6713_ = _7054_ ^ _7062_ /*87191*/;
assign _7060_ = _7061_ | _7063_ /*87188*/;
assign _7065_ = ~Q[56] /*87187*/;
assign _7064_ = _7065_ & D[57] /*87186*/;
assign _7067_ = _6266_ & _7064_ /*87181*/;
assign _7068_ = _6266_ ^ _7064_ /*87184*/;
assign _7069_ = _7060_ & _7068_ /*87182*/;
assign _6714_ = _7060_ ^ _7068_ /*87183*/;
assign _7066_ = _7067_ | _7069_ /*87180*/;
assign _7071_ = ~Q[56] /*87179*/;
assign _7070_ = _7071_ & D[58] /*87178*/;
assign _7073_ = _6267_ & _7070_ /*87173*/;
assign _7074_ = _6267_ ^ _7070_ /*87176*/;
assign _7075_ = _7066_ & _7074_ /*87174*/;
assign _6715_ = _7066_ ^ _7074_ /*87175*/;
assign _7072_ = _7073_ | _7075_ /*87172*/;
assign _7077_ = ~Q[56] /*87171*/;
assign _7076_ = _7077_ & D[59] /*87170*/;
assign _7079_ = _6268_ & _7076_ /*87165*/;
assign _7080_ = _6268_ ^ _7076_ /*87168*/;
assign _7081_ = _7072_ & _7080_ /*87166*/;
assign _6716_ = _7072_ ^ _7080_ /*87167*/;
assign _7078_ = _7079_ | _7081_ /*87164*/;
assign _7083_ = ~Q[56] /*87163*/;
assign _7082_ = _7083_ & D[60] /*87162*/;
assign _7085_ = _6269_ & _7082_ /*87157*/;
assign _7086_ = _6269_ ^ _7082_ /*87160*/;
assign _7087_ = _7078_ & _7086_ /*87158*/;
assign _6717_ = _7078_ ^ _7086_ /*87159*/;
assign _7084_ = _7085_ | _7087_ /*87156*/;
assign _7089_ = ~Q[56] /*87155*/;
assign _7088_ = _7089_ & D[61] /*87154*/;
assign _7091_ = _6270_ & _7088_ /*87149*/;
assign _7092_ = _6270_ ^ _7088_ /*87152*/;
assign _7093_ = _7084_ & _7092_ /*87150*/;
assign _6718_ = _7084_ ^ _7092_ /*87151*/;
assign _7090_ = _7091_ | _7093_ /*87148*/;
assign _7095_ = ~Q[56] /*87147*/;
assign _7094_ = _7095_ & D[62] /*87146*/;
assign _7097_ = _6271_ & _7094_ /*87141*/;
assign _7098_ = _6271_ ^ _7094_ /*87144*/;
assign _7099_ = _7090_ & _7098_ /*87142*/;
assign _6719_ = _7090_ ^ _7098_ /*87143*/;
assign _7096_ = _7097_ | _7099_ /*87140*/;
assign _7101_ = ~Q[56] /*87139*/;
assign _7100_ = _7101_ & zeroWire /*87138*/;
assign _7102_ = _6272_ ^ _7100_ /*87136*/;
assign _6720_ = _7102_ ^ _7096_ /*87135*/;
assign _7173_ = ~D[0] /*86881*/;
assign _7170_ = R_0[55] & _7173_ /*86877*/;
assign _7171_ = R_0[55] ^ _7173_ /*86880*/;
assign _7172_ = oneWire & _7171_ /*86878*/;
assign _7105_ = oneWire ^ _7171_ /*86879*/;
assign _7169_ = _7170_ | _7172_ /*86876*/;
assign _7178_ = ~D[1] /*86875*/;
assign _7175_ = _6657_ & _7178_ /*86871*/;
assign _7176_ = _6657_ ^ _7178_ /*86874*/;
assign _7177_ = _7169_ & _7176_ /*86872*/;
assign _7106_ = _7169_ ^ _7176_ /*86873*/;
assign _7174_ = _7175_ | _7177_ /*86870*/;
assign _7183_ = ~D[2] /*86869*/;
assign _7180_ = _6658_ & _7183_ /*86865*/;
assign _7181_ = _6658_ ^ _7183_ /*86868*/;
assign _7182_ = _7174_ & _7181_ /*86866*/;
assign _7107_ = _7174_ ^ _7181_ /*86867*/;
assign _7179_ = _7180_ | _7182_ /*86864*/;
assign _7188_ = ~D[3] /*86863*/;
assign _7185_ = _6659_ & _7188_ /*86859*/;
assign _7186_ = _6659_ ^ _7188_ /*86862*/;
assign _7187_ = _7179_ & _7186_ /*86860*/;
assign _7108_ = _7179_ ^ _7186_ /*86861*/;
assign _7184_ = _7185_ | _7187_ /*86858*/;
assign _7193_ = ~D[4] /*86857*/;
assign _7190_ = _6660_ & _7193_ /*86853*/;
assign _7191_ = _6660_ ^ _7193_ /*86856*/;
assign _7192_ = _7184_ & _7191_ /*86854*/;
assign _7109_ = _7184_ ^ _7191_ /*86855*/;
assign _7189_ = _7190_ | _7192_ /*86852*/;
assign _7198_ = ~D[5] /*86851*/;
assign _7195_ = _6661_ & _7198_ /*86847*/;
assign _7196_ = _6661_ ^ _7198_ /*86850*/;
assign _7197_ = _7189_ & _7196_ /*86848*/;
assign _7110_ = _7189_ ^ _7196_ /*86849*/;
assign _7194_ = _7195_ | _7197_ /*86846*/;
assign _7203_ = ~D[6] /*86845*/;
assign _7200_ = _6662_ & _7203_ /*86841*/;
assign _7201_ = _6662_ ^ _7203_ /*86844*/;
assign _7202_ = _7194_ & _7201_ /*86842*/;
assign _7111_ = _7194_ ^ _7201_ /*86843*/;
assign _7199_ = _7200_ | _7202_ /*86840*/;
assign _7208_ = ~D[7] /*86839*/;
assign _7205_ = _6663_ & _7208_ /*86835*/;
assign _7206_ = _6663_ ^ _7208_ /*86838*/;
assign _7207_ = _7199_ & _7206_ /*86836*/;
assign _7112_ = _7199_ ^ _7206_ /*86837*/;
assign _7204_ = _7205_ | _7207_ /*86834*/;
assign _7213_ = ~D[8] /*86833*/;
assign _7210_ = _6664_ & _7213_ /*86829*/;
assign _7211_ = _6664_ ^ _7213_ /*86832*/;
assign _7212_ = _7204_ & _7211_ /*86830*/;
assign _7113_ = _7204_ ^ _7211_ /*86831*/;
assign _7209_ = _7210_ | _7212_ /*86828*/;
assign _7218_ = ~D[9] /*86827*/;
assign _7215_ = _6665_ & _7218_ /*86823*/;
assign _7216_ = _6665_ ^ _7218_ /*86826*/;
assign _7217_ = _7209_ & _7216_ /*86824*/;
assign _7114_ = _7209_ ^ _7216_ /*86825*/;
assign _7214_ = _7215_ | _7217_ /*86822*/;
assign _7223_ = ~D[10] /*86821*/;
assign _7220_ = _6666_ & _7223_ /*86817*/;
assign _7221_ = _6666_ ^ _7223_ /*86820*/;
assign _7222_ = _7214_ & _7221_ /*86818*/;
assign _7115_ = _7214_ ^ _7221_ /*86819*/;
assign _7219_ = _7220_ | _7222_ /*86816*/;
assign _7228_ = ~D[11] /*86815*/;
assign _7225_ = _6667_ & _7228_ /*86811*/;
assign _7226_ = _6667_ ^ _7228_ /*86814*/;
assign _7227_ = _7219_ & _7226_ /*86812*/;
assign _7116_ = _7219_ ^ _7226_ /*86813*/;
assign _7224_ = _7225_ | _7227_ /*86810*/;
assign _7233_ = ~D[12] /*86809*/;
assign _7230_ = _6668_ & _7233_ /*86805*/;
assign _7231_ = _6668_ ^ _7233_ /*86808*/;
assign _7232_ = _7224_ & _7231_ /*86806*/;
assign _7117_ = _7224_ ^ _7231_ /*86807*/;
assign _7229_ = _7230_ | _7232_ /*86804*/;
assign _7238_ = ~D[13] /*86803*/;
assign _7235_ = _6669_ & _7238_ /*86799*/;
assign _7236_ = _6669_ ^ _7238_ /*86802*/;
assign _7237_ = _7229_ & _7236_ /*86800*/;
assign _7118_ = _7229_ ^ _7236_ /*86801*/;
assign _7234_ = _7235_ | _7237_ /*86798*/;
assign _7243_ = ~D[14] /*86797*/;
assign _7240_ = _6670_ & _7243_ /*86793*/;
assign _7241_ = _6670_ ^ _7243_ /*86796*/;
assign _7242_ = _7234_ & _7241_ /*86794*/;
assign _7119_ = _7234_ ^ _7241_ /*86795*/;
assign _7239_ = _7240_ | _7242_ /*86792*/;
assign _7248_ = ~D[15] /*86791*/;
assign _7245_ = _6671_ & _7248_ /*86787*/;
assign _7246_ = _6671_ ^ _7248_ /*86790*/;
assign _7247_ = _7239_ & _7246_ /*86788*/;
assign _7120_ = _7239_ ^ _7246_ /*86789*/;
assign _7244_ = _7245_ | _7247_ /*86786*/;
assign _7253_ = ~D[16] /*86785*/;
assign _7250_ = _6672_ & _7253_ /*86781*/;
assign _7251_ = _6672_ ^ _7253_ /*86784*/;
assign _7252_ = _7244_ & _7251_ /*86782*/;
assign _7121_ = _7244_ ^ _7251_ /*86783*/;
assign _7249_ = _7250_ | _7252_ /*86780*/;
assign _7258_ = ~D[17] /*86779*/;
assign _7255_ = _6673_ & _7258_ /*86775*/;
assign _7256_ = _6673_ ^ _7258_ /*86778*/;
assign _7257_ = _7249_ & _7256_ /*86776*/;
assign _7122_ = _7249_ ^ _7256_ /*86777*/;
assign _7254_ = _7255_ | _7257_ /*86774*/;
assign _7263_ = ~D[18] /*86773*/;
assign _7260_ = _6674_ & _7263_ /*86769*/;
assign _7261_ = _6674_ ^ _7263_ /*86772*/;
assign _7262_ = _7254_ & _7261_ /*86770*/;
assign _7123_ = _7254_ ^ _7261_ /*86771*/;
assign _7259_ = _7260_ | _7262_ /*86768*/;
assign _7268_ = ~D[19] /*86767*/;
assign _7265_ = _6675_ & _7268_ /*86763*/;
assign _7266_ = _6675_ ^ _7268_ /*86766*/;
assign _7267_ = _7259_ & _7266_ /*86764*/;
assign _7124_ = _7259_ ^ _7266_ /*86765*/;
assign _7264_ = _7265_ | _7267_ /*86762*/;
assign _7273_ = ~D[20] /*86761*/;
assign _7270_ = _6676_ & _7273_ /*86757*/;
assign _7271_ = _6676_ ^ _7273_ /*86760*/;
assign _7272_ = _7264_ & _7271_ /*86758*/;
assign _7125_ = _7264_ ^ _7271_ /*86759*/;
assign _7269_ = _7270_ | _7272_ /*86756*/;
assign _7278_ = ~D[21] /*86755*/;
assign _7275_ = _6677_ & _7278_ /*86751*/;
assign _7276_ = _6677_ ^ _7278_ /*86754*/;
assign _7277_ = _7269_ & _7276_ /*86752*/;
assign _7126_ = _7269_ ^ _7276_ /*86753*/;
assign _7274_ = _7275_ | _7277_ /*86750*/;
assign _7283_ = ~D[22] /*86749*/;
assign _7280_ = _6678_ & _7283_ /*86745*/;
assign _7281_ = _6678_ ^ _7283_ /*86748*/;
assign _7282_ = _7274_ & _7281_ /*86746*/;
assign _7127_ = _7274_ ^ _7281_ /*86747*/;
assign _7279_ = _7280_ | _7282_ /*86744*/;
assign _7288_ = ~D[23] /*86743*/;
assign _7285_ = _6679_ & _7288_ /*86739*/;
assign _7286_ = _6679_ ^ _7288_ /*86742*/;
assign _7287_ = _7279_ & _7286_ /*86740*/;
assign _7128_ = _7279_ ^ _7286_ /*86741*/;
assign _7284_ = _7285_ | _7287_ /*86738*/;
assign _7293_ = ~D[24] /*86737*/;
assign _7290_ = _6680_ & _7293_ /*86733*/;
assign _7291_ = _6680_ ^ _7293_ /*86736*/;
assign _7292_ = _7284_ & _7291_ /*86734*/;
assign _7129_ = _7284_ ^ _7291_ /*86735*/;
assign _7289_ = _7290_ | _7292_ /*86732*/;
assign _7298_ = ~D[25] /*86731*/;
assign _7295_ = _6681_ & _7298_ /*86727*/;
assign _7296_ = _6681_ ^ _7298_ /*86730*/;
assign _7297_ = _7289_ & _7296_ /*86728*/;
assign _7130_ = _7289_ ^ _7296_ /*86729*/;
assign _7294_ = _7295_ | _7297_ /*86726*/;
assign _7303_ = ~D[26] /*86725*/;
assign _7300_ = _6682_ & _7303_ /*86721*/;
assign _7301_ = _6682_ ^ _7303_ /*86724*/;
assign _7302_ = _7294_ & _7301_ /*86722*/;
assign _7131_ = _7294_ ^ _7301_ /*86723*/;
assign _7299_ = _7300_ | _7302_ /*86720*/;
assign _7308_ = ~D[27] /*86719*/;
assign _7305_ = _6683_ & _7308_ /*86715*/;
assign _7306_ = _6683_ ^ _7308_ /*86718*/;
assign _7307_ = _7299_ & _7306_ /*86716*/;
assign _7132_ = _7299_ ^ _7306_ /*86717*/;
assign _7304_ = _7305_ | _7307_ /*86714*/;
assign _7313_ = ~D[28] /*86713*/;
assign _7310_ = _6684_ & _7313_ /*86709*/;
assign _7311_ = _6684_ ^ _7313_ /*86712*/;
assign _7312_ = _7304_ & _7311_ /*86710*/;
assign _7133_ = _7304_ ^ _7311_ /*86711*/;
assign _7309_ = _7310_ | _7312_ /*86708*/;
assign _7318_ = ~D[29] /*86707*/;
assign _7315_ = _6685_ & _7318_ /*86703*/;
assign _7316_ = _6685_ ^ _7318_ /*86706*/;
assign _7317_ = _7309_ & _7316_ /*86704*/;
assign _7134_ = _7309_ ^ _7316_ /*86705*/;
assign _7314_ = _7315_ | _7317_ /*86702*/;
assign _7323_ = ~D[30] /*86701*/;
assign _7320_ = _6686_ & _7323_ /*86697*/;
assign _7321_ = _6686_ ^ _7323_ /*86700*/;
assign _7322_ = _7314_ & _7321_ /*86698*/;
assign _7135_ = _7314_ ^ _7321_ /*86699*/;
assign _7319_ = _7320_ | _7322_ /*86696*/;
assign _7328_ = ~D[31] /*86695*/;
assign _7325_ = _6687_ & _7328_ /*86691*/;
assign _7326_ = _6687_ ^ _7328_ /*86694*/;
assign _7327_ = _7319_ & _7326_ /*86692*/;
assign _7136_ = _7319_ ^ _7326_ /*86693*/;
assign _7324_ = _7325_ | _7327_ /*86690*/;
assign _7333_ = ~D[32] /*86689*/;
assign _7330_ = _6688_ & _7333_ /*86685*/;
assign _7331_ = _6688_ ^ _7333_ /*86688*/;
assign _7332_ = _7324_ & _7331_ /*86686*/;
assign _7137_ = _7324_ ^ _7331_ /*86687*/;
assign _7329_ = _7330_ | _7332_ /*86684*/;
assign _7338_ = ~D[33] /*86683*/;
assign _7335_ = _6689_ & _7338_ /*86679*/;
assign _7336_ = _6689_ ^ _7338_ /*86682*/;
assign _7337_ = _7329_ & _7336_ /*86680*/;
assign _7138_ = _7329_ ^ _7336_ /*86681*/;
assign _7334_ = _7335_ | _7337_ /*86678*/;
assign _7343_ = ~D[34] /*86677*/;
assign _7340_ = _6690_ & _7343_ /*86673*/;
assign _7341_ = _6690_ ^ _7343_ /*86676*/;
assign _7342_ = _7334_ & _7341_ /*86674*/;
assign _7139_ = _7334_ ^ _7341_ /*86675*/;
assign _7339_ = _7340_ | _7342_ /*86672*/;
assign _7348_ = ~D[35] /*86671*/;
assign _7345_ = _6691_ & _7348_ /*86667*/;
assign _7346_ = _6691_ ^ _7348_ /*86670*/;
assign _7347_ = _7339_ & _7346_ /*86668*/;
assign _7140_ = _7339_ ^ _7346_ /*86669*/;
assign _7344_ = _7345_ | _7347_ /*86666*/;
assign _7353_ = ~D[36] /*86665*/;
assign _7350_ = _6692_ & _7353_ /*86661*/;
assign _7351_ = _6692_ ^ _7353_ /*86664*/;
assign _7352_ = _7344_ & _7351_ /*86662*/;
assign _7141_ = _7344_ ^ _7351_ /*86663*/;
assign _7349_ = _7350_ | _7352_ /*86660*/;
assign _7358_ = ~D[37] /*86659*/;
assign _7355_ = _6693_ & _7358_ /*86655*/;
assign _7356_ = _6693_ ^ _7358_ /*86658*/;
assign _7357_ = _7349_ & _7356_ /*86656*/;
assign _7142_ = _7349_ ^ _7356_ /*86657*/;
assign _7354_ = _7355_ | _7357_ /*86654*/;
assign _7363_ = ~D[38] /*86653*/;
assign _7360_ = _6694_ & _7363_ /*86649*/;
assign _7361_ = _6694_ ^ _7363_ /*86652*/;
assign _7362_ = _7354_ & _7361_ /*86650*/;
assign _7143_ = _7354_ ^ _7361_ /*86651*/;
assign _7359_ = _7360_ | _7362_ /*86648*/;
assign _7368_ = ~D[39] /*86647*/;
assign _7365_ = _6695_ & _7368_ /*86643*/;
assign _7366_ = _6695_ ^ _7368_ /*86646*/;
assign _7367_ = _7359_ & _7366_ /*86644*/;
assign _7144_ = _7359_ ^ _7366_ /*86645*/;
assign _7364_ = _7365_ | _7367_ /*86642*/;
assign _7373_ = ~D[40] /*86641*/;
assign _7370_ = _6696_ & _7373_ /*86637*/;
assign _7371_ = _6696_ ^ _7373_ /*86640*/;
assign _7372_ = _7364_ & _7371_ /*86638*/;
assign _7145_ = _7364_ ^ _7371_ /*86639*/;
assign _7369_ = _7370_ | _7372_ /*86636*/;
assign _7378_ = ~D[41] /*86635*/;
assign _7375_ = _6697_ & _7378_ /*86631*/;
assign _7376_ = _6697_ ^ _7378_ /*86634*/;
assign _7377_ = _7369_ & _7376_ /*86632*/;
assign _7146_ = _7369_ ^ _7376_ /*86633*/;
assign _7374_ = _7375_ | _7377_ /*86630*/;
assign _7383_ = ~D[42] /*86629*/;
assign _7380_ = _6698_ & _7383_ /*86625*/;
assign _7381_ = _6698_ ^ _7383_ /*86628*/;
assign _7382_ = _7374_ & _7381_ /*86626*/;
assign _7147_ = _7374_ ^ _7381_ /*86627*/;
assign _7379_ = _7380_ | _7382_ /*86624*/;
assign _7388_ = ~D[43] /*86623*/;
assign _7385_ = _6699_ & _7388_ /*86619*/;
assign _7386_ = _6699_ ^ _7388_ /*86622*/;
assign _7387_ = _7379_ & _7386_ /*86620*/;
assign _7148_ = _7379_ ^ _7386_ /*86621*/;
assign _7384_ = _7385_ | _7387_ /*86618*/;
assign _7393_ = ~D[44] /*86617*/;
assign _7390_ = _6700_ & _7393_ /*86613*/;
assign _7391_ = _6700_ ^ _7393_ /*86616*/;
assign _7392_ = _7384_ & _7391_ /*86614*/;
assign _7149_ = _7384_ ^ _7391_ /*86615*/;
assign _7389_ = _7390_ | _7392_ /*86612*/;
assign _7398_ = ~D[45] /*86611*/;
assign _7395_ = _6701_ & _7398_ /*86607*/;
assign _7396_ = _6701_ ^ _7398_ /*86610*/;
assign _7397_ = _7389_ & _7396_ /*86608*/;
assign _7150_ = _7389_ ^ _7396_ /*86609*/;
assign _7394_ = _7395_ | _7397_ /*86606*/;
assign _7403_ = ~D[46] /*86605*/;
assign _7400_ = _6702_ & _7403_ /*86601*/;
assign _7401_ = _6702_ ^ _7403_ /*86604*/;
assign _7402_ = _7394_ & _7401_ /*86602*/;
assign _7151_ = _7394_ ^ _7401_ /*86603*/;
assign _7399_ = _7400_ | _7402_ /*86600*/;
assign _7408_ = ~D[47] /*86599*/;
assign _7405_ = _6703_ & _7408_ /*86595*/;
assign _7406_ = _6703_ ^ _7408_ /*86598*/;
assign _7407_ = _7399_ & _7406_ /*86596*/;
assign _7152_ = _7399_ ^ _7406_ /*86597*/;
assign _7404_ = _7405_ | _7407_ /*86594*/;
assign _7413_ = ~D[48] /*86593*/;
assign _7410_ = _6704_ & _7413_ /*86589*/;
assign _7411_ = _6704_ ^ _7413_ /*86592*/;
assign _7412_ = _7404_ & _7411_ /*86590*/;
assign _7153_ = _7404_ ^ _7411_ /*86591*/;
assign _7409_ = _7410_ | _7412_ /*86588*/;
assign _7418_ = ~D[49] /*86587*/;
assign _7415_ = _6705_ & _7418_ /*86583*/;
assign _7416_ = _6705_ ^ _7418_ /*86586*/;
assign _7417_ = _7409_ & _7416_ /*86584*/;
assign _7154_ = _7409_ ^ _7416_ /*86585*/;
assign _7414_ = _7415_ | _7417_ /*86582*/;
assign _7423_ = ~D[50] /*86581*/;
assign _7420_ = _6706_ & _7423_ /*86577*/;
assign _7421_ = _6706_ ^ _7423_ /*86580*/;
assign _7422_ = _7414_ & _7421_ /*86578*/;
assign _7155_ = _7414_ ^ _7421_ /*86579*/;
assign _7419_ = _7420_ | _7422_ /*86576*/;
assign _7428_ = ~D[51] /*86575*/;
assign _7425_ = _6707_ & _7428_ /*86571*/;
assign _7426_ = _6707_ ^ _7428_ /*86574*/;
assign _7427_ = _7419_ & _7426_ /*86572*/;
assign _7156_ = _7419_ ^ _7426_ /*86573*/;
assign _7424_ = _7425_ | _7427_ /*86570*/;
assign _7433_ = ~D[52] /*86569*/;
assign _7430_ = _6708_ & _7433_ /*86565*/;
assign _7431_ = _6708_ ^ _7433_ /*86568*/;
assign _7432_ = _7424_ & _7431_ /*86566*/;
assign _7157_ = _7424_ ^ _7431_ /*86567*/;
assign _7429_ = _7430_ | _7432_ /*86564*/;
assign _7438_ = ~D[53] /*86563*/;
assign _7435_ = _6709_ & _7438_ /*86559*/;
assign _7436_ = _6709_ ^ _7438_ /*86562*/;
assign _7437_ = _7429_ & _7436_ /*86560*/;
assign _7158_ = _7429_ ^ _7436_ /*86561*/;
assign _7434_ = _7435_ | _7437_ /*86558*/;
assign _7443_ = ~D[54] /*86557*/;
assign _7440_ = _6710_ & _7443_ /*86553*/;
assign _7441_ = _6710_ ^ _7443_ /*86556*/;
assign _7442_ = _7434_ & _7441_ /*86554*/;
assign _7159_ = _7434_ ^ _7441_ /*86555*/;
assign _7439_ = _7440_ | _7442_ /*86552*/;
assign _7448_ = ~D[55] /*86551*/;
assign _7445_ = _6711_ & _7448_ /*86547*/;
assign _7446_ = _6711_ ^ _7448_ /*86550*/;
assign _7447_ = _7439_ & _7446_ /*86548*/;
assign _7160_ = _7439_ ^ _7446_ /*86549*/;
assign _7444_ = _7445_ | _7447_ /*86546*/;
assign _7453_ = ~D[56] /*86545*/;
assign _7450_ = _6712_ & _7453_ /*86541*/;
assign _7451_ = _6712_ ^ _7453_ /*86544*/;
assign _7452_ = _7444_ & _7451_ /*86542*/;
assign _7161_ = _7444_ ^ _7451_ /*86543*/;
assign _7449_ = _7450_ | _7452_ /*86540*/;
assign _7458_ = ~D[57] /*86539*/;
assign _7455_ = _6713_ & _7458_ /*86535*/;
assign _7456_ = _6713_ ^ _7458_ /*86538*/;
assign _7457_ = _7449_ & _7456_ /*86536*/;
assign _7162_ = _7449_ ^ _7456_ /*86537*/;
assign _7454_ = _7455_ | _7457_ /*86534*/;
assign _7463_ = ~D[58] /*86533*/;
assign _7460_ = _6714_ & _7463_ /*86529*/;
assign _7461_ = _6714_ ^ _7463_ /*86532*/;
assign _7462_ = _7454_ & _7461_ /*86530*/;
assign _7163_ = _7454_ ^ _7461_ /*86531*/;
assign _7459_ = _7460_ | _7462_ /*86528*/;
assign _7468_ = ~D[59] /*86527*/;
assign _7465_ = _6715_ & _7468_ /*86523*/;
assign _7466_ = _6715_ ^ _7468_ /*86526*/;
assign _7467_ = _7459_ & _7466_ /*86524*/;
assign _7164_ = _7459_ ^ _7466_ /*86525*/;
assign _7464_ = _7465_ | _7467_ /*86522*/;
assign _7473_ = ~D[60] /*86521*/;
assign _7470_ = _6716_ & _7473_ /*86517*/;
assign _7471_ = _6716_ ^ _7473_ /*86520*/;
assign _7472_ = _7464_ & _7471_ /*86518*/;
assign _7165_ = _7464_ ^ _7471_ /*86519*/;
assign _7469_ = _7470_ | _7472_ /*86516*/;
assign _7478_ = ~D[61] /*86515*/;
assign _7475_ = _6717_ & _7478_ /*86511*/;
assign _7476_ = _6717_ ^ _7478_ /*86514*/;
assign _7477_ = _7469_ & _7476_ /*86512*/;
assign _7166_ = _7469_ ^ _7476_ /*86513*/;
assign _7474_ = _7475_ | _7477_ /*86510*/;
assign _7483_ = ~D[62] /*86509*/;
assign _7480_ = _6718_ & _7483_ /*86505*/;
assign _7481_ = _6718_ ^ _7483_ /*86508*/;
assign _7482_ = _7474_ & _7481_ /*86506*/;
assign _7167_ = _7474_ ^ _7481_ /*86507*/;
assign _7479_ = _7480_ | _7482_ /*86504*/;
assign _7484_ = _6719_ & oneWire /*86499*/;
assign _7485_ = _6719_ ^ oneWire /*86502*/;
assign _7486_ = _7479_ & _7485_ /*86500*/;
assign _7168_ = _7479_ ^ _7485_ /*86501*/;
assign Q[55] = _7484_ | _7486_ /*86498*/;
assign _7619_ = ~Q[55] /*86113*/;
assign _7618_ = _7619_ & D[0] /*86112*/;
assign _7621_ = _7105_ & _7618_ /*86107*/;
assign _7622_ = _7105_ ^ _7618_ /*86110*/;
assign _7623_ = zeroWire & _7622_ /*86108*/;
assign _7553_ = zeroWire ^ _7622_ /*86109*/;
assign _7620_ = _7621_ | _7623_ /*86106*/;
assign _7625_ = ~Q[55] /*86105*/;
assign _7624_ = _7625_ & D[1] /*86104*/;
assign _7627_ = _7106_ & _7624_ /*86099*/;
assign _7628_ = _7106_ ^ _7624_ /*86102*/;
assign _7629_ = _7620_ & _7628_ /*86100*/;
assign _7554_ = _7620_ ^ _7628_ /*86101*/;
assign _7626_ = _7627_ | _7629_ /*86098*/;
assign _7631_ = ~Q[55] /*86097*/;
assign _7630_ = _7631_ & D[2] /*86096*/;
assign _7633_ = _7107_ & _7630_ /*86091*/;
assign _7634_ = _7107_ ^ _7630_ /*86094*/;
assign _7635_ = _7626_ & _7634_ /*86092*/;
assign _7555_ = _7626_ ^ _7634_ /*86093*/;
assign _7632_ = _7633_ | _7635_ /*86090*/;
assign _7637_ = ~Q[55] /*86089*/;
assign _7636_ = _7637_ & D[3] /*86088*/;
assign _7639_ = _7108_ & _7636_ /*86083*/;
assign _7640_ = _7108_ ^ _7636_ /*86086*/;
assign _7641_ = _7632_ & _7640_ /*86084*/;
assign _7556_ = _7632_ ^ _7640_ /*86085*/;
assign _7638_ = _7639_ | _7641_ /*86082*/;
assign _7643_ = ~Q[55] /*86081*/;
assign _7642_ = _7643_ & D[4] /*86080*/;
assign _7645_ = _7109_ & _7642_ /*86075*/;
assign _7646_ = _7109_ ^ _7642_ /*86078*/;
assign _7647_ = _7638_ & _7646_ /*86076*/;
assign _7557_ = _7638_ ^ _7646_ /*86077*/;
assign _7644_ = _7645_ | _7647_ /*86074*/;
assign _7649_ = ~Q[55] /*86073*/;
assign _7648_ = _7649_ & D[5] /*86072*/;
assign _7651_ = _7110_ & _7648_ /*86067*/;
assign _7652_ = _7110_ ^ _7648_ /*86070*/;
assign _7653_ = _7644_ & _7652_ /*86068*/;
assign _7558_ = _7644_ ^ _7652_ /*86069*/;
assign _7650_ = _7651_ | _7653_ /*86066*/;
assign _7655_ = ~Q[55] /*86065*/;
assign _7654_ = _7655_ & D[6] /*86064*/;
assign _7657_ = _7111_ & _7654_ /*86059*/;
assign _7658_ = _7111_ ^ _7654_ /*86062*/;
assign _7659_ = _7650_ & _7658_ /*86060*/;
assign _7559_ = _7650_ ^ _7658_ /*86061*/;
assign _7656_ = _7657_ | _7659_ /*86058*/;
assign _7661_ = ~Q[55] /*86057*/;
assign _7660_ = _7661_ & D[7] /*86056*/;
assign _7663_ = _7112_ & _7660_ /*86051*/;
assign _7664_ = _7112_ ^ _7660_ /*86054*/;
assign _7665_ = _7656_ & _7664_ /*86052*/;
assign _7560_ = _7656_ ^ _7664_ /*86053*/;
assign _7662_ = _7663_ | _7665_ /*86050*/;
assign _7667_ = ~Q[55] /*86049*/;
assign _7666_ = _7667_ & D[8] /*86048*/;
assign _7669_ = _7113_ & _7666_ /*86043*/;
assign _7670_ = _7113_ ^ _7666_ /*86046*/;
assign _7671_ = _7662_ & _7670_ /*86044*/;
assign _7561_ = _7662_ ^ _7670_ /*86045*/;
assign _7668_ = _7669_ | _7671_ /*86042*/;
assign _7673_ = ~Q[55] /*86041*/;
assign _7672_ = _7673_ & D[9] /*86040*/;
assign _7675_ = _7114_ & _7672_ /*86035*/;
assign _7676_ = _7114_ ^ _7672_ /*86038*/;
assign _7677_ = _7668_ & _7676_ /*86036*/;
assign _7562_ = _7668_ ^ _7676_ /*86037*/;
assign _7674_ = _7675_ | _7677_ /*86034*/;
assign _7679_ = ~Q[55] /*86033*/;
assign _7678_ = _7679_ & D[10] /*86032*/;
assign _7681_ = _7115_ & _7678_ /*86027*/;
assign _7682_ = _7115_ ^ _7678_ /*86030*/;
assign _7683_ = _7674_ & _7682_ /*86028*/;
assign _7563_ = _7674_ ^ _7682_ /*86029*/;
assign _7680_ = _7681_ | _7683_ /*86026*/;
assign _7685_ = ~Q[55] /*86025*/;
assign _7684_ = _7685_ & D[11] /*86024*/;
assign _7687_ = _7116_ & _7684_ /*86019*/;
assign _7688_ = _7116_ ^ _7684_ /*86022*/;
assign _7689_ = _7680_ & _7688_ /*86020*/;
assign _7564_ = _7680_ ^ _7688_ /*86021*/;
assign _7686_ = _7687_ | _7689_ /*86018*/;
assign _7691_ = ~Q[55] /*86017*/;
assign _7690_ = _7691_ & D[12] /*86016*/;
assign _7693_ = _7117_ & _7690_ /*86011*/;
assign _7694_ = _7117_ ^ _7690_ /*86014*/;
assign _7695_ = _7686_ & _7694_ /*86012*/;
assign _7565_ = _7686_ ^ _7694_ /*86013*/;
assign _7692_ = _7693_ | _7695_ /*86010*/;
assign _7697_ = ~Q[55] /*86009*/;
assign _7696_ = _7697_ & D[13] /*86008*/;
assign _7699_ = _7118_ & _7696_ /*86003*/;
assign _7700_ = _7118_ ^ _7696_ /*86006*/;
assign _7701_ = _7692_ & _7700_ /*86004*/;
assign _7566_ = _7692_ ^ _7700_ /*86005*/;
assign _7698_ = _7699_ | _7701_ /*86002*/;
assign _7703_ = ~Q[55] /*86001*/;
assign _7702_ = _7703_ & D[14] /*86000*/;
assign _7705_ = _7119_ & _7702_ /*85995*/;
assign _7706_ = _7119_ ^ _7702_ /*85998*/;
assign _7707_ = _7698_ & _7706_ /*85996*/;
assign _7567_ = _7698_ ^ _7706_ /*85997*/;
assign _7704_ = _7705_ | _7707_ /*85994*/;
assign _7709_ = ~Q[55] /*85993*/;
assign _7708_ = _7709_ & D[15] /*85992*/;
assign _7711_ = _7120_ & _7708_ /*85987*/;
assign _7712_ = _7120_ ^ _7708_ /*85990*/;
assign _7713_ = _7704_ & _7712_ /*85988*/;
assign _7568_ = _7704_ ^ _7712_ /*85989*/;
assign _7710_ = _7711_ | _7713_ /*85986*/;
assign _7715_ = ~Q[55] /*85985*/;
assign _7714_ = _7715_ & D[16] /*85984*/;
assign _7717_ = _7121_ & _7714_ /*85979*/;
assign _7718_ = _7121_ ^ _7714_ /*85982*/;
assign _7719_ = _7710_ & _7718_ /*85980*/;
assign _7569_ = _7710_ ^ _7718_ /*85981*/;
assign _7716_ = _7717_ | _7719_ /*85978*/;
assign _7721_ = ~Q[55] /*85977*/;
assign _7720_ = _7721_ & D[17] /*85976*/;
assign _7723_ = _7122_ & _7720_ /*85971*/;
assign _7724_ = _7122_ ^ _7720_ /*85974*/;
assign _7725_ = _7716_ & _7724_ /*85972*/;
assign _7570_ = _7716_ ^ _7724_ /*85973*/;
assign _7722_ = _7723_ | _7725_ /*85970*/;
assign _7727_ = ~Q[55] /*85969*/;
assign _7726_ = _7727_ & D[18] /*85968*/;
assign _7729_ = _7123_ & _7726_ /*85963*/;
assign _7730_ = _7123_ ^ _7726_ /*85966*/;
assign _7731_ = _7722_ & _7730_ /*85964*/;
assign _7571_ = _7722_ ^ _7730_ /*85965*/;
assign _7728_ = _7729_ | _7731_ /*85962*/;
assign _7733_ = ~Q[55] /*85961*/;
assign _7732_ = _7733_ & D[19] /*85960*/;
assign _7735_ = _7124_ & _7732_ /*85955*/;
assign _7736_ = _7124_ ^ _7732_ /*85958*/;
assign _7737_ = _7728_ & _7736_ /*85956*/;
assign _7572_ = _7728_ ^ _7736_ /*85957*/;
assign _7734_ = _7735_ | _7737_ /*85954*/;
assign _7739_ = ~Q[55] /*85953*/;
assign _7738_ = _7739_ & D[20] /*85952*/;
assign _7741_ = _7125_ & _7738_ /*85947*/;
assign _7742_ = _7125_ ^ _7738_ /*85950*/;
assign _7743_ = _7734_ & _7742_ /*85948*/;
assign _7573_ = _7734_ ^ _7742_ /*85949*/;
assign _7740_ = _7741_ | _7743_ /*85946*/;
assign _7745_ = ~Q[55] /*85945*/;
assign _7744_ = _7745_ & D[21] /*85944*/;
assign _7747_ = _7126_ & _7744_ /*85939*/;
assign _7748_ = _7126_ ^ _7744_ /*85942*/;
assign _7749_ = _7740_ & _7748_ /*85940*/;
assign _7574_ = _7740_ ^ _7748_ /*85941*/;
assign _7746_ = _7747_ | _7749_ /*85938*/;
assign _7751_ = ~Q[55] /*85937*/;
assign _7750_ = _7751_ & D[22] /*85936*/;
assign _7753_ = _7127_ & _7750_ /*85931*/;
assign _7754_ = _7127_ ^ _7750_ /*85934*/;
assign _7755_ = _7746_ & _7754_ /*85932*/;
assign _7575_ = _7746_ ^ _7754_ /*85933*/;
assign _7752_ = _7753_ | _7755_ /*85930*/;
assign _7757_ = ~Q[55] /*85929*/;
assign _7756_ = _7757_ & D[23] /*85928*/;
assign _7759_ = _7128_ & _7756_ /*85923*/;
assign _7760_ = _7128_ ^ _7756_ /*85926*/;
assign _7761_ = _7752_ & _7760_ /*85924*/;
assign _7576_ = _7752_ ^ _7760_ /*85925*/;
assign _7758_ = _7759_ | _7761_ /*85922*/;
assign _7763_ = ~Q[55] /*85921*/;
assign _7762_ = _7763_ & D[24] /*85920*/;
assign _7765_ = _7129_ & _7762_ /*85915*/;
assign _7766_ = _7129_ ^ _7762_ /*85918*/;
assign _7767_ = _7758_ & _7766_ /*85916*/;
assign _7577_ = _7758_ ^ _7766_ /*85917*/;
assign _7764_ = _7765_ | _7767_ /*85914*/;
assign _7769_ = ~Q[55] /*85913*/;
assign _7768_ = _7769_ & D[25] /*85912*/;
assign _7771_ = _7130_ & _7768_ /*85907*/;
assign _7772_ = _7130_ ^ _7768_ /*85910*/;
assign _7773_ = _7764_ & _7772_ /*85908*/;
assign _7578_ = _7764_ ^ _7772_ /*85909*/;
assign _7770_ = _7771_ | _7773_ /*85906*/;
assign _7775_ = ~Q[55] /*85905*/;
assign _7774_ = _7775_ & D[26] /*85904*/;
assign _7777_ = _7131_ & _7774_ /*85899*/;
assign _7778_ = _7131_ ^ _7774_ /*85902*/;
assign _7779_ = _7770_ & _7778_ /*85900*/;
assign _7579_ = _7770_ ^ _7778_ /*85901*/;
assign _7776_ = _7777_ | _7779_ /*85898*/;
assign _7781_ = ~Q[55] /*85897*/;
assign _7780_ = _7781_ & D[27] /*85896*/;
assign _7783_ = _7132_ & _7780_ /*85891*/;
assign _7784_ = _7132_ ^ _7780_ /*85894*/;
assign _7785_ = _7776_ & _7784_ /*85892*/;
assign _7580_ = _7776_ ^ _7784_ /*85893*/;
assign _7782_ = _7783_ | _7785_ /*85890*/;
assign _7787_ = ~Q[55] /*85889*/;
assign _7786_ = _7787_ & D[28] /*85888*/;
assign _7789_ = _7133_ & _7786_ /*85883*/;
assign _7790_ = _7133_ ^ _7786_ /*85886*/;
assign _7791_ = _7782_ & _7790_ /*85884*/;
assign _7581_ = _7782_ ^ _7790_ /*85885*/;
assign _7788_ = _7789_ | _7791_ /*85882*/;
assign _7793_ = ~Q[55] /*85881*/;
assign _7792_ = _7793_ & D[29] /*85880*/;
assign _7795_ = _7134_ & _7792_ /*85875*/;
assign _7796_ = _7134_ ^ _7792_ /*85878*/;
assign _7797_ = _7788_ & _7796_ /*85876*/;
assign _7582_ = _7788_ ^ _7796_ /*85877*/;
assign _7794_ = _7795_ | _7797_ /*85874*/;
assign _7799_ = ~Q[55] /*85873*/;
assign _7798_ = _7799_ & D[30] /*85872*/;
assign _7801_ = _7135_ & _7798_ /*85867*/;
assign _7802_ = _7135_ ^ _7798_ /*85870*/;
assign _7803_ = _7794_ & _7802_ /*85868*/;
assign _7583_ = _7794_ ^ _7802_ /*85869*/;
assign _7800_ = _7801_ | _7803_ /*85866*/;
assign _7805_ = ~Q[55] /*85865*/;
assign _7804_ = _7805_ & D[31] /*85864*/;
assign _7807_ = _7136_ & _7804_ /*85859*/;
assign _7808_ = _7136_ ^ _7804_ /*85862*/;
assign _7809_ = _7800_ & _7808_ /*85860*/;
assign _7584_ = _7800_ ^ _7808_ /*85861*/;
assign _7806_ = _7807_ | _7809_ /*85858*/;
assign _7811_ = ~Q[55] /*85857*/;
assign _7810_ = _7811_ & D[32] /*85856*/;
assign _7813_ = _7137_ & _7810_ /*85851*/;
assign _7814_ = _7137_ ^ _7810_ /*85854*/;
assign _7815_ = _7806_ & _7814_ /*85852*/;
assign _7585_ = _7806_ ^ _7814_ /*85853*/;
assign _7812_ = _7813_ | _7815_ /*85850*/;
assign _7817_ = ~Q[55] /*85849*/;
assign _7816_ = _7817_ & D[33] /*85848*/;
assign _7819_ = _7138_ & _7816_ /*85843*/;
assign _7820_ = _7138_ ^ _7816_ /*85846*/;
assign _7821_ = _7812_ & _7820_ /*85844*/;
assign _7586_ = _7812_ ^ _7820_ /*85845*/;
assign _7818_ = _7819_ | _7821_ /*85842*/;
assign _7823_ = ~Q[55] /*85841*/;
assign _7822_ = _7823_ & D[34] /*85840*/;
assign _7825_ = _7139_ & _7822_ /*85835*/;
assign _7826_ = _7139_ ^ _7822_ /*85838*/;
assign _7827_ = _7818_ & _7826_ /*85836*/;
assign _7587_ = _7818_ ^ _7826_ /*85837*/;
assign _7824_ = _7825_ | _7827_ /*85834*/;
assign _7829_ = ~Q[55] /*85833*/;
assign _7828_ = _7829_ & D[35] /*85832*/;
assign _7831_ = _7140_ & _7828_ /*85827*/;
assign _7832_ = _7140_ ^ _7828_ /*85830*/;
assign _7833_ = _7824_ & _7832_ /*85828*/;
assign _7588_ = _7824_ ^ _7832_ /*85829*/;
assign _7830_ = _7831_ | _7833_ /*85826*/;
assign _7835_ = ~Q[55] /*85825*/;
assign _7834_ = _7835_ & D[36] /*85824*/;
assign _7837_ = _7141_ & _7834_ /*85819*/;
assign _7838_ = _7141_ ^ _7834_ /*85822*/;
assign _7839_ = _7830_ & _7838_ /*85820*/;
assign _7589_ = _7830_ ^ _7838_ /*85821*/;
assign _7836_ = _7837_ | _7839_ /*85818*/;
assign _7841_ = ~Q[55] /*85817*/;
assign _7840_ = _7841_ & D[37] /*85816*/;
assign _7843_ = _7142_ & _7840_ /*85811*/;
assign _7844_ = _7142_ ^ _7840_ /*85814*/;
assign _7845_ = _7836_ & _7844_ /*85812*/;
assign _7590_ = _7836_ ^ _7844_ /*85813*/;
assign _7842_ = _7843_ | _7845_ /*85810*/;
assign _7847_ = ~Q[55] /*85809*/;
assign _7846_ = _7847_ & D[38] /*85808*/;
assign _7849_ = _7143_ & _7846_ /*85803*/;
assign _7850_ = _7143_ ^ _7846_ /*85806*/;
assign _7851_ = _7842_ & _7850_ /*85804*/;
assign _7591_ = _7842_ ^ _7850_ /*85805*/;
assign _7848_ = _7849_ | _7851_ /*85802*/;
assign _7853_ = ~Q[55] /*85801*/;
assign _7852_ = _7853_ & D[39] /*85800*/;
assign _7855_ = _7144_ & _7852_ /*85795*/;
assign _7856_ = _7144_ ^ _7852_ /*85798*/;
assign _7857_ = _7848_ & _7856_ /*85796*/;
assign _7592_ = _7848_ ^ _7856_ /*85797*/;
assign _7854_ = _7855_ | _7857_ /*85794*/;
assign _7859_ = ~Q[55] /*85793*/;
assign _7858_ = _7859_ & D[40] /*85792*/;
assign _7861_ = _7145_ & _7858_ /*85787*/;
assign _7862_ = _7145_ ^ _7858_ /*85790*/;
assign _7863_ = _7854_ & _7862_ /*85788*/;
assign _7593_ = _7854_ ^ _7862_ /*85789*/;
assign _7860_ = _7861_ | _7863_ /*85786*/;
assign _7865_ = ~Q[55] /*85785*/;
assign _7864_ = _7865_ & D[41] /*85784*/;
assign _7867_ = _7146_ & _7864_ /*85779*/;
assign _7868_ = _7146_ ^ _7864_ /*85782*/;
assign _7869_ = _7860_ & _7868_ /*85780*/;
assign _7594_ = _7860_ ^ _7868_ /*85781*/;
assign _7866_ = _7867_ | _7869_ /*85778*/;
assign _7871_ = ~Q[55] /*85777*/;
assign _7870_ = _7871_ & D[42] /*85776*/;
assign _7873_ = _7147_ & _7870_ /*85771*/;
assign _7874_ = _7147_ ^ _7870_ /*85774*/;
assign _7875_ = _7866_ & _7874_ /*85772*/;
assign _7595_ = _7866_ ^ _7874_ /*85773*/;
assign _7872_ = _7873_ | _7875_ /*85770*/;
assign _7877_ = ~Q[55] /*85769*/;
assign _7876_ = _7877_ & D[43] /*85768*/;
assign _7879_ = _7148_ & _7876_ /*85763*/;
assign _7880_ = _7148_ ^ _7876_ /*85766*/;
assign _7881_ = _7872_ & _7880_ /*85764*/;
assign _7596_ = _7872_ ^ _7880_ /*85765*/;
assign _7878_ = _7879_ | _7881_ /*85762*/;
assign _7883_ = ~Q[55] /*85761*/;
assign _7882_ = _7883_ & D[44] /*85760*/;
assign _7885_ = _7149_ & _7882_ /*85755*/;
assign _7886_ = _7149_ ^ _7882_ /*85758*/;
assign _7887_ = _7878_ & _7886_ /*85756*/;
assign _7597_ = _7878_ ^ _7886_ /*85757*/;
assign _7884_ = _7885_ | _7887_ /*85754*/;
assign _7889_ = ~Q[55] /*85753*/;
assign _7888_ = _7889_ & D[45] /*85752*/;
assign _7891_ = _7150_ & _7888_ /*85747*/;
assign _7892_ = _7150_ ^ _7888_ /*85750*/;
assign _7893_ = _7884_ & _7892_ /*85748*/;
assign _7598_ = _7884_ ^ _7892_ /*85749*/;
assign _7890_ = _7891_ | _7893_ /*85746*/;
assign _7895_ = ~Q[55] /*85745*/;
assign _7894_ = _7895_ & D[46] /*85744*/;
assign _7897_ = _7151_ & _7894_ /*85739*/;
assign _7898_ = _7151_ ^ _7894_ /*85742*/;
assign _7899_ = _7890_ & _7898_ /*85740*/;
assign _7599_ = _7890_ ^ _7898_ /*85741*/;
assign _7896_ = _7897_ | _7899_ /*85738*/;
assign _7901_ = ~Q[55] /*85737*/;
assign _7900_ = _7901_ & D[47] /*85736*/;
assign _7903_ = _7152_ & _7900_ /*85731*/;
assign _7904_ = _7152_ ^ _7900_ /*85734*/;
assign _7905_ = _7896_ & _7904_ /*85732*/;
assign _7600_ = _7896_ ^ _7904_ /*85733*/;
assign _7902_ = _7903_ | _7905_ /*85730*/;
assign _7907_ = ~Q[55] /*85729*/;
assign _7906_ = _7907_ & D[48] /*85728*/;
assign _7909_ = _7153_ & _7906_ /*85723*/;
assign _7910_ = _7153_ ^ _7906_ /*85726*/;
assign _7911_ = _7902_ & _7910_ /*85724*/;
assign _7601_ = _7902_ ^ _7910_ /*85725*/;
assign _7908_ = _7909_ | _7911_ /*85722*/;
assign _7913_ = ~Q[55] /*85721*/;
assign _7912_ = _7913_ & D[49] /*85720*/;
assign _7915_ = _7154_ & _7912_ /*85715*/;
assign _7916_ = _7154_ ^ _7912_ /*85718*/;
assign _7917_ = _7908_ & _7916_ /*85716*/;
assign _7602_ = _7908_ ^ _7916_ /*85717*/;
assign _7914_ = _7915_ | _7917_ /*85714*/;
assign _7919_ = ~Q[55] /*85713*/;
assign _7918_ = _7919_ & D[50] /*85712*/;
assign _7921_ = _7155_ & _7918_ /*85707*/;
assign _7922_ = _7155_ ^ _7918_ /*85710*/;
assign _7923_ = _7914_ & _7922_ /*85708*/;
assign _7603_ = _7914_ ^ _7922_ /*85709*/;
assign _7920_ = _7921_ | _7923_ /*85706*/;
assign _7925_ = ~Q[55] /*85705*/;
assign _7924_ = _7925_ & D[51] /*85704*/;
assign _7927_ = _7156_ & _7924_ /*85699*/;
assign _7928_ = _7156_ ^ _7924_ /*85702*/;
assign _7929_ = _7920_ & _7928_ /*85700*/;
assign _7604_ = _7920_ ^ _7928_ /*85701*/;
assign _7926_ = _7927_ | _7929_ /*85698*/;
assign _7931_ = ~Q[55] /*85697*/;
assign _7930_ = _7931_ & D[52] /*85696*/;
assign _7933_ = _7157_ & _7930_ /*85691*/;
assign _7934_ = _7157_ ^ _7930_ /*85694*/;
assign _7935_ = _7926_ & _7934_ /*85692*/;
assign _7605_ = _7926_ ^ _7934_ /*85693*/;
assign _7932_ = _7933_ | _7935_ /*85690*/;
assign _7937_ = ~Q[55] /*85689*/;
assign _7936_ = _7937_ & D[53] /*85688*/;
assign _7939_ = _7158_ & _7936_ /*85683*/;
assign _7940_ = _7158_ ^ _7936_ /*85686*/;
assign _7941_ = _7932_ & _7940_ /*85684*/;
assign _7606_ = _7932_ ^ _7940_ /*85685*/;
assign _7938_ = _7939_ | _7941_ /*85682*/;
assign _7943_ = ~Q[55] /*85681*/;
assign _7942_ = _7943_ & D[54] /*85680*/;
assign _7945_ = _7159_ & _7942_ /*85675*/;
assign _7946_ = _7159_ ^ _7942_ /*85678*/;
assign _7947_ = _7938_ & _7946_ /*85676*/;
assign _7607_ = _7938_ ^ _7946_ /*85677*/;
assign _7944_ = _7945_ | _7947_ /*85674*/;
assign _7949_ = ~Q[55] /*85673*/;
assign _7948_ = _7949_ & D[55] /*85672*/;
assign _7951_ = _7160_ & _7948_ /*85667*/;
assign _7952_ = _7160_ ^ _7948_ /*85670*/;
assign _7953_ = _7944_ & _7952_ /*85668*/;
assign _7608_ = _7944_ ^ _7952_ /*85669*/;
assign _7950_ = _7951_ | _7953_ /*85666*/;
assign _7955_ = ~Q[55] /*85665*/;
assign _7954_ = _7955_ & D[56] /*85664*/;
assign _7957_ = _7161_ & _7954_ /*85659*/;
assign _7958_ = _7161_ ^ _7954_ /*85662*/;
assign _7959_ = _7950_ & _7958_ /*85660*/;
assign _7609_ = _7950_ ^ _7958_ /*85661*/;
assign _7956_ = _7957_ | _7959_ /*85658*/;
assign _7961_ = ~Q[55] /*85657*/;
assign _7960_ = _7961_ & D[57] /*85656*/;
assign _7963_ = _7162_ & _7960_ /*85651*/;
assign _7964_ = _7162_ ^ _7960_ /*85654*/;
assign _7965_ = _7956_ & _7964_ /*85652*/;
assign _7610_ = _7956_ ^ _7964_ /*85653*/;
assign _7962_ = _7963_ | _7965_ /*85650*/;
assign _7967_ = ~Q[55] /*85649*/;
assign _7966_ = _7967_ & D[58] /*85648*/;
assign _7969_ = _7163_ & _7966_ /*85643*/;
assign _7970_ = _7163_ ^ _7966_ /*85646*/;
assign _7971_ = _7962_ & _7970_ /*85644*/;
assign _7611_ = _7962_ ^ _7970_ /*85645*/;
assign _7968_ = _7969_ | _7971_ /*85642*/;
assign _7973_ = ~Q[55] /*85641*/;
assign _7972_ = _7973_ & D[59] /*85640*/;
assign _7975_ = _7164_ & _7972_ /*85635*/;
assign _7976_ = _7164_ ^ _7972_ /*85638*/;
assign _7977_ = _7968_ & _7976_ /*85636*/;
assign _7612_ = _7968_ ^ _7976_ /*85637*/;
assign _7974_ = _7975_ | _7977_ /*85634*/;
assign _7979_ = ~Q[55] /*85633*/;
assign _7978_ = _7979_ & D[60] /*85632*/;
assign _7981_ = _7165_ & _7978_ /*85627*/;
assign _7982_ = _7165_ ^ _7978_ /*85630*/;
assign _7983_ = _7974_ & _7982_ /*85628*/;
assign _7613_ = _7974_ ^ _7982_ /*85629*/;
assign _7980_ = _7981_ | _7983_ /*85626*/;
assign _7985_ = ~Q[55] /*85625*/;
assign _7984_ = _7985_ & D[61] /*85624*/;
assign _7987_ = _7166_ & _7984_ /*85619*/;
assign _7988_ = _7166_ ^ _7984_ /*85622*/;
assign _7989_ = _7980_ & _7988_ /*85620*/;
assign _7614_ = _7980_ ^ _7988_ /*85621*/;
assign _7986_ = _7987_ | _7989_ /*85618*/;
assign _7991_ = ~Q[55] /*85617*/;
assign _7990_ = _7991_ & D[62] /*85616*/;
assign _7993_ = _7167_ & _7990_ /*85611*/;
assign _7994_ = _7167_ ^ _7990_ /*85614*/;
assign _7995_ = _7986_ & _7994_ /*85612*/;
assign _7615_ = _7986_ ^ _7994_ /*85613*/;
assign _7992_ = _7993_ | _7995_ /*85610*/;
assign _7997_ = ~Q[55] /*85609*/;
assign _7996_ = _7997_ & zeroWire /*85608*/;
assign _7998_ = _7168_ ^ _7996_ /*85606*/;
assign _7616_ = _7998_ ^ _7992_ /*85605*/;
assign _8069_ = ~D[0] /*85351*/;
assign _8066_ = R_0[54] & _8069_ /*85347*/;
assign _8067_ = R_0[54] ^ _8069_ /*85350*/;
assign _8068_ = oneWire & _8067_ /*85348*/;
assign _8001_ = oneWire ^ _8067_ /*85349*/;
assign _8065_ = _8066_ | _8068_ /*85346*/;
assign _8074_ = ~D[1] /*85345*/;
assign _8071_ = _7553_ & _8074_ /*85341*/;
assign _8072_ = _7553_ ^ _8074_ /*85344*/;
assign _8073_ = _8065_ & _8072_ /*85342*/;
assign _8002_ = _8065_ ^ _8072_ /*85343*/;
assign _8070_ = _8071_ | _8073_ /*85340*/;
assign _8079_ = ~D[2] /*85339*/;
assign _8076_ = _7554_ & _8079_ /*85335*/;
assign _8077_ = _7554_ ^ _8079_ /*85338*/;
assign _8078_ = _8070_ & _8077_ /*85336*/;
assign _8003_ = _8070_ ^ _8077_ /*85337*/;
assign _8075_ = _8076_ | _8078_ /*85334*/;
assign _8084_ = ~D[3] /*85333*/;
assign _8081_ = _7555_ & _8084_ /*85329*/;
assign _8082_ = _7555_ ^ _8084_ /*85332*/;
assign _8083_ = _8075_ & _8082_ /*85330*/;
assign _8004_ = _8075_ ^ _8082_ /*85331*/;
assign _8080_ = _8081_ | _8083_ /*85328*/;
assign _8089_ = ~D[4] /*85327*/;
assign _8086_ = _7556_ & _8089_ /*85323*/;
assign _8087_ = _7556_ ^ _8089_ /*85326*/;
assign _8088_ = _8080_ & _8087_ /*85324*/;
assign _8005_ = _8080_ ^ _8087_ /*85325*/;
assign _8085_ = _8086_ | _8088_ /*85322*/;
assign _8094_ = ~D[5] /*85321*/;
assign _8091_ = _7557_ & _8094_ /*85317*/;
assign _8092_ = _7557_ ^ _8094_ /*85320*/;
assign _8093_ = _8085_ & _8092_ /*85318*/;
assign _8006_ = _8085_ ^ _8092_ /*85319*/;
assign _8090_ = _8091_ | _8093_ /*85316*/;
assign _8099_ = ~D[6] /*85315*/;
assign _8096_ = _7558_ & _8099_ /*85311*/;
assign _8097_ = _7558_ ^ _8099_ /*85314*/;
assign _8098_ = _8090_ & _8097_ /*85312*/;
assign _8007_ = _8090_ ^ _8097_ /*85313*/;
assign _8095_ = _8096_ | _8098_ /*85310*/;
assign _8104_ = ~D[7] /*85309*/;
assign _8101_ = _7559_ & _8104_ /*85305*/;
assign _8102_ = _7559_ ^ _8104_ /*85308*/;
assign _8103_ = _8095_ & _8102_ /*85306*/;
assign _8008_ = _8095_ ^ _8102_ /*85307*/;
assign _8100_ = _8101_ | _8103_ /*85304*/;
assign _8109_ = ~D[8] /*85303*/;
assign _8106_ = _7560_ & _8109_ /*85299*/;
assign _8107_ = _7560_ ^ _8109_ /*85302*/;
assign _8108_ = _8100_ & _8107_ /*85300*/;
assign _8009_ = _8100_ ^ _8107_ /*85301*/;
assign _8105_ = _8106_ | _8108_ /*85298*/;
assign _8114_ = ~D[9] /*85297*/;
assign _8111_ = _7561_ & _8114_ /*85293*/;
assign _8112_ = _7561_ ^ _8114_ /*85296*/;
assign _8113_ = _8105_ & _8112_ /*85294*/;
assign _8010_ = _8105_ ^ _8112_ /*85295*/;
assign _8110_ = _8111_ | _8113_ /*85292*/;
assign _8119_ = ~D[10] /*85291*/;
assign _8116_ = _7562_ & _8119_ /*85287*/;
assign _8117_ = _7562_ ^ _8119_ /*85290*/;
assign _8118_ = _8110_ & _8117_ /*85288*/;
assign _8011_ = _8110_ ^ _8117_ /*85289*/;
assign _8115_ = _8116_ | _8118_ /*85286*/;
assign _8124_ = ~D[11] /*85285*/;
assign _8121_ = _7563_ & _8124_ /*85281*/;
assign _8122_ = _7563_ ^ _8124_ /*85284*/;
assign _8123_ = _8115_ & _8122_ /*85282*/;
assign _8012_ = _8115_ ^ _8122_ /*85283*/;
assign _8120_ = _8121_ | _8123_ /*85280*/;
assign _8129_ = ~D[12] /*85279*/;
assign _8126_ = _7564_ & _8129_ /*85275*/;
assign _8127_ = _7564_ ^ _8129_ /*85278*/;
assign _8128_ = _8120_ & _8127_ /*85276*/;
assign _8013_ = _8120_ ^ _8127_ /*85277*/;
assign _8125_ = _8126_ | _8128_ /*85274*/;
assign _8134_ = ~D[13] /*85273*/;
assign _8131_ = _7565_ & _8134_ /*85269*/;
assign _8132_ = _7565_ ^ _8134_ /*85272*/;
assign _8133_ = _8125_ & _8132_ /*85270*/;
assign _8014_ = _8125_ ^ _8132_ /*85271*/;
assign _8130_ = _8131_ | _8133_ /*85268*/;
assign _8139_ = ~D[14] /*85267*/;
assign _8136_ = _7566_ & _8139_ /*85263*/;
assign _8137_ = _7566_ ^ _8139_ /*85266*/;
assign _8138_ = _8130_ & _8137_ /*85264*/;
assign _8015_ = _8130_ ^ _8137_ /*85265*/;
assign _8135_ = _8136_ | _8138_ /*85262*/;
assign _8144_ = ~D[15] /*85261*/;
assign _8141_ = _7567_ & _8144_ /*85257*/;
assign _8142_ = _7567_ ^ _8144_ /*85260*/;
assign _8143_ = _8135_ & _8142_ /*85258*/;
assign _8016_ = _8135_ ^ _8142_ /*85259*/;
assign _8140_ = _8141_ | _8143_ /*85256*/;
assign _8149_ = ~D[16] /*85255*/;
assign _8146_ = _7568_ & _8149_ /*85251*/;
assign _8147_ = _7568_ ^ _8149_ /*85254*/;
assign _8148_ = _8140_ & _8147_ /*85252*/;
assign _8017_ = _8140_ ^ _8147_ /*85253*/;
assign _8145_ = _8146_ | _8148_ /*85250*/;
assign _8154_ = ~D[17] /*85249*/;
assign _8151_ = _7569_ & _8154_ /*85245*/;
assign _8152_ = _7569_ ^ _8154_ /*85248*/;
assign _8153_ = _8145_ & _8152_ /*85246*/;
assign _8018_ = _8145_ ^ _8152_ /*85247*/;
assign _8150_ = _8151_ | _8153_ /*85244*/;
assign _8159_ = ~D[18] /*85243*/;
assign _8156_ = _7570_ & _8159_ /*85239*/;
assign _8157_ = _7570_ ^ _8159_ /*85242*/;
assign _8158_ = _8150_ & _8157_ /*85240*/;
assign _8019_ = _8150_ ^ _8157_ /*85241*/;
assign _8155_ = _8156_ | _8158_ /*85238*/;
assign _8164_ = ~D[19] /*85237*/;
assign _8161_ = _7571_ & _8164_ /*85233*/;
assign _8162_ = _7571_ ^ _8164_ /*85236*/;
assign _8163_ = _8155_ & _8162_ /*85234*/;
assign _8020_ = _8155_ ^ _8162_ /*85235*/;
assign _8160_ = _8161_ | _8163_ /*85232*/;
assign _8169_ = ~D[20] /*85231*/;
assign _8166_ = _7572_ & _8169_ /*85227*/;
assign _8167_ = _7572_ ^ _8169_ /*85230*/;
assign _8168_ = _8160_ & _8167_ /*85228*/;
assign _8021_ = _8160_ ^ _8167_ /*85229*/;
assign _8165_ = _8166_ | _8168_ /*85226*/;
assign _8174_ = ~D[21] /*85225*/;
assign _8171_ = _7573_ & _8174_ /*85221*/;
assign _8172_ = _7573_ ^ _8174_ /*85224*/;
assign _8173_ = _8165_ & _8172_ /*85222*/;
assign _8022_ = _8165_ ^ _8172_ /*85223*/;
assign _8170_ = _8171_ | _8173_ /*85220*/;
assign _8179_ = ~D[22] /*85219*/;
assign _8176_ = _7574_ & _8179_ /*85215*/;
assign _8177_ = _7574_ ^ _8179_ /*85218*/;
assign _8178_ = _8170_ & _8177_ /*85216*/;
assign _8023_ = _8170_ ^ _8177_ /*85217*/;
assign _8175_ = _8176_ | _8178_ /*85214*/;
assign _8184_ = ~D[23] /*85213*/;
assign _8181_ = _7575_ & _8184_ /*85209*/;
assign _8182_ = _7575_ ^ _8184_ /*85212*/;
assign _8183_ = _8175_ & _8182_ /*85210*/;
assign _8024_ = _8175_ ^ _8182_ /*85211*/;
assign _8180_ = _8181_ | _8183_ /*85208*/;
assign _8189_ = ~D[24] /*85207*/;
assign _8186_ = _7576_ & _8189_ /*85203*/;
assign _8187_ = _7576_ ^ _8189_ /*85206*/;
assign _8188_ = _8180_ & _8187_ /*85204*/;
assign _8025_ = _8180_ ^ _8187_ /*85205*/;
assign _8185_ = _8186_ | _8188_ /*85202*/;
assign _8194_ = ~D[25] /*85201*/;
assign _8191_ = _7577_ & _8194_ /*85197*/;
assign _8192_ = _7577_ ^ _8194_ /*85200*/;
assign _8193_ = _8185_ & _8192_ /*85198*/;
assign _8026_ = _8185_ ^ _8192_ /*85199*/;
assign _8190_ = _8191_ | _8193_ /*85196*/;
assign _8199_ = ~D[26] /*85195*/;
assign _8196_ = _7578_ & _8199_ /*85191*/;
assign _8197_ = _7578_ ^ _8199_ /*85194*/;
assign _8198_ = _8190_ & _8197_ /*85192*/;
assign _8027_ = _8190_ ^ _8197_ /*85193*/;
assign _8195_ = _8196_ | _8198_ /*85190*/;
assign _8204_ = ~D[27] /*85189*/;
assign _8201_ = _7579_ & _8204_ /*85185*/;
assign _8202_ = _7579_ ^ _8204_ /*85188*/;
assign _8203_ = _8195_ & _8202_ /*85186*/;
assign _8028_ = _8195_ ^ _8202_ /*85187*/;
assign _8200_ = _8201_ | _8203_ /*85184*/;
assign _8209_ = ~D[28] /*85183*/;
assign _8206_ = _7580_ & _8209_ /*85179*/;
assign _8207_ = _7580_ ^ _8209_ /*85182*/;
assign _8208_ = _8200_ & _8207_ /*85180*/;
assign _8029_ = _8200_ ^ _8207_ /*85181*/;
assign _8205_ = _8206_ | _8208_ /*85178*/;
assign _8214_ = ~D[29] /*85177*/;
assign _8211_ = _7581_ & _8214_ /*85173*/;
assign _8212_ = _7581_ ^ _8214_ /*85176*/;
assign _8213_ = _8205_ & _8212_ /*85174*/;
assign _8030_ = _8205_ ^ _8212_ /*85175*/;
assign _8210_ = _8211_ | _8213_ /*85172*/;
assign _8219_ = ~D[30] /*85171*/;
assign _8216_ = _7582_ & _8219_ /*85167*/;
assign _8217_ = _7582_ ^ _8219_ /*85170*/;
assign _8218_ = _8210_ & _8217_ /*85168*/;
assign _8031_ = _8210_ ^ _8217_ /*85169*/;
assign _8215_ = _8216_ | _8218_ /*85166*/;
assign _8224_ = ~D[31] /*85165*/;
assign _8221_ = _7583_ & _8224_ /*85161*/;
assign _8222_ = _7583_ ^ _8224_ /*85164*/;
assign _8223_ = _8215_ & _8222_ /*85162*/;
assign _8032_ = _8215_ ^ _8222_ /*85163*/;
assign _8220_ = _8221_ | _8223_ /*85160*/;
assign _8229_ = ~D[32] /*85159*/;
assign _8226_ = _7584_ & _8229_ /*85155*/;
assign _8227_ = _7584_ ^ _8229_ /*85158*/;
assign _8228_ = _8220_ & _8227_ /*85156*/;
assign _8033_ = _8220_ ^ _8227_ /*85157*/;
assign _8225_ = _8226_ | _8228_ /*85154*/;
assign _8234_ = ~D[33] /*85153*/;
assign _8231_ = _7585_ & _8234_ /*85149*/;
assign _8232_ = _7585_ ^ _8234_ /*85152*/;
assign _8233_ = _8225_ & _8232_ /*85150*/;
assign _8034_ = _8225_ ^ _8232_ /*85151*/;
assign _8230_ = _8231_ | _8233_ /*85148*/;
assign _8239_ = ~D[34] /*85147*/;
assign _8236_ = _7586_ & _8239_ /*85143*/;
assign _8237_ = _7586_ ^ _8239_ /*85146*/;
assign _8238_ = _8230_ & _8237_ /*85144*/;
assign _8035_ = _8230_ ^ _8237_ /*85145*/;
assign _8235_ = _8236_ | _8238_ /*85142*/;
assign _8244_ = ~D[35] /*85141*/;
assign _8241_ = _7587_ & _8244_ /*85137*/;
assign _8242_ = _7587_ ^ _8244_ /*85140*/;
assign _8243_ = _8235_ & _8242_ /*85138*/;
assign _8036_ = _8235_ ^ _8242_ /*85139*/;
assign _8240_ = _8241_ | _8243_ /*85136*/;
assign _8249_ = ~D[36] /*85135*/;
assign _8246_ = _7588_ & _8249_ /*85131*/;
assign _8247_ = _7588_ ^ _8249_ /*85134*/;
assign _8248_ = _8240_ & _8247_ /*85132*/;
assign _8037_ = _8240_ ^ _8247_ /*85133*/;
assign _8245_ = _8246_ | _8248_ /*85130*/;
assign _8254_ = ~D[37] /*85129*/;
assign _8251_ = _7589_ & _8254_ /*85125*/;
assign _8252_ = _7589_ ^ _8254_ /*85128*/;
assign _8253_ = _8245_ & _8252_ /*85126*/;
assign _8038_ = _8245_ ^ _8252_ /*85127*/;
assign _8250_ = _8251_ | _8253_ /*85124*/;
assign _8259_ = ~D[38] /*85123*/;
assign _8256_ = _7590_ & _8259_ /*85119*/;
assign _8257_ = _7590_ ^ _8259_ /*85122*/;
assign _8258_ = _8250_ & _8257_ /*85120*/;
assign _8039_ = _8250_ ^ _8257_ /*85121*/;
assign _8255_ = _8256_ | _8258_ /*85118*/;
assign _8264_ = ~D[39] /*85117*/;
assign _8261_ = _7591_ & _8264_ /*85113*/;
assign _8262_ = _7591_ ^ _8264_ /*85116*/;
assign _8263_ = _8255_ & _8262_ /*85114*/;
assign _8040_ = _8255_ ^ _8262_ /*85115*/;
assign _8260_ = _8261_ | _8263_ /*85112*/;
assign _8269_ = ~D[40] /*85111*/;
assign _8266_ = _7592_ & _8269_ /*85107*/;
assign _8267_ = _7592_ ^ _8269_ /*85110*/;
assign _8268_ = _8260_ & _8267_ /*85108*/;
assign _8041_ = _8260_ ^ _8267_ /*85109*/;
assign _8265_ = _8266_ | _8268_ /*85106*/;
assign _8274_ = ~D[41] /*85105*/;
assign _8271_ = _7593_ & _8274_ /*85101*/;
assign _8272_ = _7593_ ^ _8274_ /*85104*/;
assign _8273_ = _8265_ & _8272_ /*85102*/;
assign _8042_ = _8265_ ^ _8272_ /*85103*/;
assign _8270_ = _8271_ | _8273_ /*85100*/;
assign _8279_ = ~D[42] /*85099*/;
assign _8276_ = _7594_ & _8279_ /*85095*/;
assign _8277_ = _7594_ ^ _8279_ /*85098*/;
assign _8278_ = _8270_ & _8277_ /*85096*/;
assign _8043_ = _8270_ ^ _8277_ /*85097*/;
assign _8275_ = _8276_ | _8278_ /*85094*/;
assign _8284_ = ~D[43] /*85093*/;
assign _8281_ = _7595_ & _8284_ /*85089*/;
assign _8282_ = _7595_ ^ _8284_ /*85092*/;
assign _8283_ = _8275_ & _8282_ /*85090*/;
assign _8044_ = _8275_ ^ _8282_ /*85091*/;
assign _8280_ = _8281_ | _8283_ /*85088*/;
assign _8289_ = ~D[44] /*85087*/;
assign _8286_ = _7596_ & _8289_ /*85083*/;
assign _8287_ = _7596_ ^ _8289_ /*85086*/;
assign _8288_ = _8280_ & _8287_ /*85084*/;
assign _8045_ = _8280_ ^ _8287_ /*85085*/;
assign _8285_ = _8286_ | _8288_ /*85082*/;
assign _8294_ = ~D[45] /*85081*/;
assign _8291_ = _7597_ & _8294_ /*85077*/;
assign _8292_ = _7597_ ^ _8294_ /*85080*/;
assign _8293_ = _8285_ & _8292_ /*85078*/;
assign _8046_ = _8285_ ^ _8292_ /*85079*/;
assign _8290_ = _8291_ | _8293_ /*85076*/;
assign _8299_ = ~D[46] /*85075*/;
assign _8296_ = _7598_ & _8299_ /*85071*/;
assign _8297_ = _7598_ ^ _8299_ /*85074*/;
assign _8298_ = _8290_ & _8297_ /*85072*/;
assign _8047_ = _8290_ ^ _8297_ /*85073*/;
assign _8295_ = _8296_ | _8298_ /*85070*/;
assign _8304_ = ~D[47] /*85069*/;
assign _8301_ = _7599_ & _8304_ /*85065*/;
assign _8302_ = _7599_ ^ _8304_ /*85068*/;
assign _8303_ = _8295_ & _8302_ /*85066*/;
assign _8048_ = _8295_ ^ _8302_ /*85067*/;
assign _8300_ = _8301_ | _8303_ /*85064*/;
assign _8309_ = ~D[48] /*85063*/;
assign _8306_ = _7600_ & _8309_ /*85059*/;
assign _8307_ = _7600_ ^ _8309_ /*85062*/;
assign _8308_ = _8300_ & _8307_ /*85060*/;
assign _8049_ = _8300_ ^ _8307_ /*85061*/;
assign _8305_ = _8306_ | _8308_ /*85058*/;
assign _8314_ = ~D[49] /*85057*/;
assign _8311_ = _7601_ & _8314_ /*85053*/;
assign _8312_ = _7601_ ^ _8314_ /*85056*/;
assign _8313_ = _8305_ & _8312_ /*85054*/;
assign _8050_ = _8305_ ^ _8312_ /*85055*/;
assign _8310_ = _8311_ | _8313_ /*85052*/;
assign _8319_ = ~D[50] /*85051*/;
assign _8316_ = _7602_ & _8319_ /*85047*/;
assign _8317_ = _7602_ ^ _8319_ /*85050*/;
assign _8318_ = _8310_ & _8317_ /*85048*/;
assign _8051_ = _8310_ ^ _8317_ /*85049*/;
assign _8315_ = _8316_ | _8318_ /*85046*/;
assign _8324_ = ~D[51] /*85045*/;
assign _8321_ = _7603_ & _8324_ /*85041*/;
assign _8322_ = _7603_ ^ _8324_ /*85044*/;
assign _8323_ = _8315_ & _8322_ /*85042*/;
assign _8052_ = _8315_ ^ _8322_ /*85043*/;
assign _8320_ = _8321_ | _8323_ /*85040*/;
assign _8329_ = ~D[52] /*85039*/;
assign _8326_ = _7604_ & _8329_ /*85035*/;
assign _8327_ = _7604_ ^ _8329_ /*85038*/;
assign _8328_ = _8320_ & _8327_ /*85036*/;
assign _8053_ = _8320_ ^ _8327_ /*85037*/;
assign _8325_ = _8326_ | _8328_ /*85034*/;
assign _8334_ = ~D[53] /*85033*/;
assign _8331_ = _7605_ & _8334_ /*85029*/;
assign _8332_ = _7605_ ^ _8334_ /*85032*/;
assign _8333_ = _8325_ & _8332_ /*85030*/;
assign _8054_ = _8325_ ^ _8332_ /*85031*/;
assign _8330_ = _8331_ | _8333_ /*85028*/;
assign _8339_ = ~D[54] /*85027*/;
assign _8336_ = _7606_ & _8339_ /*85023*/;
assign _8337_ = _7606_ ^ _8339_ /*85026*/;
assign _8338_ = _8330_ & _8337_ /*85024*/;
assign _8055_ = _8330_ ^ _8337_ /*85025*/;
assign _8335_ = _8336_ | _8338_ /*85022*/;
assign _8344_ = ~D[55] /*85021*/;
assign _8341_ = _7607_ & _8344_ /*85017*/;
assign _8342_ = _7607_ ^ _8344_ /*85020*/;
assign _8343_ = _8335_ & _8342_ /*85018*/;
assign _8056_ = _8335_ ^ _8342_ /*85019*/;
assign _8340_ = _8341_ | _8343_ /*85016*/;
assign _8349_ = ~D[56] /*85015*/;
assign _8346_ = _7608_ & _8349_ /*85011*/;
assign _8347_ = _7608_ ^ _8349_ /*85014*/;
assign _8348_ = _8340_ & _8347_ /*85012*/;
assign _8057_ = _8340_ ^ _8347_ /*85013*/;
assign _8345_ = _8346_ | _8348_ /*85010*/;
assign _8354_ = ~D[57] /*85009*/;
assign _8351_ = _7609_ & _8354_ /*85005*/;
assign _8352_ = _7609_ ^ _8354_ /*85008*/;
assign _8353_ = _8345_ & _8352_ /*85006*/;
assign _8058_ = _8345_ ^ _8352_ /*85007*/;
assign _8350_ = _8351_ | _8353_ /*85004*/;
assign _8359_ = ~D[58] /*85003*/;
assign _8356_ = _7610_ & _8359_ /*84999*/;
assign _8357_ = _7610_ ^ _8359_ /*85002*/;
assign _8358_ = _8350_ & _8357_ /*85000*/;
assign _8059_ = _8350_ ^ _8357_ /*85001*/;
assign _8355_ = _8356_ | _8358_ /*84998*/;
assign _8364_ = ~D[59] /*84997*/;
assign _8361_ = _7611_ & _8364_ /*84993*/;
assign _8362_ = _7611_ ^ _8364_ /*84996*/;
assign _8363_ = _8355_ & _8362_ /*84994*/;
assign _8060_ = _8355_ ^ _8362_ /*84995*/;
assign _8360_ = _8361_ | _8363_ /*84992*/;
assign _8369_ = ~D[60] /*84991*/;
assign _8366_ = _7612_ & _8369_ /*84987*/;
assign _8367_ = _7612_ ^ _8369_ /*84990*/;
assign _8368_ = _8360_ & _8367_ /*84988*/;
assign _8061_ = _8360_ ^ _8367_ /*84989*/;
assign _8365_ = _8366_ | _8368_ /*84986*/;
assign _8374_ = ~D[61] /*84985*/;
assign _8371_ = _7613_ & _8374_ /*84981*/;
assign _8372_ = _7613_ ^ _8374_ /*84984*/;
assign _8373_ = _8365_ & _8372_ /*84982*/;
assign _8062_ = _8365_ ^ _8372_ /*84983*/;
assign _8370_ = _8371_ | _8373_ /*84980*/;
assign _8379_ = ~D[62] /*84979*/;
assign _8376_ = _7614_ & _8379_ /*84975*/;
assign _8377_ = _7614_ ^ _8379_ /*84978*/;
assign _8378_ = _8370_ & _8377_ /*84976*/;
assign _8063_ = _8370_ ^ _8377_ /*84977*/;
assign _8375_ = _8376_ | _8378_ /*84974*/;
assign _8380_ = _7615_ & oneWire /*84969*/;
assign _8381_ = _7615_ ^ oneWire /*84972*/;
assign _8382_ = _8375_ & _8381_ /*84970*/;
assign _8064_ = _8375_ ^ _8381_ /*84971*/;
assign Q[54] = _8380_ | _8382_ /*84968*/;
assign _8515_ = ~Q[54] /*84583*/;
assign _8514_ = _8515_ & D[0] /*84582*/;
assign _8517_ = _8001_ & _8514_ /*84577*/;
assign _8518_ = _8001_ ^ _8514_ /*84580*/;
assign _8519_ = zeroWire & _8518_ /*84578*/;
assign _8449_ = zeroWire ^ _8518_ /*84579*/;
assign _8516_ = _8517_ | _8519_ /*84576*/;
assign _8521_ = ~Q[54] /*84575*/;
assign _8520_ = _8521_ & D[1] /*84574*/;
assign _8523_ = _8002_ & _8520_ /*84569*/;
assign _8524_ = _8002_ ^ _8520_ /*84572*/;
assign _8525_ = _8516_ & _8524_ /*84570*/;
assign _8450_ = _8516_ ^ _8524_ /*84571*/;
assign _8522_ = _8523_ | _8525_ /*84568*/;
assign _8527_ = ~Q[54] /*84567*/;
assign _8526_ = _8527_ & D[2] /*84566*/;
assign _8529_ = _8003_ & _8526_ /*84561*/;
assign _8530_ = _8003_ ^ _8526_ /*84564*/;
assign _8531_ = _8522_ & _8530_ /*84562*/;
assign _8451_ = _8522_ ^ _8530_ /*84563*/;
assign _8528_ = _8529_ | _8531_ /*84560*/;
assign _8533_ = ~Q[54] /*84559*/;
assign _8532_ = _8533_ & D[3] /*84558*/;
assign _8535_ = _8004_ & _8532_ /*84553*/;
assign _8536_ = _8004_ ^ _8532_ /*84556*/;
assign _8537_ = _8528_ & _8536_ /*84554*/;
assign _8452_ = _8528_ ^ _8536_ /*84555*/;
assign _8534_ = _8535_ | _8537_ /*84552*/;
assign _8539_ = ~Q[54] /*84551*/;
assign _8538_ = _8539_ & D[4] /*84550*/;
assign _8541_ = _8005_ & _8538_ /*84545*/;
assign _8542_ = _8005_ ^ _8538_ /*84548*/;
assign _8543_ = _8534_ & _8542_ /*84546*/;
assign _8453_ = _8534_ ^ _8542_ /*84547*/;
assign _8540_ = _8541_ | _8543_ /*84544*/;
assign _8545_ = ~Q[54] /*84543*/;
assign _8544_ = _8545_ & D[5] /*84542*/;
assign _8547_ = _8006_ & _8544_ /*84537*/;
assign _8548_ = _8006_ ^ _8544_ /*84540*/;
assign _8549_ = _8540_ & _8548_ /*84538*/;
assign _8454_ = _8540_ ^ _8548_ /*84539*/;
assign _8546_ = _8547_ | _8549_ /*84536*/;
assign _8551_ = ~Q[54] /*84535*/;
assign _8550_ = _8551_ & D[6] /*84534*/;
assign _8553_ = _8007_ & _8550_ /*84529*/;
assign _8554_ = _8007_ ^ _8550_ /*84532*/;
assign _8555_ = _8546_ & _8554_ /*84530*/;
assign _8455_ = _8546_ ^ _8554_ /*84531*/;
assign _8552_ = _8553_ | _8555_ /*84528*/;
assign _8557_ = ~Q[54] /*84527*/;
assign _8556_ = _8557_ & D[7] /*84526*/;
assign _8559_ = _8008_ & _8556_ /*84521*/;
assign _8560_ = _8008_ ^ _8556_ /*84524*/;
assign _8561_ = _8552_ & _8560_ /*84522*/;
assign _8456_ = _8552_ ^ _8560_ /*84523*/;
assign _8558_ = _8559_ | _8561_ /*84520*/;
assign _8563_ = ~Q[54] /*84519*/;
assign _8562_ = _8563_ & D[8] /*84518*/;
assign _8565_ = _8009_ & _8562_ /*84513*/;
assign _8566_ = _8009_ ^ _8562_ /*84516*/;
assign _8567_ = _8558_ & _8566_ /*84514*/;
assign _8457_ = _8558_ ^ _8566_ /*84515*/;
assign _8564_ = _8565_ | _8567_ /*84512*/;
assign _8569_ = ~Q[54] /*84511*/;
assign _8568_ = _8569_ & D[9] /*84510*/;
assign _8571_ = _8010_ & _8568_ /*84505*/;
assign _8572_ = _8010_ ^ _8568_ /*84508*/;
assign _8573_ = _8564_ & _8572_ /*84506*/;
assign _8458_ = _8564_ ^ _8572_ /*84507*/;
assign _8570_ = _8571_ | _8573_ /*84504*/;
assign _8575_ = ~Q[54] /*84503*/;
assign _8574_ = _8575_ & D[10] /*84502*/;
assign _8577_ = _8011_ & _8574_ /*84497*/;
assign _8578_ = _8011_ ^ _8574_ /*84500*/;
assign _8579_ = _8570_ & _8578_ /*84498*/;
assign _8459_ = _8570_ ^ _8578_ /*84499*/;
assign _8576_ = _8577_ | _8579_ /*84496*/;
assign _8581_ = ~Q[54] /*84495*/;
assign _8580_ = _8581_ & D[11] /*84494*/;
assign _8583_ = _8012_ & _8580_ /*84489*/;
assign _8584_ = _8012_ ^ _8580_ /*84492*/;
assign _8585_ = _8576_ & _8584_ /*84490*/;
assign _8460_ = _8576_ ^ _8584_ /*84491*/;
assign _8582_ = _8583_ | _8585_ /*84488*/;
assign _8587_ = ~Q[54] /*84487*/;
assign _8586_ = _8587_ & D[12] /*84486*/;
assign _8589_ = _8013_ & _8586_ /*84481*/;
assign _8590_ = _8013_ ^ _8586_ /*84484*/;
assign _8591_ = _8582_ & _8590_ /*84482*/;
assign _8461_ = _8582_ ^ _8590_ /*84483*/;
assign _8588_ = _8589_ | _8591_ /*84480*/;
assign _8593_ = ~Q[54] /*84479*/;
assign _8592_ = _8593_ & D[13] /*84478*/;
assign _8595_ = _8014_ & _8592_ /*84473*/;
assign _8596_ = _8014_ ^ _8592_ /*84476*/;
assign _8597_ = _8588_ & _8596_ /*84474*/;
assign _8462_ = _8588_ ^ _8596_ /*84475*/;
assign _8594_ = _8595_ | _8597_ /*84472*/;
assign _8599_ = ~Q[54] /*84471*/;
assign _8598_ = _8599_ & D[14] /*84470*/;
assign _8601_ = _8015_ & _8598_ /*84465*/;
assign _8602_ = _8015_ ^ _8598_ /*84468*/;
assign _8603_ = _8594_ & _8602_ /*84466*/;
assign _8463_ = _8594_ ^ _8602_ /*84467*/;
assign _8600_ = _8601_ | _8603_ /*84464*/;
assign _8605_ = ~Q[54] /*84463*/;
assign _8604_ = _8605_ & D[15] /*84462*/;
assign _8607_ = _8016_ & _8604_ /*84457*/;
assign _8608_ = _8016_ ^ _8604_ /*84460*/;
assign _8609_ = _8600_ & _8608_ /*84458*/;
assign _8464_ = _8600_ ^ _8608_ /*84459*/;
assign _8606_ = _8607_ | _8609_ /*84456*/;
assign _8611_ = ~Q[54] /*84455*/;
assign _8610_ = _8611_ & D[16] /*84454*/;
assign _8613_ = _8017_ & _8610_ /*84449*/;
assign _8614_ = _8017_ ^ _8610_ /*84452*/;
assign _8615_ = _8606_ & _8614_ /*84450*/;
assign _8465_ = _8606_ ^ _8614_ /*84451*/;
assign _8612_ = _8613_ | _8615_ /*84448*/;
assign _8617_ = ~Q[54] /*84447*/;
assign _8616_ = _8617_ & D[17] /*84446*/;
assign _8619_ = _8018_ & _8616_ /*84441*/;
assign _8620_ = _8018_ ^ _8616_ /*84444*/;
assign _8621_ = _8612_ & _8620_ /*84442*/;
assign _8466_ = _8612_ ^ _8620_ /*84443*/;
assign _8618_ = _8619_ | _8621_ /*84440*/;
assign _8623_ = ~Q[54] /*84439*/;
assign _8622_ = _8623_ & D[18] /*84438*/;
assign _8625_ = _8019_ & _8622_ /*84433*/;
assign _8626_ = _8019_ ^ _8622_ /*84436*/;
assign _8627_ = _8618_ & _8626_ /*84434*/;
assign _8467_ = _8618_ ^ _8626_ /*84435*/;
assign _8624_ = _8625_ | _8627_ /*84432*/;
assign _8629_ = ~Q[54] /*84431*/;
assign _8628_ = _8629_ & D[19] /*84430*/;
assign _8631_ = _8020_ & _8628_ /*84425*/;
assign _8632_ = _8020_ ^ _8628_ /*84428*/;
assign _8633_ = _8624_ & _8632_ /*84426*/;
assign _8468_ = _8624_ ^ _8632_ /*84427*/;
assign _8630_ = _8631_ | _8633_ /*84424*/;
assign _8635_ = ~Q[54] /*84423*/;
assign _8634_ = _8635_ & D[20] /*84422*/;
assign _8637_ = _8021_ & _8634_ /*84417*/;
assign _8638_ = _8021_ ^ _8634_ /*84420*/;
assign _8639_ = _8630_ & _8638_ /*84418*/;
assign _8469_ = _8630_ ^ _8638_ /*84419*/;
assign _8636_ = _8637_ | _8639_ /*84416*/;
assign _8641_ = ~Q[54] /*84415*/;
assign _8640_ = _8641_ & D[21] /*84414*/;
assign _8643_ = _8022_ & _8640_ /*84409*/;
assign _8644_ = _8022_ ^ _8640_ /*84412*/;
assign _8645_ = _8636_ & _8644_ /*84410*/;
assign _8470_ = _8636_ ^ _8644_ /*84411*/;
assign _8642_ = _8643_ | _8645_ /*84408*/;
assign _8647_ = ~Q[54] /*84407*/;
assign _8646_ = _8647_ & D[22] /*84406*/;
assign _8649_ = _8023_ & _8646_ /*84401*/;
assign _8650_ = _8023_ ^ _8646_ /*84404*/;
assign _8651_ = _8642_ & _8650_ /*84402*/;
assign _8471_ = _8642_ ^ _8650_ /*84403*/;
assign _8648_ = _8649_ | _8651_ /*84400*/;
assign _8653_ = ~Q[54] /*84399*/;
assign _8652_ = _8653_ & D[23] /*84398*/;
assign _8655_ = _8024_ & _8652_ /*84393*/;
assign _8656_ = _8024_ ^ _8652_ /*84396*/;
assign _8657_ = _8648_ & _8656_ /*84394*/;
assign _8472_ = _8648_ ^ _8656_ /*84395*/;
assign _8654_ = _8655_ | _8657_ /*84392*/;
assign _8659_ = ~Q[54] /*84391*/;
assign _8658_ = _8659_ & D[24] /*84390*/;
assign _8661_ = _8025_ & _8658_ /*84385*/;
assign _8662_ = _8025_ ^ _8658_ /*84388*/;
assign _8663_ = _8654_ & _8662_ /*84386*/;
assign _8473_ = _8654_ ^ _8662_ /*84387*/;
assign _8660_ = _8661_ | _8663_ /*84384*/;
assign _8665_ = ~Q[54] /*84383*/;
assign _8664_ = _8665_ & D[25] /*84382*/;
assign _8667_ = _8026_ & _8664_ /*84377*/;
assign _8668_ = _8026_ ^ _8664_ /*84380*/;
assign _8669_ = _8660_ & _8668_ /*84378*/;
assign _8474_ = _8660_ ^ _8668_ /*84379*/;
assign _8666_ = _8667_ | _8669_ /*84376*/;
assign _8671_ = ~Q[54] /*84375*/;
assign _8670_ = _8671_ & D[26] /*84374*/;
assign _8673_ = _8027_ & _8670_ /*84369*/;
assign _8674_ = _8027_ ^ _8670_ /*84372*/;
assign _8675_ = _8666_ & _8674_ /*84370*/;
assign _8475_ = _8666_ ^ _8674_ /*84371*/;
assign _8672_ = _8673_ | _8675_ /*84368*/;
assign _8677_ = ~Q[54] /*84367*/;
assign _8676_ = _8677_ & D[27] /*84366*/;
assign _8679_ = _8028_ & _8676_ /*84361*/;
assign _8680_ = _8028_ ^ _8676_ /*84364*/;
assign _8681_ = _8672_ & _8680_ /*84362*/;
assign _8476_ = _8672_ ^ _8680_ /*84363*/;
assign _8678_ = _8679_ | _8681_ /*84360*/;
assign _8683_ = ~Q[54] /*84359*/;
assign _8682_ = _8683_ & D[28] /*84358*/;
assign _8685_ = _8029_ & _8682_ /*84353*/;
assign _8686_ = _8029_ ^ _8682_ /*84356*/;
assign _8687_ = _8678_ & _8686_ /*84354*/;
assign _8477_ = _8678_ ^ _8686_ /*84355*/;
assign _8684_ = _8685_ | _8687_ /*84352*/;
assign _8689_ = ~Q[54] /*84351*/;
assign _8688_ = _8689_ & D[29] /*84350*/;
assign _8691_ = _8030_ & _8688_ /*84345*/;
assign _8692_ = _8030_ ^ _8688_ /*84348*/;
assign _8693_ = _8684_ & _8692_ /*84346*/;
assign _8478_ = _8684_ ^ _8692_ /*84347*/;
assign _8690_ = _8691_ | _8693_ /*84344*/;
assign _8695_ = ~Q[54] /*84343*/;
assign _8694_ = _8695_ & D[30] /*84342*/;
assign _8697_ = _8031_ & _8694_ /*84337*/;
assign _8698_ = _8031_ ^ _8694_ /*84340*/;
assign _8699_ = _8690_ & _8698_ /*84338*/;
assign _8479_ = _8690_ ^ _8698_ /*84339*/;
assign _8696_ = _8697_ | _8699_ /*84336*/;
assign _8701_ = ~Q[54] /*84335*/;
assign _8700_ = _8701_ & D[31] /*84334*/;
assign _8703_ = _8032_ & _8700_ /*84329*/;
assign _8704_ = _8032_ ^ _8700_ /*84332*/;
assign _8705_ = _8696_ & _8704_ /*84330*/;
assign _8480_ = _8696_ ^ _8704_ /*84331*/;
assign _8702_ = _8703_ | _8705_ /*84328*/;
assign _8707_ = ~Q[54] /*84327*/;
assign _8706_ = _8707_ & D[32] /*84326*/;
assign _8709_ = _8033_ & _8706_ /*84321*/;
assign _8710_ = _8033_ ^ _8706_ /*84324*/;
assign _8711_ = _8702_ & _8710_ /*84322*/;
assign _8481_ = _8702_ ^ _8710_ /*84323*/;
assign _8708_ = _8709_ | _8711_ /*84320*/;
assign _8713_ = ~Q[54] /*84319*/;
assign _8712_ = _8713_ & D[33] /*84318*/;
assign _8715_ = _8034_ & _8712_ /*84313*/;
assign _8716_ = _8034_ ^ _8712_ /*84316*/;
assign _8717_ = _8708_ & _8716_ /*84314*/;
assign _8482_ = _8708_ ^ _8716_ /*84315*/;
assign _8714_ = _8715_ | _8717_ /*84312*/;
assign _8719_ = ~Q[54] /*84311*/;
assign _8718_ = _8719_ & D[34] /*84310*/;
assign _8721_ = _8035_ & _8718_ /*84305*/;
assign _8722_ = _8035_ ^ _8718_ /*84308*/;
assign _8723_ = _8714_ & _8722_ /*84306*/;
assign _8483_ = _8714_ ^ _8722_ /*84307*/;
assign _8720_ = _8721_ | _8723_ /*84304*/;
assign _8725_ = ~Q[54] /*84303*/;
assign _8724_ = _8725_ & D[35] /*84302*/;
assign _8727_ = _8036_ & _8724_ /*84297*/;
assign _8728_ = _8036_ ^ _8724_ /*84300*/;
assign _8729_ = _8720_ & _8728_ /*84298*/;
assign _8484_ = _8720_ ^ _8728_ /*84299*/;
assign _8726_ = _8727_ | _8729_ /*84296*/;
assign _8731_ = ~Q[54] /*84295*/;
assign _8730_ = _8731_ & D[36] /*84294*/;
assign _8733_ = _8037_ & _8730_ /*84289*/;
assign _8734_ = _8037_ ^ _8730_ /*84292*/;
assign _8735_ = _8726_ & _8734_ /*84290*/;
assign _8485_ = _8726_ ^ _8734_ /*84291*/;
assign _8732_ = _8733_ | _8735_ /*84288*/;
assign _8737_ = ~Q[54] /*84287*/;
assign _8736_ = _8737_ & D[37] /*84286*/;
assign _8739_ = _8038_ & _8736_ /*84281*/;
assign _8740_ = _8038_ ^ _8736_ /*84284*/;
assign _8741_ = _8732_ & _8740_ /*84282*/;
assign _8486_ = _8732_ ^ _8740_ /*84283*/;
assign _8738_ = _8739_ | _8741_ /*84280*/;
assign _8743_ = ~Q[54] /*84279*/;
assign _8742_ = _8743_ & D[38] /*84278*/;
assign _8745_ = _8039_ & _8742_ /*84273*/;
assign _8746_ = _8039_ ^ _8742_ /*84276*/;
assign _8747_ = _8738_ & _8746_ /*84274*/;
assign _8487_ = _8738_ ^ _8746_ /*84275*/;
assign _8744_ = _8745_ | _8747_ /*84272*/;
assign _8749_ = ~Q[54] /*84271*/;
assign _8748_ = _8749_ & D[39] /*84270*/;
assign _8751_ = _8040_ & _8748_ /*84265*/;
assign _8752_ = _8040_ ^ _8748_ /*84268*/;
assign _8753_ = _8744_ & _8752_ /*84266*/;
assign _8488_ = _8744_ ^ _8752_ /*84267*/;
assign _8750_ = _8751_ | _8753_ /*84264*/;
assign _8755_ = ~Q[54] /*84263*/;
assign _8754_ = _8755_ & D[40] /*84262*/;
assign _8757_ = _8041_ & _8754_ /*84257*/;
assign _8758_ = _8041_ ^ _8754_ /*84260*/;
assign _8759_ = _8750_ & _8758_ /*84258*/;
assign _8489_ = _8750_ ^ _8758_ /*84259*/;
assign _8756_ = _8757_ | _8759_ /*84256*/;
assign _8761_ = ~Q[54] /*84255*/;
assign _8760_ = _8761_ & D[41] /*84254*/;
assign _8763_ = _8042_ & _8760_ /*84249*/;
assign _8764_ = _8042_ ^ _8760_ /*84252*/;
assign _8765_ = _8756_ & _8764_ /*84250*/;
assign _8490_ = _8756_ ^ _8764_ /*84251*/;
assign _8762_ = _8763_ | _8765_ /*84248*/;
assign _8767_ = ~Q[54] /*84247*/;
assign _8766_ = _8767_ & D[42] /*84246*/;
assign _8769_ = _8043_ & _8766_ /*84241*/;
assign _8770_ = _8043_ ^ _8766_ /*84244*/;
assign _8771_ = _8762_ & _8770_ /*84242*/;
assign _8491_ = _8762_ ^ _8770_ /*84243*/;
assign _8768_ = _8769_ | _8771_ /*84240*/;
assign _8773_ = ~Q[54] /*84239*/;
assign _8772_ = _8773_ & D[43] /*84238*/;
assign _8775_ = _8044_ & _8772_ /*84233*/;
assign _8776_ = _8044_ ^ _8772_ /*84236*/;
assign _8777_ = _8768_ & _8776_ /*84234*/;
assign _8492_ = _8768_ ^ _8776_ /*84235*/;
assign _8774_ = _8775_ | _8777_ /*84232*/;
assign _8779_ = ~Q[54] /*84231*/;
assign _8778_ = _8779_ & D[44] /*84230*/;
assign _8781_ = _8045_ & _8778_ /*84225*/;
assign _8782_ = _8045_ ^ _8778_ /*84228*/;
assign _8783_ = _8774_ & _8782_ /*84226*/;
assign _8493_ = _8774_ ^ _8782_ /*84227*/;
assign _8780_ = _8781_ | _8783_ /*84224*/;
assign _8785_ = ~Q[54] /*84223*/;
assign _8784_ = _8785_ & D[45] /*84222*/;
assign _8787_ = _8046_ & _8784_ /*84217*/;
assign _8788_ = _8046_ ^ _8784_ /*84220*/;
assign _8789_ = _8780_ & _8788_ /*84218*/;
assign _8494_ = _8780_ ^ _8788_ /*84219*/;
assign _8786_ = _8787_ | _8789_ /*84216*/;
assign _8791_ = ~Q[54] /*84215*/;
assign _8790_ = _8791_ & D[46] /*84214*/;
assign _8793_ = _8047_ & _8790_ /*84209*/;
assign _8794_ = _8047_ ^ _8790_ /*84212*/;
assign _8795_ = _8786_ & _8794_ /*84210*/;
assign _8495_ = _8786_ ^ _8794_ /*84211*/;
assign _8792_ = _8793_ | _8795_ /*84208*/;
assign _8797_ = ~Q[54] /*84207*/;
assign _8796_ = _8797_ & D[47] /*84206*/;
assign _8799_ = _8048_ & _8796_ /*84201*/;
assign _8800_ = _8048_ ^ _8796_ /*84204*/;
assign _8801_ = _8792_ & _8800_ /*84202*/;
assign _8496_ = _8792_ ^ _8800_ /*84203*/;
assign _8798_ = _8799_ | _8801_ /*84200*/;
assign _8803_ = ~Q[54] /*84199*/;
assign _8802_ = _8803_ & D[48] /*84198*/;
assign _8805_ = _8049_ & _8802_ /*84193*/;
assign _8806_ = _8049_ ^ _8802_ /*84196*/;
assign _8807_ = _8798_ & _8806_ /*84194*/;
assign _8497_ = _8798_ ^ _8806_ /*84195*/;
assign _8804_ = _8805_ | _8807_ /*84192*/;
assign _8809_ = ~Q[54] /*84191*/;
assign _8808_ = _8809_ & D[49] /*84190*/;
assign _8811_ = _8050_ & _8808_ /*84185*/;
assign _8812_ = _8050_ ^ _8808_ /*84188*/;
assign _8813_ = _8804_ & _8812_ /*84186*/;
assign _8498_ = _8804_ ^ _8812_ /*84187*/;
assign _8810_ = _8811_ | _8813_ /*84184*/;
assign _8815_ = ~Q[54] /*84183*/;
assign _8814_ = _8815_ & D[50] /*84182*/;
assign _8817_ = _8051_ & _8814_ /*84177*/;
assign _8818_ = _8051_ ^ _8814_ /*84180*/;
assign _8819_ = _8810_ & _8818_ /*84178*/;
assign _8499_ = _8810_ ^ _8818_ /*84179*/;
assign _8816_ = _8817_ | _8819_ /*84176*/;
assign _8821_ = ~Q[54] /*84175*/;
assign _8820_ = _8821_ & D[51] /*84174*/;
assign _8823_ = _8052_ & _8820_ /*84169*/;
assign _8824_ = _8052_ ^ _8820_ /*84172*/;
assign _8825_ = _8816_ & _8824_ /*84170*/;
assign _8500_ = _8816_ ^ _8824_ /*84171*/;
assign _8822_ = _8823_ | _8825_ /*84168*/;
assign _8827_ = ~Q[54] /*84167*/;
assign _8826_ = _8827_ & D[52] /*84166*/;
assign _8829_ = _8053_ & _8826_ /*84161*/;
assign _8830_ = _8053_ ^ _8826_ /*84164*/;
assign _8831_ = _8822_ & _8830_ /*84162*/;
assign _8501_ = _8822_ ^ _8830_ /*84163*/;
assign _8828_ = _8829_ | _8831_ /*84160*/;
assign _8833_ = ~Q[54] /*84159*/;
assign _8832_ = _8833_ & D[53] /*84158*/;
assign _8835_ = _8054_ & _8832_ /*84153*/;
assign _8836_ = _8054_ ^ _8832_ /*84156*/;
assign _8837_ = _8828_ & _8836_ /*84154*/;
assign _8502_ = _8828_ ^ _8836_ /*84155*/;
assign _8834_ = _8835_ | _8837_ /*84152*/;
assign _8839_ = ~Q[54] /*84151*/;
assign _8838_ = _8839_ & D[54] /*84150*/;
assign _8841_ = _8055_ & _8838_ /*84145*/;
assign _8842_ = _8055_ ^ _8838_ /*84148*/;
assign _8843_ = _8834_ & _8842_ /*84146*/;
assign _8503_ = _8834_ ^ _8842_ /*84147*/;
assign _8840_ = _8841_ | _8843_ /*84144*/;
assign _8845_ = ~Q[54] /*84143*/;
assign _8844_ = _8845_ & D[55] /*84142*/;
assign _8847_ = _8056_ & _8844_ /*84137*/;
assign _8848_ = _8056_ ^ _8844_ /*84140*/;
assign _8849_ = _8840_ & _8848_ /*84138*/;
assign _8504_ = _8840_ ^ _8848_ /*84139*/;
assign _8846_ = _8847_ | _8849_ /*84136*/;
assign _8851_ = ~Q[54] /*84135*/;
assign _8850_ = _8851_ & D[56] /*84134*/;
assign _8853_ = _8057_ & _8850_ /*84129*/;
assign _8854_ = _8057_ ^ _8850_ /*84132*/;
assign _8855_ = _8846_ & _8854_ /*84130*/;
assign _8505_ = _8846_ ^ _8854_ /*84131*/;
assign _8852_ = _8853_ | _8855_ /*84128*/;
assign _8857_ = ~Q[54] /*84127*/;
assign _8856_ = _8857_ & D[57] /*84126*/;
assign _8859_ = _8058_ & _8856_ /*84121*/;
assign _8860_ = _8058_ ^ _8856_ /*84124*/;
assign _8861_ = _8852_ & _8860_ /*84122*/;
assign _8506_ = _8852_ ^ _8860_ /*84123*/;
assign _8858_ = _8859_ | _8861_ /*84120*/;
assign _8863_ = ~Q[54] /*84119*/;
assign _8862_ = _8863_ & D[58] /*84118*/;
assign _8865_ = _8059_ & _8862_ /*84113*/;
assign _8866_ = _8059_ ^ _8862_ /*84116*/;
assign _8867_ = _8858_ & _8866_ /*84114*/;
assign _8507_ = _8858_ ^ _8866_ /*84115*/;
assign _8864_ = _8865_ | _8867_ /*84112*/;
assign _8869_ = ~Q[54] /*84111*/;
assign _8868_ = _8869_ & D[59] /*84110*/;
assign _8871_ = _8060_ & _8868_ /*84105*/;
assign _8872_ = _8060_ ^ _8868_ /*84108*/;
assign _8873_ = _8864_ & _8872_ /*84106*/;
assign _8508_ = _8864_ ^ _8872_ /*84107*/;
assign _8870_ = _8871_ | _8873_ /*84104*/;
assign _8875_ = ~Q[54] /*84103*/;
assign _8874_ = _8875_ & D[60] /*84102*/;
assign _8877_ = _8061_ & _8874_ /*84097*/;
assign _8878_ = _8061_ ^ _8874_ /*84100*/;
assign _8879_ = _8870_ & _8878_ /*84098*/;
assign _8509_ = _8870_ ^ _8878_ /*84099*/;
assign _8876_ = _8877_ | _8879_ /*84096*/;
assign _8881_ = ~Q[54] /*84095*/;
assign _8880_ = _8881_ & D[61] /*84094*/;
assign _8883_ = _8062_ & _8880_ /*84089*/;
assign _8884_ = _8062_ ^ _8880_ /*84092*/;
assign _8885_ = _8876_ & _8884_ /*84090*/;
assign _8510_ = _8876_ ^ _8884_ /*84091*/;
assign _8882_ = _8883_ | _8885_ /*84088*/;
assign _8887_ = ~Q[54] /*84087*/;
assign _8886_ = _8887_ & D[62] /*84086*/;
assign _8889_ = _8063_ & _8886_ /*84081*/;
assign _8890_ = _8063_ ^ _8886_ /*84084*/;
assign _8891_ = _8882_ & _8890_ /*84082*/;
assign _8511_ = _8882_ ^ _8890_ /*84083*/;
assign _8888_ = _8889_ | _8891_ /*84080*/;
assign _8893_ = ~Q[54] /*84079*/;
assign _8892_ = _8893_ & zeroWire /*84078*/;
assign _8894_ = _8064_ ^ _8892_ /*84076*/;
assign _8512_ = _8894_ ^ _8888_ /*84075*/;
assign _8965_ = ~D[0] /*83821*/;
assign _8962_ = R_0[53] & _8965_ /*83817*/;
assign _8963_ = R_0[53] ^ _8965_ /*83820*/;
assign _8964_ = oneWire & _8963_ /*83818*/;
assign _8897_ = oneWire ^ _8963_ /*83819*/;
assign _8961_ = _8962_ | _8964_ /*83816*/;
assign _8970_ = ~D[1] /*83815*/;
assign _8967_ = _8449_ & _8970_ /*83811*/;
assign _8968_ = _8449_ ^ _8970_ /*83814*/;
assign _8969_ = _8961_ & _8968_ /*83812*/;
assign _8898_ = _8961_ ^ _8968_ /*83813*/;
assign _8966_ = _8967_ | _8969_ /*83810*/;
assign _8975_ = ~D[2] /*83809*/;
assign _8972_ = _8450_ & _8975_ /*83805*/;
assign _8973_ = _8450_ ^ _8975_ /*83808*/;
assign _8974_ = _8966_ & _8973_ /*83806*/;
assign _8899_ = _8966_ ^ _8973_ /*83807*/;
assign _8971_ = _8972_ | _8974_ /*83804*/;
assign _8980_ = ~D[3] /*83803*/;
assign _8977_ = _8451_ & _8980_ /*83799*/;
assign _8978_ = _8451_ ^ _8980_ /*83802*/;
assign _8979_ = _8971_ & _8978_ /*83800*/;
assign _8900_ = _8971_ ^ _8978_ /*83801*/;
assign _8976_ = _8977_ | _8979_ /*83798*/;
assign _8985_ = ~D[4] /*83797*/;
assign _8982_ = _8452_ & _8985_ /*83793*/;
assign _8983_ = _8452_ ^ _8985_ /*83796*/;
assign _8984_ = _8976_ & _8983_ /*83794*/;
assign _8901_ = _8976_ ^ _8983_ /*83795*/;
assign _8981_ = _8982_ | _8984_ /*83792*/;
assign _8990_ = ~D[5] /*83791*/;
assign _8987_ = _8453_ & _8990_ /*83787*/;
assign _8988_ = _8453_ ^ _8990_ /*83790*/;
assign _8989_ = _8981_ & _8988_ /*83788*/;
assign _8902_ = _8981_ ^ _8988_ /*83789*/;
assign _8986_ = _8987_ | _8989_ /*83786*/;
assign _8995_ = ~D[6] /*83785*/;
assign _8992_ = _8454_ & _8995_ /*83781*/;
assign _8993_ = _8454_ ^ _8995_ /*83784*/;
assign _8994_ = _8986_ & _8993_ /*83782*/;
assign _8903_ = _8986_ ^ _8993_ /*83783*/;
assign _8991_ = _8992_ | _8994_ /*83780*/;
assign _9000_ = ~D[7] /*83779*/;
assign _8997_ = _8455_ & _9000_ /*83775*/;
assign _8998_ = _8455_ ^ _9000_ /*83778*/;
assign _8999_ = _8991_ & _8998_ /*83776*/;
assign _8904_ = _8991_ ^ _8998_ /*83777*/;
assign _8996_ = _8997_ | _8999_ /*83774*/;
assign _9005_ = ~D[8] /*83773*/;
assign _9002_ = _8456_ & _9005_ /*83769*/;
assign _9003_ = _8456_ ^ _9005_ /*83772*/;
assign _9004_ = _8996_ & _9003_ /*83770*/;
assign _8905_ = _8996_ ^ _9003_ /*83771*/;
assign _9001_ = _9002_ | _9004_ /*83768*/;
assign _9010_ = ~D[9] /*83767*/;
assign _9007_ = _8457_ & _9010_ /*83763*/;
assign _9008_ = _8457_ ^ _9010_ /*83766*/;
assign _9009_ = _9001_ & _9008_ /*83764*/;
assign _8906_ = _9001_ ^ _9008_ /*83765*/;
assign _9006_ = _9007_ | _9009_ /*83762*/;
assign _9015_ = ~D[10] /*83761*/;
assign _9012_ = _8458_ & _9015_ /*83757*/;
assign _9013_ = _8458_ ^ _9015_ /*83760*/;
assign _9014_ = _9006_ & _9013_ /*83758*/;
assign _8907_ = _9006_ ^ _9013_ /*83759*/;
assign _9011_ = _9012_ | _9014_ /*83756*/;
assign _9020_ = ~D[11] /*83755*/;
assign _9017_ = _8459_ & _9020_ /*83751*/;
assign _9018_ = _8459_ ^ _9020_ /*83754*/;
assign _9019_ = _9011_ & _9018_ /*83752*/;
assign _8908_ = _9011_ ^ _9018_ /*83753*/;
assign _9016_ = _9017_ | _9019_ /*83750*/;
assign _9025_ = ~D[12] /*83749*/;
assign _9022_ = _8460_ & _9025_ /*83745*/;
assign _9023_ = _8460_ ^ _9025_ /*83748*/;
assign _9024_ = _9016_ & _9023_ /*83746*/;
assign _8909_ = _9016_ ^ _9023_ /*83747*/;
assign _9021_ = _9022_ | _9024_ /*83744*/;
assign _9030_ = ~D[13] /*83743*/;
assign _9027_ = _8461_ & _9030_ /*83739*/;
assign _9028_ = _8461_ ^ _9030_ /*83742*/;
assign _9029_ = _9021_ & _9028_ /*83740*/;
assign _8910_ = _9021_ ^ _9028_ /*83741*/;
assign _9026_ = _9027_ | _9029_ /*83738*/;
assign _9035_ = ~D[14] /*83737*/;
assign _9032_ = _8462_ & _9035_ /*83733*/;
assign _9033_ = _8462_ ^ _9035_ /*83736*/;
assign _9034_ = _9026_ & _9033_ /*83734*/;
assign _8911_ = _9026_ ^ _9033_ /*83735*/;
assign _9031_ = _9032_ | _9034_ /*83732*/;
assign _9040_ = ~D[15] /*83731*/;
assign _9037_ = _8463_ & _9040_ /*83727*/;
assign _9038_ = _8463_ ^ _9040_ /*83730*/;
assign _9039_ = _9031_ & _9038_ /*83728*/;
assign _8912_ = _9031_ ^ _9038_ /*83729*/;
assign _9036_ = _9037_ | _9039_ /*83726*/;
assign _9045_ = ~D[16] /*83725*/;
assign _9042_ = _8464_ & _9045_ /*83721*/;
assign _9043_ = _8464_ ^ _9045_ /*83724*/;
assign _9044_ = _9036_ & _9043_ /*83722*/;
assign _8913_ = _9036_ ^ _9043_ /*83723*/;
assign _9041_ = _9042_ | _9044_ /*83720*/;
assign _9050_ = ~D[17] /*83719*/;
assign _9047_ = _8465_ & _9050_ /*83715*/;
assign _9048_ = _8465_ ^ _9050_ /*83718*/;
assign _9049_ = _9041_ & _9048_ /*83716*/;
assign _8914_ = _9041_ ^ _9048_ /*83717*/;
assign _9046_ = _9047_ | _9049_ /*83714*/;
assign _9055_ = ~D[18] /*83713*/;
assign _9052_ = _8466_ & _9055_ /*83709*/;
assign _9053_ = _8466_ ^ _9055_ /*83712*/;
assign _9054_ = _9046_ & _9053_ /*83710*/;
assign _8915_ = _9046_ ^ _9053_ /*83711*/;
assign _9051_ = _9052_ | _9054_ /*83708*/;
assign _9060_ = ~D[19] /*83707*/;
assign _9057_ = _8467_ & _9060_ /*83703*/;
assign _9058_ = _8467_ ^ _9060_ /*83706*/;
assign _9059_ = _9051_ & _9058_ /*83704*/;
assign _8916_ = _9051_ ^ _9058_ /*83705*/;
assign _9056_ = _9057_ | _9059_ /*83702*/;
assign _9065_ = ~D[20] /*83701*/;
assign _9062_ = _8468_ & _9065_ /*83697*/;
assign _9063_ = _8468_ ^ _9065_ /*83700*/;
assign _9064_ = _9056_ & _9063_ /*83698*/;
assign _8917_ = _9056_ ^ _9063_ /*83699*/;
assign _9061_ = _9062_ | _9064_ /*83696*/;
assign _9070_ = ~D[21] /*83695*/;
assign _9067_ = _8469_ & _9070_ /*83691*/;
assign _9068_ = _8469_ ^ _9070_ /*83694*/;
assign _9069_ = _9061_ & _9068_ /*83692*/;
assign _8918_ = _9061_ ^ _9068_ /*83693*/;
assign _9066_ = _9067_ | _9069_ /*83690*/;
assign _9075_ = ~D[22] /*83689*/;
assign _9072_ = _8470_ & _9075_ /*83685*/;
assign _9073_ = _8470_ ^ _9075_ /*83688*/;
assign _9074_ = _9066_ & _9073_ /*83686*/;
assign _8919_ = _9066_ ^ _9073_ /*83687*/;
assign _9071_ = _9072_ | _9074_ /*83684*/;
assign _9080_ = ~D[23] /*83683*/;
assign _9077_ = _8471_ & _9080_ /*83679*/;
assign _9078_ = _8471_ ^ _9080_ /*83682*/;
assign _9079_ = _9071_ & _9078_ /*83680*/;
assign _8920_ = _9071_ ^ _9078_ /*83681*/;
assign _9076_ = _9077_ | _9079_ /*83678*/;
assign _9085_ = ~D[24] /*83677*/;
assign _9082_ = _8472_ & _9085_ /*83673*/;
assign _9083_ = _8472_ ^ _9085_ /*83676*/;
assign _9084_ = _9076_ & _9083_ /*83674*/;
assign _8921_ = _9076_ ^ _9083_ /*83675*/;
assign _9081_ = _9082_ | _9084_ /*83672*/;
assign _9090_ = ~D[25] /*83671*/;
assign _9087_ = _8473_ & _9090_ /*83667*/;
assign _9088_ = _8473_ ^ _9090_ /*83670*/;
assign _9089_ = _9081_ & _9088_ /*83668*/;
assign _8922_ = _9081_ ^ _9088_ /*83669*/;
assign _9086_ = _9087_ | _9089_ /*83666*/;
assign _9095_ = ~D[26] /*83665*/;
assign _9092_ = _8474_ & _9095_ /*83661*/;
assign _9093_ = _8474_ ^ _9095_ /*83664*/;
assign _9094_ = _9086_ & _9093_ /*83662*/;
assign _8923_ = _9086_ ^ _9093_ /*83663*/;
assign _9091_ = _9092_ | _9094_ /*83660*/;
assign _9100_ = ~D[27] /*83659*/;
assign _9097_ = _8475_ & _9100_ /*83655*/;
assign _9098_ = _8475_ ^ _9100_ /*83658*/;
assign _9099_ = _9091_ & _9098_ /*83656*/;
assign _8924_ = _9091_ ^ _9098_ /*83657*/;
assign _9096_ = _9097_ | _9099_ /*83654*/;
assign _9105_ = ~D[28] /*83653*/;
assign _9102_ = _8476_ & _9105_ /*83649*/;
assign _9103_ = _8476_ ^ _9105_ /*83652*/;
assign _9104_ = _9096_ & _9103_ /*83650*/;
assign _8925_ = _9096_ ^ _9103_ /*83651*/;
assign _9101_ = _9102_ | _9104_ /*83648*/;
assign _9110_ = ~D[29] /*83647*/;
assign _9107_ = _8477_ & _9110_ /*83643*/;
assign _9108_ = _8477_ ^ _9110_ /*83646*/;
assign _9109_ = _9101_ & _9108_ /*83644*/;
assign _8926_ = _9101_ ^ _9108_ /*83645*/;
assign _9106_ = _9107_ | _9109_ /*83642*/;
assign _9115_ = ~D[30] /*83641*/;
assign _9112_ = _8478_ & _9115_ /*83637*/;
assign _9113_ = _8478_ ^ _9115_ /*83640*/;
assign _9114_ = _9106_ & _9113_ /*83638*/;
assign _8927_ = _9106_ ^ _9113_ /*83639*/;
assign _9111_ = _9112_ | _9114_ /*83636*/;
assign _9120_ = ~D[31] /*83635*/;
assign _9117_ = _8479_ & _9120_ /*83631*/;
assign _9118_ = _8479_ ^ _9120_ /*83634*/;
assign _9119_ = _9111_ & _9118_ /*83632*/;
assign _8928_ = _9111_ ^ _9118_ /*83633*/;
assign _9116_ = _9117_ | _9119_ /*83630*/;
assign _9125_ = ~D[32] /*83629*/;
assign _9122_ = _8480_ & _9125_ /*83625*/;
assign _9123_ = _8480_ ^ _9125_ /*83628*/;
assign _9124_ = _9116_ & _9123_ /*83626*/;
assign _8929_ = _9116_ ^ _9123_ /*83627*/;
assign _9121_ = _9122_ | _9124_ /*83624*/;
assign _9130_ = ~D[33] /*83623*/;
assign _9127_ = _8481_ & _9130_ /*83619*/;
assign _9128_ = _8481_ ^ _9130_ /*83622*/;
assign _9129_ = _9121_ & _9128_ /*83620*/;
assign _8930_ = _9121_ ^ _9128_ /*83621*/;
assign _9126_ = _9127_ | _9129_ /*83618*/;
assign _9135_ = ~D[34] /*83617*/;
assign _9132_ = _8482_ & _9135_ /*83613*/;
assign _9133_ = _8482_ ^ _9135_ /*83616*/;
assign _9134_ = _9126_ & _9133_ /*83614*/;
assign _8931_ = _9126_ ^ _9133_ /*83615*/;
assign _9131_ = _9132_ | _9134_ /*83612*/;
assign _9140_ = ~D[35] /*83611*/;
assign _9137_ = _8483_ & _9140_ /*83607*/;
assign _9138_ = _8483_ ^ _9140_ /*83610*/;
assign _9139_ = _9131_ & _9138_ /*83608*/;
assign _8932_ = _9131_ ^ _9138_ /*83609*/;
assign _9136_ = _9137_ | _9139_ /*83606*/;
assign _9145_ = ~D[36] /*83605*/;
assign _9142_ = _8484_ & _9145_ /*83601*/;
assign _9143_ = _8484_ ^ _9145_ /*83604*/;
assign _9144_ = _9136_ & _9143_ /*83602*/;
assign _8933_ = _9136_ ^ _9143_ /*83603*/;
assign _9141_ = _9142_ | _9144_ /*83600*/;
assign _9150_ = ~D[37] /*83599*/;
assign _9147_ = _8485_ & _9150_ /*83595*/;
assign _9148_ = _8485_ ^ _9150_ /*83598*/;
assign _9149_ = _9141_ & _9148_ /*83596*/;
assign _8934_ = _9141_ ^ _9148_ /*83597*/;
assign _9146_ = _9147_ | _9149_ /*83594*/;
assign _9155_ = ~D[38] /*83593*/;
assign _9152_ = _8486_ & _9155_ /*83589*/;
assign _9153_ = _8486_ ^ _9155_ /*83592*/;
assign _9154_ = _9146_ & _9153_ /*83590*/;
assign _8935_ = _9146_ ^ _9153_ /*83591*/;
assign _9151_ = _9152_ | _9154_ /*83588*/;
assign _9160_ = ~D[39] /*83587*/;
assign _9157_ = _8487_ & _9160_ /*83583*/;
assign _9158_ = _8487_ ^ _9160_ /*83586*/;
assign _9159_ = _9151_ & _9158_ /*83584*/;
assign _8936_ = _9151_ ^ _9158_ /*83585*/;
assign _9156_ = _9157_ | _9159_ /*83582*/;
assign _9165_ = ~D[40] /*83581*/;
assign _9162_ = _8488_ & _9165_ /*83577*/;
assign _9163_ = _8488_ ^ _9165_ /*83580*/;
assign _9164_ = _9156_ & _9163_ /*83578*/;
assign _8937_ = _9156_ ^ _9163_ /*83579*/;
assign _9161_ = _9162_ | _9164_ /*83576*/;
assign _9170_ = ~D[41] /*83575*/;
assign _9167_ = _8489_ & _9170_ /*83571*/;
assign _9168_ = _8489_ ^ _9170_ /*83574*/;
assign _9169_ = _9161_ & _9168_ /*83572*/;
assign _8938_ = _9161_ ^ _9168_ /*83573*/;
assign _9166_ = _9167_ | _9169_ /*83570*/;
assign _9175_ = ~D[42] /*83569*/;
assign _9172_ = _8490_ & _9175_ /*83565*/;
assign _9173_ = _8490_ ^ _9175_ /*83568*/;
assign _9174_ = _9166_ & _9173_ /*83566*/;
assign _8939_ = _9166_ ^ _9173_ /*83567*/;
assign _9171_ = _9172_ | _9174_ /*83564*/;
assign _9180_ = ~D[43] /*83563*/;
assign _9177_ = _8491_ & _9180_ /*83559*/;
assign _9178_ = _8491_ ^ _9180_ /*83562*/;
assign _9179_ = _9171_ & _9178_ /*83560*/;
assign _8940_ = _9171_ ^ _9178_ /*83561*/;
assign _9176_ = _9177_ | _9179_ /*83558*/;
assign _9185_ = ~D[44] /*83557*/;
assign _9182_ = _8492_ & _9185_ /*83553*/;
assign _9183_ = _8492_ ^ _9185_ /*83556*/;
assign _9184_ = _9176_ & _9183_ /*83554*/;
assign _8941_ = _9176_ ^ _9183_ /*83555*/;
assign _9181_ = _9182_ | _9184_ /*83552*/;
assign _9190_ = ~D[45] /*83551*/;
assign _9187_ = _8493_ & _9190_ /*83547*/;
assign _9188_ = _8493_ ^ _9190_ /*83550*/;
assign _9189_ = _9181_ & _9188_ /*83548*/;
assign _8942_ = _9181_ ^ _9188_ /*83549*/;
assign _9186_ = _9187_ | _9189_ /*83546*/;
assign _9195_ = ~D[46] /*83545*/;
assign _9192_ = _8494_ & _9195_ /*83541*/;
assign _9193_ = _8494_ ^ _9195_ /*83544*/;
assign _9194_ = _9186_ & _9193_ /*83542*/;
assign _8943_ = _9186_ ^ _9193_ /*83543*/;
assign _9191_ = _9192_ | _9194_ /*83540*/;
assign _9200_ = ~D[47] /*83539*/;
assign _9197_ = _8495_ & _9200_ /*83535*/;
assign _9198_ = _8495_ ^ _9200_ /*83538*/;
assign _9199_ = _9191_ & _9198_ /*83536*/;
assign _8944_ = _9191_ ^ _9198_ /*83537*/;
assign _9196_ = _9197_ | _9199_ /*83534*/;
assign _9205_ = ~D[48] /*83533*/;
assign _9202_ = _8496_ & _9205_ /*83529*/;
assign _9203_ = _8496_ ^ _9205_ /*83532*/;
assign _9204_ = _9196_ & _9203_ /*83530*/;
assign _8945_ = _9196_ ^ _9203_ /*83531*/;
assign _9201_ = _9202_ | _9204_ /*83528*/;
assign _9210_ = ~D[49] /*83527*/;
assign _9207_ = _8497_ & _9210_ /*83523*/;
assign _9208_ = _8497_ ^ _9210_ /*83526*/;
assign _9209_ = _9201_ & _9208_ /*83524*/;
assign _8946_ = _9201_ ^ _9208_ /*83525*/;
assign _9206_ = _9207_ | _9209_ /*83522*/;
assign _9215_ = ~D[50] /*83521*/;
assign _9212_ = _8498_ & _9215_ /*83517*/;
assign _9213_ = _8498_ ^ _9215_ /*83520*/;
assign _9214_ = _9206_ & _9213_ /*83518*/;
assign _8947_ = _9206_ ^ _9213_ /*83519*/;
assign _9211_ = _9212_ | _9214_ /*83516*/;
assign _9220_ = ~D[51] /*83515*/;
assign _9217_ = _8499_ & _9220_ /*83511*/;
assign _9218_ = _8499_ ^ _9220_ /*83514*/;
assign _9219_ = _9211_ & _9218_ /*83512*/;
assign _8948_ = _9211_ ^ _9218_ /*83513*/;
assign _9216_ = _9217_ | _9219_ /*83510*/;
assign _9225_ = ~D[52] /*83509*/;
assign _9222_ = _8500_ & _9225_ /*83505*/;
assign _9223_ = _8500_ ^ _9225_ /*83508*/;
assign _9224_ = _9216_ & _9223_ /*83506*/;
assign _8949_ = _9216_ ^ _9223_ /*83507*/;
assign _9221_ = _9222_ | _9224_ /*83504*/;
assign _9230_ = ~D[53] /*83503*/;
assign _9227_ = _8501_ & _9230_ /*83499*/;
assign _9228_ = _8501_ ^ _9230_ /*83502*/;
assign _9229_ = _9221_ & _9228_ /*83500*/;
assign _8950_ = _9221_ ^ _9228_ /*83501*/;
assign _9226_ = _9227_ | _9229_ /*83498*/;
assign _9235_ = ~D[54] /*83497*/;
assign _9232_ = _8502_ & _9235_ /*83493*/;
assign _9233_ = _8502_ ^ _9235_ /*83496*/;
assign _9234_ = _9226_ & _9233_ /*83494*/;
assign _8951_ = _9226_ ^ _9233_ /*83495*/;
assign _9231_ = _9232_ | _9234_ /*83492*/;
assign _9240_ = ~D[55] /*83491*/;
assign _9237_ = _8503_ & _9240_ /*83487*/;
assign _9238_ = _8503_ ^ _9240_ /*83490*/;
assign _9239_ = _9231_ & _9238_ /*83488*/;
assign _8952_ = _9231_ ^ _9238_ /*83489*/;
assign _9236_ = _9237_ | _9239_ /*83486*/;
assign _9245_ = ~D[56] /*83485*/;
assign _9242_ = _8504_ & _9245_ /*83481*/;
assign _9243_ = _8504_ ^ _9245_ /*83484*/;
assign _9244_ = _9236_ & _9243_ /*83482*/;
assign _8953_ = _9236_ ^ _9243_ /*83483*/;
assign _9241_ = _9242_ | _9244_ /*83480*/;
assign _9250_ = ~D[57] /*83479*/;
assign _9247_ = _8505_ & _9250_ /*83475*/;
assign _9248_ = _8505_ ^ _9250_ /*83478*/;
assign _9249_ = _9241_ & _9248_ /*83476*/;
assign _8954_ = _9241_ ^ _9248_ /*83477*/;
assign _9246_ = _9247_ | _9249_ /*83474*/;
assign _9255_ = ~D[58] /*83473*/;
assign _9252_ = _8506_ & _9255_ /*83469*/;
assign _9253_ = _8506_ ^ _9255_ /*83472*/;
assign _9254_ = _9246_ & _9253_ /*83470*/;
assign _8955_ = _9246_ ^ _9253_ /*83471*/;
assign _9251_ = _9252_ | _9254_ /*83468*/;
assign _9260_ = ~D[59] /*83467*/;
assign _9257_ = _8507_ & _9260_ /*83463*/;
assign _9258_ = _8507_ ^ _9260_ /*83466*/;
assign _9259_ = _9251_ & _9258_ /*83464*/;
assign _8956_ = _9251_ ^ _9258_ /*83465*/;
assign _9256_ = _9257_ | _9259_ /*83462*/;
assign _9265_ = ~D[60] /*83461*/;
assign _9262_ = _8508_ & _9265_ /*83457*/;
assign _9263_ = _8508_ ^ _9265_ /*83460*/;
assign _9264_ = _9256_ & _9263_ /*83458*/;
assign _8957_ = _9256_ ^ _9263_ /*83459*/;
assign _9261_ = _9262_ | _9264_ /*83456*/;
assign _9270_ = ~D[61] /*83455*/;
assign _9267_ = _8509_ & _9270_ /*83451*/;
assign _9268_ = _8509_ ^ _9270_ /*83454*/;
assign _9269_ = _9261_ & _9268_ /*83452*/;
assign _8958_ = _9261_ ^ _9268_ /*83453*/;
assign _9266_ = _9267_ | _9269_ /*83450*/;
assign _9275_ = ~D[62] /*83449*/;
assign _9272_ = _8510_ & _9275_ /*83445*/;
assign _9273_ = _8510_ ^ _9275_ /*83448*/;
assign _9274_ = _9266_ & _9273_ /*83446*/;
assign _8959_ = _9266_ ^ _9273_ /*83447*/;
assign _9271_ = _9272_ | _9274_ /*83444*/;
assign _9276_ = _8511_ & oneWire /*83439*/;
assign _9277_ = _8511_ ^ oneWire /*83442*/;
assign _9278_ = _9271_ & _9277_ /*83440*/;
assign _8960_ = _9271_ ^ _9277_ /*83441*/;
assign Q[53] = _9276_ | _9278_ /*83438*/;
assign _9411_ = ~Q[53] /*83053*/;
assign _9410_ = _9411_ & D[0] /*83052*/;
assign _9413_ = _8897_ & _9410_ /*83047*/;
assign _9414_ = _8897_ ^ _9410_ /*83050*/;
assign _9415_ = zeroWire & _9414_ /*83048*/;
assign _9345_ = zeroWire ^ _9414_ /*83049*/;
assign _9412_ = _9413_ | _9415_ /*83046*/;
assign _9417_ = ~Q[53] /*83045*/;
assign _9416_ = _9417_ & D[1] /*83044*/;
assign _9419_ = _8898_ & _9416_ /*83039*/;
assign _9420_ = _8898_ ^ _9416_ /*83042*/;
assign _9421_ = _9412_ & _9420_ /*83040*/;
assign _9346_ = _9412_ ^ _9420_ /*83041*/;
assign _9418_ = _9419_ | _9421_ /*83038*/;
assign _9423_ = ~Q[53] /*83037*/;
assign _9422_ = _9423_ & D[2] /*83036*/;
assign _9425_ = _8899_ & _9422_ /*83031*/;
assign _9426_ = _8899_ ^ _9422_ /*83034*/;
assign _9427_ = _9418_ & _9426_ /*83032*/;
assign _9347_ = _9418_ ^ _9426_ /*83033*/;
assign _9424_ = _9425_ | _9427_ /*83030*/;
assign _9429_ = ~Q[53] /*83029*/;
assign _9428_ = _9429_ & D[3] /*83028*/;
assign _9431_ = _8900_ & _9428_ /*83023*/;
assign _9432_ = _8900_ ^ _9428_ /*83026*/;
assign _9433_ = _9424_ & _9432_ /*83024*/;
assign _9348_ = _9424_ ^ _9432_ /*83025*/;
assign _9430_ = _9431_ | _9433_ /*83022*/;
assign _9435_ = ~Q[53] /*83021*/;
assign _9434_ = _9435_ & D[4] /*83020*/;
assign _9437_ = _8901_ & _9434_ /*83015*/;
assign _9438_ = _8901_ ^ _9434_ /*83018*/;
assign _9439_ = _9430_ & _9438_ /*83016*/;
assign _9349_ = _9430_ ^ _9438_ /*83017*/;
assign _9436_ = _9437_ | _9439_ /*83014*/;
assign _9441_ = ~Q[53] /*83013*/;
assign _9440_ = _9441_ & D[5] /*83012*/;
assign _9443_ = _8902_ & _9440_ /*83007*/;
assign _9444_ = _8902_ ^ _9440_ /*83010*/;
assign _9445_ = _9436_ & _9444_ /*83008*/;
assign _9350_ = _9436_ ^ _9444_ /*83009*/;
assign _9442_ = _9443_ | _9445_ /*83006*/;
assign _9447_ = ~Q[53] /*83005*/;
assign _9446_ = _9447_ & D[6] /*83004*/;
assign _9449_ = _8903_ & _9446_ /*82999*/;
assign _9450_ = _8903_ ^ _9446_ /*83002*/;
assign _9451_ = _9442_ & _9450_ /*83000*/;
assign _9351_ = _9442_ ^ _9450_ /*83001*/;
assign _9448_ = _9449_ | _9451_ /*82998*/;
assign _9453_ = ~Q[53] /*82997*/;
assign _9452_ = _9453_ & D[7] /*82996*/;
assign _9455_ = _8904_ & _9452_ /*82991*/;
assign _9456_ = _8904_ ^ _9452_ /*82994*/;
assign _9457_ = _9448_ & _9456_ /*82992*/;
assign _9352_ = _9448_ ^ _9456_ /*82993*/;
assign _9454_ = _9455_ | _9457_ /*82990*/;
assign _9459_ = ~Q[53] /*82989*/;
assign _9458_ = _9459_ & D[8] /*82988*/;
assign _9461_ = _8905_ & _9458_ /*82983*/;
assign _9462_ = _8905_ ^ _9458_ /*82986*/;
assign _9463_ = _9454_ & _9462_ /*82984*/;
assign _9353_ = _9454_ ^ _9462_ /*82985*/;
assign _9460_ = _9461_ | _9463_ /*82982*/;
assign _9465_ = ~Q[53] /*82981*/;
assign _9464_ = _9465_ & D[9] /*82980*/;
assign _9467_ = _8906_ & _9464_ /*82975*/;
assign _9468_ = _8906_ ^ _9464_ /*82978*/;
assign _9469_ = _9460_ & _9468_ /*82976*/;
assign _9354_ = _9460_ ^ _9468_ /*82977*/;
assign _9466_ = _9467_ | _9469_ /*82974*/;
assign _9471_ = ~Q[53] /*82973*/;
assign _9470_ = _9471_ & D[10] /*82972*/;
assign _9473_ = _8907_ & _9470_ /*82967*/;
assign _9474_ = _8907_ ^ _9470_ /*82970*/;
assign _9475_ = _9466_ & _9474_ /*82968*/;
assign _9355_ = _9466_ ^ _9474_ /*82969*/;
assign _9472_ = _9473_ | _9475_ /*82966*/;
assign _9477_ = ~Q[53] /*82965*/;
assign _9476_ = _9477_ & D[11] /*82964*/;
assign _9479_ = _8908_ & _9476_ /*82959*/;
assign _9480_ = _8908_ ^ _9476_ /*82962*/;
assign _9481_ = _9472_ & _9480_ /*82960*/;
assign _9356_ = _9472_ ^ _9480_ /*82961*/;
assign _9478_ = _9479_ | _9481_ /*82958*/;
assign _9483_ = ~Q[53] /*82957*/;
assign _9482_ = _9483_ & D[12] /*82956*/;
assign _9485_ = _8909_ & _9482_ /*82951*/;
assign _9486_ = _8909_ ^ _9482_ /*82954*/;
assign _9487_ = _9478_ & _9486_ /*82952*/;
assign _9357_ = _9478_ ^ _9486_ /*82953*/;
assign _9484_ = _9485_ | _9487_ /*82950*/;
assign _9489_ = ~Q[53] /*82949*/;
assign _9488_ = _9489_ & D[13] /*82948*/;
assign _9491_ = _8910_ & _9488_ /*82943*/;
assign _9492_ = _8910_ ^ _9488_ /*82946*/;
assign _9493_ = _9484_ & _9492_ /*82944*/;
assign _9358_ = _9484_ ^ _9492_ /*82945*/;
assign _9490_ = _9491_ | _9493_ /*82942*/;
assign _9495_ = ~Q[53] /*82941*/;
assign _9494_ = _9495_ & D[14] /*82940*/;
assign _9497_ = _8911_ & _9494_ /*82935*/;
assign _9498_ = _8911_ ^ _9494_ /*82938*/;
assign _9499_ = _9490_ & _9498_ /*82936*/;
assign _9359_ = _9490_ ^ _9498_ /*82937*/;
assign _9496_ = _9497_ | _9499_ /*82934*/;
assign _9501_ = ~Q[53] /*82933*/;
assign _9500_ = _9501_ & D[15] /*82932*/;
assign _9503_ = _8912_ & _9500_ /*82927*/;
assign _9504_ = _8912_ ^ _9500_ /*82930*/;
assign _9505_ = _9496_ & _9504_ /*82928*/;
assign _9360_ = _9496_ ^ _9504_ /*82929*/;
assign _9502_ = _9503_ | _9505_ /*82926*/;
assign _9507_ = ~Q[53] /*82925*/;
assign _9506_ = _9507_ & D[16] /*82924*/;
assign _9509_ = _8913_ & _9506_ /*82919*/;
assign _9510_ = _8913_ ^ _9506_ /*82922*/;
assign _9511_ = _9502_ & _9510_ /*82920*/;
assign _9361_ = _9502_ ^ _9510_ /*82921*/;
assign _9508_ = _9509_ | _9511_ /*82918*/;
assign _9513_ = ~Q[53] /*82917*/;
assign _9512_ = _9513_ & D[17] /*82916*/;
assign _9515_ = _8914_ & _9512_ /*82911*/;
assign _9516_ = _8914_ ^ _9512_ /*82914*/;
assign _9517_ = _9508_ & _9516_ /*82912*/;
assign _9362_ = _9508_ ^ _9516_ /*82913*/;
assign _9514_ = _9515_ | _9517_ /*82910*/;
assign _9519_ = ~Q[53] /*82909*/;
assign _9518_ = _9519_ & D[18] /*82908*/;
assign _9521_ = _8915_ & _9518_ /*82903*/;
assign _9522_ = _8915_ ^ _9518_ /*82906*/;
assign _9523_ = _9514_ & _9522_ /*82904*/;
assign _9363_ = _9514_ ^ _9522_ /*82905*/;
assign _9520_ = _9521_ | _9523_ /*82902*/;
assign _9525_ = ~Q[53] /*82901*/;
assign _9524_ = _9525_ & D[19] /*82900*/;
assign _9527_ = _8916_ & _9524_ /*82895*/;
assign _9528_ = _8916_ ^ _9524_ /*82898*/;
assign _9529_ = _9520_ & _9528_ /*82896*/;
assign _9364_ = _9520_ ^ _9528_ /*82897*/;
assign _9526_ = _9527_ | _9529_ /*82894*/;
assign _9531_ = ~Q[53] /*82893*/;
assign _9530_ = _9531_ & D[20] /*82892*/;
assign _9533_ = _8917_ & _9530_ /*82887*/;
assign _9534_ = _8917_ ^ _9530_ /*82890*/;
assign _9535_ = _9526_ & _9534_ /*82888*/;
assign _9365_ = _9526_ ^ _9534_ /*82889*/;
assign _9532_ = _9533_ | _9535_ /*82886*/;
assign _9537_ = ~Q[53] /*82885*/;
assign _9536_ = _9537_ & D[21] /*82884*/;
assign _9539_ = _8918_ & _9536_ /*82879*/;
assign _9540_ = _8918_ ^ _9536_ /*82882*/;
assign _9541_ = _9532_ & _9540_ /*82880*/;
assign _9366_ = _9532_ ^ _9540_ /*82881*/;
assign _9538_ = _9539_ | _9541_ /*82878*/;
assign _9543_ = ~Q[53] /*82877*/;
assign _9542_ = _9543_ & D[22] /*82876*/;
assign _9545_ = _8919_ & _9542_ /*82871*/;
assign _9546_ = _8919_ ^ _9542_ /*82874*/;
assign _9547_ = _9538_ & _9546_ /*82872*/;
assign _9367_ = _9538_ ^ _9546_ /*82873*/;
assign _9544_ = _9545_ | _9547_ /*82870*/;
assign _9549_ = ~Q[53] /*82869*/;
assign _9548_ = _9549_ & D[23] /*82868*/;
assign _9551_ = _8920_ & _9548_ /*82863*/;
assign _9552_ = _8920_ ^ _9548_ /*82866*/;
assign _9553_ = _9544_ & _9552_ /*82864*/;
assign _9368_ = _9544_ ^ _9552_ /*82865*/;
assign _9550_ = _9551_ | _9553_ /*82862*/;
assign _9555_ = ~Q[53] /*82861*/;
assign _9554_ = _9555_ & D[24] /*82860*/;
assign _9557_ = _8921_ & _9554_ /*82855*/;
assign _9558_ = _8921_ ^ _9554_ /*82858*/;
assign _9559_ = _9550_ & _9558_ /*82856*/;
assign _9369_ = _9550_ ^ _9558_ /*82857*/;
assign _9556_ = _9557_ | _9559_ /*82854*/;
assign _9561_ = ~Q[53] /*82853*/;
assign _9560_ = _9561_ & D[25] /*82852*/;
assign _9563_ = _8922_ & _9560_ /*82847*/;
assign _9564_ = _8922_ ^ _9560_ /*82850*/;
assign _9565_ = _9556_ & _9564_ /*82848*/;
assign _9370_ = _9556_ ^ _9564_ /*82849*/;
assign _9562_ = _9563_ | _9565_ /*82846*/;
assign _9567_ = ~Q[53] /*82845*/;
assign _9566_ = _9567_ & D[26] /*82844*/;
assign _9569_ = _8923_ & _9566_ /*82839*/;
assign _9570_ = _8923_ ^ _9566_ /*82842*/;
assign _9571_ = _9562_ & _9570_ /*82840*/;
assign _9371_ = _9562_ ^ _9570_ /*82841*/;
assign _9568_ = _9569_ | _9571_ /*82838*/;
assign _9573_ = ~Q[53] /*82837*/;
assign _9572_ = _9573_ & D[27] /*82836*/;
assign _9575_ = _8924_ & _9572_ /*82831*/;
assign _9576_ = _8924_ ^ _9572_ /*82834*/;
assign _9577_ = _9568_ & _9576_ /*82832*/;
assign _9372_ = _9568_ ^ _9576_ /*82833*/;
assign _9574_ = _9575_ | _9577_ /*82830*/;
assign _9579_ = ~Q[53] /*82829*/;
assign _9578_ = _9579_ & D[28] /*82828*/;
assign _9581_ = _8925_ & _9578_ /*82823*/;
assign _9582_ = _8925_ ^ _9578_ /*82826*/;
assign _9583_ = _9574_ & _9582_ /*82824*/;
assign _9373_ = _9574_ ^ _9582_ /*82825*/;
assign _9580_ = _9581_ | _9583_ /*82822*/;
assign _9585_ = ~Q[53] /*82821*/;
assign _9584_ = _9585_ & D[29] /*82820*/;
assign _9587_ = _8926_ & _9584_ /*82815*/;
assign _9588_ = _8926_ ^ _9584_ /*82818*/;
assign _9589_ = _9580_ & _9588_ /*82816*/;
assign _9374_ = _9580_ ^ _9588_ /*82817*/;
assign _9586_ = _9587_ | _9589_ /*82814*/;
assign _9591_ = ~Q[53] /*82813*/;
assign _9590_ = _9591_ & D[30] /*82812*/;
assign _9593_ = _8927_ & _9590_ /*82807*/;
assign _9594_ = _8927_ ^ _9590_ /*82810*/;
assign _9595_ = _9586_ & _9594_ /*82808*/;
assign _9375_ = _9586_ ^ _9594_ /*82809*/;
assign _9592_ = _9593_ | _9595_ /*82806*/;
assign _9597_ = ~Q[53] /*82805*/;
assign _9596_ = _9597_ & D[31] /*82804*/;
assign _9599_ = _8928_ & _9596_ /*82799*/;
assign _9600_ = _8928_ ^ _9596_ /*82802*/;
assign _9601_ = _9592_ & _9600_ /*82800*/;
assign _9376_ = _9592_ ^ _9600_ /*82801*/;
assign _9598_ = _9599_ | _9601_ /*82798*/;
assign _9603_ = ~Q[53] /*82797*/;
assign _9602_ = _9603_ & D[32] /*82796*/;
assign _9605_ = _8929_ & _9602_ /*82791*/;
assign _9606_ = _8929_ ^ _9602_ /*82794*/;
assign _9607_ = _9598_ & _9606_ /*82792*/;
assign _9377_ = _9598_ ^ _9606_ /*82793*/;
assign _9604_ = _9605_ | _9607_ /*82790*/;
assign _9609_ = ~Q[53] /*82789*/;
assign _9608_ = _9609_ & D[33] /*82788*/;
assign _9611_ = _8930_ & _9608_ /*82783*/;
assign _9612_ = _8930_ ^ _9608_ /*82786*/;
assign _9613_ = _9604_ & _9612_ /*82784*/;
assign _9378_ = _9604_ ^ _9612_ /*82785*/;
assign _9610_ = _9611_ | _9613_ /*82782*/;
assign _9615_ = ~Q[53] /*82781*/;
assign _9614_ = _9615_ & D[34] /*82780*/;
assign _9617_ = _8931_ & _9614_ /*82775*/;
assign _9618_ = _8931_ ^ _9614_ /*82778*/;
assign _9619_ = _9610_ & _9618_ /*82776*/;
assign _9379_ = _9610_ ^ _9618_ /*82777*/;
assign _9616_ = _9617_ | _9619_ /*82774*/;
assign _9621_ = ~Q[53] /*82773*/;
assign _9620_ = _9621_ & D[35] /*82772*/;
assign _9623_ = _8932_ & _9620_ /*82767*/;
assign _9624_ = _8932_ ^ _9620_ /*82770*/;
assign _9625_ = _9616_ & _9624_ /*82768*/;
assign _9380_ = _9616_ ^ _9624_ /*82769*/;
assign _9622_ = _9623_ | _9625_ /*82766*/;
assign _9627_ = ~Q[53] /*82765*/;
assign _9626_ = _9627_ & D[36] /*82764*/;
assign _9629_ = _8933_ & _9626_ /*82759*/;
assign _9630_ = _8933_ ^ _9626_ /*82762*/;
assign _9631_ = _9622_ & _9630_ /*82760*/;
assign _9381_ = _9622_ ^ _9630_ /*82761*/;
assign _9628_ = _9629_ | _9631_ /*82758*/;
assign _9633_ = ~Q[53] /*82757*/;
assign _9632_ = _9633_ & D[37] /*82756*/;
assign _9635_ = _8934_ & _9632_ /*82751*/;
assign _9636_ = _8934_ ^ _9632_ /*82754*/;
assign _9637_ = _9628_ & _9636_ /*82752*/;
assign _9382_ = _9628_ ^ _9636_ /*82753*/;
assign _9634_ = _9635_ | _9637_ /*82750*/;
assign _9639_ = ~Q[53] /*82749*/;
assign _9638_ = _9639_ & D[38] /*82748*/;
assign _9641_ = _8935_ & _9638_ /*82743*/;
assign _9642_ = _8935_ ^ _9638_ /*82746*/;
assign _9643_ = _9634_ & _9642_ /*82744*/;
assign _9383_ = _9634_ ^ _9642_ /*82745*/;
assign _9640_ = _9641_ | _9643_ /*82742*/;
assign _9645_ = ~Q[53] /*82741*/;
assign _9644_ = _9645_ & D[39] /*82740*/;
assign _9647_ = _8936_ & _9644_ /*82735*/;
assign _9648_ = _8936_ ^ _9644_ /*82738*/;
assign _9649_ = _9640_ & _9648_ /*82736*/;
assign _9384_ = _9640_ ^ _9648_ /*82737*/;
assign _9646_ = _9647_ | _9649_ /*82734*/;
assign _9651_ = ~Q[53] /*82733*/;
assign _9650_ = _9651_ & D[40] /*82732*/;
assign _9653_ = _8937_ & _9650_ /*82727*/;
assign _9654_ = _8937_ ^ _9650_ /*82730*/;
assign _9655_ = _9646_ & _9654_ /*82728*/;
assign _9385_ = _9646_ ^ _9654_ /*82729*/;
assign _9652_ = _9653_ | _9655_ /*82726*/;
assign _9657_ = ~Q[53] /*82725*/;
assign _9656_ = _9657_ & D[41] /*82724*/;
assign _9659_ = _8938_ & _9656_ /*82719*/;
assign _9660_ = _8938_ ^ _9656_ /*82722*/;
assign _9661_ = _9652_ & _9660_ /*82720*/;
assign _9386_ = _9652_ ^ _9660_ /*82721*/;
assign _9658_ = _9659_ | _9661_ /*82718*/;
assign _9663_ = ~Q[53] /*82717*/;
assign _9662_ = _9663_ & D[42] /*82716*/;
assign _9665_ = _8939_ & _9662_ /*82711*/;
assign _9666_ = _8939_ ^ _9662_ /*82714*/;
assign _9667_ = _9658_ & _9666_ /*82712*/;
assign _9387_ = _9658_ ^ _9666_ /*82713*/;
assign _9664_ = _9665_ | _9667_ /*82710*/;
assign _9669_ = ~Q[53] /*82709*/;
assign _9668_ = _9669_ & D[43] /*82708*/;
assign _9671_ = _8940_ & _9668_ /*82703*/;
assign _9672_ = _8940_ ^ _9668_ /*82706*/;
assign _9673_ = _9664_ & _9672_ /*82704*/;
assign _9388_ = _9664_ ^ _9672_ /*82705*/;
assign _9670_ = _9671_ | _9673_ /*82702*/;
assign _9675_ = ~Q[53] /*82701*/;
assign _9674_ = _9675_ & D[44] /*82700*/;
assign _9677_ = _8941_ & _9674_ /*82695*/;
assign _9678_ = _8941_ ^ _9674_ /*82698*/;
assign _9679_ = _9670_ & _9678_ /*82696*/;
assign _9389_ = _9670_ ^ _9678_ /*82697*/;
assign _9676_ = _9677_ | _9679_ /*82694*/;
assign _9681_ = ~Q[53] /*82693*/;
assign _9680_ = _9681_ & D[45] /*82692*/;
assign _9683_ = _8942_ & _9680_ /*82687*/;
assign _9684_ = _8942_ ^ _9680_ /*82690*/;
assign _9685_ = _9676_ & _9684_ /*82688*/;
assign _9390_ = _9676_ ^ _9684_ /*82689*/;
assign _9682_ = _9683_ | _9685_ /*82686*/;
assign _9687_ = ~Q[53] /*82685*/;
assign _9686_ = _9687_ & D[46] /*82684*/;
assign _9689_ = _8943_ & _9686_ /*82679*/;
assign _9690_ = _8943_ ^ _9686_ /*82682*/;
assign _9691_ = _9682_ & _9690_ /*82680*/;
assign _9391_ = _9682_ ^ _9690_ /*82681*/;
assign _9688_ = _9689_ | _9691_ /*82678*/;
assign _9693_ = ~Q[53] /*82677*/;
assign _9692_ = _9693_ & D[47] /*82676*/;
assign _9695_ = _8944_ & _9692_ /*82671*/;
assign _9696_ = _8944_ ^ _9692_ /*82674*/;
assign _9697_ = _9688_ & _9696_ /*82672*/;
assign _9392_ = _9688_ ^ _9696_ /*82673*/;
assign _9694_ = _9695_ | _9697_ /*82670*/;
assign _9699_ = ~Q[53] /*82669*/;
assign _9698_ = _9699_ & D[48] /*82668*/;
assign _9701_ = _8945_ & _9698_ /*82663*/;
assign _9702_ = _8945_ ^ _9698_ /*82666*/;
assign _9703_ = _9694_ & _9702_ /*82664*/;
assign _9393_ = _9694_ ^ _9702_ /*82665*/;
assign _9700_ = _9701_ | _9703_ /*82662*/;
assign _9705_ = ~Q[53] /*82661*/;
assign _9704_ = _9705_ & D[49] /*82660*/;
assign _9707_ = _8946_ & _9704_ /*82655*/;
assign _9708_ = _8946_ ^ _9704_ /*82658*/;
assign _9709_ = _9700_ & _9708_ /*82656*/;
assign _9394_ = _9700_ ^ _9708_ /*82657*/;
assign _9706_ = _9707_ | _9709_ /*82654*/;
assign _9711_ = ~Q[53] /*82653*/;
assign _9710_ = _9711_ & D[50] /*82652*/;
assign _9713_ = _8947_ & _9710_ /*82647*/;
assign _9714_ = _8947_ ^ _9710_ /*82650*/;
assign _9715_ = _9706_ & _9714_ /*82648*/;
assign _9395_ = _9706_ ^ _9714_ /*82649*/;
assign _9712_ = _9713_ | _9715_ /*82646*/;
assign _9717_ = ~Q[53] /*82645*/;
assign _9716_ = _9717_ & D[51] /*82644*/;
assign _9719_ = _8948_ & _9716_ /*82639*/;
assign _9720_ = _8948_ ^ _9716_ /*82642*/;
assign _9721_ = _9712_ & _9720_ /*82640*/;
assign _9396_ = _9712_ ^ _9720_ /*82641*/;
assign _9718_ = _9719_ | _9721_ /*82638*/;
assign _9723_ = ~Q[53] /*82637*/;
assign _9722_ = _9723_ & D[52] /*82636*/;
assign _9725_ = _8949_ & _9722_ /*82631*/;
assign _9726_ = _8949_ ^ _9722_ /*82634*/;
assign _9727_ = _9718_ & _9726_ /*82632*/;
assign _9397_ = _9718_ ^ _9726_ /*82633*/;
assign _9724_ = _9725_ | _9727_ /*82630*/;
assign _9729_ = ~Q[53] /*82629*/;
assign _9728_ = _9729_ & D[53] /*82628*/;
assign _9731_ = _8950_ & _9728_ /*82623*/;
assign _9732_ = _8950_ ^ _9728_ /*82626*/;
assign _9733_ = _9724_ & _9732_ /*82624*/;
assign _9398_ = _9724_ ^ _9732_ /*82625*/;
assign _9730_ = _9731_ | _9733_ /*82622*/;
assign _9735_ = ~Q[53] /*82621*/;
assign _9734_ = _9735_ & D[54] /*82620*/;
assign _9737_ = _8951_ & _9734_ /*82615*/;
assign _9738_ = _8951_ ^ _9734_ /*82618*/;
assign _9739_ = _9730_ & _9738_ /*82616*/;
assign _9399_ = _9730_ ^ _9738_ /*82617*/;
assign _9736_ = _9737_ | _9739_ /*82614*/;
assign _9741_ = ~Q[53] /*82613*/;
assign _9740_ = _9741_ & D[55] /*82612*/;
assign _9743_ = _8952_ & _9740_ /*82607*/;
assign _9744_ = _8952_ ^ _9740_ /*82610*/;
assign _9745_ = _9736_ & _9744_ /*82608*/;
assign _9400_ = _9736_ ^ _9744_ /*82609*/;
assign _9742_ = _9743_ | _9745_ /*82606*/;
assign _9747_ = ~Q[53] /*82605*/;
assign _9746_ = _9747_ & D[56] /*82604*/;
assign _9749_ = _8953_ & _9746_ /*82599*/;
assign _9750_ = _8953_ ^ _9746_ /*82602*/;
assign _9751_ = _9742_ & _9750_ /*82600*/;
assign _9401_ = _9742_ ^ _9750_ /*82601*/;
assign _9748_ = _9749_ | _9751_ /*82598*/;
assign _9753_ = ~Q[53] /*82597*/;
assign _9752_ = _9753_ & D[57] /*82596*/;
assign _9755_ = _8954_ & _9752_ /*82591*/;
assign _9756_ = _8954_ ^ _9752_ /*82594*/;
assign _9757_ = _9748_ & _9756_ /*82592*/;
assign _9402_ = _9748_ ^ _9756_ /*82593*/;
assign _9754_ = _9755_ | _9757_ /*82590*/;
assign _9759_ = ~Q[53] /*82589*/;
assign _9758_ = _9759_ & D[58] /*82588*/;
assign _9761_ = _8955_ & _9758_ /*82583*/;
assign _9762_ = _8955_ ^ _9758_ /*82586*/;
assign _9763_ = _9754_ & _9762_ /*82584*/;
assign _9403_ = _9754_ ^ _9762_ /*82585*/;
assign _9760_ = _9761_ | _9763_ /*82582*/;
assign _9765_ = ~Q[53] /*82581*/;
assign _9764_ = _9765_ & D[59] /*82580*/;
assign _9767_ = _8956_ & _9764_ /*82575*/;
assign _9768_ = _8956_ ^ _9764_ /*82578*/;
assign _9769_ = _9760_ & _9768_ /*82576*/;
assign _9404_ = _9760_ ^ _9768_ /*82577*/;
assign _9766_ = _9767_ | _9769_ /*82574*/;
assign _9771_ = ~Q[53] /*82573*/;
assign _9770_ = _9771_ & D[60] /*82572*/;
assign _9773_ = _8957_ & _9770_ /*82567*/;
assign _9774_ = _8957_ ^ _9770_ /*82570*/;
assign _9775_ = _9766_ & _9774_ /*82568*/;
assign _9405_ = _9766_ ^ _9774_ /*82569*/;
assign _9772_ = _9773_ | _9775_ /*82566*/;
assign _9777_ = ~Q[53] /*82565*/;
assign _9776_ = _9777_ & D[61] /*82564*/;
assign _9779_ = _8958_ & _9776_ /*82559*/;
assign _9780_ = _8958_ ^ _9776_ /*82562*/;
assign _9781_ = _9772_ & _9780_ /*82560*/;
assign _9406_ = _9772_ ^ _9780_ /*82561*/;
assign _9778_ = _9779_ | _9781_ /*82558*/;
assign _9783_ = ~Q[53] /*82557*/;
assign _9782_ = _9783_ & D[62] /*82556*/;
assign _9785_ = _8959_ & _9782_ /*82551*/;
assign _9786_ = _8959_ ^ _9782_ /*82554*/;
assign _9787_ = _9778_ & _9786_ /*82552*/;
assign _9407_ = _9778_ ^ _9786_ /*82553*/;
assign _9784_ = _9785_ | _9787_ /*82550*/;
assign _9789_ = ~Q[53] /*82549*/;
assign _9788_ = _9789_ & zeroWire /*82548*/;
assign _9790_ = _8960_ ^ _9788_ /*82546*/;
assign _9408_ = _9790_ ^ _9784_ /*82545*/;
assign _9861_ = ~D[0] /*82291*/;
assign _9858_ = R_0[52] & _9861_ /*82287*/;
assign _9859_ = R_0[52] ^ _9861_ /*82290*/;
assign _9860_ = oneWire & _9859_ /*82288*/;
assign _9793_ = oneWire ^ _9859_ /*82289*/;
assign _9857_ = _9858_ | _9860_ /*82286*/;
assign _9866_ = ~D[1] /*82285*/;
assign _9863_ = _9345_ & _9866_ /*82281*/;
assign _9864_ = _9345_ ^ _9866_ /*82284*/;
assign _9865_ = _9857_ & _9864_ /*82282*/;
assign _9794_ = _9857_ ^ _9864_ /*82283*/;
assign _9862_ = _9863_ | _9865_ /*82280*/;
assign _9871_ = ~D[2] /*82279*/;
assign _9868_ = _9346_ & _9871_ /*82275*/;
assign _9869_ = _9346_ ^ _9871_ /*82278*/;
assign _9870_ = _9862_ & _9869_ /*82276*/;
assign _9795_ = _9862_ ^ _9869_ /*82277*/;
assign _9867_ = _9868_ | _9870_ /*82274*/;
assign _9876_ = ~D[3] /*82273*/;
assign _9873_ = _9347_ & _9876_ /*82269*/;
assign _9874_ = _9347_ ^ _9876_ /*82272*/;
assign _9875_ = _9867_ & _9874_ /*82270*/;
assign _9796_ = _9867_ ^ _9874_ /*82271*/;
assign _9872_ = _9873_ | _9875_ /*82268*/;
assign _9881_ = ~D[4] /*82267*/;
assign _9878_ = _9348_ & _9881_ /*82263*/;
assign _9879_ = _9348_ ^ _9881_ /*82266*/;
assign _9880_ = _9872_ & _9879_ /*82264*/;
assign _9797_ = _9872_ ^ _9879_ /*82265*/;
assign _9877_ = _9878_ | _9880_ /*82262*/;
assign _9886_ = ~D[5] /*82261*/;
assign _9883_ = _9349_ & _9886_ /*82257*/;
assign _9884_ = _9349_ ^ _9886_ /*82260*/;
assign _9885_ = _9877_ & _9884_ /*82258*/;
assign _9798_ = _9877_ ^ _9884_ /*82259*/;
assign _9882_ = _9883_ | _9885_ /*82256*/;
assign _9891_ = ~D[6] /*82255*/;
assign _9888_ = _9350_ & _9891_ /*82251*/;
assign _9889_ = _9350_ ^ _9891_ /*82254*/;
assign _9890_ = _9882_ & _9889_ /*82252*/;
assign _9799_ = _9882_ ^ _9889_ /*82253*/;
assign _9887_ = _9888_ | _9890_ /*82250*/;
assign _9896_ = ~D[7] /*82249*/;
assign _9893_ = _9351_ & _9896_ /*82245*/;
assign _9894_ = _9351_ ^ _9896_ /*82248*/;
assign _9895_ = _9887_ & _9894_ /*82246*/;
assign _9800_ = _9887_ ^ _9894_ /*82247*/;
assign _9892_ = _9893_ | _9895_ /*82244*/;
assign _9901_ = ~D[8] /*82243*/;
assign _9898_ = _9352_ & _9901_ /*82239*/;
assign _9899_ = _9352_ ^ _9901_ /*82242*/;
assign _9900_ = _9892_ & _9899_ /*82240*/;
assign _9801_ = _9892_ ^ _9899_ /*82241*/;
assign _9897_ = _9898_ | _9900_ /*82238*/;
assign _9906_ = ~D[9] /*82237*/;
assign _9903_ = _9353_ & _9906_ /*82233*/;
assign _9904_ = _9353_ ^ _9906_ /*82236*/;
assign _9905_ = _9897_ & _9904_ /*82234*/;
assign _9802_ = _9897_ ^ _9904_ /*82235*/;
assign _9902_ = _9903_ | _9905_ /*82232*/;
assign _9911_ = ~D[10] /*82231*/;
assign _9908_ = _9354_ & _9911_ /*82227*/;
assign _9909_ = _9354_ ^ _9911_ /*82230*/;
assign _9910_ = _9902_ & _9909_ /*82228*/;
assign _9803_ = _9902_ ^ _9909_ /*82229*/;
assign _9907_ = _9908_ | _9910_ /*82226*/;
assign _9916_ = ~D[11] /*82225*/;
assign _9913_ = _9355_ & _9916_ /*82221*/;
assign _9914_ = _9355_ ^ _9916_ /*82224*/;
assign _9915_ = _9907_ & _9914_ /*82222*/;
assign _9804_ = _9907_ ^ _9914_ /*82223*/;
assign _9912_ = _9913_ | _9915_ /*82220*/;
assign _9921_ = ~D[12] /*82219*/;
assign _9918_ = _9356_ & _9921_ /*82215*/;
assign _9919_ = _9356_ ^ _9921_ /*82218*/;
assign _9920_ = _9912_ & _9919_ /*82216*/;
assign _9805_ = _9912_ ^ _9919_ /*82217*/;
assign _9917_ = _9918_ | _9920_ /*82214*/;
assign _9926_ = ~D[13] /*82213*/;
assign _9923_ = _9357_ & _9926_ /*82209*/;
assign _9924_ = _9357_ ^ _9926_ /*82212*/;
assign _9925_ = _9917_ & _9924_ /*82210*/;
assign _9806_ = _9917_ ^ _9924_ /*82211*/;
assign _9922_ = _9923_ | _9925_ /*82208*/;
assign _9931_ = ~D[14] /*82207*/;
assign _9928_ = _9358_ & _9931_ /*82203*/;
assign _9929_ = _9358_ ^ _9931_ /*82206*/;
assign _9930_ = _9922_ & _9929_ /*82204*/;
assign _9807_ = _9922_ ^ _9929_ /*82205*/;
assign _9927_ = _9928_ | _9930_ /*82202*/;
assign _9936_ = ~D[15] /*82201*/;
assign _9933_ = _9359_ & _9936_ /*82197*/;
assign _9934_ = _9359_ ^ _9936_ /*82200*/;
assign _9935_ = _9927_ & _9934_ /*82198*/;
assign _9808_ = _9927_ ^ _9934_ /*82199*/;
assign _9932_ = _9933_ | _9935_ /*82196*/;
assign _9941_ = ~D[16] /*82195*/;
assign _9938_ = _9360_ & _9941_ /*82191*/;
assign _9939_ = _9360_ ^ _9941_ /*82194*/;
assign _9940_ = _9932_ & _9939_ /*82192*/;
assign _9809_ = _9932_ ^ _9939_ /*82193*/;
assign _9937_ = _9938_ | _9940_ /*82190*/;
assign _9946_ = ~D[17] /*82189*/;
assign _9943_ = _9361_ & _9946_ /*82185*/;
assign _9944_ = _9361_ ^ _9946_ /*82188*/;
assign _9945_ = _9937_ & _9944_ /*82186*/;
assign _9810_ = _9937_ ^ _9944_ /*82187*/;
assign _9942_ = _9943_ | _9945_ /*82184*/;
assign _9951_ = ~D[18] /*82183*/;
assign _9948_ = _9362_ & _9951_ /*82179*/;
assign _9949_ = _9362_ ^ _9951_ /*82182*/;
assign _9950_ = _9942_ & _9949_ /*82180*/;
assign _9811_ = _9942_ ^ _9949_ /*82181*/;
assign _9947_ = _9948_ | _9950_ /*82178*/;
assign _9956_ = ~D[19] /*82177*/;
assign _9953_ = _9363_ & _9956_ /*82173*/;
assign _9954_ = _9363_ ^ _9956_ /*82176*/;
assign _9955_ = _9947_ & _9954_ /*82174*/;
assign _9812_ = _9947_ ^ _9954_ /*82175*/;
assign _9952_ = _9953_ | _9955_ /*82172*/;
assign _9961_ = ~D[20] /*82171*/;
assign _9958_ = _9364_ & _9961_ /*82167*/;
assign _9959_ = _9364_ ^ _9961_ /*82170*/;
assign _9960_ = _9952_ & _9959_ /*82168*/;
assign _9813_ = _9952_ ^ _9959_ /*82169*/;
assign _9957_ = _9958_ | _9960_ /*82166*/;
assign _9966_ = ~D[21] /*82165*/;
assign _9963_ = _9365_ & _9966_ /*82161*/;
assign _9964_ = _9365_ ^ _9966_ /*82164*/;
assign _9965_ = _9957_ & _9964_ /*82162*/;
assign _9814_ = _9957_ ^ _9964_ /*82163*/;
assign _9962_ = _9963_ | _9965_ /*82160*/;
assign _9971_ = ~D[22] /*82159*/;
assign _9968_ = _9366_ & _9971_ /*82155*/;
assign _9969_ = _9366_ ^ _9971_ /*82158*/;
assign _9970_ = _9962_ & _9969_ /*82156*/;
assign _9815_ = _9962_ ^ _9969_ /*82157*/;
assign _9967_ = _9968_ | _9970_ /*82154*/;
assign _9976_ = ~D[23] /*82153*/;
assign _9973_ = _9367_ & _9976_ /*82149*/;
assign _9974_ = _9367_ ^ _9976_ /*82152*/;
assign _9975_ = _9967_ & _9974_ /*82150*/;
assign _9816_ = _9967_ ^ _9974_ /*82151*/;
assign _9972_ = _9973_ | _9975_ /*82148*/;
assign _9981_ = ~D[24] /*82147*/;
assign _9978_ = _9368_ & _9981_ /*82143*/;
assign _9979_ = _9368_ ^ _9981_ /*82146*/;
assign _9980_ = _9972_ & _9979_ /*82144*/;
assign _9817_ = _9972_ ^ _9979_ /*82145*/;
assign _9977_ = _9978_ | _9980_ /*82142*/;
assign _9986_ = ~D[25] /*82141*/;
assign _9983_ = _9369_ & _9986_ /*82137*/;
assign _9984_ = _9369_ ^ _9986_ /*82140*/;
assign _9985_ = _9977_ & _9984_ /*82138*/;
assign _9818_ = _9977_ ^ _9984_ /*82139*/;
assign _9982_ = _9983_ | _9985_ /*82136*/;
assign _9991_ = ~D[26] /*82135*/;
assign _9988_ = _9370_ & _9991_ /*82131*/;
assign _9989_ = _9370_ ^ _9991_ /*82134*/;
assign _9990_ = _9982_ & _9989_ /*82132*/;
assign _9819_ = _9982_ ^ _9989_ /*82133*/;
assign _9987_ = _9988_ | _9990_ /*82130*/;
assign _9996_ = ~D[27] /*82129*/;
assign _9993_ = _9371_ & _9996_ /*82125*/;
assign _9994_ = _9371_ ^ _9996_ /*82128*/;
assign _9995_ = _9987_ & _9994_ /*82126*/;
assign _9820_ = _9987_ ^ _9994_ /*82127*/;
assign _9992_ = _9993_ | _9995_ /*82124*/;
assign _10001_ = ~D[28] /*82123*/;
assign _9998_ = _9372_ & _10001_ /*82119*/;
assign _9999_ = _9372_ ^ _10001_ /*82122*/;
assign _10000_ = _9992_ & _9999_ /*82120*/;
assign _9821_ = _9992_ ^ _9999_ /*82121*/;
assign _9997_ = _9998_ | _10000_ /*82118*/;
assign _10006_ = ~D[29] /*82117*/;
assign _10003_ = _9373_ & _10006_ /*82113*/;
assign _10004_ = _9373_ ^ _10006_ /*82116*/;
assign _10005_ = _9997_ & _10004_ /*82114*/;
assign _9822_ = _9997_ ^ _10004_ /*82115*/;
assign _10002_ = _10003_ | _10005_ /*82112*/;
assign _10011_ = ~D[30] /*82111*/;
assign _10008_ = _9374_ & _10011_ /*82107*/;
assign _10009_ = _9374_ ^ _10011_ /*82110*/;
assign _10010_ = _10002_ & _10009_ /*82108*/;
assign _9823_ = _10002_ ^ _10009_ /*82109*/;
assign _10007_ = _10008_ | _10010_ /*82106*/;
assign _10016_ = ~D[31] /*82105*/;
assign _10013_ = _9375_ & _10016_ /*82101*/;
assign _10014_ = _9375_ ^ _10016_ /*82104*/;
assign _10015_ = _10007_ & _10014_ /*82102*/;
assign _9824_ = _10007_ ^ _10014_ /*82103*/;
assign _10012_ = _10013_ | _10015_ /*82100*/;
assign _10021_ = ~D[32] /*82099*/;
assign _10018_ = _9376_ & _10021_ /*82095*/;
assign _10019_ = _9376_ ^ _10021_ /*82098*/;
assign _10020_ = _10012_ & _10019_ /*82096*/;
assign _9825_ = _10012_ ^ _10019_ /*82097*/;
assign _10017_ = _10018_ | _10020_ /*82094*/;
assign _10026_ = ~D[33] /*82093*/;
assign _10023_ = _9377_ & _10026_ /*82089*/;
assign _10024_ = _9377_ ^ _10026_ /*82092*/;
assign _10025_ = _10017_ & _10024_ /*82090*/;
assign _9826_ = _10017_ ^ _10024_ /*82091*/;
assign _10022_ = _10023_ | _10025_ /*82088*/;
assign _10031_ = ~D[34] /*82087*/;
assign _10028_ = _9378_ & _10031_ /*82083*/;
assign _10029_ = _9378_ ^ _10031_ /*82086*/;
assign _10030_ = _10022_ & _10029_ /*82084*/;
assign _9827_ = _10022_ ^ _10029_ /*82085*/;
assign _10027_ = _10028_ | _10030_ /*82082*/;
assign _10036_ = ~D[35] /*82081*/;
assign _10033_ = _9379_ & _10036_ /*82077*/;
assign _10034_ = _9379_ ^ _10036_ /*82080*/;
assign _10035_ = _10027_ & _10034_ /*82078*/;
assign _9828_ = _10027_ ^ _10034_ /*82079*/;
assign _10032_ = _10033_ | _10035_ /*82076*/;
assign _10041_ = ~D[36] /*82075*/;
assign _10038_ = _9380_ & _10041_ /*82071*/;
assign _10039_ = _9380_ ^ _10041_ /*82074*/;
assign _10040_ = _10032_ & _10039_ /*82072*/;
assign _9829_ = _10032_ ^ _10039_ /*82073*/;
assign _10037_ = _10038_ | _10040_ /*82070*/;
assign _10046_ = ~D[37] /*82069*/;
assign _10043_ = _9381_ & _10046_ /*82065*/;
assign _10044_ = _9381_ ^ _10046_ /*82068*/;
assign _10045_ = _10037_ & _10044_ /*82066*/;
assign _9830_ = _10037_ ^ _10044_ /*82067*/;
assign _10042_ = _10043_ | _10045_ /*82064*/;
assign _10051_ = ~D[38] /*82063*/;
assign _10048_ = _9382_ & _10051_ /*82059*/;
assign _10049_ = _9382_ ^ _10051_ /*82062*/;
assign _10050_ = _10042_ & _10049_ /*82060*/;
assign _9831_ = _10042_ ^ _10049_ /*82061*/;
assign _10047_ = _10048_ | _10050_ /*82058*/;
assign _10056_ = ~D[39] /*82057*/;
assign _10053_ = _9383_ & _10056_ /*82053*/;
assign _10054_ = _9383_ ^ _10056_ /*82056*/;
assign _10055_ = _10047_ & _10054_ /*82054*/;
assign _9832_ = _10047_ ^ _10054_ /*82055*/;
assign _10052_ = _10053_ | _10055_ /*82052*/;
assign _10061_ = ~D[40] /*82051*/;
assign _10058_ = _9384_ & _10061_ /*82047*/;
assign _10059_ = _9384_ ^ _10061_ /*82050*/;
assign _10060_ = _10052_ & _10059_ /*82048*/;
assign _9833_ = _10052_ ^ _10059_ /*82049*/;
assign _10057_ = _10058_ | _10060_ /*82046*/;
assign _10066_ = ~D[41] /*82045*/;
assign _10063_ = _9385_ & _10066_ /*82041*/;
assign _10064_ = _9385_ ^ _10066_ /*82044*/;
assign _10065_ = _10057_ & _10064_ /*82042*/;
assign _9834_ = _10057_ ^ _10064_ /*82043*/;
assign _10062_ = _10063_ | _10065_ /*82040*/;
assign _10071_ = ~D[42] /*82039*/;
assign _10068_ = _9386_ & _10071_ /*82035*/;
assign _10069_ = _9386_ ^ _10071_ /*82038*/;
assign _10070_ = _10062_ & _10069_ /*82036*/;
assign _9835_ = _10062_ ^ _10069_ /*82037*/;
assign _10067_ = _10068_ | _10070_ /*82034*/;
assign _10076_ = ~D[43] /*82033*/;
assign _10073_ = _9387_ & _10076_ /*82029*/;
assign _10074_ = _9387_ ^ _10076_ /*82032*/;
assign _10075_ = _10067_ & _10074_ /*82030*/;
assign _9836_ = _10067_ ^ _10074_ /*82031*/;
assign _10072_ = _10073_ | _10075_ /*82028*/;
assign _10081_ = ~D[44] /*82027*/;
assign _10078_ = _9388_ & _10081_ /*82023*/;
assign _10079_ = _9388_ ^ _10081_ /*82026*/;
assign _10080_ = _10072_ & _10079_ /*82024*/;
assign _9837_ = _10072_ ^ _10079_ /*82025*/;
assign _10077_ = _10078_ | _10080_ /*82022*/;
assign _10086_ = ~D[45] /*82021*/;
assign _10083_ = _9389_ & _10086_ /*82017*/;
assign _10084_ = _9389_ ^ _10086_ /*82020*/;
assign _10085_ = _10077_ & _10084_ /*82018*/;
assign _9838_ = _10077_ ^ _10084_ /*82019*/;
assign _10082_ = _10083_ | _10085_ /*82016*/;
assign _10091_ = ~D[46] /*82015*/;
assign _10088_ = _9390_ & _10091_ /*82011*/;
assign _10089_ = _9390_ ^ _10091_ /*82014*/;
assign _10090_ = _10082_ & _10089_ /*82012*/;
assign _9839_ = _10082_ ^ _10089_ /*82013*/;
assign _10087_ = _10088_ | _10090_ /*82010*/;
assign _10096_ = ~D[47] /*82009*/;
assign _10093_ = _9391_ & _10096_ /*82005*/;
assign _10094_ = _9391_ ^ _10096_ /*82008*/;
assign _10095_ = _10087_ & _10094_ /*82006*/;
assign _9840_ = _10087_ ^ _10094_ /*82007*/;
assign _10092_ = _10093_ | _10095_ /*82004*/;
assign _10101_ = ~D[48] /*82003*/;
assign _10098_ = _9392_ & _10101_ /*81999*/;
assign _10099_ = _9392_ ^ _10101_ /*82002*/;
assign _10100_ = _10092_ & _10099_ /*82000*/;
assign _9841_ = _10092_ ^ _10099_ /*82001*/;
assign _10097_ = _10098_ | _10100_ /*81998*/;
assign _10106_ = ~D[49] /*81997*/;
assign _10103_ = _9393_ & _10106_ /*81993*/;
assign _10104_ = _9393_ ^ _10106_ /*81996*/;
assign _10105_ = _10097_ & _10104_ /*81994*/;
assign _9842_ = _10097_ ^ _10104_ /*81995*/;
assign _10102_ = _10103_ | _10105_ /*81992*/;
assign _10111_ = ~D[50] /*81991*/;
assign _10108_ = _9394_ & _10111_ /*81987*/;
assign _10109_ = _9394_ ^ _10111_ /*81990*/;
assign _10110_ = _10102_ & _10109_ /*81988*/;
assign _9843_ = _10102_ ^ _10109_ /*81989*/;
assign _10107_ = _10108_ | _10110_ /*81986*/;
assign _10116_ = ~D[51] /*81985*/;
assign _10113_ = _9395_ & _10116_ /*81981*/;
assign _10114_ = _9395_ ^ _10116_ /*81984*/;
assign _10115_ = _10107_ & _10114_ /*81982*/;
assign _9844_ = _10107_ ^ _10114_ /*81983*/;
assign _10112_ = _10113_ | _10115_ /*81980*/;
assign _10121_ = ~D[52] /*81979*/;
assign _10118_ = _9396_ & _10121_ /*81975*/;
assign _10119_ = _9396_ ^ _10121_ /*81978*/;
assign _10120_ = _10112_ & _10119_ /*81976*/;
assign _9845_ = _10112_ ^ _10119_ /*81977*/;
assign _10117_ = _10118_ | _10120_ /*81974*/;
assign _10126_ = ~D[53] /*81973*/;
assign _10123_ = _9397_ & _10126_ /*81969*/;
assign _10124_ = _9397_ ^ _10126_ /*81972*/;
assign _10125_ = _10117_ & _10124_ /*81970*/;
assign _9846_ = _10117_ ^ _10124_ /*81971*/;
assign _10122_ = _10123_ | _10125_ /*81968*/;
assign _10131_ = ~D[54] /*81967*/;
assign _10128_ = _9398_ & _10131_ /*81963*/;
assign _10129_ = _9398_ ^ _10131_ /*81966*/;
assign _10130_ = _10122_ & _10129_ /*81964*/;
assign _9847_ = _10122_ ^ _10129_ /*81965*/;
assign _10127_ = _10128_ | _10130_ /*81962*/;
assign _10136_ = ~D[55] /*81961*/;
assign _10133_ = _9399_ & _10136_ /*81957*/;
assign _10134_ = _9399_ ^ _10136_ /*81960*/;
assign _10135_ = _10127_ & _10134_ /*81958*/;
assign _9848_ = _10127_ ^ _10134_ /*81959*/;
assign _10132_ = _10133_ | _10135_ /*81956*/;
assign _10141_ = ~D[56] /*81955*/;
assign _10138_ = _9400_ & _10141_ /*81951*/;
assign _10139_ = _9400_ ^ _10141_ /*81954*/;
assign _10140_ = _10132_ & _10139_ /*81952*/;
assign _9849_ = _10132_ ^ _10139_ /*81953*/;
assign _10137_ = _10138_ | _10140_ /*81950*/;
assign _10146_ = ~D[57] /*81949*/;
assign _10143_ = _9401_ & _10146_ /*81945*/;
assign _10144_ = _9401_ ^ _10146_ /*81948*/;
assign _10145_ = _10137_ & _10144_ /*81946*/;
assign _9850_ = _10137_ ^ _10144_ /*81947*/;
assign _10142_ = _10143_ | _10145_ /*81944*/;
assign _10151_ = ~D[58] /*81943*/;
assign _10148_ = _9402_ & _10151_ /*81939*/;
assign _10149_ = _9402_ ^ _10151_ /*81942*/;
assign _10150_ = _10142_ & _10149_ /*81940*/;
assign _9851_ = _10142_ ^ _10149_ /*81941*/;
assign _10147_ = _10148_ | _10150_ /*81938*/;
assign _10156_ = ~D[59] /*81937*/;
assign _10153_ = _9403_ & _10156_ /*81933*/;
assign _10154_ = _9403_ ^ _10156_ /*81936*/;
assign _10155_ = _10147_ & _10154_ /*81934*/;
assign _9852_ = _10147_ ^ _10154_ /*81935*/;
assign _10152_ = _10153_ | _10155_ /*81932*/;
assign _10161_ = ~D[60] /*81931*/;
assign _10158_ = _9404_ & _10161_ /*81927*/;
assign _10159_ = _9404_ ^ _10161_ /*81930*/;
assign _10160_ = _10152_ & _10159_ /*81928*/;
assign _9853_ = _10152_ ^ _10159_ /*81929*/;
assign _10157_ = _10158_ | _10160_ /*81926*/;
assign _10166_ = ~D[61] /*81925*/;
assign _10163_ = _9405_ & _10166_ /*81921*/;
assign _10164_ = _9405_ ^ _10166_ /*81924*/;
assign _10165_ = _10157_ & _10164_ /*81922*/;
assign _9854_ = _10157_ ^ _10164_ /*81923*/;
assign _10162_ = _10163_ | _10165_ /*81920*/;
assign _10171_ = ~D[62] /*81919*/;
assign _10168_ = _9406_ & _10171_ /*81915*/;
assign _10169_ = _9406_ ^ _10171_ /*81918*/;
assign _10170_ = _10162_ & _10169_ /*81916*/;
assign _9855_ = _10162_ ^ _10169_ /*81917*/;
assign _10167_ = _10168_ | _10170_ /*81914*/;
assign _10172_ = _9407_ & oneWire /*81909*/;
assign _10173_ = _9407_ ^ oneWire /*81912*/;
assign _10174_ = _10167_ & _10173_ /*81910*/;
assign _9856_ = _10167_ ^ _10173_ /*81911*/;
assign Q[52] = _10172_ | _10174_ /*81908*/;
assign _10307_ = ~Q[52] /*81523*/;
assign _10306_ = _10307_ & D[0] /*81522*/;
assign _10309_ = _9793_ & _10306_ /*81517*/;
assign _10310_ = _9793_ ^ _10306_ /*81520*/;
assign _10311_ = zeroWire & _10310_ /*81518*/;
assign _10241_ = zeroWire ^ _10310_ /*81519*/;
assign _10308_ = _10309_ | _10311_ /*81516*/;
assign _10313_ = ~Q[52] /*81515*/;
assign _10312_ = _10313_ & D[1] /*81514*/;
assign _10315_ = _9794_ & _10312_ /*81509*/;
assign _10316_ = _9794_ ^ _10312_ /*81512*/;
assign _10317_ = _10308_ & _10316_ /*81510*/;
assign _10242_ = _10308_ ^ _10316_ /*81511*/;
assign _10314_ = _10315_ | _10317_ /*81508*/;
assign _10319_ = ~Q[52] /*81507*/;
assign _10318_ = _10319_ & D[2] /*81506*/;
assign _10321_ = _9795_ & _10318_ /*81501*/;
assign _10322_ = _9795_ ^ _10318_ /*81504*/;
assign _10323_ = _10314_ & _10322_ /*81502*/;
assign _10243_ = _10314_ ^ _10322_ /*81503*/;
assign _10320_ = _10321_ | _10323_ /*81500*/;
assign _10325_ = ~Q[52] /*81499*/;
assign _10324_ = _10325_ & D[3] /*81498*/;
assign _10327_ = _9796_ & _10324_ /*81493*/;
assign _10328_ = _9796_ ^ _10324_ /*81496*/;
assign _10329_ = _10320_ & _10328_ /*81494*/;
assign _10244_ = _10320_ ^ _10328_ /*81495*/;
assign _10326_ = _10327_ | _10329_ /*81492*/;
assign _10331_ = ~Q[52] /*81491*/;
assign _10330_ = _10331_ & D[4] /*81490*/;
assign _10333_ = _9797_ & _10330_ /*81485*/;
assign _10334_ = _9797_ ^ _10330_ /*81488*/;
assign _10335_ = _10326_ & _10334_ /*81486*/;
assign _10245_ = _10326_ ^ _10334_ /*81487*/;
assign _10332_ = _10333_ | _10335_ /*81484*/;
assign _10337_ = ~Q[52] /*81483*/;
assign _10336_ = _10337_ & D[5] /*81482*/;
assign _10339_ = _9798_ & _10336_ /*81477*/;
assign _10340_ = _9798_ ^ _10336_ /*81480*/;
assign _10341_ = _10332_ & _10340_ /*81478*/;
assign _10246_ = _10332_ ^ _10340_ /*81479*/;
assign _10338_ = _10339_ | _10341_ /*81476*/;
assign _10343_ = ~Q[52] /*81475*/;
assign _10342_ = _10343_ & D[6] /*81474*/;
assign _10345_ = _9799_ & _10342_ /*81469*/;
assign _10346_ = _9799_ ^ _10342_ /*81472*/;
assign _10347_ = _10338_ & _10346_ /*81470*/;
assign _10247_ = _10338_ ^ _10346_ /*81471*/;
assign _10344_ = _10345_ | _10347_ /*81468*/;
assign _10349_ = ~Q[52] /*81467*/;
assign _10348_ = _10349_ & D[7] /*81466*/;
assign _10351_ = _9800_ & _10348_ /*81461*/;
assign _10352_ = _9800_ ^ _10348_ /*81464*/;
assign _10353_ = _10344_ & _10352_ /*81462*/;
assign _10248_ = _10344_ ^ _10352_ /*81463*/;
assign _10350_ = _10351_ | _10353_ /*81460*/;
assign _10355_ = ~Q[52] /*81459*/;
assign _10354_ = _10355_ & D[8] /*81458*/;
assign _10357_ = _9801_ & _10354_ /*81453*/;
assign _10358_ = _9801_ ^ _10354_ /*81456*/;
assign _10359_ = _10350_ & _10358_ /*81454*/;
assign _10249_ = _10350_ ^ _10358_ /*81455*/;
assign _10356_ = _10357_ | _10359_ /*81452*/;
assign _10361_ = ~Q[52] /*81451*/;
assign _10360_ = _10361_ & D[9] /*81450*/;
assign _10363_ = _9802_ & _10360_ /*81445*/;
assign _10364_ = _9802_ ^ _10360_ /*81448*/;
assign _10365_ = _10356_ & _10364_ /*81446*/;
assign _10250_ = _10356_ ^ _10364_ /*81447*/;
assign _10362_ = _10363_ | _10365_ /*81444*/;
assign _10367_ = ~Q[52] /*81443*/;
assign _10366_ = _10367_ & D[10] /*81442*/;
assign _10369_ = _9803_ & _10366_ /*81437*/;
assign _10370_ = _9803_ ^ _10366_ /*81440*/;
assign _10371_ = _10362_ & _10370_ /*81438*/;
assign _10251_ = _10362_ ^ _10370_ /*81439*/;
assign _10368_ = _10369_ | _10371_ /*81436*/;
assign _10373_ = ~Q[52] /*81435*/;
assign _10372_ = _10373_ & D[11] /*81434*/;
assign _10375_ = _9804_ & _10372_ /*81429*/;
assign _10376_ = _9804_ ^ _10372_ /*81432*/;
assign _10377_ = _10368_ & _10376_ /*81430*/;
assign _10252_ = _10368_ ^ _10376_ /*81431*/;
assign _10374_ = _10375_ | _10377_ /*81428*/;
assign _10379_ = ~Q[52] /*81427*/;
assign _10378_ = _10379_ & D[12] /*81426*/;
assign _10381_ = _9805_ & _10378_ /*81421*/;
assign _10382_ = _9805_ ^ _10378_ /*81424*/;
assign _10383_ = _10374_ & _10382_ /*81422*/;
assign _10253_ = _10374_ ^ _10382_ /*81423*/;
assign _10380_ = _10381_ | _10383_ /*81420*/;
assign _10385_ = ~Q[52] /*81419*/;
assign _10384_ = _10385_ & D[13] /*81418*/;
assign _10387_ = _9806_ & _10384_ /*81413*/;
assign _10388_ = _9806_ ^ _10384_ /*81416*/;
assign _10389_ = _10380_ & _10388_ /*81414*/;
assign _10254_ = _10380_ ^ _10388_ /*81415*/;
assign _10386_ = _10387_ | _10389_ /*81412*/;
assign _10391_ = ~Q[52] /*81411*/;
assign _10390_ = _10391_ & D[14] /*81410*/;
assign _10393_ = _9807_ & _10390_ /*81405*/;
assign _10394_ = _9807_ ^ _10390_ /*81408*/;
assign _10395_ = _10386_ & _10394_ /*81406*/;
assign _10255_ = _10386_ ^ _10394_ /*81407*/;
assign _10392_ = _10393_ | _10395_ /*81404*/;
assign _10397_ = ~Q[52] /*81403*/;
assign _10396_ = _10397_ & D[15] /*81402*/;
assign _10399_ = _9808_ & _10396_ /*81397*/;
assign _10400_ = _9808_ ^ _10396_ /*81400*/;
assign _10401_ = _10392_ & _10400_ /*81398*/;
assign _10256_ = _10392_ ^ _10400_ /*81399*/;
assign _10398_ = _10399_ | _10401_ /*81396*/;
assign _10403_ = ~Q[52] /*81395*/;
assign _10402_ = _10403_ & D[16] /*81394*/;
assign _10405_ = _9809_ & _10402_ /*81389*/;
assign _10406_ = _9809_ ^ _10402_ /*81392*/;
assign _10407_ = _10398_ & _10406_ /*81390*/;
assign _10257_ = _10398_ ^ _10406_ /*81391*/;
assign _10404_ = _10405_ | _10407_ /*81388*/;
assign _10409_ = ~Q[52] /*81387*/;
assign _10408_ = _10409_ & D[17] /*81386*/;
assign _10411_ = _9810_ & _10408_ /*81381*/;
assign _10412_ = _9810_ ^ _10408_ /*81384*/;
assign _10413_ = _10404_ & _10412_ /*81382*/;
assign _10258_ = _10404_ ^ _10412_ /*81383*/;
assign _10410_ = _10411_ | _10413_ /*81380*/;
assign _10415_ = ~Q[52] /*81379*/;
assign _10414_ = _10415_ & D[18] /*81378*/;
assign _10417_ = _9811_ & _10414_ /*81373*/;
assign _10418_ = _9811_ ^ _10414_ /*81376*/;
assign _10419_ = _10410_ & _10418_ /*81374*/;
assign _10259_ = _10410_ ^ _10418_ /*81375*/;
assign _10416_ = _10417_ | _10419_ /*81372*/;
assign _10421_ = ~Q[52] /*81371*/;
assign _10420_ = _10421_ & D[19] /*81370*/;
assign _10423_ = _9812_ & _10420_ /*81365*/;
assign _10424_ = _9812_ ^ _10420_ /*81368*/;
assign _10425_ = _10416_ & _10424_ /*81366*/;
assign _10260_ = _10416_ ^ _10424_ /*81367*/;
assign _10422_ = _10423_ | _10425_ /*81364*/;
assign _10427_ = ~Q[52] /*81363*/;
assign _10426_ = _10427_ & D[20] /*81362*/;
assign _10429_ = _9813_ & _10426_ /*81357*/;
assign _10430_ = _9813_ ^ _10426_ /*81360*/;
assign _10431_ = _10422_ & _10430_ /*81358*/;
assign _10261_ = _10422_ ^ _10430_ /*81359*/;
assign _10428_ = _10429_ | _10431_ /*81356*/;
assign _10433_ = ~Q[52] /*81355*/;
assign _10432_ = _10433_ & D[21] /*81354*/;
assign _10435_ = _9814_ & _10432_ /*81349*/;
assign _10436_ = _9814_ ^ _10432_ /*81352*/;
assign _10437_ = _10428_ & _10436_ /*81350*/;
assign _10262_ = _10428_ ^ _10436_ /*81351*/;
assign _10434_ = _10435_ | _10437_ /*81348*/;
assign _10439_ = ~Q[52] /*81347*/;
assign _10438_ = _10439_ & D[22] /*81346*/;
assign _10441_ = _9815_ & _10438_ /*81341*/;
assign _10442_ = _9815_ ^ _10438_ /*81344*/;
assign _10443_ = _10434_ & _10442_ /*81342*/;
assign _10263_ = _10434_ ^ _10442_ /*81343*/;
assign _10440_ = _10441_ | _10443_ /*81340*/;
assign _10445_ = ~Q[52] /*81339*/;
assign _10444_ = _10445_ & D[23] /*81338*/;
assign _10447_ = _9816_ & _10444_ /*81333*/;
assign _10448_ = _9816_ ^ _10444_ /*81336*/;
assign _10449_ = _10440_ & _10448_ /*81334*/;
assign _10264_ = _10440_ ^ _10448_ /*81335*/;
assign _10446_ = _10447_ | _10449_ /*81332*/;
assign _10451_ = ~Q[52] /*81331*/;
assign _10450_ = _10451_ & D[24] /*81330*/;
assign _10453_ = _9817_ & _10450_ /*81325*/;
assign _10454_ = _9817_ ^ _10450_ /*81328*/;
assign _10455_ = _10446_ & _10454_ /*81326*/;
assign _10265_ = _10446_ ^ _10454_ /*81327*/;
assign _10452_ = _10453_ | _10455_ /*81324*/;
assign _10457_ = ~Q[52] /*81323*/;
assign _10456_ = _10457_ & D[25] /*81322*/;
assign _10459_ = _9818_ & _10456_ /*81317*/;
assign _10460_ = _9818_ ^ _10456_ /*81320*/;
assign _10461_ = _10452_ & _10460_ /*81318*/;
assign _10266_ = _10452_ ^ _10460_ /*81319*/;
assign _10458_ = _10459_ | _10461_ /*81316*/;
assign _10463_ = ~Q[52] /*81315*/;
assign _10462_ = _10463_ & D[26] /*81314*/;
assign _10465_ = _9819_ & _10462_ /*81309*/;
assign _10466_ = _9819_ ^ _10462_ /*81312*/;
assign _10467_ = _10458_ & _10466_ /*81310*/;
assign _10267_ = _10458_ ^ _10466_ /*81311*/;
assign _10464_ = _10465_ | _10467_ /*81308*/;
assign _10469_ = ~Q[52] /*81307*/;
assign _10468_ = _10469_ & D[27] /*81306*/;
assign _10471_ = _9820_ & _10468_ /*81301*/;
assign _10472_ = _9820_ ^ _10468_ /*81304*/;
assign _10473_ = _10464_ & _10472_ /*81302*/;
assign _10268_ = _10464_ ^ _10472_ /*81303*/;
assign _10470_ = _10471_ | _10473_ /*81300*/;
assign _10475_ = ~Q[52] /*81299*/;
assign _10474_ = _10475_ & D[28] /*81298*/;
assign _10477_ = _9821_ & _10474_ /*81293*/;
assign _10478_ = _9821_ ^ _10474_ /*81296*/;
assign _10479_ = _10470_ & _10478_ /*81294*/;
assign _10269_ = _10470_ ^ _10478_ /*81295*/;
assign _10476_ = _10477_ | _10479_ /*81292*/;
assign _10481_ = ~Q[52] /*81291*/;
assign _10480_ = _10481_ & D[29] /*81290*/;
assign _10483_ = _9822_ & _10480_ /*81285*/;
assign _10484_ = _9822_ ^ _10480_ /*81288*/;
assign _10485_ = _10476_ & _10484_ /*81286*/;
assign _10270_ = _10476_ ^ _10484_ /*81287*/;
assign _10482_ = _10483_ | _10485_ /*81284*/;
assign _10487_ = ~Q[52] /*81283*/;
assign _10486_ = _10487_ & D[30] /*81282*/;
assign _10489_ = _9823_ & _10486_ /*81277*/;
assign _10490_ = _9823_ ^ _10486_ /*81280*/;
assign _10491_ = _10482_ & _10490_ /*81278*/;
assign _10271_ = _10482_ ^ _10490_ /*81279*/;
assign _10488_ = _10489_ | _10491_ /*81276*/;
assign _10493_ = ~Q[52] /*81275*/;
assign _10492_ = _10493_ & D[31] /*81274*/;
assign _10495_ = _9824_ & _10492_ /*81269*/;
assign _10496_ = _9824_ ^ _10492_ /*81272*/;
assign _10497_ = _10488_ & _10496_ /*81270*/;
assign _10272_ = _10488_ ^ _10496_ /*81271*/;
assign _10494_ = _10495_ | _10497_ /*81268*/;
assign _10499_ = ~Q[52] /*81267*/;
assign _10498_ = _10499_ & D[32] /*81266*/;
assign _10501_ = _9825_ & _10498_ /*81261*/;
assign _10502_ = _9825_ ^ _10498_ /*81264*/;
assign _10503_ = _10494_ & _10502_ /*81262*/;
assign _10273_ = _10494_ ^ _10502_ /*81263*/;
assign _10500_ = _10501_ | _10503_ /*81260*/;
assign _10505_ = ~Q[52] /*81259*/;
assign _10504_ = _10505_ & D[33] /*81258*/;
assign _10507_ = _9826_ & _10504_ /*81253*/;
assign _10508_ = _9826_ ^ _10504_ /*81256*/;
assign _10509_ = _10500_ & _10508_ /*81254*/;
assign _10274_ = _10500_ ^ _10508_ /*81255*/;
assign _10506_ = _10507_ | _10509_ /*81252*/;
assign _10511_ = ~Q[52] /*81251*/;
assign _10510_ = _10511_ & D[34] /*81250*/;
assign _10513_ = _9827_ & _10510_ /*81245*/;
assign _10514_ = _9827_ ^ _10510_ /*81248*/;
assign _10515_ = _10506_ & _10514_ /*81246*/;
assign _10275_ = _10506_ ^ _10514_ /*81247*/;
assign _10512_ = _10513_ | _10515_ /*81244*/;
assign _10517_ = ~Q[52] /*81243*/;
assign _10516_ = _10517_ & D[35] /*81242*/;
assign _10519_ = _9828_ & _10516_ /*81237*/;
assign _10520_ = _9828_ ^ _10516_ /*81240*/;
assign _10521_ = _10512_ & _10520_ /*81238*/;
assign _10276_ = _10512_ ^ _10520_ /*81239*/;
assign _10518_ = _10519_ | _10521_ /*81236*/;
assign _10523_ = ~Q[52] /*81235*/;
assign _10522_ = _10523_ & D[36] /*81234*/;
assign _10525_ = _9829_ & _10522_ /*81229*/;
assign _10526_ = _9829_ ^ _10522_ /*81232*/;
assign _10527_ = _10518_ & _10526_ /*81230*/;
assign _10277_ = _10518_ ^ _10526_ /*81231*/;
assign _10524_ = _10525_ | _10527_ /*81228*/;
assign _10529_ = ~Q[52] /*81227*/;
assign _10528_ = _10529_ & D[37] /*81226*/;
assign _10531_ = _9830_ & _10528_ /*81221*/;
assign _10532_ = _9830_ ^ _10528_ /*81224*/;
assign _10533_ = _10524_ & _10532_ /*81222*/;
assign _10278_ = _10524_ ^ _10532_ /*81223*/;
assign _10530_ = _10531_ | _10533_ /*81220*/;
assign _10535_ = ~Q[52] /*81219*/;
assign _10534_ = _10535_ & D[38] /*81218*/;
assign _10537_ = _9831_ & _10534_ /*81213*/;
assign _10538_ = _9831_ ^ _10534_ /*81216*/;
assign _10539_ = _10530_ & _10538_ /*81214*/;
assign _10279_ = _10530_ ^ _10538_ /*81215*/;
assign _10536_ = _10537_ | _10539_ /*81212*/;
assign _10541_ = ~Q[52] /*81211*/;
assign _10540_ = _10541_ & D[39] /*81210*/;
assign _10543_ = _9832_ & _10540_ /*81205*/;
assign _10544_ = _9832_ ^ _10540_ /*81208*/;
assign _10545_ = _10536_ & _10544_ /*81206*/;
assign _10280_ = _10536_ ^ _10544_ /*81207*/;
assign _10542_ = _10543_ | _10545_ /*81204*/;
assign _10547_ = ~Q[52] /*81203*/;
assign _10546_ = _10547_ & D[40] /*81202*/;
assign _10549_ = _9833_ & _10546_ /*81197*/;
assign _10550_ = _9833_ ^ _10546_ /*81200*/;
assign _10551_ = _10542_ & _10550_ /*81198*/;
assign _10281_ = _10542_ ^ _10550_ /*81199*/;
assign _10548_ = _10549_ | _10551_ /*81196*/;
assign _10553_ = ~Q[52] /*81195*/;
assign _10552_ = _10553_ & D[41] /*81194*/;
assign _10555_ = _9834_ & _10552_ /*81189*/;
assign _10556_ = _9834_ ^ _10552_ /*81192*/;
assign _10557_ = _10548_ & _10556_ /*81190*/;
assign _10282_ = _10548_ ^ _10556_ /*81191*/;
assign _10554_ = _10555_ | _10557_ /*81188*/;
assign _10559_ = ~Q[52] /*81187*/;
assign _10558_ = _10559_ & D[42] /*81186*/;
assign _10561_ = _9835_ & _10558_ /*81181*/;
assign _10562_ = _9835_ ^ _10558_ /*81184*/;
assign _10563_ = _10554_ & _10562_ /*81182*/;
assign _10283_ = _10554_ ^ _10562_ /*81183*/;
assign _10560_ = _10561_ | _10563_ /*81180*/;
assign _10565_ = ~Q[52] /*81179*/;
assign _10564_ = _10565_ & D[43] /*81178*/;
assign _10567_ = _9836_ & _10564_ /*81173*/;
assign _10568_ = _9836_ ^ _10564_ /*81176*/;
assign _10569_ = _10560_ & _10568_ /*81174*/;
assign _10284_ = _10560_ ^ _10568_ /*81175*/;
assign _10566_ = _10567_ | _10569_ /*81172*/;
assign _10571_ = ~Q[52] /*81171*/;
assign _10570_ = _10571_ & D[44] /*81170*/;
assign _10573_ = _9837_ & _10570_ /*81165*/;
assign _10574_ = _9837_ ^ _10570_ /*81168*/;
assign _10575_ = _10566_ & _10574_ /*81166*/;
assign _10285_ = _10566_ ^ _10574_ /*81167*/;
assign _10572_ = _10573_ | _10575_ /*81164*/;
assign _10577_ = ~Q[52] /*81163*/;
assign _10576_ = _10577_ & D[45] /*81162*/;
assign _10579_ = _9838_ & _10576_ /*81157*/;
assign _10580_ = _9838_ ^ _10576_ /*81160*/;
assign _10581_ = _10572_ & _10580_ /*81158*/;
assign _10286_ = _10572_ ^ _10580_ /*81159*/;
assign _10578_ = _10579_ | _10581_ /*81156*/;
assign _10583_ = ~Q[52] /*81155*/;
assign _10582_ = _10583_ & D[46] /*81154*/;
assign _10585_ = _9839_ & _10582_ /*81149*/;
assign _10586_ = _9839_ ^ _10582_ /*81152*/;
assign _10587_ = _10578_ & _10586_ /*81150*/;
assign _10287_ = _10578_ ^ _10586_ /*81151*/;
assign _10584_ = _10585_ | _10587_ /*81148*/;
assign _10589_ = ~Q[52] /*81147*/;
assign _10588_ = _10589_ & D[47] /*81146*/;
assign _10591_ = _9840_ & _10588_ /*81141*/;
assign _10592_ = _9840_ ^ _10588_ /*81144*/;
assign _10593_ = _10584_ & _10592_ /*81142*/;
assign _10288_ = _10584_ ^ _10592_ /*81143*/;
assign _10590_ = _10591_ | _10593_ /*81140*/;
assign _10595_ = ~Q[52] /*81139*/;
assign _10594_ = _10595_ & D[48] /*81138*/;
assign _10597_ = _9841_ & _10594_ /*81133*/;
assign _10598_ = _9841_ ^ _10594_ /*81136*/;
assign _10599_ = _10590_ & _10598_ /*81134*/;
assign _10289_ = _10590_ ^ _10598_ /*81135*/;
assign _10596_ = _10597_ | _10599_ /*81132*/;
assign _10601_ = ~Q[52] /*81131*/;
assign _10600_ = _10601_ & D[49] /*81130*/;
assign _10603_ = _9842_ & _10600_ /*81125*/;
assign _10604_ = _9842_ ^ _10600_ /*81128*/;
assign _10605_ = _10596_ & _10604_ /*81126*/;
assign _10290_ = _10596_ ^ _10604_ /*81127*/;
assign _10602_ = _10603_ | _10605_ /*81124*/;
assign _10607_ = ~Q[52] /*81123*/;
assign _10606_ = _10607_ & D[50] /*81122*/;
assign _10609_ = _9843_ & _10606_ /*81117*/;
assign _10610_ = _9843_ ^ _10606_ /*81120*/;
assign _10611_ = _10602_ & _10610_ /*81118*/;
assign _10291_ = _10602_ ^ _10610_ /*81119*/;
assign _10608_ = _10609_ | _10611_ /*81116*/;
assign _10613_ = ~Q[52] /*81115*/;
assign _10612_ = _10613_ & D[51] /*81114*/;
assign _10615_ = _9844_ & _10612_ /*81109*/;
assign _10616_ = _9844_ ^ _10612_ /*81112*/;
assign _10617_ = _10608_ & _10616_ /*81110*/;
assign _10292_ = _10608_ ^ _10616_ /*81111*/;
assign _10614_ = _10615_ | _10617_ /*81108*/;
assign _10619_ = ~Q[52] /*81107*/;
assign _10618_ = _10619_ & D[52] /*81106*/;
assign _10621_ = _9845_ & _10618_ /*81101*/;
assign _10622_ = _9845_ ^ _10618_ /*81104*/;
assign _10623_ = _10614_ & _10622_ /*81102*/;
assign _10293_ = _10614_ ^ _10622_ /*81103*/;
assign _10620_ = _10621_ | _10623_ /*81100*/;
assign _10625_ = ~Q[52] /*81099*/;
assign _10624_ = _10625_ & D[53] /*81098*/;
assign _10627_ = _9846_ & _10624_ /*81093*/;
assign _10628_ = _9846_ ^ _10624_ /*81096*/;
assign _10629_ = _10620_ & _10628_ /*81094*/;
assign _10294_ = _10620_ ^ _10628_ /*81095*/;
assign _10626_ = _10627_ | _10629_ /*81092*/;
assign _10631_ = ~Q[52] /*81091*/;
assign _10630_ = _10631_ & D[54] /*81090*/;
assign _10633_ = _9847_ & _10630_ /*81085*/;
assign _10634_ = _9847_ ^ _10630_ /*81088*/;
assign _10635_ = _10626_ & _10634_ /*81086*/;
assign _10295_ = _10626_ ^ _10634_ /*81087*/;
assign _10632_ = _10633_ | _10635_ /*81084*/;
assign _10637_ = ~Q[52] /*81083*/;
assign _10636_ = _10637_ & D[55] /*81082*/;
assign _10639_ = _9848_ & _10636_ /*81077*/;
assign _10640_ = _9848_ ^ _10636_ /*81080*/;
assign _10641_ = _10632_ & _10640_ /*81078*/;
assign _10296_ = _10632_ ^ _10640_ /*81079*/;
assign _10638_ = _10639_ | _10641_ /*81076*/;
assign _10643_ = ~Q[52] /*81075*/;
assign _10642_ = _10643_ & D[56] /*81074*/;
assign _10645_ = _9849_ & _10642_ /*81069*/;
assign _10646_ = _9849_ ^ _10642_ /*81072*/;
assign _10647_ = _10638_ & _10646_ /*81070*/;
assign _10297_ = _10638_ ^ _10646_ /*81071*/;
assign _10644_ = _10645_ | _10647_ /*81068*/;
assign _10649_ = ~Q[52] /*81067*/;
assign _10648_ = _10649_ & D[57] /*81066*/;
assign _10651_ = _9850_ & _10648_ /*81061*/;
assign _10652_ = _9850_ ^ _10648_ /*81064*/;
assign _10653_ = _10644_ & _10652_ /*81062*/;
assign _10298_ = _10644_ ^ _10652_ /*81063*/;
assign _10650_ = _10651_ | _10653_ /*81060*/;
assign _10655_ = ~Q[52] /*81059*/;
assign _10654_ = _10655_ & D[58] /*81058*/;
assign _10657_ = _9851_ & _10654_ /*81053*/;
assign _10658_ = _9851_ ^ _10654_ /*81056*/;
assign _10659_ = _10650_ & _10658_ /*81054*/;
assign _10299_ = _10650_ ^ _10658_ /*81055*/;
assign _10656_ = _10657_ | _10659_ /*81052*/;
assign _10661_ = ~Q[52] /*81051*/;
assign _10660_ = _10661_ & D[59] /*81050*/;
assign _10663_ = _9852_ & _10660_ /*81045*/;
assign _10664_ = _9852_ ^ _10660_ /*81048*/;
assign _10665_ = _10656_ & _10664_ /*81046*/;
assign _10300_ = _10656_ ^ _10664_ /*81047*/;
assign _10662_ = _10663_ | _10665_ /*81044*/;
assign _10667_ = ~Q[52] /*81043*/;
assign _10666_ = _10667_ & D[60] /*81042*/;
assign _10669_ = _9853_ & _10666_ /*81037*/;
assign _10670_ = _9853_ ^ _10666_ /*81040*/;
assign _10671_ = _10662_ & _10670_ /*81038*/;
assign _10301_ = _10662_ ^ _10670_ /*81039*/;
assign _10668_ = _10669_ | _10671_ /*81036*/;
assign _10673_ = ~Q[52] /*81035*/;
assign _10672_ = _10673_ & D[61] /*81034*/;
assign _10675_ = _9854_ & _10672_ /*81029*/;
assign _10676_ = _9854_ ^ _10672_ /*81032*/;
assign _10677_ = _10668_ & _10676_ /*81030*/;
assign _10302_ = _10668_ ^ _10676_ /*81031*/;
assign _10674_ = _10675_ | _10677_ /*81028*/;
assign _10679_ = ~Q[52] /*81027*/;
assign _10678_ = _10679_ & D[62] /*81026*/;
assign _10681_ = _9855_ & _10678_ /*81021*/;
assign _10682_ = _9855_ ^ _10678_ /*81024*/;
assign _10683_ = _10674_ & _10682_ /*81022*/;
assign _10303_ = _10674_ ^ _10682_ /*81023*/;
assign _10680_ = _10681_ | _10683_ /*81020*/;
assign _10685_ = ~Q[52] /*81019*/;
assign _10684_ = _10685_ & zeroWire /*81018*/;
assign _10686_ = _9856_ ^ _10684_ /*81016*/;
assign _10304_ = _10686_ ^ _10680_ /*81015*/;
assign _10757_ = ~D[0] /*80761*/;
assign _10754_ = R_0[51] & _10757_ /*80757*/;
assign _10755_ = R_0[51] ^ _10757_ /*80760*/;
assign _10756_ = oneWire & _10755_ /*80758*/;
assign _10689_ = oneWire ^ _10755_ /*80759*/;
assign _10753_ = _10754_ | _10756_ /*80756*/;
assign _10762_ = ~D[1] /*80755*/;
assign _10759_ = _10241_ & _10762_ /*80751*/;
assign _10760_ = _10241_ ^ _10762_ /*80754*/;
assign _10761_ = _10753_ & _10760_ /*80752*/;
assign _10690_ = _10753_ ^ _10760_ /*80753*/;
assign _10758_ = _10759_ | _10761_ /*80750*/;
assign _10767_ = ~D[2] /*80749*/;
assign _10764_ = _10242_ & _10767_ /*80745*/;
assign _10765_ = _10242_ ^ _10767_ /*80748*/;
assign _10766_ = _10758_ & _10765_ /*80746*/;
assign _10691_ = _10758_ ^ _10765_ /*80747*/;
assign _10763_ = _10764_ | _10766_ /*80744*/;
assign _10772_ = ~D[3] /*80743*/;
assign _10769_ = _10243_ & _10772_ /*80739*/;
assign _10770_ = _10243_ ^ _10772_ /*80742*/;
assign _10771_ = _10763_ & _10770_ /*80740*/;
assign _10692_ = _10763_ ^ _10770_ /*80741*/;
assign _10768_ = _10769_ | _10771_ /*80738*/;
assign _10777_ = ~D[4] /*80737*/;
assign _10774_ = _10244_ & _10777_ /*80733*/;
assign _10775_ = _10244_ ^ _10777_ /*80736*/;
assign _10776_ = _10768_ & _10775_ /*80734*/;
assign _10693_ = _10768_ ^ _10775_ /*80735*/;
assign _10773_ = _10774_ | _10776_ /*80732*/;
assign _10782_ = ~D[5] /*80731*/;
assign _10779_ = _10245_ & _10782_ /*80727*/;
assign _10780_ = _10245_ ^ _10782_ /*80730*/;
assign _10781_ = _10773_ & _10780_ /*80728*/;
assign _10694_ = _10773_ ^ _10780_ /*80729*/;
assign _10778_ = _10779_ | _10781_ /*80726*/;
assign _10787_ = ~D[6] /*80725*/;
assign _10784_ = _10246_ & _10787_ /*80721*/;
assign _10785_ = _10246_ ^ _10787_ /*80724*/;
assign _10786_ = _10778_ & _10785_ /*80722*/;
assign _10695_ = _10778_ ^ _10785_ /*80723*/;
assign _10783_ = _10784_ | _10786_ /*80720*/;
assign _10792_ = ~D[7] /*80719*/;
assign _10789_ = _10247_ & _10792_ /*80715*/;
assign _10790_ = _10247_ ^ _10792_ /*80718*/;
assign _10791_ = _10783_ & _10790_ /*80716*/;
assign _10696_ = _10783_ ^ _10790_ /*80717*/;
assign _10788_ = _10789_ | _10791_ /*80714*/;
assign _10797_ = ~D[8] /*80713*/;
assign _10794_ = _10248_ & _10797_ /*80709*/;
assign _10795_ = _10248_ ^ _10797_ /*80712*/;
assign _10796_ = _10788_ & _10795_ /*80710*/;
assign _10697_ = _10788_ ^ _10795_ /*80711*/;
assign _10793_ = _10794_ | _10796_ /*80708*/;
assign _10802_ = ~D[9] /*80707*/;
assign _10799_ = _10249_ & _10802_ /*80703*/;
assign _10800_ = _10249_ ^ _10802_ /*80706*/;
assign _10801_ = _10793_ & _10800_ /*80704*/;
assign _10698_ = _10793_ ^ _10800_ /*80705*/;
assign _10798_ = _10799_ | _10801_ /*80702*/;
assign _10807_ = ~D[10] /*80701*/;
assign _10804_ = _10250_ & _10807_ /*80697*/;
assign _10805_ = _10250_ ^ _10807_ /*80700*/;
assign _10806_ = _10798_ & _10805_ /*80698*/;
assign _10699_ = _10798_ ^ _10805_ /*80699*/;
assign _10803_ = _10804_ | _10806_ /*80696*/;
assign _10812_ = ~D[11] /*80695*/;
assign _10809_ = _10251_ & _10812_ /*80691*/;
assign _10810_ = _10251_ ^ _10812_ /*80694*/;
assign _10811_ = _10803_ & _10810_ /*80692*/;
assign _10700_ = _10803_ ^ _10810_ /*80693*/;
assign _10808_ = _10809_ | _10811_ /*80690*/;
assign _10817_ = ~D[12] /*80689*/;
assign _10814_ = _10252_ & _10817_ /*80685*/;
assign _10815_ = _10252_ ^ _10817_ /*80688*/;
assign _10816_ = _10808_ & _10815_ /*80686*/;
assign _10701_ = _10808_ ^ _10815_ /*80687*/;
assign _10813_ = _10814_ | _10816_ /*80684*/;
assign _10822_ = ~D[13] /*80683*/;
assign _10819_ = _10253_ & _10822_ /*80679*/;
assign _10820_ = _10253_ ^ _10822_ /*80682*/;
assign _10821_ = _10813_ & _10820_ /*80680*/;
assign _10702_ = _10813_ ^ _10820_ /*80681*/;
assign _10818_ = _10819_ | _10821_ /*80678*/;
assign _10827_ = ~D[14] /*80677*/;
assign _10824_ = _10254_ & _10827_ /*80673*/;
assign _10825_ = _10254_ ^ _10827_ /*80676*/;
assign _10826_ = _10818_ & _10825_ /*80674*/;
assign _10703_ = _10818_ ^ _10825_ /*80675*/;
assign _10823_ = _10824_ | _10826_ /*80672*/;
assign _10832_ = ~D[15] /*80671*/;
assign _10829_ = _10255_ & _10832_ /*80667*/;
assign _10830_ = _10255_ ^ _10832_ /*80670*/;
assign _10831_ = _10823_ & _10830_ /*80668*/;
assign _10704_ = _10823_ ^ _10830_ /*80669*/;
assign _10828_ = _10829_ | _10831_ /*80666*/;
assign _10837_ = ~D[16] /*80665*/;
assign _10834_ = _10256_ & _10837_ /*80661*/;
assign _10835_ = _10256_ ^ _10837_ /*80664*/;
assign _10836_ = _10828_ & _10835_ /*80662*/;
assign _10705_ = _10828_ ^ _10835_ /*80663*/;
assign _10833_ = _10834_ | _10836_ /*80660*/;
assign _10842_ = ~D[17] /*80659*/;
assign _10839_ = _10257_ & _10842_ /*80655*/;
assign _10840_ = _10257_ ^ _10842_ /*80658*/;
assign _10841_ = _10833_ & _10840_ /*80656*/;
assign _10706_ = _10833_ ^ _10840_ /*80657*/;
assign _10838_ = _10839_ | _10841_ /*80654*/;
assign _10847_ = ~D[18] /*80653*/;
assign _10844_ = _10258_ & _10847_ /*80649*/;
assign _10845_ = _10258_ ^ _10847_ /*80652*/;
assign _10846_ = _10838_ & _10845_ /*80650*/;
assign _10707_ = _10838_ ^ _10845_ /*80651*/;
assign _10843_ = _10844_ | _10846_ /*80648*/;
assign _10852_ = ~D[19] /*80647*/;
assign _10849_ = _10259_ & _10852_ /*80643*/;
assign _10850_ = _10259_ ^ _10852_ /*80646*/;
assign _10851_ = _10843_ & _10850_ /*80644*/;
assign _10708_ = _10843_ ^ _10850_ /*80645*/;
assign _10848_ = _10849_ | _10851_ /*80642*/;
assign _10857_ = ~D[20] /*80641*/;
assign _10854_ = _10260_ & _10857_ /*80637*/;
assign _10855_ = _10260_ ^ _10857_ /*80640*/;
assign _10856_ = _10848_ & _10855_ /*80638*/;
assign _10709_ = _10848_ ^ _10855_ /*80639*/;
assign _10853_ = _10854_ | _10856_ /*80636*/;
assign _10862_ = ~D[21] /*80635*/;
assign _10859_ = _10261_ & _10862_ /*80631*/;
assign _10860_ = _10261_ ^ _10862_ /*80634*/;
assign _10861_ = _10853_ & _10860_ /*80632*/;
assign _10710_ = _10853_ ^ _10860_ /*80633*/;
assign _10858_ = _10859_ | _10861_ /*80630*/;
assign _10867_ = ~D[22] /*80629*/;
assign _10864_ = _10262_ & _10867_ /*80625*/;
assign _10865_ = _10262_ ^ _10867_ /*80628*/;
assign _10866_ = _10858_ & _10865_ /*80626*/;
assign _10711_ = _10858_ ^ _10865_ /*80627*/;
assign _10863_ = _10864_ | _10866_ /*80624*/;
assign _10872_ = ~D[23] /*80623*/;
assign _10869_ = _10263_ & _10872_ /*80619*/;
assign _10870_ = _10263_ ^ _10872_ /*80622*/;
assign _10871_ = _10863_ & _10870_ /*80620*/;
assign _10712_ = _10863_ ^ _10870_ /*80621*/;
assign _10868_ = _10869_ | _10871_ /*80618*/;
assign _10877_ = ~D[24] /*80617*/;
assign _10874_ = _10264_ & _10877_ /*80613*/;
assign _10875_ = _10264_ ^ _10877_ /*80616*/;
assign _10876_ = _10868_ & _10875_ /*80614*/;
assign _10713_ = _10868_ ^ _10875_ /*80615*/;
assign _10873_ = _10874_ | _10876_ /*80612*/;
assign _10882_ = ~D[25] /*80611*/;
assign _10879_ = _10265_ & _10882_ /*80607*/;
assign _10880_ = _10265_ ^ _10882_ /*80610*/;
assign _10881_ = _10873_ & _10880_ /*80608*/;
assign _10714_ = _10873_ ^ _10880_ /*80609*/;
assign _10878_ = _10879_ | _10881_ /*80606*/;
assign _10887_ = ~D[26] /*80605*/;
assign _10884_ = _10266_ & _10887_ /*80601*/;
assign _10885_ = _10266_ ^ _10887_ /*80604*/;
assign _10886_ = _10878_ & _10885_ /*80602*/;
assign _10715_ = _10878_ ^ _10885_ /*80603*/;
assign _10883_ = _10884_ | _10886_ /*80600*/;
assign _10892_ = ~D[27] /*80599*/;
assign _10889_ = _10267_ & _10892_ /*80595*/;
assign _10890_ = _10267_ ^ _10892_ /*80598*/;
assign _10891_ = _10883_ & _10890_ /*80596*/;
assign _10716_ = _10883_ ^ _10890_ /*80597*/;
assign _10888_ = _10889_ | _10891_ /*80594*/;
assign _10897_ = ~D[28] /*80593*/;
assign _10894_ = _10268_ & _10897_ /*80589*/;
assign _10895_ = _10268_ ^ _10897_ /*80592*/;
assign _10896_ = _10888_ & _10895_ /*80590*/;
assign _10717_ = _10888_ ^ _10895_ /*80591*/;
assign _10893_ = _10894_ | _10896_ /*80588*/;
assign _10902_ = ~D[29] /*80587*/;
assign _10899_ = _10269_ & _10902_ /*80583*/;
assign _10900_ = _10269_ ^ _10902_ /*80586*/;
assign _10901_ = _10893_ & _10900_ /*80584*/;
assign _10718_ = _10893_ ^ _10900_ /*80585*/;
assign _10898_ = _10899_ | _10901_ /*80582*/;
assign _10907_ = ~D[30] /*80581*/;
assign _10904_ = _10270_ & _10907_ /*80577*/;
assign _10905_ = _10270_ ^ _10907_ /*80580*/;
assign _10906_ = _10898_ & _10905_ /*80578*/;
assign _10719_ = _10898_ ^ _10905_ /*80579*/;
assign _10903_ = _10904_ | _10906_ /*80576*/;
assign _10912_ = ~D[31] /*80575*/;
assign _10909_ = _10271_ & _10912_ /*80571*/;
assign _10910_ = _10271_ ^ _10912_ /*80574*/;
assign _10911_ = _10903_ & _10910_ /*80572*/;
assign _10720_ = _10903_ ^ _10910_ /*80573*/;
assign _10908_ = _10909_ | _10911_ /*80570*/;
assign _10917_ = ~D[32] /*80569*/;
assign _10914_ = _10272_ & _10917_ /*80565*/;
assign _10915_ = _10272_ ^ _10917_ /*80568*/;
assign _10916_ = _10908_ & _10915_ /*80566*/;
assign _10721_ = _10908_ ^ _10915_ /*80567*/;
assign _10913_ = _10914_ | _10916_ /*80564*/;
assign _10922_ = ~D[33] /*80563*/;
assign _10919_ = _10273_ & _10922_ /*80559*/;
assign _10920_ = _10273_ ^ _10922_ /*80562*/;
assign _10921_ = _10913_ & _10920_ /*80560*/;
assign _10722_ = _10913_ ^ _10920_ /*80561*/;
assign _10918_ = _10919_ | _10921_ /*80558*/;
assign _10927_ = ~D[34] /*80557*/;
assign _10924_ = _10274_ & _10927_ /*80553*/;
assign _10925_ = _10274_ ^ _10927_ /*80556*/;
assign _10926_ = _10918_ & _10925_ /*80554*/;
assign _10723_ = _10918_ ^ _10925_ /*80555*/;
assign _10923_ = _10924_ | _10926_ /*80552*/;
assign _10932_ = ~D[35] /*80551*/;
assign _10929_ = _10275_ & _10932_ /*80547*/;
assign _10930_ = _10275_ ^ _10932_ /*80550*/;
assign _10931_ = _10923_ & _10930_ /*80548*/;
assign _10724_ = _10923_ ^ _10930_ /*80549*/;
assign _10928_ = _10929_ | _10931_ /*80546*/;
assign _10937_ = ~D[36] /*80545*/;
assign _10934_ = _10276_ & _10937_ /*80541*/;
assign _10935_ = _10276_ ^ _10937_ /*80544*/;
assign _10936_ = _10928_ & _10935_ /*80542*/;
assign _10725_ = _10928_ ^ _10935_ /*80543*/;
assign _10933_ = _10934_ | _10936_ /*80540*/;
assign _10942_ = ~D[37] /*80539*/;
assign _10939_ = _10277_ & _10942_ /*80535*/;
assign _10940_ = _10277_ ^ _10942_ /*80538*/;
assign _10941_ = _10933_ & _10940_ /*80536*/;
assign _10726_ = _10933_ ^ _10940_ /*80537*/;
assign _10938_ = _10939_ | _10941_ /*80534*/;
assign _10947_ = ~D[38] /*80533*/;
assign _10944_ = _10278_ & _10947_ /*80529*/;
assign _10945_ = _10278_ ^ _10947_ /*80532*/;
assign _10946_ = _10938_ & _10945_ /*80530*/;
assign _10727_ = _10938_ ^ _10945_ /*80531*/;
assign _10943_ = _10944_ | _10946_ /*80528*/;
assign _10952_ = ~D[39] /*80527*/;
assign _10949_ = _10279_ & _10952_ /*80523*/;
assign _10950_ = _10279_ ^ _10952_ /*80526*/;
assign _10951_ = _10943_ & _10950_ /*80524*/;
assign _10728_ = _10943_ ^ _10950_ /*80525*/;
assign _10948_ = _10949_ | _10951_ /*80522*/;
assign _10957_ = ~D[40] /*80521*/;
assign _10954_ = _10280_ & _10957_ /*80517*/;
assign _10955_ = _10280_ ^ _10957_ /*80520*/;
assign _10956_ = _10948_ & _10955_ /*80518*/;
assign _10729_ = _10948_ ^ _10955_ /*80519*/;
assign _10953_ = _10954_ | _10956_ /*80516*/;
assign _10962_ = ~D[41] /*80515*/;
assign _10959_ = _10281_ & _10962_ /*80511*/;
assign _10960_ = _10281_ ^ _10962_ /*80514*/;
assign _10961_ = _10953_ & _10960_ /*80512*/;
assign _10730_ = _10953_ ^ _10960_ /*80513*/;
assign _10958_ = _10959_ | _10961_ /*80510*/;
assign _10967_ = ~D[42] /*80509*/;
assign _10964_ = _10282_ & _10967_ /*80505*/;
assign _10965_ = _10282_ ^ _10967_ /*80508*/;
assign _10966_ = _10958_ & _10965_ /*80506*/;
assign _10731_ = _10958_ ^ _10965_ /*80507*/;
assign _10963_ = _10964_ | _10966_ /*80504*/;
assign _10972_ = ~D[43] /*80503*/;
assign _10969_ = _10283_ & _10972_ /*80499*/;
assign _10970_ = _10283_ ^ _10972_ /*80502*/;
assign _10971_ = _10963_ & _10970_ /*80500*/;
assign _10732_ = _10963_ ^ _10970_ /*80501*/;
assign _10968_ = _10969_ | _10971_ /*80498*/;
assign _10977_ = ~D[44] /*80497*/;
assign _10974_ = _10284_ & _10977_ /*80493*/;
assign _10975_ = _10284_ ^ _10977_ /*80496*/;
assign _10976_ = _10968_ & _10975_ /*80494*/;
assign _10733_ = _10968_ ^ _10975_ /*80495*/;
assign _10973_ = _10974_ | _10976_ /*80492*/;
assign _10982_ = ~D[45] /*80491*/;
assign _10979_ = _10285_ & _10982_ /*80487*/;
assign _10980_ = _10285_ ^ _10982_ /*80490*/;
assign _10981_ = _10973_ & _10980_ /*80488*/;
assign _10734_ = _10973_ ^ _10980_ /*80489*/;
assign _10978_ = _10979_ | _10981_ /*80486*/;
assign _10987_ = ~D[46] /*80485*/;
assign _10984_ = _10286_ & _10987_ /*80481*/;
assign _10985_ = _10286_ ^ _10987_ /*80484*/;
assign _10986_ = _10978_ & _10985_ /*80482*/;
assign _10735_ = _10978_ ^ _10985_ /*80483*/;
assign _10983_ = _10984_ | _10986_ /*80480*/;
assign _10992_ = ~D[47] /*80479*/;
assign _10989_ = _10287_ & _10992_ /*80475*/;
assign _10990_ = _10287_ ^ _10992_ /*80478*/;
assign _10991_ = _10983_ & _10990_ /*80476*/;
assign _10736_ = _10983_ ^ _10990_ /*80477*/;
assign _10988_ = _10989_ | _10991_ /*80474*/;
assign _10997_ = ~D[48] /*80473*/;
assign _10994_ = _10288_ & _10997_ /*80469*/;
assign _10995_ = _10288_ ^ _10997_ /*80472*/;
assign _10996_ = _10988_ & _10995_ /*80470*/;
assign _10737_ = _10988_ ^ _10995_ /*80471*/;
assign _10993_ = _10994_ | _10996_ /*80468*/;
assign _11002_ = ~D[49] /*80467*/;
assign _10999_ = _10289_ & _11002_ /*80463*/;
assign _11000_ = _10289_ ^ _11002_ /*80466*/;
assign _11001_ = _10993_ & _11000_ /*80464*/;
assign _10738_ = _10993_ ^ _11000_ /*80465*/;
assign _10998_ = _10999_ | _11001_ /*80462*/;
assign _11007_ = ~D[50] /*80461*/;
assign _11004_ = _10290_ & _11007_ /*80457*/;
assign _11005_ = _10290_ ^ _11007_ /*80460*/;
assign _11006_ = _10998_ & _11005_ /*80458*/;
assign _10739_ = _10998_ ^ _11005_ /*80459*/;
assign _11003_ = _11004_ | _11006_ /*80456*/;
assign _11012_ = ~D[51] /*80455*/;
assign _11009_ = _10291_ & _11012_ /*80451*/;
assign _11010_ = _10291_ ^ _11012_ /*80454*/;
assign _11011_ = _11003_ & _11010_ /*80452*/;
assign _10740_ = _11003_ ^ _11010_ /*80453*/;
assign _11008_ = _11009_ | _11011_ /*80450*/;
assign _11017_ = ~D[52] /*80449*/;
assign _11014_ = _10292_ & _11017_ /*80445*/;
assign _11015_ = _10292_ ^ _11017_ /*80448*/;
assign _11016_ = _11008_ & _11015_ /*80446*/;
assign _10741_ = _11008_ ^ _11015_ /*80447*/;
assign _11013_ = _11014_ | _11016_ /*80444*/;
assign _11022_ = ~D[53] /*80443*/;
assign _11019_ = _10293_ & _11022_ /*80439*/;
assign _11020_ = _10293_ ^ _11022_ /*80442*/;
assign _11021_ = _11013_ & _11020_ /*80440*/;
assign _10742_ = _11013_ ^ _11020_ /*80441*/;
assign _11018_ = _11019_ | _11021_ /*80438*/;
assign _11027_ = ~D[54] /*80437*/;
assign _11024_ = _10294_ & _11027_ /*80433*/;
assign _11025_ = _10294_ ^ _11027_ /*80436*/;
assign _11026_ = _11018_ & _11025_ /*80434*/;
assign _10743_ = _11018_ ^ _11025_ /*80435*/;
assign _11023_ = _11024_ | _11026_ /*80432*/;
assign _11032_ = ~D[55] /*80431*/;
assign _11029_ = _10295_ & _11032_ /*80427*/;
assign _11030_ = _10295_ ^ _11032_ /*80430*/;
assign _11031_ = _11023_ & _11030_ /*80428*/;
assign _10744_ = _11023_ ^ _11030_ /*80429*/;
assign _11028_ = _11029_ | _11031_ /*80426*/;
assign _11037_ = ~D[56] /*80425*/;
assign _11034_ = _10296_ & _11037_ /*80421*/;
assign _11035_ = _10296_ ^ _11037_ /*80424*/;
assign _11036_ = _11028_ & _11035_ /*80422*/;
assign _10745_ = _11028_ ^ _11035_ /*80423*/;
assign _11033_ = _11034_ | _11036_ /*80420*/;
assign _11042_ = ~D[57] /*80419*/;
assign _11039_ = _10297_ & _11042_ /*80415*/;
assign _11040_ = _10297_ ^ _11042_ /*80418*/;
assign _11041_ = _11033_ & _11040_ /*80416*/;
assign _10746_ = _11033_ ^ _11040_ /*80417*/;
assign _11038_ = _11039_ | _11041_ /*80414*/;
assign _11047_ = ~D[58] /*80413*/;
assign _11044_ = _10298_ & _11047_ /*80409*/;
assign _11045_ = _10298_ ^ _11047_ /*80412*/;
assign _11046_ = _11038_ & _11045_ /*80410*/;
assign _10747_ = _11038_ ^ _11045_ /*80411*/;
assign _11043_ = _11044_ | _11046_ /*80408*/;
assign _11052_ = ~D[59] /*80407*/;
assign _11049_ = _10299_ & _11052_ /*80403*/;
assign _11050_ = _10299_ ^ _11052_ /*80406*/;
assign _11051_ = _11043_ & _11050_ /*80404*/;
assign _10748_ = _11043_ ^ _11050_ /*80405*/;
assign _11048_ = _11049_ | _11051_ /*80402*/;
assign _11057_ = ~D[60] /*80401*/;
assign _11054_ = _10300_ & _11057_ /*80397*/;
assign _11055_ = _10300_ ^ _11057_ /*80400*/;
assign _11056_ = _11048_ & _11055_ /*80398*/;
assign _10749_ = _11048_ ^ _11055_ /*80399*/;
assign _11053_ = _11054_ | _11056_ /*80396*/;
assign _11062_ = ~D[61] /*80395*/;
assign _11059_ = _10301_ & _11062_ /*80391*/;
assign _11060_ = _10301_ ^ _11062_ /*80394*/;
assign _11061_ = _11053_ & _11060_ /*80392*/;
assign _10750_ = _11053_ ^ _11060_ /*80393*/;
assign _11058_ = _11059_ | _11061_ /*80390*/;
assign _11067_ = ~D[62] /*80389*/;
assign _11064_ = _10302_ & _11067_ /*80385*/;
assign _11065_ = _10302_ ^ _11067_ /*80388*/;
assign _11066_ = _11058_ & _11065_ /*80386*/;
assign _10751_ = _11058_ ^ _11065_ /*80387*/;
assign _11063_ = _11064_ | _11066_ /*80384*/;
assign _11068_ = _10303_ & oneWire /*80379*/;
assign _11069_ = _10303_ ^ oneWire /*80382*/;
assign _11070_ = _11063_ & _11069_ /*80380*/;
assign _10752_ = _11063_ ^ _11069_ /*80381*/;
assign Q[51] = _11068_ | _11070_ /*80378*/;
assign _11203_ = ~Q[51] /*79993*/;
assign _11202_ = _11203_ & D[0] /*79992*/;
assign _11205_ = _10689_ & _11202_ /*79987*/;
assign _11206_ = _10689_ ^ _11202_ /*79990*/;
assign _11207_ = zeroWire & _11206_ /*79988*/;
assign _11137_ = zeroWire ^ _11206_ /*79989*/;
assign _11204_ = _11205_ | _11207_ /*79986*/;
assign _11209_ = ~Q[51] /*79985*/;
assign _11208_ = _11209_ & D[1] /*79984*/;
assign _11211_ = _10690_ & _11208_ /*79979*/;
assign _11212_ = _10690_ ^ _11208_ /*79982*/;
assign _11213_ = _11204_ & _11212_ /*79980*/;
assign _11138_ = _11204_ ^ _11212_ /*79981*/;
assign _11210_ = _11211_ | _11213_ /*79978*/;
assign _11215_ = ~Q[51] /*79977*/;
assign _11214_ = _11215_ & D[2] /*79976*/;
assign _11217_ = _10691_ & _11214_ /*79971*/;
assign _11218_ = _10691_ ^ _11214_ /*79974*/;
assign _11219_ = _11210_ & _11218_ /*79972*/;
assign _11139_ = _11210_ ^ _11218_ /*79973*/;
assign _11216_ = _11217_ | _11219_ /*79970*/;
assign _11221_ = ~Q[51] /*79969*/;
assign _11220_ = _11221_ & D[3] /*79968*/;
assign _11223_ = _10692_ & _11220_ /*79963*/;
assign _11224_ = _10692_ ^ _11220_ /*79966*/;
assign _11225_ = _11216_ & _11224_ /*79964*/;
assign _11140_ = _11216_ ^ _11224_ /*79965*/;
assign _11222_ = _11223_ | _11225_ /*79962*/;
assign _11227_ = ~Q[51] /*79961*/;
assign _11226_ = _11227_ & D[4] /*79960*/;
assign _11229_ = _10693_ & _11226_ /*79955*/;
assign _11230_ = _10693_ ^ _11226_ /*79958*/;
assign _11231_ = _11222_ & _11230_ /*79956*/;
assign _11141_ = _11222_ ^ _11230_ /*79957*/;
assign _11228_ = _11229_ | _11231_ /*79954*/;
assign _11233_ = ~Q[51] /*79953*/;
assign _11232_ = _11233_ & D[5] /*79952*/;
assign _11235_ = _10694_ & _11232_ /*79947*/;
assign _11236_ = _10694_ ^ _11232_ /*79950*/;
assign _11237_ = _11228_ & _11236_ /*79948*/;
assign _11142_ = _11228_ ^ _11236_ /*79949*/;
assign _11234_ = _11235_ | _11237_ /*79946*/;
assign _11239_ = ~Q[51] /*79945*/;
assign _11238_ = _11239_ & D[6] /*79944*/;
assign _11241_ = _10695_ & _11238_ /*79939*/;
assign _11242_ = _10695_ ^ _11238_ /*79942*/;
assign _11243_ = _11234_ & _11242_ /*79940*/;
assign _11143_ = _11234_ ^ _11242_ /*79941*/;
assign _11240_ = _11241_ | _11243_ /*79938*/;
assign _11245_ = ~Q[51] /*79937*/;
assign _11244_ = _11245_ & D[7] /*79936*/;
assign _11247_ = _10696_ & _11244_ /*79931*/;
assign _11248_ = _10696_ ^ _11244_ /*79934*/;
assign _11249_ = _11240_ & _11248_ /*79932*/;
assign _11144_ = _11240_ ^ _11248_ /*79933*/;
assign _11246_ = _11247_ | _11249_ /*79930*/;
assign _11251_ = ~Q[51] /*79929*/;
assign _11250_ = _11251_ & D[8] /*79928*/;
assign _11253_ = _10697_ & _11250_ /*79923*/;
assign _11254_ = _10697_ ^ _11250_ /*79926*/;
assign _11255_ = _11246_ & _11254_ /*79924*/;
assign _11145_ = _11246_ ^ _11254_ /*79925*/;
assign _11252_ = _11253_ | _11255_ /*79922*/;
assign _11257_ = ~Q[51] /*79921*/;
assign _11256_ = _11257_ & D[9] /*79920*/;
assign _11259_ = _10698_ & _11256_ /*79915*/;
assign _11260_ = _10698_ ^ _11256_ /*79918*/;
assign _11261_ = _11252_ & _11260_ /*79916*/;
assign _11146_ = _11252_ ^ _11260_ /*79917*/;
assign _11258_ = _11259_ | _11261_ /*79914*/;
assign _11263_ = ~Q[51] /*79913*/;
assign _11262_ = _11263_ & D[10] /*79912*/;
assign _11265_ = _10699_ & _11262_ /*79907*/;
assign _11266_ = _10699_ ^ _11262_ /*79910*/;
assign _11267_ = _11258_ & _11266_ /*79908*/;
assign _11147_ = _11258_ ^ _11266_ /*79909*/;
assign _11264_ = _11265_ | _11267_ /*79906*/;
assign _11269_ = ~Q[51] /*79905*/;
assign _11268_ = _11269_ & D[11] /*79904*/;
assign _11271_ = _10700_ & _11268_ /*79899*/;
assign _11272_ = _10700_ ^ _11268_ /*79902*/;
assign _11273_ = _11264_ & _11272_ /*79900*/;
assign _11148_ = _11264_ ^ _11272_ /*79901*/;
assign _11270_ = _11271_ | _11273_ /*79898*/;
assign _11275_ = ~Q[51] /*79897*/;
assign _11274_ = _11275_ & D[12] /*79896*/;
assign _11277_ = _10701_ & _11274_ /*79891*/;
assign _11278_ = _10701_ ^ _11274_ /*79894*/;
assign _11279_ = _11270_ & _11278_ /*79892*/;
assign _11149_ = _11270_ ^ _11278_ /*79893*/;
assign _11276_ = _11277_ | _11279_ /*79890*/;
assign _11281_ = ~Q[51] /*79889*/;
assign _11280_ = _11281_ & D[13] /*79888*/;
assign _11283_ = _10702_ & _11280_ /*79883*/;
assign _11284_ = _10702_ ^ _11280_ /*79886*/;
assign _11285_ = _11276_ & _11284_ /*79884*/;
assign _11150_ = _11276_ ^ _11284_ /*79885*/;
assign _11282_ = _11283_ | _11285_ /*79882*/;
assign _11287_ = ~Q[51] /*79881*/;
assign _11286_ = _11287_ & D[14] /*79880*/;
assign _11289_ = _10703_ & _11286_ /*79875*/;
assign _11290_ = _10703_ ^ _11286_ /*79878*/;
assign _11291_ = _11282_ & _11290_ /*79876*/;
assign _11151_ = _11282_ ^ _11290_ /*79877*/;
assign _11288_ = _11289_ | _11291_ /*79874*/;
assign _11293_ = ~Q[51] /*79873*/;
assign _11292_ = _11293_ & D[15] /*79872*/;
assign _11295_ = _10704_ & _11292_ /*79867*/;
assign _11296_ = _10704_ ^ _11292_ /*79870*/;
assign _11297_ = _11288_ & _11296_ /*79868*/;
assign _11152_ = _11288_ ^ _11296_ /*79869*/;
assign _11294_ = _11295_ | _11297_ /*79866*/;
assign _11299_ = ~Q[51] /*79865*/;
assign _11298_ = _11299_ & D[16] /*79864*/;
assign _11301_ = _10705_ & _11298_ /*79859*/;
assign _11302_ = _10705_ ^ _11298_ /*79862*/;
assign _11303_ = _11294_ & _11302_ /*79860*/;
assign _11153_ = _11294_ ^ _11302_ /*79861*/;
assign _11300_ = _11301_ | _11303_ /*79858*/;
assign _11305_ = ~Q[51] /*79857*/;
assign _11304_ = _11305_ & D[17] /*79856*/;
assign _11307_ = _10706_ & _11304_ /*79851*/;
assign _11308_ = _10706_ ^ _11304_ /*79854*/;
assign _11309_ = _11300_ & _11308_ /*79852*/;
assign _11154_ = _11300_ ^ _11308_ /*79853*/;
assign _11306_ = _11307_ | _11309_ /*79850*/;
assign _11311_ = ~Q[51] /*79849*/;
assign _11310_ = _11311_ & D[18] /*79848*/;
assign _11313_ = _10707_ & _11310_ /*79843*/;
assign _11314_ = _10707_ ^ _11310_ /*79846*/;
assign _11315_ = _11306_ & _11314_ /*79844*/;
assign _11155_ = _11306_ ^ _11314_ /*79845*/;
assign _11312_ = _11313_ | _11315_ /*79842*/;
assign _11317_ = ~Q[51] /*79841*/;
assign _11316_ = _11317_ & D[19] /*79840*/;
assign _11319_ = _10708_ & _11316_ /*79835*/;
assign _11320_ = _10708_ ^ _11316_ /*79838*/;
assign _11321_ = _11312_ & _11320_ /*79836*/;
assign _11156_ = _11312_ ^ _11320_ /*79837*/;
assign _11318_ = _11319_ | _11321_ /*79834*/;
assign _11323_ = ~Q[51] /*79833*/;
assign _11322_ = _11323_ & D[20] /*79832*/;
assign _11325_ = _10709_ & _11322_ /*79827*/;
assign _11326_ = _10709_ ^ _11322_ /*79830*/;
assign _11327_ = _11318_ & _11326_ /*79828*/;
assign _11157_ = _11318_ ^ _11326_ /*79829*/;
assign _11324_ = _11325_ | _11327_ /*79826*/;
assign _11329_ = ~Q[51] /*79825*/;
assign _11328_ = _11329_ & D[21] /*79824*/;
assign _11331_ = _10710_ & _11328_ /*79819*/;
assign _11332_ = _10710_ ^ _11328_ /*79822*/;
assign _11333_ = _11324_ & _11332_ /*79820*/;
assign _11158_ = _11324_ ^ _11332_ /*79821*/;
assign _11330_ = _11331_ | _11333_ /*79818*/;
assign _11335_ = ~Q[51] /*79817*/;
assign _11334_ = _11335_ & D[22] /*79816*/;
assign _11337_ = _10711_ & _11334_ /*79811*/;
assign _11338_ = _10711_ ^ _11334_ /*79814*/;
assign _11339_ = _11330_ & _11338_ /*79812*/;
assign _11159_ = _11330_ ^ _11338_ /*79813*/;
assign _11336_ = _11337_ | _11339_ /*79810*/;
assign _11341_ = ~Q[51] /*79809*/;
assign _11340_ = _11341_ & D[23] /*79808*/;
assign _11343_ = _10712_ & _11340_ /*79803*/;
assign _11344_ = _10712_ ^ _11340_ /*79806*/;
assign _11345_ = _11336_ & _11344_ /*79804*/;
assign _11160_ = _11336_ ^ _11344_ /*79805*/;
assign _11342_ = _11343_ | _11345_ /*79802*/;
assign _11347_ = ~Q[51] /*79801*/;
assign _11346_ = _11347_ & D[24] /*79800*/;
assign _11349_ = _10713_ & _11346_ /*79795*/;
assign _11350_ = _10713_ ^ _11346_ /*79798*/;
assign _11351_ = _11342_ & _11350_ /*79796*/;
assign _11161_ = _11342_ ^ _11350_ /*79797*/;
assign _11348_ = _11349_ | _11351_ /*79794*/;
assign _11353_ = ~Q[51] /*79793*/;
assign _11352_ = _11353_ & D[25] /*79792*/;
assign _11355_ = _10714_ & _11352_ /*79787*/;
assign _11356_ = _10714_ ^ _11352_ /*79790*/;
assign _11357_ = _11348_ & _11356_ /*79788*/;
assign _11162_ = _11348_ ^ _11356_ /*79789*/;
assign _11354_ = _11355_ | _11357_ /*79786*/;
assign _11359_ = ~Q[51] /*79785*/;
assign _11358_ = _11359_ & D[26] /*79784*/;
assign _11361_ = _10715_ & _11358_ /*79779*/;
assign _11362_ = _10715_ ^ _11358_ /*79782*/;
assign _11363_ = _11354_ & _11362_ /*79780*/;
assign _11163_ = _11354_ ^ _11362_ /*79781*/;
assign _11360_ = _11361_ | _11363_ /*79778*/;
assign _11365_ = ~Q[51] /*79777*/;
assign _11364_ = _11365_ & D[27] /*79776*/;
assign _11367_ = _10716_ & _11364_ /*79771*/;
assign _11368_ = _10716_ ^ _11364_ /*79774*/;
assign _11369_ = _11360_ & _11368_ /*79772*/;
assign _11164_ = _11360_ ^ _11368_ /*79773*/;
assign _11366_ = _11367_ | _11369_ /*79770*/;
assign _11371_ = ~Q[51] /*79769*/;
assign _11370_ = _11371_ & D[28] /*79768*/;
assign _11373_ = _10717_ & _11370_ /*79763*/;
assign _11374_ = _10717_ ^ _11370_ /*79766*/;
assign _11375_ = _11366_ & _11374_ /*79764*/;
assign _11165_ = _11366_ ^ _11374_ /*79765*/;
assign _11372_ = _11373_ | _11375_ /*79762*/;
assign _11377_ = ~Q[51] /*79761*/;
assign _11376_ = _11377_ & D[29] /*79760*/;
assign _11379_ = _10718_ & _11376_ /*79755*/;
assign _11380_ = _10718_ ^ _11376_ /*79758*/;
assign _11381_ = _11372_ & _11380_ /*79756*/;
assign _11166_ = _11372_ ^ _11380_ /*79757*/;
assign _11378_ = _11379_ | _11381_ /*79754*/;
assign _11383_ = ~Q[51] /*79753*/;
assign _11382_ = _11383_ & D[30] /*79752*/;
assign _11385_ = _10719_ & _11382_ /*79747*/;
assign _11386_ = _10719_ ^ _11382_ /*79750*/;
assign _11387_ = _11378_ & _11386_ /*79748*/;
assign _11167_ = _11378_ ^ _11386_ /*79749*/;
assign _11384_ = _11385_ | _11387_ /*79746*/;
assign _11389_ = ~Q[51] /*79745*/;
assign _11388_ = _11389_ & D[31] /*79744*/;
assign _11391_ = _10720_ & _11388_ /*79739*/;
assign _11392_ = _10720_ ^ _11388_ /*79742*/;
assign _11393_ = _11384_ & _11392_ /*79740*/;
assign _11168_ = _11384_ ^ _11392_ /*79741*/;
assign _11390_ = _11391_ | _11393_ /*79738*/;
assign _11395_ = ~Q[51] /*79737*/;
assign _11394_ = _11395_ & D[32] /*79736*/;
assign _11397_ = _10721_ & _11394_ /*79731*/;
assign _11398_ = _10721_ ^ _11394_ /*79734*/;
assign _11399_ = _11390_ & _11398_ /*79732*/;
assign _11169_ = _11390_ ^ _11398_ /*79733*/;
assign _11396_ = _11397_ | _11399_ /*79730*/;
assign _11401_ = ~Q[51] /*79729*/;
assign _11400_ = _11401_ & D[33] /*79728*/;
assign _11403_ = _10722_ & _11400_ /*79723*/;
assign _11404_ = _10722_ ^ _11400_ /*79726*/;
assign _11405_ = _11396_ & _11404_ /*79724*/;
assign _11170_ = _11396_ ^ _11404_ /*79725*/;
assign _11402_ = _11403_ | _11405_ /*79722*/;
assign _11407_ = ~Q[51] /*79721*/;
assign _11406_ = _11407_ & D[34] /*79720*/;
assign _11409_ = _10723_ & _11406_ /*79715*/;
assign _11410_ = _10723_ ^ _11406_ /*79718*/;
assign _11411_ = _11402_ & _11410_ /*79716*/;
assign _11171_ = _11402_ ^ _11410_ /*79717*/;
assign _11408_ = _11409_ | _11411_ /*79714*/;
assign _11413_ = ~Q[51] /*79713*/;
assign _11412_ = _11413_ & D[35] /*79712*/;
assign _11415_ = _10724_ & _11412_ /*79707*/;
assign _11416_ = _10724_ ^ _11412_ /*79710*/;
assign _11417_ = _11408_ & _11416_ /*79708*/;
assign _11172_ = _11408_ ^ _11416_ /*79709*/;
assign _11414_ = _11415_ | _11417_ /*79706*/;
assign _11419_ = ~Q[51] /*79705*/;
assign _11418_ = _11419_ & D[36] /*79704*/;
assign _11421_ = _10725_ & _11418_ /*79699*/;
assign _11422_ = _10725_ ^ _11418_ /*79702*/;
assign _11423_ = _11414_ & _11422_ /*79700*/;
assign _11173_ = _11414_ ^ _11422_ /*79701*/;
assign _11420_ = _11421_ | _11423_ /*79698*/;
assign _11425_ = ~Q[51] /*79697*/;
assign _11424_ = _11425_ & D[37] /*79696*/;
assign _11427_ = _10726_ & _11424_ /*79691*/;
assign _11428_ = _10726_ ^ _11424_ /*79694*/;
assign _11429_ = _11420_ & _11428_ /*79692*/;
assign _11174_ = _11420_ ^ _11428_ /*79693*/;
assign _11426_ = _11427_ | _11429_ /*79690*/;
assign _11431_ = ~Q[51] /*79689*/;
assign _11430_ = _11431_ & D[38] /*79688*/;
assign _11433_ = _10727_ & _11430_ /*79683*/;
assign _11434_ = _10727_ ^ _11430_ /*79686*/;
assign _11435_ = _11426_ & _11434_ /*79684*/;
assign _11175_ = _11426_ ^ _11434_ /*79685*/;
assign _11432_ = _11433_ | _11435_ /*79682*/;
assign _11437_ = ~Q[51] /*79681*/;
assign _11436_ = _11437_ & D[39] /*79680*/;
assign _11439_ = _10728_ & _11436_ /*79675*/;
assign _11440_ = _10728_ ^ _11436_ /*79678*/;
assign _11441_ = _11432_ & _11440_ /*79676*/;
assign _11176_ = _11432_ ^ _11440_ /*79677*/;
assign _11438_ = _11439_ | _11441_ /*79674*/;
assign _11443_ = ~Q[51] /*79673*/;
assign _11442_ = _11443_ & D[40] /*79672*/;
assign _11445_ = _10729_ & _11442_ /*79667*/;
assign _11446_ = _10729_ ^ _11442_ /*79670*/;
assign _11447_ = _11438_ & _11446_ /*79668*/;
assign _11177_ = _11438_ ^ _11446_ /*79669*/;
assign _11444_ = _11445_ | _11447_ /*79666*/;
assign _11449_ = ~Q[51] /*79665*/;
assign _11448_ = _11449_ & D[41] /*79664*/;
assign _11451_ = _10730_ & _11448_ /*79659*/;
assign _11452_ = _10730_ ^ _11448_ /*79662*/;
assign _11453_ = _11444_ & _11452_ /*79660*/;
assign _11178_ = _11444_ ^ _11452_ /*79661*/;
assign _11450_ = _11451_ | _11453_ /*79658*/;
assign _11455_ = ~Q[51] /*79657*/;
assign _11454_ = _11455_ & D[42] /*79656*/;
assign _11457_ = _10731_ & _11454_ /*79651*/;
assign _11458_ = _10731_ ^ _11454_ /*79654*/;
assign _11459_ = _11450_ & _11458_ /*79652*/;
assign _11179_ = _11450_ ^ _11458_ /*79653*/;
assign _11456_ = _11457_ | _11459_ /*79650*/;
assign _11461_ = ~Q[51] /*79649*/;
assign _11460_ = _11461_ & D[43] /*79648*/;
assign _11463_ = _10732_ & _11460_ /*79643*/;
assign _11464_ = _10732_ ^ _11460_ /*79646*/;
assign _11465_ = _11456_ & _11464_ /*79644*/;
assign _11180_ = _11456_ ^ _11464_ /*79645*/;
assign _11462_ = _11463_ | _11465_ /*79642*/;
assign _11467_ = ~Q[51] /*79641*/;
assign _11466_ = _11467_ & D[44] /*79640*/;
assign _11469_ = _10733_ & _11466_ /*79635*/;
assign _11470_ = _10733_ ^ _11466_ /*79638*/;
assign _11471_ = _11462_ & _11470_ /*79636*/;
assign _11181_ = _11462_ ^ _11470_ /*79637*/;
assign _11468_ = _11469_ | _11471_ /*79634*/;
assign _11473_ = ~Q[51] /*79633*/;
assign _11472_ = _11473_ & D[45] /*79632*/;
assign _11475_ = _10734_ & _11472_ /*79627*/;
assign _11476_ = _10734_ ^ _11472_ /*79630*/;
assign _11477_ = _11468_ & _11476_ /*79628*/;
assign _11182_ = _11468_ ^ _11476_ /*79629*/;
assign _11474_ = _11475_ | _11477_ /*79626*/;
assign _11479_ = ~Q[51] /*79625*/;
assign _11478_ = _11479_ & D[46] /*79624*/;
assign _11481_ = _10735_ & _11478_ /*79619*/;
assign _11482_ = _10735_ ^ _11478_ /*79622*/;
assign _11483_ = _11474_ & _11482_ /*79620*/;
assign _11183_ = _11474_ ^ _11482_ /*79621*/;
assign _11480_ = _11481_ | _11483_ /*79618*/;
assign _11485_ = ~Q[51] /*79617*/;
assign _11484_ = _11485_ & D[47] /*79616*/;
assign _11487_ = _10736_ & _11484_ /*79611*/;
assign _11488_ = _10736_ ^ _11484_ /*79614*/;
assign _11489_ = _11480_ & _11488_ /*79612*/;
assign _11184_ = _11480_ ^ _11488_ /*79613*/;
assign _11486_ = _11487_ | _11489_ /*79610*/;
assign _11491_ = ~Q[51] /*79609*/;
assign _11490_ = _11491_ & D[48] /*79608*/;
assign _11493_ = _10737_ & _11490_ /*79603*/;
assign _11494_ = _10737_ ^ _11490_ /*79606*/;
assign _11495_ = _11486_ & _11494_ /*79604*/;
assign _11185_ = _11486_ ^ _11494_ /*79605*/;
assign _11492_ = _11493_ | _11495_ /*79602*/;
assign _11497_ = ~Q[51] /*79601*/;
assign _11496_ = _11497_ & D[49] /*79600*/;
assign _11499_ = _10738_ & _11496_ /*79595*/;
assign _11500_ = _10738_ ^ _11496_ /*79598*/;
assign _11501_ = _11492_ & _11500_ /*79596*/;
assign _11186_ = _11492_ ^ _11500_ /*79597*/;
assign _11498_ = _11499_ | _11501_ /*79594*/;
assign _11503_ = ~Q[51] /*79593*/;
assign _11502_ = _11503_ & D[50] /*79592*/;
assign _11505_ = _10739_ & _11502_ /*79587*/;
assign _11506_ = _10739_ ^ _11502_ /*79590*/;
assign _11507_ = _11498_ & _11506_ /*79588*/;
assign _11187_ = _11498_ ^ _11506_ /*79589*/;
assign _11504_ = _11505_ | _11507_ /*79586*/;
assign _11509_ = ~Q[51] /*79585*/;
assign _11508_ = _11509_ & D[51] /*79584*/;
assign _11511_ = _10740_ & _11508_ /*79579*/;
assign _11512_ = _10740_ ^ _11508_ /*79582*/;
assign _11513_ = _11504_ & _11512_ /*79580*/;
assign _11188_ = _11504_ ^ _11512_ /*79581*/;
assign _11510_ = _11511_ | _11513_ /*79578*/;
assign _11515_ = ~Q[51] /*79577*/;
assign _11514_ = _11515_ & D[52] /*79576*/;
assign _11517_ = _10741_ & _11514_ /*79571*/;
assign _11518_ = _10741_ ^ _11514_ /*79574*/;
assign _11519_ = _11510_ & _11518_ /*79572*/;
assign _11189_ = _11510_ ^ _11518_ /*79573*/;
assign _11516_ = _11517_ | _11519_ /*79570*/;
assign _11521_ = ~Q[51] /*79569*/;
assign _11520_ = _11521_ & D[53] /*79568*/;
assign _11523_ = _10742_ & _11520_ /*79563*/;
assign _11524_ = _10742_ ^ _11520_ /*79566*/;
assign _11525_ = _11516_ & _11524_ /*79564*/;
assign _11190_ = _11516_ ^ _11524_ /*79565*/;
assign _11522_ = _11523_ | _11525_ /*79562*/;
assign _11527_ = ~Q[51] /*79561*/;
assign _11526_ = _11527_ & D[54] /*79560*/;
assign _11529_ = _10743_ & _11526_ /*79555*/;
assign _11530_ = _10743_ ^ _11526_ /*79558*/;
assign _11531_ = _11522_ & _11530_ /*79556*/;
assign _11191_ = _11522_ ^ _11530_ /*79557*/;
assign _11528_ = _11529_ | _11531_ /*79554*/;
assign _11533_ = ~Q[51] /*79553*/;
assign _11532_ = _11533_ & D[55] /*79552*/;
assign _11535_ = _10744_ & _11532_ /*79547*/;
assign _11536_ = _10744_ ^ _11532_ /*79550*/;
assign _11537_ = _11528_ & _11536_ /*79548*/;
assign _11192_ = _11528_ ^ _11536_ /*79549*/;
assign _11534_ = _11535_ | _11537_ /*79546*/;
assign _11539_ = ~Q[51] /*79545*/;
assign _11538_ = _11539_ & D[56] /*79544*/;
assign _11541_ = _10745_ & _11538_ /*79539*/;
assign _11542_ = _10745_ ^ _11538_ /*79542*/;
assign _11543_ = _11534_ & _11542_ /*79540*/;
assign _11193_ = _11534_ ^ _11542_ /*79541*/;
assign _11540_ = _11541_ | _11543_ /*79538*/;
assign _11545_ = ~Q[51] /*79537*/;
assign _11544_ = _11545_ & D[57] /*79536*/;
assign _11547_ = _10746_ & _11544_ /*79531*/;
assign _11548_ = _10746_ ^ _11544_ /*79534*/;
assign _11549_ = _11540_ & _11548_ /*79532*/;
assign _11194_ = _11540_ ^ _11548_ /*79533*/;
assign _11546_ = _11547_ | _11549_ /*79530*/;
assign _11551_ = ~Q[51] /*79529*/;
assign _11550_ = _11551_ & D[58] /*79528*/;
assign _11553_ = _10747_ & _11550_ /*79523*/;
assign _11554_ = _10747_ ^ _11550_ /*79526*/;
assign _11555_ = _11546_ & _11554_ /*79524*/;
assign _11195_ = _11546_ ^ _11554_ /*79525*/;
assign _11552_ = _11553_ | _11555_ /*79522*/;
assign _11557_ = ~Q[51] /*79521*/;
assign _11556_ = _11557_ & D[59] /*79520*/;
assign _11559_ = _10748_ & _11556_ /*79515*/;
assign _11560_ = _10748_ ^ _11556_ /*79518*/;
assign _11561_ = _11552_ & _11560_ /*79516*/;
assign _11196_ = _11552_ ^ _11560_ /*79517*/;
assign _11558_ = _11559_ | _11561_ /*79514*/;
assign _11563_ = ~Q[51] /*79513*/;
assign _11562_ = _11563_ & D[60] /*79512*/;
assign _11565_ = _10749_ & _11562_ /*79507*/;
assign _11566_ = _10749_ ^ _11562_ /*79510*/;
assign _11567_ = _11558_ & _11566_ /*79508*/;
assign _11197_ = _11558_ ^ _11566_ /*79509*/;
assign _11564_ = _11565_ | _11567_ /*79506*/;
assign _11569_ = ~Q[51] /*79505*/;
assign _11568_ = _11569_ & D[61] /*79504*/;
assign _11571_ = _10750_ & _11568_ /*79499*/;
assign _11572_ = _10750_ ^ _11568_ /*79502*/;
assign _11573_ = _11564_ & _11572_ /*79500*/;
assign _11198_ = _11564_ ^ _11572_ /*79501*/;
assign _11570_ = _11571_ | _11573_ /*79498*/;
assign _11575_ = ~Q[51] /*79497*/;
assign _11574_ = _11575_ & D[62] /*79496*/;
assign _11577_ = _10751_ & _11574_ /*79491*/;
assign _11578_ = _10751_ ^ _11574_ /*79494*/;
assign _11579_ = _11570_ & _11578_ /*79492*/;
assign _11199_ = _11570_ ^ _11578_ /*79493*/;
assign _11576_ = _11577_ | _11579_ /*79490*/;
assign _11581_ = ~Q[51] /*79489*/;
assign _11580_ = _11581_ & zeroWire /*79488*/;
assign _11582_ = _10752_ ^ _11580_ /*79486*/;
assign _11200_ = _11582_ ^ _11576_ /*79485*/;
assign _11653_ = ~D[0] /*79231*/;
assign _11650_ = R_0[50] & _11653_ /*79227*/;
assign _11651_ = R_0[50] ^ _11653_ /*79230*/;
assign _11652_ = oneWire & _11651_ /*79228*/;
assign _11585_ = oneWire ^ _11651_ /*79229*/;
assign _11649_ = _11650_ | _11652_ /*79226*/;
assign _11658_ = ~D[1] /*79225*/;
assign _11655_ = _11137_ & _11658_ /*79221*/;
assign _11656_ = _11137_ ^ _11658_ /*79224*/;
assign _11657_ = _11649_ & _11656_ /*79222*/;
assign _11586_ = _11649_ ^ _11656_ /*79223*/;
assign _11654_ = _11655_ | _11657_ /*79220*/;
assign _11663_ = ~D[2] /*79219*/;
assign _11660_ = _11138_ & _11663_ /*79215*/;
assign _11661_ = _11138_ ^ _11663_ /*79218*/;
assign _11662_ = _11654_ & _11661_ /*79216*/;
assign _11587_ = _11654_ ^ _11661_ /*79217*/;
assign _11659_ = _11660_ | _11662_ /*79214*/;
assign _11668_ = ~D[3] /*79213*/;
assign _11665_ = _11139_ & _11668_ /*79209*/;
assign _11666_ = _11139_ ^ _11668_ /*79212*/;
assign _11667_ = _11659_ & _11666_ /*79210*/;
assign _11588_ = _11659_ ^ _11666_ /*79211*/;
assign _11664_ = _11665_ | _11667_ /*79208*/;
assign _11673_ = ~D[4] /*79207*/;
assign _11670_ = _11140_ & _11673_ /*79203*/;
assign _11671_ = _11140_ ^ _11673_ /*79206*/;
assign _11672_ = _11664_ & _11671_ /*79204*/;
assign _11589_ = _11664_ ^ _11671_ /*79205*/;
assign _11669_ = _11670_ | _11672_ /*79202*/;
assign _11678_ = ~D[5] /*79201*/;
assign _11675_ = _11141_ & _11678_ /*79197*/;
assign _11676_ = _11141_ ^ _11678_ /*79200*/;
assign _11677_ = _11669_ & _11676_ /*79198*/;
assign _11590_ = _11669_ ^ _11676_ /*79199*/;
assign _11674_ = _11675_ | _11677_ /*79196*/;
assign _11683_ = ~D[6] /*79195*/;
assign _11680_ = _11142_ & _11683_ /*79191*/;
assign _11681_ = _11142_ ^ _11683_ /*79194*/;
assign _11682_ = _11674_ & _11681_ /*79192*/;
assign _11591_ = _11674_ ^ _11681_ /*79193*/;
assign _11679_ = _11680_ | _11682_ /*79190*/;
assign _11688_ = ~D[7] /*79189*/;
assign _11685_ = _11143_ & _11688_ /*79185*/;
assign _11686_ = _11143_ ^ _11688_ /*79188*/;
assign _11687_ = _11679_ & _11686_ /*79186*/;
assign _11592_ = _11679_ ^ _11686_ /*79187*/;
assign _11684_ = _11685_ | _11687_ /*79184*/;
assign _11693_ = ~D[8] /*79183*/;
assign _11690_ = _11144_ & _11693_ /*79179*/;
assign _11691_ = _11144_ ^ _11693_ /*79182*/;
assign _11692_ = _11684_ & _11691_ /*79180*/;
assign _11593_ = _11684_ ^ _11691_ /*79181*/;
assign _11689_ = _11690_ | _11692_ /*79178*/;
assign _11698_ = ~D[9] /*79177*/;
assign _11695_ = _11145_ & _11698_ /*79173*/;
assign _11696_ = _11145_ ^ _11698_ /*79176*/;
assign _11697_ = _11689_ & _11696_ /*79174*/;
assign _11594_ = _11689_ ^ _11696_ /*79175*/;
assign _11694_ = _11695_ | _11697_ /*79172*/;
assign _11703_ = ~D[10] /*79171*/;
assign _11700_ = _11146_ & _11703_ /*79167*/;
assign _11701_ = _11146_ ^ _11703_ /*79170*/;
assign _11702_ = _11694_ & _11701_ /*79168*/;
assign _11595_ = _11694_ ^ _11701_ /*79169*/;
assign _11699_ = _11700_ | _11702_ /*79166*/;
assign _11708_ = ~D[11] /*79165*/;
assign _11705_ = _11147_ & _11708_ /*79161*/;
assign _11706_ = _11147_ ^ _11708_ /*79164*/;
assign _11707_ = _11699_ & _11706_ /*79162*/;
assign _11596_ = _11699_ ^ _11706_ /*79163*/;
assign _11704_ = _11705_ | _11707_ /*79160*/;
assign _11713_ = ~D[12] /*79159*/;
assign _11710_ = _11148_ & _11713_ /*79155*/;
assign _11711_ = _11148_ ^ _11713_ /*79158*/;
assign _11712_ = _11704_ & _11711_ /*79156*/;
assign _11597_ = _11704_ ^ _11711_ /*79157*/;
assign _11709_ = _11710_ | _11712_ /*79154*/;
assign _11718_ = ~D[13] /*79153*/;
assign _11715_ = _11149_ & _11718_ /*79149*/;
assign _11716_ = _11149_ ^ _11718_ /*79152*/;
assign _11717_ = _11709_ & _11716_ /*79150*/;
assign _11598_ = _11709_ ^ _11716_ /*79151*/;
assign _11714_ = _11715_ | _11717_ /*79148*/;
assign _11723_ = ~D[14] /*79147*/;
assign _11720_ = _11150_ & _11723_ /*79143*/;
assign _11721_ = _11150_ ^ _11723_ /*79146*/;
assign _11722_ = _11714_ & _11721_ /*79144*/;
assign _11599_ = _11714_ ^ _11721_ /*79145*/;
assign _11719_ = _11720_ | _11722_ /*79142*/;
assign _11728_ = ~D[15] /*79141*/;
assign _11725_ = _11151_ & _11728_ /*79137*/;
assign _11726_ = _11151_ ^ _11728_ /*79140*/;
assign _11727_ = _11719_ & _11726_ /*79138*/;
assign _11600_ = _11719_ ^ _11726_ /*79139*/;
assign _11724_ = _11725_ | _11727_ /*79136*/;
assign _11733_ = ~D[16] /*79135*/;
assign _11730_ = _11152_ & _11733_ /*79131*/;
assign _11731_ = _11152_ ^ _11733_ /*79134*/;
assign _11732_ = _11724_ & _11731_ /*79132*/;
assign _11601_ = _11724_ ^ _11731_ /*79133*/;
assign _11729_ = _11730_ | _11732_ /*79130*/;
assign _11738_ = ~D[17] /*79129*/;
assign _11735_ = _11153_ & _11738_ /*79125*/;
assign _11736_ = _11153_ ^ _11738_ /*79128*/;
assign _11737_ = _11729_ & _11736_ /*79126*/;
assign _11602_ = _11729_ ^ _11736_ /*79127*/;
assign _11734_ = _11735_ | _11737_ /*79124*/;
assign _11743_ = ~D[18] /*79123*/;
assign _11740_ = _11154_ & _11743_ /*79119*/;
assign _11741_ = _11154_ ^ _11743_ /*79122*/;
assign _11742_ = _11734_ & _11741_ /*79120*/;
assign _11603_ = _11734_ ^ _11741_ /*79121*/;
assign _11739_ = _11740_ | _11742_ /*79118*/;
assign _11748_ = ~D[19] /*79117*/;
assign _11745_ = _11155_ & _11748_ /*79113*/;
assign _11746_ = _11155_ ^ _11748_ /*79116*/;
assign _11747_ = _11739_ & _11746_ /*79114*/;
assign _11604_ = _11739_ ^ _11746_ /*79115*/;
assign _11744_ = _11745_ | _11747_ /*79112*/;
assign _11753_ = ~D[20] /*79111*/;
assign _11750_ = _11156_ & _11753_ /*79107*/;
assign _11751_ = _11156_ ^ _11753_ /*79110*/;
assign _11752_ = _11744_ & _11751_ /*79108*/;
assign _11605_ = _11744_ ^ _11751_ /*79109*/;
assign _11749_ = _11750_ | _11752_ /*79106*/;
assign _11758_ = ~D[21] /*79105*/;
assign _11755_ = _11157_ & _11758_ /*79101*/;
assign _11756_ = _11157_ ^ _11758_ /*79104*/;
assign _11757_ = _11749_ & _11756_ /*79102*/;
assign _11606_ = _11749_ ^ _11756_ /*79103*/;
assign _11754_ = _11755_ | _11757_ /*79100*/;
assign _11763_ = ~D[22] /*79099*/;
assign _11760_ = _11158_ & _11763_ /*79095*/;
assign _11761_ = _11158_ ^ _11763_ /*79098*/;
assign _11762_ = _11754_ & _11761_ /*79096*/;
assign _11607_ = _11754_ ^ _11761_ /*79097*/;
assign _11759_ = _11760_ | _11762_ /*79094*/;
assign _11768_ = ~D[23] /*79093*/;
assign _11765_ = _11159_ & _11768_ /*79089*/;
assign _11766_ = _11159_ ^ _11768_ /*79092*/;
assign _11767_ = _11759_ & _11766_ /*79090*/;
assign _11608_ = _11759_ ^ _11766_ /*79091*/;
assign _11764_ = _11765_ | _11767_ /*79088*/;
assign _11773_ = ~D[24] /*79087*/;
assign _11770_ = _11160_ & _11773_ /*79083*/;
assign _11771_ = _11160_ ^ _11773_ /*79086*/;
assign _11772_ = _11764_ & _11771_ /*79084*/;
assign _11609_ = _11764_ ^ _11771_ /*79085*/;
assign _11769_ = _11770_ | _11772_ /*79082*/;
assign _11778_ = ~D[25] /*79081*/;
assign _11775_ = _11161_ & _11778_ /*79077*/;
assign _11776_ = _11161_ ^ _11778_ /*79080*/;
assign _11777_ = _11769_ & _11776_ /*79078*/;
assign _11610_ = _11769_ ^ _11776_ /*79079*/;
assign _11774_ = _11775_ | _11777_ /*79076*/;
assign _11783_ = ~D[26] /*79075*/;
assign _11780_ = _11162_ & _11783_ /*79071*/;
assign _11781_ = _11162_ ^ _11783_ /*79074*/;
assign _11782_ = _11774_ & _11781_ /*79072*/;
assign _11611_ = _11774_ ^ _11781_ /*79073*/;
assign _11779_ = _11780_ | _11782_ /*79070*/;
assign _11788_ = ~D[27] /*79069*/;
assign _11785_ = _11163_ & _11788_ /*79065*/;
assign _11786_ = _11163_ ^ _11788_ /*79068*/;
assign _11787_ = _11779_ & _11786_ /*79066*/;
assign _11612_ = _11779_ ^ _11786_ /*79067*/;
assign _11784_ = _11785_ | _11787_ /*79064*/;
assign _11793_ = ~D[28] /*79063*/;
assign _11790_ = _11164_ & _11793_ /*79059*/;
assign _11791_ = _11164_ ^ _11793_ /*79062*/;
assign _11792_ = _11784_ & _11791_ /*79060*/;
assign _11613_ = _11784_ ^ _11791_ /*79061*/;
assign _11789_ = _11790_ | _11792_ /*79058*/;
assign _11798_ = ~D[29] /*79057*/;
assign _11795_ = _11165_ & _11798_ /*79053*/;
assign _11796_ = _11165_ ^ _11798_ /*79056*/;
assign _11797_ = _11789_ & _11796_ /*79054*/;
assign _11614_ = _11789_ ^ _11796_ /*79055*/;
assign _11794_ = _11795_ | _11797_ /*79052*/;
assign _11803_ = ~D[30] /*79051*/;
assign _11800_ = _11166_ & _11803_ /*79047*/;
assign _11801_ = _11166_ ^ _11803_ /*79050*/;
assign _11802_ = _11794_ & _11801_ /*79048*/;
assign _11615_ = _11794_ ^ _11801_ /*79049*/;
assign _11799_ = _11800_ | _11802_ /*79046*/;
assign _11808_ = ~D[31] /*79045*/;
assign _11805_ = _11167_ & _11808_ /*79041*/;
assign _11806_ = _11167_ ^ _11808_ /*79044*/;
assign _11807_ = _11799_ & _11806_ /*79042*/;
assign _11616_ = _11799_ ^ _11806_ /*79043*/;
assign _11804_ = _11805_ | _11807_ /*79040*/;
assign _11813_ = ~D[32] /*79039*/;
assign _11810_ = _11168_ & _11813_ /*79035*/;
assign _11811_ = _11168_ ^ _11813_ /*79038*/;
assign _11812_ = _11804_ & _11811_ /*79036*/;
assign _11617_ = _11804_ ^ _11811_ /*79037*/;
assign _11809_ = _11810_ | _11812_ /*79034*/;
assign _11818_ = ~D[33] /*79033*/;
assign _11815_ = _11169_ & _11818_ /*79029*/;
assign _11816_ = _11169_ ^ _11818_ /*79032*/;
assign _11817_ = _11809_ & _11816_ /*79030*/;
assign _11618_ = _11809_ ^ _11816_ /*79031*/;
assign _11814_ = _11815_ | _11817_ /*79028*/;
assign _11823_ = ~D[34] /*79027*/;
assign _11820_ = _11170_ & _11823_ /*79023*/;
assign _11821_ = _11170_ ^ _11823_ /*79026*/;
assign _11822_ = _11814_ & _11821_ /*79024*/;
assign _11619_ = _11814_ ^ _11821_ /*79025*/;
assign _11819_ = _11820_ | _11822_ /*79022*/;
assign _11828_ = ~D[35] /*79021*/;
assign _11825_ = _11171_ & _11828_ /*79017*/;
assign _11826_ = _11171_ ^ _11828_ /*79020*/;
assign _11827_ = _11819_ & _11826_ /*79018*/;
assign _11620_ = _11819_ ^ _11826_ /*79019*/;
assign _11824_ = _11825_ | _11827_ /*79016*/;
assign _11833_ = ~D[36] /*79015*/;
assign _11830_ = _11172_ & _11833_ /*79011*/;
assign _11831_ = _11172_ ^ _11833_ /*79014*/;
assign _11832_ = _11824_ & _11831_ /*79012*/;
assign _11621_ = _11824_ ^ _11831_ /*79013*/;
assign _11829_ = _11830_ | _11832_ /*79010*/;
assign _11838_ = ~D[37] /*79009*/;
assign _11835_ = _11173_ & _11838_ /*79005*/;
assign _11836_ = _11173_ ^ _11838_ /*79008*/;
assign _11837_ = _11829_ & _11836_ /*79006*/;
assign _11622_ = _11829_ ^ _11836_ /*79007*/;
assign _11834_ = _11835_ | _11837_ /*79004*/;
assign _11843_ = ~D[38] /*79003*/;
assign _11840_ = _11174_ & _11843_ /*78999*/;
assign _11841_ = _11174_ ^ _11843_ /*79002*/;
assign _11842_ = _11834_ & _11841_ /*79000*/;
assign _11623_ = _11834_ ^ _11841_ /*79001*/;
assign _11839_ = _11840_ | _11842_ /*78998*/;
assign _11848_ = ~D[39] /*78997*/;
assign _11845_ = _11175_ & _11848_ /*78993*/;
assign _11846_ = _11175_ ^ _11848_ /*78996*/;
assign _11847_ = _11839_ & _11846_ /*78994*/;
assign _11624_ = _11839_ ^ _11846_ /*78995*/;
assign _11844_ = _11845_ | _11847_ /*78992*/;
assign _11853_ = ~D[40] /*78991*/;
assign _11850_ = _11176_ & _11853_ /*78987*/;
assign _11851_ = _11176_ ^ _11853_ /*78990*/;
assign _11852_ = _11844_ & _11851_ /*78988*/;
assign _11625_ = _11844_ ^ _11851_ /*78989*/;
assign _11849_ = _11850_ | _11852_ /*78986*/;
assign _11858_ = ~D[41] /*78985*/;
assign _11855_ = _11177_ & _11858_ /*78981*/;
assign _11856_ = _11177_ ^ _11858_ /*78984*/;
assign _11857_ = _11849_ & _11856_ /*78982*/;
assign _11626_ = _11849_ ^ _11856_ /*78983*/;
assign _11854_ = _11855_ | _11857_ /*78980*/;
assign _11863_ = ~D[42] /*78979*/;
assign _11860_ = _11178_ & _11863_ /*78975*/;
assign _11861_ = _11178_ ^ _11863_ /*78978*/;
assign _11862_ = _11854_ & _11861_ /*78976*/;
assign _11627_ = _11854_ ^ _11861_ /*78977*/;
assign _11859_ = _11860_ | _11862_ /*78974*/;
assign _11868_ = ~D[43] /*78973*/;
assign _11865_ = _11179_ & _11868_ /*78969*/;
assign _11866_ = _11179_ ^ _11868_ /*78972*/;
assign _11867_ = _11859_ & _11866_ /*78970*/;
assign _11628_ = _11859_ ^ _11866_ /*78971*/;
assign _11864_ = _11865_ | _11867_ /*78968*/;
assign _11873_ = ~D[44] /*78967*/;
assign _11870_ = _11180_ & _11873_ /*78963*/;
assign _11871_ = _11180_ ^ _11873_ /*78966*/;
assign _11872_ = _11864_ & _11871_ /*78964*/;
assign _11629_ = _11864_ ^ _11871_ /*78965*/;
assign _11869_ = _11870_ | _11872_ /*78962*/;
assign _11878_ = ~D[45] /*78961*/;
assign _11875_ = _11181_ & _11878_ /*78957*/;
assign _11876_ = _11181_ ^ _11878_ /*78960*/;
assign _11877_ = _11869_ & _11876_ /*78958*/;
assign _11630_ = _11869_ ^ _11876_ /*78959*/;
assign _11874_ = _11875_ | _11877_ /*78956*/;
assign _11883_ = ~D[46] /*78955*/;
assign _11880_ = _11182_ & _11883_ /*78951*/;
assign _11881_ = _11182_ ^ _11883_ /*78954*/;
assign _11882_ = _11874_ & _11881_ /*78952*/;
assign _11631_ = _11874_ ^ _11881_ /*78953*/;
assign _11879_ = _11880_ | _11882_ /*78950*/;
assign _11888_ = ~D[47] /*78949*/;
assign _11885_ = _11183_ & _11888_ /*78945*/;
assign _11886_ = _11183_ ^ _11888_ /*78948*/;
assign _11887_ = _11879_ & _11886_ /*78946*/;
assign _11632_ = _11879_ ^ _11886_ /*78947*/;
assign _11884_ = _11885_ | _11887_ /*78944*/;
assign _11893_ = ~D[48] /*78943*/;
assign _11890_ = _11184_ & _11893_ /*78939*/;
assign _11891_ = _11184_ ^ _11893_ /*78942*/;
assign _11892_ = _11884_ & _11891_ /*78940*/;
assign _11633_ = _11884_ ^ _11891_ /*78941*/;
assign _11889_ = _11890_ | _11892_ /*78938*/;
assign _11898_ = ~D[49] /*78937*/;
assign _11895_ = _11185_ & _11898_ /*78933*/;
assign _11896_ = _11185_ ^ _11898_ /*78936*/;
assign _11897_ = _11889_ & _11896_ /*78934*/;
assign _11634_ = _11889_ ^ _11896_ /*78935*/;
assign _11894_ = _11895_ | _11897_ /*78932*/;
assign _11903_ = ~D[50] /*78931*/;
assign _11900_ = _11186_ & _11903_ /*78927*/;
assign _11901_ = _11186_ ^ _11903_ /*78930*/;
assign _11902_ = _11894_ & _11901_ /*78928*/;
assign _11635_ = _11894_ ^ _11901_ /*78929*/;
assign _11899_ = _11900_ | _11902_ /*78926*/;
assign _11908_ = ~D[51] /*78925*/;
assign _11905_ = _11187_ & _11908_ /*78921*/;
assign _11906_ = _11187_ ^ _11908_ /*78924*/;
assign _11907_ = _11899_ & _11906_ /*78922*/;
assign _11636_ = _11899_ ^ _11906_ /*78923*/;
assign _11904_ = _11905_ | _11907_ /*78920*/;
assign _11913_ = ~D[52] /*78919*/;
assign _11910_ = _11188_ & _11913_ /*78915*/;
assign _11911_ = _11188_ ^ _11913_ /*78918*/;
assign _11912_ = _11904_ & _11911_ /*78916*/;
assign _11637_ = _11904_ ^ _11911_ /*78917*/;
assign _11909_ = _11910_ | _11912_ /*78914*/;
assign _11918_ = ~D[53] /*78913*/;
assign _11915_ = _11189_ & _11918_ /*78909*/;
assign _11916_ = _11189_ ^ _11918_ /*78912*/;
assign _11917_ = _11909_ & _11916_ /*78910*/;
assign _11638_ = _11909_ ^ _11916_ /*78911*/;
assign _11914_ = _11915_ | _11917_ /*78908*/;
assign _11923_ = ~D[54] /*78907*/;
assign _11920_ = _11190_ & _11923_ /*78903*/;
assign _11921_ = _11190_ ^ _11923_ /*78906*/;
assign _11922_ = _11914_ & _11921_ /*78904*/;
assign _11639_ = _11914_ ^ _11921_ /*78905*/;
assign _11919_ = _11920_ | _11922_ /*78902*/;
assign _11928_ = ~D[55] /*78901*/;
assign _11925_ = _11191_ & _11928_ /*78897*/;
assign _11926_ = _11191_ ^ _11928_ /*78900*/;
assign _11927_ = _11919_ & _11926_ /*78898*/;
assign _11640_ = _11919_ ^ _11926_ /*78899*/;
assign _11924_ = _11925_ | _11927_ /*78896*/;
assign _11933_ = ~D[56] /*78895*/;
assign _11930_ = _11192_ & _11933_ /*78891*/;
assign _11931_ = _11192_ ^ _11933_ /*78894*/;
assign _11932_ = _11924_ & _11931_ /*78892*/;
assign _11641_ = _11924_ ^ _11931_ /*78893*/;
assign _11929_ = _11930_ | _11932_ /*78890*/;
assign _11938_ = ~D[57] /*78889*/;
assign _11935_ = _11193_ & _11938_ /*78885*/;
assign _11936_ = _11193_ ^ _11938_ /*78888*/;
assign _11937_ = _11929_ & _11936_ /*78886*/;
assign _11642_ = _11929_ ^ _11936_ /*78887*/;
assign _11934_ = _11935_ | _11937_ /*78884*/;
assign _11943_ = ~D[58] /*78883*/;
assign _11940_ = _11194_ & _11943_ /*78879*/;
assign _11941_ = _11194_ ^ _11943_ /*78882*/;
assign _11942_ = _11934_ & _11941_ /*78880*/;
assign _11643_ = _11934_ ^ _11941_ /*78881*/;
assign _11939_ = _11940_ | _11942_ /*78878*/;
assign _11948_ = ~D[59] /*78877*/;
assign _11945_ = _11195_ & _11948_ /*78873*/;
assign _11946_ = _11195_ ^ _11948_ /*78876*/;
assign _11947_ = _11939_ & _11946_ /*78874*/;
assign _11644_ = _11939_ ^ _11946_ /*78875*/;
assign _11944_ = _11945_ | _11947_ /*78872*/;
assign _11953_ = ~D[60] /*78871*/;
assign _11950_ = _11196_ & _11953_ /*78867*/;
assign _11951_ = _11196_ ^ _11953_ /*78870*/;
assign _11952_ = _11944_ & _11951_ /*78868*/;
assign _11645_ = _11944_ ^ _11951_ /*78869*/;
assign _11949_ = _11950_ | _11952_ /*78866*/;
assign _11958_ = ~D[61] /*78865*/;
assign _11955_ = _11197_ & _11958_ /*78861*/;
assign _11956_ = _11197_ ^ _11958_ /*78864*/;
assign _11957_ = _11949_ & _11956_ /*78862*/;
assign _11646_ = _11949_ ^ _11956_ /*78863*/;
assign _11954_ = _11955_ | _11957_ /*78860*/;
assign _11963_ = ~D[62] /*78859*/;
assign _11960_ = _11198_ & _11963_ /*78855*/;
assign _11961_ = _11198_ ^ _11963_ /*78858*/;
assign _11962_ = _11954_ & _11961_ /*78856*/;
assign _11647_ = _11954_ ^ _11961_ /*78857*/;
assign _11959_ = _11960_ | _11962_ /*78854*/;
assign _11964_ = _11199_ & oneWire /*78849*/;
assign _11965_ = _11199_ ^ oneWire /*78852*/;
assign _11966_ = _11959_ & _11965_ /*78850*/;
assign _11648_ = _11959_ ^ _11965_ /*78851*/;
assign Q[50] = _11964_ | _11966_ /*78848*/;
assign _12099_ = ~Q[50] /*78463*/;
assign _12098_ = _12099_ & D[0] /*78462*/;
assign _12101_ = _11585_ & _12098_ /*78457*/;
assign _12102_ = _11585_ ^ _12098_ /*78460*/;
assign _12103_ = zeroWire & _12102_ /*78458*/;
assign _12033_ = zeroWire ^ _12102_ /*78459*/;
assign _12100_ = _12101_ | _12103_ /*78456*/;
assign _12105_ = ~Q[50] /*78455*/;
assign _12104_ = _12105_ & D[1] /*78454*/;
assign _12107_ = _11586_ & _12104_ /*78449*/;
assign _12108_ = _11586_ ^ _12104_ /*78452*/;
assign _12109_ = _12100_ & _12108_ /*78450*/;
assign _12034_ = _12100_ ^ _12108_ /*78451*/;
assign _12106_ = _12107_ | _12109_ /*78448*/;
assign _12111_ = ~Q[50] /*78447*/;
assign _12110_ = _12111_ & D[2] /*78446*/;
assign _12113_ = _11587_ & _12110_ /*78441*/;
assign _12114_ = _11587_ ^ _12110_ /*78444*/;
assign _12115_ = _12106_ & _12114_ /*78442*/;
assign _12035_ = _12106_ ^ _12114_ /*78443*/;
assign _12112_ = _12113_ | _12115_ /*78440*/;
assign _12117_ = ~Q[50] /*78439*/;
assign _12116_ = _12117_ & D[3] /*78438*/;
assign _12119_ = _11588_ & _12116_ /*78433*/;
assign _12120_ = _11588_ ^ _12116_ /*78436*/;
assign _12121_ = _12112_ & _12120_ /*78434*/;
assign _12036_ = _12112_ ^ _12120_ /*78435*/;
assign _12118_ = _12119_ | _12121_ /*78432*/;
assign _12123_ = ~Q[50] /*78431*/;
assign _12122_ = _12123_ & D[4] /*78430*/;
assign _12125_ = _11589_ & _12122_ /*78425*/;
assign _12126_ = _11589_ ^ _12122_ /*78428*/;
assign _12127_ = _12118_ & _12126_ /*78426*/;
assign _12037_ = _12118_ ^ _12126_ /*78427*/;
assign _12124_ = _12125_ | _12127_ /*78424*/;
assign _12129_ = ~Q[50] /*78423*/;
assign _12128_ = _12129_ & D[5] /*78422*/;
assign _12131_ = _11590_ & _12128_ /*78417*/;
assign _12132_ = _11590_ ^ _12128_ /*78420*/;
assign _12133_ = _12124_ & _12132_ /*78418*/;
assign _12038_ = _12124_ ^ _12132_ /*78419*/;
assign _12130_ = _12131_ | _12133_ /*78416*/;
assign _12135_ = ~Q[50] /*78415*/;
assign _12134_ = _12135_ & D[6] /*78414*/;
assign _12137_ = _11591_ & _12134_ /*78409*/;
assign _12138_ = _11591_ ^ _12134_ /*78412*/;
assign _12139_ = _12130_ & _12138_ /*78410*/;
assign _12039_ = _12130_ ^ _12138_ /*78411*/;
assign _12136_ = _12137_ | _12139_ /*78408*/;
assign _12141_ = ~Q[50] /*78407*/;
assign _12140_ = _12141_ & D[7] /*78406*/;
assign _12143_ = _11592_ & _12140_ /*78401*/;
assign _12144_ = _11592_ ^ _12140_ /*78404*/;
assign _12145_ = _12136_ & _12144_ /*78402*/;
assign _12040_ = _12136_ ^ _12144_ /*78403*/;
assign _12142_ = _12143_ | _12145_ /*78400*/;
assign _12147_ = ~Q[50] /*78399*/;
assign _12146_ = _12147_ & D[8] /*78398*/;
assign _12149_ = _11593_ & _12146_ /*78393*/;
assign _12150_ = _11593_ ^ _12146_ /*78396*/;
assign _12151_ = _12142_ & _12150_ /*78394*/;
assign _12041_ = _12142_ ^ _12150_ /*78395*/;
assign _12148_ = _12149_ | _12151_ /*78392*/;
assign _12153_ = ~Q[50] /*78391*/;
assign _12152_ = _12153_ & D[9] /*78390*/;
assign _12155_ = _11594_ & _12152_ /*78385*/;
assign _12156_ = _11594_ ^ _12152_ /*78388*/;
assign _12157_ = _12148_ & _12156_ /*78386*/;
assign _12042_ = _12148_ ^ _12156_ /*78387*/;
assign _12154_ = _12155_ | _12157_ /*78384*/;
assign _12159_ = ~Q[50] /*78383*/;
assign _12158_ = _12159_ & D[10] /*78382*/;
assign _12161_ = _11595_ & _12158_ /*78377*/;
assign _12162_ = _11595_ ^ _12158_ /*78380*/;
assign _12163_ = _12154_ & _12162_ /*78378*/;
assign _12043_ = _12154_ ^ _12162_ /*78379*/;
assign _12160_ = _12161_ | _12163_ /*78376*/;
assign _12165_ = ~Q[50] /*78375*/;
assign _12164_ = _12165_ & D[11] /*78374*/;
assign _12167_ = _11596_ & _12164_ /*78369*/;
assign _12168_ = _11596_ ^ _12164_ /*78372*/;
assign _12169_ = _12160_ & _12168_ /*78370*/;
assign _12044_ = _12160_ ^ _12168_ /*78371*/;
assign _12166_ = _12167_ | _12169_ /*78368*/;
assign _12171_ = ~Q[50] /*78367*/;
assign _12170_ = _12171_ & D[12] /*78366*/;
assign _12173_ = _11597_ & _12170_ /*78361*/;
assign _12174_ = _11597_ ^ _12170_ /*78364*/;
assign _12175_ = _12166_ & _12174_ /*78362*/;
assign _12045_ = _12166_ ^ _12174_ /*78363*/;
assign _12172_ = _12173_ | _12175_ /*78360*/;
assign _12177_ = ~Q[50] /*78359*/;
assign _12176_ = _12177_ & D[13] /*78358*/;
assign _12179_ = _11598_ & _12176_ /*78353*/;
assign _12180_ = _11598_ ^ _12176_ /*78356*/;
assign _12181_ = _12172_ & _12180_ /*78354*/;
assign _12046_ = _12172_ ^ _12180_ /*78355*/;
assign _12178_ = _12179_ | _12181_ /*78352*/;
assign _12183_ = ~Q[50] /*78351*/;
assign _12182_ = _12183_ & D[14] /*78350*/;
assign _12185_ = _11599_ & _12182_ /*78345*/;
assign _12186_ = _11599_ ^ _12182_ /*78348*/;
assign _12187_ = _12178_ & _12186_ /*78346*/;
assign _12047_ = _12178_ ^ _12186_ /*78347*/;
assign _12184_ = _12185_ | _12187_ /*78344*/;
assign _12189_ = ~Q[50] /*78343*/;
assign _12188_ = _12189_ & D[15] /*78342*/;
assign _12191_ = _11600_ & _12188_ /*78337*/;
assign _12192_ = _11600_ ^ _12188_ /*78340*/;
assign _12193_ = _12184_ & _12192_ /*78338*/;
assign _12048_ = _12184_ ^ _12192_ /*78339*/;
assign _12190_ = _12191_ | _12193_ /*78336*/;
assign _12195_ = ~Q[50] /*78335*/;
assign _12194_ = _12195_ & D[16] /*78334*/;
assign _12197_ = _11601_ & _12194_ /*78329*/;
assign _12198_ = _11601_ ^ _12194_ /*78332*/;
assign _12199_ = _12190_ & _12198_ /*78330*/;
assign _12049_ = _12190_ ^ _12198_ /*78331*/;
assign _12196_ = _12197_ | _12199_ /*78328*/;
assign _12201_ = ~Q[50] /*78327*/;
assign _12200_ = _12201_ & D[17] /*78326*/;
assign _12203_ = _11602_ & _12200_ /*78321*/;
assign _12204_ = _11602_ ^ _12200_ /*78324*/;
assign _12205_ = _12196_ & _12204_ /*78322*/;
assign _12050_ = _12196_ ^ _12204_ /*78323*/;
assign _12202_ = _12203_ | _12205_ /*78320*/;
assign _12207_ = ~Q[50] /*78319*/;
assign _12206_ = _12207_ & D[18] /*78318*/;
assign _12209_ = _11603_ & _12206_ /*78313*/;
assign _12210_ = _11603_ ^ _12206_ /*78316*/;
assign _12211_ = _12202_ & _12210_ /*78314*/;
assign _12051_ = _12202_ ^ _12210_ /*78315*/;
assign _12208_ = _12209_ | _12211_ /*78312*/;
assign _12213_ = ~Q[50] /*78311*/;
assign _12212_ = _12213_ & D[19] /*78310*/;
assign _12215_ = _11604_ & _12212_ /*78305*/;
assign _12216_ = _11604_ ^ _12212_ /*78308*/;
assign _12217_ = _12208_ & _12216_ /*78306*/;
assign _12052_ = _12208_ ^ _12216_ /*78307*/;
assign _12214_ = _12215_ | _12217_ /*78304*/;
assign _12219_ = ~Q[50] /*78303*/;
assign _12218_ = _12219_ & D[20] /*78302*/;
assign _12221_ = _11605_ & _12218_ /*78297*/;
assign _12222_ = _11605_ ^ _12218_ /*78300*/;
assign _12223_ = _12214_ & _12222_ /*78298*/;
assign _12053_ = _12214_ ^ _12222_ /*78299*/;
assign _12220_ = _12221_ | _12223_ /*78296*/;
assign _12225_ = ~Q[50] /*78295*/;
assign _12224_ = _12225_ & D[21] /*78294*/;
assign _12227_ = _11606_ & _12224_ /*78289*/;
assign _12228_ = _11606_ ^ _12224_ /*78292*/;
assign _12229_ = _12220_ & _12228_ /*78290*/;
assign _12054_ = _12220_ ^ _12228_ /*78291*/;
assign _12226_ = _12227_ | _12229_ /*78288*/;
assign _12231_ = ~Q[50] /*78287*/;
assign _12230_ = _12231_ & D[22] /*78286*/;
assign _12233_ = _11607_ & _12230_ /*78281*/;
assign _12234_ = _11607_ ^ _12230_ /*78284*/;
assign _12235_ = _12226_ & _12234_ /*78282*/;
assign _12055_ = _12226_ ^ _12234_ /*78283*/;
assign _12232_ = _12233_ | _12235_ /*78280*/;
assign _12237_ = ~Q[50] /*78279*/;
assign _12236_ = _12237_ & D[23] /*78278*/;
assign _12239_ = _11608_ & _12236_ /*78273*/;
assign _12240_ = _11608_ ^ _12236_ /*78276*/;
assign _12241_ = _12232_ & _12240_ /*78274*/;
assign _12056_ = _12232_ ^ _12240_ /*78275*/;
assign _12238_ = _12239_ | _12241_ /*78272*/;
assign _12243_ = ~Q[50] /*78271*/;
assign _12242_ = _12243_ & D[24] /*78270*/;
assign _12245_ = _11609_ & _12242_ /*78265*/;
assign _12246_ = _11609_ ^ _12242_ /*78268*/;
assign _12247_ = _12238_ & _12246_ /*78266*/;
assign _12057_ = _12238_ ^ _12246_ /*78267*/;
assign _12244_ = _12245_ | _12247_ /*78264*/;
assign _12249_ = ~Q[50] /*78263*/;
assign _12248_ = _12249_ & D[25] /*78262*/;
assign _12251_ = _11610_ & _12248_ /*78257*/;
assign _12252_ = _11610_ ^ _12248_ /*78260*/;
assign _12253_ = _12244_ & _12252_ /*78258*/;
assign _12058_ = _12244_ ^ _12252_ /*78259*/;
assign _12250_ = _12251_ | _12253_ /*78256*/;
assign _12255_ = ~Q[50] /*78255*/;
assign _12254_ = _12255_ & D[26] /*78254*/;
assign _12257_ = _11611_ & _12254_ /*78249*/;
assign _12258_ = _11611_ ^ _12254_ /*78252*/;
assign _12259_ = _12250_ & _12258_ /*78250*/;
assign _12059_ = _12250_ ^ _12258_ /*78251*/;
assign _12256_ = _12257_ | _12259_ /*78248*/;
assign _12261_ = ~Q[50] /*78247*/;
assign _12260_ = _12261_ & D[27] /*78246*/;
assign _12263_ = _11612_ & _12260_ /*78241*/;
assign _12264_ = _11612_ ^ _12260_ /*78244*/;
assign _12265_ = _12256_ & _12264_ /*78242*/;
assign _12060_ = _12256_ ^ _12264_ /*78243*/;
assign _12262_ = _12263_ | _12265_ /*78240*/;
assign _12267_ = ~Q[50] /*78239*/;
assign _12266_ = _12267_ & D[28] /*78238*/;
assign _12269_ = _11613_ & _12266_ /*78233*/;
assign _12270_ = _11613_ ^ _12266_ /*78236*/;
assign _12271_ = _12262_ & _12270_ /*78234*/;
assign _12061_ = _12262_ ^ _12270_ /*78235*/;
assign _12268_ = _12269_ | _12271_ /*78232*/;
assign _12273_ = ~Q[50] /*78231*/;
assign _12272_ = _12273_ & D[29] /*78230*/;
assign _12275_ = _11614_ & _12272_ /*78225*/;
assign _12276_ = _11614_ ^ _12272_ /*78228*/;
assign _12277_ = _12268_ & _12276_ /*78226*/;
assign _12062_ = _12268_ ^ _12276_ /*78227*/;
assign _12274_ = _12275_ | _12277_ /*78224*/;
assign _12279_ = ~Q[50] /*78223*/;
assign _12278_ = _12279_ & D[30] /*78222*/;
assign _12281_ = _11615_ & _12278_ /*78217*/;
assign _12282_ = _11615_ ^ _12278_ /*78220*/;
assign _12283_ = _12274_ & _12282_ /*78218*/;
assign _12063_ = _12274_ ^ _12282_ /*78219*/;
assign _12280_ = _12281_ | _12283_ /*78216*/;
assign _12285_ = ~Q[50] /*78215*/;
assign _12284_ = _12285_ & D[31] /*78214*/;
assign _12287_ = _11616_ & _12284_ /*78209*/;
assign _12288_ = _11616_ ^ _12284_ /*78212*/;
assign _12289_ = _12280_ & _12288_ /*78210*/;
assign _12064_ = _12280_ ^ _12288_ /*78211*/;
assign _12286_ = _12287_ | _12289_ /*78208*/;
assign _12291_ = ~Q[50] /*78207*/;
assign _12290_ = _12291_ & D[32] /*78206*/;
assign _12293_ = _11617_ & _12290_ /*78201*/;
assign _12294_ = _11617_ ^ _12290_ /*78204*/;
assign _12295_ = _12286_ & _12294_ /*78202*/;
assign _12065_ = _12286_ ^ _12294_ /*78203*/;
assign _12292_ = _12293_ | _12295_ /*78200*/;
assign _12297_ = ~Q[50] /*78199*/;
assign _12296_ = _12297_ & D[33] /*78198*/;
assign _12299_ = _11618_ & _12296_ /*78193*/;
assign _12300_ = _11618_ ^ _12296_ /*78196*/;
assign _12301_ = _12292_ & _12300_ /*78194*/;
assign _12066_ = _12292_ ^ _12300_ /*78195*/;
assign _12298_ = _12299_ | _12301_ /*78192*/;
assign _12303_ = ~Q[50] /*78191*/;
assign _12302_ = _12303_ & D[34] /*78190*/;
assign _12305_ = _11619_ & _12302_ /*78185*/;
assign _12306_ = _11619_ ^ _12302_ /*78188*/;
assign _12307_ = _12298_ & _12306_ /*78186*/;
assign _12067_ = _12298_ ^ _12306_ /*78187*/;
assign _12304_ = _12305_ | _12307_ /*78184*/;
assign _12309_ = ~Q[50] /*78183*/;
assign _12308_ = _12309_ & D[35] /*78182*/;
assign _12311_ = _11620_ & _12308_ /*78177*/;
assign _12312_ = _11620_ ^ _12308_ /*78180*/;
assign _12313_ = _12304_ & _12312_ /*78178*/;
assign _12068_ = _12304_ ^ _12312_ /*78179*/;
assign _12310_ = _12311_ | _12313_ /*78176*/;
assign _12315_ = ~Q[50] /*78175*/;
assign _12314_ = _12315_ & D[36] /*78174*/;
assign _12317_ = _11621_ & _12314_ /*78169*/;
assign _12318_ = _11621_ ^ _12314_ /*78172*/;
assign _12319_ = _12310_ & _12318_ /*78170*/;
assign _12069_ = _12310_ ^ _12318_ /*78171*/;
assign _12316_ = _12317_ | _12319_ /*78168*/;
assign _12321_ = ~Q[50] /*78167*/;
assign _12320_ = _12321_ & D[37] /*78166*/;
assign _12323_ = _11622_ & _12320_ /*78161*/;
assign _12324_ = _11622_ ^ _12320_ /*78164*/;
assign _12325_ = _12316_ & _12324_ /*78162*/;
assign _12070_ = _12316_ ^ _12324_ /*78163*/;
assign _12322_ = _12323_ | _12325_ /*78160*/;
assign _12327_ = ~Q[50] /*78159*/;
assign _12326_ = _12327_ & D[38] /*78158*/;
assign _12329_ = _11623_ & _12326_ /*78153*/;
assign _12330_ = _11623_ ^ _12326_ /*78156*/;
assign _12331_ = _12322_ & _12330_ /*78154*/;
assign _12071_ = _12322_ ^ _12330_ /*78155*/;
assign _12328_ = _12329_ | _12331_ /*78152*/;
assign _12333_ = ~Q[50] /*78151*/;
assign _12332_ = _12333_ & D[39] /*78150*/;
assign _12335_ = _11624_ & _12332_ /*78145*/;
assign _12336_ = _11624_ ^ _12332_ /*78148*/;
assign _12337_ = _12328_ & _12336_ /*78146*/;
assign _12072_ = _12328_ ^ _12336_ /*78147*/;
assign _12334_ = _12335_ | _12337_ /*78144*/;
assign _12339_ = ~Q[50] /*78143*/;
assign _12338_ = _12339_ & D[40] /*78142*/;
assign _12341_ = _11625_ & _12338_ /*78137*/;
assign _12342_ = _11625_ ^ _12338_ /*78140*/;
assign _12343_ = _12334_ & _12342_ /*78138*/;
assign _12073_ = _12334_ ^ _12342_ /*78139*/;
assign _12340_ = _12341_ | _12343_ /*78136*/;
assign _12345_ = ~Q[50] /*78135*/;
assign _12344_ = _12345_ & D[41] /*78134*/;
assign _12347_ = _11626_ & _12344_ /*78129*/;
assign _12348_ = _11626_ ^ _12344_ /*78132*/;
assign _12349_ = _12340_ & _12348_ /*78130*/;
assign _12074_ = _12340_ ^ _12348_ /*78131*/;
assign _12346_ = _12347_ | _12349_ /*78128*/;
assign _12351_ = ~Q[50] /*78127*/;
assign _12350_ = _12351_ & D[42] /*78126*/;
assign _12353_ = _11627_ & _12350_ /*78121*/;
assign _12354_ = _11627_ ^ _12350_ /*78124*/;
assign _12355_ = _12346_ & _12354_ /*78122*/;
assign _12075_ = _12346_ ^ _12354_ /*78123*/;
assign _12352_ = _12353_ | _12355_ /*78120*/;
assign _12357_ = ~Q[50] /*78119*/;
assign _12356_ = _12357_ & D[43] /*78118*/;
assign _12359_ = _11628_ & _12356_ /*78113*/;
assign _12360_ = _11628_ ^ _12356_ /*78116*/;
assign _12361_ = _12352_ & _12360_ /*78114*/;
assign _12076_ = _12352_ ^ _12360_ /*78115*/;
assign _12358_ = _12359_ | _12361_ /*78112*/;
assign _12363_ = ~Q[50] /*78111*/;
assign _12362_ = _12363_ & D[44] /*78110*/;
assign _12365_ = _11629_ & _12362_ /*78105*/;
assign _12366_ = _11629_ ^ _12362_ /*78108*/;
assign _12367_ = _12358_ & _12366_ /*78106*/;
assign _12077_ = _12358_ ^ _12366_ /*78107*/;
assign _12364_ = _12365_ | _12367_ /*78104*/;
assign _12369_ = ~Q[50] /*78103*/;
assign _12368_ = _12369_ & D[45] /*78102*/;
assign _12371_ = _11630_ & _12368_ /*78097*/;
assign _12372_ = _11630_ ^ _12368_ /*78100*/;
assign _12373_ = _12364_ & _12372_ /*78098*/;
assign _12078_ = _12364_ ^ _12372_ /*78099*/;
assign _12370_ = _12371_ | _12373_ /*78096*/;
assign _12375_ = ~Q[50] /*78095*/;
assign _12374_ = _12375_ & D[46] /*78094*/;
assign _12377_ = _11631_ & _12374_ /*78089*/;
assign _12378_ = _11631_ ^ _12374_ /*78092*/;
assign _12379_ = _12370_ & _12378_ /*78090*/;
assign _12079_ = _12370_ ^ _12378_ /*78091*/;
assign _12376_ = _12377_ | _12379_ /*78088*/;
assign _12381_ = ~Q[50] /*78087*/;
assign _12380_ = _12381_ & D[47] /*78086*/;
assign _12383_ = _11632_ & _12380_ /*78081*/;
assign _12384_ = _11632_ ^ _12380_ /*78084*/;
assign _12385_ = _12376_ & _12384_ /*78082*/;
assign _12080_ = _12376_ ^ _12384_ /*78083*/;
assign _12382_ = _12383_ | _12385_ /*78080*/;
assign _12387_ = ~Q[50] /*78079*/;
assign _12386_ = _12387_ & D[48] /*78078*/;
assign _12389_ = _11633_ & _12386_ /*78073*/;
assign _12390_ = _11633_ ^ _12386_ /*78076*/;
assign _12391_ = _12382_ & _12390_ /*78074*/;
assign _12081_ = _12382_ ^ _12390_ /*78075*/;
assign _12388_ = _12389_ | _12391_ /*78072*/;
assign _12393_ = ~Q[50] /*78071*/;
assign _12392_ = _12393_ & D[49] /*78070*/;
assign _12395_ = _11634_ & _12392_ /*78065*/;
assign _12396_ = _11634_ ^ _12392_ /*78068*/;
assign _12397_ = _12388_ & _12396_ /*78066*/;
assign _12082_ = _12388_ ^ _12396_ /*78067*/;
assign _12394_ = _12395_ | _12397_ /*78064*/;
assign _12399_ = ~Q[50] /*78063*/;
assign _12398_ = _12399_ & D[50] /*78062*/;
assign _12401_ = _11635_ & _12398_ /*78057*/;
assign _12402_ = _11635_ ^ _12398_ /*78060*/;
assign _12403_ = _12394_ & _12402_ /*78058*/;
assign _12083_ = _12394_ ^ _12402_ /*78059*/;
assign _12400_ = _12401_ | _12403_ /*78056*/;
assign _12405_ = ~Q[50] /*78055*/;
assign _12404_ = _12405_ & D[51] /*78054*/;
assign _12407_ = _11636_ & _12404_ /*78049*/;
assign _12408_ = _11636_ ^ _12404_ /*78052*/;
assign _12409_ = _12400_ & _12408_ /*78050*/;
assign _12084_ = _12400_ ^ _12408_ /*78051*/;
assign _12406_ = _12407_ | _12409_ /*78048*/;
assign _12411_ = ~Q[50] /*78047*/;
assign _12410_ = _12411_ & D[52] /*78046*/;
assign _12413_ = _11637_ & _12410_ /*78041*/;
assign _12414_ = _11637_ ^ _12410_ /*78044*/;
assign _12415_ = _12406_ & _12414_ /*78042*/;
assign _12085_ = _12406_ ^ _12414_ /*78043*/;
assign _12412_ = _12413_ | _12415_ /*78040*/;
assign _12417_ = ~Q[50] /*78039*/;
assign _12416_ = _12417_ & D[53] /*78038*/;
assign _12419_ = _11638_ & _12416_ /*78033*/;
assign _12420_ = _11638_ ^ _12416_ /*78036*/;
assign _12421_ = _12412_ & _12420_ /*78034*/;
assign _12086_ = _12412_ ^ _12420_ /*78035*/;
assign _12418_ = _12419_ | _12421_ /*78032*/;
assign _12423_ = ~Q[50] /*78031*/;
assign _12422_ = _12423_ & D[54] /*78030*/;
assign _12425_ = _11639_ & _12422_ /*78025*/;
assign _12426_ = _11639_ ^ _12422_ /*78028*/;
assign _12427_ = _12418_ & _12426_ /*78026*/;
assign _12087_ = _12418_ ^ _12426_ /*78027*/;
assign _12424_ = _12425_ | _12427_ /*78024*/;
assign _12429_ = ~Q[50] /*78023*/;
assign _12428_ = _12429_ & D[55] /*78022*/;
assign _12431_ = _11640_ & _12428_ /*78017*/;
assign _12432_ = _11640_ ^ _12428_ /*78020*/;
assign _12433_ = _12424_ & _12432_ /*78018*/;
assign _12088_ = _12424_ ^ _12432_ /*78019*/;
assign _12430_ = _12431_ | _12433_ /*78016*/;
assign _12435_ = ~Q[50] /*78015*/;
assign _12434_ = _12435_ & D[56] /*78014*/;
assign _12437_ = _11641_ & _12434_ /*78009*/;
assign _12438_ = _11641_ ^ _12434_ /*78012*/;
assign _12439_ = _12430_ & _12438_ /*78010*/;
assign _12089_ = _12430_ ^ _12438_ /*78011*/;
assign _12436_ = _12437_ | _12439_ /*78008*/;
assign _12441_ = ~Q[50] /*78007*/;
assign _12440_ = _12441_ & D[57] /*78006*/;
assign _12443_ = _11642_ & _12440_ /*78001*/;
assign _12444_ = _11642_ ^ _12440_ /*78004*/;
assign _12445_ = _12436_ & _12444_ /*78002*/;
assign _12090_ = _12436_ ^ _12444_ /*78003*/;
assign _12442_ = _12443_ | _12445_ /*78000*/;
assign _12447_ = ~Q[50] /*77999*/;
assign _12446_ = _12447_ & D[58] /*77998*/;
assign _12449_ = _11643_ & _12446_ /*77993*/;
assign _12450_ = _11643_ ^ _12446_ /*77996*/;
assign _12451_ = _12442_ & _12450_ /*77994*/;
assign _12091_ = _12442_ ^ _12450_ /*77995*/;
assign _12448_ = _12449_ | _12451_ /*77992*/;
assign _12453_ = ~Q[50] /*77991*/;
assign _12452_ = _12453_ & D[59] /*77990*/;
assign _12455_ = _11644_ & _12452_ /*77985*/;
assign _12456_ = _11644_ ^ _12452_ /*77988*/;
assign _12457_ = _12448_ & _12456_ /*77986*/;
assign _12092_ = _12448_ ^ _12456_ /*77987*/;
assign _12454_ = _12455_ | _12457_ /*77984*/;
assign _12459_ = ~Q[50] /*77983*/;
assign _12458_ = _12459_ & D[60] /*77982*/;
assign _12461_ = _11645_ & _12458_ /*77977*/;
assign _12462_ = _11645_ ^ _12458_ /*77980*/;
assign _12463_ = _12454_ & _12462_ /*77978*/;
assign _12093_ = _12454_ ^ _12462_ /*77979*/;
assign _12460_ = _12461_ | _12463_ /*77976*/;
assign _12465_ = ~Q[50] /*77975*/;
assign _12464_ = _12465_ & D[61] /*77974*/;
assign _12467_ = _11646_ & _12464_ /*77969*/;
assign _12468_ = _11646_ ^ _12464_ /*77972*/;
assign _12469_ = _12460_ & _12468_ /*77970*/;
assign _12094_ = _12460_ ^ _12468_ /*77971*/;
assign _12466_ = _12467_ | _12469_ /*77968*/;
assign _12471_ = ~Q[50] /*77967*/;
assign _12470_ = _12471_ & D[62] /*77966*/;
assign _12473_ = _11647_ & _12470_ /*77961*/;
assign _12474_ = _11647_ ^ _12470_ /*77964*/;
assign _12475_ = _12466_ & _12474_ /*77962*/;
assign _12095_ = _12466_ ^ _12474_ /*77963*/;
assign _12472_ = _12473_ | _12475_ /*77960*/;
assign _12477_ = ~Q[50] /*77959*/;
assign _12476_ = _12477_ & zeroWire /*77958*/;
assign _12478_ = _11648_ ^ _12476_ /*77956*/;
assign _12096_ = _12478_ ^ _12472_ /*77955*/;
assign _12549_ = ~D[0] /*77701*/;
assign _12546_ = R_0[49] & _12549_ /*77697*/;
assign _12547_ = R_0[49] ^ _12549_ /*77700*/;
assign _12548_ = oneWire & _12547_ /*77698*/;
assign _12481_ = oneWire ^ _12547_ /*77699*/;
assign _12545_ = _12546_ | _12548_ /*77696*/;
assign _12554_ = ~D[1] /*77695*/;
assign _12551_ = _12033_ & _12554_ /*77691*/;
assign _12552_ = _12033_ ^ _12554_ /*77694*/;
assign _12553_ = _12545_ & _12552_ /*77692*/;
assign _12482_ = _12545_ ^ _12552_ /*77693*/;
assign _12550_ = _12551_ | _12553_ /*77690*/;
assign _12559_ = ~D[2] /*77689*/;
assign _12556_ = _12034_ & _12559_ /*77685*/;
assign _12557_ = _12034_ ^ _12559_ /*77688*/;
assign _12558_ = _12550_ & _12557_ /*77686*/;
assign _12483_ = _12550_ ^ _12557_ /*77687*/;
assign _12555_ = _12556_ | _12558_ /*77684*/;
assign _12564_ = ~D[3] /*77683*/;
assign _12561_ = _12035_ & _12564_ /*77679*/;
assign _12562_ = _12035_ ^ _12564_ /*77682*/;
assign _12563_ = _12555_ & _12562_ /*77680*/;
assign _12484_ = _12555_ ^ _12562_ /*77681*/;
assign _12560_ = _12561_ | _12563_ /*77678*/;
assign _12569_ = ~D[4] /*77677*/;
assign _12566_ = _12036_ & _12569_ /*77673*/;
assign _12567_ = _12036_ ^ _12569_ /*77676*/;
assign _12568_ = _12560_ & _12567_ /*77674*/;
assign _12485_ = _12560_ ^ _12567_ /*77675*/;
assign _12565_ = _12566_ | _12568_ /*77672*/;
assign _12574_ = ~D[5] /*77671*/;
assign _12571_ = _12037_ & _12574_ /*77667*/;
assign _12572_ = _12037_ ^ _12574_ /*77670*/;
assign _12573_ = _12565_ & _12572_ /*77668*/;
assign _12486_ = _12565_ ^ _12572_ /*77669*/;
assign _12570_ = _12571_ | _12573_ /*77666*/;
assign _12579_ = ~D[6] /*77665*/;
assign _12576_ = _12038_ & _12579_ /*77661*/;
assign _12577_ = _12038_ ^ _12579_ /*77664*/;
assign _12578_ = _12570_ & _12577_ /*77662*/;
assign _12487_ = _12570_ ^ _12577_ /*77663*/;
assign _12575_ = _12576_ | _12578_ /*77660*/;
assign _12584_ = ~D[7] /*77659*/;
assign _12581_ = _12039_ & _12584_ /*77655*/;
assign _12582_ = _12039_ ^ _12584_ /*77658*/;
assign _12583_ = _12575_ & _12582_ /*77656*/;
assign _12488_ = _12575_ ^ _12582_ /*77657*/;
assign _12580_ = _12581_ | _12583_ /*77654*/;
assign _12589_ = ~D[8] /*77653*/;
assign _12586_ = _12040_ & _12589_ /*77649*/;
assign _12587_ = _12040_ ^ _12589_ /*77652*/;
assign _12588_ = _12580_ & _12587_ /*77650*/;
assign _12489_ = _12580_ ^ _12587_ /*77651*/;
assign _12585_ = _12586_ | _12588_ /*77648*/;
assign _12594_ = ~D[9] /*77647*/;
assign _12591_ = _12041_ & _12594_ /*77643*/;
assign _12592_ = _12041_ ^ _12594_ /*77646*/;
assign _12593_ = _12585_ & _12592_ /*77644*/;
assign _12490_ = _12585_ ^ _12592_ /*77645*/;
assign _12590_ = _12591_ | _12593_ /*77642*/;
assign _12599_ = ~D[10] /*77641*/;
assign _12596_ = _12042_ & _12599_ /*77637*/;
assign _12597_ = _12042_ ^ _12599_ /*77640*/;
assign _12598_ = _12590_ & _12597_ /*77638*/;
assign _12491_ = _12590_ ^ _12597_ /*77639*/;
assign _12595_ = _12596_ | _12598_ /*77636*/;
assign _12604_ = ~D[11] /*77635*/;
assign _12601_ = _12043_ & _12604_ /*77631*/;
assign _12602_ = _12043_ ^ _12604_ /*77634*/;
assign _12603_ = _12595_ & _12602_ /*77632*/;
assign _12492_ = _12595_ ^ _12602_ /*77633*/;
assign _12600_ = _12601_ | _12603_ /*77630*/;
assign _12609_ = ~D[12] /*77629*/;
assign _12606_ = _12044_ & _12609_ /*77625*/;
assign _12607_ = _12044_ ^ _12609_ /*77628*/;
assign _12608_ = _12600_ & _12607_ /*77626*/;
assign _12493_ = _12600_ ^ _12607_ /*77627*/;
assign _12605_ = _12606_ | _12608_ /*77624*/;
assign _12614_ = ~D[13] /*77623*/;
assign _12611_ = _12045_ & _12614_ /*77619*/;
assign _12612_ = _12045_ ^ _12614_ /*77622*/;
assign _12613_ = _12605_ & _12612_ /*77620*/;
assign _12494_ = _12605_ ^ _12612_ /*77621*/;
assign _12610_ = _12611_ | _12613_ /*77618*/;
assign _12619_ = ~D[14] /*77617*/;
assign _12616_ = _12046_ & _12619_ /*77613*/;
assign _12617_ = _12046_ ^ _12619_ /*77616*/;
assign _12618_ = _12610_ & _12617_ /*77614*/;
assign _12495_ = _12610_ ^ _12617_ /*77615*/;
assign _12615_ = _12616_ | _12618_ /*77612*/;
assign _12624_ = ~D[15] /*77611*/;
assign _12621_ = _12047_ & _12624_ /*77607*/;
assign _12622_ = _12047_ ^ _12624_ /*77610*/;
assign _12623_ = _12615_ & _12622_ /*77608*/;
assign _12496_ = _12615_ ^ _12622_ /*77609*/;
assign _12620_ = _12621_ | _12623_ /*77606*/;
assign _12629_ = ~D[16] /*77605*/;
assign _12626_ = _12048_ & _12629_ /*77601*/;
assign _12627_ = _12048_ ^ _12629_ /*77604*/;
assign _12628_ = _12620_ & _12627_ /*77602*/;
assign _12497_ = _12620_ ^ _12627_ /*77603*/;
assign _12625_ = _12626_ | _12628_ /*77600*/;
assign _12634_ = ~D[17] /*77599*/;
assign _12631_ = _12049_ & _12634_ /*77595*/;
assign _12632_ = _12049_ ^ _12634_ /*77598*/;
assign _12633_ = _12625_ & _12632_ /*77596*/;
assign _12498_ = _12625_ ^ _12632_ /*77597*/;
assign _12630_ = _12631_ | _12633_ /*77594*/;
assign _12639_ = ~D[18] /*77593*/;
assign _12636_ = _12050_ & _12639_ /*77589*/;
assign _12637_ = _12050_ ^ _12639_ /*77592*/;
assign _12638_ = _12630_ & _12637_ /*77590*/;
assign _12499_ = _12630_ ^ _12637_ /*77591*/;
assign _12635_ = _12636_ | _12638_ /*77588*/;
assign _12644_ = ~D[19] /*77587*/;
assign _12641_ = _12051_ & _12644_ /*77583*/;
assign _12642_ = _12051_ ^ _12644_ /*77586*/;
assign _12643_ = _12635_ & _12642_ /*77584*/;
assign _12500_ = _12635_ ^ _12642_ /*77585*/;
assign _12640_ = _12641_ | _12643_ /*77582*/;
assign _12649_ = ~D[20] /*77581*/;
assign _12646_ = _12052_ & _12649_ /*77577*/;
assign _12647_ = _12052_ ^ _12649_ /*77580*/;
assign _12648_ = _12640_ & _12647_ /*77578*/;
assign _12501_ = _12640_ ^ _12647_ /*77579*/;
assign _12645_ = _12646_ | _12648_ /*77576*/;
assign _12654_ = ~D[21] /*77575*/;
assign _12651_ = _12053_ & _12654_ /*77571*/;
assign _12652_ = _12053_ ^ _12654_ /*77574*/;
assign _12653_ = _12645_ & _12652_ /*77572*/;
assign _12502_ = _12645_ ^ _12652_ /*77573*/;
assign _12650_ = _12651_ | _12653_ /*77570*/;
assign _12659_ = ~D[22] /*77569*/;
assign _12656_ = _12054_ & _12659_ /*77565*/;
assign _12657_ = _12054_ ^ _12659_ /*77568*/;
assign _12658_ = _12650_ & _12657_ /*77566*/;
assign _12503_ = _12650_ ^ _12657_ /*77567*/;
assign _12655_ = _12656_ | _12658_ /*77564*/;
assign _12664_ = ~D[23] /*77563*/;
assign _12661_ = _12055_ & _12664_ /*77559*/;
assign _12662_ = _12055_ ^ _12664_ /*77562*/;
assign _12663_ = _12655_ & _12662_ /*77560*/;
assign _12504_ = _12655_ ^ _12662_ /*77561*/;
assign _12660_ = _12661_ | _12663_ /*77558*/;
assign _12669_ = ~D[24] /*77557*/;
assign _12666_ = _12056_ & _12669_ /*77553*/;
assign _12667_ = _12056_ ^ _12669_ /*77556*/;
assign _12668_ = _12660_ & _12667_ /*77554*/;
assign _12505_ = _12660_ ^ _12667_ /*77555*/;
assign _12665_ = _12666_ | _12668_ /*77552*/;
assign _12674_ = ~D[25] /*77551*/;
assign _12671_ = _12057_ & _12674_ /*77547*/;
assign _12672_ = _12057_ ^ _12674_ /*77550*/;
assign _12673_ = _12665_ & _12672_ /*77548*/;
assign _12506_ = _12665_ ^ _12672_ /*77549*/;
assign _12670_ = _12671_ | _12673_ /*77546*/;
assign _12679_ = ~D[26] /*77545*/;
assign _12676_ = _12058_ & _12679_ /*77541*/;
assign _12677_ = _12058_ ^ _12679_ /*77544*/;
assign _12678_ = _12670_ & _12677_ /*77542*/;
assign _12507_ = _12670_ ^ _12677_ /*77543*/;
assign _12675_ = _12676_ | _12678_ /*77540*/;
assign _12684_ = ~D[27] /*77539*/;
assign _12681_ = _12059_ & _12684_ /*77535*/;
assign _12682_ = _12059_ ^ _12684_ /*77538*/;
assign _12683_ = _12675_ & _12682_ /*77536*/;
assign _12508_ = _12675_ ^ _12682_ /*77537*/;
assign _12680_ = _12681_ | _12683_ /*77534*/;
assign _12689_ = ~D[28] /*77533*/;
assign _12686_ = _12060_ & _12689_ /*77529*/;
assign _12687_ = _12060_ ^ _12689_ /*77532*/;
assign _12688_ = _12680_ & _12687_ /*77530*/;
assign _12509_ = _12680_ ^ _12687_ /*77531*/;
assign _12685_ = _12686_ | _12688_ /*77528*/;
assign _12694_ = ~D[29] /*77527*/;
assign _12691_ = _12061_ & _12694_ /*77523*/;
assign _12692_ = _12061_ ^ _12694_ /*77526*/;
assign _12693_ = _12685_ & _12692_ /*77524*/;
assign _12510_ = _12685_ ^ _12692_ /*77525*/;
assign _12690_ = _12691_ | _12693_ /*77522*/;
assign _12699_ = ~D[30] /*77521*/;
assign _12696_ = _12062_ & _12699_ /*77517*/;
assign _12697_ = _12062_ ^ _12699_ /*77520*/;
assign _12698_ = _12690_ & _12697_ /*77518*/;
assign _12511_ = _12690_ ^ _12697_ /*77519*/;
assign _12695_ = _12696_ | _12698_ /*77516*/;
assign _12704_ = ~D[31] /*77515*/;
assign _12701_ = _12063_ & _12704_ /*77511*/;
assign _12702_ = _12063_ ^ _12704_ /*77514*/;
assign _12703_ = _12695_ & _12702_ /*77512*/;
assign _12512_ = _12695_ ^ _12702_ /*77513*/;
assign _12700_ = _12701_ | _12703_ /*77510*/;
assign _12709_ = ~D[32] /*77509*/;
assign _12706_ = _12064_ & _12709_ /*77505*/;
assign _12707_ = _12064_ ^ _12709_ /*77508*/;
assign _12708_ = _12700_ & _12707_ /*77506*/;
assign _12513_ = _12700_ ^ _12707_ /*77507*/;
assign _12705_ = _12706_ | _12708_ /*77504*/;
assign _12714_ = ~D[33] /*77503*/;
assign _12711_ = _12065_ & _12714_ /*77499*/;
assign _12712_ = _12065_ ^ _12714_ /*77502*/;
assign _12713_ = _12705_ & _12712_ /*77500*/;
assign _12514_ = _12705_ ^ _12712_ /*77501*/;
assign _12710_ = _12711_ | _12713_ /*77498*/;
assign _12719_ = ~D[34] /*77497*/;
assign _12716_ = _12066_ & _12719_ /*77493*/;
assign _12717_ = _12066_ ^ _12719_ /*77496*/;
assign _12718_ = _12710_ & _12717_ /*77494*/;
assign _12515_ = _12710_ ^ _12717_ /*77495*/;
assign _12715_ = _12716_ | _12718_ /*77492*/;
assign _12724_ = ~D[35] /*77491*/;
assign _12721_ = _12067_ & _12724_ /*77487*/;
assign _12722_ = _12067_ ^ _12724_ /*77490*/;
assign _12723_ = _12715_ & _12722_ /*77488*/;
assign _12516_ = _12715_ ^ _12722_ /*77489*/;
assign _12720_ = _12721_ | _12723_ /*77486*/;
assign _12729_ = ~D[36] /*77485*/;
assign _12726_ = _12068_ & _12729_ /*77481*/;
assign _12727_ = _12068_ ^ _12729_ /*77484*/;
assign _12728_ = _12720_ & _12727_ /*77482*/;
assign _12517_ = _12720_ ^ _12727_ /*77483*/;
assign _12725_ = _12726_ | _12728_ /*77480*/;
assign _12734_ = ~D[37] /*77479*/;
assign _12731_ = _12069_ & _12734_ /*77475*/;
assign _12732_ = _12069_ ^ _12734_ /*77478*/;
assign _12733_ = _12725_ & _12732_ /*77476*/;
assign _12518_ = _12725_ ^ _12732_ /*77477*/;
assign _12730_ = _12731_ | _12733_ /*77474*/;
assign _12739_ = ~D[38] /*77473*/;
assign _12736_ = _12070_ & _12739_ /*77469*/;
assign _12737_ = _12070_ ^ _12739_ /*77472*/;
assign _12738_ = _12730_ & _12737_ /*77470*/;
assign _12519_ = _12730_ ^ _12737_ /*77471*/;
assign _12735_ = _12736_ | _12738_ /*77468*/;
assign _12744_ = ~D[39] /*77467*/;
assign _12741_ = _12071_ & _12744_ /*77463*/;
assign _12742_ = _12071_ ^ _12744_ /*77466*/;
assign _12743_ = _12735_ & _12742_ /*77464*/;
assign _12520_ = _12735_ ^ _12742_ /*77465*/;
assign _12740_ = _12741_ | _12743_ /*77462*/;
assign _12749_ = ~D[40] /*77461*/;
assign _12746_ = _12072_ & _12749_ /*77457*/;
assign _12747_ = _12072_ ^ _12749_ /*77460*/;
assign _12748_ = _12740_ & _12747_ /*77458*/;
assign _12521_ = _12740_ ^ _12747_ /*77459*/;
assign _12745_ = _12746_ | _12748_ /*77456*/;
assign _12754_ = ~D[41] /*77455*/;
assign _12751_ = _12073_ & _12754_ /*77451*/;
assign _12752_ = _12073_ ^ _12754_ /*77454*/;
assign _12753_ = _12745_ & _12752_ /*77452*/;
assign _12522_ = _12745_ ^ _12752_ /*77453*/;
assign _12750_ = _12751_ | _12753_ /*77450*/;
assign _12759_ = ~D[42] /*77449*/;
assign _12756_ = _12074_ & _12759_ /*77445*/;
assign _12757_ = _12074_ ^ _12759_ /*77448*/;
assign _12758_ = _12750_ & _12757_ /*77446*/;
assign _12523_ = _12750_ ^ _12757_ /*77447*/;
assign _12755_ = _12756_ | _12758_ /*77444*/;
assign _12764_ = ~D[43] /*77443*/;
assign _12761_ = _12075_ & _12764_ /*77439*/;
assign _12762_ = _12075_ ^ _12764_ /*77442*/;
assign _12763_ = _12755_ & _12762_ /*77440*/;
assign _12524_ = _12755_ ^ _12762_ /*77441*/;
assign _12760_ = _12761_ | _12763_ /*77438*/;
assign _12769_ = ~D[44] /*77437*/;
assign _12766_ = _12076_ & _12769_ /*77433*/;
assign _12767_ = _12076_ ^ _12769_ /*77436*/;
assign _12768_ = _12760_ & _12767_ /*77434*/;
assign _12525_ = _12760_ ^ _12767_ /*77435*/;
assign _12765_ = _12766_ | _12768_ /*77432*/;
assign _12774_ = ~D[45] /*77431*/;
assign _12771_ = _12077_ & _12774_ /*77427*/;
assign _12772_ = _12077_ ^ _12774_ /*77430*/;
assign _12773_ = _12765_ & _12772_ /*77428*/;
assign _12526_ = _12765_ ^ _12772_ /*77429*/;
assign _12770_ = _12771_ | _12773_ /*77426*/;
assign _12779_ = ~D[46] /*77425*/;
assign _12776_ = _12078_ & _12779_ /*77421*/;
assign _12777_ = _12078_ ^ _12779_ /*77424*/;
assign _12778_ = _12770_ & _12777_ /*77422*/;
assign _12527_ = _12770_ ^ _12777_ /*77423*/;
assign _12775_ = _12776_ | _12778_ /*77420*/;
assign _12784_ = ~D[47] /*77419*/;
assign _12781_ = _12079_ & _12784_ /*77415*/;
assign _12782_ = _12079_ ^ _12784_ /*77418*/;
assign _12783_ = _12775_ & _12782_ /*77416*/;
assign _12528_ = _12775_ ^ _12782_ /*77417*/;
assign _12780_ = _12781_ | _12783_ /*77414*/;
assign _12789_ = ~D[48] /*77413*/;
assign _12786_ = _12080_ & _12789_ /*77409*/;
assign _12787_ = _12080_ ^ _12789_ /*77412*/;
assign _12788_ = _12780_ & _12787_ /*77410*/;
assign _12529_ = _12780_ ^ _12787_ /*77411*/;
assign _12785_ = _12786_ | _12788_ /*77408*/;
assign _12794_ = ~D[49] /*77407*/;
assign _12791_ = _12081_ & _12794_ /*77403*/;
assign _12792_ = _12081_ ^ _12794_ /*77406*/;
assign _12793_ = _12785_ & _12792_ /*77404*/;
assign _12530_ = _12785_ ^ _12792_ /*77405*/;
assign _12790_ = _12791_ | _12793_ /*77402*/;
assign _12799_ = ~D[50] /*77401*/;
assign _12796_ = _12082_ & _12799_ /*77397*/;
assign _12797_ = _12082_ ^ _12799_ /*77400*/;
assign _12798_ = _12790_ & _12797_ /*77398*/;
assign _12531_ = _12790_ ^ _12797_ /*77399*/;
assign _12795_ = _12796_ | _12798_ /*77396*/;
assign _12804_ = ~D[51] /*77395*/;
assign _12801_ = _12083_ & _12804_ /*77391*/;
assign _12802_ = _12083_ ^ _12804_ /*77394*/;
assign _12803_ = _12795_ & _12802_ /*77392*/;
assign _12532_ = _12795_ ^ _12802_ /*77393*/;
assign _12800_ = _12801_ | _12803_ /*77390*/;
assign _12809_ = ~D[52] /*77389*/;
assign _12806_ = _12084_ & _12809_ /*77385*/;
assign _12807_ = _12084_ ^ _12809_ /*77388*/;
assign _12808_ = _12800_ & _12807_ /*77386*/;
assign _12533_ = _12800_ ^ _12807_ /*77387*/;
assign _12805_ = _12806_ | _12808_ /*77384*/;
assign _12814_ = ~D[53] /*77383*/;
assign _12811_ = _12085_ & _12814_ /*77379*/;
assign _12812_ = _12085_ ^ _12814_ /*77382*/;
assign _12813_ = _12805_ & _12812_ /*77380*/;
assign _12534_ = _12805_ ^ _12812_ /*77381*/;
assign _12810_ = _12811_ | _12813_ /*77378*/;
assign _12819_ = ~D[54] /*77377*/;
assign _12816_ = _12086_ & _12819_ /*77373*/;
assign _12817_ = _12086_ ^ _12819_ /*77376*/;
assign _12818_ = _12810_ & _12817_ /*77374*/;
assign _12535_ = _12810_ ^ _12817_ /*77375*/;
assign _12815_ = _12816_ | _12818_ /*77372*/;
assign _12824_ = ~D[55] /*77371*/;
assign _12821_ = _12087_ & _12824_ /*77367*/;
assign _12822_ = _12087_ ^ _12824_ /*77370*/;
assign _12823_ = _12815_ & _12822_ /*77368*/;
assign _12536_ = _12815_ ^ _12822_ /*77369*/;
assign _12820_ = _12821_ | _12823_ /*77366*/;
assign _12829_ = ~D[56] /*77365*/;
assign _12826_ = _12088_ & _12829_ /*77361*/;
assign _12827_ = _12088_ ^ _12829_ /*77364*/;
assign _12828_ = _12820_ & _12827_ /*77362*/;
assign _12537_ = _12820_ ^ _12827_ /*77363*/;
assign _12825_ = _12826_ | _12828_ /*77360*/;
assign _12834_ = ~D[57] /*77359*/;
assign _12831_ = _12089_ & _12834_ /*77355*/;
assign _12832_ = _12089_ ^ _12834_ /*77358*/;
assign _12833_ = _12825_ & _12832_ /*77356*/;
assign _12538_ = _12825_ ^ _12832_ /*77357*/;
assign _12830_ = _12831_ | _12833_ /*77354*/;
assign _12839_ = ~D[58] /*77353*/;
assign _12836_ = _12090_ & _12839_ /*77349*/;
assign _12837_ = _12090_ ^ _12839_ /*77352*/;
assign _12838_ = _12830_ & _12837_ /*77350*/;
assign _12539_ = _12830_ ^ _12837_ /*77351*/;
assign _12835_ = _12836_ | _12838_ /*77348*/;
assign _12844_ = ~D[59] /*77347*/;
assign _12841_ = _12091_ & _12844_ /*77343*/;
assign _12842_ = _12091_ ^ _12844_ /*77346*/;
assign _12843_ = _12835_ & _12842_ /*77344*/;
assign _12540_ = _12835_ ^ _12842_ /*77345*/;
assign _12840_ = _12841_ | _12843_ /*77342*/;
assign _12849_ = ~D[60] /*77341*/;
assign _12846_ = _12092_ & _12849_ /*77337*/;
assign _12847_ = _12092_ ^ _12849_ /*77340*/;
assign _12848_ = _12840_ & _12847_ /*77338*/;
assign _12541_ = _12840_ ^ _12847_ /*77339*/;
assign _12845_ = _12846_ | _12848_ /*77336*/;
assign _12854_ = ~D[61] /*77335*/;
assign _12851_ = _12093_ & _12854_ /*77331*/;
assign _12852_ = _12093_ ^ _12854_ /*77334*/;
assign _12853_ = _12845_ & _12852_ /*77332*/;
assign _12542_ = _12845_ ^ _12852_ /*77333*/;
assign _12850_ = _12851_ | _12853_ /*77330*/;
assign _12859_ = ~D[62] /*77329*/;
assign _12856_ = _12094_ & _12859_ /*77325*/;
assign _12857_ = _12094_ ^ _12859_ /*77328*/;
assign _12858_ = _12850_ & _12857_ /*77326*/;
assign _12543_ = _12850_ ^ _12857_ /*77327*/;
assign _12855_ = _12856_ | _12858_ /*77324*/;
assign _12860_ = _12095_ & oneWire /*77319*/;
assign _12861_ = _12095_ ^ oneWire /*77322*/;
assign _12862_ = _12855_ & _12861_ /*77320*/;
assign _12544_ = _12855_ ^ _12861_ /*77321*/;
assign Q[49] = _12860_ | _12862_ /*77318*/;
assign _12995_ = ~Q[49] /*76933*/;
assign _12994_ = _12995_ & D[0] /*76932*/;
assign _12997_ = _12481_ & _12994_ /*76927*/;
assign _12998_ = _12481_ ^ _12994_ /*76930*/;
assign _12999_ = zeroWire & _12998_ /*76928*/;
assign _12929_ = zeroWire ^ _12998_ /*76929*/;
assign _12996_ = _12997_ | _12999_ /*76926*/;
assign _13001_ = ~Q[49] /*76925*/;
assign _13000_ = _13001_ & D[1] /*76924*/;
assign _13003_ = _12482_ & _13000_ /*76919*/;
assign _13004_ = _12482_ ^ _13000_ /*76922*/;
assign _13005_ = _12996_ & _13004_ /*76920*/;
assign _12930_ = _12996_ ^ _13004_ /*76921*/;
assign _13002_ = _13003_ | _13005_ /*76918*/;
assign _13007_ = ~Q[49] /*76917*/;
assign _13006_ = _13007_ & D[2] /*76916*/;
assign _13009_ = _12483_ & _13006_ /*76911*/;
assign _13010_ = _12483_ ^ _13006_ /*76914*/;
assign _13011_ = _13002_ & _13010_ /*76912*/;
assign _12931_ = _13002_ ^ _13010_ /*76913*/;
assign _13008_ = _13009_ | _13011_ /*76910*/;
assign _13013_ = ~Q[49] /*76909*/;
assign _13012_ = _13013_ & D[3] /*76908*/;
assign _13015_ = _12484_ & _13012_ /*76903*/;
assign _13016_ = _12484_ ^ _13012_ /*76906*/;
assign _13017_ = _13008_ & _13016_ /*76904*/;
assign _12932_ = _13008_ ^ _13016_ /*76905*/;
assign _13014_ = _13015_ | _13017_ /*76902*/;
assign _13019_ = ~Q[49] /*76901*/;
assign _13018_ = _13019_ & D[4] /*76900*/;
assign _13021_ = _12485_ & _13018_ /*76895*/;
assign _13022_ = _12485_ ^ _13018_ /*76898*/;
assign _13023_ = _13014_ & _13022_ /*76896*/;
assign _12933_ = _13014_ ^ _13022_ /*76897*/;
assign _13020_ = _13021_ | _13023_ /*76894*/;
assign _13025_ = ~Q[49] /*76893*/;
assign _13024_ = _13025_ & D[5] /*76892*/;
assign _13027_ = _12486_ & _13024_ /*76887*/;
assign _13028_ = _12486_ ^ _13024_ /*76890*/;
assign _13029_ = _13020_ & _13028_ /*76888*/;
assign _12934_ = _13020_ ^ _13028_ /*76889*/;
assign _13026_ = _13027_ | _13029_ /*76886*/;
assign _13031_ = ~Q[49] /*76885*/;
assign _13030_ = _13031_ & D[6] /*76884*/;
assign _13033_ = _12487_ & _13030_ /*76879*/;
assign _13034_ = _12487_ ^ _13030_ /*76882*/;
assign _13035_ = _13026_ & _13034_ /*76880*/;
assign _12935_ = _13026_ ^ _13034_ /*76881*/;
assign _13032_ = _13033_ | _13035_ /*76878*/;
assign _13037_ = ~Q[49] /*76877*/;
assign _13036_ = _13037_ & D[7] /*76876*/;
assign _13039_ = _12488_ & _13036_ /*76871*/;
assign _13040_ = _12488_ ^ _13036_ /*76874*/;
assign _13041_ = _13032_ & _13040_ /*76872*/;
assign _12936_ = _13032_ ^ _13040_ /*76873*/;
assign _13038_ = _13039_ | _13041_ /*76870*/;
assign _13043_ = ~Q[49] /*76869*/;
assign _13042_ = _13043_ & D[8] /*76868*/;
assign _13045_ = _12489_ & _13042_ /*76863*/;
assign _13046_ = _12489_ ^ _13042_ /*76866*/;
assign _13047_ = _13038_ & _13046_ /*76864*/;
assign _12937_ = _13038_ ^ _13046_ /*76865*/;
assign _13044_ = _13045_ | _13047_ /*76862*/;
assign _13049_ = ~Q[49] /*76861*/;
assign _13048_ = _13049_ & D[9] /*76860*/;
assign _13051_ = _12490_ & _13048_ /*76855*/;
assign _13052_ = _12490_ ^ _13048_ /*76858*/;
assign _13053_ = _13044_ & _13052_ /*76856*/;
assign _12938_ = _13044_ ^ _13052_ /*76857*/;
assign _13050_ = _13051_ | _13053_ /*76854*/;
assign _13055_ = ~Q[49] /*76853*/;
assign _13054_ = _13055_ & D[10] /*76852*/;
assign _13057_ = _12491_ & _13054_ /*76847*/;
assign _13058_ = _12491_ ^ _13054_ /*76850*/;
assign _13059_ = _13050_ & _13058_ /*76848*/;
assign _12939_ = _13050_ ^ _13058_ /*76849*/;
assign _13056_ = _13057_ | _13059_ /*76846*/;
assign _13061_ = ~Q[49] /*76845*/;
assign _13060_ = _13061_ & D[11] /*76844*/;
assign _13063_ = _12492_ & _13060_ /*76839*/;
assign _13064_ = _12492_ ^ _13060_ /*76842*/;
assign _13065_ = _13056_ & _13064_ /*76840*/;
assign _12940_ = _13056_ ^ _13064_ /*76841*/;
assign _13062_ = _13063_ | _13065_ /*76838*/;
assign _13067_ = ~Q[49] /*76837*/;
assign _13066_ = _13067_ & D[12] /*76836*/;
assign _13069_ = _12493_ & _13066_ /*76831*/;
assign _13070_ = _12493_ ^ _13066_ /*76834*/;
assign _13071_ = _13062_ & _13070_ /*76832*/;
assign _12941_ = _13062_ ^ _13070_ /*76833*/;
assign _13068_ = _13069_ | _13071_ /*76830*/;
assign _13073_ = ~Q[49] /*76829*/;
assign _13072_ = _13073_ & D[13] /*76828*/;
assign _13075_ = _12494_ & _13072_ /*76823*/;
assign _13076_ = _12494_ ^ _13072_ /*76826*/;
assign _13077_ = _13068_ & _13076_ /*76824*/;
assign _12942_ = _13068_ ^ _13076_ /*76825*/;
assign _13074_ = _13075_ | _13077_ /*76822*/;
assign _13079_ = ~Q[49] /*76821*/;
assign _13078_ = _13079_ & D[14] /*76820*/;
assign _13081_ = _12495_ & _13078_ /*76815*/;
assign _13082_ = _12495_ ^ _13078_ /*76818*/;
assign _13083_ = _13074_ & _13082_ /*76816*/;
assign _12943_ = _13074_ ^ _13082_ /*76817*/;
assign _13080_ = _13081_ | _13083_ /*76814*/;
assign _13085_ = ~Q[49] /*76813*/;
assign _13084_ = _13085_ & D[15] /*76812*/;
assign _13087_ = _12496_ & _13084_ /*76807*/;
assign _13088_ = _12496_ ^ _13084_ /*76810*/;
assign _13089_ = _13080_ & _13088_ /*76808*/;
assign _12944_ = _13080_ ^ _13088_ /*76809*/;
assign _13086_ = _13087_ | _13089_ /*76806*/;
assign _13091_ = ~Q[49] /*76805*/;
assign _13090_ = _13091_ & D[16] /*76804*/;
assign _13093_ = _12497_ & _13090_ /*76799*/;
assign _13094_ = _12497_ ^ _13090_ /*76802*/;
assign _13095_ = _13086_ & _13094_ /*76800*/;
assign _12945_ = _13086_ ^ _13094_ /*76801*/;
assign _13092_ = _13093_ | _13095_ /*76798*/;
assign _13097_ = ~Q[49] /*76797*/;
assign _13096_ = _13097_ & D[17] /*76796*/;
assign _13099_ = _12498_ & _13096_ /*76791*/;
assign _13100_ = _12498_ ^ _13096_ /*76794*/;
assign _13101_ = _13092_ & _13100_ /*76792*/;
assign _12946_ = _13092_ ^ _13100_ /*76793*/;
assign _13098_ = _13099_ | _13101_ /*76790*/;
assign _13103_ = ~Q[49] /*76789*/;
assign _13102_ = _13103_ & D[18] /*76788*/;
assign _13105_ = _12499_ & _13102_ /*76783*/;
assign _13106_ = _12499_ ^ _13102_ /*76786*/;
assign _13107_ = _13098_ & _13106_ /*76784*/;
assign _12947_ = _13098_ ^ _13106_ /*76785*/;
assign _13104_ = _13105_ | _13107_ /*76782*/;
assign _13109_ = ~Q[49] /*76781*/;
assign _13108_ = _13109_ & D[19] /*76780*/;
assign _13111_ = _12500_ & _13108_ /*76775*/;
assign _13112_ = _12500_ ^ _13108_ /*76778*/;
assign _13113_ = _13104_ & _13112_ /*76776*/;
assign _12948_ = _13104_ ^ _13112_ /*76777*/;
assign _13110_ = _13111_ | _13113_ /*76774*/;
assign _13115_ = ~Q[49] /*76773*/;
assign _13114_ = _13115_ & D[20] /*76772*/;
assign _13117_ = _12501_ & _13114_ /*76767*/;
assign _13118_ = _12501_ ^ _13114_ /*76770*/;
assign _13119_ = _13110_ & _13118_ /*76768*/;
assign _12949_ = _13110_ ^ _13118_ /*76769*/;
assign _13116_ = _13117_ | _13119_ /*76766*/;
assign _13121_ = ~Q[49] /*76765*/;
assign _13120_ = _13121_ & D[21] /*76764*/;
assign _13123_ = _12502_ & _13120_ /*76759*/;
assign _13124_ = _12502_ ^ _13120_ /*76762*/;
assign _13125_ = _13116_ & _13124_ /*76760*/;
assign _12950_ = _13116_ ^ _13124_ /*76761*/;
assign _13122_ = _13123_ | _13125_ /*76758*/;
assign _13127_ = ~Q[49] /*76757*/;
assign _13126_ = _13127_ & D[22] /*76756*/;
assign _13129_ = _12503_ & _13126_ /*76751*/;
assign _13130_ = _12503_ ^ _13126_ /*76754*/;
assign _13131_ = _13122_ & _13130_ /*76752*/;
assign _12951_ = _13122_ ^ _13130_ /*76753*/;
assign _13128_ = _13129_ | _13131_ /*76750*/;
assign _13133_ = ~Q[49] /*76749*/;
assign _13132_ = _13133_ & D[23] /*76748*/;
assign _13135_ = _12504_ & _13132_ /*76743*/;
assign _13136_ = _12504_ ^ _13132_ /*76746*/;
assign _13137_ = _13128_ & _13136_ /*76744*/;
assign _12952_ = _13128_ ^ _13136_ /*76745*/;
assign _13134_ = _13135_ | _13137_ /*76742*/;
assign _13139_ = ~Q[49] /*76741*/;
assign _13138_ = _13139_ & D[24] /*76740*/;
assign _13141_ = _12505_ & _13138_ /*76735*/;
assign _13142_ = _12505_ ^ _13138_ /*76738*/;
assign _13143_ = _13134_ & _13142_ /*76736*/;
assign _12953_ = _13134_ ^ _13142_ /*76737*/;
assign _13140_ = _13141_ | _13143_ /*76734*/;
assign _13145_ = ~Q[49] /*76733*/;
assign _13144_ = _13145_ & D[25] /*76732*/;
assign _13147_ = _12506_ & _13144_ /*76727*/;
assign _13148_ = _12506_ ^ _13144_ /*76730*/;
assign _13149_ = _13140_ & _13148_ /*76728*/;
assign _12954_ = _13140_ ^ _13148_ /*76729*/;
assign _13146_ = _13147_ | _13149_ /*76726*/;
assign _13151_ = ~Q[49] /*76725*/;
assign _13150_ = _13151_ & D[26] /*76724*/;
assign _13153_ = _12507_ & _13150_ /*76719*/;
assign _13154_ = _12507_ ^ _13150_ /*76722*/;
assign _13155_ = _13146_ & _13154_ /*76720*/;
assign _12955_ = _13146_ ^ _13154_ /*76721*/;
assign _13152_ = _13153_ | _13155_ /*76718*/;
assign _13157_ = ~Q[49] /*76717*/;
assign _13156_ = _13157_ & D[27] /*76716*/;
assign _13159_ = _12508_ & _13156_ /*76711*/;
assign _13160_ = _12508_ ^ _13156_ /*76714*/;
assign _13161_ = _13152_ & _13160_ /*76712*/;
assign _12956_ = _13152_ ^ _13160_ /*76713*/;
assign _13158_ = _13159_ | _13161_ /*76710*/;
assign _13163_ = ~Q[49] /*76709*/;
assign _13162_ = _13163_ & D[28] /*76708*/;
assign _13165_ = _12509_ & _13162_ /*76703*/;
assign _13166_ = _12509_ ^ _13162_ /*76706*/;
assign _13167_ = _13158_ & _13166_ /*76704*/;
assign _12957_ = _13158_ ^ _13166_ /*76705*/;
assign _13164_ = _13165_ | _13167_ /*76702*/;
assign _13169_ = ~Q[49] /*76701*/;
assign _13168_ = _13169_ & D[29] /*76700*/;
assign _13171_ = _12510_ & _13168_ /*76695*/;
assign _13172_ = _12510_ ^ _13168_ /*76698*/;
assign _13173_ = _13164_ & _13172_ /*76696*/;
assign _12958_ = _13164_ ^ _13172_ /*76697*/;
assign _13170_ = _13171_ | _13173_ /*76694*/;
assign _13175_ = ~Q[49] /*76693*/;
assign _13174_ = _13175_ & D[30] /*76692*/;
assign _13177_ = _12511_ & _13174_ /*76687*/;
assign _13178_ = _12511_ ^ _13174_ /*76690*/;
assign _13179_ = _13170_ & _13178_ /*76688*/;
assign _12959_ = _13170_ ^ _13178_ /*76689*/;
assign _13176_ = _13177_ | _13179_ /*76686*/;
assign _13181_ = ~Q[49] /*76685*/;
assign _13180_ = _13181_ & D[31] /*76684*/;
assign _13183_ = _12512_ & _13180_ /*76679*/;
assign _13184_ = _12512_ ^ _13180_ /*76682*/;
assign _13185_ = _13176_ & _13184_ /*76680*/;
assign _12960_ = _13176_ ^ _13184_ /*76681*/;
assign _13182_ = _13183_ | _13185_ /*76678*/;
assign _13187_ = ~Q[49] /*76677*/;
assign _13186_ = _13187_ & D[32] /*76676*/;
assign _13189_ = _12513_ & _13186_ /*76671*/;
assign _13190_ = _12513_ ^ _13186_ /*76674*/;
assign _13191_ = _13182_ & _13190_ /*76672*/;
assign _12961_ = _13182_ ^ _13190_ /*76673*/;
assign _13188_ = _13189_ | _13191_ /*76670*/;
assign _13193_ = ~Q[49] /*76669*/;
assign _13192_ = _13193_ & D[33] /*76668*/;
assign _13195_ = _12514_ & _13192_ /*76663*/;
assign _13196_ = _12514_ ^ _13192_ /*76666*/;
assign _13197_ = _13188_ & _13196_ /*76664*/;
assign _12962_ = _13188_ ^ _13196_ /*76665*/;
assign _13194_ = _13195_ | _13197_ /*76662*/;
assign _13199_ = ~Q[49] /*76661*/;
assign _13198_ = _13199_ & D[34] /*76660*/;
assign _13201_ = _12515_ & _13198_ /*76655*/;
assign _13202_ = _12515_ ^ _13198_ /*76658*/;
assign _13203_ = _13194_ & _13202_ /*76656*/;
assign _12963_ = _13194_ ^ _13202_ /*76657*/;
assign _13200_ = _13201_ | _13203_ /*76654*/;
assign _13205_ = ~Q[49] /*76653*/;
assign _13204_ = _13205_ & D[35] /*76652*/;
assign _13207_ = _12516_ & _13204_ /*76647*/;
assign _13208_ = _12516_ ^ _13204_ /*76650*/;
assign _13209_ = _13200_ & _13208_ /*76648*/;
assign _12964_ = _13200_ ^ _13208_ /*76649*/;
assign _13206_ = _13207_ | _13209_ /*76646*/;
assign _13211_ = ~Q[49] /*76645*/;
assign _13210_ = _13211_ & D[36] /*76644*/;
assign _13213_ = _12517_ & _13210_ /*76639*/;
assign _13214_ = _12517_ ^ _13210_ /*76642*/;
assign _13215_ = _13206_ & _13214_ /*76640*/;
assign _12965_ = _13206_ ^ _13214_ /*76641*/;
assign _13212_ = _13213_ | _13215_ /*76638*/;
assign _13217_ = ~Q[49] /*76637*/;
assign _13216_ = _13217_ & D[37] /*76636*/;
assign _13219_ = _12518_ & _13216_ /*76631*/;
assign _13220_ = _12518_ ^ _13216_ /*76634*/;
assign _13221_ = _13212_ & _13220_ /*76632*/;
assign _12966_ = _13212_ ^ _13220_ /*76633*/;
assign _13218_ = _13219_ | _13221_ /*76630*/;
assign _13223_ = ~Q[49] /*76629*/;
assign _13222_ = _13223_ & D[38] /*76628*/;
assign _13225_ = _12519_ & _13222_ /*76623*/;
assign _13226_ = _12519_ ^ _13222_ /*76626*/;
assign _13227_ = _13218_ & _13226_ /*76624*/;
assign _12967_ = _13218_ ^ _13226_ /*76625*/;
assign _13224_ = _13225_ | _13227_ /*76622*/;
assign _13229_ = ~Q[49] /*76621*/;
assign _13228_ = _13229_ & D[39] /*76620*/;
assign _13231_ = _12520_ & _13228_ /*76615*/;
assign _13232_ = _12520_ ^ _13228_ /*76618*/;
assign _13233_ = _13224_ & _13232_ /*76616*/;
assign _12968_ = _13224_ ^ _13232_ /*76617*/;
assign _13230_ = _13231_ | _13233_ /*76614*/;
assign _13235_ = ~Q[49] /*76613*/;
assign _13234_ = _13235_ & D[40] /*76612*/;
assign _13237_ = _12521_ & _13234_ /*76607*/;
assign _13238_ = _12521_ ^ _13234_ /*76610*/;
assign _13239_ = _13230_ & _13238_ /*76608*/;
assign _12969_ = _13230_ ^ _13238_ /*76609*/;
assign _13236_ = _13237_ | _13239_ /*76606*/;
assign _13241_ = ~Q[49] /*76605*/;
assign _13240_ = _13241_ & D[41] /*76604*/;
assign _13243_ = _12522_ & _13240_ /*76599*/;
assign _13244_ = _12522_ ^ _13240_ /*76602*/;
assign _13245_ = _13236_ & _13244_ /*76600*/;
assign _12970_ = _13236_ ^ _13244_ /*76601*/;
assign _13242_ = _13243_ | _13245_ /*76598*/;
assign _13247_ = ~Q[49] /*76597*/;
assign _13246_ = _13247_ & D[42] /*76596*/;
assign _13249_ = _12523_ & _13246_ /*76591*/;
assign _13250_ = _12523_ ^ _13246_ /*76594*/;
assign _13251_ = _13242_ & _13250_ /*76592*/;
assign _12971_ = _13242_ ^ _13250_ /*76593*/;
assign _13248_ = _13249_ | _13251_ /*76590*/;
assign _13253_ = ~Q[49] /*76589*/;
assign _13252_ = _13253_ & D[43] /*76588*/;
assign _13255_ = _12524_ & _13252_ /*76583*/;
assign _13256_ = _12524_ ^ _13252_ /*76586*/;
assign _13257_ = _13248_ & _13256_ /*76584*/;
assign _12972_ = _13248_ ^ _13256_ /*76585*/;
assign _13254_ = _13255_ | _13257_ /*76582*/;
assign _13259_ = ~Q[49] /*76581*/;
assign _13258_ = _13259_ & D[44] /*76580*/;
assign _13261_ = _12525_ & _13258_ /*76575*/;
assign _13262_ = _12525_ ^ _13258_ /*76578*/;
assign _13263_ = _13254_ & _13262_ /*76576*/;
assign _12973_ = _13254_ ^ _13262_ /*76577*/;
assign _13260_ = _13261_ | _13263_ /*76574*/;
assign _13265_ = ~Q[49] /*76573*/;
assign _13264_ = _13265_ & D[45] /*76572*/;
assign _13267_ = _12526_ & _13264_ /*76567*/;
assign _13268_ = _12526_ ^ _13264_ /*76570*/;
assign _13269_ = _13260_ & _13268_ /*76568*/;
assign _12974_ = _13260_ ^ _13268_ /*76569*/;
assign _13266_ = _13267_ | _13269_ /*76566*/;
assign _13271_ = ~Q[49] /*76565*/;
assign _13270_ = _13271_ & D[46] /*76564*/;
assign _13273_ = _12527_ & _13270_ /*76559*/;
assign _13274_ = _12527_ ^ _13270_ /*76562*/;
assign _13275_ = _13266_ & _13274_ /*76560*/;
assign _12975_ = _13266_ ^ _13274_ /*76561*/;
assign _13272_ = _13273_ | _13275_ /*76558*/;
assign _13277_ = ~Q[49] /*76557*/;
assign _13276_ = _13277_ & D[47] /*76556*/;
assign _13279_ = _12528_ & _13276_ /*76551*/;
assign _13280_ = _12528_ ^ _13276_ /*76554*/;
assign _13281_ = _13272_ & _13280_ /*76552*/;
assign _12976_ = _13272_ ^ _13280_ /*76553*/;
assign _13278_ = _13279_ | _13281_ /*76550*/;
assign _13283_ = ~Q[49] /*76549*/;
assign _13282_ = _13283_ & D[48] /*76548*/;
assign _13285_ = _12529_ & _13282_ /*76543*/;
assign _13286_ = _12529_ ^ _13282_ /*76546*/;
assign _13287_ = _13278_ & _13286_ /*76544*/;
assign _12977_ = _13278_ ^ _13286_ /*76545*/;
assign _13284_ = _13285_ | _13287_ /*76542*/;
assign _13289_ = ~Q[49] /*76541*/;
assign _13288_ = _13289_ & D[49] /*76540*/;
assign _13291_ = _12530_ & _13288_ /*76535*/;
assign _13292_ = _12530_ ^ _13288_ /*76538*/;
assign _13293_ = _13284_ & _13292_ /*76536*/;
assign _12978_ = _13284_ ^ _13292_ /*76537*/;
assign _13290_ = _13291_ | _13293_ /*76534*/;
assign _13295_ = ~Q[49] /*76533*/;
assign _13294_ = _13295_ & D[50] /*76532*/;
assign _13297_ = _12531_ & _13294_ /*76527*/;
assign _13298_ = _12531_ ^ _13294_ /*76530*/;
assign _13299_ = _13290_ & _13298_ /*76528*/;
assign _12979_ = _13290_ ^ _13298_ /*76529*/;
assign _13296_ = _13297_ | _13299_ /*76526*/;
assign _13301_ = ~Q[49] /*76525*/;
assign _13300_ = _13301_ & D[51] /*76524*/;
assign _13303_ = _12532_ & _13300_ /*76519*/;
assign _13304_ = _12532_ ^ _13300_ /*76522*/;
assign _13305_ = _13296_ & _13304_ /*76520*/;
assign _12980_ = _13296_ ^ _13304_ /*76521*/;
assign _13302_ = _13303_ | _13305_ /*76518*/;
assign _13307_ = ~Q[49] /*76517*/;
assign _13306_ = _13307_ & D[52] /*76516*/;
assign _13309_ = _12533_ & _13306_ /*76511*/;
assign _13310_ = _12533_ ^ _13306_ /*76514*/;
assign _13311_ = _13302_ & _13310_ /*76512*/;
assign _12981_ = _13302_ ^ _13310_ /*76513*/;
assign _13308_ = _13309_ | _13311_ /*76510*/;
assign _13313_ = ~Q[49] /*76509*/;
assign _13312_ = _13313_ & D[53] /*76508*/;
assign _13315_ = _12534_ & _13312_ /*76503*/;
assign _13316_ = _12534_ ^ _13312_ /*76506*/;
assign _13317_ = _13308_ & _13316_ /*76504*/;
assign _12982_ = _13308_ ^ _13316_ /*76505*/;
assign _13314_ = _13315_ | _13317_ /*76502*/;
assign _13319_ = ~Q[49] /*76501*/;
assign _13318_ = _13319_ & D[54] /*76500*/;
assign _13321_ = _12535_ & _13318_ /*76495*/;
assign _13322_ = _12535_ ^ _13318_ /*76498*/;
assign _13323_ = _13314_ & _13322_ /*76496*/;
assign _12983_ = _13314_ ^ _13322_ /*76497*/;
assign _13320_ = _13321_ | _13323_ /*76494*/;
assign _13325_ = ~Q[49] /*76493*/;
assign _13324_ = _13325_ & D[55] /*76492*/;
assign _13327_ = _12536_ & _13324_ /*76487*/;
assign _13328_ = _12536_ ^ _13324_ /*76490*/;
assign _13329_ = _13320_ & _13328_ /*76488*/;
assign _12984_ = _13320_ ^ _13328_ /*76489*/;
assign _13326_ = _13327_ | _13329_ /*76486*/;
assign _13331_ = ~Q[49] /*76485*/;
assign _13330_ = _13331_ & D[56] /*76484*/;
assign _13333_ = _12537_ & _13330_ /*76479*/;
assign _13334_ = _12537_ ^ _13330_ /*76482*/;
assign _13335_ = _13326_ & _13334_ /*76480*/;
assign _12985_ = _13326_ ^ _13334_ /*76481*/;
assign _13332_ = _13333_ | _13335_ /*76478*/;
assign _13337_ = ~Q[49] /*76477*/;
assign _13336_ = _13337_ & D[57] /*76476*/;
assign _13339_ = _12538_ & _13336_ /*76471*/;
assign _13340_ = _12538_ ^ _13336_ /*76474*/;
assign _13341_ = _13332_ & _13340_ /*76472*/;
assign _12986_ = _13332_ ^ _13340_ /*76473*/;
assign _13338_ = _13339_ | _13341_ /*76470*/;
assign _13343_ = ~Q[49] /*76469*/;
assign _13342_ = _13343_ & D[58] /*76468*/;
assign _13345_ = _12539_ & _13342_ /*76463*/;
assign _13346_ = _12539_ ^ _13342_ /*76466*/;
assign _13347_ = _13338_ & _13346_ /*76464*/;
assign _12987_ = _13338_ ^ _13346_ /*76465*/;
assign _13344_ = _13345_ | _13347_ /*76462*/;
assign _13349_ = ~Q[49] /*76461*/;
assign _13348_ = _13349_ & D[59] /*76460*/;
assign _13351_ = _12540_ & _13348_ /*76455*/;
assign _13352_ = _12540_ ^ _13348_ /*76458*/;
assign _13353_ = _13344_ & _13352_ /*76456*/;
assign _12988_ = _13344_ ^ _13352_ /*76457*/;
assign _13350_ = _13351_ | _13353_ /*76454*/;
assign _13355_ = ~Q[49] /*76453*/;
assign _13354_ = _13355_ & D[60] /*76452*/;
assign _13357_ = _12541_ & _13354_ /*76447*/;
assign _13358_ = _12541_ ^ _13354_ /*76450*/;
assign _13359_ = _13350_ & _13358_ /*76448*/;
assign _12989_ = _13350_ ^ _13358_ /*76449*/;
assign _13356_ = _13357_ | _13359_ /*76446*/;
assign _13361_ = ~Q[49] /*76445*/;
assign _13360_ = _13361_ & D[61] /*76444*/;
assign _13363_ = _12542_ & _13360_ /*76439*/;
assign _13364_ = _12542_ ^ _13360_ /*76442*/;
assign _13365_ = _13356_ & _13364_ /*76440*/;
assign _12990_ = _13356_ ^ _13364_ /*76441*/;
assign _13362_ = _13363_ | _13365_ /*76438*/;
assign _13367_ = ~Q[49] /*76437*/;
assign _13366_ = _13367_ & D[62] /*76436*/;
assign _13369_ = _12543_ & _13366_ /*76431*/;
assign _13370_ = _12543_ ^ _13366_ /*76434*/;
assign _13371_ = _13362_ & _13370_ /*76432*/;
assign _12991_ = _13362_ ^ _13370_ /*76433*/;
assign _13368_ = _13369_ | _13371_ /*76430*/;
assign _13373_ = ~Q[49] /*76429*/;
assign _13372_ = _13373_ & zeroWire /*76428*/;
assign _13374_ = _12544_ ^ _13372_ /*76426*/;
assign _12992_ = _13374_ ^ _13368_ /*76425*/;
assign _13445_ = ~D[0] /*76171*/;
assign _13442_ = R_0[48] & _13445_ /*76167*/;
assign _13443_ = R_0[48] ^ _13445_ /*76170*/;
assign _13444_ = oneWire & _13443_ /*76168*/;
assign _13377_ = oneWire ^ _13443_ /*76169*/;
assign _13441_ = _13442_ | _13444_ /*76166*/;
assign _13450_ = ~D[1] /*76165*/;
assign _13447_ = _12929_ & _13450_ /*76161*/;
assign _13448_ = _12929_ ^ _13450_ /*76164*/;
assign _13449_ = _13441_ & _13448_ /*76162*/;
assign _13378_ = _13441_ ^ _13448_ /*76163*/;
assign _13446_ = _13447_ | _13449_ /*76160*/;
assign _13455_ = ~D[2] /*76159*/;
assign _13452_ = _12930_ & _13455_ /*76155*/;
assign _13453_ = _12930_ ^ _13455_ /*76158*/;
assign _13454_ = _13446_ & _13453_ /*76156*/;
assign _13379_ = _13446_ ^ _13453_ /*76157*/;
assign _13451_ = _13452_ | _13454_ /*76154*/;
assign _13460_ = ~D[3] /*76153*/;
assign _13457_ = _12931_ & _13460_ /*76149*/;
assign _13458_ = _12931_ ^ _13460_ /*76152*/;
assign _13459_ = _13451_ & _13458_ /*76150*/;
assign _13380_ = _13451_ ^ _13458_ /*76151*/;
assign _13456_ = _13457_ | _13459_ /*76148*/;
assign _13465_ = ~D[4] /*76147*/;
assign _13462_ = _12932_ & _13465_ /*76143*/;
assign _13463_ = _12932_ ^ _13465_ /*76146*/;
assign _13464_ = _13456_ & _13463_ /*76144*/;
assign _13381_ = _13456_ ^ _13463_ /*76145*/;
assign _13461_ = _13462_ | _13464_ /*76142*/;
assign _13470_ = ~D[5] /*76141*/;
assign _13467_ = _12933_ & _13470_ /*76137*/;
assign _13468_ = _12933_ ^ _13470_ /*76140*/;
assign _13469_ = _13461_ & _13468_ /*76138*/;
assign _13382_ = _13461_ ^ _13468_ /*76139*/;
assign _13466_ = _13467_ | _13469_ /*76136*/;
assign _13475_ = ~D[6] /*76135*/;
assign _13472_ = _12934_ & _13475_ /*76131*/;
assign _13473_ = _12934_ ^ _13475_ /*76134*/;
assign _13474_ = _13466_ & _13473_ /*76132*/;
assign _13383_ = _13466_ ^ _13473_ /*76133*/;
assign _13471_ = _13472_ | _13474_ /*76130*/;
assign _13480_ = ~D[7] /*76129*/;
assign _13477_ = _12935_ & _13480_ /*76125*/;
assign _13478_ = _12935_ ^ _13480_ /*76128*/;
assign _13479_ = _13471_ & _13478_ /*76126*/;
assign _13384_ = _13471_ ^ _13478_ /*76127*/;
assign _13476_ = _13477_ | _13479_ /*76124*/;
assign _13485_ = ~D[8] /*76123*/;
assign _13482_ = _12936_ & _13485_ /*76119*/;
assign _13483_ = _12936_ ^ _13485_ /*76122*/;
assign _13484_ = _13476_ & _13483_ /*76120*/;
assign _13385_ = _13476_ ^ _13483_ /*76121*/;
assign _13481_ = _13482_ | _13484_ /*76118*/;
assign _13490_ = ~D[9] /*76117*/;
assign _13487_ = _12937_ & _13490_ /*76113*/;
assign _13488_ = _12937_ ^ _13490_ /*76116*/;
assign _13489_ = _13481_ & _13488_ /*76114*/;
assign _13386_ = _13481_ ^ _13488_ /*76115*/;
assign _13486_ = _13487_ | _13489_ /*76112*/;
assign _13495_ = ~D[10] /*76111*/;
assign _13492_ = _12938_ & _13495_ /*76107*/;
assign _13493_ = _12938_ ^ _13495_ /*76110*/;
assign _13494_ = _13486_ & _13493_ /*76108*/;
assign _13387_ = _13486_ ^ _13493_ /*76109*/;
assign _13491_ = _13492_ | _13494_ /*76106*/;
assign _13500_ = ~D[11] /*76105*/;
assign _13497_ = _12939_ & _13500_ /*76101*/;
assign _13498_ = _12939_ ^ _13500_ /*76104*/;
assign _13499_ = _13491_ & _13498_ /*76102*/;
assign _13388_ = _13491_ ^ _13498_ /*76103*/;
assign _13496_ = _13497_ | _13499_ /*76100*/;
assign _13505_ = ~D[12] /*76099*/;
assign _13502_ = _12940_ & _13505_ /*76095*/;
assign _13503_ = _12940_ ^ _13505_ /*76098*/;
assign _13504_ = _13496_ & _13503_ /*76096*/;
assign _13389_ = _13496_ ^ _13503_ /*76097*/;
assign _13501_ = _13502_ | _13504_ /*76094*/;
assign _13510_ = ~D[13] /*76093*/;
assign _13507_ = _12941_ & _13510_ /*76089*/;
assign _13508_ = _12941_ ^ _13510_ /*76092*/;
assign _13509_ = _13501_ & _13508_ /*76090*/;
assign _13390_ = _13501_ ^ _13508_ /*76091*/;
assign _13506_ = _13507_ | _13509_ /*76088*/;
assign _13515_ = ~D[14] /*76087*/;
assign _13512_ = _12942_ & _13515_ /*76083*/;
assign _13513_ = _12942_ ^ _13515_ /*76086*/;
assign _13514_ = _13506_ & _13513_ /*76084*/;
assign _13391_ = _13506_ ^ _13513_ /*76085*/;
assign _13511_ = _13512_ | _13514_ /*76082*/;
assign _13520_ = ~D[15] /*76081*/;
assign _13517_ = _12943_ & _13520_ /*76077*/;
assign _13518_ = _12943_ ^ _13520_ /*76080*/;
assign _13519_ = _13511_ & _13518_ /*76078*/;
assign _13392_ = _13511_ ^ _13518_ /*76079*/;
assign _13516_ = _13517_ | _13519_ /*76076*/;
assign _13525_ = ~D[16] /*76075*/;
assign _13522_ = _12944_ & _13525_ /*76071*/;
assign _13523_ = _12944_ ^ _13525_ /*76074*/;
assign _13524_ = _13516_ & _13523_ /*76072*/;
assign _13393_ = _13516_ ^ _13523_ /*76073*/;
assign _13521_ = _13522_ | _13524_ /*76070*/;
assign _13530_ = ~D[17] /*76069*/;
assign _13527_ = _12945_ & _13530_ /*76065*/;
assign _13528_ = _12945_ ^ _13530_ /*76068*/;
assign _13529_ = _13521_ & _13528_ /*76066*/;
assign _13394_ = _13521_ ^ _13528_ /*76067*/;
assign _13526_ = _13527_ | _13529_ /*76064*/;
assign _13535_ = ~D[18] /*76063*/;
assign _13532_ = _12946_ & _13535_ /*76059*/;
assign _13533_ = _12946_ ^ _13535_ /*76062*/;
assign _13534_ = _13526_ & _13533_ /*76060*/;
assign _13395_ = _13526_ ^ _13533_ /*76061*/;
assign _13531_ = _13532_ | _13534_ /*76058*/;
assign _13540_ = ~D[19] /*76057*/;
assign _13537_ = _12947_ & _13540_ /*76053*/;
assign _13538_ = _12947_ ^ _13540_ /*76056*/;
assign _13539_ = _13531_ & _13538_ /*76054*/;
assign _13396_ = _13531_ ^ _13538_ /*76055*/;
assign _13536_ = _13537_ | _13539_ /*76052*/;
assign _13545_ = ~D[20] /*76051*/;
assign _13542_ = _12948_ & _13545_ /*76047*/;
assign _13543_ = _12948_ ^ _13545_ /*76050*/;
assign _13544_ = _13536_ & _13543_ /*76048*/;
assign _13397_ = _13536_ ^ _13543_ /*76049*/;
assign _13541_ = _13542_ | _13544_ /*76046*/;
assign _13550_ = ~D[21] /*76045*/;
assign _13547_ = _12949_ & _13550_ /*76041*/;
assign _13548_ = _12949_ ^ _13550_ /*76044*/;
assign _13549_ = _13541_ & _13548_ /*76042*/;
assign _13398_ = _13541_ ^ _13548_ /*76043*/;
assign _13546_ = _13547_ | _13549_ /*76040*/;
assign _13555_ = ~D[22] /*76039*/;
assign _13552_ = _12950_ & _13555_ /*76035*/;
assign _13553_ = _12950_ ^ _13555_ /*76038*/;
assign _13554_ = _13546_ & _13553_ /*76036*/;
assign _13399_ = _13546_ ^ _13553_ /*76037*/;
assign _13551_ = _13552_ | _13554_ /*76034*/;
assign _13560_ = ~D[23] /*76033*/;
assign _13557_ = _12951_ & _13560_ /*76029*/;
assign _13558_ = _12951_ ^ _13560_ /*76032*/;
assign _13559_ = _13551_ & _13558_ /*76030*/;
assign _13400_ = _13551_ ^ _13558_ /*76031*/;
assign _13556_ = _13557_ | _13559_ /*76028*/;
assign _13565_ = ~D[24] /*76027*/;
assign _13562_ = _12952_ & _13565_ /*76023*/;
assign _13563_ = _12952_ ^ _13565_ /*76026*/;
assign _13564_ = _13556_ & _13563_ /*76024*/;
assign _13401_ = _13556_ ^ _13563_ /*76025*/;
assign _13561_ = _13562_ | _13564_ /*76022*/;
assign _13570_ = ~D[25] /*76021*/;
assign _13567_ = _12953_ & _13570_ /*76017*/;
assign _13568_ = _12953_ ^ _13570_ /*76020*/;
assign _13569_ = _13561_ & _13568_ /*76018*/;
assign _13402_ = _13561_ ^ _13568_ /*76019*/;
assign _13566_ = _13567_ | _13569_ /*76016*/;
assign _13575_ = ~D[26] /*76015*/;
assign _13572_ = _12954_ & _13575_ /*76011*/;
assign _13573_ = _12954_ ^ _13575_ /*76014*/;
assign _13574_ = _13566_ & _13573_ /*76012*/;
assign _13403_ = _13566_ ^ _13573_ /*76013*/;
assign _13571_ = _13572_ | _13574_ /*76010*/;
assign _13580_ = ~D[27] /*76009*/;
assign _13577_ = _12955_ & _13580_ /*76005*/;
assign _13578_ = _12955_ ^ _13580_ /*76008*/;
assign _13579_ = _13571_ & _13578_ /*76006*/;
assign _13404_ = _13571_ ^ _13578_ /*76007*/;
assign _13576_ = _13577_ | _13579_ /*76004*/;
assign _13585_ = ~D[28] /*76003*/;
assign _13582_ = _12956_ & _13585_ /*75999*/;
assign _13583_ = _12956_ ^ _13585_ /*76002*/;
assign _13584_ = _13576_ & _13583_ /*76000*/;
assign _13405_ = _13576_ ^ _13583_ /*76001*/;
assign _13581_ = _13582_ | _13584_ /*75998*/;
assign _13590_ = ~D[29] /*75997*/;
assign _13587_ = _12957_ & _13590_ /*75993*/;
assign _13588_ = _12957_ ^ _13590_ /*75996*/;
assign _13589_ = _13581_ & _13588_ /*75994*/;
assign _13406_ = _13581_ ^ _13588_ /*75995*/;
assign _13586_ = _13587_ | _13589_ /*75992*/;
assign _13595_ = ~D[30] /*75991*/;
assign _13592_ = _12958_ & _13595_ /*75987*/;
assign _13593_ = _12958_ ^ _13595_ /*75990*/;
assign _13594_ = _13586_ & _13593_ /*75988*/;
assign _13407_ = _13586_ ^ _13593_ /*75989*/;
assign _13591_ = _13592_ | _13594_ /*75986*/;
assign _13600_ = ~D[31] /*75985*/;
assign _13597_ = _12959_ & _13600_ /*75981*/;
assign _13598_ = _12959_ ^ _13600_ /*75984*/;
assign _13599_ = _13591_ & _13598_ /*75982*/;
assign _13408_ = _13591_ ^ _13598_ /*75983*/;
assign _13596_ = _13597_ | _13599_ /*75980*/;
assign _13605_ = ~D[32] /*75979*/;
assign _13602_ = _12960_ & _13605_ /*75975*/;
assign _13603_ = _12960_ ^ _13605_ /*75978*/;
assign _13604_ = _13596_ & _13603_ /*75976*/;
assign _13409_ = _13596_ ^ _13603_ /*75977*/;
assign _13601_ = _13602_ | _13604_ /*75974*/;
assign _13610_ = ~D[33] /*75973*/;
assign _13607_ = _12961_ & _13610_ /*75969*/;
assign _13608_ = _12961_ ^ _13610_ /*75972*/;
assign _13609_ = _13601_ & _13608_ /*75970*/;
assign _13410_ = _13601_ ^ _13608_ /*75971*/;
assign _13606_ = _13607_ | _13609_ /*75968*/;
assign _13615_ = ~D[34] /*75967*/;
assign _13612_ = _12962_ & _13615_ /*75963*/;
assign _13613_ = _12962_ ^ _13615_ /*75966*/;
assign _13614_ = _13606_ & _13613_ /*75964*/;
assign _13411_ = _13606_ ^ _13613_ /*75965*/;
assign _13611_ = _13612_ | _13614_ /*75962*/;
assign _13620_ = ~D[35] /*75961*/;
assign _13617_ = _12963_ & _13620_ /*75957*/;
assign _13618_ = _12963_ ^ _13620_ /*75960*/;
assign _13619_ = _13611_ & _13618_ /*75958*/;
assign _13412_ = _13611_ ^ _13618_ /*75959*/;
assign _13616_ = _13617_ | _13619_ /*75956*/;
assign _13625_ = ~D[36] /*75955*/;
assign _13622_ = _12964_ & _13625_ /*75951*/;
assign _13623_ = _12964_ ^ _13625_ /*75954*/;
assign _13624_ = _13616_ & _13623_ /*75952*/;
assign _13413_ = _13616_ ^ _13623_ /*75953*/;
assign _13621_ = _13622_ | _13624_ /*75950*/;
assign _13630_ = ~D[37] /*75949*/;
assign _13627_ = _12965_ & _13630_ /*75945*/;
assign _13628_ = _12965_ ^ _13630_ /*75948*/;
assign _13629_ = _13621_ & _13628_ /*75946*/;
assign _13414_ = _13621_ ^ _13628_ /*75947*/;
assign _13626_ = _13627_ | _13629_ /*75944*/;
assign _13635_ = ~D[38] /*75943*/;
assign _13632_ = _12966_ & _13635_ /*75939*/;
assign _13633_ = _12966_ ^ _13635_ /*75942*/;
assign _13634_ = _13626_ & _13633_ /*75940*/;
assign _13415_ = _13626_ ^ _13633_ /*75941*/;
assign _13631_ = _13632_ | _13634_ /*75938*/;
assign _13640_ = ~D[39] /*75937*/;
assign _13637_ = _12967_ & _13640_ /*75933*/;
assign _13638_ = _12967_ ^ _13640_ /*75936*/;
assign _13639_ = _13631_ & _13638_ /*75934*/;
assign _13416_ = _13631_ ^ _13638_ /*75935*/;
assign _13636_ = _13637_ | _13639_ /*75932*/;
assign _13645_ = ~D[40] /*75931*/;
assign _13642_ = _12968_ & _13645_ /*75927*/;
assign _13643_ = _12968_ ^ _13645_ /*75930*/;
assign _13644_ = _13636_ & _13643_ /*75928*/;
assign _13417_ = _13636_ ^ _13643_ /*75929*/;
assign _13641_ = _13642_ | _13644_ /*75926*/;
assign _13650_ = ~D[41] /*75925*/;
assign _13647_ = _12969_ & _13650_ /*75921*/;
assign _13648_ = _12969_ ^ _13650_ /*75924*/;
assign _13649_ = _13641_ & _13648_ /*75922*/;
assign _13418_ = _13641_ ^ _13648_ /*75923*/;
assign _13646_ = _13647_ | _13649_ /*75920*/;
assign _13655_ = ~D[42] /*75919*/;
assign _13652_ = _12970_ & _13655_ /*75915*/;
assign _13653_ = _12970_ ^ _13655_ /*75918*/;
assign _13654_ = _13646_ & _13653_ /*75916*/;
assign _13419_ = _13646_ ^ _13653_ /*75917*/;
assign _13651_ = _13652_ | _13654_ /*75914*/;
assign _13660_ = ~D[43] /*75913*/;
assign _13657_ = _12971_ & _13660_ /*75909*/;
assign _13658_ = _12971_ ^ _13660_ /*75912*/;
assign _13659_ = _13651_ & _13658_ /*75910*/;
assign _13420_ = _13651_ ^ _13658_ /*75911*/;
assign _13656_ = _13657_ | _13659_ /*75908*/;
assign _13665_ = ~D[44] /*75907*/;
assign _13662_ = _12972_ & _13665_ /*75903*/;
assign _13663_ = _12972_ ^ _13665_ /*75906*/;
assign _13664_ = _13656_ & _13663_ /*75904*/;
assign _13421_ = _13656_ ^ _13663_ /*75905*/;
assign _13661_ = _13662_ | _13664_ /*75902*/;
assign _13670_ = ~D[45] /*75901*/;
assign _13667_ = _12973_ & _13670_ /*75897*/;
assign _13668_ = _12973_ ^ _13670_ /*75900*/;
assign _13669_ = _13661_ & _13668_ /*75898*/;
assign _13422_ = _13661_ ^ _13668_ /*75899*/;
assign _13666_ = _13667_ | _13669_ /*75896*/;
assign _13675_ = ~D[46] /*75895*/;
assign _13672_ = _12974_ & _13675_ /*75891*/;
assign _13673_ = _12974_ ^ _13675_ /*75894*/;
assign _13674_ = _13666_ & _13673_ /*75892*/;
assign _13423_ = _13666_ ^ _13673_ /*75893*/;
assign _13671_ = _13672_ | _13674_ /*75890*/;
assign _13680_ = ~D[47] /*75889*/;
assign _13677_ = _12975_ & _13680_ /*75885*/;
assign _13678_ = _12975_ ^ _13680_ /*75888*/;
assign _13679_ = _13671_ & _13678_ /*75886*/;
assign _13424_ = _13671_ ^ _13678_ /*75887*/;
assign _13676_ = _13677_ | _13679_ /*75884*/;
assign _13685_ = ~D[48] /*75883*/;
assign _13682_ = _12976_ & _13685_ /*75879*/;
assign _13683_ = _12976_ ^ _13685_ /*75882*/;
assign _13684_ = _13676_ & _13683_ /*75880*/;
assign _13425_ = _13676_ ^ _13683_ /*75881*/;
assign _13681_ = _13682_ | _13684_ /*75878*/;
assign _13690_ = ~D[49] /*75877*/;
assign _13687_ = _12977_ & _13690_ /*75873*/;
assign _13688_ = _12977_ ^ _13690_ /*75876*/;
assign _13689_ = _13681_ & _13688_ /*75874*/;
assign _13426_ = _13681_ ^ _13688_ /*75875*/;
assign _13686_ = _13687_ | _13689_ /*75872*/;
assign _13695_ = ~D[50] /*75871*/;
assign _13692_ = _12978_ & _13695_ /*75867*/;
assign _13693_ = _12978_ ^ _13695_ /*75870*/;
assign _13694_ = _13686_ & _13693_ /*75868*/;
assign _13427_ = _13686_ ^ _13693_ /*75869*/;
assign _13691_ = _13692_ | _13694_ /*75866*/;
assign _13700_ = ~D[51] /*75865*/;
assign _13697_ = _12979_ & _13700_ /*75861*/;
assign _13698_ = _12979_ ^ _13700_ /*75864*/;
assign _13699_ = _13691_ & _13698_ /*75862*/;
assign _13428_ = _13691_ ^ _13698_ /*75863*/;
assign _13696_ = _13697_ | _13699_ /*75860*/;
assign _13705_ = ~D[52] /*75859*/;
assign _13702_ = _12980_ & _13705_ /*75855*/;
assign _13703_ = _12980_ ^ _13705_ /*75858*/;
assign _13704_ = _13696_ & _13703_ /*75856*/;
assign _13429_ = _13696_ ^ _13703_ /*75857*/;
assign _13701_ = _13702_ | _13704_ /*75854*/;
assign _13710_ = ~D[53] /*75853*/;
assign _13707_ = _12981_ & _13710_ /*75849*/;
assign _13708_ = _12981_ ^ _13710_ /*75852*/;
assign _13709_ = _13701_ & _13708_ /*75850*/;
assign _13430_ = _13701_ ^ _13708_ /*75851*/;
assign _13706_ = _13707_ | _13709_ /*75848*/;
assign _13715_ = ~D[54] /*75847*/;
assign _13712_ = _12982_ & _13715_ /*75843*/;
assign _13713_ = _12982_ ^ _13715_ /*75846*/;
assign _13714_ = _13706_ & _13713_ /*75844*/;
assign _13431_ = _13706_ ^ _13713_ /*75845*/;
assign _13711_ = _13712_ | _13714_ /*75842*/;
assign _13720_ = ~D[55] /*75841*/;
assign _13717_ = _12983_ & _13720_ /*75837*/;
assign _13718_ = _12983_ ^ _13720_ /*75840*/;
assign _13719_ = _13711_ & _13718_ /*75838*/;
assign _13432_ = _13711_ ^ _13718_ /*75839*/;
assign _13716_ = _13717_ | _13719_ /*75836*/;
assign _13725_ = ~D[56] /*75835*/;
assign _13722_ = _12984_ & _13725_ /*75831*/;
assign _13723_ = _12984_ ^ _13725_ /*75834*/;
assign _13724_ = _13716_ & _13723_ /*75832*/;
assign _13433_ = _13716_ ^ _13723_ /*75833*/;
assign _13721_ = _13722_ | _13724_ /*75830*/;
assign _13730_ = ~D[57] /*75829*/;
assign _13727_ = _12985_ & _13730_ /*75825*/;
assign _13728_ = _12985_ ^ _13730_ /*75828*/;
assign _13729_ = _13721_ & _13728_ /*75826*/;
assign _13434_ = _13721_ ^ _13728_ /*75827*/;
assign _13726_ = _13727_ | _13729_ /*75824*/;
assign _13735_ = ~D[58] /*75823*/;
assign _13732_ = _12986_ & _13735_ /*75819*/;
assign _13733_ = _12986_ ^ _13735_ /*75822*/;
assign _13734_ = _13726_ & _13733_ /*75820*/;
assign _13435_ = _13726_ ^ _13733_ /*75821*/;
assign _13731_ = _13732_ | _13734_ /*75818*/;
assign _13740_ = ~D[59] /*75817*/;
assign _13737_ = _12987_ & _13740_ /*75813*/;
assign _13738_ = _12987_ ^ _13740_ /*75816*/;
assign _13739_ = _13731_ & _13738_ /*75814*/;
assign _13436_ = _13731_ ^ _13738_ /*75815*/;
assign _13736_ = _13737_ | _13739_ /*75812*/;
assign _13745_ = ~D[60] /*75811*/;
assign _13742_ = _12988_ & _13745_ /*75807*/;
assign _13743_ = _12988_ ^ _13745_ /*75810*/;
assign _13744_ = _13736_ & _13743_ /*75808*/;
assign _13437_ = _13736_ ^ _13743_ /*75809*/;
assign _13741_ = _13742_ | _13744_ /*75806*/;
assign _13750_ = ~D[61] /*75805*/;
assign _13747_ = _12989_ & _13750_ /*75801*/;
assign _13748_ = _12989_ ^ _13750_ /*75804*/;
assign _13749_ = _13741_ & _13748_ /*75802*/;
assign _13438_ = _13741_ ^ _13748_ /*75803*/;
assign _13746_ = _13747_ | _13749_ /*75800*/;
assign _13755_ = ~D[62] /*75799*/;
assign _13752_ = _12990_ & _13755_ /*75795*/;
assign _13753_ = _12990_ ^ _13755_ /*75798*/;
assign _13754_ = _13746_ & _13753_ /*75796*/;
assign _13439_ = _13746_ ^ _13753_ /*75797*/;
assign _13751_ = _13752_ | _13754_ /*75794*/;
assign _13756_ = _12991_ & oneWire /*75789*/;
assign _13757_ = _12991_ ^ oneWire /*75792*/;
assign _13758_ = _13751_ & _13757_ /*75790*/;
assign _13440_ = _13751_ ^ _13757_ /*75791*/;
assign Q[48] = _13756_ | _13758_ /*75788*/;
assign _13891_ = ~Q[48] /*75403*/;
assign _13890_ = _13891_ & D[0] /*75402*/;
assign _13893_ = _13377_ & _13890_ /*75397*/;
assign _13894_ = _13377_ ^ _13890_ /*75400*/;
assign _13895_ = zeroWire & _13894_ /*75398*/;
assign _13825_ = zeroWire ^ _13894_ /*75399*/;
assign _13892_ = _13893_ | _13895_ /*75396*/;
assign _13897_ = ~Q[48] /*75395*/;
assign _13896_ = _13897_ & D[1] /*75394*/;
assign _13899_ = _13378_ & _13896_ /*75389*/;
assign _13900_ = _13378_ ^ _13896_ /*75392*/;
assign _13901_ = _13892_ & _13900_ /*75390*/;
assign _13826_ = _13892_ ^ _13900_ /*75391*/;
assign _13898_ = _13899_ | _13901_ /*75388*/;
assign _13903_ = ~Q[48] /*75387*/;
assign _13902_ = _13903_ & D[2] /*75386*/;
assign _13905_ = _13379_ & _13902_ /*75381*/;
assign _13906_ = _13379_ ^ _13902_ /*75384*/;
assign _13907_ = _13898_ & _13906_ /*75382*/;
assign _13827_ = _13898_ ^ _13906_ /*75383*/;
assign _13904_ = _13905_ | _13907_ /*75380*/;
assign _13909_ = ~Q[48] /*75379*/;
assign _13908_ = _13909_ & D[3] /*75378*/;
assign _13911_ = _13380_ & _13908_ /*75373*/;
assign _13912_ = _13380_ ^ _13908_ /*75376*/;
assign _13913_ = _13904_ & _13912_ /*75374*/;
assign _13828_ = _13904_ ^ _13912_ /*75375*/;
assign _13910_ = _13911_ | _13913_ /*75372*/;
assign _13915_ = ~Q[48] /*75371*/;
assign _13914_ = _13915_ & D[4] /*75370*/;
assign _13917_ = _13381_ & _13914_ /*75365*/;
assign _13918_ = _13381_ ^ _13914_ /*75368*/;
assign _13919_ = _13910_ & _13918_ /*75366*/;
assign _13829_ = _13910_ ^ _13918_ /*75367*/;
assign _13916_ = _13917_ | _13919_ /*75364*/;
assign _13921_ = ~Q[48] /*75363*/;
assign _13920_ = _13921_ & D[5] /*75362*/;
assign _13923_ = _13382_ & _13920_ /*75357*/;
assign _13924_ = _13382_ ^ _13920_ /*75360*/;
assign _13925_ = _13916_ & _13924_ /*75358*/;
assign _13830_ = _13916_ ^ _13924_ /*75359*/;
assign _13922_ = _13923_ | _13925_ /*75356*/;
assign _13927_ = ~Q[48] /*75355*/;
assign _13926_ = _13927_ & D[6] /*75354*/;
assign _13929_ = _13383_ & _13926_ /*75349*/;
assign _13930_ = _13383_ ^ _13926_ /*75352*/;
assign _13931_ = _13922_ & _13930_ /*75350*/;
assign _13831_ = _13922_ ^ _13930_ /*75351*/;
assign _13928_ = _13929_ | _13931_ /*75348*/;
assign _13933_ = ~Q[48] /*75347*/;
assign _13932_ = _13933_ & D[7] /*75346*/;
assign _13935_ = _13384_ & _13932_ /*75341*/;
assign _13936_ = _13384_ ^ _13932_ /*75344*/;
assign _13937_ = _13928_ & _13936_ /*75342*/;
assign _13832_ = _13928_ ^ _13936_ /*75343*/;
assign _13934_ = _13935_ | _13937_ /*75340*/;
assign _13939_ = ~Q[48] /*75339*/;
assign _13938_ = _13939_ & D[8] /*75338*/;
assign _13941_ = _13385_ & _13938_ /*75333*/;
assign _13942_ = _13385_ ^ _13938_ /*75336*/;
assign _13943_ = _13934_ & _13942_ /*75334*/;
assign _13833_ = _13934_ ^ _13942_ /*75335*/;
assign _13940_ = _13941_ | _13943_ /*75332*/;
assign _13945_ = ~Q[48] /*75331*/;
assign _13944_ = _13945_ & D[9] /*75330*/;
assign _13947_ = _13386_ & _13944_ /*75325*/;
assign _13948_ = _13386_ ^ _13944_ /*75328*/;
assign _13949_ = _13940_ & _13948_ /*75326*/;
assign _13834_ = _13940_ ^ _13948_ /*75327*/;
assign _13946_ = _13947_ | _13949_ /*75324*/;
assign _13951_ = ~Q[48] /*75323*/;
assign _13950_ = _13951_ & D[10] /*75322*/;
assign _13953_ = _13387_ & _13950_ /*75317*/;
assign _13954_ = _13387_ ^ _13950_ /*75320*/;
assign _13955_ = _13946_ & _13954_ /*75318*/;
assign _13835_ = _13946_ ^ _13954_ /*75319*/;
assign _13952_ = _13953_ | _13955_ /*75316*/;
assign _13957_ = ~Q[48] /*75315*/;
assign _13956_ = _13957_ & D[11] /*75314*/;
assign _13959_ = _13388_ & _13956_ /*75309*/;
assign _13960_ = _13388_ ^ _13956_ /*75312*/;
assign _13961_ = _13952_ & _13960_ /*75310*/;
assign _13836_ = _13952_ ^ _13960_ /*75311*/;
assign _13958_ = _13959_ | _13961_ /*75308*/;
assign _13963_ = ~Q[48] /*75307*/;
assign _13962_ = _13963_ & D[12] /*75306*/;
assign _13965_ = _13389_ & _13962_ /*75301*/;
assign _13966_ = _13389_ ^ _13962_ /*75304*/;
assign _13967_ = _13958_ & _13966_ /*75302*/;
assign _13837_ = _13958_ ^ _13966_ /*75303*/;
assign _13964_ = _13965_ | _13967_ /*75300*/;
assign _13969_ = ~Q[48] /*75299*/;
assign _13968_ = _13969_ & D[13] /*75298*/;
assign _13971_ = _13390_ & _13968_ /*75293*/;
assign _13972_ = _13390_ ^ _13968_ /*75296*/;
assign _13973_ = _13964_ & _13972_ /*75294*/;
assign _13838_ = _13964_ ^ _13972_ /*75295*/;
assign _13970_ = _13971_ | _13973_ /*75292*/;
assign _13975_ = ~Q[48] /*75291*/;
assign _13974_ = _13975_ & D[14] /*75290*/;
assign _13977_ = _13391_ & _13974_ /*75285*/;
assign _13978_ = _13391_ ^ _13974_ /*75288*/;
assign _13979_ = _13970_ & _13978_ /*75286*/;
assign _13839_ = _13970_ ^ _13978_ /*75287*/;
assign _13976_ = _13977_ | _13979_ /*75284*/;
assign _13981_ = ~Q[48] /*75283*/;
assign _13980_ = _13981_ & D[15] /*75282*/;
assign _13983_ = _13392_ & _13980_ /*75277*/;
assign _13984_ = _13392_ ^ _13980_ /*75280*/;
assign _13985_ = _13976_ & _13984_ /*75278*/;
assign _13840_ = _13976_ ^ _13984_ /*75279*/;
assign _13982_ = _13983_ | _13985_ /*75276*/;
assign _13987_ = ~Q[48] /*75275*/;
assign _13986_ = _13987_ & D[16] /*75274*/;
assign _13989_ = _13393_ & _13986_ /*75269*/;
assign _13990_ = _13393_ ^ _13986_ /*75272*/;
assign _13991_ = _13982_ & _13990_ /*75270*/;
assign _13841_ = _13982_ ^ _13990_ /*75271*/;
assign _13988_ = _13989_ | _13991_ /*75268*/;
assign _13993_ = ~Q[48] /*75267*/;
assign _13992_ = _13993_ & D[17] /*75266*/;
assign _13995_ = _13394_ & _13992_ /*75261*/;
assign _13996_ = _13394_ ^ _13992_ /*75264*/;
assign _13997_ = _13988_ & _13996_ /*75262*/;
assign _13842_ = _13988_ ^ _13996_ /*75263*/;
assign _13994_ = _13995_ | _13997_ /*75260*/;
assign _13999_ = ~Q[48] /*75259*/;
assign _13998_ = _13999_ & D[18] /*75258*/;
assign _14001_ = _13395_ & _13998_ /*75253*/;
assign _14002_ = _13395_ ^ _13998_ /*75256*/;
assign _14003_ = _13994_ & _14002_ /*75254*/;
assign _13843_ = _13994_ ^ _14002_ /*75255*/;
assign _14000_ = _14001_ | _14003_ /*75252*/;
assign _14005_ = ~Q[48] /*75251*/;
assign _14004_ = _14005_ & D[19] /*75250*/;
assign _14007_ = _13396_ & _14004_ /*75245*/;
assign _14008_ = _13396_ ^ _14004_ /*75248*/;
assign _14009_ = _14000_ & _14008_ /*75246*/;
assign _13844_ = _14000_ ^ _14008_ /*75247*/;
assign _14006_ = _14007_ | _14009_ /*75244*/;
assign _14011_ = ~Q[48] /*75243*/;
assign _14010_ = _14011_ & D[20] /*75242*/;
assign _14013_ = _13397_ & _14010_ /*75237*/;
assign _14014_ = _13397_ ^ _14010_ /*75240*/;
assign _14015_ = _14006_ & _14014_ /*75238*/;
assign _13845_ = _14006_ ^ _14014_ /*75239*/;
assign _14012_ = _14013_ | _14015_ /*75236*/;
assign _14017_ = ~Q[48] /*75235*/;
assign _14016_ = _14017_ & D[21] /*75234*/;
assign _14019_ = _13398_ & _14016_ /*75229*/;
assign _14020_ = _13398_ ^ _14016_ /*75232*/;
assign _14021_ = _14012_ & _14020_ /*75230*/;
assign _13846_ = _14012_ ^ _14020_ /*75231*/;
assign _14018_ = _14019_ | _14021_ /*75228*/;
assign _14023_ = ~Q[48] /*75227*/;
assign _14022_ = _14023_ & D[22] /*75226*/;
assign _14025_ = _13399_ & _14022_ /*75221*/;
assign _14026_ = _13399_ ^ _14022_ /*75224*/;
assign _14027_ = _14018_ & _14026_ /*75222*/;
assign _13847_ = _14018_ ^ _14026_ /*75223*/;
assign _14024_ = _14025_ | _14027_ /*75220*/;
assign _14029_ = ~Q[48] /*75219*/;
assign _14028_ = _14029_ & D[23] /*75218*/;
assign _14031_ = _13400_ & _14028_ /*75213*/;
assign _14032_ = _13400_ ^ _14028_ /*75216*/;
assign _14033_ = _14024_ & _14032_ /*75214*/;
assign _13848_ = _14024_ ^ _14032_ /*75215*/;
assign _14030_ = _14031_ | _14033_ /*75212*/;
assign _14035_ = ~Q[48] /*75211*/;
assign _14034_ = _14035_ & D[24] /*75210*/;
assign _14037_ = _13401_ & _14034_ /*75205*/;
assign _14038_ = _13401_ ^ _14034_ /*75208*/;
assign _14039_ = _14030_ & _14038_ /*75206*/;
assign _13849_ = _14030_ ^ _14038_ /*75207*/;
assign _14036_ = _14037_ | _14039_ /*75204*/;
assign _14041_ = ~Q[48] /*75203*/;
assign _14040_ = _14041_ & D[25] /*75202*/;
assign _14043_ = _13402_ & _14040_ /*75197*/;
assign _14044_ = _13402_ ^ _14040_ /*75200*/;
assign _14045_ = _14036_ & _14044_ /*75198*/;
assign _13850_ = _14036_ ^ _14044_ /*75199*/;
assign _14042_ = _14043_ | _14045_ /*75196*/;
assign _14047_ = ~Q[48] /*75195*/;
assign _14046_ = _14047_ & D[26] /*75194*/;
assign _14049_ = _13403_ & _14046_ /*75189*/;
assign _14050_ = _13403_ ^ _14046_ /*75192*/;
assign _14051_ = _14042_ & _14050_ /*75190*/;
assign _13851_ = _14042_ ^ _14050_ /*75191*/;
assign _14048_ = _14049_ | _14051_ /*75188*/;
assign _14053_ = ~Q[48] /*75187*/;
assign _14052_ = _14053_ & D[27] /*75186*/;
assign _14055_ = _13404_ & _14052_ /*75181*/;
assign _14056_ = _13404_ ^ _14052_ /*75184*/;
assign _14057_ = _14048_ & _14056_ /*75182*/;
assign _13852_ = _14048_ ^ _14056_ /*75183*/;
assign _14054_ = _14055_ | _14057_ /*75180*/;
assign _14059_ = ~Q[48] /*75179*/;
assign _14058_ = _14059_ & D[28] /*75178*/;
assign _14061_ = _13405_ & _14058_ /*75173*/;
assign _14062_ = _13405_ ^ _14058_ /*75176*/;
assign _14063_ = _14054_ & _14062_ /*75174*/;
assign _13853_ = _14054_ ^ _14062_ /*75175*/;
assign _14060_ = _14061_ | _14063_ /*75172*/;
assign _14065_ = ~Q[48] /*75171*/;
assign _14064_ = _14065_ & D[29] /*75170*/;
assign _14067_ = _13406_ & _14064_ /*75165*/;
assign _14068_ = _13406_ ^ _14064_ /*75168*/;
assign _14069_ = _14060_ & _14068_ /*75166*/;
assign _13854_ = _14060_ ^ _14068_ /*75167*/;
assign _14066_ = _14067_ | _14069_ /*75164*/;
assign _14071_ = ~Q[48] /*75163*/;
assign _14070_ = _14071_ & D[30] /*75162*/;
assign _14073_ = _13407_ & _14070_ /*75157*/;
assign _14074_ = _13407_ ^ _14070_ /*75160*/;
assign _14075_ = _14066_ & _14074_ /*75158*/;
assign _13855_ = _14066_ ^ _14074_ /*75159*/;
assign _14072_ = _14073_ | _14075_ /*75156*/;
assign _14077_ = ~Q[48] /*75155*/;
assign _14076_ = _14077_ & D[31] /*75154*/;
assign _14079_ = _13408_ & _14076_ /*75149*/;
assign _14080_ = _13408_ ^ _14076_ /*75152*/;
assign _14081_ = _14072_ & _14080_ /*75150*/;
assign _13856_ = _14072_ ^ _14080_ /*75151*/;
assign _14078_ = _14079_ | _14081_ /*75148*/;
assign _14083_ = ~Q[48] /*75147*/;
assign _14082_ = _14083_ & D[32] /*75146*/;
assign _14085_ = _13409_ & _14082_ /*75141*/;
assign _14086_ = _13409_ ^ _14082_ /*75144*/;
assign _14087_ = _14078_ & _14086_ /*75142*/;
assign _13857_ = _14078_ ^ _14086_ /*75143*/;
assign _14084_ = _14085_ | _14087_ /*75140*/;
assign _14089_ = ~Q[48] /*75139*/;
assign _14088_ = _14089_ & D[33] /*75138*/;
assign _14091_ = _13410_ & _14088_ /*75133*/;
assign _14092_ = _13410_ ^ _14088_ /*75136*/;
assign _14093_ = _14084_ & _14092_ /*75134*/;
assign _13858_ = _14084_ ^ _14092_ /*75135*/;
assign _14090_ = _14091_ | _14093_ /*75132*/;
assign _14095_ = ~Q[48] /*75131*/;
assign _14094_ = _14095_ & D[34] /*75130*/;
assign _14097_ = _13411_ & _14094_ /*75125*/;
assign _14098_ = _13411_ ^ _14094_ /*75128*/;
assign _14099_ = _14090_ & _14098_ /*75126*/;
assign _13859_ = _14090_ ^ _14098_ /*75127*/;
assign _14096_ = _14097_ | _14099_ /*75124*/;
assign _14101_ = ~Q[48] /*75123*/;
assign _14100_ = _14101_ & D[35] /*75122*/;
assign _14103_ = _13412_ & _14100_ /*75117*/;
assign _14104_ = _13412_ ^ _14100_ /*75120*/;
assign _14105_ = _14096_ & _14104_ /*75118*/;
assign _13860_ = _14096_ ^ _14104_ /*75119*/;
assign _14102_ = _14103_ | _14105_ /*75116*/;
assign _14107_ = ~Q[48] /*75115*/;
assign _14106_ = _14107_ & D[36] /*75114*/;
assign _14109_ = _13413_ & _14106_ /*75109*/;
assign _14110_ = _13413_ ^ _14106_ /*75112*/;
assign _14111_ = _14102_ & _14110_ /*75110*/;
assign _13861_ = _14102_ ^ _14110_ /*75111*/;
assign _14108_ = _14109_ | _14111_ /*75108*/;
assign _14113_ = ~Q[48] /*75107*/;
assign _14112_ = _14113_ & D[37] /*75106*/;
assign _14115_ = _13414_ & _14112_ /*75101*/;
assign _14116_ = _13414_ ^ _14112_ /*75104*/;
assign _14117_ = _14108_ & _14116_ /*75102*/;
assign _13862_ = _14108_ ^ _14116_ /*75103*/;
assign _14114_ = _14115_ | _14117_ /*75100*/;
assign _14119_ = ~Q[48] /*75099*/;
assign _14118_ = _14119_ & D[38] /*75098*/;
assign _14121_ = _13415_ & _14118_ /*75093*/;
assign _14122_ = _13415_ ^ _14118_ /*75096*/;
assign _14123_ = _14114_ & _14122_ /*75094*/;
assign _13863_ = _14114_ ^ _14122_ /*75095*/;
assign _14120_ = _14121_ | _14123_ /*75092*/;
assign _14125_ = ~Q[48] /*75091*/;
assign _14124_ = _14125_ & D[39] /*75090*/;
assign _14127_ = _13416_ & _14124_ /*75085*/;
assign _14128_ = _13416_ ^ _14124_ /*75088*/;
assign _14129_ = _14120_ & _14128_ /*75086*/;
assign _13864_ = _14120_ ^ _14128_ /*75087*/;
assign _14126_ = _14127_ | _14129_ /*75084*/;
assign _14131_ = ~Q[48] /*75083*/;
assign _14130_ = _14131_ & D[40] /*75082*/;
assign _14133_ = _13417_ & _14130_ /*75077*/;
assign _14134_ = _13417_ ^ _14130_ /*75080*/;
assign _14135_ = _14126_ & _14134_ /*75078*/;
assign _13865_ = _14126_ ^ _14134_ /*75079*/;
assign _14132_ = _14133_ | _14135_ /*75076*/;
assign _14137_ = ~Q[48] /*75075*/;
assign _14136_ = _14137_ & D[41] /*75074*/;
assign _14139_ = _13418_ & _14136_ /*75069*/;
assign _14140_ = _13418_ ^ _14136_ /*75072*/;
assign _14141_ = _14132_ & _14140_ /*75070*/;
assign _13866_ = _14132_ ^ _14140_ /*75071*/;
assign _14138_ = _14139_ | _14141_ /*75068*/;
assign _14143_ = ~Q[48] /*75067*/;
assign _14142_ = _14143_ & D[42] /*75066*/;
assign _14145_ = _13419_ & _14142_ /*75061*/;
assign _14146_ = _13419_ ^ _14142_ /*75064*/;
assign _14147_ = _14138_ & _14146_ /*75062*/;
assign _13867_ = _14138_ ^ _14146_ /*75063*/;
assign _14144_ = _14145_ | _14147_ /*75060*/;
assign _14149_ = ~Q[48] /*75059*/;
assign _14148_ = _14149_ & D[43] /*75058*/;
assign _14151_ = _13420_ & _14148_ /*75053*/;
assign _14152_ = _13420_ ^ _14148_ /*75056*/;
assign _14153_ = _14144_ & _14152_ /*75054*/;
assign _13868_ = _14144_ ^ _14152_ /*75055*/;
assign _14150_ = _14151_ | _14153_ /*75052*/;
assign _14155_ = ~Q[48] /*75051*/;
assign _14154_ = _14155_ & D[44] /*75050*/;
assign _14157_ = _13421_ & _14154_ /*75045*/;
assign _14158_ = _13421_ ^ _14154_ /*75048*/;
assign _14159_ = _14150_ & _14158_ /*75046*/;
assign _13869_ = _14150_ ^ _14158_ /*75047*/;
assign _14156_ = _14157_ | _14159_ /*75044*/;
assign _14161_ = ~Q[48] /*75043*/;
assign _14160_ = _14161_ & D[45] /*75042*/;
assign _14163_ = _13422_ & _14160_ /*75037*/;
assign _14164_ = _13422_ ^ _14160_ /*75040*/;
assign _14165_ = _14156_ & _14164_ /*75038*/;
assign _13870_ = _14156_ ^ _14164_ /*75039*/;
assign _14162_ = _14163_ | _14165_ /*75036*/;
assign _14167_ = ~Q[48] /*75035*/;
assign _14166_ = _14167_ & D[46] /*75034*/;
assign _14169_ = _13423_ & _14166_ /*75029*/;
assign _14170_ = _13423_ ^ _14166_ /*75032*/;
assign _14171_ = _14162_ & _14170_ /*75030*/;
assign _13871_ = _14162_ ^ _14170_ /*75031*/;
assign _14168_ = _14169_ | _14171_ /*75028*/;
assign _14173_ = ~Q[48] /*75027*/;
assign _14172_ = _14173_ & D[47] /*75026*/;
assign _14175_ = _13424_ & _14172_ /*75021*/;
assign _14176_ = _13424_ ^ _14172_ /*75024*/;
assign _14177_ = _14168_ & _14176_ /*75022*/;
assign _13872_ = _14168_ ^ _14176_ /*75023*/;
assign _14174_ = _14175_ | _14177_ /*75020*/;
assign _14179_ = ~Q[48] /*75019*/;
assign _14178_ = _14179_ & D[48] /*75018*/;
assign _14181_ = _13425_ & _14178_ /*75013*/;
assign _14182_ = _13425_ ^ _14178_ /*75016*/;
assign _14183_ = _14174_ & _14182_ /*75014*/;
assign _13873_ = _14174_ ^ _14182_ /*75015*/;
assign _14180_ = _14181_ | _14183_ /*75012*/;
assign _14185_ = ~Q[48] /*75011*/;
assign _14184_ = _14185_ & D[49] /*75010*/;
assign _14187_ = _13426_ & _14184_ /*75005*/;
assign _14188_ = _13426_ ^ _14184_ /*75008*/;
assign _14189_ = _14180_ & _14188_ /*75006*/;
assign _13874_ = _14180_ ^ _14188_ /*75007*/;
assign _14186_ = _14187_ | _14189_ /*75004*/;
assign _14191_ = ~Q[48] /*75003*/;
assign _14190_ = _14191_ & D[50] /*75002*/;
assign _14193_ = _13427_ & _14190_ /*74997*/;
assign _14194_ = _13427_ ^ _14190_ /*75000*/;
assign _14195_ = _14186_ & _14194_ /*74998*/;
assign _13875_ = _14186_ ^ _14194_ /*74999*/;
assign _14192_ = _14193_ | _14195_ /*74996*/;
assign _14197_ = ~Q[48] /*74995*/;
assign _14196_ = _14197_ & D[51] /*74994*/;
assign _14199_ = _13428_ & _14196_ /*74989*/;
assign _14200_ = _13428_ ^ _14196_ /*74992*/;
assign _14201_ = _14192_ & _14200_ /*74990*/;
assign _13876_ = _14192_ ^ _14200_ /*74991*/;
assign _14198_ = _14199_ | _14201_ /*74988*/;
assign _14203_ = ~Q[48] /*74987*/;
assign _14202_ = _14203_ & D[52] /*74986*/;
assign _14205_ = _13429_ & _14202_ /*74981*/;
assign _14206_ = _13429_ ^ _14202_ /*74984*/;
assign _14207_ = _14198_ & _14206_ /*74982*/;
assign _13877_ = _14198_ ^ _14206_ /*74983*/;
assign _14204_ = _14205_ | _14207_ /*74980*/;
assign _14209_ = ~Q[48] /*74979*/;
assign _14208_ = _14209_ & D[53] /*74978*/;
assign _14211_ = _13430_ & _14208_ /*74973*/;
assign _14212_ = _13430_ ^ _14208_ /*74976*/;
assign _14213_ = _14204_ & _14212_ /*74974*/;
assign _13878_ = _14204_ ^ _14212_ /*74975*/;
assign _14210_ = _14211_ | _14213_ /*74972*/;
assign _14215_ = ~Q[48] /*74971*/;
assign _14214_ = _14215_ & D[54] /*74970*/;
assign _14217_ = _13431_ & _14214_ /*74965*/;
assign _14218_ = _13431_ ^ _14214_ /*74968*/;
assign _14219_ = _14210_ & _14218_ /*74966*/;
assign _13879_ = _14210_ ^ _14218_ /*74967*/;
assign _14216_ = _14217_ | _14219_ /*74964*/;
assign _14221_ = ~Q[48] /*74963*/;
assign _14220_ = _14221_ & D[55] /*74962*/;
assign _14223_ = _13432_ & _14220_ /*74957*/;
assign _14224_ = _13432_ ^ _14220_ /*74960*/;
assign _14225_ = _14216_ & _14224_ /*74958*/;
assign _13880_ = _14216_ ^ _14224_ /*74959*/;
assign _14222_ = _14223_ | _14225_ /*74956*/;
assign _14227_ = ~Q[48] /*74955*/;
assign _14226_ = _14227_ & D[56] /*74954*/;
assign _14229_ = _13433_ & _14226_ /*74949*/;
assign _14230_ = _13433_ ^ _14226_ /*74952*/;
assign _14231_ = _14222_ & _14230_ /*74950*/;
assign _13881_ = _14222_ ^ _14230_ /*74951*/;
assign _14228_ = _14229_ | _14231_ /*74948*/;
assign _14233_ = ~Q[48] /*74947*/;
assign _14232_ = _14233_ & D[57] /*74946*/;
assign _14235_ = _13434_ & _14232_ /*74941*/;
assign _14236_ = _13434_ ^ _14232_ /*74944*/;
assign _14237_ = _14228_ & _14236_ /*74942*/;
assign _13882_ = _14228_ ^ _14236_ /*74943*/;
assign _14234_ = _14235_ | _14237_ /*74940*/;
assign _14239_ = ~Q[48] /*74939*/;
assign _14238_ = _14239_ & D[58] /*74938*/;
assign _14241_ = _13435_ & _14238_ /*74933*/;
assign _14242_ = _13435_ ^ _14238_ /*74936*/;
assign _14243_ = _14234_ & _14242_ /*74934*/;
assign _13883_ = _14234_ ^ _14242_ /*74935*/;
assign _14240_ = _14241_ | _14243_ /*74932*/;
assign _14245_ = ~Q[48] /*74931*/;
assign _14244_ = _14245_ & D[59] /*74930*/;
assign _14247_ = _13436_ & _14244_ /*74925*/;
assign _14248_ = _13436_ ^ _14244_ /*74928*/;
assign _14249_ = _14240_ & _14248_ /*74926*/;
assign _13884_ = _14240_ ^ _14248_ /*74927*/;
assign _14246_ = _14247_ | _14249_ /*74924*/;
assign _14251_ = ~Q[48] /*74923*/;
assign _14250_ = _14251_ & D[60] /*74922*/;
assign _14253_ = _13437_ & _14250_ /*74917*/;
assign _14254_ = _13437_ ^ _14250_ /*74920*/;
assign _14255_ = _14246_ & _14254_ /*74918*/;
assign _13885_ = _14246_ ^ _14254_ /*74919*/;
assign _14252_ = _14253_ | _14255_ /*74916*/;
assign _14257_ = ~Q[48] /*74915*/;
assign _14256_ = _14257_ & D[61] /*74914*/;
assign _14259_ = _13438_ & _14256_ /*74909*/;
assign _14260_ = _13438_ ^ _14256_ /*74912*/;
assign _14261_ = _14252_ & _14260_ /*74910*/;
assign _13886_ = _14252_ ^ _14260_ /*74911*/;
assign _14258_ = _14259_ | _14261_ /*74908*/;
assign _14263_ = ~Q[48] /*74907*/;
assign _14262_ = _14263_ & D[62] /*74906*/;
assign _14265_ = _13439_ & _14262_ /*74901*/;
assign _14266_ = _13439_ ^ _14262_ /*74904*/;
assign _14267_ = _14258_ & _14266_ /*74902*/;
assign _13887_ = _14258_ ^ _14266_ /*74903*/;
assign _14264_ = _14265_ | _14267_ /*74900*/;
assign _14269_ = ~Q[48] /*74899*/;
assign _14268_ = _14269_ & zeroWire /*74898*/;
assign _14270_ = _13440_ ^ _14268_ /*74896*/;
assign _13888_ = _14270_ ^ _14264_ /*74895*/;
assign _14341_ = ~D[0] /*74641*/;
assign _14338_ = R_0[47] & _14341_ /*74637*/;
assign _14339_ = R_0[47] ^ _14341_ /*74640*/;
assign _14340_ = oneWire & _14339_ /*74638*/;
assign _14273_ = oneWire ^ _14339_ /*74639*/;
assign _14337_ = _14338_ | _14340_ /*74636*/;
assign _14346_ = ~D[1] /*74635*/;
assign _14343_ = _13825_ & _14346_ /*74631*/;
assign _14344_ = _13825_ ^ _14346_ /*74634*/;
assign _14345_ = _14337_ & _14344_ /*74632*/;
assign _14274_ = _14337_ ^ _14344_ /*74633*/;
assign _14342_ = _14343_ | _14345_ /*74630*/;
assign _14351_ = ~D[2] /*74629*/;
assign _14348_ = _13826_ & _14351_ /*74625*/;
assign _14349_ = _13826_ ^ _14351_ /*74628*/;
assign _14350_ = _14342_ & _14349_ /*74626*/;
assign _14275_ = _14342_ ^ _14349_ /*74627*/;
assign _14347_ = _14348_ | _14350_ /*74624*/;
assign _14356_ = ~D[3] /*74623*/;
assign _14353_ = _13827_ & _14356_ /*74619*/;
assign _14354_ = _13827_ ^ _14356_ /*74622*/;
assign _14355_ = _14347_ & _14354_ /*74620*/;
assign _14276_ = _14347_ ^ _14354_ /*74621*/;
assign _14352_ = _14353_ | _14355_ /*74618*/;
assign _14361_ = ~D[4] /*74617*/;
assign _14358_ = _13828_ & _14361_ /*74613*/;
assign _14359_ = _13828_ ^ _14361_ /*74616*/;
assign _14360_ = _14352_ & _14359_ /*74614*/;
assign _14277_ = _14352_ ^ _14359_ /*74615*/;
assign _14357_ = _14358_ | _14360_ /*74612*/;
assign _14366_ = ~D[5] /*74611*/;
assign _14363_ = _13829_ & _14366_ /*74607*/;
assign _14364_ = _13829_ ^ _14366_ /*74610*/;
assign _14365_ = _14357_ & _14364_ /*74608*/;
assign _14278_ = _14357_ ^ _14364_ /*74609*/;
assign _14362_ = _14363_ | _14365_ /*74606*/;
assign _14371_ = ~D[6] /*74605*/;
assign _14368_ = _13830_ & _14371_ /*74601*/;
assign _14369_ = _13830_ ^ _14371_ /*74604*/;
assign _14370_ = _14362_ & _14369_ /*74602*/;
assign _14279_ = _14362_ ^ _14369_ /*74603*/;
assign _14367_ = _14368_ | _14370_ /*74600*/;
assign _14376_ = ~D[7] /*74599*/;
assign _14373_ = _13831_ & _14376_ /*74595*/;
assign _14374_ = _13831_ ^ _14376_ /*74598*/;
assign _14375_ = _14367_ & _14374_ /*74596*/;
assign _14280_ = _14367_ ^ _14374_ /*74597*/;
assign _14372_ = _14373_ | _14375_ /*74594*/;
assign _14381_ = ~D[8] /*74593*/;
assign _14378_ = _13832_ & _14381_ /*74589*/;
assign _14379_ = _13832_ ^ _14381_ /*74592*/;
assign _14380_ = _14372_ & _14379_ /*74590*/;
assign _14281_ = _14372_ ^ _14379_ /*74591*/;
assign _14377_ = _14378_ | _14380_ /*74588*/;
assign _14386_ = ~D[9] /*74587*/;
assign _14383_ = _13833_ & _14386_ /*74583*/;
assign _14384_ = _13833_ ^ _14386_ /*74586*/;
assign _14385_ = _14377_ & _14384_ /*74584*/;
assign _14282_ = _14377_ ^ _14384_ /*74585*/;
assign _14382_ = _14383_ | _14385_ /*74582*/;
assign _14391_ = ~D[10] /*74581*/;
assign _14388_ = _13834_ & _14391_ /*74577*/;
assign _14389_ = _13834_ ^ _14391_ /*74580*/;
assign _14390_ = _14382_ & _14389_ /*74578*/;
assign _14283_ = _14382_ ^ _14389_ /*74579*/;
assign _14387_ = _14388_ | _14390_ /*74576*/;
assign _14396_ = ~D[11] /*74575*/;
assign _14393_ = _13835_ & _14396_ /*74571*/;
assign _14394_ = _13835_ ^ _14396_ /*74574*/;
assign _14395_ = _14387_ & _14394_ /*74572*/;
assign _14284_ = _14387_ ^ _14394_ /*74573*/;
assign _14392_ = _14393_ | _14395_ /*74570*/;
assign _14401_ = ~D[12] /*74569*/;
assign _14398_ = _13836_ & _14401_ /*74565*/;
assign _14399_ = _13836_ ^ _14401_ /*74568*/;
assign _14400_ = _14392_ & _14399_ /*74566*/;
assign _14285_ = _14392_ ^ _14399_ /*74567*/;
assign _14397_ = _14398_ | _14400_ /*74564*/;
assign _14406_ = ~D[13] /*74563*/;
assign _14403_ = _13837_ & _14406_ /*74559*/;
assign _14404_ = _13837_ ^ _14406_ /*74562*/;
assign _14405_ = _14397_ & _14404_ /*74560*/;
assign _14286_ = _14397_ ^ _14404_ /*74561*/;
assign _14402_ = _14403_ | _14405_ /*74558*/;
assign _14411_ = ~D[14] /*74557*/;
assign _14408_ = _13838_ & _14411_ /*74553*/;
assign _14409_ = _13838_ ^ _14411_ /*74556*/;
assign _14410_ = _14402_ & _14409_ /*74554*/;
assign _14287_ = _14402_ ^ _14409_ /*74555*/;
assign _14407_ = _14408_ | _14410_ /*74552*/;
assign _14416_ = ~D[15] /*74551*/;
assign _14413_ = _13839_ & _14416_ /*74547*/;
assign _14414_ = _13839_ ^ _14416_ /*74550*/;
assign _14415_ = _14407_ & _14414_ /*74548*/;
assign _14288_ = _14407_ ^ _14414_ /*74549*/;
assign _14412_ = _14413_ | _14415_ /*74546*/;
assign _14421_ = ~D[16] /*74545*/;
assign _14418_ = _13840_ & _14421_ /*74541*/;
assign _14419_ = _13840_ ^ _14421_ /*74544*/;
assign _14420_ = _14412_ & _14419_ /*74542*/;
assign _14289_ = _14412_ ^ _14419_ /*74543*/;
assign _14417_ = _14418_ | _14420_ /*74540*/;
assign _14426_ = ~D[17] /*74539*/;
assign _14423_ = _13841_ & _14426_ /*74535*/;
assign _14424_ = _13841_ ^ _14426_ /*74538*/;
assign _14425_ = _14417_ & _14424_ /*74536*/;
assign _14290_ = _14417_ ^ _14424_ /*74537*/;
assign _14422_ = _14423_ | _14425_ /*74534*/;
assign _14431_ = ~D[18] /*74533*/;
assign _14428_ = _13842_ & _14431_ /*74529*/;
assign _14429_ = _13842_ ^ _14431_ /*74532*/;
assign _14430_ = _14422_ & _14429_ /*74530*/;
assign _14291_ = _14422_ ^ _14429_ /*74531*/;
assign _14427_ = _14428_ | _14430_ /*74528*/;
assign _14436_ = ~D[19] /*74527*/;
assign _14433_ = _13843_ & _14436_ /*74523*/;
assign _14434_ = _13843_ ^ _14436_ /*74526*/;
assign _14435_ = _14427_ & _14434_ /*74524*/;
assign _14292_ = _14427_ ^ _14434_ /*74525*/;
assign _14432_ = _14433_ | _14435_ /*74522*/;
assign _14441_ = ~D[20] /*74521*/;
assign _14438_ = _13844_ & _14441_ /*74517*/;
assign _14439_ = _13844_ ^ _14441_ /*74520*/;
assign _14440_ = _14432_ & _14439_ /*74518*/;
assign _14293_ = _14432_ ^ _14439_ /*74519*/;
assign _14437_ = _14438_ | _14440_ /*74516*/;
assign _14446_ = ~D[21] /*74515*/;
assign _14443_ = _13845_ & _14446_ /*74511*/;
assign _14444_ = _13845_ ^ _14446_ /*74514*/;
assign _14445_ = _14437_ & _14444_ /*74512*/;
assign _14294_ = _14437_ ^ _14444_ /*74513*/;
assign _14442_ = _14443_ | _14445_ /*74510*/;
assign _14451_ = ~D[22] /*74509*/;
assign _14448_ = _13846_ & _14451_ /*74505*/;
assign _14449_ = _13846_ ^ _14451_ /*74508*/;
assign _14450_ = _14442_ & _14449_ /*74506*/;
assign _14295_ = _14442_ ^ _14449_ /*74507*/;
assign _14447_ = _14448_ | _14450_ /*74504*/;
assign _14456_ = ~D[23] /*74503*/;
assign _14453_ = _13847_ & _14456_ /*74499*/;
assign _14454_ = _13847_ ^ _14456_ /*74502*/;
assign _14455_ = _14447_ & _14454_ /*74500*/;
assign _14296_ = _14447_ ^ _14454_ /*74501*/;
assign _14452_ = _14453_ | _14455_ /*74498*/;
assign _14461_ = ~D[24] /*74497*/;
assign _14458_ = _13848_ & _14461_ /*74493*/;
assign _14459_ = _13848_ ^ _14461_ /*74496*/;
assign _14460_ = _14452_ & _14459_ /*74494*/;
assign _14297_ = _14452_ ^ _14459_ /*74495*/;
assign _14457_ = _14458_ | _14460_ /*74492*/;
assign _14466_ = ~D[25] /*74491*/;
assign _14463_ = _13849_ & _14466_ /*74487*/;
assign _14464_ = _13849_ ^ _14466_ /*74490*/;
assign _14465_ = _14457_ & _14464_ /*74488*/;
assign _14298_ = _14457_ ^ _14464_ /*74489*/;
assign _14462_ = _14463_ | _14465_ /*74486*/;
assign _14471_ = ~D[26] /*74485*/;
assign _14468_ = _13850_ & _14471_ /*74481*/;
assign _14469_ = _13850_ ^ _14471_ /*74484*/;
assign _14470_ = _14462_ & _14469_ /*74482*/;
assign _14299_ = _14462_ ^ _14469_ /*74483*/;
assign _14467_ = _14468_ | _14470_ /*74480*/;
assign _14476_ = ~D[27] /*74479*/;
assign _14473_ = _13851_ & _14476_ /*74475*/;
assign _14474_ = _13851_ ^ _14476_ /*74478*/;
assign _14475_ = _14467_ & _14474_ /*74476*/;
assign _14300_ = _14467_ ^ _14474_ /*74477*/;
assign _14472_ = _14473_ | _14475_ /*74474*/;
assign _14481_ = ~D[28] /*74473*/;
assign _14478_ = _13852_ & _14481_ /*74469*/;
assign _14479_ = _13852_ ^ _14481_ /*74472*/;
assign _14480_ = _14472_ & _14479_ /*74470*/;
assign _14301_ = _14472_ ^ _14479_ /*74471*/;
assign _14477_ = _14478_ | _14480_ /*74468*/;
assign _14486_ = ~D[29] /*74467*/;
assign _14483_ = _13853_ & _14486_ /*74463*/;
assign _14484_ = _13853_ ^ _14486_ /*74466*/;
assign _14485_ = _14477_ & _14484_ /*74464*/;
assign _14302_ = _14477_ ^ _14484_ /*74465*/;
assign _14482_ = _14483_ | _14485_ /*74462*/;
assign _14491_ = ~D[30] /*74461*/;
assign _14488_ = _13854_ & _14491_ /*74457*/;
assign _14489_ = _13854_ ^ _14491_ /*74460*/;
assign _14490_ = _14482_ & _14489_ /*74458*/;
assign _14303_ = _14482_ ^ _14489_ /*74459*/;
assign _14487_ = _14488_ | _14490_ /*74456*/;
assign _14496_ = ~D[31] /*74455*/;
assign _14493_ = _13855_ & _14496_ /*74451*/;
assign _14494_ = _13855_ ^ _14496_ /*74454*/;
assign _14495_ = _14487_ & _14494_ /*74452*/;
assign _14304_ = _14487_ ^ _14494_ /*74453*/;
assign _14492_ = _14493_ | _14495_ /*74450*/;
assign _14501_ = ~D[32] /*74449*/;
assign _14498_ = _13856_ & _14501_ /*74445*/;
assign _14499_ = _13856_ ^ _14501_ /*74448*/;
assign _14500_ = _14492_ & _14499_ /*74446*/;
assign _14305_ = _14492_ ^ _14499_ /*74447*/;
assign _14497_ = _14498_ | _14500_ /*74444*/;
assign _14506_ = ~D[33] /*74443*/;
assign _14503_ = _13857_ & _14506_ /*74439*/;
assign _14504_ = _13857_ ^ _14506_ /*74442*/;
assign _14505_ = _14497_ & _14504_ /*74440*/;
assign _14306_ = _14497_ ^ _14504_ /*74441*/;
assign _14502_ = _14503_ | _14505_ /*74438*/;
assign _14511_ = ~D[34] /*74437*/;
assign _14508_ = _13858_ & _14511_ /*74433*/;
assign _14509_ = _13858_ ^ _14511_ /*74436*/;
assign _14510_ = _14502_ & _14509_ /*74434*/;
assign _14307_ = _14502_ ^ _14509_ /*74435*/;
assign _14507_ = _14508_ | _14510_ /*74432*/;
assign _14516_ = ~D[35] /*74431*/;
assign _14513_ = _13859_ & _14516_ /*74427*/;
assign _14514_ = _13859_ ^ _14516_ /*74430*/;
assign _14515_ = _14507_ & _14514_ /*74428*/;
assign _14308_ = _14507_ ^ _14514_ /*74429*/;
assign _14512_ = _14513_ | _14515_ /*74426*/;
assign _14521_ = ~D[36] /*74425*/;
assign _14518_ = _13860_ & _14521_ /*74421*/;
assign _14519_ = _13860_ ^ _14521_ /*74424*/;
assign _14520_ = _14512_ & _14519_ /*74422*/;
assign _14309_ = _14512_ ^ _14519_ /*74423*/;
assign _14517_ = _14518_ | _14520_ /*74420*/;
assign _14526_ = ~D[37] /*74419*/;
assign _14523_ = _13861_ & _14526_ /*74415*/;
assign _14524_ = _13861_ ^ _14526_ /*74418*/;
assign _14525_ = _14517_ & _14524_ /*74416*/;
assign _14310_ = _14517_ ^ _14524_ /*74417*/;
assign _14522_ = _14523_ | _14525_ /*74414*/;
assign _14531_ = ~D[38] /*74413*/;
assign _14528_ = _13862_ & _14531_ /*74409*/;
assign _14529_ = _13862_ ^ _14531_ /*74412*/;
assign _14530_ = _14522_ & _14529_ /*74410*/;
assign _14311_ = _14522_ ^ _14529_ /*74411*/;
assign _14527_ = _14528_ | _14530_ /*74408*/;
assign _14536_ = ~D[39] /*74407*/;
assign _14533_ = _13863_ & _14536_ /*74403*/;
assign _14534_ = _13863_ ^ _14536_ /*74406*/;
assign _14535_ = _14527_ & _14534_ /*74404*/;
assign _14312_ = _14527_ ^ _14534_ /*74405*/;
assign _14532_ = _14533_ | _14535_ /*74402*/;
assign _14541_ = ~D[40] /*74401*/;
assign _14538_ = _13864_ & _14541_ /*74397*/;
assign _14539_ = _13864_ ^ _14541_ /*74400*/;
assign _14540_ = _14532_ & _14539_ /*74398*/;
assign _14313_ = _14532_ ^ _14539_ /*74399*/;
assign _14537_ = _14538_ | _14540_ /*74396*/;
assign _14546_ = ~D[41] /*74395*/;
assign _14543_ = _13865_ & _14546_ /*74391*/;
assign _14544_ = _13865_ ^ _14546_ /*74394*/;
assign _14545_ = _14537_ & _14544_ /*74392*/;
assign _14314_ = _14537_ ^ _14544_ /*74393*/;
assign _14542_ = _14543_ | _14545_ /*74390*/;
assign _14551_ = ~D[42] /*74389*/;
assign _14548_ = _13866_ & _14551_ /*74385*/;
assign _14549_ = _13866_ ^ _14551_ /*74388*/;
assign _14550_ = _14542_ & _14549_ /*74386*/;
assign _14315_ = _14542_ ^ _14549_ /*74387*/;
assign _14547_ = _14548_ | _14550_ /*74384*/;
assign _14556_ = ~D[43] /*74383*/;
assign _14553_ = _13867_ & _14556_ /*74379*/;
assign _14554_ = _13867_ ^ _14556_ /*74382*/;
assign _14555_ = _14547_ & _14554_ /*74380*/;
assign _14316_ = _14547_ ^ _14554_ /*74381*/;
assign _14552_ = _14553_ | _14555_ /*74378*/;
assign _14561_ = ~D[44] /*74377*/;
assign _14558_ = _13868_ & _14561_ /*74373*/;
assign _14559_ = _13868_ ^ _14561_ /*74376*/;
assign _14560_ = _14552_ & _14559_ /*74374*/;
assign _14317_ = _14552_ ^ _14559_ /*74375*/;
assign _14557_ = _14558_ | _14560_ /*74372*/;
assign _14566_ = ~D[45] /*74371*/;
assign _14563_ = _13869_ & _14566_ /*74367*/;
assign _14564_ = _13869_ ^ _14566_ /*74370*/;
assign _14565_ = _14557_ & _14564_ /*74368*/;
assign _14318_ = _14557_ ^ _14564_ /*74369*/;
assign _14562_ = _14563_ | _14565_ /*74366*/;
assign _14571_ = ~D[46] /*74365*/;
assign _14568_ = _13870_ & _14571_ /*74361*/;
assign _14569_ = _13870_ ^ _14571_ /*74364*/;
assign _14570_ = _14562_ & _14569_ /*74362*/;
assign _14319_ = _14562_ ^ _14569_ /*74363*/;
assign _14567_ = _14568_ | _14570_ /*74360*/;
assign _14576_ = ~D[47] /*74359*/;
assign _14573_ = _13871_ & _14576_ /*74355*/;
assign _14574_ = _13871_ ^ _14576_ /*74358*/;
assign _14575_ = _14567_ & _14574_ /*74356*/;
assign _14320_ = _14567_ ^ _14574_ /*74357*/;
assign _14572_ = _14573_ | _14575_ /*74354*/;
assign _14581_ = ~D[48] /*74353*/;
assign _14578_ = _13872_ & _14581_ /*74349*/;
assign _14579_ = _13872_ ^ _14581_ /*74352*/;
assign _14580_ = _14572_ & _14579_ /*74350*/;
assign _14321_ = _14572_ ^ _14579_ /*74351*/;
assign _14577_ = _14578_ | _14580_ /*74348*/;
assign _14586_ = ~D[49] /*74347*/;
assign _14583_ = _13873_ & _14586_ /*74343*/;
assign _14584_ = _13873_ ^ _14586_ /*74346*/;
assign _14585_ = _14577_ & _14584_ /*74344*/;
assign _14322_ = _14577_ ^ _14584_ /*74345*/;
assign _14582_ = _14583_ | _14585_ /*74342*/;
assign _14591_ = ~D[50] /*74341*/;
assign _14588_ = _13874_ & _14591_ /*74337*/;
assign _14589_ = _13874_ ^ _14591_ /*74340*/;
assign _14590_ = _14582_ & _14589_ /*74338*/;
assign _14323_ = _14582_ ^ _14589_ /*74339*/;
assign _14587_ = _14588_ | _14590_ /*74336*/;
assign _14596_ = ~D[51] /*74335*/;
assign _14593_ = _13875_ & _14596_ /*74331*/;
assign _14594_ = _13875_ ^ _14596_ /*74334*/;
assign _14595_ = _14587_ & _14594_ /*74332*/;
assign _14324_ = _14587_ ^ _14594_ /*74333*/;
assign _14592_ = _14593_ | _14595_ /*74330*/;
assign _14601_ = ~D[52] /*74329*/;
assign _14598_ = _13876_ & _14601_ /*74325*/;
assign _14599_ = _13876_ ^ _14601_ /*74328*/;
assign _14600_ = _14592_ & _14599_ /*74326*/;
assign _14325_ = _14592_ ^ _14599_ /*74327*/;
assign _14597_ = _14598_ | _14600_ /*74324*/;
assign _14606_ = ~D[53] /*74323*/;
assign _14603_ = _13877_ & _14606_ /*74319*/;
assign _14604_ = _13877_ ^ _14606_ /*74322*/;
assign _14605_ = _14597_ & _14604_ /*74320*/;
assign _14326_ = _14597_ ^ _14604_ /*74321*/;
assign _14602_ = _14603_ | _14605_ /*74318*/;
assign _14611_ = ~D[54] /*74317*/;
assign _14608_ = _13878_ & _14611_ /*74313*/;
assign _14609_ = _13878_ ^ _14611_ /*74316*/;
assign _14610_ = _14602_ & _14609_ /*74314*/;
assign _14327_ = _14602_ ^ _14609_ /*74315*/;
assign _14607_ = _14608_ | _14610_ /*74312*/;
assign _14616_ = ~D[55] /*74311*/;
assign _14613_ = _13879_ & _14616_ /*74307*/;
assign _14614_ = _13879_ ^ _14616_ /*74310*/;
assign _14615_ = _14607_ & _14614_ /*74308*/;
assign _14328_ = _14607_ ^ _14614_ /*74309*/;
assign _14612_ = _14613_ | _14615_ /*74306*/;
assign _14621_ = ~D[56] /*74305*/;
assign _14618_ = _13880_ & _14621_ /*74301*/;
assign _14619_ = _13880_ ^ _14621_ /*74304*/;
assign _14620_ = _14612_ & _14619_ /*74302*/;
assign _14329_ = _14612_ ^ _14619_ /*74303*/;
assign _14617_ = _14618_ | _14620_ /*74300*/;
assign _14626_ = ~D[57] /*74299*/;
assign _14623_ = _13881_ & _14626_ /*74295*/;
assign _14624_ = _13881_ ^ _14626_ /*74298*/;
assign _14625_ = _14617_ & _14624_ /*74296*/;
assign _14330_ = _14617_ ^ _14624_ /*74297*/;
assign _14622_ = _14623_ | _14625_ /*74294*/;
assign _14631_ = ~D[58] /*74293*/;
assign _14628_ = _13882_ & _14631_ /*74289*/;
assign _14629_ = _13882_ ^ _14631_ /*74292*/;
assign _14630_ = _14622_ & _14629_ /*74290*/;
assign _14331_ = _14622_ ^ _14629_ /*74291*/;
assign _14627_ = _14628_ | _14630_ /*74288*/;
assign _14636_ = ~D[59] /*74287*/;
assign _14633_ = _13883_ & _14636_ /*74283*/;
assign _14634_ = _13883_ ^ _14636_ /*74286*/;
assign _14635_ = _14627_ & _14634_ /*74284*/;
assign _14332_ = _14627_ ^ _14634_ /*74285*/;
assign _14632_ = _14633_ | _14635_ /*74282*/;
assign _14641_ = ~D[60] /*74281*/;
assign _14638_ = _13884_ & _14641_ /*74277*/;
assign _14639_ = _13884_ ^ _14641_ /*74280*/;
assign _14640_ = _14632_ & _14639_ /*74278*/;
assign _14333_ = _14632_ ^ _14639_ /*74279*/;
assign _14637_ = _14638_ | _14640_ /*74276*/;
assign _14646_ = ~D[61] /*74275*/;
assign _14643_ = _13885_ & _14646_ /*74271*/;
assign _14644_ = _13885_ ^ _14646_ /*74274*/;
assign _14645_ = _14637_ & _14644_ /*74272*/;
assign _14334_ = _14637_ ^ _14644_ /*74273*/;
assign _14642_ = _14643_ | _14645_ /*74270*/;
assign _14651_ = ~D[62] /*74269*/;
assign _14648_ = _13886_ & _14651_ /*74265*/;
assign _14649_ = _13886_ ^ _14651_ /*74268*/;
assign _14650_ = _14642_ & _14649_ /*74266*/;
assign _14335_ = _14642_ ^ _14649_ /*74267*/;
assign _14647_ = _14648_ | _14650_ /*74264*/;
assign _14652_ = _13887_ & oneWire /*74259*/;
assign _14653_ = _13887_ ^ oneWire /*74262*/;
assign _14654_ = _14647_ & _14653_ /*74260*/;
assign _14336_ = _14647_ ^ _14653_ /*74261*/;
assign Q[47] = _14652_ | _14654_ /*74258*/;
assign _14787_ = ~Q[47] /*73873*/;
assign _14786_ = _14787_ & D[0] /*73872*/;
assign _14789_ = _14273_ & _14786_ /*73867*/;
assign _14790_ = _14273_ ^ _14786_ /*73870*/;
assign _14791_ = zeroWire & _14790_ /*73868*/;
assign _14721_ = zeroWire ^ _14790_ /*73869*/;
assign _14788_ = _14789_ | _14791_ /*73866*/;
assign _14793_ = ~Q[47] /*73865*/;
assign _14792_ = _14793_ & D[1] /*73864*/;
assign _14795_ = _14274_ & _14792_ /*73859*/;
assign _14796_ = _14274_ ^ _14792_ /*73862*/;
assign _14797_ = _14788_ & _14796_ /*73860*/;
assign _14722_ = _14788_ ^ _14796_ /*73861*/;
assign _14794_ = _14795_ | _14797_ /*73858*/;
assign _14799_ = ~Q[47] /*73857*/;
assign _14798_ = _14799_ & D[2] /*73856*/;
assign _14801_ = _14275_ & _14798_ /*73851*/;
assign _14802_ = _14275_ ^ _14798_ /*73854*/;
assign _14803_ = _14794_ & _14802_ /*73852*/;
assign _14723_ = _14794_ ^ _14802_ /*73853*/;
assign _14800_ = _14801_ | _14803_ /*73850*/;
assign _14805_ = ~Q[47] /*73849*/;
assign _14804_ = _14805_ & D[3] /*73848*/;
assign _14807_ = _14276_ & _14804_ /*73843*/;
assign _14808_ = _14276_ ^ _14804_ /*73846*/;
assign _14809_ = _14800_ & _14808_ /*73844*/;
assign _14724_ = _14800_ ^ _14808_ /*73845*/;
assign _14806_ = _14807_ | _14809_ /*73842*/;
assign _14811_ = ~Q[47] /*73841*/;
assign _14810_ = _14811_ & D[4] /*73840*/;
assign _14813_ = _14277_ & _14810_ /*73835*/;
assign _14814_ = _14277_ ^ _14810_ /*73838*/;
assign _14815_ = _14806_ & _14814_ /*73836*/;
assign _14725_ = _14806_ ^ _14814_ /*73837*/;
assign _14812_ = _14813_ | _14815_ /*73834*/;
assign _14817_ = ~Q[47] /*73833*/;
assign _14816_ = _14817_ & D[5] /*73832*/;
assign _14819_ = _14278_ & _14816_ /*73827*/;
assign _14820_ = _14278_ ^ _14816_ /*73830*/;
assign _14821_ = _14812_ & _14820_ /*73828*/;
assign _14726_ = _14812_ ^ _14820_ /*73829*/;
assign _14818_ = _14819_ | _14821_ /*73826*/;
assign _14823_ = ~Q[47] /*73825*/;
assign _14822_ = _14823_ & D[6] /*73824*/;
assign _14825_ = _14279_ & _14822_ /*73819*/;
assign _14826_ = _14279_ ^ _14822_ /*73822*/;
assign _14827_ = _14818_ & _14826_ /*73820*/;
assign _14727_ = _14818_ ^ _14826_ /*73821*/;
assign _14824_ = _14825_ | _14827_ /*73818*/;
assign _14829_ = ~Q[47] /*73817*/;
assign _14828_ = _14829_ & D[7] /*73816*/;
assign _14831_ = _14280_ & _14828_ /*73811*/;
assign _14832_ = _14280_ ^ _14828_ /*73814*/;
assign _14833_ = _14824_ & _14832_ /*73812*/;
assign _14728_ = _14824_ ^ _14832_ /*73813*/;
assign _14830_ = _14831_ | _14833_ /*73810*/;
assign _14835_ = ~Q[47] /*73809*/;
assign _14834_ = _14835_ & D[8] /*73808*/;
assign _14837_ = _14281_ & _14834_ /*73803*/;
assign _14838_ = _14281_ ^ _14834_ /*73806*/;
assign _14839_ = _14830_ & _14838_ /*73804*/;
assign _14729_ = _14830_ ^ _14838_ /*73805*/;
assign _14836_ = _14837_ | _14839_ /*73802*/;
assign _14841_ = ~Q[47] /*73801*/;
assign _14840_ = _14841_ & D[9] /*73800*/;
assign _14843_ = _14282_ & _14840_ /*73795*/;
assign _14844_ = _14282_ ^ _14840_ /*73798*/;
assign _14845_ = _14836_ & _14844_ /*73796*/;
assign _14730_ = _14836_ ^ _14844_ /*73797*/;
assign _14842_ = _14843_ | _14845_ /*73794*/;
assign _14847_ = ~Q[47] /*73793*/;
assign _14846_ = _14847_ & D[10] /*73792*/;
assign _14849_ = _14283_ & _14846_ /*73787*/;
assign _14850_ = _14283_ ^ _14846_ /*73790*/;
assign _14851_ = _14842_ & _14850_ /*73788*/;
assign _14731_ = _14842_ ^ _14850_ /*73789*/;
assign _14848_ = _14849_ | _14851_ /*73786*/;
assign _14853_ = ~Q[47] /*73785*/;
assign _14852_ = _14853_ & D[11] /*73784*/;
assign _14855_ = _14284_ & _14852_ /*73779*/;
assign _14856_ = _14284_ ^ _14852_ /*73782*/;
assign _14857_ = _14848_ & _14856_ /*73780*/;
assign _14732_ = _14848_ ^ _14856_ /*73781*/;
assign _14854_ = _14855_ | _14857_ /*73778*/;
assign _14859_ = ~Q[47] /*73777*/;
assign _14858_ = _14859_ & D[12] /*73776*/;
assign _14861_ = _14285_ & _14858_ /*73771*/;
assign _14862_ = _14285_ ^ _14858_ /*73774*/;
assign _14863_ = _14854_ & _14862_ /*73772*/;
assign _14733_ = _14854_ ^ _14862_ /*73773*/;
assign _14860_ = _14861_ | _14863_ /*73770*/;
assign _14865_ = ~Q[47] /*73769*/;
assign _14864_ = _14865_ & D[13] /*73768*/;
assign _14867_ = _14286_ & _14864_ /*73763*/;
assign _14868_ = _14286_ ^ _14864_ /*73766*/;
assign _14869_ = _14860_ & _14868_ /*73764*/;
assign _14734_ = _14860_ ^ _14868_ /*73765*/;
assign _14866_ = _14867_ | _14869_ /*73762*/;
assign _14871_ = ~Q[47] /*73761*/;
assign _14870_ = _14871_ & D[14] /*73760*/;
assign _14873_ = _14287_ & _14870_ /*73755*/;
assign _14874_ = _14287_ ^ _14870_ /*73758*/;
assign _14875_ = _14866_ & _14874_ /*73756*/;
assign _14735_ = _14866_ ^ _14874_ /*73757*/;
assign _14872_ = _14873_ | _14875_ /*73754*/;
assign _14877_ = ~Q[47] /*73753*/;
assign _14876_ = _14877_ & D[15] /*73752*/;
assign _14879_ = _14288_ & _14876_ /*73747*/;
assign _14880_ = _14288_ ^ _14876_ /*73750*/;
assign _14881_ = _14872_ & _14880_ /*73748*/;
assign _14736_ = _14872_ ^ _14880_ /*73749*/;
assign _14878_ = _14879_ | _14881_ /*73746*/;
assign _14883_ = ~Q[47] /*73745*/;
assign _14882_ = _14883_ & D[16] /*73744*/;
assign _14885_ = _14289_ & _14882_ /*73739*/;
assign _14886_ = _14289_ ^ _14882_ /*73742*/;
assign _14887_ = _14878_ & _14886_ /*73740*/;
assign _14737_ = _14878_ ^ _14886_ /*73741*/;
assign _14884_ = _14885_ | _14887_ /*73738*/;
assign _14889_ = ~Q[47] /*73737*/;
assign _14888_ = _14889_ & D[17] /*73736*/;
assign _14891_ = _14290_ & _14888_ /*73731*/;
assign _14892_ = _14290_ ^ _14888_ /*73734*/;
assign _14893_ = _14884_ & _14892_ /*73732*/;
assign _14738_ = _14884_ ^ _14892_ /*73733*/;
assign _14890_ = _14891_ | _14893_ /*73730*/;
assign _14895_ = ~Q[47] /*73729*/;
assign _14894_ = _14895_ & D[18] /*73728*/;
assign _14897_ = _14291_ & _14894_ /*73723*/;
assign _14898_ = _14291_ ^ _14894_ /*73726*/;
assign _14899_ = _14890_ & _14898_ /*73724*/;
assign _14739_ = _14890_ ^ _14898_ /*73725*/;
assign _14896_ = _14897_ | _14899_ /*73722*/;
assign _14901_ = ~Q[47] /*73721*/;
assign _14900_ = _14901_ & D[19] /*73720*/;
assign _14903_ = _14292_ & _14900_ /*73715*/;
assign _14904_ = _14292_ ^ _14900_ /*73718*/;
assign _14905_ = _14896_ & _14904_ /*73716*/;
assign _14740_ = _14896_ ^ _14904_ /*73717*/;
assign _14902_ = _14903_ | _14905_ /*73714*/;
assign _14907_ = ~Q[47] /*73713*/;
assign _14906_ = _14907_ & D[20] /*73712*/;
assign _14909_ = _14293_ & _14906_ /*73707*/;
assign _14910_ = _14293_ ^ _14906_ /*73710*/;
assign _14911_ = _14902_ & _14910_ /*73708*/;
assign _14741_ = _14902_ ^ _14910_ /*73709*/;
assign _14908_ = _14909_ | _14911_ /*73706*/;
assign _14913_ = ~Q[47] /*73705*/;
assign _14912_ = _14913_ & D[21] /*73704*/;
assign _14915_ = _14294_ & _14912_ /*73699*/;
assign _14916_ = _14294_ ^ _14912_ /*73702*/;
assign _14917_ = _14908_ & _14916_ /*73700*/;
assign _14742_ = _14908_ ^ _14916_ /*73701*/;
assign _14914_ = _14915_ | _14917_ /*73698*/;
assign _14919_ = ~Q[47] /*73697*/;
assign _14918_ = _14919_ & D[22] /*73696*/;
assign _14921_ = _14295_ & _14918_ /*73691*/;
assign _14922_ = _14295_ ^ _14918_ /*73694*/;
assign _14923_ = _14914_ & _14922_ /*73692*/;
assign _14743_ = _14914_ ^ _14922_ /*73693*/;
assign _14920_ = _14921_ | _14923_ /*73690*/;
assign _14925_ = ~Q[47] /*73689*/;
assign _14924_ = _14925_ & D[23] /*73688*/;
assign _14927_ = _14296_ & _14924_ /*73683*/;
assign _14928_ = _14296_ ^ _14924_ /*73686*/;
assign _14929_ = _14920_ & _14928_ /*73684*/;
assign _14744_ = _14920_ ^ _14928_ /*73685*/;
assign _14926_ = _14927_ | _14929_ /*73682*/;
assign _14931_ = ~Q[47] /*73681*/;
assign _14930_ = _14931_ & D[24] /*73680*/;
assign _14933_ = _14297_ & _14930_ /*73675*/;
assign _14934_ = _14297_ ^ _14930_ /*73678*/;
assign _14935_ = _14926_ & _14934_ /*73676*/;
assign _14745_ = _14926_ ^ _14934_ /*73677*/;
assign _14932_ = _14933_ | _14935_ /*73674*/;
assign _14937_ = ~Q[47] /*73673*/;
assign _14936_ = _14937_ & D[25] /*73672*/;
assign _14939_ = _14298_ & _14936_ /*73667*/;
assign _14940_ = _14298_ ^ _14936_ /*73670*/;
assign _14941_ = _14932_ & _14940_ /*73668*/;
assign _14746_ = _14932_ ^ _14940_ /*73669*/;
assign _14938_ = _14939_ | _14941_ /*73666*/;
assign _14943_ = ~Q[47] /*73665*/;
assign _14942_ = _14943_ & D[26] /*73664*/;
assign _14945_ = _14299_ & _14942_ /*73659*/;
assign _14946_ = _14299_ ^ _14942_ /*73662*/;
assign _14947_ = _14938_ & _14946_ /*73660*/;
assign _14747_ = _14938_ ^ _14946_ /*73661*/;
assign _14944_ = _14945_ | _14947_ /*73658*/;
assign _14949_ = ~Q[47] /*73657*/;
assign _14948_ = _14949_ & D[27] /*73656*/;
assign _14951_ = _14300_ & _14948_ /*73651*/;
assign _14952_ = _14300_ ^ _14948_ /*73654*/;
assign _14953_ = _14944_ & _14952_ /*73652*/;
assign _14748_ = _14944_ ^ _14952_ /*73653*/;
assign _14950_ = _14951_ | _14953_ /*73650*/;
assign _14955_ = ~Q[47] /*73649*/;
assign _14954_ = _14955_ & D[28] /*73648*/;
assign _14957_ = _14301_ & _14954_ /*73643*/;
assign _14958_ = _14301_ ^ _14954_ /*73646*/;
assign _14959_ = _14950_ & _14958_ /*73644*/;
assign _14749_ = _14950_ ^ _14958_ /*73645*/;
assign _14956_ = _14957_ | _14959_ /*73642*/;
assign _14961_ = ~Q[47] /*73641*/;
assign _14960_ = _14961_ & D[29] /*73640*/;
assign _14963_ = _14302_ & _14960_ /*73635*/;
assign _14964_ = _14302_ ^ _14960_ /*73638*/;
assign _14965_ = _14956_ & _14964_ /*73636*/;
assign _14750_ = _14956_ ^ _14964_ /*73637*/;
assign _14962_ = _14963_ | _14965_ /*73634*/;
assign _14967_ = ~Q[47] /*73633*/;
assign _14966_ = _14967_ & D[30] /*73632*/;
assign _14969_ = _14303_ & _14966_ /*73627*/;
assign _14970_ = _14303_ ^ _14966_ /*73630*/;
assign _14971_ = _14962_ & _14970_ /*73628*/;
assign _14751_ = _14962_ ^ _14970_ /*73629*/;
assign _14968_ = _14969_ | _14971_ /*73626*/;
assign _14973_ = ~Q[47] /*73625*/;
assign _14972_ = _14973_ & D[31] /*73624*/;
assign _14975_ = _14304_ & _14972_ /*73619*/;
assign _14976_ = _14304_ ^ _14972_ /*73622*/;
assign _14977_ = _14968_ & _14976_ /*73620*/;
assign _14752_ = _14968_ ^ _14976_ /*73621*/;
assign _14974_ = _14975_ | _14977_ /*73618*/;
assign _14979_ = ~Q[47] /*73617*/;
assign _14978_ = _14979_ & D[32] /*73616*/;
assign _14981_ = _14305_ & _14978_ /*73611*/;
assign _14982_ = _14305_ ^ _14978_ /*73614*/;
assign _14983_ = _14974_ & _14982_ /*73612*/;
assign _14753_ = _14974_ ^ _14982_ /*73613*/;
assign _14980_ = _14981_ | _14983_ /*73610*/;
assign _14985_ = ~Q[47] /*73609*/;
assign _14984_ = _14985_ & D[33] /*73608*/;
assign _14987_ = _14306_ & _14984_ /*73603*/;
assign _14988_ = _14306_ ^ _14984_ /*73606*/;
assign _14989_ = _14980_ & _14988_ /*73604*/;
assign _14754_ = _14980_ ^ _14988_ /*73605*/;
assign _14986_ = _14987_ | _14989_ /*73602*/;
assign _14991_ = ~Q[47] /*73601*/;
assign _14990_ = _14991_ & D[34] /*73600*/;
assign _14993_ = _14307_ & _14990_ /*73595*/;
assign _14994_ = _14307_ ^ _14990_ /*73598*/;
assign _14995_ = _14986_ & _14994_ /*73596*/;
assign _14755_ = _14986_ ^ _14994_ /*73597*/;
assign _14992_ = _14993_ | _14995_ /*73594*/;
assign _14997_ = ~Q[47] /*73593*/;
assign _14996_ = _14997_ & D[35] /*73592*/;
assign _14999_ = _14308_ & _14996_ /*73587*/;
assign _15000_ = _14308_ ^ _14996_ /*73590*/;
assign _15001_ = _14992_ & _15000_ /*73588*/;
assign _14756_ = _14992_ ^ _15000_ /*73589*/;
assign _14998_ = _14999_ | _15001_ /*73586*/;
assign _15003_ = ~Q[47] /*73585*/;
assign _15002_ = _15003_ & D[36] /*73584*/;
assign _15005_ = _14309_ & _15002_ /*73579*/;
assign _15006_ = _14309_ ^ _15002_ /*73582*/;
assign _15007_ = _14998_ & _15006_ /*73580*/;
assign _14757_ = _14998_ ^ _15006_ /*73581*/;
assign _15004_ = _15005_ | _15007_ /*73578*/;
assign _15009_ = ~Q[47] /*73577*/;
assign _15008_ = _15009_ & D[37] /*73576*/;
assign _15011_ = _14310_ & _15008_ /*73571*/;
assign _15012_ = _14310_ ^ _15008_ /*73574*/;
assign _15013_ = _15004_ & _15012_ /*73572*/;
assign _14758_ = _15004_ ^ _15012_ /*73573*/;
assign _15010_ = _15011_ | _15013_ /*73570*/;
assign _15015_ = ~Q[47] /*73569*/;
assign _15014_ = _15015_ & D[38] /*73568*/;
assign _15017_ = _14311_ & _15014_ /*73563*/;
assign _15018_ = _14311_ ^ _15014_ /*73566*/;
assign _15019_ = _15010_ & _15018_ /*73564*/;
assign _14759_ = _15010_ ^ _15018_ /*73565*/;
assign _15016_ = _15017_ | _15019_ /*73562*/;
assign _15021_ = ~Q[47] /*73561*/;
assign _15020_ = _15021_ & D[39] /*73560*/;
assign _15023_ = _14312_ & _15020_ /*73555*/;
assign _15024_ = _14312_ ^ _15020_ /*73558*/;
assign _15025_ = _15016_ & _15024_ /*73556*/;
assign _14760_ = _15016_ ^ _15024_ /*73557*/;
assign _15022_ = _15023_ | _15025_ /*73554*/;
assign _15027_ = ~Q[47] /*73553*/;
assign _15026_ = _15027_ & D[40] /*73552*/;
assign _15029_ = _14313_ & _15026_ /*73547*/;
assign _15030_ = _14313_ ^ _15026_ /*73550*/;
assign _15031_ = _15022_ & _15030_ /*73548*/;
assign _14761_ = _15022_ ^ _15030_ /*73549*/;
assign _15028_ = _15029_ | _15031_ /*73546*/;
assign _15033_ = ~Q[47] /*73545*/;
assign _15032_ = _15033_ & D[41] /*73544*/;
assign _15035_ = _14314_ & _15032_ /*73539*/;
assign _15036_ = _14314_ ^ _15032_ /*73542*/;
assign _15037_ = _15028_ & _15036_ /*73540*/;
assign _14762_ = _15028_ ^ _15036_ /*73541*/;
assign _15034_ = _15035_ | _15037_ /*73538*/;
assign _15039_ = ~Q[47] /*73537*/;
assign _15038_ = _15039_ & D[42] /*73536*/;
assign _15041_ = _14315_ & _15038_ /*73531*/;
assign _15042_ = _14315_ ^ _15038_ /*73534*/;
assign _15043_ = _15034_ & _15042_ /*73532*/;
assign _14763_ = _15034_ ^ _15042_ /*73533*/;
assign _15040_ = _15041_ | _15043_ /*73530*/;
assign _15045_ = ~Q[47] /*73529*/;
assign _15044_ = _15045_ & D[43] /*73528*/;
assign _15047_ = _14316_ & _15044_ /*73523*/;
assign _15048_ = _14316_ ^ _15044_ /*73526*/;
assign _15049_ = _15040_ & _15048_ /*73524*/;
assign _14764_ = _15040_ ^ _15048_ /*73525*/;
assign _15046_ = _15047_ | _15049_ /*73522*/;
assign _15051_ = ~Q[47] /*73521*/;
assign _15050_ = _15051_ & D[44] /*73520*/;
assign _15053_ = _14317_ & _15050_ /*73515*/;
assign _15054_ = _14317_ ^ _15050_ /*73518*/;
assign _15055_ = _15046_ & _15054_ /*73516*/;
assign _14765_ = _15046_ ^ _15054_ /*73517*/;
assign _15052_ = _15053_ | _15055_ /*73514*/;
assign _15057_ = ~Q[47] /*73513*/;
assign _15056_ = _15057_ & D[45] /*73512*/;
assign _15059_ = _14318_ & _15056_ /*73507*/;
assign _15060_ = _14318_ ^ _15056_ /*73510*/;
assign _15061_ = _15052_ & _15060_ /*73508*/;
assign _14766_ = _15052_ ^ _15060_ /*73509*/;
assign _15058_ = _15059_ | _15061_ /*73506*/;
assign _15063_ = ~Q[47] /*73505*/;
assign _15062_ = _15063_ & D[46] /*73504*/;
assign _15065_ = _14319_ & _15062_ /*73499*/;
assign _15066_ = _14319_ ^ _15062_ /*73502*/;
assign _15067_ = _15058_ & _15066_ /*73500*/;
assign _14767_ = _15058_ ^ _15066_ /*73501*/;
assign _15064_ = _15065_ | _15067_ /*73498*/;
assign _15069_ = ~Q[47] /*73497*/;
assign _15068_ = _15069_ & D[47] /*73496*/;
assign _15071_ = _14320_ & _15068_ /*73491*/;
assign _15072_ = _14320_ ^ _15068_ /*73494*/;
assign _15073_ = _15064_ & _15072_ /*73492*/;
assign _14768_ = _15064_ ^ _15072_ /*73493*/;
assign _15070_ = _15071_ | _15073_ /*73490*/;
assign _15075_ = ~Q[47] /*73489*/;
assign _15074_ = _15075_ & D[48] /*73488*/;
assign _15077_ = _14321_ & _15074_ /*73483*/;
assign _15078_ = _14321_ ^ _15074_ /*73486*/;
assign _15079_ = _15070_ & _15078_ /*73484*/;
assign _14769_ = _15070_ ^ _15078_ /*73485*/;
assign _15076_ = _15077_ | _15079_ /*73482*/;
assign _15081_ = ~Q[47] /*73481*/;
assign _15080_ = _15081_ & D[49] /*73480*/;
assign _15083_ = _14322_ & _15080_ /*73475*/;
assign _15084_ = _14322_ ^ _15080_ /*73478*/;
assign _15085_ = _15076_ & _15084_ /*73476*/;
assign _14770_ = _15076_ ^ _15084_ /*73477*/;
assign _15082_ = _15083_ | _15085_ /*73474*/;
assign _15087_ = ~Q[47] /*73473*/;
assign _15086_ = _15087_ & D[50] /*73472*/;
assign _15089_ = _14323_ & _15086_ /*73467*/;
assign _15090_ = _14323_ ^ _15086_ /*73470*/;
assign _15091_ = _15082_ & _15090_ /*73468*/;
assign _14771_ = _15082_ ^ _15090_ /*73469*/;
assign _15088_ = _15089_ | _15091_ /*73466*/;
assign _15093_ = ~Q[47] /*73465*/;
assign _15092_ = _15093_ & D[51] /*73464*/;
assign _15095_ = _14324_ & _15092_ /*73459*/;
assign _15096_ = _14324_ ^ _15092_ /*73462*/;
assign _15097_ = _15088_ & _15096_ /*73460*/;
assign _14772_ = _15088_ ^ _15096_ /*73461*/;
assign _15094_ = _15095_ | _15097_ /*73458*/;
assign _15099_ = ~Q[47] /*73457*/;
assign _15098_ = _15099_ & D[52] /*73456*/;
assign _15101_ = _14325_ & _15098_ /*73451*/;
assign _15102_ = _14325_ ^ _15098_ /*73454*/;
assign _15103_ = _15094_ & _15102_ /*73452*/;
assign _14773_ = _15094_ ^ _15102_ /*73453*/;
assign _15100_ = _15101_ | _15103_ /*73450*/;
assign _15105_ = ~Q[47] /*73449*/;
assign _15104_ = _15105_ & D[53] /*73448*/;
assign _15107_ = _14326_ & _15104_ /*73443*/;
assign _15108_ = _14326_ ^ _15104_ /*73446*/;
assign _15109_ = _15100_ & _15108_ /*73444*/;
assign _14774_ = _15100_ ^ _15108_ /*73445*/;
assign _15106_ = _15107_ | _15109_ /*73442*/;
assign _15111_ = ~Q[47] /*73441*/;
assign _15110_ = _15111_ & D[54] /*73440*/;
assign _15113_ = _14327_ & _15110_ /*73435*/;
assign _15114_ = _14327_ ^ _15110_ /*73438*/;
assign _15115_ = _15106_ & _15114_ /*73436*/;
assign _14775_ = _15106_ ^ _15114_ /*73437*/;
assign _15112_ = _15113_ | _15115_ /*73434*/;
assign _15117_ = ~Q[47] /*73433*/;
assign _15116_ = _15117_ & D[55] /*73432*/;
assign _15119_ = _14328_ & _15116_ /*73427*/;
assign _15120_ = _14328_ ^ _15116_ /*73430*/;
assign _15121_ = _15112_ & _15120_ /*73428*/;
assign _14776_ = _15112_ ^ _15120_ /*73429*/;
assign _15118_ = _15119_ | _15121_ /*73426*/;
assign _15123_ = ~Q[47] /*73425*/;
assign _15122_ = _15123_ & D[56] /*73424*/;
assign _15125_ = _14329_ & _15122_ /*73419*/;
assign _15126_ = _14329_ ^ _15122_ /*73422*/;
assign _15127_ = _15118_ & _15126_ /*73420*/;
assign _14777_ = _15118_ ^ _15126_ /*73421*/;
assign _15124_ = _15125_ | _15127_ /*73418*/;
assign _15129_ = ~Q[47] /*73417*/;
assign _15128_ = _15129_ & D[57] /*73416*/;
assign _15131_ = _14330_ & _15128_ /*73411*/;
assign _15132_ = _14330_ ^ _15128_ /*73414*/;
assign _15133_ = _15124_ & _15132_ /*73412*/;
assign _14778_ = _15124_ ^ _15132_ /*73413*/;
assign _15130_ = _15131_ | _15133_ /*73410*/;
assign _15135_ = ~Q[47] /*73409*/;
assign _15134_ = _15135_ & D[58] /*73408*/;
assign _15137_ = _14331_ & _15134_ /*73403*/;
assign _15138_ = _14331_ ^ _15134_ /*73406*/;
assign _15139_ = _15130_ & _15138_ /*73404*/;
assign _14779_ = _15130_ ^ _15138_ /*73405*/;
assign _15136_ = _15137_ | _15139_ /*73402*/;
assign _15141_ = ~Q[47] /*73401*/;
assign _15140_ = _15141_ & D[59] /*73400*/;
assign _15143_ = _14332_ & _15140_ /*73395*/;
assign _15144_ = _14332_ ^ _15140_ /*73398*/;
assign _15145_ = _15136_ & _15144_ /*73396*/;
assign _14780_ = _15136_ ^ _15144_ /*73397*/;
assign _15142_ = _15143_ | _15145_ /*73394*/;
assign _15147_ = ~Q[47] /*73393*/;
assign _15146_ = _15147_ & D[60] /*73392*/;
assign _15149_ = _14333_ & _15146_ /*73387*/;
assign _15150_ = _14333_ ^ _15146_ /*73390*/;
assign _15151_ = _15142_ & _15150_ /*73388*/;
assign _14781_ = _15142_ ^ _15150_ /*73389*/;
assign _15148_ = _15149_ | _15151_ /*73386*/;
assign _15153_ = ~Q[47] /*73385*/;
assign _15152_ = _15153_ & D[61] /*73384*/;
assign _15155_ = _14334_ & _15152_ /*73379*/;
assign _15156_ = _14334_ ^ _15152_ /*73382*/;
assign _15157_ = _15148_ & _15156_ /*73380*/;
assign _14782_ = _15148_ ^ _15156_ /*73381*/;
assign _15154_ = _15155_ | _15157_ /*73378*/;
assign _15159_ = ~Q[47] /*73377*/;
assign _15158_ = _15159_ & D[62] /*73376*/;
assign _15161_ = _14335_ & _15158_ /*73371*/;
assign _15162_ = _14335_ ^ _15158_ /*73374*/;
assign _15163_ = _15154_ & _15162_ /*73372*/;
assign _14783_ = _15154_ ^ _15162_ /*73373*/;
assign _15160_ = _15161_ | _15163_ /*73370*/;
assign _15165_ = ~Q[47] /*73369*/;
assign _15164_ = _15165_ & zeroWire /*73368*/;
assign _15166_ = _14336_ ^ _15164_ /*73366*/;
assign _14784_ = _15166_ ^ _15160_ /*73365*/;
assign _15237_ = ~D[0] /*73111*/;
assign _15234_ = R_0[46] & _15237_ /*73107*/;
assign _15235_ = R_0[46] ^ _15237_ /*73110*/;
assign _15236_ = oneWire & _15235_ /*73108*/;
assign _15169_ = oneWire ^ _15235_ /*73109*/;
assign _15233_ = _15234_ | _15236_ /*73106*/;
assign _15242_ = ~D[1] /*73105*/;
assign _15239_ = _14721_ & _15242_ /*73101*/;
assign _15240_ = _14721_ ^ _15242_ /*73104*/;
assign _15241_ = _15233_ & _15240_ /*73102*/;
assign _15170_ = _15233_ ^ _15240_ /*73103*/;
assign _15238_ = _15239_ | _15241_ /*73100*/;
assign _15247_ = ~D[2] /*73099*/;
assign _15244_ = _14722_ & _15247_ /*73095*/;
assign _15245_ = _14722_ ^ _15247_ /*73098*/;
assign _15246_ = _15238_ & _15245_ /*73096*/;
assign _15171_ = _15238_ ^ _15245_ /*73097*/;
assign _15243_ = _15244_ | _15246_ /*73094*/;
assign _15252_ = ~D[3] /*73093*/;
assign _15249_ = _14723_ & _15252_ /*73089*/;
assign _15250_ = _14723_ ^ _15252_ /*73092*/;
assign _15251_ = _15243_ & _15250_ /*73090*/;
assign _15172_ = _15243_ ^ _15250_ /*73091*/;
assign _15248_ = _15249_ | _15251_ /*73088*/;
assign _15257_ = ~D[4] /*73087*/;
assign _15254_ = _14724_ & _15257_ /*73083*/;
assign _15255_ = _14724_ ^ _15257_ /*73086*/;
assign _15256_ = _15248_ & _15255_ /*73084*/;
assign _15173_ = _15248_ ^ _15255_ /*73085*/;
assign _15253_ = _15254_ | _15256_ /*73082*/;
assign _15262_ = ~D[5] /*73081*/;
assign _15259_ = _14725_ & _15262_ /*73077*/;
assign _15260_ = _14725_ ^ _15262_ /*73080*/;
assign _15261_ = _15253_ & _15260_ /*73078*/;
assign _15174_ = _15253_ ^ _15260_ /*73079*/;
assign _15258_ = _15259_ | _15261_ /*73076*/;
assign _15267_ = ~D[6] /*73075*/;
assign _15264_ = _14726_ & _15267_ /*73071*/;
assign _15265_ = _14726_ ^ _15267_ /*73074*/;
assign _15266_ = _15258_ & _15265_ /*73072*/;
assign _15175_ = _15258_ ^ _15265_ /*73073*/;
assign _15263_ = _15264_ | _15266_ /*73070*/;
assign _15272_ = ~D[7] /*73069*/;
assign _15269_ = _14727_ & _15272_ /*73065*/;
assign _15270_ = _14727_ ^ _15272_ /*73068*/;
assign _15271_ = _15263_ & _15270_ /*73066*/;
assign _15176_ = _15263_ ^ _15270_ /*73067*/;
assign _15268_ = _15269_ | _15271_ /*73064*/;
assign _15277_ = ~D[8] /*73063*/;
assign _15274_ = _14728_ & _15277_ /*73059*/;
assign _15275_ = _14728_ ^ _15277_ /*73062*/;
assign _15276_ = _15268_ & _15275_ /*73060*/;
assign _15177_ = _15268_ ^ _15275_ /*73061*/;
assign _15273_ = _15274_ | _15276_ /*73058*/;
assign _15282_ = ~D[9] /*73057*/;
assign _15279_ = _14729_ & _15282_ /*73053*/;
assign _15280_ = _14729_ ^ _15282_ /*73056*/;
assign _15281_ = _15273_ & _15280_ /*73054*/;
assign _15178_ = _15273_ ^ _15280_ /*73055*/;
assign _15278_ = _15279_ | _15281_ /*73052*/;
assign _15287_ = ~D[10] /*73051*/;
assign _15284_ = _14730_ & _15287_ /*73047*/;
assign _15285_ = _14730_ ^ _15287_ /*73050*/;
assign _15286_ = _15278_ & _15285_ /*73048*/;
assign _15179_ = _15278_ ^ _15285_ /*73049*/;
assign _15283_ = _15284_ | _15286_ /*73046*/;
assign _15292_ = ~D[11] /*73045*/;
assign _15289_ = _14731_ & _15292_ /*73041*/;
assign _15290_ = _14731_ ^ _15292_ /*73044*/;
assign _15291_ = _15283_ & _15290_ /*73042*/;
assign _15180_ = _15283_ ^ _15290_ /*73043*/;
assign _15288_ = _15289_ | _15291_ /*73040*/;
assign _15297_ = ~D[12] /*73039*/;
assign _15294_ = _14732_ & _15297_ /*73035*/;
assign _15295_ = _14732_ ^ _15297_ /*73038*/;
assign _15296_ = _15288_ & _15295_ /*73036*/;
assign _15181_ = _15288_ ^ _15295_ /*73037*/;
assign _15293_ = _15294_ | _15296_ /*73034*/;
assign _15302_ = ~D[13] /*73033*/;
assign _15299_ = _14733_ & _15302_ /*73029*/;
assign _15300_ = _14733_ ^ _15302_ /*73032*/;
assign _15301_ = _15293_ & _15300_ /*73030*/;
assign _15182_ = _15293_ ^ _15300_ /*73031*/;
assign _15298_ = _15299_ | _15301_ /*73028*/;
assign _15307_ = ~D[14] /*73027*/;
assign _15304_ = _14734_ & _15307_ /*73023*/;
assign _15305_ = _14734_ ^ _15307_ /*73026*/;
assign _15306_ = _15298_ & _15305_ /*73024*/;
assign _15183_ = _15298_ ^ _15305_ /*73025*/;
assign _15303_ = _15304_ | _15306_ /*73022*/;
assign _15312_ = ~D[15] /*73021*/;
assign _15309_ = _14735_ & _15312_ /*73017*/;
assign _15310_ = _14735_ ^ _15312_ /*73020*/;
assign _15311_ = _15303_ & _15310_ /*73018*/;
assign _15184_ = _15303_ ^ _15310_ /*73019*/;
assign _15308_ = _15309_ | _15311_ /*73016*/;
assign _15317_ = ~D[16] /*73015*/;
assign _15314_ = _14736_ & _15317_ /*73011*/;
assign _15315_ = _14736_ ^ _15317_ /*73014*/;
assign _15316_ = _15308_ & _15315_ /*73012*/;
assign _15185_ = _15308_ ^ _15315_ /*73013*/;
assign _15313_ = _15314_ | _15316_ /*73010*/;
assign _15322_ = ~D[17] /*73009*/;
assign _15319_ = _14737_ & _15322_ /*73005*/;
assign _15320_ = _14737_ ^ _15322_ /*73008*/;
assign _15321_ = _15313_ & _15320_ /*73006*/;
assign _15186_ = _15313_ ^ _15320_ /*73007*/;
assign _15318_ = _15319_ | _15321_ /*73004*/;
assign _15327_ = ~D[18] /*73003*/;
assign _15324_ = _14738_ & _15327_ /*72999*/;
assign _15325_ = _14738_ ^ _15327_ /*73002*/;
assign _15326_ = _15318_ & _15325_ /*73000*/;
assign _15187_ = _15318_ ^ _15325_ /*73001*/;
assign _15323_ = _15324_ | _15326_ /*72998*/;
assign _15332_ = ~D[19] /*72997*/;
assign _15329_ = _14739_ & _15332_ /*72993*/;
assign _15330_ = _14739_ ^ _15332_ /*72996*/;
assign _15331_ = _15323_ & _15330_ /*72994*/;
assign _15188_ = _15323_ ^ _15330_ /*72995*/;
assign _15328_ = _15329_ | _15331_ /*72992*/;
assign _15337_ = ~D[20] /*72991*/;
assign _15334_ = _14740_ & _15337_ /*72987*/;
assign _15335_ = _14740_ ^ _15337_ /*72990*/;
assign _15336_ = _15328_ & _15335_ /*72988*/;
assign _15189_ = _15328_ ^ _15335_ /*72989*/;
assign _15333_ = _15334_ | _15336_ /*72986*/;
assign _15342_ = ~D[21] /*72985*/;
assign _15339_ = _14741_ & _15342_ /*72981*/;
assign _15340_ = _14741_ ^ _15342_ /*72984*/;
assign _15341_ = _15333_ & _15340_ /*72982*/;
assign _15190_ = _15333_ ^ _15340_ /*72983*/;
assign _15338_ = _15339_ | _15341_ /*72980*/;
assign _15347_ = ~D[22] /*72979*/;
assign _15344_ = _14742_ & _15347_ /*72975*/;
assign _15345_ = _14742_ ^ _15347_ /*72978*/;
assign _15346_ = _15338_ & _15345_ /*72976*/;
assign _15191_ = _15338_ ^ _15345_ /*72977*/;
assign _15343_ = _15344_ | _15346_ /*72974*/;
assign _15352_ = ~D[23] /*72973*/;
assign _15349_ = _14743_ & _15352_ /*72969*/;
assign _15350_ = _14743_ ^ _15352_ /*72972*/;
assign _15351_ = _15343_ & _15350_ /*72970*/;
assign _15192_ = _15343_ ^ _15350_ /*72971*/;
assign _15348_ = _15349_ | _15351_ /*72968*/;
assign _15357_ = ~D[24] /*72967*/;
assign _15354_ = _14744_ & _15357_ /*72963*/;
assign _15355_ = _14744_ ^ _15357_ /*72966*/;
assign _15356_ = _15348_ & _15355_ /*72964*/;
assign _15193_ = _15348_ ^ _15355_ /*72965*/;
assign _15353_ = _15354_ | _15356_ /*72962*/;
assign _15362_ = ~D[25] /*72961*/;
assign _15359_ = _14745_ & _15362_ /*72957*/;
assign _15360_ = _14745_ ^ _15362_ /*72960*/;
assign _15361_ = _15353_ & _15360_ /*72958*/;
assign _15194_ = _15353_ ^ _15360_ /*72959*/;
assign _15358_ = _15359_ | _15361_ /*72956*/;
assign _15367_ = ~D[26] /*72955*/;
assign _15364_ = _14746_ & _15367_ /*72951*/;
assign _15365_ = _14746_ ^ _15367_ /*72954*/;
assign _15366_ = _15358_ & _15365_ /*72952*/;
assign _15195_ = _15358_ ^ _15365_ /*72953*/;
assign _15363_ = _15364_ | _15366_ /*72950*/;
assign _15372_ = ~D[27] /*72949*/;
assign _15369_ = _14747_ & _15372_ /*72945*/;
assign _15370_ = _14747_ ^ _15372_ /*72948*/;
assign _15371_ = _15363_ & _15370_ /*72946*/;
assign _15196_ = _15363_ ^ _15370_ /*72947*/;
assign _15368_ = _15369_ | _15371_ /*72944*/;
assign _15377_ = ~D[28] /*72943*/;
assign _15374_ = _14748_ & _15377_ /*72939*/;
assign _15375_ = _14748_ ^ _15377_ /*72942*/;
assign _15376_ = _15368_ & _15375_ /*72940*/;
assign _15197_ = _15368_ ^ _15375_ /*72941*/;
assign _15373_ = _15374_ | _15376_ /*72938*/;
assign _15382_ = ~D[29] /*72937*/;
assign _15379_ = _14749_ & _15382_ /*72933*/;
assign _15380_ = _14749_ ^ _15382_ /*72936*/;
assign _15381_ = _15373_ & _15380_ /*72934*/;
assign _15198_ = _15373_ ^ _15380_ /*72935*/;
assign _15378_ = _15379_ | _15381_ /*72932*/;
assign _15387_ = ~D[30] /*72931*/;
assign _15384_ = _14750_ & _15387_ /*72927*/;
assign _15385_ = _14750_ ^ _15387_ /*72930*/;
assign _15386_ = _15378_ & _15385_ /*72928*/;
assign _15199_ = _15378_ ^ _15385_ /*72929*/;
assign _15383_ = _15384_ | _15386_ /*72926*/;
assign _15392_ = ~D[31] /*72925*/;
assign _15389_ = _14751_ & _15392_ /*72921*/;
assign _15390_ = _14751_ ^ _15392_ /*72924*/;
assign _15391_ = _15383_ & _15390_ /*72922*/;
assign _15200_ = _15383_ ^ _15390_ /*72923*/;
assign _15388_ = _15389_ | _15391_ /*72920*/;
assign _15397_ = ~D[32] /*72919*/;
assign _15394_ = _14752_ & _15397_ /*72915*/;
assign _15395_ = _14752_ ^ _15397_ /*72918*/;
assign _15396_ = _15388_ & _15395_ /*72916*/;
assign _15201_ = _15388_ ^ _15395_ /*72917*/;
assign _15393_ = _15394_ | _15396_ /*72914*/;
assign _15402_ = ~D[33] /*72913*/;
assign _15399_ = _14753_ & _15402_ /*72909*/;
assign _15400_ = _14753_ ^ _15402_ /*72912*/;
assign _15401_ = _15393_ & _15400_ /*72910*/;
assign _15202_ = _15393_ ^ _15400_ /*72911*/;
assign _15398_ = _15399_ | _15401_ /*72908*/;
assign _15407_ = ~D[34] /*72907*/;
assign _15404_ = _14754_ & _15407_ /*72903*/;
assign _15405_ = _14754_ ^ _15407_ /*72906*/;
assign _15406_ = _15398_ & _15405_ /*72904*/;
assign _15203_ = _15398_ ^ _15405_ /*72905*/;
assign _15403_ = _15404_ | _15406_ /*72902*/;
assign _15412_ = ~D[35] /*72901*/;
assign _15409_ = _14755_ & _15412_ /*72897*/;
assign _15410_ = _14755_ ^ _15412_ /*72900*/;
assign _15411_ = _15403_ & _15410_ /*72898*/;
assign _15204_ = _15403_ ^ _15410_ /*72899*/;
assign _15408_ = _15409_ | _15411_ /*72896*/;
assign _15417_ = ~D[36] /*72895*/;
assign _15414_ = _14756_ & _15417_ /*72891*/;
assign _15415_ = _14756_ ^ _15417_ /*72894*/;
assign _15416_ = _15408_ & _15415_ /*72892*/;
assign _15205_ = _15408_ ^ _15415_ /*72893*/;
assign _15413_ = _15414_ | _15416_ /*72890*/;
assign _15422_ = ~D[37] /*72889*/;
assign _15419_ = _14757_ & _15422_ /*72885*/;
assign _15420_ = _14757_ ^ _15422_ /*72888*/;
assign _15421_ = _15413_ & _15420_ /*72886*/;
assign _15206_ = _15413_ ^ _15420_ /*72887*/;
assign _15418_ = _15419_ | _15421_ /*72884*/;
assign _15427_ = ~D[38] /*72883*/;
assign _15424_ = _14758_ & _15427_ /*72879*/;
assign _15425_ = _14758_ ^ _15427_ /*72882*/;
assign _15426_ = _15418_ & _15425_ /*72880*/;
assign _15207_ = _15418_ ^ _15425_ /*72881*/;
assign _15423_ = _15424_ | _15426_ /*72878*/;
assign _15432_ = ~D[39] /*72877*/;
assign _15429_ = _14759_ & _15432_ /*72873*/;
assign _15430_ = _14759_ ^ _15432_ /*72876*/;
assign _15431_ = _15423_ & _15430_ /*72874*/;
assign _15208_ = _15423_ ^ _15430_ /*72875*/;
assign _15428_ = _15429_ | _15431_ /*72872*/;
assign _15437_ = ~D[40] /*72871*/;
assign _15434_ = _14760_ & _15437_ /*72867*/;
assign _15435_ = _14760_ ^ _15437_ /*72870*/;
assign _15436_ = _15428_ & _15435_ /*72868*/;
assign _15209_ = _15428_ ^ _15435_ /*72869*/;
assign _15433_ = _15434_ | _15436_ /*72866*/;
assign _15442_ = ~D[41] /*72865*/;
assign _15439_ = _14761_ & _15442_ /*72861*/;
assign _15440_ = _14761_ ^ _15442_ /*72864*/;
assign _15441_ = _15433_ & _15440_ /*72862*/;
assign _15210_ = _15433_ ^ _15440_ /*72863*/;
assign _15438_ = _15439_ | _15441_ /*72860*/;
assign _15447_ = ~D[42] /*72859*/;
assign _15444_ = _14762_ & _15447_ /*72855*/;
assign _15445_ = _14762_ ^ _15447_ /*72858*/;
assign _15446_ = _15438_ & _15445_ /*72856*/;
assign _15211_ = _15438_ ^ _15445_ /*72857*/;
assign _15443_ = _15444_ | _15446_ /*72854*/;
assign _15452_ = ~D[43] /*72853*/;
assign _15449_ = _14763_ & _15452_ /*72849*/;
assign _15450_ = _14763_ ^ _15452_ /*72852*/;
assign _15451_ = _15443_ & _15450_ /*72850*/;
assign _15212_ = _15443_ ^ _15450_ /*72851*/;
assign _15448_ = _15449_ | _15451_ /*72848*/;
assign _15457_ = ~D[44] /*72847*/;
assign _15454_ = _14764_ & _15457_ /*72843*/;
assign _15455_ = _14764_ ^ _15457_ /*72846*/;
assign _15456_ = _15448_ & _15455_ /*72844*/;
assign _15213_ = _15448_ ^ _15455_ /*72845*/;
assign _15453_ = _15454_ | _15456_ /*72842*/;
assign _15462_ = ~D[45] /*72841*/;
assign _15459_ = _14765_ & _15462_ /*72837*/;
assign _15460_ = _14765_ ^ _15462_ /*72840*/;
assign _15461_ = _15453_ & _15460_ /*72838*/;
assign _15214_ = _15453_ ^ _15460_ /*72839*/;
assign _15458_ = _15459_ | _15461_ /*72836*/;
assign _15467_ = ~D[46] /*72835*/;
assign _15464_ = _14766_ & _15467_ /*72831*/;
assign _15465_ = _14766_ ^ _15467_ /*72834*/;
assign _15466_ = _15458_ & _15465_ /*72832*/;
assign _15215_ = _15458_ ^ _15465_ /*72833*/;
assign _15463_ = _15464_ | _15466_ /*72830*/;
assign _15472_ = ~D[47] /*72829*/;
assign _15469_ = _14767_ & _15472_ /*72825*/;
assign _15470_ = _14767_ ^ _15472_ /*72828*/;
assign _15471_ = _15463_ & _15470_ /*72826*/;
assign _15216_ = _15463_ ^ _15470_ /*72827*/;
assign _15468_ = _15469_ | _15471_ /*72824*/;
assign _15477_ = ~D[48] /*72823*/;
assign _15474_ = _14768_ & _15477_ /*72819*/;
assign _15475_ = _14768_ ^ _15477_ /*72822*/;
assign _15476_ = _15468_ & _15475_ /*72820*/;
assign _15217_ = _15468_ ^ _15475_ /*72821*/;
assign _15473_ = _15474_ | _15476_ /*72818*/;
assign _15482_ = ~D[49] /*72817*/;
assign _15479_ = _14769_ & _15482_ /*72813*/;
assign _15480_ = _14769_ ^ _15482_ /*72816*/;
assign _15481_ = _15473_ & _15480_ /*72814*/;
assign _15218_ = _15473_ ^ _15480_ /*72815*/;
assign _15478_ = _15479_ | _15481_ /*72812*/;
assign _15487_ = ~D[50] /*72811*/;
assign _15484_ = _14770_ & _15487_ /*72807*/;
assign _15485_ = _14770_ ^ _15487_ /*72810*/;
assign _15486_ = _15478_ & _15485_ /*72808*/;
assign _15219_ = _15478_ ^ _15485_ /*72809*/;
assign _15483_ = _15484_ | _15486_ /*72806*/;
assign _15492_ = ~D[51] /*72805*/;
assign _15489_ = _14771_ & _15492_ /*72801*/;
assign _15490_ = _14771_ ^ _15492_ /*72804*/;
assign _15491_ = _15483_ & _15490_ /*72802*/;
assign _15220_ = _15483_ ^ _15490_ /*72803*/;
assign _15488_ = _15489_ | _15491_ /*72800*/;
assign _15497_ = ~D[52] /*72799*/;
assign _15494_ = _14772_ & _15497_ /*72795*/;
assign _15495_ = _14772_ ^ _15497_ /*72798*/;
assign _15496_ = _15488_ & _15495_ /*72796*/;
assign _15221_ = _15488_ ^ _15495_ /*72797*/;
assign _15493_ = _15494_ | _15496_ /*72794*/;
assign _15502_ = ~D[53] /*72793*/;
assign _15499_ = _14773_ & _15502_ /*72789*/;
assign _15500_ = _14773_ ^ _15502_ /*72792*/;
assign _15501_ = _15493_ & _15500_ /*72790*/;
assign _15222_ = _15493_ ^ _15500_ /*72791*/;
assign _15498_ = _15499_ | _15501_ /*72788*/;
assign _15507_ = ~D[54] /*72787*/;
assign _15504_ = _14774_ & _15507_ /*72783*/;
assign _15505_ = _14774_ ^ _15507_ /*72786*/;
assign _15506_ = _15498_ & _15505_ /*72784*/;
assign _15223_ = _15498_ ^ _15505_ /*72785*/;
assign _15503_ = _15504_ | _15506_ /*72782*/;
assign _15512_ = ~D[55] /*72781*/;
assign _15509_ = _14775_ & _15512_ /*72777*/;
assign _15510_ = _14775_ ^ _15512_ /*72780*/;
assign _15511_ = _15503_ & _15510_ /*72778*/;
assign _15224_ = _15503_ ^ _15510_ /*72779*/;
assign _15508_ = _15509_ | _15511_ /*72776*/;
assign _15517_ = ~D[56] /*72775*/;
assign _15514_ = _14776_ & _15517_ /*72771*/;
assign _15515_ = _14776_ ^ _15517_ /*72774*/;
assign _15516_ = _15508_ & _15515_ /*72772*/;
assign _15225_ = _15508_ ^ _15515_ /*72773*/;
assign _15513_ = _15514_ | _15516_ /*72770*/;
assign _15522_ = ~D[57] /*72769*/;
assign _15519_ = _14777_ & _15522_ /*72765*/;
assign _15520_ = _14777_ ^ _15522_ /*72768*/;
assign _15521_ = _15513_ & _15520_ /*72766*/;
assign _15226_ = _15513_ ^ _15520_ /*72767*/;
assign _15518_ = _15519_ | _15521_ /*72764*/;
assign _15527_ = ~D[58] /*72763*/;
assign _15524_ = _14778_ & _15527_ /*72759*/;
assign _15525_ = _14778_ ^ _15527_ /*72762*/;
assign _15526_ = _15518_ & _15525_ /*72760*/;
assign _15227_ = _15518_ ^ _15525_ /*72761*/;
assign _15523_ = _15524_ | _15526_ /*72758*/;
assign _15532_ = ~D[59] /*72757*/;
assign _15529_ = _14779_ & _15532_ /*72753*/;
assign _15530_ = _14779_ ^ _15532_ /*72756*/;
assign _15531_ = _15523_ & _15530_ /*72754*/;
assign _15228_ = _15523_ ^ _15530_ /*72755*/;
assign _15528_ = _15529_ | _15531_ /*72752*/;
assign _15537_ = ~D[60] /*72751*/;
assign _15534_ = _14780_ & _15537_ /*72747*/;
assign _15535_ = _14780_ ^ _15537_ /*72750*/;
assign _15536_ = _15528_ & _15535_ /*72748*/;
assign _15229_ = _15528_ ^ _15535_ /*72749*/;
assign _15533_ = _15534_ | _15536_ /*72746*/;
assign _15542_ = ~D[61] /*72745*/;
assign _15539_ = _14781_ & _15542_ /*72741*/;
assign _15540_ = _14781_ ^ _15542_ /*72744*/;
assign _15541_ = _15533_ & _15540_ /*72742*/;
assign _15230_ = _15533_ ^ _15540_ /*72743*/;
assign _15538_ = _15539_ | _15541_ /*72740*/;
assign _15547_ = ~D[62] /*72739*/;
assign _15544_ = _14782_ & _15547_ /*72735*/;
assign _15545_ = _14782_ ^ _15547_ /*72738*/;
assign _15546_ = _15538_ & _15545_ /*72736*/;
assign _15231_ = _15538_ ^ _15545_ /*72737*/;
assign _15543_ = _15544_ | _15546_ /*72734*/;
assign _15548_ = _14783_ & oneWire /*72729*/;
assign _15549_ = _14783_ ^ oneWire /*72732*/;
assign _15550_ = _15543_ & _15549_ /*72730*/;
assign _15232_ = _15543_ ^ _15549_ /*72731*/;
assign Q[46] = _15548_ | _15550_ /*72728*/;
assign _15683_ = ~Q[46] /*72343*/;
assign _15682_ = _15683_ & D[0] /*72342*/;
assign _15685_ = _15169_ & _15682_ /*72337*/;
assign _15686_ = _15169_ ^ _15682_ /*72340*/;
assign _15687_ = zeroWire & _15686_ /*72338*/;
assign _15617_ = zeroWire ^ _15686_ /*72339*/;
assign _15684_ = _15685_ | _15687_ /*72336*/;
assign _15689_ = ~Q[46] /*72335*/;
assign _15688_ = _15689_ & D[1] /*72334*/;
assign _15691_ = _15170_ & _15688_ /*72329*/;
assign _15692_ = _15170_ ^ _15688_ /*72332*/;
assign _15693_ = _15684_ & _15692_ /*72330*/;
assign _15618_ = _15684_ ^ _15692_ /*72331*/;
assign _15690_ = _15691_ | _15693_ /*72328*/;
assign _15695_ = ~Q[46] /*72327*/;
assign _15694_ = _15695_ & D[2] /*72326*/;
assign _15697_ = _15171_ & _15694_ /*72321*/;
assign _15698_ = _15171_ ^ _15694_ /*72324*/;
assign _15699_ = _15690_ & _15698_ /*72322*/;
assign _15619_ = _15690_ ^ _15698_ /*72323*/;
assign _15696_ = _15697_ | _15699_ /*72320*/;
assign _15701_ = ~Q[46] /*72319*/;
assign _15700_ = _15701_ & D[3] /*72318*/;
assign _15703_ = _15172_ & _15700_ /*72313*/;
assign _15704_ = _15172_ ^ _15700_ /*72316*/;
assign _15705_ = _15696_ & _15704_ /*72314*/;
assign _15620_ = _15696_ ^ _15704_ /*72315*/;
assign _15702_ = _15703_ | _15705_ /*72312*/;
assign _15707_ = ~Q[46] /*72311*/;
assign _15706_ = _15707_ & D[4] /*72310*/;
assign _15709_ = _15173_ & _15706_ /*72305*/;
assign _15710_ = _15173_ ^ _15706_ /*72308*/;
assign _15711_ = _15702_ & _15710_ /*72306*/;
assign _15621_ = _15702_ ^ _15710_ /*72307*/;
assign _15708_ = _15709_ | _15711_ /*72304*/;
assign _15713_ = ~Q[46] /*72303*/;
assign _15712_ = _15713_ & D[5] /*72302*/;
assign _15715_ = _15174_ & _15712_ /*72297*/;
assign _15716_ = _15174_ ^ _15712_ /*72300*/;
assign _15717_ = _15708_ & _15716_ /*72298*/;
assign _15622_ = _15708_ ^ _15716_ /*72299*/;
assign _15714_ = _15715_ | _15717_ /*72296*/;
assign _15719_ = ~Q[46] /*72295*/;
assign _15718_ = _15719_ & D[6] /*72294*/;
assign _15721_ = _15175_ & _15718_ /*72289*/;
assign _15722_ = _15175_ ^ _15718_ /*72292*/;
assign _15723_ = _15714_ & _15722_ /*72290*/;
assign _15623_ = _15714_ ^ _15722_ /*72291*/;
assign _15720_ = _15721_ | _15723_ /*72288*/;
assign _15725_ = ~Q[46] /*72287*/;
assign _15724_ = _15725_ & D[7] /*72286*/;
assign _15727_ = _15176_ & _15724_ /*72281*/;
assign _15728_ = _15176_ ^ _15724_ /*72284*/;
assign _15729_ = _15720_ & _15728_ /*72282*/;
assign _15624_ = _15720_ ^ _15728_ /*72283*/;
assign _15726_ = _15727_ | _15729_ /*72280*/;
assign _15731_ = ~Q[46] /*72279*/;
assign _15730_ = _15731_ & D[8] /*72278*/;
assign _15733_ = _15177_ & _15730_ /*72273*/;
assign _15734_ = _15177_ ^ _15730_ /*72276*/;
assign _15735_ = _15726_ & _15734_ /*72274*/;
assign _15625_ = _15726_ ^ _15734_ /*72275*/;
assign _15732_ = _15733_ | _15735_ /*72272*/;
assign _15737_ = ~Q[46] /*72271*/;
assign _15736_ = _15737_ & D[9] /*72270*/;
assign _15739_ = _15178_ & _15736_ /*72265*/;
assign _15740_ = _15178_ ^ _15736_ /*72268*/;
assign _15741_ = _15732_ & _15740_ /*72266*/;
assign _15626_ = _15732_ ^ _15740_ /*72267*/;
assign _15738_ = _15739_ | _15741_ /*72264*/;
assign _15743_ = ~Q[46] /*72263*/;
assign _15742_ = _15743_ & D[10] /*72262*/;
assign _15745_ = _15179_ & _15742_ /*72257*/;
assign _15746_ = _15179_ ^ _15742_ /*72260*/;
assign _15747_ = _15738_ & _15746_ /*72258*/;
assign _15627_ = _15738_ ^ _15746_ /*72259*/;
assign _15744_ = _15745_ | _15747_ /*72256*/;
assign _15749_ = ~Q[46] /*72255*/;
assign _15748_ = _15749_ & D[11] /*72254*/;
assign _15751_ = _15180_ & _15748_ /*72249*/;
assign _15752_ = _15180_ ^ _15748_ /*72252*/;
assign _15753_ = _15744_ & _15752_ /*72250*/;
assign _15628_ = _15744_ ^ _15752_ /*72251*/;
assign _15750_ = _15751_ | _15753_ /*72248*/;
assign _15755_ = ~Q[46] /*72247*/;
assign _15754_ = _15755_ & D[12] /*72246*/;
assign _15757_ = _15181_ & _15754_ /*72241*/;
assign _15758_ = _15181_ ^ _15754_ /*72244*/;
assign _15759_ = _15750_ & _15758_ /*72242*/;
assign _15629_ = _15750_ ^ _15758_ /*72243*/;
assign _15756_ = _15757_ | _15759_ /*72240*/;
assign _15761_ = ~Q[46] /*72239*/;
assign _15760_ = _15761_ & D[13] /*72238*/;
assign _15763_ = _15182_ & _15760_ /*72233*/;
assign _15764_ = _15182_ ^ _15760_ /*72236*/;
assign _15765_ = _15756_ & _15764_ /*72234*/;
assign _15630_ = _15756_ ^ _15764_ /*72235*/;
assign _15762_ = _15763_ | _15765_ /*72232*/;
assign _15767_ = ~Q[46] /*72231*/;
assign _15766_ = _15767_ & D[14] /*72230*/;
assign _15769_ = _15183_ & _15766_ /*72225*/;
assign _15770_ = _15183_ ^ _15766_ /*72228*/;
assign _15771_ = _15762_ & _15770_ /*72226*/;
assign _15631_ = _15762_ ^ _15770_ /*72227*/;
assign _15768_ = _15769_ | _15771_ /*72224*/;
assign _15773_ = ~Q[46] /*72223*/;
assign _15772_ = _15773_ & D[15] /*72222*/;
assign _15775_ = _15184_ & _15772_ /*72217*/;
assign _15776_ = _15184_ ^ _15772_ /*72220*/;
assign _15777_ = _15768_ & _15776_ /*72218*/;
assign _15632_ = _15768_ ^ _15776_ /*72219*/;
assign _15774_ = _15775_ | _15777_ /*72216*/;
assign _15779_ = ~Q[46] /*72215*/;
assign _15778_ = _15779_ & D[16] /*72214*/;
assign _15781_ = _15185_ & _15778_ /*72209*/;
assign _15782_ = _15185_ ^ _15778_ /*72212*/;
assign _15783_ = _15774_ & _15782_ /*72210*/;
assign _15633_ = _15774_ ^ _15782_ /*72211*/;
assign _15780_ = _15781_ | _15783_ /*72208*/;
assign _15785_ = ~Q[46] /*72207*/;
assign _15784_ = _15785_ & D[17] /*72206*/;
assign _15787_ = _15186_ & _15784_ /*72201*/;
assign _15788_ = _15186_ ^ _15784_ /*72204*/;
assign _15789_ = _15780_ & _15788_ /*72202*/;
assign _15634_ = _15780_ ^ _15788_ /*72203*/;
assign _15786_ = _15787_ | _15789_ /*72200*/;
assign _15791_ = ~Q[46] /*72199*/;
assign _15790_ = _15791_ & D[18] /*72198*/;
assign _15793_ = _15187_ & _15790_ /*72193*/;
assign _15794_ = _15187_ ^ _15790_ /*72196*/;
assign _15795_ = _15786_ & _15794_ /*72194*/;
assign _15635_ = _15786_ ^ _15794_ /*72195*/;
assign _15792_ = _15793_ | _15795_ /*72192*/;
assign _15797_ = ~Q[46] /*72191*/;
assign _15796_ = _15797_ & D[19] /*72190*/;
assign _15799_ = _15188_ & _15796_ /*72185*/;
assign _15800_ = _15188_ ^ _15796_ /*72188*/;
assign _15801_ = _15792_ & _15800_ /*72186*/;
assign _15636_ = _15792_ ^ _15800_ /*72187*/;
assign _15798_ = _15799_ | _15801_ /*72184*/;
assign _15803_ = ~Q[46] /*72183*/;
assign _15802_ = _15803_ & D[20] /*72182*/;
assign _15805_ = _15189_ & _15802_ /*72177*/;
assign _15806_ = _15189_ ^ _15802_ /*72180*/;
assign _15807_ = _15798_ & _15806_ /*72178*/;
assign _15637_ = _15798_ ^ _15806_ /*72179*/;
assign _15804_ = _15805_ | _15807_ /*72176*/;
assign _15809_ = ~Q[46] /*72175*/;
assign _15808_ = _15809_ & D[21] /*72174*/;
assign _15811_ = _15190_ & _15808_ /*72169*/;
assign _15812_ = _15190_ ^ _15808_ /*72172*/;
assign _15813_ = _15804_ & _15812_ /*72170*/;
assign _15638_ = _15804_ ^ _15812_ /*72171*/;
assign _15810_ = _15811_ | _15813_ /*72168*/;
assign _15815_ = ~Q[46] /*72167*/;
assign _15814_ = _15815_ & D[22] /*72166*/;
assign _15817_ = _15191_ & _15814_ /*72161*/;
assign _15818_ = _15191_ ^ _15814_ /*72164*/;
assign _15819_ = _15810_ & _15818_ /*72162*/;
assign _15639_ = _15810_ ^ _15818_ /*72163*/;
assign _15816_ = _15817_ | _15819_ /*72160*/;
assign _15821_ = ~Q[46] /*72159*/;
assign _15820_ = _15821_ & D[23] /*72158*/;
assign _15823_ = _15192_ & _15820_ /*72153*/;
assign _15824_ = _15192_ ^ _15820_ /*72156*/;
assign _15825_ = _15816_ & _15824_ /*72154*/;
assign _15640_ = _15816_ ^ _15824_ /*72155*/;
assign _15822_ = _15823_ | _15825_ /*72152*/;
assign _15827_ = ~Q[46] /*72151*/;
assign _15826_ = _15827_ & D[24] /*72150*/;
assign _15829_ = _15193_ & _15826_ /*72145*/;
assign _15830_ = _15193_ ^ _15826_ /*72148*/;
assign _15831_ = _15822_ & _15830_ /*72146*/;
assign _15641_ = _15822_ ^ _15830_ /*72147*/;
assign _15828_ = _15829_ | _15831_ /*72144*/;
assign _15833_ = ~Q[46] /*72143*/;
assign _15832_ = _15833_ & D[25] /*72142*/;
assign _15835_ = _15194_ & _15832_ /*72137*/;
assign _15836_ = _15194_ ^ _15832_ /*72140*/;
assign _15837_ = _15828_ & _15836_ /*72138*/;
assign _15642_ = _15828_ ^ _15836_ /*72139*/;
assign _15834_ = _15835_ | _15837_ /*72136*/;
assign _15839_ = ~Q[46] /*72135*/;
assign _15838_ = _15839_ & D[26] /*72134*/;
assign _15841_ = _15195_ & _15838_ /*72129*/;
assign _15842_ = _15195_ ^ _15838_ /*72132*/;
assign _15843_ = _15834_ & _15842_ /*72130*/;
assign _15643_ = _15834_ ^ _15842_ /*72131*/;
assign _15840_ = _15841_ | _15843_ /*72128*/;
assign _15845_ = ~Q[46] /*72127*/;
assign _15844_ = _15845_ & D[27] /*72126*/;
assign _15847_ = _15196_ & _15844_ /*72121*/;
assign _15848_ = _15196_ ^ _15844_ /*72124*/;
assign _15849_ = _15840_ & _15848_ /*72122*/;
assign _15644_ = _15840_ ^ _15848_ /*72123*/;
assign _15846_ = _15847_ | _15849_ /*72120*/;
assign _15851_ = ~Q[46] /*72119*/;
assign _15850_ = _15851_ & D[28] /*72118*/;
assign _15853_ = _15197_ & _15850_ /*72113*/;
assign _15854_ = _15197_ ^ _15850_ /*72116*/;
assign _15855_ = _15846_ & _15854_ /*72114*/;
assign _15645_ = _15846_ ^ _15854_ /*72115*/;
assign _15852_ = _15853_ | _15855_ /*72112*/;
assign _15857_ = ~Q[46] /*72111*/;
assign _15856_ = _15857_ & D[29] /*72110*/;
assign _15859_ = _15198_ & _15856_ /*72105*/;
assign _15860_ = _15198_ ^ _15856_ /*72108*/;
assign _15861_ = _15852_ & _15860_ /*72106*/;
assign _15646_ = _15852_ ^ _15860_ /*72107*/;
assign _15858_ = _15859_ | _15861_ /*72104*/;
assign _15863_ = ~Q[46] /*72103*/;
assign _15862_ = _15863_ & D[30] /*72102*/;
assign _15865_ = _15199_ & _15862_ /*72097*/;
assign _15866_ = _15199_ ^ _15862_ /*72100*/;
assign _15867_ = _15858_ & _15866_ /*72098*/;
assign _15647_ = _15858_ ^ _15866_ /*72099*/;
assign _15864_ = _15865_ | _15867_ /*72096*/;
assign _15869_ = ~Q[46] /*72095*/;
assign _15868_ = _15869_ & D[31] /*72094*/;
assign _15871_ = _15200_ & _15868_ /*72089*/;
assign _15872_ = _15200_ ^ _15868_ /*72092*/;
assign _15873_ = _15864_ & _15872_ /*72090*/;
assign _15648_ = _15864_ ^ _15872_ /*72091*/;
assign _15870_ = _15871_ | _15873_ /*72088*/;
assign _15875_ = ~Q[46] /*72087*/;
assign _15874_ = _15875_ & D[32] /*72086*/;
assign _15877_ = _15201_ & _15874_ /*72081*/;
assign _15878_ = _15201_ ^ _15874_ /*72084*/;
assign _15879_ = _15870_ & _15878_ /*72082*/;
assign _15649_ = _15870_ ^ _15878_ /*72083*/;
assign _15876_ = _15877_ | _15879_ /*72080*/;
assign _15881_ = ~Q[46] /*72079*/;
assign _15880_ = _15881_ & D[33] /*72078*/;
assign _15883_ = _15202_ & _15880_ /*72073*/;
assign _15884_ = _15202_ ^ _15880_ /*72076*/;
assign _15885_ = _15876_ & _15884_ /*72074*/;
assign _15650_ = _15876_ ^ _15884_ /*72075*/;
assign _15882_ = _15883_ | _15885_ /*72072*/;
assign _15887_ = ~Q[46] /*72071*/;
assign _15886_ = _15887_ & D[34] /*72070*/;
assign _15889_ = _15203_ & _15886_ /*72065*/;
assign _15890_ = _15203_ ^ _15886_ /*72068*/;
assign _15891_ = _15882_ & _15890_ /*72066*/;
assign _15651_ = _15882_ ^ _15890_ /*72067*/;
assign _15888_ = _15889_ | _15891_ /*72064*/;
assign _15893_ = ~Q[46] /*72063*/;
assign _15892_ = _15893_ & D[35] /*72062*/;
assign _15895_ = _15204_ & _15892_ /*72057*/;
assign _15896_ = _15204_ ^ _15892_ /*72060*/;
assign _15897_ = _15888_ & _15896_ /*72058*/;
assign _15652_ = _15888_ ^ _15896_ /*72059*/;
assign _15894_ = _15895_ | _15897_ /*72056*/;
assign _15899_ = ~Q[46] /*72055*/;
assign _15898_ = _15899_ & D[36] /*72054*/;
assign _15901_ = _15205_ & _15898_ /*72049*/;
assign _15902_ = _15205_ ^ _15898_ /*72052*/;
assign _15903_ = _15894_ & _15902_ /*72050*/;
assign _15653_ = _15894_ ^ _15902_ /*72051*/;
assign _15900_ = _15901_ | _15903_ /*72048*/;
assign _15905_ = ~Q[46] /*72047*/;
assign _15904_ = _15905_ & D[37] /*72046*/;
assign _15907_ = _15206_ & _15904_ /*72041*/;
assign _15908_ = _15206_ ^ _15904_ /*72044*/;
assign _15909_ = _15900_ & _15908_ /*72042*/;
assign _15654_ = _15900_ ^ _15908_ /*72043*/;
assign _15906_ = _15907_ | _15909_ /*72040*/;
assign _15911_ = ~Q[46] /*72039*/;
assign _15910_ = _15911_ & D[38] /*72038*/;
assign _15913_ = _15207_ & _15910_ /*72033*/;
assign _15914_ = _15207_ ^ _15910_ /*72036*/;
assign _15915_ = _15906_ & _15914_ /*72034*/;
assign _15655_ = _15906_ ^ _15914_ /*72035*/;
assign _15912_ = _15913_ | _15915_ /*72032*/;
assign _15917_ = ~Q[46] /*72031*/;
assign _15916_ = _15917_ & D[39] /*72030*/;
assign _15919_ = _15208_ & _15916_ /*72025*/;
assign _15920_ = _15208_ ^ _15916_ /*72028*/;
assign _15921_ = _15912_ & _15920_ /*72026*/;
assign _15656_ = _15912_ ^ _15920_ /*72027*/;
assign _15918_ = _15919_ | _15921_ /*72024*/;
assign _15923_ = ~Q[46] /*72023*/;
assign _15922_ = _15923_ & D[40] /*72022*/;
assign _15925_ = _15209_ & _15922_ /*72017*/;
assign _15926_ = _15209_ ^ _15922_ /*72020*/;
assign _15927_ = _15918_ & _15926_ /*72018*/;
assign _15657_ = _15918_ ^ _15926_ /*72019*/;
assign _15924_ = _15925_ | _15927_ /*72016*/;
assign _15929_ = ~Q[46] /*72015*/;
assign _15928_ = _15929_ & D[41] /*72014*/;
assign _15931_ = _15210_ & _15928_ /*72009*/;
assign _15932_ = _15210_ ^ _15928_ /*72012*/;
assign _15933_ = _15924_ & _15932_ /*72010*/;
assign _15658_ = _15924_ ^ _15932_ /*72011*/;
assign _15930_ = _15931_ | _15933_ /*72008*/;
assign _15935_ = ~Q[46] /*72007*/;
assign _15934_ = _15935_ & D[42] /*72006*/;
assign _15937_ = _15211_ & _15934_ /*72001*/;
assign _15938_ = _15211_ ^ _15934_ /*72004*/;
assign _15939_ = _15930_ & _15938_ /*72002*/;
assign _15659_ = _15930_ ^ _15938_ /*72003*/;
assign _15936_ = _15937_ | _15939_ /*72000*/;
assign _15941_ = ~Q[46] /*71999*/;
assign _15940_ = _15941_ & D[43] /*71998*/;
assign _15943_ = _15212_ & _15940_ /*71993*/;
assign _15944_ = _15212_ ^ _15940_ /*71996*/;
assign _15945_ = _15936_ & _15944_ /*71994*/;
assign _15660_ = _15936_ ^ _15944_ /*71995*/;
assign _15942_ = _15943_ | _15945_ /*71992*/;
assign _15947_ = ~Q[46] /*71991*/;
assign _15946_ = _15947_ & D[44] /*71990*/;
assign _15949_ = _15213_ & _15946_ /*71985*/;
assign _15950_ = _15213_ ^ _15946_ /*71988*/;
assign _15951_ = _15942_ & _15950_ /*71986*/;
assign _15661_ = _15942_ ^ _15950_ /*71987*/;
assign _15948_ = _15949_ | _15951_ /*71984*/;
assign _15953_ = ~Q[46] /*71983*/;
assign _15952_ = _15953_ & D[45] /*71982*/;
assign _15955_ = _15214_ & _15952_ /*71977*/;
assign _15956_ = _15214_ ^ _15952_ /*71980*/;
assign _15957_ = _15948_ & _15956_ /*71978*/;
assign _15662_ = _15948_ ^ _15956_ /*71979*/;
assign _15954_ = _15955_ | _15957_ /*71976*/;
assign _15959_ = ~Q[46] /*71975*/;
assign _15958_ = _15959_ & D[46] /*71974*/;
assign _15961_ = _15215_ & _15958_ /*71969*/;
assign _15962_ = _15215_ ^ _15958_ /*71972*/;
assign _15963_ = _15954_ & _15962_ /*71970*/;
assign _15663_ = _15954_ ^ _15962_ /*71971*/;
assign _15960_ = _15961_ | _15963_ /*71968*/;
assign _15965_ = ~Q[46] /*71967*/;
assign _15964_ = _15965_ & D[47] /*71966*/;
assign _15967_ = _15216_ & _15964_ /*71961*/;
assign _15968_ = _15216_ ^ _15964_ /*71964*/;
assign _15969_ = _15960_ & _15968_ /*71962*/;
assign _15664_ = _15960_ ^ _15968_ /*71963*/;
assign _15966_ = _15967_ | _15969_ /*71960*/;
assign _15971_ = ~Q[46] /*71959*/;
assign _15970_ = _15971_ & D[48] /*71958*/;
assign _15973_ = _15217_ & _15970_ /*71953*/;
assign _15974_ = _15217_ ^ _15970_ /*71956*/;
assign _15975_ = _15966_ & _15974_ /*71954*/;
assign _15665_ = _15966_ ^ _15974_ /*71955*/;
assign _15972_ = _15973_ | _15975_ /*71952*/;
assign _15977_ = ~Q[46] /*71951*/;
assign _15976_ = _15977_ & D[49] /*71950*/;
assign _15979_ = _15218_ & _15976_ /*71945*/;
assign _15980_ = _15218_ ^ _15976_ /*71948*/;
assign _15981_ = _15972_ & _15980_ /*71946*/;
assign _15666_ = _15972_ ^ _15980_ /*71947*/;
assign _15978_ = _15979_ | _15981_ /*71944*/;
assign _15983_ = ~Q[46] /*71943*/;
assign _15982_ = _15983_ & D[50] /*71942*/;
assign _15985_ = _15219_ & _15982_ /*71937*/;
assign _15986_ = _15219_ ^ _15982_ /*71940*/;
assign _15987_ = _15978_ & _15986_ /*71938*/;
assign _15667_ = _15978_ ^ _15986_ /*71939*/;
assign _15984_ = _15985_ | _15987_ /*71936*/;
assign _15989_ = ~Q[46] /*71935*/;
assign _15988_ = _15989_ & D[51] /*71934*/;
assign _15991_ = _15220_ & _15988_ /*71929*/;
assign _15992_ = _15220_ ^ _15988_ /*71932*/;
assign _15993_ = _15984_ & _15992_ /*71930*/;
assign _15668_ = _15984_ ^ _15992_ /*71931*/;
assign _15990_ = _15991_ | _15993_ /*71928*/;
assign _15995_ = ~Q[46] /*71927*/;
assign _15994_ = _15995_ & D[52] /*71926*/;
assign _15997_ = _15221_ & _15994_ /*71921*/;
assign _15998_ = _15221_ ^ _15994_ /*71924*/;
assign _15999_ = _15990_ & _15998_ /*71922*/;
assign _15669_ = _15990_ ^ _15998_ /*71923*/;
assign _15996_ = _15997_ | _15999_ /*71920*/;
assign _16001_ = ~Q[46] /*71919*/;
assign _16000_ = _16001_ & D[53] /*71918*/;
assign _16003_ = _15222_ & _16000_ /*71913*/;
assign _16004_ = _15222_ ^ _16000_ /*71916*/;
assign _16005_ = _15996_ & _16004_ /*71914*/;
assign _15670_ = _15996_ ^ _16004_ /*71915*/;
assign _16002_ = _16003_ | _16005_ /*71912*/;
assign _16007_ = ~Q[46] /*71911*/;
assign _16006_ = _16007_ & D[54] /*71910*/;
assign _16009_ = _15223_ & _16006_ /*71905*/;
assign _16010_ = _15223_ ^ _16006_ /*71908*/;
assign _16011_ = _16002_ & _16010_ /*71906*/;
assign _15671_ = _16002_ ^ _16010_ /*71907*/;
assign _16008_ = _16009_ | _16011_ /*71904*/;
assign _16013_ = ~Q[46] /*71903*/;
assign _16012_ = _16013_ & D[55] /*71902*/;
assign _16015_ = _15224_ & _16012_ /*71897*/;
assign _16016_ = _15224_ ^ _16012_ /*71900*/;
assign _16017_ = _16008_ & _16016_ /*71898*/;
assign _15672_ = _16008_ ^ _16016_ /*71899*/;
assign _16014_ = _16015_ | _16017_ /*71896*/;
assign _16019_ = ~Q[46] /*71895*/;
assign _16018_ = _16019_ & D[56] /*71894*/;
assign _16021_ = _15225_ & _16018_ /*71889*/;
assign _16022_ = _15225_ ^ _16018_ /*71892*/;
assign _16023_ = _16014_ & _16022_ /*71890*/;
assign _15673_ = _16014_ ^ _16022_ /*71891*/;
assign _16020_ = _16021_ | _16023_ /*71888*/;
assign _16025_ = ~Q[46] /*71887*/;
assign _16024_ = _16025_ & D[57] /*71886*/;
assign _16027_ = _15226_ & _16024_ /*71881*/;
assign _16028_ = _15226_ ^ _16024_ /*71884*/;
assign _16029_ = _16020_ & _16028_ /*71882*/;
assign _15674_ = _16020_ ^ _16028_ /*71883*/;
assign _16026_ = _16027_ | _16029_ /*71880*/;
assign _16031_ = ~Q[46] /*71879*/;
assign _16030_ = _16031_ & D[58] /*71878*/;
assign _16033_ = _15227_ & _16030_ /*71873*/;
assign _16034_ = _15227_ ^ _16030_ /*71876*/;
assign _16035_ = _16026_ & _16034_ /*71874*/;
assign _15675_ = _16026_ ^ _16034_ /*71875*/;
assign _16032_ = _16033_ | _16035_ /*71872*/;
assign _16037_ = ~Q[46] /*71871*/;
assign _16036_ = _16037_ & D[59] /*71870*/;
assign _16039_ = _15228_ & _16036_ /*71865*/;
assign _16040_ = _15228_ ^ _16036_ /*71868*/;
assign _16041_ = _16032_ & _16040_ /*71866*/;
assign _15676_ = _16032_ ^ _16040_ /*71867*/;
assign _16038_ = _16039_ | _16041_ /*71864*/;
assign _16043_ = ~Q[46] /*71863*/;
assign _16042_ = _16043_ & D[60] /*71862*/;
assign _16045_ = _15229_ & _16042_ /*71857*/;
assign _16046_ = _15229_ ^ _16042_ /*71860*/;
assign _16047_ = _16038_ & _16046_ /*71858*/;
assign _15677_ = _16038_ ^ _16046_ /*71859*/;
assign _16044_ = _16045_ | _16047_ /*71856*/;
assign _16049_ = ~Q[46] /*71855*/;
assign _16048_ = _16049_ & D[61] /*71854*/;
assign _16051_ = _15230_ & _16048_ /*71849*/;
assign _16052_ = _15230_ ^ _16048_ /*71852*/;
assign _16053_ = _16044_ & _16052_ /*71850*/;
assign _15678_ = _16044_ ^ _16052_ /*71851*/;
assign _16050_ = _16051_ | _16053_ /*71848*/;
assign _16055_ = ~Q[46] /*71847*/;
assign _16054_ = _16055_ & D[62] /*71846*/;
assign _16057_ = _15231_ & _16054_ /*71841*/;
assign _16058_ = _15231_ ^ _16054_ /*71844*/;
assign _16059_ = _16050_ & _16058_ /*71842*/;
assign _15679_ = _16050_ ^ _16058_ /*71843*/;
assign _16056_ = _16057_ | _16059_ /*71840*/;
assign _16061_ = ~Q[46] /*71839*/;
assign _16060_ = _16061_ & zeroWire /*71838*/;
assign _16062_ = _15232_ ^ _16060_ /*71836*/;
assign _15680_ = _16062_ ^ _16056_ /*71835*/;
assign _16133_ = ~D[0] /*71581*/;
assign _16130_ = R_0[45] & _16133_ /*71577*/;
assign _16131_ = R_0[45] ^ _16133_ /*71580*/;
assign _16132_ = oneWire & _16131_ /*71578*/;
assign _16065_ = oneWire ^ _16131_ /*71579*/;
assign _16129_ = _16130_ | _16132_ /*71576*/;
assign _16138_ = ~D[1] /*71575*/;
assign _16135_ = _15617_ & _16138_ /*71571*/;
assign _16136_ = _15617_ ^ _16138_ /*71574*/;
assign _16137_ = _16129_ & _16136_ /*71572*/;
assign _16066_ = _16129_ ^ _16136_ /*71573*/;
assign _16134_ = _16135_ | _16137_ /*71570*/;
assign _16143_ = ~D[2] /*71569*/;
assign _16140_ = _15618_ & _16143_ /*71565*/;
assign _16141_ = _15618_ ^ _16143_ /*71568*/;
assign _16142_ = _16134_ & _16141_ /*71566*/;
assign _16067_ = _16134_ ^ _16141_ /*71567*/;
assign _16139_ = _16140_ | _16142_ /*71564*/;
assign _16148_ = ~D[3] /*71563*/;
assign _16145_ = _15619_ & _16148_ /*71559*/;
assign _16146_ = _15619_ ^ _16148_ /*71562*/;
assign _16147_ = _16139_ & _16146_ /*71560*/;
assign _16068_ = _16139_ ^ _16146_ /*71561*/;
assign _16144_ = _16145_ | _16147_ /*71558*/;
assign _16153_ = ~D[4] /*71557*/;
assign _16150_ = _15620_ & _16153_ /*71553*/;
assign _16151_ = _15620_ ^ _16153_ /*71556*/;
assign _16152_ = _16144_ & _16151_ /*71554*/;
assign _16069_ = _16144_ ^ _16151_ /*71555*/;
assign _16149_ = _16150_ | _16152_ /*71552*/;
assign _16158_ = ~D[5] /*71551*/;
assign _16155_ = _15621_ & _16158_ /*71547*/;
assign _16156_ = _15621_ ^ _16158_ /*71550*/;
assign _16157_ = _16149_ & _16156_ /*71548*/;
assign _16070_ = _16149_ ^ _16156_ /*71549*/;
assign _16154_ = _16155_ | _16157_ /*71546*/;
assign _16163_ = ~D[6] /*71545*/;
assign _16160_ = _15622_ & _16163_ /*71541*/;
assign _16161_ = _15622_ ^ _16163_ /*71544*/;
assign _16162_ = _16154_ & _16161_ /*71542*/;
assign _16071_ = _16154_ ^ _16161_ /*71543*/;
assign _16159_ = _16160_ | _16162_ /*71540*/;
assign _16168_ = ~D[7] /*71539*/;
assign _16165_ = _15623_ & _16168_ /*71535*/;
assign _16166_ = _15623_ ^ _16168_ /*71538*/;
assign _16167_ = _16159_ & _16166_ /*71536*/;
assign _16072_ = _16159_ ^ _16166_ /*71537*/;
assign _16164_ = _16165_ | _16167_ /*71534*/;
assign _16173_ = ~D[8] /*71533*/;
assign _16170_ = _15624_ & _16173_ /*71529*/;
assign _16171_ = _15624_ ^ _16173_ /*71532*/;
assign _16172_ = _16164_ & _16171_ /*71530*/;
assign _16073_ = _16164_ ^ _16171_ /*71531*/;
assign _16169_ = _16170_ | _16172_ /*71528*/;
assign _16178_ = ~D[9] /*71527*/;
assign _16175_ = _15625_ & _16178_ /*71523*/;
assign _16176_ = _15625_ ^ _16178_ /*71526*/;
assign _16177_ = _16169_ & _16176_ /*71524*/;
assign _16074_ = _16169_ ^ _16176_ /*71525*/;
assign _16174_ = _16175_ | _16177_ /*71522*/;
assign _16183_ = ~D[10] /*71521*/;
assign _16180_ = _15626_ & _16183_ /*71517*/;
assign _16181_ = _15626_ ^ _16183_ /*71520*/;
assign _16182_ = _16174_ & _16181_ /*71518*/;
assign _16075_ = _16174_ ^ _16181_ /*71519*/;
assign _16179_ = _16180_ | _16182_ /*71516*/;
assign _16188_ = ~D[11] /*71515*/;
assign _16185_ = _15627_ & _16188_ /*71511*/;
assign _16186_ = _15627_ ^ _16188_ /*71514*/;
assign _16187_ = _16179_ & _16186_ /*71512*/;
assign _16076_ = _16179_ ^ _16186_ /*71513*/;
assign _16184_ = _16185_ | _16187_ /*71510*/;
assign _16193_ = ~D[12] /*71509*/;
assign _16190_ = _15628_ & _16193_ /*71505*/;
assign _16191_ = _15628_ ^ _16193_ /*71508*/;
assign _16192_ = _16184_ & _16191_ /*71506*/;
assign _16077_ = _16184_ ^ _16191_ /*71507*/;
assign _16189_ = _16190_ | _16192_ /*71504*/;
assign _16198_ = ~D[13] /*71503*/;
assign _16195_ = _15629_ & _16198_ /*71499*/;
assign _16196_ = _15629_ ^ _16198_ /*71502*/;
assign _16197_ = _16189_ & _16196_ /*71500*/;
assign _16078_ = _16189_ ^ _16196_ /*71501*/;
assign _16194_ = _16195_ | _16197_ /*71498*/;
assign _16203_ = ~D[14] /*71497*/;
assign _16200_ = _15630_ & _16203_ /*71493*/;
assign _16201_ = _15630_ ^ _16203_ /*71496*/;
assign _16202_ = _16194_ & _16201_ /*71494*/;
assign _16079_ = _16194_ ^ _16201_ /*71495*/;
assign _16199_ = _16200_ | _16202_ /*71492*/;
assign _16208_ = ~D[15] /*71491*/;
assign _16205_ = _15631_ & _16208_ /*71487*/;
assign _16206_ = _15631_ ^ _16208_ /*71490*/;
assign _16207_ = _16199_ & _16206_ /*71488*/;
assign _16080_ = _16199_ ^ _16206_ /*71489*/;
assign _16204_ = _16205_ | _16207_ /*71486*/;
assign _16213_ = ~D[16] /*71485*/;
assign _16210_ = _15632_ & _16213_ /*71481*/;
assign _16211_ = _15632_ ^ _16213_ /*71484*/;
assign _16212_ = _16204_ & _16211_ /*71482*/;
assign _16081_ = _16204_ ^ _16211_ /*71483*/;
assign _16209_ = _16210_ | _16212_ /*71480*/;
assign _16218_ = ~D[17] /*71479*/;
assign _16215_ = _15633_ & _16218_ /*71475*/;
assign _16216_ = _15633_ ^ _16218_ /*71478*/;
assign _16217_ = _16209_ & _16216_ /*71476*/;
assign _16082_ = _16209_ ^ _16216_ /*71477*/;
assign _16214_ = _16215_ | _16217_ /*71474*/;
assign _16223_ = ~D[18] /*71473*/;
assign _16220_ = _15634_ & _16223_ /*71469*/;
assign _16221_ = _15634_ ^ _16223_ /*71472*/;
assign _16222_ = _16214_ & _16221_ /*71470*/;
assign _16083_ = _16214_ ^ _16221_ /*71471*/;
assign _16219_ = _16220_ | _16222_ /*71468*/;
assign _16228_ = ~D[19] /*71467*/;
assign _16225_ = _15635_ & _16228_ /*71463*/;
assign _16226_ = _15635_ ^ _16228_ /*71466*/;
assign _16227_ = _16219_ & _16226_ /*71464*/;
assign _16084_ = _16219_ ^ _16226_ /*71465*/;
assign _16224_ = _16225_ | _16227_ /*71462*/;
assign _16233_ = ~D[20] /*71461*/;
assign _16230_ = _15636_ & _16233_ /*71457*/;
assign _16231_ = _15636_ ^ _16233_ /*71460*/;
assign _16232_ = _16224_ & _16231_ /*71458*/;
assign _16085_ = _16224_ ^ _16231_ /*71459*/;
assign _16229_ = _16230_ | _16232_ /*71456*/;
assign _16238_ = ~D[21] /*71455*/;
assign _16235_ = _15637_ & _16238_ /*71451*/;
assign _16236_ = _15637_ ^ _16238_ /*71454*/;
assign _16237_ = _16229_ & _16236_ /*71452*/;
assign _16086_ = _16229_ ^ _16236_ /*71453*/;
assign _16234_ = _16235_ | _16237_ /*71450*/;
assign _16243_ = ~D[22] /*71449*/;
assign _16240_ = _15638_ & _16243_ /*71445*/;
assign _16241_ = _15638_ ^ _16243_ /*71448*/;
assign _16242_ = _16234_ & _16241_ /*71446*/;
assign _16087_ = _16234_ ^ _16241_ /*71447*/;
assign _16239_ = _16240_ | _16242_ /*71444*/;
assign _16248_ = ~D[23] /*71443*/;
assign _16245_ = _15639_ & _16248_ /*71439*/;
assign _16246_ = _15639_ ^ _16248_ /*71442*/;
assign _16247_ = _16239_ & _16246_ /*71440*/;
assign _16088_ = _16239_ ^ _16246_ /*71441*/;
assign _16244_ = _16245_ | _16247_ /*71438*/;
assign _16253_ = ~D[24] /*71437*/;
assign _16250_ = _15640_ & _16253_ /*71433*/;
assign _16251_ = _15640_ ^ _16253_ /*71436*/;
assign _16252_ = _16244_ & _16251_ /*71434*/;
assign _16089_ = _16244_ ^ _16251_ /*71435*/;
assign _16249_ = _16250_ | _16252_ /*71432*/;
assign _16258_ = ~D[25] /*71431*/;
assign _16255_ = _15641_ & _16258_ /*71427*/;
assign _16256_ = _15641_ ^ _16258_ /*71430*/;
assign _16257_ = _16249_ & _16256_ /*71428*/;
assign _16090_ = _16249_ ^ _16256_ /*71429*/;
assign _16254_ = _16255_ | _16257_ /*71426*/;
assign _16263_ = ~D[26] /*71425*/;
assign _16260_ = _15642_ & _16263_ /*71421*/;
assign _16261_ = _15642_ ^ _16263_ /*71424*/;
assign _16262_ = _16254_ & _16261_ /*71422*/;
assign _16091_ = _16254_ ^ _16261_ /*71423*/;
assign _16259_ = _16260_ | _16262_ /*71420*/;
assign _16268_ = ~D[27] /*71419*/;
assign _16265_ = _15643_ & _16268_ /*71415*/;
assign _16266_ = _15643_ ^ _16268_ /*71418*/;
assign _16267_ = _16259_ & _16266_ /*71416*/;
assign _16092_ = _16259_ ^ _16266_ /*71417*/;
assign _16264_ = _16265_ | _16267_ /*71414*/;
assign _16273_ = ~D[28] /*71413*/;
assign _16270_ = _15644_ & _16273_ /*71409*/;
assign _16271_ = _15644_ ^ _16273_ /*71412*/;
assign _16272_ = _16264_ & _16271_ /*71410*/;
assign _16093_ = _16264_ ^ _16271_ /*71411*/;
assign _16269_ = _16270_ | _16272_ /*71408*/;
assign _16278_ = ~D[29] /*71407*/;
assign _16275_ = _15645_ & _16278_ /*71403*/;
assign _16276_ = _15645_ ^ _16278_ /*71406*/;
assign _16277_ = _16269_ & _16276_ /*71404*/;
assign _16094_ = _16269_ ^ _16276_ /*71405*/;
assign _16274_ = _16275_ | _16277_ /*71402*/;
assign _16283_ = ~D[30] /*71401*/;
assign _16280_ = _15646_ & _16283_ /*71397*/;
assign _16281_ = _15646_ ^ _16283_ /*71400*/;
assign _16282_ = _16274_ & _16281_ /*71398*/;
assign _16095_ = _16274_ ^ _16281_ /*71399*/;
assign _16279_ = _16280_ | _16282_ /*71396*/;
assign _16288_ = ~D[31] /*71395*/;
assign _16285_ = _15647_ & _16288_ /*71391*/;
assign _16286_ = _15647_ ^ _16288_ /*71394*/;
assign _16287_ = _16279_ & _16286_ /*71392*/;
assign _16096_ = _16279_ ^ _16286_ /*71393*/;
assign _16284_ = _16285_ | _16287_ /*71390*/;
assign _16293_ = ~D[32] /*71389*/;
assign _16290_ = _15648_ & _16293_ /*71385*/;
assign _16291_ = _15648_ ^ _16293_ /*71388*/;
assign _16292_ = _16284_ & _16291_ /*71386*/;
assign _16097_ = _16284_ ^ _16291_ /*71387*/;
assign _16289_ = _16290_ | _16292_ /*71384*/;
assign _16298_ = ~D[33] /*71383*/;
assign _16295_ = _15649_ & _16298_ /*71379*/;
assign _16296_ = _15649_ ^ _16298_ /*71382*/;
assign _16297_ = _16289_ & _16296_ /*71380*/;
assign _16098_ = _16289_ ^ _16296_ /*71381*/;
assign _16294_ = _16295_ | _16297_ /*71378*/;
assign _16303_ = ~D[34] /*71377*/;
assign _16300_ = _15650_ & _16303_ /*71373*/;
assign _16301_ = _15650_ ^ _16303_ /*71376*/;
assign _16302_ = _16294_ & _16301_ /*71374*/;
assign _16099_ = _16294_ ^ _16301_ /*71375*/;
assign _16299_ = _16300_ | _16302_ /*71372*/;
assign _16308_ = ~D[35] /*71371*/;
assign _16305_ = _15651_ & _16308_ /*71367*/;
assign _16306_ = _15651_ ^ _16308_ /*71370*/;
assign _16307_ = _16299_ & _16306_ /*71368*/;
assign _16100_ = _16299_ ^ _16306_ /*71369*/;
assign _16304_ = _16305_ | _16307_ /*71366*/;
assign _16313_ = ~D[36] /*71365*/;
assign _16310_ = _15652_ & _16313_ /*71361*/;
assign _16311_ = _15652_ ^ _16313_ /*71364*/;
assign _16312_ = _16304_ & _16311_ /*71362*/;
assign _16101_ = _16304_ ^ _16311_ /*71363*/;
assign _16309_ = _16310_ | _16312_ /*71360*/;
assign _16318_ = ~D[37] /*71359*/;
assign _16315_ = _15653_ & _16318_ /*71355*/;
assign _16316_ = _15653_ ^ _16318_ /*71358*/;
assign _16317_ = _16309_ & _16316_ /*71356*/;
assign _16102_ = _16309_ ^ _16316_ /*71357*/;
assign _16314_ = _16315_ | _16317_ /*71354*/;
assign _16323_ = ~D[38] /*71353*/;
assign _16320_ = _15654_ & _16323_ /*71349*/;
assign _16321_ = _15654_ ^ _16323_ /*71352*/;
assign _16322_ = _16314_ & _16321_ /*71350*/;
assign _16103_ = _16314_ ^ _16321_ /*71351*/;
assign _16319_ = _16320_ | _16322_ /*71348*/;
assign _16328_ = ~D[39] /*71347*/;
assign _16325_ = _15655_ & _16328_ /*71343*/;
assign _16326_ = _15655_ ^ _16328_ /*71346*/;
assign _16327_ = _16319_ & _16326_ /*71344*/;
assign _16104_ = _16319_ ^ _16326_ /*71345*/;
assign _16324_ = _16325_ | _16327_ /*71342*/;
assign _16333_ = ~D[40] /*71341*/;
assign _16330_ = _15656_ & _16333_ /*71337*/;
assign _16331_ = _15656_ ^ _16333_ /*71340*/;
assign _16332_ = _16324_ & _16331_ /*71338*/;
assign _16105_ = _16324_ ^ _16331_ /*71339*/;
assign _16329_ = _16330_ | _16332_ /*71336*/;
assign _16338_ = ~D[41] /*71335*/;
assign _16335_ = _15657_ & _16338_ /*71331*/;
assign _16336_ = _15657_ ^ _16338_ /*71334*/;
assign _16337_ = _16329_ & _16336_ /*71332*/;
assign _16106_ = _16329_ ^ _16336_ /*71333*/;
assign _16334_ = _16335_ | _16337_ /*71330*/;
assign _16343_ = ~D[42] /*71329*/;
assign _16340_ = _15658_ & _16343_ /*71325*/;
assign _16341_ = _15658_ ^ _16343_ /*71328*/;
assign _16342_ = _16334_ & _16341_ /*71326*/;
assign _16107_ = _16334_ ^ _16341_ /*71327*/;
assign _16339_ = _16340_ | _16342_ /*71324*/;
assign _16348_ = ~D[43] /*71323*/;
assign _16345_ = _15659_ & _16348_ /*71319*/;
assign _16346_ = _15659_ ^ _16348_ /*71322*/;
assign _16347_ = _16339_ & _16346_ /*71320*/;
assign _16108_ = _16339_ ^ _16346_ /*71321*/;
assign _16344_ = _16345_ | _16347_ /*71318*/;
assign _16353_ = ~D[44] /*71317*/;
assign _16350_ = _15660_ & _16353_ /*71313*/;
assign _16351_ = _15660_ ^ _16353_ /*71316*/;
assign _16352_ = _16344_ & _16351_ /*71314*/;
assign _16109_ = _16344_ ^ _16351_ /*71315*/;
assign _16349_ = _16350_ | _16352_ /*71312*/;
assign _16358_ = ~D[45] /*71311*/;
assign _16355_ = _15661_ & _16358_ /*71307*/;
assign _16356_ = _15661_ ^ _16358_ /*71310*/;
assign _16357_ = _16349_ & _16356_ /*71308*/;
assign _16110_ = _16349_ ^ _16356_ /*71309*/;
assign _16354_ = _16355_ | _16357_ /*71306*/;
assign _16363_ = ~D[46] /*71305*/;
assign _16360_ = _15662_ & _16363_ /*71301*/;
assign _16361_ = _15662_ ^ _16363_ /*71304*/;
assign _16362_ = _16354_ & _16361_ /*71302*/;
assign _16111_ = _16354_ ^ _16361_ /*71303*/;
assign _16359_ = _16360_ | _16362_ /*71300*/;
assign _16368_ = ~D[47] /*71299*/;
assign _16365_ = _15663_ & _16368_ /*71295*/;
assign _16366_ = _15663_ ^ _16368_ /*71298*/;
assign _16367_ = _16359_ & _16366_ /*71296*/;
assign _16112_ = _16359_ ^ _16366_ /*71297*/;
assign _16364_ = _16365_ | _16367_ /*71294*/;
assign _16373_ = ~D[48] /*71293*/;
assign _16370_ = _15664_ & _16373_ /*71289*/;
assign _16371_ = _15664_ ^ _16373_ /*71292*/;
assign _16372_ = _16364_ & _16371_ /*71290*/;
assign _16113_ = _16364_ ^ _16371_ /*71291*/;
assign _16369_ = _16370_ | _16372_ /*71288*/;
assign _16378_ = ~D[49] /*71287*/;
assign _16375_ = _15665_ & _16378_ /*71283*/;
assign _16376_ = _15665_ ^ _16378_ /*71286*/;
assign _16377_ = _16369_ & _16376_ /*71284*/;
assign _16114_ = _16369_ ^ _16376_ /*71285*/;
assign _16374_ = _16375_ | _16377_ /*71282*/;
assign _16383_ = ~D[50] /*71281*/;
assign _16380_ = _15666_ & _16383_ /*71277*/;
assign _16381_ = _15666_ ^ _16383_ /*71280*/;
assign _16382_ = _16374_ & _16381_ /*71278*/;
assign _16115_ = _16374_ ^ _16381_ /*71279*/;
assign _16379_ = _16380_ | _16382_ /*71276*/;
assign _16388_ = ~D[51] /*71275*/;
assign _16385_ = _15667_ & _16388_ /*71271*/;
assign _16386_ = _15667_ ^ _16388_ /*71274*/;
assign _16387_ = _16379_ & _16386_ /*71272*/;
assign _16116_ = _16379_ ^ _16386_ /*71273*/;
assign _16384_ = _16385_ | _16387_ /*71270*/;
assign _16393_ = ~D[52] /*71269*/;
assign _16390_ = _15668_ & _16393_ /*71265*/;
assign _16391_ = _15668_ ^ _16393_ /*71268*/;
assign _16392_ = _16384_ & _16391_ /*71266*/;
assign _16117_ = _16384_ ^ _16391_ /*71267*/;
assign _16389_ = _16390_ | _16392_ /*71264*/;
assign _16398_ = ~D[53] /*71263*/;
assign _16395_ = _15669_ & _16398_ /*71259*/;
assign _16396_ = _15669_ ^ _16398_ /*71262*/;
assign _16397_ = _16389_ & _16396_ /*71260*/;
assign _16118_ = _16389_ ^ _16396_ /*71261*/;
assign _16394_ = _16395_ | _16397_ /*71258*/;
assign _16403_ = ~D[54] /*71257*/;
assign _16400_ = _15670_ & _16403_ /*71253*/;
assign _16401_ = _15670_ ^ _16403_ /*71256*/;
assign _16402_ = _16394_ & _16401_ /*71254*/;
assign _16119_ = _16394_ ^ _16401_ /*71255*/;
assign _16399_ = _16400_ | _16402_ /*71252*/;
assign _16408_ = ~D[55] /*71251*/;
assign _16405_ = _15671_ & _16408_ /*71247*/;
assign _16406_ = _15671_ ^ _16408_ /*71250*/;
assign _16407_ = _16399_ & _16406_ /*71248*/;
assign _16120_ = _16399_ ^ _16406_ /*71249*/;
assign _16404_ = _16405_ | _16407_ /*71246*/;
assign _16413_ = ~D[56] /*71245*/;
assign _16410_ = _15672_ & _16413_ /*71241*/;
assign _16411_ = _15672_ ^ _16413_ /*71244*/;
assign _16412_ = _16404_ & _16411_ /*71242*/;
assign _16121_ = _16404_ ^ _16411_ /*71243*/;
assign _16409_ = _16410_ | _16412_ /*71240*/;
assign _16418_ = ~D[57] /*71239*/;
assign _16415_ = _15673_ & _16418_ /*71235*/;
assign _16416_ = _15673_ ^ _16418_ /*71238*/;
assign _16417_ = _16409_ & _16416_ /*71236*/;
assign _16122_ = _16409_ ^ _16416_ /*71237*/;
assign _16414_ = _16415_ | _16417_ /*71234*/;
assign _16423_ = ~D[58] /*71233*/;
assign _16420_ = _15674_ & _16423_ /*71229*/;
assign _16421_ = _15674_ ^ _16423_ /*71232*/;
assign _16422_ = _16414_ & _16421_ /*71230*/;
assign _16123_ = _16414_ ^ _16421_ /*71231*/;
assign _16419_ = _16420_ | _16422_ /*71228*/;
assign _16428_ = ~D[59] /*71227*/;
assign _16425_ = _15675_ & _16428_ /*71223*/;
assign _16426_ = _15675_ ^ _16428_ /*71226*/;
assign _16427_ = _16419_ & _16426_ /*71224*/;
assign _16124_ = _16419_ ^ _16426_ /*71225*/;
assign _16424_ = _16425_ | _16427_ /*71222*/;
assign _16433_ = ~D[60] /*71221*/;
assign _16430_ = _15676_ & _16433_ /*71217*/;
assign _16431_ = _15676_ ^ _16433_ /*71220*/;
assign _16432_ = _16424_ & _16431_ /*71218*/;
assign _16125_ = _16424_ ^ _16431_ /*71219*/;
assign _16429_ = _16430_ | _16432_ /*71216*/;
assign _16438_ = ~D[61] /*71215*/;
assign _16435_ = _15677_ & _16438_ /*71211*/;
assign _16436_ = _15677_ ^ _16438_ /*71214*/;
assign _16437_ = _16429_ & _16436_ /*71212*/;
assign _16126_ = _16429_ ^ _16436_ /*71213*/;
assign _16434_ = _16435_ | _16437_ /*71210*/;
assign _16443_ = ~D[62] /*71209*/;
assign _16440_ = _15678_ & _16443_ /*71205*/;
assign _16441_ = _15678_ ^ _16443_ /*71208*/;
assign _16442_ = _16434_ & _16441_ /*71206*/;
assign _16127_ = _16434_ ^ _16441_ /*71207*/;
assign _16439_ = _16440_ | _16442_ /*71204*/;
assign _16444_ = _15679_ & oneWire /*71199*/;
assign _16445_ = _15679_ ^ oneWire /*71202*/;
assign _16446_ = _16439_ & _16445_ /*71200*/;
assign _16128_ = _16439_ ^ _16445_ /*71201*/;
assign Q[45] = _16444_ | _16446_ /*71198*/;
assign _16579_ = ~Q[45] /*70813*/;
assign _16578_ = _16579_ & D[0] /*70812*/;
assign _16581_ = _16065_ & _16578_ /*70807*/;
assign _16582_ = _16065_ ^ _16578_ /*70810*/;
assign _16583_ = zeroWire & _16582_ /*70808*/;
assign _16513_ = zeroWire ^ _16582_ /*70809*/;
assign _16580_ = _16581_ | _16583_ /*70806*/;
assign _16585_ = ~Q[45] /*70805*/;
assign _16584_ = _16585_ & D[1] /*70804*/;
assign _16587_ = _16066_ & _16584_ /*70799*/;
assign _16588_ = _16066_ ^ _16584_ /*70802*/;
assign _16589_ = _16580_ & _16588_ /*70800*/;
assign _16514_ = _16580_ ^ _16588_ /*70801*/;
assign _16586_ = _16587_ | _16589_ /*70798*/;
assign _16591_ = ~Q[45] /*70797*/;
assign _16590_ = _16591_ & D[2] /*70796*/;
assign _16593_ = _16067_ & _16590_ /*70791*/;
assign _16594_ = _16067_ ^ _16590_ /*70794*/;
assign _16595_ = _16586_ & _16594_ /*70792*/;
assign _16515_ = _16586_ ^ _16594_ /*70793*/;
assign _16592_ = _16593_ | _16595_ /*70790*/;
assign _16597_ = ~Q[45] /*70789*/;
assign _16596_ = _16597_ & D[3] /*70788*/;
assign _16599_ = _16068_ & _16596_ /*70783*/;
assign _16600_ = _16068_ ^ _16596_ /*70786*/;
assign _16601_ = _16592_ & _16600_ /*70784*/;
assign _16516_ = _16592_ ^ _16600_ /*70785*/;
assign _16598_ = _16599_ | _16601_ /*70782*/;
assign _16603_ = ~Q[45] /*70781*/;
assign _16602_ = _16603_ & D[4] /*70780*/;
assign _16605_ = _16069_ & _16602_ /*70775*/;
assign _16606_ = _16069_ ^ _16602_ /*70778*/;
assign _16607_ = _16598_ & _16606_ /*70776*/;
assign _16517_ = _16598_ ^ _16606_ /*70777*/;
assign _16604_ = _16605_ | _16607_ /*70774*/;
assign _16609_ = ~Q[45] /*70773*/;
assign _16608_ = _16609_ & D[5] /*70772*/;
assign _16611_ = _16070_ & _16608_ /*70767*/;
assign _16612_ = _16070_ ^ _16608_ /*70770*/;
assign _16613_ = _16604_ & _16612_ /*70768*/;
assign _16518_ = _16604_ ^ _16612_ /*70769*/;
assign _16610_ = _16611_ | _16613_ /*70766*/;
assign _16615_ = ~Q[45] /*70765*/;
assign _16614_ = _16615_ & D[6] /*70764*/;
assign _16617_ = _16071_ & _16614_ /*70759*/;
assign _16618_ = _16071_ ^ _16614_ /*70762*/;
assign _16619_ = _16610_ & _16618_ /*70760*/;
assign _16519_ = _16610_ ^ _16618_ /*70761*/;
assign _16616_ = _16617_ | _16619_ /*70758*/;
assign _16621_ = ~Q[45] /*70757*/;
assign _16620_ = _16621_ & D[7] /*70756*/;
assign _16623_ = _16072_ & _16620_ /*70751*/;
assign _16624_ = _16072_ ^ _16620_ /*70754*/;
assign _16625_ = _16616_ & _16624_ /*70752*/;
assign _16520_ = _16616_ ^ _16624_ /*70753*/;
assign _16622_ = _16623_ | _16625_ /*70750*/;
assign _16627_ = ~Q[45] /*70749*/;
assign _16626_ = _16627_ & D[8] /*70748*/;
assign _16629_ = _16073_ & _16626_ /*70743*/;
assign _16630_ = _16073_ ^ _16626_ /*70746*/;
assign _16631_ = _16622_ & _16630_ /*70744*/;
assign _16521_ = _16622_ ^ _16630_ /*70745*/;
assign _16628_ = _16629_ | _16631_ /*70742*/;
assign _16633_ = ~Q[45] /*70741*/;
assign _16632_ = _16633_ & D[9] /*70740*/;
assign _16635_ = _16074_ & _16632_ /*70735*/;
assign _16636_ = _16074_ ^ _16632_ /*70738*/;
assign _16637_ = _16628_ & _16636_ /*70736*/;
assign _16522_ = _16628_ ^ _16636_ /*70737*/;
assign _16634_ = _16635_ | _16637_ /*70734*/;
assign _16639_ = ~Q[45] /*70733*/;
assign _16638_ = _16639_ & D[10] /*70732*/;
assign _16641_ = _16075_ & _16638_ /*70727*/;
assign _16642_ = _16075_ ^ _16638_ /*70730*/;
assign _16643_ = _16634_ & _16642_ /*70728*/;
assign _16523_ = _16634_ ^ _16642_ /*70729*/;
assign _16640_ = _16641_ | _16643_ /*70726*/;
assign _16645_ = ~Q[45] /*70725*/;
assign _16644_ = _16645_ & D[11] /*70724*/;
assign _16647_ = _16076_ & _16644_ /*70719*/;
assign _16648_ = _16076_ ^ _16644_ /*70722*/;
assign _16649_ = _16640_ & _16648_ /*70720*/;
assign _16524_ = _16640_ ^ _16648_ /*70721*/;
assign _16646_ = _16647_ | _16649_ /*70718*/;
assign _16651_ = ~Q[45] /*70717*/;
assign _16650_ = _16651_ & D[12] /*70716*/;
assign _16653_ = _16077_ & _16650_ /*70711*/;
assign _16654_ = _16077_ ^ _16650_ /*70714*/;
assign _16655_ = _16646_ & _16654_ /*70712*/;
assign _16525_ = _16646_ ^ _16654_ /*70713*/;
assign _16652_ = _16653_ | _16655_ /*70710*/;
assign _16657_ = ~Q[45] /*70709*/;
assign _16656_ = _16657_ & D[13] /*70708*/;
assign _16659_ = _16078_ & _16656_ /*70703*/;
assign _16660_ = _16078_ ^ _16656_ /*70706*/;
assign _16661_ = _16652_ & _16660_ /*70704*/;
assign _16526_ = _16652_ ^ _16660_ /*70705*/;
assign _16658_ = _16659_ | _16661_ /*70702*/;
assign _16663_ = ~Q[45] /*70701*/;
assign _16662_ = _16663_ & D[14] /*70700*/;
assign _16665_ = _16079_ & _16662_ /*70695*/;
assign _16666_ = _16079_ ^ _16662_ /*70698*/;
assign _16667_ = _16658_ & _16666_ /*70696*/;
assign _16527_ = _16658_ ^ _16666_ /*70697*/;
assign _16664_ = _16665_ | _16667_ /*70694*/;
assign _16669_ = ~Q[45] /*70693*/;
assign _16668_ = _16669_ & D[15] /*70692*/;
assign _16671_ = _16080_ & _16668_ /*70687*/;
assign _16672_ = _16080_ ^ _16668_ /*70690*/;
assign _16673_ = _16664_ & _16672_ /*70688*/;
assign _16528_ = _16664_ ^ _16672_ /*70689*/;
assign _16670_ = _16671_ | _16673_ /*70686*/;
assign _16675_ = ~Q[45] /*70685*/;
assign _16674_ = _16675_ & D[16] /*70684*/;
assign _16677_ = _16081_ & _16674_ /*70679*/;
assign _16678_ = _16081_ ^ _16674_ /*70682*/;
assign _16679_ = _16670_ & _16678_ /*70680*/;
assign _16529_ = _16670_ ^ _16678_ /*70681*/;
assign _16676_ = _16677_ | _16679_ /*70678*/;
assign _16681_ = ~Q[45] /*70677*/;
assign _16680_ = _16681_ & D[17] /*70676*/;
assign _16683_ = _16082_ & _16680_ /*70671*/;
assign _16684_ = _16082_ ^ _16680_ /*70674*/;
assign _16685_ = _16676_ & _16684_ /*70672*/;
assign _16530_ = _16676_ ^ _16684_ /*70673*/;
assign _16682_ = _16683_ | _16685_ /*70670*/;
assign _16687_ = ~Q[45] /*70669*/;
assign _16686_ = _16687_ & D[18] /*70668*/;
assign _16689_ = _16083_ & _16686_ /*70663*/;
assign _16690_ = _16083_ ^ _16686_ /*70666*/;
assign _16691_ = _16682_ & _16690_ /*70664*/;
assign _16531_ = _16682_ ^ _16690_ /*70665*/;
assign _16688_ = _16689_ | _16691_ /*70662*/;
assign _16693_ = ~Q[45] /*70661*/;
assign _16692_ = _16693_ & D[19] /*70660*/;
assign _16695_ = _16084_ & _16692_ /*70655*/;
assign _16696_ = _16084_ ^ _16692_ /*70658*/;
assign _16697_ = _16688_ & _16696_ /*70656*/;
assign _16532_ = _16688_ ^ _16696_ /*70657*/;
assign _16694_ = _16695_ | _16697_ /*70654*/;
assign _16699_ = ~Q[45] /*70653*/;
assign _16698_ = _16699_ & D[20] /*70652*/;
assign _16701_ = _16085_ & _16698_ /*70647*/;
assign _16702_ = _16085_ ^ _16698_ /*70650*/;
assign _16703_ = _16694_ & _16702_ /*70648*/;
assign _16533_ = _16694_ ^ _16702_ /*70649*/;
assign _16700_ = _16701_ | _16703_ /*70646*/;
assign _16705_ = ~Q[45] /*70645*/;
assign _16704_ = _16705_ & D[21] /*70644*/;
assign _16707_ = _16086_ & _16704_ /*70639*/;
assign _16708_ = _16086_ ^ _16704_ /*70642*/;
assign _16709_ = _16700_ & _16708_ /*70640*/;
assign _16534_ = _16700_ ^ _16708_ /*70641*/;
assign _16706_ = _16707_ | _16709_ /*70638*/;
assign _16711_ = ~Q[45] /*70637*/;
assign _16710_ = _16711_ & D[22] /*70636*/;
assign _16713_ = _16087_ & _16710_ /*70631*/;
assign _16714_ = _16087_ ^ _16710_ /*70634*/;
assign _16715_ = _16706_ & _16714_ /*70632*/;
assign _16535_ = _16706_ ^ _16714_ /*70633*/;
assign _16712_ = _16713_ | _16715_ /*70630*/;
assign _16717_ = ~Q[45] /*70629*/;
assign _16716_ = _16717_ & D[23] /*70628*/;
assign _16719_ = _16088_ & _16716_ /*70623*/;
assign _16720_ = _16088_ ^ _16716_ /*70626*/;
assign _16721_ = _16712_ & _16720_ /*70624*/;
assign _16536_ = _16712_ ^ _16720_ /*70625*/;
assign _16718_ = _16719_ | _16721_ /*70622*/;
assign _16723_ = ~Q[45] /*70621*/;
assign _16722_ = _16723_ & D[24] /*70620*/;
assign _16725_ = _16089_ & _16722_ /*70615*/;
assign _16726_ = _16089_ ^ _16722_ /*70618*/;
assign _16727_ = _16718_ & _16726_ /*70616*/;
assign _16537_ = _16718_ ^ _16726_ /*70617*/;
assign _16724_ = _16725_ | _16727_ /*70614*/;
assign _16729_ = ~Q[45] /*70613*/;
assign _16728_ = _16729_ & D[25] /*70612*/;
assign _16731_ = _16090_ & _16728_ /*70607*/;
assign _16732_ = _16090_ ^ _16728_ /*70610*/;
assign _16733_ = _16724_ & _16732_ /*70608*/;
assign _16538_ = _16724_ ^ _16732_ /*70609*/;
assign _16730_ = _16731_ | _16733_ /*70606*/;
assign _16735_ = ~Q[45] /*70605*/;
assign _16734_ = _16735_ & D[26] /*70604*/;
assign _16737_ = _16091_ & _16734_ /*70599*/;
assign _16738_ = _16091_ ^ _16734_ /*70602*/;
assign _16739_ = _16730_ & _16738_ /*70600*/;
assign _16539_ = _16730_ ^ _16738_ /*70601*/;
assign _16736_ = _16737_ | _16739_ /*70598*/;
assign _16741_ = ~Q[45] /*70597*/;
assign _16740_ = _16741_ & D[27] /*70596*/;
assign _16743_ = _16092_ & _16740_ /*70591*/;
assign _16744_ = _16092_ ^ _16740_ /*70594*/;
assign _16745_ = _16736_ & _16744_ /*70592*/;
assign _16540_ = _16736_ ^ _16744_ /*70593*/;
assign _16742_ = _16743_ | _16745_ /*70590*/;
assign _16747_ = ~Q[45] /*70589*/;
assign _16746_ = _16747_ & D[28] /*70588*/;
assign _16749_ = _16093_ & _16746_ /*70583*/;
assign _16750_ = _16093_ ^ _16746_ /*70586*/;
assign _16751_ = _16742_ & _16750_ /*70584*/;
assign _16541_ = _16742_ ^ _16750_ /*70585*/;
assign _16748_ = _16749_ | _16751_ /*70582*/;
assign _16753_ = ~Q[45] /*70581*/;
assign _16752_ = _16753_ & D[29] /*70580*/;
assign _16755_ = _16094_ & _16752_ /*70575*/;
assign _16756_ = _16094_ ^ _16752_ /*70578*/;
assign _16757_ = _16748_ & _16756_ /*70576*/;
assign _16542_ = _16748_ ^ _16756_ /*70577*/;
assign _16754_ = _16755_ | _16757_ /*70574*/;
assign _16759_ = ~Q[45] /*70573*/;
assign _16758_ = _16759_ & D[30] /*70572*/;
assign _16761_ = _16095_ & _16758_ /*70567*/;
assign _16762_ = _16095_ ^ _16758_ /*70570*/;
assign _16763_ = _16754_ & _16762_ /*70568*/;
assign _16543_ = _16754_ ^ _16762_ /*70569*/;
assign _16760_ = _16761_ | _16763_ /*70566*/;
assign _16765_ = ~Q[45] /*70565*/;
assign _16764_ = _16765_ & D[31] /*70564*/;
assign _16767_ = _16096_ & _16764_ /*70559*/;
assign _16768_ = _16096_ ^ _16764_ /*70562*/;
assign _16769_ = _16760_ & _16768_ /*70560*/;
assign _16544_ = _16760_ ^ _16768_ /*70561*/;
assign _16766_ = _16767_ | _16769_ /*70558*/;
assign _16771_ = ~Q[45] /*70557*/;
assign _16770_ = _16771_ & D[32] /*70556*/;
assign _16773_ = _16097_ & _16770_ /*70551*/;
assign _16774_ = _16097_ ^ _16770_ /*70554*/;
assign _16775_ = _16766_ & _16774_ /*70552*/;
assign _16545_ = _16766_ ^ _16774_ /*70553*/;
assign _16772_ = _16773_ | _16775_ /*70550*/;
assign _16777_ = ~Q[45] /*70549*/;
assign _16776_ = _16777_ & D[33] /*70548*/;
assign _16779_ = _16098_ & _16776_ /*70543*/;
assign _16780_ = _16098_ ^ _16776_ /*70546*/;
assign _16781_ = _16772_ & _16780_ /*70544*/;
assign _16546_ = _16772_ ^ _16780_ /*70545*/;
assign _16778_ = _16779_ | _16781_ /*70542*/;
assign _16783_ = ~Q[45] /*70541*/;
assign _16782_ = _16783_ & D[34] /*70540*/;
assign _16785_ = _16099_ & _16782_ /*70535*/;
assign _16786_ = _16099_ ^ _16782_ /*70538*/;
assign _16787_ = _16778_ & _16786_ /*70536*/;
assign _16547_ = _16778_ ^ _16786_ /*70537*/;
assign _16784_ = _16785_ | _16787_ /*70534*/;
assign _16789_ = ~Q[45] /*70533*/;
assign _16788_ = _16789_ & D[35] /*70532*/;
assign _16791_ = _16100_ & _16788_ /*70527*/;
assign _16792_ = _16100_ ^ _16788_ /*70530*/;
assign _16793_ = _16784_ & _16792_ /*70528*/;
assign _16548_ = _16784_ ^ _16792_ /*70529*/;
assign _16790_ = _16791_ | _16793_ /*70526*/;
assign _16795_ = ~Q[45] /*70525*/;
assign _16794_ = _16795_ & D[36] /*70524*/;
assign _16797_ = _16101_ & _16794_ /*70519*/;
assign _16798_ = _16101_ ^ _16794_ /*70522*/;
assign _16799_ = _16790_ & _16798_ /*70520*/;
assign _16549_ = _16790_ ^ _16798_ /*70521*/;
assign _16796_ = _16797_ | _16799_ /*70518*/;
assign _16801_ = ~Q[45] /*70517*/;
assign _16800_ = _16801_ & D[37] /*70516*/;
assign _16803_ = _16102_ & _16800_ /*70511*/;
assign _16804_ = _16102_ ^ _16800_ /*70514*/;
assign _16805_ = _16796_ & _16804_ /*70512*/;
assign _16550_ = _16796_ ^ _16804_ /*70513*/;
assign _16802_ = _16803_ | _16805_ /*70510*/;
assign _16807_ = ~Q[45] /*70509*/;
assign _16806_ = _16807_ & D[38] /*70508*/;
assign _16809_ = _16103_ & _16806_ /*70503*/;
assign _16810_ = _16103_ ^ _16806_ /*70506*/;
assign _16811_ = _16802_ & _16810_ /*70504*/;
assign _16551_ = _16802_ ^ _16810_ /*70505*/;
assign _16808_ = _16809_ | _16811_ /*70502*/;
assign _16813_ = ~Q[45] /*70501*/;
assign _16812_ = _16813_ & D[39] /*70500*/;
assign _16815_ = _16104_ & _16812_ /*70495*/;
assign _16816_ = _16104_ ^ _16812_ /*70498*/;
assign _16817_ = _16808_ & _16816_ /*70496*/;
assign _16552_ = _16808_ ^ _16816_ /*70497*/;
assign _16814_ = _16815_ | _16817_ /*70494*/;
assign _16819_ = ~Q[45] /*70493*/;
assign _16818_ = _16819_ & D[40] /*70492*/;
assign _16821_ = _16105_ & _16818_ /*70487*/;
assign _16822_ = _16105_ ^ _16818_ /*70490*/;
assign _16823_ = _16814_ & _16822_ /*70488*/;
assign _16553_ = _16814_ ^ _16822_ /*70489*/;
assign _16820_ = _16821_ | _16823_ /*70486*/;
assign _16825_ = ~Q[45] /*70485*/;
assign _16824_ = _16825_ & D[41] /*70484*/;
assign _16827_ = _16106_ & _16824_ /*70479*/;
assign _16828_ = _16106_ ^ _16824_ /*70482*/;
assign _16829_ = _16820_ & _16828_ /*70480*/;
assign _16554_ = _16820_ ^ _16828_ /*70481*/;
assign _16826_ = _16827_ | _16829_ /*70478*/;
assign _16831_ = ~Q[45] /*70477*/;
assign _16830_ = _16831_ & D[42] /*70476*/;
assign _16833_ = _16107_ & _16830_ /*70471*/;
assign _16834_ = _16107_ ^ _16830_ /*70474*/;
assign _16835_ = _16826_ & _16834_ /*70472*/;
assign _16555_ = _16826_ ^ _16834_ /*70473*/;
assign _16832_ = _16833_ | _16835_ /*70470*/;
assign _16837_ = ~Q[45] /*70469*/;
assign _16836_ = _16837_ & D[43] /*70468*/;
assign _16839_ = _16108_ & _16836_ /*70463*/;
assign _16840_ = _16108_ ^ _16836_ /*70466*/;
assign _16841_ = _16832_ & _16840_ /*70464*/;
assign _16556_ = _16832_ ^ _16840_ /*70465*/;
assign _16838_ = _16839_ | _16841_ /*70462*/;
assign _16843_ = ~Q[45] /*70461*/;
assign _16842_ = _16843_ & D[44] /*70460*/;
assign _16845_ = _16109_ & _16842_ /*70455*/;
assign _16846_ = _16109_ ^ _16842_ /*70458*/;
assign _16847_ = _16838_ & _16846_ /*70456*/;
assign _16557_ = _16838_ ^ _16846_ /*70457*/;
assign _16844_ = _16845_ | _16847_ /*70454*/;
assign _16849_ = ~Q[45] /*70453*/;
assign _16848_ = _16849_ & D[45] /*70452*/;
assign _16851_ = _16110_ & _16848_ /*70447*/;
assign _16852_ = _16110_ ^ _16848_ /*70450*/;
assign _16853_ = _16844_ & _16852_ /*70448*/;
assign _16558_ = _16844_ ^ _16852_ /*70449*/;
assign _16850_ = _16851_ | _16853_ /*70446*/;
assign _16855_ = ~Q[45] /*70445*/;
assign _16854_ = _16855_ & D[46] /*70444*/;
assign _16857_ = _16111_ & _16854_ /*70439*/;
assign _16858_ = _16111_ ^ _16854_ /*70442*/;
assign _16859_ = _16850_ & _16858_ /*70440*/;
assign _16559_ = _16850_ ^ _16858_ /*70441*/;
assign _16856_ = _16857_ | _16859_ /*70438*/;
assign _16861_ = ~Q[45] /*70437*/;
assign _16860_ = _16861_ & D[47] /*70436*/;
assign _16863_ = _16112_ & _16860_ /*70431*/;
assign _16864_ = _16112_ ^ _16860_ /*70434*/;
assign _16865_ = _16856_ & _16864_ /*70432*/;
assign _16560_ = _16856_ ^ _16864_ /*70433*/;
assign _16862_ = _16863_ | _16865_ /*70430*/;
assign _16867_ = ~Q[45] /*70429*/;
assign _16866_ = _16867_ & D[48] /*70428*/;
assign _16869_ = _16113_ & _16866_ /*70423*/;
assign _16870_ = _16113_ ^ _16866_ /*70426*/;
assign _16871_ = _16862_ & _16870_ /*70424*/;
assign _16561_ = _16862_ ^ _16870_ /*70425*/;
assign _16868_ = _16869_ | _16871_ /*70422*/;
assign _16873_ = ~Q[45] /*70421*/;
assign _16872_ = _16873_ & D[49] /*70420*/;
assign _16875_ = _16114_ & _16872_ /*70415*/;
assign _16876_ = _16114_ ^ _16872_ /*70418*/;
assign _16877_ = _16868_ & _16876_ /*70416*/;
assign _16562_ = _16868_ ^ _16876_ /*70417*/;
assign _16874_ = _16875_ | _16877_ /*70414*/;
assign _16879_ = ~Q[45] /*70413*/;
assign _16878_ = _16879_ & D[50] /*70412*/;
assign _16881_ = _16115_ & _16878_ /*70407*/;
assign _16882_ = _16115_ ^ _16878_ /*70410*/;
assign _16883_ = _16874_ & _16882_ /*70408*/;
assign _16563_ = _16874_ ^ _16882_ /*70409*/;
assign _16880_ = _16881_ | _16883_ /*70406*/;
assign _16885_ = ~Q[45] /*70405*/;
assign _16884_ = _16885_ & D[51] /*70404*/;
assign _16887_ = _16116_ & _16884_ /*70399*/;
assign _16888_ = _16116_ ^ _16884_ /*70402*/;
assign _16889_ = _16880_ & _16888_ /*70400*/;
assign _16564_ = _16880_ ^ _16888_ /*70401*/;
assign _16886_ = _16887_ | _16889_ /*70398*/;
assign _16891_ = ~Q[45] /*70397*/;
assign _16890_ = _16891_ & D[52] /*70396*/;
assign _16893_ = _16117_ & _16890_ /*70391*/;
assign _16894_ = _16117_ ^ _16890_ /*70394*/;
assign _16895_ = _16886_ & _16894_ /*70392*/;
assign _16565_ = _16886_ ^ _16894_ /*70393*/;
assign _16892_ = _16893_ | _16895_ /*70390*/;
assign _16897_ = ~Q[45] /*70389*/;
assign _16896_ = _16897_ & D[53] /*70388*/;
assign _16899_ = _16118_ & _16896_ /*70383*/;
assign _16900_ = _16118_ ^ _16896_ /*70386*/;
assign _16901_ = _16892_ & _16900_ /*70384*/;
assign _16566_ = _16892_ ^ _16900_ /*70385*/;
assign _16898_ = _16899_ | _16901_ /*70382*/;
assign _16903_ = ~Q[45] /*70381*/;
assign _16902_ = _16903_ & D[54] /*70380*/;
assign _16905_ = _16119_ & _16902_ /*70375*/;
assign _16906_ = _16119_ ^ _16902_ /*70378*/;
assign _16907_ = _16898_ & _16906_ /*70376*/;
assign _16567_ = _16898_ ^ _16906_ /*70377*/;
assign _16904_ = _16905_ | _16907_ /*70374*/;
assign _16909_ = ~Q[45] /*70373*/;
assign _16908_ = _16909_ & D[55] /*70372*/;
assign _16911_ = _16120_ & _16908_ /*70367*/;
assign _16912_ = _16120_ ^ _16908_ /*70370*/;
assign _16913_ = _16904_ & _16912_ /*70368*/;
assign _16568_ = _16904_ ^ _16912_ /*70369*/;
assign _16910_ = _16911_ | _16913_ /*70366*/;
assign _16915_ = ~Q[45] /*70365*/;
assign _16914_ = _16915_ & D[56] /*70364*/;
assign _16917_ = _16121_ & _16914_ /*70359*/;
assign _16918_ = _16121_ ^ _16914_ /*70362*/;
assign _16919_ = _16910_ & _16918_ /*70360*/;
assign _16569_ = _16910_ ^ _16918_ /*70361*/;
assign _16916_ = _16917_ | _16919_ /*70358*/;
assign _16921_ = ~Q[45] /*70357*/;
assign _16920_ = _16921_ & D[57] /*70356*/;
assign _16923_ = _16122_ & _16920_ /*70351*/;
assign _16924_ = _16122_ ^ _16920_ /*70354*/;
assign _16925_ = _16916_ & _16924_ /*70352*/;
assign _16570_ = _16916_ ^ _16924_ /*70353*/;
assign _16922_ = _16923_ | _16925_ /*70350*/;
assign _16927_ = ~Q[45] /*70349*/;
assign _16926_ = _16927_ & D[58] /*70348*/;
assign _16929_ = _16123_ & _16926_ /*70343*/;
assign _16930_ = _16123_ ^ _16926_ /*70346*/;
assign _16931_ = _16922_ & _16930_ /*70344*/;
assign _16571_ = _16922_ ^ _16930_ /*70345*/;
assign _16928_ = _16929_ | _16931_ /*70342*/;
assign _16933_ = ~Q[45] /*70341*/;
assign _16932_ = _16933_ & D[59] /*70340*/;
assign _16935_ = _16124_ & _16932_ /*70335*/;
assign _16936_ = _16124_ ^ _16932_ /*70338*/;
assign _16937_ = _16928_ & _16936_ /*70336*/;
assign _16572_ = _16928_ ^ _16936_ /*70337*/;
assign _16934_ = _16935_ | _16937_ /*70334*/;
assign _16939_ = ~Q[45] /*70333*/;
assign _16938_ = _16939_ & D[60] /*70332*/;
assign _16941_ = _16125_ & _16938_ /*70327*/;
assign _16942_ = _16125_ ^ _16938_ /*70330*/;
assign _16943_ = _16934_ & _16942_ /*70328*/;
assign _16573_ = _16934_ ^ _16942_ /*70329*/;
assign _16940_ = _16941_ | _16943_ /*70326*/;
assign _16945_ = ~Q[45] /*70325*/;
assign _16944_ = _16945_ & D[61] /*70324*/;
assign _16947_ = _16126_ & _16944_ /*70319*/;
assign _16948_ = _16126_ ^ _16944_ /*70322*/;
assign _16949_ = _16940_ & _16948_ /*70320*/;
assign _16574_ = _16940_ ^ _16948_ /*70321*/;
assign _16946_ = _16947_ | _16949_ /*70318*/;
assign _16951_ = ~Q[45] /*70317*/;
assign _16950_ = _16951_ & D[62] /*70316*/;
assign _16953_ = _16127_ & _16950_ /*70311*/;
assign _16954_ = _16127_ ^ _16950_ /*70314*/;
assign _16955_ = _16946_ & _16954_ /*70312*/;
assign _16575_ = _16946_ ^ _16954_ /*70313*/;
assign _16952_ = _16953_ | _16955_ /*70310*/;
assign _16957_ = ~Q[45] /*70309*/;
assign _16956_ = _16957_ & zeroWire /*70308*/;
assign _16958_ = _16128_ ^ _16956_ /*70306*/;
assign _16576_ = _16958_ ^ _16952_ /*70305*/;
assign _17029_ = ~D[0] /*70051*/;
assign _17026_ = R_0[44] & _17029_ /*70047*/;
assign _17027_ = R_0[44] ^ _17029_ /*70050*/;
assign _17028_ = oneWire & _17027_ /*70048*/;
assign _16961_ = oneWire ^ _17027_ /*70049*/;
assign _17025_ = _17026_ | _17028_ /*70046*/;
assign _17034_ = ~D[1] /*70045*/;
assign _17031_ = _16513_ & _17034_ /*70041*/;
assign _17032_ = _16513_ ^ _17034_ /*70044*/;
assign _17033_ = _17025_ & _17032_ /*70042*/;
assign _16962_ = _17025_ ^ _17032_ /*70043*/;
assign _17030_ = _17031_ | _17033_ /*70040*/;
assign _17039_ = ~D[2] /*70039*/;
assign _17036_ = _16514_ & _17039_ /*70035*/;
assign _17037_ = _16514_ ^ _17039_ /*70038*/;
assign _17038_ = _17030_ & _17037_ /*70036*/;
assign _16963_ = _17030_ ^ _17037_ /*70037*/;
assign _17035_ = _17036_ | _17038_ /*70034*/;
assign _17044_ = ~D[3] /*70033*/;
assign _17041_ = _16515_ & _17044_ /*70029*/;
assign _17042_ = _16515_ ^ _17044_ /*70032*/;
assign _17043_ = _17035_ & _17042_ /*70030*/;
assign _16964_ = _17035_ ^ _17042_ /*70031*/;
assign _17040_ = _17041_ | _17043_ /*70028*/;
assign _17049_ = ~D[4] /*70027*/;
assign _17046_ = _16516_ & _17049_ /*70023*/;
assign _17047_ = _16516_ ^ _17049_ /*70026*/;
assign _17048_ = _17040_ & _17047_ /*70024*/;
assign _16965_ = _17040_ ^ _17047_ /*70025*/;
assign _17045_ = _17046_ | _17048_ /*70022*/;
assign _17054_ = ~D[5] /*70021*/;
assign _17051_ = _16517_ & _17054_ /*70017*/;
assign _17052_ = _16517_ ^ _17054_ /*70020*/;
assign _17053_ = _17045_ & _17052_ /*70018*/;
assign _16966_ = _17045_ ^ _17052_ /*70019*/;
assign _17050_ = _17051_ | _17053_ /*70016*/;
assign _17059_ = ~D[6] /*70015*/;
assign _17056_ = _16518_ & _17059_ /*70011*/;
assign _17057_ = _16518_ ^ _17059_ /*70014*/;
assign _17058_ = _17050_ & _17057_ /*70012*/;
assign _16967_ = _17050_ ^ _17057_ /*70013*/;
assign _17055_ = _17056_ | _17058_ /*70010*/;
assign _17064_ = ~D[7] /*70009*/;
assign _17061_ = _16519_ & _17064_ /*70005*/;
assign _17062_ = _16519_ ^ _17064_ /*70008*/;
assign _17063_ = _17055_ & _17062_ /*70006*/;
assign _16968_ = _17055_ ^ _17062_ /*70007*/;
assign _17060_ = _17061_ | _17063_ /*70004*/;
assign _17069_ = ~D[8] /*70003*/;
assign _17066_ = _16520_ & _17069_ /*69999*/;
assign _17067_ = _16520_ ^ _17069_ /*70002*/;
assign _17068_ = _17060_ & _17067_ /*70000*/;
assign _16969_ = _17060_ ^ _17067_ /*70001*/;
assign _17065_ = _17066_ | _17068_ /*69998*/;
assign _17074_ = ~D[9] /*69997*/;
assign _17071_ = _16521_ & _17074_ /*69993*/;
assign _17072_ = _16521_ ^ _17074_ /*69996*/;
assign _17073_ = _17065_ & _17072_ /*69994*/;
assign _16970_ = _17065_ ^ _17072_ /*69995*/;
assign _17070_ = _17071_ | _17073_ /*69992*/;
assign _17079_ = ~D[10] /*69991*/;
assign _17076_ = _16522_ & _17079_ /*69987*/;
assign _17077_ = _16522_ ^ _17079_ /*69990*/;
assign _17078_ = _17070_ & _17077_ /*69988*/;
assign _16971_ = _17070_ ^ _17077_ /*69989*/;
assign _17075_ = _17076_ | _17078_ /*69986*/;
assign _17084_ = ~D[11] /*69985*/;
assign _17081_ = _16523_ & _17084_ /*69981*/;
assign _17082_ = _16523_ ^ _17084_ /*69984*/;
assign _17083_ = _17075_ & _17082_ /*69982*/;
assign _16972_ = _17075_ ^ _17082_ /*69983*/;
assign _17080_ = _17081_ | _17083_ /*69980*/;
assign _17089_ = ~D[12] /*69979*/;
assign _17086_ = _16524_ & _17089_ /*69975*/;
assign _17087_ = _16524_ ^ _17089_ /*69978*/;
assign _17088_ = _17080_ & _17087_ /*69976*/;
assign _16973_ = _17080_ ^ _17087_ /*69977*/;
assign _17085_ = _17086_ | _17088_ /*69974*/;
assign _17094_ = ~D[13] /*69973*/;
assign _17091_ = _16525_ & _17094_ /*69969*/;
assign _17092_ = _16525_ ^ _17094_ /*69972*/;
assign _17093_ = _17085_ & _17092_ /*69970*/;
assign _16974_ = _17085_ ^ _17092_ /*69971*/;
assign _17090_ = _17091_ | _17093_ /*69968*/;
assign _17099_ = ~D[14] /*69967*/;
assign _17096_ = _16526_ & _17099_ /*69963*/;
assign _17097_ = _16526_ ^ _17099_ /*69966*/;
assign _17098_ = _17090_ & _17097_ /*69964*/;
assign _16975_ = _17090_ ^ _17097_ /*69965*/;
assign _17095_ = _17096_ | _17098_ /*69962*/;
assign _17104_ = ~D[15] /*69961*/;
assign _17101_ = _16527_ & _17104_ /*69957*/;
assign _17102_ = _16527_ ^ _17104_ /*69960*/;
assign _17103_ = _17095_ & _17102_ /*69958*/;
assign _16976_ = _17095_ ^ _17102_ /*69959*/;
assign _17100_ = _17101_ | _17103_ /*69956*/;
assign _17109_ = ~D[16] /*69955*/;
assign _17106_ = _16528_ & _17109_ /*69951*/;
assign _17107_ = _16528_ ^ _17109_ /*69954*/;
assign _17108_ = _17100_ & _17107_ /*69952*/;
assign _16977_ = _17100_ ^ _17107_ /*69953*/;
assign _17105_ = _17106_ | _17108_ /*69950*/;
assign _17114_ = ~D[17] /*69949*/;
assign _17111_ = _16529_ & _17114_ /*69945*/;
assign _17112_ = _16529_ ^ _17114_ /*69948*/;
assign _17113_ = _17105_ & _17112_ /*69946*/;
assign _16978_ = _17105_ ^ _17112_ /*69947*/;
assign _17110_ = _17111_ | _17113_ /*69944*/;
assign _17119_ = ~D[18] /*69943*/;
assign _17116_ = _16530_ & _17119_ /*69939*/;
assign _17117_ = _16530_ ^ _17119_ /*69942*/;
assign _17118_ = _17110_ & _17117_ /*69940*/;
assign _16979_ = _17110_ ^ _17117_ /*69941*/;
assign _17115_ = _17116_ | _17118_ /*69938*/;
assign _17124_ = ~D[19] /*69937*/;
assign _17121_ = _16531_ & _17124_ /*69933*/;
assign _17122_ = _16531_ ^ _17124_ /*69936*/;
assign _17123_ = _17115_ & _17122_ /*69934*/;
assign _16980_ = _17115_ ^ _17122_ /*69935*/;
assign _17120_ = _17121_ | _17123_ /*69932*/;
assign _17129_ = ~D[20] /*69931*/;
assign _17126_ = _16532_ & _17129_ /*69927*/;
assign _17127_ = _16532_ ^ _17129_ /*69930*/;
assign _17128_ = _17120_ & _17127_ /*69928*/;
assign _16981_ = _17120_ ^ _17127_ /*69929*/;
assign _17125_ = _17126_ | _17128_ /*69926*/;
assign _17134_ = ~D[21] /*69925*/;
assign _17131_ = _16533_ & _17134_ /*69921*/;
assign _17132_ = _16533_ ^ _17134_ /*69924*/;
assign _17133_ = _17125_ & _17132_ /*69922*/;
assign _16982_ = _17125_ ^ _17132_ /*69923*/;
assign _17130_ = _17131_ | _17133_ /*69920*/;
assign _17139_ = ~D[22] /*69919*/;
assign _17136_ = _16534_ & _17139_ /*69915*/;
assign _17137_ = _16534_ ^ _17139_ /*69918*/;
assign _17138_ = _17130_ & _17137_ /*69916*/;
assign _16983_ = _17130_ ^ _17137_ /*69917*/;
assign _17135_ = _17136_ | _17138_ /*69914*/;
assign _17144_ = ~D[23] /*69913*/;
assign _17141_ = _16535_ & _17144_ /*69909*/;
assign _17142_ = _16535_ ^ _17144_ /*69912*/;
assign _17143_ = _17135_ & _17142_ /*69910*/;
assign _16984_ = _17135_ ^ _17142_ /*69911*/;
assign _17140_ = _17141_ | _17143_ /*69908*/;
assign _17149_ = ~D[24] /*69907*/;
assign _17146_ = _16536_ & _17149_ /*69903*/;
assign _17147_ = _16536_ ^ _17149_ /*69906*/;
assign _17148_ = _17140_ & _17147_ /*69904*/;
assign _16985_ = _17140_ ^ _17147_ /*69905*/;
assign _17145_ = _17146_ | _17148_ /*69902*/;
assign _17154_ = ~D[25] /*69901*/;
assign _17151_ = _16537_ & _17154_ /*69897*/;
assign _17152_ = _16537_ ^ _17154_ /*69900*/;
assign _17153_ = _17145_ & _17152_ /*69898*/;
assign _16986_ = _17145_ ^ _17152_ /*69899*/;
assign _17150_ = _17151_ | _17153_ /*69896*/;
assign _17159_ = ~D[26] /*69895*/;
assign _17156_ = _16538_ & _17159_ /*69891*/;
assign _17157_ = _16538_ ^ _17159_ /*69894*/;
assign _17158_ = _17150_ & _17157_ /*69892*/;
assign _16987_ = _17150_ ^ _17157_ /*69893*/;
assign _17155_ = _17156_ | _17158_ /*69890*/;
assign _17164_ = ~D[27] /*69889*/;
assign _17161_ = _16539_ & _17164_ /*69885*/;
assign _17162_ = _16539_ ^ _17164_ /*69888*/;
assign _17163_ = _17155_ & _17162_ /*69886*/;
assign _16988_ = _17155_ ^ _17162_ /*69887*/;
assign _17160_ = _17161_ | _17163_ /*69884*/;
assign _17169_ = ~D[28] /*69883*/;
assign _17166_ = _16540_ & _17169_ /*69879*/;
assign _17167_ = _16540_ ^ _17169_ /*69882*/;
assign _17168_ = _17160_ & _17167_ /*69880*/;
assign _16989_ = _17160_ ^ _17167_ /*69881*/;
assign _17165_ = _17166_ | _17168_ /*69878*/;
assign _17174_ = ~D[29] /*69877*/;
assign _17171_ = _16541_ & _17174_ /*69873*/;
assign _17172_ = _16541_ ^ _17174_ /*69876*/;
assign _17173_ = _17165_ & _17172_ /*69874*/;
assign _16990_ = _17165_ ^ _17172_ /*69875*/;
assign _17170_ = _17171_ | _17173_ /*69872*/;
assign _17179_ = ~D[30] /*69871*/;
assign _17176_ = _16542_ & _17179_ /*69867*/;
assign _17177_ = _16542_ ^ _17179_ /*69870*/;
assign _17178_ = _17170_ & _17177_ /*69868*/;
assign _16991_ = _17170_ ^ _17177_ /*69869*/;
assign _17175_ = _17176_ | _17178_ /*69866*/;
assign _17184_ = ~D[31] /*69865*/;
assign _17181_ = _16543_ & _17184_ /*69861*/;
assign _17182_ = _16543_ ^ _17184_ /*69864*/;
assign _17183_ = _17175_ & _17182_ /*69862*/;
assign _16992_ = _17175_ ^ _17182_ /*69863*/;
assign _17180_ = _17181_ | _17183_ /*69860*/;
assign _17189_ = ~D[32] /*69859*/;
assign _17186_ = _16544_ & _17189_ /*69855*/;
assign _17187_ = _16544_ ^ _17189_ /*69858*/;
assign _17188_ = _17180_ & _17187_ /*69856*/;
assign _16993_ = _17180_ ^ _17187_ /*69857*/;
assign _17185_ = _17186_ | _17188_ /*69854*/;
assign _17194_ = ~D[33] /*69853*/;
assign _17191_ = _16545_ & _17194_ /*69849*/;
assign _17192_ = _16545_ ^ _17194_ /*69852*/;
assign _17193_ = _17185_ & _17192_ /*69850*/;
assign _16994_ = _17185_ ^ _17192_ /*69851*/;
assign _17190_ = _17191_ | _17193_ /*69848*/;
assign _17199_ = ~D[34] /*69847*/;
assign _17196_ = _16546_ & _17199_ /*69843*/;
assign _17197_ = _16546_ ^ _17199_ /*69846*/;
assign _17198_ = _17190_ & _17197_ /*69844*/;
assign _16995_ = _17190_ ^ _17197_ /*69845*/;
assign _17195_ = _17196_ | _17198_ /*69842*/;
assign _17204_ = ~D[35] /*69841*/;
assign _17201_ = _16547_ & _17204_ /*69837*/;
assign _17202_ = _16547_ ^ _17204_ /*69840*/;
assign _17203_ = _17195_ & _17202_ /*69838*/;
assign _16996_ = _17195_ ^ _17202_ /*69839*/;
assign _17200_ = _17201_ | _17203_ /*69836*/;
assign _17209_ = ~D[36] /*69835*/;
assign _17206_ = _16548_ & _17209_ /*69831*/;
assign _17207_ = _16548_ ^ _17209_ /*69834*/;
assign _17208_ = _17200_ & _17207_ /*69832*/;
assign _16997_ = _17200_ ^ _17207_ /*69833*/;
assign _17205_ = _17206_ | _17208_ /*69830*/;
assign _17214_ = ~D[37] /*69829*/;
assign _17211_ = _16549_ & _17214_ /*69825*/;
assign _17212_ = _16549_ ^ _17214_ /*69828*/;
assign _17213_ = _17205_ & _17212_ /*69826*/;
assign _16998_ = _17205_ ^ _17212_ /*69827*/;
assign _17210_ = _17211_ | _17213_ /*69824*/;
assign _17219_ = ~D[38] /*69823*/;
assign _17216_ = _16550_ & _17219_ /*69819*/;
assign _17217_ = _16550_ ^ _17219_ /*69822*/;
assign _17218_ = _17210_ & _17217_ /*69820*/;
assign _16999_ = _17210_ ^ _17217_ /*69821*/;
assign _17215_ = _17216_ | _17218_ /*69818*/;
assign _17224_ = ~D[39] /*69817*/;
assign _17221_ = _16551_ & _17224_ /*69813*/;
assign _17222_ = _16551_ ^ _17224_ /*69816*/;
assign _17223_ = _17215_ & _17222_ /*69814*/;
assign _17000_ = _17215_ ^ _17222_ /*69815*/;
assign _17220_ = _17221_ | _17223_ /*69812*/;
assign _17229_ = ~D[40] /*69811*/;
assign _17226_ = _16552_ & _17229_ /*69807*/;
assign _17227_ = _16552_ ^ _17229_ /*69810*/;
assign _17228_ = _17220_ & _17227_ /*69808*/;
assign _17001_ = _17220_ ^ _17227_ /*69809*/;
assign _17225_ = _17226_ | _17228_ /*69806*/;
assign _17234_ = ~D[41] /*69805*/;
assign _17231_ = _16553_ & _17234_ /*69801*/;
assign _17232_ = _16553_ ^ _17234_ /*69804*/;
assign _17233_ = _17225_ & _17232_ /*69802*/;
assign _17002_ = _17225_ ^ _17232_ /*69803*/;
assign _17230_ = _17231_ | _17233_ /*69800*/;
assign _17239_ = ~D[42] /*69799*/;
assign _17236_ = _16554_ & _17239_ /*69795*/;
assign _17237_ = _16554_ ^ _17239_ /*69798*/;
assign _17238_ = _17230_ & _17237_ /*69796*/;
assign _17003_ = _17230_ ^ _17237_ /*69797*/;
assign _17235_ = _17236_ | _17238_ /*69794*/;
assign _17244_ = ~D[43] /*69793*/;
assign _17241_ = _16555_ & _17244_ /*69789*/;
assign _17242_ = _16555_ ^ _17244_ /*69792*/;
assign _17243_ = _17235_ & _17242_ /*69790*/;
assign _17004_ = _17235_ ^ _17242_ /*69791*/;
assign _17240_ = _17241_ | _17243_ /*69788*/;
assign _17249_ = ~D[44] /*69787*/;
assign _17246_ = _16556_ & _17249_ /*69783*/;
assign _17247_ = _16556_ ^ _17249_ /*69786*/;
assign _17248_ = _17240_ & _17247_ /*69784*/;
assign _17005_ = _17240_ ^ _17247_ /*69785*/;
assign _17245_ = _17246_ | _17248_ /*69782*/;
assign _17254_ = ~D[45] /*69781*/;
assign _17251_ = _16557_ & _17254_ /*69777*/;
assign _17252_ = _16557_ ^ _17254_ /*69780*/;
assign _17253_ = _17245_ & _17252_ /*69778*/;
assign _17006_ = _17245_ ^ _17252_ /*69779*/;
assign _17250_ = _17251_ | _17253_ /*69776*/;
assign _17259_ = ~D[46] /*69775*/;
assign _17256_ = _16558_ & _17259_ /*69771*/;
assign _17257_ = _16558_ ^ _17259_ /*69774*/;
assign _17258_ = _17250_ & _17257_ /*69772*/;
assign _17007_ = _17250_ ^ _17257_ /*69773*/;
assign _17255_ = _17256_ | _17258_ /*69770*/;
assign _17264_ = ~D[47] /*69769*/;
assign _17261_ = _16559_ & _17264_ /*69765*/;
assign _17262_ = _16559_ ^ _17264_ /*69768*/;
assign _17263_ = _17255_ & _17262_ /*69766*/;
assign _17008_ = _17255_ ^ _17262_ /*69767*/;
assign _17260_ = _17261_ | _17263_ /*69764*/;
assign _17269_ = ~D[48] /*69763*/;
assign _17266_ = _16560_ & _17269_ /*69759*/;
assign _17267_ = _16560_ ^ _17269_ /*69762*/;
assign _17268_ = _17260_ & _17267_ /*69760*/;
assign _17009_ = _17260_ ^ _17267_ /*69761*/;
assign _17265_ = _17266_ | _17268_ /*69758*/;
assign _17274_ = ~D[49] /*69757*/;
assign _17271_ = _16561_ & _17274_ /*69753*/;
assign _17272_ = _16561_ ^ _17274_ /*69756*/;
assign _17273_ = _17265_ & _17272_ /*69754*/;
assign _17010_ = _17265_ ^ _17272_ /*69755*/;
assign _17270_ = _17271_ | _17273_ /*69752*/;
assign _17279_ = ~D[50] /*69751*/;
assign _17276_ = _16562_ & _17279_ /*69747*/;
assign _17277_ = _16562_ ^ _17279_ /*69750*/;
assign _17278_ = _17270_ & _17277_ /*69748*/;
assign _17011_ = _17270_ ^ _17277_ /*69749*/;
assign _17275_ = _17276_ | _17278_ /*69746*/;
assign _17284_ = ~D[51] /*69745*/;
assign _17281_ = _16563_ & _17284_ /*69741*/;
assign _17282_ = _16563_ ^ _17284_ /*69744*/;
assign _17283_ = _17275_ & _17282_ /*69742*/;
assign _17012_ = _17275_ ^ _17282_ /*69743*/;
assign _17280_ = _17281_ | _17283_ /*69740*/;
assign _17289_ = ~D[52] /*69739*/;
assign _17286_ = _16564_ & _17289_ /*69735*/;
assign _17287_ = _16564_ ^ _17289_ /*69738*/;
assign _17288_ = _17280_ & _17287_ /*69736*/;
assign _17013_ = _17280_ ^ _17287_ /*69737*/;
assign _17285_ = _17286_ | _17288_ /*69734*/;
assign _17294_ = ~D[53] /*69733*/;
assign _17291_ = _16565_ & _17294_ /*69729*/;
assign _17292_ = _16565_ ^ _17294_ /*69732*/;
assign _17293_ = _17285_ & _17292_ /*69730*/;
assign _17014_ = _17285_ ^ _17292_ /*69731*/;
assign _17290_ = _17291_ | _17293_ /*69728*/;
assign _17299_ = ~D[54] /*69727*/;
assign _17296_ = _16566_ & _17299_ /*69723*/;
assign _17297_ = _16566_ ^ _17299_ /*69726*/;
assign _17298_ = _17290_ & _17297_ /*69724*/;
assign _17015_ = _17290_ ^ _17297_ /*69725*/;
assign _17295_ = _17296_ | _17298_ /*69722*/;
assign _17304_ = ~D[55] /*69721*/;
assign _17301_ = _16567_ & _17304_ /*69717*/;
assign _17302_ = _16567_ ^ _17304_ /*69720*/;
assign _17303_ = _17295_ & _17302_ /*69718*/;
assign _17016_ = _17295_ ^ _17302_ /*69719*/;
assign _17300_ = _17301_ | _17303_ /*69716*/;
assign _17309_ = ~D[56] /*69715*/;
assign _17306_ = _16568_ & _17309_ /*69711*/;
assign _17307_ = _16568_ ^ _17309_ /*69714*/;
assign _17308_ = _17300_ & _17307_ /*69712*/;
assign _17017_ = _17300_ ^ _17307_ /*69713*/;
assign _17305_ = _17306_ | _17308_ /*69710*/;
assign _17314_ = ~D[57] /*69709*/;
assign _17311_ = _16569_ & _17314_ /*69705*/;
assign _17312_ = _16569_ ^ _17314_ /*69708*/;
assign _17313_ = _17305_ & _17312_ /*69706*/;
assign _17018_ = _17305_ ^ _17312_ /*69707*/;
assign _17310_ = _17311_ | _17313_ /*69704*/;
assign _17319_ = ~D[58] /*69703*/;
assign _17316_ = _16570_ & _17319_ /*69699*/;
assign _17317_ = _16570_ ^ _17319_ /*69702*/;
assign _17318_ = _17310_ & _17317_ /*69700*/;
assign _17019_ = _17310_ ^ _17317_ /*69701*/;
assign _17315_ = _17316_ | _17318_ /*69698*/;
assign _17324_ = ~D[59] /*69697*/;
assign _17321_ = _16571_ & _17324_ /*69693*/;
assign _17322_ = _16571_ ^ _17324_ /*69696*/;
assign _17323_ = _17315_ & _17322_ /*69694*/;
assign _17020_ = _17315_ ^ _17322_ /*69695*/;
assign _17320_ = _17321_ | _17323_ /*69692*/;
assign _17329_ = ~D[60] /*69691*/;
assign _17326_ = _16572_ & _17329_ /*69687*/;
assign _17327_ = _16572_ ^ _17329_ /*69690*/;
assign _17328_ = _17320_ & _17327_ /*69688*/;
assign _17021_ = _17320_ ^ _17327_ /*69689*/;
assign _17325_ = _17326_ | _17328_ /*69686*/;
assign _17334_ = ~D[61] /*69685*/;
assign _17331_ = _16573_ & _17334_ /*69681*/;
assign _17332_ = _16573_ ^ _17334_ /*69684*/;
assign _17333_ = _17325_ & _17332_ /*69682*/;
assign _17022_ = _17325_ ^ _17332_ /*69683*/;
assign _17330_ = _17331_ | _17333_ /*69680*/;
assign _17339_ = ~D[62] /*69679*/;
assign _17336_ = _16574_ & _17339_ /*69675*/;
assign _17337_ = _16574_ ^ _17339_ /*69678*/;
assign _17338_ = _17330_ & _17337_ /*69676*/;
assign _17023_ = _17330_ ^ _17337_ /*69677*/;
assign _17335_ = _17336_ | _17338_ /*69674*/;
assign _17340_ = _16575_ & oneWire /*69669*/;
assign _17341_ = _16575_ ^ oneWire /*69672*/;
assign _17342_ = _17335_ & _17341_ /*69670*/;
assign _17024_ = _17335_ ^ _17341_ /*69671*/;
assign Q[44] = _17340_ | _17342_ /*69668*/;
assign _17475_ = ~Q[44] /*69283*/;
assign _17474_ = _17475_ & D[0] /*69282*/;
assign _17477_ = _16961_ & _17474_ /*69277*/;
assign _17478_ = _16961_ ^ _17474_ /*69280*/;
assign _17479_ = zeroWire & _17478_ /*69278*/;
assign _17409_ = zeroWire ^ _17478_ /*69279*/;
assign _17476_ = _17477_ | _17479_ /*69276*/;
assign _17481_ = ~Q[44] /*69275*/;
assign _17480_ = _17481_ & D[1] /*69274*/;
assign _17483_ = _16962_ & _17480_ /*69269*/;
assign _17484_ = _16962_ ^ _17480_ /*69272*/;
assign _17485_ = _17476_ & _17484_ /*69270*/;
assign _17410_ = _17476_ ^ _17484_ /*69271*/;
assign _17482_ = _17483_ | _17485_ /*69268*/;
assign _17487_ = ~Q[44] /*69267*/;
assign _17486_ = _17487_ & D[2] /*69266*/;
assign _17489_ = _16963_ & _17486_ /*69261*/;
assign _17490_ = _16963_ ^ _17486_ /*69264*/;
assign _17491_ = _17482_ & _17490_ /*69262*/;
assign _17411_ = _17482_ ^ _17490_ /*69263*/;
assign _17488_ = _17489_ | _17491_ /*69260*/;
assign _17493_ = ~Q[44] /*69259*/;
assign _17492_ = _17493_ & D[3] /*69258*/;
assign _17495_ = _16964_ & _17492_ /*69253*/;
assign _17496_ = _16964_ ^ _17492_ /*69256*/;
assign _17497_ = _17488_ & _17496_ /*69254*/;
assign _17412_ = _17488_ ^ _17496_ /*69255*/;
assign _17494_ = _17495_ | _17497_ /*69252*/;
assign _17499_ = ~Q[44] /*69251*/;
assign _17498_ = _17499_ & D[4] /*69250*/;
assign _17501_ = _16965_ & _17498_ /*69245*/;
assign _17502_ = _16965_ ^ _17498_ /*69248*/;
assign _17503_ = _17494_ & _17502_ /*69246*/;
assign _17413_ = _17494_ ^ _17502_ /*69247*/;
assign _17500_ = _17501_ | _17503_ /*69244*/;
assign _17505_ = ~Q[44] /*69243*/;
assign _17504_ = _17505_ & D[5] /*69242*/;
assign _17507_ = _16966_ & _17504_ /*69237*/;
assign _17508_ = _16966_ ^ _17504_ /*69240*/;
assign _17509_ = _17500_ & _17508_ /*69238*/;
assign _17414_ = _17500_ ^ _17508_ /*69239*/;
assign _17506_ = _17507_ | _17509_ /*69236*/;
assign _17511_ = ~Q[44] /*69235*/;
assign _17510_ = _17511_ & D[6] /*69234*/;
assign _17513_ = _16967_ & _17510_ /*69229*/;
assign _17514_ = _16967_ ^ _17510_ /*69232*/;
assign _17515_ = _17506_ & _17514_ /*69230*/;
assign _17415_ = _17506_ ^ _17514_ /*69231*/;
assign _17512_ = _17513_ | _17515_ /*69228*/;
assign _17517_ = ~Q[44] /*69227*/;
assign _17516_ = _17517_ & D[7] /*69226*/;
assign _17519_ = _16968_ & _17516_ /*69221*/;
assign _17520_ = _16968_ ^ _17516_ /*69224*/;
assign _17521_ = _17512_ & _17520_ /*69222*/;
assign _17416_ = _17512_ ^ _17520_ /*69223*/;
assign _17518_ = _17519_ | _17521_ /*69220*/;
assign _17523_ = ~Q[44] /*69219*/;
assign _17522_ = _17523_ & D[8] /*69218*/;
assign _17525_ = _16969_ & _17522_ /*69213*/;
assign _17526_ = _16969_ ^ _17522_ /*69216*/;
assign _17527_ = _17518_ & _17526_ /*69214*/;
assign _17417_ = _17518_ ^ _17526_ /*69215*/;
assign _17524_ = _17525_ | _17527_ /*69212*/;
assign _17529_ = ~Q[44] /*69211*/;
assign _17528_ = _17529_ & D[9] /*69210*/;
assign _17531_ = _16970_ & _17528_ /*69205*/;
assign _17532_ = _16970_ ^ _17528_ /*69208*/;
assign _17533_ = _17524_ & _17532_ /*69206*/;
assign _17418_ = _17524_ ^ _17532_ /*69207*/;
assign _17530_ = _17531_ | _17533_ /*69204*/;
assign _17535_ = ~Q[44] /*69203*/;
assign _17534_ = _17535_ & D[10] /*69202*/;
assign _17537_ = _16971_ & _17534_ /*69197*/;
assign _17538_ = _16971_ ^ _17534_ /*69200*/;
assign _17539_ = _17530_ & _17538_ /*69198*/;
assign _17419_ = _17530_ ^ _17538_ /*69199*/;
assign _17536_ = _17537_ | _17539_ /*69196*/;
assign _17541_ = ~Q[44] /*69195*/;
assign _17540_ = _17541_ & D[11] /*69194*/;
assign _17543_ = _16972_ & _17540_ /*69189*/;
assign _17544_ = _16972_ ^ _17540_ /*69192*/;
assign _17545_ = _17536_ & _17544_ /*69190*/;
assign _17420_ = _17536_ ^ _17544_ /*69191*/;
assign _17542_ = _17543_ | _17545_ /*69188*/;
assign _17547_ = ~Q[44] /*69187*/;
assign _17546_ = _17547_ & D[12] /*69186*/;
assign _17549_ = _16973_ & _17546_ /*69181*/;
assign _17550_ = _16973_ ^ _17546_ /*69184*/;
assign _17551_ = _17542_ & _17550_ /*69182*/;
assign _17421_ = _17542_ ^ _17550_ /*69183*/;
assign _17548_ = _17549_ | _17551_ /*69180*/;
assign _17553_ = ~Q[44] /*69179*/;
assign _17552_ = _17553_ & D[13] /*69178*/;
assign _17555_ = _16974_ & _17552_ /*69173*/;
assign _17556_ = _16974_ ^ _17552_ /*69176*/;
assign _17557_ = _17548_ & _17556_ /*69174*/;
assign _17422_ = _17548_ ^ _17556_ /*69175*/;
assign _17554_ = _17555_ | _17557_ /*69172*/;
assign _17559_ = ~Q[44] /*69171*/;
assign _17558_ = _17559_ & D[14] /*69170*/;
assign _17561_ = _16975_ & _17558_ /*69165*/;
assign _17562_ = _16975_ ^ _17558_ /*69168*/;
assign _17563_ = _17554_ & _17562_ /*69166*/;
assign _17423_ = _17554_ ^ _17562_ /*69167*/;
assign _17560_ = _17561_ | _17563_ /*69164*/;
assign _17565_ = ~Q[44] /*69163*/;
assign _17564_ = _17565_ & D[15] /*69162*/;
assign _17567_ = _16976_ & _17564_ /*69157*/;
assign _17568_ = _16976_ ^ _17564_ /*69160*/;
assign _17569_ = _17560_ & _17568_ /*69158*/;
assign _17424_ = _17560_ ^ _17568_ /*69159*/;
assign _17566_ = _17567_ | _17569_ /*69156*/;
assign _17571_ = ~Q[44] /*69155*/;
assign _17570_ = _17571_ & D[16] /*69154*/;
assign _17573_ = _16977_ & _17570_ /*69149*/;
assign _17574_ = _16977_ ^ _17570_ /*69152*/;
assign _17575_ = _17566_ & _17574_ /*69150*/;
assign _17425_ = _17566_ ^ _17574_ /*69151*/;
assign _17572_ = _17573_ | _17575_ /*69148*/;
assign _17577_ = ~Q[44] /*69147*/;
assign _17576_ = _17577_ & D[17] /*69146*/;
assign _17579_ = _16978_ & _17576_ /*69141*/;
assign _17580_ = _16978_ ^ _17576_ /*69144*/;
assign _17581_ = _17572_ & _17580_ /*69142*/;
assign _17426_ = _17572_ ^ _17580_ /*69143*/;
assign _17578_ = _17579_ | _17581_ /*69140*/;
assign _17583_ = ~Q[44] /*69139*/;
assign _17582_ = _17583_ & D[18] /*69138*/;
assign _17585_ = _16979_ & _17582_ /*69133*/;
assign _17586_ = _16979_ ^ _17582_ /*69136*/;
assign _17587_ = _17578_ & _17586_ /*69134*/;
assign _17427_ = _17578_ ^ _17586_ /*69135*/;
assign _17584_ = _17585_ | _17587_ /*69132*/;
assign _17589_ = ~Q[44] /*69131*/;
assign _17588_ = _17589_ & D[19] /*69130*/;
assign _17591_ = _16980_ & _17588_ /*69125*/;
assign _17592_ = _16980_ ^ _17588_ /*69128*/;
assign _17593_ = _17584_ & _17592_ /*69126*/;
assign _17428_ = _17584_ ^ _17592_ /*69127*/;
assign _17590_ = _17591_ | _17593_ /*69124*/;
assign _17595_ = ~Q[44] /*69123*/;
assign _17594_ = _17595_ & D[20] /*69122*/;
assign _17597_ = _16981_ & _17594_ /*69117*/;
assign _17598_ = _16981_ ^ _17594_ /*69120*/;
assign _17599_ = _17590_ & _17598_ /*69118*/;
assign _17429_ = _17590_ ^ _17598_ /*69119*/;
assign _17596_ = _17597_ | _17599_ /*69116*/;
assign _17601_ = ~Q[44] /*69115*/;
assign _17600_ = _17601_ & D[21] /*69114*/;
assign _17603_ = _16982_ & _17600_ /*69109*/;
assign _17604_ = _16982_ ^ _17600_ /*69112*/;
assign _17605_ = _17596_ & _17604_ /*69110*/;
assign _17430_ = _17596_ ^ _17604_ /*69111*/;
assign _17602_ = _17603_ | _17605_ /*69108*/;
assign _17607_ = ~Q[44] /*69107*/;
assign _17606_ = _17607_ & D[22] /*69106*/;
assign _17609_ = _16983_ & _17606_ /*69101*/;
assign _17610_ = _16983_ ^ _17606_ /*69104*/;
assign _17611_ = _17602_ & _17610_ /*69102*/;
assign _17431_ = _17602_ ^ _17610_ /*69103*/;
assign _17608_ = _17609_ | _17611_ /*69100*/;
assign _17613_ = ~Q[44] /*69099*/;
assign _17612_ = _17613_ & D[23] /*69098*/;
assign _17615_ = _16984_ & _17612_ /*69093*/;
assign _17616_ = _16984_ ^ _17612_ /*69096*/;
assign _17617_ = _17608_ & _17616_ /*69094*/;
assign _17432_ = _17608_ ^ _17616_ /*69095*/;
assign _17614_ = _17615_ | _17617_ /*69092*/;
assign _17619_ = ~Q[44] /*69091*/;
assign _17618_ = _17619_ & D[24] /*69090*/;
assign _17621_ = _16985_ & _17618_ /*69085*/;
assign _17622_ = _16985_ ^ _17618_ /*69088*/;
assign _17623_ = _17614_ & _17622_ /*69086*/;
assign _17433_ = _17614_ ^ _17622_ /*69087*/;
assign _17620_ = _17621_ | _17623_ /*69084*/;
assign _17625_ = ~Q[44] /*69083*/;
assign _17624_ = _17625_ & D[25] /*69082*/;
assign _17627_ = _16986_ & _17624_ /*69077*/;
assign _17628_ = _16986_ ^ _17624_ /*69080*/;
assign _17629_ = _17620_ & _17628_ /*69078*/;
assign _17434_ = _17620_ ^ _17628_ /*69079*/;
assign _17626_ = _17627_ | _17629_ /*69076*/;
assign _17631_ = ~Q[44] /*69075*/;
assign _17630_ = _17631_ & D[26] /*69074*/;
assign _17633_ = _16987_ & _17630_ /*69069*/;
assign _17634_ = _16987_ ^ _17630_ /*69072*/;
assign _17635_ = _17626_ & _17634_ /*69070*/;
assign _17435_ = _17626_ ^ _17634_ /*69071*/;
assign _17632_ = _17633_ | _17635_ /*69068*/;
assign _17637_ = ~Q[44] /*69067*/;
assign _17636_ = _17637_ & D[27] /*69066*/;
assign _17639_ = _16988_ & _17636_ /*69061*/;
assign _17640_ = _16988_ ^ _17636_ /*69064*/;
assign _17641_ = _17632_ & _17640_ /*69062*/;
assign _17436_ = _17632_ ^ _17640_ /*69063*/;
assign _17638_ = _17639_ | _17641_ /*69060*/;
assign _17643_ = ~Q[44] /*69059*/;
assign _17642_ = _17643_ & D[28] /*69058*/;
assign _17645_ = _16989_ & _17642_ /*69053*/;
assign _17646_ = _16989_ ^ _17642_ /*69056*/;
assign _17647_ = _17638_ & _17646_ /*69054*/;
assign _17437_ = _17638_ ^ _17646_ /*69055*/;
assign _17644_ = _17645_ | _17647_ /*69052*/;
assign _17649_ = ~Q[44] /*69051*/;
assign _17648_ = _17649_ & D[29] /*69050*/;
assign _17651_ = _16990_ & _17648_ /*69045*/;
assign _17652_ = _16990_ ^ _17648_ /*69048*/;
assign _17653_ = _17644_ & _17652_ /*69046*/;
assign _17438_ = _17644_ ^ _17652_ /*69047*/;
assign _17650_ = _17651_ | _17653_ /*69044*/;
assign _17655_ = ~Q[44] /*69043*/;
assign _17654_ = _17655_ & D[30] /*69042*/;
assign _17657_ = _16991_ & _17654_ /*69037*/;
assign _17658_ = _16991_ ^ _17654_ /*69040*/;
assign _17659_ = _17650_ & _17658_ /*69038*/;
assign _17439_ = _17650_ ^ _17658_ /*69039*/;
assign _17656_ = _17657_ | _17659_ /*69036*/;
assign _17661_ = ~Q[44] /*69035*/;
assign _17660_ = _17661_ & D[31] /*69034*/;
assign _17663_ = _16992_ & _17660_ /*69029*/;
assign _17664_ = _16992_ ^ _17660_ /*69032*/;
assign _17665_ = _17656_ & _17664_ /*69030*/;
assign _17440_ = _17656_ ^ _17664_ /*69031*/;
assign _17662_ = _17663_ | _17665_ /*69028*/;
assign _17667_ = ~Q[44] /*69027*/;
assign _17666_ = _17667_ & D[32] /*69026*/;
assign _17669_ = _16993_ & _17666_ /*69021*/;
assign _17670_ = _16993_ ^ _17666_ /*69024*/;
assign _17671_ = _17662_ & _17670_ /*69022*/;
assign _17441_ = _17662_ ^ _17670_ /*69023*/;
assign _17668_ = _17669_ | _17671_ /*69020*/;
assign _17673_ = ~Q[44] /*69019*/;
assign _17672_ = _17673_ & D[33] /*69018*/;
assign _17675_ = _16994_ & _17672_ /*69013*/;
assign _17676_ = _16994_ ^ _17672_ /*69016*/;
assign _17677_ = _17668_ & _17676_ /*69014*/;
assign _17442_ = _17668_ ^ _17676_ /*69015*/;
assign _17674_ = _17675_ | _17677_ /*69012*/;
assign _17679_ = ~Q[44] /*69011*/;
assign _17678_ = _17679_ & D[34] /*69010*/;
assign _17681_ = _16995_ & _17678_ /*69005*/;
assign _17682_ = _16995_ ^ _17678_ /*69008*/;
assign _17683_ = _17674_ & _17682_ /*69006*/;
assign _17443_ = _17674_ ^ _17682_ /*69007*/;
assign _17680_ = _17681_ | _17683_ /*69004*/;
assign _17685_ = ~Q[44] /*69003*/;
assign _17684_ = _17685_ & D[35] /*69002*/;
assign _17687_ = _16996_ & _17684_ /*68997*/;
assign _17688_ = _16996_ ^ _17684_ /*69000*/;
assign _17689_ = _17680_ & _17688_ /*68998*/;
assign _17444_ = _17680_ ^ _17688_ /*68999*/;
assign _17686_ = _17687_ | _17689_ /*68996*/;
assign _17691_ = ~Q[44] /*68995*/;
assign _17690_ = _17691_ & D[36] /*68994*/;
assign _17693_ = _16997_ & _17690_ /*68989*/;
assign _17694_ = _16997_ ^ _17690_ /*68992*/;
assign _17695_ = _17686_ & _17694_ /*68990*/;
assign _17445_ = _17686_ ^ _17694_ /*68991*/;
assign _17692_ = _17693_ | _17695_ /*68988*/;
assign _17697_ = ~Q[44] /*68987*/;
assign _17696_ = _17697_ & D[37] /*68986*/;
assign _17699_ = _16998_ & _17696_ /*68981*/;
assign _17700_ = _16998_ ^ _17696_ /*68984*/;
assign _17701_ = _17692_ & _17700_ /*68982*/;
assign _17446_ = _17692_ ^ _17700_ /*68983*/;
assign _17698_ = _17699_ | _17701_ /*68980*/;
assign _17703_ = ~Q[44] /*68979*/;
assign _17702_ = _17703_ & D[38] /*68978*/;
assign _17705_ = _16999_ & _17702_ /*68973*/;
assign _17706_ = _16999_ ^ _17702_ /*68976*/;
assign _17707_ = _17698_ & _17706_ /*68974*/;
assign _17447_ = _17698_ ^ _17706_ /*68975*/;
assign _17704_ = _17705_ | _17707_ /*68972*/;
assign _17709_ = ~Q[44] /*68971*/;
assign _17708_ = _17709_ & D[39] /*68970*/;
assign _17711_ = _17000_ & _17708_ /*68965*/;
assign _17712_ = _17000_ ^ _17708_ /*68968*/;
assign _17713_ = _17704_ & _17712_ /*68966*/;
assign _17448_ = _17704_ ^ _17712_ /*68967*/;
assign _17710_ = _17711_ | _17713_ /*68964*/;
assign _17715_ = ~Q[44] /*68963*/;
assign _17714_ = _17715_ & D[40] /*68962*/;
assign _17717_ = _17001_ & _17714_ /*68957*/;
assign _17718_ = _17001_ ^ _17714_ /*68960*/;
assign _17719_ = _17710_ & _17718_ /*68958*/;
assign _17449_ = _17710_ ^ _17718_ /*68959*/;
assign _17716_ = _17717_ | _17719_ /*68956*/;
assign _17721_ = ~Q[44] /*68955*/;
assign _17720_ = _17721_ & D[41] /*68954*/;
assign _17723_ = _17002_ & _17720_ /*68949*/;
assign _17724_ = _17002_ ^ _17720_ /*68952*/;
assign _17725_ = _17716_ & _17724_ /*68950*/;
assign _17450_ = _17716_ ^ _17724_ /*68951*/;
assign _17722_ = _17723_ | _17725_ /*68948*/;
assign _17727_ = ~Q[44] /*68947*/;
assign _17726_ = _17727_ & D[42] /*68946*/;
assign _17729_ = _17003_ & _17726_ /*68941*/;
assign _17730_ = _17003_ ^ _17726_ /*68944*/;
assign _17731_ = _17722_ & _17730_ /*68942*/;
assign _17451_ = _17722_ ^ _17730_ /*68943*/;
assign _17728_ = _17729_ | _17731_ /*68940*/;
assign _17733_ = ~Q[44] /*68939*/;
assign _17732_ = _17733_ & D[43] /*68938*/;
assign _17735_ = _17004_ & _17732_ /*68933*/;
assign _17736_ = _17004_ ^ _17732_ /*68936*/;
assign _17737_ = _17728_ & _17736_ /*68934*/;
assign _17452_ = _17728_ ^ _17736_ /*68935*/;
assign _17734_ = _17735_ | _17737_ /*68932*/;
assign _17739_ = ~Q[44] /*68931*/;
assign _17738_ = _17739_ & D[44] /*68930*/;
assign _17741_ = _17005_ & _17738_ /*68925*/;
assign _17742_ = _17005_ ^ _17738_ /*68928*/;
assign _17743_ = _17734_ & _17742_ /*68926*/;
assign _17453_ = _17734_ ^ _17742_ /*68927*/;
assign _17740_ = _17741_ | _17743_ /*68924*/;
assign _17745_ = ~Q[44] /*68923*/;
assign _17744_ = _17745_ & D[45] /*68922*/;
assign _17747_ = _17006_ & _17744_ /*68917*/;
assign _17748_ = _17006_ ^ _17744_ /*68920*/;
assign _17749_ = _17740_ & _17748_ /*68918*/;
assign _17454_ = _17740_ ^ _17748_ /*68919*/;
assign _17746_ = _17747_ | _17749_ /*68916*/;
assign _17751_ = ~Q[44] /*68915*/;
assign _17750_ = _17751_ & D[46] /*68914*/;
assign _17753_ = _17007_ & _17750_ /*68909*/;
assign _17754_ = _17007_ ^ _17750_ /*68912*/;
assign _17755_ = _17746_ & _17754_ /*68910*/;
assign _17455_ = _17746_ ^ _17754_ /*68911*/;
assign _17752_ = _17753_ | _17755_ /*68908*/;
assign _17757_ = ~Q[44] /*68907*/;
assign _17756_ = _17757_ & D[47] /*68906*/;
assign _17759_ = _17008_ & _17756_ /*68901*/;
assign _17760_ = _17008_ ^ _17756_ /*68904*/;
assign _17761_ = _17752_ & _17760_ /*68902*/;
assign _17456_ = _17752_ ^ _17760_ /*68903*/;
assign _17758_ = _17759_ | _17761_ /*68900*/;
assign _17763_ = ~Q[44] /*68899*/;
assign _17762_ = _17763_ & D[48] /*68898*/;
assign _17765_ = _17009_ & _17762_ /*68893*/;
assign _17766_ = _17009_ ^ _17762_ /*68896*/;
assign _17767_ = _17758_ & _17766_ /*68894*/;
assign _17457_ = _17758_ ^ _17766_ /*68895*/;
assign _17764_ = _17765_ | _17767_ /*68892*/;
assign _17769_ = ~Q[44] /*68891*/;
assign _17768_ = _17769_ & D[49] /*68890*/;
assign _17771_ = _17010_ & _17768_ /*68885*/;
assign _17772_ = _17010_ ^ _17768_ /*68888*/;
assign _17773_ = _17764_ & _17772_ /*68886*/;
assign _17458_ = _17764_ ^ _17772_ /*68887*/;
assign _17770_ = _17771_ | _17773_ /*68884*/;
assign _17775_ = ~Q[44] /*68883*/;
assign _17774_ = _17775_ & D[50] /*68882*/;
assign _17777_ = _17011_ & _17774_ /*68877*/;
assign _17778_ = _17011_ ^ _17774_ /*68880*/;
assign _17779_ = _17770_ & _17778_ /*68878*/;
assign _17459_ = _17770_ ^ _17778_ /*68879*/;
assign _17776_ = _17777_ | _17779_ /*68876*/;
assign _17781_ = ~Q[44] /*68875*/;
assign _17780_ = _17781_ & D[51] /*68874*/;
assign _17783_ = _17012_ & _17780_ /*68869*/;
assign _17784_ = _17012_ ^ _17780_ /*68872*/;
assign _17785_ = _17776_ & _17784_ /*68870*/;
assign _17460_ = _17776_ ^ _17784_ /*68871*/;
assign _17782_ = _17783_ | _17785_ /*68868*/;
assign _17787_ = ~Q[44] /*68867*/;
assign _17786_ = _17787_ & D[52] /*68866*/;
assign _17789_ = _17013_ & _17786_ /*68861*/;
assign _17790_ = _17013_ ^ _17786_ /*68864*/;
assign _17791_ = _17782_ & _17790_ /*68862*/;
assign _17461_ = _17782_ ^ _17790_ /*68863*/;
assign _17788_ = _17789_ | _17791_ /*68860*/;
assign _17793_ = ~Q[44] /*68859*/;
assign _17792_ = _17793_ & D[53] /*68858*/;
assign _17795_ = _17014_ & _17792_ /*68853*/;
assign _17796_ = _17014_ ^ _17792_ /*68856*/;
assign _17797_ = _17788_ & _17796_ /*68854*/;
assign _17462_ = _17788_ ^ _17796_ /*68855*/;
assign _17794_ = _17795_ | _17797_ /*68852*/;
assign _17799_ = ~Q[44] /*68851*/;
assign _17798_ = _17799_ & D[54] /*68850*/;
assign _17801_ = _17015_ & _17798_ /*68845*/;
assign _17802_ = _17015_ ^ _17798_ /*68848*/;
assign _17803_ = _17794_ & _17802_ /*68846*/;
assign _17463_ = _17794_ ^ _17802_ /*68847*/;
assign _17800_ = _17801_ | _17803_ /*68844*/;
assign _17805_ = ~Q[44] /*68843*/;
assign _17804_ = _17805_ & D[55] /*68842*/;
assign _17807_ = _17016_ & _17804_ /*68837*/;
assign _17808_ = _17016_ ^ _17804_ /*68840*/;
assign _17809_ = _17800_ & _17808_ /*68838*/;
assign _17464_ = _17800_ ^ _17808_ /*68839*/;
assign _17806_ = _17807_ | _17809_ /*68836*/;
assign _17811_ = ~Q[44] /*68835*/;
assign _17810_ = _17811_ & D[56] /*68834*/;
assign _17813_ = _17017_ & _17810_ /*68829*/;
assign _17814_ = _17017_ ^ _17810_ /*68832*/;
assign _17815_ = _17806_ & _17814_ /*68830*/;
assign _17465_ = _17806_ ^ _17814_ /*68831*/;
assign _17812_ = _17813_ | _17815_ /*68828*/;
assign _17817_ = ~Q[44] /*68827*/;
assign _17816_ = _17817_ & D[57] /*68826*/;
assign _17819_ = _17018_ & _17816_ /*68821*/;
assign _17820_ = _17018_ ^ _17816_ /*68824*/;
assign _17821_ = _17812_ & _17820_ /*68822*/;
assign _17466_ = _17812_ ^ _17820_ /*68823*/;
assign _17818_ = _17819_ | _17821_ /*68820*/;
assign _17823_ = ~Q[44] /*68819*/;
assign _17822_ = _17823_ & D[58] /*68818*/;
assign _17825_ = _17019_ & _17822_ /*68813*/;
assign _17826_ = _17019_ ^ _17822_ /*68816*/;
assign _17827_ = _17818_ & _17826_ /*68814*/;
assign _17467_ = _17818_ ^ _17826_ /*68815*/;
assign _17824_ = _17825_ | _17827_ /*68812*/;
assign _17829_ = ~Q[44] /*68811*/;
assign _17828_ = _17829_ & D[59] /*68810*/;
assign _17831_ = _17020_ & _17828_ /*68805*/;
assign _17832_ = _17020_ ^ _17828_ /*68808*/;
assign _17833_ = _17824_ & _17832_ /*68806*/;
assign _17468_ = _17824_ ^ _17832_ /*68807*/;
assign _17830_ = _17831_ | _17833_ /*68804*/;
assign _17835_ = ~Q[44] /*68803*/;
assign _17834_ = _17835_ & D[60] /*68802*/;
assign _17837_ = _17021_ & _17834_ /*68797*/;
assign _17838_ = _17021_ ^ _17834_ /*68800*/;
assign _17839_ = _17830_ & _17838_ /*68798*/;
assign _17469_ = _17830_ ^ _17838_ /*68799*/;
assign _17836_ = _17837_ | _17839_ /*68796*/;
assign _17841_ = ~Q[44] /*68795*/;
assign _17840_ = _17841_ & D[61] /*68794*/;
assign _17843_ = _17022_ & _17840_ /*68789*/;
assign _17844_ = _17022_ ^ _17840_ /*68792*/;
assign _17845_ = _17836_ & _17844_ /*68790*/;
assign _17470_ = _17836_ ^ _17844_ /*68791*/;
assign _17842_ = _17843_ | _17845_ /*68788*/;
assign _17847_ = ~Q[44] /*68787*/;
assign _17846_ = _17847_ & D[62] /*68786*/;
assign _17849_ = _17023_ & _17846_ /*68781*/;
assign _17850_ = _17023_ ^ _17846_ /*68784*/;
assign _17851_ = _17842_ & _17850_ /*68782*/;
assign _17471_ = _17842_ ^ _17850_ /*68783*/;
assign _17848_ = _17849_ | _17851_ /*68780*/;
assign _17853_ = ~Q[44] /*68779*/;
assign _17852_ = _17853_ & zeroWire /*68778*/;
assign _17854_ = _17024_ ^ _17852_ /*68776*/;
assign _17472_ = _17854_ ^ _17848_ /*68775*/;
assign _17925_ = ~D[0] /*68521*/;
assign _17922_ = R_0[43] & _17925_ /*68517*/;
assign _17923_ = R_0[43] ^ _17925_ /*68520*/;
assign _17924_ = oneWire & _17923_ /*68518*/;
assign _17857_ = oneWire ^ _17923_ /*68519*/;
assign _17921_ = _17922_ | _17924_ /*68516*/;
assign _17930_ = ~D[1] /*68515*/;
assign _17927_ = _17409_ & _17930_ /*68511*/;
assign _17928_ = _17409_ ^ _17930_ /*68514*/;
assign _17929_ = _17921_ & _17928_ /*68512*/;
assign _17858_ = _17921_ ^ _17928_ /*68513*/;
assign _17926_ = _17927_ | _17929_ /*68510*/;
assign _17935_ = ~D[2] /*68509*/;
assign _17932_ = _17410_ & _17935_ /*68505*/;
assign _17933_ = _17410_ ^ _17935_ /*68508*/;
assign _17934_ = _17926_ & _17933_ /*68506*/;
assign _17859_ = _17926_ ^ _17933_ /*68507*/;
assign _17931_ = _17932_ | _17934_ /*68504*/;
assign _17940_ = ~D[3] /*68503*/;
assign _17937_ = _17411_ & _17940_ /*68499*/;
assign _17938_ = _17411_ ^ _17940_ /*68502*/;
assign _17939_ = _17931_ & _17938_ /*68500*/;
assign _17860_ = _17931_ ^ _17938_ /*68501*/;
assign _17936_ = _17937_ | _17939_ /*68498*/;
assign _17945_ = ~D[4] /*68497*/;
assign _17942_ = _17412_ & _17945_ /*68493*/;
assign _17943_ = _17412_ ^ _17945_ /*68496*/;
assign _17944_ = _17936_ & _17943_ /*68494*/;
assign _17861_ = _17936_ ^ _17943_ /*68495*/;
assign _17941_ = _17942_ | _17944_ /*68492*/;
assign _17950_ = ~D[5] /*68491*/;
assign _17947_ = _17413_ & _17950_ /*68487*/;
assign _17948_ = _17413_ ^ _17950_ /*68490*/;
assign _17949_ = _17941_ & _17948_ /*68488*/;
assign _17862_ = _17941_ ^ _17948_ /*68489*/;
assign _17946_ = _17947_ | _17949_ /*68486*/;
assign _17955_ = ~D[6] /*68485*/;
assign _17952_ = _17414_ & _17955_ /*68481*/;
assign _17953_ = _17414_ ^ _17955_ /*68484*/;
assign _17954_ = _17946_ & _17953_ /*68482*/;
assign _17863_ = _17946_ ^ _17953_ /*68483*/;
assign _17951_ = _17952_ | _17954_ /*68480*/;
assign _17960_ = ~D[7] /*68479*/;
assign _17957_ = _17415_ & _17960_ /*68475*/;
assign _17958_ = _17415_ ^ _17960_ /*68478*/;
assign _17959_ = _17951_ & _17958_ /*68476*/;
assign _17864_ = _17951_ ^ _17958_ /*68477*/;
assign _17956_ = _17957_ | _17959_ /*68474*/;
assign _17965_ = ~D[8] /*68473*/;
assign _17962_ = _17416_ & _17965_ /*68469*/;
assign _17963_ = _17416_ ^ _17965_ /*68472*/;
assign _17964_ = _17956_ & _17963_ /*68470*/;
assign _17865_ = _17956_ ^ _17963_ /*68471*/;
assign _17961_ = _17962_ | _17964_ /*68468*/;
assign _17970_ = ~D[9] /*68467*/;
assign _17967_ = _17417_ & _17970_ /*68463*/;
assign _17968_ = _17417_ ^ _17970_ /*68466*/;
assign _17969_ = _17961_ & _17968_ /*68464*/;
assign _17866_ = _17961_ ^ _17968_ /*68465*/;
assign _17966_ = _17967_ | _17969_ /*68462*/;
assign _17975_ = ~D[10] /*68461*/;
assign _17972_ = _17418_ & _17975_ /*68457*/;
assign _17973_ = _17418_ ^ _17975_ /*68460*/;
assign _17974_ = _17966_ & _17973_ /*68458*/;
assign _17867_ = _17966_ ^ _17973_ /*68459*/;
assign _17971_ = _17972_ | _17974_ /*68456*/;
assign _17980_ = ~D[11] /*68455*/;
assign _17977_ = _17419_ & _17980_ /*68451*/;
assign _17978_ = _17419_ ^ _17980_ /*68454*/;
assign _17979_ = _17971_ & _17978_ /*68452*/;
assign _17868_ = _17971_ ^ _17978_ /*68453*/;
assign _17976_ = _17977_ | _17979_ /*68450*/;
assign _17985_ = ~D[12] /*68449*/;
assign _17982_ = _17420_ & _17985_ /*68445*/;
assign _17983_ = _17420_ ^ _17985_ /*68448*/;
assign _17984_ = _17976_ & _17983_ /*68446*/;
assign _17869_ = _17976_ ^ _17983_ /*68447*/;
assign _17981_ = _17982_ | _17984_ /*68444*/;
assign _17990_ = ~D[13] /*68443*/;
assign _17987_ = _17421_ & _17990_ /*68439*/;
assign _17988_ = _17421_ ^ _17990_ /*68442*/;
assign _17989_ = _17981_ & _17988_ /*68440*/;
assign _17870_ = _17981_ ^ _17988_ /*68441*/;
assign _17986_ = _17987_ | _17989_ /*68438*/;
assign _17995_ = ~D[14] /*68437*/;
assign _17992_ = _17422_ & _17995_ /*68433*/;
assign _17993_ = _17422_ ^ _17995_ /*68436*/;
assign _17994_ = _17986_ & _17993_ /*68434*/;
assign _17871_ = _17986_ ^ _17993_ /*68435*/;
assign _17991_ = _17992_ | _17994_ /*68432*/;
assign _18000_ = ~D[15] /*68431*/;
assign _17997_ = _17423_ & _18000_ /*68427*/;
assign _17998_ = _17423_ ^ _18000_ /*68430*/;
assign _17999_ = _17991_ & _17998_ /*68428*/;
assign _17872_ = _17991_ ^ _17998_ /*68429*/;
assign _17996_ = _17997_ | _17999_ /*68426*/;
assign _18005_ = ~D[16] /*68425*/;
assign _18002_ = _17424_ & _18005_ /*68421*/;
assign _18003_ = _17424_ ^ _18005_ /*68424*/;
assign _18004_ = _17996_ & _18003_ /*68422*/;
assign _17873_ = _17996_ ^ _18003_ /*68423*/;
assign _18001_ = _18002_ | _18004_ /*68420*/;
assign _18010_ = ~D[17] /*68419*/;
assign _18007_ = _17425_ & _18010_ /*68415*/;
assign _18008_ = _17425_ ^ _18010_ /*68418*/;
assign _18009_ = _18001_ & _18008_ /*68416*/;
assign _17874_ = _18001_ ^ _18008_ /*68417*/;
assign _18006_ = _18007_ | _18009_ /*68414*/;
assign _18015_ = ~D[18] /*68413*/;
assign _18012_ = _17426_ & _18015_ /*68409*/;
assign _18013_ = _17426_ ^ _18015_ /*68412*/;
assign _18014_ = _18006_ & _18013_ /*68410*/;
assign _17875_ = _18006_ ^ _18013_ /*68411*/;
assign _18011_ = _18012_ | _18014_ /*68408*/;
assign _18020_ = ~D[19] /*68407*/;
assign _18017_ = _17427_ & _18020_ /*68403*/;
assign _18018_ = _17427_ ^ _18020_ /*68406*/;
assign _18019_ = _18011_ & _18018_ /*68404*/;
assign _17876_ = _18011_ ^ _18018_ /*68405*/;
assign _18016_ = _18017_ | _18019_ /*68402*/;
assign _18025_ = ~D[20] /*68401*/;
assign _18022_ = _17428_ & _18025_ /*68397*/;
assign _18023_ = _17428_ ^ _18025_ /*68400*/;
assign _18024_ = _18016_ & _18023_ /*68398*/;
assign _17877_ = _18016_ ^ _18023_ /*68399*/;
assign _18021_ = _18022_ | _18024_ /*68396*/;
assign _18030_ = ~D[21] /*68395*/;
assign _18027_ = _17429_ & _18030_ /*68391*/;
assign _18028_ = _17429_ ^ _18030_ /*68394*/;
assign _18029_ = _18021_ & _18028_ /*68392*/;
assign _17878_ = _18021_ ^ _18028_ /*68393*/;
assign _18026_ = _18027_ | _18029_ /*68390*/;
assign _18035_ = ~D[22] /*68389*/;
assign _18032_ = _17430_ & _18035_ /*68385*/;
assign _18033_ = _17430_ ^ _18035_ /*68388*/;
assign _18034_ = _18026_ & _18033_ /*68386*/;
assign _17879_ = _18026_ ^ _18033_ /*68387*/;
assign _18031_ = _18032_ | _18034_ /*68384*/;
assign _18040_ = ~D[23] /*68383*/;
assign _18037_ = _17431_ & _18040_ /*68379*/;
assign _18038_ = _17431_ ^ _18040_ /*68382*/;
assign _18039_ = _18031_ & _18038_ /*68380*/;
assign _17880_ = _18031_ ^ _18038_ /*68381*/;
assign _18036_ = _18037_ | _18039_ /*68378*/;
assign _18045_ = ~D[24] /*68377*/;
assign _18042_ = _17432_ & _18045_ /*68373*/;
assign _18043_ = _17432_ ^ _18045_ /*68376*/;
assign _18044_ = _18036_ & _18043_ /*68374*/;
assign _17881_ = _18036_ ^ _18043_ /*68375*/;
assign _18041_ = _18042_ | _18044_ /*68372*/;
assign _18050_ = ~D[25] /*68371*/;
assign _18047_ = _17433_ & _18050_ /*68367*/;
assign _18048_ = _17433_ ^ _18050_ /*68370*/;
assign _18049_ = _18041_ & _18048_ /*68368*/;
assign _17882_ = _18041_ ^ _18048_ /*68369*/;
assign _18046_ = _18047_ | _18049_ /*68366*/;
assign _18055_ = ~D[26] /*68365*/;
assign _18052_ = _17434_ & _18055_ /*68361*/;
assign _18053_ = _17434_ ^ _18055_ /*68364*/;
assign _18054_ = _18046_ & _18053_ /*68362*/;
assign _17883_ = _18046_ ^ _18053_ /*68363*/;
assign _18051_ = _18052_ | _18054_ /*68360*/;
assign _18060_ = ~D[27] /*68359*/;
assign _18057_ = _17435_ & _18060_ /*68355*/;
assign _18058_ = _17435_ ^ _18060_ /*68358*/;
assign _18059_ = _18051_ & _18058_ /*68356*/;
assign _17884_ = _18051_ ^ _18058_ /*68357*/;
assign _18056_ = _18057_ | _18059_ /*68354*/;
assign _18065_ = ~D[28] /*68353*/;
assign _18062_ = _17436_ & _18065_ /*68349*/;
assign _18063_ = _17436_ ^ _18065_ /*68352*/;
assign _18064_ = _18056_ & _18063_ /*68350*/;
assign _17885_ = _18056_ ^ _18063_ /*68351*/;
assign _18061_ = _18062_ | _18064_ /*68348*/;
assign _18070_ = ~D[29] /*68347*/;
assign _18067_ = _17437_ & _18070_ /*68343*/;
assign _18068_ = _17437_ ^ _18070_ /*68346*/;
assign _18069_ = _18061_ & _18068_ /*68344*/;
assign _17886_ = _18061_ ^ _18068_ /*68345*/;
assign _18066_ = _18067_ | _18069_ /*68342*/;
assign _18075_ = ~D[30] /*68341*/;
assign _18072_ = _17438_ & _18075_ /*68337*/;
assign _18073_ = _17438_ ^ _18075_ /*68340*/;
assign _18074_ = _18066_ & _18073_ /*68338*/;
assign _17887_ = _18066_ ^ _18073_ /*68339*/;
assign _18071_ = _18072_ | _18074_ /*68336*/;
assign _18080_ = ~D[31] /*68335*/;
assign _18077_ = _17439_ & _18080_ /*68331*/;
assign _18078_ = _17439_ ^ _18080_ /*68334*/;
assign _18079_ = _18071_ & _18078_ /*68332*/;
assign _17888_ = _18071_ ^ _18078_ /*68333*/;
assign _18076_ = _18077_ | _18079_ /*68330*/;
assign _18085_ = ~D[32] /*68329*/;
assign _18082_ = _17440_ & _18085_ /*68325*/;
assign _18083_ = _17440_ ^ _18085_ /*68328*/;
assign _18084_ = _18076_ & _18083_ /*68326*/;
assign _17889_ = _18076_ ^ _18083_ /*68327*/;
assign _18081_ = _18082_ | _18084_ /*68324*/;
assign _18090_ = ~D[33] /*68323*/;
assign _18087_ = _17441_ & _18090_ /*68319*/;
assign _18088_ = _17441_ ^ _18090_ /*68322*/;
assign _18089_ = _18081_ & _18088_ /*68320*/;
assign _17890_ = _18081_ ^ _18088_ /*68321*/;
assign _18086_ = _18087_ | _18089_ /*68318*/;
assign _18095_ = ~D[34] /*68317*/;
assign _18092_ = _17442_ & _18095_ /*68313*/;
assign _18093_ = _17442_ ^ _18095_ /*68316*/;
assign _18094_ = _18086_ & _18093_ /*68314*/;
assign _17891_ = _18086_ ^ _18093_ /*68315*/;
assign _18091_ = _18092_ | _18094_ /*68312*/;
assign _18100_ = ~D[35] /*68311*/;
assign _18097_ = _17443_ & _18100_ /*68307*/;
assign _18098_ = _17443_ ^ _18100_ /*68310*/;
assign _18099_ = _18091_ & _18098_ /*68308*/;
assign _17892_ = _18091_ ^ _18098_ /*68309*/;
assign _18096_ = _18097_ | _18099_ /*68306*/;
assign _18105_ = ~D[36] /*68305*/;
assign _18102_ = _17444_ & _18105_ /*68301*/;
assign _18103_ = _17444_ ^ _18105_ /*68304*/;
assign _18104_ = _18096_ & _18103_ /*68302*/;
assign _17893_ = _18096_ ^ _18103_ /*68303*/;
assign _18101_ = _18102_ | _18104_ /*68300*/;
assign _18110_ = ~D[37] /*68299*/;
assign _18107_ = _17445_ & _18110_ /*68295*/;
assign _18108_ = _17445_ ^ _18110_ /*68298*/;
assign _18109_ = _18101_ & _18108_ /*68296*/;
assign _17894_ = _18101_ ^ _18108_ /*68297*/;
assign _18106_ = _18107_ | _18109_ /*68294*/;
assign _18115_ = ~D[38] /*68293*/;
assign _18112_ = _17446_ & _18115_ /*68289*/;
assign _18113_ = _17446_ ^ _18115_ /*68292*/;
assign _18114_ = _18106_ & _18113_ /*68290*/;
assign _17895_ = _18106_ ^ _18113_ /*68291*/;
assign _18111_ = _18112_ | _18114_ /*68288*/;
assign _18120_ = ~D[39] /*68287*/;
assign _18117_ = _17447_ & _18120_ /*68283*/;
assign _18118_ = _17447_ ^ _18120_ /*68286*/;
assign _18119_ = _18111_ & _18118_ /*68284*/;
assign _17896_ = _18111_ ^ _18118_ /*68285*/;
assign _18116_ = _18117_ | _18119_ /*68282*/;
assign _18125_ = ~D[40] /*68281*/;
assign _18122_ = _17448_ & _18125_ /*68277*/;
assign _18123_ = _17448_ ^ _18125_ /*68280*/;
assign _18124_ = _18116_ & _18123_ /*68278*/;
assign _17897_ = _18116_ ^ _18123_ /*68279*/;
assign _18121_ = _18122_ | _18124_ /*68276*/;
assign _18130_ = ~D[41] /*68275*/;
assign _18127_ = _17449_ & _18130_ /*68271*/;
assign _18128_ = _17449_ ^ _18130_ /*68274*/;
assign _18129_ = _18121_ & _18128_ /*68272*/;
assign _17898_ = _18121_ ^ _18128_ /*68273*/;
assign _18126_ = _18127_ | _18129_ /*68270*/;
assign _18135_ = ~D[42] /*68269*/;
assign _18132_ = _17450_ & _18135_ /*68265*/;
assign _18133_ = _17450_ ^ _18135_ /*68268*/;
assign _18134_ = _18126_ & _18133_ /*68266*/;
assign _17899_ = _18126_ ^ _18133_ /*68267*/;
assign _18131_ = _18132_ | _18134_ /*68264*/;
assign _18140_ = ~D[43] /*68263*/;
assign _18137_ = _17451_ & _18140_ /*68259*/;
assign _18138_ = _17451_ ^ _18140_ /*68262*/;
assign _18139_ = _18131_ & _18138_ /*68260*/;
assign _17900_ = _18131_ ^ _18138_ /*68261*/;
assign _18136_ = _18137_ | _18139_ /*68258*/;
assign _18145_ = ~D[44] /*68257*/;
assign _18142_ = _17452_ & _18145_ /*68253*/;
assign _18143_ = _17452_ ^ _18145_ /*68256*/;
assign _18144_ = _18136_ & _18143_ /*68254*/;
assign _17901_ = _18136_ ^ _18143_ /*68255*/;
assign _18141_ = _18142_ | _18144_ /*68252*/;
assign _18150_ = ~D[45] /*68251*/;
assign _18147_ = _17453_ & _18150_ /*68247*/;
assign _18148_ = _17453_ ^ _18150_ /*68250*/;
assign _18149_ = _18141_ & _18148_ /*68248*/;
assign _17902_ = _18141_ ^ _18148_ /*68249*/;
assign _18146_ = _18147_ | _18149_ /*68246*/;
assign _18155_ = ~D[46] /*68245*/;
assign _18152_ = _17454_ & _18155_ /*68241*/;
assign _18153_ = _17454_ ^ _18155_ /*68244*/;
assign _18154_ = _18146_ & _18153_ /*68242*/;
assign _17903_ = _18146_ ^ _18153_ /*68243*/;
assign _18151_ = _18152_ | _18154_ /*68240*/;
assign _18160_ = ~D[47] /*68239*/;
assign _18157_ = _17455_ & _18160_ /*68235*/;
assign _18158_ = _17455_ ^ _18160_ /*68238*/;
assign _18159_ = _18151_ & _18158_ /*68236*/;
assign _17904_ = _18151_ ^ _18158_ /*68237*/;
assign _18156_ = _18157_ | _18159_ /*68234*/;
assign _18165_ = ~D[48] /*68233*/;
assign _18162_ = _17456_ & _18165_ /*68229*/;
assign _18163_ = _17456_ ^ _18165_ /*68232*/;
assign _18164_ = _18156_ & _18163_ /*68230*/;
assign _17905_ = _18156_ ^ _18163_ /*68231*/;
assign _18161_ = _18162_ | _18164_ /*68228*/;
assign _18170_ = ~D[49] /*68227*/;
assign _18167_ = _17457_ & _18170_ /*68223*/;
assign _18168_ = _17457_ ^ _18170_ /*68226*/;
assign _18169_ = _18161_ & _18168_ /*68224*/;
assign _17906_ = _18161_ ^ _18168_ /*68225*/;
assign _18166_ = _18167_ | _18169_ /*68222*/;
assign _18175_ = ~D[50] /*68221*/;
assign _18172_ = _17458_ & _18175_ /*68217*/;
assign _18173_ = _17458_ ^ _18175_ /*68220*/;
assign _18174_ = _18166_ & _18173_ /*68218*/;
assign _17907_ = _18166_ ^ _18173_ /*68219*/;
assign _18171_ = _18172_ | _18174_ /*68216*/;
assign _18180_ = ~D[51] /*68215*/;
assign _18177_ = _17459_ & _18180_ /*68211*/;
assign _18178_ = _17459_ ^ _18180_ /*68214*/;
assign _18179_ = _18171_ & _18178_ /*68212*/;
assign _17908_ = _18171_ ^ _18178_ /*68213*/;
assign _18176_ = _18177_ | _18179_ /*68210*/;
assign _18185_ = ~D[52] /*68209*/;
assign _18182_ = _17460_ & _18185_ /*68205*/;
assign _18183_ = _17460_ ^ _18185_ /*68208*/;
assign _18184_ = _18176_ & _18183_ /*68206*/;
assign _17909_ = _18176_ ^ _18183_ /*68207*/;
assign _18181_ = _18182_ | _18184_ /*68204*/;
assign _18190_ = ~D[53] /*68203*/;
assign _18187_ = _17461_ & _18190_ /*68199*/;
assign _18188_ = _17461_ ^ _18190_ /*68202*/;
assign _18189_ = _18181_ & _18188_ /*68200*/;
assign _17910_ = _18181_ ^ _18188_ /*68201*/;
assign _18186_ = _18187_ | _18189_ /*68198*/;
assign _18195_ = ~D[54] /*68197*/;
assign _18192_ = _17462_ & _18195_ /*68193*/;
assign _18193_ = _17462_ ^ _18195_ /*68196*/;
assign _18194_ = _18186_ & _18193_ /*68194*/;
assign _17911_ = _18186_ ^ _18193_ /*68195*/;
assign _18191_ = _18192_ | _18194_ /*68192*/;
assign _18200_ = ~D[55] /*68191*/;
assign _18197_ = _17463_ & _18200_ /*68187*/;
assign _18198_ = _17463_ ^ _18200_ /*68190*/;
assign _18199_ = _18191_ & _18198_ /*68188*/;
assign _17912_ = _18191_ ^ _18198_ /*68189*/;
assign _18196_ = _18197_ | _18199_ /*68186*/;
assign _18205_ = ~D[56] /*68185*/;
assign _18202_ = _17464_ & _18205_ /*68181*/;
assign _18203_ = _17464_ ^ _18205_ /*68184*/;
assign _18204_ = _18196_ & _18203_ /*68182*/;
assign _17913_ = _18196_ ^ _18203_ /*68183*/;
assign _18201_ = _18202_ | _18204_ /*68180*/;
assign _18210_ = ~D[57] /*68179*/;
assign _18207_ = _17465_ & _18210_ /*68175*/;
assign _18208_ = _17465_ ^ _18210_ /*68178*/;
assign _18209_ = _18201_ & _18208_ /*68176*/;
assign _17914_ = _18201_ ^ _18208_ /*68177*/;
assign _18206_ = _18207_ | _18209_ /*68174*/;
assign _18215_ = ~D[58] /*68173*/;
assign _18212_ = _17466_ & _18215_ /*68169*/;
assign _18213_ = _17466_ ^ _18215_ /*68172*/;
assign _18214_ = _18206_ & _18213_ /*68170*/;
assign _17915_ = _18206_ ^ _18213_ /*68171*/;
assign _18211_ = _18212_ | _18214_ /*68168*/;
assign _18220_ = ~D[59] /*68167*/;
assign _18217_ = _17467_ & _18220_ /*68163*/;
assign _18218_ = _17467_ ^ _18220_ /*68166*/;
assign _18219_ = _18211_ & _18218_ /*68164*/;
assign _17916_ = _18211_ ^ _18218_ /*68165*/;
assign _18216_ = _18217_ | _18219_ /*68162*/;
assign _18225_ = ~D[60] /*68161*/;
assign _18222_ = _17468_ & _18225_ /*68157*/;
assign _18223_ = _17468_ ^ _18225_ /*68160*/;
assign _18224_ = _18216_ & _18223_ /*68158*/;
assign _17917_ = _18216_ ^ _18223_ /*68159*/;
assign _18221_ = _18222_ | _18224_ /*68156*/;
assign _18230_ = ~D[61] /*68155*/;
assign _18227_ = _17469_ & _18230_ /*68151*/;
assign _18228_ = _17469_ ^ _18230_ /*68154*/;
assign _18229_ = _18221_ & _18228_ /*68152*/;
assign _17918_ = _18221_ ^ _18228_ /*68153*/;
assign _18226_ = _18227_ | _18229_ /*68150*/;
assign _18235_ = ~D[62] /*68149*/;
assign _18232_ = _17470_ & _18235_ /*68145*/;
assign _18233_ = _17470_ ^ _18235_ /*68148*/;
assign _18234_ = _18226_ & _18233_ /*68146*/;
assign _17919_ = _18226_ ^ _18233_ /*68147*/;
assign _18231_ = _18232_ | _18234_ /*68144*/;
assign _18236_ = _17471_ & oneWire /*68139*/;
assign _18237_ = _17471_ ^ oneWire /*68142*/;
assign _18238_ = _18231_ & _18237_ /*68140*/;
assign _17920_ = _18231_ ^ _18237_ /*68141*/;
assign Q[43] = _18236_ | _18238_ /*68138*/;
assign _18371_ = ~Q[43] /*67753*/;
assign _18370_ = _18371_ & D[0] /*67752*/;
assign _18373_ = _17857_ & _18370_ /*67747*/;
assign _18374_ = _17857_ ^ _18370_ /*67750*/;
assign _18375_ = zeroWire & _18374_ /*67748*/;
assign _18305_ = zeroWire ^ _18374_ /*67749*/;
assign _18372_ = _18373_ | _18375_ /*67746*/;
assign _18377_ = ~Q[43] /*67745*/;
assign _18376_ = _18377_ & D[1] /*67744*/;
assign _18379_ = _17858_ & _18376_ /*67739*/;
assign _18380_ = _17858_ ^ _18376_ /*67742*/;
assign _18381_ = _18372_ & _18380_ /*67740*/;
assign _18306_ = _18372_ ^ _18380_ /*67741*/;
assign _18378_ = _18379_ | _18381_ /*67738*/;
assign _18383_ = ~Q[43] /*67737*/;
assign _18382_ = _18383_ & D[2] /*67736*/;
assign _18385_ = _17859_ & _18382_ /*67731*/;
assign _18386_ = _17859_ ^ _18382_ /*67734*/;
assign _18387_ = _18378_ & _18386_ /*67732*/;
assign _18307_ = _18378_ ^ _18386_ /*67733*/;
assign _18384_ = _18385_ | _18387_ /*67730*/;
assign _18389_ = ~Q[43] /*67729*/;
assign _18388_ = _18389_ & D[3] /*67728*/;
assign _18391_ = _17860_ & _18388_ /*67723*/;
assign _18392_ = _17860_ ^ _18388_ /*67726*/;
assign _18393_ = _18384_ & _18392_ /*67724*/;
assign _18308_ = _18384_ ^ _18392_ /*67725*/;
assign _18390_ = _18391_ | _18393_ /*67722*/;
assign _18395_ = ~Q[43] /*67721*/;
assign _18394_ = _18395_ & D[4] /*67720*/;
assign _18397_ = _17861_ & _18394_ /*67715*/;
assign _18398_ = _17861_ ^ _18394_ /*67718*/;
assign _18399_ = _18390_ & _18398_ /*67716*/;
assign _18309_ = _18390_ ^ _18398_ /*67717*/;
assign _18396_ = _18397_ | _18399_ /*67714*/;
assign _18401_ = ~Q[43] /*67713*/;
assign _18400_ = _18401_ & D[5] /*67712*/;
assign _18403_ = _17862_ & _18400_ /*67707*/;
assign _18404_ = _17862_ ^ _18400_ /*67710*/;
assign _18405_ = _18396_ & _18404_ /*67708*/;
assign _18310_ = _18396_ ^ _18404_ /*67709*/;
assign _18402_ = _18403_ | _18405_ /*67706*/;
assign _18407_ = ~Q[43] /*67705*/;
assign _18406_ = _18407_ & D[6] /*67704*/;
assign _18409_ = _17863_ & _18406_ /*67699*/;
assign _18410_ = _17863_ ^ _18406_ /*67702*/;
assign _18411_ = _18402_ & _18410_ /*67700*/;
assign _18311_ = _18402_ ^ _18410_ /*67701*/;
assign _18408_ = _18409_ | _18411_ /*67698*/;
assign _18413_ = ~Q[43] /*67697*/;
assign _18412_ = _18413_ & D[7] /*67696*/;
assign _18415_ = _17864_ & _18412_ /*67691*/;
assign _18416_ = _17864_ ^ _18412_ /*67694*/;
assign _18417_ = _18408_ & _18416_ /*67692*/;
assign _18312_ = _18408_ ^ _18416_ /*67693*/;
assign _18414_ = _18415_ | _18417_ /*67690*/;
assign _18419_ = ~Q[43] /*67689*/;
assign _18418_ = _18419_ & D[8] /*67688*/;
assign _18421_ = _17865_ & _18418_ /*67683*/;
assign _18422_ = _17865_ ^ _18418_ /*67686*/;
assign _18423_ = _18414_ & _18422_ /*67684*/;
assign _18313_ = _18414_ ^ _18422_ /*67685*/;
assign _18420_ = _18421_ | _18423_ /*67682*/;
assign _18425_ = ~Q[43] /*67681*/;
assign _18424_ = _18425_ & D[9] /*67680*/;
assign _18427_ = _17866_ & _18424_ /*67675*/;
assign _18428_ = _17866_ ^ _18424_ /*67678*/;
assign _18429_ = _18420_ & _18428_ /*67676*/;
assign _18314_ = _18420_ ^ _18428_ /*67677*/;
assign _18426_ = _18427_ | _18429_ /*67674*/;
assign _18431_ = ~Q[43] /*67673*/;
assign _18430_ = _18431_ & D[10] /*67672*/;
assign _18433_ = _17867_ & _18430_ /*67667*/;
assign _18434_ = _17867_ ^ _18430_ /*67670*/;
assign _18435_ = _18426_ & _18434_ /*67668*/;
assign _18315_ = _18426_ ^ _18434_ /*67669*/;
assign _18432_ = _18433_ | _18435_ /*67666*/;
assign _18437_ = ~Q[43] /*67665*/;
assign _18436_ = _18437_ & D[11] /*67664*/;
assign _18439_ = _17868_ & _18436_ /*67659*/;
assign _18440_ = _17868_ ^ _18436_ /*67662*/;
assign _18441_ = _18432_ & _18440_ /*67660*/;
assign _18316_ = _18432_ ^ _18440_ /*67661*/;
assign _18438_ = _18439_ | _18441_ /*67658*/;
assign _18443_ = ~Q[43] /*67657*/;
assign _18442_ = _18443_ & D[12] /*67656*/;
assign _18445_ = _17869_ & _18442_ /*67651*/;
assign _18446_ = _17869_ ^ _18442_ /*67654*/;
assign _18447_ = _18438_ & _18446_ /*67652*/;
assign _18317_ = _18438_ ^ _18446_ /*67653*/;
assign _18444_ = _18445_ | _18447_ /*67650*/;
assign _18449_ = ~Q[43] /*67649*/;
assign _18448_ = _18449_ & D[13] /*67648*/;
assign _18451_ = _17870_ & _18448_ /*67643*/;
assign _18452_ = _17870_ ^ _18448_ /*67646*/;
assign _18453_ = _18444_ & _18452_ /*67644*/;
assign _18318_ = _18444_ ^ _18452_ /*67645*/;
assign _18450_ = _18451_ | _18453_ /*67642*/;
assign _18455_ = ~Q[43] /*67641*/;
assign _18454_ = _18455_ & D[14] /*67640*/;
assign _18457_ = _17871_ & _18454_ /*67635*/;
assign _18458_ = _17871_ ^ _18454_ /*67638*/;
assign _18459_ = _18450_ & _18458_ /*67636*/;
assign _18319_ = _18450_ ^ _18458_ /*67637*/;
assign _18456_ = _18457_ | _18459_ /*67634*/;
assign _18461_ = ~Q[43] /*67633*/;
assign _18460_ = _18461_ & D[15] /*67632*/;
assign _18463_ = _17872_ & _18460_ /*67627*/;
assign _18464_ = _17872_ ^ _18460_ /*67630*/;
assign _18465_ = _18456_ & _18464_ /*67628*/;
assign _18320_ = _18456_ ^ _18464_ /*67629*/;
assign _18462_ = _18463_ | _18465_ /*67626*/;
assign _18467_ = ~Q[43] /*67625*/;
assign _18466_ = _18467_ & D[16] /*67624*/;
assign _18469_ = _17873_ & _18466_ /*67619*/;
assign _18470_ = _17873_ ^ _18466_ /*67622*/;
assign _18471_ = _18462_ & _18470_ /*67620*/;
assign _18321_ = _18462_ ^ _18470_ /*67621*/;
assign _18468_ = _18469_ | _18471_ /*67618*/;
assign _18473_ = ~Q[43] /*67617*/;
assign _18472_ = _18473_ & D[17] /*67616*/;
assign _18475_ = _17874_ & _18472_ /*67611*/;
assign _18476_ = _17874_ ^ _18472_ /*67614*/;
assign _18477_ = _18468_ & _18476_ /*67612*/;
assign _18322_ = _18468_ ^ _18476_ /*67613*/;
assign _18474_ = _18475_ | _18477_ /*67610*/;
assign _18479_ = ~Q[43] /*67609*/;
assign _18478_ = _18479_ & D[18] /*67608*/;
assign _18481_ = _17875_ & _18478_ /*67603*/;
assign _18482_ = _17875_ ^ _18478_ /*67606*/;
assign _18483_ = _18474_ & _18482_ /*67604*/;
assign _18323_ = _18474_ ^ _18482_ /*67605*/;
assign _18480_ = _18481_ | _18483_ /*67602*/;
assign _18485_ = ~Q[43] /*67601*/;
assign _18484_ = _18485_ & D[19] /*67600*/;
assign _18487_ = _17876_ & _18484_ /*67595*/;
assign _18488_ = _17876_ ^ _18484_ /*67598*/;
assign _18489_ = _18480_ & _18488_ /*67596*/;
assign _18324_ = _18480_ ^ _18488_ /*67597*/;
assign _18486_ = _18487_ | _18489_ /*67594*/;
assign _18491_ = ~Q[43] /*67593*/;
assign _18490_ = _18491_ & D[20] /*67592*/;
assign _18493_ = _17877_ & _18490_ /*67587*/;
assign _18494_ = _17877_ ^ _18490_ /*67590*/;
assign _18495_ = _18486_ & _18494_ /*67588*/;
assign _18325_ = _18486_ ^ _18494_ /*67589*/;
assign _18492_ = _18493_ | _18495_ /*67586*/;
assign _18497_ = ~Q[43] /*67585*/;
assign _18496_ = _18497_ & D[21] /*67584*/;
assign _18499_ = _17878_ & _18496_ /*67579*/;
assign _18500_ = _17878_ ^ _18496_ /*67582*/;
assign _18501_ = _18492_ & _18500_ /*67580*/;
assign _18326_ = _18492_ ^ _18500_ /*67581*/;
assign _18498_ = _18499_ | _18501_ /*67578*/;
assign _18503_ = ~Q[43] /*67577*/;
assign _18502_ = _18503_ & D[22] /*67576*/;
assign _18505_ = _17879_ & _18502_ /*67571*/;
assign _18506_ = _17879_ ^ _18502_ /*67574*/;
assign _18507_ = _18498_ & _18506_ /*67572*/;
assign _18327_ = _18498_ ^ _18506_ /*67573*/;
assign _18504_ = _18505_ | _18507_ /*67570*/;
assign _18509_ = ~Q[43] /*67569*/;
assign _18508_ = _18509_ & D[23] /*67568*/;
assign _18511_ = _17880_ & _18508_ /*67563*/;
assign _18512_ = _17880_ ^ _18508_ /*67566*/;
assign _18513_ = _18504_ & _18512_ /*67564*/;
assign _18328_ = _18504_ ^ _18512_ /*67565*/;
assign _18510_ = _18511_ | _18513_ /*67562*/;
assign _18515_ = ~Q[43] /*67561*/;
assign _18514_ = _18515_ & D[24] /*67560*/;
assign _18517_ = _17881_ & _18514_ /*67555*/;
assign _18518_ = _17881_ ^ _18514_ /*67558*/;
assign _18519_ = _18510_ & _18518_ /*67556*/;
assign _18329_ = _18510_ ^ _18518_ /*67557*/;
assign _18516_ = _18517_ | _18519_ /*67554*/;
assign _18521_ = ~Q[43] /*67553*/;
assign _18520_ = _18521_ & D[25] /*67552*/;
assign _18523_ = _17882_ & _18520_ /*67547*/;
assign _18524_ = _17882_ ^ _18520_ /*67550*/;
assign _18525_ = _18516_ & _18524_ /*67548*/;
assign _18330_ = _18516_ ^ _18524_ /*67549*/;
assign _18522_ = _18523_ | _18525_ /*67546*/;
assign _18527_ = ~Q[43] /*67545*/;
assign _18526_ = _18527_ & D[26] /*67544*/;
assign _18529_ = _17883_ & _18526_ /*67539*/;
assign _18530_ = _17883_ ^ _18526_ /*67542*/;
assign _18531_ = _18522_ & _18530_ /*67540*/;
assign _18331_ = _18522_ ^ _18530_ /*67541*/;
assign _18528_ = _18529_ | _18531_ /*67538*/;
assign _18533_ = ~Q[43] /*67537*/;
assign _18532_ = _18533_ & D[27] /*67536*/;
assign _18535_ = _17884_ & _18532_ /*67531*/;
assign _18536_ = _17884_ ^ _18532_ /*67534*/;
assign _18537_ = _18528_ & _18536_ /*67532*/;
assign _18332_ = _18528_ ^ _18536_ /*67533*/;
assign _18534_ = _18535_ | _18537_ /*67530*/;
assign _18539_ = ~Q[43] /*67529*/;
assign _18538_ = _18539_ & D[28] /*67528*/;
assign _18541_ = _17885_ & _18538_ /*67523*/;
assign _18542_ = _17885_ ^ _18538_ /*67526*/;
assign _18543_ = _18534_ & _18542_ /*67524*/;
assign _18333_ = _18534_ ^ _18542_ /*67525*/;
assign _18540_ = _18541_ | _18543_ /*67522*/;
assign _18545_ = ~Q[43] /*67521*/;
assign _18544_ = _18545_ & D[29] /*67520*/;
assign _18547_ = _17886_ & _18544_ /*67515*/;
assign _18548_ = _17886_ ^ _18544_ /*67518*/;
assign _18549_ = _18540_ & _18548_ /*67516*/;
assign _18334_ = _18540_ ^ _18548_ /*67517*/;
assign _18546_ = _18547_ | _18549_ /*67514*/;
assign _18551_ = ~Q[43] /*67513*/;
assign _18550_ = _18551_ & D[30] /*67512*/;
assign _18553_ = _17887_ & _18550_ /*67507*/;
assign _18554_ = _17887_ ^ _18550_ /*67510*/;
assign _18555_ = _18546_ & _18554_ /*67508*/;
assign _18335_ = _18546_ ^ _18554_ /*67509*/;
assign _18552_ = _18553_ | _18555_ /*67506*/;
assign _18557_ = ~Q[43] /*67505*/;
assign _18556_ = _18557_ & D[31] /*67504*/;
assign _18559_ = _17888_ & _18556_ /*67499*/;
assign _18560_ = _17888_ ^ _18556_ /*67502*/;
assign _18561_ = _18552_ & _18560_ /*67500*/;
assign _18336_ = _18552_ ^ _18560_ /*67501*/;
assign _18558_ = _18559_ | _18561_ /*67498*/;
assign _18563_ = ~Q[43] /*67497*/;
assign _18562_ = _18563_ & D[32] /*67496*/;
assign _18565_ = _17889_ & _18562_ /*67491*/;
assign _18566_ = _17889_ ^ _18562_ /*67494*/;
assign _18567_ = _18558_ & _18566_ /*67492*/;
assign _18337_ = _18558_ ^ _18566_ /*67493*/;
assign _18564_ = _18565_ | _18567_ /*67490*/;
assign _18569_ = ~Q[43] /*67489*/;
assign _18568_ = _18569_ & D[33] /*67488*/;
assign _18571_ = _17890_ & _18568_ /*67483*/;
assign _18572_ = _17890_ ^ _18568_ /*67486*/;
assign _18573_ = _18564_ & _18572_ /*67484*/;
assign _18338_ = _18564_ ^ _18572_ /*67485*/;
assign _18570_ = _18571_ | _18573_ /*67482*/;
assign _18575_ = ~Q[43] /*67481*/;
assign _18574_ = _18575_ & D[34] /*67480*/;
assign _18577_ = _17891_ & _18574_ /*67475*/;
assign _18578_ = _17891_ ^ _18574_ /*67478*/;
assign _18579_ = _18570_ & _18578_ /*67476*/;
assign _18339_ = _18570_ ^ _18578_ /*67477*/;
assign _18576_ = _18577_ | _18579_ /*67474*/;
assign _18581_ = ~Q[43] /*67473*/;
assign _18580_ = _18581_ & D[35] /*67472*/;
assign _18583_ = _17892_ & _18580_ /*67467*/;
assign _18584_ = _17892_ ^ _18580_ /*67470*/;
assign _18585_ = _18576_ & _18584_ /*67468*/;
assign _18340_ = _18576_ ^ _18584_ /*67469*/;
assign _18582_ = _18583_ | _18585_ /*67466*/;
assign _18587_ = ~Q[43] /*67465*/;
assign _18586_ = _18587_ & D[36] /*67464*/;
assign _18589_ = _17893_ & _18586_ /*67459*/;
assign _18590_ = _17893_ ^ _18586_ /*67462*/;
assign _18591_ = _18582_ & _18590_ /*67460*/;
assign _18341_ = _18582_ ^ _18590_ /*67461*/;
assign _18588_ = _18589_ | _18591_ /*67458*/;
assign _18593_ = ~Q[43] /*67457*/;
assign _18592_ = _18593_ & D[37] /*67456*/;
assign _18595_ = _17894_ & _18592_ /*67451*/;
assign _18596_ = _17894_ ^ _18592_ /*67454*/;
assign _18597_ = _18588_ & _18596_ /*67452*/;
assign _18342_ = _18588_ ^ _18596_ /*67453*/;
assign _18594_ = _18595_ | _18597_ /*67450*/;
assign _18599_ = ~Q[43] /*67449*/;
assign _18598_ = _18599_ & D[38] /*67448*/;
assign _18601_ = _17895_ & _18598_ /*67443*/;
assign _18602_ = _17895_ ^ _18598_ /*67446*/;
assign _18603_ = _18594_ & _18602_ /*67444*/;
assign _18343_ = _18594_ ^ _18602_ /*67445*/;
assign _18600_ = _18601_ | _18603_ /*67442*/;
assign _18605_ = ~Q[43] /*67441*/;
assign _18604_ = _18605_ & D[39] /*67440*/;
assign _18607_ = _17896_ & _18604_ /*67435*/;
assign _18608_ = _17896_ ^ _18604_ /*67438*/;
assign _18609_ = _18600_ & _18608_ /*67436*/;
assign _18344_ = _18600_ ^ _18608_ /*67437*/;
assign _18606_ = _18607_ | _18609_ /*67434*/;
assign _18611_ = ~Q[43] /*67433*/;
assign _18610_ = _18611_ & D[40] /*67432*/;
assign _18613_ = _17897_ & _18610_ /*67427*/;
assign _18614_ = _17897_ ^ _18610_ /*67430*/;
assign _18615_ = _18606_ & _18614_ /*67428*/;
assign _18345_ = _18606_ ^ _18614_ /*67429*/;
assign _18612_ = _18613_ | _18615_ /*67426*/;
assign _18617_ = ~Q[43] /*67425*/;
assign _18616_ = _18617_ & D[41] /*67424*/;
assign _18619_ = _17898_ & _18616_ /*67419*/;
assign _18620_ = _17898_ ^ _18616_ /*67422*/;
assign _18621_ = _18612_ & _18620_ /*67420*/;
assign _18346_ = _18612_ ^ _18620_ /*67421*/;
assign _18618_ = _18619_ | _18621_ /*67418*/;
assign _18623_ = ~Q[43] /*67417*/;
assign _18622_ = _18623_ & D[42] /*67416*/;
assign _18625_ = _17899_ & _18622_ /*67411*/;
assign _18626_ = _17899_ ^ _18622_ /*67414*/;
assign _18627_ = _18618_ & _18626_ /*67412*/;
assign _18347_ = _18618_ ^ _18626_ /*67413*/;
assign _18624_ = _18625_ | _18627_ /*67410*/;
assign _18629_ = ~Q[43] /*67409*/;
assign _18628_ = _18629_ & D[43] /*67408*/;
assign _18631_ = _17900_ & _18628_ /*67403*/;
assign _18632_ = _17900_ ^ _18628_ /*67406*/;
assign _18633_ = _18624_ & _18632_ /*67404*/;
assign _18348_ = _18624_ ^ _18632_ /*67405*/;
assign _18630_ = _18631_ | _18633_ /*67402*/;
assign _18635_ = ~Q[43] /*67401*/;
assign _18634_ = _18635_ & D[44] /*67400*/;
assign _18637_ = _17901_ & _18634_ /*67395*/;
assign _18638_ = _17901_ ^ _18634_ /*67398*/;
assign _18639_ = _18630_ & _18638_ /*67396*/;
assign _18349_ = _18630_ ^ _18638_ /*67397*/;
assign _18636_ = _18637_ | _18639_ /*67394*/;
assign _18641_ = ~Q[43] /*67393*/;
assign _18640_ = _18641_ & D[45] /*67392*/;
assign _18643_ = _17902_ & _18640_ /*67387*/;
assign _18644_ = _17902_ ^ _18640_ /*67390*/;
assign _18645_ = _18636_ & _18644_ /*67388*/;
assign _18350_ = _18636_ ^ _18644_ /*67389*/;
assign _18642_ = _18643_ | _18645_ /*67386*/;
assign _18647_ = ~Q[43] /*67385*/;
assign _18646_ = _18647_ & D[46] /*67384*/;
assign _18649_ = _17903_ & _18646_ /*67379*/;
assign _18650_ = _17903_ ^ _18646_ /*67382*/;
assign _18651_ = _18642_ & _18650_ /*67380*/;
assign _18351_ = _18642_ ^ _18650_ /*67381*/;
assign _18648_ = _18649_ | _18651_ /*67378*/;
assign _18653_ = ~Q[43] /*67377*/;
assign _18652_ = _18653_ & D[47] /*67376*/;
assign _18655_ = _17904_ & _18652_ /*67371*/;
assign _18656_ = _17904_ ^ _18652_ /*67374*/;
assign _18657_ = _18648_ & _18656_ /*67372*/;
assign _18352_ = _18648_ ^ _18656_ /*67373*/;
assign _18654_ = _18655_ | _18657_ /*67370*/;
assign _18659_ = ~Q[43] /*67369*/;
assign _18658_ = _18659_ & D[48] /*67368*/;
assign _18661_ = _17905_ & _18658_ /*67363*/;
assign _18662_ = _17905_ ^ _18658_ /*67366*/;
assign _18663_ = _18654_ & _18662_ /*67364*/;
assign _18353_ = _18654_ ^ _18662_ /*67365*/;
assign _18660_ = _18661_ | _18663_ /*67362*/;
assign _18665_ = ~Q[43] /*67361*/;
assign _18664_ = _18665_ & D[49] /*67360*/;
assign _18667_ = _17906_ & _18664_ /*67355*/;
assign _18668_ = _17906_ ^ _18664_ /*67358*/;
assign _18669_ = _18660_ & _18668_ /*67356*/;
assign _18354_ = _18660_ ^ _18668_ /*67357*/;
assign _18666_ = _18667_ | _18669_ /*67354*/;
assign _18671_ = ~Q[43] /*67353*/;
assign _18670_ = _18671_ & D[50] /*67352*/;
assign _18673_ = _17907_ & _18670_ /*67347*/;
assign _18674_ = _17907_ ^ _18670_ /*67350*/;
assign _18675_ = _18666_ & _18674_ /*67348*/;
assign _18355_ = _18666_ ^ _18674_ /*67349*/;
assign _18672_ = _18673_ | _18675_ /*67346*/;
assign _18677_ = ~Q[43] /*67345*/;
assign _18676_ = _18677_ & D[51] /*67344*/;
assign _18679_ = _17908_ & _18676_ /*67339*/;
assign _18680_ = _17908_ ^ _18676_ /*67342*/;
assign _18681_ = _18672_ & _18680_ /*67340*/;
assign _18356_ = _18672_ ^ _18680_ /*67341*/;
assign _18678_ = _18679_ | _18681_ /*67338*/;
assign _18683_ = ~Q[43] /*67337*/;
assign _18682_ = _18683_ & D[52] /*67336*/;
assign _18685_ = _17909_ & _18682_ /*67331*/;
assign _18686_ = _17909_ ^ _18682_ /*67334*/;
assign _18687_ = _18678_ & _18686_ /*67332*/;
assign _18357_ = _18678_ ^ _18686_ /*67333*/;
assign _18684_ = _18685_ | _18687_ /*67330*/;
assign _18689_ = ~Q[43] /*67329*/;
assign _18688_ = _18689_ & D[53] /*67328*/;
assign _18691_ = _17910_ & _18688_ /*67323*/;
assign _18692_ = _17910_ ^ _18688_ /*67326*/;
assign _18693_ = _18684_ & _18692_ /*67324*/;
assign _18358_ = _18684_ ^ _18692_ /*67325*/;
assign _18690_ = _18691_ | _18693_ /*67322*/;
assign _18695_ = ~Q[43] /*67321*/;
assign _18694_ = _18695_ & D[54] /*67320*/;
assign _18697_ = _17911_ & _18694_ /*67315*/;
assign _18698_ = _17911_ ^ _18694_ /*67318*/;
assign _18699_ = _18690_ & _18698_ /*67316*/;
assign _18359_ = _18690_ ^ _18698_ /*67317*/;
assign _18696_ = _18697_ | _18699_ /*67314*/;
assign _18701_ = ~Q[43] /*67313*/;
assign _18700_ = _18701_ & D[55] /*67312*/;
assign _18703_ = _17912_ & _18700_ /*67307*/;
assign _18704_ = _17912_ ^ _18700_ /*67310*/;
assign _18705_ = _18696_ & _18704_ /*67308*/;
assign _18360_ = _18696_ ^ _18704_ /*67309*/;
assign _18702_ = _18703_ | _18705_ /*67306*/;
assign _18707_ = ~Q[43] /*67305*/;
assign _18706_ = _18707_ & D[56] /*67304*/;
assign _18709_ = _17913_ & _18706_ /*67299*/;
assign _18710_ = _17913_ ^ _18706_ /*67302*/;
assign _18711_ = _18702_ & _18710_ /*67300*/;
assign _18361_ = _18702_ ^ _18710_ /*67301*/;
assign _18708_ = _18709_ | _18711_ /*67298*/;
assign _18713_ = ~Q[43] /*67297*/;
assign _18712_ = _18713_ & D[57] /*67296*/;
assign _18715_ = _17914_ & _18712_ /*67291*/;
assign _18716_ = _17914_ ^ _18712_ /*67294*/;
assign _18717_ = _18708_ & _18716_ /*67292*/;
assign _18362_ = _18708_ ^ _18716_ /*67293*/;
assign _18714_ = _18715_ | _18717_ /*67290*/;
assign _18719_ = ~Q[43] /*67289*/;
assign _18718_ = _18719_ & D[58] /*67288*/;
assign _18721_ = _17915_ & _18718_ /*67283*/;
assign _18722_ = _17915_ ^ _18718_ /*67286*/;
assign _18723_ = _18714_ & _18722_ /*67284*/;
assign _18363_ = _18714_ ^ _18722_ /*67285*/;
assign _18720_ = _18721_ | _18723_ /*67282*/;
assign _18725_ = ~Q[43] /*67281*/;
assign _18724_ = _18725_ & D[59] /*67280*/;
assign _18727_ = _17916_ & _18724_ /*67275*/;
assign _18728_ = _17916_ ^ _18724_ /*67278*/;
assign _18729_ = _18720_ & _18728_ /*67276*/;
assign _18364_ = _18720_ ^ _18728_ /*67277*/;
assign _18726_ = _18727_ | _18729_ /*67274*/;
assign _18731_ = ~Q[43] /*67273*/;
assign _18730_ = _18731_ & D[60] /*67272*/;
assign _18733_ = _17917_ & _18730_ /*67267*/;
assign _18734_ = _17917_ ^ _18730_ /*67270*/;
assign _18735_ = _18726_ & _18734_ /*67268*/;
assign _18365_ = _18726_ ^ _18734_ /*67269*/;
assign _18732_ = _18733_ | _18735_ /*67266*/;
assign _18737_ = ~Q[43] /*67265*/;
assign _18736_ = _18737_ & D[61] /*67264*/;
assign _18739_ = _17918_ & _18736_ /*67259*/;
assign _18740_ = _17918_ ^ _18736_ /*67262*/;
assign _18741_ = _18732_ & _18740_ /*67260*/;
assign _18366_ = _18732_ ^ _18740_ /*67261*/;
assign _18738_ = _18739_ | _18741_ /*67258*/;
assign _18743_ = ~Q[43] /*67257*/;
assign _18742_ = _18743_ & D[62] /*67256*/;
assign _18745_ = _17919_ & _18742_ /*67251*/;
assign _18746_ = _17919_ ^ _18742_ /*67254*/;
assign _18747_ = _18738_ & _18746_ /*67252*/;
assign _18367_ = _18738_ ^ _18746_ /*67253*/;
assign _18744_ = _18745_ | _18747_ /*67250*/;
assign _18749_ = ~Q[43] /*67249*/;
assign _18748_ = _18749_ & zeroWire /*67248*/;
assign _18750_ = _17920_ ^ _18748_ /*67246*/;
assign _18368_ = _18750_ ^ _18744_ /*67245*/;
assign _18821_ = ~D[0] /*66991*/;
assign _18818_ = R_0[42] & _18821_ /*66987*/;
assign _18819_ = R_0[42] ^ _18821_ /*66990*/;
assign _18820_ = oneWire & _18819_ /*66988*/;
assign _18753_ = oneWire ^ _18819_ /*66989*/;
assign _18817_ = _18818_ | _18820_ /*66986*/;
assign _18826_ = ~D[1] /*66985*/;
assign _18823_ = _18305_ & _18826_ /*66981*/;
assign _18824_ = _18305_ ^ _18826_ /*66984*/;
assign _18825_ = _18817_ & _18824_ /*66982*/;
assign _18754_ = _18817_ ^ _18824_ /*66983*/;
assign _18822_ = _18823_ | _18825_ /*66980*/;
assign _18831_ = ~D[2] /*66979*/;
assign _18828_ = _18306_ & _18831_ /*66975*/;
assign _18829_ = _18306_ ^ _18831_ /*66978*/;
assign _18830_ = _18822_ & _18829_ /*66976*/;
assign _18755_ = _18822_ ^ _18829_ /*66977*/;
assign _18827_ = _18828_ | _18830_ /*66974*/;
assign _18836_ = ~D[3] /*66973*/;
assign _18833_ = _18307_ & _18836_ /*66969*/;
assign _18834_ = _18307_ ^ _18836_ /*66972*/;
assign _18835_ = _18827_ & _18834_ /*66970*/;
assign _18756_ = _18827_ ^ _18834_ /*66971*/;
assign _18832_ = _18833_ | _18835_ /*66968*/;
assign _18841_ = ~D[4] /*66967*/;
assign _18838_ = _18308_ & _18841_ /*66963*/;
assign _18839_ = _18308_ ^ _18841_ /*66966*/;
assign _18840_ = _18832_ & _18839_ /*66964*/;
assign _18757_ = _18832_ ^ _18839_ /*66965*/;
assign _18837_ = _18838_ | _18840_ /*66962*/;
assign _18846_ = ~D[5] /*66961*/;
assign _18843_ = _18309_ & _18846_ /*66957*/;
assign _18844_ = _18309_ ^ _18846_ /*66960*/;
assign _18845_ = _18837_ & _18844_ /*66958*/;
assign _18758_ = _18837_ ^ _18844_ /*66959*/;
assign _18842_ = _18843_ | _18845_ /*66956*/;
assign _18851_ = ~D[6] /*66955*/;
assign _18848_ = _18310_ & _18851_ /*66951*/;
assign _18849_ = _18310_ ^ _18851_ /*66954*/;
assign _18850_ = _18842_ & _18849_ /*66952*/;
assign _18759_ = _18842_ ^ _18849_ /*66953*/;
assign _18847_ = _18848_ | _18850_ /*66950*/;
assign _18856_ = ~D[7] /*66949*/;
assign _18853_ = _18311_ & _18856_ /*66945*/;
assign _18854_ = _18311_ ^ _18856_ /*66948*/;
assign _18855_ = _18847_ & _18854_ /*66946*/;
assign _18760_ = _18847_ ^ _18854_ /*66947*/;
assign _18852_ = _18853_ | _18855_ /*66944*/;
assign _18861_ = ~D[8] /*66943*/;
assign _18858_ = _18312_ & _18861_ /*66939*/;
assign _18859_ = _18312_ ^ _18861_ /*66942*/;
assign _18860_ = _18852_ & _18859_ /*66940*/;
assign _18761_ = _18852_ ^ _18859_ /*66941*/;
assign _18857_ = _18858_ | _18860_ /*66938*/;
assign _18866_ = ~D[9] /*66937*/;
assign _18863_ = _18313_ & _18866_ /*66933*/;
assign _18864_ = _18313_ ^ _18866_ /*66936*/;
assign _18865_ = _18857_ & _18864_ /*66934*/;
assign _18762_ = _18857_ ^ _18864_ /*66935*/;
assign _18862_ = _18863_ | _18865_ /*66932*/;
assign _18871_ = ~D[10] /*66931*/;
assign _18868_ = _18314_ & _18871_ /*66927*/;
assign _18869_ = _18314_ ^ _18871_ /*66930*/;
assign _18870_ = _18862_ & _18869_ /*66928*/;
assign _18763_ = _18862_ ^ _18869_ /*66929*/;
assign _18867_ = _18868_ | _18870_ /*66926*/;
assign _18876_ = ~D[11] /*66925*/;
assign _18873_ = _18315_ & _18876_ /*66921*/;
assign _18874_ = _18315_ ^ _18876_ /*66924*/;
assign _18875_ = _18867_ & _18874_ /*66922*/;
assign _18764_ = _18867_ ^ _18874_ /*66923*/;
assign _18872_ = _18873_ | _18875_ /*66920*/;
assign _18881_ = ~D[12] /*66919*/;
assign _18878_ = _18316_ & _18881_ /*66915*/;
assign _18879_ = _18316_ ^ _18881_ /*66918*/;
assign _18880_ = _18872_ & _18879_ /*66916*/;
assign _18765_ = _18872_ ^ _18879_ /*66917*/;
assign _18877_ = _18878_ | _18880_ /*66914*/;
assign _18886_ = ~D[13] /*66913*/;
assign _18883_ = _18317_ & _18886_ /*66909*/;
assign _18884_ = _18317_ ^ _18886_ /*66912*/;
assign _18885_ = _18877_ & _18884_ /*66910*/;
assign _18766_ = _18877_ ^ _18884_ /*66911*/;
assign _18882_ = _18883_ | _18885_ /*66908*/;
assign _18891_ = ~D[14] /*66907*/;
assign _18888_ = _18318_ & _18891_ /*66903*/;
assign _18889_ = _18318_ ^ _18891_ /*66906*/;
assign _18890_ = _18882_ & _18889_ /*66904*/;
assign _18767_ = _18882_ ^ _18889_ /*66905*/;
assign _18887_ = _18888_ | _18890_ /*66902*/;
assign _18896_ = ~D[15] /*66901*/;
assign _18893_ = _18319_ & _18896_ /*66897*/;
assign _18894_ = _18319_ ^ _18896_ /*66900*/;
assign _18895_ = _18887_ & _18894_ /*66898*/;
assign _18768_ = _18887_ ^ _18894_ /*66899*/;
assign _18892_ = _18893_ | _18895_ /*66896*/;
assign _18901_ = ~D[16] /*66895*/;
assign _18898_ = _18320_ & _18901_ /*66891*/;
assign _18899_ = _18320_ ^ _18901_ /*66894*/;
assign _18900_ = _18892_ & _18899_ /*66892*/;
assign _18769_ = _18892_ ^ _18899_ /*66893*/;
assign _18897_ = _18898_ | _18900_ /*66890*/;
assign _18906_ = ~D[17] /*66889*/;
assign _18903_ = _18321_ & _18906_ /*66885*/;
assign _18904_ = _18321_ ^ _18906_ /*66888*/;
assign _18905_ = _18897_ & _18904_ /*66886*/;
assign _18770_ = _18897_ ^ _18904_ /*66887*/;
assign _18902_ = _18903_ | _18905_ /*66884*/;
assign _18911_ = ~D[18] /*66883*/;
assign _18908_ = _18322_ & _18911_ /*66879*/;
assign _18909_ = _18322_ ^ _18911_ /*66882*/;
assign _18910_ = _18902_ & _18909_ /*66880*/;
assign _18771_ = _18902_ ^ _18909_ /*66881*/;
assign _18907_ = _18908_ | _18910_ /*66878*/;
assign _18916_ = ~D[19] /*66877*/;
assign _18913_ = _18323_ & _18916_ /*66873*/;
assign _18914_ = _18323_ ^ _18916_ /*66876*/;
assign _18915_ = _18907_ & _18914_ /*66874*/;
assign _18772_ = _18907_ ^ _18914_ /*66875*/;
assign _18912_ = _18913_ | _18915_ /*66872*/;
assign _18921_ = ~D[20] /*66871*/;
assign _18918_ = _18324_ & _18921_ /*66867*/;
assign _18919_ = _18324_ ^ _18921_ /*66870*/;
assign _18920_ = _18912_ & _18919_ /*66868*/;
assign _18773_ = _18912_ ^ _18919_ /*66869*/;
assign _18917_ = _18918_ | _18920_ /*66866*/;
assign _18926_ = ~D[21] /*66865*/;
assign _18923_ = _18325_ & _18926_ /*66861*/;
assign _18924_ = _18325_ ^ _18926_ /*66864*/;
assign _18925_ = _18917_ & _18924_ /*66862*/;
assign _18774_ = _18917_ ^ _18924_ /*66863*/;
assign _18922_ = _18923_ | _18925_ /*66860*/;
assign _18931_ = ~D[22] /*66859*/;
assign _18928_ = _18326_ & _18931_ /*66855*/;
assign _18929_ = _18326_ ^ _18931_ /*66858*/;
assign _18930_ = _18922_ & _18929_ /*66856*/;
assign _18775_ = _18922_ ^ _18929_ /*66857*/;
assign _18927_ = _18928_ | _18930_ /*66854*/;
assign _18936_ = ~D[23] /*66853*/;
assign _18933_ = _18327_ & _18936_ /*66849*/;
assign _18934_ = _18327_ ^ _18936_ /*66852*/;
assign _18935_ = _18927_ & _18934_ /*66850*/;
assign _18776_ = _18927_ ^ _18934_ /*66851*/;
assign _18932_ = _18933_ | _18935_ /*66848*/;
assign _18941_ = ~D[24] /*66847*/;
assign _18938_ = _18328_ & _18941_ /*66843*/;
assign _18939_ = _18328_ ^ _18941_ /*66846*/;
assign _18940_ = _18932_ & _18939_ /*66844*/;
assign _18777_ = _18932_ ^ _18939_ /*66845*/;
assign _18937_ = _18938_ | _18940_ /*66842*/;
assign _18946_ = ~D[25] /*66841*/;
assign _18943_ = _18329_ & _18946_ /*66837*/;
assign _18944_ = _18329_ ^ _18946_ /*66840*/;
assign _18945_ = _18937_ & _18944_ /*66838*/;
assign _18778_ = _18937_ ^ _18944_ /*66839*/;
assign _18942_ = _18943_ | _18945_ /*66836*/;
assign _18951_ = ~D[26] /*66835*/;
assign _18948_ = _18330_ & _18951_ /*66831*/;
assign _18949_ = _18330_ ^ _18951_ /*66834*/;
assign _18950_ = _18942_ & _18949_ /*66832*/;
assign _18779_ = _18942_ ^ _18949_ /*66833*/;
assign _18947_ = _18948_ | _18950_ /*66830*/;
assign _18956_ = ~D[27] /*66829*/;
assign _18953_ = _18331_ & _18956_ /*66825*/;
assign _18954_ = _18331_ ^ _18956_ /*66828*/;
assign _18955_ = _18947_ & _18954_ /*66826*/;
assign _18780_ = _18947_ ^ _18954_ /*66827*/;
assign _18952_ = _18953_ | _18955_ /*66824*/;
assign _18961_ = ~D[28] /*66823*/;
assign _18958_ = _18332_ & _18961_ /*66819*/;
assign _18959_ = _18332_ ^ _18961_ /*66822*/;
assign _18960_ = _18952_ & _18959_ /*66820*/;
assign _18781_ = _18952_ ^ _18959_ /*66821*/;
assign _18957_ = _18958_ | _18960_ /*66818*/;
assign _18966_ = ~D[29] /*66817*/;
assign _18963_ = _18333_ & _18966_ /*66813*/;
assign _18964_ = _18333_ ^ _18966_ /*66816*/;
assign _18965_ = _18957_ & _18964_ /*66814*/;
assign _18782_ = _18957_ ^ _18964_ /*66815*/;
assign _18962_ = _18963_ | _18965_ /*66812*/;
assign _18971_ = ~D[30] /*66811*/;
assign _18968_ = _18334_ & _18971_ /*66807*/;
assign _18969_ = _18334_ ^ _18971_ /*66810*/;
assign _18970_ = _18962_ & _18969_ /*66808*/;
assign _18783_ = _18962_ ^ _18969_ /*66809*/;
assign _18967_ = _18968_ | _18970_ /*66806*/;
assign _18976_ = ~D[31] /*66805*/;
assign _18973_ = _18335_ & _18976_ /*66801*/;
assign _18974_ = _18335_ ^ _18976_ /*66804*/;
assign _18975_ = _18967_ & _18974_ /*66802*/;
assign _18784_ = _18967_ ^ _18974_ /*66803*/;
assign _18972_ = _18973_ | _18975_ /*66800*/;
assign _18981_ = ~D[32] /*66799*/;
assign _18978_ = _18336_ & _18981_ /*66795*/;
assign _18979_ = _18336_ ^ _18981_ /*66798*/;
assign _18980_ = _18972_ & _18979_ /*66796*/;
assign _18785_ = _18972_ ^ _18979_ /*66797*/;
assign _18977_ = _18978_ | _18980_ /*66794*/;
assign _18986_ = ~D[33] /*66793*/;
assign _18983_ = _18337_ & _18986_ /*66789*/;
assign _18984_ = _18337_ ^ _18986_ /*66792*/;
assign _18985_ = _18977_ & _18984_ /*66790*/;
assign _18786_ = _18977_ ^ _18984_ /*66791*/;
assign _18982_ = _18983_ | _18985_ /*66788*/;
assign _18991_ = ~D[34] /*66787*/;
assign _18988_ = _18338_ & _18991_ /*66783*/;
assign _18989_ = _18338_ ^ _18991_ /*66786*/;
assign _18990_ = _18982_ & _18989_ /*66784*/;
assign _18787_ = _18982_ ^ _18989_ /*66785*/;
assign _18987_ = _18988_ | _18990_ /*66782*/;
assign _18996_ = ~D[35] /*66781*/;
assign _18993_ = _18339_ & _18996_ /*66777*/;
assign _18994_ = _18339_ ^ _18996_ /*66780*/;
assign _18995_ = _18987_ & _18994_ /*66778*/;
assign _18788_ = _18987_ ^ _18994_ /*66779*/;
assign _18992_ = _18993_ | _18995_ /*66776*/;
assign _19001_ = ~D[36] /*66775*/;
assign _18998_ = _18340_ & _19001_ /*66771*/;
assign _18999_ = _18340_ ^ _19001_ /*66774*/;
assign _19000_ = _18992_ & _18999_ /*66772*/;
assign _18789_ = _18992_ ^ _18999_ /*66773*/;
assign _18997_ = _18998_ | _19000_ /*66770*/;
assign _19006_ = ~D[37] /*66769*/;
assign _19003_ = _18341_ & _19006_ /*66765*/;
assign _19004_ = _18341_ ^ _19006_ /*66768*/;
assign _19005_ = _18997_ & _19004_ /*66766*/;
assign _18790_ = _18997_ ^ _19004_ /*66767*/;
assign _19002_ = _19003_ | _19005_ /*66764*/;
assign _19011_ = ~D[38] /*66763*/;
assign _19008_ = _18342_ & _19011_ /*66759*/;
assign _19009_ = _18342_ ^ _19011_ /*66762*/;
assign _19010_ = _19002_ & _19009_ /*66760*/;
assign _18791_ = _19002_ ^ _19009_ /*66761*/;
assign _19007_ = _19008_ | _19010_ /*66758*/;
assign _19016_ = ~D[39] /*66757*/;
assign _19013_ = _18343_ & _19016_ /*66753*/;
assign _19014_ = _18343_ ^ _19016_ /*66756*/;
assign _19015_ = _19007_ & _19014_ /*66754*/;
assign _18792_ = _19007_ ^ _19014_ /*66755*/;
assign _19012_ = _19013_ | _19015_ /*66752*/;
assign _19021_ = ~D[40] /*66751*/;
assign _19018_ = _18344_ & _19021_ /*66747*/;
assign _19019_ = _18344_ ^ _19021_ /*66750*/;
assign _19020_ = _19012_ & _19019_ /*66748*/;
assign _18793_ = _19012_ ^ _19019_ /*66749*/;
assign _19017_ = _19018_ | _19020_ /*66746*/;
assign _19026_ = ~D[41] /*66745*/;
assign _19023_ = _18345_ & _19026_ /*66741*/;
assign _19024_ = _18345_ ^ _19026_ /*66744*/;
assign _19025_ = _19017_ & _19024_ /*66742*/;
assign _18794_ = _19017_ ^ _19024_ /*66743*/;
assign _19022_ = _19023_ | _19025_ /*66740*/;
assign _19031_ = ~D[42] /*66739*/;
assign _19028_ = _18346_ & _19031_ /*66735*/;
assign _19029_ = _18346_ ^ _19031_ /*66738*/;
assign _19030_ = _19022_ & _19029_ /*66736*/;
assign _18795_ = _19022_ ^ _19029_ /*66737*/;
assign _19027_ = _19028_ | _19030_ /*66734*/;
assign _19036_ = ~D[43] /*66733*/;
assign _19033_ = _18347_ & _19036_ /*66729*/;
assign _19034_ = _18347_ ^ _19036_ /*66732*/;
assign _19035_ = _19027_ & _19034_ /*66730*/;
assign _18796_ = _19027_ ^ _19034_ /*66731*/;
assign _19032_ = _19033_ | _19035_ /*66728*/;
assign _19041_ = ~D[44] /*66727*/;
assign _19038_ = _18348_ & _19041_ /*66723*/;
assign _19039_ = _18348_ ^ _19041_ /*66726*/;
assign _19040_ = _19032_ & _19039_ /*66724*/;
assign _18797_ = _19032_ ^ _19039_ /*66725*/;
assign _19037_ = _19038_ | _19040_ /*66722*/;
assign _19046_ = ~D[45] /*66721*/;
assign _19043_ = _18349_ & _19046_ /*66717*/;
assign _19044_ = _18349_ ^ _19046_ /*66720*/;
assign _19045_ = _19037_ & _19044_ /*66718*/;
assign _18798_ = _19037_ ^ _19044_ /*66719*/;
assign _19042_ = _19043_ | _19045_ /*66716*/;
assign _19051_ = ~D[46] /*66715*/;
assign _19048_ = _18350_ & _19051_ /*66711*/;
assign _19049_ = _18350_ ^ _19051_ /*66714*/;
assign _19050_ = _19042_ & _19049_ /*66712*/;
assign _18799_ = _19042_ ^ _19049_ /*66713*/;
assign _19047_ = _19048_ | _19050_ /*66710*/;
assign _19056_ = ~D[47] /*66709*/;
assign _19053_ = _18351_ & _19056_ /*66705*/;
assign _19054_ = _18351_ ^ _19056_ /*66708*/;
assign _19055_ = _19047_ & _19054_ /*66706*/;
assign _18800_ = _19047_ ^ _19054_ /*66707*/;
assign _19052_ = _19053_ | _19055_ /*66704*/;
assign _19061_ = ~D[48] /*66703*/;
assign _19058_ = _18352_ & _19061_ /*66699*/;
assign _19059_ = _18352_ ^ _19061_ /*66702*/;
assign _19060_ = _19052_ & _19059_ /*66700*/;
assign _18801_ = _19052_ ^ _19059_ /*66701*/;
assign _19057_ = _19058_ | _19060_ /*66698*/;
assign _19066_ = ~D[49] /*66697*/;
assign _19063_ = _18353_ & _19066_ /*66693*/;
assign _19064_ = _18353_ ^ _19066_ /*66696*/;
assign _19065_ = _19057_ & _19064_ /*66694*/;
assign _18802_ = _19057_ ^ _19064_ /*66695*/;
assign _19062_ = _19063_ | _19065_ /*66692*/;
assign _19071_ = ~D[50] /*66691*/;
assign _19068_ = _18354_ & _19071_ /*66687*/;
assign _19069_ = _18354_ ^ _19071_ /*66690*/;
assign _19070_ = _19062_ & _19069_ /*66688*/;
assign _18803_ = _19062_ ^ _19069_ /*66689*/;
assign _19067_ = _19068_ | _19070_ /*66686*/;
assign _19076_ = ~D[51] /*66685*/;
assign _19073_ = _18355_ & _19076_ /*66681*/;
assign _19074_ = _18355_ ^ _19076_ /*66684*/;
assign _19075_ = _19067_ & _19074_ /*66682*/;
assign _18804_ = _19067_ ^ _19074_ /*66683*/;
assign _19072_ = _19073_ | _19075_ /*66680*/;
assign _19081_ = ~D[52] /*66679*/;
assign _19078_ = _18356_ & _19081_ /*66675*/;
assign _19079_ = _18356_ ^ _19081_ /*66678*/;
assign _19080_ = _19072_ & _19079_ /*66676*/;
assign _18805_ = _19072_ ^ _19079_ /*66677*/;
assign _19077_ = _19078_ | _19080_ /*66674*/;
assign _19086_ = ~D[53] /*66673*/;
assign _19083_ = _18357_ & _19086_ /*66669*/;
assign _19084_ = _18357_ ^ _19086_ /*66672*/;
assign _19085_ = _19077_ & _19084_ /*66670*/;
assign _18806_ = _19077_ ^ _19084_ /*66671*/;
assign _19082_ = _19083_ | _19085_ /*66668*/;
assign _19091_ = ~D[54] /*66667*/;
assign _19088_ = _18358_ & _19091_ /*66663*/;
assign _19089_ = _18358_ ^ _19091_ /*66666*/;
assign _19090_ = _19082_ & _19089_ /*66664*/;
assign _18807_ = _19082_ ^ _19089_ /*66665*/;
assign _19087_ = _19088_ | _19090_ /*66662*/;
assign _19096_ = ~D[55] /*66661*/;
assign _19093_ = _18359_ & _19096_ /*66657*/;
assign _19094_ = _18359_ ^ _19096_ /*66660*/;
assign _19095_ = _19087_ & _19094_ /*66658*/;
assign _18808_ = _19087_ ^ _19094_ /*66659*/;
assign _19092_ = _19093_ | _19095_ /*66656*/;
assign _19101_ = ~D[56] /*66655*/;
assign _19098_ = _18360_ & _19101_ /*66651*/;
assign _19099_ = _18360_ ^ _19101_ /*66654*/;
assign _19100_ = _19092_ & _19099_ /*66652*/;
assign _18809_ = _19092_ ^ _19099_ /*66653*/;
assign _19097_ = _19098_ | _19100_ /*66650*/;
assign _19106_ = ~D[57] /*66649*/;
assign _19103_ = _18361_ & _19106_ /*66645*/;
assign _19104_ = _18361_ ^ _19106_ /*66648*/;
assign _19105_ = _19097_ & _19104_ /*66646*/;
assign _18810_ = _19097_ ^ _19104_ /*66647*/;
assign _19102_ = _19103_ | _19105_ /*66644*/;
assign _19111_ = ~D[58] /*66643*/;
assign _19108_ = _18362_ & _19111_ /*66639*/;
assign _19109_ = _18362_ ^ _19111_ /*66642*/;
assign _19110_ = _19102_ & _19109_ /*66640*/;
assign _18811_ = _19102_ ^ _19109_ /*66641*/;
assign _19107_ = _19108_ | _19110_ /*66638*/;
assign _19116_ = ~D[59] /*66637*/;
assign _19113_ = _18363_ & _19116_ /*66633*/;
assign _19114_ = _18363_ ^ _19116_ /*66636*/;
assign _19115_ = _19107_ & _19114_ /*66634*/;
assign _18812_ = _19107_ ^ _19114_ /*66635*/;
assign _19112_ = _19113_ | _19115_ /*66632*/;
assign _19121_ = ~D[60] /*66631*/;
assign _19118_ = _18364_ & _19121_ /*66627*/;
assign _19119_ = _18364_ ^ _19121_ /*66630*/;
assign _19120_ = _19112_ & _19119_ /*66628*/;
assign _18813_ = _19112_ ^ _19119_ /*66629*/;
assign _19117_ = _19118_ | _19120_ /*66626*/;
assign _19126_ = ~D[61] /*66625*/;
assign _19123_ = _18365_ & _19126_ /*66621*/;
assign _19124_ = _18365_ ^ _19126_ /*66624*/;
assign _19125_ = _19117_ & _19124_ /*66622*/;
assign _18814_ = _19117_ ^ _19124_ /*66623*/;
assign _19122_ = _19123_ | _19125_ /*66620*/;
assign _19131_ = ~D[62] /*66619*/;
assign _19128_ = _18366_ & _19131_ /*66615*/;
assign _19129_ = _18366_ ^ _19131_ /*66618*/;
assign _19130_ = _19122_ & _19129_ /*66616*/;
assign _18815_ = _19122_ ^ _19129_ /*66617*/;
assign _19127_ = _19128_ | _19130_ /*66614*/;
assign _19132_ = _18367_ & oneWire /*66609*/;
assign _19133_ = _18367_ ^ oneWire /*66612*/;
assign _19134_ = _19127_ & _19133_ /*66610*/;
assign _18816_ = _19127_ ^ _19133_ /*66611*/;
assign Q[42] = _19132_ | _19134_ /*66608*/;
assign _19267_ = ~Q[42] /*66223*/;
assign _19266_ = _19267_ & D[0] /*66222*/;
assign _19269_ = _18753_ & _19266_ /*66217*/;
assign _19270_ = _18753_ ^ _19266_ /*66220*/;
assign _19271_ = zeroWire & _19270_ /*66218*/;
assign _19201_ = zeroWire ^ _19270_ /*66219*/;
assign _19268_ = _19269_ | _19271_ /*66216*/;
assign _19273_ = ~Q[42] /*66215*/;
assign _19272_ = _19273_ & D[1] /*66214*/;
assign _19275_ = _18754_ & _19272_ /*66209*/;
assign _19276_ = _18754_ ^ _19272_ /*66212*/;
assign _19277_ = _19268_ & _19276_ /*66210*/;
assign _19202_ = _19268_ ^ _19276_ /*66211*/;
assign _19274_ = _19275_ | _19277_ /*66208*/;
assign _19279_ = ~Q[42] /*66207*/;
assign _19278_ = _19279_ & D[2] /*66206*/;
assign _19281_ = _18755_ & _19278_ /*66201*/;
assign _19282_ = _18755_ ^ _19278_ /*66204*/;
assign _19283_ = _19274_ & _19282_ /*66202*/;
assign _19203_ = _19274_ ^ _19282_ /*66203*/;
assign _19280_ = _19281_ | _19283_ /*66200*/;
assign _19285_ = ~Q[42] /*66199*/;
assign _19284_ = _19285_ & D[3] /*66198*/;
assign _19287_ = _18756_ & _19284_ /*66193*/;
assign _19288_ = _18756_ ^ _19284_ /*66196*/;
assign _19289_ = _19280_ & _19288_ /*66194*/;
assign _19204_ = _19280_ ^ _19288_ /*66195*/;
assign _19286_ = _19287_ | _19289_ /*66192*/;
assign _19291_ = ~Q[42] /*66191*/;
assign _19290_ = _19291_ & D[4] /*66190*/;
assign _19293_ = _18757_ & _19290_ /*66185*/;
assign _19294_ = _18757_ ^ _19290_ /*66188*/;
assign _19295_ = _19286_ & _19294_ /*66186*/;
assign _19205_ = _19286_ ^ _19294_ /*66187*/;
assign _19292_ = _19293_ | _19295_ /*66184*/;
assign _19297_ = ~Q[42] /*66183*/;
assign _19296_ = _19297_ & D[5] /*66182*/;
assign _19299_ = _18758_ & _19296_ /*66177*/;
assign _19300_ = _18758_ ^ _19296_ /*66180*/;
assign _19301_ = _19292_ & _19300_ /*66178*/;
assign _19206_ = _19292_ ^ _19300_ /*66179*/;
assign _19298_ = _19299_ | _19301_ /*66176*/;
assign _19303_ = ~Q[42] /*66175*/;
assign _19302_ = _19303_ & D[6] /*66174*/;
assign _19305_ = _18759_ & _19302_ /*66169*/;
assign _19306_ = _18759_ ^ _19302_ /*66172*/;
assign _19307_ = _19298_ & _19306_ /*66170*/;
assign _19207_ = _19298_ ^ _19306_ /*66171*/;
assign _19304_ = _19305_ | _19307_ /*66168*/;
assign _19309_ = ~Q[42] /*66167*/;
assign _19308_ = _19309_ & D[7] /*66166*/;
assign _19311_ = _18760_ & _19308_ /*66161*/;
assign _19312_ = _18760_ ^ _19308_ /*66164*/;
assign _19313_ = _19304_ & _19312_ /*66162*/;
assign _19208_ = _19304_ ^ _19312_ /*66163*/;
assign _19310_ = _19311_ | _19313_ /*66160*/;
assign _19315_ = ~Q[42] /*66159*/;
assign _19314_ = _19315_ & D[8] /*66158*/;
assign _19317_ = _18761_ & _19314_ /*66153*/;
assign _19318_ = _18761_ ^ _19314_ /*66156*/;
assign _19319_ = _19310_ & _19318_ /*66154*/;
assign _19209_ = _19310_ ^ _19318_ /*66155*/;
assign _19316_ = _19317_ | _19319_ /*66152*/;
assign _19321_ = ~Q[42] /*66151*/;
assign _19320_ = _19321_ & D[9] /*66150*/;
assign _19323_ = _18762_ & _19320_ /*66145*/;
assign _19324_ = _18762_ ^ _19320_ /*66148*/;
assign _19325_ = _19316_ & _19324_ /*66146*/;
assign _19210_ = _19316_ ^ _19324_ /*66147*/;
assign _19322_ = _19323_ | _19325_ /*66144*/;
assign _19327_ = ~Q[42] /*66143*/;
assign _19326_ = _19327_ & D[10] /*66142*/;
assign _19329_ = _18763_ & _19326_ /*66137*/;
assign _19330_ = _18763_ ^ _19326_ /*66140*/;
assign _19331_ = _19322_ & _19330_ /*66138*/;
assign _19211_ = _19322_ ^ _19330_ /*66139*/;
assign _19328_ = _19329_ | _19331_ /*66136*/;
assign _19333_ = ~Q[42] /*66135*/;
assign _19332_ = _19333_ & D[11] /*66134*/;
assign _19335_ = _18764_ & _19332_ /*66129*/;
assign _19336_ = _18764_ ^ _19332_ /*66132*/;
assign _19337_ = _19328_ & _19336_ /*66130*/;
assign _19212_ = _19328_ ^ _19336_ /*66131*/;
assign _19334_ = _19335_ | _19337_ /*66128*/;
assign _19339_ = ~Q[42] /*66127*/;
assign _19338_ = _19339_ & D[12] /*66126*/;
assign _19341_ = _18765_ & _19338_ /*66121*/;
assign _19342_ = _18765_ ^ _19338_ /*66124*/;
assign _19343_ = _19334_ & _19342_ /*66122*/;
assign _19213_ = _19334_ ^ _19342_ /*66123*/;
assign _19340_ = _19341_ | _19343_ /*66120*/;
assign _19345_ = ~Q[42] /*66119*/;
assign _19344_ = _19345_ & D[13] /*66118*/;
assign _19347_ = _18766_ & _19344_ /*66113*/;
assign _19348_ = _18766_ ^ _19344_ /*66116*/;
assign _19349_ = _19340_ & _19348_ /*66114*/;
assign _19214_ = _19340_ ^ _19348_ /*66115*/;
assign _19346_ = _19347_ | _19349_ /*66112*/;
assign _19351_ = ~Q[42] /*66111*/;
assign _19350_ = _19351_ & D[14] /*66110*/;
assign _19353_ = _18767_ & _19350_ /*66105*/;
assign _19354_ = _18767_ ^ _19350_ /*66108*/;
assign _19355_ = _19346_ & _19354_ /*66106*/;
assign _19215_ = _19346_ ^ _19354_ /*66107*/;
assign _19352_ = _19353_ | _19355_ /*66104*/;
assign _19357_ = ~Q[42] /*66103*/;
assign _19356_ = _19357_ & D[15] /*66102*/;
assign _19359_ = _18768_ & _19356_ /*66097*/;
assign _19360_ = _18768_ ^ _19356_ /*66100*/;
assign _19361_ = _19352_ & _19360_ /*66098*/;
assign _19216_ = _19352_ ^ _19360_ /*66099*/;
assign _19358_ = _19359_ | _19361_ /*66096*/;
assign _19363_ = ~Q[42] /*66095*/;
assign _19362_ = _19363_ & D[16] /*66094*/;
assign _19365_ = _18769_ & _19362_ /*66089*/;
assign _19366_ = _18769_ ^ _19362_ /*66092*/;
assign _19367_ = _19358_ & _19366_ /*66090*/;
assign _19217_ = _19358_ ^ _19366_ /*66091*/;
assign _19364_ = _19365_ | _19367_ /*66088*/;
assign _19369_ = ~Q[42] /*66087*/;
assign _19368_ = _19369_ & D[17] /*66086*/;
assign _19371_ = _18770_ & _19368_ /*66081*/;
assign _19372_ = _18770_ ^ _19368_ /*66084*/;
assign _19373_ = _19364_ & _19372_ /*66082*/;
assign _19218_ = _19364_ ^ _19372_ /*66083*/;
assign _19370_ = _19371_ | _19373_ /*66080*/;
assign _19375_ = ~Q[42] /*66079*/;
assign _19374_ = _19375_ & D[18] /*66078*/;
assign _19377_ = _18771_ & _19374_ /*66073*/;
assign _19378_ = _18771_ ^ _19374_ /*66076*/;
assign _19379_ = _19370_ & _19378_ /*66074*/;
assign _19219_ = _19370_ ^ _19378_ /*66075*/;
assign _19376_ = _19377_ | _19379_ /*66072*/;
assign _19381_ = ~Q[42] /*66071*/;
assign _19380_ = _19381_ & D[19] /*66070*/;
assign _19383_ = _18772_ & _19380_ /*66065*/;
assign _19384_ = _18772_ ^ _19380_ /*66068*/;
assign _19385_ = _19376_ & _19384_ /*66066*/;
assign _19220_ = _19376_ ^ _19384_ /*66067*/;
assign _19382_ = _19383_ | _19385_ /*66064*/;
assign _19387_ = ~Q[42] /*66063*/;
assign _19386_ = _19387_ & D[20] /*66062*/;
assign _19389_ = _18773_ & _19386_ /*66057*/;
assign _19390_ = _18773_ ^ _19386_ /*66060*/;
assign _19391_ = _19382_ & _19390_ /*66058*/;
assign _19221_ = _19382_ ^ _19390_ /*66059*/;
assign _19388_ = _19389_ | _19391_ /*66056*/;
assign _19393_ = ~Q[42] /*66055*/;
assign _19392_ = _19393_ & D[21] /*66054*/;
assign _19395_ = _18774_ & _19392_ /*66049*/;
assign _19396_ = _18774_ ^ _19392_ /*66052*/;
assign _19397_ = _19388_ & _19396_ /*66050*/;
assign _19222_ = _19388_ ^ _19396_ /*66051*/;
assign _19394_ = _19395_ | _19397_ /*66048*/;
assign _19399_ = ~Q[42] /*66047*/;
assign _19398_ = _19399_ & D[22] /*66046*/;
assign _19401_ = _18775_ & _19398_ /*66041*/;
assign _19402_ = _18775_ ^ _19398_ /*66044*/;
assign _19403_ = _19394_ & _19402_ /*66042*/;
assign _19223_ = _19394_ ^ _19402_ /*66043*/;
assign _19400_ = _19401_ | _19403_ /*66040*/;
assign _19405_ = ~Q[42] /*66039*/;
assign _19404_ = _19405_ & D[23] /*66038*/;
assign _19407_ = _18776_ & _19404_ /*66033*/;
assign _19408_ = _18776_ ^ _19404_ /*66036*/;
assign _19409_ = _19400_ & _19408_ /*66034*/;
assign _19224_ = _19400_ ^ _19408_ /*66035*/;
assign _19406_ = _19407_ | _19409_ /*66032*/;
assign _19411_ = ~Q[42] /*66031*/;
assign _19410_ = _19411_ & D[24] /*66030*/;
assign _19413_ = _18777_ & _19410_ /*66025*/;
assign _19414_ = _18777_ ^ _19410_ /*66028*/;
assign _19415_ = _19406_ & _19414_ /*66026*/;
assign _19225_ = _19406_ ^ _19414_ /*66027*/;
assign _19412_ = _19413_ | _19415_ /*66024*/;
assign _19417_ = ~Q[42] /*66023*/;
assign _19416_ = _19417_ & D[25] /*66022*/;
assign _19419_ = _18778_ & _19416_ /*66017*/;
assign _19420_ = _18778_ ^ _19416_ /*66020*/;
assign _19421_ = _19412_ & _19420_ /*66018*/;
assign _19226_ = _19412_ ^ _19420_ /*66019*/;
assign _19418_ = _19419_ | _19421_ /*66016*/;
assign _19423_ = ~Q[42] /*66015*/;
assign _19422_ = _19423_ & D[26] /*66014*/;
assign _19425_ = _18779_ & _19422_ /*66009*/;
assign _19426_ = _18779_ ^ _19422_ /*66012*/;
assign _19427_ = _19418_ & _19426_ /*66010*/;
assign _19227_ = _19418_ ^ _19426_ /*66011*/;
assign _19424_ = _19425_ | _19427_ /*66008*/;
assign _19429_ = ~Q[42] /*66007*/;
assign _19428_ = _19429_ & D[27] /*66006*/;
assign _19431_ = _18780_ & _19428_ /*66001*/;
assign _19432_ = _18780_ ^ _19428_ /*66004*/;
assign _19433_ = _19424_ & _19432_ /*66002*/;
assign _19228_ = _19424_ ^ _19432_ /*66003*/;
assign _19430_ = _19431_ | _19433_ /*66000*/;
assign _19435_ = ~Q[42] /*65999*/;
assign _19434_ = _19435_ & D[28] /*65998*/;
assign _19437_ = _18781_ & _19434_ /*65993*/;
assign _19438_ = _18781_ ^ _19434_ /*65996*/;
assign _19439_ = _19430_ & _19438_ /*65994*/;
assign _19229_ = _19430_ ^ _19438_ /*65995*/;
assign _19436_ = _19437_ | _19439_ /*65992*/;
assign _19441_ = ~Q[42] /*65991*/;
assign _19440_ = _19441_ & D[29] /*65990*/;
assign _19443_ = _18782_ & _19440_ /*65985*/;
assign _19444_ = _18782_ ^ _19440_ /*65988*/;
assign _19445_ = _19436_ & _19444_ /*65986*/;
assign _19230_ = _19436_ ^ _19444_ /*65987*/;
assign _19442_ = _19443_ | _19445_ /*65984*/;
assign _19447_ = ~Q[42] /*65983*/;
assign _19446_ = _19447_ & D[30] /*65982*/;
assign _19449_ = _18783_ & _19446_ /*65977*/;
assign _19450_ = _18783_ ^ _19446_ /*65980*/;
assign _19451_ = _19442_ & _19450_ /*65978*/;
assign _19231_ = _19442_ ^ _19450_ /*65979*/;
assign _19448_ = _19449_ | _19451_ /*65976*/;
assign _19453_ = ~Q[42] /*65975*/;
assign _19452_ = _19453_ & D[31] /*65974*/;
assign _19455_ = _18784_ & _19452_ /*65969*/;
assign _19456_ = _18784_ ^ _19452_ /*65972*/;
assign _19457_ = _19448_ & _19456_ /*65970*/;
assign _19232_ = _19448_ ^ _19456_ /*65971*/;
assign _19454_ = _19455_ | _19457_ /*65968*/;
assign _19459_ = ~Q[42] /*65967*/;
assign _19458_ = _19459_ & D[32] /*65966*/;
assign _19461_ = _18785_ & _19458_ /*65961*/;
assign _19462_ = _18785_ ^ _19458_ /*65964*/;
assign _19463_ = _19454_ & _19462_ /*65962*/;
assign _19233_ = _19454_ ^ _19462_ /*65963*/;
assign _19460_ = _19461_ | _19463_ /*65960*/;
assign _19465_ = ~Q[42] /*65959*/;
assign _19464_ = _19465_ & D[33] /*65958*/;
assign _19467_ = _18786_ & _19464_ /*65953*/;
assign _19468_ = _18786_ ^ _19464_ /*65956*/;
assign _19469_ = _19460_ & _19468_ /*65954*/;
assign _19234_ = _19460_ ^ _19468_ /*65955*/;
assign _19466_ = _19467_ | _19469_ /*65952*/;
assign _19471_ = ~Q[42] /*65951*/;
assign _19470_ = _19471_ & D[34] /*65950*/;
assign _19473_ = _18787_ & _19470_ /*65945*/;
assign _19474_ = _18787_ ^ _19470_ /*65948*/;
assign _19475_ = _19466_ & _19474_ /*65946*/;
assign _19235_ = _19466_ ^ _19474_ /*65947*/;
assign _19472_ = _19473_ | _19475_ /*65944*/;
assign _19477_ = ~Q[42] /*65943*/;
assign _19476_ = _19477_ & D[35] /*65942*/;
assign _19479_ = _18788_ & _19476_ /*65937*/;
assign _19480_ = _18788_ ^ _19476_ /*65940*/;
assign _19481_ = _19472_ & _19480_ /*65938*/;
assign _19236_ = _19472_ ^ _19480_ /*65939*/;
assign _19478_ = _19479_ | _19481_ /*65936*/;
assign _19483_ = ~Q[42] /*65935*/;
assign _19482_ = _19483_ & D[36] /*65934*/;
assign _19485_ = _18789_ & _19482_ /*65929*/;
assign _19486_ = _18789_ ^ _19482_ /*65932*/;
assign _19487_ = _19478_ & _19486_ /*65930*/;
assign _19237_ = _19478_ ^ _19486_ /*65931*/;
assign _19484_ = _19485_ | _19487_ /*65928*/;
assign _19489_ = ~Q[42] /*65927*/;
assign _19488_ = _19489_ & D[37] /*65926*/;
assign _19491_ = _18790_ & _19488_ /*65921*/;
assign _19492_ = _18790_ ^ _19488_ /*65924*/;
assign _19493_ = _19484_ & _19492_ /*65922*/;
assign _19238_ = _19484_ ^ _19492_ /*65923*/;
assign _19490_ = _19491_ | _19493_ /*65920*/;
assign _19495_ = ~Q[42] /*65919*/;
assign _19494_ = _19495_ & D[38] /*65918*/;
assign _19497_ = _18791_ & _19494_ /*65913*/;
assign _19498_ = _18791_ ^ _19494_ /*65916*/;
assign _19499_ = _19490_ & _19498_ /*65914*/;
assign _19239_ = _19490_ ^ _19498_ /*65915*/;
assign _19496_ = _19497_ | _19499_ /*65912*/;
assign _19501_ = ~Q[42] /*65911*/;
assign _19500_ = _19501_ & D[39] /*65910*/;
assign _19503_ = _18792_ & _19500_ /*65905*/;
assign _19504_ = _18792_ ^ _19500_ /*65908*/;
assign _19505_ = _19496_ & _19504_ /*65906*/;
assign _19240_ = _19496_ ^ _19504_ /*65907*/;
assign _19502_ = _19503_ | _19505_ /*65904*/;
assign _19507_ = ~Q[42] /*65903*/;
assign _19506_ = _19507_ & D[40] /*65902*/;
assign _19509_ = _18793_ & _19506_ /*65897*/;
assign _19510_ = _18793_ ^ _19506_ /*65900*/;
assign _19511_ = _19502_ & _19510_ /*65898*/;
assign _19241_ = _19502_ ^ _19510_ /*65899*/;
assign _19508_ = _19509_ | _19511_ /*65896*/;
assign _19513_ = ~Q[42] /*65895*/;
assign _19512_ = _19513_ & D[41] /*65894*/;
assign _19515_ = _18794_ & _19512_ /*65889*/;
assign _19516_ = _18794_ ^ _19512_ /*65892*/;
assign _19517_ = _19508_ & _19516_ /*65890*/;
assign _19242_ = _19508_ ^ _19516_ /*65891*/;
assign _19514_ = _19515_ | _19517_ /*65888*/;
assign _19519_ = ~Q[42] /*65887*/;
assign _19518_ = _19519_ & D[42] /*65886*/;
assign _19521_ = _18795_ & _19518_ /*65881*/;
assign _19522_ = _18795_ ^ _19518_ /*65884*/;
assign _19523_ = _19514_ & _19522_ /*65882*/;
assign _19243_ = _19514_ ^ _19522_ /*65883*/;
assign _19520_ = _19521_ | _19523_ /*65880*/;
assign _19525_ = ~Q[42] /*65879*/;
assign _19524_ = _19525_ & D[43] /*65878*/;
assign _19527_ = _18796_ & _19524_ /*65873*/;
assign _19528_ = _18796_ ^ _19524_ /*65876*/;
assign _19529_ = _19520_ & _19528_ /*65874*/;
assign _19244_ = _19520_ ^ _19528_ /*65875*/;
assign _19526_ = _19527_ | _19529_ /*65872*/;
assign _19531_ = ~Q[42] /*65871*/;
assign _19530_ = _19531_ & D[44] /*65870*/;
assign _19533_ = _18797_ & _19530_ /*65865*/;
assign _19534_ = _18797_ ^ _19530_ /*65868*/;
assign _19535_ = _19526_ & _19534_ /*65866*/;
assign _19245_ = _19526_ ^ _19534_ /*65867*/;
assign _19532_ = _19533_ | _19535_ /*65864*/;
assign _19537_ = ~Q[42] /*65863*/;
assign _19536_ = _19537_ & D[45] /*65862*/;
assign _19539_ = _18798_ & _19536_ /*65857*/;
assign _19540_ = _18798_ ^ _19536_ /*65860*/;
assign _19541_ = _19532_ & _19540_ /*65858*/;
assign _19246_ = _19532_ ^ _19540_ /*65859*/;
assign _19538_ = _19539_ | _19541_ /*65856*/;
assign _19543_ = ~Q[42] /*65855*/;
assign _19542_ = _19543_ & D[46] /*65854*/;
assign _19545_ = _18799_ & _19542_ /*65849*/;
assign _19546_ = _18799_ ^ _19542_ /*65852*/;
assign _19547_ = _19538_ & _19546_ /*65850*/;
assign _19247_ = _19538_ ^ _19546_ /*65851*/;
assign _19544_ = _19545_ | _19547_ /*65848*/;
assign _19549_ = ~Q[42] /*65847*/;
assign _19548_ = _19549_ & D[47] /*65846*/;
assign _19551_ = _18800_ & _19548_ /*65841*/;
assign _19552_ = _18800_ ^ _19548_ /*65844*/;
assign _19553_ = _19544_ & _19552_ /*65842*/;
assign _19248_ = _19544_ ^ _19552_ /*65843*/;
assign _19550_ = _19551_ | _19553_ /*65840*/;
assign _19555_ = ~Q[42] /*65839*/;
assign _19554_ = _19555_ & D[48] /*65838*/;
assign _19557_ = _18801_ & _19554_ /*65833*/;
assign _19558_ = _18801_ ^ _19554_ /*65836*/;
assign _19559_ = _19550_ & _19558_ /*65834*/;
assign _19249_ = _19550_ ^ _19558_ /*65835*/;
assign _19556_ = _19557_ | _19559_ /*65832*/;
assign _19561_ = ~Q[42] /*65831*/;
assign _19560_ = _19561_ & D[49] /*65830*/;
assign _19563_ = _18802_ & _19560_ /*65825*/;
assign _19564_ = _18802_ ^ _19560_ /*65828*/;
assign _19565_ = _19556_ & _19564_ /*65826*/;
assign _19250_ = _19556_ ^ _19564_ /*65827*/;
assign _19562_ = _19563_ | _19565_ /*65824*/;
assign _19567_ = ~Q[42] /*65823*/;
assign _19566_ = _19567_ & D[50] /*65822*/;
assign _19569_ = _18803_ & _19566_ /*65817*/;
assign _19570_ = _18803_ ^ _19566_ /*65820*/;
assign _19571_ = _19562_ & _19570_ /*65818*/;
assign _19251_ = _19562_ ^ _19570_ /*65819*/;
assign _19568_ = _19569_ | _19571_ /*65816*/;
assign _19573_ = ~Q[42] /*65815*/;
assign _19572_ = _19573_ & D[51] /*65814*/;
assign _19575_ = _18804_ & _19572_ /*65809*/;
assign _19576_ = _18804_ ^ _19572_ /*65812*/;
assign _19577_ = _19568_ & _19576_ /*65810*/;
assign _19252_ = _19568_ ^ _19576_ /*65811*/;
assign _19574_ = _19575_ | _19577_ /*65808*/;
assign _19579_ = ~Q[42] /*65807*/;
assign _19578_ = _19579_ & D[52] /*65806*/;
assign _19581_ = _18805_ & _19578_ /*65801*/;
assign _19582_ = _18805_ ^ _19578_ /*65804*/;
assign _19583_ = _19574_ & _19582_ /*65802*/;
assign _19253_ = _19574_ ^ _19582_ /*65803*/;
assign _19580_ = _19581_ | _19583_ /*65800*/;
assign _19585_ = ~Q[42] /*65799*/;
assign _19584_ = _19585_ & D[53] /*65798*/;
assign _19587_ = _18806_ & _19584_ /*65793*/;
assign _19588_ = _18806_ ^ _19584_ /*65796*/;
assign _19589_ = _19580_ & _19588_ /*65794*/;
assign _19254_ = _19580_ ^ _19588_ /*65795*/;
assign _19586_ = _19587_ | _19589_ /*65792*/;
assign _19591_ = ~Q[42] /*65791*/;
assign _19590_ = _19591_ & D[54] /*65790*/;
assign _19593_ = _18807_ & _19590_ /*65785*/;
assign _19594_ = _18807_ ^ _19590_ /*65788*/;
assign _19595_ = _19586_ & _19594_ /*65786*/;
assign _19255_ = _19586_ ^ _19594_ /*65787*/;
assign _19592_ = _19593_ | _19595_ /*65784*/;
assign _19597_ = ~Q[42] /*65783*/;
assign _19596_ = _19597_ & D[55] /*65782*/;
assign _19599_ = _18808_ & _19596_ /*65777*/;
assign _19600_ = _18808_ ^ _19596_ /*65780*/;
assign _19601_ = _19592_ & _19600_ /*65778*/;
assign _19256_ = _19592_ ^ _19600_ /*65779*/;
assign _19598_ = _19599_ | _19601_ /*65776*/;
assign _19603_ = ~Q[42] /*65775*/;
assign _19602_ = _19603_ & D[56] /*65774*/;
assign _19605_ = _18809_ & _19602_ /*65769*/;
assign _19606_ = _18809_ ^ _19602_ /*65772*/;
assign _19607_ = _19598_ & _19606_ /*65770*/;
assign _19257_ = _19598_ ^ _19606_ /*65771*/;
assign _19604_ = _19605_ | _19607_ /*65768*/;
assign _19609_ = ~Q[42] /*65767*/;
assign _19608_ = _19609_ & D[57] /*65766*/;
assign _19611_ = _18810_ & _19608_ /*65761*/;
assign _19612_ = _18810_ ^ _19608_ /*65764*/;
assign _19613_ = _19604_ & _19612_ /*65762*/;
assign _19258_ = _19604_ ^ _19612_ /*65763*/;
assign _19610_ = _19611_ | _19613_ /*65760*/;
assign _19615_ = ~Q[42] /*65759*/;
assign _19614_ = _19615_ & D[58] /*65758*/;
assign _19617_ = _18811_ & _19614_ /*65753*/;
assign _19618_ = _18811_ ^ _19614_ /*65756*/;
assign _19619_ = _19610_ & _19618_ /*65754*/;
assign _19259_ = _19610_ ^ _19618_ /*65755*/;
assign _19616_ = _19617_ | _19619_ /*65752*/;
assign _19621_ = ~Q[42] /*65751*/;
assign _19620_ = _19621_ & D[59] /*65750*/;
assign _19623_ = _18812_ & _19620_ /*65745*/;
assign _19624_ = _18812_ ^ _19620_ /*65748*/;
assign _19625_ = _19616_ & _19624_ /*65746*/;
assign _19260_ = _19616_ ^ _19624_ /*65747*/;
assign _19622_ = _19623_ | _19625_ /*65744*/;
assign _19627_ = ~Q[42] /*65743*/;
assign _19626_ = _19627_ & D[60] /*65742*/;
assign _19629_ = _18813_ & _19626_ /*65737*/;
assign _19630_ = _18813_ ^ _19626_ /*65740*/;
assign _19631_ = _19622_ & _19630_ /*65738*/;
assign _19261_ = _19622_ ^ _19630_ /*65739*/;
assign _19628_ = _19629_ | _19631_ /*65736*/;
assign _19633_ = ~Q[42] /*65735*/;
assign _19632_ = _19633_ & D[61] /*65734*/;
assign _19635_ = _18814_ & _19632_ /*65729*/;
assign _19636_ = _18814_ ^ _19632_ /*65732*/;
assign _19637_ = _19628_ & _19636_ /*65730*/;
assign _19262_ = _19628_ ^ _19636_ /*65731*/;
assign _19634_ = _19635_ | _19637_ /*65728*/;
assign _19639_ = ~Q[42] /*65727*/;
assign _19638_ = _19639_ & D[62] /*65726*/;
assign _19641_ = _18815_ & _19638_ /*65721*/;
assign _19642_ = _18815_ ^ _19638_ /*65724*/;
assign _19643_ = _19634_ & _19642_ /*65722*/;
assign _19263_ = _19634_ ^ _19642_ /*65723*/;
assign _19640_ = _19641_ | _19643_ /*65720*/;
assign _19645_ = ~Q[42] /*65719*/;
assign _19644_ = _19645_ & zeroWire /*65718*/;
assign _19646_ = _18816_ ^ _19644_ /*65716*/;
assign _19264_ = _19646_ ^ _19640_ /*65715*/;
assign _19717_ = ~D[0] /*65461*/;
assign _19714_ = R_0[41] & _19717_ /*65457*/;
assign _19715_ = R_0[41] ^ _19717_ /*65460*/;
assign _19716_ = oneWire & _19715_ /*65458*/;
assign _19649_ = oneWire ^ _19715_ /*65459*/;
assign _19713_ = _19714_ | _19716_ /*65456*/;
assign _19722_ = ~D[1] /*65455*/;
assign _19719_ = _19201_ & _19722_ /*65451*/;
assign _19720_ = _19201_ ^ _19722_ /*65454*/;
assign _19721_ = _19713_ & _19720_ /*65452*/;
assign _19650_ = _19713_ ^ _19720_ /*65453*/;
assign _19718_ = _19719_ | _19721_ /*65450*/;
assign _19727_ = ~D[2] /*65449*/;
assign _19724_ = _19202_ & _19727_ /*65445*/;
assign _19725_ = _19202_ ^ _19727_ /*65448*/;
assign _19726_ = _19718_ & _19725_ /*65446*/;
assign _19651_ = _19718_ ^ _19725_ /*65447*/;
assign _19723_ = _19724_ | _19726_ /*65444*/;
assign _19732_ = ~D[3] /*65443*/;
assign _19729_ = _19203_ & _19732_ /*65439*/;
assign _19730_ = _19203_ ^ _19732_ /*65442*/;
assign _19731_ = _19723_ & _19730_ /*65440*/;
assign _19652_ = _19723_ ^ _19730_ /*65441*/;
assign _19728_ = _19729_ | _19731_ /*65438*/;
assign _19737_ = ~D[4] /*65437*/;
assign _19734_ = _19204_ & _19737_ /*65433*/;
assign _19735_ = _19204_ ^ _19737_ /*65436*/;
assign _19736_ = _19728_ & _19735_ /*65434*/;
assign _19653_ = _19728_ ^ _19735_ /*65435*/;
assign _19733_ = _19734_ | _19736_ /*65432*/;
assign _19742_ = ~D[5] /*65431*/;
assign _19739_ = _19205_ & _19742_ /*65427*/;
assign _19740_ = _19205_ ^ _19742_ /*65430*/;
assign _19741_ = _19733_ & _19740_ /*65428*/;
assign _19654_ = _19733_ ^ _19740_ /*65429*/;
assign _19738_ = _19739_ | _19741_ /*65426*/;
assign _19747_ = ~D[6] /*65425*/;
assign _19744_ = _19206_ & _19747_ /*65421*/;
assign _19745_ = _19206_ ^ _19747_ /*65424*/;
assign _19746_ = _19738_ & _19745_ /*65422*/;
assign _19655_ = _19738_ ^ _19745_ /*65423*/;
assign _19743_ = _19744_ | _19746_ /*65420*/;
assign _19752_ = ~D[7] /*65419*/;
assign _19749_ = _19207_ & _19752_ /*65415*/;
assign _19750_ = _19207_ ^ _19752_ /*65418*/;
assign _19751_ = _19743_ & _19750_ /*65416*/;
assign _19656_ = _19743_ ^ _19750_ /*65417*/;
assign _19748_ = _19749_ | _19751_ /*65414*/;
assign _19757_ = ~D[8] /*65413*/;
assign _19754_ = _19208_ & _19757_ /*65409*/;
assign _19755_ = _19208_ ^ _19757_ /*65412*/;
assign _19756_ = _19748_ & _19755_ /*65410*/;
assign _19657_ = _19748_ ^ _19755_ /*65411*/;
assign _19753_ = _19754_ | _19756_ /*65408*/;
assign _19762_ = ~D[9] /*65407*/;
assign _19759_ = _19209_ & _19762_ /*65403*/;
assign _19760_ = _19209_ ^ _19762_ /*65406*/;
assign _19761_ = _19753_ & _19760_ /*65404*/;
assign _19658_ = _19753_ ^ _19760_ /*65405*/;
assign _19758_ = _19759_ | _19761_ /*65402*/;
assign _19767_ = ~D[10] /*65401*/;
assign _19764_ = _19210_ & _19767_ /*65397*/;
assign _19765_ = _19210_ ^ _19767_ /*65400*/;
assign _19766_ = _19758_ & _19765_ /*65398*/;
assign _19659_ = _19758_ ^ _19765_ /*65399*/;
assign _19763_ = _19764_ | _19766_ /*65396*/;
assign _19772_ = ~D[11] /*65395*/;
assign _19769_ = _19211_ & _19772_ /*65391*/;
assign _19770_ = _19211_ ^ _19772_ /*65394*/;
assign _19771_ = _19763_ & _19770_ /*65392*/;
assign _19660_ = _19763_ ^ _19770_ /*65393*/;
assign _19768_ = _19769_ | _19771_ /*65390*/;
assign _19777_ = ~D[12] /*65389*/;
assign _19774_ = _19212_ & _19777_ /*65385*/;
assign _19775_ = _19212_ ^ _19777_ /*65388*/;
assign _19776_ = _19768_ & _19775_ /*65386*/;
assign _19661_ = _19768_ ^ _19775_ /*65387*/;
assign _19773_ = _19774_ | _19776_ /*65384*/;
assign _19782_ = ~D[13] /*65383*/;
assign _19779_ = _19213_ & _19782_ /*65379*/;
assign _19780_ = _19213_ ^ _19782_ /*65382*/;
assign _19781_ = _19773_ & _19780_ /*65380*/;
assign _19662_ = _19773_ ^ _19780_ /*65381*/;
assign _19778_ = _19779_ | _19781_ /*65378*/;
assign _19787_ = ~D[14] /*65377*/;
assign _19784_ = _19214_ & _19787_ /*65373*/;
assign _19785_ = _19214_ ^ _19787_ /*65376*/;
assign _19786_ = _19778_ & _19785_ /*65374*/;
assign _19663_ = _19778_ ^ _19785_ /*65375*/;
assign _19783_ = _19784_ | _19786_ /*65372*/;
assign _19792_ = ~D[15] /*65371*/;
assign _19789_ = _19215_ & _19792_ /*65367*/;
assign _19790_ = _19215_ ^ _19792_ /*65370*/;
assign _19791_ = _19783_ & _19790_ /*65368*/;
assign _19664_ = _19783_ ^ _19790_ /*65369*/;
assign _19788_ = _19789_ | _19791_ /*65366*/;
assign _19797_ = ~D[16] /*65365*/;
assign _19794_ = _19216_ & _19797_ /*65361*/;
assign _19795_ = _19216_ ^ _19797_ /*65364*/;
assign _19796_ = _19788_ & _19795_ /*65362*/;
assign _19665_ = _19788_ ^ _19795_ /*65363*/;
assign _19793_ = _19794_ | _19796_ /*65360*/;
assign _19802_ = ~D[17] /*65359*/;
assign _19799_ = _19217_ & _19802_ /*65355*/;
assign _19800_ = _19217_ ^ _19802_ /*65358*/;
assign _19801_ = _19793_ & _19800_ /*65356*/;
assign _19666_ = _19793_ ^ _19800_ /*65357*/;
assign _19798_ = _19799_ | _19801_ /*65354*/;
assign _19807_ = ~D[18] /*65353*/;
assign _19804_ = _19218_ & _19807_ /*65349*/;
assign _19805_ = _19218_ ^ _19807_ /*65352*/;
assign _19806_ = _19798_ & _19805_ /*65350*/;
assign _19667_ = _19798_ ^ _19805_ /*65351*/;
assign _19803_ = _19804_ | _19806_ /*65348*/;
assign _19812_ = ~D[19] /*65347*/;
assign _19809_ = _19219_ & _19812_ /*65343*/;
assign _19810_ = _19219_ ^ _19812_ /*65346*/;
assign _19811_ = _19803_ & _19810_ /*65344*/;
assign _19668_ = _19803_ ^ _19810_ /*65345*/;
assign _19808_ = _19809_ | _19811_ /*65342*/;
assign _19817_ = ~D[20] /*65341*/;
assign _19814_ = _19220_ & _19817_ /*65337*/;
assign _19815_ = _19220_ ^ _19817_ /*65340*/;
assign _19816_ = _19808_ & _19815_ /*65338*/;
assign _19669_ = _19808_ ^ _19815_ /*65339*/;
assign _19813_ = _19814_ | _19816_ /*65336*/;
assign _19822_ = ~D[21] /*65335*/;
assign _19819_ = _19221_ & _19822_ /*65331*/;
assign _19820_ = _19221_ ^ _19822_ /*65334*/;
assign _19821_ = _19813_ & _19820_ /*65332*/;
assign _19670_ = _19813_ ^ _19820_ /*65333*/;
assign _19818_ = _19819_ | _19821_ /*65330*/;
assign _19827_ = ~D[22] /*65329*/;
assign _19824_ = _19222_ & _19827_ /*65325*/;
assign _19825_ = _19222_ ^ _19827_ /*65328*/;
assign _19826_ = _19818_ & _19825_ /*65326*/;
assign _19671_ = _19818_ ^ _19825_ /*65327*/;
assign _19823_ = _19824_ | _19826_ /*65324*/;
assign _19832_ = ~D[23] /*65323*/;
assign _19829_ = _19223_ & _19832_ /*65319*/;
assign _19830_ = _19223_ ^ _19832_ /*65322*/;
assign _19831_ = _19823_ & _19830_ /*65320*/;
assign _19672_ = _19823_ ^ _19830_ /*65321*/;
assign _19828_ = _19829_ | _19831_ /*65318*/;
assign _19837_ = ~D[24] /*65317*/;
assign _19834_ = _19224_ & _19837_ /*65313*/;
assign _19835_ = _19224_ ^ _19837_ /*65316*/;
assign _19836_ = _19828_ & _19835_ /*65314*/;
assign _19673_ = _19828_ ^ _19835_ /*65315*/;
assign _19833_ = _19834_ | _19836_ /*65312*/;
assign _19842_ = ~D[25] /*65311*/;
assign _19839_ = _19225_ & _19842_ /*65307*/;
assign _19840_ = _19225_ ^ _19842_ /*65310*/;
assign _19841_ = _19833_ & _19840_ /*65308*/;
assign _19674_ = _19833_ ^ _19840_ /*65309*/;
assign _19838_ = _19839_ | _19841_ /*65306*/;
assign _19847_ = ~D[26] /*65305*/;
assign _19844_ = _19226_ & _19847_ /*65301*/;
assign _19845_ = _19226_ ^ _19847_ /*65304*/;
assign _19846_ = _19838_ & _19845_ /*65302*/;
assign _19675_ = _19838_ ^ _19845_ /*65303*/;
assign _19843_ = _19844_ | _19846_ /*65300*/;
assign _19852_ = ~D[27] /*65299*/;
assign _19849_ = _19227_ & _19852_ /*65295*/;
assign _19850_ = _19227_ ^ _19852_ /*65298*/;
assign _19851_ = _19843_ & _19850_ /*65296*/;
assign _19676_ = _19843_ ^ _19850_ /*65297*/;
assign _19848_ = _19849_ | _19851_ /*65294*/;
assign _19857_ = ~D[28] /*65293*/;
assign _19854_ = _19228_ & _19857_ /*65289*/;
assign _19855_ = _19228_ ^ _19857_ /*65292*/;
assign _19856_ = _19848_ & _19855_ /*65290*/;
assign _19677_ = _19848_ ^ _19855_ /*65291*/;
assign _19853_ = _19854_ | _19856_ /*65288*/;
assign _19862_ = ~D[29] /*65287*/;
assign _19859_ = _19229_ & _19862_ /*65283*/;
assign _19860_ = _19229_ ^ _19862_ /*65286*/;
assign _19861_ = _19853_ & _19860_ /*65284*/;
assign _19678_ = _19853_ ^ _19860_ /*65285*/;
assign _19858_ = _19859_ | _19861_ /*65282*/;
assign _19867_ = ~D[30] /*65281*/;
assign _19864_ = _19230_ & _19867_ /*65277*/;
assign _19865_ = _19230_ ^ _19867_ /*65280*/;
assign _19866_ = _19858_ & _19865_ /*65278*/;
assign _19679_ = _19858_ ^ _19865_ /*65279*/;
assign _19863_ = _19864_ | _19866_ /*65276*/;
assign _19872_ = ~D[31] /*65275*/;
assign _19869_ = _19231_ & _19872_ /*65271*/;
assign _19870_ = _19231_ ^ _19872_ /*65274*/;
assign _19871_ = _19863_ & _19870_ /*65272*/;
assign _19680_ = _19863_ ^ _19870_ /*65273*/;
assign _19868_ = _19869_ | _19871_ /*65270*/;
assign _19877_ = ~D[32] /*65269*/;
assign _19874_ = _19232_ & _19877_ /*65265*/;
assign _19875_ = _19232_ ^ _19877_ /*65268*/;
assign _19876_ = _19868_ & _19875_ /*65266*/;
assign _19681_ = _19868_ ^ _19875_ /*65267*/;
assign _19873_ = _19874_ | _19876_ /*65264*/;
assign _19882_ = ~D[33] /*65263*/;
assign _19879_ = _19233_ & _19882_ /*65259*/;
assign _19880_ = _19233_ ^ _19882_ /*65262*/;
assign _19881_ = _19873_ & _19880_ /*65260*/;
assign _19682_ = _19873_ ^ _19880_ /*65261*/;
assign _19878_ = _19879_ | _19881_ /*65258*/;
assign _19887_ = ~D[34] /*65257*/;
assign _19884_ = _19234_ & _19887_ /*65253*/;
assign _19885_ = _19234_ ^ _19887_ /*65256*/;
assign _19886_ = _19878_ & _19885_ /*65254*/;
assign _19683_ = _19878_ ^ _19885_ /*65255*/;
assign _19883_ = _19884_ | _19886_ /*65252*/;
assign _19892_ = ~D[35] /*65251*/;
assign _19889_ = _19235_ & _19892_ /*65247*/;
assign _19890_ = _19235_ ^ _19892_ /*65250*/;
assign _19891_ = _19883_ & _19890_ /*65248*/;
assign _19684_ = _19883_ ^ _19890_ /*65249*/;
assign _19888_ = _19889_ | _19891_ /*65246*/;
assign _19897_ = ~D[36] /*65245*/;
assign _19894_ = _19236_ & _19897_ /*65241*/;
assign _19895_ = _19236_ ^ _19897_ /*65244*/;
assign _19896_ = _19888_ & _19895_ /*65242*/;
assign _19685_ = _19888_ ^ _19895_ /*65243*/;
assign _19893_ = _19894_ | _19896_ /*65240*/;
assign _19902_ = ~D[37] /*65239*/;
assign _19899_ = _19237_ & _19902_ /*65235*/;
assign _19900_ = _19237_ ^ _19902_ /*65238*/;
assign _19901_ = _19893_ & _19900_ /*65236*/;
assign _19686_ = _19893_ ^ _19900_ /*65237*/;
assign _19898_ = _19899_ | _19901_ /*65234*/;
assign _19907_ = ~D[38] /*65233*/;
assign _19904_ = _19238_ & _19907_ /*65229*/;
assign _19905_ = _19238_ ^ _19907_ /*65232*/;
assign _19906_ = _19898_ & _19905_ /*65230*/;
assign _19687_ = _19898_ ^ _19905_ /*65231*/;
assign _19903_ = _19904_ | _19906_ /*65228*/;
assign _19912_ = ~D[39] /*65227*/;
assign _19909_ = _19239_ & _19912_ /*65223*/;
assign _19910_ = _19239_ ^ _19912_ /*65226*/;
assign _19911_ = _19903_ & _19910_ /*65224*/;
assign _19688_ = _19903_ ^ _19910_ /*65225*/;
assign _19908_ = _19909_ | _19911_ /*65222*/;
assign _19917_ = ~D[40] /*65221*/;
assign _19914_ = _19240_ & _19917_ /*65217*/;
assign _19915_ = _19240_ ^ _19917_ /*65220*/;
assign _19916_ = _19908_ & _19915_ /*65218*/;
assign _19689_ = _19908_ ^ _19915_ /*65219*/;
assign _19913_ = _19914_ | _19916_ /*65216*/;
assign _19922_ = ~D[41] /*65215*/;
assign _19919_ = _19241_ & _19922_ /*65211*/;
assign _19920_ = _19241_ ^ _19922_ /*65214*/;
assign _19921_ = _19913_ & _19920_ /*65212*/;
assign _19690_ = _19913_ ^ _19920_ /*65213*/;
assign _19918_ = _19919_ | _19921_ /*65210*/;
assign _19927_ = ~D[42] /*65209*/;
assign _19924_ = _19242_ & _19927_ /*65205*/;
assign _19925_ = _19242_ ^ _19927_ /*65208*/;
assign _19926_ = _19918_ & _19925_ /*65206*/;
assign _19691_ = _19918_ ^ _19925_ /*65207*/;
assign _19923_ = _19924_ | _19926_ /*65204*/;
assign _19932_ = ~D[43] /*65203*/;
assign _19929_ = _19243_ & _19932_ /*65199*/;
assign _19930_ = _19243_ ^ _19932_ /*65202*/;
assign _19931_ = _19923_ & _19930_ /*65200*/;
assign _19692_ = _19923_ ^ _19930_ /*65201*/;
assign _19928_ = _19929_ | _19931_ /*65198*/;
assign _19937_ = ~D[44] /*65197*/;
assign _19934_ = _19244_ & _19937_ /*65193*/;
assign _19935_ = _19244_ ^ _19937_ /*65196*/;
assign _19936_ = _19928_ & _19935_ /*65194*/;
assign _19693_ = _19928_ ^ _19935_ /*65195*/;
assign _19933_ = _19934_ | _19936_ /*65192*/;
assign _19942_ = ~D[45] /*65191*/;
assign _19939_ = _19245_ & _19942_ /*65187*/;
assign _19940_ = _19245_ ^ _19942_ /*65190*/;
assign _19941_ = _19933_ & _19940_ /*65188*/;
assign _19694_ = _19933_ ^ _19940_ /*65189*/;
assign _19938_ = _19939_ | _19941_ /*65186*/;
assign _19947_ = ~D[46] /*65185*/;
assign _19944_ = _19246_ & _19947_ /*65181*/;
assign _19945_ = _19246_ ^ _19947_ /*65184*/;
assign _19946_ = _19938_ & _19945_ /*65182*/;
assign _19695_ = _19938_ ^ _19945_ /*65183*/;
assign _19943_ = _19944_ | _19946_ /*65180*/;
assign _19952_ = ~D[47] /*65179*/;
assign _19949_ = _19247_ & _19952_ /*65175*/;
assign _19950_ = _19247_ ^ _19952_ /*65178*/;
assign _19951_ = _19943_ & _19950_ /*65176*/;
assign _19696_ = _19943_ ^ _19950_ /*65177*/;
assign _19948_ = _19949_ | _19951_ /*65174*/;
assign _19957_ = ~D[48] /*65173*/;
assign _19954_ = _19248_ & _19957_ /*65169*/;
assign _19955_ = _19248_ ^ _19957_ /*65172*/;
assign _19956_ = _19948_ & _19955_ /*65170*/;
assign _19697_ = _19948_ ^ _19955_ /*65171*/;
assign _19953_ = _19954_ | _19956_ /*65168*/;
assign _19962_ = ~D[49] /*65167*/;
assign _19959_ = _19249_ & _19962_ /*65163*/;
assign _19960_ = _19249_ ^ _19962_ /*65166*/;
assign _19961_ = _19953_ & _19960_ /*65164*/;
assign _19698_ = _19953_ ^ _19960_ /*65165*/;
assign _19958_ = _19959_ | _19961_ /*65162*/;
assign _19967_ = ~D[50] /*65161*/;
assign _19964_ = _19250_ & _19967_ /*65157*/;
assign _19965_ = _19250_ ^ _19967_ /*65160*/;
assign _19966_ = _19958_ & _19965_ /*65158*/;
assign _19699_ = _19958_ ^ _19965_ /*65159*/;
assign _19963_ = _19964_ | _19966_ /*65156*/;
assign _19972_ = ~D[51] /*65155*/;
assign _19969_ = _19251_ & _19972_ /*65151*/;
assign _19970_ = _19251_ ^ _19972_ /*65154*/;
assign _19971_ = _19963_ & _19970_ /*65152*/;
assign _19700_ = _19963_ ^ _19970_ /*65153*/;
assign _19968_ = _19969_ | _19971_ /*65150*/;
assign _19977_ = ~D[52] /*65149*/;
assign _19974_ = _19252_ & _19977_ /*65145*/;
assign _19975_ = _19252_ ^ _19977_ /*65148*/;
assign _19976_ = _19968_ & _19975_ /*65146*/;
assign _19701_ = _19968_ ^ _19975_ /*65147*/;
assign _19973_ = _19974_ | _19976_ /*65144*/;
assign _19982_ = ~D[53] /*65143*/;
assign _19979_ = _19253_ & _19982_ /*65139*/;
assign _19980_ = _19253_ ^ _19982_ /*65142*/;
assign _19981_ = _19973_ & _19980_ /*65140*/;
assign _19702_ = _19973_ ^ _19980_ /*65141*/;
assign _19978_ = _19979_ | _19981_ /*65138*/;
assign _19987_ = ~D[54] /*65137*/;
assign _19984_ = _19254_ & _19987_ /*65133*/;
assign _19985_ = _19254_ ^ _19987_ /*65136*/;
assign _19986_ = _19978_ & _19985_ /*65134*/;
assign _19703_ = _19978_ ^ _19985_ /*65135*/;
assign _19983_ = _19984_ | _19986_ /*65132*/;
assign _19992_ = ~D[55] /*65131*/;
assign _19989_ = _19255_ & _19992_ /*65127*/;
assign _19990_ = _19255_ ^ _19992_ /*65130*/;
assign _19991_ = _19983_ & _19990_ /*65128*/;
assign _19704_ = _19983_ ^ _19990_ /*65129*/;
assign _19988_ = _19989_ | _19991_ /*65126*/;
assign _19997_ = ~D[56] /*65125*/;
assign _19994_ = _19256_ & _19997_ /*65121*/;
assign _19995_ = _19256_ ^ _19997_ /*65124*/;
assign _19996_ = _19988_ & _19995_ /*65122*/;
assign _19705_ = _19988_ ^ _19995_ /*65123*/;
assign _19993_ = _19994_ | _19996_ /*65120*/;
assign _20002_ = ~D[57] /*65119*/;
assign _19999_ = _19257_ & _20002_ /*65115*/;
assign _20000_ = _19257_ ^ _20002_ /*65118*/;
assign _20001_ = _19993_ & _20000_ /*65116*/;
assign _19706_ = _19993_ ^ _20000_ /*65117*/;
assign _19998_ = _19999_ | _20001_ /*65114*/;
assign _20007_ = ~D[58] /*65113*/;
assign _20004_ = _19258_ & _20007_ /*65109*/;
assign _20005_ = _19258_ ^ _20007_ /*65112*/;
assign _20006_ = _19998_ & _20005_ /*65110*/;
assign _19707_ = _19998_ ^ _20005_ /*65111*/;
assign _20003_ = _20004_ | _20006_ /*65108*/;
assign _20012_ = ~D[59] /*65107*/;
assign _20009_ = _19259_ & _20012_ /*65103*/;
assign _20010_ = _19259_ ^ _20012_ /*65106*/;
assign _20011_ = _20003_ & _20010_ /*65104*/;
assign _19708_ = _20003_ ^ _20010_ /*65105*/;
assign _20008_ = _20009_ | _20011_ /*65102*/;
assign _20017_ = ~D[60] /*65101*/;
assign _20014_ = _19260_ & _20017_ /*65097*/;
assign _20015_ = _19260_ ^ _20017_ /*65100*/;
assign _20016_ = _20008_ & _20015_ /*65098*/;
assign _19709_ = _20008_ ^ _20015_ /*65099*/;
assign _20013_ = _20014_ | _20016_ /*65096*/;
assign _20022_ = ~D[61] /*65095*/;
assign _20019_ = _19261_ & _20022_ /*65091*/;
assign _20020_ = _19261_ ^ _20022_ /*65094*/;
assign _20021_ = _20013_ & _20020_ /*65092*/;
assign _19710_ = _20013_ ^ _20020_ /*65093*/;
assign _20018_ = _20019_ | _20021_ /*65090*/;
assign _20027_ = ~D[62] /*65089*/;
assign _20024_ = _19262_ & _20027_ /*65085*/;
assign _20025_ = _19262_ ^ _20027_ /*65088*/;
assign _20026_ = _20018_ & _20025_ /*65086*/;
assign _19711_ = _20018_ ^ _20025_ /*65087*/;
assign _20023_ = _20024_ | _20026_ /*65084*/;
assign _20028_ = _19263_ & oneWire /*65079*/;
assign _20029_ = _19263_ ^ oneWire /*65082*/;
assign _20030_ = _20023_ & _20029_ /*65080*/;
assign _19712_ = _20023_ ^ _20029_ /*65081*/;
assign Q[41] = _20028_ | _20030_ /*65078*/;
assign _20163_ = ~Q[41] /*64693*/;
assign _20162_ = _20163_ & D[0] /*64692*/;
assign _20165_ = _19649_ & _20162_ /*64687*/;
assign _20166_ = _19649_ ^ _20162_ /*64690*/;
assign _20167_ = zeroWire & _20166_ /*64688*/;
assign _20097_ = zeroWire ^ _20166_ /*64689*/;
assign _20164_ = _20165_ | _20167_ /*64686*/;
assign _20169_ = ~Q[41] /*64685*/;
assign _20168_ = _20169_ & D[1] /*64684*/;
assign _20171_ = _19650_ & _20168_ /*64679*/;
assign _20172_ = _19650_ ^ _20168_ /*64682*/;
assign _20173_ = _20164_ & _20172_ /*64680*/;
assign _20098_ = _20164_ ^ _20172_ /*64681*/;
assign _20170_ = _20171_ | _20173_ /*64678*/;
assign _20175_ = ~Q[41] /*64677*/;
assign _20174_ = _20175_ & D[2] /*64676*/;
assign _20177_ = _19651_ & _20174_ /*64671*/;
assign _20178_ = _19651_ ^ _20174_ /*64674*/;
assign _20179_ = _20170_ & _20178_ /*64672*/;
assign _20099_ = _20170_ ^ _20178_ /*64673*/;
assign _20176_ = _20177_ | _20179_ /*64670*/;
assign _20181_ = ~Q[41] /*64669*/;
assign _20180_ = _20181_ & D[3] /*64668*/;
assign _20183_ = _19652_ & _20180_ /*64663*/;
assign _20184_ = _19652_ ^ _20180_ /*64666*/;
assign _20185_ = _20176_ & _20184_ /*64664*/;
assign _20100_ = _20176_ ^ _20184_ /*64665*/;
assign _20182_ = _20183_ | _20185_ /*64662*/;
assign _20187_ = ~Q[41] /*64661*/;
assign _20186_ = _20187_ & D[4] /*64660*/;
assign _20189_ = _19653_ & _20186_ /*64655*/;
assign _20190_ = _19653_ ^ _20186_ /*64658*/;
assign _20191_ = _20182_ & _20190_ /*64656*/;
assign _20101_ = _20182_ ^ _20190_ /*64657*/;
assign _20188_ = _20189_ | _20191_ /*64654*/;
assign _20193_ = ~Q[41] /*64653*/;
assign _20192_ = _20193_ & D[5] /*64652*/;
assign _20195_ = _19654_ & _20192_ /*64647*/;
assign _20196_ = _19654_ ^ _20192_ /*64650*/;
assign _20197_ = _20188_ & _20196_ /*64648*/;
assign _20102_ = _20188_ ^ _20196_ /*64649*/;
assign _20194_ = _20195_ | _20197_ /*64646*/;
assign _20199_ = ~Q[41] /*64645*/;
assign _20198_ = _20199_ & D[6] /*64644*/;
assign _20201_ = _19655_ & _20198_ /*64639*/;
assign _20202_ = _19655_ ^ _20198_ /*64642*/;
assign _20203_ = _20194_ & _20202_ /*64640*/;
assign _20103_ = _20194_ ^ _20202_ /*64641*/;
assign _20200_ = _20201_ | _20203_ /*64638*/;
assign _20205_ = ~Q[41] /*64637*/;
assign _20204_ = _20205_ & D[7] /*64636*/;
assign _20207_ = _19656_ & _20204_ /*64631*/;
assign _20208_ = _19656_ ^ _20204_ /*64634*/;
assign _20209_ = _20200_ & _20208_ /*64632*/;
assign _20104_ = _20200_ ^ _20208_ /*64633*/;
assign _20206_ = _20207_ | _20209_ /*64630*/;
assign _20211_ = ~Q[41] /*64629*/;
assign _20210_ = _20211_ & D[8] /*64628*/;
assign _20213_ = _19657_ & _20210_ /*64623*/;
assign _20214_ = _19657_ ^ _20210_ /*64626*/;
assign _20215_ = _20206_ & _20214_ /*64624*/;
assign _20105_ = _20206_ ^ _20214_ /*64625*/;
assign _20212_ = _20213_ | _20215_ /*64622*/;
assign _20217_ = ~Q[41] /*64621*/;
assign _20216_ = _20217_ & D[9] /*64620*/;
assign _20219_ = _19658_ & _20216_ /*64615*/;
assign _20220_ = _19658_ ^ _20216_ /*64618*/;
assign _20221_ = _20212_ & _20220_ /*64616*/;
assign _20106_ = _20212_ ^ _20220_ /*64617*/;
assign _20218_ = _20219_ | _20221_ /*64614*/;
assign _20223_ = ~Q[41] /*64613*/;
assign _20222_ = _20223_ & D[10] /*64612*/;
assign _20225_ = _19659_ & _20222_ /*64607*/;
assign _20226_ = _19659_ ^ _20222_ /*64610*/;
assign _20227_ = _20218_ & _20226_ /*64608*/;
assign _20107_ = _20218_ ^ _20226_ /*64609*/;
assign _20224_ = _20225_ | _20227_ /*64606*/;
assign _20229_ = ~Q[41] /*64605*/;
assign _20228_ = _20229_ & D[11] /*64604*/;
assign _20231_ = _19660_ & _20228_ /*64599*/;
assign _20232_ = _19660_ ^ _20228_ /*64602*/;
assign _20233_ = _20224_ & _20232_ /*64600*/;
assign _20108_ = _20224_ ^ _20232_ /*64601*/;
assign _20230_ = _20231_ | _20233_ /*64598*/;
assign _20235_ = ~Q[41] /*64597*/;
assign _20234_ = _20235_ & D[12] /*64596*/;
assign _20237_ = _19661_ & _20234_ /*64591*/;
assign _20238_ = _19661_ ^ _20234_ /*64594*/;
assign _20239_ = _20230_ & _20238_ /*64592*/;
assign _20109_ = _20230_ ^ _20238_ /*64593*/;
assign _20236_ = _20237_ | _20239_ /*64590*/;
assign _20241_ = ~Q[41] /*64589*/;
assign _20240_ = _20241_ & D[13] /*64588*/;
assign _20243_ = _19662_ & _20240_ /*64583*/;
assign _20244_ = _19662_ ^ _20240_ /*64586*/;
assign _20245_ = _20236_ & _20244_ /*64584*/;
assign _20110_ = _20236_ ^ _20244_ /*64585*/;
assign _20242_ = _20243_ | _20245_ /*64582*/;
assign _20247_ = ~Q[41] /*64581*/;
assign _20246_ = _20247_ & D[14] /*64580*/;
assign _20249_ = _19663_ & _20246_ /*64575*/;
assign _20250_ = _19663_ ^ _20246_ /*64578*/;
assign _20251_ = _20242_ & _20250_ /*64576*/;
assign _20111_ = _20242_ ^ _20250_ /*64577*/;
assign _20248_ = _20249_ | _20251_ /*64574*/;
assign _20253_ = ~Q[41] /*64573*/;
assign _20252_ = _20253_ & D[15] /*64572*/;
assign _20255_ = _19664_ & _20252_ /*64567*/;
assign _20256_ = _19664_ ^ _20252_ /*64570*/;
assign _20257_ = _20248_ & _20256_ /*64568*/;
assign _20112_ = _20248_ ^ _20256_ /*64569*/;
assign _20254_ = _20255_ | _20257_ /*64566*/;
assign _20259_ = ~Q[41] /*64565*/;
assign _20258_ = _20259_ & D[16] /*64564*/;
assign _20261_ = _19665_ & _20258_ /*64559*/;
assign _20262_ = _19665_ ^ _20258_ /*64562*/;
assign _20263_ = _20254_ & _20262_ /*64560*/;
assign _20113_ = _20254_ ^ _20262_ /*64561*/;
assign _20260_ = _20261_ | _20263_ /*64558*/;
assign _20265_ = ~Q[41] /*64557*/;
assign _20264_ = _20265_ & D[17] /*64556*/;
assign _20267_ = _19666_ & _20264_ /*64551*/;
assign _20268_ = _19666_ ^ _20264_ /*64554*/;
assign _20269_ = _20260_ & _20268_ /*64552*/;
assign _20114_ = _20260_ ^ _20268_ /*64553*/;
assign _20266_ = _20267_ | _20269_ /*64550*/;
assign _20271_ = ~Q[41] /*64549*/;
assign _20270_ = _20271_ & D[18] /*64548*/;
assign _20273_ = _19667_ & _20270_ /*64543*/;
assign _20274_ = _19667_ ^ _20270_ /*64546*/;
assign _20275_ = _20266_ & _20274_ /*64544*/;
assign _20115_ = _20266_ ^ _20274_ /*64545*/;
assign _20272_ = _20273_ | _20275_ /*64542*/;
assign _20277_ = ~Q[41] /*64541*/;
assign _20276_ = _20277_ & D[19] /*64540*/;
assign _20279_ = _19668_ & _20276_ /*64535*/;
assign _20280_ = _19668_ ^ _20276_ /*64538*/;
assign _20281_ = _20272_ & _20280_ /*64536*/;
assign _20116_ = _20272_ ^ _20280_ /*64537*/;
assign _20278_ = _20279_ | _20281_ /*64534*/;
assign _20283_ = ~Q[41] /*64533*/;
assign _20282_ = _20283_ & D[20] /*64532*/;
assign _20285_ = _19669_ & _20282_ /*64527*/;
assign _20286_ = _19669_ ^ _20282_ /*64530*/;
assign _20287_ = _20278_ & _20286_ /*64528*/;
assign _20117_ = _20278_ ^ _20286_ /*64529*/;
assign _20284_ = _20285_ | _20287_ /*64526*/;
assign _20289_ = ~Q[41] /*64525*/;
assign _20288_ = _20289_ & D[21] /*64524*/;
assign _20291_ = _19670_ & _20288_ /*64519*/;
assign _20292_ = _19670_ ^ _20288_ /*64522*/;
assign _20293_ = _20284_ & _20292_ /*64520*/;
assign _20118_ = _20284_ ^ _20292_ /*64521*/;
assign _20290_ = _20291_ | _20293_ /*64518*/;
assign _20295_ = ~Q[41] /*64517*/;
assign _20294_ = _20295_ & D[22] /*64516*/;
assign _20297_ = _19671_ & _20294_ /*64511*/;
assign _20298_ = _19671_ ^ _20294_ /*64514*/;
assign _20299_ = _20290_ & _20298_ /*64512*/;
assign _20119_ = _20290_ ^ _20298_ /*64513*/;
assign _20296_ = _20297_ | _20299_ /*64510*/;
assign _20301_ = ~Q[41] /*64509*/;
assign _20300_ = _20301_ & D[23] /*64508*/;
assign _20303_ = _19672_ & _20300_ /*64503*/;
assign _20304_ = _19672_ ^ _20300_ /*64506*/;
assign _20305_ = _20296_ & _20304_ /*64504*/;
assign _20120_ = _20296_ ^ _20304_ /*64505*/;
assign _20302_ = _20303_ | _20305_ /*64502*/;
assign _20307_ = ~Q[41] /*64501*/;
assign _20306_ = _20307_ & D[24] /*64500*/;
assign _20309_ = _19673_ & _20306_ /*64495*/;
assign _20310_ = _19673_ ^ _20306_ /*64498*/;
assign _20311_ = _20302_ & _20310_ /*64496*/;
assign _20121_ = _20302_ ^ _20310_ /*64497*/;
assign _20308_ = _20309_ | _20311_ /*64494*/;
assign _20313_ = ~Q[41] /*64493*/;
assign _20312_ = _20313_ & D[25] /*64492*/;
assign _20315_ = _19674_ & _20312_ /*64487*/;
assign _20316_ = _19674_ ^ _20312_ /*64490*/;
assign _20317_ = _20308_ & _20316_ /*64488*/;
assign _20122_ = _20308_ ^ _20316_ /*64489*/;
assign _20314_ = _20315_ | _20317_ /*64486*/;
assign _20319_ = ~Q[41] /*64485*/;
assign _20318_ = _20319_ & D[26] /*64484*/;
assign _20321_ = _19675_ & _20318_ /*64479*/;
assign _20322_ = _19675_ ^ _20318_ /*64482*/;
assign _20323_ = _20314_ & _20322_ /*64480*/;
assign _20123_ = _20314_ ^ _20322_ /*64481*/;
assign _20320_ = _20321_ | _20323_ /*64478*/;
assign _20325_ = ~Q[41] /*64477*/;
assign _20324_ = _20325_ & D[27] /*64476*/;
assign _20327_ = _19676_ & _20324_ /*64471*/;
assign _20328_ = _19676_ ^ _20324_ /*64474*/;
assign _20329_ = _20320_ & _20328_ /*64472*/;
assign _20124_ = _20320_ ^ _20328_ /*64473*/;
assign _20326_ = _20327_ | _20329_ /*64470*/;
assign _20331_ = ~Q[41] /*64469*/;
assign _20330_ = _20331_ & D[28] /*64468*/;
assign _20333_ = _19677_ & _20330_ /*64463*/;
assign _20334_ = _19677_ ^ _20330_ /*64466*/;
assign _20335_ = _20326_ & _20334_ /*64464*/;
assign _20125_ = _20326_ ^ _20334_ /*64465*/;
assign _20332_ = _20333_ | _20335_ /*64462*/;
assign _20337_ = ~Q[41] /*64461*/;
assign _20336_ = _20337_ & D[29] /*64460*/;
assign _20339_ = _19678_ & _20336_ /*64455*/;
assign _20340_ = _19678_ ^ _20336_ /*64458*/;
assign _20341_ = _20332_ & _20340_ /*64456*/;
assign _20126_ = _20332_ ^ _20340_ /*64457*/;
assign _20338_ = _20339_ | _20341_ /*64454*/;
assign _20343_ = ~Q[41] /*64453*/;
assign _20342_ = _20343_ & D[30] /*64452*/;
assign _20345_ = _19679_ & _20342_ /*64447*/;
assign _20346_ = _19679_ ^ _20342_ /*64450*/;
assign _20347_ = _20338_ & _20346_ /*64448*/;
assign _20127_ = _20338_ ^ _20346_ /*64449*/;
assign _20344_ = _20345_ | _20347_ /*64446*/;
assign _20349_ = ~Q[41] /*64445*/;
assign _20348_ = _20349_ & D[31] /*64444*/;
assign _20351_ = _19680_ & _20348_ /*64439*/;
assign _20352_ = _19680_ ^ _20348_ /*64442*/;
assign _20353_ = _20344_ & _20352_ /*64440*/;
assign _20128_ = _20344_ ^ _20352_ /*64441*/;
assign _20350_ = _20351_ | _20353_ /*64438*/;
assign _20355_ = ~Q[41] /*64437*/;
assign _20354_ = _20355_ & D[32] /*64436*/;
assign _20357_ = _19681_ & _20354_ /*64431*/;
assign _20358_ = _19681_ ^ _20354_ /*64434*/;
assign _20359_ = _20350_ & _20358_ /*64432*/;
assign _20129_ = _20350_ ^ _20358_ /*64433*/;
assign _20356_ = _20357_ | _20359_ /*64430*/;
assign _20361_ = ~Q[41] /*64429*/;
assign _20360_ = _20361_ & D[33] /*64428*/;
assign _20363_ = _19682_ & _20360_ /*64423*/;
assign _20364_ = _19682_ ^ _20360_ /*64426*/;
assign _20365_ = _20356_ & _20364_ /*64424*/;
assign _20130_ = _20356_ ^ _20364_ /*64425*/;
assign _20362_ = _20363_ | _20365_ /*64422*/;
assign _20367_ = ~Q[41] /*64421*/;
assign _20366_ = _20367_ & D[34] /*64420*/;
assign _20369_ = _19683_ & _20366_ /*64415*/;
assign _20370_ = _19683_ ^ _20366_ /*64418*/;
assign _20371_ = _20362_ & _20370_ /*64416*/;
assign _20131_ = _20362_ ^ _20370_ /*64417*/;
assign _20368_ = _20369_ | _20371_ /*64414*/;
assign _20373_ = ~Q[41] /*64413*/;
assign _20372_ = _20373_ & D[35] /*64412*/;
assign _20375_ = _19684_ & _20372_ /*64407*/;
assign _20376_ = _19684_ ^ _20372_ /*64410*/;
assign _20377_ = _20368_ & _20376_ /*64408*/;
assign _20132_ = _20368_ ^ _20376_ /*64409*/;
assign _20374_ = _20375_ | _20377_ /*64406*/;
assign _20379_ = ~Q[41] /*64405*/;
assign _20378_ = _20379_ & D[36] /*64404*/;
assign _20381_ = _19685_ & _20378_ /*64399*/;
assign _20382_ = _19685_ ^ _20378_ /*64402*/;
assign _20383_ = _20374_ & _20382_ /*64400*/;
assign _20133_ = _20374_ ^ _20382_ /*64401*/;
assign _20380_ = _20381_ | _20383_ /*64398*/;
assign _20385_ = ~Q[41] /*64397*/;
assign _20384_ = _20385_ & D[37] /*64396*/;
assign _20387_ = _19686_ & _20384_ /*64391*/;
assign _20388_ = _19686_ ^ _20384_ /*64394*/;
assign _20389_ = _20380_ & _20388_ /*64392*/;
assign _20134_ = _20380_ ^ _20388_ /*64393*/;
assign _20386_ = _20387_ | _20389_ /*64390*/;
assign _20391_ = ~Q[41] /*64389*/;
assign _20390_ = _20391_ & D[38] /*64388*/;
assign _20393_ = _19687_ & _20390_ /*64383*/;
assign _20394_ = _19687_ ^ _20390_ /*64386*/;
assign _20395_ = _20386_ & _20394_ /*64384*/;
assign _20135_ = _20386_ ^ _20394_ /*64385*/;
assign _20392_ = _20393_ | _20395_ /*64382*/;
assign _20397_ = ~Q[41] /*64381*/;
assign _20396_ = _20397_ & D[39] /*64380*/;
assign _20399_ = _19688_ & _20396_ /*64375*/;
assign _20400_ = _19688_ ^ _20396_ /*64378*/;
assign _20401_ = _20392_ & _20400_ /*64376*/;
assign _20136_ = _20392_ ^ _20400_ /*64377*/;
assign _20398_ = _20399_ | _20401_ /*64374*/;
assign _20403_ = ~Q[41] /*64373*/;
assign _20402_ = _20403_ & D[40] /*64372*/;
assign _20405_ = _19689_ & _20402_ /*64367*/;
assign _20406_ = _19689_ ^ _20402_ /*64370*/;
assign _20407_ = _20398_ & _20406_ /*64368*/;
assign _20137_ = _20398_ ^ _20406_ /*64369*/;
assign _20404_ = _20405_ | _20407_ /*64366*/;
assign _20409_ = ~Q[41] /*64365*/;
assign _20408_ = _20409_ & D[41] /*64364*/;
assign _20411_ = _19690_ & _20408_ /*64359*/;
assign _20412_ = _19690_ ^ _20408_ /*64362*/;
assign _20413_ = _20404_ & _20412_ /*64360*/;
assign _20138_ = _20404_ ^ _20412_ /*64361*/;
assign _20410_ = _20411_ | _20413_ /*64358*/;
assign _20415_ = ~Q[41] /*64357*/;
assign _20414_ = _20415_ & D[42] /*64356*/;
assign _20417_ = _19691_ & _20414_ /*64351*/;
assign _20418_ = _19691_ ^ _20414_ /*64354*/;
assign _20419_ = _20410_ & _20418_ /*64352*/;
assign _20139_ = _20410_ ^ _20418_ /*64353*/;
assign _20416_ = _20417_ | _20419_ /*64350*/;
assign _20421_ = ~Q[41] /*64349*/;
assign _20420_ = _20421_ & D[43] /*64348*/;
assign _20423_ = _19692_ & _20420_ /*64343*/;
assign _20424_ = _19692_ ^ _20420_ /*64346*/;
assign _20425_ = _20416_ & _20424_ /*64344*/;
assign _20140_ = _20416_ ^ _20424_ /*64345*/;
assign _20422_ = _20423_ | _20425_ /*64342*/;
assign _20427_ = ~Q[41] /*64341*/;
assign _20426_ = _20427_ & D[44] /*64340*/;
assign _20429_ = _19693_ & _20426_ /*64335*/;
assign _20430_ = _19693_ ^ _20426_ /*64338*/;
assign _20431_ = _20422_ & _20430_ /*64336*/;
assign _20141_ = _20422_ ^ _20430_ /*64337*/;
assign _20428_ = _20429_ | _20431_ /*64334*/;
assign _20433_ = ~Q[41] /*64333*/;
assign _20432_ = _20433_ & D[45] /*64332*/;
assign _20435_ = _19694_ & _20432_ /*64327*/;
assign _20436_ = _19694_ ^ _20432_ /*64330*/;
assign _20437_ = _20428_ & _20436_ /*64328*/;
assign _20142_ = _20428_ ^ _20436_ /*64329*/;
assign _20434_ = _20435_ | _20437_ /*64326*/;
assign _20439_ = ~Q[41] /*64325*/;
assign _20438_ = _20439_ & D[46] /*64324*/;
assign _20441_ = _19695_ & _20438_ /*64319*/;
assign _20442_ = _19695_ ^ _20438_ /*64322*/;
assign _20443_ = _20434_ & _20442_ /*64320*/;
assign _20143_ = _20434_ ^ _20442_ /*64321*/;
assign _20440_ = _20441_ | _20443_ /*64318*/;
assign _20445_ = ~Q[41] /*64317*/;
assign _20444_ = _20445_ & D[47] /*64316*/;
assign _20447_ = _19696_ & _20444_ /*64311*/;
assign _20448_ = _19696_ ^ _20444_ /*64314*/;
assign _20449_ = _20440_ & _20448_ /*64312*/;
assign _20144_ = _20440_ ^ _20448_ /*64313*/;
assign _20446_ = _20447_ | _20449_ /*64310*/;
assign _20451_ = ~Q[41] /*64309*/;
assign _20450_ = _20451_ & D[48] /*64308*/;
assign _20453_ = _19697_ & _20450_ /*64303*/;
assign _20454_ = _19697_ ^ _20450_ /*64306*/;
assign _20455_ = _20446_ & _20454_ /*64304*/;
assign _20145_ = _20446_ ^ _20454_ /*64305*/;
assign _20452_ = _20453_ | _20455_ /*64302*/;
assign _20457_ = ~Q[41] /*64301*/;
assign _20456_ = _20457_ & D[49] /*64300*/;
assign _20459_ = _19698_ & _20456_ /*64295*/;
assign _20460_ = _19698_ ^ _20456_ /*64298*/;
assign _20461_ = _20452_ & _20460_ /*64296*/;
assign _20146_ = _20452_ ^ _20460_ /*64297*/;
assign _20458_ = _20459_ | _20461_ /*64294*/;
assign _20463_ = ~Q[41] /*64293*/;
assign _20462_ = _20463_ & D[50] /*64292*/;
assign _20465_ = _19699_ & _20462_ /*64287*/;
assign _20466_ = _19699_ ^ _20462_ /*64290*/;
assign _20467_ = _20458_ & _20466_ /*64288*/;
assign _20147_ = _20458_ ^ _20466_ /*64289*/;
assign _20464_ = _20465_ | _20467_ /*64286*/;
assign _20469_ = ~Q[41] /*64285*/;
assign _20468_ = _20469_ & D[51] /*64284*/;
assign _20471_ = _19700_ & _20468_ /*64279*/;
assign _20472_ = _19700_ ^ _20468_ /*64282*/;
assign _20473_ = _20464_ & _20472_ /*64280*/;
assign _20148_ = _20464_ ^ _20472_ /*64281*/;
assign _20470_ = _20471_ | _20473_ /*64278*/;
assign _20475_ = ~Q[41] /*64277*/;
assign _20474_ = _20475_ & D[52] /*64276*/;
assign _20477_ = _19701_ & _20474_ /*64271*/;
assign _20478_ = _19701_ ^ _20474_ /*64274*/;
assign _20479_ = _20470_ & _20478_ /*64272*/;
assign _20149_ = _20470_ ^ _20478_ /*64273*/;
assign _20476_ = _20477_ | _20479_ /*64270*/;
assign _20481_ = ~Q[41] /*64269*/;
assign _20480_ = _20481_ & D[53] /*64268*/;
assign _20483_ = _19702_ & _20480_ /*64263*/;
assign _20484_ = _19702_ ^ _20480_ /*64266*/;
assign _20485_ = _20476_ & _20484_ /*64264*/;
assign _20150_ = _20476_ ^ _20484_ /*64265*/;
assign _20482_ = _20483_ | _20485_ /*64262*/;
assign _20487_ = ~Q[41] /*64261*/;
assign _20486_ = _20487_ & D[54] /*64260*/;
assign _20489_ = _19703_ & _20486_ /*64255*/;
assign _20490_ = _19703_ ^ _20486_ /*64258*/;
assign _20491_ = _20482_ & _20490_ /*64256*/;
assign _20151_ = _20482_ ^ _20490_ /*64257*/;
assign _20488_ = _20489_ | _20491_ /*64254*/;
assign _20493_ = ~Q[41] /*64253*/;
assign _20492_ = _20493_ & D[55] /*64252*/;
assign _20495_ = _19704_ & _20492_ /*64247*/;
assign _20496_ = _19704_ ^ _20492_ /*64250*/;
assign _20497_ = _20488_ & _20496_ /*64248*/;
assign _20152_ = _20488_ ^ _20496_ /*64249*/;
assign _20494_ = _20495_ | _20497_ /*64246*/;
assign _20499_ = ~Q[41] /*64245*/;
assign _20498_ = _20499_ & D[56] /*64244*/;
assign _20501_ = _19705_ & _20498_ /*64239*/;
assign _20502_ = _19705_ ^ _20498_ /*64242*/;
assign _20503_ = _20494_ & _20502_ /*64240*/;
assign _20153_ = _20494_ ^ _20502_ /*64241*/;
assign _20500_ = _20501_ | _20503_ /*64238*/;
assign _20505_ = ~Q[41] /*64237*/;
assign _20504_ = _20505_ & D[57] /*64236*/;
assign _20507_ = _19706_ & _20504_ /*64231*/;
assign _20508_ = _19706_ ^ _20504_ /*64234*/;
assign _20509_ = _20500_ & _20508_ /*64232*/;
assign _20154_ = _20500_ ^ _20508_ /*64233*/;
assign _20506_ = _20507_ | _20509_ /*64230*/;
assign _20511_ = ~Q[41] /*64229*/;
assign _20510_ = _20511_ & D[58] /*64228*/;
assign _20513_ = _19707_ & _20510_ /*64223*/;
assign _20514_ = _19707_ ^ _20510_ /*64226*/;
assign _20515_ = _20506_ & _20514_ /*64224*/;
assign _20155_ = _20506_ ^ _20514_ /*64225*/;
assign _20512_ = _20513_ | _20515_ /*64222*/;
assign _20517_ = ~Q[41] /*64221*/;
assign _20516_ = _20517_ & D[59] /*64220*/;
assign _20519_ = _19708_ & _20516_ /*64215*/;
assign _20520_ = _19708_ ^ _20516_ /*64218*/;
assign _20521_ = _20512_ & _20520_ /*64216*/;
assign _20156_ = _20512_ ^ _20520_ /*64217*/;
assign _20518_ = _20519_ | _20521_ /*64214*/;
assign _20523_ = ~Q[41] /*64213*/;
assign _20522_ = _20523_ & D[60] /*64212*/;
assign _20525_ = _19709_ & _20522_ /*64207*/;
assign _20526_ = _19709_ ^ _20522_ /*64210*/;
assign _20527_ = _20518_ & _20526_ /*64208*/;
assign _20157_ = _20518_ ^ _20526_ /*64209*/;
assign _20524_ = _20525_ | _20527_ /*64206*/;
assign _20529_ = ~Q[41] /*64205*/;
assign _20528_ = _20529_ & D[61] /*64204*/;
assign _20531_ = _19710_ & _20528_ /*64199*/;
assign _20532_ = _19710_ ^ _20528_ /*64202*/;
assign _20533_ = _20524_ & _20532_ /*64200*/;
assign _20158_ = _20524_ ^ _20532_ /*64201*/;
assign _20530_ = _20531_ | _20533_ /*64198*/;
assign _20535_ = ~Q[41] /*64197*/;
assign _20534_ = _20535_ & D[62] /*64196*/;
assign _20537_ = _19711_ & _20534_ /*64191*/;
assign _20538_ = _19711_ ^ _20534_ /*64194*/;
assign _20539_ = _20530_ & _20538_ /*64192*/;
assign _20159_ = _20530_ ^ _20538_ /*64193*/;
assign _20536_ = _20537_ | _20539_ /*64190*/;
assign _20541_ = ~Q[41] /*64189*/;
assign _20540_ = _20541_ & zeroWire /*64188*/;
assign _20542_ = _19712_ ^ _20540_ /*64186*/;
assign _20160_ = _20542_ ^ _20536_ /*64185*/;
assign _20613_ = ~D[0] /*63931*/;
assign _20610_ = R_0[40] & _20613_ /*63927*/;
assign _20611_ = R_0[40] ^ _20613_ /*63930*/;
assign _20612_ = oneWire & _20611_ /*63928*/;
assign _20545_ = oneWire ^ _20611_ /*63929*/;
assign _20609_ = _20610_ | _20612_ /*63926*/;
assign _20618_ = ~D[1] /*63925*/;
assign _20615_ = _20097_ & _20618_ /*63921*/;
assign _20616_ = _20097_ ^ _20618_ /*63924*/;
assign _20617_ = _20609_ & _20616_ /*63922*/;
assign _20546_ = _20609_ ^ _20616_ /*63923*/;
assign _20614_ = _20615_ | _20617_ /*63920*/;
assign _20623_ = ~D[2] /*63919*/;
assign _20620_ = _20098_ & _20623_ /*63915*/;
assign _20621_ = _20098_ ^ _20623_ /*63918*/;
assign _20622_ = _20614_ & _20621_ /*63916*/;
assign _20547_ = _20614_ ^ _20621_ /*63917*/;
assign _20619_ = _20620_ | _20622_ /*63914*/;
assign _20628_ = ~D[3] /*63913*/;
assign _20625_ = _20099_ & _20628_ /*63909*/;
assign _20626_ = _20099_ ^ _20628_ /*63912*/;
assign _20627_ = _20619_ & _20626_ /*63910*/;
assign _20548_ = _20619_ ^ _20626_ /*63911*/;
assign _20624_ = _20625_ | _20627_ /*63908*/;
assign _20633_ = ~D[4] /*63907*/;
assign _20630_ = _20100_ & _20633_ /*63903*/;
assign _20631_ = _20100_ ^ _20633_ /*63906*/;
assign _20632_ = _20624_ & _20631_ /*63904*/;
assign _20549_ = _20624_ ^ _20631_ /*63905*/;
assign _20629_ = _20630_ | _20632_ /*63902*/;
assign _20638_ = ~D[5] /*63901*/;
assign _20635_ = _20101_ & _20638_ /*63897*/;
assign _20636_ = _20101_ ^ _20638_ /*63900*/;
assign _20637_ = _20629_ & _20636_ /*63898*/;
assign _20550_ = _20629_ ^ _20636_ /*63899*/;
assign _20634_ = _20635_ | _20637_ /*63896*/;
assign _20643_ = ~D[6] /*63895*/;
assign _20640_ = _20102_ & _20643_ /*63891*/;
assign _20641_ = _20102_ ^ _20643_ /*63894*/;
assign _20642_ = _20634_ & _20641_ /*63892*/;
assign _20551_ = _20634_ ^ _20641_ /*63893*/;
assign _20639_ = _20640_ | _20642_ /*63890*/;
assign _20648_ = ~D[7] /*63889*/;
assign _20645_ = _20103_ & _20648_ /*63885*/;
assign _20646_ = _20103_ ^ _20648_ /*63888*/;
assign _20647_ = _20639_ & _20646_ /*63886*/;
assign _20552_ = _20639_ ^ _20646_ /*63887*/;
assign _20644_ = _20645_ | _20647_ /*63884*/;
assign _20653_ = ~D[8] /*63883*/;
assign _20650_ = _20104_ & _20653_ /*63879*/;
assign _20651_ = _20104_ ^ _20653_ /*63882*/;
assign _20652_ = _20644_ & _20651_ /*63880*/;
assign _20553_ = _20644_ ^ _20651_ /*63881*/;
assign _20649_ = _20650_ | _20652_ /*63878*/;
assign _20658_ = ~D[9] /*63877*/;
assign _20655_ = _20105_ & _20658_ /*63873*/;
assign _20656_ = _20105_ ^ _20658_ /*63876*/;
assign _20657_ = _20649_ & _20656_ /*63874*/;
assign _20554_ = _20649_ ^ _20656_ /*63875*/;
assign _20654_ = _20655_ | _20657_ /*63872*/;
assign _20663_ = ~D[10] /*63871*/;
assign _20660_ = _20106_ & _20663_ /*63867*/;
assign _20661_ = _20106_ ^ _20663_ /*63870*/;
assign _20662_ = _20654_ & _20661_ /*63868*/;
assign _20555_ = _20654_ ^ _20661_ /*63869*/;
assign _20659_ = _20660_ | _20662_ /*63866*/;
assign _20668_ = ~D[11] /*63865*/;
assign _20665_ = _20107_ & _20668_ /*63861*/;
assign _20666_ = _20107_ ^ _20668_ /*63864*/;
assign _20667_ = _20659_ & _20666_ /*63862*/;
assign _20556_ = _20659_ ^ _20666_ /*63863*/;
assign _20664_ = _20665_ | _20667_ /*63860*/;
assign _20673_ = ~D[12] /*63859*/;
assign _20670_ = _20108_ & _20673_ /*63855*/;
assign _20671_ = _20108_ ^ _20673_ /*63858*/;
assign _20672_ = _20664_ & _20671_ /*63856*/;
assign _20557_ = _20664_ ^ _20671_ /*63857*/;
assign _20669_ = _20670_ | _20672_ /*63854*/;
assign _20678_ = ~D[13] /*63853*/;
assign _20675_ = _20109_ & _20678_ /*63849*/;
assign _20676_ = _20109_ ^ _20678_ /*63852*/;
assign _20677_ = _20669_ & _20676_ /*63850*/;
assign _20558_ = _20669_ ^ _20676_ /*63851*/;
assign _20674_ = _20675_ | _20677_ /*63848*/;
assign _20683_ = ~D[14] /*63847*/;
assign _20680_ = _20110_ & _20683_ /*63843*/;
assign _20681_ = _20110_ ^ _20683_ /*63846*/;
assign _20682_ = _20674_ & _20681_ /*63844*/;
assign _20559_ = _20674_ ^ _20681_ /*63845*/;
assign _20679_ = _20680_ | _20682_ /*63842*/;
assign _20688_ = ~D[15] /*63841*/;
assign _20685_ = _20111_ & _20688_ /*63837*/;
assign _20686_ = _20111_ ^ _20688_ /*63840*/;
assign _20687_ = _20679_ & _20686_ /*63838*/;
assign _20560_ = _20679_ ^ _20686_ /*63839*/;
assign _20684_ = _20685_ | _20687_ /*63836*/;
assign _20693_ = ~D[16] /*63835*/;
assign _20690_ = _20112_ & _20693_ /*63831*/;
assign _20691_ = _20112_ ^ _20693_ /*63834*/;
assign _20692_ = _20684_ & _20691_ /*63832*/;
assign _20561_ = _20684_ ^ _20691_ /*63833*/;
assign _20689_ = _20690_ | _20692_ /*63830*/;
assign _20698_ = ~D[17] /*63829*/;
assign _20695_ = _20113_ & _20698_ /*63825*/;
assign _20696_ = _20113_ ^ _20698_ /*63828*/;
assign _20697_ = _20689_ & _20696_ /*63826*/;
assign _20562_ = _20689_ ^ _20696_ /*63827*/;
assign _20694_ = _20695_ | _20697_ /*63824*/;
assign _20703_ = ~D[18] /*63823*/;
assign _20700_ = _20114_ & _20703_ /*63819*/;
assign _20701_ = _20114_ ^ _20703_ /*63822*/;
assign _20702_ = _20694_ & _20701_ /*63820*/;
assign _20563_ = _20694_ ^ _20701_ /*63821*/;
assign _20699_ = _20700_ | _20702_ /*63818*/;
assign _20708_ = ~D[19] /*63817*/;
assign _20705_ = _20115_ & _20708_ /*63813*/;
assign _20706_ = _20115_ ^ _20708_ /*63816*/;
assign _20707_ = _20699_ & _20706_ /*63814*/;
assign _20564_ = _20699_ ^ _20706_ /*63815*/;
assign _20704_ = _20705_ | _20707_ /*63812*/;
assign _20713_ = ~D[20] /*63811*/;
assign _20710_ = _20116_ & _20713_ /*63807*/;
assign _20711_ = _20116_ ^ _20713_ /*63810*/;
assign _20712_ = _20704_ & _20711_ /*63808*/;
assign _20565_ = _20704_ ^ _20711_ /*63809*/;
assign _20709_ = _20710_ | _20712_ /*63806*/;
assign _20718_ = ~D[21] /*63805*/;
assign _20715_ = _20117_ & _20718_ /*63801*/;
assign _20716_ = _20117_ ^ _20718_ /*63804*/;
assign _20717_ = _20709_ & _20716_ /*63802*/;
assign _20566_ = _20709_ ^ _20716_ /*63803*/;
assign _20714_ = _20715_ | _20717_ /*63800*/;
assign _20723_ = ~D[22] /*63799*/;
assign _20720_ = _20118_ & _20723_ /*63795*/;
assign _20721_ = _20118_ ^ _20723_ /*63798*/;
assign _20722_ = _20714_ & _20721_ /*63796*/;
assign _20567_ = _20714_ ^ _20721_ /*63797*/;
assign _20719_ = _20720_ | _20722_ /*63794*/;
assign _20728_ = ~D[23] /*63793*/;
assign _20725_ = _20119_ & _20728_ /*63789*/;
assign _20726_ = _20119_ ^ _20728_ /*63792*/;
assign _20727_ = _20719_ & _20726_ /*63790*/;
assign _20568_ = _20719_ ^ _20726_ /*63791*/;
assign _20724_ = _20725_ | _20727_ /*63788*/;
assign _20733_ = ~D[24] /*63787*/;
assign _20730_ = _20120_ & _20733_ /*63783*/;
assign _20731_ = _20120_ ^ _20733_ /*63786*/;
assign _20732_ = _20724_ & _20731_ /*63784*/;
assign _20569_ = _20724_ ^ _20731_ /*63785*/;
assign _20729_ = _20730_ | _20732_ /*63782*/;
assign _20738_ = ~D[25] /*63781*/;
assign _20735_ = _20121_ & _20738_ /*63777*/;
assign _20736_ = _20121_ ^ _20738_ /*63780*/;
assign _20737_ = _20729_ & _20736_ /*63778*/;
assign _20570_ = _20729_ ^ _20736_ /*63779*/;
assign _20734_ = _20735_ | _20737_ /*63776*/;
assign _20743_ = ~D[26] /*63775*/;
assign _20740_ = _20122_ & _20743_ /*63771*/;
assign _20741_ = _20122_ ^ _20743_ /*63774*/;
assign _20742_ = _20734_ & _20741_ /*63772*/;
assign _20571_ = _20734_ ^ _20741_ /*63773*/;
assign _20739_ = _20740_ | _20742_ /*63770*/;
assign _20748_ = ~D[27] /*63769*/;
assign _20745_ = _20123_ & _20748_ /*63765*/;
assign _20746_ = _20123_ ^ _20748_ /*63768*/;
assign _20747_ = _20739_ & _20746_ /*63766*/;
assign _20572_ = _20739_ ^ _20746_ /*63767*/;
assign _20744_ = _20745_ | _20747_ /*63764*/;
assign _20753_ = ~D[28] /*63763*/;
assign _20750_ = _20124_ & _20753_ /*63759*/;
assign _20751_ = _20124_ ^ _20753_ /*63762*/;
assign _20752_ = _20744_ & _20751_ /*63760*/;
assign _20573_ = _20744_ ^ _20751_ /*63761*/;
assign _20749_ = _20750_ | _20752_ /*63758*/;
assign _20758_ = ~D[29] /*63757*/;
assign _20755_ = _20125_ & _20758_ /*63753*/;
assign _20756_ = _20125_ ^ _20758_ /*63756*/;
assign _20757_ = _20749_ & _20756_ /*63754*/;
assign _20574_ = _20749_ ^ _20756_ /*63755*/;
assign _20754_ = _20755_ | _20757_ /*63752*/;
assign _20763_ = ~D[30] /*63751*/;
assign _20760_ = _20126_ & _20763_ /*63747*/;
assign _20761_ = _20126_ ^ _20763_ /*63750*/;
assign _20762_ = _20754_ & _20761_ /*63748*/;
assign _20575_ = _20754_ ^ _20761_ /*63749*/;
assign _20759_ = _20760_ | _20762_ /*63746*/;
assign _20768_ = ~D[31] /*63745*/;
assign _20765_ = _20127_ & _20768_ /*63741*/;
assign _20766_ = _20127_ ^ _20768_ /*63744*/;
assign _20767_ = _20759_ & _20766_ /*63742*/;
assign _20576_ = _20759_ ^ _20766_ /*63743*/;
assign _20764_ = _20765_ | _20767_ /*63740*/;
assign _20773_ = ~D[32] /*63739*/;
assign _20770_ = _20128_ & _20773_ /*63735*/;
assign _20771_ = _20128_ ^ _20773_ /*63738*/;
assign _20772_ = _20764_ & _20771_ /*63736*/;
assign _20577_ = _20764_ ^ _20771_ /*63737*/;
assign _20769_ = _20770_ | _20772_ /*63734*/;
assign _20778_ = ~D[33] /*63733*/;
assign _20775_ = _20129_ & _20778_ /*63729*/;
assign _20776_ = _20129_ ^ _20778_ /*63732*/;
assign _20777_ = _20769_ & _20776_ /*63730*/;
assign _20578_ = _20769_ ^ _20776_ /*63731*/;
assign _20774_ = _20775_ | _20777_ /*63728*/;
assign _20783_ = ~D[34] /*63727*/;
assign _20780_ = _20130_ & _20783_ /*63723*/;
assign _20781_ = _20130_ ^ _20783_ /*63726*/;
assign _20782_ = _20774_ & _20781_ /*63724*/;
assign _20579_ = _20774_ ^ _20781_ /*63725*/;
assign _20779_ = _20780_ | _20782_ /*63722*/;
assign _20788_ = ~D[35] /*63721*/;
assign _20785_ = _20131_ & _20788_ /*63717*/;
assign _20786_ = _20131_ ^ _20788_ /*63720*/;
assign _20787_ = _20779_ & _20786_ /*63718*/;
assign _20580_ = _20779_ ^ _20786_ /*63719*/;
assign _20784_ = _20785_ | _20787_ /*63716*/;
assign _20793_ = ~D[36] /*63715*/;
assign _20790_ = _20132_ & _20793_ /*63711*/;
assign _20791_ = _20132_ ^ _20793_ /*63714*/;
assign _20792_ = _20784_ & _20791_ /*63712*/;
assign _20581_ = _20784_ ^ _20791_ /*63713*/;
assign _20789_ = _20790_ | _20792_ /*63710*/;
assign _20798_ = ~D[37] /*63709*/;
assign _20795_ = _20133_ & _20798_ /*63705*/;
assign _20796_ = _20133_ ^ _20798_ /*63708*/;
assign _20797_ = _20789_ & _20796_ /*63706*/;
assign _20582_ = _20789_ ^ _20796_ /*63707*/;
assign _20794_ = _20795_ | _20797_ /*63704*/;
assign _20803_ = ~D[38] /*63703*/;
assign _20800_ = _20134_ & _20803_ /*63699*/;
assign _20801_ = _20134_ ^ _20803_ /*63702*/;
assign _20802_ = _20794_ & _20801_ /*63700*/;
assign _20583_ = _20794_ ^ _20801_ /*63701*/;
assign _20799_ = _20800_ | _20802_ /*63698*/;
assign _20808_ = ~D[39] /*63697*/;
assign _20805_ = _20135_ & _20808_ /*63693*/;
assign _20806_ = _20135_ ^ _20808_ /*63696*/;
assign _20807_ = _20799_ & _20806_ /*63694*/;
assign _20584_ = _20799_ ^ _20806_ /*63695*/;
assign _20804_ = _20805_ | _20807_ /*63692*/;
assign _20813_ = ~D[40] /*63691*/;
assign _20810_ = _20136_ & _20813_ /*63687*/;
assign _20811_ = _20136_ ^ _20813_ /*63690*/;
assign _20812_ = _20804_ & _20811_ /*63688*/;
assign _20585_ = _20804_ ^ _20811_ /*63689*/;
assign _20809_ = _20810_ | _20812_ /*63686*/;
assign _20818_ = ~D[41] /*63685*/;
assign _20815_ = _20137_ & _20818_ /*63681*/;
assign _20816_ = _20137_ ^ _20818_ /*63684*/;
assign _20817_ = _20809_ & _20816_ /*63682*/;
assign _20586_ = _20809_ ^ _20816_ /*63683*/;
assign _20814_ = _20815_ | _20817_ /*63680*/;
assign _20823_ = ~D[42] /*63679*/;
assign _20820_ = _20138_ & _20823_ /*63675*/;
assign _20821_ = _20138_ ^ _20823_ /*63678*/;
assign _20822_ = _20814_ & _20821_ /*63676*/;
assign _20587_ = _20814_ ^ _20821_ /*63677*/;
assign _20819_ = _20820_ | _20822_ /*63674*/;
assign _20828_ = ~D[43] /*63673*/;
assign _20825_ = _20139_ & _20828_ /*63669*/;
assign _20826_ = _20139_ ^ _20828_ /*63672*/;
assign _20827_ = _20819_ & _20826_ /*63670*/;
assign _20588_ = _20819_ ^ _20826_ /*63671*/;
assign _20824_ = _20825_ | _20827_ /*63668*/;
assign _20833_ = ~D[44] /*63667*/;
assign _20830_ = _20140_ & _20833_ /*63663*/;
assign _20831_ = _20140_ ^ _20833_ /*63666*/;
assign _20832_ = _20824_ & _20831_ /*63664*/;
assign _20589_ = _20824_ ^ _20831_ /*63665*/;
assign _20829_ = _20830_ | _20832_ /*63662*/;
assign _20838_ = ~D[45] /*63661*/;
assign _20835_ = _20141_ & _20838_ /*63657*/;
assign _20836_ = _20141_ ^ _20838_ /*63660*/;
assign _20837_ = _20829_ & _20836_ /*63658*/;
assign _20590_ = _20829_ ^ _20836_ /*63659*/;
assign _20834_ = _20835_ | _20837_ /*63656*/;
assign _20843_ = ~D[46] /*63655*/;
assign _20840_ = _20142_ & _20843_ /*63651*/;
assign _20841_ = _20142_ ^ _20843_ /*63654*/;
assign _20842_ = _20834_ & _20841_ /*63652*/;
assign _20591_ = _20834_ ^ _20841_ /*63653*/;
assign _20839_ = _20840_ | _20842_ /*63650*/;
assign _20848_ = ~D[47] /*63649*/;
assign _20845_ = _20143_ & _20848_ /*63645*/;
assign _20846_ = _20143_ ^ _20848_ /*63648*/;
assign _20847_ = _20839_ & _20846_ /*63646*/;
assign _20592_ = _20839_ ^ _20846_ /*63647*/;
assign _20844_ = _20845_ | _20847_ /*63644*/;
assign _20853_ = ~D[48] /*63643*/;
assign _20850_ = _20144_ & _20853_ /*63639*/;
assign _20851_ = _20144_ ^ _20853_ /*63642*/;
assign _20852_ = _20844_ & _20851_ /*63640*/;
assign _20593_ = _20844_ ^ _20851_ /*63641*/;
assign _20849_ = _20850_ | _20852_ /*63638*/;
assign _20858_ = ~D[49] /*63637*/;
assign _20855_ = _20145_ & _20858_ /*63633*/;
assign _20856_ = _20145_ ^ _20858_ /*63636*/;
assign _20857_ = _20849_ & _20856_ /*63634*/;
assign _20594_ = _20849_ ^ _20856_ /*63635*/;
assign _20854_ = _20855_ | _20857_ /*63632*/;
assign _20863_ = ~D[50] /*63631*/;
assign _20860_ = _20146_ & _20863_ /*63627*/;
assign _20861_ = _20146_ ^ _20863_ /*63630*/;
assign _20862_ = _20854_ & _20861_ /*63628*/;
assign _20595_ = _20854_ ^ _20861_ /*63629*/;
assign _20859_ = _20860_ | _20862_ /*63626*/;
assign _20868_ = ~D[51] /*63625*/;
assign _20865_ = _20147_ & _20868_ /*63621*/;
assign _20866_ = _20147_ ^ _20868_ /*63624*/;
assign _20867_ = _20859_ & _20866_ /*63622*/;
assign _20596_ = _20859_ ^ _20866_ /*63623*/;
assign _20864_ = _20865_ | _20867_ /*63620*/;
assign _20873_ = ~D[52] /*63619*/;
assign _20870_ = _20148_ & _20873_ /*63615*/;
assign _20871_ = _20148_ ^ _20873_ /*63618*/;
assign _20872_ = _20864_ & _20871_ /*63616*/;
assign _20597_ = _20864_ ^ _20871_ /*63617*/;
assign _20869_ = _20870_ | _20872_ /*63614*/;
assign _20878_ = ~D[53] /*63613*/;
assign _20875_ = _20149_ & _20878_ /*63609*/;
assign _20876_ = _20149_ ^ _20878_ /*63612*/;
assign _20877_ = _20869_ & _20876_ /*63610*/;
assign _20598_ = _20869_ ^ _20876_ /*63611*/;
assign _20874_ = _20875_ | _20877_ /*63608*/;
assign _20883_ = ~D[54] /*63607*/;
assign _20880_ = _20150_ & _20883_ /*63603*/;
assign _20881_ = _20150_ ^ _20883_ /*63606*/;
assign _20882_ = _20874_ & _20881_ /*63604*/;
assign _20599_ = _20874_ ^ _20881_ /*63605*/;
assign _20879_ = _20880_ | _20882_ /*63602*/;
assign _20888_ = ~D[55] /*63601*/;
assign _20885_ = _20151_ & _20888_ /*63597*/;
assign _20886_ = _20151_ ^ _20888_ /*63600*/;
assign _20887_ = _20879_ & _20886_ /*63598*/;
assign _20600_ = _20879_ ^ _20886_ /*63599*/;
assign _20884_ = _20885_ | _20887_ /*63596*/;
assign _20893_ = ~D[56] /*63595*/;
assign _20890_ = _20152_ & _20893_ /*63591*/;
assign _20891_ = _20152_ ^ _20893_ /*63594*/;
assign _20892_ = _20884_ & _20891_ /*63592*/;
assign _20601_ = _20884_ ^ _20891_ /*63593*/;
assign _20889_ = _20890_ | _20892_ /*63590*/;
assign _20898_ = ~D[57] /*63589*/;
assign _20895_ = _20153_ & _20898_ /*63585*/;
assign _20896_ = _20153_ ^ _20898_ /*63588*/;
assign _20897_ = _20889_ & _20896_ /*63586*/;
assign _20602_ = _20889_ ^ _20896_ /*63587*/;
assign _20894_ = _20895_ | _20897_ /*63584*/;
assign _20903_ = ~D[58] /*63583*/;
assign _20900_ = _20154_ & _20903_ /*63579*/;
assign _20901_ = _20154_ ^ _20903_ /*63582*/;
assign _20902_ = _20894_ & _20901_ /*63580*/;
assign _20603_ = _20894_ ^ _20901_ /*63581*/;
assign _20899_ = _20900_ | _20902_ /*63578*/;
assign _20908_ = ~D[59] /*63577*/;
assign _20905_ = _20155_ & _20908_ /*63573*/;
assign _20906_ = _20155_ ^ _20908_ /*63576*/;
assign _20907_ = _20899_ & _20906_ /*63574*/;
assign _20604_ = _20899_ ^ _20906_ /*63575*/;
assign _20904_ = _20905_ | _20907_ /*63572*/;
assign _20913_ = ~D[60] /*63571*/;
assign _20910_ = _20156_ & _20913_ /*63567*/;
assign _20911_ = _20156_ ^ _20913_ /*63570*/;
assign _20912_ = _20904_ & _20911_ /*63568*/;
assign _20605_ = _20904_ ^ _20911_ /*63569*/;
assign _20909_ = _20910_ | _20912_ /*63566*/;
assign _20918_ = ~D[61] /*63565*/;
assign _20915_ = _20157_ & _20918_ /*63561*/;
assign _20916_ = _20157_ ^ _20918_ /*63564*/;
assign _20917_ = _20909_ & _20916_ /*63562*/;
assign _20606_ = _20909_ ^ _20916_ /*63563*/;
assign _20914_ = _20915_ | _20917_ /*63560*/;
assign _20923_ = ~D[62] /*63559*/;
assign _20920_ = _20158_ & _20923_ /*63555*/;
assign _20921_ = _20158_ ^ _20923_ /*63558*/;
assign _20922_ = _20914_ & _20921_ /*63556*/;
assign _20607_ = _20914_ ^ _20921_ /*63557*/;
assign _20919_ = _20920_ | _20922_ /*63554*/;
assign _20924_ = _20159_ & oneWire /*63549*/;
assign _20925_ = _20159_ ^ oneWire /*63552*/;
assign _20926_ = _20919_ & _20925_ /*63550*/;
assign _20608_ = _20919_ ^ _20925_ /*63551*/;
assign Q[40] = _20924_ | _20926_ /*63548*/;
assign _21059_ = ~Q[40] /*63163*/;
assign _21058_ = _21059_ & D[0] /*63162*/;
assign _21061_ = _20545_ & _21058_ /*63157*/;
assign _21062_ = _20545_ ^ _21058_ /*63160*/;
assign _21063_ = zeroWire & _21062_ /*63158*/;
assign _20993_ = zeroWire ^ _21062_ /*63159*/;
assign _21060_ = _21061_ | _21063_ /*63156*/;
assign _21065_ = ~Q[40] /*63155*/;
assign _21064_ = _21065_ & D[1] /*63154*/;
assign _21067_ = _20546_ & _21064_ /*63149*/;
assign _21068_ = _20546_ ^ _21064_ /*63152*/;
assign _21069_ = _21060_ & _21068_ /*63150*/;
assign _20994_ = _21060_ ^ _21068_ /*63151*/;
assign _21066_ = _21067_ | _21069_ /*63148*/;
assign _21071_ = ~Q[40] /*63147*/;
assign _21070_ = _21071_ & D[2] /*63146*/;
assign _21073_ = _20547_ & _21070_ /*63141*/;
assign _21074_ = _20547_ ^ _21070_ /*63144*/;
assign _21075_ = _21066_ & _21074_ /*63142*/;
assign _20995_ = _21066_ ^ _21074_ /*63143*/;
assign _21072_ = _21073_ | _21075_ /*63140*/;
assign _21077_ = ~Q[40] /*63139*/;
assign _21076_ = _21077_ & D[3] /*63138*/;
assign _21079_ = _20548_ & _21076_ /*63133*/;
assign _21080_ = _20548_ ^ _21076_ /*63136*/;
assign _21081_ = _21072_ & _21080_ /*63134*/;
assign _20996_ = _21072_ ^ _21080_ /*63135*/;
assign _21078_ = _21079_ | _21081_ /*63132*/;
assign _21083_ = ~Q[40] /*63131*/;
assign _21082_ = _21083_ & D[4] /*63130*/;
assign _21085_ = _20549_ & _21082_ /*63125*/;
assign _21086_ = _20549_ ^ _21082_ /*63128*/;
assign _21087_ = _21078_ & _21086_ /*63126*/;
assign _20997_ = _21078_ ^ _21086_ /*63127*/;
assign _21084_ = _21085_ | _21087_ /*63124*/;
assign _21089_ = ~Q[40] /*63123*/;
assign _21088_ = _21089_ & D[5] /*63122*/;
assign _21091_ = _20550_ & _21088_ /*63117*/;
assign _21092_ = _20550_ ^ _21088_ /*63120*/;
assign _21093_ = _21084_ & _21092_ /*63118*/;
assign _20998_ = _21084_ ^ _21092_ /*63119*/;
assign _21090_ = _21091_ | _21093_ /*63116*/;
assign _21095_ = ~Q[40] /*63115*/;
assign _21094_ = _21095_ & D[6] /*63114*/;
assign _21097_ = _20551_ & _21094_ /*63109*/;
assign _21098_ = _20551_ ^ _21094_ /*63112*/;
assign _21099_ = _21090_ & _21098_ /*63110*/;
assign _20999_ = _21090_ ^ _21098_ /*63111*/;
assign _21096_ = _21097_ | _21099_ /*63108*/;
assign _21101_ = ~Q[40] /*63107*/;
assign _21100_ = _21101_ & D[7] /*63106*/;
assign _21103_ = _20552_ & _21100_ /*63101*/;
assign _21104_ = _20552_ ^ _21100_ /*63104*/;
assign _21105_ = _21096_ & _21104_ /*63102*/;
assign _21000_ = _21096_ ^ _21104_ /*63103*/;
assign _21102_ = _21103_ | _21105_ /*63100*/;
assign _21107_ = ~Q[40] /*63099*/;
assign _21106_ = _21107_ & D[8] /*63098*/;
assign _21109_ = _20553_ & _21106_ /*63093*/;
assign _21110_ = _20553_ ^ _21106_ /*63096*/;
assign _21111_ = _21102_ & _21110_ /*63094*/;
assign _21001_ = _21102_ ^ _21110_ /*63095*/;
assign _21108_ = _21109_ | _21111_ /*63092*/;
assign _21113_ = ~Q[40] /*63091*/;
assign _21112_ = _21113_ & D[9] /*63090*/;
assign _21115_ = _20554_ & _21112_ /*63085*/;
assign _21116_ = _20554_ ^ _21112_ /*63088*/;
assign _21117_ = _21108_ & _21116_ /*63086*/;
assign _21002_ = _21108_ ^ _21116_ /*63087*/;
assign _21114_ = _21115_ | _21117_ /*63084*/;
assign _21119_ = ~Q[40] /*63083*/;
assign _21118_ = _21119_ & D[10] /*63082*/;
assign _21121_ = _20555_ & _21118_ /*63077*/;
assign _21122_ = _20555_ ^ _21118_ /*63080*/;
assign _21123_ = _21114_ & _21122_ /*63078*/;
assign _21003_ = _21114_ ^ _21122_ /*63079*/;
assign _21120_ = _21121_ | _21123_ /*63076*/;
assign _21125_ = ~Q[40] /*63075*/;
assign _21124_ = _21125_ & D[11] /*63074*/;
assign _21127_ = _20556_ & _21124_ /*63069*/;
assign _21128_ = _20556_ ^ _21124_ /*63072*/;
assign _21129_ = _21120_ & _21128_ /*63070*/;
assign _21004_ = _21120_ ^ _21128_ /*63071*/;
assign _21126_ = _21127_ | _21129_ /*63068*/;
assign _21131_ = ~Q[40] /*63067*/;
assign _21130_ = _21131_ & D[12] /*63066*/;
assign _21133_ = _20557_ & _21130_ /*63061*/;
assign _21134_ = _20557_ ^ _21130_ /*63064*/;
assign _21135_ = _21126_ & _21134_ /*63062*/;
assign _21005_ = _21126_ ^ _21134_ /*63063*/;
assign _21132_ = _21133_ | _21135_ /*63060*/;
assign _21137_ = ~Q[40] /*63059*/;
assign _21136_ = _21137_ & D[13] /*63058*/;
assign _21139_ = _20558_ & _21136_ /*63053*/;
assign _21140_ = _20558_ ^ _21136_ /*63056*/;
assign _21141_ = _21132_ & _21140_ /*63054*/;
assign _21006_ = _21132_ ^ _21140_ /*63055*/;
assign _21138_ = _21139_ | _21141_ /*63052*/;
assign _21143_ = ~Q[40] /*63051*/;
assign _21142_ = _21143_ & D[14] /*63050*/;
assign _21145_ = _20559_ & _21142_ /*63045*/;
assign _21146_ = _20559_ ^ _21142_ /*63048*/;
assign _21147_ = _21138_ & _21146_ /*63046*/;
assign _21007_ = _21138_ ^ _21146_ /*63047*/;
assign _21144_ = _21145_ | _21147_ /*63044*/;
assign _21149_ = ~Q[40] /*63043*/;
assign _21148_ = _21149_ & D[15] /*63042*/;
assign _21151_ = _20560_ & _21148_ /*63037*/;
assign _21152_ = _20560_ ^ _21148_ /*63040*/;
assign _21153_ = _21144_ & _21152_ /*63038*/;
assign _21008_ = _21144_ ^ _21152_ /*63039*/;
assign _21150_ = _21151_ | _21153_ /*63036*/;
assign _21155_ = ~Q[40] /*63035*/;
assign _21154_ = _21155_ & D[16] /*63034*/;
assign _21157_ = _20561_ & _21154_ /*63029*/;
assign _21158_ = _20561_ ^ _21154_ /*63032*/;
assign _21159_ = _21150_ & _21158_ /*63030*/;
assign _21009_ = _21150_ ^ _21158_ /*63031*/;
assign _21156_ = _21157_ | _21159_ /*63028*/;
assign _21161_ = ~Q[40] /*63027*/;
assign _21160_ = _21161_ & D[17] /*63026*/;
assign _21163_ = _20562_ & _21160_ /*63021*/;
assign _21164_ = _20562_ ^ _21160_ /*63024*/;
assign _21165_ = _21156_ & _21164_ /*63022*/;
assign _21010_ = _21156_ ^ _21164_ /*63023*/;
assign _21162_ = _21163_ | _21165_ /*63020*/;
assign _21167_ = ~Q[40] /*63019*/;
assign _21166_ = _21167_ & D[18] /*63018*/;
assign _21169_ = _20563_ & _21166_ /*63013*/;
assign _21170_ = _20563_ ^ _21166_ /*63016*/;
assign _21171_ = _21162_ & _21170_ /*63014*/;
assign _21011_ = _21162_ ^ _21170_ /*63015*/;
assign _21168_ = _21169_ | _21171_ /*63012*/;
assign _21173_ = ~Q[40] /*63011*/;
assign _21172_ = _21173_ & D[19] /*63010*/;
assign _21175_ = _20564_ & _21172_ /*63005*/;
assign _21176_ = _20564_ ^ _21172_ /*63008*/;
assign _21177_ = _21168_ & _21176_ /*63006*/;
assign _21012_ = _21168_ ^ _21176_ /*63007*/;
assign _21174_ = _21175_ | _21177_ /*63004*/;
assign _21179_ = ~Q[40] /*63003*/;
assign _21178_ = _21179_ & D[20] /*63002*/;
assign _21181_ = _20565_ & _21178_ /*62997*/;
assign _21182_ = _20565_ ^ _21178_ /*63000*/;
assign _21183_ = _21174_ & _21182_ /*62998*/;
assign _21013_ = _21174_ ^ _21182_ /*62999*/;
assign _21180_ = _21181_ | _21183_ /*62996*/;
assign _21185_ = ~Q[40] /*62995*/;
assign _21184_ = _21185_ & D[21] /*62994*/;
assign _21187_ = _20566_ & _21184_ /*62989*/;
assign _21188_ = _20566_ ^ _21184_ /*62992*/;
assign _21189_ = _21180_ & _21188_ /*62990*/;
assign _21014_ = _21180_ ^ _21188_ /*62991*/;
assign _21186_ = _21187_ | _21189_ /*62988*/;
assign _21191_ = ~Q[40] /*62987*/;
assign _21190_ = _21191_ & D[22] /*62986*/;
assign _21193_ = _20567_ & _21190_ /*62981*/;
assign _21194_ = _20567_ ^ _21190_ /*62984*/;
assign _21195_ = _21186_ & _21194_ /*62982*/;
assign _21015_ = _21186_ ^ _21194_ /*62983*/;
assign _21192_ = _21193_ | _21195_ /*62980*/;
assign _21197_ = ~Q[40] /*62979*/;
assign _21196_ = _21197_ & D[23] /*62978*/;
assign _21199_ = _20568_ & _21196_ /*62973*/;
assign _21200_ = _20568_ ^ _21196_ /*62976*/;
assign _21201_ = _21192_ & _21200_ /*62974*/;
assign _21016_ = _21192_ ^ _21200_ /*62975*/;
assign _21198_ = _21199_ | _21201_ /*62972*/;
assign _21203_ = ~Q[40] /*62971*/;
assign _21202_ = _21203_ & D[24] /*62970*/;
assign _21205_ = _20569_ & _21202_ /*62965*/;
assign _21206_ = _20569_ ^ _21202_ /*62968*/;
assign _21207_ = _21198_ & _21206_ /*62966*/;
assign _21017_ = _21198_ ^ _21206_ /*62967*/;
assign _21204_ = _21205_ | _21207_ /*62964*/;
assign _21209_ = ~Q[40] /*62963*/;
assign _21208_ = _21209_ & D[25] /*62962*/;
assign _21211_ = _20570_ & _21208_ /*62957*/;
assign _21212_ = _20570_ ^ _21208_ /*62960*/;
assign _21213_ = _21204_ & _21212_ /*62958*/;
assign _21018_ = _21204_ ^ _21212_ /*62959*/;
assign _21210_ = _21211_ | _21213_ /*62956*/;
assign _21215_ = ~Q[40] /*62955*/;
assign _21214_ = _21215_ & D[26] /*62954*/;
assign _21217_ = _20571_ & _21214_ /*62949*/;
assign _21218_ = _20571_ ^ _21214_ /*62952*/;
assign _21219_ = _21210_ & _21218_ /*62950*/;
assign _21019_ = _21210_ ^ _21218_ /*62951*/;
assign _21216_ = _21217_ | _21219_ /*62948*/;
assign _21221_ = ~Q[40] /*62947*/;
assign _21220_ = _21221_ & D[27] /*62946*/;
assign _21223_ = _20572_ & _21220_ /*62941*/;
assign _21224_ = _20572_ ^ _21220_ /*62944*/;
assign _21225_ = _21216_ & _21224_ /*62942*/;
assign _21020_ = _21216_ ^ _21224_ /*62943*/;
assign _21222_ = _21223_ | _21225_ /*62940*/;
assign _21227_ = ~Q[40] /*62939*/;
assign _21226_ = _21227_ & D[28] /*62938*/;
assign _21229_ = _20573_ & _21226_ /*62933*/;
assign _21230_ = _20573_ ^ _21226_ /*62936*/;
assign _21231_ = _21222_ & _21230_ /*62934*/;
assign _21021_ = _21222_ ^ _21230_ /*62935*/;
assign _21228_ = _21229_ | _21231_ /*62932*/;
assign _21233_ = ~Q[40] /*62931*/;
assign _21232_ = _21233_ & D[29] /*62930*/;
assign _21235_ = _20574_ & _21232_ /*62925*/;
assign _21236_ = _20574_ ^ _21232_ /*62928*/;
assign _21237_ = _21228_ & _21236_ /*62926*/;
assign _21022_ = _21228_ ^ _21236_ /*62927*/;
assign _21234_ = _21235_ | _21237_ /*62924*/;
assign _21239_ = ~Q[40] /*62923*/;
assign _21238_ = _21239_ & D[30] /*62922*/;
assign _21241_ = _20575_ & _21238_ /*62917*/;
assign _21242_ = _20575_ ^ _21238_ /*62920*/;
assign _21243_ = _21234_ & _21242_ /*62918*/;
assign _21023_ = _21234_ ^ _21242_ /*62919*/;
assign _21240_ = _21241_ | _21243_ /*62916*/;
assign _21245_ = ~Q[40] /*62915*/;
assign _21244_ = _21245_ & D[31] /*62914*/;
assign _21247_ = _20576_ & _21244_ /*62909*/;
assign _21248_ = _20576_ ^ _21244_ /*62912*/;
assign _21249_ = _21240_ & _21248_ /*62910*/;
assign _21024_ = _21240_ ^ _21248_ /*62911*/;
assign _21246_ = _21247_ | _21249_ /*62908*/;
assign _21251_ = ~Q[40] /*62907*/;
assign _21250_ = _21251_ & D[32] /*62906*/;
assign _21253_ = _20577_ & _21250_ /*62901*/;
assign _21254_ = _20577_ ^ _21250_ /*62904*/;
assign _21255_ = _21246_ & _21254_ /*62902*/;
assign _21025_ = _21246_ ^ _21254_ /*62903*/;
assign _21252_ = _21253_ | _21255_ /*62900*/;
assign _21257_ = ~Q[40] /*62899*/;
assign _21256_ = _21257_ & D[33] /*62898*/;
assign _21259_ = _20578_ & _21256_ /*62893*/;
assign _21260_ = _20578_ ^ _21256_ /*62896*/;
assign _21261_ = _21252_ & _21260_ /*62894*/;
assign _21026_ = _21252_ ^ _21260_ /*62895*/;
assign _21258_ = _21259_ | _21261_ /*62892*/;
assign _21263_ = ~Q[40] /*62891*/;
assign _21262_ = _21263_ & D[34] /*62890*/;
assign _21265_ = _20579_ & _21262_ /*62885*/;
assign _21266_ = _20579_ ^ _21262_ /*62888*/;
assign _21267_ = _21258_ & _21266_ /*62886*/;
assign _21027_ = _21258_ ^ _21266_ /*62887*/;
assign _21264_ = _21265_ | _21267_ /*62884*/;
assign _21269_ = ~Q[40] /*62883*/;
assign _21268_ = _21269_ & D[35] /*62882*/;
assign _21271_ = _20580_ & _21268_ /*62877*/;
assign _21272_ = _20580_ ^ _21268_ /*62880*/;
assign _21273_ = _21264_ & _21272_ /*62878*/;
assign _21028_ = _21264_ ^ _21272_ /*62879*/;
assign _21270_ = _21271_ | _21273_ /*62876*/;
assign _21275_ = ~Q[40] /*62875*/;
assign _21274_ = _21275_ & D[36] /*62874*/;
assign _21277_ = _20581_ & _21274_ /*62869*/;
assign _21278_ = _20581_ ^ _21274_ /*62872*/;
assign _21279_ = _21270_ & _21278_ /*62870*/;
assign _21029_ = _21270_ ^ _21278_ /*62871*/;
assign _21276_ = _21277_ | _21279_ /*62868*/;
assign _21281_ = ~Q[40] /*62867*/;
assign _21280_ = _21281_ & D[37] /*62866*/;
assign _21283_ = _20582_ & _21280_ /*62861*/;
assign _21284_ = _20582_ ^ _21280_ /*62864*/;
assign _21285_ = _21276_ & _21284_ /*62862*/;
assign _21030_ = _21276_ ^ _21284_ /*62863*/;
assign _21282_ = _21283_ | _21285_ /*62860*/;
assign _21287_ = ~Q[40] /*62859*/;
assign _21286_ = _21287_ & D[38] /*62858*/;
assign _21289_ = _20583_ & _21286_ /*62853*/;
assign _21290_ = _20583_ ^ _21286_ /*62856*/;
assign _21291_ = _21282_ & _21290_ /*62854*/;
assign _21031_ = _21282_ ^ _21290_ /*62855*/;
assign _21288_ = _21289_ | _21291_ /*62852*/;
assign _21293_ = ~Q[40] /*62851*/;
assign _21292_ = _21293_ & D[39] /*62850*/;
assign _21295_ = _20584_ & _21292_ /*62845*/;
assign _21296_ = _20584_ ^ _21292_ /*62848*/;
assign _21297_ = _21288_ & _21296_ /*62846*/;
assign _21032_ = _21288_ ^ _21296_ /*62847*/;
assign _21294_ = _21295_ | _21297_ /*62844*/;
assign _21299_ = ~Q[40] /*62843*/;
assign _21298_ = _21299_ & D[40] /*62842*/;
assign _21301_ = _20585_ & _21298_ /*62837*/;
assign _21302_ = _20585_ ^ _21298_ /*62840*/;
assign _21303_ = _21294_ & _21302_ /*62838*/;
assign _21033_ = _21294_ ^ _21302_ /*62839*/;
assign _21300_ = _21301_ | _21303_ /*62836*/;
assign _21305_ = ~Q[40] /*62835*/;
assign _21304_ = _21305_ & D[41] /*62834*/;
assign _21307_ = _20586_ & _21304_ /*62829*/;
assign _21308_ = _20586_ ^ _21304_ /*62832*/;
assign _21309_ = _21300_ & _21308_ /*62830*/;
assign _21034_ = _21300_ ^ _21308_ /*62831*/;
assign _21306_ = _21307_ | _21309_ /*62828*/;
assign _21311_ = ~Q[40] /*62827*/;
assign _21310_ = _21311_ & D[42] /*62826*/;
assign _21313_ = _20587_ & _21310_ /*62821*/;
assign _21314_ = _20587_ ^ _21310_ /*62824*/;
assign _21315_ = _21306_ & _21314_ /*62822*/;
assign _21035_ = _21306_ ^ _21314_ /*62823*/;
assign _21312_ = _21313_ | _21315_ /*62820*/;
assign _21317_ = ~Q[40] /*62819*/;
assign _21316_ = _21317_ & D[43] /*62818*/;
assign _21319_ = _20588_ & _21316_ /*62813*/;
assign _21320_ = _20588_ ^ _21316_ /*62816*/;
assign _21321_ = _21312_ & _21320_ /*62814*/;
assign _21036_ = _21312_ ^ _21320_ /*62815*/;
assign _21318_ = _21319_ | _21321_ /*62812*/;
assign _21323_ = ~Q[40] /*62811*/;
assign _21322_ = _21323_ & D[44] /*62810*/;
assign _21325_ = _20589_ & _21322_ /*62805*/;
assign _21326_ = _20589_ ^ _21322_ /*62808*/;
assign _21327_ = _21318_ & _21326_ /*62806*/;
assign _21037_ = _21318_ ^ _21326_ /*62807*/;
assign _21324_ = _21325_ | _21327_ /*62804*/;
assign _21329_ = ~Q[40] /*62803*/;
assign _21328_ = _21329_ & D[45] /*62802*/;
assign _21331_ = _20590_ & _21328_ /*62797*/;
assign _21332_ = _20590_ ^ _21328_ /*62800*/;
assign _21333_ = _21324_ & _21332_ /*62798*/;
assign _21038_ = _21324_ ^ _21332_ /*62799*/;
assign _21330_ = _21331_ | _21333_ /*62796*/;
assign _21335_ = ~Q[40] /*62795*/;
assign _21334_ = _21335_ & D[46] /*62794*/;
assign _21337_ = _20591_ & _21334_ /*62789*/;
assign _21338_ = _20591_ ^ _21334_ /*62792*/;
assign _21339_ = _21330_ & _21338_ /*62790*/;
assign _21039_ = _21330_ ^ _21338_ /*62791*/;
assign _21336_ = _21337_ | _21339_ /*62788*/;
assign _21341_ = ~Q[40] /*62787*/;
assign _21340_ = _21341_ & D[47] /*62786*/;
assign _21343_ = _20592_ & _21340_ /*62781*/;
assign _21344_ = _20592_ ^ _21340_ /*62784*/;
assign _21345_ = _21336_ & _21344_ /*62782*/;
assign _21040_ = _21336_ ^ _21344_ /*62783*/;
assign _21342_ = _21343_ | _21345_ /*62780*/;
assign _21347_ = ~Q[40] /*62779*/;
assign _21346_ = _21347_ & D[48] /*62778*/;
assign _21349_ = _20593_ & _21346_ /*62773*/;
assign _21350_ = _20593_ ^ _21346_ /*62776*/;
assign _21351_ = _21342_ & _21350_ /*62774*/;
assign _21041_ = _21342_ ^ _21350_ /*62775*/;
assign _21348_ = _21349_ | _21351_ /*62772*/;
assign _21353_ = ~Q[40] /*62771*/;
assign _21352_ = _21353_ & D[49] /*62770*/;
assign _21355_ = _20594_ & _21352_ /*62765*/;
assign _21356_ = _20594_ ^ _21352_ /*62768*/;
assign _21357_ = _21348_ & _21356_ /*62766*/;
assign _21042_ = _21348_ ^ _21356_ /*62767*/;
assign _21354_ = _21355_ | _21357_ /*62764*/;
assign _21359_ = ~Q[40] /*62763*/;
assign _21358_ = _21359_ & D[50] /*62762*/;
assign _21361_ = _20595_ & _21358_ /*62757*/;
assign _21362_ = _20595_ ^ _21358_ /*62760*/;
assign _21363_ = _21354_ & _21362_ /*62758*/;
assign _21043_ = _21354_ ^ _21362_ /*62759*/;
assign _21360_ = _21361_ | _21363_ /*62756*/;
assign _21365_ = ~Q[40] /*62755*/;
assign _21364_ = _21365_ & D[51] /*62754*/;
assign _21367_ = _20596_ & _21364_ /*62749*/;
assign _21368_ = _20596_ ^ _21364_ /*62752*/;
assign _21369_ = _21360_ & _21368_ /*62750*/;
assign _21044_ = _21360_ ^ _21368_ /*62751*/;
assign _21366_ = _21367_ | _21369_ /*62748*/;
assign _21371_ = ~Q[40] /*62747*/;
assign _21370_ = _21371_ & D[52] /*62746*/;
assign _21373_ = _20597_ & _21370_ /*62741*/;
assign _21374_ = _20597_ ^ _21370_ /*62744*/;
assign _21375_ = _21366_ & _21374_ /*62742*/;
assign _21045_ = _21366_ ^ _21374_ /*62743*/;
assign _21372_ = _21373_ | _21375_ /*62740*/;
assign _21377_ = ~Q[40] /*62739*/;
assign _21376_ = _21377_ & D[53] /*62738*/;
assign _21379_ = _20598_ & _21376_ /*62733*/;
assign _21380_ = _20598_ ^ _21376_ /*62736*/;
assign _21381_ = _21372_ & _21380_ /*62734*/;
assign _21046_ = _21372_ ^ _21380_ /*62735*/;
assign _21378_ = _21379_ | _21381_ /*62732*/;
assign _21383_ = ~Q[40] /*62731*/;
assign _21382_ = _21383_ & D[54] /*62730*/;
assign _21385_ = _20599_ & _21382_ /*62725*/;
assign _21386_ = _20599_ ^ _21382_ /*62728*/;
assign _21387_ = _21378_ & _21386_ /*62726*/;
assign _21047_ = _21378_ ^ _21386_ /*62727*/;
assign _21384_ = _21385_ | _21387_ /*62724*/;
assign _21389_ = ~Q[40] /*62723*/;
assign _21388_ = _21389_ & D[55] /*62722*/;
assign _21391_ = _20600_ & _21388_ /*62717*/;
assign _21392_ = _20600_ ^ _21388_ /*62720*/;
assign _21393_ = _21384_ & _21392_ /*62718*/;
assign _21048_ = _21384_ ^ _21392_ /*62719*/;
assign _21390_ = _21391_ | _21393_ /*62716*/;
assign _21395_ = ~Q[40] /*62715*/;
assign _21394_ = _21395_ & D[56] /*62714*/;
assign _21397_ = _20601_ & _21394_ /*62709*/;
assign _21398_ = _20601_ ^ _21394_ /*62712*/;
assign _21399_ = _21390_ & _21398_ /*62710*/;
assign _21049_ = _21390_ ^ _21398_ /*62711*/;
assign _21396_ = _21397_ | _21399_ /*62708*/;
assign _21401_ = ~Q[40] /*62707*/;
assign _21400_ = _21401_ & D[57] /*62706*/;
assign _21403_ = _20602_ & _21400_ /*62701*/;
assign _21404_ = _20602_ ^ _21400_ /*62704*/;
assign _21405_ = _21396_ & _21404_ /*62702*/;
assign _21050_ = _21396_ ^ _21404_ /*62703*/;
assign _21402_ = _21403_ | _21405_ /*62700*/;
assign _21407_ = ~Q[40] /*62699*/;
assign _21406_ = _21407_ & D[58] /*62698*/;
assign _21409_ = _20603_ & _21406_ /*62693*/;
assign _21410_ = _20603_ ^ _21406_ /*62696*/;
assign _21411_ = _21402_ & _21410_ /*62694*/;
assign _21051_ = _21402_ ^ _21410_ /*62695*/;
assign _21408_ = _21409_ | _21411_ /*62692*/;
assign _21413_ = ~Q[40] /*62691*/;
assign _21412_ = _21413_ & D[59] /*62690*/;
assign _21415_ = _20604_ & _21412_ /*62685*/;
assign _21416_ = _20604_ ^ _21412_ /*62688*/;
assign _21417_ = _21408_ & _21416_ /*62686*/;
assign _21052_ = _21408_ ^ _21416_ /*62687*/;
assign _21414_ = _21415_ | _21417_ /*62684*/;
assign _21419_ = ~Q[40] /*62683*/;
assign _21418_ = _21419_ & D[60] /*62682*/;
assign _21421_ = _20605_ & _21418_ /*62677*/;
assign _21422_ = _20605_ ^ _21418_ /*62680*/;
assign _21423_ = _21414_ & _21422_ /*62678*/;
assign _21053_ = _21414_ ^ _21422_ /*62679*/;
assign _21420_ = _21421_ | _21423_ /*62676*/;
assign _21425_ = ~Q[40] /*62675*/;
assign _21424_ = _21425_ & D[61] /*62674*/;
assign _21427_ = _20606_ & _21424_ /*62669*/;
assign _21428_ = _20606_ ^ _21424_ /*62672*/;
assign _21429_ = _21420_ & _21428_ /*62670*/;
assign _21054_ = _21420_ ^ _21428_ /*62671*/;
assign _21426_ = _21427_ | _21429_ /*62668*/;
assign _21431_ = ~Q[40] /*62667*/;
assign _21430_ = _21431_ & D[62] /*62666*/;
assign _21433_ = _20607_ & _21430_ /*62661*/;
assign _21434_ = _20607_ ^ _21430_ /*62664*/;
assign _21435_ = _21426_ & _21434_ /*62662*/;
assign _21055_ = _21426_ ^ _21434_ /*62663*/;
assign _21432_ = _21433_ | _21435_ /*62660*/;
assign _21437_ = ~Q[40] /*62659*/;
assign _21436_ = _21437_ & zeroWire /*62658*/;
assign _21438_ = _20608_ ^ _21436_ /*62656*/;
assign _21056_ = _21438_ ^ _21432_ /*62655*/;
assign _21509_ = ~D[0] /*62401*/;
assign _21506_ = R_0[39] & _21509_ /*62397*/;
assign _21507_ = R_0[39] ^ _21509_ /*62400*/;
assign _21508_ = oneWire & _21507_ /*62398*/;
assign _21441_ = oneWire ^ _21507_ /*62399*/;
assign _21505_ = _21506_ | _21508_ /*62396*/;
assign _21514_ = ~D[1] /*62395*/;
assign _21511_ = _20993_ & _21514_ /*62391*/;
assign _21512_ = _20993_ ^ _21514_ /*62394*/;
assign _21513_ = _21505_ & _21512_ /*62392*/;
assign _21442_ = _21505_ ^ _21512_ /*62393*/;
assign _21510_ = _21511_ | _21513_ /*62390*/;
assign _21519_ = ~D[2] /*62389*/;
assign _21516_ = _20994_ & _21519_ /*62385*/;
assign _21517_ = _20994_ ^ _21519_ /*62388*/;
assign _21518_ = _21510_ & _21517_ /*62386*/;
assign _21443_ = _21510_ ^ _21517_ /*62387*/;
assign _21515_ = _21516_ | _21518_ /*62384*/;
assign _21524_ = ~D[3] /*62383*/;
assign _21521_ = _20995_ & _21524_ /*62379*/;
assign _21522_ = _20995_ ^ _21524_ /*62382*/;
assign _21523_ = _21515_ & _21522_ /*62380*/;
assign _21444_ = _21515_ ^ _21522_ /*62381*/;
assign _21520_ = _21521_ | _21523_ /*62378*/;
assign _21529_ = ~D[4] /*62377*/;
assign _21526_ = _20996_ & _21529_ /*62373*/;
assign _21527_ = _20996_ ^ _21529_ /*62376*/;
assign _21528_ = _21520_ & _21527_ /*62374*/;
assign _21445_ = _21520_ ^ _21527_ /*62375*/;
assign _21525_ = _21526_ | _21528_ /*62372*/;
assign _21534_ = ~D[5] /*62371*/;
assign _21531_ = _20997_ & _21534_ /*62367*/;
assign _21532_ = _20997_ ^ _21534_ /*62370*/;
assign _21533_ = _21525_ & _21532_ /*62368*/;
assign _21446_ = _21525_ ^ _21532_ /*62369*/;
assign _21530_ = _21531_ | _21533_ /*62366*/;
assign _21539_ = ~D[6] /*62365*/;
assign _21536_ = _20998_ & _21539_ /*62361*/;
assign _21537_ = _20998_ ^ _21539_ /*62364*/;
assign _21538_ = _21530_ & _21537_ /*62362*/;
assign _21447_ = _21530_ ^ _21537_ /*62363*/;
assign _21535_ = _21536_ | _21538_ /*62360*/;
assign _21544_ = ~D[7] /*62359*/;
assign _21541_ = _20999_ & _21544_ /*62355*/;
assign _21542_ = _20999_ ^ _21544_ /*62358*/;
assign _21543_ = _21535_ & _21542_ /*62356*/;
assign _21448_ = _21535_ ^ _21542_ /*62357*/;
assign _21540_ = _21541_ | _21543_ /*62354*/;
assign _21549_ = ~D[8] /*62353*/;
assign _21546_ = _21000_ & _21549_ /*62349*/;
assign _21547_ = _21000_ ^ _21549_ /*62352*/;
assign _21548_ = _21540_ & _21547_ /*62350*/;
assign _21449_ = _21540_ ^ _21547_ /*62351*/;
assign _21545_ = _21546_ | _21548_ /*62348*/;
assign _21554_ = ~D[9] /*62347*/;
assign _21551_ = _21001_ & _21554_ /*62343*/;
assign _21552_ = _21001_ ^ _21554_ /*62346*/;
assign _21553_ = _21545_ & _21552_ /*62344*/;
assign _21450_ = _21545_ ^ _21552_ /*62345*/;
assign _21550_ = _21551_ | _21553_ /*62342*/;
assign _21559_ = ~D[10] /*62341*/;
assign _21556_ = _21002_ & _21559_ /*62337*/;
assign _21557_ = _21002_ ^ _21559_ /*62340*/;
assign _21558_ = _21550_ & _21557_ /*62338*/;
assign _21451_ = _21550_ ^ _21557_ /*62339*/;
assign _21555_ = _21556_ | _21558_ /*62336*/;
assign _21564_ = ~D[11] /*62335*/;
assign _21561_ = _21003_ & _21564_ /*62331*/;
assign _21562_ = _21003_ ^ _21564_ /*62334*/;
assign _21563_ = _21555_ & _21562_ /*62332*/;
assign _21452_ = _21555_ ^ _21562_ /*62333*/;
assign _21560_ = _21561_ | _21563_ /*62330*/;
assign _21569_ = ~D[12] /*62329*/;
assign _21566_ = _21004_ & _21569_ /*62325*/;
assign _21567_ = _21004_ ^ _21569_ /*62328*/;
assign _21568_ = _21560_ & _21567_ /*62326*/;
assign _21453_ = _21560_ ^ _21567_ /*62327*/;
assign _21565_ = _21566_ | _21568_ /*62324*/;
assign _21574_ = ~D[13] /*62323*/;
assign _21571_ = _21005_ & _21574_ /*62319*/;
assign _21572_ = _21005_ ^ _21574_ /*62322*/;
assign _21573_ = _21565_ & _21572_ /*62320*/;
assign _21454_ = _21565_ ^ _21572_ /*62321*/;
assign _21570_ = _21571_ | _21573_ /*62318*/;
assign _21579_ = ~D[14] /*62317*/;
assign _21576_ = _21006_ & _21579_ /*62313*/;
assign _21577_ = _21006_ ^ _21579_ /*62316*/;
assign _21578_ = _21570_ & _21577_ /*62314*/;
assign _21455_ = _21570_ ^ _21577_ /*62315*/;
assign _21575_ = _21576_ | _21578_ /*62312*/;
assign _21584_ = ~D[15] /*62311*/;
assign _21581_ = _21007_ & _21584_ /*62307*/;
assign _21582_ = _21007_ ^ _21584_ /*62310*/;
assign _21583_ = _21575_ & _21582_ /*62308*/;
assign _21456_ = _21575_ ^ _21582_ /*62309*/;
assign _21580_ = _21581_ | _21583_ /*62306*/;
assign _21589_ = ~D[16] /*62305*/;
assign _21586_ = _21008_ & _21589_ /*62301*/;
assign _21587_ = _21008_ ^ _21589_ /*62304*/;
assign _21588_ = _21580_ & _21587_ /*62302*/;
assign _21457_ = _21580_ ^ _21587_ /*62303*/;
assign _21585_ = _21586_ | _21588_ /*62300*/;
assign _21594_ = ~D[17] /*62299*/;
assign _21591_ = _21009_ & _21594_ /*62295*/;
assign _21592_ = _21009_ ^ _21594_ /*62298*/;
assign _21593_ = _21585_ & _21592_ /*62296*/;
assign _21458_ = _21585_ ^ _21592_ /*62297*/;
assign _21590_ = _21591_ | _21593_ /*62294*/;
assign _21599_ = ~D[18] /*62293*/;
assign _21596_ = _21010_ & _21599_ /*62289*/;
assign _21597_ = _21010_ ^ _21599_ /*62292*/;
assign _21598_ = _21590_ & _21597_ /*62290*/;
assign _21459_ = _21590_ ^ _21597_ /*62291*/;
assign _21595_ = _21596_ | _21598_ /*62288*/;
assign _21604_ = ~D[19] /*62287*/;
assign _21601_ = _21011_ & _21604_ /*62283*/;
assign _21602_ = _21011_ ^ _21604_ /*62286*/;
assign _21603_ = _21595_ & _21602_ /*62284*/;
assign _21460_ = _21595_ ^ _21602_ /*62285*/;
assign _21600_ = _21601_ | _21603_ /*62282*/;
assign _21609_ = ~D[20] /*62281*/;
assign _21606_ = _21012_ & _21609_ /*62277*/;
assign _21607_ = _21012_ ^ _21609_ /*62280*/;
assign _21608_ = _21600_ & _21607_ /*62278*/;
assign _21461_ = _21600_ ^ _21607_ /*62279*/;
assign _21605_ = _21606_ | _21608_ /*62276*/;
assign _21614_ = ~D[21] /*62275*/;
assign _21611_ = _21013_ & _21614_ /*62271*/;
assign _21612_ = _21013_ ^ _21614_ /*62274*/;
assign _21613_ = _21605_ & _21612_ /*62272*/;
assign _21462_ = _21605_ ^ _21612_ /*62273*/;
assign _21610_ = _21611_ | _21613_ /*62270*/;
assign _21619_ = ~D[22] /*62269*/;
assign _21616_ = _21014_ & _21619_ /*62265*/;
assign _21617_ = _21014_ ^ _21619_ /*62268*/;
assign _21618_ = _21610_ & _21617_ /*62266*/;
assign _21463_ = _21610_ ^ _21617_ /*62267*/;
assign _21615_ = _21616_ | _21618_ /*62264*/;
assign _21624_ = ~D[23] /*62263*/;
assign _21621_ = _21015_ & _21624_ /*62259*/;
assign _21622_ = _21015_ ^ _21624_ /*62262*/;
assign _21623_ = _21615_ & _21622_ /*62260*/;
assign _21464_ = _21615_ ^ _21622_ /*62261*/;
assign _21620_ = _21621_ | _21623_ /*62258*/;
assign _21629_ = ~D[24] /*62257*/;
assign _21626_ = _21016_ & _21629_ /*62253*/;
assign _21627_ = _21016_ ^ _21629_ /*62256*/;
assign _21628_ = _21620_ & _21627_ /*62254*/;
assign _21465_ = _21620_ ^ _21627_ /*62255*/;
assign _21625_ = _21626_ | _21628_ /*62252*/;
assign _21634_ = ~D[25] /*62251*/;
assign _21631_ = _21017_ & _21634_ /*62247*/;
assign _21632_ = _21017_ ^ _21634_ /*62250*/;
assign _21633_ = _21625_ & _21632_ /*62248*/;
assign _21466_ = _21625_ ^ _21632_ /*62249*/;
assign _21630_ = _21631_ | _21633_ /*62246*/;
assign _21639_ = ~D[26] /*62245*/;
assign _21636_ = _21018_ & _21639_ /*62241*/;
assign _21637_ = _21018_ ^ _21639_ /*62244*/;
assign _21638_ = _21630_ & _21637_ /*62242*/;
assign _21467_ = _21630_ ^ _21637_ /*62243*/;
assign _21635_ = _21636_ | _21638_ /*62240*/;
assign _21644_ = ~D[27] /*62239*/;
assign _21641_ = _21019_ & _21644_ /*62235*/;
assign _21642_ = _21019_ ^ _21644_ /*62238*/;
assign _21643_ = _21635_ & _21642_ /*62236*/;
assign _21468_ = _21635_ ^ _21642_ /*62237*/;
assign _21640_ = _21641_ | _21643_ /*62234*/;
assign _21649_ = ~D[28] /*62233*/;
assign _21646_ = _21020_ & _21649_ /*62229*/;
assign _21647_ = _21020_ ^ _21649_ /*62232*/;
assign _21648_ = _21640_ & _21647_ /*62230*/;
assign _21469_ = _21640_ ^ _21647_ /*62231*/;
assign _21645_ = _21646_ | _21648_ /*62228*/;
assign _21654_ = ~D[29] /*62227*/;
assign _21651_ = _21021_ & _21654_ /*62223*/;
assign _21652_ = _21021_ ^ _21654_ /*62226*/;
assign _21653_ = _21645_ & _21652_ /*62224*/;
assign _21470_ = _21645_ ^ _21652_ /*62225*/;
assign _21650_ = _21651_ | _21653_ /*62222*/;
assign _21659_ = ~D[30] /*62221*/;
assign _21656_ = _21022_ & _21659_ /*62217*/;
assign _21657_ = _21022_ ^ _21659_ /*62220*/;
assign _21658_ = _21650_ & _21657_ /*62218*/;
assign _21471_ = _21650_ ^ _21657_ /*62219*/;
assign _21655_ = _21656_ | _21658_ /*62216*/;
assign _21664_ = ~D[31] /*62215*/;
assign _21661_ = _21023_ & _21664_ /*62211*/;
assign _21662_ = _21023_ ^ _21664_ /*62214*/;
assign _21663_ = _21655_ & _21662_ /*62212*/;
assign _21472_ = _21655_ ^ _21662_ /*62213*/;
assign _21660_ = _21661_ | _21663_ /*62210*/;
assign _21669_ = ~D[32] /*62209*/;
assign _21666_ = _21024_ & _21669_ /*62205*/;
assign _21667_ = _21024_ ^ _21669_ /*62208*/;
assign _21668_ = _21660_ & _21667_ /*62206*/;
assign _21473_ = _21660_ ^ _21667_ /*62207*/;
assign _21665_ = _21666_ | _21668_ /*62204*/;
assign _21674_ = ~D[33] /*62203*/;
assign _21671_ = _21025_ & _21674_ /*62199*/;
assign _21672_ = _21025_ ^ _21674_ /*62202*/;
assign _21673_ = _21665_ & _21672_ /*62200*/;
assign _21474_ = _21665_ ^ _21672_ /*62201*/;
assign _21670_ = _21671_ | _21673_ /*62198*/;
assign _21679_ = ~D[34] /*62197*/;
assign _21676_ = _21026_ & _21679_ /*62193*/;
assign _21677_ = _21026_ ^ _21679_ /*62196*/;
assign _21678_ = _21670_ & _21677_ /*62194*/;
assign _21475_ = _21670_ ^ _21677_ /*62195*/;
assign _21675_ = _21676_ | _21678_ /*62192*/;
assign _21684_ = ~D[35] /*62191*/;
assign _21681_ = _21027_ & _21684_ /*62187*/;
assign _21682_ = _21027_ ^ _21684_ /*62190*/;
assign _21683_ = _21675_ & _21682_ /*62188*/;
assign _21476_ = _21675_ ^ _21682_ /*62189*/;
assign _21680_ = _21681_ | _21683_ /*62186*/;
assign _21689_ = ~D[36] /*62185*/;
assign _21686_ = _21028_ & _21689_ /*62181*/;
assign _21687_ = _21028_ ^ _21689_ /*62184*/;
assign _21688_ = _21680_ & _21687_ /*62182*/;
assign _21477_ = _21680_ ^ _21687_ /*62183*/;
assign _21685_ = _21686_ | _21688_ /*62180*/;
assign _21694_ = ~D[37] /*62179*/;
assign _21691_ = _21029_ & _21694_ /*62175*/;
assign _21692_ = _21029_ ^ _21694_ /*62178*/;
assign _21693_ = _21685_ & _21692_ /*62176*/;
assign _21478_ = _21685_ ^ _21692_ /*62177*/;
assign _21690_ = _21691_ | _21693_ /*62174*/;
assign _21699_ = ~D[38] /*62173*/;
assign _21696_ = _21030_ & _21699_ /*62169*/;
assign _21697_ = _21030_ ^ _21699_ /*62172*/;
assign _21698_ = _21690_ & _21697_ /*62170*/;
assign _21479_ = _21690_ ^ _21697_ /*62171*/;
assign _21695_ = _21696_ | _21698_ /*62168*/;
assign _21704_ = ~D[39] /*62167*/;
assign _21701_ = _21031_ & _21704_ /*62163*/;
assign _21702_ = _21031_ ^ _21704_ /*62166*/;
assign _21703_ = _21695_ & _21702_ /*62164*/;
assign _21480_ = _21695_ ^ _21702_ /*62165*/;
assign _21700_ = _21701_ | _21703_ /*62162*/;
assign _21709_ = ~D[40] /*62161*/;
assign _21706_ = _21032_ & _21709_ /*62157*/;
assign _21707_ = _21032_ ^ _21709_ /*62160*/;
assign _21708_ = _21700_ & _21707_ /*62158*/;
assign _21481_ = _21700_ ^ _21707_ /*62159*/;
assign _21705_ = _21706_ | _21708_ /*62156*/;
assign _21714_ = ~D[41] /*62155*/;
assign _21711_ = _21033_ & _21714_ /*62151*/;
assign _21712_ = _21033_ ^ _21714_ /*62154*/;
assign _21713_ = _21705_ & _21712_ /*62152*/;
assign _21482_ = _21705_ ^ _21712_ /*62153*/;
assign _21710_ = _21711_ | _21713_ /*62150*/;
assign _21719_ = ~D[42] /*62149*/;
assign _21716_ = _21034_ & _21719_ /*62145*/;
assign _21717_ = _21034_ ^ _21719_ /*62148*/;
assign _21718_ = _21710_ & _21717_ /*62146*/;
assign _21483_ = _21710_ ^ _21717_ /*62147*/;
assign _21715_ = _21716_ | _21718_ /*62144*/;
assign _21724_ = ~D[43] /*62143*/;
assign _21721_ = _21035_ & _21724_ /*62139*/;
assign _21722_ = _21035_ ^ _21724_ /*62142*/;
assign _21723_ = _21715_ & _21722_ /*62140*/;
assign _21484_ = _21715_ ^ _21722_ /*62141*/;
assign _21720_ = _21721_ | _21723_ /*62138*/;
assign _21729_ = ~D[44] /*62137*/;
assign _21726_ = _21036_ & _21729_ /*62133*/;
assign _21727_ = _21036_ ^ _21729_ /*62136*/;
assign _21728_ = _21720_ & _21727_ /*62134*/;
assign _21485_ = _21720_ ^ _21727_ /*62135*/;
assign _21725_ = _21726_ | _21728_ /*62132*/;
assign _21734_ = ~D[45] /*62131*/;
assign _21731_ = _21037_ & _21734_ /*62127*/;
assign _21732_ = _21037_ ^ _21734_ /*62130*/;
assign _21733_ = _21725_ & _21732_ /*62128*/;
assign _21486_ = _21725_ ^ _21732_ /*62129*/;
assign _21730_ = _21731_ | _21733_ /*62126*/;
assign _21739_ = ~D[46] /*62125*/;
assign _21736_ = _21038_ & _21739_ /*62121*/;
assign _21737_ = _21038_ ^ _21739_ /*62124*/;
assign _21738_ = _21730_ & _21737_ /*62122*/;
assign _21487_ = _21730_ ^ _21737_ /*62123*/;
assign _21735_ = _21736_ | _21738_ /*62120*/;
assign _21744_ = ~D[47] /*62119*/;
assign _21741_ = _21039_ & _21744_ /*62115*/;
assign _21742_ = _21039_ ^ _21744_ /*62118*/;
assign _21743_ = _21735_ & _21742_ /*62116*/;
assign _21488_ = _21735_ ^ _21742_ /*62117*/;
assign _21740_ = _21741_ | _21743_ /*62114*/;
assign _21749_ = ~D[48] /*62113*/;
assign _21746_ = _21040_ & _21749_ /*62109*/;
assign _21747_ = _21040_ ^ _21749_ /*62112*/;
assign _21748_ = _21740_ & _21747_ /*62110*/;
assign _21489_ = _21740_ ^ _21747_ /*62111*/;
assign _21745_ = _21746_ | _21748_ /*62108*/;
assign _21754_ = ~D[49] /*62107*/;
assign _21751_ = _21041_ & _21754_ /*62103*/;
assign _21752_ = _21041_ ^ _21754_ /*62106*/;
assign _21753_ = _21745_ & _21752_ /*62104*/;
assign _21490_ = _21745_ ^ _21752_ /*62105*/;
assign _21750_ = _21751_ | _21753_ /*62102*/;
assign _21759_ = ~D[50] /*62101*/;
assign _21756_ = _21042_ & _21759_ /*62097*/;
assign _21757_ = _21042_ ^ _21759_ /*62100*/;
assign _21758_ = _21750_ & _21757_ /*62098*/;
assign _21491_ = _21750_ ^ _21757_ /*62099*/;
assign _21755_ = _21756_ | _21758_ /*62096*/;
assign _21764_ = ~D[51] /*62095*/;
assign _21761_ = _21043_ & _21764_ /*62091*/;
assign _21762_ = _21043_ ^ _21764_ /*62094*/;
assign _21763_ = _21755_ & _21762_ /*62092*/;
assign _21492_ = _21755_ ^ _21762_ /*62093*/;
assign _21760_ = _21761_ | _21763_ /*62090*/;
assign _21769_ = ~D[52] /*62089*/;
assign _21766_ = _21044_ & _21769_ /*62085*/;
assign _21767_ = _21044_ ^ _21769_ /*62088*/;
assign _21768_ = _21760_ & _21767_ /*62086*/;
assign _21493_ = _21760_ ^ _21767_ /*62087*/;
assign _21765_ = _21766_ | _21768_ /*62084*/;
assign _21774_ = ~D[53] /*62083*/;
assign _21771_ = _21045_ & _21774_ /*62079*/;
assign _21772_ = _21045_ ^ _21774_ /*62082*/;
assign _21773_ = _21765_ & _21772_ /*62080*/;
assign _21494_ = _21765_ ^ _21772_ /*62081*/;
assign _21770_ = _21771_ | _21773_ /*62078*/;
assign _21779_ = ~D[54] /*62077*/;
assign _21776_ = _21046_ & _21779_ /*62073*/;
assign _21777_ = _21046_ ^ _21779_ /*62076*/;
assign _21778_ = _21770_ & _21777_ /*62074*/;
assign _21495_ = _21770_ ^ _21777_ /*62075*/;
assign _21775_ = _21776_ | _21778_ /*62072*/;
assign _21784_ = ~D[55] /*62071*/;
assign _21781_ = _21047_ & _21784_ /*62067*/;
assign _21782_ = _21047_ ^ _21784_ /*62070*/;
assign _21783_ = _21775_ & _21782_ /*62068*/;
assign _21496_ = _21775_ ^ _21782_ /*62069*/;
assign _21780_ = _21781_ | _21783_ /*62066*/;
assign _21789_ = ~D[56] /*62065*/;
assign _21786_ = _21048_ & _21789_ /*62061*/;
assign _21787_ = _21048_ ^ _21789_ /*62064*/;
assign _21788_ = _21780_ & _21787_ /*62062*/;
assign _21497_ = _21780_ ^ _21787_ /*62063*/;
assign _21785_ = _21786_ | _21788_ /*62060*/;
assign _21794_ = ~D[57] /*62059*/;
assign _21791_ = _21049_ & _21794_ /*62055*/;
assign _21792_ = _21049_ ^ _21794_ /*62058*/;
assign _21793_ = _21785_ & _21792_ /*62056*/;
assign _21498_ = _21785_ ^ _21792_ /*62057*/;
assign _21790_ = _21791_ | _21793_ /*62054*/;
assign _21799_ = ~D[58] /*62053*/;
assign _21796_ = _21050_ & _21799_ /*62049*/;
assign _21797_ = _21050_ ^ _21799_ /*62052*/;
assign _21798_ = _21790_ & _21797_ /*62050*/;
assign _21499_ = _21790_ ^ _21797_ /*62051*/;
assign _21795_ = _21796_ | _21798_ /*62048*/;
assign _21804_ = ~D[59] /*62047*/;
assign _21801_ = _21051_ & _21804_ /*62043*/;
assign _21802_ = _21051_ ^ _21804_ /*62046*/;
assign _21803_ = _21795_ & _21802_ /*62044*/;
assign _21500_ = _21795_ ^ _21802_ /*62045*/;
assign _21800_ = _21801_ | _21803_ /*62042*/;
assign _21809_ = ~D[60] /*62041*/;
assign _21806_ = _21052_ & _21809_ /*62037*/;
assign _21807_ = _21052_ ^ _21809_ /*62040*/;
assign _21808_ = _21800_ & _21807_ /*62038*/;
assign _21501_ = _21800_ ^ _21807_ /*62039*/;
assign _21805_ = _21806_ | _21808_ /*62036*/;
assign _21814_ = ~D[61] /*62035*/;
assign _21811_ = _21053_ & _21814_ /*62031*/;
assign _21812_ = _21053_ ^ _21814_ /*62034*/;
assign _21813_ = _21805_ & _21812_ /*62032*/;
assign _21502_ = _21805_ ^ _21812_ /*62033*/;
assign _21810_ = _21811_ | _21813_ /*62030*/;
assign _21819_ = ~D[62] /*62029*/;
assign _21816_ = _21054_ & _21819_ /*62025*/;
assign _21817_ = _21054_ ^ _21819_ /*62028*/;
assign _21818_ = _21810_ & _21817_ /*62026*/;
assign _21503_ = _21810_ ^ _21817_ /*62027*/;
assign _21815_ = _21816_ | _21818_ /*62024*/;
assign _21820_ = _21055_ & oneWire /*62019*/;
assign _21821_ = _21055_ ^ oneWire /*62022*/;
assign _21822_ = _21815_ & _21821_ /*62020*/;
assign _21504_ = _21815_ ^ _21821_ /*62021*/;
assign Q[39] = _21820_ | _21822_ /*62018*/;
assign _21955_ = ~Q[39] /*61633*/;
assign _21954_ = _21955_ & D[0] /*61632*/;
assign _21957_ = _21441_ & _21954_ /*61627*/;
assign _21958_ = _21441_ ^ _21954_ /*61630*/;
assign _21959_ = zeroWire & _21958_ /*61628*/;
assign _21889_ = zeroWire ^ _21958_ /*61629*/;
assign _21956_ = _21957_ | _21959_ /*61626*/;
assign _21961_ = ~Q[39] /*61625*/;
assign _21960_ = _21961_ & D[1] /*61624*/;
assign _21963_ = _21442_ & _21960_ /*61619*/;
assign _21964_ = _21442_ ^ _21960_ /*61622*/;
assign _21965_ = _21956_ & _21964_ /*61620*/;
assign _21890_ = _21956_ ^ _21964_ /*61621*/;
assign _21962_ = _21963_ | _21965_ /*61618*/;
assign _21967_ = ~Q[39] /*61617*/;
assign _21966_ = _21967_ & D[2] /*61616*/;
assign _21969_ = _21443_ & _21966_ /*61611*/;
assign _21970_ = _21443_ ^ _21966_ /*61614*/;
assign _21971_ = _21962_ & _21970_ /*61612*/;
assign _21891_ = _21962_ ^ _21970_ /*61613*/;
assign _21968_ = _21969_ | _21971_ /*61610*/;
assign _21973_ = ~Q[39] /*61609*/;
assign _21972_ = _21973_ & D[3] /*61608*/;
assign _21975_ = _21444_ & _21972_ /*61603*/;
assign _21976_ = _21444_ ^ _21972_ /*61606*/;
assign _21977_ = _21968_ & _21976_ /*61604*/;
assign _21892_ = _21968_ ^ _21976_ /*61605*/;
assign _21974_ = _21975_ | _21977_ /*61602*/;
assign _21979_ = ~Q[39] /*61601*/;
assign _21978_ = _21979_ & D[4] /*61600*/;
assign _21981_ = _21445_ & _21978_ /*61595*/;
assign _21982_ = _21445_ ^ _21978_ /*61598*/;
assign _21983_ = _21974_ & _21982_ /*61596*/;
assign _21893_ = _21974_ ^ _21982_ /*61597*/;
assign _21980_ = _21981_ | _21983_ /*61594*/;
assign _21985_ = ~Q[39] /*61593*/;
assign _21984_ = _21985_ & D[5] /*61592*/;
assign _21987_ = _21446_ & _21984_ /*61587*/;
assign _21988_ = _21446_ ^ _21984_ /*61590*/;
assign _21989_ = _21980_ & _21988_ /*61588*/;
assign _21894_ = _21980_ ^ _21988_ /*61589*/;
assign _21986_ = _21987_ | _21989_ /*61586*/;
assign _21991_ = ~Q[39] /*61585*/;
assign _21990_ = _21991_ & D[6] /*61584*/;
assign _21993_ = _21447_ & _21990_ /*61579*/;
assign _21994_ = _21447_ ^ _21990_ /*61582*/;
assign _21995_ = _21986_ & _21994_ /*61580*/;
assign _21895_ = _21986_ ^ _21994_ /*61581*/;
assign _21992_ = _21993_ | _21995_ /*61578*/;
assign _21997_ = ~Q[39] /*61577*/;
assign _21996_ = _21997_ & D[7] /*61576*/;
assign _21999_ = _21448_ & _21996_ /*61571*/;
assign _22000_ = _21448_ ^ _21996_ /*61574*/;
assign _22001_ = _21992_ & _22000_ /*61572*/;
assign _21896_ = _21992_ ^ _22000_ /*61573*/;
assign _21998_ = _21999_ | _22001_ /*61570*/;
assign _22003_ = ~Q[39] /*61569*/;
assign _22002_ = _22003_ & D[8] /*61568*/;
assign _22005_ = _21449_ & _22002_ /*61563*/;
assign _22006_ = _21449_ ^ _22002_ /*61566*/;
assign _22007_ = _21998_ & _22006_ /*61564*/;
assign _21897_ = _21998_ ^ _22006_ /*61565*/;
assign _22004_ = _22005_ | _22007_ /*61562*/;
assign _22009_ = ~Q[39] /*61561*/;
assign _22008_ = _22009_ & D[9] /*61560*/;
assign _22011_ = _21450_ & _22008_ /*61555*/;
assign _22012_ = _21450_ ^ _22008_ /*61558*/;
assign _22013_ = _22004_ & _22012_ /*61556*/;
assign _21898_ = _22004_ ^ _22012_ /*61557*/;
assign _22010_ = _22011_ | _22013_ /*61554*/;
assign _22015_ = ~Q[39] /*61553*/;
assign _22014_ = _22015_ & D[10] /*61552*/;
assign _22017_ = _21451_ & _22014_ /*61547*/;
assign _22018_ = _21451_ ^ _22014_ /*61550*/;
assign _22019_ = _22010_ & _22018_ /*61548*/;
assign _21899_ = _22010_ ^ _22018_ /*61549*/;
assign _22016_ = _22017_ | _22019_ /*61546*/;
assign _22021_ = ~Q[39] /*61545*/;
assign _22020_ = _22021_ & D[11] /*61544*/;
assign _22023_ = _21452_ & _22020_ /*61539*/;
assign _22024_ = _21452_ ^ _22020_ /*61542*/;
assign _22025_ = _22016_ & _22024_ /*61540*/;
assign _21900_ = _22016_ ^ _22024_ /*61541*/;
assign _22022_ = _22023_ | _22025_ /*61538*/;
assign _22027_ = ~Q[39] /*61537*/;
assign _22026_ = _22027_ & D[12] /*61536*/;
assign _22029_ = _21453_ & _22026_ /*61531*/;
assign _22030_ = _21453_ ^ _22026_ /*61534*/;
assign _22031_ = _22022_ & _22030_ /*61532*/;
assign _21901_ = _22022_ ^ _22030_ /*61533*/;
assign _22028_ = _22029_ | _22031_ /*61530*/;
assign _22033_ = ~Q[39] /*61529*/;
assign _22032_ = _22033_ & D[13] /*61528*/;
assign _22035_ = _21454_ & _22032_ /*61523*/;
assign _22036_ = _21454_ ^ _22032_ /*61526*/;
assign _22037_ = _22028_ & _22036_ /*61524*/;
assign _21902_ = _22028_ ^ _22036_ /*61525*/;
assign _22034_ = _22035_ | _22037_ /*61522*/;
assign _22039_ = ~Q[39] /*61521*/;
assign _22038_ = _22039_ & D[14] /*61520*/;
assign _22041_ = _21455_ & _22038_ /*61515*/;
assign _22042_ = _21455_ ^ _22038_ /*61518*/;
assign _22043_ = _22034_ & _22042_ /*61516*/;
assign _21903_ = _22034_ ^ _22042_ /*61517*/;
assign _22040_ = _22041_ | _22043_ /*61514*/;
assign _22045_ = ~Q[39] /*61513*/;
assign _22044_ = _22045_ & D[15] /*61512*/;
assign _22047_ = _21456_ & _22044_ /*61507*/;
assign _22048_ = _21456_ ^ _22044_ /*61510*/;
assign _22049_ = _22040_ & _22048_ /*61508*/;
assign _21904_ = _22040_ ^ _22048_ /*61509*/;
assign _22046_ = _22047_ | _22049_ /*61506*/;
assign _22051_ = ~Q[39] /*61505*/;
assign _22050_ = _22051_ & D[16] /*61504*/;
assign _22053_ = _21457_ & _22050_ /*61499*/;
assign _22054_ = _21457_ ^ _22050_ /*61502*/;
assign _22055_ = _22046_ & _22054_ /*61500*/;
assign _21905_ = _22046_ ^ _22054_ /*61501*/;
assign _22052_ = _22053_ | _22055_ /*61498*/;
assign _22057_ = ~Q[39] /*61497*/;
assign _22056_ = _22057_ & D[17] /*61496*/;
assign _22059_ = _21458_ & _22056_ /*61491*/;
assign _22060_ = _21458_ ^ _22056_ /*61494*/;
assign _22061_ = _22052_ & _22060_ /*61492*/;
assign _21906_ = _22052_ ^ _22060_ /*61493*/;
assign _22058_ = _22059_ | _22061_ /*61490*/;
assign _22063_ = ~Q[39] /*61489*/;
assign _22062_ = _22063_ & D[18] /*61488*/;
assign _22065_ = _21459_ & _22062_ /*61483*/;
assign _22066_ = _21459_ ^ _22062_ /*61486*/;
assign _22067_ = _22058_ & _22066_ /*61484*/;
assign _21907_ = _22058_ ^ _22066_ /*61485*/;
assign _22064_ = _22065_ | _22067_ /*61482*/;
assign _22069_ = ~Q[39] /*61481*/;
assign _22068_ = _22069_ & D[19] /*61480*/;
assign _22071_ = _21460_ & _22068_ /*61475*/;
assign _22072_ = _21460_ ^ _22068_ /*61478*/;
assign _22073_ = _22064_ & _22072_ /*61476*/;
assign _21908_ = _22064_ ^ _22072_ /*61477*/;
assign _22070_ = _22071_ | _22073_ /*61474*/;
assign _22075_ = ~Q[39] /*61473*/;
assign _22074_ = _22075_ & D[20] /*61472*/;
assign _22077_ = _21461_ & _22074_ /*61467*/;
assign _22078_ = _21461_ ^ _22074_ /*61470*/;
assign _22079_ = _22070_ & _22078_ /*61468*/;
assign _21909_ = _22070_ ^ _22078_ /*61469*/;
assign _22076_ = _22077_ | _22079_ /*61466*/;
assign _22081_ = ~Q[39] /*61465*/;
assign _22080_ = _22081_ & D[21] /*61464*/;
assign _22083_ = _21462_ & _22080_ /*61459*/;
assign _22084_ = _21462_ ^ _22080_ /*61462*/;
assign _22085_ = _22076_ & _22084_ /*61460*/;
assign _21910_ = _22076_ ^ _22084_ /*61461*/;
assign _22082_ = _22083_ | _22085_ /*61458*/;
assign _22087_ = ~Q[39] /*61457*/;
assign _22086_ = _22087_ & D[22] /*61456*/;
assign _22089_ = _21463_ & _22086_ /*61451*/;
assign _22090_ = _21463_ ^ _22086_ /*61454*/;
assign _22091_ = _22082_ & _22090_ /*61452*/;
assign _21911_ = _22082_ ^ _22090_ /*61453*/;
assign _22088_ = _22089_ | _22091_ /*61450*/;
assign _22093_ = ~Q[39] /*61449*/;
assign _22092_ = _22093_ & D[23] /*61448*/;
assign _22095_ = _21464_ & _22092_ /*61443*/;
assign _22096_ = _21464_ ^ _22092_ /*61446*/;
assign _22097_ = _22088_ & _22096_ /*61444*/;
assign _21912_ = _22088_ ^ _22096_ /*61445*/;
assign _22094_ = _22095_ | _22097_ /*61442*/;
assign _22099_ = ~Q[39] /*61441*/;
assign _22098_ = _22099_ & D[24] /*61440*/;
assign _22101_ = _21465_ & _22098_ /*61435*/;
assign _22102_ = _21465_ ^ _22098_ /*61438*/;
assign _22103_ = _22094_ & _22102_ /*61436*/;
assign _21913_ = _22094_ ^ _22102_ /*61437*/;
assign _22100_ = _22101_ | _22103_ /*61434*/;
assign _22105_ = ~Q[39] /*61433*/;
assign _22104_ = _22105_ & D[25] /*61432*/;
assign _22107_ = _21466_ & _22104_ /*61427*/;
assign _22108_ = _21466_ ^ _22104_ /*61430*/;
assign _22109_ = _22100_ & _22108_ /*61428*/;
assign _21914_ = _22100_ ^ _22108_ /*61429*/;
assign _22106_ = _22107_ | _22109_ /*61426*/;
assign _22111_ = ~Q[39] /*61425*/;
assign _22110_ = _22111_ & D[26] /*61424*/;
assign _22113_ = _21467_ & _22110_ /*61419*/;
assign _22114_ = _21467_ ^ _22110_ /*61422*/;
assign _22115_ = _22106_ & _22114_ /*61420*/;
assign _21915_ = _22106_ ^ _22114_ /*61421*/;
assign _22112_ = _22113_ | _22115_ /*61418*/;
assign _22117_ = ~Q[39] /*61417*/;
assign _22116_ = _22117_ & D[27] /*61416*/;
assign _22119_ = _21468_ & _22116_ /*61411*/;
assign _22120_ = _21468_ ^ _22116_ /*61414*/;
assign _22121_ = _22112_ & _22120_ /*61412*/;
assign _21916_ = _22112_ ^ _22120_ /*61413*/;
assign _22118_ = _22119_ | _22121_ /*61410*/;
assign _22123_ = ~Q[39] /*61409*/;
assign _22122_ = _22123_ & D[28] /*61408*/;
assign _22125_ = _21469_ & _22122_ /*61403*/;
assign _22126_ = _21469_ ^ _22122_ /*61406*/;
assign _22127_ = _22118_ & _22126_ /*61404*/;
assign _21917_ = _22118_ ^ _22126_ /*61405*/;
assign _22124_ = _22125_ | _22127_ /*61402*/;
assign _22129_ = ~Q[39] /*61401*/;
assign _22128_ = _22129_ & D[29] /*61400*/;
assign _22131_ = _21470_ & _22128_ /*61395*/;
assign _22132_ = _21470_ ^ _22128_ /*61398*/;
assign _22133_ = _22124_ & _22132_ /*61396*/;
assign _21918_ = _22124_ ^ _22132_ /*61397*/;
assign _22130_ = _22131_ | _22133_ /*61394*/;
assign _22135_ = ~Q[39] /*61393*/;
assign _22134_ = _22135_ & D[30] /*61392*/;
assign _22137_ = _21471_ & _22134_ /*61387*/;
assign _22138_ = _21471_ ^ _22134_ /*61390*/;
assign _22139_ = _22130_ & _22138_ /*61388*/;
assign _21919_ = _22130_ ^ _22138_ /*61389*/;
assign _22136_ = _22137_ | _22139_ /*61386*/;
assign _22141_ = ~Q[39] /*61385*/;
assign _22140_ = _22141_ & D[31] /*61384*/;
assign _22143_ = _21472_ & _22140_ /*61379*/;
assign _22144_ = _21472_ ^ _22140_ /*61382*/;
assign _22145_ = _22136_ & _22144_ /*61380*/;
assign _21920_ = _22136_ ^ _22144_ /*61381*/;
assign _22142_ = _22143_ | _22145_ /*61378*/;
assign _22147_ = ~Q[39] /*61377*/;
assign _22146_ = _22147_ & D[32] /*61376*/;
assign _22149_ = _21473_ & _22146_ /*61371*/;
assign _22150_ = _21473_ ^ _22146_ /*61374*/;
assign _22151_ = _22142_ & _22150_ /*61372*/;
assign _21921_ = _22142_ ^ _22150_ /*61373*/;
assign _22148_ = _22149_ | _22151_ /*61370*/;
assign _22153_ = ~Q[39] /*61369*/;
assign _22152_ = _22153_ & D[33] /*61368*/;
assign _22155_ = _21474_ & _22152_ /*61363*/;
assign _22156_ = _21474_ ^ _22152_ /*61366*/;
assign _22157_ = _22148_ & _22156_ /*61364*/;
assign _21922_ = _22148_ ^ _22156_ /*61365*/;
assign _22154_ = _22155_ | _22157_ /*61362*/;
assign _22159_ = ~Q[39] /*61361*/;
assign _22158_ = _22159_ & D[34] /*61360*/;
assign _22161_ = _21475_ & _22158_ /*61355*/;
assign _22162_ = _21475_ ^ _22158_ /*61358*/;
assign _22163_ = _22154_ & _22162_ /*61356*/;
assign _21923_ = _22154_ ^ _22162_ /*61357*/;
assign _22160_ = _22161_ | _22163_ /*61354*/;
assign _22165_ = ~Q[39] /*61353*/;
assign _22164_ = _22165_ & D[35] /*61352*/;
assign _22167_ = _21476_ & _22164_ /*61347*/;
assign _22168_ = _21476_ ^ _22164_ /*61350*/;
assign _22169_ = _22160_ & _22168_ /*61348*/;
assign _21924_ = _22160_ ^ _22168_ /*61349*/;
assign _22166_ = _22167_ | _22169_ /*61346*/;
assign _22171_ = ~Q[39] /*61345*/;
assign _22170_ = _22171_ & D[36] /*61344*/;
assign _22173_ = _21477_ & _22170_ /*61339*/;
assign _22174_ = _21477_ ^ _22170_ /*61342*/;
assign _22175_ = _22166_ & _22174_ /*61340*/;
assign _21925_ = _22166_ ^ _22174_ /*61341*/;
assign _22172_ = _22173_ | _22175_ /*61338*/;
assign _22177_ = ~Q[39] /*61337*/;
assign _22176_ = _22177_ & D[37] /*61336*/;
assign _22179_ = _21478_ & _22176_ /*61331*/;
assign _22180_ = _21478_ ^ _22176_ /*61334*/;
assign _22181_ = _22172_ & _22180_ /*61332*/;
assign _21926_ = _22172_ ^ _22180_ /*61333*/;
assign _22178_ = _22179_ | _22181_ /*61330*/;
assign _22183_ = ~Q[39] /*61329*/;
assign _22182_ = _22183_ & D[38] /*61328*/;
assign _22185_ = _21479_ & _22182_ /*61323*/;
assign _22186_ = _21479_ ^ _22182_ /*61326*/;
assign _22187_ = _22178_ & _22186_ /*61324*/;
assign _21927_ = _22178_ ^ _22186_ /*61325*/;
assign _22184_ = _22185_ | _22187_ /*61322*/;
assign _22189_ = ~Q[39] /*61321*/;
assign _22188_ = _22189_ & D[39] /*61320*/;
assign _22191_ = _21480_ & _22188_ /*61315*/;
assign _22192_ = _21480_ ^ _22188_ /*61318*/;
assign _22193_ = _22184_ & _22192_ /*61316*/;
assign _21928_ = _22184_ ^ _22192_ /*61317*/;
assign _22190_ = _22191_ | _22193_ /*61314*/;
assign _22195_ = ~Q[39] /*61313*/;
assign _22194_ = _22195_ & D[40] /*61312*/;
assign _22197_ = _21481_ & _22194_ /*61307*/;
assign _22198_ = _21481_ ^ _22194_ /*61310*/;
assign _22199_ = _22190_ & _22198_ /*61308*/;
assign _21929_ = _22190_ ^ _22198_ /*61309*/;
assign _22196_ = _22197_ | _22199_ /*61306*/;
assign _22201_ = ~Q[39] /*61305*/;
assign _22200_ = _22201_ & D[41] /*61304*/;
assign _22203_ = _21482_ & _22200_ /*61299*/;
assign _22204_ = _21482_ ^ _22200_ /*61302*/;
assign _22205_ = _22196_ & _22204_ /*61300*/;
assign _21930_ = _22196_ ^ _22204_ /*61301*/;
assign _22202_ = _22203_ | _22205_ /*61298*/;
assign _22207_ = ~Q[39] /*61297*/;
assign _22206_ = _22207_ & D[42] /*61296*/;
assign _22209_ = _21483_ & _22206_ /*61291*/;
assign _22210_ = _21483_ ^ _22206_ /*61294*/;
assign _22211_ = _22202_ & _22210_ /*61292*/;
assign _21931_ = _22202_ ^ _22210_ /*61293*/;
assign _22208_ = _22209_ | _22211_ /*61290*/;
assign _22213_ = ~Q[39] /*61289*/;
assign _22212_ = _22213_ & D[43] /*61288*/;
assign _22215_ = _21484_ & _22212_ /*61283*/;
assign _22216_ = _21484_ ^ _22212_ /*61286*/;
assign _22217_ = _22208_ & _22216_ /*61284*/;
assign _21932_ = _22208_ ^ _22216_ /*61285*/;
assign _22214_ = _22215_ | _22217_ /*61282*/;
assign _22219_ = ~Q[39] /*61281*/;
assign _22218_ = _22219_ & D[44] /*61280*/;
assign _22221_ = _21485_ & _22218_ /*61275*/;
assign _22222_ = _21485_ ^ _22218_ /*61278*/;
assign _22223_ = _22214_ & _22222_ /*61276*/;
assign _21933_ = _22214_ ^ _22222_ /*61277*/;
assign _22220_ = _22221_ | _22223_ /*61274*/;
assign _22225_ = ~Q[39] /*61273*/;
assign _22224_ = _22225_ & D[45] /*61272*/;
assign _22227_ = _21486_ & _22224_ /*61267*/;
assign _22228_ = _21486_ ^ _22224_ /*61270*/;
assign _22229_ = _22220_ & _22228_ /*61268*/;
assign _21934_ = _22220_ ^ _22228_ /*61269*/;
assign _22226_ = _22227_ | _22229_ /*61266*/;
assign _22231_ = ~Q[39] /*61265*/;
assign _22230_ = _22231_ & D[46] /*61264*/;
assign _22233_ = _21487_ & _22230_ /*61259*/;
assign _22234_ = _21487_ ^ _22230_ /*61262*/;
assign _22235_ = _22226_ & _22234_ /*61260*/;
assign _21935_ = _22226_ ^ _22234_ /*61261*/;
assign _22232_ = _22233_ | _22235_ /*61258*/;
assign _22237_ = ~Q[39] /*61257*/;
assign _22236_ = _22237_ & D[47] /*61256*/;
assign _22239_ = _21488_ & _22236_ /*61251*/;
assign _22240_ = _21488_ ^ _22236_ /*61254*/;
assign _22241_ = _22232_ & _22240_ /*61252*/;
assign _21936_ = _22232_ ^ _22240_ /*61253*/;
assign _22238_ = _22239_ | _22241_ /*61250*/;
assign _22243_ = ~Q[39] /*61249*/;
assign _22242_ = _22243_ & D[48] /*61248*/;
assign _22245_ = _21489_ & _22242_ /*61243*/;
assign _22246_ = _21489_ ^ _22242_ /*61246*/;
assign _22247_ = _22238_ & _22246_ /*61244*/;
assign _21937_ = _22238_ ^ _22246_ /*61245*/;
assign _22244_ = _22245_ | _22247_ /*61242*/;
assign _22249_ = ~Q[39] /*61241*/;
assign _22248_ = _22249_ & D[49] /*61240*/;
assign _22251_ = _21490_ & _22248_ /*61235*/;
assign _22252_ = _21490_ ^ _22248_ /*61238*/;
assign _22253_ = _22244_ & _22252_ /*61236*/;
assign _21938_ = _22244_ ^ _22252_ /*61237*/;
assign _22250_ = _22251_ | _22253_ /*61234*/;
assign _22255_ = ~Q[39] /*61233*/;
assign _22254_ = _22255_ & D[50] /*61232*/;
assign _22257_ = _21491_ & _22254_ /*61227*/;
assign _22258_ = _21491_ ^ _22254_ /*61230*/;
assign _22259_ = _22250_ & _22258_ /*61228*/;
assign _21939_ = _22250_ ^ _22258_ /*61229*/;
assign _22256_ = _22257_ | _22259_ /*61226*/;
assign _22261_ = ~Q[39] /*61225*/;
assign _22260_ = _22261_ & D[51] /*61224*/;
assign _22263_ = _21492_ & _22260_ /*61219*/;
assign _22264_ = _21492_ ^ _22260_ /*61222*/;
assign _22265_ = _22256_ & _22264_ /*61220*/;
assign _21940_ = _22256_ ^ _22264_ /*61221*/;
assign _22262_ = _22263_ | _22265_ /*61218*/;
assign _22267_ = ~Q[39] /*61217*/;
assign _22266_ = _22267_ & D[52] /*61216*/;
assign _22269_ = _21493_ & _22266_ /*61211*/;
assign _22270_ = _21493_ ^ _22266_ /*61214*/;
assign _22271_ = _22262_ & _22270_ /*61212*/;
assign _21941_ = _22262_ ^ _22270_ /*61213*/;
assign _22268_ = _22269_ | _22271_ /*61210*/;
assign _22273_ = ~Q[39] /*61209*/;
assign _22272_ = _22273_ & D[53] /*61208*/;
assign _22275_ = _21494_ & _22272_ /*61203*/;
assign _22276_ = _21494_ ^ _22272_ /*61206*/;
assign _22277_ = _22268_ & _22276_ /*61204*/;
assign _21942_ = _22268_ ^ _22276_ /*61205*/;
assign _22274_ = _22275_ | _22277_ /*61202*/;
assign _22279_ = ~Q[39] /*61201*/;
assign _22278_ = _22279_ & D[54] /*61200*/;
assign _22281_ = _21495_ & _22278_ /*61195*/;
assign _22282_ = _21495_ ^ _22278_ /*61198*/;
assign _22283_ = _22274_ & _22282_ /*61196*/;
assign _21943_ = _22274_ ^ _22282_ /*61197*/;
assign _22280_ = _22281_ | _22283_ /*61194*/;
assign _22285_ = ~Q[39] /*61193*/;
assign _22284_ = _22285_ & D[55] /*61192*/;
assign _22287_ = _21496_ & _22284_ /*61187*/;
assign _22288_ = _21496_ ^ _22284_ /*61190*/;
assign _22289_ = _22280_ & _22288_ /*61188*/;
assign _21944_ = _22280_ ^ _22288_ /*61189*/;
assign _22286_ = _22287_ | _22289_ /*61186*/;
assign _22291_ = ~Q[39] /*61185*/;
assign _22290_ = _22291_ & D[56] /*61184*/;
assign _22293_ = _21497_ & _22290_ /*61179*/;
assign _22294_ = _21497_ ^ _22290_ /*61182*/;
assign _22295_ = _22286_ & _22294_ /*61180*/;
assign _21945_ = _22286_ ^ _22294_ /*61181*/;
assign _22292_ = _22293_ | _22295_ /*61178*/;
assign _22297_ = ~Q[39] /*61177*/;
assign _22296_ = _22297_ & D[57] /*61176*/;
assign _22299_ = _21498_ & _22296_ /*61171*/;
assign _22300_ = _21498_ ^ _22296_ /*61174*/;
assign _22301_ = _22292_ & _22300_ /*61172*/;
assign _21946_ = _22292_ ^ _22300_ /*61173*/;
assign _22298_ = _22299_ | _22301_ /*61170*/;
assign _22303_ = ~Q[39] /*61169*/;
assign _22302_ = _22303_ & D[58] /*61168*/;
assign _22305_ = _21499_ & _22302_ /*61163*/;
assign _22306_ = _21499_ ^ _22302_ /*61166*/;
assign _22307_ = _22298_ & _22306_ /*61164*/;
assign _21947_ = _22298_ ^ _22306_ /*61165*/;
assign _22304_ = _22305_ | _22307_ /*61162*/;
assign _22309_ = ~Q[39] /*61161*/;
assign _22308_ = _22309_ & D[59] /*61160*/;
assign _22311_ = _21500_ & _22308_ /*61155*/;
assign _22312_ = _21500_ ^ _22308_ /*61158*/;
assign _22313_ = _22304_ & _22312_ /*61156*/;
assign _21948_ = _22304_ ^ _22312_ /*61157*/;
assign _22310_ = _22311_ | _22313_ /*61154*/;
assign _22315_ = ~Q[39] /*61153*/;
assign _22314_ = _22315_ & D[60] /*61152*/;
assign _22317_ = _21501_ & _22314_ /*61147*/;
assign _22318_ = _21501_ ^ _22314_ /*61150*/;
assign _22319_ = _22310_ & _22318_ /*61148*/;
assign _21949_ = _22310_ ^ _22318_ /*61149*/;
assign _22316_ = _22317_ | _22319_ /*61146*/;
assign _22321_ = ~Q[39] /*61145*/;
assign _22320_ = _22321_ & D[61] /*61144*/;
assign _22323_ = _21502_ & _22320_ /*61139*/;
assign _22324_ = _21502_ ^ _22320_ /*61142*/;
assign _22325_ = _22316_ & _22324_ /*61140*/;
assign _21950_ = _22316_ ^ _22324_ /*61141*/;
assign _22322_ = _22323_ | _22325_ /*61138*/;
assign _22327_ = ~Q[39] /*61137*/;
assign _22326_ = _22327_ & D[62] /*61136*/;
assign _22329_ = _21503_ & _22326_ /*61131*/;
assign _22330_ = _21503_ ^ _22326_ /*61134*/;
assign _22331_ = _22322_ & _22330_ /*61132*/;
assign _21951_ = _22322_ ^ _22330_ /*61133*/;
assign _22328_ = _22329_ | _22331_ /*61130*/;
assign _22333_ = ~Q[39] /*61129*/;
assign _22332_ = _22333_ & zeroWire /*61128*/;
assign _22334_ = _21504_ ^ _22332_ /*61126*/;
assign _21952_ = _22334_ ^ _22328_ /*61125*/;
assign _22405_ = ~D[0] /*60871*/;
assign _22402_ = R_0[38] & _22405_ /*60867*/;
assign _22403_ = R_0[38] ^ _22405_ /*60870*/;
assign _22404_ = oneWire & _22403_ /*60868*/;
assign _22337_ = oneWire ^ _22403_ /*60869*/;
assign _22401_ = _22402_ | _22404_ /*60866*/;
assign _22410_ = ~D[1] /*60865*/;
assign _22407_ = _21889_ & _22410_ /*60861*/;
assign _22408_ = _21889_ ^ _22410_ /*60864*/;
assign _22409_ = _22401_ & _22408_ /*60862*/;
assign _22338_ = _22401_ ^ _22408_ /*60863*/;
assign _22406_ = _22407_ | _22409_ /*60860*/;
assign _22415_ = ~D[2] /*60859*/;
assign _22412_ = _21890_ & _22415_ /*60855*/;
assign _22413_ = _21890_ ^ _22415_ /*60858*/;
assign _22414_ = _22406_ & _22413_ /*60856*/;
assign _22339_ = _22406_ ^ _22413_ /*60857*/;
assign _22411_ = _22412_ | _22414_ /*60854*/;
assign _22420_ = ~D[3] /*60853*/;
assign _22417_ = _21891_ & _22420_ /*60849*/;
assign _22418_ = _21891_ ^ _22420_ /*60852*/;
assign _22419_ = _22411_ & _22418_ /*60850*/;
assign _22340_ = _22411_ ^ _22418_ /*60851*/;
assign _22416_ = _22417_ | _22419_ /*60848*/;
assign _22425_ = ~D[4] /*60847*/;
assign _22422_ = _21892_ & _22425_ /*60843*/;
assign _22423_ = _21892_ ^ _22425_ /*60846*/;
assign _22424_ = _22416_ & _22423_ /*60844*/;
assign _22341_ = _22416_ ^ _22423_ /*60845*/;
assign _22421_ = _22422_ | _22424_ /*60842*/;
assign _22430_ = ~D[5] /*60841*/;
assign _22427_ = _21893_ & _22430_ /*60837*/;
assign _22428_ = _21893_ ^ _22430_ /*60840*/;
assign _22429_ = _22421_ & _22428_ /*60838*/;
assign _22342_ = _22421_ ^ _22428_ /*60839*/;
assign _22426_ = _22427_ | _22429_ /*60836*/;
assign _22435_ = ~D[6] /*60835*/;
assign _22432_ = _21894_ & _22435_ /*60831*/;
assign _22433_ = _21894_ ^ _22435_ /*60834*/;
assign _22434_ = _22426_ & _22433_ /*60832*/;
assign _22343_ = _22426_ ^ _22433_ /*60833*/;
assign _22431_ = _22432_ | _22434_ /*60830*/;
assign _22440_ = ~D[7] /*60829*/;
assign _22437_ = _21895_ & _22440_ /*60825*/;
assign _22438_ = _21895_ ^ _22440_ /*60828*/;
assign _22439_ = _22431_ & _22438_ /*60826*/;
assign _22344_ = _22431_ ^ _22438_ /*60827*/;
assign _22436_ = _22437_ | _22439_ /*60824*/;
assign _22445_ = ~D[8] /*60823*/;
assign _22442_ = _21896_ & _22445_ /*60819*/;
assign _22443_ = _21896_ ^ _22445_ /*60822*/;
assign _22444_ = _22436_ & _22443_ /*60820*/;
assign _22345_ = _22436_ ^ _22443_ /*60821*/;
assign _22441_ = _22442_ | _22444_ /*60818*/;
assign _22450_ = ~D[9] /*60817*/;
assign _22447_ = _21897_ & _22450_ /*60813*/;
assign _22448_ = _21897_ ^ _22450_ /*60816*/;
assign _22449_ = _22441_ & _22448_ /*60814*/;
assign _22346_ = _22441_ ^ _22448_ /*60815*/;
assign _22446_ = _22447_ | _22449_ /*60812*/;
assign _22455_ = ~D[10] /*60811*/;
assign _22452_ = _21898_ & _22455_ /*60807*/;
assign _22453_ = _21898_ ^ _22455_ /*60810*/;
assign _22454_ = _22446_ & _22453_ /*60808*/;
assign _22347_ = _22446_ ^ _22453_ /*60809*/;
assign _22451_ = _22452_ | _22454_ /*60806*/;
assign _22460_ = ~D[11] /*60805*/;
assign _22457_ = _21899_ & _22460_ /*60801*/;
assign _22458_ = _21899_ ^ _22460_ /*60804*/;
assign _22459_ = _22451_ & _22458_ /*60802*/;
assign _22348_ = _22451_ ^ _22458_ /*60803*/;
assign _22456_ = _22457_ | _22459_ /*60800*/;
assign _22465_ = ~D[12] /*60799*/;
assign _22462_ = _21900_ & _22465_ /*60795*/;
assign _22463_ = _21900_ ^ _22465_ /*60798*/;
assign _22464_ = _22456_ & _22463_ /*60796*/;
assign _22349_ = _22456_ ^ _22463_ /*60797*/;
assign _22461_ = _22462_ | _22464_ /*60794*/;
assign _22470_ = ~D[13] /*60793*/;
assign _22467_ = _21901_ & _22470_ /*60789*/;
assign _22468_ = _21901_ ^ _22470_ /*60792*/;
assign _22469_ = _22461_ & _22468_ /*60790*/;
assign _22350_ = _22461_ ^ _22468_ /*60791*/;
assign _22466_ = _22467_ | _22469_ /*60788*/;
assign _22475_ = ~D[14] /*60787*/;
assign _22472_ = _21902_ & _22475_ /*60783*/;
assign _22473_ = _21902_ ^ _22475_ /*60786*/;
assign _22474_ = _22466_ & _22473_ /*60784*/;
assign _22351_ = _22466_ ^ _22473_ /*60785*/;
assign _22471_ = _22472_ | _22474_ /*60782*/;
assign _22480_ = ~D[15] /*60781*/;
assign _22477_ = _21903_ & _22480_ /*60777*/;
assign _22478_ = _21903_ ^ _22480_ /*60780*/;
assign _22479_ = _22471_ & _22478_ /*60778*/;
assign _22352_ = _22471_ ^ _22478_ /*60779*/;
assign _22476_ = _22477_ | _22479_ /*60776*/;
assign _22485_ = ~D[16] /*60775*/;
assign _22482_ = _21904_ & _22485_ /*60771*/;
assign _22483_ = _21904_ ^ _22485_ /*60774*/;
assign _22484_ = _22476_ & _22483_ /*60772*/;
assign _22353_ = _22476_ ^ _22483_ /*60773*/;
assign _22481_ = _22482_ | _22484_ /*60770*/;
assign _22490_ = ~D[17] /*60769*/;
assign _22487_ = _21905_ & _22490_ /*60765*/;
assign _22488_ = _21905_ ^ _22490_ /*60768*/;
assign _22489_ = _22481_ & _22488_ /*60766*/;
assign _22354_ = _22481_ ^ _22488_ /*60767*/;
assign _22486_ = _22487_ | _22489_ /*60764*/;
assign _22495_ = ~D[18] /*60763*/;
assign _22492_ = _21906_ & _22495_ /*60759*/;
assign _22493_ = _21906_ ^ _22495_ /*60762*/;
assign _22494_ = _22486_ & _22493_ /*60760*/;
assign _22355_ = _22486_ ^ _22493_ /*60761*/;
assign _22491_ = _22492_ | _22494_ /*60758*/;
assign _22500_ = ~D[19] /*60757*/;
assign _22497_ = _21907_ & _22500_ /*60753*/;
assign _22498_ = _21907_ ^ _22500_ /*60756*/;
assign _22499_ = _22491_ & _22498_ /*60754*/;
assign _22356_ = _22491_ ^ _22498_ /*60755*/;
assign _22496_ = _22497_ | _22499_ /*60752*/;
assign _22505_ = ~D[20] /*60751*/;
assign _22502_ = _21908_ & _22505_ /*60747*/;
assign _22503_ = _21908_ ^ _22505_ /*60750*/;
assign _22504_ = _22496_ & _22503_ /*60748*/;
assign _22357_ = _22496_ ^ _22503_ /*60749*/;
assign _22501_ = _22502_ | _22504_ /*60746*/;
assign _22510_ = ~D[21] /*60745*/;
assign _22507_ = _21909_ & _22510_ /*60741*/;
assign _22508_ = _21909_ ^ _22510_ /*60744*/;
assign _22509_ = _22501_ & _22508_ /*60742*/;
assign _22358_ = _22501_ ^ _22508_ /*60743*/;
assign _22506_ = _22507_ | _22509_ /*60740*/;
assign _22515_ = ~D[22] /*60739*/;
assign _22512_ = _21910_ & _22515_ /*60735*/;
assign _22513_ = _21910_ ^ _22515_ /*60738*/;
assign _22514_ = _22506_ & _22513_ /*60736*/;
assign _22359_ = _22506_ ^ _22513_ /*60737*/;
assign _22511_ = _22512_ | _22514_ /*60734*/;
assign _22520_ = ~D[23] /*60733*/;
assign _22517_ = _21911_ & _22520_ /*60729*/;
assign _22518_ = _21911_ ^ _22520_ /*60732*/;
assign _22519_ = _22511_ & _22518_ /*60730*/;
assign _22360_ = _22511_ ^ _22518_ /*60731*/;
assign _22516_ = _22517_ | _22519_ /*60728*/;
assign _22525_ = ~D[24] /*60727*/;
assign _22522_ = _21912_ & _22525_ /*60723*/;
assign _22523_ = _21912_ ^ _22525_ /*60726*/;
assign _22524_ = _22516_ & _22523_ /*60724*/;
assign _22361_ = _22516_ ^ _22523_ /*60725*/;
assign _22521_ = _22522_ | _22524_ /*60722*/;
assign _22530_ = ~D[25] /*60721*/;
assign _22527_ = _21913_ & _22530_ /*60717*/;
assign _22528_ = _21913_ ^ _22530_ /*60720*/;
assign _22529_ = _22521_ & _22528_ /*60718*/;
assign _22362_ = _22521_ ^ _22528_ /*60719*/;
assign _22526_ = _22527_ | _22529_ /*60716*/;
assign _22535_ = ~D[26] /*60715*/;
assign _22532_ = _21914_ & _22535_ /*60711*/;
assign _22533_ = _21914_ ^ _22535_ /*60714*/;
assign _22534_ = _22526_ & _22533_ /*60712*/;
assign _22363_ = _22526_ ^ _22533_ /*60713*/;
assign _22531_ = _22532_ | _22534_ /*60710*/;
assign _22540_ = ~D[27] /*60709*/;
assign _22537_ = _21915_ & _22540_ /*60705*/;
assign _22538_ = _21915_ ^ _22540_ /*60708*/;
assign _22539_ = _22531_ & _22538_ /*60706*/;
assign _22364_ = _22531_ ^ _22538_ /*60707*/;
assign _22536_ = _22537_ | _22539_ /*60704*/;
assign _22545_ = ~D[28] /*60703*/;
assign _22542_ = _21916_ & _22545_ /*60699*/;
assign _22543_ = _21916_ ^ _22545_ /*60702*/;
assign _22544_ = _22536_ & _22543_ /*60700*/;
assign _22365_ = _22536_ ^ _22543_ /*60701*/;
assign _22541_ = _22542_ | _22544_ /*60698*/;
assign _22550_ = ~D[29] /*60697*/;
assign _22547_ = _21917_ & _22550_ /*60693*/;
assign _22548_ = _21917_ ^ _22550_ /*60696*/;
assign _22549_ = _22541_ & _22548_ /*60694*/;
assign _22366_ = _22541_ ^ _22548_ /*60695*/;
assign _22546_ = _22547_ | _22549_ /*60692*/;
assign _22555_ = ~D[30] /*60691*/;
assign _22552_ = _21918_ & _22555_ /*60687*/;
assign _22553_ = _21918_ ^ _22555_ /*60690*/;
assign _22554_ = _22546_ & _22553_ /*60688*/;
assign _22367_ = _22546_ ^ _22553_ /*60689*/;
assign _22551_ = _22552_ | _22554_ /*60686*/;
assign _22560_ = ~D[31] /*60685*/;
assign _22557_ = _21919_ & _22560_ /*60681*/;
assign _22558_ = _21919_ ^ _22560_ /*60684*/;
assign _22559_ = _22551_ & _22558_ /*60682*/;
assign _22368_ = _22551_ ^ _22558_ /*60683*/;
assign _22556_ = _22557_ | _22559_ /*60680*/;
assign _22565_ = ~D[32] /*60679*/;
assign _22562_ = _21920_ & _22565_ /*60675*/;
assign _22563_ = _21920_ ^ _22565_ /*60678*/;
assign _22564_ = _22556_ & _22563_ /*60676*/;
assign _22369_ = _22556_ ^ _22563_ /*60677*/;
assign _22561_ = _22562_ | _22564_ /*60674*/;
assign _22570_ = ~D[33] /*60673*/;
assign _22567_ = _21921_ & _22570_ /*60669*/;
assign _22568_ = _21921_ ^ _22570_ /*60672*/;
assign _22569_ = _22561_ & _22568_ /*60670*/;
assign _22370_ = _22561_ ^ _22568_ /*60671*/;
assign _22566_ = _22567_ | _22569_ /*60668*/;
assign _22575_ = ~D[34] /*60667*/;
assign _22572_ = _21922_ & _22575_ /*60663*/;
assign _22573_ = _21922_ ^ _22575_ /*60666*/;
assign _22574_ = _22566_ & _22573_ /*60664*/;
assign _22371_ = _22566_ ^ _22573_ /*60665*/;
assign _22571_ = _22572_ | _22574_ /*60662*/;
assign _22580_ = ~D[35] /*60661*/;
assign _22577_ = _21923_ & _22580_ /*60657*/;
assign _22578_ = _21923_ ^ _22580_ /*60660*/;
assign _22579_ = _22571_ & _22578_ /*60658*/;
assign _22372_ = _22571_ ^ _22578_ /*60659*/;
assign _22576_ = _22577_ | _22579_ /*60656*/;
assign _22585_ = ~D[36] /*60655*/;
assign _22582_ = _21924_ & _22585_ /*60651*/;
assign _22583_ = _21924_ ^ _22585_ /*60654*/;
assign _22584_ = _22576_ & _22583_ /*60652*/;
assign _22373_ = _22576_ ^ _22583_ /*60653*/;
assign _22581_ = _22582_ | _22584_ /*60650*/;
assign _22590_ = ~D[37] /*60649*/;
assign _22587_ = _21925_ & _22590_ /*60645*/;
assign _22588_ = _21925_ ^ _22590_ /*60648*/;
assign _22589_ = _22581_ & _22588_ /*60646*/;
assign _22374_ = _22581_ ^ _22588_ /*60647*/;
assign _22586_ = _22587_ | _22589_ /*60644*/;
assign _22595_ = ~D[38] /*60643*/;
assign _22592_ = _21926_ & _22595_ /*60639*/;
assign _22593_ = _21926_ ^ _22595_ /*60642*/;
assign _22594_ = _22586_ & _22593_ /*60640*/;
assign _22375_ = _22586_ ^ _22593_ /*60641*/;
assign _22591_ = _22592_ | _22594_ /*60638*/;
assign _22600_ = ~D[39] /*60637*/;
assign _22597_ = _21927_ & _22600_ /*60633*/;
assign _22598_ = _21927_ ^ _22600_ /*60636*/;
assign _22599_ = _22591_ & _22598_ /*60634*/;
assign _22376_ = _22591_ ^ _22598_ /*60635*/;
assign _22596_ = _22597_ | _22599_ /*60632*/;
assign _22605_ = ~D[40] /*60631*/;
assign _22602_ = _21928_ & _22605_ /*60627*/;
assign _22603_ = _21928_ ^ _22605_ /*60630*/;
assign _22604_ = _22596_ & _22603_ /*60628*/;
assign _22377_ = _22596_ ^ _22603_ /*60629*/;
assign _22601_ = _22602_ | _22604_ /*60626*/;
assign _22610_ = ~D[41] /*60625*/;
assign _22607_ = _21929_ & _22610_ /*60621*/;
assign _22608_ = _21929_ ^ _22610_ /*60624*/;
assign _22609_ = _22601_ & _22608_ /*60622*/;
assign _22378_ = _22601_ ^ _22608_ /*60623*/;
assign _22606_ = _22607_ | _22609_ /*60620*/;
assign _22615_ = ~D[42] /*60619*/;
assign _22612_ = _21930_ & _22615_ /*60615*/;
assign _22613_ = _21930_ ^ _22615_ /*60618*/;
assign _22614_ = _22606_ & _22613_ /*60616*/;
assign _22379_ = _22606_ ^ _22613_ /*60617*/;
assign _22611_ = _22612_ | _22614_ /*60614*/;
assign _22620_ = ~D[43] /*60613*/;
assign _22617_ = _21931_ & _22620_ /*60609*/;
assign _22618_ = _21931_ ^ _22620_ /*60612*/;
assign _22619_ = _22611_ & _22618_ /*60610*/;
assign _22380_ = _22611_ ^ _22618_ /*60611*/;
assign _22616_ = _22617_ | _22619_ /*60608*/;
assign _22625_ = ~D[44] /*60607*/;
assign _22622_ = _21932_ & _22625_ /*60603*/;
assign _22623_ = _21932_ ^ _22625_ /*60606*/;
assign _22624_ = _22616_ & _22623_ /*60604*/;
assign _22381_ = _22616_ ^ _22623_ /*60605*/;
assign _22621_ = _22622_ | _22624_ /*60602*/;
assign _22630_ = ~D[45] /*60601*/;
assign _22627_ = _21933_ & _22630_ /*60597*/;
assign _22628_ = _21933_ ^ _22630_ /*60600*/;
assign _22629_ = _22621_ & _22628_ /*60598*/;
assign _22382_ = _22621_ ^ _22628_ /*60599*/;
assign _22626_ = _22627_ | _22629_ /*60596*/;
assign _22635_ = ~D[46] /*60595*/;
assign _22632_ = _21934_ & _22635_ /*60591*/;
assign _22633_ = _21934_ ^ _22635_ /*60594*/;
assign _22634_ = _22626_ & _22633_ /*60592*/;
assign _22383_ = _22626_ ^ _22633_ /*60593*/;
assign _22631_ = _22632_ | _22634_ /*60590*/;
assign _22640_ = ~D[47] /*60589*/;
assign _22637_ = _21935_ & _22640_ /*60585*/;
assign _22638_ = _21935_ ^ _22640_ /*60588*/;
assign _22639_ = _22631_ & _22638_ /*60586*/;
assign _22384_ = _22631_ ^ _22638_ /*60587*/;
assign _22636_ = _22637_ | _22639_ /*60584*/;
assign _22645_ = ~D[48] /*60583*/;
assign _22642_ = _21936_ & _22645_ /*60579*/;
assign _22643_ = _21936_ ^ _22645_ /*60582*/;
assign _22644_ = _22636_ & _22643_ /*60580*/;
assign _22385_ = _22636_ ^ _22643_ /*60581*/;
assign _22641_ = _22642_ | _22644_ /*60578*/;
assign _22650_ = ~D[49] /*60577*/;
assign _22647_ = _21937_ & _22650_ /*60573*/;
assign _22648_ = _21937_ ^ _22650_ /*60576*/;
assign _22649_ = _22641_ & _22648_ /*60574*/;
assign _22386_ = _22641_ ^ _22648_ /*60575*/;
assign _22646_ = _22647_ | _22649_ /*60572*/;
assign _22655_ = ~D[50] /*60571*/;
assign _22652_ = _21938_ & _22655_ /*60567*/;
assign _22653_ = _21938_ ^ _22655_ /*60570*/;
assign _22654_ = _22646_ & _22653_ /*60568*/;
assign _22387_ = _22646_ ^ _22653_ /*60569*/;
assign _22651_ = _22652_ | _22654_ /*60566*/;
assign _22660_ = ~D[51] /*60565*/;
assign _22657_ = _21939_ & _22660_ /*60561*/;
assign _22658_ = _21939_ ^ _22660_ /*60564*/;
assign _22659_ = _22651_ & _22658_ /*60562*/;
assign _22388_ = _22651_ ^ _22658_ /*60563*/;
assign _22656_ = _22657_ | _22659_ /*60560*/;
assign _22665_ = ~D[52] /*60559*/;
assign _22662_ = _21940_ & _22665_ /*60555*/;
assign _22663_ = _21940_ ^ _22665_ /*60558*/;
assign _22664_ = _22656_ & _22663_ /*60556*/;
assign _22389_ = _22656_ ^ _22663_ /*60557*/;
assign _22661_ = _22662_ | _22664_ /*60554*/;
assign _22670_ = ~D[53] /*60553*/;
assign _22667_ = _21941_ & _22670_ /*60549*/;
assign _22668_ = _21941_ ^ _22670_ /*60552*/;
assign _22669_ = _22661_ & _22668_ /*60550*/;
assign _22390_ = _22661_ ^ _22668_ /*60551*/;
assign _22666_ = _22667_ | _22669_ /*60548*/;
assign _22675_ = ~D[54] /*60547*/;
assign _22672_ = _21942_ & _22675_ /*60543*/;
assign _22673_ = _21942_ ^ _22675_ /*60546*/;
assign _22674_ = _22666_ & _22673_ /*60544*/;
assign _22391_ = _22666_ ^ _22673_ /*60545*/;
assign _22671_ = _22672_ | _22674_ /*60542*/;
assign _22680_ = ~D[55] /*60541*/;
assign _22677_ = _21943_ & _22680_ /*60537*/;
assign _22678_ = _21943_ ^ _22680_ /*60540*/;
assign _22679_ = _22671_ & _22678_ /*60538*/;
assign _22392_ = _22671_ ^ _22678_ /*60539*/;
assign _22676_ = _22677_ | _22679_ /*60536*/;
assign _22685_ = ~D[56] /*60535*/;
assign _22682_ = _21944_ & _22685_ /*60531*/;
assign _22683_ = _21944_ ^ _22685_ /*60534*/;
assign _22684_ = _22676_ & _22683_ /*60532*/;
assign _22393_ = _22676_ ^ _22683_ /*60533*/;
assign _22681_ = _22682_ | _22684_ /*60530*/;
assign _22690_ = ~D[57] /*60529*/;
assign _22687_ = _21945_ & _22690_ /*60525*/;
assign _22688_ = _21945_ ^ _22690_ /*60528*/;
assign _22689_ = _22681_ & _22688_ /*60526*/;
assign _22394_ = _22681_ ^ _22688_ /*60527*/;
assign _22686_ = _22687_ | _22689_ /*60524*/;
assign _22695_ = ~D[58] /*60523*/;
assign _22692_ = _21946_ & _22695_ /*60519*/;
assign _22693_ = _21946_ ^ _22695_ /*60522*/;
assign _22694_ = _22686_ & _22693_ /*60520*/;
assign _22395_ = _22686_ ^ _22693_ /*60521*/;
assign _22691_ = _22692_ | _22694_ /*60518*/;
assign _22700_ = ~D[59] /*60517*/;
assign _22697_ = _21947_ & _22700_ /*60513*/;
assign _22698_ = _21947_ ^ _22700_ /*60516*/;
assign _22699_ = _22691_ & _22698_ /*60514*/;
assign _22396_ = _22691_ ^ _22698_ /*60515*/;
assign _22696_ = _22697_ | _22699_ /*60512*/;
assign _22705_ = ~D[60] /*60511*/;
assign _22702_ = _21948_ & _22705_ /*60507*/;
assign _22703_ = _21948_ ^ _22705_ /*60510*/;
assign _22704_ = _22696_ & _22703_ /*60508*/;
assign _22397_ = _22696_ ^ _22703_ /*60509*/;
assign _22701_ = _22702_ | _22704_ /*60506*/;
assign _22710_ = ~D[61] /*60505*/;
assign _22707_ = _21949_ & _22710_ /*60501*/;
assign _22708_ = _21949_ ^ _22710_ /*60504*/;
assign _22709_ = _22701_ & _22708_ /*60502*/;
assign _22398_ = _22701_ ^ _22708_ /*60503*/;
assign _22706_ = _22707_ | _22709_ /*60500*/;
assign _22715_ = ~D[62] /*60499*/;
assign _22712_ = _21950_ & _22715_ /*60495*/;
assign _22713_ = _21950_ ^ _22715_ /*60498*/;
assign _22714_ = _22706_ & _22713_ /*60496*/;
assign _22399_ = _22706_ ^ _22713_ /*60497*/;
assign _22711_ = _22712_ | _22714_ /*60494*/;
assign _22716_ = _21951_ & oneWire /*60489*/;
assign _22717_ = _21951_ ^ oneWire /*60492*/;
assign _22718_ = _22711_ & _22717_ /*60490*/;
assign _22400_ = _22711_ ^ _22717_ /*60491*/;
assign Q[38] = _22716_ | _22718_ /*60488*/;
assign _22851_ = ~Q[38] /*60103*/;
assign _22850_ = _22851_ & D[0] /*60102*/;
assign _22853_ = _22337_ & _22850_ /*60097*/;
assign _22854_ = _22337_ ^ _22850_ /*60100*/;
assign _22855_ = zeroWire & _22854_ /*60098*/;
assign _22785_ = zeroWire ^ _22854_ /*60099*/;
assign _22852_ = _22853_ | _22855_ /*60096*/;
assign _22857_ = ~Q[38] /*60095*/;
assign _22856_ = _22857_ & D[1] /*60094*/;
assign _22859_ = _22338_ & _22856_ /*60089*/;
assign _22860_ = _22338_ ^ _22856_ /*60092*/;
assign _22861_ = _22852_ & _22860_ /*60090*/;
assign _22786_ = _22852_ ^ _22860_ /*60091*/;
assign _22858_ = _22859_ | _22861_ /*60088*/;
assign _22863_ = ~Q[38] /*60087*/;
assign _22862_ = _22863_ & D[2] /*60086*/;
assign _22865_ = _22339_ & _22862_ /*60081*/;
assign _22866_ = _22339_ ^ _22862_ /*60084*/;
assign _22867_ = _22858_ & _22866_ /*60082*/;
assign _22787_ = _22858_ ^ _22866_ /*60083*/;
assign _22864_ = _22865_ | _22867_ /*60080*/;
assign _22869_ = ~Q[38] /*60079*/;
assign _22868_ = _22869_ & D[3] /*60078*/;
assign _22871_ = _22340_ & _22868_ /*60073*/;
assign _22872_ = _22340_ ^ _22868_ /*60076*/;
assign _22873_ = _22864_ & _22872_ /*60074*/;
assign _22788_ = _22864_ ^ _22872_ /*60075*/;
assign _22870_ = _22871_ | _22873_ /*60072*/;
assign _22875_ = ~Q[38] /*60071*/;
assign _22874_ = _22875_ & D[4] /*60070*/;
assign _22877_ = _22341_ & _22874_ /*60065*/;
assign _22878_ = _22341_ ^ _22874_ /*60068*/;
assign _22879_ = _22870_ & _22878_ /*60066*/;
assign _22789_ = _22870_ ^ _22878_ /*60067*/;
assign _22876_ = _22877_ | _22879_ /*60064*/;
assign _22881_ = ~Q[38] /*60063*/;
assign _22880_ = _22881_ & D[5] /*60062*/;
assign _22883_ = _22342_ & _22880_ /*60057*/;
assign _22884_ = _22342_ ^ _22880_ /*60060*/;
assign _22885_ = _22876_ & _22884_ /*60058*/;
assign _22790_ = _22876_ ^ _22884_ /*60059*/;
assign _22882_ = _22883_ | _22885_ /*60056*/;
assign _22887_ = ~Q[38] /*60055*/;
assign _22886_ = _22887_ & D[6] /*60054*/;
assign _22889_ = _22343_ & _22886_ /*60049*/;
assign _22890_ = _22343_ ^ _22886_ /*60052*/;
assign _22891_ = _22882_ & _22890_ /*60050*/;
assign _22791_ = _22882_ ^ _22890_ /*60051*/;
assign _22888_ = _22889_ | _22891_ /*60048*/;
assign _22893_ = ~Q[38] /*60047*/;
assign _22892_ = _22893_ & D[7] /*60046*/;
assign _22895_ = _22344_ & _22892_ /*60041*/;
assign _22896_ = _22344_ ^ _22892_ /*60044*/;
assign _22897_ = _22888_ & _22896_ /*60042*/;
assign _22792_ = _22888_ ^ _22896_ /*60043*/;
assign _22894_ = _22895_ | _22897_ /*60040*/;
assign _22899_ = ~Q[38] /*60039*/;
assign _22898_ = _22899_ & D[8] /*60038*/;
assign _22901_ = _22345_ & _22898_ /*60033*/;
assign _22902_ = _22345_ ^ _22898_ /*60036*/;
assign _22903_ = _22894_ & _22902_ /*60034*/;
assign _22793_ = _22894_ ^ _22902_ /*60035*/;
assign _22900_ = _22901_ | _22903_ /*60032*/;
assign _22905_ = ~Q[38] /*60031*/;
assign _22904_ = _22905_ & D[9] /*60030*/;
assign _22907_ = _22346_ & _22904_ /*60025*/;
assign _22908_ = _22346_ ^ _22904_ /*60028*/;
assign _22909_ = _22900_ & _22908_ /*60026*/;
assign _22794_ = _22900_ ^ _22908_ /*60027*/;
assign _22906_ = _22907_ | _22909_ /*60024*/;
assign _22911_ = ~Q[38] /*60023*/;
assign _22910_ = _22911_ & D[10] /*60022*/;
assign _22913_ = _22347_ & _22910_ /*60017*/;
assign _22914_ = _22347_ ^ _22910_ /*60020*/;
assign _22915_ = _22906_ & _22914_ /*60018*/;
assign _22795_ = _22906_ ^ _22914_ /*60019*/;
assign _22912_ = _22913_ | _22915_ /*60016*/;
assign _22917_ = ~Q[38] /*60015*/;
assign _22916_ = _22917_ & D[11] /*60014*/;
assign _22919_ = _22348_ & _22916_ /*60009*/;
assign _22920_ = _22348_ ^ _22916_ /*60012*/;
assign _22921_ = _22912_ & _22920_ /*60010*/;
assign _22796_ = _22912_ ^ _22920_ /*60011*/;
assign _22918_ = _22919_ | _22921_ /*60008*/;
assign _22923_ = ~Q[38] /*60007*/;
assign _22922_ = _22923_ & D[12] /*60006*/;
assign _22925_ = _22349_ & _22922_ /*60001*/;
assign _22926_ = _22349_ ^ _22922_ /*60004*/;
assign _22927_ = _22918_ & _22926_ /*60002*/;
assign _22797_ = _22918_ ^ _22926_ /*60003*/;
assign _22924_ = _22925_ | _22927_ /*60000*/;
assign _22929_ = ~Q[38] /*59999*/;
assign _22928_ = _22929_ & D[13] /*59998*/;
assign _22931_ = _22350_ & _22928_ /*59993*/;
assign _22932_ = _22350_ ^ _22928_ /*59996*/;
assign _22933_ = _22924_ & _22932_ /*59994*/;
assign _22798_ = _22924_ ^ _22932_ /*59995*/;
assign _22930_ = _22931_ | _22933_ /*59992*/;
assign _22935_ = ~Q[38] /*59991*/;
assign _22934_ = _22935_ & D[14] /*59990*/;
assign _22937_ = _22351_ & _22934_ /*59985*/;
assign _22938_ = _22351_ ^ _22934_ /*59988*/;
assign _22939_ = _22930_ & _22938_ /*59986*/;
assign _22799_ = _22930_ ^ _22938_ /*59987*/;
assign _22936_ = _22937_ | _22939_ /*59984*/;
assign _22941_ = ~Q[38] /*59983*/;
assign _22940_ = _22941_ & D[15] /*59982*/;
assign _22943_ = _22352_ & _22940_ /*59977*/;
assign _22944_ = _22352_ ^ _22940_ /*59980*/;
assign _22945_ = _22936_ & _22944_ /*59978*/;
assign _22800_ = _22936_ ^ _22944_ /*59979*/;
assign _22942_ = _22943_ | _22945_ /*59976*/;
assign _22947_ = ~Q[38] /*59975*/;
assign _22946_ = _22947_ & D[16] /*59974*/;
assign _22949_ = _22353_ & _22946_ /*59969*/;
assign _22950_ = _22353_ ^ _22946_ /*59972*/;
assign _22951_ = _22942_ & _22950_ /*59970*/;
assign _22801_ = _22942_ ^ _22950_ /*59971*/;
assign _22948_ = _22949_ | _22951_ /*59968*/;
assign _22953_ = ~Q[38] /*59967*/;
assign _22952_ = _22953_ & D[17] /*59966*/;
assign _22955_ = _22354_ & _22952_ /*59961*/;
assign _22956_ = _22354_ ^ _22952_ /*59964*/;
assign _22957_ = _22948_ & _22956_ /*59962*/;
assign _22802_ = _22948_ ^ _22956_ /*59963*/;
assign _22954_ = _22955_ | _22957_ /*59960*/;
assign _22959_ = ~Q[38] /*59959*/;
assign _22958_ = _22959_ & D[18] /*59958*/;
assign _22961_ = _22355_ & _22958_ /*59953*/;
assign _22962_ = _22355_ ^ _22958_ /*59956*/;
assign _22963_ = _22954_ & _22962_ /*59954*/;
assign _22803_ = _22954_ ^ _22962_ /*59955*/;
assign _22960_ = _22961_ | _22963_ /*59952*/;
assign _22965_ = ~Q[38] /*59951*/;
assign _22964_ = _22965_ & D[19] /*59950*/;
assign _22967_ = _22356_ & _22964_ /*59945*/;
assign _22968_ = _22356_ ^ _22964_ /*59948*/;
assign _22969_ = _22960_ & _22968_ /*59946*/;
assign _22804_ = _22960_ ^ _22968_ /*59947*/;
assign _22966_ = _22967_ | _22969_ /*59944*/;
assign _22971_ = ~Q[38] /*59943*/;
assign _22970_ = _22971_ & D[20] /*59942*/;
assign _22973_ = _22357_ & _22970_ /*59937*/;
assign _22974_ = _22357_ ^ _22970_ /*59940*/;
assign _22975_ = _22966_ & _22974_ /*59938*/;
assign _22805_ = _22966_ ^ _22974_ /*59939*/;
assign _22972_ = _22973_ | _22975_ /*59936*/;
assign _22977_ = ~Q[38] /*59935*/;
assign _22976_ = _22977_ & D[21] /*59934*/;
assign _22979_ = _22358_ & _22976_ /*59929*/;
assign _22980_ = _22358_ ^ _22976_ /*59932*/;
assign _22981_ = _22972_ & _22980_ /*59930*/;
assign _22806_ = _22972_ ^ _22980_ /*59931*/;
assign _22978_ = _22979_ | _22981_ /*59928*/;
assign _22983_ = ~Q[38] /*59927*/;
assign _22982_ = _22983_ & D[22] /*59926*/;
assign _22985_ = _22359_ & _22982_ /*59921*/;
assign _22986_ = _22359_ ^ _22982_ /*59924*/;
assign _22987_ = _22978_ & _22986_ /*59922*/;
assign _22807_ = _22978_ ^ _22986_ /*59923*/;
assign _22984_ = _22985_ | _22987_ /*59920*/;
assign _22989_ = ~Q[38] /*59919*/;
assign _22988_ = _22989_ & D[23] /*59918*/;
assign _22991_ = _22360_ & _22988_ /*59913*/;
assign _22992_ = _22360_ ^ _22988_ /*59916*/;
assign _22993_ = _22984_ & _22992_ /*59914*/;
assign _22808_ = _22984_ ^ _22992_ /*59915*/;
assign _22990_ = _22991_ | _22993_ /*59912*/;
assign _22995_ = ~Q[38] /*59911*/;
assign _22994_ = _22995_ & D[24] /*59910*/;
assign _22997_ = _22361_ & _22994_ /*59905*/;
assign _22998_ = _22361_ ^ _22994_ /*59908*/;
assign _22999_ = _22990_ & _22998_ /*59906*/;
assign _22809_ = _22990_ ^ _22998_ /*59907*/;
assign _22996_ = _22997_ | _22999_ /*59904*/;
assign _23001_ = ~Q[38] /*59903*/;
assign _23000_ = _23001_ & D[25] /*59902*/;
assign _23003_ = _22362_ & _23000_ /*59897*/;
assign _23004_ = _22362_ ^ _23000_ /*59900*/;
assign _23005_ = _22996_ & _23004_ /*59898*/;
assign _22810_ = _22996_ ^ _23004_ /*59899*/;
assign _23002_ = _23003_ | _23005_ /*59896*/;
assign _23007_ = ~Q[38] /*59895*/;
assign _23006_ = _23007_ & D[26] /*59894*/;
assign _23009_ = _22363_ & _23006_ /*59889*/;
assign _23010_ = _22363_ ^ _23006_ /*59892*/;
assign _23011_ = _23002_ & _23010_ /*59890*/;
assign _22811_ = _23002_ ^ _23010_ /*59891*/;
assign _23008_ = _23009_ | _23011_ /*59888*/;
assign _23013_ = ~Q[38] /*59887*/;
assign _23012_ = _23013_ & D[27] /*59886*/;
assign _23015_ = _22364_ & _23012_ /*59881*/;
assign _23016_ = _22364_ ^ _23012_ /*59884*/;
assign _23017_ = _23008_ & _23016_ /*59882*/;
assign _22812_ = _23008_ ^ _23016_ /*59883*/;
assign _23014_ = _23015_ | _23017_ /*59880*/;
assign _23019_ = ~Q[38] /*59879*/;
assign _23018_ = _23019_ & D[28] /*59878*/;
assign _23021_ = _22365_ & _23018_ /*59873*/;
assign _23022_ = _22365_ ^ _23018_ /*59876*/;
assign _23023_ = _23014_ & _23022_ /*59874*/;
assign _22813_ = _23014_ ^ _23022_ /*59875*/;
assign _23020_ = _23021_ | _23023_ /*59872*/;
assign _23025_ = ~Q[38] /*59871*/;
assign _23024_ = _23025_ & D[29] /*59870*/;
assign _23027_ = _22366_ & _23024_ /*59865*/;
assign _23028_ = _22366_ ^ _23024_ /*59868*/;
assign _23029_ = _23020_ & _23028_ /*59866*/;
assign _22814_ = _23020_ ^ _23028_ /*59867*/;
assign _23026_ = _23027_ | _23029_ /*59864*/;
assign _23031_ = ~Q[38] /*59863*/;
assign _23030_ = _23031_ & D[30] /*59862*/;
assign _23033_ = _22367_ & _23030_ /*59857*/;
assign _23034_ = _22367_ ^ _23030_ /*59860*/;
assign _23035_ = _23026_ & _23034_ /*59858*/;
assign _22815_ = _23026_ ^ _23034_ /*59859*/;
assign _23032_ = _23033_ | _23035_ /*59856*/;
assign _23037_ = ~Q[38] /*59855*/;
assign _23036_ = _23037_ & D[31] /*59854*/;
assign _23039_ = _22368_ & _23036_ /*59849*/;
assign _23040_ = _22368_ ^ _23036_ /*59852*/;
assign _23041_ = _23032_ & _23040_ /*59850*/;
assign _22816_ = _23032_ ^ _23040_ /*59851*/;
assign _23038_ = _23039_ | _23041_ /*59848*/;
assign _23043_ = ~Q[38] /*59847*/;
assign _23042_ = _23043_ & D[32] /*59846*/;
assign _23045_ = _22369_ & _23042_ /*59841*/;
assign _23046_ = _22369_ ^ _23042_ /*59844*/;
assign _23047_ = _23038_ & _23046_ /*59842*/;
assign _22817_ = _23038_ ^ _23046_ /*59843*/;
assign _23044_ = _23045_ | _23047_ /*59840*/;
assign _23049_ = ~Q[38] /*59839*/;
assign _23048_ = _23049_ & D[33] /*59838*/;
assign _23051_ = _22370_ & _23048_ /*59833*/;
assign _23052_ = _22370_ ^ _23048_ /*59836*/;
assign _23053_ = _23044_ & _23052_ /*59834*/;
assign _22818_ = _23044_ ^ _23052_ /*59835*/;
assign _23050_ = _23051_ | _23053_ /*59832*/;
assign _23055_ = ~Q[38] /*59831*/;
assign _23054_ = _23055_ & D[34] /*59830*/;
assign _23057_ = _22371_ & _23054_ /*59825*/;
assign _23058_ = _22371_ ^ _23054_ /*59828*/;
assign _23059_ = _23050_ & _23058_ /*59826*/;
assign _22819_ = _23050_ ^ _23058_ /*59827*/;
assign _23056_ = _23057_ | _23059_ /*59824*/;
assign _23061_ = ~Q[38] /*59823*/;
assign _23060_ = _23061_ & D[35] /*59822*/;
assign _23063_ = _22372_ & _23060_ /*59817*/;
assign _23064_ = _22372_ ^ _23060_ /*59820*/;
assign _23065_ = _23056_ & _23064_ /*59818*/;
assign _22820_ = _23056_ ^ _23064_ /*59819*/;
assign _23062_ = _23063_ | _23065_ /*59816*/;
assign _23067_ = ~Q[38] /*59815*/;
assign _23066_ = _23067_ & D[36] /*59814*/;
assign _23069_ = _22373_ & _23066_ /*59809*/;
assign _23070_ = _22373_ ^ _23066_ /*59812*/;
assign _23071_ = _23062_ & _23070_ /*59810*/;
assign _22821_ = _23062_ ^ _23070_ /*59811*/;
assign _23068_ = _23069_ | _23071_ /*59808*/;
assign _23073_ = ~Q[38] /*59807*/;
assign _23072_ = _23073_ & D[37] /*59806*/;
assign _23075_ = _22374_ & _23072_ /*59801*/;
assign _23076_ = _22374_ ^ _23072_ /*59804*/;
assign _23077_ = _23068_ & _23076_ /*59802*/;
assign _22822_ = _23068_ ^ _23076_ /*59803*/;
assign _23074_ = _23075_ | _23077_ /*59800*/;
assign _23079_ = ~Q[38] /*59799*/;
assign _23078_ = _23079_ & D[38] /*59798*/;
assign _23081_ = _22375_ & _23078_ /*59793*/;
assign _23082_ = _22375_ ^ _23078_ /*59796*/;
assign _23083_ = _23074_ & _23082_ /*59794*/;
assign _22823_ = _23074_ ^ _23082_ /*59795*/;
assign _23080_ = _23081_ | _23083_ /*59792*/;
assign _23085_ = ~Q[38] /*59791*/;
assign _23084_ = _23085_ & D[39] /*59790*/;
assign _23087_ = _22376_ & _23084_ /*59785*/;
assign _23088_ = _22376_ ^ _23084_ /*59788*/;
assign _23089_ = _23080_ & _23088_ /*59786*/;
assign _22824_ = _23080_ ^ _23088_ /*59787*/;
assign _23086_ = _23087_ | _23089_ /*59784*/;
assign _23091_ = ~Q[38] /*59783*/;
assign _23090_ = _23091_ & D[40] /*59782*/;
assign _23093_ = _22377_ & _23090_ /*59777*/;
assign _23094_ = _22377_ ^ _23090_ /*59780*/;
assign _23095_ = _23086_ & _23094_ /*59778*/;
assign _22825_ = _23086_ ^ _23094_ /*59779*/;
assign _23092_ = _23093_ | _23095_ /*59776*/;
assign _23097_ = ~Q[38] /*59775*/;
assign _23096_ = _23097_ & D[41] /*59774*/;
assign _23099_ = _22378_ & _23096_ /*59769*/;
assign _23100_ = _22378_ ^ _23096_ /*59772*/;
assign _23101_ = _23092_ & _23100_ /*59770*/;
assign _22826_ = _23092_ ^ _23100_ /*59771*/;
assign _23098_ = _23099_ | _23101_ /*59768*/;
assign _23103_ = ~Q[38] /*59767*/;
assign _23102_ = _23103_ & D[42] /*59766*/;
assign _23105_ = _22379_ & _23102_ /*59761*/;
assign _23106_ = _22379_ ^ _23102_ /*59764*/;
assign _23107_ = _23098_ & _23106_ /*59762*/;
assign _22827_ = _23098_ ^ _23106_ /*59763*/;
assign _23104_ = _23105_ | _23107_ /*59760*/;
assign _23109_ = ~Q[38] /*59759*/;
assign _23108_ = _23109_ & D[43] /*59758*/;
assign _23111_ = _22380_ & _23108_ /*59753*/;
assign _23112_ = _22380_ ^ _23108_ /*59756*/;
assign _23113_ = _23104_ & _23112_ /*59754*/;
assign _22828_ = _23104_ ^ _23112_ /*59755*/;
assign _23110_ = _23111_ | _23113_ /*59752*/;
assign _23115_ = ~Q[38] /*59751*/;
assign _23114_ = _23115_ & D[44] /*59750*/;
assign _23117_ = _22381_ & _23114_ /*59745*/;
assign _23118_ = _22381_ ^ _23114_ /*59748*/;
assign _23119_ = _23110_ & _23118_ /*59746*/;
assign _22829_ = _23110_ ^ _23118_ /*59747*/;
assign _23116_ = _23117_ | _23119_ /*59744*/;
assign _23121_ = ~Q[38] /*59743*/;
assign _23120_ = _23121_ & D[45] /*59742*/;
assign _23123_ = _22382_ & _23120_ /*59737*/;
assign _23124_ = _22382_ ^ _23120_ /*59740*/;
assign _23125_ = _23116_ & _23124_ /*59738*/;
assign _22830_ = _23116_ ^ _23124_ /*59739*/;
assign _23122_ = _23123_ | _23125_ /*59736*/;
assign _23127_ = ~Q[38] /*59735*/;
assign _23126_ = _23127_ & D[46] /*59734*/;
assign _23129_ = _22383_ & _23126_ /*59729*/;
assign _23130_ = _22383_ ^ _23126_ /*59732*/;
assign _23131_ = _23122_ & _23130_ /*59730*/;
assign _22831_ = _23122_ ^ _23130_ /*59731*/;
assign _23128_ = _23129_ | _23131_ /*59728*/;
assign _23133_ = ~Q[38] /*59727*/;
assign _23132_ = _23133_ & D[47] /*59726*/;
assign _23135_ = _22384_ & _23132_ /*59721*/;
assign _23136_ = _22384_ ^ _23132_ /*59724*/;
assign _23137_ = _23128_ & _23136_ /*59722*/;
assign _22832_ = _23128_ ^ _23136_ /*59723*/;
assign _23134_ = _23135_ | _23137_ /*59720*/;
assign _23139_ = ~Q[38] /*59719*/;
assign _23138_ = _23139_ & D[48] /*59718*/;
assign _23141_ = _22385_ & _23138_ /*59713*/;
assign _23142_ = _22385_ ^ _23138_ /*59716*/;
assign _23143_ = _23134_ & _23142_ /*59714*/;
assign _22833_ = _23134_ ^ _23142_ /*59715*/;
assign _23140_ = _23141_ | _23143_ /*59712*/;
assign _23145_ = ~Q[38] /*59711*/;
assign _23144_ = _23145_ & D[49] /*59710*/;
assign _23147_ = _22386_ & _23144_ /*59705*/;
assign _23148_ = _22386_ ^ _23144_ /*59708*/;
assign _23149_ = _23140_ & _23148_ /*59706*/;
assign _22834_ = _23140_ ^ _23148_ /*59707*/;
assign _23146_ = _23147_ | _23149_ /*59704*/;
assign _23151_ = ~Q[38] /*59703*/;
assign _23150_ = _23151_ & D[50] /*59702*/;
assign _23153_ = _22387_ & _23150_ /*59697*/;
assign _23154_ = _22387_ ^ _23150_ /*59700*/;
assign _23155_ = _23146_ & _23154_ /*59698*/;
assign _22835_ = _23146_ ^ _23154_ /*59699*/;
assign _23152_ = _23153_ | _23155_ /*59696*/;
assign _23157_ = ~Q[38] /*59695*/;
assign _23156_ = _23157_ & D[51] /*59694*/;
assign _23159_ = _22388_ & _23156_ /*59689*/;
assign _23160_ = _22388_ ^ _23156_ /*59692*/;
assign _23161_ = _23152_ & _23160_ /*59690*/;
assign _22836_ = _23152_ ^ _23160_ /*59691*/;
assign _23158_ = _23159_ | _23161_ /*59688*/;
assign _23163_ = ~Q[38] /*59687*/;
assign _23162_ = _23163_ & D[52] /*59686*/;
assign _23165_ = _22389_ & _23162_ /*59681*/;
assign _23166_ = _22389_ ^ _23162_ /*59684*/;
assign _23167_ = _23158_ & _23166_ /*59682*/;
assign _22837_ = _23158_ ^ _23166_ /*59683*/;
assign _23164_ = _23165_ | _23167_ /*59680*/;
assign _23169_ = ~Q[38] /*59679*/;
assign _23168_ = _23169_ & D[53] /*59678*/;
assign _23171_ = _22390_ & _23168_ /*59673*/;
assign _23172_ = _22390_ ^ _23168_ /*59676*/;
assign _23173_ = _23164_ & _23172_ /*59674*/;
assign _22838_ = _23164_ ^ _23172_ /*59675*/;
assign _23170_ = _23171_ | _23173_ /*59672*/;
assign _23175_ = ~Q[38] /*59671*/;
assign _23174_ = _23175_ & D[54] /*59670*/;
assign _23177_ = _22391_ & _23174_ /*59665*/;
assign _23178_ = _22391_ ^ _23174_ /*59668*/;
assign _23179_ = _23170_ & _23178_ /*59666*/;
assign _22839_ = _23170_ ^ _23178_ /*59667*/;
assign _23176_ = _23177_ | _23179_ /*59664*/;
assign _23181_ = ~Q[38] /*59663*/;
assign _23180_ = _23181_ & D[55] /*59662*/;
assign _23183_ = _22392_ & _23180_ /*59657*/;
assign _23184_ = _22392_ ^ _23180_ /*59660*/;
assign _23185_ = _23176_ & _23184_ /*59658*/;
assign _22840_ = _23176_ ^ _23184_ /*59659*/;
assign _23182_ = _23183_ | _23185_ /*59656*/;
assign _23187_ = ~Q[38] /*59655*/;
assign _23186_ = _23187_ & D[56] /*59654*/;
assign _23189_ = _22393_ & _23186_ /*59649*/;
assign _23190_ = _22393_ ^ _23186_ /*59652*/;
assign _23191_ = _23182_ & _23190_ /*59650*/;
assign _22841_ = _23182_ ^ _23190_ /*59651*/;
assign _23188_ = _23189_ | _23191_ /*59648*/;
assign _23193_ = ~Q[38] /*59647*/;
assign _23192_ = _23193_ & D[57] /*59646*/;
assign _23195_ = _22394_ & _23192_ /*59641*/;
assign _23196_ = _22394_ ^ _23192_ /*59644*/;
assign _23197_ = _23188_ & _23196_ /*59642*/;
assign _22842_ = _23188_ ^ _23196_ /*59643*/;
assign _23194_ = _23195_ | _23197_ /*59640*/;
assign _23199_ = ~Q[38] /*59639*/;
assign _23198_ = _23199_ & D[58] /*59638*/;
assign _23201_ = _22395_ & _23198_ /*59633*/;
assign _23202_ = _22395_ ^ _23198_ /*59636*/;
assign _23203_ = _23194_ & _23202_ /*59634*/;
assign _22843_ = _23194_ ^ _23202_ /*59635*/;
assign _23200_ = _23201_ | _23203_ /*59632*/;
assign _23205_ = ~Q[38] /*59631*/;
assign _23204_ = _23205_ & D[59] /*59630*/;
assign _23207_ = _22396_ & _23204_ /*59625*/;
assign _23208_ = _22396_ ^ _23204_ /*59628*/;
assign _23209_ = _23200_ & _23208_ /*59626*/;
assign _22844_ = _23200_ ^ _23208_ /*59627*/;
assign _23206_ = _23207_ | _23209_ /*59624*/;
assign _23211_ = ~Q[38] /*59623*/;
assign _23210_ = _23211_ & D[60] /*59622*/;
assign _23213_ = _22397_ & _23210_ /*59617*/;
assign _23214_ = _22397_ ^ _23210_ /*59620*/;
assign _23215_ = _23206_ & _23214_ /*59618*/;
assign _22845_ = _23206_ ^ _23214_ /*59619*/;
assign _23212_ = _23213_ | _23215_ /*59616*/;
assign _23217_ = ~Q[38] /*59615*/;
assign _23216_ = _23217_ & D[61] /*59614*/;
assign _23219_ = _22398_ & _23216_ /*59609*/;
assign _23220_ = _22398_ ^ _23216_ /*59612*/;
assign _23221_ = _23212_ & _23220_ /*59610*/;
assign _22846_ = _23212_ ^ _23220_ /*59611*/;
assign _23218_ = _23219_ | _23221_ /*59608*/;
assign _23223_ = ~Q[38] /*59607*/;
assign _23222_ = _23223_ & D[62] /*59606*/;
assign _23225_ = _22399_ & _23222_ /*59601*/;
assign _23226_ = _22399_ ^ _23222_ /*59604*/;
assign _23227_ = _23218_ & _23226_ /*59602*/;
assign _22847_ = _23218_ ^ _23226_ /*59603*/;
assign _23224_ = _23225_ | _23227_ /*59600*/;
assign _23229_ = ~Q[38] /*59599*/;
assign _23228_ = _23229_ & zeroWire /*59598*/;
assign _23230_ = _22400_ ^ _23228_ /*59596*/;
assign _22848_ = _23230_ ^ _23224_ /*59595*/;
assign _23301_ = ~D[0] /*59341*/;
assign _23298_ = R_0[37] & _23301_ /*59337*/;
assign _23299_ = R_0[37] ^ _23301_ /*59340*/;
assign _23300_ = oneWire & _23299_ /*59338*/;
assign _23233_ = oneWire ^ _23299_ /*59339*/;
assign _23297_ = _23298_ | _23300_ /*59336*/;
assign _23306_ = ~D[1] /*59335*/;
assign _23303_ = _22785_ & _23306_ /*59331*/;
assign _23304_ = _22785_ ^ _23306_ /*59334*/;
assign _23305_ = _23297_ & _23304_ /*59332*/;
assign _23234_ = _23297_ ^ _23304_ /*59333*/;
assign _23302_ = _23303_ | _23305_ /*59330*/;
assign _23311_ = ~D[2] /*59329*/;
assign _23308_ = _22786_ & _23311_ /*59325*/;
assign _23309_ = _22786_ ^ _23311_ /*59328*/;
assign _23310_ = _23302_ & _23309_ /*59326*/;
assign _23235_ = _23302_ ^ _23309_ /*59327*/;
assign _23307_ = _23308_ | _23310_ /*59324*/;
assign _23316_ = ~D[3] /*59323*/;
assign _23313_ = _22787_ & _23316_ /*59319*/;
assign _23314_ = _22787_ ^ _23316_ /*59322*/;
assign _23315_ = _23307_ & _23314_ /*59320*/;
assign _23236_ = _23307_ ^ _23314_ /*59321*/;
assign _23312_ = _23313_ | _23315_ /*59318*/;
assign _23321_ = ~D[4] /*59317*/;
assign _23318_ = _22788_ & _23321_ /*59313*/;
assign _23319_ = _22788_ ^ _23321_ /*59316*/;
assign _23320_ = _23312_ & _23319_ /*59314*/;
assign _23237_ = _23312_ ^ _23319_ /*59315*/;
assign _23317_ = _23318_ | _23320_ /*59312*/;
assign _23326_ = ~D[5] /*59311*/;
assign _23323_ = _22789_ & _23326_ /*59307*/;
assign _23324_ = _22789_ ^ _23326_ /*59310*/;
assign _23325_ = _23317_ & _23324_ /*59308*/;
assign _23238_ = _23317_ ^ _23324_ /*59309*/;
assign _23322_ = _23323_ | _23325_ /*59306*/;
assign _23331_ = ~D[6] /*59305*/;
assign _23328_ = _22790_ & _23331_ /*59301*/;
assign _23329_ = _22790_ ^ _23331_ /*59304*/;
assign _23330_ = _23322_ & _23329_ /*59302*/;
assign _23239_ = _23322_ ^ _23329_ /*59303*/;
assign _23327_ = _23328_ | _23330_ /*59300*/;
assign _23336_ = ~D[7] /*59299*/;
assign _23333_ = _22791_ & _23336_ /*59295*/;
assign _23334_ = _22791_ ^ _23336_ /*59298*/;
assign _23335_ = _23327_ & _23334_ /*59296*/;
assign _23240_ = _23327_ ^ _23334_ /*59297*/;
assign _23332_ = _23333_ | _23335_ /*59294*/;
assign _23341_ = ~D[8] /*59293*/;
assign _23338_ = _22792_ & _23341_ /*59289*/;
assign _23339_ = _22792_ ^ _23341_ /*59292*/;
assign _23340_ = _23332_ & _23339_ /*59290*/;
assign _23241_ = _23332_ ^ _23339_ /*59291*/;
assign _23337_ = _23338_ | _23340_ /*59288*/;
assign _23346_ = ~D[9] /*59287*/;
assign _23343_ = _22793_ & _23346_ /*59283*/;
assign _23344_ = _22793_ ^ _23346_ /*59286*/;
assign _23345_ = _23337_ & _23344_ /*59284*/;
assign _23242_ = _23337_ ^ _23344_ /*59285*/;
assign _23342_ = _23343_ | _23345_ /*59282*/;
assign _23351_ = ~D[10] /*59281*/;
assign _23348_ = _22794_ & _23351_ /*59277*/;
assign _23349_ = _22794_ ^ _23351_ /*59280*/;
assign _23350_ = _23342_ & _23349_ /*59278*/;
assign _23243_ = _23342_ ^ _23349_ /*59279*/;
assign _23347_ = _23348_ | _23350_ /*59276*/;
assign _23356_ = ~D[11] /*59275*/;
assign _23353_ = _22795_ & _23356_ /*59271*/;
assign _23354_ = _22795_ ^ _23356_ /*59274*/;
assign _23355_ = _23347_ & _23354_ /*59272*/;
assign _23244_ = _23347_ ^ _23354_ /*59273*/;
assign _23352_ = _23353_ | _23355_ /*59270*/;
assign _23361_ = ~D[12] /*59269*/;
assign _23358_ = _22796_ & _23361_ /*59265*/;
assign _23359_ = _22796_ ^ _23361_ /*59268*/;
assign _23360_ = _23352_ & _23359_ /*59266*/;
assign _23245_ = _23352_ ^ _23359_ /*59267*/;
assign _23357_ = _23358_ | _23360_ /*59264*/;
assign _23366_ = ~D[13] /*59263*/;
assign _23363_ = _22797_ & _23366_ /*59259*/;
assign _23364_ = _22797_ ^ _23366_ /*59262*/;
assign _23365_ = _23357_ & _23364_ /*59260*/;
assign _23246_ = _23357_ ^ _23364_ /*59261*/;
assign _23362_ = _23363_ | _23365_ /*59258*/;
assign _23371_ = ~D[14] /*59257*/;
assign _23368_ = _22798_ & _23371_ /*59253*/;
assign _23369_ = _22798_ ^ _23371_ /*59256*/;
assign _23370_ = _23362_ & _23369_ /*59254*/;
assign _23247_ = _23362_ ^ _23369_ /*59255*/;
assign _23367_ = _23368_ | _23370_ /*59252*/;
assign _23376_ = ~D[15] /*59251*/;
assign _23373_ = _22799_ & _23376_ /*59247*/;
assign _23374_ = _22799_ ^ _23376_ /*59250*/;
assign _23375_ = _23367_ & _23374_ /*59248*/;
assign _23248_ = _23367_ ^ _23374_ /*59249*/;
assign _23372_ = _23373_ | _23375_ /*59246*/;
assign _23381_ = ~D[16] /*59245*/;
assign _23378_ = _22800_ & _23381_ /*59241*/;
assign _23379_ = _22800_ ^ _23381_ /*59244*/;
assign _23380_ = _23372_ & _23379_ /*59242*/;
assign _23249_ = _23372_ ^ _23379_ /*59243*/;
assign _23377_ = _23378_ | _23380_ /*59240*/;
assign _23386_ = ~D[17] /*59239*/;
assign _23383_ = _22801_ & _23386_ /*59235*/;
assign _23384_ = _22801_ ^ _23386_ /*59238*/;
assign _23385_ = _23377_ & _23384_ /*59236*/;
assign _23250_ = _23377_ ^ _23384_ /*59237*/;
assign _23382_ = _23383_ | _23385_ /*59234*/;
assign _23391_ = ~D[18] /*59233*/;
assign _23388_ = _22802_ & _23391_ /*59229*/;
assign _23389_ = _22802_ ^ _23391_ /*59232*/;
assign _23390_ = _23382_ & _23389_ /*59230*/;
assign _23251_ = _23382_ ^ _23389_ /*59231*/;
assign _23387_ = _23388_ | _23390_ /*59228*/;
assign _23396_ = ~D[19] /*59227*/;
assign _23393_ = _22803_ & _23396_ /*59223*/;
assign _23394_ = _22803_ ^ _23396_ /*59226*/;
assign _23395_ = _23387_ & _23394_ /*59224*/;
assign _23252_ = _23387_ ^ _23394_ /*59225*/;
assign _23392_ = _23393_ | _23395_ /*59222*/;
assign _23401_ = ~D[20] /*59221*/;
assign _23398_ = _22804_ & _23401_ /*59217*/;
assign _23399_ = _22804_ ^ _23401_ /*59220*/;
assign _23400_ = _23392_ & _23399_ /*59218*/;
assign _23253_ = _23392_ ^ _23399_ /*59219*/;
assign _23397_ = _23398_ | _23400_ /*59216*/;
assign _23406_ = ~D[21] /*59215*/;
assign _23403_ = _22805_ & _23406_ /*59211*/;
assign _23404_ = _22805_ ^ _23406_ /*59214*/;
assign _23405_ = _23397_ & _23404_ /*59212*/;
assign _23254_ = _23397_ ^ _23404_ /*59213*/;
assign _23402_ = _23403_ | _23405_ /*59210*/;
assign _23411_ = ~D[22] /*59209*/;
assign _23408_ = _22806_ & _23411_ /*59205*/;
assign _23409_ = _22806_ ^ _23411_ /*59208*/;
assign _23410_ = _23402_ & _23409_ /*59206*/;
assign _23255_ = _23402_ ^ _23409_ /*59207*/;
assign _23407_ = _23408_ | _23410_ /*59204*/;
assign _23416_ = ~D[23] /*59203*/;
assign _23413_ = _22807_ & _23416_ /*59199*/;
assign _23414_ = _22807_ ^ _23416_ /*59202*/;
assign _23415_ = _23407_ & _23414_ /*59200*/;
assign _23256_ = _23407_ ^ _23414_ /*59201*/;
assign _23412_ = _23413_ | _23415_ /*59198*/;
assign _23421_ = ~D[24] /*59197*/;
assign _23418_ = _22808_ & _23421_ /*59193*/;
assign _23419_ = _22808_ ^ _23421_ /*59196*/;
assign _23420_ = _23412_ & _23419_ /*59194*/;
assign _23257_ = _23412_ ^ _23419_ /*59195*/;
assign _23417_ = _23418_ | _23420_ /*59192*/;
assign _23426_ = ~D[25] /*59191*/;
assign _23423_ = _22809_ & _23426_ /*59187*/;
assign _23424_ = _22809_ ^ _23426_ /*59190*/;
assign _23425_ = _23417_ & _23424_ /*59188*/;
assign _23258_ = _23417_ ^ _23424_ /*59189*/;
assign _23422_ = _23423_ | _23425_ /*59186*/;
assign _23431_ = ~D[26] /*59185*/;
assign _23428_ = _22810_ & _23431_ /*59181*/;
assign _23429_ = _22810_ ^ _23431_ /*59184*/;
assign _23430_ = _23422_ & _23429_ /*59182*/;
assign _23259_ = _23422_ ^ _23429_ /*59183*/;
assign _23427_ = _23428_ | _23430_ /*59180*/;
assign _23436_ = ~D[27] /*59179*/;
assign _23433_ = _22811_ & _23436_ /*59175*/;
assign _23434_ = _22811_ ^ _23436_ /*59178*/;
assign _23435_ = _23427_ & _23434_ /*59176*/;
assign _23260_ = _23427_ ^ _23434_ /*59177*/;
assign _23432_ = _23433_ | _23435_ /*59174*/;
assign _23441_ = ~D[28] /*59173*/;
assign _23438_ = _22812_ & _23441_ /*59169*/;
assign _23439_ = _22812_ ^ _23441_ /*59172*/;
assign _23440_ = _23432_ & _23439_ /*59170*/;
assign _23261_ = _23432_ ^ _23439_ /*59171*/;
assign _23437_ = _23438_ | _23440_ /*59168*/;
assign _23446_ = ~D[29] /*59167*/;
assign _23443_ = _22813_ & _23446_ /*59163*/;
assign _23444_ = _22813_ ^ _23446_ /*59166*/;
assign _23445_ = _23437_ & _23444_ /*59164*/;
assign _23262_ = _23437_ ^ _23444_ /*59165*/;
assign _23442_ = _23443_ | _23445_ /*59162*/;
assign _23451_ = ~D[30] /*59161*/;
assign _23448_ = _22814_ & _23451_ /*59157*/;
assign _23449_ = _22814_ ^ _23451_ /*59160*/;
assign _23450_ = _23442_ & _23449_ /*59158*/;
assign _23263_ = _23442_ ^ _23449_ /*59159*/;
assign _23447_ = _23448_ | _23450_ /*59156*/;
assign _23456_ = ~D[31] /*59155*/;
assign _23453_ = _22815_ & _23456_ /*59151*/;
assign _23454_ = _22815_ ^ _23456_ /*59154*/;
assign _23455_ = _23447_ & _23454_ /*59152*/;
assign _23264_ = _23447_ ^ _23454_ /*59153*/;
assign _23452_ = _23453_ | _23455_ /*59150*/;
assign _23461_ = ~D[32] /*59149*/;
assign _23458_ = _22816_ & _23461_ /*59145*/;
assign _23459_ = _22816_ ^ _23461_ /*59148*/;
assign _23460_ = _23452_ & _23459_ /*59146*/;
assign _23265_ = _23452_ ^ _23459_ /*59147*/;
assign _23457_ = _23458_ | _23460_ /*59144*/;
assign _23466_ = ~D[33] /*59143*/;
assign _23463_ = _22817_ & _23466_ /*59139*/;
assign _23464_ = _22817_ ^ _23466_ /*59142*/;
assign _23465_ = _23457_ & _23464_ /*59140*/;
assign _23266_ = _23457_ ^ _23464_ /*59141*/;
assign _23462_ = _23463_ | _23465_ /*59138*/;
assign _23471_ = ~D[34] /*59137*/;
assign _23468_ = _22818_ & _23471_ /*59133*/;
assign _23469_ = _22818_ ^ _23471_ /*59136*/;
assign _23470_ = _23462_ & _23469_ /*59134*/;
assign _23267_ = _23462_ ^ _23469_ /*59135*/;
assign _23467_ = _23468_ | _23470_ /*59132*/;
assign _23476_ = ~D[35] /*59131*/;
assign _23473_ = _22819_ & _23476_ /*59127*/;
assign _23474_ = _22819_ ^ _23476_ /*59130*/;
assign _23475_ = _23467_ & _23474_ /*59128*/;
assign _23268_ = _23467_ ^ _23474_ /*59129*/;
assign _23472_ = _23473_ | _23475_ /*59126*/;
assign _23481_ = ~D[36] /*59125*/;
assign _23478_ = _22820_ & _23481_ /*59121*/;
assign _23479_ = _22820_ ^ _23481_ /*59124*/;
assign _23480_ = _23472_ & _23479_ /*59122*/;
assign _23269_ = _23472_ ^ _23479_ /*59123*/;
assign _23477_ = _23478_ | _23480_ /*59120*/;
assign _23486_ = ~D[37] /*59119*/;
assign _23483_ = _22821_ & _23486_ /*59115*/;
assign _23484_ = _22821_ ^ _23486_ /*59118*/;
assign _23485_ = _23477_ & _23484_ /*59116*/;
assign _23270_ = _23477_ ^ _23484_ /*59117*/;
assign _23482_ = _23483_ | _23485_ /*59114*/;
assign _23491_ = ~D[38] /*59113*/;
assign _23488_ = _22822_ & _23491_ /*59109*/;
assign _23489_ = _22822_ ^ _23491_ /*59112*/;
assign _23490_ = _23482_ & _23489_ /*59110*/;
assign _23271_ = _23482_ ^ _23489_ /*59111*/;
assign _23487_ = _23488_ | _23490_ /*59108*/;
assign _23496_ = ~D[39] /*59107*/;
assign _23493_ = _22823_ & _23496_ /*59103*/;
assign _23494_ = _22823_ ^ _23496_ /*59106*/;
assign _23495_ = _23487_ & _23494_ /*59104*/;
assign _23272_ = _23487_ ^ _23494_ /*59105*/;
assign _23492_ = _23493_ | _23495_ /*59102*/;
assign _23501_ = ~D[40] /*59101*/;
assign _23498_ = _22824_ & _23501_ /*59097*/;
assign _23499_ = _22824_ ^ _23501_ /*59100*/;
assign _23500_ = _23492_ & _23499_ /*59098*/;
assign _23273_ = _23492_ ^ _23499_ /*59099*/;
assign _23497_ = _23498_ | _23500_ /*59096*/;
assign _23506_ = ~D[41] /*59095*/;
assign _23503_ = _22825_ & _23506_ /*59091*/;
assign _23504_ = _22825_ ^ _23506_ /*59094*/;
assign _23505_ = _23497_ & _23504_ /*59092*/;
assign _23274_ = _23497_ ^ _23504_ /*59093*/;
assign _23502_ = _23503_ | _23505_ /*59090*/;
assign _23511_ = ~D[42] /*59089*/;
assign _23508_ = _22826_ & _23511_ /*59085*/;
assign _23509_ = _22826_ ^ _23511_ /*59088*/;
assign _23510_ = _23502_ & _23509_ /*59086*/;
assign _23275_ = _23502_ ^ _23509_ /*59087*/;
assign _23507_ = _23508_ | _23510_ /*59084*/;
assign _23516_ = ~D[43] /*59083*/;
assign _23513_ = _22827_ & _23516_ /*59079*/;
assign _23514_ = _22827_ ^ _23516_ /*59082*/;
assign _23515_ = _23507_ & _23514_ /*59080*/;
assign _23276_ = _23507_ ^ _23514_ /*59081*/;
assign _23512_ = _23513_ | _23515_ /*59078*/;
assign _23521_ = ~D[44] /*59077*/;
assign _23518_ = _22828_ & _23521_ /*59073*/;
assign _23519_ = _22828_ ^ _23521_ /*59076*/;
assign _23520_ = _23512_ & _23519_ /*59074*/;
assign _23277_ = _23512_ ^ _23519_ /*59075*/;
assign _23517_ = _23518_ | _23520_ /*59072*/;
assign _23526_ = ~D[45] /*59071*/;
assign _23523_ = _22829_ & _23526_ /*59067*/;
assign _23524_ = _22829_ ^ _23526_ /*59070*/;
assign _23525_ = _23517_ & _23524_ /*59068*/;
assign _23278_ = _23517_ ^ _23524_ /*59069*/;
assign _23522_ = _23523_ | _23525_ /*59066*/;
assign _23531_ = ~D[46] /*59065*/;
assign _23528_ = _22830_ & _23531_ /*59061*/;
assign _23529_ = _22830_ ^ _23531_ /*59064*/;
assign _23530_ = _23522_ & _23529_ /*59062*/;
assign _23279_ = _23522_ ^ _23529_ /*59063*/;
assign _23527_ = _23528_ | _23530_ /*59060*/;
assign _23536_ = ~D[47] /*59059*/;
assign _23533_ = _22831_ & _23536_ /*59055*/;
assign _23534_ = _22831_ ^ _23536_ /*59058*/;
assign _23535_ = _23527_ & _23534_ /*59056*/;
assign _23280_ = _23527_ ^ _23534_ /*59057*/;
assign _23532_ = _23533_ | _23535_ /*59054*/;
assign _23541_ = ~D[48] /*59053*/;
assign _23538_ = _22832_ & _23541_ /*59049*/;
assign _23539_ = _22832_ ^ _23541_ /*59052*/;
assign _23540_ = _23532_ & _23539_ /*59050*/;
assign _23281_ = _23532_ ^ _23539_ /*59051*/;
assign _23537_ = _23538_ | _23540_ /*59048*/;
assign _23546_ = ~D[49] /*59047*/;
assign _23543_ = _22833_ & _23546_ /*59043*/;
assign _23544_ = _22833_ ^ _23546_ /*59046*/;
assign _23545_ = _23537_ & _23544_ /*59044*/;
assign _23282_ = _23537_ ^ _23544_ /*59045*/;
assign _23542_ = _23543_ | _23545_ /*59042*/;
assign _23551_ = ~D[50] /*59041*/;
assign _23548_ = _22834_ & _23551_ /*59037*/;
assign _23549_ = _22834_ ^ _23551_ /*59040*/;
assign _23550_ = _23542_ & _23549_ /*59038*/;
assign _23283_ = _23542_ ^ _23549_ /*59039*/;
assign _23547_ = _23548_ | _23550_ /*59036*/;
assign _23556_ = ~D[51] /*59035*/;
assign _23553_ = _22835_ & _23556_ /*59031*/;
assign _23554_ = _22835_ ^ _23556_ /*59034*/;
assign _23555_ = _23547_ & _23554_ /*59032*/;
assign _23284_ = _23547_ ^ _23554_ /*59033*/;
assign _23552_ = _23553_ | _23555_ /*59030*/;
assign _23561_ = ~D[52] /*59029*/;
assign _23558_ = _22836_ & _23561_ /*59025*/;
assign _23559_ = _22836_ ^ _23561_ /*59028*/;
assign _23560_ = _23552_ & _23559_ /*59026*/;
assign _23285_ = _23552_ ^ _23559_ /*59027*/;
assign _23557_ = _23558_ | _23560_ /*59024*/;
assign _23566_ = ~D[53] /*59023*/;
assign _23563_ = _22837_ & _23566_ /*59019*/;
assign _23564_ = _22837_ ^ _23566_ /*59022*/;
assign _23565_ = _23557_ & _23564_ /*59020*/;
assign _23286_ = _23557_ ^ _23564_ /*59021*/;
assign _23562_ = _23563_ | _23565_ /*59018*/;
assign _23571_ = ~D[54] /*59017*/;
assign _23568_ = _22838_ & _23571_ /*59013*/;
assign _23569_ = _22838_ ^ _23571_ /*59016*/;
assign _23570_ = _23562_ & _23569_ /*59014*/;
assign _23287_ = _23562_ ^ _23569_ /*59015*/;
assign _23567_ = _23568_ | _23570_ /*59012*/;
assign _23576_ = ~D[55] /*59011*/;
assign _23573_ = _22839_ & _23576_ /*59007*/;
assign _23574_ = _22839_ ^ _23576_ /*59010*/;
assign _23575_ = _23567_ & _23574_ /*59008*/;
assign _23288_ = _23567_ ^ _23574_ /*59009*/;
assign _23572_ = _23573_ | _23575_ /*59006*/;
assign _23581_ = ~D[56] /*59005*/;
assign _23578_ = _22840_ & _23581_ /*59001*/;
assign _23579_ = _22840_ ^ _23581_ /*59004*/;
assign _23580_ = _23572_ & _23579_ /*59002*/;
assign _23289_ = _23572_ ^ _23579_ /*59003*/;
assign _23577_ = _23578_ | _23580_ /*59000*/;
assign _23586_ = ~D[57] /*58999*/;
assign _23583_ = _22841_ & _23586_ /*58995*/;
assign _23584_ = _22841_ ^ _23586_ /*58998*/;
assign _23585_ = _23577_ & _23584_ /*58996*/;
assign _23290_ = _23577_ ^ _23584_ /*58997*/;
assign _23582_ = _23583_ | _23585_ /*58994*/;
assign _23591_ = ~D[58] /*58993*/;
assign _23588_ = _22842_ & _23591_ /*58989*/;
assign _23589_ = _22842_ ^ _23591_ /*58992*/;
assign _23590_ = _23582_ & _23589_ /*58990*/;
assign _23291_ = _23582_ ^ _23589_ /*58991*/;
assign _23587_ = _23588_ | _23590_ /*58988*/;
assign _23596_ = ~D[59] /*58987*/;
assign _23593_ = _22843_ & _23596_ /*58983*/;
assign _23594_ = _22843_ ^ _23596_ /*58986*/;
assign _23595_ = _23587_ & _23594_ /*58984*/;
assign _23292_ = _23587_ ^ _23594_ /*58985*/;
assign _23592_ = _23593_ | _23595_ /*58982*/;
assign _23601_ = ~D[60] /*58981*/;
assign _23598_ = _22844_ & _23601_ /*58977*/;
assign _23599_ = _22844_ ^ _23601_ /*58980*/;
assign _23600_ = _23592_ & _23599_ /*58978*/;
assign _23293_ = _23592_ ^ _23599_ /*58979*/;
assign _23597_ = _23598_ | _23600_ /*58976*/;
assign _23606_ = ~D[61] /*58975*/;
assign _23603_ = _22845_ & _23606_ /*58971*/;
assign _23604_ = _22845_ ^ _23606_ /*58974*/;
assign _23605_ = _23597_ & _23604_ /*58972*/;
assign _23294_ = _23597_ ^ _23604_ /*58973*/;
assign _23602_ = _23603_ | _23605_ /*58970*/;
assign _23611_ = ~D[62] /*58969*/;
assign _23608_ = _22846_ & _23611_ /*58965*/;
assign _23609_ = _22846_ ^ _23611_ /*58968*/;
assign _23610_ = _23602_ & _23609_ /*58966*/;
assign _23295_ = _23602_ ^ _23609_ /*58967*/;
assign _23607_ = _23608_ | _23610_ /*58964*/;
assign _23612_ = _22847_ & oneWire /*58959*/;
assign _23613_ = _22847_ ^ oneWire /*58962*/;
assign _23614_ = _23607_ & _23613_ /*58960*/;
assign _23296_ = _23607_ ^ _23613_ /*58961*/;
assign Q[37] = _23612_ | _23614_ /*58958*/;
assign _23747_ = ~Q[37] /*58573*/;
assign _23746_ = _23747_ & D[0] /*58572*/;
assign _23749_ = _23233_ & _23746_ /*58567*/;
assign _23750_ = _23233_ ^ _23746_ /*58570*/;
assign _23751_ = zeroWire & _23750_ /*58568*/;
assign _23681_ = zeroWire ^ _23750_ /*58569*/;
assign _23748_ = _23749_ | _23751_ /*58566*/;
assign _23753_ = ~Q[37] /*58565*/;
assign _23752_ = _23753_ & D[1] /*58564*/;
assign _23755_ = _23234_ & _23752_ /*58559*/;
assign _23756_ = _23234_ ^ _23752_ /*58562*/;
assign _23757_ = _23748_ & _23756_ /*58560*/;
assign _23682_ = _23748_ ^ _23756_ /*58561*/;
assign _23754_ = _23755_ | _23757_ /*58558*/;
assign _23759_ = ~Q[37] /*58557*/;
assign _23758_ = _23759_ & D[2] /*58556*/;
assign _23761_ = _23235_ & _23758_ /*58551*/;
assign _23762_ = _23235_ ^ _23758_ /*58554*/;
assign _23763_ = _23754_ & _23762_ /*58552*/;
assign _23683_ = _23754_ ^ _23762_ /*58553*/;
assign _23760_ = _23761_ | _23763_ /*58550*/;
assign _23765_ = ~Q[37] /*58549*/;
assign _23764_ = _23765_ & D[3] /*58548*/;
assign _23767_ = _23236_ & _23764_ /*58543*/;
assign _23768_ = _23236_ ^ _23764_ /*58546*/;
assign _23769_ = _23760_ & _23768_ /*58544*/;
assign _23684_ = _23760_ ^ _23768_ /*58545*/;
assign _23766_ = _23767_ | _23769_ /*58542*/;
assign _23771_ = ~Q[37] /*58541*/;
assign _23770_ = _23771_ & D[4] /*58540*/;
assign _23773_ = _23237_ & _23770_ /*58535*/;
assign _23774_ = _23237_ ^ _23770_ /*58538*/;
assign _23775_ = _23766_ & _23774_ /*58536*/;
assign _23685_ = _23766_ ^ _23774_ /*58537*/;
assign _23772_ = _23773_ | _23775_ /*58534*/;
assign _23777_ = ~Q[37] /*58533*/;
assign _23776_ = _23777_ & D[5] /*58532*/;
assign _23779_ = _23238_ & _23776_ /*58527*/;
assign _23780_ = _23238_ ^ _23776_ /*58530*/;
assign _23781_ = _23772_ & _23780_ /*58528*/;
assign _23686_ = _23772_ ^ _23780_ /*58529*/;
assign _23778_ = _23779_ | _23781_ /*58526*/;
assign _23783_ = ~Q[37] /*58525*/;
assign _23782_ = _23783_ & D[6] /*58524*/;
assign _23785_ = _23239_ & _23782_ /*58519*/;
assign _23786_ = _23239_ ^ _23782_ /*58522*/;
assign _23787_ = _23778_ & _23786_ /*58520*/;
assign _23687_ = _23778_ ^ _23786_ /*58521*/;
assign _23784_ = _23785_ | _23787_ /*58518*/;
assign _23789_ = ~Q[37] /*58517*/;
assign _23788_ = _23789_ & D[7] /*58516*/;
assign _23791_ = _23240_ & _23788_ /*58511*/;
assign _23792_ = _23240_ ^ _23788_ /*58514*/;
assign _23793_ = _23784_ & _23792_ /*58512*/;
assign _23688_ = _23784_ ^ _23792_ /*58513*/;
assign _23790_ = _23791_ | _23793_ /*58510*/;
assign _23795_ = ~Q[37] /*58509*/;
assign _23794_ = _23795_ & D[8] /*58508*/;
assign _23797_ = _23241_ & _23794_ /*58503*/;
assign _23798_ = _23241_ ^ _23794_ /*58506*/;
assign _23799_ = _23790_ & _23798_ /*58504*/;
assign _23689_ = _23790_ ^ _23798_ /*58505*/;
assign _23796_ = _23797_ | _23799_ /*58502*/;
assign _23801_ = ~Q[37] /*58501*/;
assign _23800_ = _23801_ & D[9] /*58500*/;
assign _23803_ = _23242_ & _23800_ /*58495*/;
assign _23804_ = _23242_ ^ _23800_ /*58498*/;
assign _23805_ = _23796_ & _23804_ /*58496*/;
assign _23690_ = _23796_ ^ _23804_ /*58497*/;
assign _23802_ = _23803_ | _23805_ /*58494*/;
assign _23807_ = ~Q[37] /*58493*/;
assign _23806_ = _23807_ & D[10] /*58492*/;
assign _23809_ = _23243_ & _23806_ /*58487*/;
assign _23810_ = _23243_ ^ _23806_ /*58490*/;
assign _23811_ = _23802_ & _23810_ /*58488*/;
assign _23691_ = _23802_ ^ _23810_ /*58489*/;
assign _23808_ = _23809_ | _23811_ /*58486*/;
assign _23813_ = ~Q[37] /*58485*/;
assign _23812_ = _23813_ & D[11] /*58484*/;
assign _23815_ = _23244_ & _23812_ /*58479*/;
assign _23816_ = _23244_ ^ _23812_ /*58482*/;
assign _23817_ = _23808_ & _23816_ /*58480*/;
assign _23692_ = _23808_ ^ _23816_ /*58481*/;
assign _23814_ = _23815_ | _23817_ /*58478*/;
assign _23819_ = ~Q[37] /*58477*/;
assign _23818_ = _23819_ & D[12] /*58476*/;
assign _23821_ = _23245_ & _23818_ /*58471*/;
assign _23822_ = _23245_ ^ _23818_ /*58474*/;
assign _23823_ = _23814_ & _23822_ /*58472*/;
assign _23693_ = _23814_ ^ _23822_ /*58473*/;
assign _23820_ = _23821_ | _23823_ /*58470*/;
assign _23825_ = ~Q[37] /*58469*/;
assign _23824_ = _23825_ & D[13] /*58468*/;
assign _23827_ = _23246_ & _23824_ /*58463*/;
assign _23828_ = _23246_ ^ _23824_ /*58466*/;
assign _23829_ = _23820_ & _23828_ /*58464*/;
assign _23694_ = _23820_ ^ _23828_ /*58465*/;
assign _23826_ = _23827_ | _23829_ /*58462*/;
assign _23831_ = ~Q[37] /*58461*/;
assign _23830_ = _23831_ & D[14] /*58460*/;
assign _23833_ = _23247_ & _23830_ /*58455*/;
assign _23834_ = _23247_ ^ _23830_ /*58458*/;
assign _23835_ = _23826_ & _23834_ /*58456*/;
assign _23695_ = _23826_ ^ _23834_ /*58457*/;
assign _23832_ = _23833_ | _23835_ /*58454*/;
assign _23837_ = ~Q[37] /*58453*/;
assign _23836_ = _23837_ & D[15] /*58452*/;
assign _23839_ = _23248_ & _23836_ /*58447*/;
assign _23840_ = _23248_ ^ _23836_ /*58450*/;
assign _23841_ = _23832_ & _23840_ /*58448*/;
assign _23696_ = _23832_ ^ _23840_ /*58449*/;
assign _23838_ = _23839_ | _23841_ /*58446*/;
assign _23843_ = ~Q[37] /*58445*/;
assign _23842_ = _23843_ & D[16] /*58444*/;
assign _23845_ = _23249_ & _23842_ /*58439*/;
assign _23846_ = _23249_ ^ _23842_ /*58442*/;
assign _23847_ = _23838_ & _23846_ /*58440*/;
assign _23697_ = _23838_ ^ _23846_ /*58441*/;
assign _23844_ = _23845_ | _23847_ /*58438*/;
assign _23849_ = ~Q[37] /*58437*/;
assign _23848_ = _23849_ & D[17] /*58436*/;
assign _23851_ = _23250_ & _23848_ /*58431*/;
assign _23852_ = _23250_ ^ _23848_ /*58434*/;
assign _23853_ = _23844_ & _23852_ /*58432*/;
assign _23698_ = _23844_ ^ _23852_ /*58433*/;
assign _23850_ = _23851_ | _23853_ /*58430*/;
assign _23855_ = ~Q[37] /*58429*/;
assign _23854_ = _23855_ & D[18] /*58428*/;
assign _23857_ = _23251_ & _23854_ /*58423*/;
assign _23858_ = _23251_ ^ _23854_ /*58426*/;
assign _23859_ = _23850_ & _23858_ /*58424*/;
assign _23699_ = _23850_ ^ _23858_ /*58425*/;
assign _23856_ = _23857_ | _23859_ /*58422*/;
assign _23861_ = ~Q[37] /*58421*/;
assign _23860_ = _23861_ & D[19] /*58420*/;
assign _23863_ = _23252_ & _23860_ /*58415*/;
assign _23864_ = _23252_ ^ _23860_ /*58418*/;
assign _23865_ = _23856_ & _23864_ /*58416*/;
assign _23700_ = _23856_ ^ _23864_ /*58417*/;
assign _23862_ = _23863_ | _23865_ /*58414*/;
assign _23867_ = ~Q[37] /*58413*/;
assign _23866_ = _23867_ & D[20] /*58412*/;
assign _23869_ = _23253_ & _23866_ /*58407*/;
assign _23870_ = _23253_ ^ _23866_ /*58410*/;
assign _23871_ = _23862_ & _23870_ /*58408*/;
assign _23701_ = _23862_ ^ _23870_ /*58409*/;
assign _23868_ = _23869_ | _23871_ /*58406*/;
assign _23873_ = ~Q[37] /*58405*/;
assign _23872_ = _23873_ & D[21] /*58404*/;
assign _23875_ = _23254_ & _23872_ /*58399*/;
assign _23876_ = _23254_ ^ _23872_ /*58402*/;
assign _23877_ = _23868_ & _23876_ /*58400*/;
assign _23702_ = _23868_ ^ _23876_ /*58401*/;
assign _23874_ = _23875_ | _23877_ /*58398*/;
assign _23879_ = ~Q[37] /*58397*/;
assign _23878_ = _23879_ & D[22] /*58396*/;
assign _23881_ = _23255_ & _23878_ /*58391*/;
assign _23882_ = _23255_ ^ _23878_ /*58394*/;
assign _23883_ = _23874_ & _23882_ /*58392*/;
assign _23703_ = _23874_ ^ _23882_ /*58393*/;
assign _23880_ = _23881_ | _23883_ /*58390*/;
assign _23885_ = ~Q[37] /*58389*/;
assign _23884_ = _23885_ & D[23] /*58388*/;
assign _23887_ = _23256_ & _23884_ /*58383*/;
assign _23888_ = _23256_ ^ _23884_ /*58386*/;
assign _23889_ = _23880_ & _23888_ /*58384*/;
assign _23704_ = _23880_ ^ _23888_ /*58385*/;
assign _23886_ = _23887_ | _23889_ /*58382*/;
assign _23891_ = ~Q[37] /*58381*/;
assign _23890_ = _23891_ & D[24] /*58380*/;
assign _23893_ = _23257_ & _23890_ /*58375*/;
assign _23894_ = _23257_ ^ _23890_ /*58378*/;
assign _23895_ = _23886_ & _23894_ /*58376*/;
assign _23705_ = _23886_ ^ _23894_ /*58377*/;
assign _23892_ = _23893_ | _23895_ /*58374*/;
assign _23897_ = ~Q[37] /*58373*/;
assign _23896_ = _23897_ & D[25] /*58372*/;
assign _23899_ = _23258_ & _23896_ /*58367*/;
assign _23900_ = _23258_ ^ _23896_ /*58370*/;
assign _23901_ = _23892_ & _23900_ /*58368*/;
assign _23706_ = _23892_ ^ _23900_ /*58369*/;
assign _23898_ = _23899_ | _23901_ /*58366*/;
assign _23903_ = ~Q[37] /*58365*/;
assign _23902_ = _23903_ & D[26] /*58364*/;
assign _23905_ = _23259_ & _23902_ /*58359*/;
assign _23906_ = _23259_ ^ _23902_ /*58362*/;
assign _23907_ = _23898_ & _23906_ /*58360*/;
assign _23707_ = _23898_ ^ _23906_ /*58361*/;
assign _23904_ = _23905_ | _23907_ /*58358*/;
assign _23909_ = ~Q[37] /*58357*/;
assign _23908_ = _23909_ & D[27] /*58356*/;
assign _23911_ = _23260_ & _23908_ /*58351*/;
assign _23912_ = _23260_ ^ _23908_ /*58354*/;
assign _23913_ = _23904_ & _23912_ /*58352*/;
assign _23708_ = _23904_ ^ _23912_ /*58353*/;
assign _23910_ = _23911_ | _23913_ /*58350*/;
assign _23915_ = ~Q[37] /*58349*/;
assign _23914_ = _23915_ & D[28] /*58348*/;
assign _23917_ = _23261_ & _23914_ /*58343*/;
assign _23918_ = _23261_ ^ _23914_ /*58346*/;
assign _23919_ = _23910_ & _23918_ /*58344*/;
assign _23709_ = _23910_ ^ _23918_ /*58345*/;
assign _23916_ = _23917_ | _23919_ /*58342*/;
assign _23921_ = ~Q[37] /*58341*/;
assign _23920_ = _23921_ & D[29] /*58340*/;
assign _23923_ = _23262_ & _23920_ /*58335*/;
assign _23924_ = _23262_ ^ _23920_ /*58338*/;
assign _23925_ = _23916_ & _23924_ /*58336*/;
assign _23710_ = _23916_ ^ _23924_ /*58337*/;
assign _23922_ = _23923_ | _23925_ /*58334*/;
assign _23927_ = ~Q[37] /*58333*/;
assign _23926_ = _23927_ & D[30] /*58332*/;
assign _23929_ = _23263_ & _23926_ /*58327*/;
assign _23930_ = _23263_ ^ _23926_ /*58330*/;
assign _23931_ = _23922_ & _23930_ /*58328*/;
assign _23711_ = _23922_ ^ _23930_ /*58329*/;
assign _23928_ = _23929_ | _23931_ /*58326*/;
assign _23933_ = ~Q[37] /*58325*/;
assign _23932_ = _23933_ & D[31] /*58324*/;
assign _23935_ = _23264_ & _23932_ /*58319*/;
assign _23936_ = _23264_ ^ _23932_ /*58322*/;
assign _23937_ = _23928_ & _23936_ /*58320*/;
assign _23712_ = _23928_ ^ _23936_ /*58321*/;
assign _23934_ = _23935_ | _23937_ /*58318*/;
assign _23939_ = ~Q[37] /*58317*/;
assign _23938_ = _23939_ & D[32] /*58316*/;
assign _23941_ = _23265_ & _23938_ /*58311*/;
assign _23942_ = _23265_ ^ _23938_ /*58314*/;
assign _23943_ = _23934_ & _23942_ /*58312*/;
assign _23713_ = _23934_ ^ _23942_ /*58313*/;
assign _23940_ = _23941_ | _23943_ /*58310*/;
assign _23945_ = ~Q[37] /*58309*/;
assign _23944_ = _23945_ & D[33] /*58308*/;
assign _23947_ = _23266_ & _23944_ /*58303*/;
assign _23948_ = _23266_ ^ _23944_ /*58306*/;
assign _23949_ = _23940_ & _23948_ /*58304*/;
assign _23714_ = _23940_ ^ _23948_ /*58305*/;
assign _23946_ = _23947_ | _23949_ /*58302*/;
assign _23951_ = ~Q[37] /*58301*/;
assign _23950_ = _23951_ & D[34] /*58300*/;
assign _23953_ = _23267_ & _23950_ /*58295*/;
assign _23954_ = _23267_ ^ _23950_ /*58298*/;
assign _23955_ = _23946_ & _23954_ /*58296*/;
assign _23715_ = _23946_ ^ _23954_ /*58297*/;
assign _23952_ = _23953_ | _23955_ /*58294*/;
assign _23957_ = ~Q[37] /*58293*/;
assign _23956_ = _23957_ & D[35] /*58292*/;
assign _23959_ = _23268_ & _23956_ /*58287*/;
assign _23960_ = _23268_ ^ _23956_ /*58290*/;
assign _23961_ = _23952_ & _23960_ /*58288*/;
assign _23716_ = _23952_ ^ _23960_ /*58289*/;
assign _23958_ = _23959_ | _23961_ /*58286*/;
assign _23963_ = ~Q[37] /*58285*/;
assign _23962_ = _23963_ & D[36] /*58284*/;
assign _23965_ = _23269_ & _23962_ /*58279*/;
assign _23966_ = _23269_ ^ _23962_ /*58282*/;
assign _23967_ = _23958_ & _23966_ /*58280*/;
assign _23717_ = _23958_ ^ _23966_ /*58281*/;
assign _23964_ = _23965_ | _23967_ /*58278*/;
assign _23969_ = ~Q[37] /*58277*/;
assign _23968_ = _23969_ & D[37] /*58276*/;
assign _23971_ = _23270_ & _23968_ /*58271*/;
assign _23972_ = _23270_ ^ _23968_ /*58274*/;
assign _23973_ = _23964_ & _23972_ /*58272*/;
assign _23718_ = _23964_ ^ _23972_ /*58273*/;
assign _23970_ = _23971_ | _23973_ /*58270*/;
assign _23975_ = ~Q[37] /*58269*/;
assign _23974_ = _23975_ & D[38] /*58268*/;
assign _23977_ = _23271_ & _23974_ /*58263*/;
assign _23978_ = _23271_ ^ _23974_ /*58266*/;
assign _23979_ = _23970_ & _23978_ /*58264*/;
assign _23719_ = _23970_ ^ _23978_ /*58265*/;
assign _23976_ = _23977_ | _23979_ /*58262*/;
assign _23981_ = ~Q[37] /*58261*/;
assign _23980_ = _23981_ & D[39] /*58260*/;
assign _23983_ = _23272_ & _23980_ /*58255*/;
assign _23984_ = _23272_ ^ _23980_ /*58258*/;
assign _23985_ = _23976_ & _23984_ /*58256*/;
assign _23720_ = _23976_ ^ _23984_ /*58257*/;
assign _23982_ = _23983_ | _23985_ /*58254*/;
assign _23987_ = ~Q[37] /*58253*/;
assign _23986_ = _23987_ & D[40] /*58252*/;
assign _23989_ = _23273_ & _23986_ /*58247*/;
assign _23990_ = _23273_ ^ _23986_ /*58250*/;
assign _23991_ = _23982_ & _23990_ /*58248*/;
assign _23721_ = _23982_ ^ _23990_ /*58249*/;
assign _23988_ = _23989_ | _23991_ /*58246*/;
assign _23993_ = ~Q[37] /*58245*/;
assign _23992_ = _23993_ & D[41] /*58244*/;
assign _23995_ = _23274_ & _23992_ /*58239*/;
assign _23996_ = _23274_ ^ _23992_ /*58242*/;
assign _23997_ = _23988_ & _23996_ /*58240*/;
assign _23722_ = _23988_ ^ _23996_ /*58241*/;
assign _23994_ = _23995_ | _23997_ /*58238*/;
assign _23999_ = ~Q[37] /*58237*/;
assign _23998_ = _23999_ & D[42] /*58236*/;
assign _24001_ = _23275_ & _23998_ /*58231*/;
assign _24002_ = _23275_ ^ _23998_ /*58234*/;
assign _24003_ = _23994_ & _24002_ /*58232*/;
assign _23723_ = _23994_ ^ _24002_ /*58233*/;
assign _24000_ = _24001_ | _24003_ /*58230*/;
assign _24005_ = ~Q[37] /*58229*/;
assign _24004_ = _24005_ & D[43] /*58228*/;
assign _24007_ = _23276_ & _24004_ /*58223*/;
assign _24008_ = _23276_ ^ _24004_ /*58226*/;
assign _24009_ = _24000_ & _24008_ /*58224*/;
assign _23724_ = _24000_ ^ _24008_ /*58225*/;
assign _24006_ = _24007_ | _24009_ /*58222*/;
assign _24011_ = ~Q[37] /*58221*/;
assign _24010_ = _24011_ & D[44] /*58220*/;
assign _24013_ = _23277_ & _24010_ /*58215*/;
assign _24014_ = _23277_ ^ _24010_ /*58218*/;
assign _24015_ = _24006_ & _24014_ /*58216*/;
assign _23725_ = _24006_ ^ _24014_ /*58217*/;
assign _24012_ = _24013_ | _24015_ /*58214*/;
assign _24017_ = ~Q[37] /*58213*/;
assign _24016_ = _24017_ & D[45] /*58212*/;
assign _24019_ = _23278_ & _24016_ /*58207*/;
assign _24020_ = _23278_ ^ _24016_ /*58210*/;
assign _24021_ = _24012_ & _24020_ /*58208*/;
assign _23726_ = _24012_ ^ _24020_ /*58209*/;
assign _24018_ = _24019_ | _24021_ /*58206*/;
assign _24023_ = ~Q[37] /*58205*/;
assign _24022_ = _24023_ & D[46] /*58204*/;
assign _24025_ = _23279_ & _24022_ /*58199*/;
assign _24026_ = _23279_ ^ _24022_ /*58202*/;
assign _24027_ = _24018_ & _24026_ /*58200*/;
assign _23727_ = _24018_ ^ _24026_ /*58201*/;
assign _24024_ = _24025_ | _24027_ /*58198*/;
assign _24029_ = ~Q[37] /*58197*/;
assign _24028_ = _24029_ & D[47] /*58196*/;
assign _24031_ = _23280_ & _24028_ /*58191*/;
assign _24032_ = _23280_ ^ _24028_ /*58194*/;
assign _24033_ = _24024_ & _24032_ /*58192*/;
assign _23728_ = _24024_ ^ _24032_ /*58193*/;
assign _24030_ = _24031_ | _24033_ /*58190*/;
assign _24035_ = ~Q[37] /*58189*/;
assign _24034_ = _24035_ & D[48] /*58188*/;
assign _24037_ = _23281_ & _24034_ /*58183*/;
assign _24038_ = _23281_ ^ _24034_ /*58186*/;
assign _24039_ = _24030_ & _24038_ /*58184*/;
assign _23729_ = _24030_ ^ _24038_ /*58185*/;
assign _24036_ = _24037_ | _24039_ /*58182*/;
assign _24041_ = ~Q[37] /*58181*/;
assign _24040_ = _24041_ & D[49] /*58180*/;
assign _24043_ = _23282_ & _24040_ /*58175*/;
assign _24044_ = _23282_ ^ _24040_ /*58178*/;
assign _24045_ = _24036_ & _24044_ /*58176*/;
assign _23730_ = _24036_ ^ _24044_ /*58177*/;
assign _24042_ = _24043_ | _24045_ /*58174*/;
assign _24047_ = ~Q[37] /*58173*/;
assign _24046_ = _24047_ & D[50] /*58172*/;
assign _24049_ = _23283_ & _24046_ /*58167*/;
assign _24050_ = _23283_ ^ _24046_ /*58170*/;
assign _24051_ = _24042_ & _24050_ /*58168*/;
assign _23731_ = _24042_ ^ _24050_ /*58169*/;
assign _24048_ = _24049_ | _24051_ /*58166*/;
assign _24053_ = ~Q[37] /*58165*/;
assign _24052_ = _24053_ & D[51] /*58164*/;
assign _24055_ = _23284_ & _24052_ /*58159*/;
assign _24056_ = _23284_ ^ _24052_ /*58162*/;
assign _24057_ = _24048_ & _24056_ /*58160*/;
assign _23732_ = _24048_ ^ _24056_ /*58161*/;
assign _24054_ = _24055_ | _24057_ /*58158*/;
assign _24059_ = ~Q[37] /*58157*/;
assign _24058_ = _24059_ & D[52] /*58156*/;
assign _24061_ = _23285_ & _24058_ /*58151*/;
assign _24062_ = _23285_ ^ _24058_ /*58154*/;
assign _24063_ = _24054_ & _24062_ /*58152*/;
assign _23733_ = _24054_ ^ _24062_ /*58153*/;
assign _24060_ = _24061_ | _24063_ /*58150*/;
assign _24065_ = ~Q[37] /*58149*/;
assign _24064_ = _24065_ & D[53] /*58148*/;
assign _24067_ = _23286_ & _24064_ /*58143*/;
assign _24068_ = _23286_ ^ _24064_ /*58146*/;
assign _24069_ = _24060_ & _24068_ /*58144*/;
assign _23734_ = _24060_ ^ _24068_ /*58145*/;
assign _24066_ = _24067_ | _24069_ /*58142*/;
assign _24071_ = ~Q[37] /*58141*/;
assign _24070_ = _24071_ & D[54] /*58140*/;
assign _24073_ = _23287_ & _24070_ /*58135*/;
assign _24074_ = _23287_ ^ _24070_ /*58138*/;
assign _24075_ = _24066_ & _24074_ /*58136*/;
assign _23735_ = _24066_ ^ _24074_ /*58137*/;
assign _24072_ = _24073_ | _24075_ /*58134*/;
assign _24077_ = ~Q[37] /*58133*/;
assign _24076_ = _24077_ & D[55] /*58132*/;
assign _24079_ = _23288_ & _24076_ /*58127*/;
assign _24080_ = _23288_ ^ _24076_ /*58130*/;
assign _24081_ = _24072_ & _24080_ /*58128*/;
assign _23736_ = _24072_ ^ _24080_ /*58129*/;
assign _24078_ = _24079_ | _24081_ /*58126*/;
assign _24083_ = ~Q[37] /*58125*/;
assign _24082_ = _24083_ & D[56] /*58124*/;
assign _24085_ = _23289_ & _24082_ /*58119*/;
assign _24086_ = _23289_ ^ _24082_ /*58122*/;
assign _24087_ = _24078_ & _24086_ /*58120*/;
assign _23737_ = _24078_ ^ _24086_ /*58121*/;
assign _24084_ = _24085_ | _24087_ /*58118*/;
assign _24089_ = ~Q[37] /*58117*/;
assign _24088_ = _24089_ & D[57] /*58116*/;
assign _24091_ = _23290_ & _24088_ /*58111*/;
assign _24092_ = _23290_ ^ _24088_ /*58114*/;
assign _24093_ = _24084_ & _24092_ /*58112*/;
assign _23738_ = _24084_ ^ _24092_ /*58113*/;
assign _24090_ = _24091_ | _24093_ /*58110*/;
assign _24095_ = ~Q[37] /*58109*/;
assign _24094_ = _24095_ & D[58] /*58108*/;
assign _24097_ = _23291_ & _24094_ /*58103*/;
assign _24098_ = _23291_ ^ _24094_ /*58106*/;
assign _24099_ = _24090_ & _24098_ /*58104*/;
assign _23739_ = _24090_ ^ _24098_ /*58105*/;
assign _24096_ = _24097_ | _24099_ /*58102*/;
assign _24101_ = ~Q[37] /*58101*/;
assign _24100_ = _24101_ & D[59] /*58100*/;
assign _24103_ = _23292_ & _24100_ /*58095*/;
assign _24104_ = _23292_ ^ _24100_ /*58098*/;
assign _24105_ = _24096_ & _24104_ /*58096*/;
assign _23740_ = _24096_ ^ _24104_ /*58097*/;
assign _24102_ = _24103_ | _24105_ /*58094*/;
assign _24107_ = ~Q[37] /*58093*/;
assign _24106_ = _24107_ & D[60] /*58092*/;
assign _24109_ = _23293_ & _24106_ /*58087*/;
assign _24110_ = _23293_ ^ _24106_ /*58090*/;
assign _24111_ = _24102_ & _24110_ /*58088*/;
assign _23741_ = _24102_ ^ _24110_ /*58089*/;
assign _24108_ = _24109_ | _24111_ /*58086*/;
assign _24113_ = ~Q[37] /*58085*/;
assign _24112_ = _24113_ & D[61] /*58084*/;
assign _24115_ = _23294_ & _24112_ /*58079*/;
assign _24116_ = _23294_ ^ _24112_ /*58082*/;
assign _24117_ = _24108_ & _24116_ /*58080*/;
assign _23742_ = _24108_ ^ _24116_ /*58081*/;
assign _24114_ = _24115_ | _24117_ /*58078*/;
assign _24119_ = ~Q[37] /*58077*/;
assign _24118_ = _24119_ & D[62] /*58076*/;
assign _24121_ = _23295_ & _24118_ /*58071*/;
assign _24122_ = _23295_ ^ _24118_ /*58074*/;
assign _24123_ = _24114_ & _24122_ /*58072*/;
assign _23743_ = _24114_ ^ _24122_ /*58073*/;
assign _24120_ = _24121_ | _24123_ /*58070*/;
assign _24125_ = ~Q[37] /*58069*/;
assign _24124_ = _24125_ & zeroWire /*58068*/;
assign _24126_ = _23296_ ^ _24124_ /*58066*/;
assign _23744_ = _24126_ ^ _24120_ /*58065*/;
assign _24197_ = ~D[0] /*57811*/;
assign _24194_ = R_0[36] & _24197_ /*57807*/;
assign _24195_ = R_0[36] ^ _24197_ /*57810*/;
assign _24196_ = oneWire & _24195_ /*57808*/;
assign _24129_ = oneWire ^ _24195_ /*57809*/;
assign _24193_ = _24194_ | _24196_ /*57806*/;
assign _24202_ = ~D[1] /*57805*/;
assign _24199_ = _23681_ & _24202_ /*57801*/;
assign _24200_ = _23681_ ^ _24202_ /*57804*/;
assign _24201_ = _24193_ & _24200_ /*57802*/;
assign _24130_ = _24193_ ^ _24200_ /*57803*/;
assign _24198_ = _24199_ | _24201_ /*57800*/;
assign _24207_ = ~D[2] /*57799*/;
assign _24204_ = _23682_ & _24207_ /*57795*/;
assign _24205_ = _23682_ ^ _24207_ /*57798*/;
assign _24206_ = _24198_ & _24205_ /*57796*/;
assign _24131_ = _24198_ ^ _24205_ /*57797*/;
assign _24203_ = _24204_ | _24206_ /*57794*/;
assign _24212_ = ~D[3] /*57793*/;
assign _24209_ = _23683_ & _24212_ /*57789*/;
assign _24210_ = _23683_ ^ _24212_ /*57792*/;
assign _24211_ = _24203_ & _24210_ /*57790*/;
assign _24132_ = _24203_ ^ _24210_ /*57791*/;
assign _24208_ = _24209_ | _24211_ /*57788*/;
assign _24217_ = ~D[4] /*57787*/;
assign _24214_ = _23684_ & _24217_ /*57783*/;
assign _24215_ = _23684_ ^ _24217_ /*57786*/;
assign _24216_ = _24208_ & _24215_ /*57784*/;
assign _24133_ = _24208_ ^ _24215_ /*57785*/;
assign _24213_ = _24214_ | _24216_ /*57782*/;
assign _24222_ = ~D[5] /*57781*/;
assign _24219_ = _23685_ & _24222_ /*57777*/;
assign _24220_ = _23685_ ^ _24222_ /*57780*/;
assign _24221_ = _24213_ & _24220_ /*57778*/;
assign _24134_ = _24213_ ^ _24220_ /*57779*/;
assign _24218_ = _24219_ | _24221_ /*57776*/;
assign _24227_ = ~D[6] /*57775*/;
assign _24224_ = _23686_ & _24227_ /*57771*/;
assign _24225_ = _23686_ ^ _24227_ /*57774*/;
assign _24226_ = _24218_ & _24225_ /*57772*/;
assign _24135_ = _24218_ ^ _24225_ /*57773*/;
assign _24223_ = _24224_ | _24226_ /*57770*/;
assign _24232_ = ~D[7] /*57769*/;
assign _24229_ = _23687_ & _24232_ /*57765*/;
assign _24230_ = _23687_ ^ _24232_ /*57768*/;
assign _24231_ = _24223_ & _24230_ /*57766*/;
assign _24136_ = _24223_ ^ _24230_ /*57767*/;
assign _24228_ = _24229_ | _24231_ /*57764*/;
assign _24237_ = ~D[8] /*57763*/;
assign _24234_ = _23688_ & _24237_ /*57759*/;
assign _24235_ = _23688_ ^ _24237_ /*57762*/;
assign _24236_ = _24228_ & _24235_ /*57760*/;
assign _24137_ = _24228_ ^ _24235_ /*57761*/;
assign _24233_ = _24234_ | _24236_ /*57758*/;
assign _24242_ = ~D[9] /*57757*/;
assign _24239_ = _23689_ & _24242_ /*57753*/;
assign _24240_ = _23689_ ^ _24242_ /*57756*/;
assign _24241_ = _24233_ & _24240_ /*57754*/;
assign _24138_ = _24233_ ^ _24240_ /*57755*/;
assign _24238_ = _24239_ | _24241_ /*57752*/;
assign _24247_ = ~D[10] /*57751*/;
assign _24244_ = _23690_ & _24247_ /*57747*/;
assign _24245_ = _23690_ ^ _24247_ /*57750*/;
assign _24246_ = _24238_ & _24245_ /*57748*/;
assign _24139_ = _24238_ ^ _24245_ /*57749*/;
assign _24243_ = _24244_ | _24246_ /*57746*/;
assign _24252_ = ~D[11] /*57745*/;
assign _24249_ = _23691_ & _24252_ /*57741*/;
assign _24250_ = _23691_ ^ _24252_ /*57744*/;
assign _24251_ = _24243_ & _24250_ /*57742*/;
assign _24140_ = _24243_ ^ _24250_ /*57743*/;
assign _24248_ = _24249_ | _24251_ /*57740*/;
assign _24257_ = ~D[12] /*57739*/;
assign _24254_ = _23692_ & _24257_ /*57735*/;
assign _24255_ = _23692_ ^ _24257_ /*57738*/;
assign _24256_ = _24248_ & _24255_ /*57736*/;
assign _24141_ = _24248_ ^ _24255_ /*57737*/;
assign _24253_ = _24254_ | _24256_ /*57734*/;
assign _24262_ = ~D[13] /*57733*/;
assign _24259_ = _23693_ & _24262_ /*57729*/;
assign _24260_ = _23693_ ^ _24262_ /*57732*/;
assign _24261_ = _24253_ & _24260_ /*57730*/;
assign _24142_ = _24253_ ^ _24260_ /*57731*/;
assign _24258_ = _24259_ | _24261_ /*57728*/;
assign _24267_ = ~D[14] /*57727*/;
assign _24264_ = _23694_ & _24267_ /*57723*/;
assign _24265_ = _23694_ ^ _24267_ /*57726*/;
assign _24266_ = _24258_ & _24265_ /*57724*/;
assign _24143_ = _24258_ ^ _24265_ /*57725*/;
assign _24263_ = _24264_ | _24266_ /*57722*/;
assign _24272_ = ~D[15] /*57721*/;
assign _24269_ = _23695_ & _24272_ /*57717*/;
assign _24270_ = _23695_ ^ _24272_ /*57720*/;
assign _24271_ = _24263_ & _24270_ /*57718*/;
assign _24144_ = _24263_ ^ _24270_ /*57719*/;
assign _24268_ = _24269_ | _24271_ /*57716*/;
assign _24277_ = ~D[16] /*57715*/;
assign _24274_ = _23696_ & _24277_ /*57711*/;
assign _24275_ = _23696_ ^ _24277_ /*57714*/;
assign _24276_ = _24268_ & _24275_ /*57712*/;
assign _24145_ = _24268_ ^ _24275_ /*57713*/;
assign _24273_ = _24274_ | _24276_ /*57710*/;
assign _24282_ = ~D[17] /*57709*/;
assign _24279_ = _23697_ & _24282_ /*57705*/;
assign _24280_ = _23697_ ^ _24282_ /*57708*/;
assign _24281_ = _24273_ & _24280_ /*57706*/;
assign _24146_ = _24273_ ^ _24280_ /*57707*/;
assign _24278_ = _24279_ | _24281_ /*57704*/;
assign _24287_ = ~D[18] /*57703*/;
assign _24284_ = _23698_ & _24287_ /*57699*/;
assign _24285_ = _23698_ ^ _24287_ /*57702*/;
assign _24286_ = _24278_ & _24285_ /*57700*/;
assign _24147_ = _24278_ ^ _24285_ /*57701*/;
assign _24283_ = _24284_ | _24286_ /*57698*/;
assign _24292_ = ~D[19] /*57697*/;
assign _24289_ = _23699_ & _24292_ /*57693*/;
assign _24290_ = _23699_ ^ _24292_ /*57696*/;
assign _24291_ = _24283_ & _24290_ /*57694*/;
assign _24148_ = _24283_ ^ _24290_ /*57695*/;
assign _24288_ = _24289_ | _24291_ /*57692*/;
assign _24297_ = ~D[20] /*57691*/;
assign _24294_ = _23700_ & _24297_ /*57687*/;
assign _24295_ = _23700_ ^ _24297_ /*57690*/;
assign _24296_ = _24288_ & _24295_ /*57688*/;
assign _24149_ = _24288_ ^ _24295_ /*57689*/;
assign _24293_ = _24294_ | _24296_ /*57686*/;
assign _24302_ = ~D[21] /*57685*/;
assign _24299_ = _23701_ & _24302_ /*57681*/;
assign _24300_ = _23701_ ^ _24302_ /*57684*/;
assign _24301_ = _24293_ & _24300_ /*57682*/;
assign _24150_ = _24293_ ^ _24300_ /*57683*/;
assign _24298_ = _24299_ | _24301_ /*57680*/;
assign _24307_ = ~D[22] /*57679*/;
assign _24304_ = _23702_ & _24307_ /*57675*/;
assign _24305_ = _23702_ ^ _24307_ /*57678*/;
assign _24306_ = _24298_ & _24305_ /*57676*/;
assign _24151_ = _24298_ ^ _24305_ /*57677*/;
assign _24303_ = _24304_ | _24306_ /*57674*/;
assign _24312_ = ~D[23] /*57673*/;
assign _24309_ = _23703_ & _24312_ /*57669*/;
assign _24310_ = _23703_ ^ _24312_ /*57672*/;
assign _24311_ = _24303_ & _24310_ /*57670*/;
assign _24152_ = _24303_ ^ _24310_ /*57671*/;
assign _24308_ = _24309_ | _24311_ /*57668*/;
assign _24317_ = ~D[24] /*57667*/;
assign _24314_ = _23704_ & _24317_ /*57663*/;
assign _24315_ = _23704_ ^ _24317_ /*57666*/;
assign _24316_ = _24308_ & _24315_ /*57664*/;
assign _24153_ = _24308_ ^ _24315_ /*57665*/;
assign _24313_ = _24314_ | _24316_ /*57662*/;
assign _24322_ = ~D[25] /*57661*/;
assign _24319_ = _23705_ & _24322_ /*57657*/;
assign _24320_ = _23705_ ^ _24322_ /*57660*/;
assign _24321_ = _24313_ & _24320_ /*57658*/;
assign _24154_ = _24313_ ^ _24320_ /*57659*/;
assign _24318_ = _24319_ | _24321_ /*57656*/;
assign _24327_ = ~D[26] /*57655*/;
assign _24324_ = _23706_ & _24327_ /*57651*/;
assign _24325_ = _23706_ ^ _24327_ /*57654*/;
assign _24326_ = _24318_ & _24325_ /*57652*/;
assign _24155_ = _24318_ ^ _24325_ /*57653*/;
assign _24323_ = _24324_ | _24326_ /*57650*/;
assign _24332_ = ~D[27] /*57649*/;
assign _24329_ = _23707_ & _24332_ /*57645*/;
assign _24330_ = _23707_ ^ _24332_ /*57648*/;
assign _24331_ = _24323_ & _24330_ /*57646*/;
assign _24156_ = _24323_ ^ _24330_ /*57647*/;
assign _24328_ = _24329_ | _24331_ /*57644*/;
assign _24337_ = ~D[28] /*57643*/;
assign _24334_ = _23708_ & _24337_ /*57639*/;
assign _24335_ = _23708_ ^ _24337_ /*57642*/;
assign _24336_ = _24328_ & _24335_ /*57640*/;
assign _24157_ = _24328_ ^ _24335_ /*57641*/;
assign _24333_ = _24334_ | _24336_ /*57638*/;
assign _24342_ = ~D[29] /*57637*/;
assign _24339_ = _23709_ & _24342_ /*57633*/;
assign _24340_ = _23709_ ^ _24342_ /*57636*/;
assign _24341_ = _24333_ & _24340_ /*57634*/;
assign _24158_ = _24333_ ^ _24340_ /*57635*/;
assign _24338_ = _24339_ | _24341_ /*57632*/;
assign _24347_ = ~D[30] /*57631*/;
assign _24344_ = _23710_ & _24347_ /*57627*/;
assign _24345_ = _23710_ ^ _24347_ /*57630*/;
assign _24346_ = _24338_ & _24345_ /*57628*/;
assign _24159_ = _24338_ ^ _24345_ /*57629*/;
assign _24343_ = _24344_ | _24346_ /*57626*/;
assign _24352_ = ~D[31] /*57625*/;
assign _24349_ = _23711_ & _24352_ /*57621*/;
assign _24350_ = _23711_ ^ _24352_ /*57624*/;
assign _24351_ = _24343_ & _24350_ /*57622*/;
assign _24160_ = _24343_ ^ _24350_ /*57623*/;
assign _24348_ = _24349_ | _24351_ /*57620*/;
assign _24357_ = ~D[32] /*57619*/;
assign _24354_ = _23712_ & _24357_ /*57615*/;
assign _24355_ = _23712_ ^ _24357_ /*57618*/;
assign _24356_ = _24348_ & _24355_ /*57616*/;
assign _24161_ = _24348_ ^ _24355_ /*57617*/;
assign _24353_ = _24354_ | _24356_ /*57614*/;
assign _24362_ = ~D[33] /*57613*/;
assign _24359_ = _23713_ & _24362_ /*57609*/;
assign _24360_ = _23713_ ^ _24362_ /*57612*/;
assign _24361_ = _24353_ & _24360_ /*57610*/;
assign _24162_ = _24353_ ^ _24360_ /*57611*/;
assign _24358_ = _24359_ | _24361_ /*57608*/;
assign _24367_ = ~D[34] /*57607*/;
assign _24364_ = _23714_ & _24367_ /*57603*/;
assign _24365_ = _23714_ ^ _24367_ /*57606*/;
assign _24366_ = _24358_ & _24365_ /*57604*/;
assign _24163_ = _24358_ ^ _24365_ /*57605*/;
assign _24363_ = _24364_ | _24366_ /*57602*/;
assign _24372_ = ~D[35] /*57601*/;
assign _24369_ = _23715_ & _24372_ /*57597*/;
assign _24370_ = _23715_ ^ _24372_ /*57600*/;
assign _24371_ = _24363_ & _24370_ /*57598*/;
assign _24164_ = _24363_ ^ _24370_ /*57599*/;
assign _24368_ = _24369_ | _24371_ /*57596*/;
assign _24377_ = ~D[36] /*57595*/;
assign _24374_ = _23716_ & _24377_ /*57591*/;
assign _24375_ = _23716_ ^ _24377_ /*57594*/;
assign _24376_ = _24368_ & _24375_ /*57592*/;
assign _24165_ = _24368_ ^ _24375_ /*57593*/;
assign _24373_ = _24374_ | _24376_ /*57590*/;
assign _24382_ = ~D[37] /*57589*/;
assign _24379_ = _23717_ & _24382_ /*57585*/;
assign _24380_ = _23717_ ^ _24382_ /*57588*/;
assign _24381_ = _24373_ & _24380_ /*57586*/;
assign _24166_ = _24373_ ^ _24380_ /*57587*/;
assign _24378_ = _24379_ | _24381_ /*57584*/;
assign _24387_ = ~D[38] /*57583*/;
assign _24384_ = _23718_ & _24387_ /*57579*/;
assign _24385_ = _23718_ ^ _24387_ /*57582*/;
assign _24386_ = _24378_ & _24385_ /*57580*/;
assign _24167_ = _24378_ ^ _24385_ /*57581*/;
assign _24383_ = _24384_ | _24386_ /*57578*/;
assign _24392_ = ~D[39] /*57577*/;
assign _24389_ = _23719_ & _24392_ /*57573*/;
assign _24390_ = _23719_ ^ _24392_ /*57576*/;
assign _24391_ = _24383_ & _24390_ /*57574*/;
assign _24168_ = _24383_ ^ _24390_ /*57575*/;
assign _24388_ = _24389_ | _24391_ /*57572*/;
assign _24397_ = ~D[40] /*57571*/;
assign _24394_ = _23720_ & _24397_ /*57567*/;
assign _24395_ = _23720_ ^ _24397_ /*57570*/;
assign _24396_ = _24388_ & _24395_ /*57568*/;
assign _24169_ = _24388_ ^ _24395_ /*57569*/;
assign _24393_ = _24394_ | _24396_ /*57566*/;
assign _24402_ = ~D[41] /*57565*/;
assign _24399_ = _23721_ & _24402_ /*57561*/;
assign _24400_ = _23721_ ^ _24402_ /*57564*/;
assign _24401_ = _24393_ & _24400_ /*57562*/;
assign _24170_ = _24393_ ^ _24400_ /*57563*/;
assign _24398_ = _24399_ | _24401_ /*57560*/;
assign _24407_ = ~D[42] /*57559*/;
assign _24404_ = _23722_ & _24407_ /*57555*/;
assign _24405_ = _23722_ ^ _24407_ /*57558*/;
assign _24406_ = _24398_ & _24405_ /*57556*/;
assign _24171_ = _24398_ ^ _24405_ /*57557*/;
assign _24403_ = _24404_ | _24406_ /*57554*/;
assign _24412_ = ~D[43] /*57553*/;
assign _24409_ = _23723_ & _24412_ /*57549*/;
assign _24410_ = _23723_ ^ _24412_ /*57552*/;
assign _24411_ = _24403_ & _24410_ /*57550*/;
assign _24172_ = _24403_ ^ _24410_ /*57551*/;
assign _24408_ = _24409_ | _24411_ /*57548*/;
assign _24417_ = ~D[44] /*57547*/;
assign _24414_ = _23724_ & _24417_ /*57543*/;
assign _24415_ = _23724_ ^ _24417_ /*57546*/;
assign _24416_ = _24408_ & _24415_ /*57544*/;
assign _24173_ = _24408_ ^ _24415_ /*57545*/;
assign _24413_ = _24414_ | _24416_ /*57542*/;
assign _24422_ = ~D[45] /*57541*/;
assign _24419_ = _23725_ & _24422_ /*57537*/;
assign _24420_ = _23725_ ^ _24422_ /*57540*/;
assign _24421_ = _24413_ & _24420_ /*57538*/;
assign _24174_ = _24413_ ^ _24420_ /*57539*/;
assign _24418_ = _24419_ | _24421_ /*57536*/;
assign _24427_ = ~D[46] /*57535*/;
assign _24424_ = _23726_ & _24427_ /*57531*/;
assign _24425_ = _23726_ ^ _24427_ /*57534*/;
assign _24426_ = _24418_ & _24425_ /*57532*/;
assign _24175_ = _24418_ ^ _24425_ /*57533*/;
assign _24423_ = _24424_ | _24426_ /*57530*/;
assign _24432_ = ~D[47] /*57529*/;
assign _24429_ = _23727_ & _24432_ /*57525*/;
assign _24430_ = _23727_ ^ _24432_ /*57528*/;
assign _24431_ = _24423_ & _24430_ /*57526*/;
assign _24176_ = _24423_ ^ _24430_ /*57527*/;
assign _24428_ = _24429_ | _24431_ /*57524*/;
assign _24437_ = ~D[48] /*57523*/;
assign _24434_ = _23728_ & _24437_ /*57519*/;
assign _24435_ = _23728_ ^ _24437_ /*57522*/;
assign _24436_ = _24428_ & _24435_ /*57520*/;
assign _24177_ = _24428_ ^ _24435_ /*57521*/;
assign _24433_ = _24434_ | _24436_ /*57518*/;
assign _24442_ = ~D[49] /*57517*/;
assign _24439_ = _23729_ & _24442_ /*57513*/;
assign _24440_ = _23729_ ^ _24442_ /*57516*/;
assign _24441_ = _24433_ & _24440_ /*57514*/;
assign _24178_ = _24433_ ^ _24440_ /*57515*/;
assign _24438_ = _24439_ | _24441_ /*57512*/;
assign _24447_ = ~D[50] /*57511*/;
assign _24444_ = _23730_ & _24447_ /*57507*/;
assign _24445_ = _23730_ ^ _24447_ /*57510*/;
assign _24446_ = _24438_ & _24445_ /*57508*/;
assign _24179_ = _24438_ ^ _24445_ /*57509*/;
assign _24443_ = _24444_ | _24446_ /*57506*/;
assign _24452_ = ~D[51] /*57505*/;
assign _24449_ = _23731_ & _24452_ /*57501*/;
assign _24450_ = _23731_ ^ _24452_ /*57504*/;
assign _24451_ = _24443_ & _24450_ /*57502*/;
assign _24180_ = _24443_ ^ _24450_ /*57503*/;
assign _24448_ = _24449_ | _24451_ /*57500*/;
assign _24457_ = ~D[52] /*57499*/;
assign _24454_ = _23732_ & _24457_ /*57495*/;
assign _24455_ = _23732_ ^ _24457_ /*57498*/;
assign _24456_ = _24448_ & _24455_ /*57496*/;
assign _24181_ = _24448_ ^ _24455_ /*57497*/;
assign _24453_ = _24454_ | _24456_ /*57494*/;
assign _24462_ = ~D[53] /*57493*/;
assign _24459_ = _23733_ & _24462_ /*57489*/;
assign _24460_ = _23733_ ^ _24462_ /*57492*/;
assign _24461_ = _24453_ & _24460_ /*57490*/;
assign _24182_ = _24453_ ^ _24460_ /*57491*/;
assign _24458_ = _24459_ | _24461_ /*57488*/;
assign _24467_ = ~D[54] /*57487*/;
assign _24464_ = _23734_ & _24467_ /*57483*/;
assign _24465_ = _23734_ ^ _24467_ /*57486*/;
assign _24466_ = _24458_ & _24465_ /*57484*/;
assign _24183_ = _24458_ ^ _24465_ /*57485*/;
assign _24463_ = _24464_ | _24466_ /*57482*/;
assign _24472_ = ~D[55] /*57481*/;
assign _24469_ = _23735_ & _24472_ /*57477*/;
assign _24470_ = _23735_ ^ _24472_ /*57480*/;
assign _24471_ = _24463_ & _24470_ /*57478*/;
assign _24184_ = _24463_ ^ _24470_ /*57479*/;
assign _24468_ = _24469_ | _24471_ /*57476*/;
assign _24477_ = ~D[56] /*57475*/;
assign _24474_ = _23736_ & _24477_ /*57471*/;
assign _24475_ = _23736_ ^ _24477_ /*57474*/;
assign _24476_ = _24468_ & _24475_ /*57472*/;
assign _24185_ = _24468_ ^ _24475_ /*57473*/;
assign _24473_ = _24474_ | _24476_ /*57470*/;
assign _24482_ = ~D[57] /*57469*/;
assign _24479_ = _23737_ & _24482_ /*57465*/;
assign _24480_ = _23737_ ^ _24482_ /*57468*/;
assign _24481_ = _24473_ & _24480_ /*57466*/;
assign _24186_ = _24473_ ^ _24480_ /*57467*/;
assign _24478_ = _24479_ | _24481_ /*57464*/;
assign _24487_ = ~D[58] /*57463*/;
assign _24484_ = _23738_ & _24487_ /*57459*/;
assign _24485_ = _23738_ ^ _24487_ /*57462*/;
assign _24486_ = _24478_ & _24485_ /*57460*/;
assign _24187_ = _24478_ ^ _24485_ /*57461*/;
assign _24483_ = _24484_ | _24486_ /*57458*/;
assign _24492_ = ~D[59] /*57457*/;
assign _24489_ = _23739_ & _24492_ /*57453*/;
assign _24490_ = _23739_ ^ _24492_ /*57456*/;
assign _24491_ = _24483_ & _24490_ /*57454*/;
assign _24188_ = _24483_ ^ _24490_ /*57455*/;
assign _24488_ = _24489_ | _24491_ /*57452*/;
assign _24497_ = ~D[60] /*57451*/;
assign _24494_ = _23740_ & _24497_ /*57447*/;
assign _24495_ = _23740_ ^ _24497_ /*57450*/;
assign _24496_ = _24488_ & _24495_ /*57448*/;
assign _24189_ = _24488_ ^ _24495_ /*57449*/;
assign _24493_ = _24494_ | _24496_ /*57446*/;
assign _24502_ = ~D[61] /*57445*/;
assign _24499_ = _23741_ & _24502_ /*57441*/;
assign _24500_ = _23741_ ^ _24502_ /*57444*/;
assign _24501_ = _24493_ & _24500_ /*57442*/;
assign _24190_ = _24493_ ^ _24500_ /*57443*/;
assign _24498_ = _24499_ | _24501_ /*57440*/;
assign _24507_ = ~D[62] /*57439*/;
assign _24504_ = _23742_ & _24507_ /*57435*/;
assign _24505_ = _23742_ ^ _24507_ /*57438*/;
assign _24506_ = _24498_ & _24505_ /*57436*/;
assign _24191_ = _24498_ ^ _24505_ /*57437*/;
assign _24503_ = _24504_ | _24506_ /*57434*/;
assign _24508_ = _23743_ & oneWire /*57429*/;
assign _24509_ = _23743_ ^ oneWire /*57432*/;
assign _24510_ = _24503_ & _24509_ /*57430*/;
assign _24192_ = _24503_ ^ _24509_ /*57431*/;
assign Q[36] = _24508_ | _24510_ /*57428*/;
assign _24643_ = ~Q[36] /*57043*/;
assign _24642_ = _24643_ & D[0] /*57042*/;
assign _24645_ = _24129_ & _24642_ /*57037*/;
assign _24646_ = _24129_ ^ _24642_ /*57040*/;
assign _24647_ = zeroWire & _24646_ /*57038*/;
assign _24577_ = zeroWire ^ _24646_ /*57039*/;
assign _24644_ = _24645_ | _24647_ /*57036*/;
assign _24649_ = ~Q[36] /*57035*/;
assign _24648_ = _24649_ & D[1] /*57034*/;
assign _24651_ = _24130_ & _24648_ /*57029*/;
assign _24652_ = _24130_ ^ _24648_ /*57032*/;
assign _24653_ = _24644_ & _24652_ /*57030*/;
assign _24578_ = _24644_ ^ _24652_ /*57031*/;
assign _24650_ = _24651_ | _24653_ /*57028*/;
assign _24655_ = ~Q[36] /*57027*/;
assign _24654_ = _24655_ & D[2] /*57026*/;
assign _24657_ = _24131_ & _24654_ /*57021*/;
assign _24658_ = _24131_ ^ _24654_ /*57024*/;
assign _24659_ = _24650_ & _24658_ /*57022*/;
assign _24579_ = _24650_ ^ _24658_ /*57023*/;
assign _24656_ = _24657_ | _24659_ /*57020*/;
assign _24661_ = ~Q[36] /*57019*/;
assign _24660_ = _24661_ & D[3] /*57018*/;
assign _24663_ = _24132_ & _24660_ /*57013*/;
assign _24664_ = _24132_ ^ _24660_ /*57016*/;
assign _24665_ = _24656_ & _24664_ /*57014*/;
assign _24580_ = _24656_ ^ _24664_ /*57015*/;
assign _24662_ = _24663_ | _24665_ /*57012*/;
assign _24667_ = ~Q[36] /*57011*/;
assign _24666_ = _24667_ & D[4] /*57010*/;
assign _24669_ = _24133_ & _24666_ /*57005*/;
assign _24670_ = _24133_ ^ _24666_ /*57008*/;
assign _24671_ = _24662_ & _24670_ /*57006*/;
assign _24581_ = _24662_ ^ _24670_ /*57007*/;
assign _24668_ = _24669_ | _24671_ /*57004*/;
assign _24673_ = ~Q[36] /*57003*/;
assign _24672_ = _24673_ & D[5] /*57002*/;
assign _24675_ = _24134_ & _24672_ /*56997*/;
assign _24676_ = _24134_ ^ _24672_ /*57000*/;
assign _24677_ = _24668_ & _24676_ /*56998*/;
assign _24582_ = _24668_ ^ _24676_ /*56999*/;
assign _24674_ = _24675_ | _24677_ /*56996*/;
assign _24679_ = ~Q[36] /*56995*/;
assign _24678_ = _24679_ & D[6] /*56994*/;
assign _24681_ = _24135_ & _24678_ /*56989*/;
assign _24682_ = _24135_ ^ _24678_ /*56992*/;
assign _24683_ = _24674_ & _24682_ /*56990*/;
assign _24583_ = _24674_ ^ _24682_ /*56991*/;
assign _24680_ = _24681_ | _24683_ /*56988*/;
assign _24685_ = ~Q[36] /*56987*/;
assign _24684_ = _24685_ & D[7] /*56986*/;
assign _24687_ = _24136_ & _24684_ /*56981*/;
assign _24688_ = _24136_ ^ _24684_ /*56984*/;
assign _24689_ = _24680_ & _24688_ /*56982*/;
assign _24584_ = _24680_ ^ _24688_ /*56983*/;
assign _24686_ = _24687_ | _24689_ /*56980*/;
assign _24691_ = ~Q[36] /*56979*/;
assign _24690_ = _24691_ & D[8] /*56978*/;
assign _24693_ = _24137_ & _24690_ /*56973*/;
assign _24694_ = _24137_ ^ _24690_ /*56976*/;
assign _24695_ = _24686_ & _24694_ /*56974*/;
assign _24585_ = _24686_ ^ _24694_ /*56975*/;
assign _24692_ = _24693_ | _24695_ /*56972*/;
assign _24697_ = ~Q[36] /*56971*/;
assign _24696_ = _24697_ & D[9] /*56970*/;
assign _24699_ = _24138_ & _24696_ /*56965*/;
assign _24700_ = _24138_ ^ _24696_ /*56968*/;
assign _24701_ = _24692_ & _24700_ /*56966*/;
assign _24586_ = _24692_ ^ _24700_ /*56967*/;
assign _24698_ = _24699_ | _24701_ /*56964*/;
assign _24703_ = ~Q[36] /*56963*/;
assign _24702_ = _24703_ & D[10] /*56962*/;
assign _24705_ = _24139_ & _24702_ /*56957*/;
assign _24706_ = _24139_ ^ _24702_ /*56960*/;
assign _24707_ = _24698_ & _24706_ /*56958*/;
assign _24587_ = _24698_ ^ _24706_ /*56959*/;
assign _24704_ = _24705_ | _24707_ /*56956*/;
assign _24709_ = ~Q[36] /*56955*/;
assign _24708_ = _24709_ & D[11] /*56954*/;
assign _24711_ = _24140_ & _24708_ /*56949*/;
assign _24712_ = _24140_ ^ _24708_ /*56952*/;
assign _24713_ = _24704_ & _24712_ /*56950*/;
assign _24588_ = _24704_ ^ _24712_ /*56951*/;
assign _24710_ = _24711_ | _24713_ /*56948*/;
assign _24715_ = ~Q[36] /*56947*/;
assign _24714_ = _24715_ & D[12] /*56946*/;
assign _24717_ = _24141_ & _24714_ /*56941*/;
assign _24718_ = _24141_ ^ _24714_ /*56944*/;
assign _24719_ = _24710_ & _24718_ /*56942*/;
assign _24589_ = _24710_ ^ _24718_ /*56943*/;
assign _24716_ = _24717_ | _24719_ /*56940*/;
assign _24721_ = ~Q[36] /*56939*/;
assign _24720_ = _24721_ & D[13] /*56938*/;
assign _24723_ = _24142_ & _24720_ /*56933*/;
assign _24724_ = _24142_ ^ _24720_ /*56936*/;
assign _24725_ = _24716_ & _24724_ /*56934*/;
assign _24590_ = _24716_ ^ _24724_ /*56935*/;
assign _24722_ = _24723_ | _24725_ /*56932*/;
assign _24727_ = ~Q[36] /*56931*/;
assign _24726_ = _24727_ & D[14] /*56930*/;
assign _24729_ = _24143_ & _24726_ /*56925*/;
assign _24730_ = _24143_ ^ _24726_ /*56928*/;
assign _24731_ = _24722_ & _24730_ /*56926*/;
assign _24591_ = _24722_ ^ _24730_ /*56927*/;
assign _24728_ = _24729_ | _24731_ /*56924*/;
assign _24733_ = ~Q[36] /*56923*/;
assign _24732_ = _24733_ & D[15] /*56922*/;
assign _24735_ = _24144_ & _24732_ /*56917*/;
assign _24736_ = _24144_ ^ _24732_ /*56920*/;
assign _24737_ = _24728_ & _24736_ /*56918*/;
assign _24592_ = _24728_ ^ _24736_ /*56919*/;
assign _24734_ = _24735_ | _24737_ /*56916*/;
assign _24739_ = ~Q[36] /*56915*/;
assign _24738_ = _24739_ & D[16] /*56914*/;
assign _24741_ = _24145_ & _24738_ /*56909*/;
assign _24742_ = _24145_ ^ _24738_ /*56912*/;
assign _24743_ = _24734_ & _24742_ /*56910*/;
assign _24593_ = _24734_ ^ _24742_ /*56911*/;
assign _24740_ = _24741_ | _24743_ /*56908*/;
assign _24745_ = ~Q[36] /*56907*/;
assign _24744_ = _24745_ & D[17] /*56906*/;
assign _24747_ = _24146_ & _24744_ /*56901*/;
assign _24748_ = _24146_ ^ _24744_ /*56904*/;
assign _24749_ = _24740_ & _24748_ /*56902*/;
assign _24594_ = _24740_ ^ _24748_ /*56903*/;
assign _24746_ = _24747_ | _24749_ /*56900*/;
assign _24751_ = ~Q[36] /*56899*/;
assign _24750_ = _24751_ & D[18] /*56898*/;
assign _24753_ = _24147_ & _24750_ /*56893*/;
assign _24754_ = _24147_ ^ _24750_ /*56896*/;
assign _24755_ = _24746_ & _24754_ /*56894*/;
assign _24595_ = _24746_ ^ _24754_ /*56895*/;
assign _24752_ = _24753_ | _24755_ /*56892*/;
assign _24757_ = ~Q[36] /*56891*/;
assign _24756_ = _24757_ & D[19] /*56890*/;
assign _24759_ = _24148_ & _24756_ /*56885*/;
assign _24760_ = _24148_ ^ _24756_ /*56888*/;
assign _24761_ = _24752_ & _24760_ /*56886*/;
assign _24596_ = _24752_ ^ _24760_ /*56887*/;
assign _24758_ = _24759_ | _24761_ /*56884*/;
assign _24763_ = ~Q[36] /*56883*/;
assign _24762_ = _24763_ & D[20] /*56882*/;
assign _24765_ = _24149_ & _24762_ /*56877*/;
assign _24766_ = _24149_ ^ _24762_ /*56880*/;
assign _24767_ = _24758_ & _24766_ /*56878*/;
assign _24597_ = _24758_ ^ _24766_ /*56879*/;
assign _24764_ = _24765_ | _24767_ /*56876*/;
assign _24769_ = ~Q[36] /*56875*/;
assign _24768_ = _24769_ & D[21] /*56874*/;
assign _24771_ = _24150_ & _24768_ /*56869*/;
assign _24772_ = _24150_ ^ _24768_ /*56872*/;
assign _24773_ = _24764_ & _24772_ /*56870*/;
assign _24598_ = _24764_ ^ _24772_ /*56871*/;
assign _24770_ = _24771_ | _24773_ /*56868*/;
assign _24775_ = ~Q[36] /*56867*/;
assign _24774_ = _24775_ & D[22] /*56866*/;
assign _24777_ = _24151_ & _24774_ /*56861*/;
assign _24778_ = _24151_ ^ _24774_ /*56864*/;
assign _24779_ = _24770_ & _24778_ /*56862*/;
assign _24599_ = _24770_ ^ _24778_ /*56863*/;
assign _24776_ = _24777_ | _24779_ /*56860*/;
assign _24781_ = ~Q[36] /*56859*/;
assign _24780_ = _24781_ & D[23] /*56858*/;
assign _24783_ = _24152_ & _24780_ /*56853*/;
assign _24784_ = _24152_ ^ _24780_ /*56856*/;
assign _24785_ = _24776_ & _24784_ /*56854*/;
assign _24600_ = _24776_ ^ _24784_ /*56855*/;
assign _24782_ = _24783_ | _24785_ /*56852*/;
assign _24787_ = ~Q[36] /*56851*/;
assign _24786_ = _24787_ & D[24] /*56850*/;
assign _24789_ = _24153_ & _24786_ /*56845*/;
assign _24790_ = _24153_ ^ _24786_ /*56848*/;
assign _24791_ = _24782_ & _24790_ /*56846*/;
assign _24601_ = _24782_ ^ _24790_ /*56847*/;
assign _24788_ = _24789_ | _24791_ /*56844*/;
assign _24793_ = ~Q[36] /*56843*/;
assign _24792_ = _24793_ & D[25] /*56842*/;
assign _24795_ = _24154_ & _24792_ /*56837*/;
assign _24796_ = _24154_ ^ _24792_ /*56840*/;
assign _24797_ = _24788_ & _24796_ /*56838*/;
assign _24602_ = _24788_ ^ _24796_ /*56839*/;
assign _24794_ = _24795_ | _24797_ /*56836*/;
assign _24799_ = ~Q[36] /*56835*/;
assign _24798_ = _24799_ & D[26] /*56834*/;
assign _24801_ = _24155_ & _24798_ /*56829*/;
assign _24802_ = _24155_ ^ _24798_ /*56832*/;
assign _24803_ = _24794_ & _24802_ /*56830*/;
assign _24603_ = _24794_ ^ _24802_ /*56831*/;
assign _24800_ = _24801_ | _24803_ /*56828*/;
assign _24805_ = ~Q[36] /*56827*/;
assign _24804_ = _24805_ & D[27] /*56826*/;
assign _24807_ = _24156_ & _24804_ /*56821*/;
assign _24808_ = _24156_ ^ _24804_ /*56824*/;
assign _24809_ = _24800_ & _24808_ /*56822*/;
assign _24604_ = _24800_ ^ _24808_ /*56823*/;
assign _24806_ = _24807_ | _24809_ /*56820*/;
assign _24811_ = ~Q[36] /*56819*/;
assign _24810_ = _24811_ & D[28] /*56818*/;
assign _24813_ = _24157_ & _24810_ /*56813*/;
assign _24814_ = _24157_ ^ _24810_ /*56816*/;
assign _24815_ = _24806_ & _24814_ /*56814*/;
assign _24605_ = _24806_ ^ _24814_ /*56815*/;
assign _24812_ = _24813_ | _24815_ /*56812*/;
assign _24817_ = ~Q[36] /*56811*/;
assign _24816_ = _24817_ & D[29] /*56810*/;
assign _24819_ = _24158_ & _24816_ /*56805*/;
assign _24820_ = _24158_ ^ _24816_ /*56808*/;
assign _24821_ = _24812_ & _24820_ /*56806*/;
assign _24606_ = _24812_ ^ _24820_ /*56807*/;
assign _24818_ = _24819_ | _24821_ /*56804*/;
assign _24823_ = ~Q[36] /*56803*/;
assign _24822_ = _24823_ & D[30] /*56802*/;
assign _24825_ = _24159_ & _24822_ /*56797*/;
assign _24826_ = _24159_ ^ _24822_ /*56800*/;
assign _24827_ = _24818_ & _24826_ /*56798*/;
assign _24607_ = _24818_ ^ _24826_ /*56799*/;
assign _24824_ = _24825_ | _24827_ /*56796*/;
assign _24829_ = ~Q[36] /*56795*/;
assign _24828_ = _24829_ & D[31] /*56794*/;
assign _24831_ = _24160_ & _24828_ /*56789*/;
assign _24832_ = _24160_ ^ _24828_ /*56792*/;
assign _24833_ = _24824_ & _24832_ /*56790*/;
assign _24608_ = _24824_ ^ _24832_ /*56791*/;
assign _24830_ = _24831_ | _24833_ /*56788*/;
assign _24835_ = ~Q[36] /*56787*/;
assign _24834_ = _24835_ & D[32] /*56786*/;
assign _24837_ = _24161_ & _24834_ /*56781*/;
assign _24838_ = _24161_ ^ _24834_ /*56784*/;
assign _24839_ = _24830_ & _24838_ /*56782*/;
assign _24609_ = _24830_ ^ _24838_ /*56783*/;
assign _24836_ = _24837_ | _24839_ /*56780*/;
assign _24841_ = ~Q[36] /*56779*/;
assign _24840_ = _24841_ & D[33] /*56778*/;
assign _24843_ = _24162_ & _24840_ /*56773*/;
assign _24844_ = _24162_ ^ _24840_ /*56776*/;
assign _24845_ = _24836_ & _24844_ /*56774*/;
assign _24610_ = _24836_ ^ _24844_ /*56775*/;
assign _24842_ = _24843_ | _24845_ /*56772*/;
assign _24847_ = ~Q[36] /*56771*/;
assign _24846_ = _24847_ & D[34] /*56770*/;
assign _24849_ = _24163_ & _24846_ /*56765*/;
assign _24850_ = _24163_ ^ _24846_ /*56768*/;
assign _24851_ = _24842_ & _24850_ /*56766*/;
assign _24611_ = _24842_ ^ _24850_ /*56767*/;
assign _24848_ = _24849_ | _24851_ /*56764*/;
assign _24853_ = ~Q[36] /*56763*/;
assign _24852_ = _24853_ & D[35] /*56762*/;
assign _24855_ = _24164_ & _24852_ /*56757*/;
assign _24856_ = _24164_ ^ _24852_ /*56760*/;
assign _24857_ = _24848_ & _24856_ /*56758*/;
assign _24612_ = _24848_ ^ _24856_ /*56759*/;
assign _24854_ = _24855_ | _24857_ /*56756*/;
assign _24859_ = ~Q[36] /*56755*/;
assign _24858_ = _24859_ & D[36] /*56754*/;
assign _24861_ = _24165_ & _24858_ /*56749*/;
assign _24862_ = _24165_ ^ _24858_ /*56752*/;
assign _24863_ = _24854_ & _24862_ /*56750*/;
assign _24613_ = _24854_ ^ _24862_ /*56751*/;
assign _24860_ = _24861_ | _24863_ /*56748*/;
assign _24865_ = ~Q[36] /*56747*/;
assign _24864_ = _24865_ & D[37] /*56746*/;
assign _24867_ = _24166_ & _24864_ /*56741*/;
assign _24868_ = _24166_ ^ _24864_ /*56744*/;
assign _24869_ = _24860_ & _24868_ /*56742*/;
assign _24614_ = _24860_ ^ _24868_ /*56743*/;
assign _24866_ = _24867_ | _24869_ /*56740*/;
assign _24871_ = ~Q[36] /*56739*/;
assign _24870_ = _24871_ & D[38] /*56738*/;
assign _24873_ = _24167_ & _24870_ /*56733*/;
assign _24874_ = _24167_ ^ _24870_ /*56736*/;
assign _24875_ = _24866_ & _24874_ /*56734*/;
assign _24615_ = _24866_ ^ _24874_ /*56735*/;
assign _24872_ = _24873_ | _24875_ /*56732*/;
assign _24877_ = ~Q[36] /*56731*/;
assign _24876_ = _24877_ & D[39] /*56730*/;
assign _24879_ = _24168_ & _24876_ /*56725*/;
assign _24880_ = _24168_ ^ _24876_ /*56728*/;
assign _24881_ = _24872_ & _24880_ /*56726*/;
assign _24616_ = _24872_ ^ _24880_ /*56727*/;
assign _24878_ = _24879_ | _24881_ /*56724*/;
assign _24883_ = ~Q[36] /*56723*/;
assign _24882_ = _24883_ & D[40] /*56722*/;
assign _24885_ = _24169_ & _24882_ /*56717*/;
assign _24886_ = _24169_ ^ _24882_ /*56720*/;
assign _24887_ = _24878_ & _24886_ /*56718*/;
assign _24617_ = _24878_ ^ _24886_ /*56719*/;
assign _24884_ = _24885_ | _24887_ /*56716*/;
assign _24889_ = ~Q[36] /*56715*/;
assign _24888_ = _24889_ & D[41] /*56714*/;
assign _24891_ = _24170_ & _24888_ /*56709*/;
assign _24892_ = _24170_ ^ _24888_ /*56712*/;
assign _24893_ = _24884_ & _24892_ /*56710*/;
assign _24618_ = _24884_ ^ _24892_ /*56711*/;
assign _24890_ = _24891_ | _24893_ /*56708*/;
assign _24895_ = ~Q[36] /*56707*/;
assign _24894_ = _24895_ & D[42] /*56706*/;
assign _24897_ = _24171_ & _24894_ /*56701*/;
assign _24898_ = _24171_ ^ _24894_ /*56704*/;
assign _24899_ = _24890_ & _24898_ /*56702*/;
assign _24619_ = _24890_ ^ _24898_ /*56703*/;
assign _24896_ = _24897_ | _24899_ /*56700*/;
assign _24901_ = ~Q[36] /*56699*/;
assign _24900_ = _24901_ & D[43] /*56698*/;
assign _24903_ = _24172_ & _24900_ /*56693*/;
assign _24904_ = _24172_ ^ _24900_ /*56696*/;
assign _24905_ = _24896_ & _24904_ /*56694*/;
assign _24620_ = _24896_ ^ _24904_ /*56695*/;
assign _24902_ = _24903_ | _24905_ /*56692*/;
assign _24907_ = ~Q[36] /*56691*/;
assign _24906_ = _24907_ & D[44] /*56690*/;
assign _24909_ = _24173_ & _24906_ /*56685*/;
assign _24910_ = _24173_ ^ _24906_ /*56688*/;
assign _24911_ = _24902_ & _24910_ /*56686*/;
assign _24621_ = _24902_ ^ _24910_ /*56687*/;
assign _24908_ = _24909_ | _24911_ /*56684*/;
assign _24913_ = ~Q[36] /*56683*/;
assign _24912_ = _24913_ & D[45] /*56682*/;
assign _24915_ = _24174_ & _24912_ /*56677*/;
assign _24916_ = _24174_ ^ _24912_ /*56680*/;
assign _24917_ = _24908_ & _24916_ /*56678*/;
assign _24622_ = _24908_ ^ _24916_ /*56679*/;
assign _24914_ = _24915_ | _24917_ /*56676*/;
assign _24919_ = ~Q[36] /*56675*/;
assign _24918_ = _24919_ & D[46] /*56674*/;
assign _24921_ = _24175_ & _24918_ /*56669*/;
assign _24922_ = _24175_ ^ _24918_ /*56672*/;
assign _24923_ = _24914_ & _24922_ /*56670*/;
assign _24623_ = _24914_ ^ _24922_ /*56671*/;
assign _24920_ = _24921_ | _24923_ /*56668*/;
assign _24925_ = ~Q[36] /*56667*/;
assign _24924_ = _24925_ & D[47] /*56666*/;
assign _24927_ = _24176_ & _24924_ /*56661*/;
assign _24928_ = _24176_ ^ _24924_ /*56664*/;
assign _24929_ = _24920_ & _24928_ /*56662*/;
assign _24624_ = _24920_ ^ _24928_ /*56663*/;
assign _24926_ = _24927_ | _24929_ /*56660*/;
assign _24931_ = ~Q[36] /*56659*/;
assign _24930_ = _24931_ & D[48] /*56658*/;
assign _24933_ = _24177_ & _24930_ /*56653*/;
assign _24934_ = _24177_ ^ _24930_ /*56656*/;
assign _24935_ = _24926_ & _24934_ /*56654*/;
assign _24625_ = _24926_ ^ _24934_ /*56655*/;
assign _24932_ = _24933_ | _24935_ /*56652*/;
assign _24937_ = ~Q[36] /*56651*/;
assign _24936_ = _24937_ & D[49] /*56650*/;
assign _24939_ = _24178_ & _24936_ /*56645*/;
assign _24940_ = _24178_ ^ _24936_ /*56648*/;
assign _24941_ = _24932_ & _24940_ /*56646*/;
assign _24626_ = _24932_ ^ _24940_ /*56647*/;
assign _24938_ = _24939_ | _24941_ /*56644*/;
assign _24943_ = ~Q[36] /*56643*/;
assign _24942_ = _24943_ & D[50] /*56642*/;
assign _24945_ = _24179_ & _24942_ /*56637*/;
assign _24946_ = _24179_ ^ _24942_ /*56640*/;
assign _24947_ = _24938_ & _24946_ /*56638*/;
assign _24627_ = _24938_ ^ _24946_ /*56639*/;
assign _24944_ = _24945_ | _24947_ /*56636*/;
assign _24949_ = ~Q[36] /*56635*/;
assign _24948_ = _24949_ & D[51] /*56634*/;
assign _24951_ = _24180_ & _24948_ /*56629*/;
assign _24952_ = _24180_ ^ _24948_ /*56632*/;
assign _24953_ = _24944_ & _24952_ /*56630*/;
assign _24628_ = _24944_ ^ _24952_ /*56631*/;
assign _24950_ = _24951_ | _24953_ /*56628*/;
assign _24955_ = ~Q[36] /*56627*/;
assign _24954_ = _24955_ & D[52] /*56626*/;
assign _24957_ = _24181_ & _24954_ /*56621*/;
assign _24958_ = _24181_ ^ _24954_ /*56624*/;
assign _24959_ = _24950_ & _24958_ /*56622*/;
assign _24629_ = _24950_ ^ _24958_ /*56623*/;
assign _24956_ = _24957_ | _24959_ /*56620*/;
assign _24961_ = ~Q[36] /*56619*/;
assign _24960_ = _24961_ & D[53] /*56618*/;
assign _24963_ = _24182_ & _24960_ /*56613*/;
assign _24964_ = _24182_ ^ _24960_ /*56616*/;
assign _24965_ = _24956_ & _24964_ /*56614*/;
assign _24630_ = _24956_ ^ _24964_ /*56615*/;
assign _24962_ = _24963_ | _24965_ /*56612*/;
assign _24967_ = ~Q[36] /*56611*/;
assign _24966_ = _24967_ & D[54] /*56610*/;
assign _24969_ = _24183_ & _24966_ /*56605*/;
assign _24970_ = _24183_ ^ _24966_ /*56608*/;
assign _24971_ = _24962_ & _24970_ /*56606*/;
assign _24631_ = _24962_ ^ _24970_ /*56607*/;
assign _24968_ = _24969_ | _24971_ /*56604*/;
assign _24973_ = ~Q[36] /*56603*/;
assign _24972_ = _24973_ & D[55] /*56602*/;
assign _24975_ = _24184_ & _24972_ /*56597*/;
assign _24976_ = _24184_ ^ _24972_ /*56600*/;
assign _24977_ = _24968_ & _24976_ /*56598*/;
assign _24632_ = _24968_ ^ _24976_ /*56599*/;
assign _24974_ = _24975_ | _24977_ /*56596*/;
assign _24979_ = ~Q[36] /*56595*/;
assign _24978_ = _24979_ & D[56] /*56594*/;
assign _24981_ = _24185_ & _24978_ /*56589*/;
assign _24982_ = _24185_ ^ _24978_ /*56592*/;
assign _24983_ = _24974_ & _24982_ /*56590*/;
assign _24633_ = _24974_ ^ _24982_ /*56591*/;
assign _24980_ = _24981_ | _24983_ /*56588*/;
assign _24985_ = ~Q[36] /*56587*/;
assign _24984_ = _24985_ & D[57] /*56586*/;
assign _24987_ = _24186_ & _24984_ /*56581*/;
assign _24988_ = _24186_ ^ _24984_ /*56584*/;
assign _24989_ = _24980_ & _24988_ /*56582*/;
assign _24634_ = _24980_ ^ _24988_ /*56583*/;
assign _24986_ = _24987_ | _24989_ /*56580*/;
assign _24991_ = ~Q[36] /*56579*/;
assign _24990_ = _24991_ & D[58] /*56578*/;
assign _24993_ = _24187_ & _24990_ /*56573*/;
assign _24994_ = _24187_ ^ _24990_ /*56576*/;
assign _24995_ = _24986_ & _24994_ /*56574*/;
assign _24635_ = _24986_ ^ _24994_ /*56575*/;
assign _24992_ = _24993_ | _24995_ /*56572*/;
assign _24997_ = ~Q[36] /*56571*/;
assign _24996_ = _24997_ & D[59] /*56570*/;
assign _24999_ = _24188_ & _24996_ /*56565*/;
assign _25000_ = _24188_ ^ _24996_ /*56568*/;
assign _25001_ = _24992_ & _25000_ /*56566*/;
assign _24636_ = _24992_ ^ _25000_ /*56567*/;
assign _24998_ = _24999_ | _25001_ /*56564*/;
assign _25003_ = ~Q[36] /*56563*/;
assign _25002_ = _25003_ & D[60] /*56562*/;
assign _25005_ = _24189_ & _25002_ /*56557*/;
assign _25006_ = _24189_ ^ _25002_ /*56560*/;
assign _25007_ = _24998_ & _25006_ /*56558*/;
assign _24637_ = _24998_ ^ _25006_ /*56559*/;
assign _25004_ = _25005_ | _25007_ /*56556*/;
assign _25009_ = ~Q[36] /*56555*/;
assign _25008_ = _25009_ & D[61] /*56554*/;
assign _25011_ = _24190_ & _25008_ /*56549*/;
assign _25012_ = _24190_ ^ _25008_ /*56552*/;
assign _25013_ = _25004_ & _25012_ /*56550*/;
assign _24638_ = _25004_ ^ _25012_ /*56551*/;
assign _25010_ = _25011_ | _25013_ /*56548*/;
assign _25015_ = ~Q[36] /*56547*/;
assign _25014_ = _25015_ & D[62] /*56546*/;
assign _25017_ = _24191_ & _25014_ /*56541*/;
assign _25018_ = _24191_ ^ _25014_ /*56544*/;
assign _25019_ = _25010_ & _25018_ /*56542*/;
assign _24639_ = _25010_ ^ _25018_ /*56543*/;
assign _25016_ = _25017_ | _25019_ /*56540*/;
assign _25021_ = ~Q[36] /*56539*/;
assign _25020_ = _25021_ & zeroWire /*56538*/;
assign _25022_ = _24192_ ^ _25020_ /*56536*/;
assign _24640_ = _25022_ ^ _25016_ /*56535*/;
assign _25093_ = ~D[0] /*56281*/;
assign _25090_ = R_0[35] & _25093_ /*56277*/;
assign _25091_ = R_0[35] ^ _25093_ /*56280*/;
assign _25092_ = oneWire & _25091_ /*56278*/;
assign _25025_ = oneWire ^ _25091_ /*56279*/;
assign _25089_ = _25090_ | _25092_ /*56276*/;
assign _25098_ = ~D[1] /*56275*/;
assign _25095_ = _24577_ & _25098_ /*56271*/;
assign _25096_ = _24577_ ^ _25098_ /*56274*/;
assign _25097_ = _25089_ & _25096_ /*56272*/;
assign _25026_ = _25089_ ^ _25096_ /*56273*/;
assign _25094_ = _25095_ | _25097_ /*56270*/;
assign _25103_ = ~D[2] /*56269*/;
assign _25100_ = _24578_ & _25103_ /*56265*/;
assign _25101_ = _24578_ ^ _25103_ /*56268*/;
assign _25102_ = _25094_ & _25101_ /*56266*/;
assign _25027_ = _25094_ ^ _25101_ /*56267*/;
assign _25099_ = _25100_ | _25102_ /*56264*/;
assign _25108_ = ~D[3] /*56263*/;
assign _25105_ = _24579_ & _25108_ /*56259*/;
assign _25106_ = _24579_ ^ _25108_ /*56262*/;
assign _25107_ = _25099_ & _25106_ /*56260*/;
assign _25028_ = _25099_ ^ _25106_ /*56261*/;
assign _25104_ = _25105_ | _25107_ /*56258*/;
assign _25113_ = ~D[4] /*56257*/;
assign _25110_ = _24580_ & _25113_ /*56253*/;
assign _25111_ = _24580_ ^ _25113_ /*56256*/;
assign _25112_ = _25104_ & _25111_ /*56254*/;
assign _25029_ = _25104_ ^ _25111_ /*56255*/;
assign _25109_ = _25110_ | _25112_ /*56252*/;
assign _25118_ = ~D[5] /*56251*/;
assign _25115_ = _24581_ & _25118_ /*56247*/;
assign _25116_ = _24581_ ^ _25118_ /*56250*/;
assign _25117_ = _25109_ & _25116_ /*56248*/;
assign _25030_ = _25109_ ^ _25116_ /*56249*/;
assign _25114_ = _25115_ | _25117_ /*56246*/;
assign _25123_ = ~D[6] /*56245*/;
assign _25120_ = _24582_ & _25123_ /*56241*/;
assign _25121_ = _24582_ ^ _25123_ /*56244*/;
assign _25122_ = _25114_ & _25121_ /*56242*/;
assign _25031_ = _25114_ ^ _25121_ /*56243*/;
assign _25119_ = _25120_ | _25122_ /*56240*/;
assign _25128_ = ~D[7] /*56239*/;
assign _25125_ = _24583_ & _25128_ /*56235*/;
assign _25126_ = _24583_ ^ _25128_ /*56238*/;
assign _25127_ = _25119_ & _25126_ /*56236*/;
assign _25032_ = _25119_ ^ _25126_ /*56237*/;
assign _25124_ = _25125_ | _25127_ /*56234*/;
assign _25133_ = ~D[8] /*56233*/;
assign _25130_ = _24584_ & _25133_ /*56229*/;
assign _25131_ = _24584_ ^ _25133_ /*56232*/;
assign _25132_ = _25124_ & _25131_ /*56230*/;
assign _25033_ = _25124_ ^ _25131_ /*56231*/;
assign _25129_ = _25130_ | _25132_ /*56228*/;
assign _25138_ = ~D[9] /*56227*/;
assign _25135_ = _24585_ & _25138_ /*56223*/;
assign _25136_ = _24585_ ^ _25138_ /*56226*/;
assign _25137_ = _25129_ & _25136_ /*56224*/;
assign _25034_ = _25129_ ^ _25136_ /*56225*/;
assign _25134_ = _25135_ | _25137_ /*56222*/;
assign _25143_ = ~D[10] /*56221*/;
assign _25140_ = _24586_ & _25143_ /*56217*/;
assign _25141_ = _24586_ ^ _25143_ /*56220*/;
assign _25142_ = _25134_ & _25141_ /*56218*/;
assign _25035_ = _25134_ ^ _25141_ /*56219*/;
assign _25139_ = _25140_ | _25142_ /*56216*/;
assign _25148_ = ~D[11] /*56215*/;
assign _25145_ = _24587_ & _25148_ /*56211*/;
assign _25146_ = _24587_ ^ _25148_ /*56214*/;
assign _25147_ = _25139_ & _25146_ /*56212*/;
assign _25036_ = _25139_ ^ _25146_ /*56213*/;
assign _25144_ = _25145_ | _25147_ /*56210*/;
assign _25153_ = ~D[12] /*56209*/;
assign _25150_ = _24588_ & _25153_ /*56205*/;
assign _25151_ = _24588_ ^ _25153_ /*56208*/;
assign _25152_ = _25144_ & _25151_ /*56206*/;
assign _25037_ = _25144_ ^ _25151_ /*56207*/;
assign _25149_ = _25150_ | _25152_ /*56204*/;
assign _25158_ = ~D[13] /*56203*/;
assign _25155_ = _24589_ & _25158_ /*56199*/;
assign _25156_ = _24589_ ^ _25158_ /*56202*/;
assign _25157_ = _25149_ & _25156_ /*56200*/;
assign _25038_ = _25149_ ^ _25156_ /*56201*/;
assign _25154_ = _25155_ | _25157_ /*56198*/;
assign _25163_ = ~D[14] /*56197*/;
assign _25160_ = _24590_ & _25163_ /*56193*/;
assign _25161_ = _24590_ ^ _25163_ /*56196*/;
assign _25162_ = _25154_ & _25161_ /*56194*/;
assign _25039_ = _25154_ ^ _25161_ /*56195*/;
assign _25159_ = _25160_ | _25162_ /*56192*/;
assign _25168_ = ~D[15] /*56191*/;
assign _25165_ = _24591_ & _25168_ /*56187*/;
assign _25166_ = _24591_ ^ _25168_ /*56190*/;
assign _25167_ = _25159_ & _25166_ /*56188*/;
assign _25040_ = _25159_ ^ _25166_ /*56189*/;
assign _25164_ = _25165_ | _25167_ /*56186*/;
assign _25173_ = ~D[16] /*56185*/;
assign _25170_ = _24592_ & _25173_ /*56181*/;
assign _25171_ = _24592_ ^ _25173_ /*56184*/;
assign _25172_ = _25164_ & _25171_ /*56182*/;
assign _25041_ = _25164_ ^ _25171_ /*56183*/;
assign _25169_ = _25170_ | _25172_ /*56180*/;
assign _25178_ = ~D[17] /*56179*/;
assign _25175_ = _24593_ & _25178_ /*56175*/;
assign _25176_ = _24593_ ^ _25178_ /*56178*/;
assign _25177_ = _25169_ & _25176_ /*56176*/;
assign _25042_ = _25169_ ^ _25176_ /*56177*/;
assign _25174_ = _25175_ | _25177_ /*56174*/;
assign _25183_ = ~D[18] /*56173*/;
assign _25180_ = _24594_ & _25183_ /*56169*/;
assign _25181_ = _24594_ ^ _25183_ /*56172*/;
assign _25182_ = _25174_ & _25181_ /*56170*/;
assign _25043_ = _25174_ ^ _25181_ /*56171*/;
assign _25179_ = _25180_ | _25182_ /*56168*/;
assign _25188_ = ~D[19] /*56167*/;
assign _25185_ = _24595_ & _25188_ /*56163*/;
assign _25186_ = _24595_ ^ _25188_ /*56166*/;
assign _25187_ = _25179_ & _25186_ /*56164*/;
assign _25044_ = _25179_ ^ _25186_ /*56165*/;
assign _25184_ = _25185_ | _25187_ /*56162*/;
assign _25193_ = ~D[20] /*56161*/;
assign _25190_ = _24596_ & _25193_ /*56157*/;
assign _25191_ = _24596_ ^ _25193_ /*56160*/;
assign _25192_ = _25184_ & _25191_ /*56158*/;
assign _25045_ = _25184_ ^ _25191_ /*56159*/;
assign _25189_ = _25190_ | _25192_ /*56156*/;
assign _25198_ = ~D[21] /*56155*/;
assign _25195_ = _24597_ & _25198_ /*56151*/;
assign _25196_ = _24597_ ^ _25198_ /*56154*/;
assign _25197_ = _25189_ & _25196_ /*56152*/;
assign _25046_ = _25189_ ^ _25196_ /*56153*/;
assign _25194_ = _25195_ | _25197_ /*56150*/;
assign _25203_ = ~D[22] /*56149*/;
assign _25200_ = _24598_ & _25203_ /*56145*/;
assign _25201_ = _24598_ ^ _25203_ /*56148*/;
assign _25202_ = _25194_ & _25201_ /*56146*/;
assign _25047_ = _25194_ ^ _25201_ /*56147*/;
assign _25199_ = _25200_ | _25202_ /*56144*/;
assign _25208_ = ~D[23] /*56143*/;
assign _25205_ = _24599_ & _25208_ /*56139*/;
assign _25206_ = _24599_ ^ _25208_ /*56142*/;
assign _25207_ = _25199_ & _25206_ /*56140*/;
assign _25048_ = _25199_ ^ _25206_ /*56141*/;
assign _25204_ = _25205_ | _25207_ /*56138*/;
assign _25213_ = ~D[24] /*56137*/;
assign _25210_ = _24600_ & _25213_ /*56133*/;
assign _25211_ = _24600_ ^ _25213_ /*56136*/;
assign _25212_ = _25204_ & _25211_ /*56134*/;
assign _25049_ = _25204_ ^ _25211_ /*56135*/;
assign _25209_ = _25210_ | _25212_ /*56132*/;
assign _25218_ = ~D[25] /*56131*/;
assign _25215_ = _24601_ & _25218_ /*56127*/;
assign _25216_ = _24601_ ^ _25218_ /*56130*/;
assign _25217_ = _25209_ & _25216_ /*56128*/;
assign _25050_ = _25209_ ^ _25216_ /*56129*/;
assign _25214_ = _25215_ | _25217_ /*56126*/;
assign _25223_ = ~D[26] /*56125*/;
assign _25220_ = _24602_ & _25223_ /*56121*/;
assign _25221_ = _24602_ ^ _25223_ /*56124*/;
assign _25222_ = _25214_ & _25221_ /*56122*/;
assign _25051_ = _25214_ ^ _25221_ /*56123*/;
assign _25219_ = _25220_ | _25222_ /*56120*/;
assign _25228_ = ~D[27] /*56119*/;
assign _25225_ = _24603_ & _25228_ /*56115*/;
assign _25226_ = _24603_ ^ _25228_ /*56118*/;
assign _25227_ = _25219_ & _25226_ /*56116*/;
assign _25052_ = _25219_ ^ _25226_ /*56117*/;
assign _25224_ = _25225_ | _25227_ /*56114*/;
assign _25233_ = ~D[28] /*56113*/;
assign _25230_ = _24604_ & _25233_ /*56109*/;
assign _25231_ = _24604_ ^ _25233_ /*56112*/;
assign _25232_ = _25224_ & _25231_ /*56110*/;
assign _25053_ = _25224_ ^ _25231_ /*56111*/;
assign _25229_ = _25230_ | _25232_ /*56108*/;
assign _25238_ = ~D[29] /*56107*/;
assign _25235_ = _24605_ & _25238_ /*56103*/;
assign _25236_ = _24605_ ^ _25238_ /*56106*/;
assign _25237_ = _25229_ & _25236_ /*56104*/;
assign _25054_ = _25229_ ^ _25236_ /*56105*/;
assign _25234_ = _25235_ | _25237_ /*56102*/;
assign _25243_ = ~D[30] /*56101*/;
assign _25240_ = _24606_ & _25243_ /*56097*/;
assign _25241_ = _24606_ ^ _25243_ /*56100*/;
assign _25242_ = _25234_ & _25241_ /*56098*/;
assign _25055_ = _25234_ ^ _25241_ /*56099*/;
assign _25239_ = _25240_ | _25242_ /*56096*/;
assign _25248_ = ~D[31] /*56095*/;
assign _25245_ = _24607_ & _25248_ /*56091*/;
assign _25246_ = _24607_ ^ _25248_ /*56094*/;
assign _25247_ = _25239_ & _25246_ /*56092*/;
assign _25056_ = _25239_ ^ _25246_ /*56093*/;
assign _25244_ = _25245_ | _25247_ /*56090*/;
assign _25253_ = ~D[32] /*56089*/;
assign _25250_ = _24608_ & _25253_ /*56085*/;
assign _25251_ = _24608_ ^ _25253_ /*56088*/;
assign _25252_ = _25244_ & _25251_ /*56086*/;
assign _25057_ = _25244_ ^ _25251_ /*56087*/;
assign _25249_ = _25250_ | _25252_ /*56084*/;
assign _25258_ = ~D[33] /*56083*/;
assign _25255_ = _24609_ & _25258_ /*56079*/;
assign _25256_ = _24609_ ^ _25258_ /*56082*/;
assign _25257_ = _25249_ & _25256_ /*56080*/;
assign _25058_ = _25249_ ^ _25256_ /*56081*/;
assign _25254_ = _25255_ | _25257_ /*56078*/;
assign _25263_ = ~D[34] /*56077*/;
assign _25260_ = _24610_ & _25263_ /*56073*/;
assign _25261_ = _24610_ ^ _25263_ /*56076*/;
assign _25262_ = _25254_ & _25261_ /*56074*/;
assign _25059_ = _25254_ ^ _25261_ /*56075*/;
assign _25259_ = _25260_ | _25262_ /*56072*/;
assign _25268_ = ~D[35] /*56071*/;
assign _25265_ = _24611_ & _25268_ /*56067*/;
assign _25266_ = _24611_ ^ _25268_ /*56070*/;
assign _25267_ = _25259_ & _25266_ /*56068*/;
assign _25060_ = _25259_ ^ _25266_ /*56069*/;
assign _25264_ = _25265_ | _25267_ /*56066*/;
assign _25273_ = ~D[36] /*56065*/;
assign _25270_ = _24612_ & _25273_ /*56061*/;
assign _25271_ = _24612_ ^ _25273_ /*56064*/;
assign _25272_ = _25264_ & _25271_ /*56062*/;
assign _25061_ = _25264_ ^ _25271_ /*56063*/;
assign _25269_ = _25270_ | _25272_ /*56060*/;
assign _25278_ = ~D[37] /*56059*/;
assign _25275_ = _24613_ & _25278_ /*56055*/;
assign _25276_ = _24613_ ^ _25278_ /*56058*/;
assign _25277_ = _25269_ & _25276_ /*56056*/;
assign _25062_ = _25269_ ^ _25276_ /*56057*/;
assign _25274_ = _25275_ | _25277_ /*56054*/;
assign _25283_ = ~D[38] /*56053*/;
assign _25280_ = _24614_ & _25283_ /*56049*/;
assign _25281_ = _24614_ ^ _25283_ /*56052*/;
assign _25282_ = _25274_ & _25281_ /*56050*/;
assign _25063_ = _25274_ ^ _25281_ /*56051*/;
assign _25279_ = _25280_ | _25282_ /*56048*/;
assign _25288_ = ~D[39] /*56047*/;
assign _25285_ = _24615_ & _25288_ /*56043*/;
assign _25286_ = _24615_ ^ _25288_ /*56046*/;
assign _25287_ = _25279_ & _25286_ /*56044*/;
assign _25064_ = _25279_ ^ _25286_ /*56045*/;
assign _25284_ = _25285_ | _25287_ /*56042*/;
assign _25293_ = ~D[40] /*56041*/;
assign _25290_ = _24616_ & _25293_ /*56037*/;
assign _25291_ = _24616_ ^ _25293_ /*56040*/;
assign _25292_ = _25284_ & _25291_ /*56038*/;
assign _25065_ = _25284_ ^ _25291_ /*56039*/;
assign _25289_ = _25290_ | _25292_ /*56036*/;
assign _25298_ = ~D[41] /*56035*/;
assign _25295_ = _24617_ & _25298_ /*56031*/;
assign _25296_ = _24617_ ^ _25298_ /*56034*/;
assign _25297_ = _25289_ & _25296_ /*56032*/;
assign _25066_ = _25289_ ^ _25296_ /*56033*/;
assign _25294_ = _25295_ | _25297_ /*56030*/;
assign _25303_ = ~D[42] /*56029*/;
assign _25300_ = _24618_ & _25303_ /*56025*/;
assign _25301_ = _24618_ ^ _25303_ /*56028*/;
assign _25302_ = _25294_ & _25301_ /*56026*/;
assign _25067_ = _25294_ ^ _25301_ /*56027*/;
assign _25299_ = _25300_ | _25302_ /*56024*/;
assign _25308_ = ~D[43] /*56023*/;
assign _25305_ = _24619_ & _25308_ /*56019*/;
assign _25306_ = _24619_ ^ _25308_ /*56022*/;
assign _25307_ = _25299_ & _25306_ /*56020*/;
assign _25068_ = _25299_ ^ _25306_ /*56021*/;
assign _25304_ = _25305_ | _25307_ /*56018*/;
assign _25313_ = ~D[44] /*56017*/;
assign _25310_ = _24620_ & _25313_ /*56013*/;
assign _25311_ = _24620_ ^ _25313_ /*56016*/;
assign _25312_ = _25304_ & _25311_ /*56014*/;
assign _25069_ = _25304_ ^ _25311_ /*56015*/;
assign _25309_ = _25310_ | _25312_ /*56012*/;
assign _25318_ = ~D[45] /*56011*/;
assign _25315_ = _24621_ & _25318_ /*56007*/;
assign _25316_ = _24621_ ^ _25318_ /*56010*/;
assign _25317_ = _25309_ & _25316_ /*56008*/;
assign _25070_ = _25309_ ^ _25316_ /*56009*/;
assign _25314_ = _25315_ | _25317_ /*56006*/;
assign _25323_ = ~D[46] /*56005*/;
assign _25320_ = _24622_ & _25323_ /*56001*/;
assign _25321_ = _24622_ ^ _25323_ /*56004*/;
assign _25322_ = _25314_ & _25321_ /*56002*/;
assign _25071_ = _25314_ ^ _25321_ /*56003*/;
assign _25319_ = _25320_ | _25322_ /*56000*/;
assign _25328_ = ~D[47] /*55999*/;
assign _25325_ = _24623_ & _25328_ /*55995*/;
assign _25326_ = _24623_ ^ _25328_ /*55998*/;
assign _25327_ = _25319_ & _25326_ /*55996*/;
assign _25072_ = _25319_ ^ _25326_ /*55997*/;
assign _25324_ = _25325_ | _25327_ /*55994*/;
assign _25333_ = ~D[48] /*55993*/;
assign _25330_ = _24624_ & _25333_ /*55989*/;
assign _25331_ = _24624_ ^ _25333_ /*55992*/;
assign _25332_ = _25324_ & _25331_ /*55990*/;
assign _25073_ = _25324_ ^ _25331_ /*55991*/;
assign _25329_ = _25330_ | _25332_ /*55988*/;
assign _25338_ = ~D[49] /*55987*/;
assign _25335_ = _24625_ & _25338_ /*55983*/;
assign _25336_ = _24625_ ^ _25338_ /*55986*/;
assign _25337_ = _25329_ & _25336_ /*55984*/;
assign _25074_ = _25329_ ^ _25336_ /*55985*/;
assign _25334_ = _25335_ | _25337_ /*55982*/;
assign _25343_ = ~D[50] /*55981*/;
assign _25340_ = _24626_ & _25343_ /*55977*/;
assign _25341_ = _24626_ ^ _25343_ /*55980*/;
assign _25342_ = _25334_ & _25341_ /*55978*/;
assign _25075_ = _25334_ ^ _25341_ /*55979*/;
assign _25339_ = _25340_ | _25342_ /*55976*/;
assign _25348_ = ~D[51] /*55975*/;
assign _25345_ = _24627_ & _25348_ /*55971*/;
assign _25346_ = _24627_ ^ _25348_ /*55974*/;
assign _25347_ = _25339_ & _25346_ /*55972*/;
assign _25076_ = _25339_ ^ _25346_ /*55973*/;
assign _25344_ = _25345_ | _25347_ /*55970*/;
assign _25353_ = ~D[52] /*55969*/;
assign _25350_ = _24628_ & _25353_ /*55965*/;
assign _25351_ = _24628_ ^ _25353_ /*55968*/;
assign _25352_ = _25344_ & _25351_ /*55966*/;
assign _25077_ = _25344_ ^ _25351_ /*55967*/;
assign _25349_ = _25350_ | _25352_ /*55964*/;
assign _25358_ = ~D[53] /*55963*/;
assign _25355_ = _24629_ & _25358_ /*55959*/;
assign _25356_ = _24629_ ^ _25358_ /*55962*/;
assign _25357_ = _25349_ & _25356_ /*55960*/;
assign _25078_ = _25349_ ^ _25356_ /*55961*/;
assign _25354_ = _25355_ | _25357_ /*55958*/;
assign _25363_ = ~D[54] /*55957*/;
assign _25360_ = _24630_ & _25363_ /*55953*/;
assign _25361_ = _24630_ ^ _25363_ /*55956*/;
assign _25362_ = _25354_ & _25361_ /*55954*/;
assign _25079_ = _25354_ ^ _25361_ /*55955*/;
assign _25359_ = _25360_ | _25362_ /*55952*/;
assign _25368_ = ~D[55] /*55951*/;
assign _25365_ = _24631_ & _25368_ /*55947*/;
assign _25366_ = _24631_ ^ _25368_ /*55950*/;
assign _25367_ = _25359_ & _25366_ /*55948*/;
assign _25080_ = _25359_ ^ _25366_ /*55949*/;
assign _25364_ = _25365_ | _25367_ /*55946*/;
assign _25373_ = ~D[56] /*55945*/;
assign _25370_ = _24632_ & _25373_ /*55941*/;
assign _25371_ = _24632_ ^ _25373_ /*55944*/;
assign _25372_ = _25364_ & _25371_ /*55942*/;
assign _25081_ = _25364_ ^ _25371_ /*55943*/;
assign _25369_ = _25370_ | _25372_ /*55940*/;
assign _25378_ = ~D[57] /*55939*/;
assign _25375_ = _24633_ & _25378_ /*55935*/;
assign _25376_ = _24633_ ^ _25378_ /*55938*/;
assign _25377_ = _25369_ & _25376_ /*55936*/;
assign _25082_ = _25369_ ^ _25376_ /*55937*/;
assign _25374_ = _25375_ | _25377_ /*55934*/;
assign _25383_ = ~D[58] /*55933*/;
assign _25380_ = _24634_ & _25383_ /*55929*/;
assign _25381_ = _24634_ ^ _25383_ /*55932*/;
assign _25382_ = _25374_ & _25381_ /*55930*/;
assign _25083_ = _25374_ ^ _25381_ /*55931*/;
assign _25379_ = _25380_ | _25382_ /*55928*/;
assign _25388_ = ~D[59] /*55927*/;
assign _25385_ = _24635_ & _25388_ /*55923*/;
assign _25386_ = _24635_ ^ _25388_ /*55926*/;
assign _25387_ = _25379_ & _25386_ /*55924*/;
assign _25084_ = _25379_ ^ _25386_ /*55925*/;
assign _25384_ = _25385_ | _25387_ /*55922*/;
assign _25393_ = ~D[60] /*55921*/;
assign _25390_ = _24636_ & _25393_ /*55917*/;
assign _25391_ = _24636_ ^ _25393_ /*55920*/;
assign _25392_ = _25384_ & _25391_ /*55918*/;
assign _25085_ = _25384_ ^ _25391_ /*55919*/;
assign _25389_ = _25390_ | _25392_ /*55916*/;
assign _25398_ = ~D[61] /*55915*/;
assign _25395_ = _24637_ & _25398_ /*55911*/;
assign _25396_ = _24637_ ^ _25398_ /*55914*/;
assign _25397_ = _25389_ & _25396_ /*55912*/;
assign _25086_ = _25389_ ^ _25396_ /*55913*/;
assign _25394_ = _25395_ | _25397_ /*55910*/;
assign _25403_ = ~D[62] /*55909*/;
assign _25400_ = _24638_ & _25403_ /*55905*/;
assign _25401_ = _24638_ ^ _25403_ /*55908*/;
assign _25402_ = _25394_ & _25401_ /*55906*/;
assign _25087_ = _25394_ ^ _25401_ /*55907*/;
assign _25399_ = _25400_ | _25402_ /*55904*/;
assign _25404_ = _24639_ & oneWire /*55899*/;
assign _25405_ = _24639_ ^ oneWire /*55902*/;
assign _25406_ = _25399_ & _25405_ /*55900*/;
assign _25088_ = _25399_ ^ _25405_ /*55901*/;
assign Q[35] = _25404_ | _25406_ /*55898*/;
assign _25539_ = ~Q[35] /*55513*/;
assign _25538_ = _25539_ & D[0] /*55512*/;
assign _25541_ = _25025_ & _25538_ /*55507*/;
assign _25542_ = _25025_ ^ _25538_ /*55510*/;
assign _25543_ = zeroWire & _25542_ /*55508*/;
assign _25473_ = zeroWire ^ _25542_ /*55509*/;
assign _25540_ = _25541_ | _25543_ /*55506*/;
assign _25545_ = ~Q[35] /*55505*/;
assign _25544_ = _25545_ & D[1] /*55504*/;
assign _25547_ = _25026_ & _25544_ /*55499*/;
assign _25548_ = _25026_ ^ _25544_ /*55502*/;
assign _25549_ = _25540_ & _25548_ /*55500*/;
assign _25474_ = _25540_ ^ _25548_ /*55501*/;
assign _25546_ = _25547_ | _25549_ /*55498*/;
assign _25551_ = ~Q[35] /*55497*/;
assign _25550_ = _25551_ & D[2] /*55496*/;
assign _25553_ = _25027_ & _25550_ /*55491*/;
assign _25554_ = _25027_ ^ _25550_ /*55494*/;
assign _25555_ = _25546_ & _25554_ /*55492*/;
assign _25475_ = _25546_ ^ _25554_ /*55493*/;
assign _25552_ = _25553_ | _25555_ /*55490*/;
assign _25557_ = ~Q[35] /*55489*/;
assign _25556_ = _25557_ & D[3] /*55488*/;
assign _25559_ = _25028_ & _25556_ /*55483*/;
assign _25560_ = _25028_ ^ _25556_ /*55486*/;
assign _25561_ = _25552_ & _25560_ /*55484*/;
assign _25476_ = _25552_ ^ _25560_ /*55485*/;
assign _25558_ = _25559_ | _25561_ /*55482*/;
assign _25563_ = ~Q[35] /*55481*/;
assign _25562_ = _25563_ & D[4] /*55480*/;
assign _25565_ = _25029_ & _25562_ /*55475*/;
assign _25566_ = _25029_ ^ _25562_ /*55478*/;
assign _25567_ = _25558_ & _25566_ /*55476*/;
assign _25477_ = _25558_ ^ _25566_ /*55477*/;
assign _25564_ = _25565_ | _25567_ /*55474*/;
assign _25569_ = ~Q[35] /*55473*/;
assign _25568_ = _25569_ & D[5] /*55472*/;
assign _25571_ = _25030_ & _25568_ /*55467*/;
assign _25572_ = _25030_ ^ _25568_ /*55470*/;
assign _25573_ = _25564_ & _25572_ /*55468*/;
assign _25478_ = _25564_ ^ _25572_ /*55469*/;
assign _25570_ = _25571_ | _25573_ /*55466*/;
assign _25575_ = ~Q[35] /*55465*/;
assign _25574_ = _25575_ & D[6] /*55464*/;
assign _25577_ = _25031_ & _25574_ /*55459*/;
assign _25578_ = _25031_ ^ _25574_ /*55462*/;
assign _25579_ = _25570_ & _25578_ /*55460*/;
assign _25479_ = _25570_ ^ _25578_ /*55461*/;
assign _25576_ = _25577_ | _25579_ /*55458*/;
assign _25581_ = ~Q[35] /*55457*/;
assign _25580_ = _25581_ & D[7] /*55456*/;
assign _25583_ = _25032_ & _25580_ /*55451*/;
assign _25584_ = _25032_ ^ _25580_ /*55454*/;
assign _25585_ = _25576_ & _25584_ /*55452*/;
assign _25480_ = _25576_ ^ _25584_ /*55453*/;
assign _25582_ = _25583_ | _25585_ /*55450*/;
assign _25587_ = ~Q[35] /*55449*/;
assign _25586_ = _25587_ & D[8] /*55448*/;
assign _25589_ = _25033_ & _25586_ /*55443*/;
assign _25590_ = _25033_ ^ _25586_ /*55446*/;
assign _25591_ = _25582_ & _25590_ /*55444*/;
assign _25481_ = _25582_ ^ _25590_ /*55445*/;
assign _25588_ = _25589_ | _25591_ /*55442*/;
assign _25593_ = ~Q[35] /*55441*/;
assign _25592_ = _25593_ & D[9] /*55440*/;
assign _25595_ = _25034_ & _25592_ /*55435*/;
assign _25596_ = _25034_ ^ _25592_ /*55438*/;
assign _25597_ = _25588_ & _25596_ /*55436*/;
assign _25482_ = _25588_ ^ _25596_ /*55437*/;
assign _25594_ = _25595_ | _25597_ /*55434*/;
assign _25599_ = ~Q[35] /*55433*/;
assign _25598_ = _25599_ & D[10] /*55432*/;
assign _25601_ = _25035_ & _25598_ /*55427*/;
assign _25602_ = _25035_ ^ _25598_ /*55430*/;
assign _25603_ = _25594_ & _25602_ /*55428*/;
assign _25483_ = _25594_ ^ _25602_ /*55429*/;
assign _25600_ = _25601_ | _25603_ /*55426*/;
assign _25605_ = ~Q[35] /*55425*/;
assign _25604_ = _25605_ & D[11] /*55424*/;
assign _25607_ = _25036_ & _25604_ /*55419*/;
assign _25608_ = _25036_ ^ _25604_ /*55422*/;
assign _25609_ = _25600_ & _25608_ /*55420*/;
assign _25484_ = _25600_ ^ _25608_ /*55421*/;
assign _25606_ = _25607_ | _25609_ /*55418*/;
assign _25611_ = ~Q[35] /*55417*/;
assign _25610_ = _25611_ & D[12] /*55416*/;
assign _25613_ = _25037_ & _25610_ /*55411*/;
assign _25614_ = _25037_ ^ _25610_ /*55414*/;
assign _25615_ = _25606_ & _25614_ /*55412*/;
assign _25485_ = _25606_ ^ _25614_ /*55413*/;
assign _25612_ = _25613_ | _25615_ /*55410*/;
assign _25617_ = ~Q[35] /*55409*/;
assign _25616_ = _25617_ & D[13] /*55408*/;
assign _25619_ = _25038_ & _25616_ /*55403*/;
assign _25620_ = _25038_ ^ _25616_ /*55406*/;
assign _25621_ = _25612_ & _25620_ /*55404*/;
assign _25486_ = _25612_ ^ _25620_ /*55405*/;
assign _25618_ = _25619_ | _25621_ /*55402*/;
assign _25623_ = ~Q[35] /*55401*/;
assign _25622_ = _25623_ & D[14] /*55400*/;
assign _25625_ = _25039_ & _25622_ /*55395*/;
assign _25626_ = _25039_ ^ _25622_ /*55398*/;
assign _25627_ = _25618_ & _25626_ /*55396*/;
assign _25487_ = _25618_ ^ _25626_ /*55397*/;
assign _25624_ = _25625_ | _25627_ /*55394*/;
assign _25629_ = ~Q[35] /*55393*/;
assign _25628_ = _25629_ & D[15] /*55392*/;
assign _25631_ = _25040_ & _25628_ /*55387*/;
assign _25632_ = _25040_ ^ _25628_ /*55390*/;
assign _25633_ = _25624_ & _25632_ /*55388*/;
assign _25488_ = _25624_ ^ _25632_ /*55389*/;
assign _25630_ = _25631_ | _25633_ /*55386*/;
assign _25635_ = ~Q[35] /*55385*/;
assign _25634_ = _25635_ & D[16] /*55384*/;
assign _25637_ = _25041_ & _25634_ /*55379*/;
assign _25638_ = _25041_ ^ _25634_ /*55382*/;
assign _25639_ = _25630_ & _25638_ /*55380*/;
assign _25489_ = _25630_ ^ _25638_ /*55381*/;
assign _25636_ = _25637_ | _25639_ /*55378*/;
assign _25641_ = ~Q[35] /*55377*/;
assign _25640_ = _25641_ & D[17] /*55376*/;
assign _25643_ = _25042_ & _25640_ /*55371*/;
assign _25644_ = _25042_ ^ _25640_ /*55374*/;
assign _25645_ = _25636_ & _25644_ /*55372*/;
assign _25490_ = _25636_ ^ _25644_ /*55373*/;
assign _25642_ = _25643_ | _25645_ /*55370*/;
assign _25647_ = ~Q[35] /*55369*/;
assign _25646_ = _25647_ & D[18] /*55368*/;
assign _25649_ = _25043_ & _25646_ /*55363*/;
assign _25650_ = _25043_ ^ _25646_ /*55366*/;
assign _25651_ = _25642_ & _25650_ /*55364*/;
assign _25491_ = _25642_ ^ _25650_ /*55365*/;
assign _25648_ = _25649_ | _25651_ /*55362*/;
assign _25653_ = ~Q[35] /*55361*/;
assign _25652_ = _25653_ & D[19] /*55360*/;
assign _25655_ = _25044_ & _25652_ /*55355*/;
assign _25656_ = _25044_ ^ _25652_ /*55358*/;
assign _25657_ = _25648_ & _25656_ /*55356*/;
assign _25492_ = _25648_ ^ _25656_ /*55357*/;
assign _25654_ = _25655_ | _25657_ /*55354*/;
assign _25659_ = ~Q[35] /*55353*/;
assign _25658_ = _25659_ & D[20] /*55352*/;
assign _25661_ = _25045_ & _25658_ /*55347*/;
assign _25662_ = _25045_ ^ _25658_ /*55350*/;
assign _25663_ = _25654_ & _25662_ /*55348*/;
assign _25493_ = _25654_ ^ _25662_ /*55349*/;
assign _25660_ = _25661_ | _25663_ /*55346*/;
assign _25665_ = ~Q[35] /*55345*/;
assign _25664_ = _25665_ & D[21] /*55344*/;
assign _25667_ = _25046_ & _25664_ /*55339*/;
assign _25668_ = _25046_ ^ _25664_ /*55342*/;
assign _25669_ = _25660_ & _25668_ /*55340*/;
assign _25494_ = _25660_ ^ _25668_ /*55341*/;
assign _25666_ = _25667_ | _25669_ /*55338*/;
assign _25671_ = ~Q[35] /*55337*/;
assign _25670_ = _25671_ & D[22] /*55336*/;
assign _25673_ = _25047_ & _25670_ /*55331*/;
assign _25674_ = _25047_ ^ _25670_ /*55334*/;
assign _25675_ = _25666_ & _25674_ /*55332*/;
assign _25495_ = _25666_ ^ _25674_ /*55333*/;
assign _25672_ = _25673_ | _25675_ /*55330*/;
assign _25677_ = ~Q[35] /*55329*/;
assign _25676_ = _25677_ & D[23] /*55328*/;
assign _25679_ = _25048_ & _25676_ /*55323*/;
assign _25680_ = _25048_ ^ _25676_ /*55326*/;
assign _25681_ = _25672_ & _25680_ /*55324*/;
assign _25496_ = _25672_ ^ _25680_ /*55325*/;
assign _25678_ = _25679_ | _25681_ /*55322*/;
assign _25683_ = ~Q[35] /*55321*/;
assign _25682_ = _25683_ & D[24] /*55320*/;
assign _25685_ = _25049_ & _25682_ /*55315*/;
assign _25686_ = _25049_ ^ _25682_ /*55318*/;
assign _25687_ = _25678_ & _25686_ /*55316*/;
assign _25497_ = _25678_ ^ _25686_ /*55317*/;
assign _25684_ = _25685_ | _25687_ /*55314*/;
assign _25689_ = ~Q[35] /*55313*/;
assign _25688_ = _25689_ & D[25] /*55312*/;
assign _25691_ = _25050_ & _25688_ /*55307*/;
assign _25692_ = _25050_ ^ _25688_ /*55310*/;
assign _25693_ = _25684_ & _25692_ /*55308*/;
assign _25498_ = _25684_ ^ _25692_ /*55309*/;
assign _25690_ = _25691_ | _25693_ /*55306*/;
assign _25695_ = ~Q[35] /*55305*/;
assign _25694_ = _25695_ & D[26] /*55304*/;
assign _25697_ = _25051_ & _25694_ /*55299*/;
assign _25698_ = _25051_ ^ _25694_ /*55302*/;
assign _25699_ = _25690_ & _25698_ /*55300*/;
assign _25499_ = _25690_ ^ _25698_ /*55301*/;
assign _25696_ = _25697_ | _25699_ /*55298*/;
assign _25701_ = ~Q[35] /*55297*/;
assign _25700_ = _25701_ & D[27] /*55296*/;
assign _25703_ = _25052_ & _25700_ /*55291*/;
assign _25704_ = _25052_ ^ _25700_ /*55294*/;
assign _25705_ = _25696_ & _25704_ /*55292*/;
assign _25500_ = _25696_ ^ _25704_ /*55293*/;
assign _25702_ = _25703_ | _25705_ /*55290*/;
assign _25707_ = ~Q[35] /*55289*/;
assign _25706_ = _25707_ & D[28] /*55288*/;
assign _25709_ = _25053_ & _25706_ /*55283*/;
assign _25710_ = _25053_ ^ _25706_ /*55286*/;
assign _25711_ = _25702_ & _25710_ /*55284*/;
assign _25501_ = _25702_ ^ _25710_ /*55285*/;
assign _25708_ = _25709_ | _25711_ /*55282*/;
assign _25713_ = ~Q[35] /*55281*/;
assign _25712_ = _25713_ & D[29] /*55280*/;
assign _25715_ = _25054_ & _25712_ /*55275*/;
assign _25716_ = _25054_ ^ _25712_ /*55278*/;
assign _25717_ = _25708_ & _25716_ /*55276*/;
assign _25502_ = _25708_ ^ _25716_ /*55277*/;
assign _25714_ = _25715_ | _25717_ /*55274*/;
assign _25719_ = ~Q[35] /*55273*/;
assign _25718_ = _25719_ & D[30] /*55272*/;
assign _25721_ = _25055_ & _25718_ /*55267*/;
assign _25722_ = _25055_ ^ _25718_ /*55270*/;
assign _25723_ = _25714_ & _25722_ /*55268*/;
assign _25503_ = _25714_ ^ _25722_ /*55269*/;
assign _25720_ = _25721_ | _25723_ /*55266*/;
assign _25725_ = ~Q[35] /*55265*/;
assign _25724_ = _25725_ & D[31] /*55264*/;
assign _25727_ = _25056_ & _25724_ /*55259*/;
assign _25728_ = _25056_ ^ _25724_ /*55262*/;
assign _25729_ = _25720_ & _25728_ /*55260*/;
assign _25504_ = _25720_ ^ _25728_ /*55261*/;
assign _25726_ = _25727_ | _25729_ /*55258*/;
assign _25731_ = ~Q[35] /*55257*/;
assign _25730_ = _25731_ & D[32] /*55256*/;
assign _25733_ = _25057_ & _25730_ /*55251*/;
assign _25734_ = _25057_ ^ _25730_ /*55254*/;
assign _25735_ = _25726_ & _25734_ /*55252*/;
assign _25505_ = _25726_ ^ _25734_ /*55253*/;
assign _25732_ = _25733_ | _25735_ /*55250*/;
assign _25737_ = ~Q[35] /*55249*/;
assign _25736_ = _25737_ & D[33] /*55248*/;
assign _25739_ = _25058_ & _25736_ /*55243*/;
assign _25740_ = _25058_ ^ _25736_ /*55246*/;
assign _25741_ = _25732_ & _25740_ /*55244*/;
assign _25506_ = _25732_ ^ _25740_ /*55245*/;
assign _25738_ = _25739_ | _25741_ /*55242*/;
assign _25743_ = ~Q[35] /*55241*/;
assign _25742_ = _25743_ & D[34] /*55240*/;
assign _25745_ = _25059_ & _25742_ /*55235*/;
assign _25746_ = _25059_ ^ _25742_ /*55238*/;
assign _25747_ = _25738_ & _25746_ /*55236*/;
assign _25507_ = _25738_ ^ _25746_ /*55237*/;
assign _25744_ = _25745_ | _25747_ /*55234*/;
assign _25749_ = ~Q[35] /*55233*/;
assign _25748_ = _25749_ & D[35] /*55232*/;
assign _25751_ = _25060_ & _25748_ /*55227*/;
assign _25752_ = _25060_ ^ _25748_ /*55230*/;
assign _25753_ = _25744_ & _25752_ /*55228*/;
assign _25508_ = _25744_ ^ _25752_ /*55229*/;
assign _25750_ = _25751_ | _25753_ /*55226*/;
assign _25755_ = ~Q[35] /*55225*/;
assign _25754_ = _25755_ & D[36] /*55224*/;
assign _25757_ = _25061_ & _25754_ /*55219*/;
assign _25758_ = _25061_ ^ _25754_ /*55222*/;
assign _25759_ = _25750_ & _25758_ /*55220*/;
assign _25509_ = _25750_ ^ _25758_ /*55221*/;
assign _25756_ = _25757_ | _25759_ /*55218*/;
assign _25761_ = ~Q[35] /*55217*/;
assign _25760_ = _25761_ & D[37] /*55216*/;
assign _25763_ = _25062_ & _25760_ /*55211*/;
assign _25764_ = _25062_ ^ _25760_ /*55214*/;
assign _25765_ = _25756_ & _25764_ /*55212*/;
assign _25510_ = _25756_ ^ _25764_ /*55213*/;
assign _25762_ = _25763_ | _25765_ /*55210*/;
assign _25767_ = ~Q[35] /*55209*/;
assign _25766_ = _25767_ & D[38] /*55208*/;
assign _25769_ = _25063_ & _25766_ /*55203*/;
assign _25770_ = _25063_ ^ _25766_ /*55206*/;
assign _25771_ = _25762_ & _25770_ /*55204*/;
assign _25511_ = _25762_ ^ _25770_ /*55205*/;
assign _25768_ = _25769_ | _25771_ /*55202*/;
assign _25773_ = ~Q[35] /*55201*/;
assign _25772_ = _25773_ & D[39] /*55200*/;
assign _25775_ = _25064_ & _25772_ /*55195*/;
assign _25776_ = _25064_ ^ _25772_ /*55198*/;
assign _25777_ = _25768_ & _25776_ /*55196*/;
assign _25512_ = _25768_ ^ _25776_ /*55197*/;
assign _25774_ = _25775_ | _25777_ /*55194*/;
assign _25779_ = ~Q[35] /*55193*/;
assign _25778_ = _25779_ & D[40] /*55192*/;
assign _25781_ = _25065_ & _25778_ /*55187*/;
assign _25782_ = _25065_ ^ _25778_ /*55190*/;
assign _25783_ = _25774_ & _25782_ /*55188*/;
assign _25513_ = _25774_ ^ _25782_ /*55189*/;
assign _25780_ = _25781_ | _25783_ /*55186*/;
assign _25785_ = ~Q[35] /*55185*/;
assign _25784_ = _25785_ & D[41] /*55184*/;
assign _25787_ = _25066_ & _25784_ /*55179*/;
assign _25788_ = _25066_ ^ _25784_ /*55182*/;
assign _25789_ = _25780_ & _25788_ /*55180*/;
assign _25514_ = _25780_ ^ _25788_ /*55181*/;
assign _25786_ = _25787_ | _25789_ /*55178*/;
assign _25791_ = ~Q[35] /*55177*/;
assign _25790_ = _25791_ & D[42] /*55176*/;
assign _25793_ = _25067_ & _25790_ /*55171*/;
assign _25794_ = _25067_ ^ _25790_ /*55174*/;
assign _25795_ = _25786_ & _25794_ /*55172*/;
assign _25515_ = _25786_ ^ _25794_ /*55173*/;
assign _25792_ = _25793_ | _25795_ /*55170*/;
assign _25797_ = ~Q[35] /*55169*/;
assign _25796_ = _25797_ & D[43] /*55168*/;
assign _25799_ = _25068_ & _25796_ /*55163*/;
assign _25800_ = _25068_ ^ _25796_ /*55166*/;
assign _25801_ = _25792_ & _25800_ /*55164*/;
assign _25516_ = _25792_ ^ _25800_ /*55165*/;
assign _25798_ = _25799_ | _25801_ /*55162*/;
assign _25803_ = ~Q[35] /*55161*/;
assign _25802_ = _25803_ & D[44] /*55160*/;
assign _25805_ = _25069_ & _25802_ /*55155*/;
assign _25806_ = _25069_ ^ _25802_ /*55158*/;
assign _25807_ = _25798_ & _25806_ /*55156*/;
assign _25517_ = _25798_ ^ _25806_ /*55157*/;
assign _25804_ = _25805_ | _25807_ /*55154*/;
assign _25809_ = ~Q[35] /*55153*/;
assign _25808_ = _25809_ & D[45] /*55152*/;
assign _25811_ = _25070_ & _25808_ /*55147*/;
assign _25812_ = _25070_ ^ _25808_ /*55150*/;
assign _25813_ = _25804_ & _25812_ /*55148*/;
assign _25518_ = _25804_ ^ _25812_ /*55149*/;
assign _25810_ = _25811_ | _25813_ /*55146*/;
assign _25815_ = ~Q[35] /*55145*/;
assign _25814_ = _25815_ & D[46] /*55144*/;
assign _25817_ = _25071_ & _25814_ /*55139*/;
assign _25818_ = _25071_ ^ _25814_ /*55142*/;
assign _25819_ = _25810_ & _25818_ /*55140*/;
assign _25519_ = _25810_ ^ _25818_ /*55141*/;
assign _25816_ = _25817_ | _25819_ /*55138*/;
assign _25821_ = ~Q[35] /*55137*/;
assign _25820_ = _25821_ & D[47] /*55136*/;
assign _25823_ = _25072_ & _25820_ /*55131*/;
assign _25824_ = _25072_ ^ _25820_ /*55134*/;
assign _25825_ = _25816_ & _25824_ /*55132*/;
assign _25520_ = _25816_ ^ _25824_ /*55133*/;
assign _25822_ = _25823_ | _25825_ /*55130*/;
assign _25827_ = ~Q[35] /*55129*/;
assign _25826_ = _25827_ & D[48] /*55128*/;
assign _25829_ = _25073_ & _25826_ /*55123*/;
assign _25830_ = _25073_ ^ _25826_ /*55126*/;
assign _25831_ = _25822_ & _25830_ /*55124*/;
assign _25521_ = _25822_ ^ _25830_ /*55125*/;
assign _25828_ = _25829_ | _25831_ /*55122*/;
assign _25833_ = ~Q[35] /*55121*/;
assign _25832_ = _25833_ & D[49] /*55120*/;
assign _25835_ = _25074_ & _25832_ /*55115*/;
assign _25836_ = _25074_ ^ _25832_ /*55118*/;
assign _25837_ = _25828_ & _25836_ /*55116*/;
assign _25522_ = _25828_ ^ _25836_ /*55117*/;
assign _25834_ = _25835_ | _25837_ /*55114*/;
assign _25839_ = ~Q[35] /*55113*/;
assign _25838_ = _25839_ & D[50] /*55112*/;
assign _25841_ = _25075_ & _25838_ /*55107*/;
assign _25842_ = _25075_ ^ _25838_ /*55110*/;
assign _25843_ = _25834_ & _25842_ /*55108*/;
assign _25523_ = _25834_ ^ _25842_ /*55109*/;
assign _25840_ = _25841_ | _25843_ /*55106*/;
assign _25845_ = ~Q[35] /*55105*/;
assign _25844_ = _25845_ & D[51] /*55104*/;
assign _25847_ = _25076_ & _25844_ /*55099*/;
assign _25848_ = _25076_ ^ _25844_ /*55102*/;
assign _25849_ = _25840_ & _25848_ /*55100*/;
assign _25524_ = _25840_ ^ _25848_ /*55101*/;
assign _25846_ = _25847_ | _25849_ /*55098*/;
assign _25851_ = ~Q[35] /*55097*/;
assign _25850_ = _25851_ & D[52] /*55096*/;
assign _25853_ = _25077_ & _25850_ /*55091*/;
assign _25854_ = _25077_ ^ _25850_ /*55094*/;
assign _25855_ = _25846_ & _25854_ /*55092*/;
assign _25525_ = _25846_ ^ _25854_ /*55093*/;
assign _25852_ = _25853_ | _25855_ /*55090*/;
assign _25857_ = ~Q[35] /*55089*/;
assign _25856_ = _25857_ & D[53] /*55088*/;
assign _25859_ = _25078_ & _25856_ /*55083*/;
assign _25860_ = _25078_ ^ _25856_ /*55086*/;
assign _25861_ = _25852_ & _25860_ /*55084*/;
assign _25526_ = _25852_ ^ _25860_ /*55085*/;
assign _25858_ = _25859_ | _25861_ /*55082*/;
assign _25863_ = ~Q[35] /*55081*/;
assign _25862_ = _25863_ & D[54] /*55080*/;
assign _25865_ = _25079_ & _25862_ /*55075*/;
assign _25866_ = _25079_ ^ _25862_ /*55078*/;
assign _25867_ = _25858_ & _25866_ /*55076*/;
assign _25527_ = _25858_ ^ _25866_ /*55077*/;
assign _25864_ = _25865_ | _25867_ /*55074*/;
assign _25869_ = ~Q[35] /*55073*/;
assign _25868_ = _25869_ & D[55] /*55072*/;
assign _25871_ = _25080_ & _25868_ /*55067*/;
assign _25872_ = _25080_ ^ _25868_ /*55070*/;
assign _25873_ = _25864_ & _25872_ /*55068*/;
assign _25528_ = _25864_ ^ _25872_ /*55069*/;
assign _25870_ = _25871_ | _25873_ /*55066*/;
assign _25875_ = ~Q[35] /*55065*/;
assign _25874_ = _25875_ & D[56] /*55064*/;
assign _25877_ = _25081_ & _25874_ /*55059*/;
assign _25878_ = _25081_ ^ _25874_ /*55062*/;
assign _25879_ = _25870_ & _25878_ /*55060*/;
assign _25529_ = _25870_ ^ _25878_ /*55061*/;
assign _25876_ = _25877_ | _25879_ /*55058*/;
assign _25881_ = ~Q[35] /*55057*/;
assign _25880_ = _25881_ & D[57] /*55056*/;
assign _25883_ = _25082_ & _25880_ /*55051*/;
assign _25884_ = _25082_ ^ _25880_ /*55054*/;
assign _25885_ = _25876_ & _25884_ /*55052*/;
assign _25530_ = _25876_ ^ _25884_ /*55053*/;
assign _25882_ = _25883_ | _25885_ /*55050*/;
assign _25887_ = ~Q[35] /*55049*/;
assign _25886_ = _25887_ & D[58] /*55048*/;
assign _25889_ = _25083_ & _25886_ /*55043*/;
assign _25890_ = _25083_ ^ _25886_ /*55046*/;
assign _25891_ = _25882_ & _25890_ /*55044*/;
assign _25531_ = _25882_ ^ _25890_ /*55045*/;
assign _25888_ = _25889_ | _25891_ /*55042*/;
assign _25893_ = ~Q[35] /*55041*/;
assign _25892_ = _25893_ & D[59] /*55040*/;
assign _25895_ = _25084_ & _25892_ /*55035*/;
assign _25896_ = _25084_ ^ _25892_ /*55038*/;
assign _25897_ = _25888_ & _25896_ /*55036*/;
assign _25532_ = _25888_ ^ _25896_ /*55037*/;
assign _25894_ = _25895_ | _25897_ /*55034*/;
assign _25899_ = ~Q[35] /*55033*/;
assign _25898_ = _25899_ & D[60] /*55032*/;
assign _25901_ = _25085_ & _25898_ /*55027*/;
assign _25902_ = _25085_ ^ _25898_ /*55030*/;
assign _25903_ = _25894_ & _25902_ /*55028*/;
assign _25533_ = _25894_ ^ _25902_ /*55029*/;
assign _25900_ = _25901_ | _25903_ /*55026*/;
assign _25905_ = ~Q[35] /*55025*/;
assign _25904_ = _25905_ & D[61] /*55024*/;
assign _25907_ = _25086_ & _25904_ /*55019*/;
assign _25908_ = _25086_ ^ _25904_ /*55022*/;
assign _25909_ = _25900_ & _25908_ /*55020*/;
assign _25534_ = _25900_ ^ _25908_ /*55021*/;
assign _25906_ = _25907_ | _25909_ /*55018*/;
assign _25911_ = ~Q[35] /*55017*/;
assign _25910_ = _25911_ & D[62] /*55016*/;
assign _25913_ = _25087_ & _25910_ /*55011*/;
assign _25914_ = _25087_ ^ _25910_ /*55014*/;
assign _25915_ = _25906_ & _25914_ /*55012*/;
assign _25535_ = _25906_ ^ _25914_ /*55013*/;
assign _25912_ = _25913_ | _25915_ /*55010*/;
assign _25917_ = ~Q[35] /*55009*/;
assign _25916_ = _25917_ & zeroWire /*55008*/;
assign _25918_ = _25088_ ^ _25916_ /*55006*/;
assign _25536_ = _25918_ ^ _25912_ /*55005*/;
assign _25989_ = ~D[0] /*54751*/;
assign _25986_ = R_0[34] & _25989_ /*54747*/;
assign _25987_ = R_0[34] ^ _25989_ /*54750*/;
assign _25988_ = oneWire & _25987_ /*54748*/;
assign _25921_ = oneWire ^ _25987_ /*54749*/;
assign _25985_ = _25986_ | _25988_ /*54746*/;
assign _25994_ = ~D[1] /*54745*/;
assign _25991_ = _25473_ & _25994_ /*54741*/;
assign _25992_ = _25473_ ^ _25994_ /*54744*/;
assign _25993_ = _25985_ & _25992_ /*54742*/;
assign _25922_ = _25985_ ^ _25992_ /*54743*/;
assign _25990_ = _25991_ | _25993_ /*54740*/;
assign _25999_ = ~D[2] /*54739*/;
assign _25996_ = _25474_ & _25999_ /*54735*/;
assign _25997_ = _25474_ ^ _25999_ /*54738*/;
assign _25998_ = _25990_ & _25997_ /*54736*/;
assign _25923_ = _25990_ ^ _25997_ /*54737*/;
assign _25995_ = _25996_ | _25998_ /*54734*/;
assign _26004_ = ~D[3] /*54733*/;
assign _26001_ = _25475_ & _26004_ /*54729*/;
assign _26002_ = _25475_ ^ _26004_ /*54732*/;
assign _26003_ = _25995_ & _26002_ /*54730*/;
assign _25924_ = _25995_ ^ _26002_ /*54731*/;
assign _26000_ = _26001_ | _26003_ /*54728*/;
assign _26009_ = ~D[4] /*54727*/;
assign _26006_ = _25476_ & _26009_ /*54723*/;
assign _26007_ = _25476_ ^ _26009_ /*54726*/;
assign _26008_ = _26000_ & _26007_ /*54724*/;
assign _25925_ = _26000_ ^ _26007_ /*54725*/;
assign _26005_ = _26006_ | _26008_ /*54722*/;
assign _26014_ = ~D[5] /*54721*/;
assign _26011_ = _25477_ & _26014_ /*54717*/;
assign _26012_ = _25477_ ^ _26014_ /*54720*/;
assign _26013_ = _26005_ & _26012_ /*54718*/;
assign _25926_ = _26005_ ^ _26012_ /*54719*/;
assign _26010_ = _26011_ | _26013_ /*54716*/;
assign _26019_ = ~D[6] /*54715*/;
assign _26016_ = _25478_ & _26019_ /*54711*/;
assign _26017_ = _25478_ ^ _26019_ /*54714*/;
assign _26018_ = _26010_ & _26017_ /*54712*/;
assign _25927_ = _26010_ ^ _26017_ /*54713*/;
assign _26015_ = _26016_ | _26018_ /*54710*/;
assign _26024_ = ~D[7] /*54709*/;
assign _26021_ = _25479_ & _26024_ /*54705*/;
assign _26022_ = _25479_ ^ _26024_ /*54708*/;
assign _26023_ = _26015_ & _26022_ /*54706*/;
assign _25928_ = _26015_ ^ _26022_ /*54707*/;
assign _26020_ = _26021_ | _26023_ /*54704*/;
assign _26029_ = ~D[8] /*54703*/;
assign _26026_ = _25480_ & _26029_ /*54699*/;
assign _26027_ = _25480_ ^ _26029_ /*54702*/;
assign _26028_ = _26020_ & _26027_ /*54700*/;
assign _25929_ = _26020_ ^ _26027_ /*54701*/;
assign _26025_ = _26026_ | _26028_ /*54698*/;
assign _26034_ = ~D[9] /*54697*/;
assign _26031_ = _25481_ & _26034_ /*54693*/;
assign _26032_ = _25481_ ^ _26034_ /*54696*/;
assign _26033_ = _26025_ & _26032_ /*54694*/;
assign _25930_ = _26025_ ^ _26032_ /*54695*/;
assign _26030_ = _26031_ | _26033_ /*54692*/;
assign _26039_ = ~D[10] /*54691*/;
assign _26036_ = _25482_ & _26039_ /*54687*/;
assign _26037_ = _25482_ ^ _26039_ /*54690*/;
assign _26038_ = _26030_ & _26037_ /*54688*/;
assign _25931_ = _26030_ ^ _26037_ /*54689*/;
assign _26035_ = _26036_ | _26038_ /*54686*/;
assign _26044_ = ~D[11] /*54685*/;
assign _26041_ = _25483_ & _26044_ /*54681*/;
assign _26042_ = _25483_ ^ _26044_ /*54684*/;
assign _26043_ = _26035_ & _26042_ /*54682*/;
assign _25932_ = _26035_ ^ _26042_ /*54683*/;
assign _26040_ = _26041_ | _26043_ /*54680*/;
assign _26049_ = ~D[12] /*54679*/;
assign _26046_ = _25484_ & _26049_ /*54675*/;
assign _26047_ = _25484_ ^ _26049_ /*54678*/;
assign _26048_ = _26040_ & _26047_ /*54676*/;
assign _25933_ = _26040_ ^ _26047_ /*54677*/;
assign _26045_ = _26046_ | _26048_ /*54674*/;
assign _26054_ = ~D[13] /*54673*/;
assign _26051_ = _25485_ & _26054_ /*54669*/;
assign _26052_ = _25485_ ^ _26054_ /*54672*/;
assign _26053_ = _26045_ & _26052_ /*54670*/;
assign _25934_ = _26045_ ^ _26052_ /*54671*/;
assign _26050_ = _26051_ | _26053_ /*54668*/;
assign _26059_ = ~D[14] /*54667*/;
assign _26056_ = _25486_ & _26059_ /*54663*/;
assign _26057_ = _25486_ ^ _26059_ /*54666*/;
assign _26058_ = _26050_ & _26057_ /*54664*/;
assign _25935_ = _26050_ ^ _26057_ /*54665*/;
assign _26055_ = _26056_ | _26058_ /*54662*/;
assign _26064_ = ~D[15] /*54661*/;
assign _26061_ = _25487_ & _26064_ /*54657*/;
assign _26062_ = _25487_ ^ _26064_ /*54660*/;
assign _26063_ = _26055_ & _26062_ /*54658*/;
assign _25936_ = _26055_ ^ _26062_ /*54659*/;
assign _26060_ = _26061_ | _26063_ /*54656*/;
assign _26069_ = ~D[16] /*54655*/;
assign _26066_ = _25488_ & _26069_ /*54651*/;
assign _26067_ = _25488_ ^ _26069_ /*54654*/;
assign _26068_ = _26060_ & _26067_ /*54652*/;
assign _25937_ = _26060_ ^ _26067_ /*54653*/;
assign _26065_ = _26066_ | _26068_ /*54650*/;
assign _26074_ = ~D[17] /*54649*/;
assign _26071_ = _25489_ & _26074_ /*54645*/;
assign _26072_ = _25489_ ^ _26074_ /*54648*/;
assign _26073_ = _26065_ & _26072_ /*54646*/;
assign _25938_ = _26065_ ^ _26072_ /*54647*/;
assign _26070_ = _26071_ | _26073_ /*54644*/;
assign _26079_ = ~D[18] /*54643*/;
assign _26076_ = _25490_ & _26079_ /*54639*/;
assign _26077_ = _25490_ ^ _26079_ /*54642*/;
assign _26078_ = _26070_ & _26077_ /*54640*/;
assign _25939_ = _26070_ ^ _26077_ /*54641*/;
assign _26075_ = _26076_ | _26078_ /*54638*/;
assign _26084_ = ~D[19] /*54637*/;
assign _26081_ = _25491_ & _26084_ /*54633*/;
assign _26082_ = _25491_ ^ _26084_ /*54636*/;
assign _26083_ = _26075_ & _26082_ /*54634*/;
assign _25940_ = _26075_ ^ _26082_ /*54635*/;
assign _26080_ = _26081_ | _26083_ /*54632*/;
assign _26089_ = ~D[20] /*54631*/;
assign _26086_ = _25492_ & _26089_ /*54627*/;
assign _26087_ = _25492_ ^ _26089_ /*54630*/;
assign _26088_ = _26080_ & _26087_ /*54628*/;
assign _25941_ = _26080_ ^ _26087_ /*54629*/;
assign _26085_ = _26086_ | _26088_ /*54626*/;
assign _26094_ = ~D[21] /*54625*/;
assign _26091_ = _25493_ & _26094_ /*54621*/;
assign _26092_ = _25493_ ^ _26094_ /*54624*/;
assign _26093_ = _26085_ & _26092_ /*54622*/;
assign _25942_ = _26085_ ^ _26092_ /*54623*/;
assign _26090_ = _26091_ | _26093_ /*54620*/;
assign _26099_ = ~D[22] /*54619*/;
assign _26096_ = _25494_ & _26099_ /*54615*/;
assign _26097_ = _25494_ ^ _26099_ /*54618*/;
assign _26098_ = _26090_ & _26097_ /*54616*/;
assign _25943_ = _26090_ ^ _26097_ /*54617*/;
assign _26095_ = _26096_ | _26098_ /*54614*/;
assign _26104_ = ~D[23] /*54613*/;
assign _26101_ = _25495_ & _26104_ /*54609*/;
assign _26102_ = _25495_ ^ _26104_ /*54612*/;
assign _26103_ = _26095_ & _26102_ /*54610*/;
assign _25944_ = _26095_ ^ _26102_ /*54611*/;
assign _26100_ = _26101_ | _26103_ /*54608*/;
assign _26109_ = ~D[24] /*54607*/;
assign _26106_ = _25496_ & _26109_ /*54603*/;
assign _26107_ = _25496_ ^ _26109_ /*54606*/;
assign _26108_ = _26100_ & _26107_ /*54604*/;
assign _25945_ = _26100_ ^ _26107_ /*54605*/;
assign _26105_ = _26106_ | _26108_ /*54602*/;
assign _26114_ = ~D[25] /*54601*/;
assign _26111_ = _25497_ & _26114_ /*54597*/;
assign _26112_ = _25497_ ^ _26114_ /*54600*/;
assign _26113_ = _26105_ & _26112_ /*54598*/;
assign _25946_ = _26105_ ^ _26112_ /*54599*/;
assign _26110_ = _26111_ | _26113_ /*54596*/;
assign _26119_ = ~D[26] /*54595*/;
assign _26116_ = _25498_ & _26119_ /*54591*/;
assign _26117_ = _25498_ ^ _26119_ /*54594*/;
assign _26118_ = _26110_ & _26117_ /*54592*/;
assign _25947_ = _26110_ ^ _26117_ /*54593*/;
assign _26115_ = _26116_ | _26118_ /*54590*/;
assign _26124_ = ~D[27] /*54589*/;
assign _26121_ = _25499_ & _26124_ /*54585*/;
assign _26122_ = _25499_ ^ _26124_ /*54588*/;
assign _26123_ = _26115_ & _26122_ /*54586*/;
assign _25948_ = _26115_ ^ _26122_ /*54587*/;
assign _26120_ = _26121_ | _26123_ /*54584*/;
assign _26129_ = ~D[28] /*54583*/;
assign _26126_ = _25500_ & _26129_ /*54579*/;
assign _26127_ = _25500_ ^ _26129_ /*54582*/;
assign _26128_ = _26120_ & _26127_ /*54580*/;
assign _25949_ = _26120_ ^ _26127_ /*54581*/;
assign _26125_ = _26126_ | _26128_ /*54578*/;
assign _26134_ = ~D[29] /*54577*/;
assign _26131_ = _25501_ & _26134_ /*54573*/;
assign _26132_ = _25501_ ^ _26134_ /*54576*/;
assign _26133_ = _26125_ & _26132_ /*54574*/;
assign _25950_ = _26125_ ^ _26132_ /*54575*/;
assign _26130_ = _26131_ | _26133_ /*54572*/;
assign _26139_ = ~D[30] /*54571*/;
assign _26136_ = _25502_ & _26139_ /*54567*/;
assign _26137_ = _25502_ ^ _26139_ /*54570*/;
assign _26138_ = _26130_ & _26137_ /*54568*/;
assign _25951_ = _26130_ ^ _26137_ /*54569*/;
assign _26135_ = _26136_ | _26138_ /*54566*/;
assign _26144_ = ~D[31] /*54565*/;
assign _26141_ = _25503_ & _26144_ /*54561*/;
assign _26142_ = _25503_ ^ _26144_ /*54564*/;
assign _26143_ = _26135_ & _26142_ /*54562*/;
assign _25952_ = _26135_ ^ _26142_ /*54563*/;
assign _26140_ = _26141_ | _26143_ /*54560*/;
assign _26149_ = ~D[32] /*54559*/;
assign _26146_ = _25504_ & _26149_ /*54555*/;
assign _26147_ = _25504_ ^ _26149_ /*54558*/;
assign _26148_ = _26140_ & _26147_ /*54556*/;
assign _25953_ = _26140_ ^ _26147_ /*54557*/;
assign _26145_ = _26146_ | _26148_ /*54554*/;
assign _26154_ = ~D[33] /*54553*/;
assign _26151_ = _25505_ & _26154_ /*54549*/;
assign _26152_ = _25505_ ^ _26154_ /*54552*/;
assign _26153_ = _26145_ & _26152_ /*54550*/;
assign _25954_ = _26145_ ^ _26152_ /*54551*/;
assign _26150_ = _26151_ | _26153_ /*54548*/;
assign _26159_ = ~D[34] /*54547*/;
assign _26156_ = _25506_ & _26159_ /*54543*/;
assign _26157_ = _25506_ ^ _26159_ /*54546*/;
assign _26158_ = _26150_ & _26157_ /*54544*/;
assign _25955_ = _26150_ ^ _26157_ /*54545*/;
assign _26155_ = _26156_ | _26158_ /*54542*/;
assign _26164_ = ~D[35] /*54541*/;
assign _26161_ = _25507_ & _26164_ /*54537*/;
assign _26162_ = _25507_ ^ _26164_ /*54540*/;
assign _26163_ = _26155_ & _26162_ /*54538*/;
assign _25956_ = _26155_ ^ _26162_ /*54539*/;
assign _26160_ = _26161_ | _26163_ /*54536*/;
assign _26169_ = ~D[36] /*54535*/;
assign _26166_ = _25508_ & _26169_ /*54531*/;
assign _26167_ = _25508_ ^ _26169_ /*54534*/;
assign _26168_ = _26160_ & _26167_ /*54532*/;
assign _25957_ = _26160_ ^ _26167_ /*54533*/;
assign _26165_ = _26166_ | _26168_ /*54530*/;
assign _26174_ = ~D[37] /*54529*/;
assign _26171_ = _25509_ & _26174_ /*54525*/;
assign _26172_ = _25509_ ^ _26174_ /*54528*/;
assign _26173_ = _26165_ & _26172_ /*54526*/;
assign _25958_ = _26165_ ^ _26172_ /*54527*/;
assign _26170_ = _26171_ | _26173_ /*54524*/;
assign _26179_ = ~D[38] /*54523*/;
assign _26176_ = _25510_ & _26179_ /*54519*/;
assign _26177_ = _25510_ ^ _26179_ /*54522*/;
assign _26178_ = _26170_ & _26177_ /*54520*/;
assign _25959_ = _26170_ ^ _26177_ /*54521*/;
assign _26175_ = _26176_ | _26178_ /*54518*/;
assign _26184_ = ~D[39] /*54517*/;
assign _26181_ = _25511_ & _26184_ /*54513*/;
assign _26182_ = _25511_ ^ _26184_ /*54516*/;
assign _26183_ = _26175_ & _26182_ /*54514*/;
assign _25960_ = _26175_ ^ _26182_ /*54515*/;
assign _26180_ = _26181_ | _26183_ /*54512*/;
assign _26189_ = ~D[40] /*54511*/;
assign _26186_ = _25512_ & _26189_ /*54507*/;
assign _26187_ = _25512_ ^ _26189_ /*54510*/;
assign _26188_ = _26180_ & _26187_ /*54508*/;
assign _25961_ = _26180_ ^ _26187_ /*54509*/;
assign _26185_ = _26186_ | _26188_ /*54506*/;
assign _26194_ = ~D[41] /*54505*/;
assign _26191_ = _25513_ & _26194_ /*54501*/;
assign _26192_ = _25513_ ^ _26194_ /*54504*/;
assign _26193_ = _26185_ & _26192_ /*54502*/;
assign _25962_ = _26185_ ^ _26192_ /*54503*/;
assign _26190_ = _26191_ | _26193_ /*54500*/;
assign _26199_ = ~D[42] /*54499*/;
assign _26196_ = _25514_ & _26199_ /*54495*/;
assign _26197_ = _25514_ ^ _26199_ /*54498*/;
assign _26198_ = _26190_ & _26197_ /*54496*/;
assign _25963_ = _26190_ ^ _26197_ /*54497*/;
assign _26195_ = _26196_ | _26198_ /*54494*/;
assign _26204_ = ~D[43] /*54493*/;
assign _26201_ = _25515_ & _26204_ /*54489*/;
assign _26202_ = _25515_ ^ _26204_ /*54492*/;
assign _26203_ = _26195_ & _26202_ /*54490*/;
assign _25964_ = _26195_ ^ _26202_ /*54491*/;
assign _26200_ = _26201_ | _26203_ /*54488*/;
assign _26209_ = ~D[44] /*54487*/;
assign _26206_ = _25516_ & _26209_ /*54483*/;
assign _26207_ = _25516_ ^ _26209_ /*54486*/;
assign _26208_ = _26200_ & _26207_ /*54484*/;
assign _25965_ = _26200_ ^ _26207_ /*54485*/;
assign _26205_ = _26206_ | _26208_ /*54482*/;
assign _26214_ = ~D[45] /*54481*/;
assign _26211_ = _25517_ & _26214_ /*54477*/;
assign _26212_ = _25517_ ^ _26214_ /*54480*/;
assign _26213_ = _26205_ & _26212_ /*54478*/;
assign _25966_ = _26205_ ^ _26212_ /*54479*/;
assign _26210_ = _26211_ | _26213_ /*54476*/;
assign _26219_ = ~D[46] /*54475*/;
assign _26216_ = _25518_ & _26219_ /*54471*/;
assign _26217_ = _25518_ ^ _26219_ /*54474*/;
assign _26218_ = _26210_ & _26217_ /*54472*/;
assign _25967_ = _26210_ ^ _26217_ /*54473*/;
assign _26215_ = _26216_ | _26218_ /*54470*/;
assign _26224_ = ~D[47] /*54469*/;
assign _26221_ = _25519_ & _26224_ /*54465*/;
assign _26222_ = _25519_ ^ _26224_ /*54468*/;
assign _26223_ = _26215_ & _26222_ /*54466*/;
assign _25968_ = _26215_ ^ _26222_ /*54467*/;
assign _26220_ = _26221_ | _26223_ /*54464*/;
assign _26229_ = ~D[48] /*54463*/;
assign _26226_ = _25520_ & _26229_ /*54459*/;
assign _26227_ = _25520_ ^ _26229_ /*54462*/;
assign _26228_ = _26220_ & _26227_ /*54460*/;
assign _25969_ = _26220_ ^ _26227_ /*54461*/;
assign _26225_ = _26226_ | _26228_ /*54458*/;
assign _26234_ = ~D[49] /*54457*/;
assign _26231_ = _25521_ & _26234_ /*54453*/;
assign _26232_ = _25521_ ^ _26234_ /*54456*/;
assign _26233_ = _26225_ & _26232_ /*54454*/;
assign _25970_ = _26225_ ^ _26232_ /*54455*/;
assign _26230_ = _26231_ | _26233_ /*54452*/;
assign _26239_ = ~D[50] /*54451*/;
assign _26236_ = _25522_ & _26239_ /*54447*/;
assign _26237_ = _25522_ ^ _26239_ /*54450*/;
assign _26238_ = _26230_ & _26237_ /*54448*/;
assign _25971_ = _26230_ ^ _26237_ /*54449*/;
assign _26235_ = _26236_ | _26238_ /*54446*/;
assign _26244_ = ~D[51] /*54445*/;
assign _26241_ = _25523_ & _26244_ /*54441*/;
assign _26242_ = _25523_ ^ _26244_ /*54444*/;
assign _26243_ = _26235_ & _26242_ /*54442*/;
assign _25972_ = _26235_ ^ _26242_ /*54443*/;
assign _26240_ = _26241_ | _26243_ /*54440*/;
assign _26249_ = ~D[52] /*54439*/;
assign _26246_ = _25524_ & _26249_ /*54435*/;
assign _26247_ = _25524_ ^ _26249_ /*54438*/;
assign _26248_ = _26240_ & _26247_ /*54436*/;
assign _25973_ = _26240_ ^ _26247_ /*54437*/;
assign _26245_ = _26246_ | _26248_ /*54434*/;
assign _26254_ = ~D[53] /*54433*/;
assign _26251_ = _25525_ & _26254_ /*54429*/;
assign _26252_ = _25525_ ^ _26254_ /*54432*/;
assign _26253_ = _26245_ & _26252_ /*54430*/;
assign _25974_ = _26245_ ^ _26252_ /*54431*/;
assign _26250_ = _26251_ | _26253_ /*54428*/;
assign _26259_ = ~D[54] /*54427*/;
assign _26256_ = _25526_ & _26259_ /*54423*/;
assign _26257_ = _25526_ ^ _26259_ /*54426*/;
assign _26258_ = _26250_ & _26257_ /*54424*/;
assign _25975_ = _26250_ ^ _26257_ /*54425*/;
assign _26255_ = _26256_ | _26258_ /*54422*/;
assign _26264_ = ~D[55] /*54421*/;
assign _26261_ = _25527_ & _26264_ /*54417*/;
assign _26262_ = _25527_ ^ _26264_ /*54420*/;
assign _26263_ = _26255_ & _26262_ /*54418*/;
assign _25976_ = _26255_ ^ _26262_ /*54419*/;
assign _26260_ = _26261_ | _26263_ /*54416*/;
assign _26269_ = ~D[56] /*54415*/;
assign _26266_ = _25528_ & _26269_ /*54411*/;
assign _26267_ = _25528_ ^ _26269_ /*54414*/;
assign _26268_ = _26260_ & _26267_ /*54412*/;
assign _25977_ = _26260_ ^ _26267_ /*54413*/;
assign _26265_ = _26266_ | _26268_ /*54410*/;
assign _26274_ = ~D[57] /*54409*/;
assign _26271_ = _25529_ & _26274_ /*54405*/;
assign _26272_ = _25529_ ^ _26274_ /*54408*/;
assign _26273_ = _26265_ & _26272_ /*54406*/;
assign _25978_ = _26265_ ^ _26272_ /*54407*/;
assign _26270_ = _26271_ | _26273_ /*54404*/;
assign _26279_ = ~D[58] /*54403*/;
assign _26276_ = _25530_ & _26279_ /*54399*/;
assign _26277_ = _25530_ ^ _26279_ /*54402*/;
assign _26278_ = _26270_ & _26277_ /*54400*/;
assign _25979_ = _26270_ ^ _26277_ /*54401*/;
assign _26275_ = _26276_ | _26278_ /*54398*/;
assign _26284_ = ~D[59] /*54397*/;
assign _26281_ = _25531_ & _26284_ /*54393*/;
assign _26282_ = _25531_ ^ _26284_ /*54396*/;
assign _26283_ = _26275_ & _26282_ /*54394*/;
assign _25980_ = _26275_ ^ _26282_ /*54395*/;
assign _26280_ = _26281_ | _26283_ /*54392*/;
assign _26289_ = ~D[60] /*54391*/;
assign _26286_ = _25532_ & _26289_ /*54387*/;
assign _26287_ = _25532_ ^ _26289_ /*54390*/;
assign _26288_ = _26280_ & _26287_ /*54388*/;
assign _25981_ = _26280_ ^ _26287_ /*54389*/;
assign _26285_ = _26286_ | _26288_ /*54386*/;
assign _26294_ = ~D[61] /*54385*/;
assign _26291_ = _25533_ & _26294_ /*54381*/;
assign _26292_ = _25533_ ^ _26294_ /*54384*/;
assign _26293_ = _26285_ & _26292_ /*54382*/;
assign _25982_ = _26285_ ^ _26292_ /*54383*/;
assign _26290_ = _26291_ | _26293_ /*54380*/;
assign _26299_ = ~D[62] /*54379*/;
assign _26296_ = _25534_ & _26299_ /*54375*/;
assign _26297_ = _25534_ ^ _26299_ /*54378*/;
assign _26298_ = _26290_ & _26297_ /*54376*/;
assign _25983_ = _26290_ ^ _26297_ /*54377*/;
assign _26295_ = _26296_ | _26298_ /*54374*/;
assign _26300_ = _25535_ & oneWire /*54369*/;
assign _26301_ = _25535_ ^ oneWire /*54372*/;
assign _26302_ = _26295_ & _26301_ /*54370*/;
assign _25984_ = _26295_ ^ _26301_ /*54371*/;
assign Q[34] = _26300_ | _26302_ /*54368*/;
assign _26435_ = ~Q[34] /*53983*/;
assign _26434_ = _26435_ & D[0] /*53982*/;
assign _26437_ = _25921_ & _26434_ /*53977*/;
assign _26438_ = _25921_ ^ _26434_ /*53980*/;
assign _26439_ = zeroWire & _26438_ /*53978*/;
assign _26369_ = zeroWire ^ _26438_ /*53979*/;
assign _26436_ = _26437_ | _26439_ /*53976*/;
assign _26441_ = ~Q[34] /*53975*/;
assign _26440_ = _26441_ & D[1] /*53974*/;
assign _26443_ = _25922_ & _26440_ /*53969*/;
assign _26444_ = _25922_ ^ _26440_ /*53972*/;
assign _26445_ = _26436_ & _26444_ /*53970*/;
assign _26370_ = _26436_ ^ _26444_ /*53971*/;
assign _26442_ = _26443_ | _26445_ /*53968*/;
assign _26447_ = ~Q[34] /*53967*/;
assign _26446_ = _26447_ & D[2] /*53966*/;
assign _26449_ = _25923_ & _26446_ /*53961*/;
assign _26450_ = _25923_ ^ _26446_ /*53964*/;
assign _26451_ = _26442_ & _26450_ /*53962*/;
assign _26371_ = _26442_ ^ _26450_ /*53963*/;
assign _26448_ = _26449_ | _26451_ /*53960*/;
assign _26453_ = ~Q[34] /*53959*/;
assign _26452_ = _26453_ & D[3] /*53958*/;
assign _26455_ = _25924_ & _26452_ /*53953*/;
assign _26456_ = _25924_ ^ _26452_ /*53956*/;
assign _26457_ = _26448_ & _26456_ /*53954*/;
assign _26372_ = _26448_ ^ _26456_ /*53955*/;
assign _26454_ = _26455_ | _26457_ /*53952*/;
assign _26459_ = ~Q[34] /*53951*/;
assign _26458_ = _26459_ & D[4] /*53950*/;
assign _26461_ = _25925_ & _26458_ /*53945*/;
assign _26462_ = _25925_ ^ _26458_ /*53948*/;
assign _26463_ = _26454_ & _26462_ /*53946*/;
assign _26373_ = _26454_ ^ _26462_ /*53947*/;
assign _26460_ = _26461_ | _26463_ /*53944*/;
assign _26465_ = ~Q[34] /*53943*/;
assign _26464_ = _26465_ & D[5] /*53942*/;
assign _26467_ = _25926_ & _26464_ /*53937*/;
assign _26468_ = _25926_ ^ _26464_ /*53940*/;
assign _26469_ = _26460_ & _26468_ /*53938*/;
assign _26374_ = _26460_ ^ _26468_ /*53939*/;
assign _26466_ = _26467_ | _26469_ /*53936*/;
assign _26471_ = ~Q[34] /*53935*/;
assign _26470_ = _26471_ & D[6] /*53934*/;
assign _26473_ = _25927_ & _26470_ /*53929*/;
assign _26474_ = _25927_ ^ _26470_ /*53932*/;
assign _26475_ = _26466_ & _26474_ /*53930*/;
assign _26375_ = _26466_ ^ _26474_ /*53931*/;
assign _26472_ = _26473_ | _26475_ /*53928*/;
assign _26477_ = ~Q[34] /*53927*/;
assign _26476_ = _26477_ & D[7] /*53926*/;
assign _26479_ = _25928_ & _26476_ /*53921*/;
assign _26480_ = _25928_ ^ _26476_ /*53924*/;
assign _26481_ = _26472_ & _26480_ /*53922*/;
assign _26376_ = _26472_ ^ _26480_ /*53923*/;
assign _26478_ = _26479_ | _26481_ /*53920*/;
assign _26483_ = ~Q[34] /*53919*/;
assign _26482_ = _26483_ & D[8] /*53918*/;
assign _26485_ = _25929_ & _26482_ /*53913*/;
assign _26486_ = _25929_ ^ _26482_ /*53916*/;
assign _26487_ = _26478_ & _26486_ /*53914*/;
assign _26377_ = _26478_ ^ _26486_ /*53915*/;
assign _26484_ = _26485_ | _26487_ /*53912*/;
assign _26489_ = ~Q[34] /*53911*/;
assign _26488_ = _26489_ & D[9] /*53910*/;
assign _26491_ = _25930_ & _26488_ /*53905*/;
assign _26492_ = _25930_ ^ _26488_ /*53908*/;
assign _26493_ = _26484_ & _26492_ /*53906*/;
assign _26378_ = _26484_ ^ _26492_ /*53907*/;
assign _26490_ = _26491_ | _26493_ /*53904*/;
assign _26495_ = ~Q[34] /*53903*/;
assign _26494_ = _26495_ & D[10] /*53902*/;
assign _26497_ = _25931_ & _26494_ /*53897*/;
assign _26498_ = _25931_ ^ _26494_ /*53900*/;
assign _26499_ = _26490_ & _26498_ /*53898*/;
assign _26379_ = _26490_ ^ _26498_ /*53899*/;
assign _26496_ = _26497_ | _26499_ /*53896*/;
assign _26501_ = ~Q[34] /*53895*/;
assign _26500_ = _26501_ & D[11] /*53894*/;
assign _26503_ = _25932_ & _26500_ /*53889*/;
assign _26504_ = _25932_ ^ _26500_ /*53892*/;
assign _26505_ = _26496_ & _26504_ /*53890*/;
assign _26380_ = _26496_ ^ _26504_ /*53891*/;
assign _26502_ = _26503_ | _26505_ /*53888*/;
assign _26507_ = ~Q[34] /*53887*/;
assign _26506_ = _26507_ & D[12] /*53886*/;
assign _26509_ = _25933_ & _26506_ /*53881*/;
assign _26510_ = _25933_ ^ _26506_ /*53884*/;
assign _26511_ = _26502_ & _26510_ /*53882*/;
assign _26381_ = _26502_ ^ _26510_ /*53883*/;
assign _26508_ = _26509_ | _26511_ /*53880*/;
assign _26513_ = ~Q[34] /*53879*/;
assign _26512_ = _26513_ & D[13] /*53878*/;
assign _26515_ = _25934_ & _26512_ /*53873*/;
assign _26516_ = _25934_ ^ _26512_ /*53876*/;
assign _26517_ = _26508_ & _26516_ /*53874*/;
assign _26382_ = _26508_ ^ _26516_ /*53875*/;
assign _26514_ = _26515_ | _26517_ /*53872*/;
assign _26519_ = ~Q[34] /*53871*/;
assign _26518_ = _26519_ & D[14] /*53870*/;
assign _26521_ = _25935_ & _26518_ /*53865*/;
assign _26522_ = _25935_ ^ _26518_ /*53868*/;
assign _26523_ = _26514_ & _26522_ /*53866*/;
assign _26383_ = _26514_ ^ _26522_ /*53867*/;
assign _26520_ = _26521_ | _26523_ /*53864*/;
assign _26525_ = ~Q[34] /*53863*/;
assign _26524_ = _26525_ & D[15] /*53862*/;
assign _26527_ = _25936_ & _26524_ /*53857*/;
assign _26528_ = _25936_ ^ _26524_ /*53860*/;
assign _26529_ = _26520_ & _26528_ /*53858*/;
assign _26384_ = _26520_ ^ _26528_ /*53859*/;
assign _26526_ = _26527_ | _26529_ /*53856*/;
assign _26531_ = ~Q[34] /*53855*/;
assign _26530_ = _26531_ & D[16] /*53854*/;
assign _26533_ = _25937_ & _26530_ /*53849*/;
assign _26534_ = _25937_ ^ _26530_ /*53852*/;
assign _26535_ = _26526_ & _26534_ /*53850*/;
assign _26385_ = _26526_ ^ _26534_ /*53851*/;
assign _26532_ = _26533_ | _26535_ /*53848*/;
assign _26537_ = ~Q[34] /*53847*/;
assign _26536_ = _26537_ & D[17] /*53846*/;
assign _26539_ = _25938_ & _26536_ /*53841*/;
assign _26540_ = _25938_ ^ _26536_ /*53844*/;
assign _26541_ = _26532_ & _26540_ /*53842*/;
assign _26386_ = _26532_ ^ _26540_ /*53843*/;
assign _26538_ = _26539_ | _26541_ /*53840*/;
assign _26543_ = ~Q[34] /*53839*/;
assign _26542_ = _26543_ & D[18] /*53838*/;
assign _26545_ = _25939_ & _26542_ /*53833*/;
assign _26546_ = _25939_ ^ _26542_ /*53836*/;
assign _26547_ = _26538_ & _26546_ /*53834*/;
assign _26387_ = _26538_ ^ _26546_ /*53835*/;
assign _26544_ = _26545_ | _26547_ /*53832*/;
assign _26549_ = ~Q[34] /*53831*/;
assign _26548_ = _26549_ & D[19] /*53830*/;
assign _26551_ = _25940_ & _26548_ /*53825*/;
assign _26552_ = _25940_ ^ _26548_ /*53828*/;
assign _26553_ = _26544_ & _26552_ /*53826*/;
assign _26388_ = _26544_ ^ _26552_ /*53827*/;
assign _26550_ = _26551_ | _26553_ /*53824*/;
assign _26555_ = ~Q[34] /*53823*/;
assign _26554_ = _26555_ & D[20] /*53822*/;
assign _26557_ = _25941_ & _26554_ /*53817*/;
assign _26558_ = _25941_ ^ _26554_ /*53820*/;
assign _26559_ = _26550_ & _26558_ /*53818*/;
assign _26389_ = _26550_ ^ _26558_ /*53819*/;
assign _26556_ = _26557_ | _26559_ /*53816*/;
assign _26561_ = ~Q[34] /*53815*/;
assign _26560_ = _26561_ & D[21] /*53814*/;
assign _26563_ = _25942_ & _26560_ /*53809*/;
assign _26564_ = _25942_ ^ _26560_ /*53812*/;
assign _26565_ = _26556_ & _26564_ /*53810*/;
assign _26390_ = _26556_ ^ _26564_ /*53811*/;
assign _26562_ = _26563_ | _26565_ /*53808*/;
assign _26567_ = ~Q[34] /*53807*/;
assign _26566_ = _26567_ & D[22] /*53806*/;
assign _26569_ = _25943_ & _26566_ /*53801*/;
assign _26570_ = _25943_ ^ _26566_ /*53804*/;
assign _26571_ = _26562_ & _26570_ /*53802*/;
assign _26391_ = _26562_ ^ _26570_ /*53803*/;
assign _26568_ = _26569_ | _26571_ /*53800*/;
assign _26573_ = ~Q[34] /*53799*/;
assign _26572_ = _26573_ & D[23] /*53798*/;
assign _26575_ = _25944_ & _26572_ /*53793*/;
assign _26576_ = _25944_ ^ _26572_ /*53796*/;
assign _26577_ = _26568_ & _26576_ /*53794*/;
assign _26392_ = _26568_ ^ _26576_ /*53795*/;
assign _26574_ = _26575_ | _26577_ /*53792*/;
assign _26579_ = ~Q[34] /*53791*/;
assign _26578_ = _26579_ & D[24] /*53790*/;
assign _26581_ = _25945_ & _26578_ /*53785*/;
assign _26582_ = _25945_ ^ _26578_ /*53788*/;
assign _26583_ = _26574_ & _26582_ /*53786*/;
assign _26393_ = _26574_ ^ _26582_ /*53787*/;
assign _26580_ = _26581_ | _26583_ /*53784*/;
assign _26585_ = ~Q[34] /*53783*/;
assign _26584_ = _26585_ & D[25] /*53782*/;
assign _26587_ = _25946_ & _26584_ /*53777*/;
assign _26588_ = _25946_ ^ _26584_ /*53780*/;
assign _26589_ = _26580_ & _26588_ /*53778*/;
assign _26394_ = _26580_ ^ _26588_ /*53779*/;
assign _26586_ = _26587_ | _26589_ /*53776*/;
assign _26591_ = ~Q[34] /*53775*/;
assign _26590_ = _26591_ & D[26] /*53774*/;
assign _26593_ = _25947_ & _26590_ /*53769*/;
assign _26594_ = _25947_ ^ _26590_ /*53772*/;
assign _26595_ = _26586_ & _26594_ /*53770*/;
assign _26395_ = _26586_ ^ _26594_ /*53771*/;
assign _26592_ = _26593_ | _26595_ /*53768*/;
assign _26597_ = ~Q[34] /*53767*/;
assign _26596_ = _26597_ & D[27] /*53766*/;
assign _26599_ = _25948_ & _26596_ /*53761*/;
assign _26600_ = _25948_ ^ _26596_ /*53764*/;
assign _26601_ = _26592_ & _26600_ /*53762*/;
assign _26396_ = _26592_ ^ _26600_ /*53763*/;
assign _26598_ = _26599_ | _26601_ /*53760*/;
assign _26603_ = ~Q[34] /*53759*/;
assign _26602_ = _26603_ & D[28] /*53758*/;
assign _26605_ = _25949_ & _26602_ /*53753*/;
assign _26606_ = _25949_ ^ _26602_ /*53756*/;
assign _26607_ = _26598_ & _26606_ /*53754*/;
assign _26397_ = _26598_ ^ _26606_ /*53755*/;
assign _26604_ = _26605_ | _26607_ /*53752*/;
assign _26609_ = ~Q[34] /*53751*/;
assign _26608_ = _26609_ & D[29] /*53750*/;
assign _26611_ = _25950_ & _26608_ /*53745*/;
assign _26612_ = _25950_ ^ _26608_ /*53748*/;
assign _26613_ = _26604_ & _26612_ /*53746*/;
assign _26398_ = _26604_ ^ _26612_ /*53747*/;
assign _26610_ = _26611_ | _26613_ /*53744*/;
assign _26615_ = ~Q[34] /*53743*/;
assign _26614_ = _26615_ & D[30] /*53742*/;
assign _26617_ = _25951_ & _26614_ /*53737*/;
assign _26618_ = _25951_ ^ _26614_ /*53740*/;
assign _26619_ = _26610_ & _26618_ /*53738*/;
assign _26399_ = _26610_ ^ _26618_ /*53739*/;
assign _26616_ = _26617_ | _26619_ /*53736*/;
assign _26621_ = ~Q[34] /*53735*/;
assign _26620_ = _26621_ & D[31] /*53734*/;
assign _26623_ = _25952_ & _26620_ /*53729*/;
assign _26624_ = _25952_ ^ _26620_ /*53732*/;
assign _26625_ = _26616_ & _26624_ /*53730*/;
assign _26400_ = _26616_ ^ _26624_ /*53731*/;
assign _26622_ = _26623_ | _26625_ /*53728*/;
assign _26627_ = ~Q[34] /*53727*/;
assign _26626_ = _26627_ & D[32] /*53726*/;
assign _26629_ = _25953_ & _26626_ /*53721*/;
assign _26630_ = _25953_ ^ _26626_ /*53724*/;
assign _26631_ = _26622_ & _26630_ /*53722*/;
assign _26401_ = _26622_ ^ _26630_ /*53723*/;
assign _26628_ = _26629_ | _26631_ /*53720*/;
assign _26633_ = ~Q[34] /*53719*/;
assign _26632_ = _26633_ & D[33] /*53718*/;
assign _26635_ = _25954_ & _26632_ /*53713*/;
assign _26636_ = _25954_ ^ _26632_ /*53716*/;
assign _26637_ = _26628_ & _26636_ /*53714*/;
assign _26402_ = _26628_ ^ _26636_ /*53715*/;
assign _26634_ = _26635_ | _26637_ /*53712*/;
assign _26639_ = ~Q[34] /*53711*/;
assign _26638_ = _26639_ & D[34] /*53710*/;
assign _26641_ = _25955_ & _26638_ /*53705*/;
assign _26642_ = _25955_ ^ _26638_ /*53708*/;
assign _26643_ = _26634_ & _26642_ /*53706*/;
assign _26403_ = _26634_ ^ _26642_ /*53707*/;
assign _26640_ = _26641_ | _26643_ /*53704*/;
assign _26645_ = ~Q[34] /*53703*/;
assign _26644_ = _26645_ & D[35] /*53702*/;
assign _26647_ = _25956_ & _26644_ /*53697*/;
assign _26648_ = _25956_ ^ _26644_ /*53700*/;
assign _26649_ = _26640_ & _26648_ /*53698*/;
assign _26404_ = _26640_ ^ _26648_ /*53699*/;
assign _26646_ = _26647_ | _26649_ /*53696*/;
assign _26651_ = ~Q[34] /*53695*/;
assign _26650_ = _26651_ & D[36] /*53694*/;
assign _26653_ = _25957_ & _26650_ /*53689*/;
assign _26654_ = _25957_ ^ _26650_ /*53692*/;
assign _26655_ = _26646_ & _26654_ /*53690*/;
assign _26405_ = _26646_ ^ _26654_ /*53691*/;
assign _26652_ = _26653_ | _26655_ /*53688*/;
assign _26657_ = ~Q[34] /*53687*/;
assign _26656_ = _26657_ & D[37] /*53686*/;
assign _26659_ = _25958_ & _26656_ /*53681*/;
assign _26660_ = _25958_ ^ _26656_ /*53684*/;
assign _26661_ = _26652_ & _26660_ /*53682*/;
assign _26406_ = _26652_ ^ _26660_ /*53683*/;
assign _26658_ = _26659_ | _26661_ /*53680*/;
assign _26663_ = ~Q[34] /*53679*/;
assign _26662_ = _26663_ & D[38] /*53678*/;
assign _26665_ = _25959_ & _26662_ /*53673*/;
assign _26666_ = _25959_ ^ _26662_ /*53676*/;
assign _26667_ = _26658_ & _26666_ /*53674*/;
assign _26407_ = _26658_ ^ _26666_ /*53675*/;
assign _26664_ = _26665_ | _26667_ /*53672*/;
assign _26669_ = ~Q[34] /*53671*/;
assign _26668_ = _26669_ & D[39] /*53670*/;
assign _26671_ = _25960_ & _26668_ /*53665*/;
assign _26672_ = _25960_ ^ _26668_ /*53668*/;
assign _26673_ = _26664_ & _26672_ /*53666*/;
assign _26408_ = _26664_ ^ _26672_ /*53667*/;
assign _26670_ = _26671_ | _26673_ /*53664*/;
assign _26675_ = ~Q[34] /*53663*/;
assign _26674_ = _26675_ & D[40] /*53662*/;
assign _26677_ = _25961_ & _26674_ /*53657*/;
assign _26678_ = _25961_ ^ _26674_ /*53660*/;
assign _26679_ = _26670_ & _26678_ /*53658*/;
assign _26409_ = _26670_ ^ _26678_ /*53659*/;
assign _26676_ = _26677_ | _26679_ /*53656*/;
assign _26681_ = ~Q[34] /*53655*/;
assign _26680_ = _26681_ & D[41] /*53654*/;
assign _26683_ = _25962_ & _26680_ /*53649*/;
assign _26684_ = _25962_ ^ _26680_ /*53652*/;
assign _26685_ = _26676_ & _26684_ /*53650*/;
assign _26410_ = _26676_ ^ _26684_ /*53651*/;
assign _26682_ = _26683_ | _26685_ /*53648*/;
assign _26687_ = ~Q[34] /*53647*/;
assign _26686_ = _26687_ & D[42] /*53646*/;
assign _26689_ = _25963_ & _26686_ /*53641*/;
assign _26690_ = _25963_ ^ _26686_ /*53644*/;
assign _26691_ = _26682_ & _26690_ /*53642*/;
assign _26411_ = _26682_ ^ _26690_ /*53643*/;
assign _26688_ = _26689_ | _26691_ /*53640*/;
assign _26693_ = ~Q[34] /*53639*/;
assign _26692_ = _26693_ & D[43] /*53638*/;
assign _26695_ = _25964_ & _26692_ /*53633*/;
assign _26696_ = _25964_ ^ _26692_ /*53636*/;
assign _26697_ = _26688_ & _26696_ /*53634*/;
assign _26412_ = _26688_ ^ _26696_ /*53635*/;
assign _26694_ = _26695_ | _26697_ /*53632*/;
assign _26699_ = ~Q[34] /*53631*/;
assign _26698_ = _26699_ & D[44] /*53630*/;
assign _26701_ = _25965_ & _26698_ /*53625*/;
assign _26702_ = _25965_ ^ _26698_ /*53628*/;
assign _26703_ = _26694_ & _26702_ /*53626*/;
assign _26413_ = _26694_ ^ _26702_ /*53627*/;
assign _26700_ = _26701_ | _26703_ /*53624*/;
assign _26705_ = ~Q[34] /*53623*/;
assign _26704_ = _26705_ & D[45] /*53622*/;
assign _26707_ = _25966_ & _26704_ /*53617*/;
assign _26708_ = _25966_ ^ _26704_ /*53620*/;
assign _26709_ = _26700_ & _26708_ /*53618*/;
assign _26414_ = _26700_ ^ _26708_ /*53619*/;
assign _26706_ = _26707_ | _26709_ /*53616*/;
assign _26711_ = ~Q[34] /*53615*/;
assign _26710_ = _26711_ & D[46] /*53614*/;
assign _26713_ = _25967_ & _26710_ /*53609*/;
assign _26714_ = _25967_ ^ _26710_ /*53612*/;
assign _26715_ = _26706_ & _26714_ /*53610*/;
assign _26415_ = _26706_ ^ _26714_ /*53611*/;
assign _26712_ = _26713_ | _26715_ /*53608*/;
assign _26717_ = ~Q[34] /*53607*/;
assign _26716_ = _26717_ & D[47] /*53606*/;
assign _26719_ = _25968_ & _26716_ /*53601*/;
assign _26720_ = _25968_ ^ _26716_ /*53604*/;
assign _26721_ = _26712_ & _26720_ /*53602*/;
assign _26416_ = _26712_ ^ _26720_ /*53603*/;
assign _26718_ = _26719_ | _26721_ /*53600*/;
assign _26723_ = ~Q[34] /*53599*/;
assign _26722_ = _26723_ & D[48] /*53598*/;
assign _26725_ = _25969_ & _26722_ /*53593*/;
assign _26726_ = _25969_ ^ _26722_ /*53596*/;
assign _26727_ = _26718_ & _26726_ /*53594*/;
assign _26417_ = _26718_ ^ _26726_ /*53595*/;
assign _26724_ = _26725_ | _26727_ /*53592*/;
assign _26729_ = ~Q[34] /*53591*/;
assign _26728_ = _26729_ & D[49] /*53590*/;
assign _26731_ = _25970_ & _26728_ /*53585*/;
assign _26732_ = _25970_ ^ _26728_ /*53588*/;
assign _26733_ = _26724_ & _26732_ /*53586*/;
assign _26418_ = _26724_ ^ _26732_ /*53587*/;
assign _26730_ = _26731_ | _26733_ /*53584*/;
assign _26735_ = ~Q[34] /*53583*/;
assign _26734_ = _26735_ & D[50] /*53582*/;
assign _26737_ = _25971_ & _26734_ /*53577*/;
assign _26738_ = _25971_ ^ _26734_ /*53580*/;
assign _26739_ = _26730_ & _26738_ /*53578*/;
assign _26419_ = _26730_ ^ _26738_ /*53579*/;
assign _26736_ = _26737_ | _26739_ /*53576*/;
assign _26741_ = ~Q[34] /*53575*/;
assign _26740_ = _26741_ & D[51] /*53574*/;
assign _26743_ = _25972_ & _26740_ /*53569*/;
assign _26744_ = _25972_ ^ _26740_ /*53572*/;
assign _26745_ = _26736_ & _26744_ /*53570*/;
assign _26420_ = _26736_ ^ _26744_ /*53571*/;
assign _26742_ = _26743_ | _26745_ /*53568*/;
assign _26747_ = ~Q[34] /*53567*/;
assign _26746_ = _26747_ & D[52] /*53566*/;
assign _26749_ = _25973_ & _26746_ /*53561*/;
assign _26750_ = _25973_ ^ _26746_ /*53564*/;
assign _26751_ = _26742_ & _26750_ /*53562*/;
assign _26421_ = _26742_ ^ _26750_ /*53563*/;
assign _26748_ = _26749_ | _26751_ /*53560*/;
assign _26753_ = ~Q[34] /*53559*/;
assign _26752_ = _26753_ & D[53] /*53558*/;
assign _26755_ = _25974_ & _26752_ /*53553*/;
assign _26756_ = _25974_ ^ _26752_ /*53556*/;
assign _26757_ = _26748_ & _26756_ /*53554*/;
assign _26422_ = _26748_ ^ _26756_ /*53555*/;
assign _26754_ = _26755_ | _26757_ /*53552*/;
assign _26759_ = ~Q[34] /*53551*/;
assign _26758_ = _26759_ & D[54] /*53550*/;
assign _26761_ = _25975_ & _26758_ /*53545*/;
assign _26762_ = _25975_ ^ _26758_ /*53548*/;
assign _26763_ = _26754_ & _26762_ /*53546*/;
assign _26423_ = _26754_ ^ _26762_ /*53547*/;
assign _26760_ = _26761_ | _26763_ /*53544*/;
assign _26765_ = ~Q[34] /*53543*/;
assign _26764_ = _26765_ & D[55] /*53542*/;
assign _26767_ = _25976_ & _26764_ /*53537*/;
assign _26768_ = _25976_ ^ _26764_ /*53540*/;
assign _26769_ = _26760_ & _26768_ /*53538*/;
assign _26424_ = _26760_ ^ _26768_ /*53539*/;
assign _26766_ = _26767_ | _26769_ /*53536*/;
assign _26771_ = ~Q[34] /*53535*/;
assign _26770_ = _26771_ & D[56] /*53534*/;
assign _26773_ = _25977_ & _26770_ /*53529*/;
assign _26774_ = _25977_ ^ _26770_ /*53532*/;
assign _26775_ = _26766_ & _26774_ /*53530*/;
assign _26425_ = _26766_ ^ _26774_ /*53531*/;
assign _26772_ = _26773_ | _26775_ /*53528*/;
assign _26777_ = ~Q[34] /*53527*/;
assign _26776_ = _26777_ & D[57] /*53526*/;
assign _26779_ = _25978_ & _26776_ /*53521*/;
assign _26780_ = _25978_ ^ _26776_ /*53524*/;
assign _26781_ = _26772_ & _26780_ /*53522*/;
assign _26426_ = _26772_ ^ _26780_ /*53523*/;
assign _26778_ = _26779_ | _26781_ /*53520*/;
assign _26783_ = ~Q[34] /*53519*/;
assign _26782_ = _26783_ & D[58] /*53518*/;
assign _26785_ = _25979_ & _26782_ /*53513*/;
assign _26786_ = _25979_ ^ _26782_ /*53516*/;
assign _26787_ = _26778_ & _26786_ /*53514*/;
assign _26427_ = _26778_ ^ _26786_ /*53515*/;
assign _26784_ = _26785_ | _26787_ /*53512*/;
assign _26789_ = ~Q[34] /*53511*/;
assign _26788_ = _26789_ & D[59] /*53510*/;
assign _26791_ = _25980_ & _26788_ /*53505*/;
assign _26792_ = _25980_ ^ _26788_ /*53508*/;
assign _26793_ = _26784_ & _26792_ /*53506*/;
assign _26428_ = _26784_ ^ _26792_ /*53507*/;
assign _26790_ = _26791_ | _26793_ /*53504*/;
assign _26795_ = ~Q[34] /*53503*/;
assign _26794_ = _26795_ & D[60] /*53502*/;
assign _26797_ = _25981_ & _26794_ /*53497*/;
assign _26798_ = _25981_ ^ _26794_ /*53500*/;
assign _26799_ = _26790_ & _26798_ /*53498*/;
assign _26429_ = _26790_ ^ _26798_ /*53499*/;
assign _26796_ = _26797_ | _26799_ /*53496*/;
assign _26801_ = ~Q[34] /*53495*/;
assign _26800_ = _26801_ & D[61] /*53494*/;
assign _26803_ = _25982_ & _26800_ /*53489*/;
assign _26804_ = _25982_ ^ _26800_ /*53492*/;
assign _26805_ = _26796_ & _26804_ /*53490*/;
assign _26430_ = _26796_ ^ _26804_ /*53491*/;
assign _26802_ = _26803_ | _26805_ /*53488*/;
assign _26807_ = ~Q[34] /*53487*/;
assign _26806_ = _26807_ & D[62] /*53486*/;
assign _26809_ = _25983_ & _26806_ /*53481*/;
assign _26810_ = _25983_ ^ _26806_ /*53484*/;
assign _26811_ = _26802_ & _26810_ /*53482*/;
assign _26431_ = _26802_ ^ _26810_ /*53483*/;
assign _26808_ = _26809_ | _26811_ /*53480*/;
assign _26813_ = ~Q[34] /*53479*/;
assign _26812_ = _26813_ & zeroWire /*53478*/;
assign _26814_ = _25984_ ^ _26812_ /*53476*/;
assign _26432_ = _26814_ ^ _26808_ /*53475*/;
assign _26885_ = ~D[0] /*53221*/;
assign _26882_ = R_0[33] & _26885_ /*53217*/;
assign _26883_ = R_0[33] ^ _26885_ /*53220*/;
assign _26884_ = oneWire & _26883_ /*53218*/;
assign _26817_ = oneWire ^ _26883_ /*53219*/;
assign _26881_ = _26882_ | _26884_ /*53216*/;
assign _26890_ = ~D[1] /*53215*/;
assign _26887_ = _26369_ & _26890_ /*53211*/;
assign _26888_ = _26369_ ^ _26890_ /*53214*/;
assign _26889_ = _26881_ & _26888_ /*53212*/;
assign _26818_ = _26881_ ^ _26888_ /*53213*/;
assign _26886_ = _26887_ | _26889_ /*53210*/;
assign _26895_ = ~D[2] /*53209*/;
assign _26892_ = _26370_ & _26895_ /*53205*/;
assign _26893_ = _26370_ ^ _26895_ /*53208*/;
assign _26894_ = _26886_ & _26893_ /*53206*/;
assign _26819_ = _26886_ ^ _26893_ /*53207*/;
assign _26891_ = _26892_ | _26894_ /*53204*/;
assign _26900_ = ~D[3] /*53203*/;
assign _26897_ = _26371_ & _26900_ /*53199*/;
assign _26898_ = _26371_ ^ _26900_ /*53202*/;
assign _26899_ = _26891_ & _26898_ /*53200*/;
assign _26820_ = _26891_ ^ _26898_ /*53201*/;
assign _26896_ = _26897_ | _26899_ /*53198*/;
assign _26905_ = ~D[4] /*53197*/;
assign _26902_ = _26372_ & _26905_ /*53193*/;
assign _26903_ = _26372_ ^ _26905_ /*53196*/;
assign _26904_ = _26896_ & _26903_ /*53194*/;
assign _26821_ = _26896_ ^ _26903_ /*53195*/;
assign _26901_ = _26902_ | _26904_ /*53192*/;
assign _26910_ = ~D[5] /*53191*/;
assign _26907_ = _26373_ & _26910_ /*53187*/;
assign _26908_ = _26373_ ^ _26910_ /*53190*/;
assign _26909_ = _26901_ & _26908_ /*53188*/;
assign _26822_ = _26901_ ^ _26908_ /*53189*/;
assign _26906_ = _26907_ | _26909_ /*53186*/;
assign _26915_ = ~D[6] /*53185*/;
assign _26912_ = _26374_ & _26915_ /*53181*/;
assign _26913_ = _26374_ ^ _26915_ /*53184*/;
assign _26914_ = _26906_ & _26913_ /*53182*/;
assign _26823_ = _26906_ ^ _26913_ /*53183*/;
assign _26911_ = _26912_ | _26914_ /*53180*/;
assign _26920_ = ~D[7] /*53179*/;
assign _26917_ = _26375_ & _26920_ /*53175*/;
assign _26918_ = _26375_ ^ _26920_ /*53178*/;
assign _26919_ = _26911_ & _26918_ /*53176*/;
assign _26824_ = _26911_ ^ _26918_ /*53177*/;
assign _26916_ = _26917_ | _26919_ /*53174*/;
assign _26925_ = ~D[8] /*53173*/;
assign _26922_ = _26376_ & _26925_ /*53169*/;
assign _26923_ = _26376_ ^ _26925_ /*53172*/;
assign _26924_ = _26916_ & _26923_ /*53170*/;
assign _26825_ = _26916_ ^ _26923_ /*53171*/;
assign _26921_ = _26922_ | _26924_ /*53168*/;
assign _26930_ = ~D[9] /*53167*/;
assign _26927_ = _26377_ & _26930_ /*53163*/;
assign _26928_ = _26377_ ^ _26930_ /*53166*/;
assign _26929_ = _26921_ & _26928_ /*53164*/;
assign _26826_ = _26921_ ^ _26928_ /*53165*/;
assign _26926_ = _26927_ | _26929_ /*53162*/;
assign _26935_ = ~D[10] /*53161*/;
assign _26932_ = _26378_ & _26935_ /*53157*/;
assign _26933_ = _26378_ ^ _26935_ /*53160*/;
assign _26934_ = _26926_ & _26933_ /*53158*/;
assign _26827_ = _26926_ ^ _26933_ /*53159*/;
assign _26931_ = _26932_ | _26934_ /*53156*/;
assign _26940_ = ~D[11] /*53155*/;
assign _26937_ = _26379_ & _26940_ /*53151*/;
assign _26938_ = _26379_ ^ _26940_ /*53154*/;
assign _26939_ = _26931_ & _26938_ /*53152*/;
assign _26828_ = _26931_ ^ _26938_ /*53153*/;
assign _26936_ = _26937_ | _26939_ /*53150*/;
assign _26945_ = ~D[12] /*53149*/;
assign _26942_ = _26380_ & _26945_ /*53145*/;
assign _26943_ = _26380_ ^ _26945_ /*53148*/;
assign _26944_ = _26936_ & _26943_ /*53146*/;
assign _26829_ = _26936_ ^ _26943_ /*53147*/;
assign _26941_ = _26942_ | _26944_ /*53144*/;
assign _26950_ = ~D[13] /*53143*/;
assign _26947_ = _26381_ & _26950_ /*53139*/;
assign _26948_ = _26381_ ^ _26950_ /*53142*/;
assign _26949_ = _26941_ & _26948_ /*53140*/;
assign _26830_ = _26941_ ^ _26948_ /*53141*/;
assign _26946_ = _26947_ | _26949_ /*53138*/;
assign _26955_ = ~D[14] /*53137*/;
assign _26952_ = _26382_ & _26955_ /*53133*/;
assign _26953_ = _26382_ ^ _26955_ /*53136*/;
assign _26954_ = _26946_ & _26953_ /*53134*/;
assign _26831_ = _26946_ ^ _26953_ /*53135*/;
assign _26951_ = _26952_ | _26954_ /*53132*/;
assign _26960_ = ~D[15] /*53131*/;
assign _26957_ = _26383_ & _26960_ /*53127*/;
assign _26958_ = _26383_ ^ _26960_ /*53130*/;
assign _26959_ = _26951_ & _26958_ /*53128*/;
assign _26832_ = _26951_ ^ _26958_ /*53129*/;
assign _26956_ = _26957_ | _26959_ /*53126*/;
assign _26965_ = ~D[16] /*53125*/;
assign _26962_ = _26384_ & _26965_ /*53121*/;
assign _26963_ = _26384_ ^ _26965_ /*53124*/;
assign _26964_ = _26956_ & _26963_ /*53122*/;
assign _26833_ = _26956_ ^ _26963_ /*53123*/;
assign _26961_ = _26962_ | _26964_ /*53120*/;
assign _26970_ = ~D[17] /*53119*/;
assign _26967_ = _26385_ & _26970_ /*53115*/;
assign _26968_ = _26385_ ^ _26970_ /*53118*/;
assign _26969_ = _26961_ & _26968_ /*53116*/;
assign _26834_ = _26961_ ^ _26968_ /*53117*/;
assign _26966_ = _26967_ | _26969_ /*53114*/;
assign _26975_ = ~D[18] /*53113*/;
assign _26972_ = _26386_ & _26975_ /*53109*/;
assign _26973_ = _26386_ ^ _26975_ /*53112*/;
assign _26974_ = _26966_ & _26973_ /*53110*/;
assign _26835_ = _26966_ ^ _26973_ /*53111*/;
assign _26971_ = _26972_ | _26974_ /*53108*/;
assign _26980_ = ~D[19] /*53107*/;
assign _26977_ = _26387_ & _26980_ /*53103*/;
assign _26978_ = _26387_ ^ _26980_ /*53106*/;
assign _26979_ = _26971_ & _26978_ /*53104*/;
assign _26836_ = _26971_ ^ _26978_ /*53105*/;
assign _26976_ = _26977_ | _26979_ /*53102*/;
assign _26985_ = ~D[20] /*53101*/;
assign _26982_ = _26388_ & _26985_ /*53097*/;
assign _26983_ = _26388_ ^ _26985_ /*53100*/;
assign _26984_ = _26976_ & _26983_ /*53098*/;
assign _26837_ = _26976_ ^ _26983_ /*53099*/;
assign _26981_ = _26982_ | _26984_ /*53096*/;
assign _26990_ = ~D[21] /*53095*/;
assign _26987_ = _26389_ & _26990_ /*53091*/;
assign _26988_ = _26389_ ^ _26990_ /*53094*/;
assign _26989_ = _26981_ & _26988_ /*53092*/;
assign _26838_ = _26981_ ^ _26988_ /*53093*/;
assign _26986_ = _26987_ | _26989_ /*53090*/;
assign _26995_ = ~D[22] /*53089*/;
assign _26992_ = _26390_ & _26995_ /*53085*/;
assign _26993_ = _26390_ ^ _26995_ /*53088*/;
assign _26994_ = _26986_ & _26993_ /*53086*/;
assign _26839_ = _26986_ ^ _26993_ /*53087*/;
assign _26991_ = _26992_ | _26994_ /*53084*/;
assign _27000_ = ~D[23] /*53083*/;
assign _26997_ = _26391_ & _27000_ /*53079*/;
assign _26998_ = _26391_ ^ _27000_ /*53082*/;
assign _26999_ = _26991_ & _26998_ /*53080*/;
assign _26840_ = _26991_ ^ _26998_ /*53081*/;
assign _26996_ = _26997_ | _26999_ /*53078*/;
assign _27005_ = ~D[24] /*53077*/;
assign _27002_ = _26392_ & _27005_ /*53073*/;
assign _27003_ = _26392_ ^ _27005_ /*53076*/;
assign _27004_ = _26996_ & _27003_ /*53074*/;
assign _26841_ = _26996_ ^ _27003_ /*53075*/;
assign _27001_ = _27002_ | _27004_ /*53072*/;
assign _27010_ = ~D[25] /*53071*/;
assign _27007_ = _26393_ & _27010_ /*53067*/;
assign _27008_ = _26393_ ^ _27010_ /*53070*/;
assign _27009_ = _27001_ & _27008_ /*53068*/;
assign _26842_ = _27001_ ^ _27008_ /*53069*/;
assign _27006_ = _27007_ | _27009_ /*53066*/;
assign _27015_ = ~D[26] /*53065*/;
assign _27012_ = _26394_ & _27015_ /*53061*/;
assign _27013_ = _26394_ ^ _27015_ /*53064*/;
assign _27014_ = _27006_ & _27013_ /*53062*/;
assign _26843_ = _27006_ ^ _27013_ /*53063*/;
assign _27011_ = _27012_ | _27014_ /*53060*/;
assign _27020_ = ~D[27] /*53059*/;
assign _27017_ = _26395_ & _27020_ /*53055*/;
assign _27018_ = _26395_ ^ _27020_ /*53058*/;
assign _27019_ = _27011_ & _27018_ /*53056*/;
assign _26844_ = _27011_ ^ _27018_ /*53057*/;
assign _27016_ = _27017_ | _27019_ /*53054*/;
assign _27025_ = ~D[28] /*53053*/;
assign _27022_ = _26396_ & _27025_ /*53049*/;
assign _27023_ = _26396_ ^ _27025_ /*53052*/;
assign _27024_ = _27016_ & _27023_ /*53050*/;
assign _26845_ = _27016_ ^ _27023_ /*53051*/;
assign _27021_ = _27022_ | _27024_ /*53048*/;
assign _27030_ = ~D[29] /*53047*/;
assign _27027_ = _26397_ & _27030_ /*53043*/;
assign _27028_ = _26397_ ^ _27030_ /*53046*/;
assign _27029_ = _27021_ & _27028_ /*53044*/;
assign _26846_ = _27021_ ^ _27028_ /*53045*/;
assign _27026_ = _27027_ | _27029_ /*53042*/;
assign _27035_ = ~D[30] /*53041*/;
assign _27032_ = _26398_ & _27035_ /*53037*/;
assign _27033_ = _26398_ ^ _27035_ /*53040*/;
assign _27034_ = _27026_ & _27033_ /*53038*/;
assign _26847_ = _27026_ ^ _27033_ /*53039*/;
assign _27031_ = _27032_ | _27034_ /*53036*/;
assign _27040_ = ~D[31] /*53035*/;
assign _27037_ = _26399_ & _27040_ /*53031*/;
assign _27038_ = _26399_ ^ _27040_ /*53034*/;
assign _27039_ = _27031_ & _27038_ /*53032*/;
assign _26848_ = _27031_ ^ _27038_ /*53033*/;
assign _27036_ = _27037_ | _27039_ /*53030*/;
assign _27045_ = ~D[32] /*53029*/;
assign _27042_ = _26400_ & _27045_ /*53025*/;
assign _27043_ = _26400_ ^ _27045_ /*53028*/;
assign _27044_ = _27036_ & _27043_ /*53026*/;
assign _26849_ = _27036_ ^ _27043_ /*53027*/;
assign _27041_ = _27042_ | _27044_ /*53024*/;
assign _27050_ = ~D[33] /*53023*/;
assign _27047_ = _26401_ & _27050_ /*53019*/;
assign _27048_ = _26401_ ^ _27050_ /*53022*/;
assign _27049_ = _27041_ & _27048_ /*53020*/;
assign _26850_ = _27041_ ^ _27048_ /*53021*/;
assign _27046_ = _27047_ | _27049_ /*53018*/;
assign _27055_ = ~D[34] /*53017*/;
assign _27052_ = _26402_ & _27055_ /*53013*/;
assign _27053_ = _26402_ ^ _27055_ /*53016*/;
assign _27054_ = _27046_ & _27053_ /*53014*/;
assign _26851_ = _27046_ ^ _27053_ /*53015*/;
assign _27051_ = _27052_ | _27054_ /*53012*/;
assign _27060_ = ~D[35] /*53011*/;
assign _27057_ = _26403_ & _27060_ /*53007*/;
assign _27058_ = _26403_ ^ _27060_ /*53010*/;
assign _27059_ = _27051_ & _27058_ /*53008*/;
assign _26852_ = _27051_ ^ _27058_ /*53009*/;
assign _27056_ = _27057_ | _27059_ /*53006*/;
assign _27065_ = ~D[36] /*53005*/;
assign _27062_ = _26404_ & _27065_ /*53001*/;
assign _27063_ = _26404_ ^ _27065_ /*53004*/;
assign _27064_ = _27056_ & _27063_ /*53002*/;
assign _26853_ = _27056_ ^ _27063_ /*53003*/;
assign _27061_ = _27062_ | _27064_ /*53000*/;
assign _27070_ = ~D[37] /*52999*/;
assign _27067_ = _26405_ & _27070_ /*52995*/;
assign _27068_ = _26405_ ^ _27070_ /*52998*/;
assign _27069_ = _27061_ & _27068_ /*52996*/;
assign _26854_ = _27061_ ^ _27068_ /*52997*/;
assign _27066_ = _27067_ | _27069_ /*52994*/;
assign _27075_ = ~D[38] /*52993*/;
assign _27072_ = _26406_ & _27075_ /*52989*/;
assign _27073_ = _26406_ ^ _27075_ /*52992*/;
assign _27074_ = _27066_ & _27073_ /*52990*/;
assign _26855_ = _27066_ ^ _27073_ /*52991*/;
assign _27071_ = _27072_ | _27074_ /*52988*/;
assign _27080_ = ~D[39] /*52987*/;
assign _27077_ = _26407_ & _27080_ /*52983*/;
assign _27078_ = _26407_ ^ _27080_ /*52986*/;
assign _27079_ = _27071_ & _27078_ /*52984*/;
assign _26856_ = _27071_ ^ _27078_ /*52985*/;
assign _27076_ = _27077_ | _27079_ /*52982*/;
assign _27085_ = ~D[40] /*52981*/;
assign _27082_ = _26408_ & _27085_ /*52977*/;
assign _27083_ = _26408_ ^ _27085_ /*52980*/;
assign _27084_ = _27076_ & _27083_ /*52978*/;
assign _26857_ = _27076_ ^ _27083_ /*52979*/;
assign _27081_ = _27082_ | _27084_ /*52976*/;
assign _27090_ = ~D[41] /*52975*/;
assign _27087_ = _26409_ & _27090_ /*52971*/;
assign _27088_ = _26409_ ^ _27090_ /*52974*/;
assign _27089_ = _27081_ & _27088_ /*52972*/;
assign _26858_ = _27081_ ^ _27088_ /*52973*/;
assign _27086_ = _27087_ | _27089_ /*52970*/;
assign _27095_ = ~D[42] /*52969*/;
assign _27092_ = _26410_ & _27095_ /*52965*/;
assign _27093_ = _26410_ ^ _27095_ /*52968*/;
assign _27094_ = _27086_ & _27093_ /*52966*/;
assign _26859_ = _27086_ ^ _27093_ /*52967*/;
assign _27091_ = _27092_ | _27094_ /*52964*/;
assign _27100_ = ~D[43] /*52963*/;
assign _27097_ = _26411_ & _27100_ /*52959*/;
assign _27098_ = _26411_ ^ _27100_ /*52962*/;
assign _27099_ = _27091_ & _27098_ /*52960*/;
assign _26860_ = _27091_ ^ _27098_ /*52961*/;
assign _27096_ = _27097_ | _27099_ /*52958*/;
assign _27105_ = ~D[44] /*52957*/;
assign _27102_ = _26412_ & _27105_ /*52953*/;
assign _27103_ = _26412_ ^ _27105_ /*52956*/;
assign _27104_ = _27096_ & _27103_ /*52954*/;
assign _26861_ = _27096_ ^ _27103_ /*52955*/;
assign _27101_ = _27102_ | _27104_ /*52952*/;
assign _27110_ = ~D[45] /*52951*/;
assign _27107_ = _26413_ & _27110_ /*52947*/;
assign _27108_ = _26413_ ^ _27110_ /*52950*/;
assign _27109_ = _27101_ & _27108_ /*52948*/;
assign _26862_ = _27101_ ^ _27108_ /*52949*/;
assign _27106_ = _27107_ | _27109_ /*52946*/;
assign _27115_ = ~D[46] /*52945*/;
assign _27112_ = _26414_ & _27115_ /*52941*/;
assign _27113_ = _26414_ ^ _27115_ /*52944*/;
assign _27114_ = _27106_ & _27113_ /*52942*/;
assign _26863_ = _27106_ ^ _27113_ /*52943*/;
assign _27111_ = _27112_ | _27114_ /*52940*/;
assign _27120_ = ~D[47] /*52939*/;
assign _27117_ = _26415_ & _27120_ /*52935*/;
assign _27118_ = _26415_ ^ _27120_ /*52938*/;
assign _27119_ = _27111_ & _27118_ /*52936*/;
assign _26864_ = _27111_ ^ _27118_ /*52937*/;
assign _27116_ = _27117_ | _27119_ /*52934*/;
assign _27125_ = ~D[48] /*52933*/;
assign _27122_ = _26416_ & _27125_ /*52929*/;
assign _27123_ = _26416_ ^ _27125_ /*52932*/;
assign _27124_ = _27116_ & _27123_ /*52930*/;
assign _26865_ = _27116_ ^ _27123_ /*52931*/;
assign _27121_ = _27122_ | _27124_ /*52928*/;
assign _27130_ = ~D[49] /*52927*/;
assign _27127_ = _26417_ & _27130_ /*52923*/;
assign _27128_ = _26417_ ^ _27130_ /*52926*/;
assign _27129_ = _27121_ & _27128_ /*52924*/;
assign _26866_ = _27121_ ^ _27128_ /*52925*/;
assign _27126_ = _27127_ | _27129_ /*52922*/;
assign _27135_ = ~D[50] /*52921*/;
assign _27132_ = _26418_ & _27135_ /*52917*/;
assign _27133_ = _26418_ ^ _27135_ /*52920*/;
assign _27134_ = _27126_ & _27133_ /*52918*/;
assign _26867_ = _27126_ ^ _27133_ /*52919*/;
assign _27131_ = _27132_ | _27134_ /*52916*/;
assign _27140_ = ~D[51] /*52915*/;
assign _27137_ = _26419_ & _27140_ /*52911*/;
assign _27138_ = _26419_ ^ _27140_ /*52914*/;
assign _27139_ = _27131_ & _27138_ /*52912*/;
assign _26868_ = _27131_ ^ _27138_ /*52913*/;
assign _27136_ = _27137_ | _27139_ /*52910*/;
assign _27145_ = ~D[52] /*52909*/;
assign _27142_ = _26420_ & _27145_ /*52905*/;
assign _27143_ = _26420_ ^ _27145_ /*52908*/;
assign _27144_ = _27136_ & _27143_ /*52906*/;
assign _26869_ = _27136_ ^ _27143_ /*52907*/;
assign _27141_ = _27142_ | _27144_ /*52904*/;
assign _27150_ = ~D[53] /*52903*/;
assign _27147_ = _26421_ & _27150_ /*52899*/;
assign _27148_ = _26421_ ^ _27150_ /*52902*/;
assign _27149_ = _27141_ & _27148_ /*52900*/;
assign _26870_ = _27141_ ^ _27148_ /*52901*/;
assign _27146_ = _27147_ | _27149_ /*52898*/;
assign _27155_ = ~D[54] /*52897*/;
assign _27152_ = _26422_ & _27155_ /*52893*/;
assign _27153_ = _26422_ ^ _27155_ /*52896*/;
assign _27154_ = _27146_ & _27153_ /*52894*/;
assign _26871_ = _27146_ ^ _27153_ /*52895*/;
assign _27151_ = _27152_ | _27154_ /*52892*/;
assign _27160_ = ~D[55] /*52891*/;
assign _27157_ = _26423_ & _27160_ /*52887*/;
assign _27158_ = _26423_ ^ _27160_ /*52890*/;
assign _27159_ = _27151_ & _27158_ /*52888*/;
assign _26872_ = _27151_ ^ _27158_ /*52889*/;
assign _27156_ = _27157_ | _27159_ /*52886*/;
assign _27165_ = ~D[56] /*52885*/;
assign _27162_ = _26424_ & _27165_ /*52881*/;
assign _27163_ = _26424_ ^ _27165_ /*52884*/;
assign _27164_ = _27156_ & _27163_ /*52882*/;
assign _26873_ = _27156_ ^ _27163_ /*52883*/;
assign _27161_ = _27162_ | _27164_ /*52880*/;
assign _27170_ = ~D[57] /*52879*/;
assign _27167_ = _26425_ & _27170_ /*52875*/;
assign _27168_ = _26425_ ^ _27170_ /*52878*/;
assign _27169_ = _27161_ & _27168_ /*52876*/;
assign _26874_ = _27161_ ^ _27168_ /*52877*/;
assign _27166_ = _27167_ | _27169_ /*52874*/;
assign _27175_ = ~D[58] /*52873*/;
assign _27172_ = _26426_ & _27175_ /*52869*/;
assign _27173_ = _26426_ ^ _27175_ /*52872*/;
assign _27174_ = _27166_ & _27173_ /*52870*/;
assign _26875_ = _27166_ ^ _27173_ /*52871*/;
assign _27171_ = _27172_ | _27174_ /*52868*/;
assign _27180_ = ~D[59] /*52867*/;
assign _27177_ = _26427_ & _27180_ /*52863*/;
assign _27178_ = _26427_ ^ _27180_ /*52866*/;
assign _27179_ = _27171_ & _27178_ /*52864*/;
assign _26876_ = _27171_ ^ _27178_ /*52865*/;
assign _27176_ = _27177_ | _27179_ /*52862*/;
assign _27185_ = ~D[60] /*52861*/;
assign _27182_ = _26428_ & _27185_ /*52857*/;
assign _27183_ = _26428_ ^ _27185_ /*52860*/;
assign _27184_ = _27176_ & _27183_ /*52858*/;
assign _26877_ = _27176_ ^ _27183_ /*52859*/;
assign _27181_ = _27182_ | _27184_ /*52856*/;
assign _27190_ = ~D[61] /*52855*/;
assign _27187_ = _26429_ & _27190_ /*52851*/;
assign _27188_ = _26429_ ^ _27190_ /*52854*/;
assign _27189_ = _27181_ & _27188_ /*52852*/;
assign _26878_ = _27181_ ^ _27188_ /*52853*/;
assign _27186_ = _27187_ | _27189_ /*52850*/;
assign _27195_ = ~D[62] /*52849*/;
assign _27192_ = _26430_ & _27195_ /*52845*/;
assign _27193_ = _26430_ ^ _27195_ /*52848*/;
assign _27194_ = _27186_ & _27193_ /*52846*/;
assign _26879_ = _27186_ ^ _27193_ /*52847*/;
assign _27191_ = _27192_ | _27194_ /*52844*/;
assign _27196_ = _26431_ & oneWire /*52839*/;
assign _27197_ = _26431_ ^ oneWire /*52842*/;
assign _27198_ = _27191_ & _27197_ /*52840*/;
assign _26880_ = _27191_ ^ _27197_ /*52841*/;
assign Q[33] = _27196_ | _27198_ /*52838*/;
assign _27331_ = ~Q[33] /*52453*/;
assign _27330_ = _27331_ & D[0] /*52452*/;
assign _27333_ = _26817_ & _27330_ /*52447*/;
assign _27334_ = _26817_ ^ _27330_ /*52450*/;
assign _27335_ = zeroWire & _27334_ /*52448*/;
assign _27265_ = zeroWire ^ _27334_ /*52449*/;
assign _27332_ = _27333_ | _27335_ /*52446*/;
assign _27337_ = ~Q[33] /*52445*/;
assign _27336_ = _27337_ & D[1] /*52444*/;
assign _27339_ = _26818_ & _27336_ /*52439*/;
assign _27340_ = _26818_ ^ _27336_ /*52442*/;
assign _27341_ = _27332_ & _27340_ /*52440*/;
assign _27266_ = _27332_ ^ _27340_ /*52441*/;
assign _27338_ = _27339_ | _27341_ /*52438*/;
assign _27343_ = ~Q[33] /*52437*/;
assign _27342_ = _27343_ & D[2] /*52436*/;
assign _27345_ = _26819_ & _27342_ /*52431*/;
assign _27346_ = _26819_ ^ _27342_ /*52434*/;
assign _27347_ = _27338_ & _27346_ /*52432*/;
assign _27267_ = _27338_ ^ _27346_ /*52433*/;
assign _27344_ = _27345_ | _27347_ /*52430*/;
assign _27349_ = ~Q[33] /*52429*/;
assign _27348_ = _27349_ & D[3] /*52428*/;
assign _27351_ = _26820_ & _27348_ /*52423*/;
assign _27352_ = _26820_ ^ _27348_ /*52426*/;
assign _27353_ = _27344_ & _27352_ /*52424*/;
assign _27268_ = _27344_ ^ _27352_ /*52425*/;
assign _27350_ = _27351_ | _27353_ /*52422*/;
assign _27355_ = ~Q[33] /*52421*/;
assign _27354_ = _27355_ & D[4] /*52420*/;
assign _27357_ = _26821_ & _27354_ /*52415*/;
assign _27358_ = _26821_ ^ _27354_ /*52418*/;
assign _27359_ = _27350_ & _27358_ /*52416*/;
assign _27269_ = _27350_ ^ _27358_ /*52417*/;
assign _27356_ = _27357_ | _27359_ /*52414*/;
assign _27361_ = ~Q[33] /*52413*/;
assign _27360_ = _27361_ & D[5] /*52412*/;
assign _27363_ = _26822_ & _27360_ /*52407*/;
assign _27364_ = _26822_ ^ _27360_ /*52410*/;
assign _27365_ = _27356_ & _27364_ /*52408*/;
assign _27270_ = _27356_ ^ _27364_ /*52409*/;
assign _27362_ = _27363_ | _27365_ /*52406*/;
assign _27367_ = ~Q[33] /*52405*/;
assign _27366_ = _27367_ & D[6] /*52404*/;
assign _27369_ = _26823_ & _27366_ /*52399*/;
assign _27370_ = _26823_ ^ _27366_ /*52402*/;
assign _27371_ = _27362_ & _27370_ /*52400*/;
assign _27271_ = _27362_ ^ _27370_ /*52401*/;
assign _27368_ = _27369_ | _27371_ /*52398*/;
assign _27373_ = ~Q[33] /*52397*/;
assign _27372_ = _27373_ & D[7] /*52396*/;
assign _27375_ = _26824_ & _27372_ /*52391*/;
assign _27376_ = _26824_ ^ _27372_ /*52394*/;
assign _27377_ = _27368_ & _27376_ /*52392*/;
assign _27272_ = _27368_ ^ _27376_ /*52393*/;
assign _27374_ = _27375_ | _27377_ /*52390*/;
assign _27379_ = ~Q[33] /*52389*/;
assign _27378_ = _27379_ & D[8] /*52388*/;
assign _27381_ = _26825_ & _27378_ /*52383*/;
assign _27382_ = _26825_ ^ _27378_ /*52386*/;
assign _27383_ = _27374_ & _27382_ /*52384*/;
assign _27273_ = _27374_ ^ _27382_ /*52385*/;
assign _27380_ = _27381_ | _27383_ /*52382*/;
assign _27385_ = ~Q[33] /*52381*/;
assign _27384_ = _27385_ & D[9] /*52380*/;
assign _27387_ = _26826_ & _27384_ /*52375*/;
assign _27388_ = _26826_ ^ _27384_ /*52378*/;
assign _27389_ = _27380_ & _27388_ /*52376*/;
assign _27274_ = _27380_ ^ _27388_ /*52377*/;
assign _27386_ = _27387_ | _27389_ /*52374*/;
assign _27391_ = ~Q[33] /*52373*/;
assign _27390_ = _27391_ & D[10] /*52372*/;
assign _27393_ = _26827_ & _27390_ /*52367*/;
assign _27394_ = _26827_ ^ _27390_ /*52370*/;
assign _27395_ = _27386_ & _27394_ /*52368*/;
assign _27275_ = _27386_ ^ _27394_ /*52369*/;
assign _27392_ = _27393_ | _27395_ /*52366*/;
assign _27397_ = ~Q[33] /*52365*/;
assign _27396_ = _27397_ & D[11] /*52364*/;
assign _27399_ = _26828_ & _27396_ /*52359*/;
assign _27400_ = _26828_ ^ _27396_ /*52362*/;
assign _27401_ = _27392_ & _27400_ /*52360*/;
assign _27276_ = _27392_ ^ _27400_ /*52361*/;
assign _27398_ = _27399_ | _27401_ /*52358*/;
assign _27403_ = ~Q[33] /*52357*/;
assign _27402_ = _27403_ & D[12] /*52356*/;
assign _27405_ = _26829_ & _27402_ /*52351*/;
assign _27406_ = _26829_ ^ _27402_ /*52354*/;
assign _27407_ = _27398_ & _27406_ /*52352*/;
assign _27277_ = _27398_ ^ _27406_ /*52353*/;
assign _27404_ = _27405_ | _27407_ /*52350*/;
assign _27409_ = ~Q[33] /*52349*/;
assign _27408_ = _27409_ & D[13] /*52348*/;
assign _27411_ = _26830_ & _27408_ /*52343*/;
assign _27412_ = _26830_ ^ _27408_ /*52346*/;
assign _27413_ = _27404_ & _27412_ /*52344*/;
assign _27278_ = _27404_ ^ _27412_ /*52345*/;
assign _27410_ = _27411_ | _27413_ /*52342*/;
assign _27415_ = ~Q[33] /*52341*/;
assign _27414_ = _27415_ & D[14] /*52340*/;
assign _27417_ = _26831_ & _27414_ /*52335*/;
assign _27418_ = _26831_ ^ _27414_ /*52338*/;
assign _27419_ = _27410_ & _27418_ /*52336*/;
assign _27279_ = _27410_ ^ _27418_ /*52337*/;
assign _27416_ = _27417_ | _27419_ /*52334*/;
assign _27421_ = ~Q[33] /*52333*/;
assign _27420_ = _27421_ & D[15] /*52332*/;
assign _27423_ = _26832_ & _27420_ /*52327*/;
assign _27424_ = _26832_ ^ _27420_ /*52330*/;
assign _27425_ = _27416_ & _27424_ /*52328*/;
assign _27280_ = _27416_ ^ _27424_ /*52329*/;
assign _27422_ = _27423_ | _27425_ /*52326*/;
assign _27427_ = ~Q[33] /*52325*/;
assign _27426_ = _27427_ & D[16] /*52324*/;
assign _27429_ = _26833_ & _27426_ /*52319*/;
assign _27430_ = _26833_ ^ _27426_ /*52322*/;
assign _27431_ = _27422_ & _27430_ /*52320*/;
assign _27281_ = _27422_ ^ _27430_ /*52321*/;
assign _27428_ = _27429_ | _27431_ /*52318*/;
assign _27433_ = ~Q[33] /*52317*/;
assign _27432_ = _27433_ & D[17] /*52316*/;
assign _27435_ = _26834_ & _27432_ /*52311*/;
assign _27436_ = _26834_ ^ _27432_ /*52314*/;
assign _27437_ = _27428_ & _27436_ /*52312*/;
assign _27282_ = _27428_ ^ _27436_ /*52313*/;
assign _27434_ = _27435_ | _27437_ /*52310*/;
assign _27439_ = ~Q[33] /*52309*/;
assign _27438_ = _27439_ & D[18] /*52308*/;
assign _27441_ = _26835_ & _27438_ /*52303*/;
assign _27442_ = _26835_ ^ _27438_ /*52306*/;
assign _27443_ = _27434_ & _27442_ /*52304*/;
assign _27283_ = _27434_ ^ _27442_ /*52305*/;
assign _27440_ = _27441_ | _27443_ /*52302*/;
assign _27445_ = ~Q[33] /*52301*/;
assign _27444_ = _27445_ & D[19] /*52300*/;
assign _27447_ = _26836_ & _27444_ /*52295*/;
assign _27448_ = _26836_ ^ _27444_ /*52298*/;
assign _27449_ = _27440_ & _27448_ /*52296*/;
assign _27284_ = _27440_ ^ _27448_ /*52297*/;
assign _27446_ = _27447_ | _27449_ /*52294*/;
assign _27451_ = ~Q[33] /*52293*/;
assign _27450_ = _27451_ & D[20] /*52292*/;
assign _27453_ = _26837_ & _27450_ /*52287*/;
assign _27454_ = _26837_ ^ _27450_ /*52290*/;
assign _27455_ = _27446_ & _27454_ /*52288*/;
assign _27285_ = _27446_ ^ _27454_ /*52289*/;
assign _27452_ = _27453_ | _27455_ /*52286*/;
assign _27457_ = ~Q[33] /*52285*/;
assign _27456_ = _27457_ & D[21] /*52284*/;
assign _27459_ = _26838_ & _27456_ /*52279*/;
assign _27460_ = _26838_ ^ _27456_ /*52282*/;
assign _27461_ = _27452_ & _27460_ /*52280*/;
assign _27286_ = _27452_ ^ _27460_ /*52281*/;
assign _27458_ = _27459_ | _27461_ /*52278*/;
assign _27463_ = ~Q[33] /*52277*/;
assign _27462_ = _27463_ & D[22] /*52276*/;
assign _27465_ = _26839_ & _27462_ /*52271*/;
assign _27466_ = _26839_ ^ _27462_ /*52274*/;
assign _27467_ = _27458_ & _27466_ /*52272*/;
assign _27287_ = _27458_ ^ _27466_ /*52273*/;
assign _27464_ = _27465_ | _27467_ /*52270*/;
assign _27469_ = ~Q[33] /*52269*/;
assign _27468_ = _27469_ & D[23] /*52268*/;
assign _27471_ = _26840_ & _27468_ /*52263*/;
assign _27472_ = _26840_ ^ _27468_ /*52266*/;
assign _27473_ = _27464_ & _27472_ /*52264*/;
assign _27288_ = _27464_ ^ _27472_ /*52265*/;
assign _27470_ = _27471_ | _27473_ /*52262*/;
assign _27475_ = ~Q[33] /*52261*/;
assign _27474_ = _27475_ & D[24] /*52260*/;
assign _27477_ = _26841_ & _27474_ /*52255*/;
assign _27478_ = _26841_ ^ _27474_ /*52258*/;
assign _27479_ = _27470_ & _27478_ /*52256*/;
assign _27289_ = _27470_ ^ _27478_ /*52257*/;
assign _27476_ = _27477_ | _27479_ /*52254*/;
assign _27481_ = ~Q[33] /*52253*/;
assign _27480_ = _27481_ & D[25] /*52252*/;
assign _27483_ = _26842_ & _27480_ /*52247*/;
assign _27484_ = _26842_ ^ _27480_ /*52250*/;
assign _27485_ = _27476_ & _27484_ /*52248*/;
assign _27290_ = _27476_ ^ _27484_ /*52249*/;
assign _27482_ = _27483_ | _27485_ /*52246*/;
assign _27487_ = ~Q[33] /*52245*/;
assign _27486_ = _27487_ & D[26] /*52244*/;
assign _27489_ = _26843_ & _27486_ /*52239*/;
assign _27490_ = _26843_ ^ _27486_ /*52242*/;
assign _27491_ = _27482_ & _27490_ /*52240*/;
assign _27291_ = _27482_ ^ _27490_ /*52241*/;
assign _27488_ = _27489_ | _27491_ /*52238*/;
assign _27493_ = ~Q[33] /*52237*/;
assign _27492_ = _27493_ & D[27] /*52236*/;
assign _27495_ = _26844_ & _27492_ /*52231*/;
assign _27496_ = _26844_ ^ _27492_ /*52234*/;
assign _27497_ = _27488_ & _27496_ /*52232*/;
assign _27292_ = _27488_ ^ _27496_ /*52233*/;
assign _27494_ = _27495_ | _27497_ /*52230*/;
assign _27499_ = ~Q[33] /*52229*/;
assign _27498_ = _27499_ & D[28] /*52228*/;
assign _27501_ = _26845_ & _27498_ /*52223*/;
assign _27502_ = _26845_ ^ _27498_ /*52226*/;
assign _27503_ = _27494_ & _27502_ /*52224*/;
assign _27293_ = _27494_ ^ _27502_ /*52225*/;
assign _27500_ = _27501_ | _27503_ /*52222*/;
assign _27505_ = ~Q[33] /*52221*/;
assign _27504_ = _27505_ & D[29] /*52220*/;
assign _27507_ = _26846_ & _27504_ /*52215*/;
assign _27508_ = _26846_ ^ _27504_ /*52218*/;
assign _27509_ = _27500_ & _27508_ /*52216*/;
assign _27294_ = _27500_ ^ _27508_ /*52217*/;
assign _27506_ = _27507_ | _27509_ /*52214*/;
assign _27511_ = ~Q[33] /*52213*/;
assign _27510_ = _27511_ & D[30] /*52212*/;
assign _27513_ = _26847_ & _27510_ /*52207*/;
assign _27514_ = _26847_ ^ _27510_ /*52210*/;
assign _27515_ = _27506_ & _27514_ /*52208*/;
assign _27295_ = _27506_ ^ _27514_ /*52209*/;
assign _27512_ = _27513_ | _27515_ /*52206*/;
assign _27517_ = ~Q[33] /*52205*/;
assign _27516_ = _27517_ & D[31] /*52204*/;
assign _27519_ = _26848_ & _27516_ /*52199*/;
assign _27520_ = _26848_ ^ _27516_ /*52202*/;
assign _27521_ = _27512_ & _27520_ /*52200*/;
assign _27296_ = _27512_ ^ _27520_ /*52201*/;
assign _27518_ = _27519_ | _27521_ /*52198*/;
assign _27523_ = ~Q[33] /*52197*/;
assign _27522_ = _27523_ & D[32] /*52196*/;
assign _27525_ = _26849_ & _27522_ /*52191*/;
assign _27526_ = _26849_ ^ _27522_ /*52194*/;
assign _27527_ = _27518_ & _27526_ /*52192*/;
assign _27297_ = _27518_ ^ _27526_ /*52193*/;
assign _27524_ = _27525_ | _27527_ /*52190*/;
assign _27529_ = ~Q[33] /*52189*/;
assign _27528_ = _27529_ & D[33] /*52188*/;
assign _27531_ = _26850_ & _27528_ /*52183*/;
assign _27532_ = _26850_ ^ _27528_ /*52186*/;
assign _27533_ = _27524_ & _27532_ /*52184*/;
assign _27298_ = _27524_ ^ _27532_ /*52185*/;
assign _27530_ = _27531_ | _27533_ /*52182*/;
assign _27535_ = ~Q[33] /*52181*/;
assign _27534_ = _27535_ & D[34] /*52180*/;
assign _27537_ = _26851_ & _27534_ /*52175*/;
assign _27538_ = _26851_ ^ _27534_ /*52178*/;
assign _27539_ = _27530_ & _27538_ /*52176*/;
assign _27299_ = _27530_ ^ _27538_ /*52177*/;
assign _27536_ = _27537_ | _27539_ /*52174*/;
assign _27541_ = ~Q[33] /*52173*/;
assign _27540_ = _27541_ & D[35] /*52172*/;
assign _27543_ = _26852_ & _27540_ /*52167*/;
assign _27544_ = _26852_ ^ _27540_ /*52170*/;
assign _27545_ = _27536_ & _27544_ /*52168*/;
assign _27300_ = _27536_ ^ _27544_ /*52169*/;
assign _27542_ = _27543_ | _27545_ /*52166*/;
assign _27547_ = ~Q[33] /*52165*/;
assign _27546_ = _27547_ & D[36] /*52164*/;
assign _27549_ = _26853_ & _27546_ /*52159*/;
assign _27550_ = _26853_ ^ _27546_ /*52162*/;
assign _27551_ = _27542_ & _27550_ /*52160*/;
assign _27301_ = _27542_ ^ _27550_ /*52161*/;
assign _27548_ = _27549_ | _27551_ /*52158*/;
assign _27553_ = ~Q[33] /*52157*/;
assign _27552_ = _27553_ & D[37] /*52156*/;
assign _27555_ = _26854_ & _27552_ /*52151*/;
assign _27556_ = _26854_ ^ _27552_ /*52154*/;
assign _27557_ = _27548_ & _27556_ /*52152*/;
assign _27302_ = _27548_ ^ _27556_ /*52153*/;
assign _27554_ = _27555_ | _27557_ /*52150*/;
assign _27559_ = ~Q[33] /*52149*/;
assign _27558_ = _27559_ & D[38] /*52148*/;
assign _27561_ = _26855_ & _27558_ /*52143*/;
assign _27562_ = _26855_ ^ _27558_ /*52146*/;
assign _27563_ = _27554_ & _27562_ /*52144*/;
assign _27303_ = _27554_ ^ _27562_ /*52145*/;
assign _27560_ = _27561_ | _27563_ /*52142*/;
assign _27565_ = ~Q[33] /*52141*/;
assign _27564_ = _27565_ & D[39] /*52140*/;
assign _27567_ = _26856_ & _27564_ /*52135*/;
assign _27568_ = _26856_ ^ _27564_ /*52138*/;
assign _27569_ = _27560_ & _27568_ /*52136*/;
assign _27304_ = _27560_ ^ _27568_ /*52137*/;
assign _27566_ = _27567_ | _27569_ /*52134*/;
assign _27571_ = ~Q[33] /*52133*/;
assign _27570_ = _27571_ & D[40] /*52132*/;
assign _27573_ = _26857_ & _27570_ /*52127*/;
assign _27574_ = _26857_ ^ _27570_ /*52130*/;
assign _27575_ = _27566_ & _27574_ /*52128*/;
assign _27305_ = _27566_ ^ _27574_ /*52129*/;
assign _27572_ = _27573_ | _27575_ /*52126*/;
assign _27577_ = ~Q[33] /*52125*/;
assign _27576_ = _27577_ & D[41] /*52124*/;
assign _27579_ = _26858_ & _27576_ /*52119*/;
assign _27580_ = _26858_ ^ _27576_ /*52122*/;
assign _27581_ = _27572_ & _27580_ /*52120*/;
assign _27306_ = _27572_ ^ _27580_ /*52121*/;
assign _27578_ = _27579_ | _27581_ /*52118*/;
assign _27583_ = ~Q[33] /*52117*/;
assign _27582_ = _27583_ & D[42] /*52116*/;
assign _27585_ = _26859_ & _27582_ /*52111*/;
assign _27586_ = _26859_ ^ _27582_ /*52114*/;
assign _27587_ = _27578_ & _27586_ /*52112*/;
assign _27307_ = _27578_ ^ _27586_ /*52113*/;
assign _27584_ = _27585_ | _27587_ /*52110*/;
assign _27589_ = ~Q[33] /*52109*/;
assign _27588_ = _27589_ & D[43] /*52108*/;
assign _27591_ = _26860_ & _27588_ /*52103*/;
assign _27592_ = _26860_ ^ _27588_ /*52106*/;
assign _27593_ = _27584_ & _27592_ /*52104*/;
assign _27308_ = _27584_ ^ _27592_ /*52105*/;
assign _27590_ = _27591_ | _27593_ /*52102*/;
assign _27595_ = ~Q[33] /*52101*/;
assign _27594_ = _27595_ & D[44] /*52100*/;
assign _27597_ = _26861_ & _27594_ /*52095*/;
assign _27598_ = _26861_ ^ _27594_ /*52098*/;
assign _27599_ = _27590_ & _27598_ /*52096*/;
assign _27309_ = _27590_ ^ _27598_ /*52097*/;
assign _27596_ = _27597_ | _27599_ /*52094*/;
assign _27601_ = ~Q[33] /*52093*/;
assign _27600_ = _27601_ & D[45] /*52092*/;
assign _27603_ = _26862_ & _27600_ /*52087*/;
assign _27604_ = _26862_ ^ _27600_ /*52090*/;
assign _27605_ = _27596_ & _27604_ /*52088*/;
assign _27310_ = _27596_ ^ _27604_ /*52089*/;
assign _27602_ = _27603_ | _27605_ /*52086*/;
assign _27607_ = ~Q[33] /*52085*/;
assign _27606_ = _27607_ & D[46] /*52084*/;
assign _27609_ = _26863_ & _27606_ /*52079*/;
assign _27610_ = _26863_ ^ _27606_ /*52082*/;
assign _27611_ = _27602_ & _27610_ /*52080*/;
assign _27311_ = _27602_ ^ _27610_ /*52081*/;
assign _27608_ = _27609_ | _27611_ /*52078*/;
assign _27613_ = ~Q[33] /*52077*/;
assign _27612_ = _27613_ & D[47] /*52076*/;
assign _27615_ = _26864_ & _27612_ /*52071*/;
assign _27616_ = _26864_ ^ _27612_ /*52074*/;
assign _27617_ = _27608_ & _27616_ /*52072*/;
assign _27312_ = _27608_ ^ _27616_ /*52073*/;
assign _27614_ = _27615_ | _27617_ /*52070*/;
assign _27619_ = ~Q[33] /*52069*/;
assign _27618_ = _27619_ & D[48] /*52068*/;
assign _27621_ = _26865_ & _27618_ /*52063*/;
assign _27622_ = _26865_ ^ _27618_ /*52066*/;
assign _27623_ = _27614_ & _27622_ /*52064*/;
assign _27313_ = _27614_ ^ _27622_ /*52065*/;
assign _27620_ = _27621_ | _27623_ /*52062*/;
assign _27625_ = ~Q[33] /*52061*/;
assign _27624_ = _27625_ & D[49] /*52060*/;
assign _27627_ = _26866_ & _27624_ /*52055*/;
assign _27628_ = _26866_ ^ _27624_ /*52058*/;
assign _27629_ = _27620_ & _27628_ /*52056*/;
assign _27314_ = _27620_ ^ _27628_ /*52057*/;
assign _27626_ = _27627_ | _27629_ /*52054*/;
assign _27631_ = ~Q[33] /*52053*/;
assign _27630_ = _27631_ & D[50] /*52052*/;
assign _27633_ = _26867_ & _27630_ /*52047*/;
assign _27634_ = _26867_ ^ _27630_ /*52050*/;
assign _27635_ = _27626_ & _27634_ /*52048*/;
assign _27315_ = _27626_ ^ _27634_ /*52049*/;
assign _27632_ = _27633_ | _27635_ /*52046*/;
assign _27637_ = ~Q[33] /*52045*/;
assign _27636_ = _27637_ & D[51] /*52044*/;
assign _27639_ = _26868_ & _27636_ /*52039*/;
assign _27640_ = _26868_ ^ _27636_ /*52042*/;
assign _27641_ = _27632_ & _27640_ /*52040*/;
assign _27316_ = _27632_ ^ _27640_ /*52041*/;
assign _27638_ = _27639_ | _27641_ /*52038*/;
assign _27643_ = ~Q[33] /*52037*/;
assign _27642_ = _27643_ & D[52] /*52036*/;
assign _27645_ = _26869_ & _27642_ /*52031*/;
assign _27646_ = _26869_ ^ _27642_ /*52034*/;
assign _27647_ = _27638_ & _27646_ /*52032*/;
assign _27317_ = _27638_ ^ _27646_ /*52033*/;
assign _27644_ = _27645_ | _27647_ /*52030*/;
assign _27649_ = ~Q[33] /*52029*/;
assign _27648_ = _27649_ & D[53] /*52028*/;
assign _27651_ = _26870_ & _27648_ /*52023*/;
assign _27652_ = _26870_ ^ _27648_ /*52026*/;
assign _27653_ = _27644_ & _27652_ /*52024*/;
assign _27318_ = _27644_ ^ _27652_ /*52025*/;
assign _27650_ = _27651_ | _27653_ /*52022*/;
assign _27655_ = ~Q[33] /*52021*/;
assign _27654_ = _27655_ & D[54] /*52020*/;
assign _27657_ = _26871_ & _27654_ /*52015*/;
assign _27658_ = _26871_ ^ _27654_ /*52018*/;
assign _27659_ = _27650_ & _27658_ /*52016*/;
assign _27319_ = _27650_ ^ _27658_ /*52017*/;
assign _27656_ = _27657_ | _27659_ /*52014*/;
assign _27661_ = ~Q[33] /*52013*/;
assign _27660_ = _27661_ & D[55] /*52012*/;
assign _27663_ = _26872_ & _27660_ /*52007*/;
assign _27664_ = _26872_ ^ _27660_ /*52010*/;
assign _27665_ = _27656_ & _27664_ /*52008*/;
assign _27320_ = _27656_ ^ _27664_ /*52009*/;
assign _27662_ = _27663_ | _27665_ /*52006*/;
assign _27667_ = ~Q[33] /*52005*/;
assign _27666_ = _27667_ & D[56] /*52004*/;
assign _27669_ = _26873_ & _27666_ /*51999*/;
assign _27670_ = _26873_ ^ _27666_ /*52002*/;
assign _27671_ = _27662_ & _27670_ /*52000*/;
assign _27321_ = _27662_ ^ _27670_ /*52001*/;
assign _27668_ = _27669_ | _27671_ /*51998*/;
assign _27673_ = ~Q[33] /*51997*/;
assign _27672_ = _27673_ & D[57] /*51996*/;
assign _27675_ = _26874_ & _27672_ /*51991*/;
assign _27676_ = _26874_ ^ _27672_ /*51994*/;
assign _27677_ = _27668_ & _27676_ /*51992*/;
assign _27322_ = _27668_ ^ _27676_ /*51993*/;
assign _27674_ = _27675_ | _27677_ /*51990*/;
assign _27679_ = ~Q[33] /*51989*/;
assign _27678_ = _27679_ & D[58] /*51988*/;
assign _27681_ = _26875_ & _27678_ /*51983*/;
assign _27682_ = _26875_ ^ _27678_ /*51986*/;
assign _27683_ = _27674_ & _27682_ /*51984*/;
assign _27323_ = _27674_ ^ _27682_ /*51985*/;
assign _27680_ = _27681_ | _27683_ /*51982*/;
assign _27685_ = ~Q[33] /*51981*/;
assign _27684_ = _27685_ & D[59] /*51980*/;
assign _27687_ = _26876_ & _27684_ /*51975*/;
assign _27688_ = _26876_ ^ _27684_ /*51978*/;
assign _27689_ = _27680_ & _27688_ /*51976*/;
assign _27324_ = _27680_ ^ _27688_ /*51977*/;
assign _27686_ = _27687_ | _27689_ /*51974*/;
assign _27691_ = ~Q[33] /*51973*/;
assign _27690_ = _27691_ & D[60] /*51972*/;
assign _27693_ = _26877_ & _27690_ /*51967*/;
assign _27694_ = _26877_ ^ _27690_ /*51970*/;
assign _27695_ = _27686_ & _27694_ /*51968*/;
assign _27325_ = _27686_ ^ _27694_ /*51969*/;
assign _27692_ = _27693_ | _27695_ /*51966*/;
assign _27697_ = ~Q[33] /*51965*/;
assign _27696_ = _27697_ & D[61] /*51964*/;
assign _27699_ = _26878_ & _27696_ /*51959*/;
assign _27700_ = _26878_ ^ _27696_ /*51962*/;
assign _27701_ = _27692_ & _27700_ /*51960*/;
assign _27326_ = _27692_ ^ _27700_ /*51961*/;
assign _27698_ = _27699_ | _27701_ /*51958*/;
assign _27703_ = ~Q[33] /*51957*/;
assign _27702_ = _27703_ & D[62] /*51956*/;
assign _27705_ = _26879_ & _27702_ /*51951*/;
assign _27706_ = _26879_ ^ _27702_ /*51954*/;
assign _27707_ = _27698_ & _27706_ /*51952*/;
assign _27327_ = _27698_ ^ _27706_ /*51953*/;
assign _27704_ = _27705_ | _27707_ /*51950*/;
assign _27709_ = ~Q[33] /*51949*/;
assign _27708_ = _27709_ & zeroWire /*51948*/;
assign _27710_ = _26880_ ^ _27708_ /*51946*/;
assign _27328_ = _27710_ ^ _27704_ /*51945*/;
assign _27781_ = ~D[0] /*51691*/;
assign _27778_ = R_0[32] & _27781_ /*51687*/;
assign _27779_ = R_0[32] ^ _27781_ /*51690*/;
assign _27780_ = oneWire & _27779_ /*51688*/;
assign _27713_ = oneWire ^ _27779_ /*51689*/;
assign _27777_ = _27778_ | _27780_ /*51686*/;
assign _27786_ = ~D[1] /*51685*/;
assign _27783_ = _27265_ & _27786_ /*51681*/;
assign _27784_ = _27265_ ^ _27786_ /*51684*/;
assign _27785_ = _27777_ & _27784_ /*51682*/;
assign _27714_ = _27777_ ^ _27784_ /*51683*/;
assign _27782_ = _27783_ | _27785_ /*51680*/;
assign _27791_ = ~D[2] /*51679*/;
assign _27788_ = _27266_ & _27791_ /*51675*/;
assign _27789_ = _27266_ ^ _27791_ /*51678*/;
assign _27790_ = _27782_ & _27789_ /*51676*/;
assign _27715_ = _27782_ ^ _27789_ /*51677*/;
assign _27787_ = _27788_ | _27790_ /*51674*/;
assign _27796_ = ~D[3] /*51673*/;
assign _27793_ = _27267_ & _27796_ /*51669*/;
assign _27794_ = _27267_ ^ _27796_ /*51672*/;
assign _27795_ = _27787_ & _27794_ /*51670*/;
assign _27716_ = _27787_ ^ _27794_ /*51671*/;
assign _27792_ = _27793_ | _27795_ /*51668*/;
assign _27801_ = ~D[4] /*51667*/;
assign _27798_ = _27268_ & _27801_ /*51663*/;
assign _27799_ = _27268_ ^ _27801_ /*51666*/;
assign _27800_ = _27792_ & _27799_ /*51664*/;
assign _27717_ = _27792_ ^ _27799_ /*51665*/;
assign _27797_ = _27798_ | _27800_ /*51662*/;
assign _27806_ = ~D[5] /*51661*/;
assign _27803_ = _27269_ & _27806_ /*51657*/;
assign _27804_ = _27269_ ^ _27806_ /*51660*/;
assign _27805_ = _27797_ & _27804_ /*51658*/;
assign _27718_ = _27797_ ^ _27804_ /*51659*/;
assign _27802_ = _27803_ | _27805_ /*51656*/;
assign _27811_ = ~D[6] /*51655*/;
assign _27808_ = _27270_ & _27811_ /*51651*/;
assign _27809_ = _27270_ ^ _27811_ /*51654*/;
assign _27810_ = _27802_ & _27809_ /*51652*/;
assign _27719_ = _27802_ ^ _27809_ /*51653*/;
assign _27807_ = _27808_ | _27810_ /*51650*/;
assign _27816_ = ~D[7] /*51649*/;
assign _27813_ = _27271_ & _27816_ /*51645*/;
assign _27814_ = _27271_ ^ _27816_ /*51648*/;
assign _27815_ = _27807_ & _27814_ /*51646*/;
assign _27720_ = _27807_ ^ _27814_ /*51647*/;
assign _27812_ = _27813_ | _27815_ /*51644*/;
assign _27821_ = ~D[8] /*51643*/;
assign _27818_ = _27272_ & _27821_ /*51639*/;
assign _27819_ = _27272_ ^ _27821_ /*51642*/;
assign _27820_ = _27812_ & _27819_ /*51640*/;
assign _27721_ = _27812_ ^ _27819_ /*51641*/;
assign _27817_ = _27818_ | _27820_ /*51638*/;
assign _27826_ = ~D[9] /*51637*/;
assign _27823_ = _27273_ & _27826_ /*51633*/;
assign _27824_ = _27273_ ^ _27826_ /*51636*/;
assign _27825_ = _27817_ & _27824_ /*51634*/;
assign _27722_ = _27817_ ^ _27824_ /*51635*/;
assign _27822_ = _27823_ | _27825_ /*51632*/;
assign _27831_ = ~D[10] /*51631*/;
assign _27828_ = _27274_ & _27831_ /*51627*/;
assign _27829_ = _27274_ ^ _27831_ /*51630*/;
assign _27830_ = _27822_ & _27829_ /*51628*/;
assign _27723_ = _27822_ ^ _27829_ /*51629*/;
assign _27827_ = _27828_ | _27830_ /*51626*/;
assign _27836_ = ~D[11] /*51625*/;
assign _27833_ = _27275_ & _27836_ /*51621*/;
assign _27834_ = _27275_ ^ _27836_ /*51624*/;
assign _27835_ = _27827_ & _27834_ /*51622*/;
assign _27724_ = _27827_ ^ _27834_ /*51623*/;
assign _27832_ = _27833_ | _27835_ /*51620*/;
assign _27841_ = ~D[12] /*51619*/;
assign _27838_ = _27276_ & _27841_ /*51615*/;
assign _27839_ = _27276_ ^ _27841_ /*51618*/;
assign _27840_ = _27832_ & _27839_ /*51616*/;
assign _27725_ = _27832_ ^ _27839_ /*51617*/;
assign _27837_ = _27838_ | _27840_ /*51614*/;
assign _27846_ = ~D[13] /*51613*/;
assign _27843_ = _27277_ & _27846_ /*51609*/;
assign _27844_ = _27277_ ^ _27846_ /*51612*/;
assign _27845_ = _27837_ & _27844_ /*51610*/;
assign _27726_ = _27837_ ^ _27844_ /*51611*/;
assign _27842_ = _27843_ | _27845_ /*51608*/;
assign _27851_ = ~D[14] /*51607*/;
assign _27848_ = _27278_ & _27851_ /*51603*/;
assign _27849_ = _27278_ ^ _27851_ /*51606*/;
assign _27850_ = _27842_ & _27849_ /*51604*/;
assign _27727_ = _27842_ ^ _27849_ /*51605*/;
assign _27847_ = _27848_ | _27850_ /*51602*/;
assign _27856_ = ~D[15] /*51601*/;
assign _27853_ = _27279_ & _27856_ /*51597*/;
assign _27854_ = _27279_ ^ _27856_ /*51600*/;
assign _27855_ = _27847_ & _27854_ /*51598*/;
assign _27728_ = _27847_ ^ _27854_ /*51599*/;
assign _27852_ = _27853_ | _27855_ /*51596*/;
assign _27861_ = ~D[16] /*51595*/;
assign _27858_ = _27280_ & _27861_ /*51591*/;
assign _27859_ = _27280_ ^ _27861_ /*51594*/;
assign _27860_ = _27852_ & _27859_ /*51592*/;
assign _27729_ = _27852_ ^ _27859_ /*51593*/;
assign _27857_ = _27858_ | _27860_ /*51590*/;
assign _27866_ = ~D[17] /*51589*/;
assign _27863_ = _27281_ & _27866_ /*51585*/;
assign _27864_ = _27281_ ^ _27866_ /*51588*/;
assign _27865_ = _27857_ & _27864_ /*51586*/;
assign _27730_ = _27857_ ^ _27864_ /*51587*/;
assign _27862_ = _27863_ | _27865_ /*51584*/;
assign _27871_ = ~D[18] /*51583*/;
assign _27868_ = _27282_ & _27871_ /*51579*/;
assign _27869_ = _27282_ ^ _27871_ /*51582*/;
assign _27870_ = _27862_ & _27869_ /*51580*/;
assign _27731_ = _27862_ ^ _27869_ /*51581*/;
assign _27867_ = _27868_ | _27870_ /*51578*/;
assign _27876_ = ~D[19] /*51577*/;
assign _27873_ = _27283_ & _27876_ /*51573*/;
assign _27874_ = _27283_ ^ _27876_ /*51576*/;
assign _27875_ = _27867_ & _27874_ /*51574*/;
assign _27732_ = _27867_ ^ _27874_ /*51575*/;
assign _27872_ = _27873_ | _27875_ /*51572*/;
assign _27881_ = ~D[20] /*51571*/;
assign _27878_ = _27284_ & _27881_ /*51567*/;
assign _27879_ = _27284_ ^ _27881_ /*51570*/;
assign _27880_ = _27872_ & _27879_ /*51568*/;
assign _27733_ = _27872_ ^ _27879_ /*51569*/;
assign _27877_ = _27878_ | _27880_ /*51566*/;
assign _27886_ = ~D[21] /*51565*/;
assign _27883_ = _27285_ & _27886_ /*51561*/;
assign _27884_ = _27285_ ^ _27886_ /*51564*/;
assign _27885_ = _27877_ & _27884_ /*51562*/;
assign _27734_ = _27877_ ^ _27884_ /*51563*/;
assign _27882_ = _27883_ | _27885_ /*51560*/;
assign _27891_ = ~D[22] /*51559*/;
assign _27888_ = _27286_ & _27891_ /*51555*/;
assign _27889_ = _27286_ ^ _27891_ /*51558*/;
assign _27890_ = _27882_ & _27889_ /*51556*/;
assign _27735_ = _27882_ ^ _27889_ /*51557*/;
assign _27887_ = _27888_ | _27890_ /*51554*/;
assign _27896_ = ~D[23] /*51553*/;
assign _27893_ = _27287_ & _27896_ /*51549*/;
assign _27894_ = _27287_ ^ _27896_ /*51552*/;
assign _27895_ = _27887_ & _27894_ /*51550*/;
assign _27736_ = _27887_ ^ _27894_ /*51551*/;
assign _27892_ = _27893_ | _27895_ /*51548*/;
assign _27901_ = ~D[24] /*51547*/;
assign _27898_ = _27288_ & _27901_ /*51543*/;
assign _27899_ = _27288_ ^ _27901_ /*51546*/;
assign _27900_ = _27892_ & _27899_ /*51544*/;
assign _27737_ = _27892_ ^ _27899_ /*51545*/;
assign _27897_ = _27898_ | _27900_ /*51542*/;
assign _27906_ = ~D[25] /*51541*/;
assign _27903_ = _27289_ & _27906_ /*51537*/;
assign _27904_ = _27289_ ^ _27906_ /*51540*/;
assign _27905_ = _27897_ & _27904_ /*51538*/;
assign _27738_ = _27897_ ^ _27904_ /*51539*/;
assign _27902_ = _27903_ | _27905_ /*51536*/;
assign _27911_ = ~D[26] /*51535*/;
assign _27908_ = _27290_ & _27911_ /*51531*/;
assign _27909_ = _27290_ ^ _27911_ /*51534*/;
assign _27910_ = _27902_ & _27909_ /*51532*/;
assign _27739_ = _27902_ ^ _27909_ /*51533*/;
assign _27907_ = _27908_ | _27910_ /*51530*/;
assign _27916_ = ~D[27] /*51529*/;
assign _27913_ = _27291_ & _27916_ /*51525*/;
assign _27914_ = _27291_ ^ _27916_ /*51528*/;
assign _27915_ = _27907_ & _27914_ /*51526*/;
assign _27740_ = _27907_ ^ _27914_ /*51527*/;
assign _27912_ = _27913_ | _27915_ /*51524*/;
assign _27921_ = ~D[28] /*51523*/;
assign _27918_ = _27292_ & _27921_ /*51519*/;
assign _27919_ = _27292_ ^ _27921_ /*51522*/;
assign _27920_ = _27912_ & _27919_ /*51520*/;
assign _27741_ = _27912_ ^ _27919_ /*51521*/;
assign _27917_ = _27918_ | _27920_ /*51518*/;
assign _27926_ = ~D[29] /*51517*/;
assign _27923_ = _27293_ & _27926_ /*51513*/;
assign _27924_ = _27293_ ^ _27926_ /*51516*/;
assign _27925_ = _27917_ & _27924_ /*51514*/;
assign _27742_ = _27917_ ^ _27924_ /*51515*/;
assign _27922_ = _27923_ | _27925_ /*51512*/;
assign _27931_ = ~D[30] /*51511*/;
assign _27928_ = _27294_ & _27931_ /*51507*/;
assign _27929_ = _27294_ ^ _27931_ /*51510*/;
assign _27930_ = _27922_ & _27929_ /*51508*/;
assign _27743_ = _27922_ ^ _27929_ /*51509*/;
assign _27927_ = _27928_ | _27930_ /*51506*/;
assign _27936_ = ~D[31] /*51505*/;
assign _27933_ = _27295_ & _27936_ /*51501*/;
assign _27934_ = _27295_ ^ _27936_ /*51504*/;
assign _27935_ = _27927_ & _27934_ /*51502*/;
assign _27744_ = _27927_ ^ _27934_ /*51503*/;
assign _27932_ = _27933_ | _27935_ /*51500*/;
assign _27941_ = ~D[32] /*51499*/;
assign _27938_ = _27296_ & _27941_ /*51495*/;
assign _27939_ = _27296_ ^ _27941_ /*51498*/;
assign _27940_ = _27932_ & _27939_ /*51496*/;
assign _27745_ = _27932_ ^ _27939_ /*51497*/;
assign _27937_ = _27938_ | _27940_ /*51494*/;
assign _27946_ = ~D[33] /*51493*/;
assign _27943_ = _27297_ & _27946_ /*51489*/;
assign _27944_ = _27297_ ^ _27946_ /*51492*/;
assign _27945_ = _27937_ & _27944_ /*51490*/;
assign _27746_ = _27937_ ^ _27944_ /*51491*/;
assign _27942_ = _27943_ | _27945_ /*51488*/;
assign _27951_ = ~D[34] /*51487*/;
assign _27948_ = _27298_ & _27951_ /*51483*/;
assign _27949_ = _27298_ ^ _27951_ /*51486*/;
assign _27950_ = _27942_ & _27949_ /*51484*/;
assign _27747_ = _27942_ ^ _27949_ /*51485*/;
assign _27947_ = _27948_ | _27950_ /*51482*/;
assign _27956_ = ~D[35] /*51481*/;
assign _27953_ = _27299_ & _27956_ /*51477*/;
assign _27954_ = _27299_ ^ _27956_ /*51480*/;
assign _27955_ = _27947_ & _27954_ /*51478*/;
assign _27748_ = _27947_ ^ _27954_ /*51479*/;
assign _27952_ = _27953_ | _27955_ /*51476*/;
assign _27961_ = ~D[36] /*51475*/;
assign _27958_ = _27300_ & _27961_ /*51471*/;
assign _27959_ = _27300_ ^ _27961_ /*51474*/;
assign _27960_ = _27952_ & _27959_ /*51472*/;
assign _27749_ = _27952_ ^ _27959_ /*51473*/;
assign _27957_ = _27958_ | _27960_ /*51470*/;
assign _27966_ = ~D[37] /*51469*/;
assign _27963_ = _27301_ & _27966_ /*51465*/;
assign _27964_ = _27301_ ^ _27966_ /*51468*/;
assign _27965_ = _27957_ & _27964_ /*51466*/;
assign _27750_ = _27957_ ^ _27964_ /*51467*/;
assign _27962_ = _27963_ | _27965_ /*51464*/;
assign _27971_ = ~D[38] /*51463*/;
assign _27968_ = _27302_ & _27971_ /*51459*/;
assign _27969_ = _27302_ ^ _27971_ /*51462*/;
assign _27970_ = _27962_ & _27969_ /*51460*/;
assign _27751_ = _27962_ ^ _27969_ /*51461*/;
assign _27967_ = _27968_ | _27970_ /*51458*/;
assign _27976_ = ~D[39] /*51457*/;
assign _27973_ = _27303_ & _27976_ /*51453*/;
assign _27974_ = _27303_ ^ _27976_ /*51456*/;
assign _27975_ = _27967_ & _27974_ /*51454*/;
assign _27752_ = _27967_ ^ _27974_ /*51455*/;
assign _27972_ = _27973_ | _27975_ /*51452*/;
assign _27981_ = ~D[40] /*51451*/;
assign _27978_ = _27304_ & _27981_ /*51447*/;
assign _27979_ = _27304_ ^ _27981_ /*51450*/;
assign _27980_ = _27972_ & _27979_ /*51448*/;
assign _27753_ = _27972_ ^ _27979_ /*51449*/;
assign _27977_ = _27978_ | _27980_ /*51446*/;
assign _27986_ = ~D[41] /*51445*/;
assign _27983_ = _27305_ & _27986_ /*51441*/;
assign _27984_ = _27305_ ^ _27986_ /*51444*/;
assign _27985_ = _27977_ & _27984_ /*51442*/;
assign _27754_ = _27977_ ^ _27984_ /*51443*/;
assign _27982_ = _27983_ | _27985_ /*51440*/;
assign _27991_ = ~D[42] /*51439*/;
assign _27988_ = _27306_ & _27991_ /*51435*/;
assign _27989_ = _27306_ ^ _27991_ /*51438*/;
assign _27990_ = _27982_ & _27989_ /*51436*/;
assign _27755_ = _27982_ ^ _27989_ /*51437*/;
assign _27987_ = _27988_ | _27990_ /*51434*/;
assign _27996_ = ~D[43] /*51433*/;
assign _27993_ = _27307_ & _27996_ /*51429*/;
assign _27994_ = _27307_ ^ _27996_ /*51432*/;
assign _27995_ = _27987_ & _27994_ /*51430*/;
assign _27756_ = _27987_ ^ _27994_ /*51431*/;
assign _27992_ = _27993_ | _27995_ /*51428*/;
assign _28001_ = ~D[44] /*51427*/;
assign _27998_ = _27308_ & _28001_ /*51423*/;
assign _27999_ = _27308_ ^ _28001_ /*51426*/;
assign _28000_ = _27992_ & _27999_ /*51424*/;
assign _27757_ = _27992_ ^ _27999_ /*51425*/;
assign _27997_ = _27998_ | _28000_ /*51422*/;
assign _28006_ = ~D[45] /*51421*/;
assign _28003_ = _27309_ & _28006_ /*51417*/;
assign _28004_ = _27309_ ^ _28006_ /*51420*/;
assign _28005_ = _27997_ & _28004_ /*51418*/;
assign _27758_ = _27997_ ^ _28004_ /*51419*/;
assign _28002_ = _28003_ | _28005_ /*51416*/;
assign _28011_ = ~D[46] /*51415*/;
assign _28008_ = _27310_ & _28011_ /*51411*/;
assign _28009_ = _27310_ ^ _28011_ /*51414*/;
assign _28010_ = _28002_ & _28009_ /*51412*/;
assign _27759_ = _28002_ ^ _28009_ /*51413*/;
assign _28007_ = _28008_ | _28010_ /*51410*/;
assign _28016_ = ~D[47] /*51409*/;
assign _28013_ = _27311_ & _28016_ /*51405*/;
assign _28014_ = _27311_ ^ _28016_ /*51408*/;
assign _28015_ = _28007_ & _28014_ /*51406*/;
assign _27760_ = _28007_ ^ _28014_ /*51407*/;
assign _28012_ = _28013_ | _28015_ /*51404*/;
assign _28021_ = ~D[48] /*51403*/;
assign _28018_ = _27312_ & _28021_ /*51399*/;
assign _28019_ = _27312_ ^ _28021_ /*51402*/;
assign _28020_ = _28012_ & _28019_ /*51400*/;
assign _27761_ = _28012_ ^ _28019_ /*51401*/;
assign _28017_ = _28018_ | _28020_ /*51398*/;
assign _28026_ = ~D[49] /*51397*/;
assign _28023_ = _27313_ & _28026_ /*51393*/;
assign _28024_ = _27313_ ^ _28026_ /*51396*/;
assign _28025_ = _28017_ & _28024_ /*51394*/;
assign _27762_ = _28017_ ^ _28024_ /*51395*/;
assign _28022_ = _28023_ | _28025_ /*51392*/;
assign _28031_ = ~D[50] /*51391*/;
assign _28028_ = _27314_ & _28031_ /*51387*/;
assign _28029_ = _27314_ ^ _28031_ /*51390*/;
assign _28030_ = _28022_ & _28029_ /*51388*/;
assign _27763_ = _28022_ ^ _28029_ /*51389*/;
assign _28027_ = _28028_ | _28030_ /*51386*/;
assign _28036_ = ~D[51] /*51385*/;
assign _28033_ = _27315_ & _28036_ /*51381*/;
assign _28034_ = _27315_ ^ _28036_ /*51384*/;
assign _28035_ = _28027_ & _28034_ /*51382*/;
assign _27764_ = _28027_ ^ _28034_ /*51383*/;
assign _28032_ = _28033_ | _28035_ /*51380*/;
assign _28041_ = ~D[52] /*51379*/;
assign _28038_ = _27316_ & _28041_ /*51375*/;
assign _28039_ = _27316_ ^ _28041_ /*51378*/;
assign _28040_ = _28032_ & _28039_ /*51376*/;
assign _27765_ = _28032_ ^ _28039_ /*51377*/;
assign _28037_ = _28038_ | _28040_ /*51374*/;
assign _28046_ = ~D[53] /*51373*/;
assign _28043_ = _27317_ & _28046_ /*51369*/;
assign _28044_ = _27317_ ^ _28046_ /*51372*/;
assign _28045_ = _28037_ & _28044_ /*51370*/;
assign _27766_ = _28037_ ^ _28044_ /*51371*/;
assign _28042_ = _28043_ | _28045_ /*51368*/;
assign _28051_ = ~D[54] /*51367*/;
assign _28048_ = _27318_ & _28051_ /*51363*/;
assign _28049_ = _27318_ ^ _28051_ /*51366*/;
assign _28050_ = _28042_ & _28049_ /*51364*/;
assign _27767_ = _28042_ ^ _28049_ /*51365*/;
assign _28047_ = _28048_ | _28050_ /*51362*/;
assign _28056_ = ~D[55] /*51361*/;
assign _28053_ = _27319_ & _28056_ /*51357*/;
assign _28054_ = _27319_ ^ _28056_ /*51360*/;
assign _28055_ = _28047_ & _28054_ /*51358*/;
assign _27768_ = _28047_ ^ _28054_ /*51359*/;
assign _28052_ = _28053_ | _28055_ /*51356*/;
assign _28061_ = ~D[56] /*51355*/;
assign _28058_ = _27320_ & _28061_ /*51351*/;
assign _28059_ = _27320_ ^ _28061_ /*51354*/;
assign _28060_ = _28052_ & _28059_ /*51352*/;
assign _27769_ = _28052_ ^ _28059_ /*51353*/;
assign _28057_ = _28058_ | _28060_ /*51350*/;
assign _28066_ = ~D[57] /*51349*/;
assign _28063_ = _27321_ & _28066_ /*51345*/;
assign _28064_ = _27321_ ^ _28066_ /*51348*/;
assign _28065_ = _28057_ & _28064_ /*51346*/;
assign _27770_ = _28057_ ^ _28064_ /*51347*/;
assign _28062_ = _28063_ | _28065_ /*51344*/;
assign _28071_ = ~D[58] /*51343*/;
assign _28068_ = _27322_ & _28071_ /*51339*/;
assign _28069_ = _27322_ ^ _28071_ /*51342*/;
assign _28070_ = _28062_ & _28069_ /*51340*/;
assign _27771_ = _28062_ ^ _28069_ /*51341*/;
assign _28067_ = _28068_ | _28070_ /*51338*/;
assign _28076_ = ~D[59] /*51337*/;
assign _28073_ = _27323_ & _28076_ /*51333*/;
assign _28074_ = _27323_ ^ _28076_ /*51336*/;
assign _28075_ = _28067_ & _28074_ /*51334*/;
assign _27772_ = _28067_ ^ _28074_ /*51335*/;
assign _28072_ = _28073_ | _28075_ /*51332*/;
assign _28081_ = ~D[60] /*51331*/;
assign _28078_ = _27324_ & _28081_ /*51327*/;
assign _28079_ = _27324_ ^ _28081_ /*51330*/;
assign _28080_ = _28072_ & _28079_ /*51328*/;
assign _27773_ = _28072_ ^ _28079_ /*51329*/;
assign _28077_ = _28078_ | _28080_ /*51326*/;
assign _28086_ = ~D[61] /*51325*/;
assign _28083_ = _27325_ & _28086_ /*51321*/;
assign _28084_ = _27325_ ^ _28086_ /*51324*/;
assign _28085_ = _28077_ & _28084_ /*51322*/;
assign _27774_ = _28077_ ^ _28084_ /*51323*/;
assign _28082_ = _28083_ | _28085_ /*51320*/;
assign _28091_ = ~D[62] /*51319*/;
assign _28088_ = _27326_ & _28091_ /*51315*/;
assign _28089_ = _27326_ ^ _28091_ /*51318*/;
assign _28090_ = _28082_ & _28089_ /*51316*/;
assign _27775_ = _28082_ ^ _28089_ /*51317*/;
assign _28087_ = _28088_ | _28090_ /*51314*/;
assign _28092_ = _27327_ & oneWire /*51309*/;
assign _28093_ = _27327_ ^ oneWire /*51312*/;
assign _28094_ = _28087_ & _28093_ /*51310*/;
assign _27776_ = _28087_ ^ _28093_ /*51311*/;
assign Q[32] = _28092_ | _28094_ /*51308*/;
assign _28227_ = ~Q[32] /*50923*/;
assign _28226_ = _28227_ & D[0] /*50922*/;
assign _28229_ = _27713_ & _28226_ /*50917*/;
assign _28230_ = _27713_ ^ _28226_ /*50920*/;
assign _28231_ = zeroWire & _28230_ /*50918*/;
assign _28161_ = zeroWire ^ _28230_ /*50919*/;
assign _28228_ = _28229_ | _28231_ /*50916*/;
assign _28233_ = ~Q[32] /*50915*/;
assign _28232_ = _28233_ & D[1] /*50914*/;
assign _28235_ = _27714_ & _28232_ /*50909*/;
assign _28236_ = _27714_ ^ _28232_ /*50912*/;
assign _28237_ = _28228_ & _28236_ /*50910*/;
assign _28162_ = _28228_ ^ _28236_ /*50911*/;
assign _28234_ = _28235_ | _28237_ /*50908*/;
assign _28239_ = ~Q[32] /*50907*/;
assign _28238_ = _28239_ & D[2] /*50906*/;
assign _28241_ = _27715_ & _28238_ /*50901*/;
assign _28242_ = _27715_ ^ _28238_ /*50904*/;
assign _28243_ = _28234_ & _28242_ /*50902*/;
assign _28163_ = _28234_ ^ _28242_ /*50903*/;
assign _28240_ = _28241_ | _28243_ /*50900*/;
assign _28245_ = ~Q[32] /*50899*/;
assign _28244_ = _28245_ & D[3] /*50898*/;
assign _28247_ = _27716_ & _28244_ /*50893*/;
assign _28248_ = _27716_ ^ _28244_ /*50896*/;
assign _28249_ = _28240_ & _28248_ /*50894*/;
assign _28164_ = _28240_ ^ _28248_ /*50895*/;
assign _28246_ = _28247_ | _28249_ /*50892*/;
assign _28251_ = ~Q[32] /*50891*/;
assign _28250_ = _28251_ & D[4] /*50890*/;
assign _28253_ = _27717_ & _28250_ /*50885*/;
assign _28254_ = _27717_ ^ _28250_ /*50888*/;
assign _28255_ = _28246_ & _28254_ /*50886*/;
assign _28165_ = _28246_ ^ _28254_ /*50887*/;
assign _28252_ = _28253_ | _28255_ /*50884*/;
assign _28257_ = ~Q[32] /*50883*/;
assign _28256_ = _28257_ & D[5] /*50882*/;
assign _28259_ = _27718_ & _28256_ /*50877*/;
assign _28260_ = _27718_ ^ _28256_ /*50880*/;
assign _28261_ = _28252_ & _28260_ /*50878*/;
assign _28166_ = _28252_ ^ _28260_ /*50879*/;
assign _28258_ = _28259_ | _28261_ /*50876*/;
assign _28263_ = ~Q[32] /*50875*/;
assign _28262_ = _28263_ & D[6] /*50874*/;
assign _28265_ = _27719_ & _28262_ /*50869*/;
assign _28266_ = _27719_ ^ _28262_ /*50872*/;
assign _28267_ = _28258_ & _28266_ /*50870*/;
assign _28167_ = _28258_ ^ _28266_ /*50871*/;
assign _28264_ = _28265_ | _28267_ /*50868*/;
assign _28269_ = ~Q[32] /*50867*/;
assign _28268_ = _28269_ & D[7] /*50866*/;
assign _28271_ = _27720_ & _28268_ /*50861*/;
assign _28272_ = _27720_ ^ _28268_ /*50864*/;
assign _28273_ = _28264_ & _28272_ /*50862*/;
assign _28168_ = _28264_ ^ _28272_ /*50863*/;
assign _28270_ = _28271_ | _28273_ /*50860*/;
assign _28275_ = ~Q[32] /*50859*/;
assign _28274_ = _28275_ & D[8] /*50858*/;
assign _28277_ = _27721_ & _28274_ /*50853*/;
assign _28278_ = _27721_ ^ _28274_ /*50856*/;
assign _28279_ = _28270_ & _28278_ /*50854*/;
assign _28169_ = _28270_ ^ _28278_ /*50855*/;
assign _28276_ = _28277_ | _28279_ /*50852*/;
assign _28281_ = ~Q[32] /*50851*/;
assign _28280_ = _28281_ & D[9] /*50850*/;
assign _28283_ = _27722_ & _28280_ /*50845*/;
assign _28284_ = _27722_ ^ _28280_ /*50848*/;
assign _28285_ = _28276_ & _28284_ /*50846*/;
assign _28170_ = _28276_ ^ _28284_ /*50847*/;
assign _28282_ = _28283_ | _28285_ /*50844*/;
assign _28287_ = ~Q[32] /*50843*/;
assign _28286_ = _28287_ & D[10] /*50842*/;
assign _28289_ = _27723_ & _28286_ /*50837*/;
assign _28290_ = _27723_ ^ _28286_ /*50840*/;
assign _28291_ = _28282_ & _28290_ /*50838*/;
assign _28171_ = _28282_ ^ _28290_ /*50839*/;
assign _28288_ = _28289_ | _28291_ /*50836*/;
assign _28293_ = ~Q[32] /*50835*/;
assign _28292_ = _28293_ & D[11] /*50834*/;
assign _28295_ = _27724_ & _28292_ /*50829*/;
assign _28296_ = _27724_ ^ _28292_ /*50832*/;
assign _28297_ = _28288_ & _28296_ /*50830*/;
assign _28172_ = _28288_ ^ _28296_ /*50831*/;
assign _28294_ = _28295_ | _28297_ /*50828*/;
assign _28299_ = ~Q[32] /*50827*/;
assign _28298_ = _28299_ & D[12] /*50826*/;
assign _28301_ = _27725_ & _28298_ /*50821*/;
assign _28302_ = _27725_ ^ _28298_ /*50824*/;
assign _28303_ = _28294_ & _28302_ /*50822*/;
assign _28173_ = _28294_ ^ _28302_ /*50823*/;
assign _28300_ = _28301_ | _28303_ /*50820*/;
assign _28305_ = ~Q[32] /*50819*/;
assign _28304_ = _28305_ & D[13] /*50818*/;
assign _28307_ = _27726_ & _28304_ /*50813*/;
assign _28308_ = _27726_ ^ _28304_ /*50816*/;
assign _28309_ = _28300_ & _28308_ /*50814*/;
assign _28174_ = _28300_ ^ _28308_ /*50815*/;
assign _28306_ = _28307_ | _28309_ /*50812*/;
assign _28311_ = ~Q[32] /*50811*/;
assign _28310_ = _28311_ & D[14] /*50810*/;
assign _28313_ = _27727_ & _28310_ /*50805*/;
assign _28314_ = _27727_ ^ _28310_ /*50808*/;
assign _28315_ = _28306_ & _28314_ /*50806*/;
assign _28175_ = _28306_ ^ _28314_ /*50807*/;
assign _28312_ = _28313_ | _28315_ /*50804*/;
assign _28317_ = ~Q[32] /*50803*/;
assign _28316_ = _28317_ & D[15] /*50802*/;
assign _28319_ = _27728_ & _28316_ /*50797*/;
assign _28320_ = _27728_ ^ _28316_ /*50800*/;
assign _28321_ = _28312_ & _28320_ /*50798*/;
assign _28176_ = _28312_ ^ _28320_ /*50799*/;
assign _28318_ = _28319_ | _28321_ /*50796*/;
assign _28323_ = ~Q[32] /*50795*/;
assign _28322_ = _28323_ & D[16] /*50794*/;
assign _28325_ = _27729_ & _28322_ /*50789*/;
assign _28326_ = _27729_ ^ _28322_ /*50792*/;
assign _28327_ = _28318_ & _28326_ /*50790*/;
assign _28177_ = _28318_ ^ _28326_ /*50791*/;
assign _28324_ = _28325_ | _28327_ /*50788*/;
assign _28329_ = ~Q[32] /*50787*/;
assign _28328_ = _28329_ & D[17] /*50786*/;
assign _28331_ = _27730_ & _28328_ /*50781*/;
assign _28332_ = _27730_ ^ _28328_ /*50784*/;
assign _28333_ = _28324_ & _28332_ /*50782*/;
assign _28178_ = _28324_ ^ _28332_ /*50783*/;
assign _28330_ = _28331_ | _28333_ /*50780*/;
assign _28335_ = ~Q[32] /*50779*/;
assign _28334_ = _28335_ & D[18] /*50778*/;
assign _28337_ = _27731_ & _28334_ /*50773*/;
assign _28338_ = _27731_ ^ _28334_ /*50776*/;
assign _28339_ = _28330_ & _28338_ /*50774*/;
assign _28179_ = _28330_ ^ _28338_ /*50775*/;
assign _28336_ = _28337_ | _28339_ /*50772*/;
assign _28341_ = ~Q[32] /*50771*/;
assign _28340_ = _28341_ & D[19] /*50770*/;
assign _28343_ = _27732_ & _28340_ /*50765*/;
assign _28344_ = _27732_ ^ _28340_ /*50768*/;
assign _28345_ = _28336_ & _28344_ /*50766*/;
assign _28180_ = _28336_ ^ _28344_ /*50767*/;
assign _28342_ = _28343_ | _28345_ /*50764*/;
assign _28347_ = ~Q[32] /*50763*/;
assign _28346_ = _28347_ & D[20] /*50762*/;
assign _28349_ = _27733_ & _28346_ /*50757*/;
assign _28350_ = _27733_ ^ _28346_ /*50760*/;
assign _28351_ = _28342_ & _28350_ /*50758*/;
assign _28181_ = _28342_ ^ _28350_ /*50759*/;
assign _28348_ = _28349_ | _28351_ /*50756*/;
assign _28353_ = ~Q[32] /*50755*/;
assign _28352_ = _28353_ & D[21] /*50754*/;
assign _28355_ = _27734_ & _28352_ /*50749*/;
assign _28356_ = _27734_ ^ _28352_ /*50752*/;
assign _28357_ = _28348_ & _28356_ /*50750*/;
assign _28182_ = _28348_ ^ _28356_ /*50751*/;
assign _28354_ = _28355_ | _28357_ /*50748*/;
assign _28359_ = ~Q[32] /*50747*/;
assign _28358_ = _28359_ & D[22] /*50746*/;
assign _28361_ = _27735_ & _28358_ /*50741*/;
assign _28362_ = _27735_ ^ _28358_ /*50744*/;
assign _28363_ = _28354_ & _28362_ /*50742*/;
assign _28183_ = _28354_ ^ _28362_ /*50743*/;
assign _28360_ = _28361_ | _28363_ /*50740*/;
assign _28365_ = ~Q[32] /*50739*/;
assign _28364_ = _28365_ & D[23] /*50738*/;
assign _28367_ = _27736_ & _28364_ /*50733*/;
assign _28368_ = _27736_ ^ _28364_ /*50736*/;
assign _28369_ = _28360_ & _28368_ /*50734*/;
assign _28184_ = _28360_ ^ _28368_ /*50735*/;
assign _28366_ = _28367_ | _28369_ /*50732*/;
assign _28371_ = ~Q[32] /*50731*/;
assign _28370_ = _28371_ & D[24] /*50730*/;
assign _28373_ = _27737_ & _28370_ /*50725*/;
assign _28374_ = _27737_ ^ _28370_ /*50728*/;
assign _28375_ = _28366_ & _28374_ /*50726*/;
assign _28185_ = _28366_ ^ _28374_ /*50727*/;
assign _28372_ = _28373_ | _28375_ /*50724*/;
assign _28377_ = ~Q[32] /*50723*/;
assign _28376_ = _28377_ & D[25] /*50722*/;
assign _28379_ = _27738_ & _28376_ /*50717*/;
assign _28380_ = _27738_ ^ _28376_ /*50720*/;
assign _28381_ = _28372_ & _28380_ /*50718*/;
assign _28186_ = _28372_ ^ _28380_ /*50719*/;
assign _28378_ = _28379_ | _28381_ /*50716*/;
assign _28383_ = ~Q[32] /*50715*/;
assign _28382_ = _28383_ & D[26] /*50714*/;
assign _28385_ = _27739_ & _28382_ /*50709*/;
assign _28386_ = _27739_ ^ _28382_ /*50712*/;
assign _28387_ = _28378_ & _28386_ /*50710*/;
assign _28187_ = _28378_ ^ _28386_ /*50711*/;
assign _28384_ = _28385_ | _28387_ /*50708*/;
assign _28389_ = ~Q[32] /*50707*/;
assign _28388_ = _28389_ & D[27] /*50706*/;
assign _28391_ = _27740_ & _28388_ /*50701*/;
assign _28392_ = _27740_ ^ _28388_ /*50704*/;
assign _28393_ = _28384_ & _28392_ /*50702*/;
assign _28188_ = _28384_ ^ _28392_ /*50703*/;
assign _28390_ = _28391_ | _28393_ /*50700*/;
assign _28395_ = ~Q[32] /*50699*/;
assign _28394_ = _28395_ & D[28] /*50698*/;
assign _28397_ = _27741_ & _28394_ /*50693*/;
assign _28398_ = _27741_ ^ _28394_ /*50696*/;
assign _28399_ = _28390_ & _28398_ /*50694*/;
assign _28189_ = _28390_ ^ _28398_ /*50695*/;
assign _28396_ = _28397_ | _28399_ /*50692*/;
assign _28401_ = ~Q[32] /*50691*/;
assign _28400_ = _28401_ & D[29] /*50690*/;
assign _28403_ = _27742_ & _28400_ /*50685*/;
assign _28404_ = _27742_ ^ _28400_ /*50688*/;
assign _28405_ = _28396_ & _28404_ /*50686*/;
assign _28190_ = _28396_ ^ _28404_ /*50687*/;
assign _28402_ = _28403_ | _28405_ /*50684*/;
assign _28407_ = ~Q[32] /*50683*/;
assign _28406_ = _28407_ & D[30] /*50682*/;
assign _28409_ = _27743_ & _28406_ /*50677*/;
assign _28410_ = _27743_ ^ _28406_ /*50680*/;
assign _28411_ = _28402_ & _28410_ /*50678*/;
assign _28191_ = _28402_ ^ _28410_ /*50679*/;
assign _28408_ = _28409_ | _28411_ /*50676*/;
assign _28413_ = ~Q[32] /*50675*/;
assign _28412_ = _28413_ & D[31] /*50674*/;
assign _28415_ = _27744_ & _28412_ /*50669*/;
assign _28416_ = _27744_ ^ _28412_ /*50672*/;
assign _28417_ = _28408_ & _28416_ /*50670*/;
assign _28192_ = _28408_ ^ _28416_ /*50671*/;
assign _28414_ = _28415_ | _28417_ /*50668*/;
assign _28419_ = ~Q[32] /*50667*/;
assign _28418_ = _28419_ & D[32] /*50666*/;
assign _28421_ = _27745_ & _28418_ /*50661*/;
assign _28422_ = _27745_ ^ _28418_ /*50664*/;
assign _28423_ = _28414_ & _28422_ /*50662*/;
assign _28193_ = _28414_ ^ _28422_ /*50663*/;
assign _28420_ = _28421_ | _28423_ /*50660*/;
assign _28425_ = ~Q[32] /*50659*/;
assign _28424_ = _28425_ & D[33] /*50658*/;
assign _28427_ = _27746_ & _28424_ /*50653*/;
assign _28428_ = _27746_ ^ _28424_ /*50656*/;
assign _28429_ = _28420_ & _28428_ /*50654*/;
assign _28194_ = _28420_ ^ _28428_ /*50655*/;
assign _28426_ = _28427_ | _28429_ /*50652*/;
assign _28431_ = ~Q[32] /*50651*/;
assign _28430_ = _28431_ & D[34] /*50650*/;
assign _28433_ = _27747_ & _28430_ /*50645*/;
assign _28434_ = _27747_ ^ _28430_ /*50648*/;
assign _28435_ = _28426_ & _28434_ /*50646*/;
assign _28195_ = _28426_ ^ _28434_ /*50647*/;
assign _28432_ = _28433_ | _28435_ /*50644*/;
assign _28437_ = ~Q[32] /*50643*/;
assign _28436_ = _28437_ & D[35] /*50642*/;
assign _28439_ = _27748_ & _28436_ /*50637*/;
assign _28440_ = _27748_ ^ _28436_ /*50640*/;
assign _28441_ = _28432_ & _28440_ /*50638*/;
assign _28196_ = _28432_ ^ _28440_ /*50639*/;
assign _28438_ = _28439_ | _28441_ /*50636*/;
assign _28443_ = ~Q[32] /*50635*/;
assign _28442_ = _28443_ & D[36] /*50634*/;
assign _28445_ = _27749_ & _28442_ /*50629*/;
assign _28446_ = _27749_ ^ _28442_ /*50632*/;
assign _28447_ = _28438_ & _28446_ /*50630*/;
assign _28197_ = _28438_ ^ _28446_ /*50631*/;
assign _28444_ = _28445_ | _28447_ /*50628*/;
assign _28449_ = ~Q[32] /*50627*/;
assign _28448_ = _28449_ & D[37] /*50626*/;
assign _28451_ = _27750_ & _28448_ /*50621*/;
assign _28452_ = _27750_ ^ _28448_ /*50624*/;
assign _28453_ = _28444_ & _28452_ /*50622*/;
assign _28198_ = _28444_ ^ _28452_ /*50623*/;
assign _28450_ = _28451_ | _28453_ /*50620*/;
assign _28455_ = ~Q[32] /*50619*/;
assign _28454_ = _28455_ & D[38] /*50618*/;
assign _28457_ = _27751_ & _28454_ /*50613*/;
assign _28458_ = _27751_ ^ _28454_ /*50616*/;
assign _28459_ = _28450_ & _28458_ /*50614*/;
assign _28199_ = _28450_ ^ _28458_ /*50615*/;
assign _28456_ = _28457_ | _28459_ /*50612*/;
assign _28461_ = ~Q[32] /*50611*/;
assign _28460_ = _28461_ & D[39] /*50610*/;
assign _28463_ = _27752_ & _28460_ /*50605*/;
assign _28464_ = _27752_ ^ _28460_ /*50608*/;
assign _28465_ = _28456_ & _28464_ /*50606*/;
assign _28200_ = _28456_ ^ _28464_ /*50607*/;
assign _28462_ = _28463_ | _28465_ /*50604*/;
assign _28467_ = ~Q[32] /*50603*/;
assign _28466_ = _28467_ & D[40] /*50602*/;
assign _28469_ = _27753_ & _28466_ /*50597*/;
assign _28470_ = _27753_ ^ _28466_ /*50600*/;
assign _28471_ = _28462_ & _28470_ /*50598*/;
assign _28201_ = _28462_ ^ _28470_ /*50599*/;
assign _28468_ = _28469_ | _28471_ /*50596*/;
assign _28473_ = ~Q[32] /*50595*/;
assign _28472_ = _28473_ & D[41] /*50594*/;
assign _28475_ = _27754_ & _28472_ /*50589*/;
assign _28476_ = _27754_ ^ _28472_ /*50592*/;
assign _28477_ = _28468_ & _28476_ /*50590*/;
assign _28202_ = _28468_ ^ _28476_ /*50591*/;
assign _28474_ = _28475_ | _28477_ /*50588*/;
assign _28479_ = ~Q[32] /*50587*/;
assign _28478_ = _28479_ & D[42] /*50586*/;
assign _28481_ = _27755_ & _28478_ /*50581*/;
assign _28482_ = _27755_ ^ _28478_ /*50584*/;
assign _28483_ = _28474_ & _28482_ /*50582*/;
assign _28203_ = _28474_ ^ _28482_ /*50583*/;
assign _28480_ = _28481_ | _28483_ /*50580*/;
assign _28485_ = ~Q[32] /*50579*/;
assign _28484_ = _28485_ & D[43] /*50578*/;
assign _28487_ = _27756_ & _28484_ /*50573*/;
assign _28488_ = _27756_ ^ _28484_ /*50576*/;
assign _28489_ = _28480_ & _28488_ /*50574*/;
assign _28204_ = _28480_ ^ _28488_ /*50575*/;
assign _28486_ = _28487_ | _28489_ /*50572*/;
assign _28491_ = ~Q[32] /*50571*/;
assign _28490_ = _28491_ & D[44] /*50570*/;
assign _28493_ = _27757_ & _28490_ /*50565*/;
assign _28494_ = _27757_ ^ _28490_ /*50568*/;
assign _28495_ = _28486_ & _28494_ /*50566*/;
assign _28205_ = _28486_ ^ _28494_ /*50567*/;
assign _28492_ = _28493_ | _28495_ /*50564*/;
assign _28497_ = ~Q[32] /*50563*/;
assign _28496_ = _28497_ & D[45] /*50562*/;
assign _28499_ = _27758_ & _28496_ /*50557*/;
assign _28500_ = _27758_ ^ _28496_ /*50560*/;
assign _28501_ = _28492_ & _28500_ /*50558*/;
assign _28206_ = _28492_ ^ _28500_ /*50559*/;
assign _28498_ = _28499_ | _28501_ /*50556*/;
assign _28503_ = ~Q[32] /*50555*/;
assign _28502_ = _28503_ & D[46] /*50554*/;
assign _28505_ = _27759_ & _28502_ /*50549*/;
assign _28506_ = _27759_ ^ _28502_ /*50552*/;
assign _28507_ = _28498_ & _28506_ /*50550*/;
assign _28207_ = _28498_ ^ _28506_ /*50551*/;
assign _28504_ = _28505_ | _28507_ /*50548*/;
assign _28509_ = ~Q[32] /*50547*/;
assign _28508_ = _28509_ & D[47] /*50546*/;
assign _28511_ = _27760_ & _28508_ /*50541*/;
assign _28512_ = _27760_ ^ _28508_ /*50544*/;
assign _28513_ = _28504_ & _28512_ /*50542*/;
assign _28208_ = _28504_ ^ _28512_ /*50543*/;
assign _28510_ = _28511_ | _28513_ /*50540*/;
assign _28515_ = ~Q[32] /*50539*/;
assign _28514_ = _28515_ & D[48] /*50538*/;
assign _28517_ = _27761_ & _28514_ /*50533*/;
assign _28518_ = _27761_ ^ _28514_ /*50536*/;
assign _28519_ = _28510_ & _28518_ /*50534*/;
assign _28209_ = _28510_ ^ _28518_ /*50535*/;
assign _28516_ = _28517_ | _28519_ /*50532*/;
assign _28521_ = ~Q[32] /*50531*/;
assign _28520_ = _28521_ & D[49] /*50530*/;
assign _28523_ = _27762_ & _28520_ /*50525*/;
assign _28524_ = _27762_ ^ _28520_ /*50528*/;
assign _28525_ = _28516_ & _28524_ /*50526*/;
assign _28210_ = _28516_ ^ _28524_ /*50527*/;
assign _28522_ = _28523_ | _28525_ /*50524*/;
assign _28527_ = ~Q[32] /*50523*/;
assign _28526_ = _28527_ & D[50] /*50522*/;
assign _28529_ = _27763_ & _28526_ /*50517*/;
assign _28530_ = _27763_ ^ _28526_ /*50520*/;
assign _28531_ = _28522_ & _28530_ /*50518*/;
assign _28211_ = _28522_ ^ _28530_ /*50519*/;
assign _28528_ = _28529_ | _28531_ /*50516*/;
assign _28533_ = ~Q[32] /*50515*/;
assign _28532_ = _28533_ & D[51] /*50514*/;
assign _28535_ = _27764_ & _28532_ /*50509*/;
assign _28536_ = _27764_ ^ _28532_ /*50512*/;
assign _28537_ = _28528_ & _28536_ /*50510*/;
assign _28212_ = _28528_ ^ _28536_ /*50511*/;
assign _28534_ = _28535_ | _28537_ /*50508*/;
assign _28539_ = ~Q[32] /*50507*/;
assign _28538_ = _28539_ & D[52] /*50506*/;
assign _28541_ = _27765_ & _28538_ /*50501*/;
assign _28542_ = _27765_ ^ _28538_ /*50504*/;
assign _28543_ = _28534_ & _28542_ /*50502*/;
assign _28213_ = _28534_ ^ _28542_ /*50503*/;
assign _28540_ = _28541_ | _28543_ /*50500*/;
assign _28545_ = ~Q[32] /*50499*/;
assign _28544_ = _28545_ & D[53] /*50498*/;
assign _28547_ = _27766_ & _28544_ /*50493*/;
assign _28548_ = _27766_ ^ _28544_ /*50496*/;
assign _28549_ = _28540_ & _28548_ /*50494*/;
assign _28214_ = _28540_ ^ _28548_ /*50495*/;
assign _28546_ = _28547_ | _28549_ /*50492*/;
assign _28551_ = ~Q[32] /*50491*/;
assign _28550_ = _28551_ & D[54] /*50490*/;
assign _28553_ = _27767_ & _28550_ /*50485*/;
assign _28554_ = _27767_ ^ _28550_ /*50488*/;
assign _28555_ = _28546_ & _28554_ /*50486*/;
assign _28215_ = _28546_ ^ _28554_ /*50487*/;
assign _28552_ = _28553_ | _28555_ /*50484*/;
assign _28557_ = ~Q[32] /*50483*/;
assign _28556_ = _28557_ & D[55] /*50482*/;
assign _28559_ = _27768_ & _28556_ /*50477*/;
assign _28560_ = _27768_ ^ _28556_ /*50480*/;
assign _28561_ = _28552_ & _28560_ /*50478*/;
assign _28216_ = _28552_ ^ _28560_ /*50479*/;
assign _28558_ = _28559_ | _28561_ /*50476*/;
assign _28563_ = ~Q[32] /*50475*/;
assign _28562_ = _28563_ & D[56] /*50474*/;
assign _28565_ = _27769_ & _28562_ /*50469*/;
assign _28566_ = _27769_ ^ _28562_ /*50472*/;
assign _28567_ = _28558_ & _28566_ /*50470*/;
assign _28217_ = _28558_ ^ _28566_ /*50471*/;
assign _28564_ = _28565_ | _28567_ /*50468*/;
assign _28569_ = ~Q[32] /*50467*/;
assign _28568_ = _28569_ & D[57] /*50466*/;
assign _28571_ = _27770_ & _28568_ /*50461*/;
assign _28572_ = _27770_ ^ _28568_ /*50464*/;
assign _28573_ = _28564_ & _28572_ /*50462*/;
assign _28218_ = _28564_ ^ _28572_ /*50463*/;
assign _28570_ = _28571_ | _28573_ /*50460*/;
assign _28575_ = ~Q[32] /*50459*/;
assign _28574_ = _28575_ & D[58] /*50458*/;
assign _28577_ = _27771_ & _28574_ /*50453*/;
assign _28578_ = _27771_ ^ _28574_ /*50456*/;
assign _28579_ = _28570_ & _28578_ /*50454*/;
assign _28219_ = _28570_ ^ _28578_ /*50455*/;
assign _28576_ = _28577_ | _28579_ /*50452*/;
assign _28581_ = ~Q[32] /*50451*/;
assign _28580_ = _28581_ & D[59] /*50450*/;
assign _28583_ = _27772_ & _28580_ /*50445*/;
assign _28584_ = _27772_ ^ _28580_ /*50448*/;
assign _28585_ = _28576_ & _28584_ /*50446*/;
assign _28220_ = _28576_ ^ _28584_ /*50447*/;
assign _28582_ = _28583_ | _28585_ /*50444*/;
assign _28587_ = ~Q[32] /*50443*/;
assign _28586_ = _28587_ & D[60] /*50442*/;
assign _28589_ = _27773_ & _28586_ /*50437*/;
assign _28590_ = _27773_ ^ _28586_ /*50440*/;
assign _28591_ = _28582_ & _28590_ /*50438*/;
assign _28221_ = _28582_ ^ _28590_ /*50439*/;
assign _28588_ = _28589_ | _28591_ /*50436*/;
assign _28593_ = ~Q[32] /*50435*/;
assign _28592_ = _28593_ & D[61] /*50434*/;
assign _28595_ = _27774_ & _28592_ /*50429*/;
assign _28596_ = _27774_ ^ _28592_ /*50432*/;
assign _28597_ = _28588_ & _28596_ /*50430*/;
assign _28222_ = _28588_ ^ _28596_ /*50431*/;
assign _28594_ = _28595_ | _28597_ /*50428*/;
assign _28599_ = ~Q[32] /*50427*/;
assign _28598_ = _28599_ & D[62] /*50426*/;
assign _28601_ = _27775_ & _28598_ /*50421*/;
assign _28602_ = _27775_ ^ _28598_ /*50424*/;
assign _28603_ = _28594_ & _28602_ /*50422*/;
assign _28223_ = _28594_ ^ _28602_ /*50423*/;
assign _28600_ = _28601_ | _28603_ /*50420*/;
assign _28605_ = ~Q[32] /*50419*/;
assign _28604_ = _28605_ & zeroWire /*50418*/;
assign _28606_ = _27776_ ^ _28604_ /*50416*/;
assign _28224_ = _28606_ ^ _28600_ /*50415*/;
assign _28677_ = ~D[0] /*50161*/;
assign _28674_ = R_0[31] & _28677_ /*50157*/;
assign _28675_ = R_0[31] ^ _28677_ /*50160*/;
assign _28676_ = oneWire & _28675_ /*50158*/;
assign _28609_ = oneWire ^ _28675_ /*50159*/;
assign _28673_ = _28674_ | _28676_ /*50156*/;
assign _28682_ = ~D[1] /*50155*/;
assign _28679_ = _28161_ & _28682_ /*50151*/;
assign _28680_ = _28161_ ^ _28682_ /*50154*/;
assign _28681_ = _28673_ & _28680_ /*50152*/;
assign _28610_ = _28673_ ^ _28680_ /*50153*/;
assign _28678_ = _28679_ | _28681_ /*50150*/;
assign _28687_ = ~D[2] /*50149*/;
assign _28684_ = _28162_ & _28687_ /*50145*/;
assign _28685_ = _28162_ ^ _28687_ /*50148*/;
assign _28686_ = _28678_ & _28685_ /*50146*/;
assign _28611_ = _28678_ ^ _28685_ /*50147*/;
assign _28683_ = _28684_ | _28686_ /*50144*/;
assign _28692_ = ~D[3] /*50143*/;
assign _28689_ = _28163_ & _28692_ /*50139*/;
assign _28690_ = _28163_ ^ _28692_ /*50142*/;
assign _28691_ = _28683_ & _28690_ /*50140*/;
assign _28612_ = _28683_ ^ _28690_ /*50141*/;
assign _28688_ = _28689_ | _28691_ /*50138*/;
assign _28697_ = ~D[4] /*50137*/;
assign _28694_ = _28164_ & _28697_ /*50133*/;
assign _28695_ = _28164_ ^ _28697_ /*50136*/;
assign _28696_ = _28688_ & _28695_ /*50134*/;
assign _28613_ = _28688_ ^ _28695_ /*50135*/;
assign _28693_ = _28694_ | _28696_ /*50132*/;
assign _28702_ = ~D[5] /*50131*/;
assign _28699_ = _28165_ & _28702_ /*50127*/;
assign _28700_ = _28165_ ^ _28702_ /*50130*/;
assign _28701_ = _28693_ & _28700_ /*50128*/;
assign _28614_ = _28693_ ^ _28700_ /*50129*/;
assign _28698_ = _28699_ | _28701_ /*50126*/;
assign _28707_ = ~D[6] /*50125*/;
assign _28704_ = _28166_ & _28707_ /*50121*/;
assign _28705_ = _28166_ ^ _28707_ /*50124*/;
assign _28706_ = _28698_ & _28705_ /*50122*/;
assign _28615_ = _28698_ ^ _28705_ /*50123*/;
assign _28703_ = _28704_ | _28706_ /*50120*/;
assign _28712_ = ~D[7] /*50119*/;
assign _28709_ = _28167_ & _28712_ /*50115*/;
assign _28710_ = _28167_ ^ _28712_ /*50118*/;
assign _28711_ = _28703_ & _28710_ /*50116*/;
assign _28616_ = _28703_ ^ _28710_ /*50117*/;
assign _28708_ = _28709_ | _28711_ /*50114*/;
assign _28717_ = ~D[8] /*50113*/;
assign _28714_ = _28168_ & _28717_ /*50109*/;
assign _28715_ = _28168_ ^ _28717_ /*50112*/;
assign _28716_ = _28708_ & _28715_ /*50110*/;
assign _28617_ = _28708_ ^ _28715_ /*50111*/;
assign _28713_ = _28714_ | _28716_ /*50108*/;
assign _28722_ = ~D[9] /*50107*/;
assign _28719_ = _28169_ & _28722_ /*50103*/;
assign _28720_ = _28169_ ^ _28722_ /*50106*/;
assign _28721_ = _28713_ & _28720_ /*50104*/;
assign _28618_ = _28713_ ^ _28720_ /*50105*/;
assign _28718_ = _28719_ | _28721_ /*50102*/;
assign _28727_ = ~D[10] /*50101*/;
assign _28724_ = _28170_ & _28727_ /*50097*/;
assign _28725_ = _28170_ ^ _28727_ /*50100*/;
assign _28726_ = _28718_ & _28725_ /*50098*/;
assign _28619_ = _28718_ ^ _28725_ /*50099*/;
assign _28723_ = _28724_ | _28726_ /*50096*/;
assign _28732_ = ~D[11] /*50095*/;
assign _28729_ = _28171_ & _28732_ /*50091*/;
assign _28730_ = _28171_ ^ _28732_ /*50094*/;
assign _28731_ = _28723_ & _28730_ /*50092*/;
assign _28620_ = _28723_ ^ _28730_ /*50093*/;
assign _28728_ = _28729_ | _28731_ /*50090*/;
assign _28737_ = ~D[12] /*50089*/;
assign _28734_ = _28172_ & _28737_ /*50085*/;
assign _28735_ = _28172_ ^ _28737_ /*50088*/;
assign _28736_ = _28728_ & _28735_ /*50086*/;
assign _28621_ = _28728_ ^ _28735_ /*50087*/;
assign _28733_ = _28734_ | _28736_ /*50084*/;
assign _28742_ = ~D[13] /*50083*/;
assign _28739_ = _28173_ & _28742_ /*50079*/;
assign _28740_ = _28173_ ^ _28742_ /*50082*/;
assign _28741_ = _28733_ & _28740_ /*50080*/;
assign _28622_ = _28733_ ^ _28740_ /*50081*/;
assign _28738_ = _28739_ | _28741_ /*50078*/;
assign _28747_ = ~D[14] /*50077*/;
assign _28744_ = _28174_ & _28747_ /*50073*/;
assign _28745_ = _28174_ ^ _28747_ /*50076*/;
assign _28746_ = _28738_ & _28745_ /*50074*/;
assign _28623_ = _28738_ ^ _28745_ /*50075*/;
assign _28743_ = _28744_ | _28746_ /*50072*/;
assign _28752_ = ~D[15] /*50071*/;
assign _28749_ = _28175_ & _28752_ /*50067*/;
assign _28750_ = _28175_ ^ _28752_ /*50070*/;
assign _28751_ = _28743_ & _28750_ /*50068*/;
assign _28624_ = _28743_ ^ _28750_ /*50069*/;
assign _28748_ = _28749_ | _28751_ /*50066*/;
assign _28757_ = ~D[16] /*50065*/;
assign _28754_ = _28176_ & _28757_ /*50061*/;
assign _28755_ = _28176_ ^ _28757_ /*50064*/;
assign _28756_ = _28748_ & _28755_ /*50062*/;
assign _28625_ = _28748_ ^ _28755_ /*50063*/;
assign _28753_ = _28754_ | _28756_ /*50060*/;
assign _28762_ = ~D[17] /*50059*/;
assign _28759_ = _28177_ & _28762_ /*50055*/;
assign _28760_ = _28177_ ^ _28762_ /*50058*/;
assign _28761_ = _28753_ & _28760_ /*50056*/;
assign _28626_ = _28753_ ^ _28760_ /*50057*/;
assign _28758_ = _28759_ | _28761_ /*50054*/;
assign _28767_ = ~D[18] /*50053*/;
assign _28764_ = _28178_ & _28767_ /*50049*/;
assign _28765_ = _28178_ ^ _28767_ /*50052*/;
assign _28766_ = _28758_ & _28765_ /*50050*/;
assign _28627_ = _28758_ ^ _28765_ /*50051*/;
assign _28763_ = _28764_ | _28766_ /*50048*/;
assign _28772_ = ~D[19] /*50047*/;
assign _28769_ = _28179_ & _28772_ /*50043*/;
assign _28770_ = _28179_ ^ _28772_ /*50046*/;
assign _28771_ = _28763_ & _28770_ /*50044*/;
assign _28628_ = _28763_ ^ _28770_ /*50045*/;
assign _28768_ = _28769_ | _28771_ /*50042*/;
assign _28777_ = ~D[20] /*50041*/;
assign _28774_ = _28180_ & _28777_ /*50037*/;
assign _28775_ = _28180_ ^ _28777_ /*50040*/;
assign _28776_ = _28768_ & _28775_ /*50038*/;
assign _28629_ = _28768_ ^ _28775_ /*50039*/;
assign _28773_ = _28774_ | _28776_ /*50036*/;
assign _28782_ = ~D[21] /*50035*/;
assign _28779_ = _28181_ & _28782_ /*50031*/;
assign _28780_ = _28181_ ^ _28782_ /*50034*/;
assign _28781_ = _28773_ & _28780_ /*50032*/;
assign _28630_ = _28773_ ^ _28780_ /*50033*/;
assign _28778_ = _28779_ | _28781_ /*50030*/;
assign _28787_ = ~D[22] /*50029*/;
assign _28784_ = _28182_ & _28787_ /*50025*/;
assign _28785_ = _28182_ ^ _28787_ /*50028*/;
assign _28786_ = _28778_ & _28785_ /*50026*/;
assign _28631_ = _28778_ ^ _28785_ /*50027*/;
assign _28783_ = _28784_ | _28786_ /*50024*/;
assign _28792_ = ~D[23] /*50023*/;
assign _28789_ = _28183_ & _28792_ /*50019*/;
assign _28790_ = _28183_ ^ _28792_ /*50022*/;
assign _28791_ = _28783_ & _28790_ /*50020*/;
assign _28632_ = _28783_ ^ _28790_ /*50021*/;
assign _28788_ = _28789_ | _28791_ /*50018*/;
assign _28797_ = ~D[24] /*50017*/;
assign _28794_ = _28184_ & _28797_ /*50013*/;
assign _28795_ = _28184_ ^ _28797_ /*50016*/;
assign _28796_ = _28788_ & _28795_ /*50014*/;
assign _28633_ = _28788_ ^ _28795_ /*50015*/;
assign _28793_ = _28794_ | _28796_ /*50012*/;
assign _28802_ = ~D[25] /*50011*/;
assign _28799_ = _28185_ & _28802_ /*50007*/;
assign _28800_ = _28185_ ^ _28802_ /*50010*/;
assign _28801_ = _28793_ & _28800_ /*50008*/;
assign _28634_ = _28793_ ^ _28800_ /*50009*/;
assign _28798_ = _28799_ | _28801_ /*50006*/;
assign _28807_ = ~D[26] /*50005*/;
assign _28804_ = _28186_ & _28807_ /*50001*/;
assign _28805_ = _28186_ ^ _28807_ /*50004*/;
assign _28806_ = _28798_ & _28805_ /*50002*/;
assign _28635_ = _28798_ ^ _28805_ /*50003*/;
assign _28803_ = _28804_ | _28806_ /*50000*/;
assign _28812_ = ~D[27] /*49999*/;
assign _28809_ = _28187_ & _28812_ /*49995*/;
assign _28810_ = _28187_ ^ _28812_ /*49998*/;
assign _28811_ = _28803_ & _28810_ /*49996*/;
assign _28636_ = _28803_ ^ _28810_ /*49997*/;
assign _28808_ = _28809_ | _28811_ /*49994*/;
assign _28817_ = ~D[28] /*49993*/;
assign _28814_ = _28188_ & _28817_ /*49989*/;
assign _28815_ = _28188_ ^ _28817_ /*49992*/;
assign _28816_ = _28808_ & _28815_ /*49990*/;
assign _28637_ = _28808_ ^ _28815_ /*49991*/;
assign _28813_ = _28814_ | _28816_ /*49988*/;
assign _28822_ = ~D[29] /*49987*/;
assign _28819_ = _28189_ & _28822_ /*49983*/;
assign _28820_ = _28189_ ^ _28822_ /*49986*/;
assign _28821_ = _28813_ & _28820_ /*49984*/;
assign _28638_ = _28813_ ^ _28820_ /*49985*/;
assign _28818_ = _28819_ | _28821_ /*49982*/;
assign _28827_ = ~D[30] /*49981*/;
assign _28824_ = _28190_ & _28827_ /*49977*/;
assign _28825_ = _28190_ ^ _28827_ /*49980*/;
assign _28826_ = _28818_ & _28825_ /*49978*/;
assign _28639_ = _28818_ ^ _28825_ /*49979*/;
assign _28823_ = _28824_ | _28826_ /*49976*/;
assign _28832_ = ~D[31] /*49975*/;
assign _28829_ = _28191_ & _28832_ /*49971*/;
assign _28830_ = _28191_ ^ _28832_ /*49974*/;
assign _28831_ = _28823_ & _28830_ /*49972*/;
assign _28640_ = _28823_ ^ _28830_ /*49973*/;
assign _28828_ = _28829_ | _28831_ /*49970*/;
assign _28837_ = ~D[32] /*49969*/;
assign _28834_ = _28192_ & _28837_ /*49965*/;
assign _28835_ = _28192_ ^ _28837_ /*49968*/;
assign _28836_ = _28828_ & _28835_ /*49966*/;
assign _28641_ = _28828_ ^ _28835_ /*49967*/;
assign _28833_ = _28834_ | _28836_ /*49964*/;
assign _28842_ = ~D[33] /*49963*/;
assign _28839_ = _28193_ & _28842_ /*49959*/;
assign _28840_ = _28193_ ^ _28842_ /*49962*/;
assign _28841_ = _28833_ & _28840_ /*49960*/;
assign _28642_ = _28833_ ^ _28840_ /*49961*/;
assign _28838_ = _28839_ | _28841_ /*49958*/;
assign _28847_ = ~D[34] /*49957*/;
assign _28844_ = _28194_ & _28847_ /*49953*/;
assign _28845_ = _28194_ ^ _28847_ /*49956*/;
assign _28846_ = _28838_ & _28845_ /*49954*/;
assign _28643_ = _28838_ ^ _28845_ /*49955*/;
assign _28843_ = _28844_ | _28846_ /*49952*/;
assign _28852_ = ~D[35] /*49951*/;
assign _28849_ = _28195_ & _28852_ /*49947*/;
assign _28850_ = _28195_ ^ _28852_ /*49950*/;
assign _28851_ = _28843_ & _28850_ /*49948*/;
assign _28644_ = _28843_ ^ _28850_ /*49949*/;
assign _28848_ = _28849_ | _28851_ /*49946*/;
assign _28857_ = ~D[36] /*49945*/;
assign _28854_ = _28196_ & _28857_ /*49941*/;
assign _28855_ = _28196_ ^ _28857_ /*49944*/;
assign _28856_ = _28848_ & _28855_ /*49942*/;
assign _28645_ = _28848_ ^ _28855_ /*49943*/;
assign _28853_ = _28854_ | _28856_ /*49940*/;
assign _28862_ = ~D[37] /*49939*/;
assign _28859_ = _28197_ & _28862_ /*49935*/;
assign _28860_ = _28197_ ^ _28862_ /*49938*/;
assign _28861_ = _28853_ & _28860_ /*49936*/;
assign _28646_ = _28853_ ^ _28860_ /*49937*/;
assign _28858_ = _28859_ | _28861_ /*49934*/;
assign _28867_ = ~D[38] /*49933*/;
assign _28864_ = _28198_ & _28867_ /*49929*/;
assign _28865_ = _28198_ ^ _28867_ /*49932*/;
assign _28866_ = _28858_ & _28865_ /*49930*/;
assign _28647_ = _28858_ ^ _28865_ /*49931*/;
assign _28863_ = _28864_ | _28866_ /*49928*/;
assign _28872_ = ~D[39] /*49927*/;
assign _28869_ = _28199_ & _28872_ /*49923*/;
assign _28870_ = _28199_ ^ _28872_ /*49926*/;
assign _28871_ = _28863_ & _28870_ /*49924*/;
assign _28648_ = _28863_ ^ _28870_ /*49925*/;
assign _28868_ = _28869_ | _28871_ /*49922*/;
assign _28877_ = ~D[40] /*49921*/;
assign _28874_ = _28200_ & _28877_ /*49917*/;
assign _28875_ = _28200_ ^ _28877_ /*49920*/;
assign _28876_ = _28868_ & _28875_ /*49918*/;
assign _28649_ = _28868_ ^ _28875_ /*49919*/;
assign _28873_ = _28874_ | _28876_ /*49916*/;
assign _28882_ = ~D[41] /*49915*/;
assign _28879_ = _28201_ & _28882_ /*49911*/;
assign _28880_ = _28201_ ^ _28882_ /*49914*/;
assign _28881_ = _28873_ & _28880_ /*49912*/;
assign _28650_ = _28873_ ^ _28880_ /*49913*/;
assign _28878_ = _28879_ | _28881_ /*49910*/;
assign _28887_ = ~D[42] /*49909*/;
assign _28884_ = _28202_ & _28887_ /*49905*/;
assign _28885_ = _28202_ ^ _28887_ /*49908*/;
assign _28886_ = _28878_ & _28885_ /*49906*/;
assign _28651_ = _28878_ ^ _28885_ /*49907*/;
assign _28883_ = _28884_ | _28886_ /*49904*/;
assign _28892_ = ~D[43] /*49903*/;
assign _28889_ = _28203_ & _28892_ /*49899*/;
assign _28890_ = _28203_ ^ _28892_ /*49902*/;
assign _28891_ = _28883_ & _28890_ /*49900*/;
assign _28652_ = _28883_ ^ _28890_ /*49901*/;
assign _28888_ = _28889_ | _28891_ /*49898*/;
assign _28897_ = ~D[44] /*49897*/;
assign _28894_ = _28204_ & _28897_ /*49893*/;
assign _28895_ = _28204_ ^ _28897_ /*49896*/;
assign _28896_ = _28888_ & _28895_ /*49894*/;
assign _28653_ = _28888_ ^ _28895_ /*49895*/;
assign _28893_ = _28894_ | _28896_ /*49892*/;
assign _28902_ = ~D[45] /*49891*/;
assign _28899_ = _28205_ & _28902_ /*49887*/;
assign _28900_ = _28205_ ^ _28902_ /*49890*/;
assign _28901_ = _28893_ & _28900_ /*49888*/;
assign _28654_ = _28893_ ^ _28900_ /*49889*/;
assign _28898_ = _28899_ | _28901_ /*49886*/;
assign _28907_ = ~D[46] /*49885*/;
assign _28904_ = _28206_ & _28907_ /*49881*/;
assign _28905_ = _28206_ ^ _28907_ /*49884*/;
assign _28906_ = _28898_ & _28905_ /*49882*/;
assign _28655_ = _28898_ ^ _28905_ /*49883*/;
assign _28903_ = _28904_ | _28906_ /*49880*/;
assign _28912_ = ~D[47] /*49879*/;
assign _28909_ = _28207_ & _28912_ /*49875*/;
assign _28910_ = _28207_ ^ _28912_ /*49878*/;
assign _28911_ = _28903_ & _28910_ /*49876*/;
assign _28656_ = _28903_ ^ _28910_ /*49877*/;
assign _28908_ = _28909_ | _28911_ /*49874*/;
assign _28917_ = ~D[48] /*49873*/;
assign _28914_ = _28208_ & _28917_ /*49869*/;
assign _28915_ = _28208_ ^ _28917_ /*49872*/;
assign _28916_ = _28908_ & _28915_ /*49870*/;
assign _28657_ = _28908_ ^ _28915_ /*49871*/;
assign _28913_ = _28914_ | _28916_ /*49868*/;
assign _28922_ = ~D[49] /*49867*/;
assign _28919_ = _28209_ & _28922_ /*49863*/;
assign _28920_ = _28209_ ^ _28922_ /*49866*/;
assign _28921_ = _28913_ & _28920_ /*49864*/;
assign _28658_ = _28913_ ^ _28920_ /*49865*/;
assign _28918_ = _28919_ | _28921_ /*49862*/;
assign _28927_ = ~D[50] /*49861*/;
assign _28924_ = _28210_ & _28927_ /*49857*/;
assign _28925_ = _28210_ ^ _28927_ /*49860*/;
assign _28926_ = _28918_ & _28925_ /*49858*/;
assign _28659_ = _28918_ ^ _28925_ /*49859*/;
assign _28923_ = _28924_ | _28926_ /*49856*/;
assign _28932_ = ~D[51] /*49855*/;
assign _28929_ = _28211_ & _28932_ /*49851*/;
assign _28930_ = _28211_ ^ _28932_ /*49854*/;
assign _28931_ = _28923_ & _28930_ /*49852*/;
assign _28660_ = _28923_ ^ _28930_ /*49853*/;
assign _28928_ = _28929_ | _28931_ /*49850*/;
assign _28937_ = ~D[52] /*49849*/;
assign _28934_ = _28212_ & _28937_ /*49845*/;
assign _28935_ = _28212_ ^ _28937_ /*49848*/;
assign _28936_ = _28928_ & _28935_ /*49846*/;
assign _28661_ = _28928_ ^ _28935_ /*49847*/;
assign _28933_ = _28934_ | _28936_ /*49844*/;
assign _28942_ = ~D[53] /*49843*/;
assign _28939_ = _28213_ & _28942_ /*49839*/;
assign _28940_ = _28213_ ^ _28942_ /*49842*/;
assign _28941_ = _28933_ & _28940_ /*49840*/;
assign _28662_ = _28933_ ^ _28940_ /*49841*/;
assign _28938_ = _28939_ | _28941_ /*49838*/;
assign _28947_ = ~D[54] /*49837*/;
assign _28944_ = _28214_ & _28947_ /*49833*/;
assign _28945_ = _28214_ ^ _28947_ /*49836*/;
assign _28946_ = _28938_ & _28945_ /*49834*/;
assign _28663_ = _28938_ ^ _28945_ /*49835*/;
assign _28943_ = _28944_ | _28946_ /*49832*/;
assign _28952_ = ~D[55] /*49831*/;
assign _28949_ = _28215_ & _28952_ /*49827*/;
assign _28950_ = _28215_ ^ _28952_ /*49830*/;
assign _28951_ = _28943_ & _28950_ /*49828*/;
assign _28664_ = _28943_ ^ _28950_ /*49829*/;
assign _28948_ = _28949_ | _28951_ /*49826*/;
assign _28957_ = ~D[56] /*49825*/;
assign _28954_ = _28216_ & _28957_ /*49821*/;
assign _28955_ = _28216_ ^ _28957_ /*49824*/;
assign _28956_ = _28948_ & _28955_ /*49822*/;
assign _28665_ = _28948_ ^ _28955_ /*49823*/;
assign _28953_ = _28954_ | _28956_ /*49820*/;
assign _28962_ = ~D[57] /*49819*/;
assign _28959_ = _28217_ & _28962_ /*49815*/;
assign _28960_ = _28217_ ^ _28962_ /*49818*/;
assign _28961_ = _28953_ & _28960_ /*49816*/;
assign _28666_ = _28953_ ^ _28960_ /*49817*/;
assign _28958_ = _28959_ | _28961_ /*49814*/;
assign _28967_ = ~D[58] /*49813*/;
assign _28964_ = _28218_ & _28967_ /*49809*/;
assign _28965_ = _28218_ ^ _28967_ /*49812*/;
assign _28966_ = _28958_ & _28965_ /*49810*/;
assign _28667_ = _28958_ ^ _28965_ /*49811*/;
assign _28963_ = _28964_ | _28966_ /*49808*/;
assign _28972_ = ~D[59] /*49807*/;
assign _28969_ = _28219_ & _28972_ /*49803*/;
assign _28970_ = _28219_ ^ _28972_ /*49806*/;
assign _28971_ = _28963_ & _28970_ /*49804*/;
assign _28668_ = _28963_ ^ _28970_ /*49805*/;
assign _28968_ = _28969_ | _28971_ /*49802*/;
assign _28977_ = ~D[60] /*49801*/;
assign _28974_ = _28220_ & _28977_ /*49797*/;
assign _28975_ = _28220_ ^ _28977_ /*49800*/;
assign _28976_ = _28968_ & _28975_ /*49798*/;
assign _28669_ = _28968_ ^ _28975_ /*49799*/;
assign _28973_ = _28974_ | _28976_ /*49796*/;
assign _28982_ = ~D[61] /*49795*/;
assign _28979_ = _28221_ & _28982_ /*49791*/;
assign _28980_ = _28221_ ^ _28982_ /*49794*/;
assign _28981_ = _28973_ & _28980_ /*49792*/;
assign _28670_ = _28973_ ^ _28980_ /*49793*/;
assign _28978_ = _28979_ | _28981_ /*49790*/;
assign _28987_ = ~D[62] /*49789*/;
assign _28984_ = _28222_ & _28987_ /*49785*/;
assign _28985_ = _28222_ ^ _28987_ /*49788*/;
assign _28986_ = _28978_ & _28985_ /*49786*/;
assign _28671_ = _28978_ ^ _28985_ /*49787*/;
assign _28983_ = _28984_ | _28986_ /*49784*/;
assign _28988_ = _28223_ & oneWire /*49779*/;
assign _28989_ = _28223_ ^ oneWire /*49782*/;
assign _28990_ = _28983_ & _28989_ /*49780*/;
assign _28672_ = _28983_ ^ _28989_ /*49781*/;
assign Q[31] = _28988_ | _28990_ /*49778*/;
assign _29123_ = ~Q[31] /*49393*/;
assign _29122_ = _29123_ & D[0] /*49392*/;
assign _29125_ = _28609_ & _29122_ /*49387*/;
assign _29126_ = _28609_ ^ _29122_ /*49390*/;
assign _29127_ = zeroWire & _29126_ /*49388*/;
assign _29057_ = zeroWire ^ _29126_ /*49389*/;
assign _29124_ = _29125_ | _29127_ /*49386*/;
assign _29129_ = ~Q[31] /*49385*/;
assign _29128_ = _29129_ & D[1] /*49384*/;
assign _29131_ = _28610_ & _29128_ /*49379*/;
assign _29132_ = _28610_ ^ _29128_ /*49382*/;
assign _29133_ = _29124_ & _29132_ /*49380*/;
assign _29058_ = _29124_ ^ _29132_ /*49381*/;
assign _29130_ = _29131_ | _29133_ /*49378*/;
assign _29135_ = ~Q[31] /*49377*/;
assign _29134_ = _29135_ & D[2] /*49376*/;
assign _29137_ = _28611_ & _29134_ /*49371*/;
assign _29138_ = _28611_ ^ _29134_ /*49374*/;
assign _29139_ = _29130_ & _29138_ /*49372*/;
assign _29059_ = _29130_ ^ _29138_ /*49373*/;
assign _29136_ = _29137_ | _29139_ /*49370*/;
assign _29141_ = ~Q[31] /*49369*/;
assign _29140_ = _29141_ & D[3] /*49368*/;
assign _29143_ = _28612_ & _29140_ /*49363*/;
assign _29144_ = _28612_ ^ _29140_ /*49366*/;
assign _29145_ = _29136_ & _29144_ /*49364*/;
assign _29060_ = _29136_ ^ _29144_ /*49365*/;
assign _29142_ = _29143_ | _29145_ /*49362*/;
assign _29147_ = ~Q[31] /*49361*/;
assign _29146_ = _29147_ & D[4] /*49360*/;
assign _29149_ = _28613_ & _29146_ /*49355*/;
assign _29150_ = _28613_ ^ _29146_ /*49358*/;
assign _29151_ = _29142_ & _29150_ /*49356*/;
assign _29061_ = _29142_ ^ _29150_ /*49357*/;
assign _29148_ = _29149_ | _29151_ /*49354*/;
assign _29153_ = ~Q[31] /*49353*/;
assign _29152_ = _29153_ & D[5] /*49352*/;
assign _29155_ = _28614_ & _29152_ /*49347*/;
assign _29156_ = _28614_ ^ _29152_ /*49350*/;
assign _29157_ = _29148_ & _29156_ /*49348*/;
assign _29062_ = _29148_ ^ _29156_ /*49349*/;
assign _29154_ = _29155_ | _29157_ /*49346*/;
assign _29159_ = ~Q[31] /*49345*/;
assign _29158_ = _29159_ & D[6] /*49344*/;
assign _29161_ = _28615_ & _29158_ /*49339*/;
assign _29162_ = _28615_ ^ _29158_ /*49342*/;
assign _29163_ = _29154_ & _29162_ /*49340*/;
assign _29063_ = _29154_ ^ _29162_ /*49341*/;
assign _29160_ = _29161_ | _29163_ /*49338*/;
assign _29165_ = ~Q[31] /*49337*/;
assign _29164_ = _29165_ & D[7] /*49336*/;
assign _29167_ = _28616_ & _29164_ /*49331*/;
assign _29168_ = _28616_ ^ _29164_ /*49334*/;
assign _29169_ = _29160_ & _29168_ /*49332*/;
assign _29064_ = _29160_ ^ _29168_ /*49333*/;
assign _29166_ = _29167_ | _29169_ /*49330*/;
assign _29171_ = ~Q[31] /*49329*/;
assign _29170_ = _29171_ & D[8] /*49328*/;
assign _29173_ = _28617_ & _29170_ /*49323*/;
assign _29174_ = _28617_ ^ _29170_ /*49326*/;
assign _29175_ = _29166_ & _29174_ /*49324*/;
assign _29065_ = _29166_ ^ _29174_ /*49325*/;
assign _29172_ = _29173_ | _29175_ /*49322*/;
assign _29177_ = ~Q[31] /*49321*/;
assign _29176_ = _29177_ & D[9] /*49320*/;
assign _29179_ = _28618_ & _29176_ /*49315*/;
assign _29180_ = _28618_ ^ _29176_ /*49318*/;
assign _29181_ = _29172_ & _29180_ /*49316*/;
assign _29066_ = _29172_ ^ _29180_ /*49317*/;
assign _29178_ = _29179_ | _29181_ /*49314*/;
assign _29183_ = ~Q[31] /*49313*/;
assign _29182_ = _29183_ & D[10] /*49312*/;
assign _29185_ = _28619_ & _29182_ /*49307*/;
assign _29186_ = _28619_ ^ _29182_ /*49310*/;
assign _29187_ = _29178_ & _29186_ /*49308*/;
assign _29067_ = _29178_ ^ _29186_ /*49309*/;
assign _29184_ = _29185_ | _29187_ /*49306*/;
assign _29189_ = ~Q[31] /*49305*/;
assign _29188_ = _29189_ & D[11] /*49304*/;
assign _29191_ = _28620_ & _29188_ /*49299*/;
assign _29192_ = _28620_ ^ _29188_ /*49302*/;
assign _29193_ = _29184_ & _29192_ /*49300*/;
assign _29068_ = _29184_ ^ _29192_ /*49301*/;
assign _29190_ = _29191_ | _29193_ /*49298*/;
assign _29195_ = ~Q[31] /*49297*/;
assign _29194_ = _29195_ & D[12] /*49296*/;
assign _29197_ = _28621_ & _29194_ /*49291*/;
assign _29198_ = _28621_ ^ _29194_ /*49294*/;
assign _29199_ = _29190_ & _29198_ /*49292*/;
assign _29069_ = _29190_ ^ _29198_ /*49293*/;
assign _29196_ = _29197_ | _29199_ /*49290*/;
assign _29201_ = ~Q[31] /*49289*/;
assign _29200_ = _29201_ & D[13] /*49288*/;
assign _29203_ = _28622_ & _29200_ /*49283*/;
assign _29204_ = _28622_ ^ _29200_ /*49286*/;
assign _29205_ = _29196_ & _29204_ /*49284*/;
assign _29070_ = _29196_ ^ _29204_ /*49285*/;
assign _29202_ = _29203_ | _29205_ /*49282*/;
assign _29207_ = ~Q[31] /*49281*/;
assign _29206_ = _29207_ & D[14] /*49280*/;
assign _29209_ = _28623_ & _29206_ /*49275*/;
assign _29210_ = _28623_ ^ _29206_ /*49278*/;
assign _29211_ = _29202_ & _29210_ /*49276*/;
assign _29071_ = _29202_ ^ _29210_ /*49277*/;
assign _29208_ = _29209_ | _29211_ /*49274*/;
assign _29213_ = ~Q[31] /*49273*/;
assign _29212_ = _29213_ & D[15] /*49272*/;
assign _29215_ = _28624_ & _29212_ /*49267*/;
assign _29216_ = _28624_ ^ _29212_ /*49270*/;
assign _29217_ = _29208_ & _29216_ /*49268*/;
assign _29072_ = _29208_ ^ _29216_ /*49269*/;
assign _29214_ = _29215_ | _29217_ /*49266*/;
assign _29219_ = ~Q[31] /*49265*/;
assign _29218_ = _29219_ & D[16] /*49264*/;
assign _29221_ = _28625_ & _29218_ /*49259*/;
assign _29222_ = _28625_ ^ _29218_ /*49262*/;
assign _29223_ = _29214_ & _29222_ /*49260*/;
assign _29073_ = _29214_ ^ _29222_ /*49261*/;
assign _29220_ = _29221_ | _29223_ /*49258*/;
assign _29225_ = ~Q[31] /*49257*/;
assign _29224_ = _29225_ & D[17] /*49256*/;
assign _29227_ = _28626_ & _29224_ /*49251*/;
assign _29228_ = _28626_ ^ _29224_ /*49254*/;
assign _29229_ = _29220_ & _29228_ /*49252*/;
assign _29074_ = _29220_ ^ _29228_ /*49253*/;
assign _29226_ = _29227_ | _29229_ /*49250*/;
assign _29231_ = ~Q[31] /*49249*/;
assign _29230_ = _29231_ & D[18] /*49248*/;
assign _29233_ = _28627_ & _29230_ /*49243*/;
assign _29234_ = _28627_ ^ _29230_ /*49246*/;
assign _29235_ = _29226_ & _29234_ /*49244*/;
assign _29075_ = _29226_ ^ _29234_ /*49245*/;
assign _29232_ = _29233_ | _29235_ /*49242*/;
assign _29237_ = ~Q[31] /*49241*/;
assign _29236_ = _29237_ & D[19] /*49240*/;
assign _29239_ = _28628_ & _29236_ /*49235*/;
assign _29240_ = _28628_ ^ _29236_ /*49238*/;
assign _29241_ = _29232_ & _29240_ /*49236*/;
assign _29076_ = _29232_ ^ _29240_ /*49237*/;
assign _29238_ = _29239_ | _29241_ /*49234*/;
assign _29243_ = ~Q[31] /*49233*/;
assign _29242_ = _29243_ & D[20] /*49232*/;
assign _29245_ = _28629_ & _29242_ /*49227*/;
assign _29246_ = _28629_ ^ _29242_ /*49230*/;
assign _29247_ = _29238_ & _29246_ /*49228*/;
assign _29077_ = _29238_ ^ _29246_ /*49229*/;
assign _29244_ = _29245_ | _29247_ /*49226*/;
assign _29249_ = ~Q[31] /*49225*/;
assign _29248_ = _29249_ & D[21] /*49224*/;
assign _29251_ = _28630_ & _29248_ /*49219*/;
assign _29252_ = _28630_ ^ _29248_ /*49222*/;
assign _29253_ = _29244_ & _29252_ /*49220*/;
assign _29078_ = _29244_ ^ _29252_ /*49221*/;
assign _29250_ = _29251_ | _29253_ /*49218*/;
assign _29255_ = ~Q[31] /*49217*/;
assign _29254_ = _29255_ & D[22] /*49216*/;
assign _29257_ = _28631_ & _29254_ /*49211*/;
assign _29258_ = _28631_ ^ _29254_ /*49214*/;
assign _29259_ = _29250_ & _29258_ /*49212*/;
assign _29079_ = _29250_ ^ _29258_ /*49213*/;
assign _29256_ = _29257_ | _29259_ /*49210*/;
assign _29261_ = ~Q[31] /*49209*/;
assign _29260_ = _29261_ & D[23] /*49208*/;
assign _29263_ = _28632_ & _29260_ /*49203*/;
assign _29264_ = _28632_ ^ _29260_ /*49206*/;
assign _29265_ = _29256_ & _29264_ /*49204*/;
assign _29080_ = _29256_ ^ _29264_ /*49205*/;
assign _29262_ = _29263_ | _29265_ /*49202*/;
assign _29267_ = ~Q[31] /*49201*/;
assign _29266_ = _29267_ & D[24] /*49200*/;
assign _29269_ = _28633_ & _29266_ /*49195*/;
assign _29270_ = _28633_ ^ _29266_ /*49198*/;
assign _29271_ = _29262_ & _29270_ /*49196*/;
assign _29081_ = _29262_ ^ _29270_ /*49197*/;
assign _29268_ = _29269_ | _29271_ /*49194*/;
assign _29273_ = ~Q[31] /*49193*/;
assign _29272_ = _29273_ & D[25] /*49192*/;
assign _29275_ = _28634_ & _29272_ /*49187*/;
assign _29276_ = _28634_ ^ _29272_ /*49190*/;
assign _29277_ = _29268_ & _29276_ /*49188*/;
assign _29082_ = _29268_ ^ _29276_ /*49189*/;
assign _29274_ = _29275_ | _29277_ /*49186*/;
assign _29279_ = ~Q[31] /*49185*/;
assign _29278_ = _29279_ & D[26] /*49184*/;
assign _29281_ = _28635_ & _29278_ /*49179*/;
assign _29282_ = _28635_ ^ _29278_ /*49182*/;
assign _29283_ = _29274_ & _29282_ /*49180*/;
assign _29083_ = _29274_ ^ _29282_ /*49181*/;
assign _29280_ = _29281_ | _29283_ /*49178*/;
assign _29285_ = ~Q[31] /*49177*/;
assign _29284_ = _29285_ & D[27] /*49176*/;
assign _29287_ = _28636_ & _29284_ /*49171*/;
assign _29288_ = _28636_ ^ _29284_ /*49174*/;
assign _29289_ = _29280_ & _29288_ /*49172*/;
assign _29084_ = _29280_ ^ _29288_ /*49173*/;
assign _29286_ = _29287_ | _29289_ /*49170*/;
assign _29291_ = ~Q[31] /*49169*/;
assign _29290_ = _29291_ & D[28] /*49168*/;
assign _29293_ = _28637_ & _29290_ /*49163*/;
assign _29294_ = _28637_ ^ _29290_ /*49166*/;
assign _29295_ = _29286_ & _29294_ /*49164*/;
assign _29085_ = _29286_ ^ _29294_ /*49165*/;
assign _29292_ = _29293_ | _29295_ /*49162*/;
assign _29297_ = ~Q[31] /*49161*/;
assign _29296_ = _29297_ & D[29] /*49160*/;
assign _29299_ = _28638_ & _29296_ /*49155*/;
assign _29300_ = _28638_ ^ _29296_ /*49158*/;
assign _29301_ = _29292_ & _29300_ /*49156*/;
assign _29086_ = _29292_ ^ _29300_ /*49157*/;
assign _29298_ = _29299_ | _29301_ /*49154*/;
assign _29303_ = ~Q[31] /*49153*/;
assign _29302_ = _29303_ & D[30] /*49152*/;
assign _29305_ = _28639_ & _29302_ /*49147*/;
assign _29306_ = _28639_ ^ _29302_ /*49150*/;
assign _29307_ = _29298_ & _29306_ /*49148*/;
assign _29087_ = _29298_ ^ _29306_ /*49149*/;
assign _29304_ = _29305_ | _29307_ /*49146*/;
assign _29309_ = ~Q[31] /*49145*/;
assign _29308_ = _29309_ & D[31] /*49144*/;
assign _29311_ = _28640_ & _29308_ /*49139*/;
assign _29312_ = _28640_ ^ _29308_ /*49142*/;
assign _29313_ = _29304_ & _29312_ /*49140*/;
assign _29088_ = _29304_ ^ _29312_ /*49141*/;
assign _29310_ = _29311_ | _29313_ /*49138*/;
assign _29315_ = ~Q[31] /*49137*/;
assign _29314_ = _29315_ & D[32] /*49136*/;
assign _29317_ = _28641_ & _29314_ /*49131*/;
assign _29318_ = _28641_ ^ _29314_ /*49134*/;
assign _29319_ = _29310_ & _29318_ /*49132*/;
assign _29089_ = _29310_ ^ _29318_ /*49133*/;
assign _29316_ = _29317_ | _29319_ /*49130*/;
assign _29321_ = ~Q[31] /*49129*/;
assign _29320_ = _29321_ & D[33] /*49128*/;
assign _29323_ = _28642_ & _29320_ /*49123*/;
assign _29324_ = _28642_ ^ _29320_ /*49126*/;
assign _29325_ = _29316_ & _29324_ /*49124*/;
assign _29090_ = _29316_ ^ _29324_ /*49125*/;
assign _29322_ = _29323_ | _29325_ /*49122*/;
assign _29327_ = ~Q[31] /*49121*/;
assign _29326_ = _29327_ & D[34] /*49120*/;
assign _29329_ = _28643_ & _29326_ /*49115*/;
assign _29330_ = _28643_ ^ _29326_ /*49118*/;
assign _29331_ = _29322_ & _29330_ /*49116*/;
assign _29091_ = _29322_ ^ _29330_ /*49117*/;
assign _29328_ = _29329_ | _29331_ /*49114*/;
assign _29333_ = ~Q[31] /*49113*/;
assign _29332_ = _29333_ & D[35] /*49112*/;
assign _29335_ = _28644_ & _29332_ /*49107*/;
assign _29336_ = _28644_ ^ _29332_ /*49110*/;
assign _29337_ = _29328_ & _29336_ /*49108*/;
assign _29092_ = _29328_ ^ _29336_ /*49109*/;
assign _29334_ = _29335_ | _29337_ /*49106*/;
assign _29339_ = ~Q[31] /*49105*/;
assign _29338_ = _29339_ & D[36] /*49104*/;
assign _29341_ = _28645_ & _29338_ /*49099*/;
assign _29342_ = _28645_ ^ _29338_ /*49102*/;
assign _29343_ = _29334_ & _29342_ /*49100*/;
assign _29093_ = _29334_ ^ _29342_ /*49101*/;
assign _29340_ = _29341_ | _29343_ /*49098*/;
assign _29345_ = ~Q[31] /*49097*/;
assign _29344_ = _29345_ & D[37] /*49096*/;
assign _29347_ = _28646_ & _29344_ /*49091*/;
assign _29348_ = _28646_ ^ _29344_ /*49094*/;
assign _29349_ = _29340_ & _29348_ /*49092*/;
assign _29094_ = _29340_ ^ _29348_ /*49093*/;
assign _29346_ = _29347_ | _29349_ /*49090*/;
assign _29351_ = ~Q[31] /*49089*/;
assign _29350_ = _29351_ & D[38] /*49088*/;
assign _29353_ = _28647_ & _29350_ /*49083*/;
assign _29354_ = _28647_ ^ _29350_ /*49086*/;
assign _29355_ = _29346_ & _29354_ /*49084*/;
assign _29095_ = _29346_ ^ _29354_ /*49085*/;
assign _29352_ = _29353_ | _29355_ /*49082*/;
assign _29357_ = ~Q[31] /*49081*/;
assign _29356_ = _29357_ & D[39] /*49080*/;
assign _29359_ = _28648_ & _29356_ /*49075*/;
assign _29360_ = _28648_ ^ _29356_ /*49078*/;
assign _29361_ = _29352_ & _29360_ /*49076*/;
assign _29096_ = _29352_ ^ _29360_ /*49077*/;
assign _29358_ = _29359_ | _29361_ /*49074*/;
assign _29363_ = ~Q[31] /*49073*/;
assign _29362_ = _29363_ & D[40] /*49072*/;
assign _29365_ = _28649_ & _29362_ /*49067*/;
assign _29366_ = _28649_ ^ _29362_ /*49070*/;
assign _29367_ = _29358_ & _29366_ /*49068*/;
assign _29097_ = _29358_ ^ _29366_ /*49069*/;
assign _29364_ = _29365_ | _29367_ /*49066*/;
assign _29369_ = ~Q[31] /*49065*/;
assign _29368_ = _29369_ & D[41] /*49064*/;
assign _29371_ = _28650_ & _29368_ /*49059*/;
assign _29372_ = _28650_ ^ _29368_ /*49062*/;
assign _29373_ = _29364_ & _29372_ /*49060*/;
assign _29098_ = _29364_ ^ _29372_ /*49061*/;
assign _29370_ = _29371_ | _29373_ /*49058*/;
assign _29375_ = ~Q[31] /*49057*/;
assign _29374_ = _29375_ & D[42] /*49056*/;
assign _29377_ = _28651_ & _29374_ /*49051*/;
assign _29378_ = _28651_ ^ _29374_ /*49054*/;
assign _29379_ = _29370_ & _29378_ /*49052*/;
assign _29099_ = _29370_ ^ _29378_ /*49053*/;
assign _29376_ = _29377_ | _29379_ /*49050*/;
assign _29381_ = ~Q[31] /*49049*/;
assign _29380_ = _29381_ & D[43] /*49048*/;
assign _29383_ = _28652_ & _29380_ /*49043*/;
assign _29384_ = _28652_ ^ _29380_ /*49046*/;
assign _29385_ = _29376_ & _29384_ /*49044*/;
assign _29100_ = _29376_ ^ _29384_ /*49045*/;
assign _29382_ = _29383_ | _29385_ /*49042*/;
assign _29387_ = ~Q[31] /*49041*/;
assign _29386_ = _29387_ & D[44] /*49040*/;
assign _29389_ = _28653_ & _29386_ /*49035*/;
assign _29390_ = _28653_ ^ _29386_ /*49038*/;
assign _29391_ = _29382_ & _29390_ /*49036*/;
assign _29101_ = _29382_ ^ _29390_ /*49037*/;
assign _29388_ = _29389_ | _29391_ /*49034*/;
assign _29393_ = ~Q[31] /*49033*/;
assign _29392_ = _29393_ & D[45] /*49032*/;
assign _29395_ = _28654_ & _29392_ /*49027*/;
assign _29396_ = _28654_ ^ _29392_ /*49030*/;
assign _29397_ = _29388_ & _29396_ /*49028*/;
assign _29102_ = _29388_ ^ _29396_ /*49029*/;
assign _29394_ = _29395_ | _29397_ /*49026*/;
assign _29399_ = ~Q[31] /*49025*/;
assign _29398_ = _29399_ & D[46] /*49024*/;
assign _29401_ = _28655_ & _29398_ /*49019*/;
assign _29402_ = _28655_ ^ _29398_ /*49022*/;
assign _29403_ = _29394_ & _29402_ /*49020*/;
assign _29103_ = _29394_ ^ _29402_ /*49021*/;
assign _29400_ = _29401_ | _29403_ /*49018*/;
assign _29405_ = ~Q[31] /*49017*/;
assign _29404_ = _29405_ & D[47] /*49016*/;
assign _29407_ = _28656_ & _29404_ /*49011*/;
assign _29408_ = _28656_ ^ _29404_ /*49014*/;
assign _29409_ = _29400_ & _29408_ /*49012*/;
assign _29104_ = _29400_ ^ _29408_ /*49013*/;
assign _29406_ = _29407_ | _29409_ /*49010*/;
assign _29411_ = ~Q[31] /*49009*/;
assign _29410_ = _29411_ & D[48] /*49008*/;
assign _29413_ = _28657_ & _29410_ /*49003*/;
assign _29414_ = _28657_ ^ _29410_ /*49006*/;
assign _29415_ = _29406_ & _29414_ /*49004*/;
assign _29105_ = _29406_ ^ _29414_ /*49005*/;
assign _29412_ = _29413_ | _29415_ /*49002*/;
assign _29417_ = ~Q[31] /*49001*/;
assign _29416_ = _29417_ & D[49] /*49000*/;
assign _29419_ = _28658_ & _29416_ /*48995*/;
assign _29420_ = _28658_ ^ _29416_ /*48998*/;
assign _29421_ = _29412_ & _29420_ /*48996*/;
assign _29106_ = _29412_ ^ _29420_ /*48997*/;
assign _29418_ = _29419_ | _29421_ /*48994*/;
assign _29423_ = ~Q[31] /*48993*/;
assign _29422_ = _29423_ & D[50] /*48992*/;
assign _29425_ = _28659_ & _29422_ /*48987*/;
assign _29426_ = _28659_ ^ _29422_ /*48990*/;
assign _29427_ = _29418_ & _29426_ /*48988*/;
assign _29107_ = _29418_ ^ _29426_ /*48989*/;
assign _29424_ = _29425_ | _29427_ /*48986*/;
assign _29429_ = ~Q[31] /*48985*/;
assign _29428_ = _29429_ & D[51] /*48984*/;
assign _29431_ = _28660_ & _29428_ /*48979*/;
assign _29432_ = _28660_ ^ _29428_ /*48982*/;
assign _29433_ = _29424_ & _29432_ /*48980*/;
assign _29108_ = _29424_ ^ _29432_ /*48981*/;
assign _29430_ = _29431_ | _29433_ /*48978*/;
assign _29435_ = ~Q[31] /*48977*/;
assign _29434_ = _29435_ & D[52] /*48976*/;
assign _29437_ = _28661_ & _29434_ /*48971*/;
assign _29438_ = _28661_ ^ _29434_ /*48974*/;
assign _29439_ = _29430_ & _29438_ /*48972*/;
assign _29109_ = _29430_ ^ _29438_ /*48973*/;
assign _29436_ = _29437_ | _29439_ /*48970*/;
assign _29441_ = ~Q[31] /*48969*/;
assign _29440_ = _29441_ & D[53] /*48968*/;
assign _29443_ = _28662_ & _29440_ /*48963*/;
assign _29444_ = _28662_ ^ _29440_ /*48966*/;
assign _29445_ = _29436_ & _29444_ /*48964*/;
assign _29110_ = _29436_ ^ _29444_ /*48965*/;
assign _29442_ = _29443_ | _29445_ /*48962*/;
assign _29447_ = ~Q[31] /*48961*/;
assign _29446_ = _29447_ & D[54] /*48960*/;
assign _29449_ = _28663_ & _29446_ /*48955*/;
assign _29450_ = _28663_ ^ _29446_ /*48958*/;
assign _29451_ = _29442_ & _29450_ /*48956*/;
assign _29111_ = _29442_ ^ _29450_ /*48957*/;
assign _29448_ = _29449_ | _29451_ /*48954*/;
assign _29453_ = ~Q[31] /*48953*/;
assign _29452_ = _29453_ & D[55] /*48952*/;
assign _29455_ = _28664_ & _29452_ /*48947*/;
assign _29456_ = _28664_ ^ _29452_ /*48950*/;
assign _29457_ = _29448_ & _29456_ /*48948*/;
assign _29112_ = _29448_ ^ _29456_ /*48949*/;
assign _29454_ = _29455_ | _29457_ /*48946*/;
assign _29459_ = ~Q[31] /*48945*/;
assign _29458_ = _29459_ & D[56] /*48944*/;
assign _29461_ = _28665_ & _29458_ /*48939*/;
assign _29462_ = _28665_ ^ _29458_ /*48942*/;
assign _29463_ = _29454_ & _29462_ /*48940*/;
assign _29113_ = _29454_ ^ _29462_ /*48941*/;
assign _29460_ = _29461_ | _29463_ /*48938*/;
assign _29465_ = ~Q[31] /*48937*/;
assign _29464_ = _29465_ & D[57] /*48936*/;
assign _29467_ = _28666_ & _29464_ /*48931*/;
assign _29468_ = _28666_ ^ _29464_ /*48934*/;
assign _29469_ = _29460_ & _29468_ /*48932*/;
assign _29114_ = _29460_ ^ _29468_ /*48933*/;
assign _29466_ = _29467_ | _29469_ /*48930*/;
assign _29471_ = ~Q[31] /*48929*/;
assign _29470_ = _29471_ & D[58] /*48928*/;
assign _29473_ = _28667_ & _29470_ /*48923*/;
assign _29474_ = _28667_ ^ _29470_ /*48926*/;
assign _29475_ = _29466_ & _29474_ /*48924*/;
assign _29115_ = _29466_ ^ _29474_ /*48925*/;
assign _29472_ = _29473_ | _29475_ /*48922*/;
assign _29477_ = ~Q[31] /*48921*/;
assign _29476_ = _29477_ & D[59] /*48920*/;
assign _29479_ = _28668_ & _29476_ /*48915*/;
assign _29480_ = _28668_ ^ _29476_ /*48918*/;
assign _29481_ = _29472_ & _29480_ /*48916*/;
assign _29116_ = _29472_ ^ _29480_ /*48917*/;
assign _29478_ = _29479_ | _29481_ /*48914*/;
assign _29483_ = ~Q[31] /*48913*/;
assign _29482_ = _29483_ & D[60] /*48912*/;
assign _29485_ = _28669_ & _29482_ /*48907*/;
assign _29486_ = _28669_ ^ _29482_ /*48910*/;
assign _29487_ = _29478_ & _29486_ /*48908*/;
assign _29117_ = _29478_ ^ _29486_ /*48909*/;
assign _29484_ = _29485_ | _29487_ /*48906*/;
assign _29489_ = ~Q[31] /*48905*/;
assign _29488_ = _29489_ & D[61] /*48904*/;
assign _29491_ = _28670_ & _29488_ /*48899*/;
assign _29492_ = _28670_ ^ _29488_ /*48902*/;
assign _29493_ = _29484_ & _29492_ /*48900*/;
assign _29118_ = _29484_ ^ _29492_ /*48901*/;
assign _29490_ = _29491_ | _29493_ /*48898*/;
assign _29495_ = ~Q[31] /*48897*/;
assign _29494_ = _29495_ & D[62] /*48896*/;
assign _29497_ = _28671_ & _29494_ /*48891*/;
assign _29498_ = _28671_ ^ _29494_ /*48894*/;
assign _29499_ = _29490_ & _29498_ /*48892*/;
assign _29119_ = _29490_ ^ _29498_ /*48893*/;
assign _29496_ = _29497_ | _29499_ /*48890*/;
assign _29501_ = ~Q[31] /*48889*/;
assign _29500_ = _29501_ & zeroWire /*48888*/;
assign _29502_ = _28672_ ^ _29500_ /*48886*/;
assign _29120_ = _29502_ ^ _29496_ /*48885*/;
assign _29573_ = ~D[0] /*48631*/;
assign _29570_ = R_0[30] & _29573_ /*48627*/;
assign _29571_ = R_0[30] ^ _29573_ /*48630*/;
assign _29572_ = oneWire & _29571_ /*48628*/;
assign _29505_ = oneWire ^ _29571_ /*48629*/;
assign _29569_ = _29570_ | _29572_ /*48626*/;
assign _29578_ = ~D[1] /*48625*/;
assign _29575_ = _29057_ & _29578_ /*48621*/;
assign _29576_ = _29057_ ^ _29578_ /*48624*/;
assign _29577_ = _29569_ & _29576_ /*48622*/;
assign _29506_ = _29569_ ^ _29576_ /*48623*/;
assign _29574_ = _29575_ | _29577_ /*48620*/;
assign _29583_ = ~D[2] /*48619*/;
assign _29580_ = _29058_ & _29583_ /*48615*/;
assign _29581_ = _29058_ ^ _29583_ /*48618*/;
assign _29582_ = _29574_ & _29581_ /*48616*/;
assign _29507_ = _29574_ ^ _29581_ /*48617*/;
assign _29579_ = _29580_ | _29582_ /*48614*/;
assign _29588_ = ~D[3] /*48613*/;
assign _29585_ = _29059_ & _29588_ /*48609*/;
assign _29586_ = _29059_ ^ _29588_ /*48612*/;
assign _29587_ = _29579_ & _29586_ /*48610*/;
assign _29508_ = _29579_ ^ _29586_ /*48611*/;
assign _29584_ = _29585_ | _29587_ /*48608*/;
assign _29593_ = ~D[4] /*48607*/;
assign _29590_ = _29060_ & _29593_ /*48603*/;
assign _29591_ = _29060_ ^ _29593_ /*48606*/;
assign _29592_ = _29584_ & _29591_ /*48604*/;
assign _29509_ = _29584_ ^ _29591_ /*48605*/;
assign _29589_ = _29590_ | _29592_ /*48602*/;
assign _29598_ = ~D[5] /*48601*/;
assign _29595_ = _29061_ & _29598_ /*48597*/;
assign _29596_ = _29061_ ^ _29598_ /*48600*/;
assign _29597_ = _29589_ & _29596_ /*48598*/;
assign _29510_ = _29589_ ^ _29596_ /*48599*/;
assign _29594_ = _29595_ | _29597_ /*48596*/;
assign _29603_ = ~D[6] /*48595*/;
assign _29600_ = _29062_ & _29603_ /*48591*/;
assign _29601_ = _29062_ ^ _29603_ /*48594*/;
assign _29602_ = _29594_ & _29601_ /*48592*/;
assign _29511_ = _29594_ ^ _29601_ /*48593*/;
assign _29599_ = _29600_ | _29602_ /*48590*/;
assign _29608_ = ~D[7] /*48589*/;
assign _29605_ = _29063_ & _29608_ /*48585*/;
assign _29606_ = _29063_ ^ _29608_ /*48588*/;
assign _29607_ = _29599_ & _29606_ /*48586*/;
assign _29512_ = _29599_ ^ _29606_ /*48587*/;
assign _29604_ = _29605_ | _29607_ /*48584*/;
assign _29613_ = ~D[8] /*48583*/;
assign _29610_ = _29064_ & _29613_ /*48579*/;
assign _29611_ = _29064_ ^ _29613_ /*48582*/;
assign _29612_ = _29604_ & _29611_ /*48580*/;
assign _29513_ = _29604_ ^ _29611_ /*48581*/;
assign _29609_ = _29610_ | _29612_ /*48578*/;
assign _29618_ = ~D[9] /*48577*/;
assign _29615_ = _29065_ & _29618_ /*48573*/;
assign _29616_ = _29065_ ^ _29618_ /*48576*/;
assign _29617_ = _29609_ & _29616_ /*48574*/;
assign _29514_ = _29609_ ^ _29616_ /*48575*/;
assign _29614_ = _29615_ | _29617_ /*48572*/;
assign _29623_ = ~D[10] /*48571*/;
assign _29620_ = _29066_ & _29623_ /*48567*/;
assign _29621_ = _29066_ ^ _29623_ /*48570*/;
assign _29622_ = _29614_ & _29621_ /*48568*/;
assign _29515_ = _29614_ ^ _29621_ /*48569*/;
assign _29619_ = _29620_ | _29622_ /*48566*/;
assign _29628_ = ~D[11] /*48565*/;
assign _29625_ = _29067_ & _29628_ /*48561*/;
assign _29626_ = _29067_ ^ _29628_ /*48564*/;
assign _29627_ = _29619_ & _29626_ /*48562*/;
assign _29516_ = _29619_ ^ _29626_ /*48563*/;
assign _29624_ = _29625_ | _29627_ /*48560*/;
assign _29633_ = ~D[12] /*48559*/;
assign _29630_ = _29068_ & _29633_ /*48555*/;
assign _29631_ = _29068_ ^ _29633_ /*48558*/;
assign _29632_ = _29624_ & _29631_ /*48556*/;
assign _29517_ = _29624_ ^ _29631_ /*48557*/;
assign _29629_ = _29630_ | _29632_ /*48554*/;
assign _29638_ = ~D[13] /*48553*/;
assign _29635_ = _29069_ & _29638_ /*48549*/;
assign _29636_ = _29069_ ^ _29638_ /*48552*/;
assign _29637_ = _29629_ & _29636_ /*48550*/;
assign _29518_ = _29629_ ^ _29636_ /*48551*/;
assign _29634_ = _29635_ | _29637_ /*48548*/;
assign _29643_ = ~D[14] /*48547*/;
assign _29640_ = _29070_ & _29643_ /*48543*/;
assign _29641_ = _29070_ ^ _29643_ /*48546*/;
assign _29642_ = _29634_ & _29641_ /*48544*/;
assign _29519_ = _29634_ ^ _29641_ /*48545*/;
assign _29639_ = _29640_ | _29642_ /*48542*/;
assign _29648_ = ~D[15] /*48541*/;
assign _29645_ = _29071_ & _29648_ /*48537*/;
assign _29646_ = _29071_ ^ _29648_ /*48540*/;
assign _29647_ = _29639_ & _29646_ /*48538*/;
assign _29520_ = _29639_ ^ _29646_ /*48539*/;
assign _29644_ = _29645_ | _29647_ /*48536*/;
assign _29653_ = ~D[16] /*48535*/;
assign _29650_ = _29072_ & _29653_ /*48531*/;
assign _29651_ = _29072_ ^ _29653_ /*48534*/;
assign _29652_ = _29644_ & _29651_ /*48532*/;
assign _29521_ = _29644_ ^ _29651_ /*48533*/;
assign _29649_ = _29650_ | _29652_ /*48530*/;
assign _29658_ = ~D[17] /*48529*/;
assign _29655_ = _29073_ & _29658_ /*48525*/;
assign _29656_ = _29073_ ^ _29658_ /*48528*/;
assign _29657_ = _29649_ & _29656_ /*48526*/;
assign _29522_ = _29649_ ^ _29656_ /*48527*/;
assign _29654_ = _29655_ | _29657_ /*48524*/;
assign _29663_ = ~D[18] /*48523*/;
assign _29660_ = _29074_ & _29663_ /*48519*/;
assign _29661_ = _29074_ ^ _29663_ /*48522*/;
assign _29662_ = _29654_ & _29661_ /*48520*/;
assign _29523_ = _29654_ ^ _29661_ /*48521*/;
assign _29659_ = _29660_ | _29662_ /*48518*/;
assign _29668_ = ~D[19] /*48517*/;
assign _29665_ = _29075_ & _29668_ /*48513*/;
assign _29666_ = _29075_ ^ _29668_ /*48516*/;
assign _29667_ = _29659_ & _29666_ /*48514*/;
assign _29524_ = _29659_ ^ _29666_ /*48515*/;
assign _29664_ = _29665_ | _29667_ /*48512*/;
assign _29673_ = ~D[20] /*48511*/;
assign _29670_ = _29076_ & _29673_ /*48507*/;
assign _29671_ = _29076_ ^ _29673_ /*48510*/;
assign _29672_ = _29664_ & _29671_ /*48508*/;
assign _29525_ = _29664_ ^ _29671_ /*48509*/;
assign _29669_ = _29670_ | _29672_ /*48506*/;
assign _29678_ = ~D[21] /*48505*/;
assign _29675_ = _29077_ & _29678_ /*48501*/;
assign _29676_ = _29077_ ^ _29678_ /*48504*/;
assign _29677_ = _29669_ & _29676_ /*48502*/;
assign _29526_ = _29669_ ^ _29676_ /*48503*/;
assign _29674_ = _29675_ | _29677_ /*48500*/;
assign _29683_ = ~D[22] /*48499*/;
assign _29680_ = _29078_ & _29683_ /*48495*/;
assign _29681_ = _29078_ ^ _29683_ /*48498*/;
assign _29682_ = _29674_ & _29681_ /*48496*/;
assign _29527_ = _29674_ ^ _29681_ /*48497*/;
assign _29679_ = _29680_ | _29682_ /*48494*/;
assign _29688_ = ~D[23] /*48493*/;
assign _29685_ = _29079_ & _29688_ /*48489*/;
assign _29686_ = _29079_ ^ _29688_ /*48492*/;
assign _29687_ = _29679_ & _29686_ /*48490*/;
assign _29528_ = _29679_ ^ _29686_ /*48491*/;
assign _29684_ = _29685_ | _29687_ /*48488*/;
assign _29693_ = ~D[24] /*48487*/;
assign _29690_ = _29080_ & _29693_ /*48483*/;
assign _29691_ = _29080_ ^ _29693_ /*48486*/;
assign _29692_ = _29684_ & _29691_ /*48484*/;
assign _29529_ = _29684_ ^ _29691_ /*48485*/;
assign _29689_ = _29690_ | _29692_ /*48482*/;
assign _29698_ = ~D[25] /*48481*/;
assign _29695_ = _29081_ & _29698_ /*48477*/;
assign _29696_ = _29081_ ^ _29698_ /*48480*/;
assign _29697_ = _29689_ & _29696_ /*48478*/;
assign _29530_ = _29689_ ^ _29696_ /*48479*/;
assign _29694_ = _29695_ | _29697_ /*48476*/;
assign _29703_ = ~D[26] /*48475*/;
assign _29700_ = _29082_ & _29703_ /*48471*/;
assign _29701_ = _29082_ ^ _29703_ /*48474*/;
assign _29702_ = _29694_ & _29701_ /*48472*/;
assign _29531_ = _29694_ ^ _29701_ /*48473*/;
assign _29699_ = _29700_ | _29702_ /*48470*/;
assign _29708_ = ~D[27] /*48469*/;
assign _29705_ = _29083_ & _29708_ /*48465*/;
assign _29706_ = _29083_ ^ _29708_ /*48468*/;
assign _29707_ = _29699_ & _29706_ /*48466*/;
assign _29532_ = _29699_ ^ _29706_ /*48467*/;
assign _29704_ = _29705_ | _29707_ /*48464*/;
assign _29713_ = ~D[28] /*48463*/;
assign _29710_ = _29084_ & _29713_ /*48459*/;
assign _29711_ = _29084_ ^ _29713_ /*48462*/;
assign _29712_ = _29704_ & _29711_ /*48460*/;
assign _29533_ = _29704_ ^ _29711_ /*48461*/;
assign _29709_ = _29710_ | _29712_ /*48458*/;
assign _29718_ = ~D[29] /*48457*/;
assign _29715_ = _29085_ & _29718_ /*48453*/;
assign _29716_ = _29085_ ^ _29718_ /*48456*/;
assign _29717_ = _29709_ & _29716_ /*48454*/;
assign _29534_ = _29709_ ^ _29716_ /*48455*/;
assign _29714_ = _29715_ | _29717_ /*48452*/;
assign _29723_ = ~D[30] /*48451*/;
assign _29720_ = _29086_ & _29723_ /*48447*/;
assign _29721_ = _29086_ ^ _29723_ /*48450*/;
assign _29722_ = _29714_ & _29721_ /*48448*/;
assign _29535_ = _29714_ ^ _29721_ /*48449*/;
assign _29719_ = _29720_ | _29722_ /*48446*/;
assign _29728_ = ~D[31] /*48445*/;
assign _29725_ = _29087_ & _29728_ /*48441*/;
assign _29726_ = _29087_ ^ _29728_ /*48444*/;
assign _29727_ = _29719_ & _29726_ /*48442*/;
assign _29536_ = _29719_ ^ _29726_ /*48443*/;
assign _29724_ = _29725_ | _29727_ /*48440*/;
assign _29733_ = ~D[32] /*48439*/;
assign _29730_ = _29088_ & _29733_ /*48435*/;
assign _29731_ = _29088_ ^ _29733_ /*48438*/;
assign _29732_ = _29724_ & _29731_ /*48436*/;
assign _29537_ = _29724_ ^ _29731_ /*48437*/;
assign _29729_ = _29730_ | _29732_ /*48434*/;
assign _29738_ = ~D[33] /*48433*/;
assign _29735_ = _29089_ & _29738_ /*48429*/;
assign _29736_ = _29089_ ^ _29738_ /*48432*/;
assign _29737_ = _29729_ & _29736_ /*48430*/;
assign _29538_ = _29729_ ^ _29736_ /*48431*/;
assign _29734_ = _29735_ | _29737_ /*48428*/;
assign _29743_ = ~D[34] /*48427*/;
assign _29740_ = _29090_ & _29743_ /*48423*/;
assign _29741_ = _29090_ ^ _29743_ /*48426*/;
assign _29742_ = _29734_ & _29741_ /*48424*/;
assign _29539_ = _29734_ ^ _29741_ /*48425*/;
assign _29739_ = _29740_ | _29742_ /*48422*/;
assign _29748_ = ~D[35] /*48421*/;
assign _29745_ = _29091_ & _29748_ /*48417*/;
assign _29746_ = _29091_ ^ _29748_ /*48420*/;
assign _29747_ = _29739_ & _29746_ /*48418*/;
assign _29540_ = _29739_ ^ _29746_ /*48419*/;
assign _29744_ = _29745_ | _29747_ /*48416*/;
assign _29753_ = ~D[36] /*48415*/;
assign _29750_ = _29092_ & _29753_ /*48411*/;
assign _29751_ = _29092_ ^ _29753_ /*48414*/;
assign _29752_ = _29744_ & _29751_ /*48412*/;
assign _29541_ = _29744_ ^ _29751_ /*48413*/;
assign _29749_ = _29750_ | _29752_ /*48410*/;
assign _29758_ = ~D[37] /*48409*/;
assign _29755_ = _29093_ & _29758_ /*48405*/;
assign _29756_ = _29093_ ^ _29758_ /*48408*/;
assign _29757_ = _29749_ & _29756_ /*48406*/;
assign _29542_ = _29749_ ^ _29756_ /*48407*/;
assign _29754_ = _29755_ | _29757_ /*48404*/;
assign _29763_ = ~D[38] /*48403*/;
assign _29760_ = _29094_ & _29763_ /*48399*/;
assign _29761_ = _29094_ ^ _29763_ /*48402*/;
assign _29762_ = _29754_ & _29761_ /*48400*/;
assign _29543_ = _29754_ ^ _29761_ /*48401*/;
assign _29759_ = _29760_ | _29762_ /*48398*/;
assign _29768_ = ~D[39] /*48397*/;
assign _29765_ = _29095_ & _29768_ /*48393*/;
assign _29766_ = _29095_ ^ _29768_ /*48396*/;
assign _29767_ = _29759_ & _29766_ /*48394*/;
assign _29544_ = _29759_ ^ _29766_ /*48395*/;
assign _29764_ = _29765_ | _29767_ /*48392*/;
assign _29773_ = ~D[40] /*48391*/;
assign _29770_ = _29096_ & _29773_ /*48387*/;
assign _29771_ = _29096_ ^ _29773_ /*48390*/;
assign _29772_ = _29764_ & _29771_ /*48388*/;
assign _29545_ = _29764_ ^ _29771_ /*48389*/;
assign _29769_ = _29770_ | _29772_ /*48386*/;
assign _29778_ = ~D[41] /*48385*/;
assign _29775_ = _29097_ & _29778_ /*48381*/;
assign _29776_ = _29097_ ^ _29778_ /*48384*/;
assign _29777_ = _29769_ & _29776_ /*48382*/;
assign _29546_ = _29769_ ^ _29776_ /*48383*/;
assign _29774_ = _29775_ | _29777_ /*48380*/;
assign _29783_ = ~D[42] /*48379*/;
assign _29780_ = _29098_ & _29783_ /*48375*/;
assign _29781_ = _29098_ ^ _29783_ /*48378*/;
assign _29782_ = _29774_ & _29781_ /*48376*/;
assign _29547_ = _29774_ ^ _29781_ /*48377*/;
assign _29779_ = _29780_ | _29782_ /*48374*/;
assign _29788_ = ~D[43] /*48373*/;
assign _29785_ = _29099_ & _29788_ /*48369*/;
assign _29786_ = _29099_ ^ _29788_ /*48372*/;
assign _29787_ = _29779_ & _29786_ /*48370*/;
assign _29548_ = _29779_ ^ _29786_ /*48371*/;
assign _29784_ = _29785_ | _29787_ /*48368*/;
assign _29793_ = ~D[44] /*48367*/;
assign _29790_ = _29100_ & _29793_ /*48363*/;
assign _29791_ = _29100_ ^ _29793_ /*48366*/;
assign _29792_ = _29784_ & _29791_ /*48364*/;
assign _29549_ = _29784_ ^ _29791_ /*48365*/;
assign _29789_ = _29790_ | _29792_ /*48362*/;
assign _29798_ = ~D[45] /*48361*/;
assign _29795_ = _29101_ & _29798_ /*48357*/;
assign _29796_ = _29101_ ^ _29798_ /*48360*/;
assign _29797_ = _29789_ & _29796_ /*48358*/;
assign _29550_ = _29789_ ^ _29796_ /*48359*/;
assign _29794_ = _29795_ | _29797_ /*48356*/;
assign _29803_ = ~D[46] /*48355*/;
assign _29800_ = _29102_ & _29803_ /*48351*/;
assign _29801_ = _29102_ ^ _29803_ /*48354*/;
assign _29802_ = _29794_ & _29801_ /*48352*/;
assign _29551_ = _29794_ ^ _29801_ /*48353*/;
assign _29799_ = _29800_ | _29802_ /*48350*/;
assign _29808_ = ~D[47] /*48349*/;
assign _29805_ = _29103_ & _29808_ /*48345*/;
assign _29806_ = _29103_ ^ _29808_ /*48348*/;
assign _29807_ = _29799_ & _29806_ /*48346*/;
assign _29552_ = _29799_ ^ _29806_ /*48347*/;
assign _29804_ = _29805_ | _29807_ /*48344*/;
assign _29813_ = ~D[48] /*48343*/;
assign _29810_ = _29104_ & _29813_ /*48339*/;
assign _29811_ = _29104_ ^ _29813_ /*48342*/;
assign _29812_ = _29804_ & _29811_ /*48340*/;
assign _29553_ = _29804_ ^ _29811_ /*48341*/;
assign _29809_ = _29810_ | _29812_ /*48338*/;
assign _29818_ = ~D[49] /*48337*/;
assign _29815_ = _29105_ & _29818_ /*48333*/;
assign _29816_ = _29105_ ^ _29818_ /*48336*/;
assign _29817_ = _29809_ & _29816_ /*48334*/;
assign _29554_ = _29809_ ^ _29816_ /*48335*/;
assign _29814_ = _29815_ | _29817_ /*48332*/;
assign _29823_ = ~D[50] /*48331*/;
assign _29820_ = _29106_ & _29823_ /*48327*/;
assign _29821_ = _29106_ ^ _29823_ /*48330*/;
assign _29822_ = _29814_ & _29821_ /*48328*/;
assign _29555_ = _29814_ ^ _29821_ /*48329*/;
assign _29819_ = _29820_ | _29822_ /*48326*/;
assign _29828_ = ~D[51] /*48325*/;
assign _29825_ = _29107_ & _29828_ /*48321*/;
assign _29826_ = _29107_ ^ _29828_ /*48324*/;
assign _29827_ = _29819_ & _29826_ /*48322*/;
assign _29556_ = _29819_ ^ _29826_ /*48323*/;
assign _29824_ = _29825_ | _29827_ /*48320*/;
assign _29833_ = ~D[52] /*48319*/;
assign _29830_ = _29108_ & _29833_ /*48315*/;
assign _29831_ = _29108_ ^ _29833_ /*48318*/;
assign _29832_ = _29824_ & _29831_ /*48316*/;
assign _29557_ = _29824_ ^ _29831_ /*48317*/;
assign _29829_ = _29830_ | _29832_ /*48314*/;
assign _29838_ = ~D[53] /*48313*/;
assign _29835_ = _29109_ & _29838_ /*48309*/;
assign _29836_ = _29109_ ^ _29838_ /*48312*/;
assign _29837_ = _29829_ & _29836_ /*48310*/;
assign _29558_ = _29829_ ^ _29836_ /*48311*/;
assign _29834_ = _29835_ | _29837_ /*48308*/;
assign _29843_ = ~D[54] /*48307*/;
assign _29840_ = _29110_ & _29843_ /*48303*/;
assign _29841_ = _29110_ ^ _29843_ /*48306*/;
assign _29842_ = _29834_ & _29841_ /*48304*/;
assign _29559_ = _29834_ ^ _29841_ /*48305*/;
assign _29839_ = _29840_ | _29842_ /*48302*/;
assign _29848_ = ~D[55] /*48301*/;
assign _29845_ = _29111_ & _29848_ /*48297*/;
assign _29846_ = _29111_ ^ _29848_ /*48300*/;
assign _29847_ = _29839_ & _29846_ /*48298*/;
assign _29560_ = _29839_ ^ _29846_ /*48299*/;
assign _29844_ = _29845_ | _29847_ /*48296*/;
assign _29853_ = ~D[56] /*48295*/;
assign _29850_ = _29112_ & _29853_ /*48291*/;
assign _29851_ = _29112_ ^ _29853_ /*48294*/;
assign _29852_ = _29844_ & _29851_ /*48292*/;
assign _29561_ = _29844_ ^ _29851_ /*48293*/;
assign _29849_ = _29850_ | _29852_ /*48290*/;
assign _29858_ = ~D[57] /*48289*/;
assign _29855_ = _29113_ & _29858_ /*48285*/;
assign _29856_ = _29113_ ^ _29858_ /*48288*/;
assign _29857_ = _29849_ & _29856_ /*48286*/;
assign _29562_ = _29849_ ^ _29856_ /*48287*/;
assign _29854_ = _29855_ | _29857_ /*48284*/;
assign _29863_ = ~D[58] /*48283*/;
assign _29860_ = _29114_ & _29863_ /*48279*/;
assign _29861_ = _29114_ ^ _29863_ /*48282*/;
assign _29862_ = _29854_ & _29861_ /*48280*/;
assign _29563_ = _29854_ ^ _29861_ /*48281*/;
assign _29859_ = _29860_ | _29862_ /*48278*/;
assign _29868_ = ~D[59] /*48277*/;
assign _29865_ = _29115_ & _29868_ /*48273*/;
assign _29866_ = _29115_ ^ _29868_ /*48276*/;
assign _29867_ = _29859_ & _29866_ /*48274*/;
assign _29564_ = _29859_ ^ _29866_ /*48275*/;
assign _29864_ = _29865_ | _29867_ /*48272*/;
assign _29873_ = ~D[60] /*48271*/;
assign _29870_ = _29116_ & _29873_ /*48267*/;
assign _29871_ = _29116_ ^ _29873_ /*48270*/;
assign _29872_ = _29864_ & _29871_ /*48268*/;
assign _29565_ = _29864_ ^ _29871_ /*48269*/;
assign _29869_ = _29870_ | _29872_ /*48266*/;
assign _29878_ = ~D[61] /*48265*/;
assign _29875_ = _29117_ & _29878_ /*48261*/;
assign _29876_ = _29117_ ^ _29878_ /*48264*/;
assign _29877_ = _29869_ & _29876_ /*48262*/;
assign _29566_ = _29869_ ^ _29876_ /*48263*/;
assign _29874_ = _29875_ | _29877_ /*48260*/;
assign _29883_ = ~D[62] /*48259*/;
assign _29880_ = _29118_ & _29883_ /*48255*/;
assign _29881_ = _29118_ ^ _29883_ /*48258*/;
assign _29882_ = _29874_ & _29881_ /*48256*/;
assign _29567_ = _29874_ ^ _29881_ /*48257*/;
assign _29879_ = _29880_ | _29882_ /*48254*/;
assign _29884_ = _29119_ & oneWire /*48249*/;
assign _29885_ = _29119_ ^ oneWire /*48252*/;
assign _29886_ = _29879_ & _29885_ /*48250*/;
assign _29568_ = _29879_ ^ _29885_ /*48251*/;
assign Q[30] = _29884_ | _29886_ /*48248*/;
assign _30019_ = ~Q[30] /*47863*/;
assign _30018_ = _30019_ & D[0] /*47862*/;
assign _30021_ = _29505_ & _30018_ /*47857*/;
assign _30022_ = _29505_ ^ _30018_ /*47860*/;
assign _30023_ = zeroWire & _30022_ /*47858*/;
assign _29953_ = zeroWire ^ _30022_ /*47859*/;
assign _30020_ = _30021_ | _30023_ /*47856*/;
assign _30025_ = ~Q[30] /*47855*/;
assign _30024_ = _30025_ & D[1] /*47854*/;
assign _30027_ = _29506_ & _30024_ /*47849*/;
assign _30028_ = _29506_ ^ _30024_ /*47852*/;
assign _30029_ = _30020_ & _30028_ /*47850*/;
assign _29954_ = _30020_ ^ _30028_ /*47851*/;
assign _30026_ = _30027_ | _30029_ /*47848*/;
assign _30031_ = ~Q[30] /*47847*/;
assign _30030_ = _30031_ & D[2] /*47846*/;
assign _30033_ = _29507_ & _30030_ /*47841*/;
assign _30034_ = _29507_ ^ _30030_ /*47844*/;
assign _30035_ = _30026_ & _30034_ /*47842*/;
assign _29955_ = _30026_ ^ _30034_ /*47843*/;
assign _30032_ = _30033_ | _30035_ /*47840*/;
assign _30037_ = ~Q[30] /*47839*/;
assign _30036_ = _30037_ & D[3] /*47838*/;
assign _30039_ = _29508_ & _30036_ /*47833*/;
assign _30040_ = _29508_ ^ _30036_ /*47836*/;
assign _30041_ = _30032_ & _30040_ /*47834*/;
assign _29956_ = _30032_ ^ _30040_ /*47835*/;
assign _30038_ = _30039_ | _30041_ /*47832*/;
assign _30043_ = ~Q[30] /*47831*/;
assign _30042_ = _30043_ & D[4] /*47830*/;
assign _30045_ = _29509_ & _30042_ /*47825*/;
assign _30046_ = _29509_ ^ _30042_ /*47828*/;
assign _30047_ = _30038_ & _30046_ /*47826*/;
assign _29957_ = _30038_ ^ _30046_ /*47827*/;
assign _30044_ = _30045_ | _30047_ /*47824*/;
assign _30049_ = ~Q[30] /*47823*/;
assign _30048_ = _30049_ & D[5] /*47822*/;
assign _30051_ = _29510_ & _30048_ /*47817*/;
assign _30052_ = _29510_ ^ _30048_ /*47820*/;
assign _30053_ = _30044_ & _30052_ /*47818*/;
assign _29958_ = _30044_ ^ _30052_ /*47819*/;
assign _30050_ = _30051_ | _30053_ /*47816*/;
assign _30055_ = ~Q[30] /*47815*/;
assign _30054_ = _30055_ & D[6] /*47814*/;
assign _30057_ = _29511_ & _30054_ /*47809*/;
assign _30058_ = _29511_ ^ _30054_ /*47812*/;
assign _30059_ = _30050_ & _30058_ /*47810*/;
assign _29959_ = _30050_ ^ _30058_ /*47811*/;
assign _30056_ = _30057_ | _30059_ /*47808*/;
assign _30061_ = ~Q[30] /*47807*/;
assign _30060_ = _30061_ & D[7] /*47806*/;
assign _30063_ = _29512_ & _30060_ /*47801*/;
assign _30064_ = _29512_ ^ _30060_ /*47804*/;
assign _30065_ = _30056_ & _30064_ /*47802*/;
assign _29960_ = _30056_ ^ _30064_ /*47803*/;
assign _30062_ = _30063_ | _30065_ /*47800*/;
assign _30067_ = ~Q[30] /*47799*/;
assign _30066_ = _30067_ & D[8] /*47798*/;
assign _30069_ = _29513_ & _30066_ /*47793*/;
assign _30070_ = _29513_ ^ _30066_ /*47796*/;
assign _30071_ = _30062_ & _30070_ /*47794*/;
assign _29961_ = _30062_ ^ _30070_ /*47795*/;
assign _30068_ = _30069_ | _30071_ /*47792*/;
assign _30073_ = ~Q[30] /*47791*/;
assign _30072_ = _30073_ & D[9] /*47790*/;
assign _30075_ = _29514_ & _30072_ /*47785*/;
assign _30076_ = _29514_ ^ _30072_ /*47788*/;
assign _30077_ = _30068_ & _30076_ /*47786*/;
assign _29962_ = _30068_ ^ _30076_ /*47787*/;
assign _30074_ = _30075_ | _30077_ /*47784*/;
assign _30079_ = ~Q[30] /*47783*/;
assign _30078_ = _30079_ & D[10] /*47782*/;
assign _30081_ = _29515_ & _30078_ /*47777*/;
assign _30082_ = _29515_ ^ _30078_ /*47780*/;
assign _30083_ = _30074_ & _30082_ /*47778*/;
assign _29963_ = _30074_ ^ _30082_ /*47779*/;
assign _30080_ = _30081_ | _30083_ /*47776*/;
assign _30085_ = ~Q[30] /*47775*/;
assign _30084_ = _30085_ & D[11] /*47774*/;
assign _30087_ = _29516_ & _30084_ /*47769*/;
assign _30088_ = _29516_ ^ _30084_ /*47772*/;
assign _30089_ = _30080_ & _30088_ /*47770*/;
assign _29964_ = _30080_ ^ _30088_ /*47771*/;
assign _30086_ = _30087_ | _30089_ /*47768*/;
assign _30091_ = ~Q[30] /*47767*/;
assign _30090_ = _30091_ & D[12] /*47766*/;
assign _30093_ = _29517_ & _30090_ /*47761*/;
assign _30094_ = _29517_ ^ _30090_ /*47764*/;
assign _30095_ = _30086_ & _30094_ /*47762*/;
assign _29965_ = _30086_ ^ _30094_ /*47763*/;
assign _30092_ = _30093_ | _30095_ /*47760*/;
assign _30097_ = ~Q[30] /*47759*/;
assign _30096_ = _30097_ & D[13] /*47758*/;
assign _30099_ = _29518_ & _30096_ /*47753*/;
assign _30100_ = _29518_ ^ _30096_ /*47756*/;
assign _30101_ = _30092_ & _30100_ /*47754*/;
assign _29966_ = _30092_ ^ _30100_ /*47755*/;
assign _30098_ = _30099_ | _30101_ /*47752*/;
assign _30103_ = ~Q[30] /*47751*/;
assign _30102_ = _30103_ & D[14] /*47750*/;
assign _30105_ = _29519_ & _30102_ /*47745*/;
assign _30106_ = _29519_ ^ _30102_ /*47748*/;
assign _30107_ = _30098_ & _30106_ /*47746*/;
assign _29967_ = _30098_ ^ _30106_ /*47747*/;
assign _30104_ = _30105_ | _30107_ /*47744*/;
assign _30109_ = ~Q[30] /*47743*/;
assign _30108_ = _30109_ & D[15] /*47742*/;
assign _30111_ = _29520_ & _30108_ /*47737*/;
assign _30112_ = _29520_ ^ _30108_ /*47740*/;
assign _30113_ = _30104_ & _30112_ /*47738*/;
assign _29968_ = _30104_ ^ _30112_ /*47739*/;
assign _30110_ = _30111_ | _30113_ /*47736*/;
assign _30115_ = ~Q[30] /*47735*/;
assign _30114_ = _30115_ & D[16] /*47734*/;
assign _30117_ = _29521_ & _30114_ /*47729*/;
assign _30118_ = _29521_ ^ _30114_ /*47732*/;
assign _30119_ = _30110_ & _30118_ /*47730*/;
assign _29969_ = _30110_ ^ _30118_ /*47731*/;
assign _30116_ = _30117_ | _30119_ /*47728*/;
assign _30121_ = ~Q[30] /*47727*/;
assign _30120_ = _30121_ & D[17] /*47726*/;
assign _30123_ = _29522_ & _30120_ /*47721*/;
assign _30124_ = _29522_ ^ _30120_ /*47724*/;
assign _30125_ = _30116_ & _30124_ /*47722*/;
assign _29970_ = _30116_ ^ _30124_ /*47723*/;
assign _30122_ = _30123_ | _30125_ /*47720*/;
assign _30127_ = ~Q[30] /*47719*/;
assign _30126_ = _30127_ & D[18] /*47718*/;
assign _30129_ = _29523_ & _30126_ /*47713*/;
assign _30130_ = _29523_ ^ _30126_ /*47716*/;
assign _30131_ = _30122_ & _30130_ /*47714*/;
assign _29971_ = _30122_ ^ _30130_ /*47715*/;
assign _30128_ = _30129_ | _30131_ /*47712*/;
assign _30133_ = ~Q[30] /*47711*/;
assign _30132_ = _30133_ & D[19] /*47710*/;
assign _30135_ = _29524_ & _30132_ /*47705*/;
assign _30136_ = _29524_ ^ _30132_ /*47708*/;
assign _30137_ = _30128_ & _30136_ /*47706*/;
assign _29972_ = _30128_ ^ _30136_ /*47707*/;
assign _30134_ = _30135_ | _30137_ /*47704*/;
assign _30139_ = ~Q[30] /*47703*/;
assign _30138_ = _30139_ & D[20] /*47702*/;
assign _30141_ = _29525_ & _30138_ /*47697*/;
assign _30142_ = _29525_ ^ _30138_ /*47700*/;
assign _30143_ = _30134_ & _30142_ /*47698*/;
assign _29973_ = _30134_ ^ _30142_ /*47699*/;
assign _30140_ = _30141_ | _30143_ /*47696*/;
assign _30145_ = ~Q[30] /*47695*/;
assign _30144_ = _30145_ & D[21] /*47694*/;
assign _30147_ = _29526_ & _30144_ /*47689*/;
assign _30148_ = _29526_ ^ _30144_ /*47692*/;
assign _30149_ = _30140_ & _30148_ /*47690*/;
assign _29974_ = _30140_ ^ _30148_ /*47691*/;
assign _30146_ = _30147_ | _30149_ /*47688*/;
assign _30151_ = ~Q[30] /*47687*/;
assign _30150_ = _30151_ & D[22] /*47686*/;
assign _30153_ = _29527_ & _30150_ /*47681*/;
assign _30154_ = _29527_ ^ _30150_ /*47684*/;
assign _30155_ = _30146_ & _30154_ /*47682*/;
assign _29975_ = _30146_ ^ _30154_ /*47683*/;
assign _30152_ = _30153_ | _30155_ /*47680*/;
assign _30157_ = ~Q[30] /*47679*/;
assign _30156_ = _30157_ & D[23] /*47678*/;
assign _30159_ = _29528_ & _30156_ /*47673*/;
assign _30160_ = _29528_ ^ _30156_ /*47676*/;
assign _30161_ = _30152_ & _30160_ /*47674*/;
assign _29976_ = _30152_ ^ _30160_ /*47675*/;
assign _30158_ = _30159_ | _30161_ /*47672*/;
assign _30163_ = ~Q[30] /*47671*/;
assign _30162_ = _30163_ & D[24] /*47670*/;
assign _30165_ = _29529_ & _30162_ /*47665*/;
assign _30166_ = _29529_ ^ _30162_ /*47668*/;
assign _30167_ = _30158_ & _30166_ /*47666*/;
assign _29977_ = _30158_ ^ _30166_ /*47667*/;
assign _30164_ = _30165_ | _30167_ /*47664*/;
assign _30169_ = ~Q[30] /*47663*/;
assign _30168_ = _30169_ & D[25] /*47662*/;
assign _30171_ = _29530_ & _30168_ /*47657*/;
assign _30172_ = _29530_ ^ _30168_ /*47660*/;
assign _30173_ = _30164_ & _30172_ /*47658*/;
assign _29978_ = _30164_ ^ _30172_ /*47659*/;
assign _30170_ = _30171_ | _30173_ /*47656*/;
assign _30175_ = ~Q[30] /*47655*/;
assign _30174_ = _30175_ & D[26] /*47654*/;
assign _30177_ = _29531_ & _30174_ /*47649*/;
assign _30178_ = _29531_ ^ _30174_ /*47652*/;
assign _30179_ = _30170_ & _30178_ /*47650*/;
assign _29979_ = _30170_ ^ _30178_ /*47651*/;
assign _30176_ = _30177_ | _30179_ /*47648*/;
assign _30181_ = ~Q[30] /*47647*/;
assign _30180_ = _30181_ & D[27] /*47646*/;
assign _30183_ = _29532_ & _30180_ /*47641*/;
assign _30184_ = _29532_ ^ _30180_ /*47644*/;
assign _30185_ = _30176_ & _30184_ /*47642*/;
assign _29980_ = _30176_ ^ _30184_ /*47643*/;
assign _30182_ = _30183_ | _30185_ /*47640*/;
assign _30187_ = ~Q[30] /*47639*/;
assign _30186_ = _30187_ & D[28] /*47638*/;
assign _30189_ = _29533_ & _30186_ /*47633*/;
assign _30190_ = _29533_ ^ _30186_ /*47636*/;
assign _30191_ = _30182_ & _30190_ /*47634*/;
assign _29981_ = _30182_ ^ _30190_ /*47635*/;
assign _30188_ = _30189_ | _30191_ /*47632*/;
assign _30193_ = ~Q[30] /*47631*/;
assign _30192_ = _30193_ & D[29] /*47630*/;
assign _30195_ = _29534_ & _30192_ /*47625*/;
assign _30196_ = _29534_ ^ _30192_ /*47628*/;
assign _30197_ = _30188_ & _30196_ /*47626*/;
assign _29982_ = _30188_ ^ _30196_ /*47627*/;
assign _30194_ = _30195_ | _30197_ /*47624*/;
assign _30199_ = ~Q[30] /*47623*/;
assign _30198_ = _30199_ & D[30] /*47622*/;
assign _30201_ = _29535_ & _30198_ /*47617*/;
assign _30202_ = _29535_ ^ _30198_ /*47620*/;
assign _30203_ = _30194_ & _30202_ /*47618*/;
assign _29983_ = _30194_ ^ _30202_ /*47619*/;
assign _30200_ = _30201_ | _30203_ /*47616*/;
assign _30205_ = ~Q[30] /*47615*/;
assign _30204_ = _30205_ & D[31] /*47614*/;
assign _30207_ = _29536_ & _30204_ /*47609*/;
assign _30208_ = _29536_ ^ _30204_ /*47612*/;
assign _30209_ = _30200_ & _30208_ /*47610*/;
assign _29984_ = _30200_ ^ _30208_ /*47611*/;
assign _30206_ = _30207_ | _30209_ /*47608*/;
assign _30211_ = ~Q[30] /*47607*/;
assign _30210_ = _30211_ & D[32] /*47606*/;
assign _30213_ = _29537_ & _30210_ /*47601*/;
assign _30214_ = _29537_ ^ _30210_ /*47604*/;
assign _30215_ = _30206_ & _30214_ /*47602*/;
assign _29985_ = _30206_ ^ _30214_ /*47603*/;
assign _30212_ = _30213_ | _30215_ /*47600*/;
assign _30217_ = ~Q[30] /*47599*/;
assign _30216_ = _30217_ & D[33] /*47598*/;
assign _30219_ = _29538_ & _30216_ /*47593*/;
assign _30220_ = _29538_ ^ _30216_ /*47596*/;
assign _30221_ = _30212_ & _30220_ /*47594*/;
assign _29986_ = _30212_ ^ _30220_ /*47595*/;
assign _30218_ = _30219_ | _30221_ /*47592*/;
assign _30223_ = ~Q[30] /*47591*/;
assign _30222_ = _30223_ & D[34] /*47590*/;
assign _30225_ = _29539_ & _30222_ /*47585*/;
assign _30226_ = _29539_ ^ _30222_ /*47588*/;
assign _30227_ = _30218_ & _30226_ /*47586*/;
assign _29987_ = _30218_ ^ _30226_ /*47587*/;
assign _30224_ = _30225_ | _30227_ /*47584*/;
assign _30229_ = ~Q[30] /*47583*/;
assign _30228_ = _30229_ & D[35] /*47582*/;
assign _30231_ = _29540_ & _30228_ /*47577*/;
assign _30232_ = _29540_ ^ _30228_ /*47580*/;
assign _30233_ = _30224_ & _30232_ /*47578*/;
assign _29988_ = _30224_ ^ _30232_ /*47579*/;
assign _30230_ = _30231_ | _30233_ /*47576*/;
assign _30235_ = ~Q[30] /*47575*/;
assign _30234_ = _30235_ & D[36] /*47574*/;
assign _30237_ = _29541_ & _30234_ /*47569*/;
assign _30238_ = _29541_ ^ _30234_ /*47572*/;
assign _30239_ = _30230_ & _30238_ /*47570*/;
assign _29989_ = _30230_ ^ _30238_ /*47571*/;
assign _30236_ = _30237_ | _30239_ /*47568*/;
assign _30241_ = ~Q[30] /*47567*/;
assign _30240_ = _30241_ & D[37] /*47566*/;
assign _30243_ = _29542_ & _30240_ /*47561*/;
assign _30244_ = _29542_ ^ _30240_ /*47564*/;
assign _30245_ = _30236_ & _30244_ /*47562*/;
assign _29990_ = _30236_ ^ _30244_ /*47563*/;
assign _30242_ = _30243_ | _30245_ /*47560*/;
assign _30247_ = ~Q[30] /*47559*/;
assign _30246_ = _30247_ & D[38] /*47558*/;
assign _30249_ = _29543_ & _30246_ /*47553*/;
assign _30250_ = _29543_ ^ _30246_ /*47556*/;
assign _30251_ = _30242_ & _30250_ /*47554*/;
assign _29991_ = _30242_ ^ _30250_ /*47555*/;
assign _30248_ = _30249_ | _30251_ /*47552*/;
assign _30253_ = ~Q[30] /*47551*/;
assign _30252_ = _30253_ & D[39] /*47550*/;
assign _30255_ = _29544_ & _30252_ /*47545*/;
assign _30256_ = _29544_ ^ _30252_ /*47548*/;
assign _30257_ = _30248_ & _30256_ /*47546*/;
assign _29992_ = _30248_ ^ _30256_ /*47547*/;
assign _30254_ = _30255_ | _30257_ /*47544*/;
assign _30259_ = ~Q[30] /*47543*/;
assign _30258_ = _30259_ & D[40] /*47542*/;
assign _30261_ = _29545_ & _30258_ /*47537*/;
assign _30262_ = _29545_ ^ _30258_ /*47540*/;
assign _30263_ = _30254_ & _30262_ /*47538*/;
assign _29993_ = _30254_ ^ _30262_ /*47539*/;
assign _30260_ = _30261_ | _30263_ /*47536*/;
assign _30265_ = ~Q[30] /*47535*/;
assign _30264_ = _30265_ & D[41] /*47534*/;
assign _30267_ = _29546_ & _30264_ /*47529*/;
assign _30268_ = _29546_ ^ _30264_ /*47532*/;
assign _30269_ = _30260_ & _30268_ /*47530*/;
assign _29994_ = _30260_ ^ _30268_ /*47531*/;
assign _30266_ = _30267_ | _30269_ /*47528*/;
assign _30271_ = ~Q[30] /*47527*/;
assign _30270_ = _30271_ & D[42] /*47526*/;
assign _30273_ = _29547_ & _30270_ /*47521*/;
assign _30274_ = _29547_ ^ _30270_ /*47524*/;
assign _30275_ = _30266_ & _30274_ /*47522*/;
assign _29995_ = _30266_ ^ _30274_ /*47523*/;
assign _30272_ = _30273_ | _30275_ /*47520*/;
assign _30277_ = ~Q[30] /*47519*/;
assign _30276_ = _30277_ & D[43] /*47518*/;
assign _30279_ = _29548_ & _30276_ /*47513*/;
assign _30280_ = _29548_ ^ _30276_ /*47516*/;
assign _30281_ = _30272_ & _30280_ /*47514*/;
assign _29996_ = _30272_ ^ _30280_ /*47515*/;
assign _30278_ = _30279_ | _30281_ /*47512*/;
assign _30283_ = ~Q[30] /*47511*/;
assign _30282_ = _30283_ & D[44] /*47510*/;
assign _30285_ = _29549_ & _30282_ /*47505*/;
assign _30286_ = _29549_ ^ _30282_ /*47508*/;
assign _30287_ = _30278_ & _30286_ /*47506*/;
assign _29997_ = _30278_ ^ _30286_ /*47507*/;
assign _30284_ = _30285_ | _30287_ /*47504*/;
assign _30289_ = ~Q[30] /*47503*/;
assign _30288_ = _30289_ & D[45] /*47502*/;
assign _30291_ = _29550_ & _30288_ /*47497*/;
assign _30292_ = _29550_ ^ _30288_ /*47500*/;
assign _30293_ = _30284_ & _30292_ /*47498*/;
assign _29998_ = _30284_ ^ _30292_ /*47499*/;
assign _30290_ = _30291_ | _30293_ /*47496*/;
assign _30295_ = ~Q[30] /*47495*/;
assign _30294_ = _30295_ & D[46] /*47494*/;
assign _30297_ = _29551_ & _30294_ /*47489*/;
assign _30298_ = _29551_ ^ _30294_ /*47492*/;
assign _30299_ = _30290_ & _30298_ /*47490*/;
assign _29999_ = _30290_ ^ _30298_ /*47491*/;
assign _30296_ = _30297_ | _30299_ /*47488*/;
assign _30301_ = ~Q[30] /*47487*/;
assign _30300_ = _30301_ & D[47] /*47486*/;
assign _30303_ = _29552_ & _30300_ /*47481*/;
assign _30304_ = _29552_ ^ _30300_ /*47484*/;
assign _30305_ = _30296_ & _30304_ /*47482*/;
assign _30000_ = _30296_ ^ _30304_ /*47483*/;
assign _30302_ = _30303_ | _30305_ /*47480*/;
assign _30307_ = ~Q[30] /*47479*/;
assign _30306_ = _30307_ & D[48] /*47478*/;
assign _30309_ = _29553_ & _30306_ /*47473*/;
assign _30310_ = _29553_ ^ _30306_ /*47476*/;
assign _30311_ = _30302_ & _30310_ /*47474*/;
assign _30001_ = _30302_ ^ _30310_ /*47475*/;
assign _30308_ = _30309_ | _30311_ /*47472*/;
assign _30313_ = ~Q[30] /*47471*/;
assign _30312_ = _30313_ & D[49] /*47470*/;
assign _30315_ = _29554_ & _30312_ /*47465*/;
assign _30316_ = _29554_ ^ _30312_ /*47468*/;
assign _30317_ = _30308_ & _30316_ /*47466*/;
assign _30002_ = _30308_ ^ _30316_ /*47467*/;
assign _30314_ = _30315_ | _30317_ /*47464*/;
assign _30319_ = ~Q[30] /*47463*/;
assign _30318_ = _30319_ & D[50] /*47462*/;
assign _30321_ = _29555_ & _30318_ /*47457*/;
assign _30322_ = _29555_ ^ _30318_ /*47460*/;
assign _30323_ = _30314_ & _30322_ /*47458*/;
assign _30003_ = _30314_ ^ _30322_ /*47459*/;
assign _30320_ = _30321_ | _30323_ /*47456*/;
assign _30325_ = ~Q[30] /*47455*/;
assign _30324_ = _30325_ & D[51] /*47454*/;
assign _30327_ = _29556_ & _30324_ /*47449*/;
assign _30328_ = _29556_ ^ _30324_ /*47452*/;
assign _30329_ = _30320_ & _30328_ /*47450*/;
assign _30004_ = _30320_ ^ _30328_ /*47451*/;
assign _30326_ = _30327_ | _30329_ /*47448*/;
assign _30331_ = ~Q[30] /*47447*/;
assign _30330_ = _30331_ & D[52] /*47446*/;
assign _30333_ = _29557_ & _30330_ /*47441*/;
assign _30334_ = _29557_ ^ _30330_ /*47444*/;
assign _30335_ = _30326_ & _30334_ /*47442*/;
assign _30005_ = _30326_ ^ _30334_ /*47443*/;
assign _30332_ = _30333_ | _30335_ /*47440*/;
assign _30337_ = ~Q[30] /*47439*/;
assign _30336_ = _30337_ & D[53] /*47438*/;
assign _30339_ = _29558_ & _30336_ /*47433*/;
assign _30340_ = _29558_ ^ _30336_ /*47436*/;
assign _30341_ = _30332_ & _30340_ /*47434*/;
assign _30006_ = _30332_ ^ _30340_ /*47435*/;
assign _30338_ = _30339_ | _30341_ /*47432*/;
assign _30343_ = ~Q[30] /*47431*/;
assign _30342_ = _30343_ & D[54] /*47430*/;
assign _30345_ = _29559_ & _30342_ /*47425*/;
assign _30346_ = _29559_ ^ _30342_ /*47428*/;
assign _30347_ = _30338_ & _30346_ /*47426*/;
assign _30007_ = _30338_ ^ _30346_ /*47427*/;
assign _30344_ = _30345_ | _30347_ /*47424*/;
assign _30349_ = ~Q[30] /*47423*/;
assign _30348_ = _30349_ & D[55] /*47422*/;
assign _30351_ = _29560_ & _30348_ /*47417*/;
assign _30352_ = _29560_ ^ _30348_ /*47420*/;
assign _30353_ = _30344_ & _30352_ /*47418*/;
assign _30008_ = _30344_ ^ _30352_ /*47419*/;
assign _30350_ = _30351_ | _30353_ /*47416*/;
assign _30355_ = ~Q[30] /*47415*/;
assign _30354_ = _30355_ & D[56] /*47414*/;
assign _30357_ = _29561_ & _30354_ /*47409*/;
assign _30358_ = _29561_ ^ _30354_ /*47412*/;
assign _30359_ = _30350_ & _30358_ /*47410*/;
assign _30009_ = _30350_ ^ _30358_ /*47411*/;
assign _30356_ = _30357_ | _30359_ /*47408*/;
assign _30361_ = ~Q[30] /*47407*/;
assign _30360_ = _30361_ & D[57] /*47406*/;
assign _30363_ = _29562_ & _30360_ /*47401*/;
assign _30364_ = _29562_ ^ _30360_ /*47404*/;
assign _30365_ = _30356_ & _30364_ /*47402*/;
assign _30010_ = _30356_ ^ _30364_ /*47403*/;
assign _30362_ = _30363_ | _30365_ /*47400*/;
assign _30367_ = ~Q[30] /*47399*/;
assign _30366_ = _30367_ & D[58] /*47398*/;
assign _30369_ = _29563_ & _30366_ /*47393*/;
assign _30370_ = _29563_ ^ _30366_ /*47396*/;
assign _30371_ = _30362_ & _30370_ /*47394*/;
assign _30011_ = _30362_ ^ _30370_ /*47395*/;
assign _30368_ = _30369_ | _30371_ /*47392*/;
assign _30373_ = ~Q[30] /*47391*/;
assign _30372_ = _30373_ & D[59] /*47390*/;
assign _30375_ = _29564_ & _30372_ /*47385*/;
assign _30376_ = _29564_ ^ _30372_ /*47388*/;
assign _30377_ = _30368_ & _30376_ /*47386*/;
assign _30012_ = _30368_ ^ _30376_ /*47387*/;
assign _30374_ = _30375_ | _30377_ /*47384*/;
assign _30379_ = ~Q[30] /*47383*/;
assign _30378_ = _30379_ & D[60] /*47382*/;
assign _30381_ = _29565_ & _30378_ /*47377*/;
assign _30382_ = _29565_ ^ _30378_ /*47380*/;
assign _30383_ = _30374_ & _30382_ /*47378*/;
assign _30013_ = _30374_ ^ _30382_ /*47379*/;
assign _30380_ = _30381_ | _30383_ /*47376*/;
assign _30385_ = ~Q[30] /*47375*/;
assign _30384_ = _30385_ & D[61] /*47374*/;
assign _30387_ = _29566_ & _30384_ /*47369*/;
assign _30388_ = _29566_ ^ _30384_ /*47372*/;
assign _30389_ = _30380_ & _30388_ /*47370*/;
assign _30014_ = _30380_ ^ _30388_ /*47371*/;
assign _30386_ = _30387_ | _30389_ /*47368*/;
assign _30391_ = ~Q[30] /*47367*/;
assign _30390_ = _30391_ & D[62] /*47366*/;
assign _30393_ = _29567_ & _30390_ /*47361*/;
assign _30394_ = _29567_ ^ _30390_ /*47364*/;
assign _30395_ = _30386_ & _30394_ /*47362*/;
assign _30015_ = _30386_ ^ _30394_ /*47363*/;
assign _30392_ = _30393_ | _30395_ /*47360*/;
assign _30397_ = ~Q[30] /*47359*/;
assign _30396_ = _30397_ & zeroWire /*47358*/;
assign _30398_ = _29568_ ^ _30396_ /*47356*/;
assign _30016_ = _30398_ ^ _30392_ /*47355*/;
assign _30469_ = ~D[0] /*47101*/;
assign _30466_ = R_0[29] & _30469_ /*47097*/;
assign _30467_ = R_0[29] ^ _30469_ /*47100*/;
assign _30468_ = oneWire & _30467_ /*47098*/;
assign _30401_ = oneWire ^ _30467_ /*47099*/;
assign _30465_ = _30466_ | _30468_ /*47096*/;
assign _30474_ = ~D[1] /*47095*/;
assign _30471_ = _29953_ & _30474_ /*47091*/;
assign _30472_ = _29953_ ^ _30474_ /*47094*/;
assign _30473_ = _30465_ & _30472_ /*47092*/;
assign _30402_ = _30465_ ^ _30472_ /*47093*/;
assign _30470_ = _30471_ | _30473_ /*47090*/;
assign _30479_ = ~D[2] /*47089*/;
assign _30476_ = _29954_ & _30479_ /*47085*/;
assign _30477_ = _29954_ ^ _30479_ /*47088*/;
assign _30478_ = _30470_ & _30477_ /*47086*/;
assign _30403_ = _30470_ ^ _30477_ /*47087*/;
assign _30475_ = _30476_ | _30478_ /*47084*/;
assign _30484_ = ~D[3] /*47083*/;
assign _30481_ = _29955_ & _30484_ /*47079*/;
assign _30482_ = _29955_ ^ _30484_ /*47082*/;
assign _30483_ = _30475_ & _30482_ /*47080*/;
assign _30404_ = _30475_ ^ _30482_ /*47081*/;
assign _30480_ = _30481_ | _30483_ /*47078*/;
assign _30489_ = ~D[4] /*47077*/;
assign _30486_ = _29956_ & _30489_ /*47073*/;
assign _30487_ = _29956_ ^ _30489_ /*47076*/;
assign _30488_ = _30480_ & _30487_ /*47074*/;
assign _30405_ = _30480_ ^ _30487_ /*47075*/;
assign _30485_ = _30486_ | _30488_ /*47072*/;
assign _30494_ = ~D[5] /*47071*/;
assign _30491_ = _29957_ & _30494_ /*47067*/;
assign _30492_ = _29957_ ^ _30494_ /*47070*/;
assign _30493_ = _30485_ & _30492_ /*47068*/;
assign _30406_ = _30485_ ^ _30492_ /*47069*/;
assign _30490_ = _30491_ | _30493_ /*47066*/;
assign _30499_ = ~D[6] /*47065*/;
assign _30496_ = _29958_ & _30499_ /*47061*/;
assign _30497_ = _29958_ ^ _30499_ /*47064*/;
assign _30498_ = _30490_ & _30497_ /*47062*/;
assign _30407_ = _30490_ ^ _30497_ /*47063*/;
assign _30495_ = _30496_ | _30498_ /*47060*/;
assign _30504_ = ~D[7] /*47059*/;
assign _30501_ = _29959_ & _30504_ /*47055*/;
assign _30502_ = _29959_ ^ _30504_ /*47058*/;
assign _30503_ = _30495_ & _30502_ /*47056*/;
assign _30408_ = _30495_ ^ _30502_ /*47057*/;
assign _30500_ = _30501_ | _30503_ /*47054*/;
assign _30509_ = ~D[8] /*47053*/;
assign _30506_ = _29960_ & _30509_ /*47049*/;
assign _30507_ = _29960_ ^ _30509_ /*47052*/;
assign _30508_ = _30500_ & _30507_ /*47050*/;
assign _30409_ = _30500_ ^ _30507_ /*47051*/;
assign _30505_ = _30506_ | _30508_ /*47048*/;
assign _30514_ = ~D[9] /*47047*/;
assign _30511_ = _29961_ & _30514_ /*47043*/;
assign _30512_ = _29961_ ^ _30514_ /*47046*/;
assign _30513_ = _30505_ & _30512_ /*47044*/;
assign _30410_ = _30505_ ^ _30512_ /*47045*/;
assign _30510_ = _30511_ | _30513_ /*47042*/;
assign _30519_ = ~D[10] /*47041*/;
assign _30516_ = _29962_ & _30519_ /*47037*/;
assign _30517_ = _29962_ ^ _30519_ /*47040*/;
assign _30518_ = _30510_ & _30517_ /*47038*/;
assign _30411_ = _30510_ ^ _30517_ /*47039*/;
assign _30515_ = _30516_ | _30518_ /*47036*/;
assign _30524_ = ~D[11] /*47035*/;
assign _30521_ = _29963_ & _30524_ /*47031*/;
assign _30522_ = _29963_ ^ _30524_ /*47034*/;
assign _30523_ = _30515_ & _30522_ /*47032*/;
assign _30412_ = _30515_ ^ _30522_ /*47033*/;
assign _30520_ = _30521_ | _30523_ /*47030*/;
assign _30529_ = ~D[12] /*47029*/;
assign _30526_ = _29964_ & _30529_ /*47025*/;
assign _30527_ = _29964_ ^ _30529_ /*47028*/;
assign _30528_ = _30520_ & _30527_ /*47026*/;
assign _30413_ = _30520_ ^ _30527_ /*47027*/;
assign _30525_ = _30526_ | _30528_ /*47024*/;
assign _30534_ = ~D[13] /*47023*/;
assign _30531_ = _29965_ & _30534_ /*47019*/;
assign _30532_ = _29965_ ^ _30534_ /*47022*/;
assign _30533_ = _30525_ & _30532_ /*47020*/;
assign _30414_ = _30525_ ^ _30532_ /*47021*/;
assign _30530_ = _30531_ | _30533_ /*47018*/;
assign _30539_ = ~D[14] /*47017*/;
assign _30536_ = _29966_ & _30539_ /*47013*/;
assign _30537_ = _29966_ ^ _30539_ /*47016*/;
assign _30538_ = _30530_ & _30537_ /*47014*/;
assign _30415_ = _30530_ ^ _30537_ /*47015*/;
assign _30535_ = _30536_ | _30538_ /*47012*/;
assign _30544_ = ~D[15] /*47011*/;
assign _30541_ = _29967_ & _30544_ /*47007*/;
assign _30542_ = _29967_ ^ _30544_ /*47010*/;
assign _30543_ = _30535_ & _30542_ /*47008*/;
assign _30416_ = _30535_ ^ _30542_ /*47009*/;
assign _30540_ = _30541_ | _30543_ /*47006*/;
assign _30549_ = ~D[16] /*47005*/;
assign _30546_ = _29968_ & _30549_ /*47001*/;
assign _30547_ = _29968_ ^ _30549_ /*47004*/;
assign _30548_ = _30540_ & _30547_ /*47002*/;
assign _30417_ = _30540_ ^ _30547_ /*47003*/;
assign _30545_ = _30546_ | _30548_ /*47000*/;
assign _30554_ = ~D[17] /*46999*/;
assign _30551_ = _29969_ & _30554_ /*46995*/;
assign _30552_ = _29969_ ^ _30554_ /*46998*/;
assign _30553_ = _30545_ & _30552_ /*46996*/;
assign _30418_ = _30545_ ^ _30552_ /*46997*/;
assign _30550_ = _30551_ | _30553_ /*46994*/;
assign _30559_ = ~D[18] /*46993*/;
assign _30556_ = _29970_ & _30559_ /*46989*/;
assign _30557_ = _29970_ ^ _30559_ /*46992*/;
assign _30558_ = _30550_ & _30557_ /*46990*/;
assign _30419_ = _30550_ ^ _30557_ /*46991*/;
assign _30555_ = _30556_ | _30558_ /*46988*/;
assign _30564_ = ~D[19] /*46987*/;
assign _30561_ = _29971_ & _30564_ /*46983*/;
assign _30562_ = _29971_ ^ _30564_ /*46986*/;
assign _30563_ = _30555_ & _30562_ /*46984*/;
assign _30420_ = _30555_ ^ _30562_ /*46985*/;
assign _30560_ = _30561_ | _30563_ /*46982*/;
assign _30569_ = ~D[20] /*46981*/;
assign _30566_ = _29972_ & _30569_ /*46977*/;
assign _30567_ = _29972_ ^ _30569_ /*46980*/;
assign _30568_ = _30560_ & _30567_ /*46978*/;
assign _30421_ = _30560_ ^ _30567_ /*46979*/;
assign _30565_ = _30566_ | _30568_ /*46976*/;
assign _30574_ = ~D[21] /*46975*/;
assign _30571_ = _29973_ & _30574_ /*46971*/;
assign _30572_ = _29973_ ^ _30574_ /*46974*/;
assign _30573_ = _30565_ & _30572_ /*46972*/;
assign _30422_ = _30565_ ^ _30572_ /*46973*/;
assign _30570_ = _30571_ | _30573_ /*46970*/;
assign _30579_ = ~D[22] /*46969*/;
assign _30576_ = _29974_ & _30579_ /*46965*/;
assign _30577_ = _29974_ ^ _30579_ /*46968*/;
assign _30578_ = _30570_ & _30577_ /*46966*/;
assign _30423_ = _30570_ ^ _30577_ /*46967*/;
assign _30575_ = _30576_ | _30578_ /*46964*/;
assign _30584_ = ~D[23] /*46963*/;
assign _30581_ = _29975_ & _30584_ /*46959*/;
assign _30582_ = _29975_ ^ _30584_ /*46962*/;
assign _30583_ = _30575_ & _30582_ /*46960*/;
assign _30424_ = _30575_ ^ _30582_ /*46961*/;
assign _30580_ = _30581_ | _30583_ /*46958*/;
assign _30589_ = ~D[24] /*46957*/;
assign _30586_ = _29976_ & _30589_ /*46953*/;
assign _30587_ = _29976_ ^ _30589_ /*46956*/;
assign _30588_ = _30580_ & _30587_ /*46954*/;
assign _30425_ = _30580_ ^ _30587_ /*46955*/;
assign _30585_ = _30586_ | _30588_ /*46952*/;
assign _30594_ = ~D[25] /*46951*/;
assign _30591_ = _29977_ & _30594_ /*46947*/;
assign _30592_ = _29977_ ^ _30594_ /*46950*/;
assign _30593_ = _30585_ & _30592_ /*46948*/;
assign _30426_ = _30585_ ^ _30592_ /*46949*/;
assign _30590_ = _30591_ | _30593_ /*46946*/;
assign _30599_ = ~D[26] /*46945*/;
assign _30596_ = _29978_ & _30599_ /*46941*/;
assign _30597_ = _29978_ ^ _30599_ /*46944*/;
assign _30598_ = _30590_ & _30597_ /*46942*/;
assign _30427_ = _30590_ ^ _30597_ /*46943*/;
assign _30595_ = _30596_ | _30598_ /*46940*/;
assign _30604_ = ~D[27] /*46939*/;
assign _30601_ = _29979_ & _30604_ /*46935*/;
assign _30602_ = _29979_ ^ _30604_ /*46938*/;
assign _30603_ = _30595_ & _30602_ /*46936*/;
assign _30428_ = _30595_ ^ _30602_ /*46937*/;
assign _30600_ = _30601_ | _30603_ /*46934*/;
assign _30609_ = ~D[28] /*46933*/;
assign _30606_ = _29980_ & _30609_ /*46929*/;
assign _30607_ = _29980_ ^ _30609_ /*46932*/;
assign _30608_ = _30600_ & _30607_ /*46930*/;
assign _30429_ = _30600_ ^ _30607_ /*46931*/;
assign _30605_ = _30606_ | _30608_ /*46928*/;
assign _30614_ = ~D[29] /*46927*/;
assign _30611_ = _29981_ & _30614_ /*46923*/;
assign _30612_ = _29981_ ^ _30614_ /*46926*/;
assign _30613_ = _30605_ & _30612_ /*46924*/;
assign _30430_ = _30605_ ^ _30612_ /*46925*/;
assign _30610_ = _30611_ | _30613_ /*46922*/;
assign _30619_ = ~D[30] /*46921*/;
assign _30616_ = _29982_ & _30619_ /*46917*/;
assign _30617_ = _29982_ ^ _30619_ /*46920*/;
assign _30618_ = _30610_ & _30617_ /*46918*/;
assign _30431_ = _30610_ ^ _30617_ /*46919*/;
assign _30615_ = _30616_ | _30618_ /*46916*/;
assign _30624_ = ~D[31] /*46915*/;
assign _30621_ = _29983_ & _30624_ /*46911*/;
assign _30622_ = _29983_ ^ _30624_ /*46914*/;
assign _30623_ = _30615_ & _30622_ /*46912*/;
assign _30432_ = _30615_ ^ _30622_ /*46913*/;
assign _30620_ = _30621_ | _30623_ /*46910*/;
assign _30629_ = ~D[32] /*46909*/;
assign _30626_ = _29984_ & _30629_ /*46905*/;
assign _30627_ = _29984_ ^ _30629_ /*46908*/;
assign _30628_ = _30620_ & _30627_ /*46906*/;
assign _30433_ = _30620_ ^ _30627_ /*46907*/;
assign _30625_ = _30626_ | _30628_ /*46904*/;
assign _30634_ = ~D[33] /*46903*/;
assign _30631_ = _29985_ & _30634_ /*46899*/;
assign _30632_ = _29985_ ^ _30634_ /*46902*/;
assign _30633_ = _30625_ & _30632_ /*46900*/;
assign _30434_ = _30625_ ^ _30632_ /*46901*/;
assign _30630_ = _30631_ | _30633_ /*46898*/;
assign _30639_ = ~D[34] /*46897*/;
assign _30636_ = _29986_ & _30639_ /*46893*/;
assign _30637_ = _29986_ ^ _30639_ /*46896*/;
assign _30638_ = _30630_ & _30637_ /*46894*/;
assign _30435_ = _30630_ ^ _30637_ /*46895*/;
assign _30635_ = _30636_ | _30638_ /*46892*/;
assign _30644_ = ~D[35] /*46891*/;
assign _30641_ = _29987_ & _30644_ /*46887*/;
assign _30642_ = _29987_ ^ _30644_ /*46890*/;
assign _30643_ = _30635_ & _30642_ /*46888*/;
assign _30436_ = _30635_ ^ _30642_ /*46889*/;
assign _30640_ = _30641_ | _30643_ /*46886*/;
assign _30649_ = ~D[36] /*46885*/;
assign _30646_ = _29988_ & _30649_ /*46881*/;
assign _30647_ = _29988_ ^ _30649_ /*46884*/;
assign _30648_ = _30640_ & _30647_ /*46882*/;
assign _30437_ = _30640_ ^ _30647_ /*46883*/;
assign _30645_ = _30646_ | _30648_ /*46880*/;
assign _30654_ = ~D[37] /*46879*/;
assign _30651_ = _29989_ & _30654_ /*46875*/;
assign _30652_ = _29989_ ^ _30654_ /*46878*/;
assign _30653_ = _30645_ & _30652_ /*46876*/;
assign _30438_ = _30645_ ^ _30652_ /*46877*/;
assign _30650_ = _30651_ | _30653_ /*46874*/;
assign _30659_ = ~D[38] /*46873*/;
assign _30656_ = _29990_ & _30659_ /*46869*/;
assign _30657_ = _29990_ ^ _30659_ /*46872*/;
assign _30658_ = _30650_ & _30657_ /*46870*/;
assign _30439_ = _30650_ ^ _30657_ /*46871*/;
assign _30655_ = _30656_ | _30658_ /*46868*/;
assign _30664_ = ~D[39] /*46867*/;
assign _30661_ = _29991_ & _30664_ /*46863*/;
assign _30662_ = _29991_ ^ _30664_ /*46866*/;
assign _30663_ = _30655_ & _30662_ /*46864*/;
assign _30440_ = _30655_ ^ _30662_ /*46865*/;
assign _30660_ = _30661_ | _30663_ /*46862*/;
assign _30669_ = ~D[40] /*46861*/;
assign _30666_ = _29992_ & _30669_ /*46857*/;
assign _30667_ = _29992_ ^ _30669_ /*46860*/;
assign _30668_ = _30660_ & _30667_ /*46858*/;
assign _30441_ = _30660_ ^ _30667_ /*46859*/;
assign _30665_ = _30666_ | _30668_ /*46856*/;
assign _30674_ = ~D[41] /*46855*/;
assign _30671_ = _29993_ & _30674_ /*46851*/;
assign _30672_ = _29993_ ^ _30674_ /*46854*/;
assign _30673_ = _30665_ & _30672_ /*46852*/;
assign _30442_ = _30665_ ^ _30672_ /*46853*/;
assign _30670_ = _30671_ | _30673_ /*46850*/;
assign _30679_ = ~D[42] /*46849*/;
assign _30676_ = _29994_ & _30679_ /*46845*/;
assign _30677_ = _29994_ ^ _30679_ /*46848*/;
assign _30678_ = _30670_ & _30677_ /*46846*/;
assign _30443_ = _30670_ ^ _30677_ /*46847*/;
assign _30675_ = _30676_ | _30678_ /*46844*/;
assign _30684_ = ~D[43] /*46843*/;
assign _30681_ = _29995_ & _30684_ /*46839*/;
assign _30682_ = _29995_ ^ _30684_ /*46842*/;
assign _30683_ = _30675_ & _30682_ /*46840*/;
assign _30444_ = _30675_ ^ _30682_ /*46841*/;
assign _30680_ = _30681_ | _30683_ /*46838*/;
assign _30689_ = ~D[44] /*46837*/;
assign _30686_ = _29996_ & _30689_ /*46833*/;
assign _30687_ = _29996_ ^ _30689_ /*46836*/;
assign _30688_ = _30680_ & _30687_ /*46834*/;
assign _30445_ = _30680_ ^ _30687_ /*46835*/;
assign _30685_ = _30686_ | _30688_ /*46832*/;
assign _30694_ = ~D[45] /*46831*/;
assign _30691_ = _29997_ & _30694_ /*46827*/;
assign _30692_ = _29997_ ^ _30694_ /*46830*/;
assign _30693_ = _30685_ & _30692_ /*46828*/;
assign _30446_ = _30685_ ^ _30692_ /*46829*/;
assign _30690_ = _30691_ | _30693_ /*46826*/;
assign _30699_ = ~D[46] /*46825*/;
assign _30696_ = _29998_ & _30699_ /*46821*/;
assign _30697_ = _29998_ ^ _30699_ /*46824*/;
assign _30698_ = _30690_ & _30697_ /*46822*/;
assign _30447_ = _30690_ ^ _30697_ /*46823*/;
assign _30695_ = _30696_ | _30698_ /*46820*/;
assign _30704_ = ~D[47] /*46819*/;
assign _30701_ = _29999_ & _30704_ /*46815*/;
assign _30702_ = _29999_ ^ _30704_ /*46818*/;
assign _30703_ = _30695_ & _30702_ /*46816*/;
assign _30448_ = _30695_ ^ _30702_ /*46817*/;
assign _30700_ = _30701_ | _30703_ /*46814*/;
assign _30709_ = ~D[48] /*46813*/;
assign _30706_ = _30000_ & _30709_ /*46809*/;
assign _30707_ = _30000_ ^ _30709_ /*46812*/;
assign _30708_ = _30700_ & _30707_ /*46810*/;
assign _30449_ = _30700_ ^ _30707_ /*46811*/;
assign _30705_ = _30706_ | _30708_ /*46808*/;
assign _30714_ = ~D[49] /*46807*/;
assign _30711_ = _30001_ & _30714_ /*46803*/;
assign _30712_ = _30001_ ^ _30714_ /*46806*/;
assign _30713_ = _30705_ & _30712_ /*46804*/;
assign _30450_ = _30705_ ^ _30712_ /*46805*/;
assign _30710_ = _30711_ | _30713_ /*46802*/;
assign _30719_ = ~D[50] /*46801*/;
assign _30716_ = _30002_ & _30719_ /*46797*/;
assign _30717_ = _30002_ ^ _30719_ /*46800*/;
assign _30718_ = _30710_ & _30717_ /*46798*/;
assign _30451_ = _30710_ ^ _30717_ /*46799*/;
assign _30715_ = _30716_ | _30718_ /*46796*/;
assign _30724_ = ~D[51] /*46795*/;
assign _30721_ = _30003_ & _30724_ /*46791*/;
assign _30722_ = _30003_ ^ _30724_ /*46794*/;
assign _30723_ = _30715_ & _30722_ /*46792*/;
assign _30452_ = _30715_ ^ _30722_ /*46793*/;
assign _30720_ = _30721_ | _30723_ /*46790*/;
assign _30729_ = ~D[52] /*46789*/;
assign _30726_ = _30004_ & _30729_ /*46785*/;
assign _30727_ = _30004_ ^ _30729_ /*46788*/;
assign _30728_ = _30720_ & _30727_ /*46786*/;
assign _30453_ = _30720_ ^ _30727_ /*46787*/;
assign _30725_ = _30726_ | _30728_ /*46784*/;
assign _30734_ = ~D[53] /*46783*/;
assign _30731_ = _30005_ & _30734_ /*46779*/;
assign _30732_ = _30005_ ^ _30734_ /*46782*/;
assign _30733_ = _30725_ & _30732_ /*46780*/;
assign _30454_ = _30725_ ^ _30732_ /*46781*/;
assign _30730_ = _30731_ | _30733_ /*46778*/;
assign _30739_ = ~D[54] /*46777*/;
assign _30736_ = _30006_ & _30739_ /*46773*/;
assign _30737_ = _30006_ ^ _30739_ /*46776*/;
assign _30738_ = _30730_ & _30737_ /*46774*/;
assign _30455_ = _30730_ ^ _30737_ /*46775*/;
assign _30735_ = _30736_ | _30738_ /*46772*/;
assign _30744_ = ~D[55] /*46771*/;
assign _30741_ = _30007_ & _30744_ /*46767*/;
assign _30742_ = _30007_ ^ _30744_ /*46770*/;
assign _30743_ = _30735_ & _30742_ /*46768*/;
assign _30456_ = _30735_ ^ _30742_ /*46769*/;
assign _30740_ = _30741_ | _30743_ /*46766*/;
assign _30749_ = ~D[56] /*46765*/;
assign _30746_ = _30008_ & _30749_ /*46761*/;
assign _30747_ = _30008_ ^ _30749_ /*46764*/;
assign _30748_ = _30740_ & _30747_ /*46762*/;
assign _30457_ = _30740_ ^ _30747_ /*46763*/;
assign _30745_ = _30746_ | _30748_ /*46760*/;
assign _30754_ = ~D[57] /*46759*/;
assign _30751_ = _30009_ & _30754_ /*46755*/;
assign _30752_ = _30009_ ^ _30754_ /*46758*/;
assign _30753_ = _30745_ & _30752_ /*46756*/;
assign _30458_ = _30745_ ^ _30752_ /*46757*/;
assign _30750_ = _30751_ | _30753_ /*46754*/;
assign _30759_ = ~D[58] /*46753*/;
assign _30756_ = _30010_ & _30759_ /*46749*/;
assign _30757_ = _30010_ ^ _30759_ /*46752*/;
assign _30758_ = _30750_ & _30757_ /*46750*/;
assign _30459_ = _30750_ ^ _30757_ /*46751*/;
assign _30755_ = _30756_ | _30758_ /*46748*/;
assign _30764_ = ~D[59] /*46747*/;
assign _30761_ = _30011_ & _30764_ /*46743*/;
assign _30762_ = _30011_ ^ _30764_ /*46746*/;
assign _30763_ = _30755_ & _30762_ /*46744*/;
assign _30460_ = _30755_ ^ _30762_ /*46745*/;
assign _30760_ = _30761_ | _30763_ /*46742*/;
assign _30769_ = ~D[60] /*46741*/;
assign _30766_ = _30012_ & _30769_ /*46737*/;
assign _30767_ = _30012_ ^ _30769_ /*46740*/;
assign _30768_ = _30760_ & _30767_ /*46738*/;
assign _30461_ = _30760_ ^ _30767_ /*46739*/;
assign _30765_ = _30766_ | _30768_ /*46736*/;
assign _30774_ = ~D[61] /*46735*/;
assign _30771_ = _30013_ & _30774_ /*46731*/;
assign _30772_ = _30013_ ^ _30774_ /*46734*/;
assign _30773_ = _30765_ & _30772_ /*46732*/;
assign _30462_ = _30765_ ^ _30772_ /*46733*/;
assign _30770_ = _30771_ | _30773_ /*46730*/;
assign _30779_ = ~D[62] /*46729*/;
assign _30776_ = _30014_ & _30779_ /*46725*/;
assign _30777_ = _30014_ ^ _30779_ /*46728*/;
assign _30778_ = _30770_ & _30777_ /*46726*/;
assign _30463_ = _30770_ ^ _30777_ /*46727*/;
assign _30775_ = _30776_ | _30778_ /*46724*/;
assign _30780_ = _30015_ & oneWire /*46719*/;
assign _30781_ = _30015_ ^ oneWire /*46722*/;
assign _30782_ = _30775_ & _30781_ /*46720*/;
assign _30464_ = _30775_ ^ _30781_ /*46721*/;
assign Q[29] = _30780_ | _30782_ /*46718*/;
assign _30915_ = ~Q[29] /*46333*/;
assign _30914_ = _30915_ & D[0] /*46332*/;
assign _30917_ = _30401_ & _30914_ /*46327*/;
assign _30918_ = _30401_ ^ _30914_ /*46330*/;
assign _30919_ = zeroWire & _30918_ /*46328*/;
assign _30849_ = zeroWire ^ _30918_ /*46329*/;
assign _30916_ = _30917_ | _30919_ /*46326*/;
assign _30921_ = ~Q[29] /*46325*/;
assign _30920_ = _30921_ & D[1] /*46324*/;
assign _30923_ = _30402_ & _30920_ /*46319*/;
assign _30924_ = _30402_ ^ _30920_ /*46322*/;
assign _30925_ = _30916_ & _30924_ /*46320*/;
assign _30850_ = _30916_ ^ _30924_ /*46321*/;
assign _30922_ = _30923_ | _30925_ /*46318*/;
assign _30927_ = ~Q[29] /*46317*/;
assign _30926_ = _30927_ & D[2] /*46316*/;
assign _30929_ = _30403_ & _30926_ /*46311*/;
assign _30930_ = _30403_ ^ _30926_ /*46314*/;
assign _30931_ = _30922_ & _30930_ /*46312*/;
assign _30851_ = _30922_ ^ _30930_ /*46313*/;
assign _30928_ = _30929_ | _30931_ /*46310*/;
assign _30933_ = ~Q[29] /*46309*/;
assign _30932_ = _30933_ & D[3] /*46308*/;
assign _30935_ = _30404_ & _30932_ /*46303*/;
assign _30936_ = _30404_ ^ _30932_ /*46306*/;
assign _30937_ = _30928_ & _30936_ /*46304*/;
assign _30852_ = _30928_ ^ _30936_ /*46305*/;
assign _30934_ = _30935_ | _30937_ /*46302*/;
assign _30939_ = ~Q[29] /*46301*/;
assign _30938_ = _30939_ & D[4] /*46300*/;
assign _30941_ = _30405_ & _30938_ /*46295*/;
assign _30942_ = _30405_ ^ _30938_ /*46298*/;
assign _30943_ = _30934_ & _30942_ /*46296*/;
assign _30853_ = _30934_ ^ _30942_ /*46297*/;
assign _30940_ = _30941_ | _30943_ /*46294*/;
assign _30945_ = ~Q[29] /*46293*/;
assign _30944_ = _30945_ & D[5] /*46292*/;
assign _30947_ = _30406_ & _30944_ /*46287*/;
assign _30948_ = _30406_ ^ _30944_ /*46290*/;
assign _30949_ = _30940_ & _30948_ /*46288*/;
assign _30854_ = _30940_ ^ _30948_ /*46289*/;
assign _30946_ = _30947_ | _30949_ /*46286*/;
assign _30951_ = ~Q[29] /*46285*/;
assign _30950_ = _30951_ & D[6] /*46284*/;
assign _30953_ = _30407_ & _30950_ /*46279*/;
assign _30954_ = _30407_ ^ _30950_ /*46282*/;
assign _30955_ = _30946_ & _30954_ /*46280*/;
assign _30855_ = _30946_ ^ _30954_ /*46281*/;
assign _30952_ = _30953_ | _30955_ /*46278*/;
assign _30957_ = ~Q[29] /*46277*/;
assign _30956_ = _30957_ & D[7] /*46276*/;
assign _30959_ = _30408_ & _30956_ /*46271*/;
assign _30960_ = _30408_ ^ _30956_ /*46274*/;
assign _30961_ = _30952_ & _30960_ /*46272*/;
assign _30856_ = _30952_ ^ _30960_ /*46273*/;
assign _30958_ = _30959_ | _30961_ /*46270*/;
assign _30963_ = ~Q[29] /*46269*/;
assign _30962_ = _30963_ & D[8] /*46268*/;
assign _30965_ = _30409_ & _30962_ /*46263*/;
assign _30966_ = _30409_ ^ _30962_ /*46266*/;
assign _30967_ = _30958_ & _30966_ /*46264*/;
assign _30857_ = _30958_ ^ _30966_ /*46265*/;
assign _30964_ = _30965_ | _30967_ /*46262*/;
assign _30969_ = ~Q[29] /*46261*/;
assign _30968_ = _30969_ & D[9] /*46260*/;
assign _30971_ = _30410_ & _30968_ /*46255*/;
assign _30972_ = _30410_ ^ _30968_ /*46258*/;
assign _30973_ = _30964_ & _30972_ /*46256*/;
assign _30858_ = _30964_ ^ _30972_ /*46257*/;
assign _30970_ = _30971_ | _30973_ /*46254*/;
assign _30975_ = ~Q[29] /*46253*/;
assign _30974_ = _30975_ & D[10] /*46252*/;
assign _30977_ = _30411_ & _30974_ /*46247*/;
assign _30978_ = _30411_ ^ _30974_ /*46250*/;
assign _30979_ = _30970_ & _30978_ /*46248*/;
assign _30859_ = _30970_ ^ _30978_ /*46249*/;
assign _30976_ = _30977_ | _30979_ /*46246*/;
assign _30981_ = ~Q[29] /*46245*/;
assign _30980_ = _30981_ & D[11] /*46244*/;
assign _30983_ = _30412_ & _30980_ /*46239*/;
assign _30984_ = _30412_ ^ _30980_ /*46242*/;
assign _30985_ = _30976_ & _30984_ /*46240*/;
assign _30860_ = _30976_ ^ _30984_ /*46241*/;
assign _30982_ = _30983_ | _30985_ /*46238*/;
assign _30987_ = ~Q[29] /*46237*/;
assign _30986_ = _30987_ & D[12] /*46236*/;
assign _30989_ = _30413_ & _30986_ /*46231*/;
assign _30990_ = _30413_ ^ _30986_ /*46234*/;
assign _30991_ = _30982_ & _30990_ /*46232*/;
assign _30861_ = _30982_ ^ _30990_ /*46233*/;
assign _30988_ = _30989_ | _30991_ /*46230*/;
assign _30993_ = ~Q[29] /*46229*/;
assign _30992_ = _30993_ & D[13] /*46228*/;
assign _30995_ = _30414_ & _30992_ /*46223*/;
assign _30996_ = _30414_ ^ _30992_ /*46226*/;
assign _30997_ = _30988_ & _30996_ /*46224*/;
assign _30862_ = _30988_ ^ _30996_ /*46225*/;
assign _30994_ = _30995_ | _30997_ /*46222*/;
assign _30999_ = ~Q[29] /*46221*/;
assign _30998_ = _30999_ & D[14] /*46220*/;
assign _31001_ = _30415_ & _30998_ /*46215*/;
assign _31002_ = _30415_ ^ _30998_ /*46218*/;
assign _31003_ = _30994_ & _31002_ /*46216*/;
assign _30863_ = _30994_ ^ _31002_ /*46217*/;
assign _31000_ = _31001_ | _31003_ /*46214*/;
assign _31005_ = ~Q[29] /*46213*/;
assign _31004_ = _31005_ & D[15] /*46212*/;
assign _31007_ = _30416_ & _31004_ /*46207*/;
assign _31008_ = _30416_ ^ _31004_ /*46210*/;
assign _31009_ = _31000_ & _31008_ /*46208*/;
assign _30864_ = _31000_ ^ _31008_ /*46209*/;
assign _31006_ = _31007_ | _31009_ /*46206*/;
assign _31011_ = ~Q[29] /*46205*/;
assign _31010_ = _31011_ & D[16] /*46204*/;
assign _31013_ = _30417_ & _31010_ /*46199*/;
assign _31014_ = _30417_ ^ _31010_ /*46202*/;
assign _31015_ = _31006_ & _31014_ /*46200*/;
assign _30865_ = _31006_ ^ _31014_ /*46201*/;
assign _31012_ = _31013_ | _31015_ /*46198*/;
assign _31017_ = ~Q[29] /*46197*/;
assign _31016_ = _31017_ & D[17] /*46196*/;
assign _31019_ = _30418_ & _31016_ /*46191*/;
assign _31020_ = _30418_ ^ _31016_ /*46194*/;
assign _31021_ = _31012_ & _31020_ /*46192*/;
assign _30866_ = _31012_ ^ _31020_ /*46193*/;
assign _31018_ = _31019_ | _31021_ /*46190*/;
assign _31023_ = ~Q[29] /*46189*/;
assign _31022_ = _31023_ & D[18] /*46188*/;
assign _31025_ = _30419_ & _31022_ /*46183*/;
assign _31026_ = _30419_ ^ _31022_ /*46186*/;
assign _31027_ = _31018_ & _31026_ /*46184*/;
assign _30867_ = _31018_ ^ _31026_ /*46185*/;
assign _31024_ = _31025_ | _31027_ /*46182*/;
assign _31029_ = ~Q[29] /*46181*/;
assign _31028_ = _31029_ & D[19] /*46180*/;
assign _31031_ = _30420_ & _31028_ /*46175*/;
assign _31032_ = _30420_ ^ _31028_ /*46178*/;
assign _31033_ = _31024_ & _31032_ /*46176*/;
assign _30868_ = _31024_ ^ _31032_ /*46177*/;
assign _31030_ = _31031_ | _31033_ /*46174*/;
assign _31035_ = ~Q[29] /*46173*/;
assign _31034_ = _31035_ & D[20] /*46172*/;
assign _31037_ = _30421_ & _31034_ /*46167*/;
assign _31038_ = _30421_ ^ _31034_ /*46170*/;
assign _31039_ = _31030_ & _31038_ /*46168*/;
assign _30869_ = _31030_ ^ _31038_ /*46169*/;
assign _31036_ = _31037_ | _31039_ /*46166*/;
assign _31041_ = ~Q[29] /*46165*/;
assign _31040_ = _31041_ & D[21] /*46164*/;
assign _31043_ = _30422_ & _31040_ /*46159*/;
assign _31044_ = _30422_ ^ _31040_ /*46162*/;
assign _31045_ = _31036_ & _31044_ /*46160*/;
assign _30870_ = _31036_ ^ _31044_ /*46161*/;
assign _31042_ = _31043_ | _31045_ /*46158*/;
assign _31047_ = ~Q[29] /*46157*/;
assign _31046_ = _31047_ & D[22] /*46156*/;
assign _31049_ = _30423_ & _31046_ /*46151*/;
assign _31050_ = _30423_ ^ _31046_ /*46154*/;
assign _31051_ = _31042_ & _31050_ /*46152*/;
assign _30871_ = _31042_ ^ _31050_ /*46153*/;
assign _31048_ = _31049_ | _31051_ /*46150*/;
assign _31053_ = ~Q[29] /*46149*/;
assign _31052_ = _31053_ & D[23] /*46148*/;
assign _31055_ = _30424_ & _31052_ /*46143*/;
assign _31056_ = _30424_ ^ _31052_ /*46146*/;
assign _31057_ = _31048_ & _31056_ /*46144*/;
assign _30872_ = _31048_ ^ _31056_ /*46145*/;
assign _31054_ = _31055_ | _31057_ /*46142*/;
assign _31059_ = ~Q[29] /*46141*/;
assign _31058_ = _31059_ & D[24] /*46140*/;
assign _31061_ = _30425_ & _31058_ /*46135*/;
assign _31062_ = _30425_ ^ _31058_ /*46138*/;
assign _31063_ = _31054_ & _31062_ /*46136*/;
assign _30873_ = _31054_ ^ _31062_ /*46137*/;
assign _31060_ = _31061_ | _31063_ /*46134*/;
assign _31065_ = ~Q[29] /*46133*/;
assign _31064_ = _31065_ & D[25] /*46132*/;
assign _31067_ = _30426_ & _31064_ /*46127*/;
assign _31068_ = _30426_ ^ _31064_ /*46130*/;
assign _31069_ = _31060_ & _31068_ /*46128*/;
assign _30874_ = _31060_ ^ _31068_ /*46129*/;
assign _31066_ = _31067_ | _31069_ /*46126*/;
assign _31071_ = ~Q[29] /*46125*/;
assign _31070_ = _31071_ & D[26] /*46124*/;
assign _31073_ = _30427_ & _31070_ /*46119*/;
assign _31074_ = _30427_ ^ _31070_ /*46122*/;
assign _31075_ = _31066_ & _31074_ /*46120*/;
assign _30875_ = _31066_ ^ _31074_ /*46121*/;
assign _31072_ = _31073_ | _31075_ /*46118*/;
assign _31077_ = ~Q[29] /*46117*/;
assign _31076_ = _31077_ & D[27] /*46116*/;
assign _31079_ = _30428_ & _31076_ /*46111*/;
assign _31080_ = _30428_ ^ _31076_ /*46114*/;
assign _31081_ = _31072_ & _31080_ /*46112*/;
assign _30876_ = _31072_ ^ _31080_ /*46113*/;
assign _31078_ = _31079_ | _31081_ /*46110*/;
assign _31083_ = ~Q[29] /*46109*/;
assign _31082_ = _31083_ & D[28] /*46108*/;
assign _31085_ = _30429_ & _31082_ /*46103*/;
assign _31086_ = _30429_ ^ _31082_ /*46106*/;
assign _31087_ = _31078_ & _31086_ /*46104*/;
assign _30877_ = _31078_ ^ _31086_ /*46105*/;
assign _31084_ = _31085_ | _31087_ /*46102*/;
assign _31089_ = ~Q[29] /*46101*/;
assign _31088_ = _31089_ & D[29] /*46100*/;
assign _31091_ = _30430_ & _31088_ /*46095*/;
assign _31092_ = _30430_ ^ _31088_ /*46098*/;
assign _31093_ = _31084_ & _31092_ /*46096*/;
assign _30878_ = _31084_ ^ _31092_ /*46097*/;
assign _31090_ = _31091_ | _31093_ /*46094*/;
assign _31095_ = ~Q[29] /*46093*/;
assign _31094_ = _31095_ & D[30] /*46092*/;
assign _31097_ = _30431_ & _31094_ /*46087*/;
assign _31098_ = _30431_ ^ _31094_ /*46090*/;
assign _31099_ = _31090_ & _31098_ /*46088*/;
assign _30879_ = _31090_ ^ _31098_ /*46089*/;
assign _31096_ = _31097_ | _31099_ /*46086*/;
assign _31101_ = ~Q[29] /*46085*/;
assign _31100_ = _31101_ & D[31] /*46084*/;
assign _31103_ = _30432_ & _31100_ /*46079*/;
assign _31104_ = _30432_ ^ _31100_ /*46082*/;
assign _31105_ = _31096_ & _31104_ /*46080*/;
assign _30880_ = _31096_ ^ _31104_ /*46081*/;
assign _31102_ = _31103_ | _31105_ /*46078*/;
assign _31107_ = ~Q[29] /*46077*/;
assign _31106_ = _31107_ & D[32] /*46076*/;
assign _31109_ = _30433_ & _31106_ /*46071*/;
assign _31110_ = _30433_ ^ _31106_ /*46074*/;
assign _31111_ = _31102_ & _31110_ /*46072*/;
assign _30881_ = _31102_ ^ _31110_ /*46073*/;
assign _31108_ = _31109_ | _31111_ /*46070*/;
assign _31113_ = ~Q[29] /*46069*/;
assign _31112_ = _31113_ & D[33] /*46068*/;
assign _31115_ = _30434_ & _31112_ /*46063*/;
assign _31116_ = _30434_ ^ _31112_ /*46066*/;
assign _31117_ = _31108_ & _31116_ /*46064*/;
assign _30882_ = _31108_ ^ _31116_ /*46065*/;
assign _31114_ = _31115_ | _31117_ /*46062*/;
assign _31119_ = ~Q[29] /*46061*/;
assign _31118_ = _31119_ & D[34] /*46060*/;
assign _31121_ = _30435_ & _31118_ /*46055*/;
assign _31122_ = _30435_ ^ _31118_ /*46058*/;
assign _31123_ = _31114_ & _31122_ /*46056*/;
assign _30883_ = _31114_ ^ _31122_ /*46057*/;
assign _31120_ = _31121_ | _31123_ /*46054*/;
assign _31125_ = ~Q[29] /*46053*/;
assign _31124_ = _31125_ & D[35] /*46052*/;
assign _31127_ = _30436_ & _31124_ /*46047*/;
assign _31128_ = _30436_ ^ _31124_ /*46050*/;
assign _31129_ = _31120_ & _31128_ /*46048*/;
assign _30884_ = _31120_ ^ _31128_ /*46049*/;
assign _31126_ = _31127_ | _31129_ /*46046*/;
assign _31131_ = ~Q[29] /*46045*/;
assign _31130_ = _31131_ & D[36] /*46044*/;
assign _31133_ = _30437_ & _31130_ /*46039*/;
assign _31134_ = _30437_ ^ _31130_ /*46042*/;
assign _31135_ = _31126_ & _31134_ /*46040*/;
assign _30885_ = _31126_ ^ _31134_ /*46041*/;
assign _31132_ = _31133_ | _31135_ /*46038*/;
assign _31137_ = ~Q[29] /*46037*/;
assign _31136_ = _31137_ & D[37] /*46036*/;
assign _31139_ = _30438_ & _31136_ /*46031*/;
assign _31140_ = _30438_ ^ _31136_ /*46034*/;
assign _31141_ = _31132_ & _31140_ /*46032*/;
assign _30886_ = _31132_ ^ _31140_ /*46033*/;
assign _31138_ = _31139_ | _31141_ /*46030*/;
assign _31143_ = ~Q[29] /*46029*/;
assign _31142_ = _31143_ & D[38] /*46028*/;
assign _31145_ = _30439_ & _31142_ /*46023*/;
assign _31146_ = _30439_ ^ _31142_ /*46026*/;
assign _31147_ = _31138_ & _31146_ /*46024*/;
assign _30887_ = _31138_ ^ _31146_ /*46025*/;
assign _31144_ = _31145_ | _31147_ /*46022*/;
assign _31149_ = ~Q[29] /*46021*/;
assign _31148_ = _31149_ & D[39] /*46020*/;
assign _31151_ = _30440_ & _31148_ /*46015*/;
assign _31152_ = _30440_ ^ _31148_ /*46018*/;
assign _31153_ = _31144_ & _31152_ /*46016*/;
assign _30888_ = _31144_ ^ _31152_ /*46017*/;
assign _31150_ = _31151_ | _31153_ /*46014*/;
assign _31155_ = ~Q[29] /*46013*/;
assign _31154_ = _31155_ & D[40] /*46012*/;
assign _31157_ = _30441_ & _31154_ /*46007*/;
assign _31158_ = _30441_ ^ _31154_ /*46010*/;
assign _31159_ = _31150_ & _31158_ /*46008*/;
assign _30889_ = _31150_ ^ _31158_ /*46009*/;
assign _31156_ = _31157_ | _31159_ /*46006*/;
assign _31161_ = ~Q[29] /*46005*/;
assign _31160_ = _31161_ & D[41] /*46004*/;
assign _31163_ = _30442_ & _31160_ /*45999*/;
assign _31164_ = _30442_ ^ _31160_ /*46002*/;
assign _31165_ = _31156_ & _31164_ /*46000*/;
assign _30890_ = _31156_ ^ _31164_ /*46001*/;
assign _31162_ = _31163_ | _31165_ /*45998*/;
assign _31167_ = ~Q[29] /*45997*/;
assign _31166_ = _31167_ & D[42] /*45996*/;
assign _31169_ = _30443_ & _31166_ /*45991*/;
assign _31170_ = _30443_ ^ _31166_ /*45994*/;
assign _31171_ = _31162_ & _31170_ /*45992*/;
assign _30891_ = _31162_ ^ _31170_ /*45993*/;
assign _31168_ = _31169_ | _31171_ /*45990*/;
assign _31173_ = ~Q[29] /*45989*/;
assign _31172_ = _31173_ & D[43] /*45988*/;
assign _31175_ = _30444_ & _31172_ /*45983*/;
assign _31176_ = _30444_ ^ _31172_ /*45986*/;
assign _31177_ = _31168_ & _31176_ /*45984*/;
assign _30892_ = _31168_ ^ _31176_ /*45985*/;
assign _31174_ = _31175_ | _31177_ /*45982*/;
assign _31179_ = ~Q[29] /*45981*/;
assign _31178_ = _31179_ & D[44] /*45980*/;
assign _31181_ = _30445_ & _31178_ /*45975*/;
assign _31182_ = _30445_ ^ _31178_ /*45978*/;
assign _31183_ = _31174_ & _31182_ /*45976*/;
assign _30893_ = _31174_ ^ _31182_ /*45977*/;
assign _31180_ = _31181_ | _31183_ /*45974*/;
assign _31185_ = ~Q[29] /*45973*/;
assign _31184_ = _31185_ & D[45] /*45972*/;
assign _31187_ = _30446_ & _31184_ /*45967*/;
assign _31188_ = _30446_ ^ _31184_ /*45970*/;
assign _31189_ = _31180_ & _31188_ /*45968*/;
assign _30894_ = _31180_ ^ _31188_ /*45969*/;
assign _31186_ = _31187_ | _31189_ /*45966*/;
assign _31191_ = ~Q[29] /*45965*/;
assign _31190_ = _31191_ & D[46] /*45964*/;
assign _31193_ = _30447_ & _31190_ /*45959*/;
assign _31194_ = _30447_ ^ _31190_ /*45962*/;
assign _31195_ = _31186_ & _31194_ /*45960*/;
assign _30895_ = _31186_ ^ _31194_ /*45961*/;
assign _31192_ = _31193_ | _31195_ /*45958*/;
assign _31197_ = ~Q[29] /*45957*/;
assign _31196_ = _31197_ & D[47] /*45956*/;
assign _31199_ = _30448_ & _31196_ /*45951*/;
assign _31200_ = _30448_ ^ _31196_ /*45954*/;
assign _31201_ = _31192_ & _31200_ /*45952*/;
assign _30896_ = _31192_ ^ _31200_ /*45953*/;
assign _31198_ = _31199_ | _31201_ /*45950*/;
assign _31203_ = ~Q[29] /*45949*/;
assign _31202_ = _31203_ & D[48] /*45948*/;
assign _31205_ = _30449_ & _31202_ /*45943*/;
assign _31206_ = _30449_ ^ _31202_ /*45946*/;
assign _31207_ = _31198_ & _31206_ /*45944*/;
assign _30897_ = _31198_ ^ _31206_ /*45945*/;
assign _31204_ = _31205_ | _31207_ /*45942*/;
assign _31209_ = ~Q[29] /*45941*/;
assign _31208_ = _31209_ & D[49] /*45940*/;
assign _31211_ = _30450_ & _31208_ /*45935*/;
assign _31212_ = _30450_ ^ _31208_ /*45938*/;
assign _31213_ = _31204_ & _31212_ /*45936*/;
assign _30898_ = _31204_ ^ _31212_ /*45937*/;
assign _31210_ = _31211_ | _31213_ /*45934*/;
assign _31215_ = ~Q[29] /*45933*/;
assign _31214_ = _31215_ & D[50] /*45932*/;
assign _31217_ = _30451_ & _31214_ /*45927*/;
assign _31218_ = _30451_ ^ _31214_ /*45930*/;
assign _31219_ = _31210_ & _31218_ /*45928*/;
assign _30899_ = _31210_ ^ _31218_ /*45929*/;
assign _31216_ = _31217_ | _31219_ /*45926*/;
assign _31221_ = ~Q[29] /*45925*/;
assign _31220_ = _31221_ & D[51] /*45924*/;
assign _31223_ = _30452_ & _31220_ /*45919*/;
assign _31224_ = _30452_ ^ _31220_ /*45922*/;
assign _31225_ = _31216_ & _31224_ /*45920*/;
assign _30900_ = _31216_ ^ _31224_ /*45921*/;
assign _31222_ = _31223_ | _31225_ /*45918*/;
assign _31227_ = ~Q[29] /*45917*/;
assign _31226_ = _31227_ & D[52] /*45916*/;
assign _31229_ = _30453_ & _31226_ /*45911*/;
assign _31230_ = _30453_ ^ _31226_ /*45914*/;
assign _31231_ = _31222_ & _31230_ /*45912*/;
assign _30901_ = _31222_ ^ _31230_ /*45913*/;
assign _31228_ = _31229_ | _31231_ /*45910*/;
assign _31233_ = ~Q[29] /*45909*/;
assign _31232_ = _31233_ & D[53] /*45908*/;
assign _31235_ = _30454_ & _31232_ /*45903*/;
assign _31236_ = _30454_ ^ _31232_ /*45906*/;
assign _31237_ = _31228_ & _31236_ /*45904*/;
assign _30902_ = _31228_ ^ _31236_ /*45905*/;
assign _31234_ = _31235_ | _31237_ /*45902*/;
assign _31239_ = ~Q[29] /*45901*/;
assign _31238_ = _31239_ & D[54] /*45900*/;
assign _31241_ = _30455_ & _31238_ /*45895*/;
assign _31242_ = _30455_ ^ _31238_ /*45898*/;
assign _31243_ = _31234_ & _31242_ /*45896*/;
assign _30903_ = _31234_ ^ _31242_ /*45897*/;
assign _31240_ = _31241_ | _31243_ /*45894*/;
assign _31245_ = ~Q[29] /*45893*/;
assign _31244_ = _31245_ & D[55] /*45892*/;
assign _31247_ = _30456_ & _31244_ /*45887*/;
assign _31248_ = _30456_ ^ _31244_ /*45890*/;
assign _31249_ = _31240_ & _31248_ /*45888*/;
assign _30904_ = _31240_ ^ _31248_ /*45889*/;
assign _31246_ = _31247_ | _31249_ /*45886*/;
assign _31251_ = ~Q[29] /*45885*/;
assign _31250_ = _31251_ & D[56] /*45884*/;
assign _31253_ = _30457_ & _31250_ /*45879*/;
assign _31254_ = _30457_ ^ _31250_ /*45882*/;
assign _31255_ = _31246_ & _31254_ /*45880*/;
assign _30905_ = _31246_ ^ _31254_ /*45881*/;
assign _31252_ = _31253_ | _31255_ /*45878*/;
assign _31257_ = ~Q[29] /*45877*/;
assign _31256_ = _31257_ & D[57] /*45876*/;
assign _31259_ = _30458_ & _31256_ /*45871*/;
assign _31260_ = _30458_ ^ _31256_ /*45874*/;
assign _31261_ = _31252_ & _31260_ /*45872*/;
assign _30906_ = _31252_ ^ _31260_ /*45873*/;
assign _31258_ = _31259_ | _31261_ /*45870*/;
assign _31263_ = ~Q[29] /*45869*/;
assign _31262_ = _31263_ & D[58] /*45868*/;
assign _31265_ = _30459_ & _31262_ /*45863*/;
assign _31266_ = _30459_ ^ _31262_ /*45866*/;
assign _31267_ = _31258_ & _31266_ /*45864*/;
assign _30907_ = _31258_ ^ _31266_ /*45865*/;
assign _31264_ = _31265_ | _31267_ /*45862*/;
assign _31269_ = ~Q[29] /*45861*/;
assign _31268_ = _31269_ & D[59] /*45860*/;
assign _31271_ = _30460_ & _31268_ /*45855*/;
assign _31272_ = _30460_ ^ _31268_ /*45858*/;
assign _31273_ = _31264_ & _31272_ /*45856*/;
assign _30908_ = _31264_ ^ _31272_ /*45857*/;
assign _31270_ = _31271_ | _31273_ /*45854*/;
assign _31275_ = ~Q[29] /*45853*/;
assign _31274_ = _31275_ & D[60] /*45852*/;
assign _31277_ = _30461_ & _31274_ /*45847*/;
assign _31278_ = _30461_ ^ _31274_ /*45850*/;
assign _31279_ = _31270_ & _31278_ /*45848*/;
assign _30909_ = _31270_ ^ _31278_ /*45849*/;
assign _31276_ = _31277_ | _31279_ /*45846*/;
assign _31281_ = ~Q[29] /*45845*/;
assign _31280_ = _31281_ & D[61] /*45844*/;
assign _31283_ = _30462_ & _31280_ /*45839*/;
assign _31284_ = _30462_ ^ _31280_ /*45842*/;
assign _31285_ = _31276_ & _31284_ /*45840*/;
assign _30910_ = _31276_ ^ _31284_ /*45841*/;
assign _31282_ = _31283_ | _31285_ /*45838*/;
assign _31287_ = ~Q[29] /*45837*/;
assign _31286_ = _31287_ & D[62] /*45836*/;
assign _31289_ = _30463_ & _31286_ /*45831*/;
assign _31290_ = _30463_ ^ _31286_ /*45834*/;
assign _31291_ = _31282_ & _31290_ /*45832*/;
assign _30911_ = _31282_ ^ _31290_ /*45833*/;
assign _31288_ = _31289_ | _31291_ /*45830*/;
assign _31293_ = ~Q[29] /*45829*/;
assign _31292_ = _31293_ & zeroWire /*45828*/;
assign _31294_ = _30464_ ^ _31292_ /*45826*/;
assign _30912_ = _31294_ ^ _31288_ /*45825*/;
assign _31365_ = ~D[0] /*45571*/;
assign _31362_ = R_0[28] & _31365_ /*45567*/;
assign _31363_ = R_0[28] ^ _31365_ /*45570*/;
assign _31364_ = oneWire & _31363_ /*45568*/;
assign _31297_ = oneWire ^ _31363_ /*45569*/;
assign _31361_ = _31362_ | _31364_ /*45566*/;
assign _31370_ = ~D[1] /*45565*/;
assign _31367_ = _30849_ & _31370_ /*45561*/;
assign _31368_ = _30849_ ^ _31370_ /*45564*/;
assign _31369_ = _31361_ & _31368_ /*45562*/;
assign _31298_ = _31361_ ^ _31368_ /*45563*/;
assign _31366_ = _31367_ | _31369_ /*45560*/;
assign _31375_ = ~D[2] /*45559*/;
assign _31372_ = _30850_ & _31375_ /*45555*/;
assign _31373_ = _30850_ ^ _31375_ /*45558*/;
assign _31374_ = _31366_ & _31373_ /*45556*/;
assign _31299_ = _31366_ ^ _31373_ /*45557*/;
assign _31371_ = _31372_ | _31374_ /*45554*/;
assign _31380_ = ~D[3] /*45553*/;
assign _31377_ = _30851_ & _31380_ /*45549*/;
assign _31378_ = _30851_ ^ _31380_ /*45552*/;
assign _31379_ = _31371_ & _31378_ /*45550*/;
assign _31300_ = _31371_ ^ _31378_ /*45551*/;
assign _31376_ = _31377_ | _31379_ /*45548*/;
assign _31385_ = ~D[4] /*45547*/;
assign _31382_ = _30852_ & _31385_ /*45543*/;
assign _31383_ = _30852_ ^ _31385_ /*45546*/;
assign _31384_ = _31376_ & _31383_ /*45544*/;
assign _31301_ = _31376_ ^ _31383_ /*45545*/;
assign _31381_ = _31382_ | _31384_ /*45542*/;
assign _31390_ = ~D[5] /*45541*/;
assign _31387_ = _30853_ & _31390_ /*45537*/;
assign _31388_ = _30853_ ^ _31390_ /*45540*/;
assign _31389_ = _31381_ & _31388_ /*45538*/;
assign _31302_ = _31381_ ^ _31388_ /*45539*/;
assign _31386_ = _31387_ | _31389_ /*45536*/;
assign _31395_ = ~D[6] /*45535*/;
assign _31392_ = _30854_ & _31395_ /*45531*/;
assign _31393_ = _30854_ ^ _31395_ /*45534*/;
assign _31394_ = _31386_ & _31393_ /*45532*/;
assign _31303_ = _31386_ ^ _31393_ /*45533*/;
assign _31391_ = _31392_ | _31394_ /*45530*/;
assign _31400_ = ~D[7] /*45529*/;
assign _31397_ = _30855_ & _31400_ /*45525*/;
assign _31398_ = _30855_ ^ _31400_ /*45528*/;
assign _31399_ = _31391_ & _31398_ /*45526*/;
assign _31304_ = _31391_ ^ _31398_ /*45527*/;
assign _31396_ = _31397_ | _31399_ /*45524*/;
assign _31405_ = ~D[8] /*45523*/;
assign _31402_ = _30856_ & _31405_ /*45519*/;
assign _31403_ = _30856_ ^ _31405_ /*45522*/;
assign _31404_ = _31396_ & _31403_ /*45520*/;
assign _31305_ = _31396_ ^ _31403_ /*45521*/;
assign _31401_ = _31402_ | _31404_ /*45518*/;
assign _31410_ = ~D[9] /*45517*/;
assign _31407_ = _30857_ & _31410_ /*45513*/;
assign _31408_ = _30857_ ^ _31410_ /*45516*/;
assign _31409_ = _31401_ & _31408_ /*45514*/;
assign _31306_ = _31401_ ^ _31408_ /*45515*/;
assign _31406_ = _31407_ | _31409_ /*45512*/;
assign _31415_ = ~D[10] /*45511*/;
assign _31412_ = _30858_ & _31415_ /*45507*/;
assign _31413_ = _30858_ ^ _31415_ /*45510*/;
assign _31414_ = _31406_ & _31413_ /*45508*/;
assign _31307_ = _31406_ ^ _31413_ /*45509*/;
assign _31411_ = _31412_ | _31414_ /*45506*/;
assign _31420_ = ~D[11] /*45505*/;
assign _31417_ = _30859_ & _31420_ /*45501*/;
assign _31418_ = _30859_ ^ _31420_ /*45504*/;
assign _31419_ = _31411_ & _31418_ /*45502*/;
assign _31308_ = _31411_ ^ _31418_ /*45503*/;
assign _31416_ = _31417_ | _31419_ /*45500*/;
assign _31425_ = ~D[12] /*45499*/;
assign _31422_ = _30860_ & _31425_ /*45495*/;
assign _31423_ = _30860_ ^ _31425_ /*45498*/;
assign _31424_ = _31416_ & _31423_ /*45496*/;
assign _31309_ = _31416_ ^ _31423_ /*45497*/;
assign _31421_ = _31422_ | _31424_ /*45494*/;
assign _31430_ = ~D[13] /*45493*/;
assign _31427_ = _30861_ & _31430_ /*45489*/;
assign _31428_ = _30861_ ^ _31430_ /*45492*/;
assign _31429_ = _31421_ & _31428_ /*45490*/;
assign _31310_ = _31421_ ^ _31428_ /*45491*/;
assign _31426_ = _31427_ | _31429_ /*45488*/;
assign _31435_ = ~D[14] /*45487*/;
assign _31432_ = _30862_ & _31435_ /*45483*/;
assign _31433_ = _30862_ ^ _31435_ /*45486*/;
assign _31434_ = _31426_ & _31433_ /*45484*/;
assign _31311_ = _31426_ ^ _31433_ /*45485*/;
assign _31431_ = _31432_ | _31434_ /*45482*/;
assign _31440_ = ~D[15] /*45481*/;
assign _31437_ = _30863_ & _31440_ /*45477*/;
assign _31438_ = _30863_ ^ _31440_ /*45480*/;
assign _31439_ = _31431_ & _31438_ /*45478*/;
assign _31312_ = _31431_ ^ _31438_ /*45479*/;
assign _31436_ = _31437_ | _31439_ /*45476*/;
assign _31445_ = ~D[16] /*45475*/;
assign _31442_ = _30864_ & _31445_ /*45471*/;
assign _31443_ = _30864_ ^ _31445_ /*45474*/;
assign _31444_ = _31436_ & _31443_ /*45472*/;
assign _31313_ = _31436_ ^ _31443_ /*45473*/;
assign _31441_ = _31442_ | _31444_ /*45470*/;
assign _31450_ = ~D[17] /*45469*/;
assign _31447_ = _30865_ & _31450_ /*45465*/;
assign _31448_ = _30865_ ^ _31450_ /*45468*/;
assign _31449_ = _31441_ & _31448_ /*45466*/;
assign _31314_ = _31441_ ^ _31448_ /*45467*/;
assign _31446_ = _31447_ | _31449_ /*45464*/;
assign _31455_ = ~D[18] /*45463*/;
assign _31452_ = _30866_ & _31455_ /*45459*/;
assign _31453_ = _30866_ ^ _31455_ /*45462*/;
assign _31454_ = _31446_ & _31453_ /*45460*/;
assign _31315_ = _31446_ ^ _31453_ /*45461*/;
assign _31451_ = _31452_ | _31454_ /*45458*/;
assign _31460_ = ~D[19] /*45457*/;
assign _31457_ = _30867_ & _31460_ /*45453*/;
assign _31458_ = _30867_ ^ _31460_ /*45456*/;
assign _31459_ = _31451_ & _31458_ /*45454*/;
assign _31316_ = _31451_ ^ _31458_ /*45455*/;
assign _31456_ = _31457_ | _31459_ /*45452*/;
assign _31465_ = ~D[20] /*45451*/;
assign _31462_ = _30868_ & _31465_ /*45447*/;
assign _31463_ = _30868_ ^ _31465_ /*45450*/;
assign _31464_ = _31456_ & _31463_ /*45448*/;
assign _31317_ = _31456_ ^ _31463_ /*45449*/;
assign _31461_ = _31462_ | _31464_ /*45446*/;
assign _31470_ = ~D[21] /*45445*/;
assign _31467_ = _30869_ & _31470_ /*45441*/;
assign _31468_ = _30869_ ^ _31470_ /*45444*/;
assign _31469_ = _31461_ & _31468_ /*45442*/;
assign _31318_ = _31461_ ^ _31468_ /*45443*/;
assign _31466_ = _31467_ | _31469_ /*45440*/;
assign _31475_ = ~D[22] /*45439*/;
assign _31472_ = _30870_ & _31475_ /*45435*/;
assign _31473_ = _30870_ ^ _31475_ /*45438*/;
assign _31474_ = _31466_ & _31473_ /*45436*/;
assign _31319_ = _31466_ ^ _31473_ /*45437*/;
assign _31471_ = _31472_ | _31474_ /*45434*/;
assign _31480_ = ~D[23] /*45433*/;
assign _31477_ = _30871_ & _31480_ /*45429*/;
assign _31478_ = _30871_ ^ _31480_ /*45432*/;
assign _31479_ = _31471_ & _31478_ /*45430*/;
assign _31320_ = _31471_ ^ _31478_ /*45431*/;
assign _31476_ = _31477_ | _31479_ /*45428*/;
assign _31485_ = ~D[24] /*45427*/;
assign _31482_ = _30872_ & _31485_ /*45423*/;
assign _31483_ = _30872_ ^ _31485_ /*45426*/;
assign _31484_ = _31476_ & _31483_ /*45424*/;
assign _31321_ = _31476_ ^ _31483_ /*45425*/;
assign _31481_ = _31482_ | _31484_ /*45422*/;
assign _31490_ = ~D[25] /*45421*/;
assign _31487_ = _30873_ & _31490_ /*45417*/;
assign _31488_ = _30873_ ^ _31490_ /*45420*/;
assign _31489_ = _31481_ & _31488_ /*45418*/;
assign _31322_ = _31481_ ^ _31488_ /*45419*/;
assign _31486_ = _31487_ | _31489_ /*45416*/;
assign _31495_ = ~D[26] /*45415*/;
assign _31492_ = _30874_ & _31495_ /*45411*/;
assign _31493_ = _30874_ ^ _31495_ /*45414*/;
assign _31494_ = _31486_ & _31493_ /*45412*/;
assign _31323_ = _31486_ ^ _31493_ /*45413*/;
assign _31491_ = _31492_ | _31494_ /*45410*/;
assign _31500_ = ~D[27] /*45409*/;
assign _31497_ = _30875_ & _31500_ /*45405*/;
assign _31498_ = _30875_ ^ _31500_ /*45408*/;
assign _31499_ = _31491_ & _31498_ /*45406*/;
assign _31324_ = _31491_ ^ _31498_ /*45407*/;
assign _31496_ = _31497_ | _31499_ /*45404*/;
assign _31505_ = ~D[28] /*45403*/;
assign _31502_ = _30876_ & _31505_ /*45399*/;
assign _31503_ = _30876_ ^ _31505_ /*45402*/;
assign _31504_ = _31496_ & _31503_ /*45400*/;
assign _31325_ = _31496_ ^ _31503_ /*45401*/;
assign _31501_ = _31502_ | _31504_ /*45398*/;
assign _31510_ = ~D[29] /*45397*/;
assign _31507_ = _30877_ & _31510_ /*45393*/;
assign _31508_ = _30877_ ^ _31510_ /*45396*/;
assign _31509_ = _31501_ & _31508_ /*45394*/;
assign _31326_ = _31501_ ^ _31508_ /*45395*/;
assign _31506_ = _31507_ | _31509_ /*45392*/;
assign _31515_ = ~D[30] /*45391*/;
assign _31512_ = _30878_ & _31515_ /*45387*/;
assign _31513_ = _30878_ ^ _31515_ /*45390*/;
assign _31514_ = _31506_ & _31513_ /*45388*/;
assign _31327_ = _31506_ ^ _31513_ /*45389*/;
assign _31511_ = _31512_ | _31514_ /*45386*/;
assign _31520_ = ~D[31] /*45385*/;
assign _31517_ = _30879_ & _31520_ /*45381*/;
assign _31518_ = _30879_ ^ _31520_ /*45384*/;
assign _31519_ = _31511_ & _31518_ /*45382*/;
assign _31328_ = _31511_ ^ _31518_ /*45383*/;
assign _31516_ = _31517_ | _31519_ /*45380*/;
assign _31525_ = ~D[32] /*45379*/;
assign _31522_ = _30880_ & _31525_ /*45375*/;
assign _31523_ = _30880_ ^ _31525_ /*45378*/;
assign _31524_ = _31516_ & _31523_ /*45376*/;
assign _31329_ = _31516_ ^ _31523_ /*45377*/;
assign _31521_ = _31522_ | _31524_ /*45374*/;
assign _31530_ = ~D[33] /*45373*/;
assign _31527_ = _30881_ & _31530_ /*45369*/;
assign _31528_ = _30881_ ^ _31530_ /*45372*/;
assign _31529_ = _31521_ & _31528_ /*45370*/;
assign _31330_ = _31521_ ^ _31528_ /*45371*/;
assign _31526_ = _31527_ | _31529_ /*45368*/;
assign _31535_ = ~D[34] /*45367*/;
assign _31532_ = _30882_ & _31535_ /*45363*/;
assign _31533_ = _30882_ ^ _31535_ /*45366*/;
assign _31534_ = _31526_ & _31533_ /*45364*/;
assign _31331_ = _31526_ ^ _31533_ /*45365*/;
assign _31531_ = _31532_ | _31534_ /*45362*/;
assign _31540_ = ~D[35] /*45361*/;
assign _31537_ = _30883_ & _31540_ /*45357*/;
assign _31538_ = _30883_ ^ _31540_ /*45360*/;
assign _31539_ = _31531_ & _31538_ /*45358*/;
assign _31332_ = _31531_ ^ _31538_ /*45359*/;
assign _31536_ = _31537_ | _31539_ /*45356*/;
assign _31545_ = ~D[36] /*45355*/;
assign _31542_ = _30884_ & _31545_ /*45351*/;
assign _31543_ = _30884_ ^ _31545_ /*45354*/;
assign _31544_ = _31536_ & _31543_ /*45352*/;
assign _31333_ = _31536_ ^ _31543_ /*45353*/;
assign _31541_ = _31542_ | _31544_ /*45350*/;
assign _31550_ = ~D[37] /*45349*/;
assign _31547_ = _30885_ & _31550_ /*45345*/;
assign _31548_ = _30885_ ^ _31550_ /*45348*/;
assign _31549_ = _31541_ & _31548_ /*45346*/;
assign _31334_ = _31541_ ^ _31548_ /*45347*/;
assign _31546_ = _31547_ | _31549_ /*45344*/;
assign _31555_ = ~D[38] /*45343*/;
assign _31552_ = _30886_ & _31555_ /*45339*/;
assign _31553_ = _30886_ ^ _31555_ /*45342*/;
assign _31554_ = _31546_ & _31553_ /*45340*/;
assign _31335_ = _31546_ ^ _31553_ /*45341*/;
assign _31551_ = _31552_ | _31554_ /*45338*/;
assign _31560_ = ~D[39] /*45337*/;
assign _31557_ = _30887_ & _31560_ /*45333*/;
assign _31558_ = _30887_ ^ _31560_ /*45336*/;
assign _31559_ = _31551_ & _31558_ /*45334*/;
assign _31336_ = _31551_ ^ _31558_ /*45335*/;
assign _31556_ = _31557_ | _31559_ /*45332*/;
assign _31565_ = ~D[40] /*45331*/;
assign _31562_ = _30888_ & _31565_ /*45327*/;
assign _31563_ = _30888_ ^ _31565_ /*45330*/;
assign _31564_ = _31556_ & _31563_ /*45328*/;
assign _31337_ = _31556_ ^ _31563_ /*45329*/;
assign _31561_ = _31562_ | _31564_ /*45326*/;
assign _31570_ = ~D[41] /*45325*/;
assign _31567_ = _30889_ & _31570_ /*45321*/;
assign _31568_ = _30889_ ^ _31570_ /*45324*/;
assign _31569_ = _31561_ & _31568_ /*45322*/;
assign _31338_ = _31561_ ^ _31568_ /*45323*/;
assign _31566_ = _31567_ | _31569_ /*45320*/;
assign _31575_ = ~D[42] /*45319*/;
assign _31572_ = _30890_ & _31575_ /*45315*/;
assign _31573_ = _30890_ ^ _31575_ /*45318*/;
assign _31574_ = _31566_ & _31573_ /*45316*/;
assign _31339_ = _31566_ ^ _31573_ /*45317*/;
assign _31571_ = _31572_ | _31574_ /*45314*/;
assign _31580_ = ~D[43] /*45313*/;
assign _31577_ = _30891_ & _31580_ /*45309*/;
assign _31578_ = _30891_ ^ _31580_ /*45312*/;
assign _31579_ = _31571_ & _31578_ /*45310*/;
assign _31340_ = _31571_ ^ _31578_ /*45311*/;
assign _31576_ = _31577_ | _31579_ /*45308*/;
assign _31585_ = ~D[44] /*45307*/;
assign _31582_ = _30892_ & _31585_ /*45303*/;
assign _31583_ = _30892_ ^ _31585_ /*45306*/;
assign _31584_ = _31576_ & _31583_ /*45304*/;
assign _31341_ = _31576_ ^ _31583_ /*45305*/;
assign _31581_ = _31582_ | _31584_ /*45302*/;
assign _31590_ = ~D[45] /*45301*/;
assign _31587_ = _30893_ & _31590_ /*45297*/;
assign _31588_ = _30893_ ^ _31590_ /*45300*/;
assign _31589_ = _31581_ & _31588_ /*45298*/;
assign _31342_ = _31581_ ^ _31588_ /*45299*/;
assign _31586_ = _31587_ | _31589_ /*45296*/;
assign _31595_ = ~D[46] /*45295*/;
assign _31592_ = _30894_ & _31595_ /*45291*/;
assign _31593_ = _30894_ ^ _31595_ /*45294*/;
assign _31594_ = _31586_ & _31593_ /*45292*/;
assign _31343_ = _31586_ ^ _31593_ /*45293*/;
assign _31591_ = _31592_ | _31594_ /*45290*/;
assign _31600_ = ~D[47] /*45289*/;
assign _31597_ = _30895_ & _31600_ /*45285*/;
assign _31598_ = _30895_ ^ _31600_ /*45288*/;
assign _31599_ = _31591_ & _31598_ /*45286*/;
assign _31344_ = _31591_ ^ _31598_ /*45287*/;
assign _31596_ = _31597_ | _31599_ /*45284*/;
assign _31605_ = ~D[48] /*45283*/;
assign _31602_ = _30896_ & _31605_ /*45279*/;
assign _31603_ = _30896_ ^ _31605_ /*45282*/;
assign _31604_ = _31596_ & _31603_ /*45280*/;
assign _31345_ = _31596_ ^ _31603_ /*45281*/;
assign _31601_ = _31602_ | _31604_ /*45278*/;
assign _31610_ = ~D[49] /*45277*/;
assign _31607_ = _30897_ & _31610_ /*45273*/;
assign _31608_ = _30897_ ^ _31610_ /*45276*/;
assign _31609_ = _31601_ & _31608_ /*45274*/;
assign _31346_ = _31601_ ^ _31608_ /*45275*/;
assign _31606_ = _31607_ | _31609_ /*45272*/;
assign _31615_ = ~D[50] /*45271*/;
assign _31612_ = _30898_ & _31615_ /*45267*/;
assign _31613_ = _30898_ ^ _31615_ /*45270*/;
assign _31614_ = _31606_ & _31613_ /*45268*/;
assign _31347_ = _31606_ ^ _31613_ /*45269*/;
assign _31611_ = _31612_ | _31614_ /*45266*/;
assign _31620_ = ~D[51] /*45265*/;
assign _31617_ = _30899_ & _31620_ /*45261*/;
assign _31618_ = _30899_ ^ _31620_ /*45264*/;
assign _31619_ = _31611_ & _31618_ /*45262*/;
assign _31348_ = _31611_ ^ _31618_ /*45263*/;
assign _31616_ = _31617_ | _31619_ /*45260*/;
assign _31625_ = ~D[52] /*45259*/;
assign _31622_ = _30900_ & _31625_ /*45255*/;
assign _31623_ = _30900_ ^ _31625_ /*45258*/;
assign _31624_ = _31616_ & _31623_ /*45256*/;
assign _31349_ = _31616_ ^ _31623_ /*45257*/;
assign _31621_ = _31622_ | _31624_ /*45254*/;
assign _31630_ = ~D[53] /*45253*/;
assign _31627_ = _30901_ & _31630_ /*45249*/;
assign _31628_ = _30901_ ^ _31630_ /*45252*/;
assign _31629_ = _31621_ & _31628_ /*45250*/;
assign _31350_ = _31621_ ^ _31628_ /*45251*/;
assign _31626_ = _31627_ | _31629_ /*45248*/;
assign _31635_ = ~D[54] /*45247*/;
assign _31632_ = _30902_ & _31635_ /*45243*/;
assign _31633_ = _30902_ ^ _31635_ /*45246*/;
assign _31634_ = _31626_ & _31633_ /*45244*/;
assign _31351_ = _31626_ ^ _31633_ /*45245*/;
assign _31631_ = _31632_ | _31634_ /*45242*/;
assign _31640_ = ~D[55] /*45241*/;
assign _31637_ = _30903_ & _31640_ /*45237*/;
assign _31638_ = _30903_ ^ _31640_ /*45240*/;
assign _31639_ = _31631_ & _31638_ /*45238*/;
assign _31352_ = _31631_ ^ _31638_ /*45239*/;
assign _31636_ = _31637_ | _31639_ /*45236*/;
assign _31645_ = ~D[56] /*45235*/;
assign _31642_ = _30904_ & _31645_ /*45231*/;
assign _31643_ = _30904_ ^ _31645_ /*45234*/;
assign _31644_ = _31636_ & _31643_ /*45232*/;
assign _31353_ = _31636_ ^ _31643_ /*45233*/;
assign _31641_ = _31642_ | _31644_ /*45230*/;
assign _31650_ = ~D[57] /*45229*/;
assign _31647_ = _30905_ & _31650_ /*45225*/;
assign _31648_ = _30905_ ^ _31650_ /*45228*/;
assign _31649_ = _31641_ & _31648_ /*45226*/;
assign _31354_ = _31641_ ^ _31648_ /*45227*/;
assign _31646_ = _31647_ | _31649_ /*45224*/;
assign _31655_ = ~D[58] /*45223*/;
assign _31652_ = _30906_ & _31655_ /*45219*/;
assign _31653_ = _30906_ ^ _31655_ /*45222*/;
assign _31654_ = _31646_ & _31653_ /*45220*/;
assign _31355_ = _31646_ ^ _31653_ /*45221*/;
assign _31651_ = _31652_ | _31654_ /*45218*/;
assign _31660_ = ~D[59] /*45217*/;
assign _31657_ = _30907_ & _31660_ /*45213*/;
assign _31658_ = _30907_ ^ _31660_ /*45216*/;
assign _31659_ = _31651_ & _31658_ /*45214*/;
assign _31356_ = _31651_ ^ _31658_ /*45215*/;
assign _31656_ = _31657_ | _31659_ /*45212*/;
assign _31665_ = ~D[60] /*45211*/;
assign _31662_ = _30908_ & _31665_ /*45207*/;
assign _31663_ = _30908_ ^ _31665_ /*45210*/;
assign _31664_ = _31656_ & _31663_ /*45208*/;
assign _31357_ = _31656_ ^ _31663_ /*45209*/;
assign _31661_ = _31662_ | _31664_ /*45206*/;
assign _31670_ = ~D[61] /*45205*/;
assign _31667_ = _30909_ & _31670_ /*45201*/;
assign _31668_ = _30909_ ^ _31670_ /*45204*/;
assign _31669_ = _31661_ & _31668_ /*45202*/;
assign _31358_ = _31661_ ^ _31668_ /*45203*/;
assign _31666_ = _31667_ | _31669_ /*45200*/;
assign _31675_ = ~D[62] /*45199*/;
assign _31672_ = _30910_ & _31675_ /*45195*/;
assign _31673_ = _30910_ ^ _31675_ /*45198*/;
assign _31674_ = _31666_ & _31673_ /*45196*/;
assign _31359_ = _31666_ ^ _31673_ /*45197*/;
assign _31671_ = _31672_ | _31674_ /*45194*/;
assign _31676_ = _30911_ & oneWire /*45189*/;
assign _31677_ = _30911_ ^ oneWire /*45192*/;
assign _31678_ = _31671_ & _31677_ /*45190*/;
assign _31360_ = _31671_ ^ _31677_ /*45191*/;
assign Q[28] = _31676_ | _31678_ /*45188*/;
assign _31811_ = ~Q[28] /*44803*/;
assign _31810_ = _31811_ & D[0] /*44802*/;
assign _31813_ = _31297_ & _31810_ /*44797*/;
assign _31814_ = _31297_ ^ _31810_ /*44800*/;
assign _31815_ = zeroWire & _31814_ /*44798*/;
assign _31745_ = zeroWire ^ _31814_ /*44799*/;
assign _31812_ = _31813_ | _31815_ /*44796*/;
assign _31817_ = ~Q[28] /*44795*/;
assign _31816_ = _31817_ & D[1] /*44794*/;
assign _31819_ = _31298_ & _31816_ /*44789*/;
assign _31820_ = _31298_ ^ _31816_ /*44792*/;
assign _31821_ = _31812_ & _31820_ /*44790*/;
assign _31746_ = _31812_ ^ _31820_ /*44791*/;
assign _31818_ = _31819_ | _31821_ /*44788*/;
assign _31823_ = ~Q[28] /*44787*/;
assign _31822_ = _31823_ & D[2] /*44786*/;
assign _31825_ = _31299_ & _31822_ /*44781*/;
assign _31826_ = _31299_ ^ _31822_ /*44784*/;
assign _31827_ = _31818_ & _31826_ /*44782*/;
assign _31747_ = _31818_ ^ _31826_ /*44783*/;
assign _31824_ = _31825_ | _31827_ /*44780*/;
assign _31829_ = ~Q[28] /*44779*/;
assign _31828_ = _31829_ & D[3] /*44778*/;
assign _31831_ = _31300_ & _31828_ /*44773*/;
assign _31832_ = _31300_ ^ _31828_ /*44776*/;
assign _31833_ = _31824_ & _31832_ /*44774*/;
assign _31748_ = _31824_ ^ _31832_ /*44775*/;
assign _31830_ = _31831_ | _31833_ /*44772*/;
assign _31835_ = ~Q[28] /*44771*/;
assign _31834_ = _31835_ & D[4] /*44770*/;
assign _31837_ = _31301_ & _31834_ /*44765*/;
assign _31838_ = _31301_ ^ _31834_ /*44768*/;
assign _31839_ = _31830_ & _31838_ /*44766*/;
assign _31749_ = _31830_ ^ _31838_ /*44767*/;
assign _31836_ = _31837_ | _31839_ /*44764*/;
assign _31841_ = ~Q[28] /*44763*/;
assign _31840_ = _31841_ & D[5] /*44762*/;
assign _31843_ = _31302_ & _31840_ /*44757*/;
assign _31844_ = _31302_ ^ _31840_ /*44760*/;
assign _31845_ = _31836_ & _31844_ /*44758*/;
assign _31750_ = _31836_ ^ _31844_ /*44759*/;
assign _31842_ = _31843_ | _31845_ /*44756*/;
assign _31847_ = ~Q[28] /*44755*/;
assign _31846_ = _31847_ & D[6] /*44754*/;
assign _31849_ = _31303_ & _31846_ /*44749*/;
assign _31850_ = _31303_ ^ _31846_ /*44752*/;
assign _31851_ = _31842_ & _31850_ /*44750*/;
assign _31751_ = _31842_ ^ _31850_ /*44751*/;
assign _31848_ = _31849_ | _31851_ /*44748*/;
assign _31853_ = ~Q[28] /*44747*/;
assign _31852_ = _31853_ & D[7] /*44746*/;
assign _31855_ = _31304_ & _31852_ /*44741*/;
assign _31856_ = _31304_ ^ _31852_ /*44744*/;
assign _31857_ = _31848_ & _31856_ /*44742*/;
assign _31752_ = _31848_ ^ _31856_ /*44743*/;
assign _31854_ = _31855_ | _31857_ /*44740*/;
assign _31859_ = ~Q[28] /*44739*/;
assign _31858_ = _31859_ & D[8] /*44738*/;
assign _31861_ = _31305_ & _31858_ /*44733*/;
assign _31862_ = _31305_ ^ _31858_ /*44736*/;
assign _31863_ = _31854_ & _31862_ /*44734*/;
assign _31753_ = _31854_ ^ _31862_ /*44735*/;
assign _31860_ = _31861_ | _31863_ /*44732*/;
assign _31865_ = ~Q[28] /*44731*/;
assign _31864_ = _31865_ & D[9] /*44730*/;
assign _31867_ = _31306_ & _31864_ /*44725*/;
assign _31868_ = _31306_ ^ _31864_ /*44728*/;
assign _31869_ = _31860_ & _31868_ /*44726*/;
assign _31754_ = _31860_ ^ _31868_ /*44727*/;
assign _31866_ = _31867_ | _31869_ /*44724*/;
assign _31871_ = ~Q[28] /*44723*/;
assign _31870_ = _31871_ & D[10] /*44722*/;
assign _31873_ = _31307_ & _31870_ /*44717*/;
assign _31874_ = _31307_ ^ _31870_ /*44720*/;
assign _31875_ = _31866_ & _31874_ /*44718*/;
assign _31755_ = _31866_ ^ _31874_ /*44719*/;
assign _31872_ = _31873_ | _31875_ /*44716*/;
assign _31877_ = ~Q[28] /*44715*/;
assign _31876_ = _31877_ & D[11] /*44714*/;
assign _31879_ = _31308_ & _31876_ /*44709*/;
assign _31880_ = _31308_ ^ _31876_ /*44712*/;
assign _31881_ = _31872_ & _31880_ /*44710*/;
assign _31756_ = _31872_ ^ _31880_ /*44711*/;
assign _31878_ = _31879_ | _31881_ /*44708*/;
assign _31883_ = ~Q[28] /*44707*/;
assign _31882_ = _31883_ & D[12] /*44706*/;
assign _31885_ = _31309_ & _31882_ /*44701*/;
assign _31886_ = _31309_ ^ _31882_ /*44704*/;
assign _31887_ = _31878_ & _31886_ /*44702*/;
assign _31757_ = _31878_ ^ _31886_ /*44703*/;
assign _31884_ = _31885_ | _31887_ /*44700*/;
assign _31889_ = ~Q[28] /*44699*/;
assign _31888_ = _31889_ & D[13] /*44698*/;
assign _31891_ = _31310_ & _31888_ /*44693*/;
assign _31892_ = _31310_ ^ _31888_ /*44696*/;
assign _31893_ = _31884_ & _31892_ /*44694*/;
assign _31758_ = _31884_ ^ _31892_ /*44695*/;
assign _31890_ = _31891_ | _31893_ /*44692*/;
assign _31895_ = ~Q[28] /*44691*/;
assign _31894_ = _31895_ & D[14] /*44690*/;
assign _31897_ = _31311_ & _31894_ /*44685*/;
assign _31898_ = _31311_ ^ _31894_ /*44688*/;
assign _31899_ = _31890_ & _31898_ /*44686*/;
assign _31759_ = _31890_ ^ _31898_ /*44687*/;
assign _31896_ = _31897_ | _31899_ /*44684*/;
assign _31901_ = ~Q[28] /*44683*/;
assign _31900_ = _31901_ & D[15] /*44682*/;
assign _31903_ = _31312_ & _31900_ /*44677*/;
assign _31904_ = _31312_ ^ _31900_ /*44680*/;
assign _31905_ = _31896_ & _31904_ /*44678*/;
assign _31760_ = _31896_ ^ _31904_ /*44679*/;
assign _31902_ = _31903_ | _31905_ /*44676*/;
assign _31907_ = ~Q[28] /*44675*/;
assign _31906_ = _31907_ & D[16] /*44674*/;
assign _31909_ = _31313_ & _31906_ /*44669*/;
assign _31910_ = _31313_ ^ _31906_ /*44672*/;
assign _31911_ = _31902_ & _31910_ /*44670*/;
assign _31761_ = _31902_ ^ _31910_ /*44671*/;
assign _31908_ = _31909_ | _31911_ /*44668*/;
assign _31913_ = ~Q[28] /*44667*/;
assign _31912_ = _31913_ & D[17] /*44666*/;
assign _31915_ = _31314_ & _31912_ /*44661*/;
assign _31916_ = _31314_ ^ _31912_ /*44664*/;
assign _31917_ = _31908_ & _31916_ /*44662*/;
assign _31762_ = _31908_ ^ _31916_ /*44663*/;
assign _31914_ = _31915_ | _31917_ /*44660*/;
assign _31919_ = ~Q[28] /*44659*/;
assign _31918_ = _31919_ & D[18] /*44658*/;
assign _31921_ = _31315_ & _31918_ /*44653*/;
assign _31922_ = _31315_ ^ _31918_ /*44656*/;
assign _31923_ = _31914_ & _31922_ /*44654*/;
assign _31763_ = _31914_ ^ _31922_ /*44655*/;
assign _31920_ = _31921_ | _31923_ /*44652*/;
assign _31925_ = ~Q[28] /*44651*/;
assign _31924_ = _31925_ & D[19] /*44650*/;
assign _31927_ = _31316_ & _31924_ /*44645*/;
assign _31928_ = _31316_ ^ _31924_ /*44648*/;
assign _31929_ = _31920_ & _31928_ /*44646*/;
assign _31764_ = _31920_ ^ _31928_ /*44647*/;
assign _31926_ = _31927_ | _31929_ /*44644*/;
assign _31931_ = ~Q[28] /*44643*/;
assign _31930_ = _31931_ & D[20] /*44642*/;
assign _31933_ = _31317_ & _31930_ /*44637*/;
assign _31934_ = _31317_ ^ _31930_ /*44640*/;
assign _31935_ = _31926_ & _31934_ /*44638*/;
assign _31765_ = _31926_ ^ _31934_ /*44639*/;
assign _31932_ = _31933_ | _31935_ /*44636*/;
assign _31937_ = ~Q[28] /*44635*/;
assign _31936_ = _31937_ & D[21] /*44634*/;
assign _31939_ = _31318_ & _31936_ /*44629*/;
assign _31940_ = _31318_ ^ _31936_ /*44632*/;
assign _31941_ = _31932_ & _31940_ /*44630*/;
assign _31766_ = _31932_ ^ _31940_ /*44631*/;
assign _31938_ = _31939_ | _31941_ /*44628*/;
assign _31943_ = ~Q[28] /*44627*/;
assign _31942_ = _31943_ & D[22] /*44626*/;
assign _31945_ = _31319_ & _31942_ /*44621*/;
assign _31946_ = _31319_ ^ _31942_ /*44624*/;
assign _31947_ = _31938_ & _31946_ /*44622*/;
assign _31767_ = _31938_ ^ _31946_ /*44623*/;
assign _31944_ = _31945_ | _31947_ /*44620*/;
assign _31949_ = ~Q[28] /*44619*/;
assign _31948_ = _31949_ & D[23] /*44618*/;
assign _31951_ = _31320_ & _31948_ /*44613*/;
assign _31952_ = _31320_ ^ _31948_ /*44616*/;
assign _31953_ = _31944_ & _31952_ /*44614*/;
assign _31768_ = _31944_ ^ _31952_ /*44615*/;
assign _31950_ = _31951_ | _31953_ /*44612*/;
assign _31955_ = ~Q[28] /*44611*/;
assign _31954_ = _31955_ & D[24] /*44610*/;
assign _31957_ = _31321_ & _31954_ /*44605*/;
assign _31958_ = _31321_ ^ _31954_ /*44608*/;
assign _31959_ = _31950_ & _31958_ /*44606*/;
assign _31769_ = _31950_ ^ _31958_ /*44607*/;
assign _31956_ = _31957_ | _31959_ /*44604*/;
assign _31961_ = ~Q[28] /*44603*/;
assign _31960_ = _31961_ & D[25] /*44602*/;
assign _31963_ = _31322_ & _31960_ /*44597*/;
assign _31964_ = _31322_ ^ _31960_ /*44600*/;
assign _31965_ = _31956_ & _31964_ /*44598*/;
assign _31770_ = _31956_ ^ _31964_ /*44599*/;
assign _31962_ = _31963_ | _31965_ /*44596*/;
assign _31967_ = ~Q[28] /*44595*/;
assign _31966_ = _31967_ & D[26] /*44594*/;
assign _31969_ = _31323_ & _31966_ /*44589*/;
assign _31970_ = _31323_ ^ _31966_ /*44592*/;
assign _31971_ = _31962_ & _31970_ /*44590*/;
assign _31771_ = _31962_ ^ _31970_ /*44591*/;
assign _31968_ = _31969_ | _31971_ /*44588*/;
assign _31973_ = ~Q[28] /*44587*/;
assign _31972_ = _31973_ & D[27] /*44586*/;
assign _31975_ = _31324_ & _31972_ /*44581*/;
assign _31976_ = _31324_ ^ _31972_ /*44584*/;
assign _31977_ = _31968_ & _31976_ /*44582*/;
assign _31772_ = _31968_ ^ _31976_ /*44583*/;
assign _31974_ = _31975_ | _31977_ /*44580*/;
assign _31979_ = ~Q[28] /*44579*/;
assign _31978_ = _31979_ & D[28] /*44578*/;
assign _31981_ = _31325_ & _31978_ /*44573*/;
assign _31982_ = _31325_ ^ _31978_ /*44576*/;
assign _31983_ = _31974_ & _31982_ /*44574*/;
assign _31773_ = _31974_ ^ _31982_ /*44575*/;
assign _31980_ = _31981_ | _31983_ /*44572*/;
assign _31985_ = ~Q[28] /*44571*/;
assign _31984_ = _31985_ & D[29] /*44570*/;
assign _31987_ = _31326_ & _31984_ /*44565*/;
assign _31988_ = _31326_ ^ _31984_ /*44568*/;
assign _31989_ = _31980_ & _31988_ /*44566*/;
assign _31774_ = _31980_ ^ _31988_ /*44567*/;
assign _31986_ = _31987_ | _31989_ /*44564*/;
assign _31991_ = ~Q[28] /*44563*/;
assign _31990_ = _31991_ & D[30] /*44562*/;
assign _31993_ = _31327_ & _31990_ /*44557*/;
assign _31994_ = _31327_ ^ _31990_ /*44560*/;
assign _31995_ = _31986_ & _31994_ /*44558*/;
assign _31775_ = _31986_ ^ _31994_ /*44559*/;
assign _31992_ = _31993_ | _31995_ /*44556*/;
assign _31997_ = ~Q[28] /*44555*/;
assign _31996_ = _31997_ & D[31] /*44554*/;
assign _31999_ = _31328_ & _31996_ /*44549*/;
assign _32000_ = _31328_ ^ _31996_ /*44552*/;
assign _32001_ = _31992_ & _32000_ /*44550*/;
assign _31776_ = _31992_ ^ _32000_ /*44551*/;
assign _31998_ = _31999_ | _32001_ /*44548*/;
assign _32003_ = ~Q[28] /*44547*/;
assign _32002_ = _32003_ & D[32] /*44546*/;
assign _32005_ = _31329_ & _32002_ /*44541*/;
assign _32006_ = _31329_ ^ _32002_ /*44544*/;
assign _32007_ = _31998_ & _32006_ /*44542*/;
assign _31777_ = _31998_ ^ _32006_ /*44543*/;
assign _32004_ = _32005_ | _32007_ /*44540*/;
assign _32009_ = ~Q[28] /*44539*/;
assign _32008_ = _32009_ & D[33] /*44538*/;
assign _32011_ = _31330_ & _32008_ /*44533*/;
assign _32012_ = _31330_ ^ _32008_ /*44536*/;
assign _32013_ = _32004_ & _32012_ /*44534*/;
assign _31778_ = _32004_ ^ _32012_ /*44535*/;
assign _32010_ = _32011_ | _32013_ /*44532*/;
assign _32015_ = ~Q[28] /*44531*/;
assign _32014_ = _32015_ & D[34] /*44530*/;
assign _32017_ = _31331_ & _32014_ /*44525*/;
assign _32018_ = _31331_ ^ _32014_ /*44528*/;
assign _32019_ = _32010_ & _32018_ /*44526*/;
assign _31779_ = _32010_ ^ _32018_ /*44527*/;
assign _32016_ = _32017_ | _32019_ /*44524*/;
assign _32021_ = ~Q[28] /*44523*/;
assign _32020_ = _32021_ & D[35] /*44522*/;
assign _32023_ = _31332_ & _32020_ /*44517*/;
assign _32024_ = _31332_ ^ _32020_ /*44520*/;
assign _32025_ = _32016_ & _32024_ /*44518*/;
assign _31780_ = _32016_ ^ _32024_ /*44519*/;
assign _32022_ = _32023_ | _32025_ /*44516*/;
assign _32027_ = ~Q[28] /*44515*/;
assign _32026_ = _32027_ & D[36] /*44514*/;
assign _32029_ = _31333_ & _32026_ /*44509*/;
assign _32030_ = _31333_ ^ _32026_ /*44512*/;
assign _32031_ = _32022_ & _32030_ /*44510*/;
assign _31781_ = _32022_ ^ _32030_ /*44511*/;
assign _32028_ = _32029_ | _32031_ /*44508*/;
assign _32033_ = ~Q[28] /*44507*/;
assign _32032_ = _32033_ & D[37] /*44506*/;
assign _32035_ = _31334_ & _32032_ /*44501*/;
assign _32036_ = _31334_ ^ _32032_ /*44504*/;
assign _32037_ = _32028_ & _32036_ /*44502*/;
assign _31782_ = _32028_ ^ _32036_ /*44503*/;
assign _32034_ = _32035_ | _32037_ /*44500*/;
assign _32039_ = ~Q[28] /*44499*/;
assign _32038_ = _32039_ & D[38] /*44498*/;
assign _32041_ = _31335_ & _32038_ /*44493*/;
assign _32042_ = _31335_ ^ _32038_ /*44496*/;
assign _32043_ = _32034_ & _32042_ /*44494*/;
assign _31783_ = _32034_ ^ _32042_ /*44495*/;
assign _32040_ = _32041_ | _32043_ /*44492*/;
assign _32045_ = ~Q[28] /*44491*/;
assign _32044_ = _32045_ & D[39] /*44490*/;
assign _32047_ = _31336_ & _32044_ /*44485*/;
assign _32048_ = _31336_ ^ _32044_ /*44488*/;
assign _32049_ = _32040_ & _32048_ /*44486*/;
assign _31784_ = _32040_ ^ _32048_ /*44487*/;
assign _32046_ = _32047_ | _32049_ /*44484*/;
assign _32051_ = ~Q[28] /*44483*/;
assign _32050_ = _32051_ & D[40] /*44482*/;
assign _32053_ = _31337_ & _32050_ /*44477*/;
assign _32054_ = _31337_ ^ _32050_ /*44480*/;
assign _32055_ = _32046_ & _32054_ /*44478*/;
assign _31785_ = _32046_ ^ _32054_ /*44479*/;
assign _32052_ = _32053_ | _32055_ /*44476*/;
assign _32057_ = ~Q[28] /*44475*/;
assign _32056_ = _32057_ & D[41] /*44474*/;
assign _32059_ = _31338_ & _32056_ /*44469*/;
assign _32060_ = _31338_ ^ _32056_ /*44472*/;
assign _32061_ = _32052_ & _32060_ /*44470*/;
assign _31786_ = _32052_ ^ _32060_ /*44471*/;
assign _32058_ = _32059_ | _32061_ /*44468*/;
assign _32063_ = ~Q[28] /*44467*/;
assign _32062_ = _32063_ & D[42] /*44466*/;
assign _32065_ = _31339_ & _32062_ /*44461*/;
assign _32066_ = _31339_ ^ _32062_ /*44464*/;
assign _32067_ = _32058_ & _32066_ /*44462*/;
assign _31787_ = _32058_ ^ _32066_ /*44463*/;
assign _32064_ = _32065_ | _32067_ /*44460*/;
assign _32069_ = ~Q[28] /*44459*/;
assign _32068_ = _32069_ & D[43] /*44458*/;
assign _32071_ = _31340_ & _32068_ /*44453*/;
assign _32072_ = _31340_ ^ _32068_ /*44456*/;
assign _32073_ = _32064_ & _32072_ /*44454*/;
assign _31788_ = _32064_ ^ _32072_ /*44455*/;
assign _32070_ = _32071_ | _32073_ /*44452*/;
assign _32075_ = ~Q[28] /*44451*/;
assign _32074_ = _32075_ & D[44] /*44450*/;
assign _32077_ = _31341_ & _32074_ /*44445*/;
assign _32078_ = _31341_ ^ _32074_ /*44448*/;
assign _32079_ = _32070_ & _32078_ /*44446*/;
assign _31789_ = _32070_ ^ _32078_ /*44447*/;
assign _32076_ = _32077_ | _32079_ /*44444*/;
assign _32081_ = ~Q[28] /*44443*/;
assign _32080_ = _32081_ & D[45] /*44442*/;
assign _32083_ = _31342_ & _32080_ /*44437*/;
assign _32084_ = _31342_ ^ _32080_ /*44440*/;
assign _32085_ = _32076_ & _32084_ /*44438*/;
assign _31790_ = _32076_ ^ _32084_ /*44439*/;
assign _32082_ = _32083_ | _32085_ /*44436*/;
assign _32087_ = ~Q[28] /*44435*/;
assign _32086_ = _32087_ & D[46] /*44434*/;
assign _32089_ = _31343_ & _32086_ /*44429*/;
assign _32090_ = _31343_ ^ _32086_ /*44432*/;
assign _32091_ = _32082_ & _32090_ /*44430*/;
assign _31791_ = _32082_ ^ _32090_ /*44431*/;
assign _32088_ = _32089_ | _32091_ /*44428*/;
assign _32093_ = ~Q[28] /*44427*/;
assign _32092_ = _32093_ & D[47] /*44426*/;
assign _32095_ = _31344_ & _32092_ /*44421*/;
assign _32096_ = _31344_ ^ _32092_ /*44424*/;
assign _32097_ = _32088_ & _32096_ /*44422*/;
assign _31792_ = _32088_ ^ _32096_ /*44423*/;
assign _32094_ = _32095_ | _32097_ /*44420*/;
assign _32099_ = ~Q[28] /*44419*/;
assign _32098_ = _32099_ & D[48] /*44418*/;
assign _32101_ = _31345_ & _32098_ /*44413*/;
assign _32102_ = _31345_ ^ _32098_ /*44416*/;
assign _32103_ = _32094_ & _32102_ /*44414*/;
assign _31793_ = _32094_ ^ _32102_ /*44415*/;
assign _32100_ = _32101_ | _32103_ /*44412*/;
assign _32105_ = ~Q[28] /*44411*/;
assign _32104_ = _32105_ & D[49] /*44410*/;
assign _32107_ = _31346_ & _32104_ /*44405*/;
assign _32108_ = _31346_ ^ _32104_ /*44408*/;
assign _32109_ = _32100_ & _32108_ /*44406*/;
assign _31794_ = _32100_ ^ _32108_ /*44407*/;
assign _32106_ = _32107_ | _32109_ /*44404*/;
assign _32111_ = ~Q[28] /*44403*/;
assign _32110_ = _32111_ & D[50] /*44402*/;
assign _32113_ = _31347_ & _32110_ /*44397*/;
assign _32114_ = _31347_ ^ _32110_ /*44400*/;
assign _32115_ = _32106_ & _32114_ /*44398*/;
assign _31795_ = _32106_ ^ _32114_ /*44399*/;
assign _32112_ = _32113_ | _32115_ /*44396*/;
assign _32117_ = ~Q[28] /*44395*/;
assign _32116_ = _32117_ & D[51] /*44394*/;
assign _32119_ = _31348_ & _32116_ /*44389*/;
assign _32120_ = _31348_ ^ _32116_ /*44392*/;
assign _32121_ = _32112_ & _32120_ /*44390*/;
assign _31796_ = _32112_ ^ _32120_ /*44391*/;
assign _32118_ = _32119_ | _32121_ /*44388*/;
assign _32123_ = ~Q[28] /*44387*/;
assign _32122_ = _32123_ & D[52] /*44386*/;
assign _32125_ = _31349_ & _32122_ /*44381*/;
assign _32126_ = _31349_ ^ _32122_ /*44384*/;
assign _32127_ = _32118_ & _32126_ /*44382*/;
assign _31797_ = _32118_ ^ _32126_ /*44383*/;
assign _32124_ = _32125_ | _32127_ /*44380*/;
assign _32129_ = ~Q[28] /*44379*/;
assign _32128_ = _32129_ & D[53] /*44378*/;
assign _32131_ = _31350_ & _32128_ /*44373*/;
assign _32132_ = _31350_ ^ _32128_ /*44376*/;
assign _32133_ = _32124_ & _32132_ /*44374*/;
assign _31798_ = _32124_ ^ _32132_ /*44375*/;
assign _32130_ = _32131_ | _32133_ /*44372*/;
assign _32135_ = ~Q[28] /*44371*/;
assign _32134_ = _32135_ & D[54] /*44370*/;
assign _32137_ = _31351_ & _32134_ /*44365*/;
assign _32138_ = _31351_ ^ _32134_ /*44368*/;
assign _32139_ = _32130_ & _32138_ /*44366*/;
assign _31799_ = _32130_ ^ _32138_ /*44367*/;
assign _32136_ = _32137_ | _32139_ /*44364*/;
assign _32141_ = ~Q[28] /*44363*/;
assign _32140_ = _32141_ & D[55] /*44362*/;
assign _32143_ = _31352_ & _32140_ /*44357*/;
assign _32144_ = _31352_ ^ _32140_ /*44360*/;
assign _32145_ = _32136_ & _32144_ /*44358*/;
assign _31800_ = _32136_ ^ _32144_ /*44359*/;
assign _32142_ = _32143_ | _32145_ /*44356*/;
assign _32147_ = ~Q[28] /*44355*/;
assign _32146_ = _32147_ & D[56] /*44354*/;
assign _32149_ = _31353_ & _32146_ /*44349*/;
assign _32150_ = _31353_ ^ _32146_ /*44352*/;
assign _32151_ = _32142_ & _32150_ /*44350*/;
assign _31801_ = _32142_ ^ _32150_ /*44351*/;
assign _32148_ = _32149_ | _32151_ /*44348*/;
assign _32153_ = ~Q[28] /*44347*/;
assign _32152_ = _32153_ & D[57] /*44346*/;
assign _32155_ = _31354_ & _32152_ /*44341*/;
assign _32156_ = _31354_ ^ _32152_ /*44344*/;
assign _32157_ = _32148_ & _32156_ /*44342*/;
assign _31802_ = _32148_ ^ _32156_ /*44343*/;
assign _32154_ = _32155_ | _32157_ /*44340*/;
assign _32159_ = ~Q[28] /*44339*/;
assign _32158_ = _32159_ & D[58] /*44338*/;
assign _32161_ = _31355_ & _32158_ /*44333*/;
assign _32162_ = _31355_ ^ _32158_ /*44336*/;
assign _32163_ = _32154_ & _32162_ /*44334*/;
assign _31803_ = _32154_ ^ _32162_ /*44335*/;
assign _32160_ = _32161_ | _32163_ /*44332*/;
assign _32165_ = ~Q[28] /*44331*/;
assign _32164_ = _32165_ & D[59] /*44330*/;
assign _32167_ = _31356_ & _32164_ /*44325*/;
assign _32168_ = _31356_ ^ _32164_ /*44328*/;
assign _32169_ = _32160_ & _32168_ /*44326*/;
assign _31804_ = _32160_ ^ _32168_ /*44327*/;
assign _32166_ = _32167_ | _32169_ /*44324*/;
assign _32171_ = ~Q[28] /*44323*/;
assign _32170_ = _32171_ & D[60] /*44322*/;
assign _32173_ = _31357_ & _32170_ /*44317*/;
assign _32174_ = _31357_ ^ _32170_ /*44320*/;
assign _32175_ = _32166_ & _32174_ /*44318*/;
assign _31805_ = _32166_ ^ _32174_ /*44319*/;
assign _32172_ = _32173_ | _32175_ /*44316*/;
assign _32177_ = ~Q[28] /*44315*/;
assign _32176_ = _32177_ & D[61] /*44314*/;
assign _32179_ = _31358_ & _32176_ /*44309*/;
assign _32180_ = _31358_ ^ _32176_ /*44312*/;
assign _32181_ = _32172_ & _32180_ /*44310*/;
assign _31806_ = _32172_ ^ _32180_ /*44311*/;
assign _32178_ = _32179_ | _32181_ /*44308*/;
assign _32183_ = ~Q[28] /*44307*/;
assign _32182_ = _32183_ & D[62] /*44306*/;
assign _32185_ = _31359_ & _32182_ /*44301*/;
assign _32186_ = _31359_ ^ _32182_ /*44304*/;
assign _32187_ = _32178_ & _32186_ /*44302*/;
assign _31807_ = _32178_ ^ _32186_ /*44303*/;
assign _32184_ = _32185_ | _32187_ /*44300*/;
assign _32189_ = ~Q[28] /*44299*/;
assign _32188_ = _32189_ & zeroWire /*44298*/;
assign _32190_ = _31360_ ^ _32188_ /*44296*/;
assign _31808_ = _32190_ ^ _32184_ /*44295*/;
assign _32261_ = ~D[0] /*44041*/;
assign _32258_ = R_0[27] & _32261_ /*44037*/;
assign _32259_ = R_0[27] ^ _32261_ /*44040*/;
assign _32260_ = oneWire & _32259_ /*44038*/;
assign _32193_ = oneWire ^ _32259_ /*44039*/;
assign _32257_ = _32258_ | _32260_ /*44036*/;
assign _32266_ = ~D[1] /*44035*/;
assign _32263_ = _31745_ & _32266_ /*44031*/;
assign _32264_ = _31745_ ^ _32266_ /*44034*/;
assign _32265_ = _32257_ & _32264_ /*44032*/;
assign _32194_ = _32257_ ^ _32264_ /*44033*/;
assign _32262_ = _32263_ | _32265_ /*44030*/;
assign _32271_ = ~D[2] /*44029*/;
assign _32268_ = _31746_ & _32271_ /*44025*/;
assign _32269_ = _31746_ ^ _32271_ /*44028*/;
assign _32270_ = _32262_ & _32269_ /*44026*/;
assign _32195_ = _32262_ ^ _32269_ /*44027*/;
assign _32267_ = _32268_ | _32270_ /*44024*/;
assign _32276_ = ~D[3] /*44023*/;
assign _32273_ = _31747_ & _32276_ /*44019*/;
assign _32274_ = _31747_ ^ _32276_ /*44022*/;
assign _32275_ = _32267_ & _32274_ /*44020*/;
assign _32196_ = _32267_ ^ _32274_ /*44021*/;
assign _32272_ = _32273_ | _32275_ /*44018*/;
assign _32281_ = ~D[4] /*44017*/;
assign _32278_ = _31748_ & _32281_ /*44013*/;
assign _32279_ = _31748_ ^ _32281_ /*44016*/;
assign _32280_ = _32272_ & _32279_ /*44014*/;
assign _32197_ = _32272_ ^ _32279_ /*44015*/;
assign _32277_ = _32278_ | _32280_ /*44012*/;
assign _32286_ = ~D[5] /*44011*/;
assign _32283_ = _31749_ & _32286_ /*44007*/;
assign _32284_ = _31749_ ^ _32286_ /*44010*/;
assign _32285_ = _32277_ & _32284_ /*44008*/;
assign _32198_ = _32277_ ^ _32284_ /*44009*/;
assign _32282_ = _32283_ | _32285_ /*44006*/;
assign _32291_ = ~D[6] /*44005*/;
assign _32288_ = _31750_ & _32291_ /*44001*/;
assign _32289_ = _31750_ ^ _32291_ /*44004*/;
assign _32290_ = _32282_ & _32289_ /*44002*/;
assign _32199_ = _32282_ ^ _32289_ /*44003*/;
assign _32287_ = _32288_ | _32290_ /*44000*/;
assign _32296_ = ~D[7] /*43999*/;
assign _32293_ = _31751_ & _32296_ /*43995*/;
assign _32294_ = _31751_ ^ _32296_ /*43998*/;
assign _32295_ = _32287_ & _32294_ /*43996*/;
assign _32200_ = _32287_ ^ _32294_ /*43997*/;
assign _32292_ = _32293_ | _32295_ /*43994*/;
assign _32301_ = ~D[8] /*43993*/;
assign _32298_ = _31752_ & _32301_ /*43989*/;
assign _32299_ = _31752_ ^ _32301_ /*43992*/;
assign _32300_ = _32292_ & _32299_ /*43990*/;
assign _32201_ = _32292_ ^ _32299_ /*43991*/;
assign _32297_ = _32298_ | _32300_ /*43988*/;
assign _32306_ = ~D[9] /*43987*/;
assign _32303_ = _31753_ & _32306_ /*43983*/;
assign _32304_ = _31753_ ^ _32306_ /*43986*/;
assign _32305_ = _32297_ & _32304_ /*43984*/;
assign _32202_ = _32297_ ^ _32304_ /*43985*/;
assign _32302_ = _32303_ | _32305_ /*43982*/;
assign _32311_ = ~D[10] /*43981*/;
assign _32308_ = _31754_ & _32311_ /*43977*/;
assign _32309_ = _31754_ ^ _32311_ /*43980*/;
assign _32310_ = _32302_ & _32309_ /*43978*/;
assign _32203_ = _32302_ ^ _32309_ /*43979*/;
assign _32307_ = _32308_ | _32310_ /*43976*/;
assign _32316_ = ~D[11] /*43975*/;
assign _32313_ = _31755_ & _32316_ /*43971*/;
assign _32314_ = _31755_ ^ _32316_ /*43974*/;
assign _32315_ = _32307_ & _32314_ /*43972*/;
assign _32204_ = _32307_ ^ _32314_ /*43973*/;
assign _32312_ = _32313_ | _32315_ /*43970*/;
assign _32321_ = ~D[12] /*43969*/;
assign _32318_ = _31756_ & _32321_ /*43965*/;
assign _32319_ = _31756_ ^ _32321_ /*43968*/;
assign _32320_ = _32312_ & _32319_ /*43966*/;
assign _32205_ = _32312_ ^ _32319_ /*43967*/;
assign _32317_ = _32318_ | _32320_ /*43964*/;
assign _32326_ = ~D[13] /*43963*/;
assign _32323_ = _31757_ & _32326_ /*43959*/;
assign _32324_ = _31757_ ^ _32326_ /*43962*/;
assign _32325_ = _32317_ & _32324_ /*43960*/;
assign _32206_ = _32317_ ^ _32324_ /*43961*/;
assign _32322_ = _32323_ | _32325_ /*43958*/;
assign _32331_ = ~D[14] /*43957*/;
assign _32328_ = _31758_ & _32331_ /*43953*/;
assign _32329_ = _31758_ ^ _32331_ /*43956*/;
assign _32330_ = _32322_ & _32329_ /*43954*/;
assign _32207_ = _32322_ ^ _32329_ /*43955*/;
assign _32327_ = _32328_ | _32330_ /*43952*/;
assign _32336_ = ~D[15] /*43951*/;
assign _32333_ = _31759_ & _32336_ /*43947*/;
assign _32334_ = _31759_ ^ _32336_ /*43950*/;
assign _32335_ = _32327_ & _32334_ /*43948*/;
assign _32208_ = _32327_ ^ _32334_ /*43949*/;
assign _32332_ = _32333_ | _32335_ /*43946*/;
assign _32341_ = ~D[16] /*43945*/;
assign _32338_ = _31760_ & _32341_ /*43941*/;
assign _32339_ = _31760_ ^ _32341_ /*43944*/;
assign _32340_ = _32332_ & _32339_ /*43942*/;
assign _32209_ = _32332_ ^ _32339_ /*43943*/;
assign _32337_ = _32338_ | _32340_ /*43940*/;
assign _32346_ = ~D[17] /*43939*/;
assign _32343_ = _31761_ & _32346_ /*43935*/;
assign _32344_ = _31761_ ^ _32346_ /*43938*/;
assign _32345_ = _32337_ & _32344_ /*43936*/;
assign _32210_ = _32337_ ^ _32344_ /*43937*/;
assign _32342_ = _32343_ | _32345_ /*43934*/;
assign _32351_ = ~D[18] /*43933*/;
assign _32348_ = _31762_ & _32351_ /*43929*/;
assign _32349_ = _31762_ ^ _32351_ /*43932*/;
assign _32350_ = _32342_ & _32349_ /*43930*/;
assign _32211_ = _32342_ ^ _32349_ /*43931*/;
assign _32347_ = _32348_ | _32350_ /*43928*/;
assign _32356_ = ~D[19] /*43927*/;
assign _32353_ = _31763_ & _32356_ /*43923*/;
assign _32354_ = _31763_ ^ _32356_ /*43926*/;
assign _32355_ = _32347_ & _32354_ /*43924*/;
assign _32212_ = _32347_ ^ _32354_ /*43925*/;
assign _32352_ = _32353_ | _32355_ /*43922*/;
assign _32361_ = ~D[20] /*43921*/;
assign _32358_ = _31764_ & _32361_ /*43917*/;
assign _32359_ = _31764_ ^ _32361_ /*43920*/;
assign _32360_ = _32352_ & _32359_ /*43918*/;
assign _32213_ = _32352_ ^ _32359_ /*43919*/;
assign _32357_ = _32358_ | _32360_ /*43916*/;
assign _32366_ = ~D[21] /*43915*/;
assign _32363_ = _31765_ & _32366_ /*43911*/;
assign _32364_ = _31765_ ^ _32366_ /*43914*/;
assign _32365_ = _32357_ & _32364_ /*43912*/;
assign _32214_ = _32357_ ^ _32364_ /*43913*/;
assign _32362_ = _32363_ | _32365_ /*43910*/;
assign _32371_ = ~D[22] /*43909*/;
assign _32368_ = _31766_ & _32371_ /*43905*/;
assign _32369_ = _31766_ ^ _32371_ /*43908*/;
assign _32370_ = _32362_ & _32369_ /*43906*/;
assign _32215_ = _32362_ ^ _32369_ /*43907*/;
assign _32367_ = _32368_ | _32370_ /*43904*/;
assign _32376_ = ~D[23] /*43903*/;
assign _32373_ = _31767_ & _32376_ /*43899*/;
assign _32374_ = _31767_ ^ _32376_ /*43902*/;
assign _32375_ = _32367_ & _32374_ /*43900*/;
assign _32216_ = _32367_ ^ _32374_ /*43901*/;
assign _32372_ = _32373_ | _32375_ /*43898*/;
assign _32381_ = ~D[24] /*43897*/;
assign _32378_ = _31768_ & _32381_ /*43893*/;
assign _32379_ = _31768_ ^ _32381_ /*43896*/;
assign _32380_ = _32372_ & _32379_ /*43894*/;
assign _32217_ = _32372_ ^ _32379_ /*43895*/;
assign _32377_ = _32378_ | _32380_ /*43892*/;
assign _32386_ = ~D[25] /*43891*/;
assign _32383_ = _31769_ & _32386_ /*43887*/;
assign _32384_ = _31769_ ^ _32386_ /*43890*/;
assign _32385_ = _32377_ & _32384_ /*43888*/;
assign _32218_ = _32377_ ^ _32384_ /*43889*/;
assign _32382_ = _32383_ | _32385_ /*43886*/;
assign _32391_ = ~D[26] /*43885*/;
assign _32388_ = _31770_ & _32391_ /*43881*/;
assign _32389_ = _31770_ ^ _32391_ /*43884*/;
assign _32390_ = _32382_ & _32389_ /*43882*/;
assign _32219_ = _32382_ ^ _32389_ /*43883*/;
assign _32387_ = _32388_ | _32390_ /*43880*/;
assign _32396_ = ~D[27] /*43879*/;
assign _32393_ = _31771_ & _32396_ /*43875*/;
assign _32394_ = _31771_ ^ _32396_ /*43878*/;
assign _32395_ = _32387_ & _32394_ /*43876*/;
assign _32220_ = _32387_ ^ _32394_ /*43877*/;
assign _32392_ = _32393_ | _32395_ /*43874*/;
assign _32401_ = ~D[28] /*43873*/;
assign _32398_ = _31772_ & _32401_ /*43869*/;
assign _32399_ = _31772_ ^ _32401_ /*43872*/;
assign _32400_ = _32392_ & _32399_ /*43870*/;
assign _32221_ = _32392_ ^ _32399_ /*43871*/;
assign _32397_ = _32398_ | _32400_ /*43868*/;
assign _32406_ = ~D[29] /*43867*/;
assign _32403_ = _31773_ & _32406_ /*43863*/;
assign _32404_ = _31773_ ^ _32406_ /*43866*/;
assign _32405_ = _32397_ & _32404_ /*43864*/;
assign _32222_ = _32397_ ^ _32404_ /*43865*/;
assign _32402_ = _32403_ | _32405_ /*43862*/;
assign _32411_ = ~D[30] /*43861*/;
assign _32408_ = _31774_ & _32411_ /*43857*/;
assign _32409_ = _31774_ ^ _32411_ /*43860*/;
assign _32410_ = _32402_ & _32409_ /*43858*/;
assign _32223_ = _32402_ ^ _32409_ /*43859*/;
assign _32407_ = _32408_ | _32410_ /*43856*/;
assign _32416_ = ~D[31] /*43855*/;
assign _32413_ = _31775_ & _32416_ /*43851*/;
assign _32414_ = _31775_ ^ _32416_ /*43854*/;
assign _32415_ = _32407_ & _32414_ /*43852*/;
assign _32224_ = _32407_ ^ _32414_ /*43853*/;
assign _32412_ = _32413_ | _32415_ /*43850*/;
assign _32421_ = ~D[32] /*43849*/;
assign _32418_ = _31776_ & _32421_ /*43845*/;
assign _32419_ = _31776_ ^ _32421_ /*43848*/;
assign _32420_ = _32412_ & _32419_ /*43846*/;
assign _32225_ = _32412_ ^ _32419_ /*43847*/;
assign _32417_ = _32418_ | _32420_ /*43844*/;
assign _32426_ = ~D[33] /*43843*/;
assign _32423_ = _31777_ & _32426_ /*43839*/;
assign _32424_ = _31777_ ^ _32426_ /*43842*/;
assign _32425_ = _32417_ & _32424_ /*43840*/;
assign _32226_ = _32417_ ^ _32424_ /*43841*/;
assign _32422_ = _32423_ | _32425_ /*43838*/;
assign _32431_ = ~D[34] /*43837*/;
assign _32428_ = _31778_ & _32431_ /*43833*/;
assign _32429_ = _31778_ ^ _32431_ /*43836*/;
assign _32430_ = _32422_ & _32429_ /*43834*/;
assign _32227_ = _32422_ ^ _32429_ /*43835*/;
assign _32427_ = _32428_ | _32430_ /*43832*/;
assign _32436_ = ~D[35] /*43831*/;
assign _32433_ = _31779_ & _32436_ /*43827*/;
assign _32434_ = _31779_ ^ _32436_ /*43830*/;
assign _32435_ = _32427_ & _32434_ /*43828*/;
assign _32228_ = _32427_ ^ _32434_ /*43829*/;
assign _32432_ = _32433_ | _32435_ /*43826*/;
assign _32441_ = ~D[36] /*43825*/;
assign _32438_ = _31780_ & _32441_ /*43821*/;
assign _32439_ = _31780_ ^ _32441_ /*43824*/;
assign _32440_ = _32432_ & _32439_ /*43822*/;
assign _32229_ = _32432_ ^ _32439_ /*43823*/;
assign _32437_ = _32438_ | _32440_ /*43820*/;
assign _32446_ = ~D[37] /*43819*/;
assign _32443_ = _31781_ & _32446_ /*43815*/;
assign _32444_ = _31781_ ^ _32446_ /*43818*/;
assign _32445_ = _32437_ & _32444_ /*43816*/;
assign _32230_ = _32437_ ^ _32444_ /*43817*/;
assign _32442_ = _32443_ | _32445_ /*43814*/;
assign _32451_ = ~D[38] /*43813*/;
assign _32448_ = _31782_ & _32451_ /*43809*/;
assign _32449_ = _31782_ ^ _32451_ /*43812*/;
assign _32450_ = _32442_ & _32449_ /*43810*/;
assign _32231_ = _32442_ ^ _32449_ /*43811*/;
assign _32447_ = _32448_ | _32450_ /*43808*/;
assign _32456_ = ~D[39] /*43807*/;
assign _32453_ = _31783_ & _32456_ /*43803*/;
assign _32454_ = _31783_ ^ _32456_ /*43806*/;
assign _32455_ = _32447_ & _32454_ /*43804*/;
assign _32232_ = _32447_ ^ _32454_ /*43805*/;
assign _32452_ = _32453_ | _32455_ /*43802*/;
assign _32461_ = ~D[40] /*43801*/;
assign _32458_ = _31784_ & _32461_ /*43797*/;
assign _32459_ = _31784_ ^ _32461_ /*43800*/;
assign _32460_ = _32452_ & _32459_ /*43798*/;
assign _32233_ = _32452_ ^ _32459_ /*43799*/;
assign _32457_ = _32458_ | _32460_ /*43796*/;
assign _32466_ = ~D[41] /*43795*/;
assign _32463_ = _31785_ & _32466_ /*43791*/;
assign _32464_ = _31785_ ^ _32466_ /*43794*/;
assign _32465_ = _32457_ & _32464_ /*43792*/;
assign _32234_ = _32457_ ^ _32464_ /*43793*/;
assign _32462_ = _32463_ | _32465_ /*43790*/;
assign _32471_ = ~D[42] /*43789*/;
assign _32468_ = _31786_ & _32471_ /*43785*/;
assign _32469_ = _31786_ ^ _32471_ /*43788*/;
assign _32470_ = _32462_ & _32469_ /*43786*/;
assign _32235_ = _32462_ ^ _32469_ /*43787*/;
assign _32467_ = _32468_ | _32470_ /*43784*/;
assign _32476_ = ~D[43] /*43783*/;
assign _32473_ = _31787_ & _32476_ /*43779*/;
assign _32474_ = _31787_ ^ _32476_ /*43782*/;
assign _32475_ = _32467_ & _32474_ /*43780*/;
assign _32236_ = _32467_ ^ _32474_ /*43781*/;
assign _32472_ = _32473_ | _32475_ /*43778*/;
assign _32481_ = ~D[44] /*43777*/;
assign _32478_ = _31788_ & _32481_ /*43773*/;
assign _32479_ = _31788_ ^ _32481_ /*43776*/;
assign _32480_ = _32472_ & _32479_ /*43774*/;
assign _32237_ = _32472_ ^ _32479_ /*43775*/;
assign _32477_ = _32478_ | _32480_ /*43772*/;
assign _32486_ = ~D[45] /*43771*/;
assign _32483_ = _31789_ & _32486_ /*43767*/;
assign _32484_ = _31789_ ^ _32486_ /*43770*/;
assign _32485_ = _32477_ & _32484_ /*43768*/;
assign _32238_ = _32477_ ^ _32484_ /*43769*/;
assign _32482_ = _32483_ | _32485_ /*43766*/;
assign _32491_ = ~D[46] /*43765*/;
assign _32488_ = _31790_ & _32491_ /*43761*/;
assign _32489_ = _31790_ ^ _32491_ /*43764*/;
assign _32490_ = _32482_ & _32489_ /*43762*/;
assign _32239_ = _32482_ ^ _32489_ /*43763*/;
assign _32487_ = _32488_ | _32490_ /*43760*/;
assign _32496_ = ~D[47] /*43759*/;
assign _32493_ = _31791_ & _32496_ /*43755*/;
assign _32494_ = _31791_ ^ _32496_ /*43758*/;
assign _32495_ = _32487_ & _32494_ /*43756*/;
assign _32240_ = _32487_ ^ _32494_ /*43757*/;
assign _32492_ = _32493_ | _32495_ /*43754*/;
assign _32501_ = ~D[48] /*43753*/;
assign _32498_ = _31792_ & _32501_ /*43749*/;
assign _32499_ = _31792_ ^ _32501_ /*43752*/;
assign _32500_ = _32492_ & _32499_ /*43750*/;
assign _32241_ = _32492_ ^ _32499_ /*43751*/;
assign _32497_ = _32498_ | _32500_ /*43748*/;
assign _32506_ = ~D[49] /*43747*/;
assign _32503_ = _31793_ & _32506_ /*43743*/;
assign _32504_ = _31793_ ^ _32506_ /*43746*/;
assign _32505_ = _32497_ & _32504_ /*43744*/;
assign _32242_ = _32497_ ^ _32504_ /*43745*/;
assign _32502_ = _32503_ | _32505_ /*43742*/;
assign _32511_ = ~D[50] /*43741*/;
assign _32508_ = _31794_ & _32511_ /*43737*/;
assign _32509_ = _31794_ ^ _32511_ /*43740*/;
assign _32510_ = _32502_ & _32509_ /*43738*/;
assign _32243_ = _32502_ ^ _32509_ /*43739*/;
assign _32507_ = _32508_ | _32510_ /*43736*/;
assign _32516_ = ~D[51] /*43735*/;
assign _32513_ = _31795_ & _32516_ /*43731*/;
assign _32514_ = _31795_ ^ _32516_ /*43734*/;
assign _32515_ = _32507_ & _32514_ /*43732*/;
assign _32244_ = _32507_ ^ _32514_ /*43733*/;
assign _32512_ = _32513_ | _32515_ /*43730*/;
assign _32521_ = ~D[52] /*43729*/;
assign _32518_ = _31796_ & _32521_ /*43725*/;
assign _32519_ = _31796_ ^ _32521_ /*43728*/;
assign _32520_ = _32512_ & _32519_ /*43726*/;
assign _32245_ = _32512_ ^ _32519_ /*43727*/;
assign _32517_ = _32518_ | _32520_ /*43724*/;
assign _32526_ = ~D[53] /*43723*/;
assign _32523_ = _31797_ & _32526_ /*43719*/;
assign _32524_ = _31797_ ^ _32526_ /*43722*/;
assign _32525_ = _32517_ & _32524_ /*43720*/;
assign _32246_ = _32517_ ^ _32524_ /*43721*/;
assign _32522_ = _32523_ | _32525_ /*43718*/;
assign _32531_ = ~D[54] /*43717*/;
assign _32528_ = _31798_ & _32531_ /*43713*/;
assign _32529_ = _31798_ ^ _32531_ /*43716*/;
assign _32530_ = _32522_ & _32529_ /*43714*/;
assign _32247_ = _32522_ ^ _32529_ /*43715*/;
assign _32527_ = _32528_ | _32530_ /*43712*/;
assign _32536_ = ~D[55] /*43711*/;
assign _32533_ = _31799_ & _32536_ /*43707*/;
assign _32534_ = _31799_ ^ _32536_ /*43710*/;
assign _32535_ = _32527_ & _32534_ /*43708*/;
assign _32248_ = _32527_ ^ _32534_ /*43709*/;
assign _32532_ = _32533_ | _32535_ /*43706*/;
assign _32541_ = ~D[56] /*43705*/;
assign _32538_ = _31800_ & _32541_ /*43701*/;
assign _32539_ = _31800_ ^ _32541_ /*43704*/;
assign _32540_ = _32532_ & _32539_ /*43702*/;
assign _32249_ = _32532_ ^ _32539_ /*43703*/;
assign _32537_ = _32538_ | _32540_ /*43700*/;
assign _32546_ = ~D[57] /*43699*/;
assign _32543_ = _31801_ & _32546_ /*43695*/;
assign _32544_ = _31801_ ^ _32546_ /*43698*/;
assign _32545_ = _32537_ & _32544_ /*43696*/;
assign _32250_ = _32537_ ^ _32544_ /*43697*/;
assign _32542_ = _32543_ | _32545_ /*43694*/;
assign _32551_ = ~D[58] /*43693*/;
assign _32548_ = _31802_ & _32551_ /*43689*/;
assign _32549_ = _31802_ ^ _32551_ /*43692*/;
assign _32550_ = _32542_ & _32549_ /*43690*/;
assign _32251_ = _32542_ ^ _32549_ /*43691*/;
assign _32547_ = _32548_ | _32550_ /*43688*/;
assign _32556_ = ~D[59] /*43687*/;
assign _32553_ = _31803_ & _32556_ /*43683*/;
assign _32554_ = _31803_ ^ _32556_ /*43686*/;
assign _32555_ = _32547_ & _32554_ /*43684*/;
assign _32252_ = _32547_ ^ _32554_ /*43685*/;
assign _32552_ = _32553_ | _32555_ /*43682*/;
assign _32561_ = ~D[60] /*43681*/;
assign _32558_ = _31804_ & _32561_ /*43677*/;
assign _32559_ = _31804_ ^ _32561_ /*43680*/;
assign _32560_ = _32552_ & _32559_ /*43678*/;
assign _32253_ = _32552_ ^ _32559_ /*43679*/;
assign _32557_ = _32558_ | _32560_ /*43676*/;
assign _32566_ = ~D[61] /*43675*/;
assign _32563_ = _31805_ & _32566_ /*43671*/;
assign _32564_ = _31805_ ^ _32566_ /*43674*/;
assign _32565_ = _32557_ & _32564_ /*43672*/;
assign _32254_ = _32557_ ^ _32564_ /*43673*/;
assign _32562_ = _32563_ | _32565_ /*43670*/;
assign _32571_ = ~D[62] /*43669*/;
assign _32568_ = _31806_ & _32571_ /*43665*/;
assign _32569_ = _31806_ ^ _32571_ /*43668*/;
assign _32570_ = _32562_ & _32569_ /*43666*/;
assign _32255_ = _32562_ ^ _32569_ /*43667*/;
assign _32567_ = _32568_ | _32570_ /*43664*/;
assign _32572_ = _31807_ & oneWire /*43659*/;
assign _32573_ = _31807_ ^ oneWire /*43662*/;
assign _32574_ = _32567_ & _32573_ /*43660*/;
assign _32256_ = _32567_ ^ _32573_ /*43661*/;
assign Q[27] = _32572_ | _32574_ /*43658*/;
assign _32707_ = ~Q[27] /*43273*/;
assign _32706_ = _32707_ & D[0] /*43272*/;
assign _32709_ = _32193_ & _32706_ /*43267*/;
assign _32710_ = _32193_ ^ _32706_ /*43270*/;
assign _32711_ = zeroWire & _32710_ /*43268*/;
assign _32641_ = zeroWire ^ _32710_ /*43269*/;
assign _32708_ = _32709_ | _32711_ /*43266*/;
assign _32713_ = ~Q[27] /*43265*/;
assign _32712_ = _32713_ & D[1] /*43264*/;
assign _32715_ = _32194_ & _32712_ /*43259*/;
assign _32716_ = _32194_ ^ _32712_ /*43262*/;
assign _32717_ = _32708_ & _32716_ /*43260*/;
assign _32642_ = _32708_ ^ _32716_ /*43261*/;
assign _32714_ = _32715_ | _32717_ /*43258*/;
assign _32719_ = ~Q[27] /*43257*/;
assign _32718_ = _32719_ & D[2] /*43256*/;
assign _32721_ = _32195_ & _32718_ /*43251*/;
assign _32722_ = _32195_ ^ _32718_ /*43254*/;
assign _32723_ = _32714_ & _32722_ /*43252*/;
assign _32643_ = _32714_ ^ _32722_ /*43253*/;
assign _32720_ = _32721_ | _32723_ /*43250*/;
assign _32725_ = ~Q[27] /*43249*/;
assign _32724_ = _32725_ & D[3] /*43248*/;
assign _32727_ = _32196_ & _32724_ /*43243*/;
assign _32728_ = _32196_ ^ _32724_ /*43246*/;
assign _32729_ = _32720_ & _32728_ /*43244*/;
assign _32644_ = _32720_ ^ _32728_ /*43245*/;
assign _32726_ = _32727_ | _32729_ /*43242*/;
assign _32731_ = ~Q[27] /*43241*/;
assign _32730_ = _32731_ & D[4] /*43240*/;
assign _32733_ = _32197_ & _32730_ /*43235*/;
assign _32734_ = _32197_ ^ _32730_ /*43238*/;
assign _32735_ = _32726_ & _32734_ /*43236*/;
assign _32645_ = _32726_ ^ _32734_ /*43237*/;
assign _32732_ = _32733_ | _32735_ /*43234*/;
assign _32737_ = ~Q[27] /*43233*/;
assign _32736_ = _32737_ & D[5] /*43232*/;
assign _32739_ = _32198_ & _32736_ /*43227*/;
assign _32740_ = _32198_ ^ _32736_ /*43230*/;
assign _32741_ = _32732_ & _32740_ /*43228*/;
assign _32646_ = _32732_ ^ _32740_ /*43229*/;
assign _32738_ = _32739_ | _32741_ /*43226*/;
assign _32743_ = ~Q[27] /*43225*/;
assign _32742_ = _32743_ & D[6] /*43224*/;
assign _32745_ = _32199_ & _32742_ /*43219*/;
assign _32746_ = _32199_ ^ _32742_ /*43222*/;
assign _32747_ = _32738_ & _32746_ /*43220*/;
assign _32647_ = _32738_ ^ _32746_ /*43221*/;
assign _32744_ = _32745_ | _32747_ /*43218*/;
assign _32749_ = ~Q[27] /*43217*/;
assign _32748_ = _32749_ & D[7] /*43216*/;
assign _32751_ = _32200_ & _32748_ /*43211*/;
assign _32752_ = _32200_ ^ _32748_ /*43214*/;
assign _32753_ = _32744_ & _32752_ /*43212*/;
assign _32648_ = _32744_ ^ _32752_ /*43213*/;
assign _32750_ = _32751_ | _32753_ /*43210*/;
assign _32755_ = ~Q[27] /*43209*/;
assign _32754_ = _32755_ & D[8] /*43208*/;
assign _32757_ = _32201_ & _32754_ /*43203*/;
assign _32758_ = _32201_ ^ _32754_ /*43206*/;
assign _32759_ = _32750_ & _32758_ /*43204*/;
assign _32649_ = _32750_ ^ _32758_ /*43205*/;
assign _32756_ = _32757_ | _32759_ /*43202*/;
assign _32761_ = ~Q[27] /*43201*/;
assign _32760_ = _32761_ & D[9] /*43200*/;
assign _32763_ = _32202_ & _32760_ /*43195*/;
assign _32764_ = _32202_ ^ _32760_ /*43198*/;
assign _32765_ = _32756_ & _32764_ /*43196*/;
assign _32650_ = _32756_ ^ _32764_ /*43197*/;
assign _32762_ = _32763_ | _32765_ /*43194*/;
assign _32767_ = ~Q[27] /*43193*/;
assign _32766_ = _32767_ & D[10] /*43192*/;
assign _32769_ = _32203_ & _32766_ /*43187*/;
assign _32770_ = _32203_ ^ _32766_ /*43190*/;
assign _32771_ = _32762_ & _32770_ /*43188*/;
assign _32651_ = _32762_ ^ _32770_ /*43189*/;
assign _32768_ = _32769_ | _32771_ /*43186*/;
assign _32773_ = ~Q[27] /*43185*/;
assign _32772_ = _32773_ & D[11] /*43184*/;
assign _32775_ = _32204_ & _32772_ /*43179*/;
assign _32776_ = _32204_ ^ _32772_ /*43182*/;
assign _32777_ = _32768_ & _32776_ /*43180*/;
assign _32652_ = _32768_ ^ _32776_ /*43181*/;
assign _32774_ = _32775_ | _32777_ /*43178*/;
assign _32779_ = ~Q[27] /*43177*/;
assign _32778_ = _32779_ & D[12] /*43176*/;
assign _32781_ = _32205_ & _32778_ /*43171*/;
assign _32782_ = _32205_ ^ _32778_ /*43174*/;
assign _32783_ = _32774_ & _32782_ /*43172*/;
assign _32653_ = _32774_ ^ _32782_ /*43173*/;
assign _32780_ = _32781_ | _32783_ /*43170*/;
assign _32785_ = ~Q[27] /*43169*/;
assign _32784_ = _32785_ & D[13] /*43168*/;
assign _32787_ = _32206_ & _32784_ /*43163*/;
assign _32788_ = _32206_ ^ _32784_ /*43166*/;
assign _32789_ = _32780_ & _32788_ /*43164*/;
assign _32654_ = _32780_ ^ _32788_ /*43165*/;
assign _32786_ = _32787_ | _32789_ /*43162*/;
assign _32791_ = ~Q[27] /*43161*/;
assign _32790_ = _32791_ & D[14] /*43160*/;
assign _32793_ = _32207_ & _32790_ /*43155*/;
assign _32794_ = _32207_ ^ _32790_ /*43158*/;
assign _32795_ = _32786_ & _32794_ /*43156*/;
assign _32655_ = _32786_ ^ _32794_ /*43157*/;
assign _32792_ = _32793_ | _32795_ /*43154*/;
assign _32797_ = ~Q[27] /*43153*/;
assign _32796_ = _32797_ & D[15] /*43152*/;
assign _32799_ = _32208_ & _32796_ /*43147*/;
assign _32800_ = _32208_ ^ _32796_ /*43150*/;
assign _32801_ = _32792_ & _32800_ /*43148*/;
assign _32656_ = _32792_ ^ _32800_ /*43149*/;
assign _32798_ = _32799_ | _32801_ /*43146*/;
assign _32803_ = ~Q[27] /*43145*/;
assign _32802_ = _32803_ & D[16] /*43144*/;
assign _32805_ = _32209_ & _32802_ /*43139*/;
assign _32806_ = _32209_ ^ _32802_ /*43142*/;
assign _32807_ = _32798_ & _32806_ /*43140*/;
assign _32657_ = _32798_ ^ _32806_ /*43141*/;
assign _32804_ = _32805_ | _32807_ /*43138*/;
assign _32809_ = ~Q[27] /*43137*/;
assign _32808_ = _32809_ & D[17] /*43136*/;
assign _32811_ = _32210_ & _32808_ /*43131*/;
assign _32812_ = _32210_ ^ _32808_ /*43134*/;
assign _32813_ = _32804_ & _32812_ /*43132*/;
assign _32658_ = _32804_ ^ _32812_ /*43133*/;
assign _32810_ = _32811_ | _32813_ /*43130*/;
assign _32815_ = ~Q[27] /*43129*/;
assign _32814_ = _32815_ & D[18] /*43128*/;
assign _32817_ = _32211_ & _32814_ /*43123*/;
assign _32818_ = _32211_ ^ _32814_ /*43126*/;
assign _32819_ = _32810_ & _32818_ /*43124*/;
assign _32659_ = _32810_ ^ _32818_ /*43125*/;
assign _32816_ = _32817_ | _32819_ /*43122*/;
assign _32821_ = ~Q[27] /*43121*/;
assign _32820_ = _32821_ & D[19] /*43120*/;
assign _32823_ = _32212_ & _32820_ /*43115*/;
assign _32824_ = _32212_ ^ _32820_ /*43118*/;
assign _32825_ = _32816_ & _32824_ /*43116*/;
assign _32660_ = _32816_ ^ _32824_ /*43117*/;
assign _32822_ = _32823_ | _32825_ /*43114*/;
assign _32827_ = ~Q[27] /*43113*/;
assign _32826_ = _32827_ & D[20] /*43112*/;
assign _32829_ = _32213_ & _32826_ /*43107*/;
assign _32830_ = _32213_ ^ _32826_ /*43110*/;
assign _32831_ = _32822_ & _32830_ /*43108*/;
assign _32661_ = _32822_ ^ _32830_ /*43109*/;
assign _32828_ = _32829_ | _32831_ /*43106*/;
assign _32833_ = ~Q[27] /*43105*/;
assign _32832_ = _32833_ & D[21] /*43104*/;
assign _32835_ = _32214_ & _32832_ /*43099*/;
assign _32836_ = _32214_ ^ _32832_ /*43102*/;
assign _32837_ = _32828_ & _32836_ /*43100*/;
assign _32662_ = _32828_ ^ _32836_ /*43101*/;
assign _32834_ = _32835_ | _32837_ /*43098*/;
assign _32839_ = ~Q[27] /*43097*/;
assign _32838_ = _32839_ & D[22] /*43096*/;
assign _32841_ = _32215_ & _32838_ /*43091*/;
assign _32842_ = _32215_ ^ _32838_ /*43094*/;
assign _32843_ = _32834_ & _32842_ /*43092*/;
assign _32663_ = _32834_ ^ _32842_ /*43093*/;
assign _32840_ = _32841_ | _32843_ /*43090*/;
assign _32845_ = ~Q[27] /*43089*/;
assign _32844_ = _32845_ & D[23] /*43088*/;
assign _32847_ = _32216_ & _32844_ /*43083*/;
assign _32848_ = _32216_ ^ _32844_ /*43086*/;
assign _32849_ = _32840_ & _32848_ /*43084*/;
assign _32664_ = _32840_ ^ _32848_ /*43085*/;
assign _32846_ = _32847_ | _32849_ /*43082*/;
assign _32851_ = ~Q[27] /*43081*/;
assign _32850_ = _32851_ & D[24] /*43080*/;
assign _32853_ = _32217_ & _32850_ /*43075*/;
assign _32854_ = _32217_ ^ _32850_ /*43078*/;
assign _32855_ = _32846_ & _32854_ /*43076*/;
assign _32665_ = _32846_ ^ _32854_ /*43077*/;
assign _32852_ = _32853_ | _32855_ /*43074*/;
assign _32857_ = ~Q[27] /*43073*/;
assign _32856_ = _32857_ & D[25] /*43072*/;
assign _32859_ = _32218_ & _32856_ /*43067*/;
assign _32860_ = _32218_ ^ _32856_ /*43070*/;
assign _32861_ = _32852_ & _32860_ /*43068*/;
assign _32666_ = _32852_ ^ _32860_ /*43069*/;
assign _32858_ = _32859_ | _32861_ /*43066*/;
assign _32863_ = ~Q[27] /*43065*/;
assign _32862_ = _32863_ & D[26] /*43064*/;
assign _32865_ = _32219_ & _32862_ /*43059*/;
assign _32866_ = _32219_ ^ _32862_ /*43062*/;
assign _32867_ = _32858_ & _32866_ /*43060*/;
assign _32667_ = _32858_ ^ _32866_ /*43061*/;
assign _32864_ = _32865_ | _32867_ /*43058*/;
assign _32869_ = ~Q[27] /*43057*/;
assign _32868_ = _32869_ & D[27] /*43056*/;
assign _32871_ = _32220_ & _32868_ /*43051*/;
assign _32872_ = _32220_ ^ _32868_ /*43054*/;
assign _32873_ = _32864_ & _32872_ /*43052*/;
assign _32668_ = _32864_ ^ _32872_ /*43053*/;
assign _32870_ = _32871_ | _32873_ /*43050*/;
assign _32875_ = ~Q[27] /*43049*/;
assign _32874_ = _32875_ & D[28] /*43048*/;
assign _32877_ = _32221_ & _32874_ /*43043*/;
assign _32878_ = _32221_ ^ _32874_ /*43046*/;
assign _32879_ = _32870_ & _32878_ /*43044*/;
assign _32669_ = _32870_ ^ _32878_ /*43045*/;
assign _32876_ = _32877_ | _32879_ /*43042*/;
assign _32881_ = ~Q[27] /*43041*/;
assign _32880_ = _32881_ & D[29] /*43040*/;
assign _32883_ = _32222_ & _32880_ /*43035*/;
assign _32884_ = _32222_ ^ _32880_ /*43038*/;
assign _32885_ = _32876_ & _32884_ /*43036*/;
assign _32670_ = _32876_ ^ _32884_ /*43037*/;
assign _32882_ = _32883_ | _32885_ /*43034*/;
assign _32887_ = ~Q[27] /*43033*/;
assign _32886_ = _32887_ & D[30] /*43032*/;
assign _32889_ = _32223_ & _32886_ /*43027*/;
assign _32890_ = _32223_ ^ _32886_ /*43030*/;
assign _32891_ = _32882_ & _32890_ /*43028*/;
assign _32671_ = _32882_ ^ _32890_ /*43029*/;
assign _32888_ = _32889_ | _32891_ /*43026*/;
assign _32893_ = ~Q[27] /*43025*/;
assign _32892_ = _32893_ & D[31] /*43024*/;
assign _32895_ = _32224_ & _32892_ /*43019*/;
assign _32896_ = _32224_ ^ _32892_ /*43022*/;
assign _32897_ = _32888_ & _32896_ /*43020*/;
assign _32672_ = _32888_ ^ _32896_ /*43021*/;
assign _32894_ = _32895_ | _32897_ /*43018*/;
assign _32899_ = ~Q[27] /*43017*/;
assign _32898_ = _32899_ & D[32] /*43016*/;
assign _32901_ = _32225_ & _32898_ /*43011*/;
assign _32902_ = _32225_ ^ _32898_ /*43014*/;
assign _32903_ = _32894_ & _32902_ /*43012*/;
assign _32673_ = _32894_ ^ _32902_ /*43013*/;
assign _32900_ = _32901_ | _32903_ /*43010*/;
assign _32905_ = ~Q[27] /*43009*/;
assign _32904_ = _32905_ & D[33] /*43008*/;
assign _32907_ = _32226_ & _32904_ /*43003*/;
assign _32908_ = _32226_ ^ _32904_ /*43006*/;
assign _32909_ = _32900_ & _32908_ /*43004*/;
assign _32674_ = _32900_ ^ _32908_ /*43005*/;
assign _32906_ = _32907_ | _32909_ /*43002*/;
assign _32911_ = ~Q[27] /*43001*/;
assign _32910_ = _32911_ & D[34] /*43000*/;
assign _32913_ = _32227_ & _32910_ /*42995*/;
assign _32914_ = _32227_ ^ _32910_ /*42998*/;
assign _32915_ = _32906_ & _32914_ /*42996*/;
assign _32675_ = _32906_ ^ _32914_ /*42997*/;
assign _32912_ = _32913_ | _32915_ /*42994*/;
assign _32917_ = ~Q[27] /*42993*/;
assign _32916_ = _32917_ & D[35] /*42992*/;
assign _32919_ = _32228_ & _32916_ /*42987*/;
assign _32920_ = _32228_ ^ _32916_ /*42990*/;
assign _32921_ = _32912_ & _32920_ /*42988*/;
assign _32676_ = _32912_ ^ _32920_ /*42989*/;
assign _32918_ = _32919_ | _32921_ /*42986*/;
assign _32923_ = ~Q[27] /*42985*/;
assign _32922_ = _32923_ & D[36] /*42984*/;
assign _32925_ = _32229_ & _32922_ /*42979*/;
assign _32926_ = _32229_ ^ _32922_ /*42982*/;
assign _32927_ = _32918_ & _32926_ /*42980*/;
assign _32677_ = _32918_ ^ _32926_ /*42981*/;
assign _32924_ = _32925_ | _32927_ /*42978*/;
assign _32929_ = ~Q[27] /*42977*/;
assign _32928_ = _32929_ & D[37] /*42976*/;
assign _32931_ = _32230_ & _32928_ /*42971*/;
assign _32932_ = _32230_ ^ _32928_ /*42974*/;
assign _32933_ = _32924_ & _32932_ /*42972*/;
assign _32678_ = _32924_ ^ _32932_ /*42973*/;
assign _32930_ = _32931_ | _32933_ /*42970*/;
assign _32935_ = ~Q[27] /*42969*/;
assign _32934_ = _32935_ & D[38] /*42968*/;
assign _32937_ = _32231_ & _32934_ /*42963*/;
assign _32938_ = _32231_ ^ _32934_ /*42966*/;
assign _32939_ = _32930_ & _32938_ /*42964*/;
assign _32679_ = _32930_ ^ _32938_ /*42965*/;
assign _32936_ = _32937_ | _32939_ /*42962*/;
assign _32941_ = ~Q[27] /*42961*/;
assign _32940_ = _32941_ & D[39] /*42960*/;
assign _32943_ = _32232_ & _32940_ /*42955*/;
assign _32944_ = _32232_ ^ _32940_ /*42958*/;
assign _32945_ = _32936_ & _32944_ /*42956*/;
assign _32680_ = _32936_ ^ _32944_ /*42957*/;
assign _32942_ = _32943_ | _32945_ /*42954*/;
assign _32947_ = ~Q[27] /*42953*/;
assign _32946_ = _32947_ & D[40] /*42952*/;
assign _32949_ = _32233_ & _32946_ /*42947*/;
assign _32950_ = _32233_ ^ _32946_ /*42950*/;
assign _32951_ = _32942_ & _32950_ /*42948*/;
assign _32681_ = _32942_ ^ _32950_ /*42949*/;
assign _32948_ = _32949_ | _32951_ /*42946*/;
assign _32953_ = ~Q[27] /*42945*/;
assign _32952_ = _32953_ & D[41] /*42944*/;
assign _32955_ = _32234_ & _32952_ /*42939*/;
assign _32956_ = _32234_ ^ _32952_ /*42942*/;
assign _32957_ = _32948_ & _32956_ /*42940*/;
assign _32682_ = _32948_ ^ _32956_ /*42941*/;
assign _32954_ = _32955_ | _32957_ /*42938*/;
assign _32959_ = ~Q[27] /*42937*/;
assign _32958_ = _32959_ & D[42] /*42936*/;
assign _32961_ = _32235_ & _32958_ /*42931*/;
assign _32962_ = _32235_ ^ _32958_ /*42934*/;
assign _32963_ = _32954_ & _32962_ /*42932*/;
assign _32683_ = _32954_ ^ _32962_ /*42933*/;
assign _32960_ = _32961_ | _32963_ /*42930*/;
assign _32965_ = ~Q[27] /*42929*/;
assign _32964_ = _32965_ & D[43] /*42928*/;
assign _32967_ = _32236_ & _32964_ /*42923*/;
assign _32968_ = _32236_ ^ _32964_ /*42926*/;
assign _32969_ = _32960_ & _32968_ /*42924*/;
assign _32684_ = _32960_ ^ _32968_ /*42925*/;
assign _32966_ = _32967_ | _32969_ /*42922*/;
assign _32971_ = ~Q[27] /*42921*/;
assign _32970_ = _32971_ & D[44] /*42920*/;
assign _32973_ = _32237_ & _32970_ /*42915*/;
assign _32974_ = _32237_ ^ _32970_ /*42918*/;
assign _32975_ = _32966_ & _32974_ /*42916*/;
assign _32685_ = _32966_ ^ _32974_ /*42917*/;
assign _32972_ = _32973_ | _32975_ /*42914*/;
assign _32977_ = ~Q[27] /*42913*/;
assign _32976_ = _32977_ & D[45] /*42912*/;
assign _32979_ = _32238_ & _32976_ /*42907*/;
assign _32980_ = _32238_ ^ _32976_ /*42910*/;
assign _32981_ = _32972_ & _32980_ /*42908*/;
assign _32686_ = _32972_ ^ _32980_ /*42909*/;
assign _32978_ = _32979_ | _32981_ /*42906*/;
assign _32983_ = ~Q[27] /*42905*/;
assign _32982_ = _32983_ & D[46] /*42904*/;
assign _32985_ = _32239_ & _32982_ /*42899*/;
assign _32986_ = _32239_ ^ _32982_ /*42902*/;
assign _32987_ = _32978_ & _32986_ /*42900*/;
assign _32687_ = _32978_ ^ _32986_ /*42901*/;
assign _32984_ = _32985_ | _32987_ /*42898*/;
assign _32989_ = ~Q[27] /*42897*/;
assign _32988_ = _32989_ & D[47] /*42896*/;
assign _32991_ = _32240_ & _32988_ /*42891*/;
assign _32992_ = _32240_ ^ _32988_ /*42894*/;
assign _32993_ = _32984_ & _32992_ /*42892*/;
assign _32688_ = _32984_ ^ _32992_ /*42893*/;
assign _32990_ = _32991_ | _32993_ /*42890*/;
assign _32995_ = ~Q[27] /*42889*/;
assign _32994_ = _32995_ & D[48] /*42888*/;
assign _32997_ = _32241_ & _32994_ /*42883*/;
assign _32998_ = _32241_ ^ _32994_ /*42886*/;
assign _32999_ = _32990_ & _32998_ /*42884*/;
assign _32689_ = _32990_ ^ _32998_ /*42885*/;
assign _32996_ = _32997_ | _32999_ /*42882*/;
assign _33001_ = ~Q[27] /*42881*/;
assign _33000_ = _33001_ & D[49] /*42880*/;
assign _33003_ = _32242_ & _33000_ /*42875*/;
assign _33004_ = _32242_ ^ _33000_ /*42878*/;
assign _33005_ = _32996_ & _33004_ /*42876*/;
assign _32690_ = _32996_ ^ _33004_ /*42877*/;
assign _33002_ = _33003_ | _33005_ /*42874*/;
assign _33007_ = ~Q[27] /*42873*/;
assign _33006_ = _33007_ & D[50] /*42872*/;
assign _33009_ = _32243_ & _33006_ /*42867*/;
assign _33010_ = _32243_ ^ _33006_ /*42870*/;
assign _33011_ = _33002_ & _33010_ /*42868*/;
assign _32691_ = _33002_ ^ _33010_ /*42869*/;
assign _33008_ = _33009_ | _33011_ /*42866*/;
assign _33013_ = ~Q[27] /*42865*/;
assign _33012_ = _33013_ & D[51] /*42864*/;
assign _33015_ = _32244_ & _33012_ /*42859*/;
assign _33016_ = _32244_ ^ _33012_ /*42862*/;
assign _33017_ = _33008_ & _33016_ /*42860*/;
assign _32692_ = _33008_ ^ _33016_ /*42861*/;
assign _33014_ = _33015_ | _33017_ /*42858*/;
assign _33019_ = ~Q[27] /*42857*/;
assign _33018_ = _33019_ & D[52] /*42856*/;
assign _33021_ = _32245_ & _33018_ /*42851*/;
assign _33022_ = _32245_ ^ _33018_ /*42854*/;
assign _33023_ = _33014_ & _33022_ /*42852*/;
assign _32693_ = _33014_ ^ _33022_ /*42853*/;
assign _33020_ = _33021_ | _33023_ /*42850*/;
assign _33025_ = ~Q[27] /*42849*/;
assign _33024_ = _33025_ & D[53] /*42848*/;
assign _33027_ = _32246_ & _33024_ /*42843*/;
assign _33028_ = _32246_ ^ _33024_ /*42846*/;
assign _33029_ = _33020_ & _33028_ /*42844*/;
assign _32694_ = _33020_ ^ _33028_ /*42845*/;
assign _33026_ = _33027_ | _33029_ /*42842*/;
assign _33031_ = ~Q[27] /*42841*/;
assign _33030_ = _33031_ & D[54] /*42840*/;
assign _33033_ = _32247_ & _33030_ /*42835*/;
assign _33034_ = _32247_ ^ _33030_ /*42838*/;
assign _33035_ = _33026_ & _33034_ /*42836*/;
assign _32695_ = _33026_ ^ _33034_ /*42837*/;
assign _33032_ = _33033_ | _33035_ /*42834*/;
assign _33037_ = ~Q[27] /*42833*/;
assign _33036_ = _33037_ & D[55] /*42832*/;
assign _33039_ = _32248_ & _33036_ /*42827*/;
assign _33040_ = _32248_ ^ _33036_ /*42830*/;
assign _33041_ = _33032_ & _33040_ /*42828*/;
assign _32696_ = _33032_ ^ _33040_ /*42829*/;
assign _33038_ = _33039_ | _33041_ /*42826*/;
assign _33043_ = ~Q[27] /*42825*/;
assign _33042_ = _33043_ & D[56] /*42824*/;
assign _33045_ = _32249_ & _33042_ /*42819*/;
assign _33046_ = _32249_ ^ _33042_ /*42822*/;
assign _33047_ = _33038_ & _33046_ /*42820*/;
assign _32697_ = _33038_ ^ _33046_ /*42821*/;
assign _33044_ = _33045_ | _33047_ /*42818*/;
assign _33049_ = ~Q[27] /*42817*/;
assign _33048_ = _33049_ & D[57] /*42816*/;
assign _33051_ = _32250_ & _33048_ /*42811*/;
assign _33052_ = _32250_ ^ _33048_ /*42814*/;
assign _33053_ = _33044_ & _33052_ /*42812*/;
assign _32698_ = _33044_ ^ _33052_ /*42813*/;
assign _33050_ = _33051_ | _33053_ /*42810*/;
assign _33055_ = ~Q[27] /*42809*/;
assign _33054_ = _33055_ & D[58] /*42808*/;
assign _33057_ = _32251_ & _33054_ /*42803*/;
assign _33058_ = _32251_ ^ _33054_ /*42806*/;
assign _33059_ = _33050_ & _33058_ /*42804*/;
assign _32699_ = _33050_ ^ _33058_ /*42805*/;
assign _33056_ = _33057_ | _33059_ /*42802*/;
assign _33061_ = ~Q[27] /*42801*/;
assign _33060_ = _33061_ & D[59] /*42800*/;
assign _33063_ = _32252_ & _33060_ /*42795*/;
assign _33064_ = _32252_ ^ _33060_ /*42798*/;
assign _33065_ = _33056_ & _33064_ /*42796*/;
assign _32700_ = _33056_ ^ _33064_ /*42797*/;
assign _33062_ = _33063_ | _33065_ /*42794*/;
assign _33067_ = ~Q[27] /*42793*/;
assign _33066_ = _33067_ & D[60] /*42792*/;
assign _33069_ = _32253_ & _33066_ /*42787*/;
assign _33070_ = _32253_ ^ _33066_ /*42790*/;
assign _33071_ = _33062_ & _33070_ /*42788*/;
assign _32701_ = _33062_ ^ _33070_ /*42789*/;
assign _33068_ = _33069_ | _33071_ /*42786*/;
assign _33073_ = ~Q[27] /*42785*/;
assign _33072_ = _33073_ & D[61] /*42784*/;
assign _33075_ = _32254_ & _33072_ /*42779*/;
assign _33076_ = _32254_ ^ _33072_ /*42782*/;
assign _33077_ = _33068_ & _33076_ /*42780*/;
assign _32702_ = _33068_ ^ _33076_ /*42781*/;
assign _33074_ = _33075_ | _33077_ /*42778*/;
assign _33079_ = ~Q[27] /*42777*/;
assign _33078_ = _33079_ & D[62] /*42776*/;
assign _33081_ = _32255_ & _33078_ /*42771*/;
assign _33082_ = _32255_ ^ _33078_ /*42774*/;
assign _33083_ = _33074_ & _33082_ /*42772*/;
assign _32703_ = _33074_ ^ _33082_ /*42773*/;
assign _33080_ = _33081_ | _33083_ /*42770*/;
assign _33085_ = ~Q[27] /*42769*/;
assign _33084_ = _33085_ & zeroWire /*42768*/;
assign _33086_ = _32256_ ^ _33084_ /*42766*/;
assign _32704_ = _33086_ ^ _33080_ /*42765*/;
assign _33157_ = ~D[0] /*42511*/;
assign _33154_ = R_0[26] & _33157_ /*42507*/;
assign _33155_ = R_0[26] ^ _33157_ /*42510*/;
assign _33156_ = oneWire & _33155_ /*42508*/;
assign _33089_ = oneWire ^ _33155_ /*42509*/;
assign _33153_ = _33154_ | _33156_ /*42506*/;
assign _33162_ = ~D[1] /*42505*/;
assign _33159_ = _32641_ & _33162_ /*42501*/;
assign _33160_ = _32641_ ^ _33162_ /*42504*/;
assign _33161_ = _33153_ & _33160_ /*42502*/;
assign _33090_ = _33153_ ^ _33160_ /*42503*/;
assign _33158_ = _33159_ | _33161_ /*42500*/;
assign _33167_ = ~D[2] /*42499*/;
assign _33164_ = _32642_ & _33167_ /*42495*/;
assign _33165_ = _32642_ ^ _33167_ /*42498*/;
assign _33166_ = _33158_ & _33165_ /*42496*/;
assign _33091_ = _33158_ ^ _33165_ /*42497*/;
assign _33163_ = _33164_ | _33166_ /*42494*/;
assign _33172_ = ~D[3] /*42493*/;
assign _33169_ = _32643_ & _33172_ /*42489*/;
assign _33170_ = _32643_ ^ _33172_ /*42492*/;
assign _33171_ = _33163_ & _33170_ /*42490*/;
assign _33092_ = _33163_ ^ _33170_ /*42491*/;
assign _33168_ = _33169_ | _33171_ /*42488*/;
assign _33177_ = ~D[4] /*42487*/;
assign _33174_ = _32644_ & _33177_ /*42483*/;
assign _33175_ = _32644_ ^ _33177_ /*42486*/;
assign _33176_ = _33168_ & _33175_ /*42484*/;
assign _33093_ = _33168_ ^ _33175_ /*42485*/;
assign _33173_ = _33174_ | _33176_ /*42482*/;
assign _33182_ = ~D[5] /*42481*/;
assign _33179_ = _32645_ & _33182_ /*42477*/;
assign _33180_ = _32645_ ^ _33182_ /*42480*/;
assign _33181_ = _33173_ & _33180_ /*42478*/;
assign _33094_ = _33173_ ^ _33180_ /*42479*/;
assign _33178_ = _33179_ | _33181_ /*42476*/;
assign _33187_ = ~D[6] /*42475*/;
assign _33184_ = _32646_ & _33187_ /*42471*/;
assign _33185_ = _32646_ ^ _33187_ /*42474*/;
assign _33186_ = _33178_ & _33185_ /*42472*/;
assign _33095_ = _33178_ ^ _33185_ /*42473*/;
assign _33183_ = _33184_ | _33186_ /*42470*/;
assign _33192_ = ~D[7] /*42469*/;
assign _33189_ = _32647_ & _33192_ /*42465*/;
assign _33190_ = _32647_ ^ _33192_ /*42468*/;
assign _33191_ = _33183_ & _33190_ /*42466*/;
assign _33096_ = _33183_ ^ _33190_ /*42467*/;
assign _33188_ = _33189_ | _33191_ /*42464*/;
assign _33197_ = ~D[8] /*42463*/;
assign _33194_ = _32648_ & _33197_ /*42459*/;
assign _33195_ = _32648_ ^ _33197_ /*42462*/;
assign _33196_ = _33188_ & _33195_ /*42460*/;
assign _33097_ = _33188_ ^ _33195_ /*42461*/;
assign _33193_ = _33194_ | _33196_ /*42458*/;
assign _33202_ = ~D[9] /*42457*/;
assign _33199_ = _32649_ & _33202_ /*42453*/;
assign _33200_ = _32649_ ^ _33202_ /*42456*/;
assign _33201_ = _33193_ & _33200_ /*42454*/;
assign _33098_ = _33193_ ^ _33200_ /*42455*/;
assign _33198_ = _33199_ | _33201_ /*42452*/;
assign _33207_ = ~D[10] /*42451*/;
assign _33204_ = _32650_ & _33207_ /*42447*/;
assign _33205_ = _32650_ ^ _33207_ /*42450*/;
assign _33206_ = _33198_ & _33205_ /*42448*/;
assign _33099_ = _33198_ ^ _33205_ /*42449*/;
assign _33203_ = _33204_ | _33206_ /*42446*/;
assign _33212_ = ~D[11] /*42445*/;
assign _33209_ = _32651_ & _33212_ /*42441*/;
assign _33210_ = _32651_ ^ _33212_ /*42444*/;
assign _33211_ = _33203_ & _33210_ /*42442*/;
assign _33100_ = _33203_ ^ _33210_ /*42443*/;
assign _33208_ = _33209_ | _33211_ /*42440*/;
assign _33217_ = ~D[12] /*42439*/;
assign _33214_ = _32652_ & _33217_ /*42435*/;
assign _33215_ = _32652_ ^ _33217_ /*42438*/;
assign _33216_ = _33208_ & _33215_ /*42436*/;
assign _33101_ = _33208_ ^ _33215_ /*42437*/;
assign _33213_ = _33214_ | _33216_ /*42434*/;
assign _33222_ = ~D[13] /*42433*/;
assign _33219_ = _32653_ & _33222_ /*42429*/;
assign _33220_ = _32653_ ^ _33222_ /*42432*/;
assign _33221_ = _33213_ & _33220_ /*42430*/;
assign _33102_ = _33213_ ^ _33220_ /*42431*/;
assign _33218_ = _33219_ | _33221_ /*42428*/;
assign _33227_ = ~D[14] /*42427*/;
assign _33224_ = _32654_ & _33227_ /*42423*/;
assign _33225_ = _32654_ ^ _33227_ /*42426*/;
assign _33226_ = _33218_ & _33225_ /*42424*/;
assign _33103_ = _33218_ ^ _33225_ /*42425*/;
assign _33223_ = _33224_ | _33226_ /*42422*/;
assign _33232_ = ~D[15] /*42421*/;
assign _33229_ = _32655_ & _33232_ /*42417*/;
assign _33230_ = _32655_ ^ _33232_ /*42420*/;
assign _33231_ = _33223_ & _33230_ /*42418*/;
assign _33104_ = _33223_ ^ _33230_ /*42419*/;
assign _33228_ = _33229_ | _33231_ /*42416*/;
assign _33237_ = ~D[16] /*42415*/;
assign _33234_ = _32656_ & _33237_ /*42411*/;
assign _33235_ = _32656_ ^ _33237_ /*42414*/;
assign _33236_ = _33228_ & _33235_ /*42412*/;
assign _33105_ = _33228_ ^ _33235_ /*42413*/;
assign _33233_ = _33234_ | _33236_ /*42410*/;
assign _33242_ = ~D[17] /*42409*/;
assign _33239_ = _32657_ & _33242_ /*42405*/;
assign _33240_ = _32657_ ^ _33242_ /*42408*/;
assign _33241_ = _33233_ & _33240_ /*42406*/;
assign _33106_ = _33233_ ^ _33240_ /*42407*/;
assign _33238_ = _33239_ | _33241_ /*42404*/;
assign _33247_ = ~D[18] /*42403*/;
assign _33244_ = _32658_ & _33247_ /*42399*/;
assign _33245_ = _32658_ ^ _33247_ /*42402*/;
assign _33246_ = _33238_ & _33245_ /*42400*/;
assign _33107_ = _33238_ ^ _33245_ /*42401*/;
assign _33243_ = _33244_ | _33246_ /*42398*/;
assign _33252_ = ~D[19] /*42397*/;
assign _33249_ = _32659_ & _33252_ /*42393*/;
assign _33250_ = _32659_ ^ _33252_ /*42396*/;
assign _33251_ = _33243_ & _33250_ /*42394*/;
assign _33108_ = _33243_ ^ _33250_ /*42395*/;
assign _33248_ = _33249_ | _33251_ /*42392*/;
assign _33257_ = ~D[20] /*42391*/;
assign _33254_ = _32660_ & _33257_ /*42387*/;
assign _33255_ = _32660_ ^ _33257_ /*42390*/;
assign _33256_ = _33248_ & _33255_ /*42388*/;
assign _33109_ = _33248_ ^ _33255_ /*42389*/;
assign _33253_ = _33254_ | _33256_ /*42386*/;
assign _33262_ = ~D[21] /*42385*/;
assign _33259_ = _32661_ & _33262_ /*42381*/;
assign _33260_ = _32661_ ^ _33262_ /*42384*/;
assign _33261_ = _33253_ & _33260_ /*42382*/;
assign _33110_ = _33253_ ^ _33260_ /*42383*/;
assign _33258_ = _33259_ | _33261_ /*42380*/;
assign _33267_ = ~D[22] /*42379*/;
assign _33264_ = _32662_ & _33267_ /*42375*/;
assign _33265_ = _32662_ ^ _33267_ /*42378*/;
assign _33266_ = _33258_ & _33265_ /*42376*/;
assign _33111_ = _33258_ ^ _33265_ /*42377*/;
assign _33263_ = _33264_ | _33266_ /*42374*/;
assign _33272_ = ~D[23] /*42373*/;
assign _33269_ = _32663_ & _33272_ /*42369*/;
assign _33270_ = _32663_ ^ _33272_ /*42372*/;
assign _33271_ = _33263_ & _33270_ /*42370*/;
assign _33112_ = _33263_ ^ _33270_ /*42371*/;
assign _33268_ = _33269_ | _33271_ /*42368*/;
assign _33277_ = ~D[24] /*42367*/;
assign _33274_ = _32664_ & _33277_ /*42363*/;
assign _33275_ = _32664_ ^ _33277_ /*42366*/;
assign _33276_ = _33268_ & _33275_ /*42364*/;
assign _33113_ = _33268_ ^ _33275_ /*42365*/;
assign _33273_ = _33274_ | _33276_ /*42362*/;
assign _33282_ = ~D[25] /*42361*/;
assign _33279_ = _32665_ & _33282_ /*42357*/;
assign _33280_ = _32665_ ^ _33282_ /*42360*/;
assign _33281_ = _33273_ & _33280_ /*42358*/;
assign _33114_ = _33273_ ^ _33280_ /*42359*/;
assign _33278_ = _33279_ | _33281_ /*42356*/;
assign _33287_ = ~D[26] /*42355*/;
assign _33284_ = _32666_ & _33287_ /*42351*/;
assign _33285_ = _32666_ ^ _33287_ /*42354*/;
assign _33286_ = _33278_ & _33285_ /*42352*/;
assign _33115_ = _33278_ ^ _33285_ /*42353*/;
assign _33283_ = _33284_ | _33286_ /*42350*/;
assign _33292_ = ~D[27] /*42349*/;
assign _33289_ = _32667_ & _33292_ /*42345*/;
assign _33290_ = _32667_ ^ _33292_ /*42348*/;
assign _33291_ = _33283_ & _33290_ /*42346*/;
assign _33116_ = _33283_ ^ _33290_ /*42347*/;
assign _33288_ = _33289_ | _33291_ /*42344*/;
assign _33297_ = ~D[28] /*42343*/;
assign _33294_ = _32668_ & _33297_ /*42339*/;
assign _33295_ = _32668_ ^ _33297_ /*42342*/;
assign _33296_ = _33288_ & _33295_ /*42340*/;
assign _33117_ = _33288_ ^ _33295_ /*42341*/;
assign _33293_ = _33294_ | _33296_ /*42338*/;
assign _33302_ = ~D[29] /*42337*/;
assign _33299_ = _32669_ & _33302_ /*42333*/;
assign _33300_ = _32669_ ^ _33302_ /*42336*/;
assign _33301_ = _33293_ & _33300_ /*42334*/;
assign _33118_ = _33293_ ^ _33300_ /*42335*/;
assign _33298_ = _33299_ | _33301_ /*42332*/;
assign _33307_ = ~D[30] /*42331*/;
assign _33304_ = _32670_ & _33307_ /*42327*/;
assign _33305_ = _32670_ ^ _33307_ /*42330*/;
assign _33306_ = _33298_ & _33305_ /*42328*/;
assign _33119_ = _33298_ ^ _33305_ /*42329*/;
assign _33303_ = _33304_ | _33306_ /*42326*/;
assign _33312_ = ~D[31] /*42325*/;
assign _33309_ = _32671_ & _33312_ /*42321*/;
assign _33310_ = _32671_ ^ _33312_ /*42324*/;
assign _33311_ = _33303_ & _33310_ /*42322*/;
assign _33120_ = _33303_ ^ _33310_ /*42323*/;
assign _33308_ = _33309_ | _33311_ /*42320*/;
assign _33317_ = ~D[32] /*42319*/;
assign _33314_ = _32672_ & _33317_ /*42315*/;
assign _33315_ = _32672_ ^ _33317_ /*42318*/;
assign _33316_ = _33308_ & _33315_ /*42316*/;
assign _33121_ = _33308_ ^ _33315_ /*42317*/;
assign _33313_ = _33314_ | _33316_ /*42314*/;
assign _33322_ = ~D[33] /*42313*/;
assign _33319_ = _32673_ & _33322_ /*42309*/;
assign _33320_ = _32673_ ^ _33322_ /*42312*/;
assign _33321_ = _33313_ & _33320_ /*42310*/;
assign _33122_ = _33313_ ^ _33320_ /*42311*/;
assign _33318_ = _33319_ | _33321_ /*42308*/;
assign _33327_ = ~D[34] /*42307*/;
assign _33324_ = _32674_ & _33327_ /*42303*/;
assign _33325_ = _32674_ ^ _33327_ /*42306*/;
assign _33326_ = _33318_ & _33325_ /*42304*/;
assign _33123_ = _33318_ ^ _33325_ /*42305*/;
assign _33323_ = _33324_ | _33326_ /*42302*/;
assign _33332_ = ~D[35] /*42301*/;
assign _33329_ = _32675_ & _33332_ /*42297*/;
assign _33330_ = _32675_ ^ _33332_ /*42300*/;
assign _33331_ = _33323_ & _33330_ /*42298*/;
assign _33124_ = _33323_ ^ _33330_ /*42299*/;
assign _33328_ = _33329_ | _33331_ /*42296*/;
assign _33337_ = ~D[36] /*42295*/;
assign _33334_ = _32676_ & _33337_ /*42291*/;
assign _33335_ = _32676_ ^ _33337_ /*42294*/;
assign _33336_ = _33328_ & _33335_ /*42292*/;
assign _33125_ = _33328_ ^ _33335_ /*42293*/;
assign _33333_ = _33334_ | _33336_ /*42290*/;
assign _33342_ = ~D[37] /*42289*/;
assign _33339_ = _32677_ & _33342_ /*42285*/;
assign _33340_ = _32677_ ^ _33342_ /*42288*/;
assign _33341_ = _33333_ & _33340_ /*42286*/;
assign _33126_ = _33333_ ^ _33340_ /*42287*/;
assign _33338_ = _33339_ | _33341_ /*42284*/;
assign _33347_ = ~D[38] /*42283*/;
assign _33344_ = _32678_ & _33347_ /*42279*/;
assign _33345_ = _32678_ ^ _33347_ /*42282*/;
assign _33346_ = _33338_ & _33345_ /*42280*/;
assign _33127_ = _33338_ ^ _33345_ /*42281*/;
assign _33343_ = _33344_ | _33346_ /*42278*/;
assign _33352_ = ~D[39] /*42277*/;
assign _33349_ = _32679_ & _33352_ /*42273*/;
assign _33350_ = _32679_ ^ _33352_ /*42276*/;
assign _33351_ = _33343_ & _33350_ /*42274*/;
assign _33128_ = _33343_ ^ _33350_ /*42275*/;
assign _33348_ = _33349_ | _33351_ /*42272*/;
assign _33357_ = ~D[40] /*42271*/;
assign _33354_ = _32680_ & _33357_ /*42267*/;
assign _33355_ = _32680_ ^ _33357_ /*42270*/;
assign _33356_ = _33348_ & _33355_ /*42268*/;
assign _33129_ = _33348_ ^ _33355_ /*42269*/;
assign _33353_ = _33354_ | _33356_ /*42266*/;
assign _33362_ = ~D[41] /*42265*/;
assign _33359_ = _32681_ & _33362_ /*42261*/;
assign _33360_ = _32681_ ^ _33362_ /*42264*/;
assign _33361_ = _33353_ & _33360_ /*42262*/;
assign _33130_ = _33353_ ^ _33360_ /*42263*/;
assign _33358_ = _33359_ | _33361_ /*42260*/;
assign _33367_ = ~D[42] /*42259*/;
assign _33364_ = _32682_ & _33367_ /*42255*/;
assign _33365_ = _32682_ ^ _33367_ /*42258*/;
assign _33366_ = _33358_ & _33365_ /*42256*/;
assign _33131_ = _33358_ ^ _33365_ /*42257*/;
assign _33363_ = _33364_ | _33366_ /*42254*/;
assign _33372_ = ~D[43] /*42253*/;
assign _33369_ = _32683_ & _33372_ /*42249*/;
assign _33370_ = _32683_ ^ _33372_ /*42252*/;
assign _33371_ = _33363_ & _33370_ /*42250*/;
assign _33132_ = _33363_ ^ _33370_ /*42251*/;
assign _33368_ = _33369_ | _33371_ /*42248*/;
assign _33377_ = ~D[44] /*42247*/;
assign _33374_ = _32684_ & _33377_ /*42243*/;
assign _33375_ = _32684_ ^ _33377_ /*42246*/;
assign _33376_ = _33368_ & _33375_ /*42244*/;
assign _33133_ = _33368_ ^ _33375_ /*42245*/;
assign _33373_ = _33374_ | _33376_ /*42242*/;
assign _33382_ = ~D[45] /*42241*/;
assign _33379_ = _32685_ & _33382_ /*42237*/;
assign _33380_ = _32685_ ^ _33382_ /*42240*/;
assign _33381_ = _33373_ & _33380_ /*42238*/;
assign _33134_ = _33373_ ^ _33380_ /*42239*/;
assign _33378_ = _33379_ | _33381_ /*42236*/;
assign _33387_ = ~D[46] /*42235*/;
assign _33384_ = _32686_ & _33387_ /*42231*/;
assign _33385_ = _32686_ ^ _33387_ /*42234*/;
assign _33386_ = _33378_ & _33385_ /*42232*/;
assign _33135_ = _33378_ ^ _33385_ /*42233*/;
assign _33383_ = _33384_ | _33386_ /*42230*/;
assign _33392_ = ~D[47] /*42229*/;
assign _33389_ = _32687_ & _33392_ /*42225*/;
assign _33390_ = _32687_ ^ _33392_ /*42228*/;
assign _33391_ = _33383_ & _33390_ /*42226*/;
assign _33136_ = _33383_ ^ _33390_ /*42227*/;
assign _33388_ = _33389_ | _33391_ /*42224*/;
assign _33397_ = ~D[48] /*42223*/;
assign _33394_ = _32688_ & _33397_ /*42219*/;
assign _33395_ = _32688_ ^ _33397_ /*42222*/;
assign _33396_ = _33388_ & _33395_ /*42220*/;
assign _33137_ = _33388_ ^ _33395_ /*42221*/;
assign _33393_ = _33394_ | _33396_ /*42218*/;
assign _33402_ = ~D[49] /*42217*/;
assign _33399_ = _32689_ & _33402_ /*42213*/;
assign _33400_ = _32689_ ^ _33402_ /*42216*/;
assign _33401_ = _33393_ & _33400_ /*42214*/;
assign _33138_ = _33393_ ^ _33400_ /*42215*/;
assign _33398_ = _33399_ | _33401_ /*42212*/;
assign _33407_ = ~D[50] /*42211*/;
assign _33404_ = _32690_ & _33407_ /*42207*/;
assign _33405_ = _32690_ ^ _33407_ /*42210*/;
assign _33406_ = _33398_ & _33405_ /*42208*/;
assign _33139_ = _33398_ ^ _33405_ /*42209*/;
assign _33403_ = _33404_ | _33406_ /*42206*/;
assign _33412_ = ~D[51] /*42205*/;
assign _33409_ = _32691_ & _33412_ /*42201*/;
assign _33410_ = _32691_ ^ _33412_ /*42204*/;
assign _33411_ = _33403_ & _33410_ /*42202*/;
assign _33140_ = _33403_ ^ _33410_ /*42203*/;
assign _33408_ = _33409_ | _33411_ /*42200*/;
assign _33417_ = ~D[52] /*42199*/;
assign _33414_ = _32692_ & _33417_ /*42195*/;
assign _33415_ = _32692_ ^ _33417_ /*42198*/;
assign _33416_ = _33408_ & _33415_ /*42196*/;
assign _33141_ = _33408_ ^ _33415_ /*42197*/;
assign _33413_ = _33414_ | _33416_ /*42194*/;
assign _33422_ = ~D[53] /*42193*/;
assign _33419_ = _32693_ & _33422_ /*42189*/;
assign _33420_ = _32693_ ^ _33422_ /*42192*/;
assign _33421_ = _33413_ & _33420_ /*42190*/;
assign _33142_ = _33413_ ^ _33420_ /*42191*/;
assign _33418_ = _33419_ | _33421_ /*42188*/;
assign _33427_ = ~D[54] /*42187*/;
assign _33424_ = _32694_ & _33427_ /*42183*/;
assign _33425_ = _32694_ ^ _33427_ /*42186*/;
assign _33426_ = _33418_ & _33425_ /*42184*/;
assign _33143_ = _33418_ ^ _33425_ /*42185*/;
assign _33423_ = _33424_ | _33426_ /*42182*/;
assign _33432_ = ~D[55] /*42181*/;
assign _33429_ = _32695_ & _33432_ /*42177*/;
assign _33430_ = _32695_ ^ _33432_ /*42180*/;
assign _33431_ = _33423_ & _33430_ /*42178*/;
assign _33144_ = _33423_ ^ _33430_ /*42179*/;
assign _33428_ = _33429_ | _33431_ /*42176*/;
assign _33437_ = ~D[56] /*42175*/;
assign _33434_ = _32696_ & _33437_ /*42171*/;
assign _33435_ = _32696_ ^ _33437_ /*42174*/;
assign _33436_ = _33428_ & _33435_ /*42172*/;
assign _33145_ = _33428_ ^ _33435_ /*42173*/;
assign _33433_ = _33434_ | _33436_ /*42170*/;
assign _33442_ = ~D[57] /*42169*/;
assign _33439_ = _32697_ & _33442_ /*42165*/;
assign _33440_ = _32697_ ^ _33442_ /*42168*/;
assign _33441_ = _33433_ & _33440_ /*42166*/;
assign _33146_ = _33433_ ^ _33440_ /*42167*/;
assign _33438_ = _33439_ | _33441_ /*42164*/;
assign _33447_ = ~D[58] /*42163*/;
assign _33444_ = _32698_ & _33447_ /*42159*/;
assign _33445_ = _32698_ ^ _33447_ /*42162*/;
assign _33446_ = _33438_ & _33445_ /*42160*/;
assign _33147_ = _33438_ ^ _33445_ /*42161*/;
assign _33443_ = _33444_ | _33446_ /*42158*/;
assign _33452_ = ~D[59] /*42157*/;
assign _33449_ = _32699_ & _33452_ /*42153*/;
assign _33450_ = _32699_ ^ _33452_ /*42156*/;
assign _33451_ = _33443_ & _33450_ /*42154*/;
assign _33148_ = _33443_ ^ _33450_ /*42155*/;
assign _33448_ = _33449_ | _33451_ /*42152*/;
assign _33457_ = ~D[60] /*42151*/;
assign _33454_ = _32700_ & _33457_ /*42147*/;
assign _33455_ = _32700_ ^ _33457_ /*42150*/;
assign _33456_ = _33448_ & _33455_ /*42148*/;
assign _33149_ = _33448_ ^ _33455_ /*42149*/;
assign _33453_ = _33454_ | _33456_ /*42146*/;
assign _33462_ = ~D[61] /*42145*/;
assign _33459_ = _32701_ & _33462_ /*42141*/;
assign _33460_ = _32701_ ^ _33462_ /*42144*/;
assign _33461_ = _33453_ & _33460_ /*42142*/;
assign _33150_ = _33453_ ^ _33460_ /*42143*/;
assign _33458_ = _33459_ | _33461_ /*42140*/;
assign _33467_ = ~D[62] /*42139*/;
assign _33464_ = _32702_ & _33467_ /*42135*/;
assign _33465_ = _32702_ ^ _33467_ /*42138*/;
assign _33466_ = _33458_ & _33465_ /*42136*/;
assign _33151_ = _33458_ ^ _33465_ /*42137*/;
assign _33463_ = _33464_ | _33466_ /*42134*/;
assign _33468_ = _32703_ & oneWire /*42129*/;
assign _33469_ = _32703_ ^ oneWire /*42132*/;
assign _33470_ = _33463_ & _33469_ /*42130*/;
assign _33152_ = _33463_ ^ _33469_ /*42131*/;
assign Q[26] = _33468_ | _33470_ /*42128*/;
assign _33603_ = ~Q[26] /*41743*/;
assign _33602_ = _33603_ & D[0] /*41742*/;
assign _33605_ = _33089_ & _33602_ /*41737*/;
assign _33606_ = _33089_ ^ _33602_ /*41740*/;
assign _33607_ = zeroWire & _33606_ /*41738*/;
assign _33537_ = zeroWire ^ _33606_ /*41739*/;
assign _33604_ = _33605_ | _33607_ /*41736*/;
assign _33609_ = ~Q[26] /*41735*/;
assign _33608_ = _33609_ & D[1] /*41734*/;
assign _33611_ = _33090_ & _33608_ /*41729*/;
assign _33612_ = _33090_ ^ _33608_ /*41732*/;
assign _33613_ = _33604_ & _33612_ /*41730*/;
assign _33538_ = _33604_ ^ _33612_ /*41731*/;
assign _33610_ = _33611_ | _33613_ /*41728*/;
assign _33615_ = ~Q[26] /*41727*/;
assign _33614_ = _33615_ & D[2] /*41726*/;
assign _33617_ = _33091_ & _33614_ /*41721*/;
assign _33618_ = _33091_ ^ _33614_ /*41724*/;
assign _33619_ = _33610_ & _33618_ /*41722*/;
assign _33539_ = _33610_ ^ _33618_ /*41723*/;
assign _33616_ = _33617_ | _33619_ /*41720*/;
assign _33621_ = ~Q[26] /*41719*/;
assign _33620_ = _33621_ & D[3] /*41718*/;
assign _33623_ = _33092_ & _33620_ /*41713*/;
assign _33624_ = _33092_ ^ _33620_ /*41716*/;
assign _33625_ = _33616_ & _33624_ /*41714*/;
assign _33540_ = _33616_ ^ _33624_ /*41715*/;
assign _33622_ = _33623_ | _33625_ /*41712*/;
assign _33627_ = ~Q[26] /*41711*/;
assign _33626_ = _33627_ & D[4] /*41710*/;
assign _33629_ = _33093_ & _33626_ /*41705*/;
assign _33630_ = _33093_ ^ _33626_ /*41708*/;
assign _33631_ = _33622_ & _33630_ /*41706*/;
assign _33541_ = _33622_ ^ _33630_ /*41707*/;
assign _33628_ = _33629_ | _33631_ /*41704*/;
assign _33633_ = ~Q[26] /*41703*/;
assign _33632_ = _33633_ & D[5] /*41702*/;
assign _33635_ = _33094_ & _33632_ /*41697*/;
assign _33636_ = _33094_ ^ _33632_ /*41700*/;
assign _33637_ = _33628_ & _33636_ /*41698*/;
assign _33542_ = _33628_ ^ _33636_ /*41699*/;
assign _33634_ = _33635_ | _33637_ /*41696*/;
assign _33639_ = ~Q[26] /*41695*/;
assign _33638_ = _33639_ & D[6] /*41694*/;
assign _33641_ = _33095_ & _33638_ /*41689*/;
assign _33642_ = _33095_ ^ _33638_ /*41692*/;
assign _33643_ = _33634_ & _33642_ /*41690*/;
assign _33543_ = _33634_ ^ _33642_ /*41691*/;
assign _33640_ = _33641_ | _33643_ /*41688*/;
assign _33645_ = ~Q[26] /*41687*/;
assign _33644_ = _33645_ & D[7] /*41686*/;
assign _33647_ = _33096_ & _33644_ /*41681*/;
assign _33648_ = _33096_ ^ _33644_ /*41684*/;
assign _33649_ = _33640_ & _33648_ /*41682*/;
assign _33544_ = _33640_ ^ _33648_ /*41683*/;
assign _33646_ = _33647_ | _33649_ /*41680*/;
assign _33651_ = ~Q[26] /*41679*/;
assign _33650_ = _33651_ & D[8] /*41678*/;
assign _33653_ = _33097_ & _33650_ /*41673*/;
assign _33654_ = _33097_ ^ _33650_ /*41676*/;
assign _33655_ = _33646_ & _33654_ /*41674*/;
assign _33545_ = _33646_ ^ _33654_ /*41675*/;
assign _33652_ = _33653_ | _33655_ /*41672*/;
assign _33657_ = ~Q[26] /*41671*/;
assign _33656_ = _33657_ & D[9] /*41670*/;
assign _33659_ = _33098_ & _33656_ /*41665*/;
assign _33660_ = _33098_ ^ _33656_ /*41668*/;
assign _33661_ = _33652_ & _33660_ /*41666*/;
assign _33546_ = _33652_ ^ _33660_ /*41667*/;
assign _33658_ = _33659_ | _33661_ /*41664*/;
assign _33663_ = ~Q[26] /*41663*/;
assign _33662_ = _33663_ & D[10] /*41662*/;
assign _33665_ = _33099_ & _33662_ /*41657*/;
assign _33666_ = _33099_ ^ _33662_ /*41660*/;
assign _33667_ = _33658_ & _33666_ /*41658*/;
assign _33547_ = _33658_ ^ _33666_ /*41659*/;
assign _33664_ = _33665_ | _33667_ /*41656*/;
assign _33669_ = ~Q[26] /*41655*/;
assign _33668_ = _33669_ & D[11] /*41654*/;
assign _33671_ = _33100_ & _33668_ /*41649*/;
assign _33672_ = _33100_ ^ _33668_ /*41652*/;
assign _33673_ = _33664_ & _33672_ /*41650*/;
assign _33548_ = _33664_ ^ _33672_ /*41651*/;
assign _33670_ = _33671_ | _33673_ /*41648*/;
assign _33675_ = ~Q[26] /*41647*/;
assign _33674_ = _33675_ & D[12] /*41646*/;
assign _33677_ = _33101_ & _33674_ /*41641*/;
assign _33678_ = _33101_ ^ _33674_ /*41644*/;
assign _33679_ = _33670_ & _33678_ /*41642*/;
assign _33549_ = _33670_ ^ _33678_ /*41643*/;
assign _33676_ = _33677_ | _33679_ /*41640*/;
assign _33681_ = ~Q[26] /*41639*/;
assign _33680_ = _33681_ & D[13] /*41638*/;
assign _33683_ = _33102_ & _33680_ /*41633*/;
assign _33684_ = _33102_ ^ _33680_ /*41636*/;
assign _33685_ = _33676_ & _33684_ /*41634*/;
assign _33550_ = _33676_ ^ _33684_ /*41635*/;
assign _33682_ = _33683_ | _33685_ /*41632*/;
assign _33687_ = ~Q[26] /*41631*/;
assign _33686_ = _33687_ & D[14] /*41630*/;
assign _33689_ = _33103_ & _33686_ /*41625*/;
assign _33690_ = _33103_ ^ _33686_ /*41628*/;
assign _33691_ = _33682_ & _33690_ /*41626*/;
assign _33551_ = _33682_ ^ _33690_ /*41627*/;
assign _33688_ = _33689_ | _33691_ /*41624*/;
assign _33693_ = ~Q[26] /*41623*/;
assign _33692_ = _33693_ & D[15] /*41622*/;
assign _33695_ = _33104_ & _33692_ /*41617*/;
assign _33696_ = _33104_ ^ _33692_ /*41620*/;
assign _33697_ = _33688_ & _33696_ /*41618*/;
assign _33552_ = _33688_ ^ _33696_ /*41619*/;
assign _33694_ = _33695_ | _33697_ /*41616*/;
assign _33699_ = ~Q[26] /*41615*/;
assign _33698_ = _33699_ & D[16] /*41614*/;
assign _33701_ = _33105_ & _33698_ /*41609*/;
assign _33702_ = _33105_ ^ _33698_ /*41612*/;
assign _33703_ = _33694_ & _33702_ /*41610*/;
assign _33553_ = _33694_ ^ _33702_ /*41611*/;
assign _33700_ = _33701_ | _33703_ /*41608*/;
assign _33705_ = ~Q[26] /*41607*/;
assign _33704_ = _33705_ & D[17] /*41606*/;
assign _33707_ = _33106_ & _33704_ /*41601*/;
assign _33708_ = _33106_ ^ _33704_ /*41604*/;
assign _33709_ = _33700_ & _33708_ /*41602*/;
assign _33554_ = _33700_ ^ _33708_ /*41603*/;
assign _33706_ = _33707_ | _33709_ /*41600*/;
assign _33711_ = ~Q[26] /*41599*/;
assign _33710_ = _33711_ & D[18] /*41598*/;
assign _33713_ = _33107_ & _33710_ /*41593*/;
assign _33714_ = _33107_ ^ _33710_ /*41596*/;
assign _33715_ = _33706_ & _33714_ /*41594*/;
assign _33555_ = _33706_ ^ _33714_ /*41595*/;
assign _33712_ = _33713_ | _33715_ /*41592*/;
assign _33717_ = ~Q[26] /*41591*/;
assign _33716_ = _33717_ & D[19] /*41590*/;
assign _33719_ = _33108_ & _33716_ /*41585*/;
assign _33720_ = _33108_ ^ _33716_ /*41588*/;
assign _33721_ = _33712_ & _33720_ /*41586*/;
assign _33556_ = _33712_ ^ _33720_ /*41587*/;
assign _33718_ = _33719_ | _33721_ /*41584*/;
assign _33723_ = ~Q[26] /*41583*/;
assign _33722_ = _33723_ & D[20] /*41582*/;
assign _33725_ = _33109_ & _33722_ /*41577*/;
assign _33726_ = _33109_ ^ _33722_ /*41580*/;
assign _33727_ = _33718_ & _33726_ /*41578*/;
assign _33557_ = _33718_ ^ _33726_ /*41579*/;
assign _33724_ = _33725_ | _33727_ /*41576*/;
assign _33729_ = ~Q[26] /*41575*/;
assign _33728_ = _33729_ & D[21] /*41574*/;
assign _33731_ = _33110_ & _33728_ /*41569*/;
assign _33732_ = _33110_ ^ _33728_ /*41572*/;
assign _33733_ = _33724_ & _33732_ /*41570*/;
assign _33558_ = _33724_ ^ _33732_ /*41571*/;
assign _33730_ = _33731_ | _33733_ /*41568*/;
assign _33735_ = ~Q[26] /*41567*/;
assign _33734_ = _33735_ & D[22] /*41566*/;
assign _33737_ = _33111_ & _33734_ /*41561*/;
assign _33738_ = _33111_ ^ _33734_ /*41564*/;
assign _33739_ = _33730_ & _33738_ /*41562*/;
assign _33559_ = _33730_ ^ _33738_ /*41563*/;
assign _33736_ = _33737_ | _33739_ /*41560*/;
assign _33741_ = ~Q[26] /*41559*/;
assign _33740_ = _33741_ & D[23] /*41558*/;
assign _33743_ = _33112_ & _33740_ /*41553*/;
assign _33744_ = _33112_ ^ _33740_ /*41556*/;
assign _33745_ = _33736_ & _33744_ /*41554*/;
assign _33560_ = _33736_ ^ _33744_ /*41555*/;
assign _33742_ = _33743_ | _33745_ /*41552*/;
assign _33747_ = ~Q[26] /*41551*/;
assign _33746_ = _33747_ & D[24] /*41550*/;
assign _33749_ = _33113_ & _33746_ /*41545*/;
assign _33750_ = _33113_ ^ _33746_ /*41548*/;
assign _33751_ = _33742_ & _33750_ /*41546*/;
assign _33561_ = _33742_ ^ _33750_ /*41547*/;
assign _33748_ = _33749_ | _33751_ /*41544*/;
assign _33753_ = ~Q[26] /*41543*/;
assign _33752_ = _33753_ & D[25] /*41542*/;
assign _33755_ = _33114_ & _33752_ /*41537*/;
assign _33756_ = _33114_ ^ _33752_ /*41540*/;
assign _33757_ = _33748_ & _33756_ /*41538*/;
assign _33562_ = _33748_ ^ _33756_ /*41539*/;
assign _33754_ = _33755_ | _33757_ /*41536*/;
assign _33759_ = ~Q[26] /*41535*/;
assign _33758_ = _33759_ & D[26] /*41534*/;
assign _33761_ = _33115_ & _33758_ /*41529*/;
assign _33762_ = _33115_ ^ _33758_ /*41532*/;
assign _33763_ = _33754_ & _33762_ /*41530*/;
assign _33563_ = _33754_ ^ _33762_ /*41531*/;
assign _33760_ = _33761_ | _33763_ /*41528*/;
assign _33765_ = ~Q[26] /*41527*/;
assign _33764_ = _33765_ & D[27] /*41526*/;
assign _33767_ = _33116_ & _33764_ /*41521*/;
assign _33768_ = _33116_ ^ _33764_ /*41524*/;
assign _33769_ = _33760_ & _33768_ /*41522*/;
assign _33564_ = _33760_ ^ _33768_ /*41523*/;
assign _33766_ = _33767_ | _33769_ /*41520*/;
assign _33771_ = ~Q[26] /*41519*/;
assign _33770_ = _33771_ & D[28] /*41518*/;
assign _33773_ = _33117_ & _33770_ /*41513*/;
assign _33774_ = _33117_ ^ _33770_ /*41516*/;
assign _33775_ = _33766_ & _33774_ /*41514*/;
assign _33565_ = _33766_ ^ _33774_ /*41515*/;
assign _33772_ = _33773_ | _33775_ /*41512*/;
assign _33777_ = ~Q[26] /*41511*/;
assign _33776_ = _33777_ & D[29] /*41510*/;
assign _33779_ = _33118_ & _33776_ /*41505*/;
assign _33780_ = _33118_ ^ _33776_ /*41508*/;
assign _33781_ = _33772_ & _33780_ /*41506*/;
assign _33566_ = _33772_ ^ _33780_ /*41507*/;
assign _33778_ = _33779_ | _33781_ /*41504*/;
assign _33783_ = ~Q[26] /*41503*/;
assign _33782_ = _33783_ & D[30] /*41502*/;
assign _33785_ = _33119_ & _33782_ /*41497*/;
assign _33786_ = _33119_ ^ _33782_ /*41500*/;
assign _33787_ = _33778_ & _33786_ /*41498*/;
assign _33567_ = _33778_ ^ _33786_ /*41499*/;
assign _33784_ = _33785_ | _33787_ /*41496*/;
assign _33789_ = ~Q[26] /*41495*/;
assign _33788_ = _33789_ & D[31] /*41494*/;
assign _33791_ = _33120_ & _33788_ /*41489*/;
assign _33792_ = _33120_ ^ _33788_ /*41492*/;
assign _33793_ = _33784_ & _33792_ /*41490*/;
assign _33568_ = _33784_ ^ _33792_ /*41491*/;
assign _33790_ = _33791_ | _33793_ /*41488*/;
assign _33795_ = ~Q[26] /*41487*/;
assign _33794_ = _33795_ & D[32] /*41486*/;
assign _33797_ = _33121_ & _33794_ /*41481*/;
assign _33798_ = _33121_ ^ _33794_ /*41484*/;
assign _33799_ = _33790_ & _33798_ /*41482*/;
assign _33569_ = _33790_ ^ _33798_ /*41483*/;
assign _33796_ = _33797_ | _33799_ /*41480*/;
assign _33801_ = ~Q[26] /*41479*/;
assign _33800_ = _33801_ & D[33] /*41478*/;
assign _33803_ = _33122_ & _33800_ /*41473*/;
assign _33804_ = _33122_ ^ _33800_ /*41476*/;
assign _33805_ = _33796_ & _33804_ /*41474*/;
assign _33570_ = _33796_ ^ _33804_ /*41475*/;
assign _33802_ = _33803_ | _33805_ /*41472*/;
assign _33807_ = ~Q[26] /*41471*/;
assign _33806_ = _33807_ & D[34] /*41470*/;
assign _33809_ = _33123_ & _33806_ /*41465*/;
assign _33810_ = _33123_ ^ _33806_ /*41468*/;
assign _33811_ = _33802_ & _33810_ /*41466*/;
assign _33571_ = _33802_ ^ _33810_ /*41467*/;
assign _33808_ = _33809_ | _33811_ /*41464*/;
assign _33813_ = ~Q[26] /*41463*/;
assign _33812_ = _33813_ & D[35] /*41462*/;
assign _33815_ = _33124_ & _33812_ /*41457*/;
assign _33816_ = _33124_ ^ _33812_ /*41460*/;
assign _33817_ = _33808_ & _33816_ /*41458*/;
assign _33572_ = _33808_ ^ _33816_ /*41459*/;
assign _33814_ = _33815_ | _33817_ /*41456*/;
assign _33819_ = ~Q[26] /*41455*/;
assign _33818_ = _33819_ & D[36] /*41454*/;
assign _33821_ = _33125_ & _33818_ /*41449*/;
assign _33822_ = _33125_ ^ _33818_ /*41452*/;
assign _33823_ = _33814_ & _33822_ /*41450*/;
assign _33573_ = _33814_ ^ _33822_ /*41451*/;
assign _33820_ = _33821_ | _33823_ /*41448*/;
assign _33825_ = ~Q[26] /*41447*/;
assign _33824_ = _33825_ & D[37] /*41446*/;
assign _33827_ = _33126_ & _33824_ /*41441*/;
assign _33828_ = _33126_ ^ _33824_ /*41444*/;
assign _33829_ = _33820_ & _33828_ /*41442*/;
assign _33574_ = _33820_ ^ _33828_ /*41443*/;
assign _33826_ = _33827_ | _33829_ /*41440*/;
assign _33831_ = ~Q[26] /*41439*/;
assign _33830_ = _33831_ & D[38] /*41438*/;
assign _33833_ = _33127_ & _33830_ /*41433*/;
assign _33834_ = _33127_ ^ _33830_ /*41436*/;
assign _33835_ = _33826_ & _33834_ /*41434*/;
assign _33575_ = _33826_ ^ _33834_ /*41435*/;
assign _33832_ = _33833_ | _33835_ /*41432*/;
assign _33837_ = ~Q[26] /*41431*/;
assign _33836_ = _33837_ & D[39] /*41430*/;
assign _33839_ = _33128_ & _33836_ /*41425*/;
assign _33840_ = _33128_ ^ _33836_ /*41428*/;
assign _33841_ = _33832_ & _33840_ /*41426*/;
assign _33576_ = _33832_ ^ _33840_ /*41427*/;
assign _33838_ = _33839_ | _33841_ /*41424*/;
assign _33843_ = ~Q[26] /*41423*/;
assign _33842_ = _33843_ & D[40] /*41422*/;
assign _33845_ = _33129_ & _33842_ /*41417*/;
assign _33846_ = _33129_ ^ _33842_ /*41420*/;
assign _33847_ = _33838_ & _33846_ /*41418*/;
assign _33577_ = _33838_ ^ _33846_ /*41419*/;
assign _33844_ = _33845_ | _33847_ /*41416*/;
assign _33849_ = ~Q[26] /*41415*/;
assign _33848_ = _33849_ & D[41] /*41414*/;
assign _33851_ = _33130_ & _33848_ /*41409*/;
assign _33852_ = _33130_ ^ _33848_ /*41412*/;
assign _33853_ = _33844_ & _33852_ /*41410*/;
assign _33578_ = _33844_ ^ _33852_ /*41411*/;
assign _33850_ = _33851_ | _33853_ /*41408*/;
assign _33855_ = ~Q[26] /*41407*/;
assign _33854_ = _33855_ & D[42] /*41406*/;
assign _33857_ = _33131_ & _33854_ /*41401*/;
assign _33858_ = _33131_ ^ _33854_ /*41404*/;
assign _33859_ = _33850_ & _33858_ /*41402*/;
assign _33579_ = _33850_ ^ _33858_ /*41403*/;
assign _33856_ = _33857_ | _33859_ /*41400*/;
assign _33861_ = ~Q[26] /*41399*/;
assign _33860_ = _33861_ & D[43] /*41398*/;
assign _33863_ = _33132_ & _33860_ /*41393*/;
assign _33864_ = _33132_ ^ _33860_ /*41396*/;
assign _33865_ = _33856_ & _33864_ /*41394*/;
assign _33580_ = _33856_ ^ _33864_ /*41395*/;
assign _33862_ = _33863_ | _33865_ /*41392*/;
assign _33867_ = ~Q[26] /*41391*/;
assign _33866_ = _33867_ & D[44] /*41390*/;
assign _33869_ = _33133_ & _33866_ /*41385*/;
assign _33870_ = _33133_ ^ _33866_ /*41388*/;
assign _33871_ = _33862_ & _33870_ /*41386*/;
assign _33581_ = _33862_ ^ _33870_ /*41387*/;
assign _33868_ = _33869_ | _33871_ /*41384*/;
assign _33873_ = ~Q[26] /*41383*/;
assign _33872_ = _33873_ & D[45] /*41382*/;
assign _33875_ = _33134_ & _33872_ /*41377*/;
assign _33876_ = _33134_ ^ _33872_ /*41380*/;
assign _33877_ = _33868_ & _33876_ /*41378*/;
assign _33582_ = _33868_ ^ _33876_ /*41379*/;
assign _33874_ = _33875_ | _33877_ /*41376*/;
assign _33879_ = ~Q[26] /*41375*/;
assign _33878_ = _33879_ & D[46] /*41374*/;
assign _33881_ = _33135_ & _33878_ /*41369*/;
assign _33882_ = _33135_ ^ _33878_ /*41372*/;
assign _33883_ = _33874_ & _33882_ /*41370*/;
assign _33583_ = _33874_ ^ _33882_ /*41371*/;
assign _33880_ = _33881_ | _33883_ /*41368*/;
assign _33885_ = ~Q[26] /*41367*/;
assign _33884_ = _33885_ & D[47] /*41366*/;
assign _33887_ = _33136_ & _33884_ /*41361*/;
assign _33888_ = _33136_ ^ _33884_ /*41364*/;
assign _33889_ = _33880_ & _33888_ /*41362*/;
assign _33584_ = _33880_ ^ _33888_ /*41363*/;
assign _33886_ = _33887_ | _33889_ /*41360*/;
assign _33891_ = ~Q[26] /*41359*/;
assign _33890_ = _33891_ & D[48] /*41358*/;
assign _33893_ = _33137_ & _33890_ /*41353*/;
assign _33894_ = _33137_ ^ _33890_ /*41356*/;
assign _33895_ = _33886_ & _33894_ /*41354*/;
assign _33585_ = _33886_ ^ _33894_ /*41355*/;
assign _33892_ = _33893_ | _33895_ /*41352*/;
assign _33897_ = ~Q[26] /*41351*/;
assign _33896_ = _33897_ & D[49] /*41350*/;
assign _33899_ = _33138_ & _33896_ /*41345*/;
assign _33900_ = _33138_ ^ _33896_ /*41348*/;
assign _33901_ = _33892_ & _33900_ /*41346*/;
assign _33586_ = _33892_ ^ _33900_ /*41347*/;
assign _33898_ = _33899_ | _33901_ /*41344*/;
assign _33903_ = ~Q[26] /*41343*/;
assign _33902_ = _33903_ & D[50] /*41342*/;
assign _33905_ = _33139_ & _33902_ /*41337*/;
assign _33906_ = _33139_ ^ _33902_ /*41340*/;
assign _33907_ = _33898_ & _33906_ /*41338*/;
assign _33587_ = _33898_ ^ _33906_ /*41339*/;
assign _33904_ = _33905_ | _33907_ /*41336*/;
assign _33909_ = ~Q[26] /*41335*/;
assign _33908_ = _33909_ & D[51] /*41334*/;
assign _33911_ = _33140_ & _33908_ /*41329*/;
assign _33912_ = _33140_ ^ _33908_ /*41332*/;
assign _33913_ = _33904_ & _33912_ /*41330*/;
assign _33588_ = _33904_ ^ _33912_ /*41331*/;
assign _33910_ = _33911_ | _33913_ /*41328*/;
assign _33915_ = ~Q[26] /*41327*/;
assign _33914_ = _33915_ & D[52] /*41326*/;
assign _33917_ = _33141_ & _33914_ /*41321*/;
assign _33918_ = _33141_ ^ _33914_ /*41324*/;
assign _33919_ = _33910_ & _33918_ /*41322*/;
assign _33589_ = _33910_ ^ _33918_ /*41323*/;
assign _33916_ = _33917_ | _33919_ /*41320*/;
assign _33921_ = ~Q[26] /*41319*/;
assign _33920_ = _33921_ & D[53] /*41318*/;
assign _33923_ = _33142_ & _33920_ /*41313*/;
assign _33924_ = _33142_ ^ _33920_ /*41316*/;
assign _33925_ = _33916_ & _33924_ /*41314*/;
assign _33590_ = _33916_ ^ _33924_ /*41315*/;
assign _33922_ = _33923_ | _33925_ /*41312*/;
assign _33927_ = ~Q[26] /*41311*/;
assign _33926_ = _33927_ & D[54] /*41310*/;
assign _33929_ = _33143_ & _33926_ /*41305*/;
assign _33930_ = _33143_ ^ _33926_ /*41308*/;
assign _33931_ = _33922_ & _33930_ /*41306*/;
assign _33591_ = _33922_ ^ _33930_ /*41307*/;
assign _33928_ = _33929_ | _33931_ /*41304*/;
assign _33933_ = ~Q[26] /*41303*/;
assign _33932_ = _33933_ & D[55] /*41302*/;
assign _33935_ = _33144_ & _33932_ /*41297*/;
assign _33936_ = _33144_ ^ _33932_ /*41300*/;
assign _33937_ = _33928_ & _33936_ /*41298*/;
assign _33592_ = _33928_ ^ _33936_ /*41299*/;
assign _33934_ = _33935_ | _33937_ /*41296*/;
assign _33939_ = ~Q[26] /*41295*/;
assign _33938_ = _33939_ & D[56] /*41294*/;
assign _33941_ = _33145_ & _33938_ /*41289*/;
assign _33942_ = _33145_ ^ _33938_ /*41292*/;
assign _33943_ = _33934_ & _33942_ /*41290*/;
assign _33593_ = _33934_ ^ _33942_ /*41291*/;
assign _33940_ = _33941_ | _33943_ /*41288*/;
assign _33945_ = ~Q[26] /*41287*/;
assign _33944_ = _33945_ & D[57] /*41286*/;
assign _33947_ = _33146_ & _33944_ /*41281*/;
assign _33948_ = _33146_ ^ _33944_ /*41284*/;
assign _33949_ = _33940_ & _33948_ /*41282*/;
assign _33594_ = _33940_ ^ _33948_ /*41283*/;
assign _33946_ = _33947_ | _33949_ /*41280*/;
assign _33951_ = ~Q[26] /*41279*/;
assign _33950_ = _33951_ & D[58] /*41278*/;
assign _33953_ = _33147_ & _33950_ /*41273*/;
assign _33954_ = _33147_ ^ _33950_ /*41276*/;
assign _33955_ = _33946_ & _33954_ /*41274*/;
assign _33595_ = _33946_ ^ _33954_ /*41275*/;
assign _33952_ = _33953_ | _33955_ /*41272*/;
assign _33957_ = ~Q[26] /*41271*/;
assign _33956_ = _33957_ & D[59] /*41270*/;
assign _33959_ = _33148_ & _33956_ /*41265*/;
assign _33960_ = _33148_ ^ _33956_ /*41268*/;
assign _33961_ = _33952_ & _33960_ /*41266*/;
assign _33596_ = _33952_ ^ _33960_ /*41267*/;
assign _33958_ = _33959_ | _33961_ /*41264*/;
assign _33963_ = ~Q[26] /*41263*/;
assign _33962_ = _33963_ & D[60] /*41262*/;
assign _33965_ = _33149_ & _33962_ /*41257*/;
assign _33966_ = _33149_ ^ _33962_ /*41260*/;
assign _33967_ = _33958_ & _33966_ /*41258*/;
assign _33597_ = _33958_ ^ _33966_ /*41259*/;
assign _33964_ = _33965_ | _33967_ /*41256*/;
assign _33969_ = ~Q[26] /*41255*/;
assign _33968_ = _33969_ & D[61] /*41254*/;
assign _33971_ = _33150_ & _33968_ /*41249*/;
assign _33972_ = _33150_ ^ _33968_ /*41252*/;
assign _33973_ = _33964_ & _33972_ /*41250*/;
assign _33598_ = _33964_ ^ _33972_ /*41251*/;
assign _33970_ = _33971_ | _33973_ /*41248*/;
assign _33975_ = ~Q[26] /*41247*/;
assign _33974_ = _33975_ & D[62] /*41246*/;
assign _33977_ = _33151_ & _33974_ /*41241*/;
assign _33978_ = _33151_ ^ _33974_ /*41244*/;
assign _33979_ = _33970_ & _33978_ /*41242*/;
assign _33599_ = _33970_ ^ _33978_ /*41243*/;
assign _33976_ = _33977_ | _33979_ /*41240*/;
assign _33981_ = ~Q[26] /*41239*/;
assign _33980_ = _33981_ & zeroWire /*41238*/;
assign _33982_ = _33152_ ^ _33980_ /*41236*/;
assign _33600_ = _33982_ ^ _33976_ /*41235*/;
assign _34053_ = ~D[0] /*40981*/;
assign _34050_ = R_0[25] & _34053_ /*40977*/;
assign _34051_ = R_0[25] ^ _34053_ /*40980*/;
assign _34052_ = oneWire & _34051_ /*40978*/;
assign _33985_ = oneWire ^ _34051_ /*40979*/;
assign _34049_ = _34050_ | _34052_ /*40976*/;
assign _34058_ = ~D[1] /*40975*/;
assign _34055_ = _33537_ & _34058_ /*40971*/;
assign _34056_ = _33537_ ^ _34058_ /*40974*/;
assign _34057_ = _34049_ & _34056_ /*40972*/;
assign _33986_ = _34049_ ^ _34056_ /*40973*/;
assign _34054_ = _34055_ | _34057_ /*40970*/;
assign _34063_ = ~D[2] /*40969*/;
assign _34060_ = _33538_ & _34063_ /*40965*/;
assign _34061_ = _33538_ ^ _34063_ /*40968*/;
assign _34062_ = _34054_ & _34061_ /*40966*/;
assign _33987_ = _34054_ ^ _34061_ /*40967*/;
assign _34059_ = _34060_ | _34062_ /*40964*/;
assign _34068_ = ~D[3] /*40963*/;
assign _34065_ = _33539_ & _34068_ /*40959*/;
assign _34066_ = _33539_ ^ _34068_ /*40962*/;
assign _34067_ = _34059_ & _34066_ /*40960*/;
assign _33988_ = _34059_ ^ _34066_ /*40961*/;
assign _34064_ = _34065_ | _34067_ /*40958*/;
assign _34073_ = ~D[4] /*40957*/;
assign _34070_ = _33540_ & _34073_ /*40953*/;
assign _34071_ = _33540_ ^ _34073_ /*40956*/;
assign _34072_ = _34064_ & _34071_ /*40954*/;
assign _33989_ = _34064_ ^ _34071_ /*40955*/;
assign _34069_ = _34070_ | _34072_ /*40952*/;
assign _34078_ = ~D[5] /*40951*/;
assign _34075_ = _33541_ & _34078_ /*40947*/;
assign _34076_ = _33541_ ^ _34078_ /*40950*/;
assign _34077_ = _34069_ & _34076_ /*40948*/;
assign _33990_ = _34069_ ^ _34076_ /*40949*/;
assign _34074_ = _34075_ | _34077_ /*40946*/;
assign _34083_ = ~D[6] /*40945*/;
assign _34080_ = _33542_ & _34083_ /*40941*/;
assign _34081_ = _33542_ ^ _34083_ /*40944*/;
assign _34082_ = _34074_ & _34081_ /*40942*/;
assign _33991_ = _34074_ ^ _34081_ /*40943*/;
assign _34079_ = _34080_ | _34082_ /*40940*/;
assign _34088_ = ~D[7] /*40939*/;
assign _34085_ = _33543_ & _34088_ /*40935*/;
assign _34086_ = _33543_ ^ _34088_ /*40938*/;
assign _34087_ = _34079_ & _34086_ /*40936*/;
assign _33992_ = _34079_ ^ _34086_ /*40937*/;
assign _34084_ = _34085_ | _34087_ /*40934*/;
assign _34093_ = ~D[8] /*40933*/;
assign _34090_ = _33544_ & _34093_ /*40929*/;
assign _34091_ = _33544_ ^ _34093_ /*40932*/;
assign _34092_ = _34084_ & _34091_ /*40930*/;
assign _33993_ = _34084_ ^ _34091_ /*40931*/;
assign _34089_ = _34090_ | _34092_ /*40928*/;
assign _34098_ = ~D[9] /*40927*/;
assign _34095_ = _33545_ & _34098_ /*40923*/;
assign _34096_ = _33545_ ^ _34098_ /*40926*/;
assign _34097_ = _34089_ & _34096_ /*40924*/;
assign _33994_ = _34089_ ^ _34096_ /*40925*/;
assign _34094_ = _34095_ | _34097_ /*40922*/;
assign _34103_ = ~D[10] /*40921*/;
assign _34100_ = _33546_ & _34103_ /*40917*/;
assign _34101_ = _33546_ ^ _34103_ /*40920*/;
assign _34102_ = _34094_ & _34101_ /*40918*/;
assign _33995_ = _34094_ ^ _34101_ /*40919*/;
assign _34099_ = _34100_ | _34102_ /*40916*/;
assign _34108_ = ~D[11] /*40915*/;
assign _34105_ = _33547_ & _34108_ /*40911*/;
assign _34106_ = _33547_ ^ _34108_ /*40914*/;
assign _34107_ = _34099_ & _34106_ /*40912*/;
assign _33996_ = _34099_ ^ _34106_ /*40913*/;
assign _34104_ = _34105_ | _34107_ /*40910*/;
assign _34113_ = ~D[12] /*40909*/;
assign _34110_ = _33548_ & _34113_ /*40905*/;
assign _34111_ = _33548_ ^ _34113_ /*40908*/;
assign _34112_ = _34104_ & _34111_ /*40906*/;
assign _33997_ = _34104_ ^ _34111_ /*40907*/;
assign _34109_ = _34110_ | _34112_ /*40904*/;
assign _34118_ = ~D[13] /*40903*/;
assign _34115_ = _33549_ & _34118_ /*40899*/;
assign _34116_ = _33549_ ^ _34118_ /*40902*/;
assign _34117_ = _34109_ & _34116_ /*40900*/;
assign _33998_ = _34109_ ^ _34116_ /*40901*/;
assign _34114_ = _34115_ | _34117_ /*40898*/;
assign _34123_ = ~D[14] /*40897*/;
assign _34120_ = _33550_ & _34123_ /*40893*/;
assign _34121_ = _33550_ ^ _34123_ /*40896*/;
assign _34122_ = _34114_ & _34121_ /*40894*/;
assign _33999_ = _34114_ ^ _34121_ /*40895*/;
assign _34119_ = _34120_ | _34122_ /*40892*/;
assign _34128_ = ~D[15] /*40891*/;
assign _34125_ = _33551_ & _34128_ /*40887*/;
assign _34126_ = _33551_ ^ _34128_ /*40890*/;
assign _34127_ = _34119_ & _34126_ /*40888*/;
assign _34000_ = _34119_ ^ _34126_ /*40889*/;
assign _34124_ = _34125_ | _34127_ /*40886*/;
assign _34133_ = ~D[16] /*40885*/;
assign _34130_ = _33552_ & _34133_ /*40881*/;
assign _34131_ = _33552_ ^ _34133_ /*40884*/;
assign _34132_ = _34124_ & _34131_ /*40882*/;
assign _34001_ = _34124_ ^ _34131_ /*40883*/;
assign _34129_ = _34130_ | _34132_ /*40880*/;
assign _34138_ = ~D[17] /*40879*/;
assign _34135_ = _33553_ & _34138_ /*40875*/;
assign _34136_ = _33553_ ^ _34138_ /*40878*/;
assign _34137_ = _34129_ & _34136_ /*40876*/;
assign _34002_ = _34129_ ^ _34136_ /*40877*/;
assign _34134_ = _34135_ | _34137_ /*40874*/;
assign _34143_ = ~D[18] /*40873*/;
assign _34140_ = _33554_ & _34143_ /*40869*/;
assign _34141_ = _33554_ ^ _34143_ /*40872*/;
assign _34142_ = _34134_ & _34141_ /*40870*/;
assign _34003_ = _34134_ ^ _34141_ /*40871*/;
assign _34139_ = _34140_ | _34142_ /*40868*/;
assign _34148_ = ~D[19] /*40867*/;
assign _34145_ = _33555_ & _34148_ /*40863*/;
assign _34146_ = _33555_ ^ _34148_ /*40866*/;
assign _34147_ = _34139_ & _34146_ /*40864*/;
assign _34004_ = _34139_ ^ _34146_ /*40865*/;
assign _34144_ = _34145_ | _34147_ /*40862*/;
assign _34153_ = ~D[20] /*40861*/;
assign _34150_ = _33556_ & _34153_ /*40857*/;
assign _34151_ = _33556_ ^ _34153_ /*40860*/;
assign _34152_ = _34144_ & _34151_ /*40858*/;
assign _34005_ = _34144_ ^ _34151_ /*40859*/;
assign _34149_ = _34150_ | _34152_ /*40856*/;
assign _34158_ = ~D[21] /*40855*/;
assign _34155_ = _33557_ & _34158_ /*40851*/;
assign _34156_ = _33557_ ^ _34158_ /*40854*/;
assign _34157_ = _34149_ & _34156_ /*40852*/;
assign _34006_ = _34149_ ^ _34156_ /*40853*/;
assign _34154_ = _34155_ | _34157_ /*40850*/;
assign _34163_ = ~D[22] /*40849*/;
assign _34160_ = _33558_ & _34163_ /*40845*/;
assign _34161_ = _33558_ ^ _34163_ /*40848*/;
assign _34162_ = _34154_ & _34161_ /*40846*/;
assign _34007_ = _34154_ ^ _34161_ /*40847*/;
assign _34159_ = _34160_ | _34162_ /*40844*/;
assign _34168_ = ~D[23] /*40843*/;
assign _34165_ = _33559_ & _34168_ /*40839*/;
assign _34166_ = _33559_ ^ _34168_ /*40842*/;
assign _34167_ = _34159_ & _34166_ /*40840*/;
assign _34008_ = _34159_ ^ _34166_ /*40841*/;
assign _34164_ = _34165_ | _34167_ /*40838*/;
assign _34173_ = ~D[24] /*40837*/;
assign _34170_ = _33560_ & _34173_ /*40833*/;
assign _34171_ = _33560_ ^ _34173_ /*40836*/;
assign _34172_ = _34164_ & _34171_ /*40834*/;
assign _34009_ = _34164_ ^ _34171_ /*40835*/;
assign _34169_ = _34170_ | _34172_ /*40832*/;
assign _34178_ = ~D[25] /*40831*/;
assign _34175_ = _33561_ & _34178_ /*40827*/;
assign _34176_ = _33561_ ^ _34178_ /*40830*/;
assign _34177_ = _34169_ & _34176_ /*40828*/;
assign _34010_ = _34169_ ^ _34176_ /*40829*/;
assign _34174_ = _34175_ | _34177_ /*40826*/;
assign _34183_ = ~D[26] /*40825*/;
assign _34180_ = _33562_ & _34183_ /*40821*/;
assign _34181_ = _33562_ ^ _34183_ /*40824*/;
assign _34182_ = _34174_ & _34181_ /*40822*/;
assign _34011_ = _34174_ ^ _34181_ /*40823*/;
assign _34179_ = _34180_ | _34182_ /*40820*/;
assign _34188_ = ~D[27] /*40819*/;
assign _34185_ = _33563_ & _34188_ /*40815*/;
assign _34186_ = _33563_ ^ _34188_ /*40818*/;
assign _34187_ = _34179_ & _34186_ /*40816*/;
assign _34012_ = _34179_ ^ _34186_ /*40817*/;
assign _34184_ = _34185_ | _34187_ /*40814*/;
assign _34193_ = ~D[28] /*40813*/;
assign _34190_ = _33564_ & _34193_ /*40809*/;
assign _34191_ = _33564_ ^ _34193_ /*40812*/;
assign _34192_ = _34184_ & _34191_ /*40810*/;
assign _34013_ = _34184_ ^ _34191_ /*40811*/;
assign _34189_ = _34190_ | _34192_ /*40808*/;
assign _34198_ = ~D[29] /*40807*/;
assign _34195_ = _33565_ & _34198_ /*40803*/;
assign _34196_ = _33565_ ^ _34198_ /*40806*/;
assign _34197_ = _34189_ & _34196_ /*40804*/;
assign _34014_ = _34189_ ^ _34196_ /*40805*/;
assign _34194_ = _34195_ | _34197_ /*40802*/;
assign _34203_ = ~D[30] /*40801*/;
assign _34200_ = _33566_ & _34203_ /*40797*/;
assign _34201_ = _33566_ ^ _34203_ /*40800*/;
assign _34202_ = _34194_ & _34201_ /*40798*/;
assign _34015_ = _34194_ ^ _34201_ /*40799*/;
assign _34199_ = _34200_ | _34202_ /*40796*/;
assign _34208_ = ~D[31] /*40795*/;
assign _34205_ = _33567_ & _34208_ /*40791*/;
assign _34206_ = _33567_ ^ _34208_ /*40794*/;
assign _34207_ = _34199_ & _34206_ /*40792*/;
assign _34016_ = _34199_ ^ _34206_ /*40793*/;
assign _34204_ = _34205_ | _34207_ /*40790*/;
assign _34213_ = ~D[32] /*40789*/;
assign _34210_ = _33568_ & _34213_ /*40785*/;
assign _34211_ = _33568_ ^ _34213_ /*40788*/;
assign _34212_ = _34204_ & _34211_ /*40786*/;
assign _34017_ = _34204_ ^ _34211_ /*40787*/;
assign _34209_ = _34210_ | _34212_ /*40784*/;
assign _34218_ = ~D[33] /*40783*/;
assign _34215_ = _33569_ & _34218_ /*40779*/;
assign _34216_ = _33569_ ^ _34218_ /*40782*/;
assign _34217_ = _34209_ & _34216_ /*40780*/;
assign _34018_ = _34209_ ^ _34216_ /*40781*/;
assign _34214_ = _34215_ | _34217_ /*40778*/;
assign _34223_ = ~D[34] /*40777*/;
assign _34220_ = _33570_ & _34223_ /*40773*/;
assign _34221_ = _33570_ ^ _34223_ /*40776*/;
assign _34222_ = _34214_ & _34221_ /*40774*/;
assign _34019_ = _34214_ ^ _34221_ /*40775*/;
assign _34219_ = _34220_ | _34222_ /*40772*/;
assign _34228_ = ~D[35] /*40771*/;
assign _34225_ = _33571_ & _34228_ /*40767*/;
assign _34226_ = _33571_ ^ _34228_ /*40770*/;
assign _34227_ = _34219_ & _34226_ /*40768*/;
assign _34020_ = _34219_ ^ _34226_ /*40769*/;
assign _34224_ = _34225_ | _34227_ /*40766*/;
assign _34233_ = ~D[36] /*40765*/;
assign _34230_ = _33572_ & _34233_ /*40761*/;
assign _34231_ = _33572_ ^ _34233_ /*40764*/;
assign _34232_ = _34224_ & _34231_ /*40762*/;
assign _34021_ = _34224_ ^ _34231_ /*40763*/;
assign _34229_ = _34230_ | _34232_ /*40760*/;
assign _34238_ = ~D[37] /*40759*/;
assign _34235_ = _33573_ & _34238_ /*40755*/;
assign _34236_ = _33573_ ^ _34238_ /*40758*/;
assign _34237_ = _34229_ & _34236_ /*40756*/;
assign _34022_ = _34229_ ^ _34236_ /*40757*/;
assign _34234_ = _34235_ | _34237_ /*40754*/;
assign _34243_ = ~D[38] /*40753*/;
assign _34240_ = _33574_ & _34243_ /*40749*/;
assign _34241_ = _33574_ ^ _34243_ /*40752*/;
assign _34242_ = _34234_ & _34241_ /*40750*/;
assign _34023_ = _34234_ ^ _34241_ /*40751*/;
assign _34239_ = _34240_ | _34242_ /*40748*/;
assign _34248_ = ~D[39] /*40747*/;
assign _34245_ = _33575_ & _34248_ /*40743*/;
assign _34246_ = _33575_ ^ _34248_ /*40746*/;
assign _34247_ = _34239_ & _34246_ /*40744*/;
assign _34024_ = _34239_ ^ _34246_ /*40745*/;
assign _34244_ = _34245_ | _34247_ /*40742*/;
assign _34253_ = ~D[40] /*40741*/;
assign _34250_ = _33576_ & _34253_ /*40737*/;
assign _34251_ = _33576_ ^ _34253_ /*40740*/;
assign _34252_ = _34244_ & _34251_ /*40738*/;
assign _34025_ = _34244_ ^ _34251_ /*40739*/;
assign _34249_ = _34250_ | _34252_ /*40736*/;
assign _34258_ = ~D[41] /*40735*/;
assign _34255_ = _33577_ & _34258_ /*40731*/;
assign _34256_ = _33577_ ^ _34258_ /*40734*/;
assign _34257_ = _34249_ & _34256_ /*40732*/;
assign _34026_ = _34249_ ^ _34256_ /*40733*/;
assign _34254_ = _34255_ | _34257_ /*40730*/;
assign _34263_ = ~D[42] /*40729*/;
assign _34260_ = _33578_ & _34263_ /*40725*/;
assign _34261_ = _33578_ ^ _34263_ /*40728*/;
assign _34262_ = _34254_ & _34261_ /*40726*/;
assign _34027_ = _34254_ ^ _34261_ /*40727*/;
assign _34259_ = _34260_ | _34262_ /*40724*/;
assign _34268_ = ~D[43] /*40723*/;
assign _34265_ = _33579_ & _34268_ /*40719*/;
assign _34266_ = _33579_ ^ _34268_ /*40722*/;
assign _34267_ = _34259_ & _34266_ /*40720*/;
assign _34028_ = _34259_ ^ _34266_ /*40721*/;
assign _34264_ = _34265_ | _34267_ /*40718*/;
assign _34273_ = ~D[44] /*40717*/;
assign _34270_ = _33580_ & _34273_ /*40713*/;
assign _34271_ = _33580_ ^ _34273_ /*40716*/;
assign _34272_ = _34264_ & _34271_ /*40714*/;
assign _34029_ = _34264_ ^ _34271_ /*40715*/;
assign _34269_ = _34270_ | _34272_ /*40712*/;
assign _34278_ = ~D[45] /*40711*/;
assign _34275_ = _33581_ & _34278_ /*40707*/;
assign _34276_ = _33581_ ^ _34278_ /*40710*/;
assign _34277_ = _34269_ & _34276_ /*40708*/;
assign _34030_ = _34269_ ^ _34276_ /*40709*/;
assign _34274_ = _34275_ | _34277_ /*40706*/;
assign _34283_ = ~D[46] /*40705*/;
assign _34280_ = _33582_ & _34283_ /*40701*/;
assign _34281_ = _33582_ ^ _34283_ /*40704*/;
assign _34282_ = _34274_ & _34281_ /*40702*/;
assign _34031_ = _34274_ ^ _34281_ /*40703*/;
assign _34279_ = _34280_ | _34282_ /*40700*/;
assign _34288_ = ~D[47] /*40699*/;
assign _34285_ = _33583_ & _34288_ /*40695*/;
assign _34286_ = _33583_ ^ _34288_ /*40698*/;
assign _34287_ = _34279_ & _34286_ /*40696*/;
assign _34032_ = _34279_ ^ _34286_ /*40697*/;
assign _34284_ = _34285_ | _34287_ /*40694*/;
assign _34293_ = ~D[48] /*40693*/;
assign _34290_ = _33584_ & _34293_ /*40689*/;
assign _34291_ = _33584_ ^ _34293_ /*40692*/;
assign _34292_ = _34284_ & _34291_ /*40690*/;
assign _34033_ = _34284_ ^ _34291_ /*40691*/;
assign _34289_ = _34290_ | _34292_ /*40688*/;
assign _34298_ = ~D[49] /*40687*/;
assign _34295_ = _33585_ & _34298_ /*40683*/;
assign _34296_ = _33585_ ^ _34298_ /*40686*/;
assign _34297_ = _34289_ & _34296_ /*40684*/;
assign _34034_ = _34289_ ^ _34296_ /*40685*/;
assign _34294_ = _34295_ | _34297_ /*40682*/;
assign _34303_ = ~D[50] /*40681*/;
assign _34300_ = _33586_ & _34303_ /*40677*/;
assign _34301_ = _33586_ ^ _34303_ /*40680*/;
assign _34302_ = _34294_ & _34301_ /*40678*/;
assign _34035_ = _34294_ ^ _34301_ /*40679*/;
assign _34299_ = _34300_ | _34302_ /*40676*/;
assign _34308_ = ~D[51] /*40675*/;
assign _34305_ = _33587_ & _34308_ /*40671*/;
assign _34306_ = _33587_ ^ _34308_ /*40674*/;
assign _34307_ = _34299_ & _34306_ /*40672*/;
assign _34036_ = _34299_ ^ _34306_ /*40673*/;
assign _34304_ = _34305_ | _34307_ /*40670*/;
assign _34313_ = ~D[52] /*40669*/;
assign _34310_ = _33588_ & _34313_ /*40665*/;
assign _34311_ = _33588_ ^ _34313_ /*40668*/;
assign _34312_ = _34304_ & _34311_ /*40666*/;
assign _34037_ = _34304_ ^ _34311_ /*40667*/;
assign _34309_ = _34310_ | _34312_ /*40664*/;
assign _34318_ = ~D[53] /*40663*/;
assign _34315_ = _33589_ & _34318_ /*40659*/;
assign _34316_ = _33589_ ^ _34318_ /*40662*/;
assign _34317_ = _34309_ & _34316_ /*40660*/;
assign _34038_ = _34309_ ^ _34316_ /*40661*/;
assign _34314_ = _34315_ | _34317_ /*40658*/;
assign _34323_ = ~D[54] /*40657*/;
assign _34320_ = _33590_ & _34323_ /*40653*/;
assign _34321_ = _33590_ ^ _34323_ /*40656*/;
assign _34322_ = _34314_ & _34321_ /*40654*/;
assign _34039_ = _34314_ ^ _34321_ /*40655*/;
assign _34319_ = _34320_ | _34322_ /*40652*/;
assign _34328_ = ~D[55] /*40651*/;
assign _34325_ = _33591_ & _34328_ /*40647*/;
assign _34326_ = _33591_ ^ _34328_ /*40650*/;
assign _34327_ = _34319_ & _34326_ /*40648*/;
assign _34040_ = _34319_ ^ _34326_ /*40649*/;
assign _34324_ = _34325_ | _34327_ /*40646*/;
assign _34333_ = ~D[56] /*40645*/;
assign _34330_ = _33592_ & _34333_ /*40641*/;
assign _34331_ = _33592_ ^ _34333_ /*40644*/;
assign _34332_ = _34324_ & _34331_ /*40642*/;
assign _34041_ = _34324_ ^ _34331_ /*40643*/;
assign _34329_ = _34330_ | _34332_ /*40640*/;
assign _34338_ = ~D[57] /*40639*/;
assign _34335_ = _33593_ & _34338_ /*40635*/;
assign _34336_ = _33593_ ^ _34338_ /*40638*/;
assign _34337_ = _34329_ & _34336_ /*40636*/;
assign _34042_ = _34329_ ^ _34336_ /*40637*/;
assign _34334_ = _34335_ | _34337_ /*40634*/;
assign _34343_ = ~D[58] /*40633*/;
assign _34340_ = _33594_ & _34343_ /*40629*/;
assign _34341_ = _33594_ ^ _34343_ /*40632*/;
assign _34342_ = _34334_ & _34341_ /*40630*/;
assign _34043_ = _34334_ ^ _34341_ /*40631*/;
assign _34339_ = _34340_ | _34342_ /*40628*/;
assign _34348_ = ~D[59] /*40627*/;
assign _34345_ = _33595_ & _34348_ /*40623*/;
assign _34346_ = _33595_ ^ _34348_ /*40626*/;
assign _34347_ = _34339_ & _34346_ /*40624*/;
assign _34044_ = _34339_ ^ _34346_ /*40625*/;
assign _34344_ = _34345_ | _34347_ /*40622*/;
assign _34353_ = ~D[60] /*40621*/;
assign _34350_ = _33596_ & _34353_ /*40617*/;
assign _34351_ = _33596_ ^ _34353_ /*40620*/;
assign _34352_ = _34344_ & _34351_ /*40618*/;
assign _34045_ = _34344_ ^ _34351_ /*40619*/;
assign _34349_ = _34350_ | _34352_ /*40616*/;
assign _34358_ = ~D[61] /*40615*/;
assign _34355_ = _33597_ & _34358_ /*40611*/;
assign _34356_ = _33597_ ^ _34358_ /*40614*/;
assign _34357_ = _34349_ & _34356_ /*40612*/;
assign _34046_ = _34349_ ^ _34356_ /*40613*/;
assign _34354_ = _34355_ | _34357_ /*40610*/;
assign _34363_ = ~D[62] /*40609*/;
assign _34360_ = _33598_ & _34363_ /*40605*/;
assign _34361_ = _33598_ ^ _34363_ /*40608*/;
assign _34362_ = _34354_ & _34361_ /*40606*/;
assign _34047_ = _34354_ ^ _34361_ /*40607*/;
assign _34359_ = _34360_ | _34362_ /*40604*/;
assign _34364_ = _33599_ & oneWire /*40599*/;
assign _34365_ = _33599_ ^ oneWire /*40602*/;
assign _34366_ = _34359_ & _34365_ /*40600*/;
assign _34048_ = _34359_ ^ _34365_ /*40601*/;
assign Q[25] = _34364_ | _34366_ /*40598*/;
assign _34499_ = ~Q[25] /*40213*/;
assign _34498_ = _34499_ & D[0] /*40212*/;
assign _34501_ = _33985_ & _34498_ /*40207*/;
assign _34502_ = _33985_ ^ _34498_ /*40210*/;
assign _34503_ = zeroWire & _34502_ /*40208*/;
assign _34433_ = zeroWire ^ _34502_ /*40209*/;
assign _34500_ = _34501_ | _34503_ /*40206*/;
assign _34505_ = ~Q[25] /*40205*/;
assign _34504_ = _34505_ & D[1] /*40204*/;
assign _34507_ = _33986_ & _34504_ /*40199*/;
assign _34508_ = _33986_ ^ _34504_ /*40202*/;
assign _34509_ = _34500_ & _34508_ /*40200*/;
assign _34434_ = _34500_ ^ _34508_ /*40201*/;
assign _34506_ = _34507_ | _34509_ /*40198*/;
assign _34511_ = ~Q[25] /*40197*/;
assign _34510_ = _34511_ & D[2] /*40196*/;
assign _34513_ = _33987_ & _34510_ /*40191*/;
assign _34514_ = _33987_ ^ _34510_ /*40194*/;
assign _34515_ = _34506_ & _34514_ /*40192*/;
assign _34435_ = _34506_ ^ _34514_ /*40193*/;
assign _34512_ = _34513_ | _34515_ /*40190*/;
assign _34517_ = ~Q[25] /*40189*/;
assign _34516_ = _34517_ & D[3] /*40188*/;
assign _34519_ = _33988_ & _34516_ /*40183*/;
assign _34520_ = _33988_ ^ _34516_ /*40186*/;
assign _34521_ = _34512_ & _34520_ /*40184*/;
assign _34436_ = _34512_ ^ _34520_ /*40185*/;
assign _34518_ = _34519_ | _34521_ /*40182*/;
assign _34523_ = ~Q[25] /*40181*/;
assign _34522_ = _34523_ & D[4] /*40180*/;
assign _34525_ = _33989_ & _34522_ /*40175*/;
assign _34526_ = _33989_ ^ _34522_ /*40178*/;
assign _34527_ = _34518_ & _34526_ /*40176*/;
assign _34437_ = _34518_ ^ _34526_ /*40177*/;
assign _34524_ = _34525_ | _34527_ /*40174*/;
assign _34529_ = ~Q[25] /*40173*/;
assign _34528_ = _34529_ & D[5] /*40172*/;
assign _34531_ = _33990_ & _34528_ /*40167*/;
assign _34532_ = _33990_ ^ _34528_ /*40170*/;
assign _34533_ = _34524_ & _34532_ /*40168*/;
assign _34438_ = _34524_ ^ _34532_ /*40169*/;
assign _34530_ = _34531_ | _34533_ /*40166*/;
assign _34535_ = ~Q[25] /*40165*/;
assign _34534_ = _34535_ & D[6] /*40164*/;
assign _34537_ = _33991_ & _34534_ /*40159*/;
assign _34538_ = _33991_ ^ _34534_ /*40162*/;
assign _34539_ = _34530_ & _34538_ /*40160*/;
assign _34439_ = _34530_ ^ _34538_ /*40161*/;
assign _34536_ = _34537_ | _34539_ /*40158*/;
assign _34541_ = ~Q[25] /*40157*/;
assign _34540_ = _34541_ & D[7] /*40156*/;
assign _34543_ = _33992_ & _34540_ /*40151*/;
assign _34544_ = _33992_ ^ _34540_ /*40154*/;
assign _34545_ = _34536_ & _34544_ /*40152*/;
assign _34440_ = _34536_ ^ _34544_ /*40153*/;
assign _34542_ = _34543_ | _34545_ /*40150*/;
assign _34547_ = ~Q[25] /*40149*/;
assign _34546_ = _34547_ & D[8] /*40148*/;
assign _34549_ = _33993_ & _34546_ /*40143*/;
assign _34550_ = _33993_ ^ _34546_ /*40146*/;
assign _34551_ = _34542_ & _34550_ /*40144*/;
assign _34441_ = _34542_ ^ _34550_ /*40145*/;
assign _34548_ = _34549_ | _34551_ /*40142*/;
assign _34553_ = ~Q[25] /*40141*/;
assign _34552_ = _34553_ & D[9] /*40140*/;
assign _34555_ = _33994_ & _34552_ /*40135*/;
assign _34556_ = _33994_ ^ _34552_ /*40138*/;
assign _34557_ = _34548_ & _34556_ /*40136*/;
assign _34442_ = _34548_ ^ _34556_ /*40137*/;
assign _34554_ = _34555_ | _34557_ /*40134*/;
assign _34559_ = ~Q[25] /*40133*/;
assign _34558_ = _34559_ & D[10] /*40132*/;
assign _34561_ = _33995_ & _34558_ /*40127*/;
assign _34562_ = _33995_ ^ _34558_ /*40130*/;
assign _34563_ = _34554_ & _34562_ /*40128*/;
assign _34443_ = _34554_ ^ _34562_ /*40129*/;
assign _34560_ = _34561_ | _34563_ /*40126*/;
assign _34565_ = ~Q[25] /*40125*/;
assign _34564_ = _34565_ & D[11] /*40124*/;
assign _34567_ = _33996_ & _34564_ /*40119*/;
assign _34568_ = _33996_ ^ _34564_ /*40122*/;
assign _34569_ = _34560_ & _34568_ /*40120*/;
assign _34444_ = _34560_ ^ _34568_ /*40121*/;
assign _34566_ = _34567_ | _34569_ /*40118*/;
assign _34571_ = ~Q[25] /*40117*/;
assign _34570_ = _34571_ & D[12] /*40116*/;
assign _34573_ = _33997_ & _34570_ /*40111*/;
assign _34574_ = _33997_ ^ _34570_ /*40114*/;
assign _34575_ = _34566_ & _34574_ /*40112*/;
assign _34445_ = _34566_ ^ _34574_ /*40113*/;
assign _34572_ = _34573_ | _34575_ /*40110*/;
assign _34577_ = ~Q[25] /*40109*/;
assign _34576_ = _34577_ & D[13] /*40108*/;
assign _34579_ = _33998_ & _34576_ /*40103*/;
assign _34580_ = _33998_ ^ _34576_ /*40106*/;
assign _34581_ = _34572_ & _34580_ /*40104*/;
assign _34446_ = _34572_ ^ _34580_ /*40105*/;
assign _34578_ = _34579_ | _34581_ /*40102*/;
assign _34583_ = ~Q[25] /*40101*/;
assign _34582_ = _34583_ & D[14] /*40100*/;
assign _34585_ = _33999_ & _34582_ /*40095*/;
assign _34586_ = _33999_ ^ _34582_ /*40098*/;
assign _34587_ = _34578_ & _34586_ /*40096*/;
assign _34447_ = _34578_ ^ _34586_ /*40097*/;
assign _34584_ = _34585_ | _34587_ /*40094*/;
assign _34589_ = ~Q[25] /*40093*/;
assign _34588_ = _34589_ & D[15] /*40092*/;
assign _34591_ = _34000_ & _34588_ /*40087*/;
assign _34592_ = _34000_ ^ _34588_ /*40090*/;
assign _34593_ = _34584_ & _34592_ /*40088*/;
assign _34448_ = _34584_ ^ _34592_ /*40089*/;
assign _34590_ = _34591_ | _34593_ /*40086*/;
assign _34595_ = ~Q[25] /*40085*/;
assign _34594_ = _34595_ & D[16] /*40084*/;
assign _34597_ = _34001_ & _34594_ /*40079*/;
assign _34598_ = _34001_ ^ _34594_ /*40082*/;
assign _34599_ = _34590_ & _34598_ /*40080*/;
assign _34449_ = _34590_ ^ _34598_ /*40081*/;
assign _34596_ = _34597_ | _34599_ /*40078*/;
assign _34601_ = ~Q[25] /*40077*/;
assign _34600_ = _34601_ & D[17] /*40076*/;
assign _34603_ = _34002_ & _34600_ /*40071*/;
assign _34604_ = _34002_ ^ _34600_ /*40074*/;
assign _34605_ = _34596_ & _34604_ /*40072*/;
assign _34450_ = _34596_ ^ _34604_ /*40073*/;
assign _34602_ = _34603_ | _34605_ /*40070*/;
assign _34607_ = ~Q[25] /*40069*/;
assign _34606_ = _34607_ & D[18] /*40068*/;
assign _34609_ = _34003_ & _34606_ /*40063*/;
assign _34610_ = _34003_ ^ _34606_ /*40066*/;
assign _34611_ = _34602_ & _34610_ /*40064*/;
assign _34451_ = _34602_ ^ _34610_ /*40065*/;
assign _34608_ = _34609_ | _34611_ /*40062*/;
assign _34613_ = ~Q[25] /*40061*/;
assign _34612_ = _34613_ & D[19] /*40060*/;
assign _34615_ = _34004_ & _34612_ /*40055*/;
assign _34616_ = _34004_ ^ _34612_ /*40058*/;
assign _34617_ = _34608_ & _34616_ /*40056*/;
assign _34452_ = _34608_ ^ _34616_ /*40057*/;
assign _34614_ = _34615_ | _34617_ /*40054*/;
assign _34619_ = ~Q[25] /*40053*/;
assign _34618_ = _34619_ & D[20] /*40052*/;
assign _34621_ = _34005_ & _34618_ /*40047*/;
assign _34622_ = _34005_ ^ _34618_ /*40050*/;
assign _34623_ = _34614_ & _34622_ /*40048*/;
assign _34453_ = _34614_ ^ _34622_ /*40049*/;
assign _34620_ = _34621_ | _34623_ /*40046*/;
assign _34625_ = ~Q[25] /*40045*/;
assign _34624_ = _34625_ & D[21] /*40044*/;
assign _34627_ = _34006_ & _34624_ /*40039*/;
assign _34628_ = _34006_ ^ _34624_ /*40042*/;
assign _34629_ = _34620_ & _34628_ /*40040*/;
assign _34454_ = _34620_ ^ _34628_ /*40041*/;
assign _34626_ = _34627_ | _34629_ /*40038*/;
assign _34631_ = ~Q[25] /*40037*/;
assign _34630_ = _34631_ & D[22] /*40036*/;
assign _34633_ = _34007_ & _34630_ /*40031*/;
assign _34634_ = _34007_ ^ _34630_ /*40034*/;
assign _34635_ = _34626_ & _34634_ /*40032*/;
assign _34455_ = _34626_ ^ _34634_ /*40033*/;
assign _34632_ = _34633_ | _34635_ /*40030*/;
assign _34637_ = ~Q[25] /*40029*/;
assign _34636_ = _34637_ & D[23] /*40028*/;
assign _34639_ = _34008_ & _34636_ /*40023*/;
assign _34640_ = _34008_ ^ _34636_ /*40026*/;
assign _34641_ = _34632_ & _34640_ /*40024*/;
assign _34456_ = _34632_ ^ _34640_ /*40025*/;
assign _34638_ = _34639_ | _34641_ /*40022*/;
assign _34643_ = ~Q[25] /*40021*/;
assign _34642_ = _34643_ & D[24] /*40020*/;
assign _34645_ = _34009_ & _34642_ /*40015*/;
assign _34646_ = _34009_ ^ _34642_ /*40018*/;
assign _34647_ = _34638_ & _34646_ /*40016*/;
assign _34457_ = _34638_ ^ _34646_ /*40017*/;
assign _34644_ = _34645_ | _34647_ /*40014*/;
assign _34649_ = ~Q[25] /*40013*/;
assign _34648_ = _34649_ & D[25] /*40012*/;
assign _34651_ = _34010_ & _34648_ /*40007*/;
assign _34652_ = _34010_ ^ _34648_ /*40010*/;
assign _34653_ = _34644_ & _34652_ /*40008*/;
assign _34458_ = _34644_ ^ _34652_ /*40009*/;
assign _34650_ = _34651_ | _34653_ /*40006*/;
assign _34655_ = ~Q[25] /*40005*/;
assign _34654_ = _34655_ & D[26] /*40004*/;
assign _34657_ = _34011_ & _34654_ /*39999*/;
assign _34658_ = _34011_ ^ _34654_ /*40002*/;
assign _34659_ = _34650_ & _34658_ /*40000*/;
assign _34459_ = _34650_ ^ _34658_ /*40001*/;
assign _34656_ = _34657_ | _34659_ /*39998*/;
assign _34661_ = ~Q[25] /*39997*/;
assign _34660_ = _34661_ & D[27] /*39996*/;
assign _34663_ = _34012_ & _34660_ /*39991*/;
assign _34664_ = _34012_ ^ _34660_ /*39994*/;
assign _34665_ = _34656_ & _34664_ /*39992*/;
assign _34460_ = _34656_ ^ _34664_ /*39993*/;
assign _34662_ = _34663_ | _34665_ /*39990*/;
assign _34667_ = ~Q[25] /*39989*/;
assign _34666_ = _34667_ & D[28] /*39988*/;
assign _34669_ = _34013_ & _34666_ /*39983*/;
assign _34670_ = _34013_ ^ _34666_ /*39986*/;
assign _34671_ = _34662_ & _34670_ /*39984*/;
assign _34461_ = _34662_ ^ _34670_ /*39985*/;
assign _34668_ = _34669_ | _34671_ /*39982*/;
assign _34673_ = ~Q[25] /*39981*/;
assign _34672_ = _34673_ & D[29] /*39980*/;
assign _34675_ = _34014_ & _34672_ /*39975*/;
assign _34676_ = _34014_ ^ _34672_ /*39978*/;
assign _34677_ = _34668_ & _34676_ /*39976*/;
assign _34462_ = _34668_ ^ _34676_ /*39977*/;
assign _34674_ = _34675_ | _34677_ /*39974*/;
assign _34679_ = ~Q[25] /*39973*/;
assign _34678_ = _34679_ & D[30] /*39972*/;
assign _34681_ = _34015_ & _34678_ /*39967*/;
assign _34682_ = _34015_ ^ _34678_ /*39970*/;
assign _34683_ = _34674_ & _34682_ /*39968*/;
assign _34463_ = _34674_ ^ _34682_ /*39969*/;
assign _34680_ = _34681_ | _34683_ /*39966*/;
assign _34685_ = ~Q[25] /*39965*/;
assign _34684_ = _34685_ & D[31] /*39964*/;
assign _34687_ = _34016_ & _34684_ /*39959*/;
assign _34688_ = _34016_ ^ _34684_ /*39962*/;
assign _34689_ = _34680_ & _34688_ /*39960*/;
assign _34464_ = _34680_ ^ _34688_ /*39961*/;
assign _34686_ = _34687_ | _34689_ /*39958*/;
assign _34691_ = ~Q[25] /*39957*/;
assign _34690_ = _34691_ & D[32] /*39956*/;
assign _34693_ = _34017_ & _34690_ /*39951*/;
assign _34694_ = _34017_ ^ _34690_ /*39954*/;
assign _34695_ = _34686_ & _34694_ /*39952*/;
assign _34465_ = _34686_ ^ _34694_ /*39953*/;
assign _34692_ = _34693_ | _34695_ /*39950*/;
assign _34697_ = ~Q[25] /*39949*/;
assign _34696_ = _34697_ & D[33] /*39948*/;
assign _34699_ = _34018_ & _34696_ /*39943*/;
assign _34700_ = _34018_ ^ _34696_ /*39946*/;
assign _34701_ = _34692_ & _34700_ /*39944*/;
assign _34466_ = _34692_ ^ _34700_ /*39945*/;
assign _34698_ = _34699_ | _34701_ /*39942*/;
assign _34703_ = ~Q[25] /*39941*/;
assign _34702_ = _34703_ & D[34] /*39940*/;
assign _34705_ = _34019_ & _34702_ /*39935*/;
assign _34706_ = _34019_ ^ _34702_ /*39938*/;
assign _34707_ = _34698_ & _34706_ /*39936*/;
assign _34467_ = _34698_ ^ _34706_ /*39937*/;
assign _34704_ = _34705_ | _34707_ /*39934*/;
assign _34709_ = ~Q[25] /*39933*/;
assign _34708_ = _34709_ & D[35] /*39932*/;
assign _34711_ = _34020_ & _34708_ /*39927*/;
assign _34712_ = _34020_ ^ _34708_ /*39930*/;
assign _34713_ = _34704_ & _34712_ /*39928*/;
assign _34468_ = _34704_ ^ _34712_ /*39929*/;
assign _34710_ = _34711_ | _34713_ /*39926*/;
assign _34715_ = ~Q[25] /*39925*/;
assign _34714_ = _34715_ & D[36] /*39924*/;
assign _34717_ = _34021_ & _34714_ /*39919*/;
assign _34718_ = _34021_ ^ _34714_ /*39922*/;
assign _34719_ = _34710_ & _34718_ /*39920*/;
assign _34469_ = _34710_ ^ _34718_ /*39921*/;
assign _34716_ = _34717_ | _34719_ /*39918*/;
assign _34721_ = ~Q[25] /*39917*/;
assign _34720_ = _34721_ & D[37] /*39916*/;
assign _34723_ = _34022_ & _34720_ /*39911*/;
assign _34724_ = _34022_ ^ _34720_ /*39914*/;
assign _34725_ = _34716_ & _34724_ /*39912*/;
assign _34470_ = _34716_ ^ _34724_ /*39913*/;
assign _34722_ = _34723_ | _34725_ /*39910*/;
assign _34727_ = ~Q[25] /*39909*/;
assign _34726_ = _34727_ & D[38] /*39908*/;
assign _34729_ = _34023_ & _34726_ /*39903*/;
assign _34730_ = _34023_ ^ _34726_ /*39906*/;
assign _34731_ = _34722_ & _34730_ /*39904*/;
assign _34471_ = _34722_ ^ _34730_ /*39905*/;
assign _34728_ = _34729_ | _34731_ /*39902*/;
assign _34733_ = ~Q[25] /*39901*/;
assign _34732_ = _34733_ & D[39] /*39900*/;
assign _34735_ = _34024_ & _34732_ /*39895*/;
assign _34736_ = _34024_ ^ _34732_ /*39898*/;
assign _34737_ = _34728_ & _34736_ /*39896*/;
assign _34472_ = _34728_ ^ _34736_ /*39897*/;
assign _34734_ = _34735_ | _34737_ /*39894*/;
assign _34739_ = ~Q[25] /*39893*/;
assign _34738_ = _34739_ & D[40] /*39892*/;
assign _34741_ = _34025_ & _34738_ /*39887*/;
assign _34742_ = _34025_ ^ _34738_ /*39890*/;
assign _34743_ = _34734_ & _34742_ /*39888*/;
assign _34473_ = _34734_ ^ _34742_ /*39889*/;
assign _34740_ = _34741_ | _34743_ /*39886*/;
assign _34745_ = ~Q[25] /*39885*/;
assign _34744_ = _34745_ & D[41] /*39884*/;
assign _34747_ = _34026_ & _34744_ /*39879*/;
assign _34748_ = _34026_ ^ _34744_ /*39882*/;
assign _34749_ = _34740_ & _34748_ /*39880*/;
assign _34474_ = _34740_ ^ _34748_ /*39881*/;
assign _34746_ = _34747_ | _34749_ /*39878*/;
assign _34751_ = ~Q[25] /*39877*/;
assign _34750_ = _34751_ & D[42] /*39876*/;
assign _34753_ = _34027_ & _34750_ /*39871*/;
assign _34754_ = _34027_ ^ _34750_ /*39874*/;
assign _34755_ = _34746_ & _34754_ /*39872*/;
assign _34475_ = _34746_ ^ _34754_ /*39873*/;
assign _34752_ = _34753_ | _34755_ /*39870*/;
assign _34757_ = ~Q[25] /*39869*/;
assign _34756_ = _34757_ & D[43] /*39868*/;
assign _34759_ = _34028_ & _34756_ /*39863*/;
assign _34760_ = _34028_ ^ _34756_ /*39866*/;
assign _34761_ = _34752_ & _34760_ /*39864*/;
assign _34476_ = _34752_ ^ _34760_ /*39865*/;
assign _34758_ = _34759_ | _34761_ /*39862*/;
assign _34763_ = ~Q[25] /*39861*/;
assign _34762_ = _34763_ & D[44] /*39860*/;
assign _34765_ = _34029_ & _34762_ /*39855*/;
assign _34766_ = _34029_ ^ _34762_ /*39858*/;
assign _34767_ = _34758_ & _34766_ /*39856*/;
assign _34477_ = _34758_ ^ _34766_ /*39857*/;
assign _34764_ = _34765_ | _34767_ /*39854*/;
assign _34769_ = ~Q[25] /*39853*/;
assign _34768_ = _34769_ & D[45] /*39852*/;
assign _34771_ = _34030_ & _34768_ /*39847*/;
assign _34772_ = _34030_ ^ _34768_ /*39850*/;
assign _34773_ = _34764_ & _34772_ /*39848*/;
assign _34478_ = _34764_ ^ _34772_ /*39849*/;
assign _34770_ = _34771_ | _34773_ /*39846*/;
assign _34775_ = ~Q[25] /*39845*/;
assign _34774_ = _34775_ & D[46] /*39844*/;
assign _34777_ = _34031_ & _34774_ /*39839*/;
assign _34778_ = _34031_ ^ _34774_ /*39842*/;
assign _34779_ = _34770_ & _34778_ /*39840*/;
assign _34479_ = _34770_ ^ _34778_ /*39841*/;
assign _34776_ = _34777_ | _34779_ /*39838*/;
assign _34781_ = ~Q[25] /*39837*/;
assign _34780_ = _34781_ & D[47] /*39836*/;
assign _34783_ = _34032_ & _34780_ /*39831*/;
assign _34784_ = _34032_ ^ _34780_ /*39834*/;
assign _34785_ = _34776_ & _34784_ /*39832*/;
assign _34480_ = _34776_ ^ _34784_ /*39833*/;
assign _34782_ = _34783_ | _34785_ /*39830*/;
assign _34787_ = ~Q[25] /*39829*/;
assign _34786_ = _34787_ & D[48] /*39828*/;
assign _34789_ = _34033_ & _34786_ /*39823*/;
assign _34790_ = _34033_ ^ _34786_ /*39826*/;
assign _34791_ = _34782_ & _34790_ /*39824*/;
assign _34481_ = _34782_ ^ _34790_ /*39825*/;
assign _34788_ = _34789_ | _34791_ /*39822*/;
assign _34793_ = ~Q[25] /*39821*/;
assign _34792_ = _34793_ & D[49] /*39820*/;
assign _34795_ = _34034_ & _34792_ /*39815*/;
assign _34796_ = _34034_ ^ _34792_ /*39818*/;
assign _34797_ = _34788_ & _34796_ /*39816*/;
assign _34482_ = _34788_ ^ _34796_ /*39817*/;
assign _34794_ = _34795_ | _34797_ /*39814*/;
assign _34799_ = ~Q[25] /*39813*/;
assign _34798_ = _34799_ & D[50] /*39812*/;
assign _34801_ = _34035_ & _34798_ /*39807*/;
assign _34802_ = _34035_ ^ _34798_ /*39810*/;
assign _34803_ = _34794_ & _34802_ /*39808*/;
assign _34483_ = _34794_ ^ _34802_ /*39809*/;
assign _34800_ = _34801_ | _34803_ /*39806*/;
assign _34805_ = ~Q[25] /*39805*/;
assign _34804_ = _34805_ & D[51] /*39804*/;
assign _34807_ = _34036_ & _34804_ /*39799*/;
assign _34808_ = _34036_ ^ _34804_ /*39802*/;
assign _34809_ = _34800_ & _34808_ /*39800*/;
assign _34484_ = _34800_ ^ _34808_ /*39801*/;
assign _34806_ = _34807_ | _34809_ /*39798*/;
assign _34811_ = ~Q[25] /*39797*/;
assign _34810_ = _34811_ & D[52] /*39796*/;
assign _34813_ = _34037_ & _34810_ /*39791*/;
assign _34814_ = _34037_ ^ _34810_ /*39794*/;
assign _34815_ = _34806_ & _34814_ /*39792*/;
assign _34485_ = _34806_ ^ _34814_ /*39793*/;
assign _34812_ = _34813_ | _34815_ /*39790*/;
assign _34817_ = ~Q[25] /*39789*/;
assign _34816_ = _34817_ & D[53] /*39788*/;
assign _34819_ = _34038_ & _34816_ /*39783*/;
assign _34820_ = _34038_ ^ _34816_ /*39786*/;
assign _34821_ = _34812_ & _34820_ /*39784*/;
assign _34486_ = _34812_ ^ _34820_ /*39785*/;
assign _34818_ = _34819_ | _34821_ /*39782*/;
assign _34823_ = ~Q[25] /*39781*/;
assign _34822_ = _34823_ & D[54] /*39780*/;
assign _34825_ = _34039_ & _34822_ /*39775*/;
assign _34826_ = _34039_ ^ _34822_ /*39778*/;
assign _34827_ = _34818_ & _34826_ /*39776*/;
assign _34487_ = _34818_ ^ _34826_ /*39777*/;
assign _34824_ = _34825_ | _34827_ /*39774*/;
assign _34829_ = ~Q[25] /*39773*/;
assign _34828_ = _34829_ & D[55] /*39772*/;
assign _34831_ = _34040_ & _34828_ /*39767*/;
assign _34832_ = _34040_ ^ _34828_ /*39770*/;
assign _34833_ = _34824_ & _34832_ /*39768*/;
assign _34488_ = _34824_ ^ _34832_ /*39769*/;
assign _34830_ = _34831_ | _34833_ /*39766*/;
assign _34835_ = ~Q[25] /*39765*/;
assign _34834_ = _34835_ & D[56] /*39764*/;
assign _34837_ = _34041_ & _34834_ /*39759*/;
assign _34838_ = _34041_ ^ _34834_ /*39762*/;
assign _34839_ = _34830_ & _34838_ /*39760*/;
assign _34489_ = _34830_ ^ _34838_ /*39761*/;
assign _34836_ = _34837_ | _34839_ /*39758*/;
assign _34841_ = ~Q[25] /*39757*/;
assign _34840_ = _34841_ & D[57] /*39756*/;
assign _34843_ = _34042_ & _34840_ /*39751*/;
assign _34844_ = _34042_ ^ _34840_ /*39754*/;
assign _34845_ = _34836_ & _34844_ /*39752*/;
assign _34490_ = _34836_ ^ _34844_ /*39753*/;
assign _34842_ = _34843_ | _34845_ /*39750*/;
assign _34847_ = ~Q[25] /*39749*/;
assign _34846_ = _34847_ & D[58] /*39748*/;
assign _34849_ = _34043_ & _34846_ /*39743*/;
assign _34850_ = _34043_ ^ _34846_ /*39746*/;
assign _34851_ = _34842_ & _34850_ /*39744*/;
assign _34491_ = _34842_ ^ _34850_ /*39745*/;
assign _34848_ = _34849_ | _34851_ /*39742*/;
assign _34853_ = ~Q[25] /*39741*/;
assign _34852_ = _34853_ & D[59] /*39740*/;
assign _34855_ = _34044_ & _34852_ /*39735*/;
assign _34856_ = _34044_ ^ _34852_ /*39738*/;
assign _34857_ = _34848_ & _34856_ /*39736*/;
assign _34492_ = _34848_ ^ _34856_ /*39737*/;
assign _34854_ = _34855_ | _34857_ /*39734*/;
assign _34859_ = ~Q[25] /*39733*/;
assign _34858_ = _34859_ & D[60] /*39732*/;
assign _34861_ = _34045_ & _34858_ /*39727*/;
assign _34862_ = _34045_ ^ _34858_ /*39730*/;
assign _34863_ = _34854_ & _34862_ /*39728*/;
assign _34493_ = _34854_ ^ _34862_ /*39729*/;
assign _34860_ = _34861_ | _34863_ /*39726*/;
assign _34865_ = ~Q[25] /*39725*/;
assign _34864_ = _34865_ & D[61] /*39724*/;
assign _34867_ = _34046_ & _34864_ /*39719*/;
assign _34868_ = _34046_ ^ _34864_ /*39722*/;
assign _34869_ = _34860_ & _34868_ /*39720*/;
assign _34494_ = _34860_ ^ _34868_ /*39721*/;
assign _34866_ = _34867_ | _34869_ /*39718*/;
assign _34871_ = ~Q[25] /*39717*/;
assign _34870_ = _34871_ & D[62] /*39716*/;
assign _34873_ = _34047_ & _34870_ /*39711*/;
assign _34874_ = _34047_ ^ _34870_ /*39714*/;
assign _34875_ = _34866_ & _34874_ /*39712*/;
assign _34495_ = _34866_ ^ _34874_ /*39713*/;
assign _34872_ = _34873_ | _34875_ /*39710*/;
assign _34877_ = ~Q[25] /*39709*/;
assign _34876_ = _34877_ & zeroWire /*39708*/;
assign _34878_ = _34048_ ^ _34876_ /*39706*/;
assign _34496_ = _34878_ ^ _34872_ /*39705*/;
assign _34949_ = ~D[0] /*39451*/;
assign _34946_ = R_0[24] & _34949_ /*39447*/;
assign _34947_ = R_0[24] ^ _34949_ /*39450*/;
assign _34948_ = oneWire & _34947_ /*39448*/;
assign _34881_ = oneWire ^ _34947_ /*39449*/;
assign _34945_ = _34946_ | _34948_ /*39446*/;
assign _34954_ = ~D[1] /*39445*/;
assign _34951_ = _34433_ & _34954_ /*39441*/;
assign _34952_ = _34433_ ^ _34954_ /*39444*/;
assign _34953_ = _34945_ & _34952_ /*39442*/;
assign _34882_ = _34945_ ^ _34952_ /*39443*/;
assign _34950_ = _34951_ | _34953_ /*39440*/;
assign _34959_ = ~D[2] /*39439*/;
assign _34956_ = _34434_ & _34959_ /*39435*/;
assign _34957_ = _34434_ ^ _34959_ /*39438*/;
assign _34958_ = _34950_ & _34957_ /*39436*/;
assign _34883_ = _34950_ ^ _34957_ /*39437*/;
assign _34955_ = _34956_ | _34958_ /*39434*/;
assign _34964_ = ~D[3] /*39433*/;
assign _34961_ = _34435_ & _34964_ /*39429*/;
assign _34962_ = _34435_ ^ _34964_ /*39432*/;
assign _34963_ = _34955_ & _34962_ /*39430*/;
assign _34884_ = _34955_ ^ _34962_ /*39431*/;
assign _34960_ = _34961_ | _34963_ /*39428*/;
assign _34969_ = ~D[4] /*39427*/;
assign _34966_ = _34436_ & _34969_ /*39423*/;
assign _34967_ = _34436_ ^ _34969_ /*39426*/;
assign _34968_ = _34960_ & _34967_ /*39424*/;
assign _34885_ = _34960_ ^ _34967_ /*39425*/;
assign _34965_ = _34966_ | _34968_ /*39422*/;
assign _34974_ = ~D[5] /*39421*/;
assign _34971_ = _34437_ & _34974_ /*39417*/;
assign _34972_ = _34437_ ^ _34974_ /*39420*/;
assign _34973_ = _34965_ & _34972_ /*39418*/;
assign _34886_ = _34965_ ^ _34972_ /*39419*/;
assign _34970_ = _34971_ | _34973_ /*39416*/;
assign _34979_ = ~D[6] /*39415*/;
assign _34976_ = _34438_ & _34979_ /*39411*/;
assign _34977_ = _34438_ ^ _34979_ /*39414*/;
assign _34978_ = _34970_ & _34977_ /*39412*/;
assign _34887_ = _34970_ ^ _34977_ /*39413*/;
assign _34975_ = _34976_ | _34978_ /*39410*/;
assign _34984_ = ~D[7] /*39409*/;
assign _34981_ = _34439_ & _34984_ /*39405*/;
assign _34982_ = _34439_ ^ _34984_ /*39408*/;
assign _34983_ = _34975_ & _34982_ /*39406*/;
assign _34888_ = _34975_ ^ _34982_ /*39407*/;
assign _34980_ = _34981_ | _34983_ /*39404*/;
assign _34989_ = ~D[8] /*39403*/;
assign _34986_ = _34440_ & _34989_ /*39399*/;
assign _34987_ = _34440_ ^ _34989_ /*39402*/;
assign _34988_ = _34980_ & _34987_ /*39400*/;
assign _34889_ = _34980_ ^ _34987_ /*39401*/;
assign _34985_ = _34986_ | _34988_ /*39398*/;
assign _34994_ = ~D[9] /*39397*/;
assign _34991_ = _34441_ & _34994_ /*39393*/;
assign _34992_ = _34441_ ^ _34994_ /*39396*/;
assign _34993_ = _34985_ & _34992_ /*39394*/;
assign _34890_ = _34985_ ^ _34992_ /*39395*/;
assign _34990_ = _34991_ | _34993_ /*39392*/;
assign _34999_ = ~D[10] /*39391*/;
assign _34996_ = _34442_ & _34999_ /*39387*/;
assign _34997_ = _34442_ ^ _34999_ /*39390*/;
assign _34998_ = _34990_ & _34997_ /*39388*/;
assign _34891_ = _34990_ ^ _34997_ /*39389*/;
assign _34995_ = _34996_ | _34998_ /*39386*/;
assign _35004_ = ~D[11] /*39385*/;
assign _35001_ = _34443_ & _35004_ /*39381*/;
assign _35002_ = _34443_ ^ _35004_ /*39384*/;
assign _35003_ = _34995_ & _35002_ /*39382*/;
assign _34892_ = _34995_ ^ _35002_ /*39383*/;
assign _35000_ = _35001_ | _35003_ /*39380*/;
assign _35009_ = ~D[12] /*39379*/;
assign _35006_ = _34444_ & _35009_ /*39375*/;
assign _35007_ = _34444_ ^ _35009_ /*39378*/;
assign _35008_ = _35000_ & _35007_ /*39376*/;
assign _34893_ = _35000_ ^ _35007_ /*39377*/;
assign _35005_ = _35006_ | _35008_ /*39374*/;
assign _35014_ = ~D[13] /*39373*/;
assign _35011_ = _34445_ & _35014_ /*39369*/;
assign _35012_ = _34445_ ^ _35014_ /*39372*/;
assign _35013_ = _35005_ & _35012_ /*39370*/;
assign _34894_ = _35005_ ^ _35012_ /*39371*/;
assign _35010_ = _35011_ | _35013_ /*39368*/;
assign _35019_ = ~D[14] /*39367*/;
assign _35016_ = _34446_ & _35019_ /*39363*/;
assign _35017_ = _34446_ ^ _35019_ /*39366*/;
assign _35018_ = _35010_ & _35017_ /*39364*/;
assign _34895_ = _35010_ ^ _35017_ /*39365*/;
assign _35015_ = _35016_ | _35018_ /*39362*/;
assign _35024_ = ~D[15] /*39361*/;
assign _35021_ = _34447_ & _35024_ /*39357*/;
assign _35022_ = _34447_ ^ _35024_ /*39360*/;
assign _35023_ = _35015_ & _35022_ /*39358*/;
assign _34896_ = _35015_ ^ _35022_ /*39359*/;
assign _35020_ = _35021_ | _35023_ /*39356*/;
assign _35029_ = ~D[16] /*39355*/;
assign _35026_ = _34448_ & _35029_ /*39351*/;
assign _35027_ = _34448_ ^ _35029_ /*39354*/;
assign _35028_ = _35020_ & _35027_ /*39352*/;
assign _34897_ = _35020_ ^ _35027_ /*39353*/;
assign _35025_ = _35026_ | _35028_ /*39350*/;
assign _35034_ = ~D[17] /*39349*/;
assign _35031_ = _34449_ & _35034_ /*39345*/;
assign _35032_ = _34449_ ^ _35034_ /*39348*/;
assign _35033_ = _35025_ & _35032_ /*39346*/;
assign _34898_ = _35025_ ^ _35032_ /*39347*/;
assign _35030_ = _35031_ | _35033_ /*39344*/;
assign _35039_ = ~D[18] /*39343*/;
assign _35036_ = _34450_ & _35039_ /*39339*/;
assign _35037_ = _34450_ ^ _35039_ /*39342*/;
assign _35038_ = _35030_ & _35037_ /*39340*/;
assign _34899_ = _35030_ ^ _35037_ /*39341*/;
assign _35035_ = _35036_ | _35038_ /*39338*/;
assign _35044_ = ~D[19] /*39337*/;
assign _35041_ = _34451_ & _35044_ /*39333*/;
assign _35042_ = _34451_ ^ _35044_ /*39336*/;
assign _35043_ = _35035_ & _35042_ /*39334*/;
assign _34900_ = _35035_ ^ _35042_ /*39335*/;
assign _35040_ = _35041_ | _35043_ /*39332*/;
assign _35049_ = ~D[20] /*39331*/;
assign _35046_ = _34452_ & _35049_ /*39327*/;
assign _35047_ = _34452_ ^ _35049_ /*39330*/;
assign _35048_ = _35040_ & _35047_ /*39328*/;
assign _34901_ = _35040_ ^ _35047_ /*39329*/;
assign _35045_ = _35046_ | _35048_ /*39326*/;
assign _35054_ = ~D[21] /*39325*/;
assign _35051_ = _34453_ & _35054_ /*39321*/;
assign _35052_ = _34453_ ^ _35054_ /*39324*/;
assign _35053_ = _35045_ & _35052_ /*39322*/;
assign _34902_ = _35045_ ^ _35052_ /*39323*/;
assign _35050_ = _35051_ | _35053_ /*39320*/;
assign _35059_ = ~D[22] /*39319*/;
assign _35056_ = _34454_ & _35059_ /*39315*/;
assign _35057_ = _34454_ ^ _35059_ /*39318*/;
assign _35058_ = _35050_ & _35057_ /*39316*/;
assign _34903_ = _35050_ ^ _35057_ /*39317*/;
assign _35055_ = _35056_ | _35058_ /*39314*/;
assign _35064_ = ~D[23] /*39313*/;
assign _35061_ = _34455_ & _35064_ /*39309*/;
assign _35062_ = _34455_ ^ _35064_ /*39312*/;
assign _35063_ = _35055_ & _35062_ /*39310*/;
assign _34904_ = _35055_ ^ _35062_ /*39311*/;
assign _35060_ = _35061_ | _35063_ /*39308*/;
assign _35069_ = ~D[24] /*39307*/;
assign _35066_ = _34456_ & _35069_ /*39303*/;
assign _35067_ = _34456_ ^ _35069_ /*39306*/;
assign _35068_ = _35060_ & _35067_ /*39304*/;
assign _34905_ = _35060_ ^ _35067_ /*39305*/;
assign _35065_ = _35066_ | _35068_ /*39302*/;
assign _35074_ = ~D[25] /*39301*/;
assign _35071_ = _34457_ & _35074_ /*39297*/;
assign _35072_ = _34457_ ^ _35074_ /*39300*/;
assign _35073_ = _35065_ & _35072_ /*39298*/;
assign _34906_ = _35065_ ^ _35072_ /*39299*/;
assign _35070_ = _35071_ | _35073_ /*39296*/;
assign _35079_ = ~D[26] /*39295*/;
assign _35076_ = _34458_ & _35079_ /*39291*/;
assign _35077_ = _34458_ ^ _35079_ /*39294*/;
assign _35078_ = _35070_ & _35077_ /*39292*/;
assign _34907_ = _35070_ ^ _35077_ /*39293*/;
assign _35075_ = _35076_ | _35078_ /*39290*/;
assign _35084_ = ~D[27] /*39289*/;
assign _35081_ = _34459_ & _35084_ /*39285*/;
assign _35082_ = _34459_ ^ _35084_ /*39288*/;
assign _35083_ = _35075_ & _35082_ /*39286*/;
assign _34908_ = _35075_ ^ _35082_ /*39287*/;
assign _35080_ = _35081_ | _35083_ /*39284*/;
assign _35089_ = ~D[28] /*39283*/;
assign _35086_ = _34460_ & _35089_ /*39279*/;
assign _35087_ = _34460_ ^ _35089_ /*39282*/;
assign _35088_ = _35080_ & _35087_ /*39280*/;
assign _34909_ = _35080_ ^ _35087_ /*39281*/;
assign _35085_ = _35086_ | _35088_ /*39278*/;
assign _35094_ = ~D[29] /*39277*/;
assign _35091_ = _34461_ & _35094_ /*39273*/;
assign _35092_ = _34461_ ^ _35094_ /*39276*/;
assign _35093_ = _35085_ & _35092_ /*39274*/;
assign _34910_ = _35085_ ^ _35092_ /*39275*/;
assign _35090_ = _35091_ | _35093_ /*39272*/;
assign _35099_ = ~D[30] /*39271*/;
assign _35096_ = _34462_ & _35099_ /*39267*/;
assign _35097_ = _34462_ ^ _35099_ /*39270*/;
assign _35098_ = _35090_ & _35097_ /*39268*/;
assign _34911_ = _35090_ ^ _35097_ /*39269*/;
assign _35095_ = _35096_ | _35098_ /*39266*/;
assign _35104_ = ~D[31] /*39265*/;
assign _35101_ = _34463_ & _35104_ /*39261*/;
assign _35102_ = _34463_ ^ _35104_ /*39264*/;
assign _35103_ = _35095_ & _35102_ /*39262*/;
assign _34912_ = _35095_ ^ _35102_ /*39263*/;
assign _35100_ = _35101_ | _35103_ /*39260*/;
assign _35109_ = ~D[32] /*39259*/;
assign _35106_ = _34464_ & _35109_ /*39255*/;
assign _35107_ = _34464_ ^ _35109_ /*39258*/;
assign _35108_ = _35100_ & _35107_ /*39256*/;
assign _34913_ = _35100_ ^ _35107_ /*39257*/;
assign _35105_ = _35106_ | _35108_ /*39254*/;
assign _35114_ = ~D[33] /*39253*/;
assign _35111_ = _34465_ & _35114_ /*39249*/;
assign _35112_ = _34465_ ^ _35114_ /*39252*/;
assign _35113_ = _35105_ & _35112_ /*39250*/;
assign _34914_ = _35105_ ^ _35112_ /*39251*/;
assign _35110_ = _35111_ | _35113_ /*39248*/;
assign _35119_ = ~D[34] /*39247*/;
assign _35116_ = _34466_ & _35119_ /*39243*/;
assign _35117_ = _34466_ ^ _35119_ /*39246*/;
assign _35118_ = _35110_ & _35117_ /*39244*/;
assign _34915_ = _35110_ ^ _35117_ /*39245*/;
assign _35115_ = _35116_ | _35118_ /*39242*/;
assign _35124_ = ~D[35] /*39241*/;
assign _35121_ = _34467_ & _35124_ /*39237*/;
assign _35122_ = _34467_ ^ _35124_ /*39240*/;
assign _35123_ = _35115_ & _35122_ /*39238*/;
assign _34916_ = _35115_ ^ _35122_ /*39239*/;
assign _35120_ = _35121_ | _35123_ /*39236*/;
assign _35129_ = ~D[36] /*39235*/;
assign _35126_ = _34468_ & _35129_ /*39231*/;
assign _35127_ = _34468_ ^ _35129_ /*39234*/;
assign _35128_ = _35120_ & _35127_ /*39232*/;
assign _34917_ = _35120_ ^ _35127_ /*39233*/;
assign _35125_ = _35126_ | _35128_ /*39230*/;
assign _35134_ = ~D[37] /*39229*/;
assign _35131_ = _34469_ & _35134_ /*39225*/;
assign _35132_ = _34469_ ^ _35134_ /*39228*/;
assign _35133_ = _35125_ & _35132_ /*39226*/;
assign _34918_ = _35125_ ^ _35132_ /*39227*/;
assign _35130_ = _35131_ | _35133_ /*39224*/;
assign _35139_ = ~D[38] /*39223*/;
assign _35136_ = _34470_ & _35139_ /*39219*/;
assign _35137_ = _34470_ ^ _35139_ /*39222*/;
assign _35138_ = _35130_ & _35137_ /*39220*/;
assign _34919_ = _35130_ ^ _35137_ /*39221*/;
assign _35135_ = _35136_ | _35138_ /*39218*/;
assign _35144_ = ~D[39] /*39217*/;
assign _35141_ = _34471_ & _35144_ /*39213*/;
assign _35142_ = _34471_ ^ _35144_ /*39216*/;
assign _35143_ = _35135_ & _35142_ /*39214*/;
assign _34920_ = _35135_ ^ _35142_ /*39215*/;
assign _35140_ = _35141_ | _35143_ /*39212*/;
assign _35149_ = ~D[40] /*39211*/;
assign _35146_ = _34472_ & _35149_ /*39207*/;
assign _35147_ = _34472_ ^ _35149_ /*39210*/;
assign _35148_ = _35140_ & _35147_ /*39208*/;
assign _34921_ = _35140_ ^ _35147_ /*39209*/;
assign _35145_ = _35146_ | _35148_ /*39206*/;
assign _35154_ = ~D[41] /*39205*/;
assign _35151_ = _34473_ & _35154_ /*39201*/;
assign _35152_ = _34473_ ^ _35154_ /*39204*/;
assign _35153_ = _35145_ & _35152_ /*39202*/;
assign _34922_ = _35145_ ^ _35152_ /*39203*/;
assign _35150_ = _35151_ | _35153_ /*39200*/;
assign _35159_ = ~D[42] /*39199*/;
assign _35156_ = _34474_ & _35159_ /*39195*/;
assign _35157_ = _34474_ ^ _35159_ /*39198*/;
assign _35158_ = _35150_ & _35157_ /*39196*/;
assign _34923_ = _35150_ ^ _35157_ /*39197*/;
assign _35155_ = _35156_ | _35158_ /*39194*/;
assign _35164_ = ~D[43] /*39193*/;
assign _35161_ = _34475_ & _35164_ /*39189*/;
assign _35162_ = _34475_ ^ _35164_ /*39192*/;
assign _35163_ = _35155_ & _35162_ /*39190*/;
assign _34924_ = _35155_ ^ _35162_ /*39191*/;
assign _35160_ = _35161_ | _35163_ /*39188*/;
assign _35169_ = ~D[44] /*39187*/;
assign _35166_ = _34476_ & _35169_ /*39183*/;
assign _35167_ = _34476_ ^ _35169_ /*39186*/;
assign _35168_ = _35160_ & _35167_ /*39184*/;
assign _34925_ = _35160_ ^ _35167_ /*39185*/;
assign _35165_ = _35166_ | _35168_ /*39182*/;
assign _35174_ = ~D[45] /*39181*/;
assign _35171_ = _34477_ & _35174_ /*39177*/;
assign _35172_ = _34477_ ^ _35174_ /*39180*/;
assign _35173_ = _35165_ & _35172_ /*39178*/;
assign _34926_ = _35165_ ^ _35172_ /*39179*/;
assign _35170_ = _35171_ | _35173_ /*39176*/;
assign _35179_ = ~D[46] /*39175*/;
assign _35176_ = _34478_ & _35179_ /*39171*/;
assign _35177_ = _34478_ ^ _35179_ /*39174*/;
assign _35178_ = _35170_ & _35177_ /*39172*/;
assign _34927_ = _35170_ ^ _35177_ /*39173*/;
assign _35175_ = _35176_ | _35178_ /*39170*/;
assign _35184_ = ~D[47] /*39169*/;
assign _35181_ = _34479_ & _35184_ /*39165*/;
assign _35182_ = _34479_ ^ _35184_ /*39168*/;
assign _35183_ = _35175_ & _35182_ /*39166*/;
assign _34928_ = _35175_ ^ _35182_ /*39167*/;
assign _35180_ = _35181_ | _35183_ /*39164*/;
assign _35189_ = ~D[48] /*39163*/;
assign _35186_ = _34480_ & _35189_ /*39159*/;
assign _35187_ = _34480_ ^ _35189_ /*39162*/;
assign _35188_ = _35180_ & _35187_ /*39160*/;
assign _34929_ = _35180_ ^ _35187_ /*39161*/;
assign _35185_ = _35186_ | _35188_ /*39158*/;
assign _35194_ = ~D[49] /*39157*/;
assign _35191_ = _34481_ & _35194_ /*39153*/;
assign _35192_ = _34481_ ^ _35194_ /*39156*/;
assign _35193_ = _35185_ & _35192_ /*39154*/;
assign _34930_ = _35185_ ^ _35192_ /*39155*/;
assign _35190_ = _35191_ | _35193_ /*39152*/;
assign _35199_ = ~D[50] /*39151*/;
assign _35196_ = _34482_ & _35199_ /*39147*/;
assign _35197_ = _34482_ ^ _35199_ /*39150*/;
assign _35198_ = _35190_ & _35197_ /*39148*/;
assign _34931_ = _35190_ ^ _35197_ /*39149*/;
assign _35195_ = _35196_ | _35198_ /*39146*/;
assign _35204_ = ~D[51] /*39145*/;
assign _35201_ = _34483_ & _35204_ /*39141*/;
assign _35202_ = _34483_ ^ _35204_ /*39144*/;
assign _35203_ = _35195_ & _35202_ /*39142*/;
assign _34932_ = _35195_ ^ _35202_ /*39143*/;
assign _35200_ = _35201_ | _35203_ /*39140*/;
assign _35209_ = ~D[52] /*39139*/;
assign _35206_ = _34484_ & _35209_ /*39135*/;
assign _35207_ = _34484_ ^ _35209_ /*39138*/;
assign _35208_ = _35200_ & _35207_ /*39136*/;
assign _34933_ = _35200_ ^ _35207_ /*39137*/;
assign _35205_ = _35206_ | _35208_ /*39134*/;
assign _35214_ = ~D[53] /*39133*/;
assign _35211_ = _34485_ & _35214_ /*39129*/;
assign _35212_ = _34485_ ^ _35214_ /*39132*/;
assign _35213_ = _35205_ & _35212_ /*39130*/;
assign _34934_ = _35205_ ^ _35212_ /*39131*/;
assign _35210_ = _35211_ | _35213_ /*39128*/;
assign _35219_ = ~D[54] /*39127*/;
assign _35216_ = _34486_ & _35219_ /*39123*/;
assign _35217_ = _34486_ ^ _35219_ /*39126*/;
assign _35218_ = _35210_ & _35217_ /*39124*/;
assign _34935_ = _35210_ ^ _35217_ /*39125*/;
assign _35215_ = _35216_ | _35218_ /*39122*/;
assign _35224_ = ~D[55] /*39121*/;
assign _35221_ = _34487_ & _35224_ /*39117*/;
assign _35222_ = _34487_ ^ _35224_ /*39120*/;
assign _35223_ = _35215_ & _35222_ /*39118*/;
assign _34936_ = _35215_ ^ _35222_ /*39119*/;
assign _35220_ = _35221_ | _35223_ /*39116*/;
assign _35229_ = ~D[56] /*39115*/;
assign _35226_ = _34488_ & _35229_ /*39111*/;
assign _35227_ = _34488_ ^ _35229_ /*39114*/;
assign _35228_ = _35220_ & _35227_ /*39112*/;
assign _34937_ = _35220_ ^ _35227_ /*39113*/;
assign _35225_ = _35226_ | _35228_ /*39110*/;
assign _35234_ = ~D[57] /*39109*/;
assign _35231_ = _34489_ & _35234_ /*39105*/;
assign _35232_ = _34489_ ^ _35234_ /*39108*/;
assign _35233_ = _35225_ & _35232_ /*39106*/;
assign _34938_ = _35225_ ^ _35232_ /*39107*/;
assign _35230_ = _35231_ | _35233_ /*39104*/;
assign _35239_ = ~D[58] /*39103*/;
assign _35236_ = _34490_ & _35239_ /*39099*/;
assign _35237_ = _34490_ ^ _35239_ /*39102*/;
assign _35238_ = _35230_ & _35237_ /*39100*/;
assign _34939_ = _35230_ ^ _35237_ /*39101*/;
assign _35235_ = _35236_ | _35238_ /*39098*/;
assign _35244_ = ~D[59] /*39097*/;
assign _35241_ = _34491_ & _35244_ /*39093*/;
assign _35242_ = _34491_ ^ _35244_ /*39096*/;
assign _35243_ = _35235_ & _35242_ /*39094*/;
assign _34940_ = _35235_ ^ _35242_ /*39095*/;
assign _35240_ = _35241_ | _35243_ /*39092*/;
assign _35249_ = ~D[60] /*39091*/;
assign _35246_ = _34492_ & _35249_ /*39087*/;
assign _35247_ = _34492_ ^ _35249_ /*39090*/;
assign _35248_ = _35240_ & _35247_ /*39088*/;
assign _34941_ = _35240_ ^ _35247_ /*39089*/;
assign _35245_ = _35246_ | _35248_ /*39086*/;
assign _35254_ = ~D[61] /*39085*/;
assign _35251_ = _34493_ & _35254_ /*39081*/;
assign _35252_ = _34493_ ^ _35254_ /*39084*/;
assign _35253_ = _35245_ & _35252_ /*39082*/;
assign _34942_ = _35245_ ^ _35252_ /*39083*/;
assign _35250_ = _35251_ | _35253_ /*39080*/;
assign _35259_ = ~D[62] /*39079*/;
assign _35256_ = _34494_ & _35259_ /*39075*/;
assign _35257_ = _34494_ ^ _35259_ /*39078*/;
assign _35258_ = _35250_ & _35257_ /*39076*/;
assign _34943_ = _35250_ ^ _35257_ /*39077*/;
assign _35255_ = _35256_ | _35258_ /*39074*/;
assign _35260_ = _34495_ & oneWire /*39069*/;
assign _35261_ = _34495_ ^ oneWire /*39072*/;
assign _35262_ = _35255_ & _35261_ /*39070*/;
assign _34944_ = _35255_ ^ _35261_ /*39071*/;
assign Q[24] = _35260_ | _35262_ /*39068*/;
assign _35395_ = ~Q[24] /*38683*/;
assign _35394_ = _35395_ & D[0] /*38682*/;
assign _35397_ = _34881_ & _35394_ /*38677*/;
assign _35398_ = _34881_ ^ _35394_ /*38680*/;
assign _35399_ = zeroWire & _35398_ /*38678*/;
assign _35329_ = zeroWire ^ _35398_ /*38679*/;
assign _35396_ = _35397_ | _35399_ /*38676*/;
assign _35401_ = ~Q[24] /*38675*/;
assign _35400_ = _35401_ & D[1] /*38674*/;
assign _35403_ = _34882_ & _35400_ /*38669*/;
assign _35404_ = _34882_ ^ _35400_ /*38672*/;
assign _35405_ = _35396_ & _35404_ /*38670*/;
assign _35330_ = _35396_ ^ _35404_ /*38671*/;
assign _35402_ = _35403_ | _35405_ /*38668*/;
assign _35407_ = ~Q[24] /*38667*/;
assign _35406_ = _35407_ & D[2] /*38666*/;
assign _35409_ = _34883_ & _35406_ /*38661*/;
assign _35410_ = _34883_ ^ _35406_ /*38664*/;
assign _35411_ = _35402_ & _35410_ /*38662*/;
assign _35331_ = _35402_ ^ _35410_ /*38663*/;
assign _35408_ = _35409_ | _35411_ /*38660*/;
assign _35413_ = ~Q[24] /*38659*/;
assign _35412_ = _35413_ & D[3] /*38658*/;
assign _35415_ = _34884_ & _35412_ /*38653*/;
assign _35416_ = _34884_ ^ _35412_ /*38656*/;
assign _35417_ = _35408_ & _35416_ /*38654*/;
assign _35332_ = _35408_ ^ _35416_ /*38655*/;
assign _35414_ = _35415_ | _35417_ /*38652*/;
assign _35419_ = ~Q[24] /*38651*/;
assign _35418_ = _35419_ & D[4] /*38650*/;
assign _35421_ = _34885_ & _35418_ /*38645*/;
assign _35422_ = _34885_ ^ _35418_ /*38648*/;
assign _35423_ = _35414_ & _35422_ /*38646*/;
assign _35333_ = _35414_ ^ _35422_ /*38647*/;
assign _35420_ = _35421_ | _35423_ /*38644*/;
assign _35425_ = ~Q[24] /*38643*/;
assign _35424_ = _35425_ & D[5] /*38642*/;
assign _35427_ = _34886_ & _35424_ /*38637*/;
assign _35428_ = _34886_ ^ _35424_ /*38640*/;
assign _35429_ = _35420_ & _35428_ /*38638*/;
assign _35334_ = _35420_ ^ _35428_ /*38639*/;
assign _35426_ = _35427_ | _35429_ /*38636*/;
assign _35431_ = ~Q[24] /*38635*/;
assign _35430_ = _35431_ & D[6] /*38634*/;
assign _35433_ = _34887_ & _35430_ /*38629*/;
assign _35434_ = _34887_ ^ _35430_ /*38632*/;
assign _35435_ = _35426_ & _35434_ /*38630*/;
assign _35335_ = _35426_ ^ _35434_ /*38631*/;
assign _35432_ = _35433_ | _35435_ /*38628*/;
assign _35437_ = ~Q[24] /*38627*/;
assign _35436_ = _35437_ & D[7] /*38626*/;
assign _35439_ = _34888_ & _35436_ /*38621*/;
assign _35440_ = _34888_ ^ _35436_ /*38624*/;
assign _35441_ = _35432_ & _35440_ /*38622*/;
assign _35336_ = _35432_ ^ _35440_ /*38623*/;
assign _35438_ = _35439_ | _35441_ /*38620*/;
assign _35443_ = ~Q[24] /*38619*/;
assign _35442_ = _35443_ & D[8] /*38618*/;
assign _35445_ = _34889_ & _35442_ /*38613*/;
assign _35446_ = _34889_ ^ _35442_ /*38616*/;
assign _35447_ = _35438_ & _35446_ /*38614*/;
assign _35337_ = _35438_ ^ _35446_ /*38615*/;
assign _35444_ = _35445_ | _35447_ /*38612*/;
assign _35449_ = ~Q[24] /*38611*/;
assign _35448_ = _35449_ & D[9] /*38610*/;
assign _35451_ = _34890_ & _35448_ /*38605*/;
assign _35452_ = _34890_ ^ _35448_ /*38608*/;
assign _35453_ = _35444_ & _35452_ /*38606*/;
assign _35338_ = _35444_ ^ _35452_ /*38607*/;
assign _35450_ = _35451_ | _35453_ /*38604*/;
assign _35455_ = ~Q[24] /*38603*/;
assign _35454_ = _35455_ & D[10] /*38602*/;
assign _35457_ = _34891_ & _35454_ /*38597*/;
assign _35458_ = _34891_ ^ _35454_ /*38600*/;
assign _35459_ = _35450_ & _35458_ /*38598*/;
assign _35339_ = _35450_ ^ _35458_ /*38599*/;
assign _35456_ = _35457_ | _35459_ /*38596*/;
assign _35461_ = ~Q[24] /*38595*/;
assign _35460_ = _35461_ & D[11] /*38594*/;
assign _35463_ = _34892_ & _35460_ /*38589*/;
assign _35464_ = _34892_ ^ _35460_ /*38592*/;
assign _35465_ = _35456_ & _35464_ /*38590*/;
assign _35340_ = _35456_ ^ _35464_ /*38591*/;
assign _35462_ = _35463_ | _35465_ /*38588*/;
assign _35467_ = ~Q[24] /*38587*/;
assign _35466_ = _35467_ & D[12] /*38586*/;
assign _35469_ = _34893_ & _35466_ /*38581*/;
assign _35470_ = _34893_ ^ _35466_ /*38584*/;
assign _35471_ = _35462_ & _35470_ /*38582*/;
assign _35341_ = _35462_ ^ _35470_ /*38583*/;
assign _35468_ = _35469_ | _35471_ /*38580*/;
assign _35473_ = ~Q[24] /*38579*/;
assign _35472_ = _35473_ & D[13] /*38578*/;
assign _35475_ = _34894_ & _35472_ /*38573*/;
assign _35476_ = _34894_ ^ _35472_ /*38576*/;
assign _35477_ = _35468_ & _35476_ /*38574*/;
assign _35342_ = _35468_ ^ _35476_ /*38575*/;
assign _35474_ = _35475_ | _35477_ /*38572*/;
assign _35479_ = ~Q[24] /*38571*/;
assign _35478_ = _35479_ & D[14] /*38570*/;
assign _35481_ = _34895_ & _35478_ /*38565*/;
assign _35482_ = _34895_ ^ _35478_ /*38568*/;
assign _35483_ = _35474_ & _35482_ /*38566*/;
assign _35343_ = _35474_ ^ _35482_ /*38567*/;
assign _35480_ = _35481_ | _35483_ /*38564*/;
assign _35485_ = ~Q[24] /*38563*/;
assign _35484_ = _35485_ & D[15] /*38562*/;
assign _35487_ = _34896_ & _35484_ /*38557*/;
assign _35488_ = _34896_ ^ _35484_ /*38560*/;
assign _35489_ = _35480_ & _35488_ /*38558*/;
assign _35344_ = _35480_ ^ _35488_ /*38559*/;
assign _35486_ = _35487_ | _35489_ /*38556*/;
assign _35491_ = ~Q[24] /*38555*/;
assign _35490_ = _35491_ & D[16] /*38554*/;
assign _35493_ = _34897_ & _35490_ /*38549*/;
assign _35494_ = _34897_ ^ _35490_ /*38552*/;
assign _35495_ = _35486_ & _35494_ /*38550*/;
assign _35345_ = _35486_ ^ _35494_ /*38551*/;
assign _35492_ = _35493_ | _35495_ /*38548*/;
assign _35497_ = ~Q[24] /*38547*/;
assign _35496_ = _35497_ & D[17] /*38546*/;
assign _35499_ = _34898_ & _35496_ /*38541*/;
assign _35500_ = _34898_ ^ _35496_ /*38544*/;
assign _35501_ = _35492_ & _35500_ /*38542*/;
assign _35346_ = _35492_ ^ _35500_ /*38543*/;
assign _35498_ = _35499_ | _35501_ /*38540*/;
assign _35503_ = ~Q[24] /*38539*/;
assign _35502_ = _35503_ & D[18] /*38538*/;
assign _35505_ = _34899_ & _35502_ /*38533*/;
assign _35506_ = _34899_ ^ _35502_ /*38536*/;
assign _35507_ = _35498_ & _35506_ /*38534*/;
assign _35347_ = _35498_ ^ _35506_ /*38535*/;
assign _35504_ = _35505_ | _35507_ /*38532*/;
assign _35509_ = ~Q[24] /*38531*/;
assign _35508_ = _35509_ & D[19] /*38530*/;
assign _35511_ = _34900_ & _35508_ /*38525*/;
assign _35512_ = _34900_ ^ _35508_ /*38528*/;
assign _35513_ = _35504_ & _35512_ /*38526*/;
assign _35348_ = _35504_ ^ _35512_ /*38527*/;
assign _35510_ = _35511_ | _35513_ /*38524*/;
assign _35515_ = ~Q[24] /*38523*/;
assign _35514_ = _35515_ & D[20] /*38522*/;
assign _35517_ = _34901_ & _35514_ /*38517*/;
assign _35518_ = _34901_ ^ _35514_ /*38520*/;
assign _35519_ = _35510_ & _35518_ /*38518*/;
assign _35349_ = _35510_ ^ _35518_ /*38519*/;
assign _35516_ = _35517_ | _35519_ /*38516*/;
assign _35521_ = ~Q[24] /*38515*/;
assign _35520_ = _35521_ & D[21] /*38514*/;
assign _35523_ = _34902_ & _35520_ /*38509*/;
assign _35524_ = _34902_ ^ _35520_ /*38512*/;
assign _35525_ = _35516_ & _35524_ /*38510*/;
assign _35350_ = _35516_ ^ _35524_ /*38511*/;
assign _35522_ = _35523_ | _35525_ /*38508*/;
assign _35527_ = ~Q[24] /*38507*/;
assign _35526_ = _35527_ & D[22] /*38506*/;
assign _35529_ = _34903_ & _35526_ /*38501*/;
assign _35530_ = _34903_ ^ _35526_ /*38504*/;
assign _35531_ = _35522_ & _35530_ /*38502*/;
assign _35351_ = _35522_ ^ _35530_ /*38503*/;
assign _35528_ = _35529_ | _35531_ /*38500*/;
assign _35533_ = ~Q[24] /*38499*/;
assign _35532_ = _35533_ & D[23] /*38498*/;
assign _35535_ = _34904_ & _35532_ /*38493*/;
assign _35536_ = _34904_ ^ _35532_ /*38496*/;
assign _35537_ = _35528_ & _35536_ /*38494*/;
assign _35352_ = _35528_ ^ _35536_ /*38495*/;
assign _35534_ = _35535_ | _35537_ /*38492*/;
assign _35539_ = ~Q[24] /*38491*/;
assign _35538_ = _35539_ & D[24] /*38490*/;
assign _35541_ = _34905_ & _35538_ /*38485*/;
assign _35542_ = _34905_ ^ _35538_ /*38488*/;
assign _35543_ = _35534_ & _35542_ /*38486*/;
assign _35353_ = _35534_ ^ _35542_ /*38487*/;
assign _35540_ = _35541_ | _35543_ /*38484*/;
assign _35545_ = ~Q[24] /*38483*/;
assign _35544_ = _35545_ & D[25] /*38482*/;
assign _35547_ = _34906_ & _35544_ /*38477*/;
assign _35548_ = _34906_ ^ _35544_ /*38480*/;
assign _35549_ = _35540_ & _35548_ /*38478*/;
assign _35354_ = _35540_ ^ _35548_ /*38479*/;
assign _35546_ = _35547_ | _35549_ /*38476*/;
assign _35551_ = ~Q[24] /*38475*/;
assign _35550_ = _35551_ & D[26] /*38474*/;
assign _35553_ = _34907_ & _35550_ /*38469*/;
assign _35554_ = _34907_ ^ _35550_ /*38472*/;
assign _35555_ = _35546_ & _35554_ /*38470*/;
assign _35355_ = _35546_ ^ _35554_ /*38471*/;
assign _35552_ = _35553_ | _35555_ /*38468*/;
assign _35557_ = ~Q[24] /*38467*/;
assign _35556_ = _35557_ & D[27] /*38466*/;
assign _35559_ = _34908_ & _35556_ /*38461*/;
assign _35560_ = _34908_ ^ _35556_ /*38464*/;
assign _35561_ = _35552_ & _35560_ /*38462*/;
assign _35356_ = _35552_ ^ _35560_ /*38463*/;
assign _35558_ = _35559_ | _35561_ /*38460*/;
assign _35563_ = ~Q[24] /*38459*/;
assign _35562_ = _35563_ & D[28] /*38458*/;
assign _35565_ = _34909_ & _35562_ /*38453*/;
assign _35566_ = _34909_ ^ _35562_ /*38456*/;
assign _35567_ = _35558_ & _35566_ /*38454*/;
assign _35357_ = _35558_ ^ _35566_ /*38455*/;
assign _35564_ = _35565_ | _35567_ /*38452*/;
assign _35569_ = ~Q[24] /*38451*/;
assign _35568_ = _35569_ & D[29] /*38450*/;
assign _35571_ = _34910_ & _35568_ /*38445*/;
assign _35572_ = _34910_ ^ _35568_ /*38448*/;
assign _35573_ = _35564_ & _35572_ /*38446*/;
assign _35358_ = _35564_ ^ _35572_ /*38447*/;
assign _35570_ = _35571_ | _35573_ /*38444*/;
assign _35575_ = ~Q[24] /*38443*/;
assign _35574_ = _35575_ & D[30] /*38442*/;
assign _35577_ = _34911_ & _35574_ /*38437*/;
assign _35578_ = _34911_ ^ _35574_ /*38440*/;
assign _35579_ = _35570_ & _35578_ /*38438*/;
assign _35359_ = _35570_ ^ _35578_ /*38439*/;
assign _35576_ = _35577_ | _35579_ /*38436*/;
assign _35581_ = ~Q[24] /*38435*/;
assign _35580_ = _35581_ & D[31] /*38434*/;
assign _35583_ = _34912_ & _35580_ /*38429*/;
assign _35584_ = _34912_ ^ _35580_ /*38432*/;
assign _35585_ = _35576_ & _35584_ /*38430*/;
assign _35360_ = _35576_ ^ _35584_ /*38431*/;
assign _35582_ = _35583_ | _35585_ /*38428*/;
assign _35587_ = ~Q[24] /*38427*/;
assign _35586_ = _35587_ & D[32] /*38426*/;
assign _35589_ = _34913_ & _35586_ /*38421*/;
assign _35590_ = _34913_ ^ _35586_ /*38424*/;
assign _35591_ = _35582_ & _35590_ /*38422*/;
assign _35361_ = _35582_ ^ _35590_ /*38423*/;
assign _35588_ = _35589_ | _35591_ /*38420*/;
assign _35593_ = ~Q[24] /*38419*/;
assign _35592_ = _35593_ & D[33] /*38418*/;
assign _35595_ = _34914_ & _35592_ /*38413*/;
assign _35596_ = _34914_ ^ _35592_ /*38416*/;
assign _35597_ = _35588_ & _35596_ /*38414*/;
assign _35362_ = _35588_ ^ _35596_ /*38415*/;
assign _35594_ = _35595_ | _35597_ /*38412*/;
assign _35599_ = ~Q[24] /*38411*/;
assign _35598_ = _35599_ & D[34] /*38410*/;
assign _35601_ = _34915_ & _35598_ /*38405*/;
assign _35602_ = _34915_ ^ _35598_ /*38408*/;
assign _35603_ = _35594_ & _35602_ /*38406*/;
assign _35363_ = _35594_ ^ _35602_ /*38407*/;
assign _35600_ = _35601_ | _35603_ /*38404*/;
assign _35605_ = ~Q[24] /*38403*/;
assign _35604_ = _35605_ & D[35] /*38402*/;
assign _35607_ = _34916_ & _35604_ /*38397*/;
assign _35608_ = _34916_ ^ _35604_ /*38400*/;
assign _35609_ = _35600_ & _35608_ /*38398*/;
assign _35364_ = _35600_ ^ _35608_ /*38399*/;
assign _35606_ = _35607_ | _35609_ /*38396*/;
assign _35611_ = ~Q[24] /*38395*/;
assign _35610_ = _35611_ & D[36] /*38394*/;
assign _35613_ = _34917_ & _35610_ /*38389*/;
assign _35614_ = _34917_ ^ _35610_ /*38392*/;
assign _35615_ = _35606_ & _35614_ /*38390*/;
assign _35365_ = _35606_ ^ _35614_ /*38391*/;
assign _35612_ = _35613_ | _35615_ /*38388*/;
assign _35617_ = ~Q[24] /*38387*/;
assign _35616_ = _35617_ & D[37] /*38386*/;
assign _35619_ = _34918_ & _35616_ /*38381*/;
assign _35620_ = _34918_ ^ _35616_ /*38384*/;
assign _35621_ = _35612_ & _35620_ /*38382*/;
assign _35366_ = _35612_ ^ _35620_ /*38383*/;
assign _35618_ = _35619_ | _35621_ /*38380*/;
assign _35623_ = ~Q[24] /*38379*/;
assign _35622_ = _35623_ & D[38] /*38378*/;
assign _35625_ = _34919_ & _35622_ /*38373*/;
assign _35626_ = _34919_ ^ _35622_ /*38376*/;
assign _35627_ = _35618_ & _35626_ /*38374*/;
assign _35367_ = _35618_ ^ _35626_ /*38375*/;
assign _35624_ = _35625_ | _35627_ /*38372*/;
assign _35629_ = ~Q[24] /*38371*/;
assign _35628_ = _35629_ & D[39] /*38370*/;
assign _35631_ = _34920_ & _35628_ /*38365*/;
assign _35632_ = _34920_ ^ _35628_ /*38368*/;
assign _35633_ = _35624_ & _35632_ /*38366*/;
assign _35368_ = _35624_ ^ _35632_ /*38367*/;
assign _35630_ = _35631_ | _35633_ /*38364*/;
assign _35635_ = ~Q[24] /*38363*/;
assign _35634_ = _35635_ & D[40] /*38362*/;
assign _35637_ = _34921_ & _35634_ /*38357*/;
assign _35638_ = _34921_ ^ _35634_ /*38360*/;
assign _35639_ = _35630_ & _35638_ /*38358*/;
assign _35369_ = _35630_ ^ _35638_ /*38359*/;
assign _35636_ = _35637_ | _35639_ /*38356*/;
assign _35641_ = ~Q[24] /*38355*/;
assign _35640_ = _35641_ & D[41] /*38354*/;
assign _35643_ = _34922_ & _35640_ /*38349*/;
assign _35644_ = _34922_ ^ _35640_ /*38352*/;
assign _35645_ = _35636_ & _35644_ /*38350*/;
assign _35370_ = _35636_ ^ _35644_ /*38351*/;
assign _35642_ = _35643_ | _35645_ /*38348*/;
assign _35647_ = ~Q[24] /*38347*/;
assign _35646_ = _35647_ & D[42] /*38346*/;
assign _35649_ = _34923_ & _35646_ /*38341*/;
assign _35650_ = _34923_ ^ _35646_ /*38344*/;
assign _35651_ = _35642_ & _35650_ /*38342*/;
assign _35371_ = _35642_ ^ _35650_ /*38343*/;
assign _35648_ = _35649_ | _35651_ /*38340*/;
assign _35653_ = ~Q[24] /*38339*/;
assign _35652_ = _35653_ & D[43] /*38338*/;
assign _35655_ = _34924_ & _35652_ /*38333*/;
assign _35656_ = _34924_ ^ _35652_ /*38336*/;
assign _35657_ = _35648_ & _35656_ /*38334*/;
assign _35372_ = _35648_ ^ _35656_ /*38335*/;
assign _35654_ = _35655_ | _35657_ /*38332*/;
assign _35659_ = ~Q[24] /*38331*/;
assign _35658_ = _35659_ & D[44] /*38330*/;
assign _35661_ = _34925_ & _35658_ /*38325*/;
assign _35662_ = _34925_ ^ _35658_ /*38328*/;
assign _35663_ = _35654_ & _35662_ /*38326*/;
assign _35373_ = _35654_ ^ _35662_ /*38327*/;
assign _35660_ = _35661_ | _35663_ /*38324*/;
assign _35665_ = ~Q[24] /*38323*/;
assign _35664_ = _35665_ & D[45] /*38322*/;
assign _35667_ = _34926_ & _35664_ /*38317*/;
assign _35668_ = _34926_ ^ _35664_ /*38320*/;
assign _35669_ = _35660_ & _35668_ /*38318*/;
assign _35374_ = _35660_ ^ _35668_ /*38319*/;
assign _35666_ = _35667_ | _35669_ /*38316*/;
assign _35671_ = ~Q[24] /*38315*/;
assign _35670_ = _35671_ & D[46] /*38314*/;
assign _35673_ = _34927_ & _35670_ /*38309*/;
assign _35674_ = _34927_ ^ _35670_ /*38312*/;
assign _35675_ = _35666_ & _35674_ /*38310*/;
assign _35375_ = _35666_ ^ _35674_ /*38311*/;
assign _35672_ = _35673_ | _35675_ /*38308*/;
assign _35677_ = ~Q[24] /*38307*/;
assign _35676_ = _35677_ & D[47] /*38306*/;
assign _35679_ = _34928_ & _35676_ /*38301*/;
assign _35680_ = _34928_ ^ _35676_ /*38304*/;
assign _35681_ = _35672_ & _35680_ /*38302*/;
assign _35376_ = _35672_ ^ _35680_ /*38303*/;
assign _35678_ = _35679_ | _35681_ /*38300*/;
assign _35683_ = ~Q[24] /*38299*/;
assign _35682_ = _35683_ & D[48] /*38298*/;
assign _35685_ = _34929_ & _35682_ /*38293*/;
assign _35686_ = _34929_ ^ _35682_ /*38296*/;
assign _35687_ = _35678_ & _35686_ /*38294*/;
assign _35377_ = _35678_ ^ _35686_ /*38295*/;
assign _35684_ = _35685_ | _35687_ /*38292*/;
assign _35689_ = ~Q[24] /*38291*/;
assign _35688_ = _35689_ & D[49] /*38290*/;
assign _35691_ = _34930_ & _35688_ /*38285*/;
assign _35692_ = _34930_ ^ _35688_ /*38288*/;
assign _35693_ = _35684_ & _35692_ /*38286*/;
assign _35378_ = _35684_ ^ _35692_ /*38287*/;
assign _35690_ = _35691_ | _35693_ /*38284*/;
assign _35695_ = ~Q[24] /*38283*/;
assign _35694_ = _35695_ & D[50] /*38282*/;
assign _35697_ = _34931_ & _35694_ /*38277*/;
assign _35698_ = _34931_ ^ _35694_ /*38280*/;
assign _35699_ = _35690_ & _35698_ /*38278*/;
assign _35379_ = _35690_ ^ _35698_ /*38279*/;
assign _35696_ = _35697_ | _35699_ /*38276*/;
assign _35701_ = ~Q[24] /*38275*/;
assign _35700_ = _35701_ & D[51] /*38274*/;
assign _35703_ = _34932_ & _35700_ /*38269*/;
assign _35704_ = _34932_ ^ _35700_ /*38272*/;
assign _35705_ = _35696_ & _35704_ /*38270*/;
assign _35380_ = _35696_ ^ _35704_ /*38271*/;
assign _35702_ = _35703_ | _35705_ /*38268*/;
assign _35707_ = ~Q[24] /*38267*/;
assign _35706_ = _35707_ & D[52] /*38266*/;
assign _35709_ = _34933_ & _35706_ /*38261*/;
assign _35710_ = _34933_ ^ _35706_ /*38264*/;
assign _35711_ = _35702_ & _35710_ /*38262*/;
assign _35381_ = _35702_ ^ _35710_ /*38263*/;
assign _35708_ = _35709_ | _35711_ /*38260*/;
assign _35713_ = ~Q[24] /*38259*/;
assign _35712_ = _35713_ & D[53] /*38258*/;
assign _35715_ = _34934_ & _35712_ /*38253*/;
assign _35716_ = _34934_ ^ _35712_ /*38256*/;
assign _35717_ = _35708_ & _35716_ /*38254*/;
assign _35382_ = _35708_ ^ _35716_ /*38255*/;
assign _35714_ = _35715_ | _35717_ /*38252*/;
assign _35719_ = ~Q[24] /*38251*/;
assign _35718_ = _35719_ & D[54] /*38250*/;
assign _35721_ = _34935_ & _35718_ /*38245*/;
assign _35722_ = _34935_ ^ _35718_ /*38248*/;
assign _35723_ = _35714_ & _35722_ /*38246*/;
assign _35383_ = _35714_ ^ _35722_ /*38247*/;
assign _35720_ = _35721_ | _35723_ /*38244*/;
assign _35725_ = ~Q[24] /*38243*/;
assign _35724_ = _35725_ & D[55] /*38242*/;
assign _35727_ = _34936_ & _35724_ /*38237*/;
assign _35728_ = _34936_ ^ _35724_ /*38240*/;
assign _35729_ = _35720_ & _35728_ /*38238*/;
assign _35384_ = _35720_ ^ _35728_ /*38239*/;
assign _35726_ = _35727_ | _35729_ /*38236*/;
assign _35731_ = ~Q[24] /*38235*/;
assign _35730_ = _35731_ & D[56] /*38234*/;
assign _35733_ = _34937_ & _35730_ /*38229*/;
assign _35734_ = _34937_ ^ _35730_ /*38232*/;
assign _35735_ = _35726_ & _35734_ /*38230*/;
assign _35385_ = _35726_ ^ _35734_ /*38231*/;
assign _35732_ = _35733_ | _35735_ /*38228*/;
assign _35737_ = ~Q[24] /*38227*/;
assign _35736_ = _35737_ & D[57] /*38226*/;
assign _35739_ = _34938_ & _35736_ /*38221*/;
assign _35740_ = _34938_ ^ _35736_ /*38224*/;
assign _35741_ = _35732_ & _35740_ /*38222*/;
assign _35386_ = _35732_ ^ _35740_ /*38223*/;
assign _35738_ = _35739_ | _35741_ /*38220*/;
assign _35743_ = ~Q[24] /*38219*/;
assign _35742_ = _35743_ & D[58] /*38218*/;
assign _35745_ = _34939_ & _35742_ /*38213*/;
assign _35746_ = _34939_ ^ _35742_ /*38216*/;
assign _35747_ = _35738_ & _35746_ /*38214*/;
assign _35387_ = _35738_ ^ _35746_ /*38215*/;
assign _35744_ = _35745_ | _35747_ /*38212*/;
assign _35749_ = ~Q[24] /*38211*/;
assign _35748_ = _35749_ & D[59] /*38210*/;
assign _35751_ = _34940_ & _35748_ /*38205*/;
assign _35752_ = _34940_ ^ _35748_ /*38208*/;
assign _35753_ = _35744_ & _35752_ /*38206*/;
assign _35388_ = _35744_ ^ _35752_ /*38207*/;
assign _35750_ = _35751_ | _35753_ /*38204*/;
assign _35755_ = ~Q[24] /*38203*/;
assign _35754_ = _35755_ & D[60] /*38202*/;
assign _35757_ = _34941_ & _35754_ /*38197*/;
assign _35758_ = _34941_ ^ _35754_ /*38200*/;
assign _35759_ = _35750_ & _35758_ /*38198*/;
assign _35389_ = _35750_ ^ _35758_ /*38199*/;
assign _35756_ = _35757_ | _35759_ /*38196*/;
assign _35761_ = ~Q[24] /*38195*/;
assign _35760_ = _35761_ & D[61] /*38194*/;
assign _35763_ = _34942_ & _35760_ /*38189*/;
assign _35764_ = _34942_ ^ _35760_ /*38192*/;
assign _35765_ = _35756_ & _35764_ /*38190*/;
assign _35390_ = _35756_ ^ _35764_ /*38191*/;
assign _35762_ = _35763_ | _35765_ /*38188*/;
assign _35767_ = ~Q[24] /*38187*/;
assign _35766_ = _35767_ & D[62] /*38186*/;
assign _35769_ = _34943_ & _35766_ /*38181*/;
assign _35770_ = _34943_ ^ _35766_ /*38184*/;
assign _35771_ = _35762_ & _35770_ /*38182*/;
assign _35391_ = _35762_ ^ _35770_ /*38183*/;
assign _35768_ = _35769_ | _35771_ /*38180*/;
assign _35773_ = ~Q[24] /*38179*/;
assign _35772_ = _35773_ & zeroWire /*38178*/;
assign _35774_ = _34944_ ^ _35772_ /*38176*/;
assign _35392_ = _35774_ ^ _35768_ /*38175*/;
assign _35845_ = ~D[0] /*37921*/;
assign _35842_ = R_0[23] & _35845_ /*37917*/;
assign _35843_ = R_0[23] ^ _35845_ /*37920*/;
assign _35844_ = oneWire & _35843_ /*37918*/;
assign _35777_ = oneWire ^ _35843_ /*37919*/;
assign _35841_ = _35842_ | _35844_ /*37916*/;
assign _35850_ = ~D[1] /*37915*/;
assign _35847_ = _35329_ & _35850_ /*37911*/;
assign _35848_ = _35329_ ^ _35850_ /*37914*/;
assign _35849_ = _35841_ & _35848_ /*37912*/;
assign _35778_ = _35841_ ^ _35848_ /*37913*/;
assign _35846_ = _35847_ | _35849_ /*37910*/;
assign _35855_ = ~D[2] /*37909*/;
assign _35852_ = _35330_ & _35855_ /*37905*/;
assign _35853_ = _35330_ ^ _35855_ /*37908*/;
assign _35854_ = _35846_ & _35853_ /*37906*/;
assign _35779_ = _35846_ ^ _35853_ /*37907*/;
assign _35851_ = _35852_ | _35854_ /*37904*/;
assign _35860_ = ~D[3] /*37903*/;
assign _35857_ = _35331_ & _35860_ /*37899*/;
assign _35858_ = _35331_ ^ _35860_ /*37902*/;
assign _35859_ = _35851_ & _35858_ /*37900*/;
assign _35780_ = _35851_ ^ _35858_ /*37901*/;
assign _35856_ = _35857_ | _35859_ /*37898*/;
assign _35865_ = ~D[4] /*37897*/;
assign _35862_ = _35332_ & _35865_ /*37893*/;
assign _35863_ = _35332_ ^ _35865_ /*37896*/;
assign _35864_ = _35856_ & _35863_ /*37894*/;
assign _35781_ = _35856_ ^ _35863_ /*37895*/;
assign _35861_ = _35862_ | _35864_ /*37892*/;
assign _35870_ = ~D[5] /*37891*/;
assign _35867_ = _35333_ & _35870_ /*37887*/;
assign _35868_ = _35333_ ^ _35870_ /*37890*/;
assign _35869_ = _35861_ & _35868_ /*37888*/;
assign _35782_ = _35861_ ^ _35868_ /*37889*/;
assign _35866_ = _35867_ | _35869_ /*37886*/;
assign _35875_ = ~D[6] /*37885*/;
assign _35872_ = _35334_ & _35875_ /*37881*/;
assign _35873_ = _35334_ ^ _35875_ /*37884*/;
assign _35874_ = _35866_ & _35873_ /*37882*/;
assign _35783_ = _35866_ ^ _35873_ /*37883*/;
assign _35871_ = _35872_ | _35874_ /*37880*/;
assign _35880_ = ~D[7] /*37879*/;
assign _35877_ = _35335_ & _35880_ /*37875*/;
assign _35878_ = _35335_ ^ _35880_ /*37878*/;
assign _35879_ = _35871_ & _35878_ /*37876*/;
assign _35784_ = _35871_ ^ _35878_ /*37877*/;
assign _35876_ = _35877_ | _35879_ /*37874*/;
assign _35885_ = ~D[8] /*37873*/;
assign _35882_ = _35336_ & _35885_ /*37869*/;
assign _35883_ = _35336_ ^ _35885_ /*37872*/;
assign _35884_ = _35876_ & _35883_ /*37870*/;
assign _35785_ = _35876_ ^ _35883_ /*37871*/;
assign _35881_ = _35882_ | _35884_ /*37868*/;
assign _35890_ = ~D[9] /*37867*/;
assign _35887_ = _35337_ & _35890_ /*37863*/;
assign _35888_ = _35337_ ^ _35890_ /*37866*/;
assign _35889_ = _35881_ & _35888_ /*37864*/;
assign _35786_ = _35881_ ^ _35888_ /*37865*/;
assign _35886_ = _35887_ | _35889_ /*37862*/;
assign _35895_ = ~D[10] /*37861*/;
assign _35892_ = _35338_ & _35895_ /*37857*/;
assign _35893_ = _35338_ ^ _35895_ /*37860*/;
assign _35894_ = _35886_ & _35893_ /*37858*/;
assign _35787_ = _35886_ ^ _35893_ /*37859*/;
assign _35891_ = _35892_ | _35894_ /*37856*/;
assign _35900_ = ~D[11] /*37855*/;
assign _35897_ = _35339_ & _35900_ /*37851*/;
assign _35898_ = _35339_ ^ _35900_ /*37854*/;
assign _35899_ = _35891_ & _35898_ /*37852*/;
assign _35788_ = _35891_ ^ _35898_ /*37853*/;
assign _35896_ = _35897_ | _35899_ /*37850*/;
assign _35905_ = ~D[12] /*37849*/;
assign _35902_ = _35340_ & _35905_ /*37845*/;
assign _35903_ = _35340_ ^ _35905_ /*37848*/;
assign _35904_ = _35896_ & _35903_ /*37846*/;
assign _35789_ = _35896_ ^ _35903_ /*37847*/;
assign _35901_ = _35902_ | _35904_ /*37844*/;
assign _35910_ = ~D[13] /*37843*/;
assign _35907_ = _35341_ & _35910_ /*37839*/;
assign _35908_ = _35341_ ^ _35910_ /*37842*/;
assign _35909_ = _35901_ & _35908_ /*37840*/;
assign _35790_ = _35901_ ^ _35908_ /*37841*/;
assign _35906_ = _35907_ | _35909_ /*37838*/;
assign _35915_ = ~D[14] /*37837*/;
assign _35912_ = _35342_ & _35915_ /*37833*/;
assign _35913_ = _35342_ ^ _35915_ /*37836*/;
assign _35914_ = _35906_ & _35913_ /*37834*/;
assign _35791_ = _35906_ ^ _35913_ /*37835*/;
assign _35911_ = _35912_ | _35914_ /*37832*/;
assign _35920_ = ~D[15] /*37831*/;
assign _35917_ = _35343_ & _35920_ /*37827*/;
assign _35918_ = _35343_ ^ _35920_ /*37830*/;
assign _35919_ = _35911_ & _35918_ /*37828*/;
assign _35792_ = _35911_ ^ _35918_ /*37829*/;
assign _35916_ = _35917_ | _35919_ /*37826*/;
assign _35925_ = ~D[16] /*37825*/;
assign _35922_ = _35344_ & _35925_ /*37821*/;
assign _35923_ = _35344_ ^ _35925_ /*37824*/;
assign _35924_ = _35916_ & _35923_ /*37822*/;
assign _35793_ = _35916_ ^ _35923_ /*37823*/;
assign _35921_ = _35922_ | _35924_ /*37820*/;
assign _35930_ = ~D[17] /*37819*/;
assign _35927_ = _35345_ & _35930_ /*37815*/;
assign _35928_ = _35345_ ^ _35930_ /*37818*/;
assign _35929_ = _35921_ & _35928_ /*37816*/;
assign _35794_ = _35921_ ^ _35928_ /*37817*/;
assign _35926_ = _35927_ | _35929_ /*37814*/;
assign _35935_ = ~D[18] /*37813*/;
assign _35932_ = _35346_ & _35935_ /*37809*/;
assign _35933_ = _35346_ ^ _35935_ /*37812*/;
assign _35934_ = _35926_ & _35933_ /*37810*/;
assign _35795_ = _35926_ ^ _35933_ /*37811*/;
assign _35931_ = _35932_ | _35934_ /*37808*/;
assign _35940_ = ~D[19] /*37807*/;
assign _35937_ = _35347_ & _35940_ /*37803*/;
assign _35938_ = _35347_ ^ _35940_ /*37806*/;
assign _35939_ = _35931_ & _35938_ /*37804*/;
assign _35796_ = _35931_ ^ _35938_ /*37805*/;
assign _35936_ = _35937_ | _35939_ /*37802*/;
assign _35945_ = ~D[20] /*37801*/;
assign _35942_ = _35348_ & _35945_ /*37797*/;
assign _35943_ = _35348_ ^ _35945_ /*37800*/;
assign _35944_ = _35936_ & _35943_ /*37798*/;
assign _35797_ = _35936_ ^ _35943_ /*37799*/;
assign _35941_ = _35942_ | _35944_ /*37796*/;
assign _35950_ = ~D[21] /*37795*/;
assign _35947_ = _35349_ & _35950_ /*37791*/;
assign _35948_ = _35349_ ^ _35950_ /*37794*/;
assign _35949_ = _35941_ & _35948_ /*37792*/;
assign _35798_ = _35941_ ^ _35948_ /*37793*/;
assign _35946_ = _35947_ | _35949_ /*37790*/;
assign _35955_ = ~D[22] /*37789*/;
assign _35952_ = _35350_ & _35955_ /*37785*/;
assign _35953_ = _35350_ ^ _35955_ /*37788*/;
assign _35954_ = _35946_ & _35953_ /*37786*/;
assign _35799_ = _35946_ ^ _35953_ /*37787*/;
assign _35951_ = _35952_ | _35954_ /*37784*/;
assign _35960_ = ~D[23] /*37783*/;
assign _35957_ = _35351_ & _35960_ /*37779*/;
assign _35958_ = _35351_ ^ _35960_ /*37782*/;
assign _35959_ = _35951_ & _35958_ /*37780*/;
assign _35800_ = _35951_ ^ _35958_ /*37781*/;
assign _35956_ = _35957_ | _35959_ /*37778*/;
assign _35965_ = ~D[24] /*37777*/;
assign _35962_ = _35352_ & _35965_ /*37773*/;
assign _35963_ = _35352_ ^ _35965_ /*37776*/;
assign _35964_ = _35956_ & _35963_ /*37774*/;
assign _35801_ = _35956_ ^ _35963_ /*37775*/;
assign _35961_ = _35962_ | _35964_ /*37772*/;
assign _35970_ = ~D[25] /*37771*/;
assign _35967_ = _35353_ & _35970_ /*37767*/;
assign _35968_ = _35353_ ^ _35970_ /*37770*/;
assign _35969_ = _35961_ & _35968_ /*37768*/;
assign _35802_ = _35961_ ^ _35968_ /*37769*/;
assign _35966_ = _35967_ | _35969_ /*37766*/;
assign _35975_ = ~D[26] /*37765*/;
assign _35972_ = _35354_ & _35975_ /*37761*/;
assign _35973_ = _35354_ ^ _35975_ /*37764*/;
assign _35974_ = _35966_ & _35973_ /*37762*/;
assign _35803_ = _35966_ ^ _35973_ /*37763*/;
assign _35971_ = _35972_ | _35974_ /*37760*/;
assign _35980_ = ~D[27] /*37759*/;
assign _35977_ = _35355_ & _35980_ /*37755*/;
assign _35978_ = _35355_ ^ _35980_ /*37758*/;
assign _35979_ = _35971_ & _35978_ /*37756*/;
assign _35804_ = _35971_ ^ _35978_ /*37757*/;
assign _35976_ = _35977_ | _35979_ /*37754*/;
assign _35985_ = ~D[28] /*37753*/;
assign _35982_ = _35356_ & _35985_ /*37749*/;
assign _35983_ = _35356_ ^ _35985_ /*37752*/;
assign _35984_ = _35976_ & _35983_ /*37750*/;
assign _35805_ = _35976_ ^ _35983_ /*37751*/;
assign _35981_ = _35982_ | _35984_ /*37748*/;
assign _35990_ = ~D[29] /*37747*/;
assign _35987_ = _35357_ & _35990_ /*37743*/;
assign _35988_ = _35357_ ^ _35990_ /*37746*/;
assign _35989_ = _35981_ & _35988_ /*37744*/;
assign _35806_ = _35981_ ^ _35988_ /*37745*/;
assign _35986_ = _35987_ | _35989_ /*37742*/;
assign _35995_ = ~D[30] /*37741*/;
assign _35992_ = _35358_ & _35995_ /*37737*/;
assign _35993_ = _35358_ ^ _35995_ /*37740*/;
assign _35994_ = _35986_ & _35993_ /*37738*/;
assign _35807_ = _35986_ ^ _35993_ /*37739*/;
assign _35991_ = _35992_ | _35994_ /*37736*/;
assign _36000_ = ~D[31] /*37735*/;
assign _35997_ = _35359_ & _36000_ /*37731*/;
assign _35998_ = _35359_ ^ _36000_ /*37734*/;
assign _35999_ = _35991_ & _35998_ /*37732*/;
assign _35808_ = _35991_ ^ _35998_ /*37733*/;
assign _35996_ = _35997_ | _35999_ /*37730*/;
assign _36005_ = ~D[32] /*37729*/;
assign _36002_ = _35360_ & _36005_ /*37725*/;
assign _36003_ = _35360_ ^ _36005_ /*37728*/;
assign _36004_ = _35996_ & _36003_ /*37726*/;
assign _35809_ = _35996_ ^ _36003_ /*37727*/;
assign _36001_ = _36002_ | _36004_ /*37724*/;
assign _36010_ = ~D[33] /*37723*/;
assign _36007_ = _35361_ & _36010_ /*37719*/;
assign _36008_ = _35361_ ^ _36010_ /*37722*/;
assign _36009_ = _36001_ & _36008_ /*37720*/;
assign _35810_ = _36001_ ^ _36008_ /*37721*/;
assign _36006_ = _36007_ | _36009_ /*37718*/;
assign _36015_ = ~D[34] /*37717*/;
assign _36012_ = _35362_ & _36015_ /*37713*/;
assign _36013_ = _35362_ ^ _36015_ /*37716*/;
assign _36014_ = _36006_ & _36013_ /*37714*/;
assign _35811_ = _36006_ ^ _36013_ /*37715*/;
assign _36011_ = _36012_ | _36014_ /*37712*/;
assign _36020_ = ~D[35] /*37711*/;
assign _36017_ = _35363_ & _36020_ /*37707*/;
assign _36018_ = _35363_ ^ _36020_ /*37710*/;
assign _36019_ = _36011_ & _36018_ /*37708*/;
assign _35812_ = _36011_ ^ _36018_ /*37709*/;
assign _36016_ = _36017_ | _36019_ /*37706*/;
assign _36025_ = ~D[36] /*37705*/;
assign _36022_ = _35364_ & _36025_ /*37701*/;
assign _36023_ = _35364_ ^ _36025_ /*37704*/;
assign _36024_ = _36016_ & _36023_ /*37702*/;
assign _35813_ = _36016_ ^ _36023_ /*37703*/;
assign _36021_ = _36022_ | _36024_ /*37700*/;
assign _36030_ = ~D[37] /*37699*/;
assign _36027_ = _35365_ & _36030_ /*37695*/;
assign _36028_ = _35365_ ^ _36030_ /*37698*/;
assign _36029_ = _36021_ & _36028_ /*37696*/;
assign _35814_ = _36021_ ^ _36028_ /*37697*/;
assign _36026_ = _36027_ | _36029_ /*37694*/;
assign _36035_ = ~D[38] /*37693*/;
assign _36032_ = _35366_ & _36035_ /*37689*/;
assign _36033_ = _35366_ ^ _36035_ /*37692*/;
assign _36034_ = _36026_ & _36033_ /*37690*/;
assign _35815_ = _36026_ ^ _36033_ /*37691*/;
assign _36031_ = _36032_ | _36034_ /*37688*/;
assign _36040_ = ~D[39] /*37687*/;
assign _36037_ = _35367_ & _36040_ /*37683*/;
assign _36038_ = _35367_ ^ _36040_ /*37686*/;
assign _36039_ = _36031_ & _36038_ /*37684*/;
assign _35816_ = _36031_ ^ _36038_ /*37685*/;
assign _36036_ = _36037_ | _36039_ /*37682*/;
assign _36045_ = ~D[40] /*37681*/;
assign _36042_ = _35368_ & _36045_ /*37677*/;
assign _36043_ = _35368_ ^ _36045_ /*37680*/;
assign _36044_ = _36036_ & _36043_ /*37678*/;
assign _35817_ = _36036_ ^ _36043_ /*37679*/;
assign _36041_ = _36042_ | _36044_ /*37676*/;
assign _36050_ = ~D[41] /*37675*/;
assign _36047_ = _35369_ & _36050_ /*37671*/;
assign _36048_ = _35369_ ^ _36050_ /*37674*/;
assign _36049_ = _36041_ & _36048_ /*37672*/;
assign _35818_ = _36041_ ^ _36048_ /*37673*/;
assign _36046_ = _36047_ | _36049_ /*37670*/;
assign _36055_ = ~D[42] /*37669*/;
assign _36052_ = _35370_ & _36055_ /*37665*/;
assign _36053_ = _35370_ ^ _36055_ /*37668*/;
assign _36054_ = _36046_ & _36053_ /*37666*/;
assign _35819_ = _36046_ ^ _36053_ /*37667*/;
assign _36051_ = _36052_ | _36054_ /*37664*/;
assign _36060_ = ~D[43] /*37663*/;
assign _36057_ = _35371_ & _36060_ /*37659*/;
assign _36058_ = _35371_ ^ _36060_ /*37662*/;
assign _36059_ = _36051_ & _36058_ /*37660*/;
assign _35820_ = _36051_ ^ _36058_ /*37661*/;
assign _36056_ = _36057_ | _36059_ /*37658*/;
assign _36065_ = ~D[44] /*37657*/;
assign _36062_ = _35372_ & _36065_ /*37653*/;
assign _36063_ = _35372_ ^ _36065_ /*37656*/;
assign _36064_ = _36056_ & _36063_ /*37654*/;
assign _35821_ = _36056_ ^ _36063_ /*37655*/;
assign _36061_ = _36062_ | _36064_ /*37652*/;
assign _36070_ = ~D[45] /*37651*/;
assign _36067_ = _35373_ & _36070_ /*37647*/;
assign _36068_ = _35373_ ^ _36070_ /*37650*/;
assign _36069_ = _36061_ & _36068_ /*37648*/;
assign _35822_ = _36061_ ^ _36068_ /*37649*/;
assign _36066_ = _36067_ | _36069_ /*37646*/;
assign _36075_ = ~D[46] /*37645*/;
assign _36072_ = _35374_ & _36075_ /*37641*/;
assign _36073_ = _35374_ ^ _36075_ /*37644*/;
assign _36074_ = _36066_ & _36073_ /*37642*/;
assign _35823_ = _36066_ ^ _36073_ /*37643*/;
assign _36071_ = _36072_ | _36074_ /*37640*/;
assign _36080_ = ~D[47] /*37639*/;
assign _36077_ = _35375_ & _36080_ /*37635*/;
assign _36078_ = _35375_ ^ _36080_ /*37638*/;
assign _36079_ = _36071_ & _36078_ /*37636*/;
assign _35824_ = _36071_ ^ _36078_ /*37637*/;
assign _36076_ = _36077_ | _36079_ /*37634*/;
assign _36085_ = ~D[48] /*37633*/;
assign _36082_ = _35376_ & _36085_ /*37629*/;
assign _36083_ = _35376_ ^ _36085_ /*37632*/;
assign _36084_ = _36076_ & _36083_ /*37630*/;
assign _35825_ = _36076_ ^ _36083_ /*37631*/;
assign _36081_ = _36082_ | _36084_ /*37628*/;
assign _36090_ = ~D[49] /*37627*/;
assign _36087_ = _35377_ & _36090_ /*37623*/;
assign _36088_ = _35377_ ^ _36090_ /*37626*/;
assign _36089_ = _36081_ & _36088_ /*37624*/;
assign _35826_ = _36081_ ^ _36088_ /*37625*/;
assign _36086_ = _36087_ | _36089_ /*37622*/;
assign _36095_ = ~D[50] /*37621*/;
assign _36092_ = _35378_ & _36095_ /*37617*/;
assign _36093_ = _35378_ ^ _36095_ /*37620*/;
assign _36094_ = _36086_ & _36093_ /*37618*/;
assign _35827_ = _36086_ ^ _36093_ /*37619*/;
assign _36091_ = _36092_ | _36094_ /*37616*/;
assign _36100_ = ~D[51] /*37615*/;
assign _36097_ = _35379_ & _36100_ /*37611*/;
assign _36098_ = _35379_ ^ _36100_ /*37614*/;
assign _36099_ = _36091_ & _36098_ /*37612*/;
assign _35828_ = _36091_ ^ _36098_ /*37613*/;
assign _36096_ = _36097_ | _36099_ /*37610*/;
assign _36105_ = ~D[52] /*37609*/;
assign _36102_ = _35380_ & _36105_ /*37605*/;
assign _36103_ = _35380_ ^ _36105_ /*37608*/;
assign _36104_ = _36096_ & _36103_ /*37606*/;
assign _35829_ = _36096_ ^ _36103_ /*37607*/;
assign _36101_ = _36102_ | _36104_ /*37604*/;
assign _36110_ = ~D[53] /*37603*/;
assign _36107_ = _35381_ & _36110_ /*37599*/;
assign _36108_ = _35381_ ^ _36110_ /*37602*/;
assign _36109_ = _36101_ & _36108_ /*37600*/;
assign _35830_ = _36101_ ^ _36108_ /*37601*/;
assign _36106_ = _36107_ | _36109_ /*37598*/;
assign _36115_ = ~D[54] /*37597*/;
assign _36112_ = _35382_ & _36115_ /*37593*/;
assign _36113_ = _35382_ ^ _36115_ /*37596*/;
assign _36114_ = _36106_ & _36113_ /*37594*/;
assign _35831_ = _36106_ ^ _36113_ /*37595*/;
assign _36111_ = _36112_ | _36114_ /*37592*/;
assign _36120_ = ~D[55] /*37591*/;
assign _36117_ = _35383_ & _36120_ /*37587*/;
assign _36118_ = _35383_ ^ _36120_ /*37590*/;
assign _36119_ = _36111_ & _36118_ /*37588*/;
assign _35832_ = _36111_ ^ _36118_ /*37589*/;
assign _36116_ = _36117_ | _36119_ /*37586*/;
assign _36125_ = ~D[56] /*37585*/;
assign _36122_ = _35384_ & _36125_ /*37581*/;
assign _36123_ = _35384_ ^ _36125_ /*37584*/;
assign _36124_ = _36116_ & _36123_ /*37582*/;
assign _35833_ = _36116_ ^ _36123_ /*37583*/;
assign _36121_ = _36122_ | _36124_ /*37580*/;
assign _36130_ = ~D[57] /*37579*/;
assign _36127_ = _35385_ & _36130_ /*37575*/;
assign _36128_ = _35385_ ^ _36130_ /*37578*/;
assign _36129_ = _36121_ & _36128_ /*37576*/;
assign _35834_ = _36121_ ^ _36128_ /*37577*/;
assign _36126_ = _36127_ | _36129_ /*37574*/;
assign _36135_ = ~D[58] /*37573*/;
assign _36132_ = _35386_ & _36135_ /*37569*/;
assign _36133_ = _35386_ ^ _36135_ /*37572*/;
assign _36134_ = _36126_ & _36133_ /*37570*/;
assign _35835_ = _36126_ ^ _36133_ /*37571*/;
assign _36131_ = _36132_ | _36134_ /*37568*/;
assign _36140_ = ~D[59] /*37567*/;
assign _36137_ = _35387_ & _36140_ /*37563*/;
assign _36138_ = _35387_ ^ _36140_ /*37566*/;
assign _36139_ = _36131_ & _36138_ /*37564*/;
assign _35836_ = _36131_ ^ _36138_ /*37565*/;
assign _36136_ = _36137_ | _36139_ /*37562*/;
assign _36145_ = ~D[60] /*37561*/;
assign _36142_ = _35388_ & _36145_ /*37557*/;
assign _36143_ = _35388_ ^ _36145_ /*37560*/;
assign _36144_ = _36136_ & _36143_ /*37558*/;
assign _35837_ = _36136_ ^ _36143_ /*37559*/;
assign _36141_ = _36142_ | _36144_ /*37556*/;
assign _36150_ = ~D[61] /*37555*/;
assign _36147_ = _35389_ & _36150_ /*37551*/;
assign _36148_ = _35389_ ^ _36150_ /*37554*/;
assign _36149_ = _36141_ & _36148_ /*37552*/;
assign _35838_ = _36141_ ^ _36148_ /*37553*/;
assign _36146_ = _36147_ | _36149_ /*37550*/;
assign _36155_ = ~D[62] /*37549*/;
assign _36152_ = _35390_ & _36155_ /*37545*/;
assign _36153_ = _35390_ ^ _36155_ /*37548*/;
assign _36154_ = _36146_ & _36153_ /*37546*/;
assign _35839_ = _36146_ ^ _36153_ /*37547*/;
assign _36151_ = _36152_ | _36154_ /*37544*/;
assign _36156_ = _35391_ & oneWire /*37539*/;
assign _36157_ = _35391_ ^ oneWire /*37542*/;
assign _36158_ = _36151_ & _36157_ /*37540*/;
assign _35840_ = _36151_ ^ _36157_ /*37541*/;
assign Q[23] = _36156_ | _36158_ /*37538*/;
assign _36291_ = ~Q[23] /*37153*/;
assign _36290_ = _36291_ & D[0] /*37152*/;
assign _36293_ = _35777_ & _36290_ /*37147*/;
assign _36294_ = _35777_ ^ _36290_ /*37150*/;
assign _36295_ = zeroWire & _36294_ /*37148*/;
assign _36225_ = zeroWire ^ _36294_ /*37149*/;
assign _36292_ = _36293_ | _36295_ /*37146*/;
assign _36297_ = ~Q[23] /*37145*/;
assign _36296_ = _36297_ & D[1] /*37144*/;
assign _36299_ = _35778_ & _36296_ /*37139*/;
assign _36300_ = _35778_ ^ _36296_ /*37142*/;
assign _36301_ = _36292_ & _36300_ /*37140*/;
assign _36226_ = _36292_ ^ _36300_ /*37141*/;
assign _36298_ = _36299_ | _36301_ /*37138*/;
assign _36303_ = ~Q[23] /*37137*/;
assign _36302_ = _36303_ & D[2] /*37136*/;
assign _36305_ = _35779_ & _36302_ /*37131*/;
assign _36306_ = _35779_ ^ _36302_ /*37134*/;
assign _36307_ = _36298_ & _36306_ /*37132*/;
assign _36227_ = _36298_ ^ _36306_ /*37133*/;
assign _36304_ = _36305_ | _36307_ /*37130*/;
assign _36309_ = ~Q[23] /*37129*/;
assign _36308_ = _36309_ & D[3] /*37128*/;
assign _36311_ = _35780_ & _36308_ /*37123*/;
assign _36312_ = _35780_ ^ _36308_ /*37126*/;
assign _36313_ = _36304_ & _36312_ /*37124*/;
assign _36228_ = _36304_ ^ _36312_ /*37125*/;
assign _36310_ = _36311_ | _36313_ /*37122*/;
assign _36315_ = ~Q[23] /*37121*/;
assign _36314_ = _36315_ & D[4] /*37120*/;
assign _36317_ = _35781_ & _36314_ /*37115*/;
assign _36318_ = _35781_ ^ _36314_ /*37118*/;
assign _36319_ = _36310_ & _36318_ /*37116*/;
assign _36229_ = _36310_ ^ _36318_ /*37117*/;
assign _36316_ = _36317_ | _36319_ /*37114*/;
assign _36321_ = ~Q[23] /*37113*/;
assign _36320_ = _36321_ & D[5] /*37112*/;
assign _36323_ = _35782_ & _36320_ /*37107*/;
assign _36324_ = _35782_ ^ _36320_ /*37110*/;
assign _36325_ = _36316_ & _36324_ /*37108*/;
assign _36230_ = _36316_ ^ _36324_ /*37109*/;
assign _36322_ = _36323_ | _36325_ /*37106*/;
assign _36327_ = ~Q[23] /*37105*/;
assign _36326_ = _36327_ & D[6] /*37104*/;
assign _36329_ = _35783_ & _36326_ /*37099*/;
assign _36330_ = _35783_ ^ _36326_ /*37102*/;
assign _36331_ = _36322_ & _36330_ /*37100*/;
assign _36231_ = _36322_ ^ _36330_ /*37101*/;
assign _36328_ = _36329_ | _36331_ /*37098*/;
assign _36333_ = ~Q[23] /*37097*/;
assign _36332_ = _36333_ & D[7] /*37096*/;
assign _36335_ = _35784_ & _36332_ /*37091*/;
assign _36336_ = _35784_ ^ _36332_ /*37094*/;
assign _36337_ = _36328_ & _36336_ /*37092*/;
assign _36232_ = _36328_ ^ _36336_ /*37093*/;
assign _36334_ = _36335_ | _36337_ /*37090*/;
assign _36339_ = ~Q[23] /*37089*/;
assign _36338_ = _36339_ & D[8] /*37088*/;
assign _36341_ = _35785_ & _36338_ /*37083*/;
assign _36342_ = _35785_ ^ _36338_ /*37086*/;
assign _36343_ = _36334_ & _36342_ /*37084*/;
assign _36233_ = _36334_ ^ _36342_ /*37085*/;
assign _36340_ = _36341_ | _36343_ /*37082*/;
assign _36345_ = ~Q[23] /*37081*/;
assign _36344_ = _36345_ & D[9] /*37080*/;
assign _36347_ = _35786_ & _36344_ /*37075*/;
assign _36348_ = _35786_ ^ _36344_ /*37078*/;
assign _36349_ = _36340_ & _36348_ /*37076*/;
assign _36234_ = _36340_ ^ _36348_ /*37077*/;
assign _36346_ = _36347_ | _36349_ /*37074*/;
assign _36351_ = ~Q[23] /*37073*/;
assign _36350_ = _36351_ & D[10] /*37072*/;
assign _36353_ = _35787_ & _36350_ /*37067*/;
assign _36354_ = _35787_ ^ _36350_ /*37070*/;
assign _36355_ = _36346_ & _36354_ /*37068*/;
assign _36235_ = _36346_ ^ _36354_ /*37069*/;
assign _36352_ = _36353_ | _36355_ /*37066*/;
assign _36357_ = ~Q[23] /*37065*/;
assign _36356_ = _36357_ & D[11] /*37064*/;
assign _36359_ = _35788_ & _36356_ /*37059*/;
assign _36360_ = _35788_ ^ _36356_ /*37062*/;
assign _36361_ = _36352_ & _36360_ /*37060*/;
assign _36236_ = _36352_ ^ _36360_ /*37061*/;
assign _36358_ = _36359_ | _36361_ /*37058*/;
assign _36363_ = ~Q[23] /*37057*/;
assign _36362_ = _36363_ & D[12] /*37056*/;
assign _36365_ = _35789_ & _36362_ /*37051*/;
assign _36366_ = _35789_ ^ _36362_ /*37054*/;
assign _36367_ = _36358_ & _36366_ /*37052*/;
assign _36237_ = _36358_ ^ _36366_ /*37053*/;
assign _36364_ = _36365_ | _36367_ /*37050*/;
assign _36369_ = ~Q[23] /*37049*/;
assign _36368_ = _36369_ & D[13] /*37048*/;
assign _36371_ = _35790_ & _36368_ /*37043*/;
assign _36372_ = _35790_ ^ _36368_ /*37046*/;
assign _36373_ = _36364_ & _36372_ /*37044*/;
assign _36238_ = _36364_ ^ _36372_ /*37045*/;
assign _36370_ = _36371_ | _36373_ /*37042*/;
assign _36375_ = ~Q[23] /*37041*/;
assign _36374_ = _36375_ & D[14] /*37040*/;
assign _36377_ = _35791_ & _36374_ /*37035*/;
assign _36378_ = _35791_ ^ _36374_ /*37038*/;
assign _36379_ = _36370_ & _36378_ /*37036*/;
assign _36239_ = _36370_ ^ _36378_ /*37037*/;
assign _36376_ = _36377_ | _36379_ /*37034*/;
assign _36381_ = ~Q[23] /*37033*/;
assign _36380_ = _36381_ & D[15] /*37032*/;
assign _36383_ = _35792_ & _36380_ /*37027*/;
assign _36384_ = _35792_ ^ _36380_ /*37030*/;
assign _36385_ = _36376_ & _36384_ /*37028*/;
assign _36240_ = _36376_ ^ _36384_ /*37029*/;
assign _36382_ = _36383_ | _36385_ /*37026*/;
assign _36387_ = ~Q[23] /*37025*/;
assign _36386_ = _36387_ & D[16] /*37024*/;
assign _36389_ = _35793_ & _36386_ /*37019*/;
assign _36390_ = _35793_ ^ _36386_ /*37022*/;
assign _36391_ = _36382_ & _36390_ /*37020*/;
assign _36241_ = _36382_ ^ _36390_ /*37021*/;
assign _36388_ = _36389_ | _36391_ /*37018*/;
assign _36393_ = ~Q[23] /*37017*/;
assign _36392_ = _36393_ & D[17] /*37016*/;
assign _36395_ = _35794_ & _36392_ /*37011*/;
assign _36396_ = _35794_ ^ _36392_ /*37014*/;
assign _36397_ = _36388_ & _36396_ /*37012*/;
assign _36242_ = _36388_ ^ _36396_ /*37013*/;
assign _36394_ = _36395_ | _36397_ /*37010*/;
assign _36399_ = ~Q[23] /*37009*/;
assign _36398_ = _36399_ & D[18] /*37008*/;
assign _36401_ = _35795_ & _36398_ /*37003*/;
assign _36402_ = _35795_ ^ _36398_ /*37006*/;
assign _36403_ = _36394_ & _36402_ /*37004*/;
assign _36243_ = _36394_ ^ _36402_ /*37005*/;
assign _36400_ = _36401_ | _36403_ /*37002*/;
assign _36405_ = ~Q[23] /*37001*/;
assign _36404_ = _36405_ & D[19] /*37000*/;
assign _36407_ = _35796_ & _36404_ /*36995*/;
assign _36408_ = _35796_ ^ _36404_ /*36998*/;
assign _36409_ = _36400_ & _36408_ /*36996*/;
assign _36244_ = _36400_ ^ _36408_ /*36997*/;
assign _36406_ = _36407_ | _36409_ /*36994*/;
assign _36411_ = ~Q[23] /*36993*/;
assign _36410_ = _36411_ & D[20] /*36992*/;
assign _36413_ = _35797_ & _36410_ /*36987*/;
assign _36414_ = _35797_ ^ _36410_ /*36990*/;
assign _36415_ = _36406_ & _36414_ /*36988*/;
assign _36245_ = _36406_ ^ _36414_ /*36989*/;
assign _36412_ = _36413_ | _36415_ /*36986*/;
assign _36417_ = ~Q[23] /*36985*/;
assign _36416_ = _36417_ & D[21] /*36984*/;
assign _36419_ = _35798_ & _36416_ /*36979*/;
assign _36420_ = _35798_ ^ _36416_ /*36982*/;
assign _36421_ = _36412_ & _36420_ /*36980*/;
assign _36246_ = _36412_ ^ _36420_ /*36981*/;
assign _36418_ = _36419_ | _36421_ /*36978*/;
assign _36423_ = ~Q[23] /*36977*/;
assign _36422_ = _36423_ & D[22] /*36976*/;
assign _36425_ = _35799_ & _36422_ /*36971*/;
assign _36426_ = _35799_ ^ _36422_ /*36974*/;
assign _36427_ = _36418_ & _36426_ /*36972*/;
assign _36247_ = _36418_ ^ _36426_ /*36973*/;
assign _36424_ = _36425_ | _36427_ /*36970*/;
assign _36429_ = ~Q[23] /*36969*/;
assign _36428_ = _36429_ & D[23] /*36968*/;
assign _36431_ = _35800_ & _36428_ /*36963*/;
assign _36432_ = _35800_ ^ _36428_ /*36966*/;
assign _36433_ = _36424_ & _36432_ /*36964*/;
assign _36248_ = _36424_ ^ _36432_ /*36965*/;
assign _36430_ = _36431_ | _36433_ /*36962*/;
assign _36435_ = ~Q[23] /*36961*/;
assign _36434_ = _36435_ & D[24] /*36960*/;
assign _36437_ = _35801_ & _36434_ /*36955*/;
assign _36438_ = _35801_ ^ _36434_ /*36958*/;
assign _36439_ = _36430_ & _36438_ /*36956*/;
assign _36249_ = _36430_ ^ _36438_ /*36957*/;
assign _36436_ = _36437_ | _36439_ /*36954*/;
assign _36441_ = ~Q[23] /*36953*/;
assign _36440_ = _36441_ & D[25] /*36952*/;
assign _36443_ = _35802_ & _36440_ /*36947*/;
assign _36444_ = _35802_ ^ _36440_ /*36950*/;
assign _36445_ = _36436_ & _36444_ /*36948*/;
assign _36250_ = _36436_ ^ _36444_ /*36949*/;
assign _36442_ = _36443_ | _36445_ /*36946*/;
assign _36447_ = ~Q[23] /*36945*/;
assign _36446_ = _36447_ & D[26] /*36944*/;
assign _36449_ = _35803_ & _36446_ /*36939*/;
assign _36450_ = _35803_ ^ _36446_ /*36942*/;
assign _36451_ = _36442_ & _36450_ /*36940*/;
assign _36251_ = _36442_ ^ _36450_ /*36941*/;
assign _36448_ = _36449_ | _36451_ /*36938*/;
assign _36453_ = ~Q[23] /*36937*/;
assign _36452_ = _36453_ & D[27] /*36936*/;
assign _36455_ = _35804_ & _36452_ /*36931*/;
assign _36456_ = _35804_ ^ _36452_ /*36934*/;
assign _36457_ = _36448_ & _36456_ /*36932*/;
assign _36252_ = _36448_ ^ _36456_ /*36933*/;
assign _36454_ = _36455_ | _36457_ /*36930*/;
assign _36459_ = ~Q[23] /*36929*/;
assign _36458_ = _36459_ & D[28] /*36928*/;
assign _36461_ = _35805_ & _36458_ /*36923*/;
assign _36462_ = _35805_ ^ _36458_ /*36926*/;
assign _36463_ = _36454_ & _36462_ /*36924*/;
assign _36253_ = _36454_ ^ _36462_ /*36925*/;
assign _36460_ = _36461_ | _36463_ /*36922*/;
assign _36465_ = ~Q[23] /*36921*/;
assign _36464_ = _36465_ & D[29] /*36920*/;
assign _36467_ = _35806_ & _36464_ /*36915*/;
assign _36468_ = _35806_ ^ _36464_ /*36918*/;
assign _36469_ = _36460_ & _36468_ /*36916*/;
assign _36254_ = _36460_ ^ _36468_ /*36917*/;
assign _36466_ = _36467_ | _36469_ /*36914*/;
assign _36471_ = ~Q[23] /*36913*/;
assign _36470_ = _36471_ & D[30] /*36912*/;
assign _36473_ = _35807_ & _36470_ /*36907*/;
assign _36474_ = _35807_ ^ _36470_ /*36910*/;
assign _36475_ = _36466_ & _36474_ /*36908*/;
assign _36255_ = _36466_ ^ _36474_ /*36909*/;
assign _36472_ = _36473_ | _36475_ /*36906*/;
assign _36477_ = ~Q[23] /*36905*/;
assign _36476_ = _36477_ & D[31] /*36904*/;
assign _36479_ = _35808_ & _36476_ /*36899*/;
assign _36480_ = _35808_ ^ _36476_ /*36902*/;
assign _36481_ = _36472_ & _36480_ /*36900*/;
assign _36256_ = _36472_ ^ _36480_ /*36901*/;
assign _36478_ = _36479_ | _36481_ /*36898*/;
assign _36483_ = ~Q[23] /*36897*/;
assign _36482_ = _36483_ & D[32] /*36896*/;
assign _36485_ = _35809_ & _36482_ /*36891*/;
assign _36486_ = _35809_ ^ _36482_ /*36894*/;
assign _36487_ = _36478_ & _36486_ /*36892*/;
assign _36257_ = _36478_ ^ _36486_ /*36893*/;
assign _36484_ = _36485_ | _36487_ /*36890*/;
assign _36489_ = ~Q[23] /*36889*/;
assign _36488_ = _36489_ & D[33] /*36888*/;
assign _36491_ = _35810_ & _36488_ /*36883*/;
assign _36492_ = _35810_ ^ _36488_ /*36886*/;
assign _36493_ = _36484_ & _36492_ /*36884*/;
assign _36258_ = _36484_ ^ _36492_ /*36885*/;
assign _36490_ = _36491_ | _36493_ /*36882*/;
assign _36495_ = ~Q[23] /*36881*/;
assign _36494_ = _36495_ & D[34] /*36880*/;
assign _36497_ = _35811_ & _36494_ /*36875*/;
assign _36498_ = _35811_ ^ _36494_ /*36878*/;
assign _36499_ = _36490_ & _36498_ /*36876*/;
assign _36259_ = _36490_ ^ _36498_ /*36877*/;
assign _36496_ = _36497_ | _36499_ /*36874*/;
assign _36501_ = ~Q[23] /*36873*/;
assign _36500_ = _36501_ & D[35] /*36872*/;
assign _36503_ = _35812_ & _36500_ /*36867*/;
assign _36504_ = _35812_ ^ _36500_ /*36870*/;
assign _36505_ = _36496_ & _36504_ /*36868*/;
assign _36260_ = _36496_ ^ _36504_ /*36869*/;
assign _36502_ = _36503_ | _36505_ /*36866*/;
assign _36507_ = ~Q[23] /*36865*/;
assign _36506_ = _36507_ & D[36] /*36864*/;
assign _36509_ = _35813_ & _36506_ /*36859*/;
assign _36510_ = _35813_ ^ _36506_ /*36862*/;
assign _36511_ = _36502_ & _36510_ /*36860*/;
assign _36261_ = _36502_ ^ _36510_ /*36861*/;
assign _36508_ = _36509_ | _36511_ /*36858*/;
assign _36513_ = ~Q[23] /*36857*/;
assign _36512_ = _36513_ & D[37] /*36856*/;
assign _36515_ = _35814_ & _36512_ /*36851*/;
assign _36516_ = _35814_ ^ _36512_ /*36854*/;
assign _36517_ = _36508_ & _36516_ /*36852*/;
assign _36262_ = _36508_ ^ _36516_ /*36853*/;
assign _36514_ = _36515_ | _36517_ /*36850*/;
assign _36519_ = ~Q[23] /*36849*/;
assign _36518_ = _36519_ & D[38] /*36848*/;
assign _36521_ = _35815_ & _36518_ /*36843*/;
assign _36522_ = _35815_ ^ _36518_ /*36846*/;
assign _36523_ = _36514_ & _36522_ /*36844*/;
assign _36263_ = _36514_ ^ _36522_ /*36845*/;
assign _36520_ = _36521_ | _36523_ /*36842*/;
assign _36525_ = ~Q[23] /*36841*/;
assign _36524_ = _36525_ & D[39] /*36840*/;
assign _36527_ = _35816_ & _36524_ /*36835*/;
assign _36528_ = _35816_ ^ _36524_ /*36838*/;
assign _36529_ = _36520_ & _36528_ /*36836*/;
assign _36264_ = _36520_ ^ _36528_ /*36837*/;
assign _36526_ = _36527_ | _36529_ /*36834*/;
assign _36531_ = ~Q[23] /*36833*/;
assign _36530_ = _36531_ & D[40] /*36832*/;
assign _36533_ = _35817_ & _36530_ /*36827*/;
assign _36534_ = _35817_ ^ _36530_ /*36830*/;
assign _36535_ = _36526_ & _36534_ /*36828*/;
assign _36265_ = _36526_ ^ _36534_ /*36829*/;
assign _36532_ = _36533_ | _36535_ /*36826*/;
assign _36537_ = ~Q[23] /*36825*/;
assign _36536_ = _36537_ & D[41] /*36824*/;
assign _36539_ = _35818_ & _36536_ /*36819*/;
assign _36540_ = _35818_ ^ _36536_ /*36822*/;
assign _36541_ = _36532_ & _36540_ /*36820*/;
assign _36266_ = _36532_ ^ _36540_ /*36821*/;
assign _36538_ = _36539_ | _36541_ /*36818*/;
assign _36543_ = ~Q[23] /*36817*/;
assign _36542_ = _36543_ & D[42] /*36816*/;
assign _36545_ = _35819_ & _36542_ /*36811*/;
assign _36546_ = _35819_ ^ _36542_ /*36814*/;
assign _36547_ = _36538_ & _36546_ /*36812*/;
assign _36267_ = _36538_ ^ _36546_ /*36813*/;
assign _36544_ = _36545_ | _36547_ /*36810*/;
assign _36549_ = ~Q[23] /*36809*/;
assign _36548_ = _36549_ & D[43] /*36808*/;
assign _36551_ = _35820_ & _36548_ /*36803*/;
assign _36552_ = _35820_ ^ _36548_ /*36806*/;
assign _36553_ = _36544_ & _36552_ /*36804*/;
assign _36268_ = _36544_ ^ _36552_ /*36805*/;
assign _36550_ = _36551_ | _36553_ /*36802*/;
assign _36555_ = ~Q[23] /*36801*/;
assign _36554_ = _36555_ & D[44] /*36800*/;
assign _36557_ = _35821_ & _36554_ /*36795*/;
assign _36558_ = _35821_ ^ _36554_ /*36798*/;
assign _36559_ = _36550_ & _36558_ /*36796*/;
assign _36269_ = _36550_ ^ _36558_ /*36797*/;
assign _36556_ = _36557_ | _36559_ /*36794*/;
assign _36561_ = ~Q[23] /*36793*/;
assign _36560_ = _36561_ & D[45] /*36792*/;
assign _36563_ = _35822_ & _36560_ /*36787*/;
assign _36564_ = _35822_ ^ _36560_ /*36790*/;
assign _36565_ = _36556_ & _36564_ /*36788*/;
assign _36270_ = _36556_ ^ _36564_ /*36789*/;
assign _36562_ = _36563_ | _36565_ /*36786*/;
assign _36567_ = ~Q[23] /*36785*/;
assign _36566_ = _36567_ & D[46] /*36784*/;
assign _36569_ = _35823_ & _36566_ /*36779*/;
assign _36570_ = _35823_ ^ _36566_ /*36782*/;
assign _36571_ = _36562_ & _36570_ /*36780*/;
assign _36271_ = _36562_ ^ _36570_ /*36781*/;
assign _36568_ = _36569_ | _36571_ /*36778*/;
assign _36573_ = ~Q[23] /*36777*/;
assign _36572_ = _36573_ & D[47] /*36776*/;
assign _36575_ = _35824_ & _36572_ /*36771*/;
assign _36576_ = _35824_ ^ _36572_ /*36774*/;
assign _36577_ = _36568_ & _36576_ /*36772*/;
assign _36272_ = _36568_ ^ _36576_ /*36773*/;
assign _36574_ = _36575_ | _36577_ /*36770*/;
assign _36579_ = ~Q[23] /*36769*/;
assign _36578_ = _36579_ & D[48] /*36768*/;
assign _36581_ = _35825_ & _36578_ /*36763*/;
assign _36582_ = _35825_ ^ _36578_ /*36766*/;
assign _36583_ = _36574_ & _36582_ /*36764*/;
assign _36273_ = _36574_ ^ _36582_ /*36765*/;
assign _36580_ = _36581_ | _36583_ /*36762*/;
assign _36585_ = ~Q[23] /*36761*/;
assign _36584_ = _36585_ & D[49] /*36760*/;
assign _36587_ = _35826_ & _36584_ /*36755*/;
assign _36588_ = _35826_ ^ _36584_ /*36758*/;
assign _36589_ = _36580_ & _36588_ /*36756*/;
assign _36274_ = _36580_ ^ _36588_ /*36757*/;
assign _36586_ = _36587_ | _36589_ /*36754*/;
assign _36591_ = ~Q[23] /*36753*/;
assign _36590_ = _36591_ & D[50] /*36752*/;
assign _36593_ = _35827_ & _36590_ /*36747*/;
assign _36594_ = _35827_ ^ _36590_ /*36750*/;
assign _36595_ = _36586_ & _36594_ /*36748*/;
assign _36275_ = _36586_ ^ _36594_ /*36749*/;
assign _36592_ = _36593_ | _36595_ /*36746*/;
assign _36597_ = ~Q[23] /*36745*/;
assign _36596_ = _36597_ & D[51] /*36744*/;
assign _36599_ = _35828_ & _36596_ /*36739*/;
assign _36600_ = _35828_ ^ _36596_ /*36742*/;
assign _36601_ = _36592_ & _36600_ /*36740*/;
assign _36276_ = _36592_ ^ _36600_ /*36741*/;
assign _36598_ = _36599_ | _36601_ /*36738*/;
assign _36603_ = ~Q[23] /*36737*/;
assign _36602_ = _36603_ & D[52] /*36736*/;
assign _36605_ = _35829_ & _36602_ /*36731*/;
assign _36606_ = _35829_ ^ _36602_ /*36734*/;
assign _36607_ = _36598_ & _36606_ /*36732*/;
assign _36277_ = _36598_ ^ _36606_ /*36733*/;
assign _36604_ = _36605_ | _36607_ /*36730*/;
assign _36609_ = ~Q[23] /*36729*/;
assign _36608_ = _36609_ & D[53] /*36728*/;
assign _36611_ = _35830_ & _36608_ /*36723*/;
assign _36612_ = _35830_ ^ _36608_ /*36726*/;
assign _36613_ = _36604_ & _36612_ /*36724*/;
assign _36278_ = _36604_ ^ _36612_ /*36725*/;
assign _36610_ = _36611_ | _36613_ /*36722*/;
assign _36615_ = ~Q[23] /*36721*/;
assign _36614_ = _36615_ & D[54] /*36720*/;
assign _36617_ = _35831_ & _36614_ /*36715*/;
assign _36618_ = _35831_ ^ _36614_ /*36718*/;
assign _36619_ = _36610_ & _36618_ /*36716*/;
assign _36279_ = _36610_ ^ _36618_ /*36717*/;
assign _36616_ = _36617_ | _36619_ /*36714*/;
assign _36621_ = ~Q[23] /*36713*/;
assign _36620_ = _36621_ & D[55] /*36712*/;
assign _36623_ = _35832_ & _36620_ /*36707*/;
assign _36624_ = _35832_ ^ _36620_ /*36710*/;
assign _36625_ = _36616_ & _36624_ /*36708*/;
assign _36280_ = _36616_ ^ _36624_ /*36709*/;
assign _36622_ = _36623_ | _36625_ /*36706*/;
assign _36627_ = ~Q[23] /*36705*/;
assign _36626_ = _36627_ & D[56] /*36704*/;
assign _36629_ = _35833_ & _36626_ /*36699*/;
assign _36630_ = _35833_ ^ _36626_ /*36702*/;
assign _36631_ = _36622_ & _36630_ /*36700*/;
assign _36281_ = _36622_ ^ _36630_ /*36701*/;
assign _36628_ = _36629_ | _36631_ /*36698*/;
assign _36633_ = ~Q[23] /*36697*/;
assign _36632_ = _36633_ & D[57] /*36696*/;
assign _36635_ = _35834_ & _36632_ /*36691*/;
assign _36636_ = _35834_ ^ _36632_ /*36694*/;
assign _36637_ = _36628_ & _36636_ /*36692*/;
assign _36282_ = _36628_ ^ _36636_ /*36693*/;
assign _36634_ = _36635_ | _36637_ /*36690*/;
assign _36639_ = ~Q[23] /*36689*/;
assign _36638_ = _36639_ & D[58] /*36688*/;
assign _36641_ = _35835_ & _36638_ /*36683*/;
assign _36642_ = _35835_ ^ _36638_ /*36686*/;
assign _36643_ = _36634_ & _36642_ /*36684*/;
assign _36283_ = _36634_ ^ _36642_ /*36685*/;
assign _36640_ = _36641_ | _36643_ /*36682*/;
assign _36645_ = ~Q[23] /*36681*/;
assign _36644_ = _36645_ & D[59] /*36680*/;
assign _36647_ = _35836_ & _36644_ /*36675*/;
assign _36648_ = _35836_ ^ _36644_ /*36678*/;
assign _36649_ = _36640_ & _36648_ /*36676*/;
assign _36284_ = _36640_ ^ _36648_ /*36677*/;
assign _36646_ = _36647_ | _36649_ /*36674*/;
assign _36651_ = ~Q[23] /*36673*/;
assign _36650_ = _36651_ & D[60] /*36672*/;
assign _36653_ = _35837_ & _36650_ /*36667*/;
assign _36654_ = _35837_ ^ _36650_ /*36670*/;
assign _36655_ = _36646_ & _36654_ /*36668*/;
assign _36285_ = _36646_ ^ _36654_ /*36669*/;
assign _36652_ = _36653_ | _36655_ /*36666*/;
assign _36657_ = ~Q[23] /*36665*/;
assign _36656_ = _36657_ & D[61] /*36664*/;
assign _36659_ = _35838_ & _36656_ /*36659*/;
assign _36660_ = _35838_ ^ _36656_ /*36662*/;
assign _36661_ = _36652_ & _36660_ /*36660*/;
assign _36286_ = _36652_ ^ _36660_ /*36661*/;
assign _36658_ = _36659_ | _36661_ /*36658*/;
assign _36663_ = ~Q[23] /*36657*/;
assign _36662_ = _36663_ & D[62] /*36656*/;
assign _36665_ = _35839_ & _36662_ /*36651*/;
assign _36666_ = _35839_ ^ _36662_ /*36654*/;
assign _36667_ = _36658_ & _36666_ /*36652*/;
assign _36287_ = _36658_ ^ _36666_ /*36653*/;
assign _36664_ = _36665_ | _36667_ /*36650*/;
assign _36669_ = ~Q[23] /*36649*/;
assign _36668_ = _36669_ & zeroWire /*36648*/;
assign _36670_ = _35840_ ^ _36668_ /*36646*/;
assign _36288_ = _36670_ ^ _36664_ /*36645*/;
assign _36741_ = ~D[0] /*36391*/;
assign _36738_ = R_0[22] & _36741_ /*36387*/;
assign _36739_ = R_0[22] ^ _36741_ /*36390*/;
assign _36740_ = oneWire & _36739_ /*36388*/;
assign _36673_ = oneWire ^ _36739_ /*36389*/;
assign _36737_ = _36738_ | _36740_ /*36386*/;
assign _36746_ = ~D[1] /*36385*/;
assign _36743_ = _36225_ & _36746_ /*36381*/;
assign _36744_ = _36225_ ^ _36746_ /*36384*/;
assign _36745_ = _36737_ & _36744_ /*36382*/;
assign _36674_ = _36737_ ^ _36744_ /*36383*/;
assign _36742_ = _36743_ | _36745_ /*36380*/;
assign _36751_ = ~D[2] /*36379*/;
assign _36748_ = _36226_ & _36751_ /*36375*/;
assign _36749_ = _36226_ ^ _36751_ /*36378*/;
assign _36750_ = _36742_ & _36749_ /*36376*/;
assign _36675_ = _36742_ ^ _36749_ /*36377*/;
assign _36747_ = _36748_ | _36750_ /*36374*/;
assign _36756_ = ~D[3] /*36373*/;
assign _36753_ = _36227_ & _36756_ /*36369*/;
assign _36754_ = _36227_ ^ _36756_ /*36372*/;
assign _36755_ = _36747_ & _36754_ /*36370*/;
assign _36676_ = _36747_ ^ _36754_ /*36371*/;
assign _36752_ = _36753_ | _36755_ /*36368*/;
assign _36761_ = ~D[4] /*36367*/;
assign _36758_ = _36228_ & _36761_ /*36363*/;
assign _36759_ = _36228_ ^ _36761_ /*36366*/;
assign _36760_ = _36752_ & _36759_ /*36364*/;
assign _36677_ = _36752_ ^ _36759_ /*36365*/;
assign _36757_ = _36758_ | _36760_ /*36362*/;
assign _36766_ = ~D[5] /*36361*/;
assign _36763_ = _36229_ & _36766_ /*36357*/;
assign _36764_ = _36229_ ^ _36766_ /*36360*/;
assign _36765_ = _36757_ & _36764_ /*36358*/;
assign _36678_ = _36757_ ^ _36764_ /*36359*/;
assign _36762_ = _36763_ | _36765_ /*36356*/;
assign _36771_ = ~D[6] /*36355*/;
assign _36768_ = _36230_ & _36771_ /*36351*/;
assign _36769_ = _36230_ ^ _36771_ /*36354*/;
assign _36770_ = _36762_ & _36769_ /*36352*/;
assign _36679_ = _36762_ ^ _36769_ /*36353*/;
assign _36767_ = _36768_ | _36770_ /*36350*/;
assign _36776_ = ~D[7] /*36349*/;
assign _36773_ = _36231_ & _36776_ /*36345*/;
assign _36774_ = _36231_ ^ _36776_ /*36348*/;
assign _36775_ = _36767_ & _36774_ /*36346*/;
assign _36680_ = _36767_ ^ _36774_ /*36347*/;
assign _36772_ = _36773_ | _36775_ /*36344*/;
assign _36781_ = ~D[8] /*36343*/;
assign _36778_ = _36232_ & _36781_ /*36339*/;
assign _36779_ = _36232_ ^ _36781_ /*36342*/;
assign _36780_ = _36772_ & _36779_ /*36340*/;
assign _36681_ = _36772_ ^ _36779_ /*36341*/;
assign _36777_ = _36778_ | _36780_ /*36338*/;
assign _36786_ = ~D[9] /*36337*/;
assign _36783_ = _36233_ & _36786_ /*36333*/;
assign _36784_ = _36233_ ^ _36786_ /*36336*/;
assign _36785_ = _36777_ & _36784_ /*36334*/;
assign _36682_ = _36777_ ^ _36784_ /*36335*/;
assign _36782_ = _36783_ | _36785_ /*36332*/;
assign _36791_ = ~D[10] /*36331*/;
assign _36788_ = _36234_ & _36791_ /*36327*/;
assign _36789_ = _36234_ ^ _36791_ /*36330*/;
assign _36790_ = _36782_ & _36789_ /*36328*/;
assign _36683_ = _36782_ ^ _36789_ /*36329*/;
assign _36787_ = _36788_ | _36790_ /*36326*/;
assign _36796_ = ~D[11] /*36325*/;
assign _36793_ = _36235_ & _36796_ /*36321*/;
assign _36794_ = _36235_ ^ _36796_ /*36324*/;
assign _36795_ = _36787_ & _36794_ /*36322*/;
assign _36684_ = _36787_ ^ _36794_ /*36323*/;
assign _36792_ = _36793_ | _36795_ /*36320*/;
assign _36801_ = ~D[12] /*36319*/;
assign _36798_ = _36236_ & _36801_ /*36315*/;
assign _36799_ = _36236_ ^ _36801_ /*36318*/;
assign _36800_ = _36792_ & _36799_ /*36316*/;
assign _36685_ = _36792_ ^ _36799_ /*36317*/;
assign _36797_ = _36798_ | _36800_ /*36314*/;
assign _36806_ = ~D[13] /*36313*/;
assign _36803_ = _36237_ & _36806_ /*36309*/;
assign _36804_ = _36237_ ^ _36806_ /*36312*/;
assign _36805_ = _36797_ & _36804_ /*36310*/;
assign _36686_ = _36797_ ^ _36804_ /*36311*/;
assign _36802_ = _36803_ | _36805_ /*36308*/;
assign _36811_ = ~D[14] /*36307*/;
assign _36808_ = _36238_ & _36811_ /*36303*/;
assign _36809_ = _36238_ ^ _36811_ /*36306*/;
assign _36810_ = _36802_ & _36809_ /*36304*/;
assign _36687_ = _36802_ ^ _36809_ /*36305*/;
assign _36807_ = _36808_ | _36810_ /*36302*/;
assign _36816_ = ~D[15] /*36301*/;
assign _36813_ = _36239_ & _36816_ /*36297*/;
assign _36814_ = _36239_ ^ _36816_ /*36300*/;
assign _36815_ = _36807_ & _36814_ /*36298*/;
assign _36688_ = _36807_ ^ _36814_ /*36299*/;
assign _36812_ = _36813_ | _36815_ /*36296*/;
assign _36821_ = ~D[16] /*36295*/;
assign _36818_ = _36240_ & _36821_ /*36291*/;
assign _36819_ = _36240_ ^ _36821_ /*36294*/;
assign _36820_ = _36812_ & _36819_ /*36292*/;
assign _36689_ = _36812_ ^ _36819_ /*36293*/;
assign _36817_ = _36818_ | _36820_ /*36290*/;
assign _36826_ = ~D[17] /*36289*/;
assign _36823_ = _36241_ & _36826_ /*36285*/;
assign _36824_ = _36241_ ^ _36826_ /*36288*/;
assign _36825_ = _36817_ & _36824_ /*36286*/;
assign _36690_ = _36817_ ^ _36824_ /*36287*/;
assign _36822_ = _36823_ | _36825_ /*36284*/;
assign _36831_ = ~D[18] /*36283*/;
assign _36828_ = _36242_ & _36831_ /*36279*/;
assign _36829_ = _36242_ ^ _36831_ /*36282*/;
assign _36830_ = _36822_ & _36829_ /*36280*/;
assign _36691_ = _36822_ ^ _36829_ /*36281*/;
assign _36827_ = _36828_ | _36830_ /*36278*/;
assign _36836_ = ~D[19] /*36277*/;
assign _36833_ = _36243_ & _36836_ /*36273*/;
assign _36834_ = _36243_ ^ _36836_ /*36276*/;
assign _36835_ = _36827_ & _36834_ /*36274*/;
assign _36692_ = _36827_ ^ _36834_ /*36275*/;
assign _36832_ = _36833_ | _36835_ /*36272*/;
assign _36841_ = ~D[20] /*36271*/;
assign _36838_ = _36244_ & _36841_ /*36267*/;
assign _36839_ = _36244_ ^ _36841_ /*36270*/;
assign _36840_ = _36832_ & _36839_ /*36268*/;
assign _36693_ = _36832_ ^ _36839_ /*36269*/;
assign _36837_ = _36838_ | _36840_ /*36266*/;
assign _36846_ = ~D[21] /*36265*/;
assign _36843_ = _36245_ & _36846_ /*36261*/;
assign _36844_ = _36245_ ^ _36846_ /*36264*/;
assign _36845_ = _36837_ & _36844_ /*36262*/;
assign _36694_ = _36837_ ^ _36844_ /*36263*/;
assign _36842_ = _36843_ | _36845_ /*36260*/;
assign _36851_ = ~D[22] /*36259*/;
assign _36848_ = _36246_ & _36851_ /*36255*/;
assign _36849_ = _36246_ ^ _36851_ /*36258*/;
assign _36850_ = _36842_ & _36849_ /*36256*/;
assign _36695_ = _36842_ ^ _36849_ /*36257*/;
assign _36847_ = _36848_ | _36850_ /*36254*/;
assign _36856_ = ~D[23] /*36253*/;
assign _36853_ = _36247_ & _36856_ /*36249*/;
assign _36854_ = _36247_ ^ _36856_ /*36252*/;
assign _36855_ = _36847_ & _36854_ /*36250*/;
assign _36696_ = _36847_ ^ _36854_ /*36251*/;
assign _36852_ = _36853_ | _36855_ /*36248*/;
assign _36861_ = ~D[24] /*36247*/;
assign _36858_ = _36248_ & _36861_ /*36243*/;
assign _36859_ = _36248_ ^ _36861_ /*36246*/;
assign _36860_ = _36852_ & _36859_ /*36244*/;
assign _36697_ = _36852_ ^ _36859_ /*36245*/;
assign _36857_ = _36858_ | _36860_ /*36242*/;
assign _36866_ = ~D[25] /*36241*/;
assign _36863_ = _36249_ & _36866_ /*36237*/;
assign _36864_ = _36249_ ^ _36866_ /*36240*/;
assign _36865_ = _36857_ & _36864_ /*36238*/;
assign _36698_ = _36857_ ^ _36864_ /*36239*/;
assign _36862_ = _36863_ | _36865_ /*36236*/;
assign _36871_ = ~D[26] /*36235*/;
assign _36868_ = _36250_ & _36871_ /*36231*/;
assign _36869_ = _36250_ ^ _36871_ /*36234*/;
assign _36870_ = _36862_ & _36869_ /*36232*/;
assign _36699_ = _36862_ ^ _36869_ /*36233*/;
assign _36867_ = _36868_ | _36870_ /*36230*/;
assign _36876_ = ~D[27] /*36229*/;
assign _36873_ = _36251_ & _36876_ /*36225*/;
assign _36874_ = _36251_ ^ _36876_ /*36228*/;
assign _36875_ = _36867_ & _36874_ /*36226*/;
assign _36700_ = _36867_ ^ _36874_ /*36227*/;
assign _36872_ = _36873_ | _36875_ /*36224*/;
assign _36881_ = ~D[28] /*36223*/;
assign _36878_ = _36252_ & _36881_ /*36219*/;
assign _36879_ = _36252_ ^ _36881_ /*36222*/;
assign _36880_ = _36872_ & _36879_ /*36220*/;
assign _36701_ = _36872_ ^ _36879_ /*36221*/;
assign _36877_ = _36878_ | _36880_ /*36218*/;
assign _36886_ = ~D[29] /*36217*/;
assign _36883_ = _36253_ & _36886_ /*36213*/;
assign _36884_ = _36253_ ^ _36886_ /*36216*/;
assign _36885_ = _36877_ & _36884_ /*36214*/;
assign _36702_ = _36877_ ^ _36884_ /*36215*/;
assign _36882_ = _36883_ | _36885_ /*36212*/;
assign _36891_ = ~D[30] /*36211*/;
assign _36888_ = _36254_ & _36891_ /*36207*/;
assign _36889_ = _36254_ ^ _36891_ /*36210*/;
assign _36890_ = _36882_ & _36889_ /*36208*/;
assign _36703_ = _36882_ ^ _36889_ /*36209*/;
assign _36887_ = _36888_ | _36890_ /*36206*/;
assign _36896_ = ~D[31] /*36205*/;
assign _36893_ = _36255_ & _36896_ /*36201*/;
assign _36894_ = _36255_ ^ _36896_ /*36204*/;
assign _36895_ = _36887_ & _36894_ /*36202*/;
assign _36704_ = _36887_ ^ _36894_ /*36203*/;
assign _36892_ = _36893_ | _36895_ /*36200*/;
assign _36901_ = ~D[32] /*36199*/;
assign _36898_ = _36256_ & _36901_ /*36195*/;
assign _36899_ = _36256_ ^ _36901_ /*36198*/;
assign _36900_ = _36892_ & _36899_ /*36196*/;
assign _36705_ = _36892_ ^ _36899_ /*36197*/;
assign _36897_ = _36898_ | _36900_ /*36194*/;
assign _36906_ = ~D[33] /*36193*/;
assign _36903_ = _36257_ & _36906_ /*36189*/;
assign _36904_ = _36257_ ^ _36906_ /*36192*/;
assign _36905_ = _36897_ & _36904_ /*36190*/;
assign _36706_ = _36897_ ^ _36904_ /*36191*/;
assign _36902_ = _36903_ | _36905_ /*36188*/;
assign _36911_ = ~D[34] /*36187*/;
assign _36908_ = _36258_ & _36911_ /*36183*/;
assign _36909_ = _36258_ ^ _36911_ /*36186*/;
assign _36910_ = _36902_ & _36909_ /*36184*/;
assign _36707_ = _36902_ ^ _36909_ /*36185*/;
assign _36907_ = _36908_ | _36910_ /*36182*/;
assign _36916_ = ~D[35] /*36181*/;
assign _36913_ = _36259_ & _36916_ /*36177*/;
assign _36914_ = _36259_ ^ _36916_ /*36180*/;
assign _36915_ = _36907_ & _36914_ /*36178*/;
assign _36708_ = _36907_ ^ _36914_ /*36179*/;
assign _36912_ = _36913_ | _36915_ /*36176*/;
assign _36921_ = ~D[36] /*36175*/;
assign _36918_ = _36260_ & _36921_ /*36171*/;
assign _36919_ = _36260_ ^ _36921_ /*36174*/;
assign _36920_ = _36912_ & _36919_ /*36172*/;
assign _36709_ = _36912_ ^ _36919_ /*36173*/;
assign _36917_ = _36918_ | _36920_ /*36170*/;
assign _36926_ = ~D[37] /*36169*/;
assign _36923_ = _36261_ & _36926_ /*36165*/;
assign _36924_ = _36261_ ^ _36926_ /*36168*/;
assign _36925_ = _36917_ & _36924_ /*36166*/;
assign _36710_ = _36917_ ^ _36924_ /*36167*/;
assign _36922_ = _36923_ | _36925_ /*36164*/;
assign _36931_ = ~D[38] /*36163*/;
assign _36928_ = _36262_ & _36931_ /*36159*/;
assign _36929_ = _36262_ ^ _36931_ /*36162*/;
assign _36930_ = _36922_ & _36929_ /*36160*/;
assign _36711_ = _36922_ ^ _36929_ /*36161*/;
assign _36927_ = _36928_ | _36930_ /*36158*/;
assign _36936_ = ~D[39] /*36157*/;
assign _36933_ = _36263_ & _36936_ /*36153*/;
assign _36934_ = _36263_ ^ _36936_ /*36156*/;
assign _36935_ = _36927_ & _36934_ /*36154*/;
assign _36712_ = _36927_ ^ _36934_ /*36155*/;
assign _36932_ = _36933_ | _36935_ /*36152*/;
assign _36941_ = ~D[40] /*36151*/;
assign _36938_ = _36264_ & _36941_ /*36147*/;
assign _36939_ = _36264_ ^ _36941_ /*36150*/;
assign _36940_ = _36932_ & _36939_ /*36148*/;
assign _36713_ = _36932_ ^ _36939_ /*36149*/;
assign _36937_ = _36938_ | _36940_ /*36146*/;
assign _36946_ = ~D[41] /*36145*/;
assign _36943_ = _36265_ & _36946_ /*36141*/;
assign _36944_ = _36265_ ^ _36946_ /*36144*/;
assign _36945_ = _36937_ & _36944_ /*36142*/;
assign _36714_ = _36937_ ^ _36944_ /*36143*/;
assign _36942_ = _36943_ | _36945_ /*36140*/;
assign _36951_ = ~D[42] /*36139*/;
assign _36948_ = _36266_ & _36951_ /*36135*/;
assign _36949_ = _36266_ ^ _36951_ /*36138*/;
assign _36950_ = _36942_ & _36949_ /*36136*/;
assign _36715_ = _36942_ ^ _36949_ /*36137*/;
assign _36947_ = _36948_ | _36950_ /*36134*/;
assign _36956_ = ~D[43] /*36133*/;
assign _36953_ = _36267_ & _36956_ /*36129*/;
assign _36954_ = _36267_ ^ _36956_ /*36132*/;
assign _36955_ = _36947_ & _36954_ /*36130*/;
assign _36716_ = _36947_ ^ _36954_ /*36131*/;
assign _36952_ = _36953_ | _36955_ /*36128*/;
assign _36961_ = ~D[44] /*36127*/;
assign _36958_ = _36268_ & _36961_ /*36123*/;
assign _36959_ = _36268_ ^ _36961_ /*36126*/;
assign _36960_ = _36952_ & _36959_ /*36124*/;
assign _36717_ = _36952_ ^ _36959_ /*36125*/;
assign _36957_ = _36958_ | _36960_ /*36122*/;
assign _36966_ = ~D[45] /*36121*/;
assign _36963_ = _36269_ & _36966_ /*36117*/;
assign _36964_ = _36269_ ^ _36966_ /*36120*/;
assign _36965_ = _36957_ & _36964_ /*36118*/;
assign _36718_ = _36957_ ^ _36964_ /*36119*/;
assign _36962_ = _36963_ | _36965_ /*36116*/;
assign _36971_ = ~D[46] /*36115*/;
assign _36968_ = _36270_ & _36971_ /*36111*/;
assign _36969_ = _36270_ ^ _36971_ /*36114*/;
assign _36970_ = _36962_ & _36969_ /*36112*/;
assign _36719_ = _36962_ ^ _36969_ /*36113*/;
assign _36967_ = _36968_ | _36970_ /*36110*/;
assign _36976_ = ~D[47] /*36109*/;
assign _36973_ = _36271_ & _36976_ /*36105*/;
assign _36974_ = _36271_ ^ _36976_ /*36108*/;
assign _36975_ = _36967_ & _36974_ /*36106*/;
assign _36720_ = _36967_ ^ _36974_ /*36107*/;
assign _36972_ = _36973_ | _36975_ /*36104*/;
assign _36981_ = ~D[48] /*36103*/;
assign _36978_ = _36272_ & _36981_ /*36099*/;
assign _36979_ = _36272_ ^ _36981_ /*36102*/;
assign _36980_ = _36972_ & _36979_ /*36100*/;
assign _36721_ = _36972_ ^ _36979_ /*36101*/;
assign _36977_ = _36978_ | _36980_ /*36098*/;
assign _36986_ = ~D[49] /*36097*/;
assign _36983_ = _36273_ & _36986_ /*36093*/;
assign _36984_ = _36273_ ^ _36986_ /*36096*/;
assign _36985_ = _36977_ & _36984_ /*36094*/;
assign _36722_ = _36977_ ^ _36984_ /*36095*/;
assign _36982_ = _36983_ | _36985_ /*36092*/;
assign _36991_ = ~D[50] /*36091*/;
assign _36988_ = _36274_ & _36991_ /*36087*/;
assign _36989_ = _36274_ ^ _36991_ /*36090*/;
assign _36990_ = _36982_ & _36989_ /*36088*/;
assign _36723_ = _36982_ ^ _36989_ /*36089*/;
assign _36987_ = _36988_ | _36990_ /*36086*/;
assign _36996_ = ~D[51] /*36085*/;
assign _36993_ = _36275_ & _36996_ /*36081*/;
assign _36994_ = _36275_ ^ _36996_ /*36084*/;
assign _36995_ = _36987_ & _36994_ /*36082*/;
assign _36724_ = _36987_ ^ _36994_ /*36083*/;
assign _36992_ = _36993_ | _36995_ /*36080*/;
assign _37001_ = ~D[52] /*36079*/;
assign _36998_ = _36276_ & _37001_ /*36075*/;
assign _36999_ = _36276_ ^ _37001_ /*36078*/;
assign _37000_ = _36992_ & _36999_ /*36076*/;
assign _36725_ = _36992_ ^ _36999_ /*36077*/;
assign _36997_ = _36998_ | _37000_ /*36074*/;
assign _37006_ = ~D[53] /*36073*/;
assign _37003_ = _36277_ & _37006_ /*36069*/;
assign _37004_ = _36277_ ^ _37006_ /*36072*/;
assign _37005_ = _36997_ & _37004_ /*36070*/;
assign _36726_ = _36997_ ^ _37004_ /*36071*/;
assign _37002_ = _37003_ | _37005_ /*36068*/;
assign _37011_ = ~D[54] /*36067*/;
assign _37008_ = _36278_ & _37011_ /*36063*/;
assign _37009_ = _36278_ ^ _37011_ /*36066*/;
assign _37010_ = _37002_ & _37009_ /*36064*/;
assign _36727_ = _37002_ ^ _37009_ /*36065*/;
assign _37007_ = _37008_ | _37010_ /*36062*/;
assign _37016_ = ~D[55] /*36061*/;
assign _37013_ = _36279_ & _37016_ /*36057*/;
assign _37014_ = _36279_ ^ _37016_ /*36060*/;
assign _37015_ = _37007_ & _37014_ /*36058*/;
assign _36728_ = _37007_ ^ _37014_ /*36059*/;
assign _37012_ = _37013_ | _37015_ /*36056*/;
assign _37021_ = ~D[56] /*36055*/;
assign _37018_ = _36280_ & _37021_ /*36051*/;
assign _37019_ = _36280_ ^ _37021_ /*36054*/;
assign _37020_ = _37012_ & _37019_ /*36052*/;
assign _36729_ = _37012_ ^ _37019_ /*36053*/;
assign _37017_ = _37018_ | _37020_ /*36050*/;
assign _37026_ = ~D[57] /*36049*/;
assign _37023_ = _36281_ & _37026_ /*36045*/;
assign _37024_ = _36281_ ^ _37026_ /*36048*/;
assign _37025_ = _37017_ & _37024_ /*36046*/;
assign _36730_ = _37017_ ^ _37024_ /*36047*/;
assign _37022_ = _37023_ | _37025_ /*36044*/;
assign _37031_ = ~D[58] /*36043*/;
assign _37028_ = _36282_ & _37031_ /*36039*/;
assign _37029_ = _36282_ ^ _37031_ /*36042*/;
assign _37030_ = _37022_ & _37029_ /*36040*/;
assign _36731_ = _37022_ ^ _37029_ /*36041*/;
assign _37027_ = _37028_ | _37030_ /*36038*/;
assign _37036_ = ~D[59] /*36037*/;
assign _37033_ = _36283_ & _37036_ /*36033*/;
assign _37034_ = _36283_ ^ _37036_ /*36036*/;
assign _37035_ = _37027_ & _37034_ /*36034*/;
assign _36732_ = _37027_ ^ _37034_ /*36035*/;
assign _37032_ = _37033_ | _37035_ /*36032*/;
assign _37041_ = ~D[60] /*36031*/;
assign _37038_ = _36284_ & _37041_ /*36027*/;
assign _37039_ = _36284_ ^ _37041_ /*36030*/;
assign _37040_ = _37032_ & _37039_ /*36028*/;
assign _36733_ = _37032_ ^ _37039_ /*36029*/;
assign _37037_ = _37038_ | _37040_ /*36026*/;
assign _37046_ = ~D[61] /*36025*/;
assign _37043_ = _36285_ & _37046_ /*36021*/;
assign _37044_ = _36285_ ^ _37046_ /*36024*/;
assign _37045_ = _37037_ & _37044_ /*36022*/;
assign _36734_ = _37037_ ^ _37044_ /*36023*/;
assign _37042_ = _37043_ | _37045_ /*36020*/;
assign _37051_ = ~D[62] /*36019*/;
assign _37048_ = _36286_ & _37051_ /*36015*/;
assign _37049_ = _36286_ ^ _37051_ /*36018*/;
assign _37050_ = _37042_ & _37049_ /*36016*/;
assign _36735_ = _37042_ ^ _37049_ /*36017*/;
assign _37047_ = _37048_ | _37050_ /*36014*/;
assign _37052_ = _36287_ & oneWire /*36009*/;
assign _37053_ = _36287_ ^ oneWire /*36012*/;
assign _37054_ = _37047_ & _37053_ /*36010*/;
assign _36736_ = _37047_ ^ _37053_ /*36011*/;
assign Q[22] = _37052_ | _37054_ /*36008*/;
assign _37187_ = ~Q[22] /*35623*/;
assign _37186_ = _37187_ & D[0] /*35622*/;
assign _37189_ = _36673_ & _37186_ /*35617*/;
assign _37190_ = _36673_ ^ _37186_ /*35620*/;
assign _37191_ = zeroWire & _37190_ /*35618*/;
assign _37121_ = zeroWire ^ _37190_ /*35619*/;
assign _37188_ = _37189_ | _37191_ /*35616*/;
assign _37193_ = ~Q[22] /*35615*/;
assign _37192_ = _37193_ & D[1] /*35614*/;
assign _37195_ = _36674_ & _37192_ /*35609*/;
assign _37196_ = _36674_ ^ _37192_ /*35612*/;
assign _37197_ = _37188_ & _37196_ /*35610*/;
assign _37122_ = _37188_ ^ _37196_ /*35611*/;
assign _37194_ = _37195_ | _37197_ /*35608*/;
assign _37199_ = ~Q[22] /*35607*/;
assign _37198_ = _37199_ & D[2] /*35606*/;
assign _37201_ = _36675_ & _37198_ /*35601*/;
assign _37202_ = _36675_ ^ _37198_ /*35604*/;
assign _37203_ = _37194_ & _37202_ /*35602*/;
assign _37123_ = _37194_ ^ _37202_ /*35603*/;
assign _37200_ = _37201_ | _37203_ /*35600*/;
assign _37205_ = ~Q[22] /*35599*/;
assign _37204_ = _37205_ & D[3] /*35598*/;
assign _37207_ = _36676_ & _37204_ /*35593*/;
assign _37208_ = _36676_ ^ _37204_ /*35596*/;
assign _37209_ = _37200_ & _37208_ /*35594*/;
assign _37124_ = _37200_ ^ _37208_ /*35595*/;
assign _37206_ = _37207_ | _37209_ /*35592*/;
assign _37211_ = ~Q[22] /*35591*/;
assign _37210_ = _37211_ & D[4] /*35590*/;
assign _37213_ = _36677_ & _37210_ /*35585*/;
assign _37214_ = _36677_ ^ _37210_ /*35588*/;
assign _37215_ = _37206_ & _37214_ /*35586*/;
assign _37125_ = _37206_ ^ _37214_ /*35587*/;
assign _37212_ = _37213_ | _37215_ /*35584*/;
assign _37217_ = ~Q[22] /*35583*/;
assign _37216_ = _37217_ & D[5] /*35582*/;
assign _37219_ = _36678_ & _37216_ /*35577*/;
assign _37220_ = _36678_ ^ _37216_ /*35580*/;
assign _37221_ = _37212_ & _37220_ /*35578*/;
assign _37126_ = _37212_ ^ _37220_ /*35579*/;
assign _37218_ = _37219_ | _37221_ /*35576*/;
assign _37223_ = ~Q[22] /*35575*/;
assign _37222_ = _37223_ & D[6] /*35574*/;
assign _37225_ = _36679_ & _37222_ /*35569*/;
assign _37226_ = _36679_ ^ _37222_ /*35572*/;
assign _37227_ = _37218_ & _37226_ /*35570*/;
assign _37127_ = _37218_ ^ _37226_ /*35571*/;
assign _37224_ = _37225_ | _37227_ /*35568*/;
assign _37229_ = ~Q[22] /*35567*/;
assign _37228_ = _37229_ & D[7] /*35566*/;
assign _37231_ = _36680_ & _37228_ /*35561*/;
assign _37232_ = _36680_ ^ _37228_ /*35564*/;
assign _37233_ = _37224_ & _37232_ /*35562*/;
assign _37128_ = _37224_ ^ _37232_ /*35563*/;
assign _37230_ = _37231_ | _37233_ /*35560*/;
assign _37235_ = ~Q[22] /*35559*/;
assign _37234_ = _37235_ & D[8] /*35558*/;
assign _37237_ = _36681_ & _37234_ /*35553*/;
assign _37238_ = _36681_ ^ _37234_ /*35556*/;
assign _37239_ = _37230_ & _37238_ /*35554*/;
assign _37129_ = _37230_ ^ _37238_ /*35555*/;
assign _37236_ = _37237_ | _37239_ /*35552*/;
assign _37241_ = ~Q[22] /*35551*/;
assign _37240_ = _37241_ & D[9] /*35550*/;
assign _37243_ = _36682_ & _37240_ /*35545*/;
assign _37244_ = _36682_ ^ _37240_ /*35548*/;
assign _37245_ = _37236_ & _37244_ /*35546*/;
assign _37130_ = _37236_ ^ _37244_ /*35547*/;
assign _37242_ = _37243_ | _37245_ /*35544*/;
assign _37247_ = ~Q[22] /*35543*/;
assign _37246_ = _37247_ & D[10] /*35542*/;
assign _37249_ = _36683_ & _37246_ /*35537*/;
assign _37250_ = _36683_ ^ _37246_ /*35540*/;
assign _37251_ = _37242_ & _37250_ /*35538*/;
assign _37131_ = _37242_ ^ _37250_ /*35539*/;
assign _37248_ = _37249_ | _37251_ /*35536*/;
assign _37253_ = ~Q[22] /*35535*/;
assign _37252_ = _37253_ & D[11] /*35534*/;
assign _37255_ = _36684_ & _37252_ /*35529*/;
assign _37256_ = _36684_ ^ _37252_ /*35532*/;
assign _37257_ = _37248_ & _37256_ /*35530*/;
assign _37132_ = _37248_ ^ _37256_ /*35531*/;
assign _37254_ = _37255_ | _37257_ /*35528*/;
assign _37259_ = ~Q[22] /*35527*/;
assign _37258_ = _37259_ & D[12] /*35526*/;
assign _37261_ = _36685_ & _37258_ /*35521*/;
assign _37262_ = _36685_ ^ _37258_ /*35524*/;
assign _37263_ = _37254_ & _37262_ /*35522*/;
assign _37133_ = _37254_ ^ _37262_ /*35523*/;
assign _37260_ = _37261_ | _37263_ /*35520*/;
assign _37265_ = ~Q[22] /*35519*/;
assign _37264_ = _37265_ & D[13] /*35518*/;
assign _37267_ = _36686_ & _37264_ /*35513*/;
assign _37268_ = _36686_ ^ _37264_ /*35516*/;
assign _37269_ = _37260_ & _37268_ /*35514*/;
assign _37134_ = _37260_ ^ _37268_ /*35515*/;
assign _37266_ = _37267_ | _37269_ /*35512*/;
assign _37271_ = ~Q[22] /*35511*/;
assign _37270_ = _37271_ & D[14] /*35510*/;
assign _37273_ = _36687_ & _37270_ /*35505*/;
assign _37274_ = _36687_ ^ _37270_ /*35508*/;
assign _37275_ = _37266_ & _37274_ /*35506*/;
assign _37135_ = _37266_ ^ _37274_ /*35507*/;
assign _37272_ = _37273_ | _37275_ /*35504*/;
assign _37277_ = ~Q[22] /*35503*/;
assign _37276_ = _37277_ & D[15] /*35502*/;
assign _37279_ = _36688_ & _37276_ /*35497*/;
assign _37280_ = _36688_ ^ _37276_ /*35500*/;
assign _37281_ = _37272_ & _37280_ /*35498*/;
assign _37136_ = _37272_ ^ _37280_ /*35499*/;
assign _37278_ = _37279_ | _37281_ /*35496*/;
assign _37283_ = ~Q[22] /*35495*/;
assign _37282_ = _37283_ & D[16] /*35494*/;
assign _37285_ = _36689_ & _37282_ /*35489*/;
assign _37286_ = _36689_ ^ _37282_ /*35492*/;
assign _37287_ = _37278_ & _37286_ /*35490*/;
assign _37137_ = _37278_ ^ _37286_ /*35491*/;
assign _37284_ = _37285_ | _37287_ /*35488*/;
assign _37289_ = ~Q[22] /*35487*/;
assign _37288_ = _37289_ & D[17] /*35486*/;
assign _37291_ = _36690_ & _37288_ /*35481*/;
assign _37292_ = _36690_ ^ _37288_ /*35484*/;
assign _37293_ = _37284_ & _37292_ /*35482*/;
assign _37138_ = _37284_ ^ _37292_ /*35483*/;
assign _37290_ = _37291_ | _37293_ /*35480*/;
assign _37295_ = ~Q[22] /*35479*/;
assign _37294_ = _37295_ & D[18] /*35478*/;
assign _37297_ = _36691_ & _37294_ /*35473*/;
assign _37298_ = _36691_ ^ _37294_ /*35476*/;
assign _37299_ = _37290_ & _37298_ /*35474*/;
assign _37139_ = _37290_ ^ _37298_ /*35475*/;
assign _37296_ = _37297_ | _37299_ /*35472*/;
assign _37301_ = ~Q[22] /*35471*/;
assign _37300_ = _37301_ & D[19] /*35470*/;
assign _37303_ = _36692_ & _37300_ /*35465*/;
assign _37304_ = _36692_ ^ _37300_ /*35468*/;
assign _37305_ = _37296_ & _37304_ /*35466*/;
assign _37140_ = _37296_ ^ _37304_ /*35467*/;
assign _37302_ = _37303_ | _37305_ /*35464*/;
assign _37307_ = ~Q[22] /*35463*/;
assign _37306_ = _37307_ & D[20] /*35462*/;
assign _37309_ = _36693_ & _37306_ /*35457*/;
assign _37310_ = _36693_ ^ _37306_ /*35460*/;
assign _37311_ = _37302_ & _37310_ /*35458*/;
assign _37141_ = _37302_ ^ _37310_ /*35459*/;
assign _37308_ = _37309_ | _37311_ /*35456*/;
assign _37313_ = ~Q[22] /*35455*/;
assign _37312_ = _37313_ & D[21] /*35454*/;
assign _37315_ = _36694_ & _37312_ /*35449*/;
assign _37316_ = _36694_ ^ _37312_ /*35452*/;
assign _37317_ = _37308_ & _37316_ /*35450*/;
assign _37142_ = _37308_ ^ _37316_ /*35451*/;
assign _37314_ = _37315_ | _37317_ /*35448*/;
assign _37319_ = ~Q[22] /*35447*/;
assign _37318_ = _37319_ & D[22] /*35446*/;
assign _37321_ = _36695_ & _37318_ /*35441*/;
assign _37322_ = _36695_ ^ _37318_ /*35444*/;
assign _37323_ = _37314_ & _37322_ /*35442*/;
assign _37143_ = _37314_ ^ _37322_ /*35443*/;
assign _37320_ = _37321_ | _37323_ /*35440*/;
assign _37325_ = ~Q[22] /*35439*/;
assign _37324_ = _37325_ & D[23] /*35438*/;
assign _37327_ = _36696_ & _37324_ /*35433*/;
assign _37328_ = _36696_ ^ _37324_ /*35436*/;
assign _37329_ = _37320_ & _37328_ /*35434*/;
assign _37144_ = _37320_ ^ _37328_ /*35435*/;
assign _37326_ = _37327_ | _37329_ /*35432*/;
assign _37331_ = ~Q[22] /*35431*/;
assign _37330_ = _37331_ & D[24] /*35430*/;
assign _37333_ = _36697_ & _37330_ /*35425*/;
assign _37334_ = _36697_ ^ _37330_ /*35428*/;
assign _37335_ = _37326_ & _37334_ /*35426*/;
assign _37145_ = _37326_ ^ _37334_ /*35427*/;
assign _37332_ = _37333_ | _37335_ /*35424*/;
assign _37337_ = ~Q[22] /*35423*/;
assign _37336_ = _37337_ & D[25] /*35422*/;
assign _37339_ = _36698_ & _37336_ /*35417*/;
assign _37340_ = _36698_ ^ _37336_ /*35420*/;
assign _37341_ = _37332_ & _37340_ /*35418*/;
assign _37146_ = _37332_ ^ _37340_ /*35419*/;
assign _37338_ = _37339_ | _37341_ /*35416*/;
assign _37343_ = ~Q[22] /*35415*/;
assign _37342_ = _37343_ & D[26] /*35414*/;
assign _37345_ = _36699_ & _37342_ /*35409*/;
assign _37346_ = _36699_ ^ _37342_ /*35412*/;
assign _37347_ = _37338_ & _37346_ /*35410*/;
assign _37147_ = _37338_ ^ _37346_ /*35411*/;
assign _37344_ = _37345_ | _37347_ /*35408*/;
assign _37349_ = ~Q[22] /*35407*/;
assign _37348_ = _37349_ & D[27] /*35406*/;
assign _37351_ = _36700_ & _37348_ /*35401*/;
assign _37352_ = _36700_ ^ _37348_ /*35404*/;
assign _37353_ = _37344_ & _37352_ /*35402*/;
assign _37148_ = _37344_ ^ _37352_ /*35403*/;
assign _37350_ = _37351_ | _37353_ /*35400*/;
assign _37355_ = ~Q[22] /*35399*/;
assign _37354_ = _37355_ & D[28] /*35398*/;
assign _37357_ = _36701_ & _37354_ /*35393*/;
assign _37358_ = _36701_ ^ _37354_ /*35396*/;
assign _37359_ = _37350_ & _37358_ /*35394*/;
assign _37149_ = _37350_ ^ _37358_ /*35395*/;
assign _37356_ = _37357_ | _37359_ /*35392*/;
assign _37361_ = ~Q[22] /*35391*/;
assign _37360_ = _37361_ & D[29] /*35390*/;
assign _37363_ = _36702_ & _37360_ /*35385*/;
assign _37364_ = _36702_ ^ _37360_ /*35388*/;
assign _37365_ = _37356_ & _37364_ /*35386*/;
assign _37150_ = _37356_ ^ _37364_ /*35387*/;
assign _37362_ = _37363_ | _37365_ /*35384*/;
assign _37367_ = ~Q[22] /*35383*/;
assign _37366_ = _37367_ & D[30] /*35382*/;
assign _37369_ = _36703_ & _37366_ /*35377*/;
assign _37370_ = _36703_ ^ _37366_ /*35380*/;
assign _37371_ = _37362_ & _37370_ /*35378*/;
assign _37151_ = _37362_ ^ _37370_ /*35379*/;
assign _37368_ = _37369_ | _37371_ /*35376*/;
assign _37373_ = ~Q[22] /*35375*/;
assign _37372_ = _37373_ & D[31] /*35374*/;
assign _37375_ = _36704_ & _37372_ /*35369*/;
assign _37376_ = _36704_ ^ _37372_ /*35372*/;
assign _37377_ = _37368_ & _37376_ /*35370*/;
assign _37152_ = _37368_ ^ _37376_ /*35371*/;
assign _37374_ = _37375_ | _37377_ /*35368*/;
assign _37379_ = ~Q[22] /*35367*/;
assign _37378_ = _37379_ & D[32] /*35366*/;
assign _37381_ = _36705_ & _37378_ /*35361*/;
assign _37382_ = _36705_ ^ _37378_ /*35364*/;
assign _37383_ = _37374_ & _37382_ /*35362*/;
assign _37153_ = _37374_ ^ _37382_ /*35363*/;
assign _37380_ = _37381_ | _37383_ /*35360*/;
assign _37385_ = ~Q[22] /*35359*/;
assign _37384_ = _37385_ & D[33] /*35358*/;
assign _37387_ = _36706_ & _37384_ /*35353*/;
assign _37388_ = _36706_ ^ _37384_ /*35356*/;
assign _37389_ = _37380_ & _37388_ /*35354*/;
assign _37154_ = _37380_ ^ _37388_ /*35355*/;
assign _37386_ = _37387_ | _37389_ /*35352*/;
assign _37391_ = ~Q[22] /*35351*/;
assign _37390_ = _37391_ & D[34] /*35350*/;
assign _37393_ = _36707_ & _37390_ /*35345*/;
assign _37394_ = _36707_ ^ _37390_ /*35348*/;
assign _37395_ = _37386_ & _37394_ /*35346*/;
assign _37155_ = _37386_ ^ _37394_ /*35347*/;
assign _37392_ = _37393_ | _37395_ /*35344*/;
assign _37397_ = ~Q[22] /*35343*/;
assign _37396_ = _37397_ & D[35] /*35342*/;
assign _37399_ = _36708_ & _37396_ /*35337*/;
assign _37400_ = _36708_ ^ _37396_ /*35340*/;
assign _37401_ = _37392_ & _37400_ /*35338*/;
assign _37156_ = _37392_ ^ _37400_ /*35339*/;
assign _37398_ = _37399_ | _37401_ /*35336*/;
assign _37403_ = ~Q[22] /*35335*/;
assign _37402_ = _37403_ & D[36] /*35334*/;
assign _37405_ = _36709_ & _37402_ /*35329*/;
assign _37406_ = _36709_ ^ _37402_ /*35332*/;
assign _37407_ = _37398_ & _37406_ /*35330*/;
assign _37157_ = _37398_ ^ _37406_ /*35331*/;
assign _37404_ = _37405_ | _37407_ /*35328*/;
assign _37409_ = ~Q[22] /*35327*/;
assign _37408_ = _37409_ & D[37] /*35326*/;
assign _37411_ = _36710_ & _37408_ /*35321*/;
assign _37412_ = _36710_ ^ _37408_ /*35324*/;
assign _37413_ = _37404_ & _37412_ /*35322*/;
assign _37158_ = _37404_ ^ _37412_ /*35323*/;
assign _37410_ = _37411_ | _37413_ /*35320*/;
assign _37415_ = ~Q[22] /*35319*/;
assign _37414_ = _37415_ & D[38] /*35318*/;
assign _37417_ = _36711_ & _37414_ /*35313*/;
assign _37418_ = _36711_ ^ _37414_ /*35316*/;
assign _37419_ = _37410_ & _37418_ /*35314*/;
assign _37159_ = _37410_ ^ _37418_ /*35315*/;
assign _37416_ = _37417_ | _37419_ /*35312*/;
assign _37421_ = ~Q[22] /*35311*/;
assign _37420_ = _37421_ & D[39] /*35310*/;
assign _37423_ = _36712_ & _37420_ /*35305*/;
assign _37424_ = _36712_ ^ _37420_ /*35308*/;
assign _37425_ = _37416_ & _37424_ /*35306*/;
assign _37160_ = _37416_ ^ _37424_ /*35307*/;
assign _37422_ = _37423_ | _37425_ /*35304*/;
assign _37427_ = ~Q[22] /*35303*/;
assign _37426_ = _37427_ & D[40] /*35302*/;
assign _37429_ = _36713_ & _37426_ /*35297*/;
assign _37430_ = _36713_ ^ _37426_ /*35300*/;
assign _37431_ = _37422_ & _37430_ /*35298*/;
assign _37161_ = _37422_ ^ _37430_ /*35299*/;
assign _37428_ = _37429_ | _37431_ /*35296*/;
assign _37433_ = ~Q[22] /*35295*/;
assign _37432_ = _37433_ & D[41] /*35294*/;
assign _37435_ = _36714_ & _37432_ /*35289*/;
assign _37436_ = _36714_ ^ _37432_ /*35292*/;
assign _37437_ = _37428_ & _37436_ /*35290*/;
assign _37162_ = _37428_ ^ _37436_ /*35291*/;
assign _37434_ = _37435_ | _37437_ /*35288*/;
assign _37439_ = ~Q[22] /*35287*/;
assign _37438_ = _37439_ & D[42] /*35286*/;
assign _37441_ = _36715_ & _37438_ /*35281*/;
assign _37442_ = _36715_ ^ _37438_ /*35284*/;
assign _37443_ = _37434_ & _37442_ /*35282*/;
assign _37163_ = _37434_ ^ _37442_ /*35283*/;
assign _37440_ = _37441_ | _37443_ /*35280*/;
assign _37445_ = ~Q[22] /*35279*/;
assign _37444_ = _37445_ & D[43] /*35278*/;
assign _37447_ = _36716_ & _37444_ /*35273*/;
assign _37448_ = _36716_ ^ _37444_ /*35276*/;
assign _37449_ = _37440_ & _37448_ /*35274*/;
assign _37164_ = _37440_ ^ _37448_ /*35275*/;
assign _37446_ = _37447_ | _37449_ /*35272*/;
assign _37451_ = ~Q[22] /*35271*/;
assign _37450_ = _37451_ & D[44] /*35270*/;
assign _37453_ = _36717_ & _37450_ /*35265*/;
assign _37454_ = _36717_ ^ _37450_ /*35268*/;
assign _37455_ = _37446_ & _37454_ /*35266*/;
assign _37165_ = _37446_ ^ _37454_ /*35267*/;
assign _37452_ = _37453_ | _37455_ /*35264*/;
assign _37457_ = ~Q[22] /*35263*/;
assign _37456_ = _37457_ & D[45] /*35262*/;
assign _37459_ = _36718_ & _37456_ /*35257*/;
assign _37460_ = _36718_ ^ _37456_ /*35260*/;
assign _37461_ = _37452_ & _37460_ /*35258*/;
assign _37166_ = _37452_ ^ _37460_ /*35259*/;
assign _37458_ = _37459_ | _37461_ /*35256*/;
assign _37463_ = ~Q[22] /*35255*/;
assign _37462_ = _37463_ & D[46] /*35254*/;
assign _37465_ = _36719_ & _37462_ /*35249*/;
assign _37466_ = _36719_ ^ _37462_ /*35252*/;
assign _37467_ = _37458_ & _37466_ /*35250*/;
assign _37167_ = _37458_ ^ _37466_ /*35251*/;
assign _37464_ = _37465_ | _37467_ /*35248*/;
assign _37469_ = ~Q[22] /*35247*/;
assign _37468_ = _37469_ & D[47] /*35246*/;
assign _37471_ = _36720_ & _37468_ /*35241*/;
assign _37472_ = _36720_ ^ _37468_ /*35244*/;
assign _37473_ = _37464_ & _37472_ /*35242*/;
assign _37168_ = _37464_ ^ _37472_ /*35243*/;
assign _37470_ = _37471_ | _37473_ /*35240*/;
assign _37475_ = ~Q[22] /*35239*/;
assign _37474_ = _37475_ & D[48] /*35238*/;
assign _37477_ = _36721_ & _37474_ /*35233*/;
assign _37478_ = _36721_ ^ _37474_ /*35236*/;
assign _37479_ = _37470_ & _37478_ /*35234*/;
assign _37169_ = _37470_ ^ _37478_ /*35235*/;
assign _37476_ = _37477_ | _37479_ /*35232*/;
assign _37481_ = ~Q[22] /*35231*/;
assign _37480_ = _37481_ & D[49] /*35230*/;
assign _37483_ = _36722_ & _37480_ /*35225*/;
assign _37484_ = _36722_ ^ _37480_ /*35228*/;
assign _37485_ = _37476_ & _37484_ /*35226*/;
assign _37170_ = _37476_ ^ _37484_ /*35227*/;
assign _37482_ = _37483_ | _37485_ /*35224*/;
assign _37487_ = ~Q[22] /*35223*/;
assign _37486_ = _37487_ & D[50] /*35222*/;
assign _37489_ = _36723_ & _37486_ /*35217*/;
assign _37490_ = _36723_ ^ _37486_ /*35220*/;
assign _37491_ = _37482_ & _37490_ /*35218*/;
assign _37171_ = _37482_ ^ _37490_ /*35219*/;
assign _37488_ = _37489_ | _37491_ /*35216*/;
assign _37493_ = ~Q[22] /*35215*/;
assign _37492_ = _37493_ & D[51] /*35214*/;
assign _37495_ = _36724_ & _37492_ /*35209*/;
assign _37496_ = _36724_ ^ _37492_ /*35212*/;
assign _37497_ = _37488_ & _37496_ /*35210*/;
assign _37172_ = _37488_ ^ _37496_ /*35211*/;
assign _37494_ = _37495_ | _37497_ /*35208*/;
assign _37499_ = ~Q[22] /*35207*/;
assign _37498_ = _37499_ & D[52] /*35206*/;
assign _37501_ = _36725_ & _37498_ /*35201*/;
assign _37502_ = _36725_ ^ _37498_ /*35204*/;
assign _37503_ = _37494_ & _37502_ /*35202*/;
assign _37173_ = _37494_ ^ _37502_ /*35203*/;
assign _37500_ = _37501_ | _37503_ /*35200*/;
assign _37505_ = ~Q[22] /*35199*/;
assign _37504_ = _37505_ & D[53] /*35198*/;
assign _37507_ = _36726_ & _37504_ /*35193*/;
assign _37508_ = _36726_ ^ _37504_ /*35196*/;
assign _37509_ = _37500_ & _37508_ /*35194*/;
assign _37174_ = _37500_ ^ _37508_ /*35195*/;
assign _37506_ = _37507_ | _37509_ /*35192*/;
assign _37511_ = ~Q[22] /*35191*/;
assign _37510_ = _37511_ & D[54] /*35190*/;
assign _37513_ = _36727_ & _37510_ /*35185*/;
assign _37514_ = _36727_ ^ _37510_ /*35188*/;
assign _37515_ = _37506_ & _37514_ /*35186*/;
assign _37175_ = _37506_ ^ _37514_ /*35187*/;
assign _37512_ = _37513_ | _37515_ /*35184*/;
assign _37517_ = ~Q[22] /*35183*/;
assign _37516_ = _37517_ & D[55] /*35182*/;
assign _37519_ = _36728_ & _37516_ /*35177*/;
assign _37520_ = _36728_ ^ _37516_ /*35180*/;
assign _37521_ = _37512_ & _37520_ /*35178*/;
assign _37176_ = _37512_ ^ _37520_ /*35179*/;
assign _37518_ = _37519_ | _37521_ /*35176*/;
assign _37523_ = ~Q[22] /*35175*/;
assign _37522_ = _37523_ & D[56] /*35174*/;
assign _37525_ = _36729_ & _37522_ /*35169*/;
assign _37526_ = _36729_ ^ _37522_ /*35172*/;
assign _37527_ = _37518_ & _37526_ /*35170*/;
assign _37177_ = _37518_ ^ _37526_ /*35171*/;
assign _37524_ = _37525_ | _37527_ /*35168*/;
assign _37529_ = ~Q[22] /*35167*/;
assign _37528_ = _37529_ & D[57] /*35166*/;
assign _37531_ = _36730_ & _37528_ /*35161*/;
assign _37532_ = _36730_ ^ _37528_ /*35164*/;
assign _37533_ = _37524_ & _37532_ /*35162*/;
assign _37178_ = _37524_ ^ _37532_ /*35163*/;
assign _37530_ = _37531_ | _37533_ /*35160*/;
assign _37535_ = ~Q[22] /*35159*/;
assign _37534_ = _37535_ & D[58] /*35158*/;
assign _37537_ = _36731_ & _37534_ /*35153*/;
assign _37538_ = _36731_ ^ _37534_ /*35156*/;
assign _37539_ = _37530_ & _37538_ /*35154*/;
assign _37179_ = _37530_ ^ _37538_ /*35155*/;
assign _37536_ = _37537_ | _37539_ /*35152*/;
assign _37541_ = ~Q[22] /*35151*/;
assign _37540_ = _37541_ & D[59] /*35150*/;
assign _37543_ = _36732_ & _37540_ /*35145*/;
assign _37544_ = _36732_ ^ _37540_ /*35148*/;
assign _37545_ = _37536_ & _37544_ /*35146*/;
assign _37180_ = _37536_ ^ _37544_ /*35147*/;
assign _37542_ = _37543_ | _37545_ /*35144*/;
assign _37547_ = ~Q[22] /*35143*/;
assign _37546_ = _37547_ & D[60] /*35142*/;
assign _37549_ = _36733_ & _37546_ /*35137*/;
assign _37550_ = _36733_ ^ _37546_ /*35140*/;
assign _37551_ = _37542_ & _37550_ /*35138*/;
assign _37181_ = _37542_ ^ _37550_ /*35139*/;
assign _37548_ = _37549_ | _37551_ /*35136*/;
assign _37553_ = ~Q[22] /*35135*/;
assign _37552_ = _37553_ & D[61] /*35134*/;
assign _37555_ = _36734_ & _37552_ /*35129*/;
assign _37556_ = _36734_ ^ _37552_ /*35132*/;
assign _37557_ = _37548_ & _37556_ /*35130*/;
assign _37182_ = _37548_ ^ _37556_ /*35131*/;
assign _37554_ = _37555_ | _37557_ /*35128*/;
assign _37559_ = ~Q[22] /*35127*/;
assign _37558_ = _37559_ & D[62] /*35126*/;
assign _37561_ = _36735_ & _37558_ /*35121*/;
assign _37562_ = _36735_ ^ _37558_ /*35124*/;
assign _37563_ = _37554_ & _37562_ /*35122*/;
assign _37183_ = _37554_ ^ _37562_ /*35123*/;
assign _37560_ = _37561_ | _37563_ /*35120*/;
assign _37565_ = ~Q[22] /*35119*/;
assign _37564_ = _37565_ & zeroWire /*35118*/;
assign _37566_ = _36736_ ^ _37564_ /*35116*/;
assign _37184_ = _37566_ ^ _37560_ /*35115*/;
assign _37637_ = ~D[0] /*34861*/;
assign _37634_ = R_0[21] & _37637_ /*34857*/;
assign _37635_ = R_0[21] ^ _37637_ /*34860*/;
assign _37636_ = oneWire & _37635_ /*34858*/;
assign _37569_ = oneWire ^ _37635_ /*34859*/;
assign _37633_ = _37634_ | _37636_ /*34856*/;
assign _37642_ = ~D[1] /*34855*/;
assign _37639_ = _37121_ & _37642_ /*34851*/;
assign _37640_ = _37121_ ^ _37642_ /*34854*/;
assign _37641_ = _37633_ & _37640_ /*34852*/;
assign _37570_ = _37633_ ^ _37640_ /*34853*/;
assign _37638_ = _37639_ | _37641_ /*34850*/;
assign _37647_ = ~D[2] /*34849*/;
assign _37644_ = _37122_ & _37647_ /*34845*/;
assign _37645_ = _37122_ ^ _37647_ /*34848*/;
assign _37646_ = _37638_ & _37645_ /*34846*/;
assign _37571_ = _37638_ ^ _37645_ /*34847*/;
assign _37643_ = _37644_ | _37646_ /*34844*/;
assign _37652_ = ~D[3] /*34843*/;
assign _37649_ = _37123_ & _37652_ /*34839*/;
assign _37650_ = _37123_ ^ _37652_ /*34842*/;
assign _37651_ = _37643_ & _37650_ /*34840*/;
assign _37572_ = _37643_ ^ _37650_ /*34841*/;
assign _37648_ = _37649_ | _37651_ /*34838*/;
assign _37657_ = ~D[4] /*34837*/;
assign _37654_ = _37124_ & _37657_ /*34833*/;
assign _37655_ = _37124_ ^ _37657_ /*34836*/;
assign _37656_ = _37648_ & _37655_ /*34834*/;
assign _37573_ = _37648_ ^ _37655_ /*34835*/;
assign _37653_ = _37654_ | _37656_ /*34832*/;
assign _37662_ = ~D[5] /*34831*/;
assign _37659_ = _37125_ & _37662_ /*34827*/;
assign _37660_ = _37125_ ^ _37662_ /*34830*/;
assign _37661_ = _37653_ & _37660_ /*34828*/;
assign _37574_ = _37653_ ^ _37660_ /*34829*/;
assign _37658_ = _37659_ | _37661_ /*34826*/;
assign _37667_ = ~D[6] /*34825*/;
assign _37664_ = _37126_ & _37667_ /*34821*/;
assign _37665_ = _37126_ ^ _37667_ /*34824*/;
assign _37666_ = _37658_ & _37665_ /*34822*/;
assign _37575_ = _37658_ ^ _37665_ /*34823*/;
assign _37663_ = _37664_ | _37666_ /*34820*/;
assign _37672_ = ~D[7] /*34819*/;
assign _37669_ = _37127_ & _37672_ /*34815*/;
assign _37670_ = _37127_ ^ _37672_ /*34818*/;
assign _37671_ = _37663_ & _37670_ /*34816*/;
assign _37576_ = _37663_ ^ _37670_ /*34817*/;
assign _37668_ = _37669_ | _37671_ /*34814*/;
assign _37677_ = ~D[8] /*34813*/;
assign _37674_ = _37128_ & _37677_ /*34809*/;
assign _37675_ = _37128_ ^ _37677_ /*34812*/;
assign _37676_ = _37668_ & _37675_ /*34810*/;
assign _37577_ = _37668_ ^ _37675_ /*34811*/;
assign _37673_ = _37674_ | _37676_ /*34808*/;
assign _37682_ = ~D[9] /*34807*/;
assign _37679_ = _37129_ & _37682_ /*34803*/;
assign _37680_ = _37129_ ^ _37682_ /*34806*/;
assign _37681_ = _37673_ & _37680_ /*34804*/;
assign _37578_ = _37673_ ^ _37680_ /*34805*/;
assign _37678_ = _37679_ | _37681_ /*34802*/;
assign _37687_ = ~D[10] /*34801*/;
assign _37684_ = _37130_ & _37687_ /*34797*/;
assign _37685_ = _37130_ ^ _37687_ /*34800*/;
assign _37686_ = _37678_ & _37685_ /*34798*/;
assign _37579_ = _37678_ ^ _37685_ /*34799*/;
assign _37683_ = _37684_ | _37686_ /*34796*/;
assign _37692_ = ~D[11] /*34795*/;
assign _37689_ = _37131_ & _37692_ /*34791*/;
assign _37690_ = _37131_ ^ _37692_ /*34794*/;
assign _37691_ = _37683_ & _37690_ /*34792*/;
assign _37580_ = _37683_ ^ _37690_ /*34793*/;
assign _37688_ = _37689_ | _37691_ /*34790*/;
assign _37697_ = ~D[12] /*34789*/;
assign _37694_ = _37132_ & _37697_ /*34785*/;
assign _37695_ = _37132_ ^ _37697_ /*34788*/;
assign _37696_ = _37688_ & _37695_ /*34786*/;
assign _37581_ = _37688_ ^ _37695_ /*34787*/;
assign _37693_ = _37694_ | _37696_ /*34784*/;
assign _37702_ = ~D[13] /*34783*/;
assign _37699_ = _37133_ & _37702_ /*34779*/;
assign _37700_ = _37133_ ^ _37702_ /*34782*/;
assign _37701_ = _37693_ & _37700_ /*34780*/;
assign _37582_ = _37693_ ^ _37700_ /*34781*/;
assign _37698_ = _37699_ | _37701_ /*34778*/;
assign _37707_ = ~D[14] /*34777*/;
assign _37704_ = _37134_ & _37707_ /*34773*/;
assign _37705_ = _37134_ ^ _37707_ /*34776*/;
assign _37706_ = _37698_ & _37705_ /*34774*/;
assign _37583_ = _37698_ ^ _37705_ /*34775*/;
assign _37703_ = _37704_ | _37706_ /*34772*/;
assign _37712_ = ~D[15] /*34771*/;
assign _37709_ = _37135_ & _37712_ /*34767*/;
assign _37710_ = _37135_ ^ _37712_ /*34770*/;
assign _37711_ = _37703_ & _37710_ /*34768*/;
assign _37584_ = _37703_ ^ _37710_ /*34769*/;
assign _37708_ = _37709_ | _37711_ /*34766*/;
assign _37717_ = ~D[16] /*34765*/;
assign _37714_ = _37136_ & _37717_ /*34761*/;
assign _37715_ = _37136_ ^ _37717_ /*34764*/;
assign _37716_ = _37708_ & _37715_ /*34762*/;
assign _37585_ = _37708_ ^ _37715_ /*34763*/;
assign _37713_ = _37714_ | _37716_ /*34760*/;
assign _37722_ = ~D[17] /*34759*/;
assign _37719_ = _37137_ & _37722_ /*34755*/;
assign _37720_ = _37137_ ^ _37722_ /*34758*/;
assign _37721_ = _37713_ & _37720_ /*34756*/;
assign _37586_ = _37713_ ^ _37720_ /*34757*/;
assign _37718_ = _37719_ | _37721_ /*34754*/;
assign _37727_ = ~D[18] /*34753*/;
assign _37724_ = _37138_ & _37727_ /*34749*/;
assign _37725_ = _37138_ ^ _37727_ /*34752*/;
assign _37726_ = _37718_ & _37725_ /*34750*/;
assign _37587_ = _37718_ ^ _37725_ /*34751*/;
assign _37723_ = _37724_ | _37726_ /*34748*/;
assign _37732_ = ~D[19] /*34747*/;
assign _37729_ = _37139_ & _37732_ /*34743*/;
assign _37730_ = _37139_ ^ _37732_ /*34746*/;
assign _37731_ = _37723_ & _37730_ /*34744*/;
assign _37588_ = _37723_ ^ _37730_ /*34745*/;
assign _37728_ = _37729_ | _37731_ /*34742*/;
assign _37737_ = ~D[20] /*34741*/;
assign _37734_ = _37140_ & _37737_ /*34737*/;
assign _37735_ = _37140_ ^ _37737_ /*34740*/;
assign _37736_ = _37728_ & _37735_ /*34738*/;
assign _37589_ = _37728_ ^ _37735_ /*34739*/;
assign _37733_ = _37734_ | _37736_ /*34736*/;
assign _37742_ = ~D[21] /*34735*/;
assign _37739_ = _37141_ & _37742_ /*34731*/;
assign _37740_ = _37141_ ^ _37742_ /*34734*/;
assign _37741_ = _37733_ & _37740_ /*34732*/;
assign _37590_ = _37733_ ^ _37740_ /*34733*/;
assign _37738_ = _37739_ | _37741_ /*34730*/;
assign _37747_ = ~D[22] /*34729*/;
assign _37744_ = _37142_ & _37747_ /*34725*/;
assign _37745_ = _37142_ ^ _37747_ /*34728*/;
assign _37746_ = _37738_ & _37745_ /*34726*/;
assign _37591_ = _37738_ ^ _37745_ /*34727*/;
assign _37743_ = _37744_ | _37746_ /*34724*/;
assign _37752_ = ~D[23] /*34723*/;
assign _37749_ = _37143_ & _37752_ /*34719*/;
assign _37750_ = _37143_ ^ _37752_ /*34722*/;
assign _37751_ = _37743_ & _37750_ /*34720*/;
assign _37592_ = _37743_ ^ _37750_ /*34721*/;
assign _37748_ = _37749_ | _37751_ /*34718*/;
assign _37757_ = ~D[24] /*34717*/;
assign _37754_ = _37144_ & _37757_ /*34713*/;
assign _37755_ = _37144_ ^ _37757_ /*34716*/;
assign _37756_ = _37748_ & _37755_ /*34714*/;
assign _37593_ = _37748_ ^ _37755_ /*34715*/;
assign _37753_ = _37754_ | _37756_ /*34712*/;
assign _37762_ = ~D[25] /*34711*/;
assign _37759_ = _37145_ & _37762_ /*34707*/;
assign _37760_ = _37145_ ^ _37762_ /*34710*/;
assign _37761_ = _37753_ & _37760_ /*34708*/;
assign _37594_ = _37753_ ^ _37760_ /*34709*/;
assign _37758_ = _37759_ | _37761_ /*34706*/;
assign _37767_ = ~D[26] /*34705*/;
assign _37764_ = _37146_ & _37767_ /*34701*/;
assign _37765_ = _37146_ ^ _37767_ /*34704*/;
assign _37766_ = _37758_ & _37765_ /*34702*/;
assign _37595_ = _37758_ ^ _37765_ /*34703*/;
assign _37763_ = _37764_ | _37766_ /*34700*/;
assign _37772_ = ~D[27] /*34699*/;
assign _37769_ = _37147_ & _37772_ /*34695*/;
assign _37770_ = _37147_ ^ _37772_ /*34698*/;
assign _37771_ = _37763_ & _37770_ /*34696*/;
assign _37596_ = _37763_ ^ _37770_ /*34697*/;
assign _37768_ = _37769_ | _37771_ /*34694*/;
assign _37777_ = ~D[28] /*34693*/;
assign _37774_ = _37148_ & _37777_ /*34689*/;
assign _37775_ = _37148_ ^ _37777_ /*34692*/;
assign _37776_ = _37768_ & _37775_ /*34690*/;
assign _37597_ = _37768_ ^ _37775_ /*34691*/;
assign _37773_ = _37774_ | _37776_ /*34688*/;
assign _37782_ = ~D[29] /*34687*/;
assign _37779_ = _37149_ & _37782_ /*34683*/;
assign _37780_ = _37149_ ^ _37782_ /*34686*/;
assign _37781_ = _37773_ & _37780_ /*34684*/;
assign _37598_ = _37773_ ^ _37780_ /*34685*/;
assign _37778_ = _37779_ | _37781_ /*34682*/;
assign _37787_ = ~D[30] /*34681*/;
assign _37784_ = _37150_ & _37787_ /*34677*/;
assign _37785_ = _37150_ ^ _37787_ /*34680*/;
assign _37786_ = _37778_ & _37785_ /*34678*/;
assign _37599_ = _37778_ ^ _37785_ /*34679*/;
assign _37783_ = _37784_ | _37786_ /*34676*/;
assign _37792_ = ~D[31] /*34675*/;
assign _37789_ = _37151_ & _37792_ /*34671*/;
assign _37790_ = _37151_ ^ _37792_ /*34674*/;
assign _37791_ = _37783_ & _37790_ /*34672*/;
assign _37600_ = _37783_ ^ _37790_ /*34673*/;
assign _37788_ = _37789_ | _37791_ /*34670*/;
assign _37797_ = ~D[32] /*34669*/;
assign _37794_ = _37152_ & _37797_ /*34665*/;
assign _37795_ = _37152_ ^ _37797_ /*34668*/;
assign _37796_ = _37788_ & _37795_ /*34666*/;
assign _37601_ = _37788_ ^ _37795_ /*34667*/;
assign _37793_ = _37794_ | _37796_ /*34664*/;
assign _37802_ = ~D[33] /*34663*/;
assign _37799_ = _37153_ & _37802_ /*34659*/;
assign _37800_ = _37153_ ^ _37802_ /*34662*/;
assign _37801_ = _37793_ & _37800_ /*34660*/;
assign _37602_ = _37793_ ^ _37800_ /*34661*/;
assign _37798_ = _37799_ | _37801_ /*34658*/;
assign _37807_ = ~D[34] /*34657*/;
assign _37804_ = _37154_ & _37807_ /*34653*/;
assign _37805_ = _37154_ ^ _37807_ /*34656*/;
assign _37806_ = _37798_ & _37805_ /*34654*/;
assign _37603_ = _37798_ ^ _37805_ /*34655*/;
assign _37803_ = _37804_ | _37806_ /*34652*/;
assign _37812_ = ~D[35] /*34651*/;
assign _37809_ = _37155_ & _37812_ /*34647*/;
assign _37810_ = _37155_ ^ _37812_ /*34650*/;
assign _37811_ = _37803_ & _37810_ /*34648*/;
assign _37604_ = _37803_ ^ _37810_ /*34649*/;
assign _37808_ = _37809_ | _37811_ /*34646*/;
assign _37817_ = ~D[36] /*34645*/;
assign _37814_ = _37156_ & _37817_ /*34641*/;
assign _37815_ = _37156_ ^ _37817_ /*34644*/;
assign _37816_ = _37808_ & _37815_ /*34642*/;
assign _37605_ = _37808_ ^ _37815_ /*34643*/;
assign _37813_ = _37814_ | _37816_ /*34640*/;
assign _37822_ = ~D[37] /*34639*/;
assign _37819_ = _37157_ & _37822_ /*34635*/;
assign _37820_ = _37157_ ^ _37822_ /*34638*/;
assign _37821_ = _37813_ & _37820_ /*34636*/;
assign _37606_ = _37813_ ^ _37820_ /*34637*/;
assign _37818_ = _37819_ | _37821_ /*34634*/;
assign _37827_ = ~D[38] /*34633*/;
assign _37824_ = _37158_ & _37827_ /*34629*/;
assign _37825_ = _37158_ ^ _37827_ /*34632*/;
assign _37826_ = _37818_ & _37825_ /*34630*/;
assign _37607_ = _37818_ ^ _37825_ /*34631*/;
assign _37823_ = _37824_ | _37826_ /*34628*/;
assign _37832_ = ~D[39] /*34627*/;
assign _37829_ = _37159_ & _37832_ /*34623*/;
assign _37830_ = _37159_ ^ _37832_ /*34626*/;
assign _37831_ = _37823_ & _37830_ /*34624*/;
assign _37608_ = _37823_ ^ _37830_ /*34625*/;
assign _37828_ = _37829_ | _37831_ /*34622*/;
assign _37837_ = ~D[40] /*34621*/;
assign _37834_ = _37160_ & _37837_ /*34617*/;
assign _37835_ = _37160_ ^ _37837_ /*34620*/;
assign _37836_ = _37828_ & _37835_ /*34618*/;
assign _37609_ = _37828_ ^ _37835_ /*34619*/;
assign _37833_ = _37834_ | _37836_ /*34616*/;
assign _37842_ = ~D[41] /*34615*/;
assign _37839_ = _37161_ & _37842_ /*34611*/;
assign _37840_ = _37161_ ^ _37842_ /*34614*/;
assign _37841_ = _37833_ & _37840_ /*34612*/;
assign _37610_ = _37833_ ^ _37840_ /*34613*/;
assign _37838_ = _37839_ | _37841_ /*34610*/;
assign _37847_ = ~D[42] /*34609*/;
assign _37844_ = _37162_ & _37847_ /*34605*/;
assign _37845_ = _37162_ ^ _37847_ /*34608*/;
assign _37846_ = _37838_ & _37845_ /*34606*/;
assign _37611_ = _37838_ ^ _37845_ /*34607*/;
assign _37843_ = _37844_ | _37846_ /*34604*/;
assign _37852_ = ~D[43] /*34603*/;
assign _37849_ = _37163_ & _37852_ /*34599*/;
assign _37850_ = _37163_ ^ _37852_ /*34602*/;
assign _37851_ = _37843_ & _37850_ /*34600*/;
assign _37612_ = _37843_ ^ _37850_ /*34601*/;
assign _37848_ = _37849_ | _37851_ /*34598*/;
assign _37857_ = ~D[44] /*34597*/;
assign _37854_ = _37164_ & _37857_ /*34593*/;
assign _37855_ = _37164_ ^ _37857_ /*34596*/;
assign _37856_ = _37848_ & _37855_ /*34594*/;
assign _37613_ = _37848_ ^ _37855_ /*34595*/;
assign _37853_ = _37854_ | _37856_ /*34592*/;
assign _37862_ = ~D[45] /*34591*/;
assign _37859_ = _37165_ & _37862_ /*34587*/;
assign _37860_ = _37165_ ^ _37862_ /*34590*/;
assign _37861_ = _37853_ & _37860_ /*34588*/;
assign _37614_ = _37853_ ^ _37860_ /*34589*/;
assign _37858_ = _37859_ | _37861_ /*34586*/;
assign _37867_ = ~D[46] /*34585*/;
assign _37864_ = _37166_ & _37867_ /*34581*/;
assign _37865_ = _37166_ ^ _37867_ /*34584*/;
assign _37866_ = _37858_ & _37865_ /*34582*/;
assign _37615_ = _37858_ ^ _37865_ /*34583*/;
assign _37863_ = _37864_ | _37866_ /*34580*/;
assign _37872_ = ~D[47] /*34579*/;
assign _37869_ = _37167_ & _37872_ /*34575*/;
assign _37870_ = _37167_ ^ _37872_ /*34578*/;
assign _37871_ = _37863_ & _37870_ /*34576*/;
assign _37616_ = _37863_ ^ _37870_ /*34577*/;
assign _37868_ = _37869_ | _37871_ /*34574*/;
assign _37877_ = ~D[48] /*34573*/;
assign _37874_ = _37168_ & _37877_ /*34569*/;
assign _37875_ = _37168_ ^ _37877_ /*34572*/;
assign _37876_ = _37868_ & _37875_ /*34570*/;
assign _37617_ = _37868_ ^ _37875_ /*34571*/;
assign _37873_ = _37874_ | _37876_ /*34568*/;
assign _37882_ = ~D[49] /*34567*/;
assign _37879_ = _37169_ & _37882_ /*34563*/;
assign _37880_ = _37169_ ^ _37882_ /*34566*/;
assign _37881_ = _37873_ & _37880_ /*34564*/;
assign _37618_ = _37873_ ^ _37880_ /*34565*/;
assign _37878_ = _37879_ | _37881_ /*34562*/;
assign _37887_ = ~D[50] /*34561*/;
assign _37884_ = _37170_ & _37887_ /*34557*/;
assign _37885_ = _37170_ ^ _37887_ /*34560*/;
assign _37886_ = _37878_ & _37885_ /*34558*/;
assign _37619_ = _37878_ ^ _37885_ /*34559*/;
assign _37883_ = _37884_ | _37886_ /*34556*/;
assign _37892_ = ~D[51] /*34555*/;
assign _37889_ = _37171_ & _37892_ /*34551*/;
assign _37890_ = _37171_ ^ _37892_ /*34554*/;
assign _37891_ = _37883_ & _37890_ /*34552*/;
assign _37620_ = _37883_ ^ _37890_ /*34553*/;
assign _37888_ = _37889_ | _37891_ /*34550*/;
assign _37897_ = ~D[52] /*34549*/;
assign _37894_ = _37172_ & _37897_ /*34545*/;
assign _37895_ = _37172_ ^ _37897_ /*34548*/;
assign _37896_ = _37888_ & _37895_ /*34546*/;
assign _37621_ = _37888_ ^ _37895_ /*34547*/;
assign _37893_ = _37894_ | _37896_ /*34544*/;
assign _37902_ = ~D[53] /*34543*/;
assign _37899_ = _37173_ & _37902_ /*34539*/;
assign _37900_ = _37173_ ^ _37902_ /*34542*/;
assign _37901_ = _37893_ & _37900_ /*34540*/;
assign _37622_ = _37893_ ^ _37900_ /*34541*/;
assign _37898_ = _37899_ | _37901_ /*34538*/;
assign _37907_ = ~D[54] /*34537*/;
assign _37904_ = _37174_ & _37907_ /*34533*/;
assign _37905_ = _37174_ ^ _37907_ /*34536*/;
assign _37906_ = _37898_ & _37905_ /*34534*/;
assign _37623_ = _37898_ ^ _37905_ /*34535*/;
assign _37903_ = _37904_ | _37906_ /*34532*/;
assign _37912_ = ~D[55] /*34531*/;
assign _37909_ = _37175_ & _37912_ /*34527*/;
assign _37910_ = _37175_ ^ _37912_ /*34530*/;
assign _37911_ = _37903_ & _37910_ /*34528*/;
assign _37624_ = _37903_ ^ _37910_ /*34529*/;
assign _37908_ = _37909_ | _37911_ /*34526*/;
assign _37917_ = ~D[56] /*34525*/;
assign _37914_ = _37176_ & _37917_ /*34521*/;
assign _37915_ = _37176_ ^ _37917_ /*34524*/;
assign _37916_ = _37908_ & _37915_ /*34522*/;
assign _37625_ = _37908_ ^ _37915_ /*34523*/;
assign _37913_ = _37914_ | _37916_ /*34520*/;
assign _37922_ = ~D[57] /*34519*/;
assign _37919_ = _37177_ & _37922_ /*34515*/;
assign _37920_ = _37177_ ^ _37922_ /*34518*/;
assign _37921_ = _37913_ & _37920_ /*34516*/;
assign _37626_ = _37913_ ^ _37920_ /*34517*/;
assign _37918_ = _37919_ | _37921_ /*34514*/;
assign _37927_ = ~D[58] /*34513*/;
assign _37924_ = _37178_ & _37927_ /*34509*/;
assign _37925_ = _37178_ ^ _37927_ /*34512*/;
assign _37926_ = _37918_ & _37925_ /*34510*/;
assign _37627_ = _37918_ ^ _37925_ /*34511*/;
assign _37923_ = _37924_ | _37926_ /*34508*/;
assign _37932_ = ~D[59] /*34507*/;
assign _37929_ = _37179_ & _37932_ /*34503*/;
assign _37930_ = _37179_ ^ _37932_ /*34506*/;
assign _37931_ = _37923_ & _37930_ /*34504*/;
assign _37628_ = _37923_ ^ _37930_ /*34505*/;
assign _37928_ = _37929_ | _37931_ /*34502*/;
assign _37937_ = ~D[60] /*34501*/;
assign _37934_ = _37180_ & _37937_ /*34497*/;
assign _37935_ = _37180_ ^ _37937_ /*34500*/;
assign _37936_ = _37928_ & _37935_ /*34498*/;
assign _37629_ = _37928_ ^ _37935_ /*34499*/;
assign _37933_ = _37934_ | _37936_ /*34496*/;
assign _37942_ = ~D[61] /*34495*/;
assign _37939_ = _37181_ & _37942_ /*34491*/;
assign _37940_ = _37181_ ^ _37942_ /*34494*/;
assign _37941_ = _37933_ & _37940_ /*34492*/;
assign _37630_ = _37933_ ^ _37940_ /*34493*/;
assign _37938_ = _37939_ | _37941_ /*34490*/;
assign _37947_ = ~D[62] /*34489*/;
assign _37944_ = _37182_ & _37947_ /*34485*/;
assign _37945_ = _37182_ ^ _37947_ /*34488*/;
assign _37946_ = _37938_ & _37945_ /*34486*/;
assign _37631_ = _37938_ ^ _37945_ /*34487*/;
assign _37943_ = _37944_ | _37946_ /*34484*/;
assign _37948_ = _37183_ & oneWire /*34479*/;
assign _37949_ = _37183_ ^ oneWire /*34482*/;
assign _37950_ = _37943_ & _37949_ /*34480*/;
assign _37632_ = _37943_ ^ _37949_ /*34481*/;
assign Q[21] = _37948_ | _37950_ /*34478*/;
assign _38083_ = ~Q[21] /*34093*/;
assign _38082_ = _38083_ & D[0] /*34092*/;
assign _38085_ = _37569_ & _38082_ /*34087*/;
assign _38086_ = _37569_ ^ _38082_ /*34090*/;
assign _38087_ = zeroWire & _38086_ /*34088*/;
assign _38017_ = zeroWire ^ _38086_ /*34089*/;
assign _38084_ = _38085_ | _38087_ /*34086*/;
assign _38089_ = ~Q[21] /*34085*/;
assign _38088_ = _38089_ & D[1] /*34084*/;
assign _38091_ = _37570_ & _38088_ /*34079*/;
assign _38092_ = _37570_ ^ _38088_ /*34082*/;
assign _38093_ = _38084_ & _38092_ /*34080*/;
assign _38018_ = _38084_ ^ _38092_ /*34081*/;
assign _38090_ = _38091_ | _38093_ /*34078*/;
assign _38095_ = ~Q[21] /*34077*/;
assign _38094_ = _38095_ & D[2] /*34076*/;
assign _38097_ = _37571_ & _38094_ /*34071*/;
assign _38098_ = _37571_ ^ _38094_ /*34074*/;
assign _38099_ = _38090_ & _38098_ /*34072*/;
assign _38019_ = _38090_ ^ _38098_ /*34073*/;
assign _38096_ = _38097_ | _38099_ /*34070*/;
assign _38101_ = ~Q[21] /*34069*/;
assign _38100_ = _38101_ & D[3] /*34068*/;
assign _38103_ = _37572_ & _38100_ /*34063*/;
assign _38104_ = _37572_ ^ _38100_ /*34066*/;
assign _38105_ = _38096_ & _38104_ /*34064*/;
assign _38020_ = _38096_ ^ _38104_ /*34065*/;
assign _38102_ = _38103_ | _38105_ /*34062*/;
assign _38107_ = ~Q[21] /*34061*/;
assign _38106_ = _38107_ & D[4] /*34060*/;
assign _38109_ = _37573_ & _38106_ /*34055*/;
assign _38110_ = _37573_ ^ _38106_ /*34058*/;
assign _38111_ = _38102_ & _38110_ /*34056*/;
assign _38021_ = _38102_ ^ _38110_ /*34057*/;
assign _38108_ = _38109_ | _38111_ /*34054*/;
assign _38113_ = ~Q[21] /*34053*/;
assign _38112_ = _38113_ & D[5] /*34052*/;
assign _38115_ = _37574_ & _38112_ /*34047*/;
assign _38116_ = _37574_ ^ _38112_ /*34050*/;
assign _38117_ = _38108_ & _38116_ /*34048*/;
assign _38022_ = _38108_ ^ _38116_ /*34049*/;
assign _38114_ = _38115_ | _38117_ /*34046*/;
assign _38119_ = ~Q[21] /*34045*/;
assign _38118_ = _38119_ & D[6] /*34044*/;
assign _38121_ = _37575_ & _38118_ /*34039*/;
assign _38122_ = _37575_ ^ _38118_ /*34042*/;
assign _38123_ = _38114_ & _38122_ /*34040*/;
assign _38023_ = _38114_ ^ _38122_ /*34041*/;
assign _38120_ = _38121_ | _38123_ /*34038*/;
assign _38125_ = ~Q[21] /*34037*/;
assign _38124_ = _38125_ & D[7] /*34036*/;
assign _38127_ = _37576_ & _38124_ /*34031*/;
assign _38128_ = _37576_ ^ _38124_ /*34034*/;
assign _38129_ = _38120_ & _38128_ /*34032*/;
assign _38024_ = _38120_ ^ _38128_ /*34033*/;
assign _38126_ = _38127_ | _38129_ /*34030*/;
assign _38131_ = ~Q[21] /*34029*/;
assign _38130_ = _38131_ & D[8] /*34028*/;
assign _38133_ = _37577_ & _38130_ /*34023*/;
assign _38134_ = _37577_ ^ _38130_ /*34026*/;
assign _38135_ = _38126_ & _38134_ /*34024*/;
assign _38025_ = _38126_ ^ _38134_ /*34025*/;
assign _38132_ = _38133_ | _38135_ /*34022*/;
assign _38137_ = ~Q[21] /*34021*/;
assign _38136_ = _38137_ & D[9] /*34020*/;
assign _38139_ = _37578_ & _38136_ /*34015*/;
assign _38140_ = _37578_ ^ _38136_ /*34018*/;
assign _38141_ = _38132_ & _38140_ /*34016*/;
assign _38026_ = _38132_ ^ _38140_ /*34017*/;
assign _38138_ = _38139_ | _38141_ /*34014*/;
assign _38143_ = ~Q[21] /*34013*/;
assign _38142_ = _38143_ & D[10] /*34012*/;
assign _38145_ = _37579_ & _38142_ /*34007*/;
assign _38146_ = _37579_ ^ _38142_ /*34010*/;
assign _38147_ = _38138_ & _38146_ /*34008*/;
assign _38027_ = _38138_ ^ _38146_ /*34009*/;
assign _38144_ = _38145_ | _38147_ /*34006*/;
assign _38149_ = ~Q[21] /*34005*/;
assign _38148_ = _38149_ & D[11] /*34004*/;
assign _38151_ = _37580_ & _38148_ /*33999*/;
assign _38152_ = _37580_ ^ _38148_ /*34002*/;
assign _38153_ = _38144_ & _38152_ /*34000*/;
assign _38028_ = _38144_ ^ _38152_ /*34001*/;
assign _38150_ = _38151_ | _38153_ /*33998*/;
assign _38155_ = ~Q[21] /*33997*/;
assign _38154_ = _38155_ & D[12] /*33996*/;
assign _38157_ = _37581_ & _38154_ /*33991*/;
assign _38158_ = _37581_ ^ _38154_ /*33994*/;
assign _38159_ = _38150_ & _38158_ /*33992*/;
assign _38029_ = _38150_ ^ _38158_ /*33993*/;
assign _38156_ = _38157_ | _38159_ /*33990*/;
assign _38161_ = ~Q[21] /*33989*/;
assign _38160_ = _38161_ & D[13] /*33988*/;
assign _38163_ = _37582_ & _38160_ /*33983*/;
assign _38164_ = _37582_ ^ _38160_ /*33986*/;
assign _38165_ = _38156_ & _38164_ /*33984*/;
assign _38030_ = _38156_ ^ _38164_ /*33985*/;
assign _38162_ = _38163_ | _38165_ /*33982*/;
assign _38167_ = ~Q[21] /*33981*/;
assign _38166_ = _38167_ & D[14] /*33980*/;
assign _38169_ = _37583_ & _38166_ /*33975*/;
assign _38170_ = _37583_ ^ _38166_ /*33978*/;
assign _38171_ = _38162_ & _38170_ /*33976*/;
assign _38031_ = _38162_ ^ _38170_ /*33977*/;
assign _38168_ = _38169_ | _38171_ /*33974*/;
assign _38173_ = ~Q[21] /*33973*/;
assign _38172_ = _38173_ & D[15] /*33972*/;
assign _38175_ = _37584_ & _38172_ /*33967*/;
assign _38176_ = _37584_ ^ _38172_ /*33970*/;
assign _38177_ = _38168_ & _38176_ /*33968*/;
assign _38032_ = _38168_ ^ _38176_ /*33969*/;
assign _38174_ = _38175_ | _38177_ /*33966*/;
assign _38179_ = ~Q[21] /*33965*/;
assign _38178_ = _38179_ & D[16] /*33964*/;
assign _38181_ = _37585_ & _38178_ /*33959*/;
assign _38182_ = _37585_ ^ _38178_ /*33962*/;
assign _38183_ = _38174_ & _38182_ /*33960*/;
assign _38033_ = _38174_ ^ _38182_ /*33961*/;
assign _38180_ = _38181_ | _38183_ /*33958*/;
assign _38185_ = ~Q[21] /*33957*/;
assign _38184_ = _38185_ & D[17] /*33956*/;
assign _38187_ = _37586_ & _38184_ /*33951*/;
assign _38188_ = _37586_ ^ _38184_ /*33954*/;
assign _38189_ = _38180_ & _38188_ /*33952*/;
assign _38034_ = _38180_ ^ _38188_ /*33953*/;
assign _38186_ = _38187_ | _38189_ /*33950*/;
assign _38191_ = ~Q[21] /*33949*/;
assign _38190_ = _38191_ & D[18] /*33948*/;
assign _38193_ = _37587_ & _38190_ /*33943*/;
assign _38194_ = _37587_ ^ _38190_ /*33946*/;
assign _38195_ = _38186_ & _38194_ /*33944*/;
assign _38035_ = _38186_ ^ _38194_ /*33945*/;
assign _38192_ = _38193_ | _38195_ /*33942*/;
assign _38197_ = ~Q[21] /*33941*/;
assign _38196_ = _38197_ & D[19] /*33940*/;
assign _38199_ = _37588_ & _38196_ /*33935*/;
assign _38200_ = _37588_ ^ _38196_ /*33938*/;
assign _38201_ = _38192_ & _38200_ /*33936*/;
assign _38036_ = _38192_ ^ _38200_ /*33937*/;
assign _38198_ = _38199_ | _38201_ /*33934*/;
assign _38203_ = ~Q[21] /*33933*/;
assign _38202_ = _38203_ & D[20] /*33932*/;
assign _38205_ = _37589_ & _38202_ /*33927*/;
assign _38206_ = _37589_ ^ _38202_ /*33930*/;
assign _38207_ = _38198_ & _38206_ /*33928*/;
assign _38037_ = _38198_ ^ _38206_ /*33929*/;
assign _38204_ = _38205_ | _38207_ /*33926*/;
assign _38209_ = ~Q[21] /*33925*/;
assign _38208_ = _38209_ & D[21] /*33924*/;
assign _38211_ = _37590_ & _38208_ /*33919*/;
assign _38212_ = _37590_ ^ _38208_ /*33922*/;
assign _38213_ = _38204_ & _38212_ /*33920*/;
assign _38038_ = _38204_ ^ _38212_ /*33921*/;
assign _38210_ = _38211_ | _38213_ /*33918*/;
assign _38215_ = ~Q[21] /*33917*/;
assign _38214_ = _38215_ & D[22] /*33916*/;
assign _38217_ = _37591_ & _38214_ /*33911*/;
assign _38218_ = _37591_ ^ _38214_ /*33914*/;
assign _38219_ = _38210_ & _38218_ /*33912*/;
assign _38039_ = _38210_ ^ _38218_ /*33913*/;
assign _38216_ = _38217_ | _38219_ /*33910*/;
assign _38221_ = ~Q[21] /*33909*/;
assign _38220_ = _38221_ & D[23] /*33908*/;
assign _38223_ = _37592_ & _38220_ /*33903*/;
assign _38224_ = _37592_ ^ _38220_ /*33906*/;
assign _38225_ = _38216_ & _38224_ /*33904*/;
assign _38040_ = _38216_ ^ _38224_ /*33905*/;
assign _38222_ = _38223_ | _38225_ /*33902*/;
assign _38227_ = ~Q[21] /*33901*/;
assign _38226_ = _38227_ & D[24] /*33900*/;
assign _38229_ = _37593_ & _38226_ /*33895*/;
assign _38230_ = _37593_ ^ _38226_ /*33898*/;
assign _38231_ = _38222_ & _38230_ /*33896*/;
assign _38041_ = _38222_ ^ _38230_ /*33897*/;
assign _38228_ = _38229_ | _38231_ /*33894*/;
assign _38233_ = ~Q[21] /*33893*/;
assign _38232_ = _38233_ & D[25] /*33892*/;
assign _38235_ = _37594_ & _38232_ /*33887*/;
assign _38236_ = _37594_ ^ _38232_ /*33890*/;
assign _38237_ = _38228_ & _38236_ /*33888*/;
assign _38042_ = _38228_ ^ _38236_ /*33889*/;
assign _38234_ = _38235_ | _38237_ /*33886*/;
assign _38239_ = ~Q[21] /*33885*/;
assign _38238_ = _38239_ & D[26] /*33884*/;
assign _38241_ = _37595_ & _38238_ /*33879*/;
assign _38242_ = _37595_ ^ _38238_ /*33882*/;
assign _38243_ = _38234_ & _38242_ /*33880*/;
assign _38043_ = _38234_ ^ _38242_ /*33881*/;
assign _38240_ = _38241_ | _38243_ /*33878*/;
assign _38245_ = ~Q[21] /*33877*/;
assign _38244_ = _38245_ & D[27] /*33876*/;
assign _38247_ = _37596_ & _38244_ /*33871*/;
assign _38248_ = _37596_ ^ _38244_ /*33874*/;
assign _38249_ = _38240_ & _38248_ /*33872*/;
assign _38044_ = _38240_ ^ _38248_ /*33873*/;
assign _38246_ = _38247_ | _38249_ /*33870*/;
assign _38251_ = ~Q[21] /*33869*/;
assign _38250_ = _38251_ & D[28] /*33868*/;
assign _38253_ = _37597_ & _38250_ /*33863*/;
assign _38254_ = _37597_ ^ _38250_ /*33866*/;
assign _38255_ = _38246_ & _38254_ /*33864*/;
assign _38045_ = _38246_ ^ _38254_ /*33865*/;
assign _38252_ = _38253_ | _38255_ /*33862*/;
assign _38257_ = ~Q[21] /*33861*/;
assign _38256_ = _38257_ & D[29] /*33860*/;
assign _38259_ = _37598_ & _38256_ /*33855*/;
assign _38260_ = _37598_ ^ _38256_ /*33858*/;
assign _38261_ = _38252_ & _38260_ /*33856*/;
assign _38046_ = _38252_ ^ _38260_ /*33857*/;
assign _38258_ = _38259_ | _38261_ /*33854*/;
assign _38263_ = ~Q[21] /*33853*/;
assign _38262_ = _38263_ & D[30] /*33852*/;
assign _38265_ = _37599_ & _38262_ /*33847*/;
assign _38266_ = _37599_ ^ _38262_ /*33850*/;
assign _38267_ = _38258_ & _38266_ /*33848*/;
assign _38047_ = _38258_ ^ _38266_ /*33849*/;
assign _38264_ = _38265_ | _38267_ /*33846*/;
assign _38269_ = ~Q[21] /*33845*/;
assign _38268_ = _38269_ & D[31] /*33844*/;
assign _38271_ = _37600_ & _38268_ /*33839*/;
assign _38272_ = _37600_ ^ _38268_ /*33842*/;
assign _38273_ = _38264_ & _38272_ /*33840*/;
assign _38048_ = _38264_ ^ _38272_ /*33841*/;
assign _38270_ = _38271_ | _38273_ /*33838*/;
assign _38275_ = ~Q[21] /*33837*/;
assign _38274_ = _38275_ & D[32] /*33836*/;
assign _38277_ = _37601_ & _38274_ /*33831*/;
assign _38278_ = _37601_ ^ _38274_ /*33834*/;
assign _38279_ = _38270_ & _38278_ /*33832*/;
assign _38049_ = _38270_ ^ _38278_ /*33833*/;
assign _38276_ = _38277_ | _38279_ /*33830*/;
assign _38281_ = ~Q[21] /*33829*/;
assign _38280_ = _38281_ & D[33] /*33828*/;
assign _38283_ = _37602_ & _38280_ /*33823*/;
assign _38284_ = _37602_ ^ _38280_ /*33826*/;
assign _38285_ = _38276_ & _38284_ /*33824*/;
assign _38050_ = _38276_ ^ _38284_ /*33825*/;
assign _38282_ = _38283_ | _38285_ /*33822*/;
assign _38287_ = ~Q[21] /*33821*/;
assign _38286_ = _38287_ & D[34] /*33820*/;
assign _38289_ = _37603_ & _38286_ /*33815*/;
assign _38290_ = _37603_ ^ _38286_ /*33818*/;
assign _38291_ = _38282_ & _38290_ /*33816*/;
assign _38051_ = _38282_ ^ _38290_ /*33817*/;
assign _38288_ = _38289_ | _38291_ /*33814*/;
assign _38293_ = ~Q[21] /*33813*/;
assign _38292_ = _38293_ & D[35] /*33812*/;
assign _38295_ = _37604_ & _38292_ /*33807*/;
assign _38296_ = _37604_ ^ _38292_ /*33810*/;
assign _38297_ = _38288_ & _38296_ /*33808*/;
assign _38052_ = _38288_ ^ _38296_ /*33809*/;
assign _38294_ = _38295_ | _38297_ /*33806*/;
assign _38299_ = ~Q[21] /*33805*/;
assign _38298_ = _38299_ & D[36] /*33804*/;
assign _38301_ = _37605_ & _38298_ /*33799*/;
assign _38302_ = _37605_ ^ _38298_ /*33802*/;
assign _38303_ = _38294_ & _38302_ /*33800*/;
assign _38053_ = _38294_ ^ _38302_ /*33801*/;
assign _38300_ = _38301_ | _38303_ /*33798*/;
assign _38305_ = ~Q[21] /*33797*/;
assign _38304_ = _38305_ & D[37] /*33796*/;
assign _38307_ = _37606_ & _38304_ /*33791*/;
assign _38308_ = _37606_ ^ _38304_ /*33794*/;
assign _38309_ = _38300_ & _38308_ /*33792*/;
assign _38054_ = _38300_ ^ _38308_ /*33793*/;
assign _38306_ = _38307_ | _38309_ /*33790*/;
assign _38311_ = ~Q[21] /*33789*/;
assign _38310_ = _38311_ & D[38] /*33788*/;
assign _38313_ = _37607_ & _38310_ /*33783*/;
assign _38314_ = _37607_ ^ _38310_ /*33786*/;
assign _38315_ = _38306_ & _38314_ /*33784*/;
assign _38055_ = _38306_ ^ _38314_ /*33785*/;
assign _38312_ = _38313_ | _38315_ /*33782*/;
assign _38317_ = ~Q[21] /*33781*/;
assign _38316_ = _38317_ & D[39] /*33780*/;
assign _38319_ = _37608_ & _38316_ /*33775*/;
assign _38320_ = _37608_ ^ _38316_ /*33778*/;
assign _38321_ = _38312_ & _38320_ /*33776*/;
assign _38056_ = _38312_ ^ _38320_ /*33777*/;
assign _38318_ = _38319_ | _38321_ /*33774*/;
assign _38323_ = ~Q[21] /*33773*/;
assign _38322_ = _38323_ & D[40] /*33772*/;
assign _38325_ = _37609_ & _38322_ /*33767*/;
assign _38326_ = _37609_ ^ _38322_ /*33770*/;
assign _38327_ = _38318_ & _38326_ /*33768*/;
assign _38057_ = _38318_ ^ _38326_ /*33769*/;
assign _38324_ = _38325_ | _38327_ /*33766*/;
assign _38329_ = ~Q[21] /*33765*/;
assign _38328_ = _38329_ & D[41] /*33764*/;
assign _38331_ = _37610_ & _38328_ /*33759*/;
assign _38332_ = _37610_ ^ _38328_ /*33762*/;
assign _38333_ = _38324_ & _38332_ /*33760*/;
assign _38058_ = _38324_ ^ _38332_ /*33761*/;
assign _38330_ = _38331_ | _38333_ /*33758*/;
assign _38335_ = ~Q[21] /*33757*/;
assign _38334_ = _38335_ & D[42] /*33756*/;
assign _38337_ = _37611_ & _38334_ /*33751*/;
assign _38338_ = _37611_ ^ _38334_ /*33754*/;
assign _38339_ = _38330_ & _38338_ /*33752*/;
assign _38059_ = _38330_ ^ _38338_ /*33753*/;
assign _38336_ = _38337_ | _38339_ /*33750*/;
assign _38341_ = ~Q[21] /*33749*/;
assign _38340_ = _38341_ & D[43] /*33748*/;
assign _38343_ = _37612_ & _38340_ /*33743*/;
assign _38344_ = _37612_ ^ _38340_ /*33746*/;
assign _38345_ = _38336_ & _38344_ /*33744*/;
assign _38060_ = _38336_ ^ _38344_ /*33745*/;
assign _38342_ = _38343_ | _38345_ /*33742*/;
assign _38347_ = ~Q[21] /*33741*/;
assign _38346_ = _38347_ & D[44] /*33740*/;
assign _38349_ = _37613_ & _38346_ /*33735*/;
assign _38350_ = _37613_ ^ _38346_ /*33738*/;
assign _38351_ = _38342_ & _38350_ /*33736*/;
assign _38061_ = _38342_ ^ _38350_ /*33737*/;
assign _38348_ = _38349_ | _38351_ /*33734*/;
assign _38353_ = ~Q[21] /*33733*/;
assign _38352_ = _38353_ & D[45] /*33732*/;
assign _38355_ = _37614_ & _38352_ /*33727*/;
assign _38356_ = _37614_ ^ _38352_ /*33730*/;
assign _38357_ = _38348_ & _38356_ /*33728*/;
assign _38062_ = _38348_ ^ _38356_ /*33729*/;
assign _38354_ = _38355_ | _38357_ /*33726*/;
assign _38359_ = ~Q[21] /*33725*/;
assign _38358_ = _38359_ & D[46] /*33724*/;
assign _38361_ = _37615_ & _38358_ /*33719*/;
assign _38362_ = _37615_ ^ _38358_ /*33722*/;
assign _38363_ = _38354_ & _38362_ /*33720*/;
assign _38063_ = _38354_ ^ _38362_ /*33721*/;
assign _38360_ = _38361_ | _38363_ /*33718*/;
assign _38365_ = ~Q[21] /*33717*/;
assign _38364_ = _38365_ & D[47] /*33716*/;
assign _38367_ = _37616_ & _38364_ /*33711*/;
assign _38368_ = _37616_ ^ _38364_ /*33714*/;
assign _38369_ = _38360_ & _38368_ /*33712*/;
assign _38064_ = _38360_ ^ _38368_ /*33713*/;
assign _38366_ = _38367_ | _38369_ /*33710*/;
assign _38371_ = ~Q[21] /*33709*/;
assign _38370_ = _38371_ & D[48] /*33708*/;
assign _38373_ = _37617_ & _38370_ /*33703*/;
assign _38374_ = _37617_ ^ _38370_ /*33706*/;
assign _38375_ = _38366_ & _38374_ /*33704*/;
assign _38065_ = _38366_ ^ _38374_ /*33705*/;
assign _38372_ = _38373_ | _38375_ /*33702*/;
assign _38377_ = ~Q[21] /*33701*/;
assign _38376_ = _38377_ & D[49] /*33700*/;
assign _38379_ = _37618_ & _38376_ /*33695*/;
assign _38380_ = _37618_ ^ _38376_ /*33698*/;
assign _38381_ = _38372_ & _38380_ /*33696*/;
assign _38066_ = _38372_ ^ _38380_ /*33697*/;
assign _38378_ = _38379_ | _38381_ /*33694*/;
assign _38383_ = ~Q[21] /*33693*/;
assign _38382_ = _38383_ & D[50] /*33692*/;
assign _38385_ = _37619_ & _38382_ /*33687*/;
assign _38386_ = _37619_ ^ _38382_ /*33690*/;
assign _38387_ = _38378_ & _38386_ /*33688*/;
assign _38067_ = _38378_ ^ _38386_ /*33689*/;
assign _38384_ = _38385_ | _38387_ /*33686*/;
assign _38389_ = ~Q[21] /*33685*/;
assign _38388_ = _38389_ & D[51] /*33684*/;
assign _38391_ = _37620_ & _38388_ /*33679*/;
assign _38392_ = _37620_ ^ _38388_ /*33682*/;
assign _38393_ = _38384_ & _38392_ /*33680*/;
assign _38068_ = _38384_ ^ _38392_ /*33681*/;
assign _38390_ = _38391_ | _38393_ /*33678*/;
assign _38395_ = ~Q[21] /*33677*/;
assign _38394_ = _38395_ & D[52] /*33676*/;
assign _38397_ = _37621_ & _38394_ /*33671*/;
assign _38398_ = _37621_ ^ _38394_ /*33674*/;
assign _38399_ = _38390_ & _38398_ /*33672*/;
assign _38069_ = _38390_ ^ _38398_ /*33673*/;
assign _38396_ = _38397_ | _38399_ /*33670*/;
assign _38401_ = ~Q[21] /*33669*/;
assign _38400_ = _38401_ & D[53] /*33668*/;
assign _38403_ = _37622_ & _38400_ /*33663*/;
assign _38404_ = _37622_ ^ _38400_ /*33666*/;
assign _38405_ = _38396_ & _38404_ /*33664*/;
assign _38070_ = _38396_ ^ _38404_ /*33665*/;
assign _38402_ = _38403_ | _38405_ /*33662*/;
assign _38407_ = ~Q[21] /*33661*/;
assign _38406_ = _38407_ & D[54] /*33660*/;
assign _38409_ = _37623_ & _38406_ /*33655*/;
assign _38410_ = _37623_ ^ _38406_ /*33658*/;
assign _38411_ = _38402_ & _38410_ /*33656*/;
assign _38071_ = _38402_ ^ _38410_ /*33657*/;
assign _38408_ = _38409_ | _38411_ /*33654*/;
assign _38413_ = ~Q[21] /*33653*/;
assign _38412_ = _38413_ & D[55] /*33652*/;
assign _38415_ = _37624_ & _38412_ /*33647*/;
assign _38416_ = _37624_ ^ _38412_ /*33650*/;
assign _38417_ = _38408_ & _38416_ /*33648*/;
assign _38072_ = _38408_ ^ _38416_ /*33649*/;
assign _38414_ = _38415_ | _38417_ /*33646*/;
assign _38419_ = ~Q[21] /*33645*/;
assign _38418_ = _38419_ & D[56] /*33644*/;
assign _38421_ = _37625_ & _38418_ /*33639*/;
assign _38422_ = _37625_ ^ _38418_ /*33642*/;
assign _38423_ = _38414_ & _38422_ /*33640*/;
assign _38073_ = _38414_ ^ _38422_ /*33641*/;
assign _38420_ = _38421_ | _38423_ /*33638*/;
assign _38425_ = ~Q[21] /*33637*/;
assign _38424_ = _38425_ & D[57] /*33636*/;
assign _38427_ = _37626_ & _38424_ /*33631*/;
assign _38428_ = _37626_ ^ _38424_ /*33634*/;
assign _38429_ = _38420_ & _38428_ /*33632*/;
assign _38074_ = _38420_ ^ _38428_ /*33633*/;
assign _38426_ = _38427_ | _38429_ /*33630*/;
assign _38431_ = ~Q[21] /*33629*/;
assign _38430_ = _38431_ & D[58] /*33628*/;
assign _38433_ = _37627_ & _38430_ /*33623*/;
assign _38434_ = _37627_ ^ _38430_ /*33626*/;
assign _38435_ = _38426_ & _38434_ /*33624*/;
assign _38075_ = _38426_ ^ _38434_ /*33625*/;
assign _38432_ = _38433_ | _38435_ /*33622*/;
assign _38437_ = ~Q[21] /*33621*/;
assign _38436_ = _38437_ & D[59] /*33620*/;
assign _38439_ = _37628_ & _38436_ /*33615*/;
assign _38440_ = _37628_ ^ _38436_ /*33618*/;
assign _38441_ = _38432_ & _38440_ /*33616*/;
assign _38076_ = _38432_ ^ _38440_ /*33617*/;
assign _38438_ = _38439_ | _38441_ /*33614*/;
assign _38443_ = ~Q[21] /*33613*/;
assign _38442_ = _38443_ & D[60] /*33612*/;
assign _38445_ = _37629_ & _38442_ /*33607*/;
assign _38446_ = _37629_ ^ _38442_ /*33610*/;
assign _38447_ = _38438_ & _38446_ /*33608*/;
assign _38077_ = _38438_ ^ _38446_ /*33609*/;
assign _38444_ = _38445_ | _38447_ /*33606*/;
assign _38449_ = ~Q[21] /*33605*/;
assign _38448_ = _38449_ & D[61] /*33604*/;
assign _38451_ = _37630_ & _38448_ /*33599*/;
assign _38452_ = _37630_ ^ _38448_ /*33602*/;
assign _38453_ = _38444_ & _38452_ /*33600*/;
assign _38078_ = _38444_ ^ _38452_ /*33601*/;
assign _38450_ = _38451_ | _38453_ /*33598*/;
assign _38455_ = ~Q[21] /*33597*/;
assign _38454_ = _38455_ & D[62] /*33596*/;
assign _38457_ = _37631_ & _38454_ /*33591*/;
assign _38458_ = _37631_ ^ _38454_ /*33594*/;
assign _38459_ = _38450_ & _38458_ /*33592*/;
assign _38079_ = _38450_ ^ _38458_ /*33593*/;
assign _38456_ = _38457_ | _38459_ /*33590*/;
assign _38461_ = ~Q[21] /*33589*/;
assign _38460_ = _38461_ & zeroWire /*33588*/;
assign _38462_ = _37632_ ^ _38460_ /*33586*/;
assign _38080_ = _38462_ ^ _38456_ /*33585*/;
assign _38533_ = ~D[0] /*33331*/;
assign _38530_ = R_0[20] & _38533_ /*33327*/;
assign _38531_ = R_0[20] ^ _38533_ /*33330*/;
assign _38532_ = oneWire & _38531_ /*33328*/;
assign _38465_ = oneWire ^ _38531_ /*33329*/;
assign _38529_ = _38530_ | _38532_ /*33326*/;
assign _38538_ = ~D[1] /*33325*/;
assign _38535_ = _38017_ & _38538_ /*33321*/;
assign _38536_ = _38017_ ^ _38538_ /*33324*/;
assign _38537_ = _38529_ & _38536_ /*33322*/;
assign _38466_ = _38529_ ^ _38536_ /*33323*/;
assign _38534_ = _38535_ | _38537_ /*33320*/;
assign _38543_ = ~D[2] /*33319*/;
assign _38540_ = _38018_ & _38543_ /*33315*/;
assign _38541_ = _38018_ ^ _38543_ /*33318*/;
assign _38542_ = _38534_ & _38541_ /*33316*/;
assign _38467_ = _38534_ ^ _38541_ /*33317*/;
assign _38539_ = _38540_ | _38542_ /*33314*/;
assign _38548_ = ~D[3] /*33313*/;
assign _38545_ = _38019_ & _38548_ /*33309*/;
assign _38546_ = _38019_ ^ _38548_ /*33312*/;
assign _38547_ = _38539_ & _38546_ /*33310*/;
assign _38468_ = _38539_ ^ _38546_ /*33311*/;
assign _38544_ = _38545_ | _38547_ /*33308*/;
assign _38553_ = ~D[4] /*33307*/;
assign _38550_ = _38020_ & _38553_ /*33303*/;
assign _38551_ = _38020_ ^ _38553_ /*33306*/;
assign _38552_ = _38544_ & _38551_ /*33304*/;
assign _38469_ = _38544_ ^ _38551_ /*33305*/;
assign _38549_ = _38550_ | _38552_ /*33302*/;
assign _38558_ = ~D[5] /*33301*/;
assign _38555_ = _38021_ & _38558_ /*33297*/;
assign _38556_ = _38021_ ^ _38558_ /*33300*/;
assign _38557_ = _38549_ & _38556_ /*33298*/;
assign _38470_ = _38549_ ^ _38556_ /*33299*/;
assign _38554_ = _38555_ | _38557_ /*33296*/;
assign _38563_ = ~D[6] /*33295*/;
assign _38560_ = _38022_ & _38563_ /*33291*/;
assign _38561_ = _38022_ ^ _38563_ /*33294*/;
assign _38562_ = _38554_ & _38561_ /*33292*/;
assign _38471_ = _38554_ ^ _38561_ /*33293*/;
assign _38559_ = _38560_ | _38562_ /*33290*/;
assign _38568_ = ~D[7] /*33289*/;
assign _38565_ = _38023_ & _38568_ /*33285*/;
assign _38566_ = _38023_ ^ _38568_ /*33288*/;
assign _38567_ = _38559_ & _38566_ /*33286*/;
assign _38472_ = _38559_ ^ _38566_ /*33287*/;
assign _38564_ = _38565_ | _38567_ /*33284*/;
assign _38573_ = ~D[8] /*33283*/;
assign _38570_ = _38024_ & _38573_ /*33279*/;
assign _38571_ = _38024_ ^ _38573_ /*33282*/;
assign _38572_ = _38564_ & _38571_ /*33280*/;
assign _38473_ = _38564_ ^ _38571_ /*33281*/;
assign _38569_ = _38570_ | _38572_ /*33278*/;
assign _38578_ = ~D[9] /*33277*/;
assign _38575_ = _38025_ & _38578_ /*33273*/;
assign _38576_ = _38025_ ^ _38578_ /*33276*/;
assign _38577_ = _38569_ & _38576_ /*33274*/;
assign _38474_ = _38569_ ^ _38576_ /*33275*/;
assign _38574_ = _38575_ | _38577_ /*33272*/;
assign _38583_ = ~D[10] /*33271*/;
assign _38580_ = _38026_ & _38583_ /*33267*/;
assign _38581_ = _38026_ ^ _38583_ /*33270*/;
assign _38582_ = _38574_ & _38581_ /*33268*/;
assign _38475_ = _38574_ ^ _38581_ /*33269*/;
assign _38579_ = _38580_ | _38582_ /*33266*/;
assign _38588_ = ~D[11] /*33265*/;
assign _38585_ = _38027_ & _38588_ /*33261*/;
assign _38586_ = _38027_ ^ _38588_ /*33264*/;
assign _38587_ = _38579_ & _38586_ /*33262*/;
assign _38476_ = _38579_ ^ _38586_ /*33263*/;
assign _38584_ = _38585_ | _38587_ /*33260*/;
assign _38593_ = ~D[12] /*33259*/;
assign _38590_ = _38028_ & _38593_ /*33255*/;
assign _38591_ = _38028_ ^ _38593_ /*33258*/;
assign _38592_ = _38584_ & _38591_ /*33256*/;
assign _38477_ = _38584_ ^ _38591_ /*33257*/;
assign _38589_ = _38590_ | _38592_ /*33254*/;
assign _38598_ = ~D[13] /*33253*/;
assign _38595_ = _38029_ & _38598_ /*33249*/;
assign _38596_ = _38029_ ^ _38598_ /*33252*/;
assign _38597_ = _38589_ & _38596_ /*33250*/;
assign _38478_ = _38589_ ^ _38596_ /*33251*/;
assign _38594_ = _38595_ | _38597_ /*33248*/;
assign _38603_ = ~D[14] /*33247*/;
assign _38600_ = _38030_ & _38603_ /*33243*/;
assign _38601_ = _38030_ ^ _38603_ /*33246*/;
assign _38602_ = _38594_ & _38601_ /*33244*/;
assign _38479_ = _38594_ ^ _38601_ /*33245*/;
assign _38599_ = _38600_ | _38602_ /*33242*/;
assign _38608_ = ~D[15] /*33241*/;
assign _38605_ = _38031_ & _38608_ /*33237*/;
assign _38606_ = _38031_ ^ _38608_ /*33240*/;
assign _38607_ = _38599_ & _38606_ /*33238*/;
assign _38480_ = _38599_ ^ _38606_ /*33239*/;
assign _38604_ = _38605_ | _38607_ /*33236*/;
assign _38613_ = ~D[16] /*33235*/;
assign _38610_ = _38032_ & _38613_ /*33231*/;
assign _38611_ = _38032_ ^ _38613_ /*33234*/;
assign _38612_ = _38604_ & _38611_ /*33232*/;
assign _38481_ = _38604_ ^ _38611_ /*33233*/;
assign _38609_ = _38610_ | _38612_ /*33230*/;
assign _38618_ = ~D[17] /*33229*/;
assign _38615_ = _38033_ & _38618_ /*33225*/;
assign _38616_ = _38033_ ^ _38618_ /*33228*/;
assign _38617_ = _38609_ & _38616_ /*33226*/;
assign _38482_ = _38609_ ^ _38616_ /*33227*/;
assign _38614_ = _38615_ | _38617_ /*33224*/;
assign _38623_ = ~D[18] /*33223*/;
assign _38620_ = _38034_ & _38623_ /*33219*/;
assign _38621_ = _38034_ ^ _38623_ /*33222*/;
assign _38622_ = _38614_ & _38621_ /*33220*/;
assign _38483_ = _38614_ ^ _38621_ /*33221*/;
assign _38619_ = _38620_ | _38622_ /*33218*/;
assign _38628_ = ~D[19] /*33217*/;
assign _38625_ = _38035_ & _38628_ /*33213*/;
assign _38626_ = _38035_ ^ _38628_ /*33216*/;
assign _38627_ = _38619_ & _38626_ /*33214*/;
assign _38484_ = _38619_ ^ _38626_ /*33215*/;
assign _38624_ = _38625_ | _38627_ /*33212*/;
assign _38633_ = ~D[20] /*33211*/;
assign _38630_ = _38036_ & _38633_ /*33207*/;
assign _38631_ = _38036_ ^ _38633_ /*33210*/;
assign _38632_ = _38624_ & _38631_ /*33208*/;
assign _38485_ = _38624_ ^ _38631_ /*33209*/;
assign _38629_ = _38630_ | _38632_ /*33206*/;
assign _38638_ = ~D[21] /*33205*/;
assign _38635_ = _38037_ & _38638_ /*33201*/;
assign _38636_ = _38037_ ^ _38638_ /*33204*/;
assign _38637_ = _38629_ & _38636_ /*33202*/;
assign _38486_ = _38629_ ^ _38636_ /*33203*/;
assign _38634_ = _38635_ | _38637_ /*33200*/;
assign _38643_ = ~D[22] /*33199*/;
assign _38640_ = _38038_ & _38643_ /*33195*/;
assign _38641_ = _38038_ ^ _38643_ /*33198*/;
assign _38642_ = _38634_ & _38641_ /*33196*/;
assign _38487_ = _38634_ ^ _38641_ /*33197*/;
assign _38639_ = _38640_ | _38642_ /*33194*/;
assign _38648_ = ~D[23] /*33193*/;
assign _38645_ = _38039_ & _38648_ /*33189*/;
assign _38646_ = _38039_ ^ _38648_ /*33192*/;
assign _38647_ = _38639_ & _38646_ /*33190*/;
assign _38488_ = _38639_ ^ _38646_ /*33191*/;
assign _38644_ = _38645_ | _38647_ /*33188*/;
assign _38653_ = ~D[24] /*33187*/;
assign _38650_ = _38040_ & _38653_ /*33183*/;
assign _38651_ = _38040_ ^ _38653_ /*33186*/;
assign _38652_ = _38644_ & _38651_ /*33184*/;
assign _38489_ = _38644_ ^ _38651_ /*33185*/;
assign _38649_ = _38650_ | _38652_ /*33182*/;
assign _38658_ = ~D[25] /*33181*/;
assign _38655_ = _38041_ & _38658_ /*33177*/;
assign _38656_ = _38041_ ^ _38658_ /*33180*/;
assign _38657_ = _38649_ & _38656_ /*33178*/;
assign _38490_ = _38649_ ^ _38656_ /*33179*/;
assign _38654_ = _38655_ | _38657_ /*33176*/;
assign _38663_ = ~D[26] /*33175*/;
assign _38660_ = _38042_ & _38663_ /*33171*/;
assign _38661_ = _38042_ ^ _38663_ /*33174*/;
assign _38662_ = _38654_ & _38661_ /*33172*/;
assign _38491_ = _38654_ ^ _38661_ /*33173*/;
assign _38659_ = _38660_ | _38662_ /*33170*/;
assign _38668_ = ~D[27] /*33169*/;
assign _38665_ = _38043_ & _38668_ /*33165*/;
assign _38666_ = _38043_ ^ _38668_ /*33168*/;
assign _38667_ = _38659_ & _38666_ /*33166*/;
assign _38492_ = _38659_ ^ _38666_ /*33167*/;
assign _38664_ = _38665_ | _38667_ /*33164*/;
assign _38673_ = ~D[28] /*33163*/;
assign _38670_ = _38044_ & _38673_ /*33159*/;
assign _38671_ = _38044_ ^ _38673_ /*33162*/;
assign _38672_ = _38664_ & _38671_ /*33160*/;
assign _38493_ = _38664_ ^ _38671_ /*33161*/;
assign _38669_ = _38670_ | _38672_ /*33158*/;
assign _38678_ = ~D[29] /*33157*/;
assign _38675_ = _38045_ & _38678_ /*33153*/;
assign _38676_ = _38045_ ^ _38678_ /*33156*/;
assign _38677_ = _38669_ & _38676_ /*33154*/;
assign _38494_ = _38669_ ^ _38676_ /*33155*/;
assign _38674_ = _38675_ | _38677_ /*33152*/;
assign _38683_ = ~D[30] /*33151*/;
assign _38680_ = _38046_ & _38683_ /*33147*/;
assign _38681_ = _38046_ ^ _38683_ /*33150*/;
assign _38682_ = _38674_ & _38681_ /*33148*/;
assign _38495_ = _38674_ ^ _38681_ /*33149*/;
assign _38679_ = _38680_ | _38682_ /*33146*/;
assign _38688_ = ~D[31] /*33145*/;
assign _38685_ = _38047_ & _38688_ /*33141*/;
assign _38686_ = _38047_ ^ _38688_ /*33144*/;
assign _38687_ = _38679_ & _38686_ /*33142*/;
assign _38496_ = _38679_ ^ _38686_ /*33143*/;
assign _38684_ = _38685_ | _38687_ /*33140*/;
assign _38693_ = ~D[32] /*33139*/;
assign _38690_ = _38048_ & _38693_ /*33135*/;
assign _38691_ = _38048_ ^ _38693_ /*33138*/;
assign _38692_ = _38684_ & _38691_ /*33136*/;
assign _38497_ = _38684_ ^ _38691_ /*33137*/;
assign _38689_ = _38690_ | _38692_ /*33134*/;
assign _38698_ = ~D[33] /*33133*/;
assign _38695_ = _38049_ & _38698_ /*33129*/;
assign _38696_ = _38049_ ^ _38698_ /*33132*/;
assign _38697_ = _38689_ & _38696_ /*33130*/;
assign _38498_ = _38689_ ^ _38696_ /*33131*/;
assign _38694_ = _38695_ | _38697_ /*33128*/;
assign _38703_ = ~D[34] /*33127*/;
assign _38700_ = _38050_ & _38703_ /*33123*/;
assign _38701_ = _38050_ ^ _38703_ /*33126*/;
assign _38702_ = _38694_ & _38701_ /*33124*/;
assign _38499_ = _38694_ ^ _38701_ /*33125*/;
assign _38699_ = _38700_ | _38702_ /*33122*/;
assign _38708_ = ~D[35] /*33121*/;
assign _38705_ = _38051_ & _38708_ /*33117*/;
assign _38706_ = _38051_ ^ _38708_ /*33120*/;
assign _38707_ = _38699_ & _38706_ /*33118*/;
assign _38500_ = _38699_ ^ _38706_ /*33119*/;
assign _38704_ = _38705_ | _38707_ /*33116*/;
assign _38713_ = ~D[36] /*33115*/;
assign _38710_ = _38052_ & _38713_ /*33111*/;
assign _38711_ = _38052_ ^ _38713_ /*33114*/;
assign _38712_ = _38704_ & _38711_ /*33112*/;
assign _38501_ = _38704_ ^ _38711_ /*33113*/;
assign _38709_ = _38710_ | _38712_ /*33110*/;
assign _38718_ = ~D[37] /*33109*/;
assign _38715_ = _38053_ & _38718_ /*33105*/;
assign _38716_ = _38053_ ^ _38718_ /*33108*/;
assign _38717_ = _38709_ & _38716_ /*33106*/;
assign _38502_ = _38709_ ^ _38716_ /*33107*/;
assign _38714_ = _38715_ | _38717_ /*33104*/;
assign _38723_ = ~D[38] /*33103*/;
assign _38720_ = _38054_ & _38723_ /*33099*/;
assign _38721_ = _38054_ ^ _38723_ /*33102*/;
assign _38722_ = _38714_ & _38721_ /*33100*/;
assign _38503_ = _38714_ ^ _38721_ /*33101*/;
assign _38719_ = _38720_ | _38722_ /*33098*/;
assign _38728_ = ~D[39] /*33097*/;
assign _38725_ = _38055_ & _38728_ /*33093*/;
assign _38726_ = _38055_ ^ _38728_ /*33096*/;
assign _38727_ = _38719_ & _38726_ /*33094*/;
assign _38504_ = _38719_ ^ _38726_ /*33095*/;
assign _38724_ = _38725_ | _38727_ /*33092*/;
assign _38733_ = ~D[40] /*33091*/;
assign _38730_ = _38056_ & _38733_ /*33087*/;
assign _38731_ = _38056_ ^ _38733_ /*33090*/;
assign _38732_ = _38724_ & _38731_ /*33088*/;
assign _38505_ = _38724_ ^ _38731_ /*33089*/;
assign _38729_ = _38730_ | _38732_ /*33086*/;
assign _38738_ = ~D[41] /*33085*/;
assign _38735_ = _38057_ & _38738_ /*33081*/;
assign _38736_ = _38057_ ^ _38738_ /*33084*/;
assign _38737_ = _38729_ & _38736_ /*33082*/;
assign _38506_ = _38729_ ^ _38736_ /*33083*/;
assign _38734_ = _38735_ | _38737_ /*33080*/;
assign _38743_ = ~D[42] /*33079*/;
assign _38740_ = _38058_ & _38743_ /*33075*/;
assign _38741_ = _38058_ ^ _38743_ /*33078*/;
assign _38742_ = _38734_ & _38741_ /*33076*/;
assign _38507_ = _38734_ ^ _38741_ /*33077*/;
assign _38739_ = _38740_ | _38742_ /*33074*/;
assign _38748_ = ~D[43] /*33073*/;
assign _38745_ = _38059_ & _38748_ /*33069*/;
assign _38746_ = _38059_ ^ _38748_ /*33072*/;
assign _38747_ = _38739_ & _38746_ /*33070*/;
assign _38508_ = _38739_ ^ _38746_ /*33071*/;
assign _38744_ = _38745_ | _38747_ /*33068*/;
assign _38753_ = ~D[44] /*33067*/;
assign _38750_ = _38060_ & _38753_ /*33063*/;
assign _38751_ = _38060_ ^ _38753_ /*33066*/;
assign _38752_ = _38744_ & _38751_ /*33064*/;
assign _38509_ = _38744_ ^ _38751_ /*33065*/;
assign _38749_ = _38750_ | _38752_ /*33062*/;
assign _38758_ = ~D[45] /*33061*/;
assign _38755_ = _38061_ & _38758_ /*33057*/;
assign _38756_ = _38061_ ^ _38758_ /*33060*/;
assign _38757_ = _38749_ & _38756_ /*33058*/;
assign _38510_ = _38749_ ^ _38756_ /*33059*/;
assign _38754_ = _38755_ | _38757_ /*33056*/;
assign _38763_ = ~D[46] /*33055*/;
assign _38760_ = _38062_ & _38763_ /*33051*/;
assign _38761_ = _38062_ ^ _38763_ /*33054*/;
assign _38762_ = _38754_ & _38761_ /*33052*/;
assign _38511_ = _38754_ ^ _38761_ /*33053*/;
assign _38759_ = _38760_ | _38762_ /*33050*/;
assign _38768_ = ~D[47] /*33049*/;
assign _38765_ = _38063_ & _38768_ /*33045*/;
assign _38766_ = _38063_ ^ _38768_ /*33048*/;
assign _38767_ = _38759_ & _38766_ /*33046*/;
assign _38512_ = _38759_ ^ _38766_ /*33047*/;
assign _38764_ = _38765_ | _38767_ /*33044*/;
assign _38773_ = ~D[48] /*33043*/;
assign _38770_ = _38064_ & _38773_ /*33039*/;
assign _38771_ = _38064_ ^ _38773_ /*33042*/;
assign _38772_ = _38764_ & _38771_ /*33040*/;
assign _38513_ = _38764_ ^ _38771_ /*33041*/;
assign _38769_ = _38770_ | _38772_ /*33038*/;
assign _38778_ = ~D[49] /*33037*/;
assign _38775_ = _38065_ & _38778_ /*33033*/;
assign _38776_ = _38065_ ^ _38778_ /*33036*/;
assign _38777_ = _38769_ & _38776_ /*33034*/;
assign _38514_ = _38769_ ^ _38776_ /*33035*/;
assign _38774_ = _38775_ | _38777_ /*33032*/;
assign _38783_ = ~D[50] /*33031*/;
assign _38780_ = _38066_ & _38783_ /*33027*/;
assign _38781_ = _38066_ ^ _38783_ /*33030*/;
assign _38782_ = _38774_ & _38781_ /*33028*/;
assign _38515_ = _38774_ ^ _38781_ /*33029*/;
assign _38779_ = _38780_ | _38782_ /*33026*/;
assign _38788_ = ~D[51] /*33025*/;
assign _38785_ = _38067_ & _38788_ /*33021*/;
assign _38786_ = _38067_ ^ _38788_ /*33024*/;
assign _38787_ = _38779_ & _38786_ /*33022*/;
assign _38516_ = _38779_ ^ _38786_ /*33023*/;
assign _38784_ = _38785_ | _38787_ /*33020*/;
assign _38793_ = ~D[52] /*33019*/;
assign _38790_ = _38068_ & _38793_ /*33015*/;
assign _38791_ = _38068_ ^ _38793_ /*33018*/;
assign _38792_ = _38784_ & _38791_ /*33016*/;
assign _38517_ = _38784_ ^ _38791_ /*33017*/;
assign _38789_ = _38790_ | _38792_ /*33014*/;
assign _38798_ = ~D[53] /*33013*/;
assign _38795_ = _38069_ & _38798_ /*33009*/;
assign _38796_ = _38069_ ^ _38798_ /*33012*/;
assign _38797_ = _38789_ & _38796_ /*33010*/;
assign _38518_ = _38789_ ^ _38796_ /*33011*/;
assign _38794_ = _38795_ | _38797_ /*33008*/;
assign _38803_ = ~D[54] /*33007*/;
assign _38800_ = _38070_ & _38803_ /*33003*/;
assign _38801_ = _38070_ ^ _38803_ /*33006*/;
assign _38802_ = _38794_ & _38801_ /*33004*/;
assign _38519_ = _38794_ ^ _38801_ /*33005*/;
assign _38799_ = _38800_ | _38802_ /*33002*/;
assign _38808_ = ~D[55] /*33001*/;
assign _38805_ = _38071_ & _38808_ /*32997*/;
assign _38806_ = _38071_ ^ _38808_ /*33000*/;
assign _38807_ = _38799_ & _38806_ /*32998*/;
assign _38520_ = _38799_ ^ _38806_ /*32999*/;
assign _38804_ = _38805_ | _38807_ /*32996*/;
assign _38813_ = ~D[56] /*32995*/;
assign _38810_ = _38072_ & _38813_ /*32991*/;
assign _38811_ = _38072_ ^ _38813_ /*32994*/;
assign _38812_ = _38804_ & _38811_ /*32992*/;
assign _38521_ = _38804_ ^ _38811_ /*32993*/;
assign _38809_ = _38810_ | _38812_ /*32990*/;
assign _38818_ = ~D[57] /*32989*/;
assign _38815_ = _38073_ & _38818_ /*32985*/;
assign _38816_ = _38073_ ^ _38818_ /*32988*/;
assign _38817_ = _38809_ & _38816_ /*32986*/;
assign _38522_ = _38809_ ^ _38816_ /*32987*/;
assign _38814_ = _38815_ | _38817_ /*32984*/;
assign _38823_ = ~D[58] /*32983*/;
assign _38820_ = _38074_ & _38823_ /*32979*/;
assign _38821_ = _38074_ ^ _38823_ /*32982*/;
assign _38822_ = _38814_ & _38821_ /*32980*/;
assign _38523_ = _38814_ ^ _38821_ /*32981*/;
assign _38819_ = _38820_ | _38822_ /*32978*/;
assign _38828_ = ~D[59] /*32977*/;
assign _38825_ = _38075_ & _38828_ /*32973*/;
assign _38826_ = _38075_ ^ _38828_ /*32976*/;
assign _38827_ = _38819_ & _38826_ /*32974*/;
assign _38524_ = _38819_ ^ _38826_ /*32975*/;
assign _38824_ = _38825_ | _38827_ /*32972*/;
assign _38833_ = ~D[60] /*32971*/;
assign _38830_ = _38076_ & _38833_ /*32967*/;
assign _38831_ = _38076_ ^ _38833_ /*32970*/;
assign _38832_ = _38824_ & _38831_ /*32968*/;
assign _38525_ = _38824_ ^ _38831_ /*32969*/;
assign _38829_ = _38830_ | _38832_ /*32966*/;
assign _38838_ = ~D[61] /*32965*/;
assign _38835_ = _38077_ & _38838_ /*32961*/;
assign _38836_ = _38077_ ^ _38838_ /*32964*/;
assign _38837_ = _38829_ & _38836_ /*32962*/;
assign _38526_ = _38829_ ^ _38836_ /*32963*/;
assign _38834_ = _38835_ | _38837_ /*32960*/;
assign _38843_ = ~D[62] /*32959*/;
assign _38840_ = _38078_ & _38843_ /*32955*/;
assign _38841_ = _38078_ ^ _38843_ /*32958*/;
assign _38842_ = _38834_ & _38841_ /*32956*/;
assign _38527_ = _38834_ ^ _38841_ /*32957*/;
assign _38839_ = _38840_ | _38842_ /*32954*/;
assign _38844_ = _38079_ & oneWire /*32949*/;
assign _38845_ = _38079_ ^ oneWire /*32952*/;
assign _38846_ = _38839_ & _38845_ /*32950*/;
assign _38528_ = _38839_ ^ _38845_ /*32951*/;
assign Q[20] = _38844_ | _38846_ /*32948*/;
assign _38979_ = ~Q[20] /*32563*/;
assign _38978_ = _38979_ & D[0] /*32562*/;
assign _38981_ = _38465_ & _38978_ /*32557*/;
assign _38982_ = _38465_ ^ _38978_ /*32560*/;
assign _38983_ = zeroWire & _38982_ /*32558*/;
assign _38913_ = zeroWire ^ _38982_ /*32559*/;
assign _38980_ = _38981_ | _38983_ /*32556*/;
assign _38985_ = ~Q[20] /*32555*/;
assign _38984_ = _38985_ & D[1] /*32554*/;
assign _38987_ = _38466_ & _38984_ /*32549*/;
assign _38988_ = _38466_ ^ _38984_ /*32552*/;
assign _38989_ = _38980_ & _38988_ /*32550*/;
assign _38914_ = _38980_ ^ _38988_ /*32551*/;
assign _38986_ = _38987_ | _38989_ /*32548*/;
assign _38991_ = ~Q[20] /*32547*/;
assign _38990_ = _38991_ & D[2] /*32546*/;
assign _38993_ = _38467_ & _38990_ /*32541*/;
assign _38994_ = _38467_ ^ _38990_ /*32544*/;
assign _38995_ = _38986_ & _38994_ /*32542*/;
assign _38915_ = _38986_ ^ _38994_ /*32543*/;
assign _38992_ = _38993_ | _38995_ /*32540*/;
assign _38997_ = ~Q[20] /*32539*/;
assign _38996_ = _38997_ & D[3] /*32538*/;
assign _38999_ = _38468_ & _38996_ /*32533*/;
assign _39000_ = _38468_ ^ _38996_ /*32536*/;
assign _39001_ = _38992_ & _39000_ /*32534*/;
assign _38916_ = _38992_ ^ _39000_ /*32535*/;
assign _38998_ = _38999_ | _39001_ /*32532*/;
assign _39003_ = ~Q[20] /*32531*/;
assign _39002_ = _39003_ & D[4] /*32530*/;
assign _39005_ = _38469_ & _39002_ /*32525*/;
assign _39006_ = _38469_ ^ _39002_ /*32528*/;
assign _39007_ = _38998_ & _39006_ /*32526*/;
assign _38917_ = _38998_ ^ _39006_ /*32527*/;
assign _39004_ = _39005_ | _39007_ /*32524*/;
assign _39009_ = ~Q[20] /*32523*/;
assign _39008_ = _39009_ & D[5] /*32522*/;
assign _39011_ = _38470_ & _39008_ /*32517*/;
assign _39012_ = _38470_ ^ _39008_ /*32520*/;
assign _39013_ = _39004_ & _39012_ /*32518*/;
assign _38918_ = _39004_ ^ _39012_ /*32519*/;
assign _39010_ = _39011_ | _39013_ /*32516*/;
assign _39015_ = ~Q[20] /*32515*/;
assign _39014_ = _39015_ & D[6] /*32514*/;
assign _39017_ = _38471_ & _39014_ /*32509*/;
assign _39018_ = _38471_ ^ _39014_ /*32512*/;
assign _39019_ = _39010_ & _39018_ /*32510*/;
assign _38919_ = _39010_ ^ _39018_ /*32511*/;
assign _39016_ = _39017_ | _39019_ /*32508*/;
assign _39021_ = ~Q[20] /*32507*/;
assign _39020_ = _39021_ & D[7] /*32506*/;
assign _39023_ = _38472_ & _39020_ /*32501*/;
assign _39024_ = _38472_ ^ _39020_ /*32504*/;
assign _39025_ = _39016_ & _39024_ /*32502*/;
assign _38920_ = _39016_ ^ _39024_ /*32503*/;
assign _39022_ = _39023_ | _39025_ /*32500*/;
assign _39027_ = ~Q[20] /*32499*/;
assign _39026_ = _39027_ & D[8] /*32498*/;
assign _39029_ = _38473_ & _39026_ /*32493*/;
assign _39030_ = _38473_ ^ _39026_ /*32496*/;
assign _39031_ = _39022_ & _39030_ /*32494*/;
assign _38921_ = _39022_ ^ _39030_ /*32495*/;
assign _39028_ = _39029_ | _39031_ /*32492*/;
assign _39033_ = ~Q[20] /*32491*/;
assign _39032_ = _39033_ & D[9] /*32490*/;
assign _39035_ = _38474_ & _39032_ /*32485*/;
assign _39036_ = _38474_ ^ _39032_ /*32488*/;
assign _39037_ = _39028_ & _39036_ /*32486*/;
assign _38922_ = _39028_ ^ _39036_ /*32487*/;
assign _39034_ = _39035_ | _39037_ /*32484*/;
assign _39039_ = ~Q[20] /*32483*/;
assign _39038_ = _39039_ & D[10] /*32482*/;
assign _39041_ = _38475_ & _39038_ /*32477*/;
assign _39042_ = _38475_ ^ _39038_ /*32480*/;
assign _39043_ = _39034_ & _39042_ /*32478*/;
assign _38923_ = _39034_ ^ _39042_ /*32479*/;
assign _39040_ = _39041_ | _39043_ /*32476*/;
assign _39045_ = ~Q[20] /*32475*/;
assign _39044_ = _39045_ & D[11] /*32474*/;
assign _39047_ = _38476_ & _39044_ /*32469*/;
assign _39048_ = _38476_ ^ _39044_ /*32472*/;
assign _39049_ = _39040_ & _39048_ /*32470*/;
assign _38924_ = _39040_ ^ _39048_ /*32471*/;
assign _39046_ = _39047_ | _39049_ /*32468*/;
assign _39051_ = ~Q[20] /*32467*/;
assign _39050_ = _39051_ & D[12] /*32466*/;
assign _39053_ = _38477_ & _39050_ /*32461*/;
assign _39054_ = _38477_ ^ _39050_ /*32464*/;
assign _39055_ = _39046_ & _39054_ /*32462*/;
assign _38925_ = _39046_ ^ _39054_ /*32463*/;
assign _39052_ = _39053_ | _39055_ /*32460*/;
assign _39057_ = ~Q[20] /*32459*/;
assign _39056_ = _39057_ & D[13] /*32458*/;
assign _39059_ = _38478_ & _39056_ /*32453*/;
assign _39060_ = _38478_ ^ _39056_ /*32456*/;
assign _39061_ = _39052_ & _39060_ /*32454*/;
assign _38926_ = _39052_ ^ _39060_ /*32455*/;
assign _39058_ = _39059_ | _39061_ /*32452*/;
assign _39063_ = ~Q[20] /*32451*/;
assign _39062_ = _39063_ & D[14] /*32450*/;
assign _39065_ = _38479_ & _39062_ /*32445*/;
assign _39066_ = _38479_ ^ _39062_ /*32448*/;
assign _39067_ = _39058_ & _39066_ /*32446*/;
assign _38927_ = _39058_ ^ _39066_ /*32447*/;
assign _39064_ = _39065_ | _39067_ /*32444*/;
assign _39069_ = ~Q[20] /*32443*/;
assign _39068_ = _39069_ & D[15] /*32442*/;
assign _39071_ = _38480_ & _39068_ /*32437*/;
assign _39072_ = _38480_ ^ _39068_ /*32440*/;
assign _39073_ = _39064_ & _39072_ /*32438*/;
assign _38928_ = _39064_ ^ _39072_ /*32439*/;
assign _39070_ = _39071_ | _39073_ /*32436*/;
assign _39075_ = ~Q[20] /*32435*/;
assign _39074_ = _39075_ & D[16] /*32434*/;
assign _39077_ = _38481_ & _39074_ /*32429*/;
assign _39078_ = _38481_ ^ _39074_ /*32432*/;
assign _39079_ = _39070_ & _39078_ /*32430*/;
assign _38929_ = _39070_ ^ _39078_ /*32431*/;
assign _39076_ = _39077_ | _39079_ /*32428*/;
assign _39081_ = ~Q[20] /*32427*/;
assign _39080_ = _39081_ & D[17] /*32426*/;
assign _39083_ = _38482_ & _39080_ /*32421*/;
assign _39084_ = _38482_ ^ _39080_ /*32424*/;
assign _39085_ = _39076_ & _39084_ /*32422*/;
assign _38930_ = _39076_ ^ _39084_ /*32423*/;
assign _39082_ = _39083_ | _39085_ /*32420*/;
assign _39087_ = ~Q[20] /*32419*/;
assign _39086_ = _39087_ & D[18] /*32418*/;
assign _39089_ = _38483_ & _39086_ /*32413*/;
assign _39090_ = _38483_ ^ _39086_ /*32416*/;
assign _39091_ = _39082_ & _39090_ /*32414*/;
assign _38931_ = _39082_ ^ _39090_ /*32415*/;
assign _39088_ = _39089_ | _39091_ /*32412*/;
assign _39093_ = ~Q[20] /*32411*/;
assign _39092_ = _39093_ & D[19] /*32410*/;
assign _39095_ = _38484_ & _39092_ /*32405*/;
assign _39096_ = _38484_ ^ _39092_ /*32408*/;
assign _39097_ = _39088_ & _39096_ /*32406*/;
assign _38932_ = _39088_ ^ _39096_ /*32407*/;
assign _39094_ = _39095_ | _39097_ /*32404*/;
assign _39099_ = ~Q[20] /*32403*/;
assign _39098_ = _39099_ & D[20] /*32402*/;
assign _39101_ = _38485_ & _39098_ /*32397*/;
assign _39102_ = _38485_ ^ _39098_ /*32400*/;
assign _39103_ = _39094_ & _39102_ /*32398*/;
assign _38933_ = _39094_ ^ _39102_ /*32399*/;
assign _39100_ = _39101_ | _39103_ /*32396*/;
assign _39105_ = ~Q[20] /*32395*/;
assign _39104_ = _39105_ & D[21] /*32394*/;
assign _39107_ = _38486_ & _39104_ /*32389*/;
assign _39108_ = _38486_ ^ _39104_ /*32392*/;
assign _39109_ = _39100_ & _39108_ /*32390*/;
assign _38934_ = _39100_ ^ _39108_ /*32391*/;
assign _39106_ = _39107_ | _39109_ /*32388*/;
assign _39111_ = ~Q[20] /*32387*/;
assign _39110_ = _39111_ & D[22] /*32386*/;
assign _39113_ = _38487_ & _39110_ /*32381*/;
assign _39114_ = _38487_ ^ _39110_ /*32384*/;
assign _39115_ = _39106_ & _39114_ /*32382*/;
assign _38935_ = _39106_ ^ _39114_ /*32383*/;
assign _39112_ = _39113_ | _39115_ /*32380*/;
assign _39117_ = ~Q[20] /*32379*/;
assign _39116_ = _39117_ & D[23] /*32378*/;
assign _39119_ = _38488_ & _39116_ /*32373*/;
assign _39120_ = _38488_ ^ _39116_ /*32376*/;
assign _39121_ = _39112_ & _39120_ /*32374*/;
assign _38936_ = _39112_ ^ _39120_ /*32375*/;
assign _39118_ = _39119_ | _39121_ /*32372*/;
assign _39123_ = ~Q[20] /*32371*/;
assign _39122_ = _39123_ & D[24] /*32370*/;
assign _39125_ = _38489_ & _39122_ /*32365*/;
assign _39126_ = _38489_ ^ _39122_ /*32368*/;
assign _39127_ = _39118_ & _39126_ /*32366*/;
assign _38937_ = _39118_ ^ _39126_ /*32367*/;
assign _39124_ = _39125_ | _39127_ /*32364*/;
assign _39129_ = ~Q[20] /*32363*/;
assign _39128_ = _39129_ & D[25] /*32362*/;
assign _39131_ = _38490_ & _39128_ /*32357*/;
assign _39132_ = _38490_ ^ _39128_ /*32360*/;
assign _39133_ = _39124_ & _39132_ /*32358*/;
assign _38938_ = _39124_ ^ _39132_ /*32359*/;
assign _39130_ = _39131_ | _39133_ /*32356*/;
assign _39135_ = ~Q[20] /*32355*/;
assign _39134_ = _39135_ & D[26] /*32354*/;
assign _39137_ = _38491_ & _39134_ /*32349*/;
assign _39138_ = _38491_ ^ _39134_ /*32352*/;
assign _39139_ = _39130_ & _39138_ /*32350*/;
assign _38939_ = _39130_ ^ _39138_ /*32351*/;
assign _39136_ = _39137_ | _39139_ /*32348*/;
assign _39141_ = ~Q[20] /*32347*/;
assign _39140_ = _39141_ & D[27] /*32346*/;
assign _39143_ = _38492_ & _39140_ /*32341*/;
assign _39144_ = _38492_ ^ _39140_ /*32344*/;
assign _39145_ = _39136_ & _39144_ /*32342*/;
assign _38940_ = _39136_ ^ _39144_ /*32343*/;
assign _39142_ = _39143_ | _39145_ /*32340*/;
assign _39147_ = ~Q[20] /*32339*/;
assign _39146_ = _39147_ & D[28] /*32338*/;
assign _39149_ = _38493_ & _39146_ /*32333*/;
assign _39150_ = _38493_ ^ _39146_ /*32336*/;
assign _39151_ = _39142_ & _39150_ /*32334*/;
assign _38941_ = _39142_ ^ _39150_ /*32335*/;
assign _39148_ = _39149_ | _39151_ /*32332*/;
assign _39153_ = ~Q[20] /*32331*/;
assign _39152_ = _39153_ & D[29] /*32330*/;
assign _39155_ = _38494_ & _39152_ /*32325*/;
assign _39156_ = _38494_ ^ _39152_ /*32328*/;
assign _39157_ = _39148_ & _39156_ /*32326*/;
assign _38942_ = _39148_ ^ _39156_ /*32327*/;
assign _39154_ = _39155_ | _39157_ /*32324*/;
assign _39159_ = ~Q[20] /*32323*/;
assign _39158_ = _39159_ & D[30] /*32322*/;
assign _39161_ = _38495_ & _39158_ /*32317*/;
assign _39162_ = _38495_ ^ _39158_ /*32320*/;
assign _39163_ = _39154_ & _39162_ /*32318*/;
assign _38943_ = _39154_ ^ _39162_ /*32319*/;
assign _39160_ = _39161_ | _39163_ /*32316*/;
assign _39165_ = ~Q[20] /*32315*/;
assign _39164_ = _39165_ & D[31] /*32314*/;
assign _39167_ = _38496_ & _39164_ /*32309*/;
assign _39168_ = _38496_ ^ _39164_ /*32312*/;
assign _39169_ = _39160_ & _39168_ /*32310*/;
assign _38944_ = _39160_ ^ _39168_ /*32311*/;
assign _39166_ = _39167_ | _39169_ /*32308*/;
assign _39171_ = ~Q[20] /*32307*/;
assign _39170_ = _39171_ & D[32] /*32306*/;
assign _39173_ = _38497_ & _39170_ /*32301*/;
assign _39174_ = _38497_ ^ _39170_ /*32304*/;
assign _39175_ = _39166_ & _39174_ /*32302*/;
assign _38945_ = _39166_ ^ _39174_ /*32303*/;
assign _39172_ = _39173_ | _39175_ /*32300*/;
assign _39177_ = ~Q[20] /*32299*/;
assign _39176_ = _39177_ & D[33] /*32298*/;
assign _39179_ = _38498_ & _39176_ /*32293*/;
assign _39180_ = _38498_ ^ _39176_ /*32296*/;
assign _39181_ = _39172_ & _39180_ /*32294*/;
assign _38946_ = _39172_ ^ _39180_ /*32295*/;
assign _39178_ = _39179_ | _39181_ /*32292*/;
assign _39183_ = ~Q[20] /*32291*/;
assign _39182_ = _39183_ & D[34] /*32290*/;
assign _39185_ = _38499_ & _39182_ /*32285*/;
assign _39186_ = _38499_ ^ _39182_ /*32288*/;
assign _39187_ = _39178_ & _39186_ /*32286*/;
assign _38947_ = _39178_ ^ _39186_ /*32287*/;
assign _39184_ = _39185_ | _39187_ /*32284*/;
assign _39189_ = ~Q[20] /*32283*/;
assign _39188_ = _39189_ & D[35] /*32282*/;
assign _39191_ = _38500_ & _39188_ /*32277*/;
assign _39192_ = _38500_ ^ _39188_ /*32280*/;
assign _39193_ = _39184_ & _39192_ /*32278*/;
assign _38948_ = _39184_ ^ _39192_ /*32279*/;
assign _39190_ = _39191_ | _39193_ /*32276*/;
assign _39195_ = ~Q[20] /*32275*/;
assign _39194_ = _39195_ & D[36] /*32274*/;
assign _39197_ = _38501_ & _39194_ /*32269*/;
assign _39198_ = _38501_ ^ _39194_ /*32272*/;
assign _39199_ = _39190_ & _39198_ /*32270*/;
assign _38949_ = _39190_ ^ _39198_ /*32271*/;
assign _39196_ = _39197_ | _39199_ /*32268*/;
assign _39201_ = ~Q[20] /*32267*/;
assign _39200_ = _39201_ & D[37] /*32266*/;
assign _39203_ = _38502_ & _39200_ /*32261*/;
assign _39204_ = _38502_ ^ _39200_ /*32264*/;
assign _39205_ = _39196_ & _39204_ /*32262*/;
assign _38950_ = _39196_ ^ _39204_ /*32263*/;
assign _39202_ = _39203_ | _39205_ /*32260*/;
assign _39207_ = ~Q[20] /*32259*/;
assign _39206_ = _39207_ & D[38] /*32258*/;
assign _39209_ = _38503_ & _39206_ /*32253*/;
assign _39210_ = _38503_ ^ _39206_ /*32256*/;
assign _39211_ = _39202_ & _39210_ /*32254*/;
assign _38951_ = _39202_ ^ _39210_ /*32255*/;
assign _39208_ = _39209_ | _39211_ /*32252*/;
assign _39213_ = ~Q[20] /*32251*/;
assign _39212_ = _39213_ & D[39] /*32250*/;
assign _39215_ = _38504_ & _39212_ /*32245*/;
assign _39216_ = _38504_ ^ _39212_ /*32248*/;
assign _39217_ = _39208_ & _39216_ /*32246*/;
assign _38952_ = _39208_ ^ _39216_ /*32247*/;
assign _39214_ = _39215_ | _39217_ /*32244*/;
assign _39219_ = ~Q[20] /*32243*/;
assign _39218_ = _39219_ & D[40] /*32242*/;
assign _39221_ = _38505_ & _39218_ /*32237*/;
assign _39222_ = _38505_ ^ _39218_ /*32240*/;
assign _39223_ = _39214_ & _39222_ /*32238*/;
assign _38953_ = _39214_ ^ _39222_ /*32239*/;
assign _39220_ = _39221_ | _39223_ /*32236*/;
assign _39225_ = ~Q[20] /*32235*/;
assign _39224_ = _39225_ & D[41] /*32234*/;
assign _39227_ = _38506_ & _39224_ /*32229*/;
assign _39228_ = _38506_ ^ _39224_ /*32232*/;
assign _39229_ = _39220_ & _39228_ /*32230*/;
assign _38954_ = _39220_ ^ _39228_ /*32231*/;
assign _39226_ = _39227_ | _39229_ /*32228*/;
assign _39231_ = ~Q[20] /*32227*/;
assign _39230_ = _39231_ & D[42] /*32226*/;
assign _39233_ = _38507_ & _39230_ /*32221*/;
assign _39234_ = _38507_ ^ _39230_ /*32224*/;
assign _39235_ = _39226_ & _39234_ /*32222*/;
assign _38955_ = _39226_ ^ _39234_ /*32223*/;
assign _39232_ = _39233_ | _39235_ /*32220*/;
assign _39237_ = ~Q[20] /*32219*/;
assign _39236_ = _39237_ & D[43] /*32218*/;
assign _39239_ = _38508_ & _39236_ /*32213*/;
assign _39240_ = _38508_ ^ _39236_ /*32216*/;
assign _39241_ = _39232_ & _39240_ /*32214*/;
assign _38956_ = _39232_ ^ _39240_ /*32215*/;
assign _39238_ = _39239_ | _39241_ /*32212*/;
assign _39243_ = ~Q[20] /*32211*/;
assign _39242_ = _39243_ & D[44] /*32210*/;
assign _39245_ = _38509_ & _39242_ /*32205*/;
assign _39246_ = _38509_ ^ _39242_ /*32208*/;
assign _39247_ = _39238_ & _39246_ /*32206*/;
assign _38957_ = _39238_ ^ _39246_ /*32207*/;
assign _39244_ = _39245_ | _39247_ /*32204*/;
assign _39249_ = ~Q[20] /*32203*/;
assign _39248_ = _39249_ & D[45] /*32202*/;
assign _39251_ = _38510_ & _39248_ /*32197*/;
assign _39252_ = _38510_ ^ _39248_ /*32200*/;
assign _39253_ = _39244_ & _39252_ /*32198*/;
assign _38958_ = _39244_ ^ _39252_ /*32199*/;
assign _39250_ = _39251_ | _39253_ /*32196*/;
assign _39255_ = ~Q[20] /*32195*/;
assign _39254_ = _39255_ & D[46] /*32194*/;
assign _39257_ = _38511_ & _39254_ /*32189*/;
assign _39258_ = _38511_ ^ _39254_ /*32192*/;
assign _39259_ = _39250_ & _39258_ /*32190*/;
assign _38959_ = _39250_ ^ _39258_ /*32191*/;
assign _39256_ = _39257_ | _39259_ /*32188*/;
assign _39261_ = ~Q[20] /*32187*/;
assign _39260_ = _39261_ & D[47] /*32186*/;
assign _39263_ = _38512_ & _39260_ /*32181*/;
assign _39264_ = _38512_ ^ _39260_ /*32184*/;
assign _39265_ = _39256_ & _39264_ /*32182*/;
assign _38960_ = _39256_ ^ _39264_ /*32183*/;
assign _39262_ = _39263_ | _39265_ /*32180*/;
assign _39267_ = ~Q[20] /*32179*/;
assign _39266_ = _39267_ & D[48] /*32178*/;
assign _39269_ = _38513_ & _39266_ /*32173*/;
assign _39270_ = _38513_ ^ _39266_ /*32176*/;
assign _39271_ = _39262_ & _39270_ /*32174*/;
assign _38961_ = _39262_ ^ _39270_ /*32175*/;
assign _39268_ = _39269_ | _39271_ /*32172*/;
assign _39273_ = ~Q[20] /*32171*/;
assign _39272_ = _39273_ & D[49] /*32170*/;
assign _39275_ = _38514_ & _39272_ /*32165*/;
assign _39276_ = _38514_ ^ _39272_ /*32168*/;
assign _39277_ = _39268_ & _39276_ /*32166*/;
assign _38962_ = _39268_ ^ _39276_ /*32167*/;
assign _39274_ = _39275_ | _39277_ /*32164*/;
assign _39279_ = ~Q[20] /*32163*/;
assign _39278_ = _39279_ & D[50] /*32162*/;
assign _39281_ = _38515_ & _39278_ /*32157*/;
assign _39282_ = _38515_ ^ _39278_ /*32160*/;
assign _39283_ = _39274_ & _39282_ /*32158*/;
assign _38963_ = _39274_ ^ _39282_ /*32159*/;
assign _39280_ = _39281_ | _39283_ /*32156*/;
assign _39285_ = ~Q[20] /*32155*/;
assign _39284_ = _39285_ & D[51] /*32154*/;
assign _39287_ = _38516_ & _39284_ /*32149*/;
assign _39288_ = _38516_ ^ _39284_ /*32152*/;
assign _39289_ = _39280_ & _39288_ /*32150*/;
assign _38964_ = _39280_ ^ _39288_ /*32151*/;
assign _39286_ = _39287_ | _39289_ /*32148*/;
assign _39291_ = ~Q[20] /*32147*/;
assign _39290_ = _39291_ & D[52] /*32146*/;
assign _39293_ = _38517_ & _39290_ /*32141*/;
assign _39294_ = _38517_ ^ _39290_ /*32144*/;
assign _39295_ = _39286_ & _39294_ /*32142*/;
assign _38965_ = _39286_ ^ _39294_ /*32143*/;
assign _39292_ = _39293_ | _39295_ /*32140*/;
assign _39297_ = ~Q[20] /*32139*/;
assign _39296_ = _39297_ & D[53] /*32138*/;
assign _39299_ = _38518_ & _39296_ /*32133*/;
assign _39300_ = _38518_ ^ _39296_ /*32136*/;
assign _39301_ = _39292_ & _39300_ /*32134*/;
assign _38966_ = _39292_ ^ _39300_ /*32135*/;
assign _39298_ = _39299_ | _39301_ /*32132*/;
assign _39303_ = ~Q[20] /*32131*/;
assign _39302_ = _39303_ & D[54] /*32130*/;
assign _39305_ = _38519_ & _39302_ /*32125*/;
assign _39306_ = _38519_ ^ _39302_ /*32128*/;
assign _39307_ = _39298_ & _39306_ /*32126*/;
assign _38967_ = _39298_ ^ _39306_ /*32127*/;
assign _39304_ = _39305_ | _39307_ /*32124*/;
assign _39309_ = ~Q[20] /*32123*/;
assign _39308_ = _39309_ & D[55] /*32122*/;
assign _39311_ = _38520_ & _39308_ /*32117*/;
assign _39312_ = _38520_ ^ _39308_ /*32120*/;
assign _39313_ = _39304_ & _39312_ /*32118*/;
assign _38968_ = _39304_ ^ _39312_ /*32119*/;
assign _39310_ = _39311_ | _39313_ /*32116*/;
assign _39315_ = ~Q[20] /*32115*/;
assign _39314_ = _39315_ & D[56] /*32114*/;
assign _39317_ = _38521_ & _39314_ /*32109*/;
assign _39318_ = _38521_ ^ _39314_ /*32112*/;
assign _39319_ = _39310_ & _39318_ /*32110*/;
assign _38969_ = _39310_ ^ _39318_ /*32111*/;
assign _39316_ = _39317_ | _39319_ /*32108*/;
assign _39321_ = ~Q[20] /*32107*/;
assign _39320_ = _39321_ & D[57] /*32106*/;
assign _39323_ = _38522_ & _39320_ /*32101*/;
assign _39324_ = _38522_ ^ _39320_ /*32104*/;
assign _39325_ = _39316_ & _39324_ /*32102*/;
assign _38970_ = _39316_ ^ _39324_ /*32103*/;
assign _39322_ = _39323_ | _39325_ /*32100*/;
assign _39327_ = ~Q[20] /*32099*/;
assign _39326_ = _39327_ & D[58] /*32098*/;
assign _39329_ = _38523_ & _39326_ /*32093*/;
assign _39330_ = _38523_ ^ _39326_ /*32096*/;
assign _39331_ = _39322_ & _39330_ /*32094*/;
assign _38971_ = _39322_ ^ _39330_ /*32095*/;
assign _39328_ = _39329_ | _39331_ /*32092*/;
assign _39333_ = ~Q[20] /*32091*/;
assign _39332_ = _39333_ & D[59] /*32090*/;
assign _39335_ = _38524_ & _39332_ /*32085*/;
assign _39336_ = _38524_ ^ _39332_ /*32088*/;
assign _39337_ = _39328_ & _39336_ /*32086*/;
assign _38972_ = _39328_ ^ _39336_ /*32087*/;
assign _39334_ = _39335_ | _39337_ /*32084*/;
assign _39339_ = ~Q[20] /*32083*/;
assign _39338_ = _39339_ & D[60] /*32082*/;
assign _39341_ = _38525_ & _39338_ /*32077*/;
assign _39342_ = _38525_ ^ _39338_ /*32080*/;
assign _39343_ = _39334_ & _39342_ /*32078*/;
assign _38973_ = _39334_ ^ _39342_ /*32079*/;
assign _39340_ = _39341_ | _39343_ /*32076*/;
assign _39345_ = ~Q[20] /*32075*/;
assign _39344_ = _39345_ & D[61] /*32074*/;
assign _39347_ = _38526_ & _39344_ /*32069*/;
assign _39348_ = _38526_ ^ _39344_ /*32072*/;
assign _39349_ = _39340_ & _39348_ /*32070*/;
assign _38974_ = _39340_ ^ _39348_ /*32071*/;
assign _39346_ = _39347_ | _39349_ /*32068*/;
assign _39351_ = ~Q[20] /*32067*/;
assign _39350_ = _39351_ & D[62] /*32066*/;
assign _39353_ = _38527_ & _39350_ /*32061*/;
assign _39354_ = _38527_ ^ _39350_ /*32064*/;
assign _39355_ = _39346_ & _39354_ /*32062*/;
assign _38975_ = _39346_ ^ _39354_ /*32063*/;
assign _39352_ = _39353_ | _39355_ /*32060*/;
assign _39357_ = ~Q[20] /*32059*/;
assign _39356_ = _39357_ & zeroWire /*32058*/;
assign _39358_ = _38528_ ^ _39356_ /*32056*/;
assign _38976_ = _39358_ ^ _39352_ /*32055*/;
assign _39429_ = ~D[0] /*31801*/;
assign _39426_ = R_0[19] & _39429_ /*31797*/;
assign _39427_ = R_0[19] ^ _39429_ /*31800*/;
assign _39428_ = oneWire & _39427_ /*31798*/;
assign _39361_ = oneWire ^ _39427_ /*31799*/;
assign _39425_ = _39426_ | _39428_ /*31796*/;
assign _39434_ = ~D[1] /*31795*/;
assign _39431_ = _38913_ & _39434_ /*31791*/;
assign _39432_ = _38913_ ^ _39434_ /*31794*/;
assign _39433_ = _39425_ & _39432_ /*31792*/;
assign _39362_ = _39425_ ^ _39432_ /*31793*/;
assign _39430_ = _39431_ | _39433_ /*31790*/;
assign _39439_ = ~D[2] /*31789*/;
assign _39436_ = _38914_ & _39439_ /*31785*/;
assign _39437_ = _38914_ ^ _39439_ /*31788*/;
assign _39438_ = _39430_ & _39437_ /*31786*/;
assign _39363_ = _39430_ ^ _39437_ /*31787*/;
assign _39435_ = _39436_ | _39438_ /*31784*/;
assign _39444_ = ~D[3] /*31783*/;
assign _39441_ = _38915_ & _39444_ /*31779*/;
assign _39442_ = _38915_ ^ _39444_ /*31782*/;
assign _39443_ = _39435_ & _39442_ /*31780*/;
assign _39364_ = _39435_ ^ _39442_ /*31781*/;
assign _39440_ = _39441_ | _39443_ /*31778*/;
assign _39449_ = ~D[4] /*31777*/;
assign _39446_ = _38916_ & _39449_ /*31773*/;
assign _39447_ = _38916_ ^ _39449_ /*31776*/;
assign _39448_ = _39440_ & _39447_ /*31774*/;
assign _39365_ = _39440_ ^ _39447_ /*31775*/;
assign _39445_ = _39446_ | _39448_ /*31772*/;
assign _39454_ = ~D[5] /*31771*/;
assign _39451_ = _38917_ & _39454_ /*31767*/;
assign _39452_ = _38917_ ^ _39454_ /*31770*/;
assign _39453_ = _39445_ & _39452_ /*31768*/;
assign _39366_ = _39445_ ^ _39452_ /*31769*/;
assign _39450_ = _39451_ | _39453_ /*31766*/;
assign _39459_ = ~D[6] /*31765*/;
assign _39456_ = _38918_ & _39459_ /*31761*/;
assign _39457_ = _38918_ ^ _39459_ /*31764*/;
assign _39458_ = _39450_ & _39457_ /*31762*/;
assign _39367_ = _39450_ ^ _39457_ /*31763*/;
assign _39455_ = _39456_ | _39458_ /*31760*/;
assign _39464_ = ~D[7] /*31759*/;
assign _39461_ = _38919_ & _39464_ /*31755*/;
assign _39462_ = _38919_ ^ _39464_ /*31758*/;
assign _39463_ = _39455_ & _39462_ /*31756*/;
assign _39368_ = _39455_ ^ _39462_ /*31757*/;
assign _39460_ = _39461_ | _39463_ /*31754*/;
assign _39469_ = ~D[8] /*31753*/;
assign _39466_ = _38920_ & _39469_ /*31749*/;
assign _39467_ = _38920_ ^ _39469_ /*31752*/;
assign _39468_ = _39460_ & _39467_ /*31750*/;
assign _39369_ = _39460_ ^ _39467_ /*31751*/;
assign _39465_ = _39466_ | _39468_ /*31748*/;
assign _39474_ = ~D[9] /*31747*/;
assign _39471_ = _38921_ & _39474_ /*31743*/;
assign _39472_ = _38921_ ^ _39474_ /*31746*/;
assign _39473_ = _39465_ & _39472_ /*31744*/;
assign _39370_ = _39465_ ^ _39472_ /*31745*/;
assign _39470_ = _39471_ | _39473_ /*31742*/;
assign _39479_ = ~D[10] /*31741*/;
assign _39476_ = _38922_ & _39479_ /*31737*/;
assign _39477_ = _38922_ ^ _39479_ /*31740*/;
assign _39478_ = _39470_ & _39477_ /*31738*/;
assign _39371_ = _39470_ ^ _39477_ /*31739*/;
assign _39475_ = _39476_ | _39478_ /*31736*/;
assign _39484_ = ~D[11] /*31735*/;
assign _39481_ = _38923_ & _39484_ /*31731*/;
assign _39482_ = _38923_ ^ _39484_ /*31734*/;
assign _39483_ = _39475_ & _39482_ /*31732*/;
assign _39372_ = _39475_ ^ _39482_ /*31733*/;
assign _39480_ = _39481_ | _39483_ /*31730*/;
assign _39489_ = ~D[12] /*31729*/;
assign _39486_ = _38924_ & _39489_ /*31725*/;
assign _39487_ = _38924_ ^ _39489_ /*31728*/;
assign _39488_ = _39480_ & _39487_ /*31726*/;
assign _39373_ = _39480_ ^ _39487_ /*31727*/;
assign _39485_ = _39486_ | _39488_ /*31724*/;
assign _39494_ = ~D[13] /*31723*/;
assign _39491_ = _38925_ & _39494_ /*31719*/;
assign _39492_ = _38925_ ^ _39494_ /*31722*/;
assign _39493_ = _39485_ & _39492_ /*31720*/;
assign _39374_ = _39485_ ^ _39492_ /*31721*/;
assign _39490_ = _39491_ | _39493_ /*31718*/;
assign _39499_ = ~D[14] /*31717*/;
assign _39496_ = _38926_ & _39499_ /*31713*/;
assign _39497_ = _38926_ ^ _39499_ /*31716*/;
assign _39498_ = _39490_ & _39497_ /*31714*/;
assign _39375_ = _39490_ ^ _39497_ /*31715*/;
assign _39495_ = _39496_ | _39498_ /*31712*/;
assign _39504_ = ~D[15] /*31711*/;
assign _39501_ = _38927_ & _39504_ /*31707*/;
assign _39502_ = _38927_ ^ _39504_ /*31710*/;
assign _39503_ = _39495_ & _39502_ /*31708*/;
assign _39376_ = _39495_ ^ _39502_ /*31709*/;
assign _39500_ = _39501_ | _39503_ /*31706*/;
assign _39509_ = ~D[16] /*31705*/;
assign _39506_ = _38928_ & _39509_ /*31701*/;
assign _39507_ = _38928_ ^ _39509_ /*31704*/;
assign _39508_ = _39500_ & _39507_ /*31702*/;
assign _39377_ = _39500_ ^ _39507_ /*31703*/;
assign _39505_ = _39506_ | _39508_ /*31700*/;
assign _39514_ = ~D[17] /*31699*/;
assign _39511_ = _38929_ & _39514_ /*31695*/;
assign _39512_ = _38929_ ^ _39514_ /*31698*/;
assign _39513_ = _39505_ & _39512_ /*31696*/;
assign _39378_ = _39505_ ^ _39512_ /*31697*/;
assign _39510_ = _39511_ | _39513_ /*31694*/;
assign _39519_ = ~D[18] /*31693*/;
assign _39516_ = _38930_ & _39519_ /*31689*/;
assign _39517_ = _38930_ ^ _39519_ /*31692*/;
assign _39518_ = _39510_ & _39517_ /*31690*/;
assign _39379_ = _39510_ ^ _39517_ /*31691*/;
assign _39515_ = _39516_ | _39518_ /*31688*/;
assign _39524_ = ~D[19] /*31687*/;
assign _39521_ = _38931_ & _39524_ /*31683*/;
assign _39522_ = _38931_ ^ _39524_ /*31686*/;
assign _39523_ = _39515_ & _39522_ /*31684*/;
assign _39380_ = _39515_ ^ _39522_ /*31685*/;
assign _39520_ = _39521_ | _39523_ /*31682*/;
assign _39529_ = ~D[20] /*31681*/;
assign _39526_ = _38932_ & _39529_ /*31677*/;
assign _39527_ = _38932_ ^ _39529_ /*31680*/;
assign _39528_ = _39520_ & _39527_ /*31678*/;
assign _39381_ = _39520_ ^ _39527_ /*31679*/;
assign _39525_ = _39526_ | _39528_ /*31676*/;
assign _39534_ = ~D[21] /*31675*/;
assign _39531_ = _38933_ & _39534_ /*31671*/;
assign _39532_ = _38933_ ^ _39534_ /*31674*/;
assign _39533_ = _39525_ & _39532_ /*31672*/;
assign _39382_ = _39525_ ^ _39532_ /*31673*/;
assign _39530_ = _39531_ | _39533_ /*31670*/;
assign _39539_ = ~D[22] /*31669*/;
assign _39536_ = _38934_ & _39539_ /*31665*/;
assign _39537_ = _38934_ ^ _39539_ /*31668*/;
assign _39538_ = _39530_ & _39537_ /*31666*/;
assign _39383_ = _39530_ ^ _39537_ /*31667*/;
assign _39535_ = _39536_ | _39538_ /*31664*/;
assign _39544_ = ~D[23] /*31663*/;
assign _39541_ = _38935_ & _39544_ /*31659*/;
assign _39542_ = _38935_ ^ _39544_ /*31662*/;
assign _39543_ = _39535_ & _39542_ /*31660*/;
assign _39384_ = _39535_ ^ _39542_ /*31661*/;
assign _39540_ = _39541_ | _39543_ /*31658*/;
assign _39549_ = ~D[24] /*31657*/;
assign _39546_ = _38936_ & _39549_ /*31653*/;
assign _39547_ = _38936_ ^ _39549_ /*31656*/;
assign _39548_ = _39540_ & _39547_ /*31654*/;
assign _39385_ = _39540_ ^ _39547_ /*31655*/;
assign _39545_ = _39546_ | _39548_ /*31652*/;
assign _39554_ = ~D[25] /*31651*/;
assign _39551_ = _38937_ & _39554_ /*31647*/;
assign _39552_ = _38937_ ^ _39554_ /*31650*/;
assign _39553_ = _39545_ & _39552_ /*31648*/;
assign _39386_ = _39545_ ^ _39552_ /*31649*/;
assign _39550_ = _39551_ | _39553_ /*31646*/;
assign _39559_ = ~D[26] /*31645*/;
assign _39556_ = _38938_ & _39559_ /*31641*/;
assign _39557_ = _38938_ ^ _39559_ /*31644*/;
assign _39558_ = _39550_ & _39557_ /*31642*/;
assign _39387_ = _39550_ ^ _39557_ /*31643*/;
assign _39555_ = _39556_ | _39558_ /*31640*/;
assign _39564_ = ~D[27] /*31639*/;
assign _39561_ = _38939_ & _39564_ /*31635*/;
assign _39562_ = _38939_ ^ _39564_ /*31638*/;
assign _39563_ = _39555_ & _39562_ /*31636*/;
assign _39388_ = _39555_ ^ _39562_ /*31637*/;
assign _39560_ = _39561_ | _39563_ /*31634*/;
assign _39569_ = ~D[28] /*31633*/;
assign _39566_ = _38940_ & _39569_ /*31629*/;
assign _39567_ = _38940_ ^ _39569_ /*31632*/;
assign _39568_ = _39560_ & _39567_ /*31630*/;
assign _39389_ = _39560_ ^ _39567_ /*31631*/;
assign _39565_ = _39566_ | _39568_ /*31628*/;
assign _39574_ = ~D[29] /*31627*/;
assign _39571_ = _38941_ & _39574_ /*31623*/;
assign _39572_ = _38941_ ^ _39574_ /*31626*/;
assign _39573_ = _39565_ & _39572_ /*31624*/;
assign _39390_ = _39565_ ^ _39572_ /*31625*/;
assign _39570_ = _39571_ | _39573_ /*31622*/;
assign _39579_ = ~D[30] /*31621*/;
assign _39576_ = _38942_ & _39579_ /*31617*/;
assign _39577_ = _38942_ ^ _39579_ /*31620*/;
assign _39578_ = _39570_ & _39577_ /*31618*/;
assign _39391_ = _39570_ ^ _39577_ /*31619*/;
assign _39575_ = _39576_ | _39578_ /*31616*/;
assign _39584_ = ~D[31] /*31615*/;
assign _39581_ = _38943_ & _39584_ /*31611*/;
assign _39582_ = _38943_ ^ _39584_ /*31614*/;
assign _39583_ = _39575_ & _39582_ /*31612*/;
assign _39392_ = _39575_ ^ _39582_ /*31613*/;
assign _39580_ = _39581_ | _39583_ /*31610*/;
assign _39589_ = ~D[32] /*31609*/;
assign _39586_ = _38944_ & _39589_ /*31605*/;
assign _39587_ = _38944_ ^ _39589_ /*31608*/;
assign _39588_ = _39580_ & _39587_ /*31606*/;
assign _39393_ = _39580_ ^ _39587_ /*31607*/;
assign _39585_ = _39586_ | _39588_ /*31604*/;
assign _39594_ = ~D[33] /*31603*/;
assign _39591_ = _38945_ & _39594_ /*31599*/;
assign _39592_ = _38945_ ^ _39594_ /*31602*/;
assign _39593_ = _39585_ & _39592_ /*31600*/;
assign _39394_ = _39585_ ^ _39592_ /*31601*/;
assign _39590_ = _39591_ | _39593_ /*31598*/;
assign _39599_ = ~D[34] /*31597*/;
assign _39596_ = _38946_ & _39599_ /*31593*/;
assign _39597_ = _38946_ ^ _39599_ /*31596*/;
assign _39598_ = _39590_ & _39597_ /*31594*/;
assign _39395_ = _39590_ ^ _39597_ /*31595*/;
assign _39595_ = _39596_ | _39598_ /*31592*/;
assign _39604_ = ~D[35] /*31591*/;
assign _39601_ = _38947_ & _39604_ /*31587*/;
assign _39602_ = _38947_ ^ _39604_ /*31590*/;
assign _39603_ = _39595_ & _39602_ /*31588*/;
assign _39396_ = _39595_ ^ _39602_ /*31589*/;
assign _39600_ = _39601_ | _39603_ /*31586*/;
assign _39609_ = ~D[36] /*31585*/;
assign _39606_ = _38948_ & _39609_ /*31581*/;
assign _39607_ = _38948_ ^ _39609_ /*31584*/;
assign _39608_ = _39600_ & _39607_ /*31582*/;
assign _39397_ = _39600_ ^ _39607_ /*31583*/;
assign _39605_ = _39606_ | _39608_ /*31580*/;
assign _39614_ = ~D[37] /*31579*/;
assign _39611_ = _38949_ & _39614_ /*31575*/;
assign _39612_ = _38949_ ^ _39614_ /*31578*/;
assign _39613_ = _39605_ & _39612_ /*31576*/;
assign _39398_ = _39605_ ^ _39612_ /*31577*/;
assign _39610_ = _39611_ | _39613_ /*31574*/;
assign _39619_ = ~D[38] /*31573*/;
assign _39616_ = _38950_ & _39619_ /*31569*/;
assign _39617_ = _38950_ ^ _39619_ /*31572*/;
assign _39618_ = _39610_ & _39617_ /*31570*/;
assign _39399_ = _39610_ ^ _39617_ /*31571*/;
assign _39615_ = _39616_ | _39618_ /*31568*/;
assign _39624_ = ~D[39] /*31567*/;
assign _39621_ = _38951_ & _39624_ /*31563*/;
assign _39622_ = _38951_ ^ _39624_ /*31566*/;
assign _39623_ = _39615_ & _39622_ /*31564*/;
assign _39400_ = _39615_ ^ _39622_ /*31565*/;
assign _39620_ = _39621_ | _39623_ /*31562*/;
assign _39629_ = ~D[40] /*31561*/;
assign _39626_ = _38952_ & _39629_ /*31557*/;
assign _39627_ = _38952_ ^ _39629_ /*31560*/;
assign _39628_ = _39620_ & _39627_ /*31558*/;
assign _39401_ = _39620_ ^ _39627_ /*31559*/;
assign _39625_ = _39626_ | _39628_ /*31556*/;
assign _39634_ = ~D[41] /*31555*/;
assign _39631_ = _38953_ & _39634_ /*31551*/;
assign _39632_ = _38953_ ^ _39634_ /*31554*/;
assign _39633_ = _39625_ & _39632_ /*31552*/;
assign _39402_ = _39625_ ^ _39632_ /*31553*/;
assign _39630_ = _39631_ | _39633_ /*31550*/;
assign _39639_ = ~D[42] /*31549*/;
assign _39636_ = _38954_ & _39639_ /*31545*/;
assign _39637_ = _38954_ ^ _39639_ /*31548*/;
assign _39638_ = _39630_ & _39637_ /*31546*/;
assign _39403_ = _39630_ ^ _39637_ /*31547*/;
assign _39635_ = _39636_ | _39638_ /*31544*/;
assign _39644_ = ~D[43] /*31543*/;
assign _39641_ = _38955_ & _39644_ /*31539*/;
assign _39642_ = _38955_ ^ _39644_ /*31542*/;
assign _39643_ = _39635_ & _39642_ /*31540*/;
assign _39404_ = _39635_ ^ _39642_ /*31541*/;
assign _39640_ = _39641_ | _39643_ /*31538*/;
assign _39649_ = ~D[44] /*31537*/;
assign _39646_ = _38956_ & _39649_ /*31533*/;
assign _39647_ = _38956_ ^ _39649_ /*31536*/;
assign _39648_ = _39640_ & _39647_ /*31534*/;
assign _39405_ = _39640_ ^ _39647_ /*31535*/;
assign _39645_ = _39646_ | _39648_ /*31532*/;
assign _39654_ = ~D[45] /*31531*/;
assign _39651_ = _38957_ & _39654_ /*31527*/;
assign _39652_ = _38957_ ^ _39654_ /*31530*/;
assign _39653_ = _39645_ & _39652_ /*31528*/;
assign _39406_ = _39645_ ^ _39652_ /*31529*/;
assign _39650_ = _39651_ | _39653_ /*31526*/;
assign _39659_ = ~D[46] /*31525*/;
assign _39656_ = _38958_ & _39659_ /*31521*/;
assign _39657_ = _38958_ ^ _39659_ /*31524*/;
assign _39658_ = _39650_ & _39657_ /*31522*/;
assign _39407_ = _39650_ ^ _39657_ /*31523*/;
assign _39655_ = _39656_ | _39658_ /*31520*/;
assign _39664_ = ~D[47] /*31519*/;
assign _39661_ = _38959_ & _39664_ /*31515*/;
assign _39662_ = _38959_ ^ _39664_ /*31518*/;
assign _39663_ = _39655_ & _39662_ /*31516*/;
assign _39408_ = _39655_ ^ _39662_ /*31517*/;
assign _39660_ = _39661_ | _39663_ /*31514*/;
assign _39669_ = ~D[48] /*31513*/;
assign _39666_ = _38960_ & _39669_ /*31509*/;
assign _39667_ = _38960_ ^ _39669_ /*31512*/;
assign _39668_ = _39660_ & _39667_ /*31510*/;
assign _39409_ = _39660_ ^ _39667_ /*31511*/;
assign _39665_ = _39666_ | _39668_ /*31508*/;
assign _39674_ = ~D[49] /*31507*/;
assign _39671_ = _38961_ & _39674_ /*31503*/;
assign _39672_ = _38961_ ^ _39674_ /*31506*/;
assign _39673_ = _39665_ & _39672_ /*31504*/;
assign _39410_ = _39665_ ^ _39672_ /*31505*/;
assign _39670_ = _39671_ | _39673_ /*31502*/;
assign _39679_ = ~D[50] /*31501*/;
assign _39676_ = _38962_ & _39679_ /*31497*/;
assign _39677_ = _38962_ ^ _39679_ /*31500*/;
assign _39678_ = _39670_ & _39677_ /*31498*/;
assign _39411_ = _39670_ ^ _39677_ /*31499*/;
assign _39675_ = _39676_ | _39678_ /*31496*/;
assign _39684_ = ~D[51] /*31495*/;
assign _39681_ = _38963_ & _39684_ /*31491*/;
assign _39682_ = _38963_ ^ _39684_ /*31494*/;
assign _39683_ = _39675_ & _39682_ /*31492*/;
assign _39412_ = _39675_ ^ _39682_ /*31493*/;
assign _39680_ = _39681_ | _39683_ /*31490*/;
assign _39689_ = ~D[52] /*31489*/;
assign _39686_ = _38964_ & _39689_ /*31485*/;
assign _39687_ = _38964_ ^ _39689_ /*31488*/;
assign _39688_ = _39680_ & _39687_ /*31486*/;
assign _39413_ = _39680_ ^ _39687_ /*31487*/;
assign _39685_ = _39686_ | _39688_ /*31484*/;
assign _39694_ = ~D[53] /*31483*/;
assign _39691_ = _38965_ & _39694_ /*31479*/;
assign _39692_ = _38965_ ^ _39694_ /*31482*/;
assign _39693_ = _39685_ & _39692_ /*31480*/;
assign _39414_ = _39685_ ^ _39692_ /*31481*/;
assign _39690_ = _39691_ | _39693_ /*31478*/;
assign _39699_ = ~D[54] /*31477*/;
assign _39696_ = _38966_ & _39699_ /*31473*/;
assign _39697_ = _38966_ ^ _39699_ /*31476*/;
assign _39698_ = _39690_ & _39697_ /*31474*/;
assign _39415_ = _39690_ ^ _39697_ /*31475*/;
assign _39695_ = _39696_ | _39698_ /*31472*/;
assign _39704_ = ~D[55] /*31471*/;
assign _39701_ = _38967_ & _39704_ /*31467*/;
assign _39702_ = _38967_ ^ _39704_ /*31470*/;
assign _39703_ = _39695_ & _39702_ /*31468*/;
assign _39416_ = _39695_ ^ _39702_ /*31469*/;
assign _39700_ = _39701_ | _39703_ /*31466*/;
assign _39709_ = ~D[56] /*31465*/;
assign _39706_ = _38968_ & _39709_ /*31461*/;
assign _39707_ = _38968_ ^ _39709_ /*31464*/;
assign _39708_ = _39700_ & _39707_ /*31462*/;
assign _39417_ = _39700_ ^ _39707_ /*31463*/;
assign _39705_ = _39706_ | _39708_ /*31460*/;
assign _39714_ = ~D[57] /*31459*/;
assign _39711_ = _38969_ & _39714_ /*31455*/;
assign _39712_ = _38969_ ^ _39714_ /*31458*/;
assign _39713_ = _39705_ & _39712_ /*31456*/;
assign _39418_ = _39705_ ^ _39712_ /*31457*/;
assign _39710_ = _39711_ | _39713_ /*31454*/;
assign _39719_ = ~D[58] /*31453*/;
assign _39716_ = _38970_ & _39719_ /*31449*/;
assign _39717_ = _38970_ ^ _39719_ /*31452*/;
assign _39718_ = _39710_ & _39717_ /*31450*/;
assign _39419_ = _39710_ ^ _39717_ /*31451*/;
assign _39715_ = _39716_ | _39718_ /*31448*/;
assign _39724_ = ~D[59] /*31447*/;
assign _39721_ = _38971_ & _39724_ /*31443*/;
assign _39722_ = _38971_ ^ _39724_ /*31446*/;
assign _39723_ = _39715_ & _39722_ /*31444*/;
assign _39420_ = _39715_ ^ _39722_ /*31445*/;
assign _39720_ = _39721_ | _39723_ /*31442*/;
assign _39729_ = ~D[60] /*31441*/;
assign _39726_ = _38972_ & _39729_ /*31437*/;
assign _39727_ = _38972_ ^ _39729_ /*31440*/;
assign _39728_ = _39720_ & _39727_ /*31438*/;
assign _39421_ = _39720_ ^ _39727_ /*31439*/;
assign _39725_ = _39726_ | _39728_ /*31436*/;
assign _39734_ = ~D[61] /*31435*/;
assign _39731_ = _38973_ & _39734_ /*31431*/;
assign _39732_ = _38973_ ^ _39734_ /*31434*/;
assign _39733_ = _39725_ & _39732_ /*31432*/;
assign _39422_ = _39725_ ^ _39732_ /*31433*/;
assign _39730_ = _39731_ | _39733_ /*31430*/;
assign _39739_ = ~D[62] /*31429*/;
assign _39736_ = _38974_ & _39739_ /*31425*/;
assign _39737_ = _38974_ ^ _39739_ /*31428*/;
assign _39738_ = _39730_ & _39737_ /*31426*/;
assign _39423_ = _39730_ ^ _39737_ /*31427*/;
assign _39735_ = _39736_ | _39738_ /*31424*/;
assign _39740_ = _38975_ & oneWire /*31419*/;
assign _39741_ = _38975_ ^ oneWire /*31422*/;
assign _39742_ = _39735_ & _39741_ /*31420*/;
assign _39424_ = _39735_ ^ _39741_ /*31421*/;
assign Q[19] = _39740_ | _39742_ /*31418*/;
assign _39875_ = ~Q[19] /*31033*/;
assign _39874_ = _39875_ & D[0] /*31032*/;
assign _39877_ = _39361_ & _39874_ /*31027*/;
assign _39878_ = _39361_ ^ _39874_ /*31030*/;
assign _39879_ = zeroWire & _39878_ /*31028*/;
assign _39809_ = zeroWire ^ _39878_ /*31029*/;
assign _39876_ = _39877_ | _39879_ /*31026*/;
assign _39881_ = ~Q[19] /*31025*/;
assign _39880_ = _39881_ & D[1] /*31024*/;
assign _39883_ = _39362_ & _39880_ /*31019*/;
assign _39884_ = _39362_ ^ _39880_ /*31022*/;
assign _39885_ = _39876_ & _39884_ /*31020*/;
assign _39810_ = _39876_ ^ _39884_ /*31021*/;
assign _39882_ = _39883_ | _39885_ /*31018*/;
assign _39887_ = ~Q[19] /*31017*/;
assign _39886_ = _39887_ & D[2] /*31016*/;
assign _39889_ = _39363_ & _39886_ /*31011*/;
assign _39890_ = _39363_ ^ _39886_ /*31014*/;
assign _39891_ = _39882_ & _39890_ /*31012*/;
assign _39811_ = _39882_ ^ _39890_ /*31013*/;
assign _39888_ = _39889_ | _39891_ /*31010*/;
assign _39893_ = ~Q[19] /*31009*/;
assign _39892_ = _39893_ & D[3] /*31008*/;
assign _39895_ = _39364_ & _39892_ /*31003*/;
assign _39896_ = _39364_ ^ _39892_ /*31006*/;
assign _39897_ = _39888_ & _39896_ /*31004*/;
assign _39812_ = _39888_ ^ _39896_ /*31005*/;
assign _39894_ = _39895_ | _39897_ /*31002*/;
assign _39899_ = ~Q[19] /*31001*/;
assign _39898_ = _39899_ & D[4] /*31000*/;
assign _39901_ = _39365_ & _39898_ /*30995*/;
assign _39902_ = _39365_ ^ _39898_ /*30998*/;
assign _39903_ = _39894_ & _39902_ /*30996*/;
assign _39813_ = _39894_ ^ _39902_ /*30997*/;
assign _39900_ = _39901_ | _39903_ /*30994*/;
assign _39905_ = ~Q[19] /*30993*/;
assign _39904_ = _39905_ & D[5] /*30992*/;
assign _39907_ = _39366_ & _39904_ /*30987*/;
assign _39908_ = _39366_ ^ _39904_ /*30990*/;
assign _39909_ = _39900_ & _39908_ /*30988*/;
assign _39814_ = _39900_ ^ _39908_ /*30989*/;
assign _39906_ = _39907_ | _39909_ /*30986*/;
assign _39911_ = ~Q[19] /*30985*/;
assign _39910_ = _39911_ & D[6] /*30984*/;
assign _39913_ = _39367_ & _39910_ /*30979*/;
assign _39914_ = _39367_ ^ _39910_ /*30982*/;
assign _39915_ = _39906_ & _39914_ /*30980*/;
assign _39815_ = _39906_ ^ _39914_ /*30981*/;
assign _39912_ = _39913_ | _39915_ /*30978*/;
assign _39917_ = ~Q[19] /*30977*/;
assign _39916_ = _39917_ & D[7] /*30976*/;
assign _39919_ = _39368_ & _39916_ /*30971*/;
assign _39920_ = _39368_ ^ _39916_ /*30974*/;
assign _39921_ = _39912_ & _39920_ /*30972*/;
assign _39816_ = _39912_ ^ _39920_ /*30973*/;
assign _39918_ = _39919_ | _39921_ /*30970*/;
assign _39923_ = ~Q[19] /*30969*/;
assign _39922_ = _39923_ & D[8] /*30968*/;
assign _39925_ = _39369_ & _39922_ /*30963*/;
assign _39926_ = _39369_ ^ _39922_ /*30966*/;
assign _39927_ = _39918_ & _39926_ /*30964*/;
assign _39817_ = _39918_ ^ _39926_ /*30965*/;
assign _39924_ = _39925_ | _39927_ /*30962*/;
assign _39929_ = ~Q[19] /*30961*/;
assign _39928_ = _39929_ & D[9] /*30960*/;
assign _39931_ = _39370_ & _39928_ /*30955*/;
assign _39932_ = _39370_ ^ _39928_ /*30958*/;
assign _39933_ = _39924_ & _39932_ /*30956*/;
assign _39818_ = _39924_ ^ _39932_ /*30957*/;
assign _39930_ = _39931_ | _39933_ /*30954*/;
assign _39935_ = ~Q[19] /*30953*/;
assign _39934_ = _39935_ & D[10] /*30952*/;
assign _39937_ = _39371_ & _39934_ /*30947*/;
assign _39938_ = _39371_ ^ _39934_ /*30950*/;
assign _39939_ = _39930_ & _39938_ /*30948*/;
assign _39819_ = _39930_ ^ _39938_ /*30949*/;
assign _39936_ = _39937_ | _39939_ /*30946*/;
assign _39941_ = ~Q[19] /*30945*/;
assign _39940_ = _39941_ & D[11] /*30944*/;
assign _39943_ = _39372_ & _39940_ /*30939*/;
assign _39944_ = _39372_ ^ _39940_ /*30942*/;
assign _39945_ = _39936_ & _39944_ /*30940*/;
assign _39820_ = _39936_ ^ _39944_ /*30941*/;
assign _39942_ = _39943_ | _39945_ /*30938*/;
assign _39947_ = ~Q[19] /*30937*/;
assign _39946_ = _39947_ & D[12] /*30936*/;
assign _39949_ = _39373_ & _39946_ /*30931*/;
assign _39950_ = _39373_ ^ _39946_ /*30934*/;
assign _39951_ = _39942_ & _39950_ /*30932*/;
assign _39821_ = _39942_ ^ _39950_ /*30933*/;
assign _39948_ = _39949_ | _39951_ /*30930*/;
assign _39953_ = ~Q[19] /*30929*/;
assign _39952_ = _39953_ & D[13] /*30928*/;
assign _39955_ = _39374_ & _39952_ /*30923*/;
assign _39956_ = _39374_ ^ _39952_ /*30926*/;
assign _39957_ = _39948_ & _39956_ /*30924*/;
assign _39822_ = _39948_ ^ _39956_ /*30925*/;
assign _39954_ = _39955_ | _39957_ /*30922*/;
assign _39959_ = ~Q[19] /*30921*/;
assign _39958_ = _39959_ & D[14] /*30920*/;
assign _39961_ = _39375_ & _39958_ /*30915*/;
assign _39962_ = _39375_ ^ _39958_ /*30918*/;
assign _39963_ = _39954_ & _39962_ /*30916*/;
assign _39823_ = _39954_ ^ _39962_ /*30917*/;
assign _39960_ = _39961_ | _39963_ /*30914*/;
assign _39965_ = ~Q[19] /*30913*/;
assign _39964_ = _39965_ & D[15] /*30912*/;
assign _39967_ = _39376_ & _39964_ /*30907*/;
assign _39968_ = _39376_ ^ _39964_ /*30910*/;
assign _39969_ = _39960_ & _39968_ /*30908*/;
assign _39824_ = _39960_ ^ _39968_ /*30909*/;
assign _39966_ = _39967_ | _39969_ /*30906*/;
assign _39971_ = ~Q[19] /*30905*/;
assign _39970_ = _39971_ & D[16] /*30904*/;
assign _39973_ = _39377_ & _39970_ /*30899*/;
assign _39974_ = _39377_ ^ _39970_ /*30902*/;
assign _39975_ = _39966_ & _39974_ /*30900*/;
assign _39825_ = _39966_ ^ _39974_ /*30901*/;
assign _39972_ = _39973_ | _39975_ /*30898*/;
assign _39977_ = ~Q[19] /*30897*/;
assign _39976_ = _39977_ & D[17] /*30896*/;
assign _39979_ = _39378_ & _39976_ /*30891*/;
assign _39980_ = _39378_ ^ _39976_ /*30894*/;
assign _39981_ = _39972_ & _39980_ /*30892*/;
assign _39826_ = _39972_ ^ _39980_ /*30893*/;
assign _39978_ = _39979_ | _39981_ /*30890*/;
assign _39983_ = ~Q[19] /*30889*/;
assign _39982_ = _39983_ & D[18] /*30888*/;
assign _39985_ = _39379_ & _39982_ /*30883*/;
assign _39986_ = _39379_ ^ _39982_ /*30886*/;
assign _39987_ = _39978_ & _39986_ /*30884*/;
assign _39827_ = _39978_ ^ _39986_ /*30885*/;
assign _39984_ = _39985_ | _39987_ /*30882*/;
assign _39989_ = ~Q[19] /*30881*/;
assign _39988_ = _39989_ & D[19] /*30880*/;
assign _39991_ = _39380_ & _39988_ /*30875*/;
assign _39992_ = _39380_ ^ _39988_ /*30878*/;
assign _39993_ = _39984_ & _39992_ /*30876*/;
assign _39828_ = _39984_ ^ _39992_ /*30877*/;
assign _39990_ = _39991_ | _39993_ /*30874*/;
assign _39995_ = ~Q[19] /*30873*/;
assign _39994_ = _39995_ & D[20] /*30872*/;
assign _39997_ = _39381_ & _39994_ /*30867*/;
assign _39998_ = _39381_ ^ _39994_ /*30870*/;
assign _39999_ = _39990_ & _39998_ /*30868*/;
assign _39829_ = _39990_ ^ _39998_ /*30869*/;
assign _39996_ = _39997_ | _39999_ /*30866*/;
assign _40001_ = ~Q[19] /*30865*/;
assign _40000_ = _40001_ & D[21] /*30864*/;
assign _40003_ = _39382_ & _40000_ /*30859*/;
assign _40004_ = _39382_ ^ _40000_ /*30862*/;
assign _40005_ = _39996_ & _40004_ /*30860*/;
assign _39830_ = _39996_ ^ _40004_ /*30861*/;
assign _40002_ = _40003_ | _40005_ /*30858*/;
assign _40007_ = ~Q[19] /*30857*/;
assign _40006_ = _40007_ & D[22] /*30856*/;
assign _40009_ = _39383_ & _40006_ /*30851*/;
assign _40010_ = _39383_ ^ _40006_ /*30854*/;
assign _40011_ = _40002_ & _40010_ /*30852*/;
assign _39831_ = _40002_ ^ _40010_ /*30853*/;
assign _40008_ = _40009_ | _40011_ /*30850*/;
assign _40013_ = ~Q[19] /*30849*/;
assign _40012_ = _40013_ & D[23] /*30848*/;
assign _40015_ = _39384_ & _40012_ /*30843*/;
assign _40016_ = _39384_ ^ _40012_ /*30846*/;
assign _40017_ = _40008_ & _40016_ /*30844*/;
assign _39832_ = _40008_ ^ _40016_ /*30845*/;
assign _40014_ = _40015_ | _40017_ /*30842*/;
assign _40019_ = ~Q[19] /*30841*/;
assign _40018_ = _40019_ & D[24] /*30840*/;
assign _40021_ = _39385_ & _40018_ /*30835*/;
assign _40022_ = _39385_ ^ _40018_ /*30838*/;
assign _40023_ = _40014_ & _40022_ /*30836*/;
assign _39833_ = _40014_ ^ _40022_ /*30837*/;
assign _40020_ = _40021_ | _40023_ /*30834*/;
assign _40025_ = ~Q[19] /*30833*/;
assign _40024_ = _40025_ & D[25] /*30832*/;
assign _40027_ = _39386_ & _40024_ /*30827*/;
assign _40028_ = _39386_ ^ _40024_ /*30830*/;
assign _40029_ = _40020_ & _40028_ /*30828*/;
assign _39834_ = _40020_ ^ _40028_ /*30829*/;
assign _40026_ = _40027_ | _40029_ /*30826*/;
assign _40031_ = ~Q[19] /*30825*/;
assign _40030_ = _40031_ & D[26] /*30824*/;
assign _40033_ = _39387_ & _40030_ /*30819*/;
assign _40034_ = _39387_ ^ _40030_ /*30822*/;
assign _40035_ = _40026_ & _40034_ /*30820*/;
assign _39835_ = _40026_ ^ _40034_ /*30821*/;
assign _40032_ = _40033_ | _40035_ /*30818*/;
assign _40037_ = ~Q[19] /*30817*/;
assign _40036_ = _40037_ & D[27] /*30816*/;
assign _40039_ = _39388_ & _40036_ /*30811*/;
assign _40040_ = _39388_ ^ _40036_ /*30814*/;
assign _40041_ = _40032_ & _40040_ /*30812*/;
assign _39836_ = _40032_ ^ _40040_ /*30813*/;
assign _40038_ = _40039_ | _40041_ /*30810*/;
assign _40043_ = ~Q[19] /*30809*/;
assign _40042_ = _40043_ & D[28] /*30808*/;
assign _40045_ = _39389_ & _40042_ /*30803*/;
assign _40046_ = _39389_ ^ _40042_ /*30806*/;
assign _40047_ = _40038_ & _40046_ /*30804*/;
assign _39837_ = _40038_ ^ _40046_ /*30805*/;
assign _40044_ = _40045_ | _40047_ /*30802*/;
assign _40049_ = ~Q[19] /*30801*/;
assign _40048_ = _40049_ & D[29] /*30800*/;
assign _40051_ = _39390_ & _40048_ /*30795*/;
assign _40052_ = _39390_ ^ _40048_ /*30798*/;
assign _40053_ = _40044_ & _40052_ /*30796*/;
assign _39838_ = _40044_ ^ _40052_ /*30797*/;
assign _40050_ = _40051_ | _40053_ /*30794*/;
assign _40055_ = ~Q[19] /*30793*/;
assign _40054_ = _40055_ & D[30] /*30792*/;
assign _40057_ = _39391_ & _40054_ /*30787*/;
assign _40058_ = _39391_ ^ _40054_ /*30790*/;
assign _40059_ = _40050_ & _40058_ /*30788*/;
assign _39839_ = _40050_ ^ _40058_ /*30789*/;
assign _40056_ = _40057_ | _40059_ /*30786*/;
assign _40061_ = ~Q[19] /*30785*/;
assign _40060_ = _40061_ & D[31] /*30784*/;
assign _40063_ = _39392_ & _40060_ /*30779*/;
assign _40064_ = _39392_ ^ _40060_ /*30782*/;
assign _40065_ = _40056_ & _40064_ /*30780*/;
assign _39840_ = _40056_ ^ _40064_ /*30781*/;
assign _40062_ = _40063_ | _40065_ /*30778*/;
assign _40067_ = ~Q[19] /*30777*/;
assign _40066_ = _40067_ & D[32] /*30776*/;
assign _40069_ = _39393_ & _40066_ /*30771*/;
assign _40070_ = _39393_ ^ _40066_ /*30774*/;
assign _40071_ = _40062_ & _40070_ /*30772*/;
assign _39841_ = _40062_ ^ _40070_ /*30773*/;
assign _40068_ = _40069_ | _40071_ /*30770*/;
assign _40073_ = ~Q[19] /*30769*/;
assign _40072_ = _40073_ & D[33] /*30768*/;
assign _40075_ = _39394_ & _40072_ /*30763*/;
assign _40076_ = _39394_ ^ _40072_ /*30766*/;
assign _40077_ = _40068_ & _40076_ /*30764*/;
assign _39842_ = _40068_ ^ _40076_ /*30765*/;
assign _40074_ = _40075_ | _40077_ /*30762*/;
assign _40079_ = ~Q[19] /*30761*/;
assign _40078_ = _40079_ & D[34] /*30760*/;
assign _40081_ = _39395_ & _40078_ /*30755*/;
assign _40082_ = _39395_ ^ _40078_ /*30758*/;
assign _40083_ = _40074_ & _40082_ /*30756*/;
assign _39843_ = _40074_ ^ _40082_ /*30757*/;
assign _40080_ = _40081_ | _40083_ /*30754*/;
assign _40085_ = ~Q[19] /*30753*/;
assign _40084_ = _40085_ & D[35] /*30752*/;
assign _40087_ = _39396_ & _40084_ /*30747*/;
assign _40088_ = _39396_ ^ _40084_ /*30750*/;
assign _40089_ = _40080_ & _40088_ /*30748*/;
assign _39844_ = _40080_ ^ _40088_ /*30749*/;
assign _40086_ = _40087_ | _40089_ /*30746*/;
assign _40091_ = ~Q[19] /*30745*/;
assign _40090_ = _40091_ & D[36] /*30744*/;
assign _40093_ = _39397_ & _40090_ /*30739*/;
assign _40094_ = _39397_ ^ _40090_ /*30742*/;
assign _40095_ = _40086_ & _40094_ /*30740*/;
assign _39845_ = _40086_ ^ _40094_ /*30741*/;
assign _40092_ = _40093_ | _40095_ /*30738*/;
assign _40097_ = ~Q[19] /*30737*/;
assign _40096_ = _40097_ & D[37] /*30736*/;
assign _40099_ = _39398_ & _40096_ /*30731*/;
assign _40100_ = _39398_ ^ _40096_ /*30734*/;
assign _40101_ = _40092_ & _40100_ /*30732*/;
assign _39846_ = _40092_ ^ _40100_ /*30733*/;
assign _40098_ = _40099_ | _40101_ /*30730*/;
assign _40103_ = ~Q[19] /*30729*/;
assign _40102_ = _40103_ & D[38] /*30728*/;
assign _40105_ = _39399_ & _40102_ /*30723*/;
assign _40106_ = _39399_ ^ _40102_ /*30726*/;
assign _40107_ = _40098_ & _40106_ /*30724*/;
assign _39847_ = _40098_ ^ _40106_ /*30725*/;
assign _40104_ = _40105_ | _40107_ /*30722*/;
assign _40109_ = ~Q[19] /*30721*/;
assign _40108_ = _40109_ & D[39] /*30720*/;
assign _40111_ = _39400_ & _40108_ /*30715*/;
assign _40112_ = _39400_ ^ _40108_ /*30718*/;
assign _40113_ = _40104_ & _40112_ /*30716*/;
assign _39848_ = _40104_ ^ _40112_ /*30717*/;
assign _40110_ = _40111_ | _40113_ /*30714*/;
assign _40115_ = ~Q[19] /*30713*/;
assign _40114_ = _40115_ & D[40] /*30712*/;
assign _40117_ = _39401_ & _40114_ /*30707*/;
assign _40118_ = _39401_ ^ _40114_ /*30710*/;
assign _40119_ = _40110_ & _40118_ /*30708*/;
assign _39849_ = _40110_ ^ _40118_ /*30709*/;
assign _40116_ = _40117_ | _40119_ /*30706*/;
assign _40121_ = ~Q[19] /*30705*/;
assign _40120_ = _40121_ & D[41] /*30704*/;
assign _40123_ = _39402_ & _40120_ /*30699*/;
assign _40124_ = _39402_ ^ _40120_ /*30702*/;
assign _40125_ = _40116_ & _40124_ /*30700*/;
assign _39850_ = _40116_ ^ _40124_ /*30701*/;
assign _40122_ = _40123_ | _40125_ /*30698*/;
assign _40127_ = ~Q[19] /*30697*/;
assign _40126_ = _40127_ & D[42] /*30696*/;
assign _40129_ = _39403_ & _40126_ /*30691*/;
assign _40130_ = _39403_ ^ _40126_ /*30694*/;
assign _40131_ = _40122_ & _40130_ /*30692*/;
assign _39851_ = _40122_ ^ _40130_ /*30693*/;
assign _40128_ = _40129_ | _40131_ /*30690*/;
assign _40133_ = ~Q[19] /*30689*/;
assign _40132_ = _40133_ & D[43] /*30688*/;
assign _40135_ = _39404_ & _40132_ /*30683*/;
assign _40136_ = _39404_ ^ _40132_ /*30686*/;
assign _40137_ = _40128_ & _40136_ /*30684*/;
assign _39852_ = _40128_ ^ _40136_ /*30685*/;
assign _40134_ = _40135_ | _40137_ /*30682*/;
assign _40139_ = ~Q[19] /*30681*/;
assign _40138_ = _40139_ & D[44] /*30680*/;
assign _40141_ = _39405_ & _40138_ /*30675*/;
assign _40142_ = _39405_ ^ _40138_ /*30678*/;
assign _40143_ = _40134_ & _40142_ /*30676*/;
assign _39853_ = _40134_ ^ _40142_ /*30677*/;
assign _40140_ = _40141_ | _40143_ /*30674*/;
assign _40145_ = ~Q[19] /*30673*/;
assign _40144_ = _40145_ & D[45] /*30672*/;
assign _40147_ = _39406_ & _40144_ /*30667*/;
assign _40148_ = _39406_ ^ _40144_ /*30670*/;
assign _40149_ = _40140_ & _40148_ /*30668*/;
assign _39854_ = _40140_ ^ _40148_ /*30669*/;
assign _40146_ = _40147_ | _40149_ /*30666*/;
assign _40151_ = ~Q[19] /*30665*/;
assign _40150_ = _40151_ & D[46] /*30664*/;
assign _40153_ = _39407_ & _40150_ /*30659*/;
assign _40154_ = _39407_ ^ _40150_ /*30662*/;
assign _40155_ = _40146_ & _40154_ /*30660*/;
assign _39855_ = _40146_ ^ _40154_ /*30661*/;
assign _40152_ = _40153_ | _40155_ /*30658*/;
assign _40157_ = ~Q[19] /*30657*/;
assign _40156_ = _40157_ & D[47] /*30656*/;
assign _40159_ = _39408_ & _40156_ /*30651*/;
assign _40160_ = _39408_ ^ _40156_ /*30654*/;
assign _40161_ = _40152_ & _40160_ /*30652*/;
assign _39856_ = _40152_ ^ _40160_ /*30653*/;
assign _40158_ = _40159_ | _40161_ /*30650*/;
assign _40163_ = ~Q[19] /*30649*/;
assign _40162_ = _40163_ & D[48] /*30648*/;
assign _40165_ = _39409_ & _40162_ /*30643*/;
assign _40166_ = _39409_ ^ _40162_ /*30646*/;
assign _40167_ = _40158_ & _40166_ /*30644*/;
assign _39857_ = _40158_ ^ _40166_ /*30645*/;
assign _40164_ = _40165_ | _40167_ /*30642*/;
assign _40169_ = ~Q[19] /*30641*/;
assign _40168_ = _40169_ & D[49] /*30640*/;
assign _40171_ = _39410_ & _40168_ /*30635*/;
assign _40172_ = _39410_ ^ _40168_ /*30638*/;
assign _40173_ = _40164_ & _40172_ /*30636*/;
assign _39858_ = _40164_ ^ _40172_ /*30637*/;
assign _40170_ = _40171_ | _40173_ /*30634*/;
assign _40175_ = ~Q[19] /*30633*/;
assign _40174_ = _40175_ & D[50] /*30632*/;
assign _40177_ = _39411_ & _40174_ /*30627*/;
assign _40178_ = _39411_ ^ _40174_ /*30630*/;
assign _40179_ = _40170_ & _40178_ /*30628*/;
assign _39859_ = _40170_ ^ _40178_ /*30629*/;
assign _40176_ = _40177_ | _40179_ /*30626*/;
assign _40181_ = ~Q[19] /*30625*/;
assign _40180_ = _40181_ & D[51] /*30624*/;
assign _40183_ = _39412_ & _40180_ /*30619*/;
assign _40184_ = _39412_ ^ _40180_ /*30622*/;
assign _40185_ = _40176_ & _40184_ /*30620*/;
assign _39860_ = _40176_ ^ _40184_ /*30621*/;
assign _40182_ = _40183_ | _40185_ /*30618*/;
assign _40187_ = ~Q[19] /*30617*/;
assign _40186_ = _40187_ & D[52] /*30616*/;
assign _40189_ = _39413_ & _40186_ /*30611*/;
assign _40190_ = _39413_ ^ _40186_ /*30614*/;
assign _40191_ = _40182_ & _40190_ /*30612*/;
assign _39861_ = _40182_ ^ _40190_ /*30613*/;
assign _40188_ = _40189_ | _40191_ /*30610*/;
assign _40193_ = ~Q[19] /*30609*/;
assign _40192_ = _40193_ & D[53] /*30608*/;
assign _40195_ = _39414_ & _40192_ /*30603*/;
assign _40196_ = _39414_ ^ _40192_ /*30606*/;
assign _40197_ = _40188_ & _40196_ /*30604*/;
assign _39862_ = _40188_ ^ _40196_ /*30605*/;
assign _40194_ = _40195_ | _40197_ /*30602*/;
assign _40199_ = ~Q[19] /*30601*/;
assign _40198_ = _40199_ & D[54] /*30600*/;
assign _40201_ = _39415_ & _40198_ /*30595*/;
assign _40202_ = _39415_ ^ _40198_ /*30598*/;
assign _40203_ = _40194_ & _40202_ /*30596*/;
assign _39863_ = _40194_ ^ _40202_ /*30597*/;
assign _40200_ = _40201_ | _40203_ /*30594*/;
assign _40205_ = ~Q[19] /*30593*/;
assign _40204_ = _40205_ & D[55] /*30592*/;
assign _40207_ = _39416_ & _40204_ /*30587*/;
assign _40208_ = _39416_ ^ _40204_ /*30590*/;
assign _40209_ = _40200_ & _40208_ /*30588*/;
assign _39864_ = _40200_ ^ _40208_ /*30589*/;
assign _40206_ = _40207_ | _40209_ /*30586*/;
assign _40211_ = ~Q[19] /*30585*/;
assign _40210_ = _40211_ & D[56] /*30584*/;
assign _40213_ = _39417_ & _40210_ /*30579*/;
assign _40214_ = _39417_ ^ _40210_ /*30582*/;
assign _40215_ = _40206_ & _40214_ /*30580*/;
assign _39865_ = _40206_ ^ _40214_ /*30581*/;
assign _40212_ = _40213_ | _40215_ /*30578*/;
assign _40217_ = ~Q[19] /*30577*/;
assign _40216_ = _40217_ & D[57] /*30576*/;
assign _40219_ = _39418_ & _40216_ /*30571*/;
assign _40220_ = _39418_ ^ _40216_ /*30574*/;
assign _40221_ = _40212_ & _40220_ /*30572*/;
assign _39866_ = _40212_ ^ _40220_ /*30573*/;
assign _40218_ = _40219_ | _40221_ /*30570*/;
assign _40223_ = ~Q[19] /*30569*/;
assign _40222_ = _40223_ & D[58] /*30568*/;
assign _40225_ = _39419_ & _40222_ /*30563*/;
assign _40226_ = _39419_ ^ _40222_ /*30566*/;
assign _40227_ = _40218_ & _40226_ /*30564*/;
assign _39867_ = _40218_ ^ _40226_ /*30565*/;
assign _40224_ = _40225_ | _40227_ /*30562*/;
assign _40229_ = ~Q[19] /*30561*/;
assign _40228_ = _40229_ & D[59] /*30560*/;
assign _40231_ = _39420_ & _40228_ /*30555*/;
assign _40232_ = _39420_ ^ _40228_ /*30558*/;
assign _40233_ = _40224_ & _40232_ /*30556*/;
assign _39868_ = _40224_ ^ _40232_ /*30557*/;
assign _40230_ = _40231_ | _40233_ /*30554*/;
assign _40235_ = ~Q[19] /*30553*/;
assign _40234_ = _40235_ & D[60] /*30552*/;
assign _40237_ = _39421_ & _40234_ /*30547*/;
assign _40238_ = _39421_ ^ _40234_ /*30550*/;
assign _40239_ = _40230_ & _40238_ /*30548*/;
assign _39869_ = _40230_ ^ _40238_ /*30549*/;
assign _40236_ = _40237_ | _40239_ /*30546*/;
assign _40241_ = ~Q[19] /*30545*/;
assign _40240_ = _40241_ & D[61] /*30544*/;
assign _40243_ = _39422_ & _40240_ /*30539*/;
assign _40244_ = _39422_ ^ _40240_ /*30542*/;
assign _40245_ = _40236_ & _40244_ /*30540*/;
assign _39870_ = _40236_ ^ _40244_ /*30541*/;
assign _40242_ = _40243_ | _40245_ /*30538*/;
assign _40247_ = ~Q[19] /*30537*/;
assign _40246_ = _40247_ & D[62] /*30536*/;
assign _40249_ = _39423_ & _40246_ /*30531*/;
assign _40250_ = _39423_ ^ _40246_ /*30534*/;
assign _40251_ = _40242_ & _40250_ /*30532*/;
assign _39871_ = _40242_ ^ _40250_ /*30533*/;
assign _40248_ = _40249_ | _40251_ /*30530*/;
assign _40253_ = ~Q[19] /*30529*/;
assign _40252_ = _40253_ & zeroWire /*30528*/;
assign _40254_ = _39424_ ^ _40252_ /*30526*/;
assign _39872_ = _40254_ ^ _40248_ /*30525*/;
assign _40325_ = ~D[0] /*30271*/;
assign _40322_ = R_0[18] & _40325_ /*30267*/;
assign _40323_ = R_0[18] ^ _40325_ /*30270*/;
assign _40324_ = oneWire & _40323_ /*30268*/;
assign _40257_ = oneWire ^ _40323_ /*30269*/;
assign _40321_ = _40322_ | _40324_ /*30266*/;
assign _40330_ = ~D[1] /*30265*/;
assign _40327_ = _39809_ & _40330_ /*30261*/;
assign _40328_ = _39809_ ^ _40330_ /*30264*/;
assign _40329_ = _40321_ & _40328_ /*30262*/;
assign _40258_ = _40321_ ^ _40328_ /*30263*/;
assign _40326_ = _40327_ | _40329_ /*30260*/;
assign _40335_ = ~D[2] /*30259*/;
assign _40332_ = _39810_ & _40335_ /*30255*/;
assign _40333_ = _39810_ ^ _40335_ /*30258*/;
assign _40334_ = _40326_ & _40333_ /*30256*/;
assign _40259_ = _40326_ ^ _40333_ /*30257*/;
assign _40331_ = _40332_ | _40334_ /*30254*/;
assign _40340_ = ~D[3] /*30253*/;
assign _40337_ = _39811_ & _40340_ /*30249*/;
assign _40338_ = _39811_ ^ _40340_ /*30252*/;
assign _40339_ = _40331_ & _40338_ /*30250*/;
assign _40260_ = _40331_ ^ _40338_ /*30251*/;
assign _40336_ = _40337_ | _40339_ /*30248*/;
assign _40345_ = ~D[4] /*30247*/;
assign _40342_ = _39812_ & _40345_ /*30243*/;
assign _40343_ = _39812_ ^ _40345_ /*30246*/;
assign _40344_ = _40336_ & _40343_ /*30244*/;
assign _40261_ = _40336_ ^ _40343_ /*30245*/;
assign _40341_ = _40342_ | _40344_ /*30242*/;
assign _40350_ = ~D[5] /*30241*/;
assign _40347_ = _39813_ & _40350_ /*30237*/;
assign _40348_ = _39813_ ^ _40350_ /*30240*/;
assign _40349_ = _40341_ & _40348_ /*30238*/;
assign _40262_ = _40341_ ^ _40348_ /*30239*/;
assign _40346_ = _40347_ | _40349_ /*30236*/;
assign _40355_ = ~D[6] /*30235*/;
assign _40352_ = _39814_ & _40355_ /*30231*/;
assign _40353_ = _39814_ ^ _40355_ /*30234*/;
assign _40354_ = _40346_ & _40353_ /*30232*/;
assign _40263_ = _40346_ ^ _40353_ /*30233*/;
assign _40351_ = _40352_ | _40354_ /*30230*/;
assign _40360_ = ~D[7] /*30229*/;
assign _40357_ = _39815_ & _40360_ /*30225*/;
assign _40358_ = _39815_ ^ _40360_ /*30228*/;
assign _40359_ = _40351_ & _40358_ /*30226*/;
assign _40264_ = _40351_ ^ _40358_ /*30227*/;
assign _40356_ = _40357_ | _40359_ /*30224*/;
assign _40365_ = ~D[8] /*30223*/;
assign _40362_ = _39816_ & _40365_ /*30219*/;
assign _40363_ = _39816_ ^ _40365_ /*30222*/;
assign _40364_ = _40356_ & _40363_ /*30220*/;
assign _40265_ = _40356_ ^ _40363_ /*30221*/;
assign _40361_ = _40362_ | _40364_ /*30218*/;
assign _40370_ = ~D[9] /*30217*/;
assign _40367_ = _39817_ & _40370_ /*30213*/;
assign _40368_ = _39817_ ^ _40370_ /*30216*/;
assign _40369_ = _40361_ & _40368_ /*30214*/;
assign _40266_ = _40361_ ^ _40368_ /*30215*/;
assign _40366_ = _40367_ | _40369_ /*30212*/;
assign _40375_ = ~D[10] /*30211*/;
assign _40372_ = _39818_ & _40375_ /*30207*/;
assign _40373_ = _39818_ ^ _40375_ /*30210*/;
assign _40374_ = _40366_ & _40373_ /*30208*/;
assign _40267_ = _40366_ ^ _40373_ /*30209*/;
assign _40371_ = _40372_ | _40374_ /*30206*/;
assign _40380_ = ~D[11] /*30205*/;
assign _40377_ = _39819_ & _40380_ /*30201*/;
assign _40378_ = _39819_ ^ _40380_ /*30204*/;
assign _40379_ = _40371_ & _40378_ /*30202*/;
assign _40268_ = _40371_ ^ _40378_ /*30203*/;
assign _40376_ = _40377_ | _40379_ /*30200*/;
assign _40385_ = ~D[12] /*30199*/;
assign _40382_ = _39820_ & _40385_ /*30195*/;
assign _40383_ = _39820_ ^ _40385_ /*30198*/;
assign _40384_ = _40376_ & _40383_ /*30196*/;
assign _40269_ = _40376_ ^ _40383_ /*30197*/;
assign _40381_ = _40382_ | _40384_ /*30194*/;
assign _40390_ = ~D[13] /*30193*/;
assign _40387_ = _39821_ & _40390_ /*30189*/;
assign _40388_ = _39821_ ^ _40390_ /*30192*/;
assign _40389_ = _40381_ & _40388_ /*30190*/;
assign _40270_ = _40381_ ^ _40388_ /*30191*/;
assign _40386_ = _40387_ | _40389_ /*30188*/;
assign _40395_ = ~D[14] /*30187*/;
assign _40392_ = _39822_ & _40395_ /*30183*/;
assign _40393_ = _39822_ ^ _40395_ /*30186*/;
assign _40394_ = _40386_ & _40393_ /*30184*/;
assign _40271_ = _40386_ ^ _40393_ /*30185*/;
assign _40391_ = _40392_ | _40394_ /*30182*/;
assign _40400_ = ~D[15] /*30181*/;
assign _40397_ = _39823_ & _40400_ /*30177*/;
assign _40398_ = _39823_ ^ _40400_ /*30180*/;
assign _40399_ = _40391_ & _40398_ /*30178*/;
assign _40272_ = _40391_ ^ _40398_ /*30179*/;
assign _40396_ = _40397_ | _40399_ /*30176*/;
assign _40405_ = ~D[16] /*30175*/;
assign _40402_ = _39824_ & _40405_ /*30171*/;
assign _40403_ = _39824_ ^ _40405_ /*30174*/;
assign _40404_ = _40396_ & _40403_ /*30172*/;
assign _40273_ = _40396_ ^ _40403_ /*30173*/;
assign _40401_ = _40402_ | _40404_ /*30170*/;
assign _40410_ = ~D[17] /*30169*/;
assign _40407_ = _39825_ & _40410_ /*30165*/;
assign _40408_ = _39825_ ^ _40410_ /*30168*/;
assign _40409_ = _40401_ & _40408_ /*30166*/;
assign _40274_ = _40401_ ^ _40408_ /*30167*/;
assign _40406_ = _40407_ | _40409_ /*30164*/;
assign _40415_ = ~D[18] /*30163*/;
assign _40412_ = _39826_ & _40415_ /*30159*/;
assign _40413_ = _39826_ ^ _40415_ /*30162*/;
assign _40414_ = _40406_ & _40413_ /*30160*/;
assign _40275_ = _40406_ ^ _40413_ /*30161*/;
assign _40411_ = _40412_ | _40414_ /*30158*/;
assign _40420_ = ~D[19] /*30157*/;
assign _40417_ = _39827_ & _40420_ /*30153*/;
assign _40418_ = _39827_ ^ _40420_ /*30156*/;
assign _40419_ = _40411_ & _40418_ /*30154*/;
assign _40276_ = _40411_ ^ _40418_ /*30155*/;
assign _40416_ = _40417_ | _40419_ /*30152*/;
assign _40425_ = ~D[20] /*30151*/;
assign _40422_ = _39828_ & _40425_ /*30147*/;
assign _40423_ = _39828_ ^ _40425_ /*30150*/;
assign _40424_ = _40416_ & _40423_ /*30148*/;
assign _40277_ = _40416_ ^ _40423_ /*30149*/;
assign _40421_ = _40422_ | _40424_ /*30146*/;
assign _40430_ = ~D[21] /*30145*/;
assign _40427_ = _39829_ & _40430_ /*30141*/;
assign _40428_ = _39829_ ^ _40430_ /*30144*/;
assign _40429_ = _40421_ & _40428_ /*30142*/;
assign _40278_ = _40421_ ^ _40428_ /*30143*/;
assign _40426_ = _40427_ | _40429_ /*30140*/;
assign _40435_ = ~D[22] /*30139*/;
assign _40432_ = _39830_ & _40435_ /*30135*/;
assign _40433_ = _39830_ ^ _40435_ /*30138*/;
assign _40434_ = _40426_ & _40433_ /*30136*/;
assign _40279_ = _40426_ ^ _40433_ /*30137*/;
assign _40431_ = _40432_ | _40434_ /*30134*/;
assign _40440_ = ~D[23] /*30133*/;
assign _40437_ = _39831_ & _40440_ /*30129*/;
assign _40438_ = _39831_ ^ _40440_ /*30132*/;
assign _40439_ = _40431_ & _40438_ /*30130*/;
assign _40280_ = _40431_ ^ _40438_ /*30131*/;
assign _40436_ = _40437_ | _40439_ /*30128*/;
assign _40445_ = ~D[24] /*30127*/;
assign _40442_ = _39832_ & _40445_ /*30123*/;
assign _40443_ = _39832_ ^ _40445_ /*30126*/;
assign _40444_ = _40436_ & _40443_ /*30124*/;
assign _40281_ = _40436_ ^ _40443_ /*30125*/;
assign _40441_ = _40442_ | _40444_ /*30122*/;
assign _40450_ = ~D[25] /*30121*/;
assign _40447_ = _39833_ & _40450_ /*30117*/;
assign _40448_ = _39833_ ^ _40450_ /*30120*/;
assign _40449_ = _40441_ & _40448_ /*30118*/;
assign _40282_ = _40441_ ^ _40448_ /*30119*/;
assign _40446_ = _40447_ | _40449_ /*30116*/;
assign _40455_ = ~D[26] /*30115*/;
assign _40452_ = _39834_ & _40455_ /*30111*/;
assign _40453_ = _39834_ ^ _40455_ /*30114*/;
assign _40454_ = _40446_ & _40453_ /*30112*/;
assign _40283_ = _40446_ ^ _40453_ /*30113*/;
assign _40451_ = _40452_ | _40454_ /*30110*/;
assign _40460_ = ~D[27] /*30109*/;
assign _40457_ = _39835_ & _40460_ /*30105*/;
assign _40458_ = _39835_ ^ _40460_ /*30108*/;
assign _40459_ = _40451_ & _40458_ /*30106*/;
assign _40284_ = _40451_ ^ _40458_ /*30107*/;
assign _40456_ = _40457_ | _40459_ /*30104*/;
assign _40465_ = ~D[28] /*30103*/;
assign _40462_ = _39836_ & _40465_ /*30099*/;
assign _40463_ = _39836_ ^ _40465_ /*30102*/;
assign _40464_ = _40456_ & _40463_ /*30100*/;
assign _40285_ = _40456_ ^ _40463_ /*30101*/;
assign _40461_ = _40462_ | _40464_ /*30098*/;
assign _40470_ = ~D[29] /*30097*/;
assign _40467_ = _39837_ & _40470_ /*30093*/;
assign _40468_ = _39837_ ^ _40470_ /*30096*/;
assign _40469_ = _40461_ & _40468_ /*30094*/;
assign _40286_ = _40461_ ^ _40468_ /*30095*/;
assign _40466_ = _40467_ | _40469_ /*30092*/;
assign _40475_ = ~D[30] /*30091*/;
assign _40472_ = _39838_ & _40475_ /*30087*/;
assign _40473_ = _39838_ ^ _40475_ /*30090*/;
assign _40474_ = _40466_ & _40473_ /*30088*/;
assign _40287_ = _40466_ ^ _40473_ /*30089*/;
assign _40471_ = _40472_ | _40474_ /*30086*/;
assign _40480_ = ~D[31] /*30085*/;
assign _40477_ = _39839_ & _40480_ /*30081*/;
assign _40478_ = _39839_ ^ _40480_ /*30084*/;
assign _40479_ = _40471_ & _40478_ /*30082*/;
assign _40288_ = _40471_ ^ _40478_ /*30083*/;
assign _40476_ = _40477_ | _40479_ /*30080*/;
assign _40485_ = ~D[32] /*30079*/;
assign _40482_ = _39840_ & _40485_ /*30075*/;
assign _40483_ = _39840_ ^ _40485_ /*30078*/;
assign _40484_ = _40476_ & _40483_ /*30076*/;
assign _40289_ = _40476_ ^ _40483_ /*30077*/;
assign _40481_ = _40482_ | _40484_ /*30074*/;
assign _40490_ = ~D[33] /*30073*/;
assign _40487_ = _39841_ & _40490_ /*30069*/;
assign _40488_ = _39841_ ^ _40490_ /*30072*/;
assign _40489_ = _40481_ & _40488_ /*30070*/;
assign _40290_ = _40481_ ^ _40488_ /*30071*/;
assign _40486_ = _40487_ | _40489_ /*30068*/;
assign _40495_ = ~D[34] /*30067*/;
assign _40492_ = _39842_ & _40495_ /*30063*/;
assign _40493_ = _39842_ ^ _40495_ /*30066*/;
assign _40494_ = _40486_ & _40493_ /*30064*/;
assign _40291_ = _40486_ ^ _40493_ /*30065*/;
assign _40491_ = _40492_ | _40494_ /*30062*/;
assign _40500_ = ~D[35] /*30061*/;
assign _40497_ = _39843_ & _40500_ /*30057*/;
assign _40498_ = _39843_ ^ _40500_ /*30060*/;
assign _40499_ = _40491_ & _40498_ /*30058*/;
assign _40292_ = _40491_ ^ _40498_ /*30059*/;
assign _40496_ = _40497_ | _40499_ /*30056*/;
assign _40505_ = ~D[36] /*30055*/;
assign _40502_ = _39844_ & _40505_ /*30051*/;
assign _40503_ = _39844_ ^ _40505_ /*30054*/;
assign _40504_ = _40496_ & _40503_ /*30052*/;
assign _40293_ = _40496_ ^ _40503_ /*30053*/;
assign _40501_ = _40502_ | _40504_ /*30050*/;
assign _40510_ = ~D[37] /*30049*/;
assign _40507_ = _39845_ & _40510_ /*30045*/;
assign _40508_ = _39845_ ^ _40510_ /*30048*/;
assign _40509_ = _40501_ & _40508_ /*30046*/;
assign _40294_ = _40501_ ^ _40508_ /*30047*/;
assign _40506_ = _40507_ | _40509_ /*30044*/;
assign _40515_ = ~D[38] /*30043*/;
assign _40512_ = _39846_ & _40515_ /*30039*/;
assign _40513_ = _39846_ ^ _40515_ /*30042*/;
assign _40514_ = _40506_ & _40513_ /*30040*/;
assign _40295_ = _40506_ ^ _40513_ /*30041*/;
assign _40511_ = _40512_ | _40514_ /*30038*/;
assign _40520_ = ~D[39] /*30037*/;
assign _40517_ = _39847_ & _40520_ /*30033*/;
assign _40518_ = _39847_ ^ _40520_ /*30036*/;
assign _40519_ = _40511_ & _40518_ /*30034*/;
assign _40296_ = _40511_ ^ _40518_ /*30035*/;
assign _40516_ = _40517_ | _40519_ /*30032*/;
assign _40525_ = ~D[40] /*30031*/;
assign _40522_ = _39848_ & _40525_ /*30027*/;
assign _40523_ = _39848_ ^ _40525_ /*30030*/;
assign _40524_ = _40516_ & _40523_ /*30028*/;
assign _40297_ = _40516_ ^ _40523_ /*30029*/;
assign _40521_ = _40522_ | _40524_ /*30026*/;
assign _40530_ = ~D[41] /*30025*/;
assign _40527_ = _39849_ & _40530_ /*30021*/;
assign _40528_ = _39849_ ^ _40530_ /*30024*/;
assign _40529_ = _40521_ & _40528_ /*30022*/;
assign _40298_ = _40521_ ^ _40528_ /*30023*/;
assign _40526_ = _40527_ | _40529_ /*30020*/;
assign _40535_ = ~D[42] /*30019*/;
assign _40532_ = _39850_ & _40535_ /*30015*/;
assign _40533_ = _39850_ ^ _40535_ /*30018*/;
assign _40534_ = _40526_ & _40533_ /*30016*/;
assign _40299_ = _40526_ ^ _40533_ /*30017*/;
assign _40531_ = _40532_ | _40534_ /*30014*/;
assign _40540_ = ~D[43] /*30013*/;
assign _40537_ = _39851_ & _40540_ /*30009*/;
assign _40538_ = _39851_ ^ _40540_ /*30012*/;
assign _40539_ = _40531_ & _40538_ /*30010*/;
assign _40300_ = _40531_ ^ _40538_ /*30011*/;
assign _40536_ = _40537_ | _40539_ /*30008*/;
assign _40545_ = ~D[44] /*30007*/;
assign _40542_ = _39852_ & _40545_ /*30003*/;
assign _40543_ = _39852_ ^ _40545_ /*30006*/;
assign _40544_ = _40536_ & _40543_ /*30004*/;
assign _40301_ = _40536_ ^ _40543_ /*30005*/;
assign _40541_ = _40542_ | _40544_ /*30002*/;
assign _40550_ = ~D[45] /*30001*/;
assign _40547_ = _39853_ & _40550_ /*29997*/;
assign _40548_ = _39853_ ^ _40550_ /*30000*/;
assign _40549_ = _40541_ & _40548_ /*29998*/;
assign _40302_ = _40541_ ^ _40548_ /*29999*/;
assign _40546_ = _40547_ | _40549_ /*29996*/;
assign _40555_ = ~D[46] /*29995*/;
assign _40552_ = _39854_ & _40555_ /*29991*/;
assign _40553_ = _39854_ ^ _40555_ /*29994*/;
assign _40554_ = _40546_ & _40553_ /*29992*/;
assign _40303_ = _40546_ ^ _40553_ /*29993*/;
assign _40551_ = _40552_ | _40554_ /*29990*/;
assign _40560_ = ~D[47] /*29989*/;
assign _40557_ = _39855_ & _40560_ /*29985*/;
assign _40558_ = _39855_ ^ _40560_ /*29988*/;
assign _40559_ = _40551_ & _40558_ /*29986*/;
assign _40304_ = _40551_ ^ _40558_ /*29987*/;
assign _40556_ = _40557_ | _40559_ /*29984*/;
assign _40565_ = ~D[48] /*29983*/;
assign _40562_ = _39856_ & _40565_ /*29979*/;
assign _40563_ = _39856_ ^ _40565_ /*29982*/;
assign _40564_ = _40556_ & _40563_ /*29980*/;
assign _40305_ = _40556_ ^ _40563_ /*29981*/;
assign _40561_ = _40562_ | _40564_ /*29978*/;
assign _40570_ = ~D[49] /*29977*/;
assign _40567_ = _39857_ & _40570_ /*29973*/;
assign _40568_ = _39857_ ^ _40570_ /*29976*/;
assign _40569_ = _40561_ & _40568_ /*29974*/;
assign _40306_ = _40561_ ^ _40568_ /*29975*/;
assign _40566_ = _40567_ | _40569_ /*29972*/;
assign _40575_ = ~D[50] /*29971*/;
assign _40572_ = _39858_ & _40575_ /*29967*/;
assign _40573_ = _39858_ ^ _40575_ /*29970*/;
assign _40574_ = _40566_ & _40573_ /*29968*/;
assign _40307_ = _40566_ ^ _40573_ /*29969*/;
assign _40571_ = _40572_ | _40574_ /*29966*/;
assign _40580_ = ~D[51] /*29965*/;
assign _40577_ = _39859_ & _40580_ /*29961*/;
assign _40578_ = _39859_ ^ _40580_ /*29964*/;
assign _40579_ = _40571_ & _40578_ /*29962*/;
assign _40308_ = _40571_ ^ _40578_ /*29963*/;
assign _40576_ = _40577_ | _40579_ /*29960*/;
assign _40585_ = ~D[52] /*29959*/;
assign _40582_ = _39860_ & _40585_ /*29955*/;
assign _40583_ = _39860_ ^ _40585_ /*29958*/;
assign _40584_ = _40576_ & _40583_ /*29956*/;
assign _40309_ = _40576_ ^ _40583_ /*29957*/;
assign _40581_ = _40582_ | _40584_ /*29954*/;
assign _40590_ = ~D[53] /*29953*/;
assign _40587_ = _39861_ & _40590_ /*29949*/;
assign _40588_ = _39861_ ^ _40590_ /*29952*/;
assign _40589_ = _40581_ & _40588_ /*29950*/;
assign _40310_ = _40581_ ^ _40588_ /*29951*/;
assign _40586_ = _40587_ | _40589_ /*29948*/;
assign _40595_ = ~D[54] /*29947*/;
assign _40592_ = _39862_ & _40595_ /*29943*/;
assign _40593_ = _39862_ ^ _40595_ /*29946*/;
assign _40594_ = _40586_ & _40593_ /*29944*/;
assign _40311_ = _40586_ ^ _40593_ /*29945*/;
assign _40591_ = _40592_ | _40594_ /*29942*/;
assign _40600_ = ~D[55] /*29941*/;
assign _40597_ = _39863_ & _40600_ /*29937*/;
assign _40598_ = _39863_ ^ _40600_ /*29940*/;
assign _40599_ = _40591_ & _40598_ /*29938*/;
assign _40312_ = _40591_ ^ _40598_ /*29939*/;
assign _40596_ = _40597_ | _40599_ /*29936*/;
assign _40605_ = ~D[56] /*29935*/;
assign _40602_ = _39864_ & _40605_ /*29931*/;
assign _40603_ = _39864_ ^ _40605_ /*29934*/;
assign _40604_ = _40596_ & _40603_ /*29932*/;
assign _40313_ = _40596_ ^ _40603_ /*29933*/;
assign _40601_ = _40602_ | _40604_ /*29930*/;
assign _40610_ = ~D[57] /*29929*/;
assign _40607_ = _39865_ & _40610_ /*29925*/;
assign _40608_ = _39865_ ^ _40610_ /*29928*/;
assign _40609_ = _40601_ & _40608_ /*29926*/;
assign _40314_ = _40601_ ^ _40608_ /*29927*/;
assign _40606_ = _40607_ | _40609_ /*29924*/;
assign _40615_ = ~D[58] /*29923*/;
assign _40612_ = _39866_ & _40615_ /*29919*/;
assign _40613_ = _39866_ ^ _40615_ /*29922*/;
assign _40614_ = _40606_ & _40613_ /*29920*/;
assign _40315_ = _40606_ ^ _40613_ /*29921*/;
assign _40611_ = _40612_ | _40614_ /*29918*/;
assign _40620_ = ~D[59] /*29917*/;
assign _40617_ = _39867_ & _40620_ /*29913*/;
assign _40618_ = _39867_ ^ _40620_ /*29916*/;
assign _40619_ = _40611_ & _40618_ /*29914*/;
assign _40316_ = _40611_ ^ _40618_ /*29915*/;
assign _40616_ = _40617_ | _40619_ /*29912*/;
assign _40625_ = ~D[60] /*29911*/;
assign _40622_ = _39868_ & _40625_ /*29907*/;
assign _40623_ = _39868_ ^ _40625_ /*29910*/;
assign _40624_ = _40616_ & _40623_ /*29908*/;
assign _40317_ = _40616_ ^ _40623_ /*29909*/;
assign _40621_ = _40622_ | _40624_ /*29906*/;
assign _40630_ = ~D[61] /*29905*/;
assign _40627_ = _39869_ & _40630_ /*29901*/;
assign _40628_ = _39869_ ^ _40630_ /*29904*/;
assign _40629_ = _40621_ & _40628_ /*29902*/;
assign _40318_ = _40621_ ^ _40628_ /*29903*/;
assign _40626_ = _40627_ | _40629_ /*29900*/;
assign _40635_ = ~D[62] /*29899*/;
assign _40632_ = _39870_ & _40635_ /*29895*/;
assign _40633_ = _39870_ ^ _40635_ /*29898*/;
assign _40634_ = _40626_ & _40633_ /*29896*/;
assign _40319_ = _40626_ ^ _40633_ /*29897*/;
assign _40631_ = _40632_ | _40634_ /*29894*/;
assign _40636_ = _39871_ & oneWire /*29889*/;
assign _40637_ = _39871_ ^ oneWire /*29892*/;
assign _40638_ = _40631_ & _40637_ /*29890*/;
assign _40320_ = _40631_ ^ _40637_ /*29891*/;
assign Q[18] = _40636_ | _40638_ /*29888*/;
assign _40771_ = ~Q[18] /*29503*/;
assign _40770_ = _40771_ & D[0] /*29502*/;
assign _40773_ = _40257_ & _40770_ /*29497*/;
assign _40774_ = _40257_ ^ _40770_ /*29500*/;
assign _40775_ = zeroWire & _40774_ /*29498*/;
assign _40705_ = zeroWire ^ _40774_ /*29499*/;
assign _40772_ = _40773_ | _40775_ /*29496*/;
assign _40777_ = ~Q[18] /*29495*/;
assign _40776_ = _40777_ & D[1] /*29494*/;
assign _40779_ = _40258_ & _40776_ /*29489*/;
assign _40780_ = _40258_ ^ _40776_ /*29492*/;
assign _40781_ = _40772_ & _40780_ /*29490*/;
assign _40706_ = _40772_ ^ _40780_ /*29491*/;
assign _40778_ = _40779_ | _40781_ /*29488*/;
assign _40783_ = ~Q[18] /*29487*/;
assign _40782_ = _40783_ & D[2] /*29486*/;
assign _40785_ = _40259_ & _40782_ /*29481*/;
assign _40786_ = _40259_ ^ _40782_ /*29484*/;
assign _40787_ = _40778_ & _40786_ /*29482*/;
assign _40707_ = _40778_ ^ _40786_ /*29483*/;
assign _40784_ = _40785_ | _40787_ /*29480*/;
assign _40789_ = ~Q[18] /*29479*/;
assign _40788_ = _40789_ & D[3] /*29478*/;
assign _40791_ = _40260_ & _40788_ /*29473*/;
assign _40792_ = _40260_ ^ _40788_ /*29476*/;
assign _40793_ = _40784_ & _40792_ /*29474*/;
assign _40708_ = _40784_ ^ _40792_ /*29475*/;
assign _40790_ = _40791_ | _40793_ /*29472*/;
assign _40795_ = ~Q[18] /*29471*/;
assign _40794_ = _40795_ & D[4] /*29470*/;
assign _40797_ = _40261_ & _40794_ /*29465*/;
assign _40798_ = _40261_ ^ _40794_ /*29468*/;
assign _40799_ = _40790_ & _40798_ /*29466*/;
assign _40709_ = _40790_ ^ _40798_ /*29467*/;
assign _40796_ = _40797_ | _40799_ /*29464*/;
assign _40801_ = ~Q[18] /*29463*/;
assign _40800_ = _40801_ & D[5] /*29462*/;
assign _40803_ = _40262_ & _40800_ /*29457*/;
assign _40804_ = _40262_ ^ _40800_ /*29460*/;
assign _40805_ = _40796_ & _40804_ /*29458*/;
assign _40710_ = _40796_ ^ _40804_ /*29459*/;
assign _40802_ = _40803_ | _40805_ /*29456*/;
assign _40807_ = ~Q[18] /*29455*/;
assign _40806_ = _40807_ & D[6] /*29454*/;
assign _40809_ = _40263_ & _40806_ /*29449*/;
assign _40810_ = _40263_ ^ _40806_ /*29452*/;
assign _40811_ = _40802_ & _40810_ /*29450*/;
assign _40711_ = _40802_ ^ _40810_ /*29451*/;
assign _40808_ = _40809_ | _40811_ /*29448*/;
assign _40813_ = ~Q[18] /*29447*/;
assign _40812_ = _40813_ & D[7] /*29446*/;
assign _40815_ = _40264_ & _40812_ /*29441*/;
assign _40816_ = _40264_ ^ _40812_ /*29444*/;
assign _40817_ = _40808_ & _40816_ /*29442*/;
assign _40712_ = _40808_ ^ _40816_ /*29443*/;
assign _40814_ = _40815_ | _40817_ /*29440*/;
assign _40819_ = ~Q[18] /*29439*/;
assign _40818_ = _40819_ & D[8] /*29438*/;
assign _40821_ = _40265_ & _40818_ /*29433*/;
assign _40822_ = _40265_ ^ _40818_ /*29436*/;
assign _40823_ = _40814_ & _40822_ /*29434*/;
assign _40713_ = _40814_ ^ _40822_ /*29435*/;
assign _40820_ = _40821_ | _40823_ /*29432*/;
assign _40825_ = ~Q[18] /*29431*/;
assign _40824_ = _40825_ & D[9] /*29430*/;
assign _40827_ = _40266_ & _40824_ /*29425*/;
assign _40828_ = _40266_ ^ _40824_ /*29428*/;
assign _40829_ = _40820_ & _40828_ /*29426*/;
assign _40714_ = _40820_ ^ _40828_ /*29427*/;
assign _40826_ = _40827_ | _40829_ /*29424*/;
assign _40831_ = ~Q[18] /*29423*/;
assign _40830_ = _40831_ & D[10] /*29422*/;
assign _40833_ = _40267_ & _40830_ /*29417*/;
assign _40834_ = _40267_ ^ _40830_ /*29420*/;
assign _40835_ = _40826_ & _40834_ /*29418*/;
assign _40715_ = _40826_ ^ _40834_ /*29419*/;
assign _40832_ = _40833_ | _40835_ /*29416*/;
assign _40837_ = ~Q[18] /*29415*/;
assign _40836_ = _40837_ & D[11] /*29414*/;
assign _40839_ = _40268_ & _40836_ /*29409*/;
assign _40840_ = _40268_ ^ _40836_ /*29412*/;
assign _40841_ = _40832_ & _40840_ /*29410*/;
assign _40716_ = _40832_ ^ _40840_ /*29411*/;
assign _40838_ = _40839_ | _40841_ /*29408*/;
assign _40843_ = ~Q[18] /*29407*/;
assign _40842_ = _40843_ & D[12] /*29406*/;
assign _40845_ = _40269_ & _40842_ /*29401*/;
assign _40846_ = _40269_ ^ _40842_ /*29404*/;
assign _40847_ = _40838_ & _40846_ /*29402*/;
assign _40717_ = _40838_ ^ _40846_ /*29403*/;
assign _40844_ = _40845_ | _40847_ /*29400*/;
assign _40849_ = ~Q[18] /*29399*/;
assign _40848_ = _40849_ & D[13] /*29398*/;
assign _40851_ = _40270_ & _40848_ /*29393*/;
assign _40852_ = _40270_ ^ _40848_ /*29396*/;
assign _40853_ = _40844_ & _40852_ /*29394*/;
assign _40718_ = _40844_ ^ _40852_ /*29395*/;
assign _40850_ = _40851_ | _40853_ /*29392*/;
assign _40855_ = ~Q[18] /*29391*/;
assign _40854_ = _40855_ & D[14] /*29390*/;
assign _40857_ = _40271_ & _40854_ /*29385*/;
assign _40858_ = _40271_ ^ _40854_ /*29388*/;
assign _40859_ = _40850_ & _40858_ /*29386*/;
assign _40719_ = _40850_ ^ _40858_ /*29387*/;
assign _40856_ = _40857_ | _40859_ /*29384*/;
assign _40861_ = ~Q[18] /*29383*/;
assign _40860_ = _40861_ & D[15] /*29382*/;
assign _40863_ = _40272_ & _40860_ /*29377*/;
assign _40864_ = _40272_ ^ _40860_ /*29380*/;
assign _40865_ = _40856_ & _40864_ /*29378*/;
assign _40720_ = _40856_ ^ _40864_ /*29379*/;
assign _40862_ = _40863_ | _40865_ /*29376*/;
assign _40867_ = ~Q[18] /*29375*/;
assign _40866_ = _40867_ & D[16] /*29374*/;
assign _40869_ = _40273_ & _40866_ /*29369*/;
assign _40870_ = _40273_ ^ _40866_ /*29372*/;
assign _40871_ = _40862_ & _40870_ /*29370*/;
assign _40721_ = _40862_ ^ _40870_ /*29371*/;
assign _40868_ = _40869_ | _40871_ /*29368*/;
assign _40873_ = ~Q[18] /*29367*/;
assign _40872_ = _40873_ & D[17] /*29366*/;
assign _40875_ = _40274_ & _40872_ /*29361*/;
assign _40876_ = _40274_ ^ _40872_ /*29364*/;
assign _40877_ = _40868_ & _40876_ /*29362*/;
assign _40722_ = _40868_ ^ _40876_ /*29363*/;
assign _40874_ = _40875_ | _40877_ /*29360*/;
assign _40879_ = ~Q[18] /*29359*/;
assign _40878_ = _40879_ & D[18] /*29358*/;
assign _40881_ = _40275_ & _40878_ /*29353*/;
assign _40882_ = _40275_ ^ _40878_ /*29356*/;
assign _40883_ = _40874_ & _40882_ /*29354*/;
assign _40723_ = _40874_ ^ _40882_ /*29355*/;
assign _40880_ = _40881_ | _40883_ /*29352*/;
assign _40885_ = ~Q[18] /*29351*/;
assign _40884_ = _40885_ & D[19] /*29350*/;
assign _40887_ = _40276_ & _40884_ /*29345*/;
assign _40888_ = _40276_ ^ _40884_ /*29348*/;
assign _40889_ = _40880_ & _40888_ /*29346*/;
assign _40724_ = _40880_ ^ _40888_ /*29347*/;
assign _40886_ = _40887_ | _40889_ /*29344*/;
assign _40891_ = ~Q[18] /*29343*/;
assign _40890_ = _40891_ & D[20] /*29342*/;
assign _40893_ = _40277_ & _40890_ /*29337*/;
assign _40894_ = _40277_ ^ _40890_ /*29340*/;
assign _40895_ = _40886_ & _40894_ /*29338*/;
assign _40725_ = _40886_ ^ _40894_ /*29339*/;
assign _40892_ = _40893_ | _40895_ /*29336*/;
assign _40897_ = ~Q[18] /*29335*/;
assign _40896_ = _40897_ & D[21] /*29334*/;
assign _40899_ = _40278_ & _40896_ /*29329*/;
assign _40900_ = _40278_ ^ _40896_ /*29332*/;
assign _40901_ = _40892_ & _40900_ /*29330*/;
assign _40726_ = _40892_ ^ _40900_ /*29331*/;
assign _40898_ = _40899_ | _40901_ /*29328*/;
assign _40903_ = ~Q[18] /*29327*/;
assign _40902_ = _40903_ & D[22] /*29326*/;
assign _40905_ = _40279_ & _40902_ /*29321*/;
assign _40906_ = _40279_ ^ _40902_ /*29324*/;
assign _40907_ = _40898_ & _40906_ /*29322*/;
assign _40727_ = _40898_ ^ _40906_ /*29323*/;
assign _40904_ = _40905_ | _40907_ /*29320*/;
assign _40909_ = ~Q[18] /*29319*/;
assign _40908_ = _40909_ & D[23] /*29318*/;
assign _40911_ = _40280_ & _40908_ /*29313*/;
assign _40912_ = _40280_ ^ _40908_ /*29316*/;
assign _40913_ = _40904_ & _40912_ /*29314*/;
assign _40728_ = _40904_ ^ _40912_ /*29315*/;
assign _40910_ = _40911_ | _40913_ /*29312*/;
assign _40915_ = ~Q[18] /*29311*/;
assign _40914_ = _40915_ & D[24] /*29310*/;
assign _40917_ = _40281_ & _40914_ /*29305*/;
assign _40918_ = _40281_ ^ _40914_ /*29308*/;
assign _40919_ = _40910_ & _40918_ /*29306*/;
assign _40729_ = _40910_ ^ _40918_ /*29307*/;
assign _40916_ = _40917_ | _40919_ /*29304*/;
assign _40921_ = ~Q[18] /*29303*/;
assign _40920_ = _40921_ & D[25] /*29302*/;
assign _40923_ = _40282_ & _40920_ /*29297*/;
assign _40924_ = _40282_ ^ _40920_ /*29300*/;
assign _40925_ = _40916_ & _40924_ /*29298*/;
assign _40730_ = _40916_ ^ _40924_ /*29299*/;
assign _40922_ = _40923_ | _40925_ /*29296*/;
assign _40927_ = ~Q[18] /*29295*/;
assign _40926_ = _40927_ & D[26] /*29294*/;
assign _40929_ = _40283_ & _40926_ /*29289*/;
assign _40930_ = _40283_ ^ _40926_ /*29292*/;
assign _40931_ = _40922_ & _40930_ /*29290*/;
assign _40731_ = _40922_ ^ _40930_ /*29291*/;
assign _40928_ = _40929_ | _40931_ /*29288*/;
assign _40933_ = ~Q[18] /*29287*/;
assign _40932_ = _40933_ & D[27] /*29286*/;
assign _40935_ = _40284_ & _40932_ /*29281*/;
assign _40936_ = _40284_ ^ _40932_ /*29284*/;
assign _40937_ = _40928_ & _40936_ /*29282*/;
assign _40732_ = _40928_ ^ _40936_ /*29283*/;
assign _40934_ = _40935_ | _40937_ /*29280*/;
assign _40939_ = ~Q[18] /*29279*/;
assign _40938_ = _40939_ & D[28] /*29278*/;
assign _40941_ = _40285_ & _40938_ /*29273*/;
assign _40942_ = _40285_ ^ _40938_ /*29276*/;
assign _40943_ = _40934_ & _40942_ /*29274*/;
assign _40733_ = _40934_ ^ _40942_ /*29275*/;
assign _40940_ = _40941_ | _40943_ /*29272*/;
assign _40945_ = ~Q[18] /*29271*/;
assign _40944_ = _40945_ & D[29] /*29270*/;
assign _40947_ = _40286_ & _40944_ /*29265*/;
assign _40948_ = _40286_ ^ _40944_ /*29268*/;
assign _40949_ = _40940_ & _40948_ /*29266*/;
assign _40734_ = _40940_ ^ _40948_ /*29267*/;
assign _40946_ = _40947_ | _40949_ /*29264*/;
assign _40951_ = ~Q[18] /*29263*/;
assign _40950_ = _40951_ & D[30] /*29262*/;
assign _40953_ = _40287_ & _40950_ /*29257*/;
assign _40954_ = _40287_ ^ _40950_ /*29260*/;
assign _40955_ = _40946_ & _40954_ /*29258*/;
assign _40735_ = _40946_ ^ _40954_ /*29259*/;
assign _40952_ = _40953_ | _40955_ /*29256*/;
assign _40957_ = ~Q[18] /*29255*/;
assign _40956_ = _40957_ & D[31] /*29254*/;
assign _40959_ = _40288_ & _40956_ /*29249*/;
assign _40960_ = _40288_ ^ _40956_ /*29252*/;
assign _40961_ = _40952_ & _40960_ /*29250*/;
assign _40736_ = _40952_ ^ _40960_ /*29251*/;
assign _40958_ = _40959_ | _40961_ /*29248*/;
assign _40963_ = ~Q[18] /*29247*/;
assign _40962_ = _40963_ & D[32] /*29246*/;
assign _40965_ = _40289_ & _40962_ /*29241*/;
assign _40966_ = _40289_ ^ _40962_ /*29244*/;
assign _40967_ = _40958_ & _40966_ /*29242*/;
assign _40737_ = _40958_ ^ _40966_ /*29243*/;
assign _40964_ = _40965_ | _40967_ /*29240*/;
assign _40969_ = ~Q[18] /*29239*/;
assign _40968_ = _40969_ & D[33] /*29238*/;
assign _40971_ = _40290_ & _40968_ /*29233*/;
assign _40972_ = _40290_ ^ _40968_ /*29236*/;
assign _40973_ = _40964_ & _40972_ /*29234*/;
assign _40738_ = _40964_ ^ _40972_ /*29235*/;
assign _40970_ = _40971_ | _40973_ /*29232*/;
assign _40975_ = ~Q[18] /*29231*/;
assign _40974_ = _40975_ & D[34] /*29230*/;
assign _40977_ = _40291_ & _40974_ /*29225*/;
assign _40978_ = _40291_ ^ _40974_ /*29228*/;
assign _40979_ = _40970_ & _40978_ /*29226*/;
assign _40739_ = _40970_ ^ _40978_ /*29227*/;
assign _40976_ = _40977_ | _40979_ /*29224*/;
assign _40981_ = ~Q[18] /*29223*/;
assign _40980_ = _40981_ & D[35] /*29222*/;
assign _40983_ = _40292_ & _40980_ /*29217*/;
assign _40984_ = _40292_ ^ _40980_ /*29220*/;
assign _40985_ = _40976_ & _40984_ /*29218*/;
assign _40740_ = _40976_ ^ _40984_ /*29219*/;
assign _40982_ = _40983_ | _40985_ /*29216*/;
assign _40987_ = ~Q[18] /*29215*/;
assign _40986_ = _40987_ & D[36] /*29214*/;
assign _40989_ = _40293_ & _40986_ /*29209*/;
assign _40990_ = _40293_ ^ _40986_ /*29212*/;
assign _40991_ = _40982_ & _40990_ /*29210*/;
assign _40741_ = _40982_ ^ _40990_ /*29211*/;
assign _40988_ = _40989_ | _40991_ /*29208*/;
assign _40993_ = ~Q[18] /*29207*/;
assign _40992_ = _40993_ & D[37] /*29206*/;
assign _40995_ = _40294_ & _40992_ /*29201*/;
assign _40996_ = _40294_ ^ _40992_ /*29204*/;
assign _40997_ = _40988_ & _40996_ /*29202*/;
assign _40742_ = _40988_ ^ _40996_ /*29203*/;
assign _40994_ = _40995_ | _40997_ /*29200*/;
assign _40999_ = ~Q[18] /*29199*/;
assign _40998_ = _40999_ & D[38] /*29198*/;
assign _41001_ = _40295_ & _40998_ /*29193*/;
assign _41002_ = _40295_ ^ _40998_ /*29196*/;
assign _41003_ = _40994_ & _41002_ /*29194*/;
assign _40743_ = _40994_ ^ _41002_ /*29195*/;
assign _41000_ = _41001_ | _41003_ /*29192*/;
assign _41005_ = ~Q[18] /*29191*/;
assign _41004_ = _41005_ & D[39] /*29190*/;
assign _41007_ = _40296_ & _41004_ /*29185*/;
assign _41008_ = _40296_ ^ _41004_ /*29188*/;
assign _41009_ = _41000_ & _41008_ /*29186*/;
assign _40744_ = _41000_ ^ _41008_ /*29187*/;
assign _41006_ = _41007_ | _41009_ /*29184*/;
assign _41011_ = ~Q[18] /*29183*/;
assign _41010_ = _41011_ & D[40] /*29182*/;
assign _41013_ = _40297_ & _41010_ /*29177*/;
assign _41014_ = _40297_ ^ _41010_ /*29180*/;
assign _41015_ = _41006_ & _41014_ /*29178*/;
assign _40745_ = _41006_ ^ _41014_ /*29179*/;
assign _41012_ = _41013_ | _41015_ /*29176*/;
assign _41017_ = ~Q[18] /*29175*/;
assign _41016_ = _41017_ & D[41] /*29174*/;
assign _41019_ = _40298_ & _41016_ /*29169*/;
assign _41020_ = _40298_ ^ _41016_ /*29172*/;
assign _41021_ = _41012_ & _41020_ /*29170*/;
assign _40746_ = _41012_ ^ _41020_ /*29171*/;
assign _41018_ = _41019_ | _41021_ /*29168*/;
assign _41023_ = ~Q[18] /*29167*/;
assign _41022_ = _41023_ & D[42] /*29166*/;
assign _41025_ = _40299_ & _41022_ /*29161*/;
assign _41026_ = _40299_ ^ _41022_ /*29164*/;
assign _41027_ = _41018_ & _41026_ /*29162*/;
assign _40747_ = _41018_ ^ _41026_ /*29163*/;
assign _41024_ = _41025_ | _41027_ /*29160*/;
assign _41029_ = ~Q[18] /*29159*/;
assign _41028_ = _41029_ & D[43] /*29158*/;
assign _41031_ = _40300_ & _41028_ /*29153*/;
assign _41032_ = _40300_ ^ _41028_ /*29156*/;
assign _41033_ = _41024_ & _41032_ /*29154*/;
assign _40748_ = _41024_ ^ _41032_ /*29155*/;
assign _41030_ = _41031_ | _41033_ /*29152*/;
assign _41035_ = ~Q[18] /*29151*/;
assign _41034_ = _41035_ & D[44] /*29150*/;
assign _41037_ = _40301_ & _41034_ /*29145*/;
assign _41038_ = _40301_ ^ _41034_ /*29148*/;
assign _41039_ = _41030_ & _41038_ /*29146*/;
assign _40749_ = _41030_ ^ _41038_ /*29147*/;
assign _41036_ = _41037_ | _41039_ /*29144*/;
assign _41041_ = ~Q[18] /*29143*/;
assign _41040_ = _41041_ & D[45] /*29142*/;
assign _41043_ = _40302_ & _41040_ /*29137*/;
assign _41044_ = _40302_ ^ _41040_ /*29140*/;
assign _41045_ = _41036_ & _41044_ /*29138*/;
assign _40750_ = _41036_ ^ _41044_ /*29139*/;
assign _41042_ = _41043_ | _41045_ /*29136*/;
assign _41047_ = ~Q[18] /*29135*/;
assign _41046_ = _41047_ & D[46] /*29134*/;
assign _41049_ = _40303_ & _41046_ /*29129*/;
assign _41050_ = _40303_ ^ _41046_ /*29132*/;
assign _41051_ = _41042_ & _41050_ /*29130*/;
assign _40751_ = _41042_ ^ _41050_ /*29131*/;
assign _41048_ = _41049_ | _41051_ /*29128*/;
assign _41053_ = ~Q[18] /*29127*/;
assign _41052_ = _41053_ & D[47] /*29126*/;
assign _41055_ = _40304_ & _41052_ /*29121*/;
assign _41056_ = _40304_ ^ _41052_ /*29124*/;
assign _41057_ = _41048_ & _41056_ /*29122*/;
assign _40752_ = _41048_ ^ _41056_ /*29123*/;
assign _41054_ = _41055_ | _41057_ /*29120*/;
assign _41059_ = ~Q[18] /*29119*/;
assign _41058_ = _41059_ & D[48] /*29118*/;
assign _41061_ = _40305_ & _41058_ /*29113*/;
assign _41062_ = _40305_ ^ _41058_ /*29116*/;
assign _41063_ = _41054_ & _41062_ /*29114*/;
assign _40753_ = _41054_ ^ _41062_ /*29115*/;
assign _41060_ = _41061_ | _41063_ /*29112*/;
assign _41065_ = ~Q[18] /*29111*/;
assign _41064_ = _41065_ & D[49] /*29110*/;
assign _41067_ = _40306_ & _41064_ /*29105*/;
assign _41068_ = _40306_ ^ _41064_ /*29108*/;
assign _41069_ = _41060_ & _41068_ /*29106*/;
assign _40754_ = _41060_ ^ _41068_ /*29107*/;
assign _41066_ = _41067_ | _41069_ /*29104*/;
assign _41071_ = ~Q[18] /*29103*/;
assign _41070_ = _41071_ & D[50] /*29102*/;
assign _41073_ = _40307_ & _41070_ /*29097*/;
assign _41074_ = _40307_ ^ _41070_ /*29100*/;
assign _41075_ = _41066_ & _41074_ /*29098*/;
assign _40755_ = _41066_ ^ _41074_ /*29099*/;
assign _41072_ = _41073_ | _41075_ /*29096*/;
assign _41077_ = ~Q[18] /*29095*/;
assign _41076_ = _41077_ & D[51] /*29094*/;
assign _41079_ = _40308_ & _41076_ /*29089*/;
assign _41080_ = _40308_ ^ _41076_ /*29092*/;
assign _41081_ = _41072_ & _41080_ /*29090*/;
assign _40756_ = _41072_ ^ _41080_ /*29091*/;
assign _41078_ = _41079_ | _41081_ /*29088*/;
assign _41083_ = ~Q[18] /*29087*/;
assign _41082_ = _41083_ & D[52] /*29086*/;
assign _41085_ = _40309_ & _41082_ /*29081*/;
assign _41086_ = _40309_ ^ _41082_ /*29084*/;
assign _41087_ = _41078_ & _41086_ /*29082*/;
assign _40757_ = _41078_ ^ _41086_ /*29083*/;
assign _41084_ = _41085_ | _41087_ /*29080*/;
assign _41089_ = ~Q[18] /*29079*/;
assign _41088_ = _41089_ & D[53] /*29078*/;
assign _41091_ = _40310_ & _41088_ /*29073*/;
assign _41092_ = _40310_ ^ _41088_ /*29076*/;
assign _41093_ = _41084_ & _41092_ /*29074*/;
assign _40758_ = _41084_ ^ _41092_ /*29075*/;
assign _41090_ = _41091_ | _41093_ /*29072*/;
assign _41095_ = ~Q[18] /*29071*/;
assign _41094_ = _41095_ & D[54] /*29070*/;
assign _41097_ = _40311_ & _41094_ /*29065*/;
assign _41098_ = _40311_ ^ _41094_ /*29068*/;
assign _41099_ = _41090_ & _41098_ /*29066*/;
assign _40759_ = _41090_ ^ _41098_ /*29067*/;
assign _41096_ = _41097_ | _41099_ /*29064*/;
assign _41101_ = ~Q[18] /*29063*/;
assign _41100_ = _41101_ & D[55] /*29062*/;
assign _41103_ = _40312_ & _41100_ /*29057*/;
assign _41104_ = _40312_ ^ _41100_ /*29060*/;
assign _41105_ = _41096_ & _41104_ /*29058*/;
assign _40760_ = _41096_ ^ _41104_ /*29059*/;
assign _41102_ = _41103_ | _41105_ /*29056*/;
assign _41107_ = ~Q[18] /*29055*/;
assign _41106_ = _41107_ & D[56] /*29054*/;
assign _41109_ = _40313_ & _41106_ /*29049*/;
assign _41110_ = _40313_ ^ _41106_ /*29052*/;
assign _41111_ = _41102_ & _41110_ /*29050*/;
assign _40761_ = _41102_ ^ _41110_ /*29051*/;
assign _41108_ = _41109_ | _41111_ /*29048*/;
assign _41113_ = ~Q[18] /*29047*/;
assign _41112_ = _41113_ & D[57] /*29046*/;
assign _41115_ = _40314_ & _41112_ /*29041*/;
assign _41116_ = _40314_ ^ _41112_ /*29044*/;
assign _41117_ = _41108_ & _41116_ /*29042*/;
assign _40762_ = _41108_ ^ _41116_ /*29043*/;
assign _41114_ = _41115_ | _41117_ /*29040*/;
assign _41119_ = ~Q[18] /*29039*/;
assign _41118_ = _41119_ & D[58] /*29038*/;
assign _41121_ = _40315_ & _41118_ /*29033*/;
assign _41122_ = _40315_ ^ _41118_ /*29036*/;
assign _41123_ = _41114_ & _41122_ /*29034*/;
assign _40763_ = _41114_ ^ _41122_ /*29035*/;
assign _41120_ = _41121_ | _41123_ /*29032*/;
assign _41125_ = ~Q[18] /*29031*/;
assign _41124_ = _41125_ & D[59] /*29030*/;
assign _41127_ = _40316_ & _41124_ /*29025*/;
assign _41128_ = _40316_ ^ _41124_ /*29028*/;
assign _41129_ = _41120_ & _41128_ /*29026*/;
assign _40764_ = _41120_ ^ _41128_ /*29027*/;
assign _41126_ = _41127_ | _41129_ /*29024*/;
assign _41131_ = ~Q[18] /*29023*/;
assign _41130_ = _41131_ & D[60] /*29022*/;
assign _41133_ = _40317_ & _41130_ /*29017*/;
assign _41134_ = _40317_ ^ _41130_ /*29020*/;
assign _41135_ = _41126_ & _41134_ /*29018*/;
assign _40765_ = _41126_ ^ _41134_ /*29019*/;
assign _41132_ = _41133_ | _41135_ /*29016*/;
assign _41137_ = ~Q[18] /*29015*/;
assign _41136_ = _41137_ & D[61] /*29014*/;
assign _41139_ = _40318_ & _41136_ /*29009*/;
assign _41140_ = _40318_ ^ _41136_ /*29012*/;
assign _41141_ = _41132_ & _41140_ /*29010*/;
assign _40766_ = _41132_ ^ _41140_ /*29011*/;
assign _41138_ = _41139_ | _41141_ /*29008*/;
assign _41143_ = ~Q[18] /*29007*/;
assign _41142_ = _41143_ & D[62] /*29006*/;
assign _41145_ = _40319_ & _41142_ /*29001*/;
assign _41146_ = _40319_ ^ _41142_ /*29004*/;
assign _41147_ = _41138_ & _41146_ /*29002*/;
assign _40767_ = _41138_ ^ _41146_ /*29003*/;
assign _41144_ = _41145_ | _41147_ /*29000*/;
assign _41149_ = ~Q[18] /*28999*/;
assign _41148_ = _41149_ & zeroWire /*28998*/;
assign _41150_ = _40320_ ^ _41148_ /*28996*/;
assign _40768_ = _41150_ ^ _41144_ /*28995*/;
assign _41221_ = ~D[0] /*28741*/;
assign _41218_ = R_0[17] & _41221_ /*28737*/;
assign _41219_ = R_0[17] ^ _41221_ /*28740*/;
assign _41220_ = oneWire & _41219_ /*28738*/;
assign _41153_ = oneWire ^ _41219_ /*28739*/;
assign _41217_ = _41218_ | _41220_ /*28736*/;
assign _41226_ = ~D[1] /*28735*/;
assign _41223_ = _40705_ & _41226_ /*28731*/;
assign _41224_ = _40705_ ^ _41226_ /*28734*/;
assign _41225_ = _41217_ & _41224_ /*28732*/;
assign _41154_ = _41217_ ^ _41224_ /*28733*/;
assign _41222_ = _41223_ | _41225_ /*28730*/;
assign _41231_ = ~D[2] /*28729*/;
assign _41228_ = _40706_ & _41231_ /*28725*/;
assign _41229_ = _40706_ ^ _41231_ /*28728*/;
assign _41230_ = _41222_ & _41229_ /*28726*/;
assign _41155_ = _41222_ ^ _41229_ /*28727*/;
assign _41227_ = _41228_ | _41230_ /*28724*/;
assign _41236_ = ~D[3] /*28723*/;
assign _41233_ = _40707_ & _41236_ /*28719*/;
assign _41234_ = _40707_ ^ _41236_ /*28722*/;
assign _41235_ = _41227_ & _41234_ /*28720*/;
assign _41156_ = _41227_ ^ _41234_ /*28721*/;
assign _41232_ = _41233_ | _41235_ /*28718*/;
assign _41241_ = ~D[4] /*28717*/;
assign _41238_ = _40708_ & _41241_ /*28713*/;
assign _41239_ = _40708_ ^ _41241_ /*28716*/;
assign _41240_ = _41232_ & _41239_ /*28714*/;
assign _41157_ = _41232_ ^ _41239_ /*28715*/;
assign _41237_ = _41238_ | _41240_ /*28712*/;
assign _41246_ = ~D[5] /*28711*/;
assign _41243_ = _40709_ & _41246_ /*28707*/;
assign _41244_ = _40709_ ^ _41246_ /*28710*/;
assign _41245_ = _41237_ & _41244_ /*28708*/;
assign _41158_ = _41237_ ^ _41244_ /*28709*/;
assign _41242_ = _41243_ | _41245_ /*28706*/;
assign _41251_ = ~D[6] /*28705*/;
assign _41248_ = _40710_ & _41251_ /*28701*/;
assign _41249_ = _40710_ ^ _41251_ /*28704*/;
assign _41250_ = _41242_ & _41249_ /*28702*/;
assign _41159_ = _41242_ ^ _41249_ /*28703*/;
assign _41247_ = _41248_ | _41250_ /*28700*/;
assign _41256_ = ~D[7] /*28699*/;
assign _41253_ = _40711_ & _41256_ /*28695*/;
assign _41254_ = _40711_ ^ _41256_ /*28698*/;
assign _41255_ = _41247_ & _41254_ /*28696*/;
assign _41160_ = _41247_ ^ _41254_ /*28697*/;
assign _41252_ = _41253_ | _41255_ /*28694*/;
assign _41261_ = ~D[8] /*28693*/;
assign _41258_ = _40712_ & _41261_ /*28689*/;
assign _41259_ = _40712_ ^ _41261_ /*28692*/;
assign _41260_ = _41252_ & _41259_ /*28690*/;
assign _41161_ = _41252_ ^ _41259_ /*28691*/;
assign _41257_ = _41258_ | _41260_ /*28688*/;
assign _41266_ = ~D[9] /*28687*/;
assign _41263_ = _40713_ & _41266_ /*28683*/;
assign _41264_ = _40713_ ^ _41266_ /*28686*/;
assign _41265_ = _41257_ & _41264_ /*28684*/;
assign _41162_ = _41257_ ^ _41264_ /*28685*/;
assign _41262_ = _41263_ | _41265_ /*28682*/;
assign _41271_ = ~D[10] /*28681*/;
assign _41268_ = _40714_ & _41271_ /*28677*/;
assign _41269_ = _40714_ ^ _41271_ /*28680*/;
assign _41270_ = _41262_ & _41269_ /*28678*/;
assign _41163_ = _41262_ ^ _41269_ /*28679*/;
assign _41267_ = _41268_ | _41270_ /*28676*/;
assign _41276_ = ~D[11] /*28675*/;
assign _41273_ = _40715_ & _41276_ /*28671*/;
assign _41274_ = _40715_ ^ _41276_ /*28674*/;
assign _41275_ = _41267_ & _41274_ /*28672*/;
assign _41164_ = _41267_ ^ _41274_ /*28673*/;
assign _41272_ = _41273_ | _41275_ /*28670*/;
assign _41281_ = ~D[12] /*28669*/;
assign _41278_ = _40716_ & _41281_ /*28665*/;
assign _41279_ = _40716_ ^ _41281_ /*28668*/;
assign _41280_ = _41272_ & _41279_ /*28666*/;
assign _41165_ = _41272_ ^ _41279_ /*28667*/;
assign _41277_ = _41278_ | _41280_ /*28664*/;
assign _41286_ = ~D[13] /*28663*/;
assign _41283_ = _40717_ & _41286_ /*28659*/;
assign _41284_ = _40717_ ^ _41286_ /*28662*/;
assign _41285_ = _41277_ & _41284_ /*28660*/;
assign _41166_ = _41277_ ^ _41284_ /*28661*/;
assign _41282_ = _41283_ | _41285_ /*28658*/;
assign _41291_ = ~D[14] /*28657*/;
assign _41288_ = _40718_ & _41291_ /*28653*/;
assign _41289_ = _40718_ ^ _41291_ /*28656*/;
assign _41290_ = _41282_ & _41289_ /*28654*/;
assign _41167_ = _41282_ ^ _41289_ /*28655*/;
assign _41287_ = _41288_ | _41290_ /*28652*/;
assign _41296_ = ~D[15] /*28651*/;
assign _41293_ = _40719_ & _41296_ /*28647*/;
assign _41294_ = _40719_ ^ _41296_ /*28650*/;
assign _41295_ = _41287_ & _41294_ /*28648*/;
assign _41168_ = _41287_ ^ _41294_ /*28649*/;
assign _41292_ = _41293_ | _41295_ /*28646*/;
assign _41301_ = ~D[16] /*28645*/;
assign _41298_ = _40720_ & _41301_ /*28641*/;
assign _41299_ = _40720_ ^ _41301_ /*28644*/;
assign _41300_ = _41292_ & _41299_ /*28642*/;
assign _41169_ = _41292_ ^ _41299_ /*28643*/;
assign _41297_ = _41298_ | _41300_ /*28640*/;
assign _41306_ = ~D[17] /*28639*/;
assign _41303_ = _40721_ & _41306_ /*28635*/;
assign _41304_ = _40721_ ^ _41306_ /*28638*/;
assign _41305_ = _41297_ & _41304_ /*28636*/;
assign _41170_ = _41297_ ^ _41304_ /*28637*/;
assign _41302_ = _41303_ | _41305_ /*28634*/;
assign _41311_ = ~D[18] /*28633*/;
assign _41308_ = _40722_ & _41311_ /*28629*/;
assign _41309_ = _40722_ ^ _41311_ /*28632*/;
assign _41310_ = _41302_ & _41309_ /*28630*/;
assign _41171_ = _41302_ ^ _41309_ /*28631*/;
assign _41307_ = _41308_ | _41310_ /*28628*/;
assign _41316_ = ~D[19] /*28627*/;
assign _41313_ = _40723_ & _41316_ /*28623*/;
assign _41314_ = _40723_ ^ _41316_ /*28626*/;
assign _41315_ = _41307_ & _41314_ /*28624*/;
assign _41172_ = _41307_ ^ _41314_ /*28625*/;
assign _41312_ = _41313_ | _41315_ /*28622*/;
assign _41321_ = ~D[20] /*28621*/;
assign _41318_ = _40724_ & _41321_ /*28617*/;
assign _41319_ = _40724_ ^ _41321_ /*28620*/;
assign _41320_ = _41312_ & _41319_ /*28618*/;
assign _41173_ = _41312_ ^ _41319_ /*28619*/;
assign _41317_ = _41318_ | _41320_ /*28616*/;
assign _41326_ = ~D[21] /*28615*/;
assign _41323_ = _40725_ & _41326_ /*28611*/;
assign _41324_ = _40725_ ^ _41326_ /*28614*/;
assign _41325_ = _41317_ & _41324_ /*28612*/;
assign _41174_ = _41317_ ^ _41324_ /*28613*/;
assign _41322_ = _41323_ | _41325_ /*28610*/;
assign _41331_ = ~D[22] /*28609*/;
assign _41328_ = _40726_ & _41331_ /*28605*/;
assign _41329_ = _40726_ ^ _41331_ /*28608*/;
assign _41330_ = _41322_ & _41329_ /*28606*/;
assign _41175_ = _41322_ ^ _41329_ /*28607*/;
assign _41327_ = _41328_ | _41330_ /*28604*/;
assign _41336_ = ~D[23] /*28603*/;
assign _41333_ = _40727_ & _41336_ /*28599*/;
assign _41334_ = _40727_ ^ _41336_ /*28602*/;
assign _41335_ = _41327_ & _41334_ /*28600*/;
assign _41176_ = _41327_ ^ _41334_ /*28601*/;
assign _41332_ = _41333_ | _41335_ /*28598*/;
assign _41341_ = ~D[24] /*28597*/;
assign _41338_ = _40728_ & _41341_ /*28593*/;
assign _41339_ = _40728_ ^ _41341_ /*28596*/;
assign _41340_ = _41332_ & _41339_ /*28594*/;
assign _41177_ = _41332_ ^ _41339_ /*28595*/;
assign _41337_ = _41338_ | _41340_ /*28592*/;
assign _41346_ = ~D[25] /*28591*/;
assign _41343_ = _40729_ & _41346_ /*28587*/;
assign _41344_ = _40729_ ^ _41346_ /*28590*/;
assign _41345_ = _41337_ & _41344_ /*28588*/;
assign _41178_ = _41337_ ^ _41344_ /*28589*/;
assign _41342_ = _41343_ | _41345_ /*28586*/;
assign _41351_ = ~D[26] /*28585*/;
assign _41348_ = _40730_ & _41351_ /*28581*/;
assign _41349_ = _40730_ ^ _41351_ /*28584*/;
assign _41350_ = _41342_ & _41349_ /*28582*/;
assign _41179_ = _41342_ ^ _41349_ /*28583*/;
assign _41347_ = _41348_ | _41350_ /*28580*/;
assign _41356_ = ~D[27] /*28579*/;
assign _41353_ = _40731_ & _41356_ /*28575*/;
assign _41354_ = _40731_ ^ _41356_ /*28578*/;
assign _41355_ = _41347_ & _41354_ /*28576*/;
assign _41180_ = _41347_ ^ _41354_ /*28577*/;
assign _41352_ = _41353_ | _41355_ /*28574*/;
assign _41361_ = ~D[28] /*28573*/;
assign _41358_ = _40732_ & _41361_ /*28569*/;
assign _41359_ = _40732_ ^ _41361_ /*28572*/;
assign _41360_ = _41352_ & _41359_ /*28570*/;
assign _41181_ = _41352_ ^ _41359_ /*28571*/;
assign _41357_ = _41358_ | _41360_ /*28568*/;
assign _41366_ = ~D[29] /*28567*/;
assign _41363_ = _40733_ & _41366_ /*28563*/;
assign _41364_ = _40733_ ^ _41366_ /*28566*/;
assign _41365_ = _41357_ & _41364_ /*28564*/;
assign _41182_ = _41357_ ^ _41364_ /*28565*/;
assign _41362_ = _41363_ | _41365_ /*28562*/;
assign _41371_ = ~D[30] /*28561*/;
assign _41368_ = _40734_ & _41371_ /*28557*/;
assign _41369_ = _40734_ ^ _41371_ /*28560*/;
assign _41370_ = _41362_ & _41369_ /*28558*/;
assign _41183_ = _41362_ ^ _41369_ /*28559*/;
assign _41367_ = _41368_ | _41370_ /*28556*/;
assign _41376_ = ~D[31] /*28555*/;
assign _41373_ = _40735_ & _41376_ /*28551*/;
assign _41374_ = _40735_ ^ _41376_ /*28554*/;
assign _41375_ = _41367_ & _41374_ /*28552*/;
assign _41184_ = _41367_ ^ _41374_ /*28553*/;
assign _41372_ = _41373_ | _41375_ /*28550*/;
assign _41381_ = ~D[32] /*28549*/;
assign _41378_ = _40736_ & _41381_ /*28545*/;
assign _41379_ = _40736_ ^ _41381_ /*28548*/;
assign _41380_ = _41372_ & _41379_ /*28546*/;
assign _41185_ = _41372_ ^ _41379_ /*28547*/;
assign _41377_ = _41378_ | _41380_ /*28544*/;
assign _41386_ = ~D[33] /*28543*/;
assign _41383_ = _40737_ & _41386_ /*28539*/;
assign _41384_ = _40737_ ^ _41386_ /*28542*/;
assign _41385_ = _41377_ & _41384_ /*28540*/;
assign _41186_ = _41377_ ^ _41384_ /*28541*/;
assign _41382_ = _41383_ | _41385_ /*28538*/;
assign _41391_ = ~D[34] /*28537*/;
assign _41388_ = _40738_ & _41391_ /*28533*/;
assign _41389_ = _40738_ ^ _41391_ /*28536*/;
assign _41390_ = _41382_ & _41389_ /*28534*/;
assign _41187_ = _41382_ ^ _41389_ /*28535*/;
assign _41387_ = _41388_ | _41390_ /*28532*/;
assign _41396_ = ~D[35] /*28531*/;
assign _41393_ = _40739_ & _41396_ /*28527*/;
assign _41394_ = _40739_ ^ _41396_ /*28530*/;
assign _41395_ = _41387_ & _41394_ /*28528*/;
assign _41188_ = _41387_ ^ _41394_ /*28529*/;
assign _41392_ = _41393_ | _41395_ /*28526*/;
assign _41401_ = ~D[36] /*28525*/;
assign _41398_ = _40740_ & _41401_ /*28521*/;
assign _41399_ = _40740_ ^ _41401_ /*28524*/;
assign _41400_ = _41392_ & _41399_ /*28522*/;
assign _41189_ = _41392_ ^ _41399_ /*28523*/;
assign _41397_ = _41398_ | _41400_ /*28520*/;
assign _41406_ = ~D[37] /*28519*/;
assign _41403_ = _40741_ & _41406_ /*28515*/;
assign _41404_ = _40741_ ^ _41406_ /*28518*/;
assign _41405_ = _41397_ & _41404_ /*28516*/;
assign _41190_ = _41397_ ^ _41404_ /*28517*/;
assign _41402_ = _41403_ | _41405_ /*28514*/;
assign _41411_ = ~D[38] /*28513*/;
assign _41408_ = _40742_ & _41411_ /*28509*/;
assign _41409_ = _40742_ ^ _41411_ /*28512*/;
assign _41410_ = _41402_ & _41409_ /*28510*/;
assign _41191_ = _41402_ ^ _41409_ /*28511*/;
assign _41407_ = _41408_ | _41410_ /*28508*/;
assign _41416_ = ~D[39] /*28507*/;
assign _41413_ = _40743_ & _41416_ /*28503*/;
assign _41414_ = _40743_ ^ _41416_ /*28506*/;
assign _41415_ = _41407_ & _41414_ /*28504*/;
assign _41192_ = _41407_ ^ _41414_ /*28505*/;
assign _41412_ = _41413_ | _41415_ /*28502*/;
assign _41421_ = ~D[40] /*28501*/;
assign _41418_ = _40744_ & _41421_ /*28497*/;
assign _41419_ = _40744_ ^ _41421_ /*28500*/;
assign _41420_ = _41412_ & _41419_ /*28498*/;
assign _41193_ = _41412_ ^ _41419_ /*28499*/;
assign _41417_ = _41418_ | _41420_ /*28496*/;
assign _41426_ = ~D[41] /*28495*/;
assign _41423_ = _40745_ & _41426_ /*28491*/;
assign _41424_ = _40745_ ^ _41426_ /*28494*/;
assign _41425_ = _41417_ & _41424_ /*28492*/;
assign _41194_ = _41417_ ^ _41424_ /*28493*/;
assign _41422_ = _41423_ | _41425_ /*28490*/;
assign _41431_ = ~D[42] /*28489*/;
assign _41428_ = _40746_ & _41431_ /*28485*/;
assign _41429_ = _40746_ ^ _41431_ /*28488*/;
assign _41430_ = _41422_ & _41429_ /*28486*/;
assign _41195_ = _41422_ ^ _41429_ /*28487*/;
assign _41427_ = _41428_ | _41430_ /*28484*/;
assign _41436_ = ~D[43] /*28483*/;
assign _41433_ = _40747_ & _41436_ /*28479*/;
assign _41434_ = _40747_ ^ _41436_ /*28482*/;
assign _41435_ = _41427_ & _41434_ /*28480*/;
assign _41196_ = _41427_ ^ _41434_ /*28481*/;
assign _41432_ = _41433_ | _41435_ /*28478*/;
assign _41441_ = ~D[44] /*28477*/;
assign _41438_ = _40748_ & _41441_ /*28473*/;
assign _41439_ = _40748_ ^ _41441_ /*28476*/;
assign _41440_ = _41432_ & _41439_ /*28474*/;
assign _41197_ = _41432_ ^ _41439_ /*28475*/;
assign _41437_ = _41438_ | _41440_ /*28472*/;
assign _41446_ = ~D[45] /*28471*/;
assign _41443_ = _40749_ & _41446_ /*28467*/;
assign _41444_ = _40749_ ^ _41446_ /*28470*/;
assign _41445_ = _41437_ & _41444_ /*28468*/;
assign _41198_ = _41437_ ^ _41444_ /*28469*/;
assign _41442_ = _41443_ | _41445_ /*28466*/;
assign _41451_ = ~D[46] /*28465*/;
assign _41448_ = _40750_ & _41451_ /*28461*/;
assign _41449_ = _40750_ ^ _41451_ /*28464*/;
assign _41450_ = _41442_ & _41449_ /*28462*/;
assign _41199_ = _41442_ ^ _41449_ /*28463*/;
assign _41447_ = _41448_ | _41450_ /*28460*/;
assign _41456_ = ~D[47] /*28459*/;
assign _41453_ = _40751_ & _41456_ /*28455*/;
assign _41454_ = _40751_ ^ _41456_ /*28458*/;
assign _41455_ = _41447_ & _41454_ /*28456*/;
assign _41200_ = _41447_ ^ _41454_ /*28457*/;
assign _41452_ = _41453_ | _41455_ /*28454*/;
assign _41461_ = ~D[48] /*28453*/;
assign _41458_ = _40752_ & _41461_ /*28449*/;
assign _41459_ = _40752_ ^ _41461_ /*28452*/;
assign _41460_ = _41452_ & _41459_ /*28450*/;
assign _41201_ = _41452_ ^ _41459_ /*28451*/;
assign _41457_ = _41458_ | _41460_ /*28448*/;
assign _41466_ = ~D[49] /*28447*/;
assign _41463_ = _40753_ & _41466_ /*28443*/;
assign _41464_ = _40753_ ^ _41466_ /*28446*/;
assign _41465_ = _41457_ & _41464_ /*28444*/;
assign _41202_ = _41457_ ^ _41464_ /*28445*/;
assign _41462_ = _41463_ | _41465_ /*28442*/;
assign _41471_ = ~D[50] /*28441*/;
assign _41468_ = _40754_ & _41471_ /*28437*/;
assign _41469_ = _40754_ ^ _41471_ /*28440*/;
assign _41470_ = _41462_ & _41469_ /*28438*/;
assign _41203_ = _41462_ ^ _41469_ /*28439*/;
assign _41467_ = _41468_ | _41470_ /*28436*/;
assign _41476_ = ~D[51] /*28435*/;
assign _41473_ = _40755_ & _41476_ /*28431*/;
assign _41474_ = _40755_ ^ _41476_ /*28434*/;
assign _41475_ = _41467_ & _41474_ /*28432*/;
assign _41204_ = _41467_ ^ _41474_ /*28433*/;
assign _41472_ = _41473_ | _41475_ /*28430*/;
assign _41481_ = ~D[52] /*28429*/;
assign _41478_ = _40756_ & _41481_ /*28425*/;
assign _41479_ = _40756_ ^ _41481_ /*28428*/;
assign _41480_ = _41472_ & _41479_ /*28426*/;
assign _41205_ = _41472_ ^ _41479_ /*28427*/;
assign _41477_ = _41478_ | _41480_ /*28424*/;
assign _41486_ = ~D[53] /*28423*/;
assign _41483_ = _40757_ & _41486_ /*28419*/;
assign _41484_ = _40757_ ^ _41486_ /*28422*/;
assign _41485_ = _41477_ & _41484_ /*28420*/;
assign _41206_ = _41477_ ^ _41484_ /*28421*/;
assign _41482_ = _41483_ | _41485_ /*28418*/;
assign _41491_ = ~D[54] /*28417*/;
assign _41488_ = _40758_ & _41491_ /*28413*/;
assign _41489_ = _40758_ ^ _41491_ /*28416*/;
assign _41490_ = _41482_ & _41489_ /*28414*/;
assign _41207_ = _41482_ ^ _41489_ /*28415*/;
assign _41487_ = _41488_ | _41490_ /*28412*/;
assign _41496_ = ~D[55] /*28411*/;
assign _41493_ = _40759_ & _41496_ /*28407*/;
assign _41494_ = _40759_ ^ _41496_ /*28410*/;
assign _41495_ = _41487_ & _41494_ /*28408*/;
assign _41208_ = _41487_ ^ _41494_ /*28409*/;
assign _41492_ = _41493_ | _41495_ /*28406*/;
assign _41501_ = ~D[56] /*28405*/;
assign _41498_ = _40760_ & _41501_ /*28401*/;
assign _41499_ = _40760_ ^ _41501_ /*28404*/;
assign _41500_ = _41492_ & _41499_ /*28402*/;
assign _41209_ = _41492_ ^ _41499_ /*28403*/;
assign _41497_ = _41498_ | _41500_ /*28400*/;
assign _41506_ = ~D[57] /*28399*/;
assign _41503_ = _40761_ & _41506_ /*28395*/;
assign _41504_ = _40761_ ^ _41506_ /*28398*/;
assign _41505_ = _41497_ & _41504_ /*28396*/;
assign _41210_ = _41497_ ^ _41504_ /*28397*/;
assign _41502_ = _41503_ | _41505_ /*28394*/;
assign _41511_ = ~D[58] /*28393*/;
assign _41508_ = _40762_ & _41511_ /*28389*/;
assign _41509_ = _40762_ ^ _41511_ /*28392*/;
assign _41510_ = _41502_ & _41509_ /*28390*/;
assign _41211_ = _41502_ ^ _41509_ /*28391*/;
assign _41507_ = _41508_ | _41510_ /*28388*/;
assign _41516_ = ~D[59] /*28387*/;
assign _41513_ = _40763_ & _41516_ /*28383*/;
assign _41514_ = _40763_ ^ _41516_ /*28386*/;
assign _41515_ = _41507_ & _41514_ /*28384*/;
assign _41212_ = _41507_ ^ _41514_ /*28385*/;
assign _41512_ = _41513_ | _41515_ /*28382*/;
assign _41521_ = ~D[60] /*28381*/;
assign _41518_ = _40764_ & _41521_ /*28377*/;
assign _41519_ = _40764_ ^ _41521_ /*28380*/;
assign _41520_ = _41512_ & _41519_ /*28378*/;
assign _41213_ = _41512_ ^ _41519_ /*28379*/;
assign _41517_ = _41518_ | _41520_ /*28376*/;
assign _41526_ = ~D[61] /*28375*/;
assign _41523_ = _40765_ & _41526_ /*28371*/;
assign _41524_ = _40765_ ^ _41526_ /*28374*/;
assign _41525_ = _41517_ & _41524_ /*28372*/;
assign _41214_ = _41517_ ^ _41524_ /*28373*/;
assign _41522_ = _41523_ | _41525_ /*28370*/;
assign _41531_ = ~D[62] /*28369*/;
assign _41528_ = _40766_ & _41531_ /*28365*/;
assign _41529_ = _40766_ ^ _41531_ /*28368*/;
assign _41530_ = _41522_ & _41529_ /*28366*/;
assign _41215_ = _41522_ ^ _41529_ /*28367*/;
assign _41527_ = _41528_ | _41530_ /*28364*/;
assign _41532_ = _40767_ & oneWire /*28359*/;
assign _41533_ = _40767_ ^ oneWire /*28362*/;
assign _41534_ = _41527_ & _41533_ /*28360*/;
assign _41216_ = _41527_ ^ _41533_ /*28361*/;
assign Q[17] = _41532_ | _41534_ /*28358*/;
assign _41667_ = ~Q[17] /*27973*/;
assign _41666_ = _41667_ & D[0] /*27972*/;
assign _41669_ = _41153_ & _41666_ /*27967*/;
assign _41670_ = _41153_ ^ _41666_ /*27970*/;
assign _41671_ = zeroWire & _41670_ /*27968*/;
assign _41601_ = zeroWire ^ _41670_ /*27969*/;
assign _41668_ = _41669_ | _41671_ /*27966*/;
assign _41673_ = ~Q[17] /*27965*/;
assign _41672_ = _41673_ & D[1] /*27964*/;
assign _41675_ = _41154_ & _41672_ /*27959*/;
assign _41676_ = _41154_ ^ _41672_ /*27962*/;
assign _41677_ = _41668_ & _41676_ /*27960*/;
assign _41602_ = _41668_ ^ _41676_ /*27961*/;
assign _41674_ = _41675_ | _41677_ /*27958*/;
assign _41679_ = ~Q[17] /*27957*/;
assign _41678_ = _41679_ & D[2] /*27956*/;
assign _41681_ = _41155_ & _41678_ /*27951*/;
assign _41682_ = _41155_ ^ _41678_ /*27954*/;
assign _41683_ = _41674_ & _41682_ /*27952*/;
assign _41603_ = _41674_ ^ _41682_ /*27953*/;
assign _41680_ = _41681_ | _41683_ /*27950*/;
assign _41685_ = ~Q[17] /*27949*/;
assign _41684_ = _41685_ & D[3] /*27948*/;
assign _41687_ = _41156_ & _41684_ /*27943*/;
assign _41688_ = _41156_ ^ _41684_ /*27946*/;
assign _41689_ = _41680_ & _41688_ /*27944*/;
assign _41604_ = _41680_ ^ _41688_ /*27945*/;
assign _41686_ = _41687_ | _41689_ /*27942*/;
assign _41691_ = ~Q[17] /*27941*/;
assign _41690_ = _41691_ & D[4] /*27940*/;
assign _41693_ = _41157_ & _41690_ /*27935*/;
assign _41694_ = _41157_ ^ _41690_ /*27938*/;
assign _41695_ = _41686_ & _41694_ /*27936*/;
assign _41605_ = _41686_ ^ _41694_ /*27937*/;
assign _41692_ = _41693_ | _41695_ /*27934*/;
assign _41697_ = ~Q[17] /*27933*/;
assign _41696_ = _41697_ & D[5] /*27932*/;
assign _41699_ = _41158_ & _41696_ /*27927*/;
assign _41700_ = _41158_ ^ _41696_ /*27930*/;
assign _41701_ = _41692_ & _41700_ /*27928*/;
assign _41606_ = _41692_ ^ _41700_ /*27929*/;
assign _41698_ = _41699_ | _41701_ /*27926*/;
assign _41703_ = ~Q[17] /*27925*/;
assign _41702_ = _41703_ & D[6] /*27924*/;
assign _41705_ = _41159_ & _41702_ /*27919*/;
assign _41706_ = _41159_ ^ _41702_ /*27922*/;
assign _41707_ = _41698_ & _41706_ /*27920*/;
assign _41607_ = _41698_ ^ _41706_ /*27921*/;
assign _41704_ = _41705_ | _41707_ /*27918*/;
assign _41709_ = ~Q[17] /*27917*/;
assign _41708_ = _41709_ & D[7] /*27916*/;
assign _41711_ = _41160_ & _41708_ /*27911*/;
assign _41712_ = _41160_ ^ _41708_ /*27914*/;
assign _41713_ = _41704_ & _41712_ /*27912*/;
assign _41608_ = _41704_ ^ _41712_ /*27913*/;
assign _41710_ = _41711_ | _41713_ /*27910*/;
assign _41715_ = ~Q[17] /*27909*/;
assign _41714_ = _41715_ & D[8] /*27908*/;
assign _41717_ = _41161_ & _41714_ /*27903*/;
assign _41718_ = _41161_ ^ _41714_ /*27906*/;
assign _41719_ = _41710_ & _41718_ /*27904*/;
assign _41609_ = _41710_ ^ _41718_ /*27905*/;
assign _41716_ = _41717_ | _41719_ /*27902*/;
assign _41721_ = ~Q[17] /*27901*/;
assign _41720_ = _41721_ & D[9] /*27900*/;
assign _41723_ = _41162_ & _41720_ /*27895*/;
assign _41724_ = _41162_ ^ _41720_ /*27898*/;
assign _41725_ = _41716_ & _41724_ /*27896*/;
assign _41610_ = _41716_ ^ _41724_ /*27897*/;
assign _41722_ = _41723_ | _41725_ /*27894*/;
assign _41727_ = ~Q[17] /*27893*/;
assign _41726_ = _41727_ & D[10] /*27892*/;
assign _41729_ = _41163_ & _41726_ /*27887*/;
assign _41730_ = _41163_ ^ _41726_ /*27890*/;
assign _41731_ = _41722_ & _41730_ /*27888*/;
assign _41611_ = _41722_ ^ _41730_ /*27889*/;
assign _41728_ = _41729_ | _41731_ /*27886*/;
assign _41733_ = ~Q[17] /*27885*/;
assign _41732_ = _41733_ & D[11] /*27884*/;
assign _41735_ = _41164_ & _41732_ /*27879*/;
assign _41736_ = _41164_ ^ _41732_ /*27882*/;
assign _41737_ = _41728_ & _41736_ /*27880*/;
assign _41612_ = _41728_ ^ _41736_ /*27881*/;
assign _41734_ = _41735_ | _41737_ /*27878*/;
assign _41739_ = ~Q[17] /*27877*/;
assign _41738_ = _41739_ & D[12] /*27876*/;
assign _41741_ = _41165_ & _41738_ /*27871*/;
assign _41742_ = _41165_ ^ _41738_ /*27874*/;
assign _41743_ = _41734_ & _41742_ /*27872*/;
assign _41613_ = _41734_ ^ _41742_ /*27873*/;
assign _41740_ = _41741_ | _41743_ /*27870*/;
assign _41745_ = ~Q[17] /*27869*/;
assign _41744_ = _41745_ & D[13] /*27868*/;
assign _41747_ = _41166_ & _41744_ /*27863*/;
assign _41748_ = _41166_ ^ _41744_ /*27866*/;
assign _41749_ = _41740_ & _41748_ /*27864*/;
assign _41614_ = _41740_ ^ _41748_ /*27865*/;
assign _41746_ = _41747_ | _41749_ /*27862*/;
assign _41751_ = ~Q[17] /*27861*/;
assign _41750_ = _41751_ & D[14] /*27860*/;
assign _41753_ = _41167_ & _41750_ /*27855*/;
assign _41754_ = _41167_ ^ _41750_ /*27858*/;
assign _41755_ = _41746_ & _41754_ /*27856*/;
assign _41615_ = _41746_ ^ _41754_ /*27857*/;
assign _41752_ = _41753_ | _41755_ /*27854*/;
assign _41757_ = ~Q[17] /*27853*/;
assign _41756_ = _41757_ & D[15] /*27852*/;
assign _41759_ = _41168_ & _41756_ /*27847*/;
assign _41760_ = _41168_ ^ _41756_ /*27850*/;
assign _41761_ = _41752_ & _41760_ /*27848*/;
assign _41616_ = _41752_ ^ _41760_ /*27849*/;
assign _41758_ = _41759_ | _41761_ /*27846*/;
assign _41763_ = ~Q[17] /*27845*/;
assign _41762_ = _41763_ & D[16] /*27844*/;
assign _41765_ = _41169_ & _41762_ /*27839*/;
assign _41766_ = _41169_ ^ _41762_ /*27842*/;
assign _41767_ = _41758_ & _41766_ /*27840*/;
assign _41617_ = _41758_ ^ _41766_ /*27841*/;
assign _41764_ = _41765_ | _41767_ /*27838*/;
assign _41769_ = ~Q[17] /*27837*/;
assign _41768_ = _41769_ & D[17] /*27836*/;
assign _41771_ = _41170_ & _41768_ /*27831*/;
assign _41772_ = _41170_ ^ _41768_ /*27834*/;
assign _41773_ = _41764_ & _41772_ /*27832*/;
assign _41618_ = _41764_ ^ _41772_ /*27833*/;
assign _41770_ = _41771_ | _41773_ /*27830*/;
assign _41775_ = ~Q[17] /*27829*/;
assign _41774_ = _41775_ & D[18] /*27828*/;
assign _41777_ = _41171_ & _41774_ /*27823*/;
assign _41778_ = _41171_ ^ _41774_ /*27826*/;
assign _41779_ = _41770_ & _41778_ /*27824*/;
assign _41619_ = _41770_ ^ _41778_ /*27825*/;
assign _41776_ = _41777_ | _41779_ /*27822*/;
assign _41781_ = ~Q[17] /*27821*/;
assign _41780_ = _41781_ & D[19] /*27820*/;
assign _41783_ = _41172_ & _41780_ /*27815*/;
assign _41784_ = _41172_ ^ _41780_ /*27818*/;
assign _41785_ = _41776_ & _41784_ /*27816*/;
assign _41620_ = _41776_ ^ _41784_ /*27817*/;
assign _41782_ = _41783_ | _41785_ /*27814*/;
assign _41787_ = ~Q[17] /*27813*/;
assign _41786_ = _41787_ & D[20] /*27812*/;
assign _41789_ = _41173_ & _41786_ /*27807*/;
assign _41790_ = _41173_ ^ _41786_ /*27810*/;
assign _41791_ = _41782_ & _41790_ /*27808*/;
assign _41621_ = _41782_ ^ _41790_ /*27809*/;
assign _41788_ = _41789_ | _41791_ /*27806*/;
assign _41793_ = ~Q[17] /*27805*/;
assign _41792_ = _41793_ & D[21] /*27804*/;
assign _41795_ = _41174_ & _41792_ /*27799*/;
assign _41796_ = _41174_ ^ _41792_ /*27802*/;
assign _41797_ = _41788_ & _41796_ /*27800*/;
assign _41622_ = _41788_ ^ _41796_ /*27801*/;
assign _41794_ = _41795_ | _41797_ /*27798*/;
assign _41799_ = ~Q[17] /*27797*/;
assign _41798_ = _41799_ & D[22] /*27796*/;
assign _41801_ = _41175_ & _41798_ /*27791*/;
assign _41802_ = _41175_ ^ _41798_ /*27794*/;
assign _41803_ = _41794_ & _41802_ /*27792*/;
assign _41623_ = _41794_ ^ _41802_ /*27793*/;
assign _41800_ = _41801_ | _41803_ /*27790*/;
assign _41805_ = ~Q[17] /*27789*/;
assign _41804_ = _41805_ & D[23] /*27788*/;
assign _41807_ = _41176_ & _41804_ /*27783*/;
assign _41808_ = _41176_ ^ _41804_ /*27786*/;
assign _41809_ = _41800_ & _41808_ /*27784*/;
assign _41624_ = _41800_ ^ _41808_ /*27785*/;
assign _41806_ = _41807_ | _41809_ /*27782*/;
assign _41811_ = ~Q[17] /*27781*/;
assign _41810_ = _41811_ & D[24] /*27780*/;
assign _41813_ = _41177_ & _41810_ /*27775*/;
assign _41814_ = _41177_ ^ _41810_ /*27778*/;
assign _41815_ = _41806_ & _41814_ /*27776*/;
assign _41625_ = _41806_ ^ _41814_ /*27777*/;
assign _41812_ = _41813_ | _41815_ /*27774*/;
assign _41817_ = ~Q[17] /*27773*/;
assign _41816_ = _41817_ & D[25] /*27772*/;
assign _41819_ = _41178_ & _41816_ /*27767*/;
assign _41820_ = _41178_ ^ _41816_ /*27770*/;
assign _41821_ = _41812_ & _41820_ /*27768*/;
assign _41626_ = _41812_ ^ _41820_ /*27769*/;
assign _41818_ = _41819_ | _41821_ /*27766*/;
assign _41823_ = ~Q[17] /*27765*/;
assign _41822_ = _41823_ & D[26] /*27764*/;
assign _41825_ = _41179_ & _41822_ /*27759*/;
assign _41826_ = _41179_ ^ _41822_ /*27762*/;
assign _41827_ = _41818_ & _41826_ /*27760*/;
assign _41627_ = _41818_ ^ _41826_ /*27761*/;
assign _41824_ = _41825_ | _41827_ /*27758*/;
assign _41829_ = ~Q[17] /*27757*/;
assign _41828_ = _41829_ & D[27] /*27756*/;
assign _41831_ = _41180_ & _41828_ /*27751*/;
assign _41832_ = _41180_ ^ _41828_ /*27754*/;
assign _41833_ = _41824_ & _41832_ /*27752*/;
assign _41628_ = _41824_ ^ _41832_ /*27753*/;
assign _41830_ = _41831_ | _41833_ /*27750*/;
assign _41835_ = ~Q[17] /*27749*/;
assign _41834_ = _41835_ & D[28] /*27748*/;
assign _41837_ = _41181_ & _41834_ /*27743*/;
assign _41838_ = _41181_ ^ _41834_ /*27746*/;
assign _41839_ = _41830_ & _41838_ /*27744*/;
assign _41629_ = _41830_ ^ _41838_ /*27745*/;
assign _41836_ = _41837_ | _41839_ /*27742*/;
assign _41841_ = ~Q[17] /*27741*/;
assign _41840_ = _41841_ & D[29] /*27740*/;
assign _41843_ = _41182_ & _41840_ /*27735*/;
assign _41844_ = _41182_ ^ _41840_ /*27738*/;
assign _41845_ = _41836_ & _41844_ /*27736*/;
assign _41630_ = _41836_ ^ _41844_ /*27737*/;
assign _41842_ = _41843_ | _41845_ /*27734*/;
assign _41847_ = ~Q[17] /*27733*/;
assign _41846_ = _41847_ & D[30] /*27732*/;
assign _41849_ = _41183_ & _41846_ /*27727*/;
assign _41850_ = _41183_ ^ _41846_ /*27730*/;
assign _41851_ = _41842_ & _41850_ /*27728*/;
assign _41631_ = _41842_ ^ _41850_ /*27729*/;
assign _41848_ = _41849_ | _41851_ /*27726*/;
assign _41853_ = ~Q[17] /*27725*/;
assign _41852_ = _41853_ & D[31] /*27724*/;
assign _41855_ = _41184_ & _41852_ /*27719*/;
assign _41856_ = _41184_ ^ _41852_ /*27722*/;
assign _41857_ = _41848_ & _41856_ /*27720*/;
assign _41632_ = _41848_ ^ _41856_ /*27721*/;
assign _41854_ = _41855_ | _41857_ /*27718*/;
assign _41859_ = ~Q[17] /*27717*/;
assign _41858_ = _41859_ & D[32] /*27716*/;
assign _41861_ = _41185_ & _41858_ /*27711*/;
assign _41862_ = _41185_ ^ _41858_ /*27714*/;
assign _41863_ = _41854_ & _41862_ /*27712*/;
assign _41633_ = _41854_ ^ _41862_ /*27713*/;
assign _41860_ = _41861_ | _41863_ /*27710*/;
assign _41865_ = ~Q[17] /*27709*/;
assign _41864_ = _41865_ & D[33] /*27708*/;
assign _41867_ = _41186_ & _41864_ /*27703*/;
assign _41868_ = _41186_ ^ _41864_ /*27706*/;
assign _41869_ = _41860_ & _41868_ /*27704*/;
assign _41634_ = _41860_ ^ _41868_ /*27705*/;
assign _41866_ = _41867_ | _41869_ /*27702*/;
assign _41871_ = ~Q[17] /*27701*/;
assign _41870_ = _41871_ & D[34] /*27700*/;
assign _41873_ = _41187_ & _41870_ /*27695*/;
assign _41874_ = _41187_ ^ _41870_ /*27698*/;
assign _41875_ = _41866_ & _41874_ /*27696*/;
assign _41635_ = _41866_ ^ _41874_ /*27697*/;
assign _41872_ = _41873_ | _41875_ /*27694*/;
assign _41877_ = ~Q[17] /*27693*/;
assign _41876_ = _41877_ & D[35] /*27692*/;
assign _41879_ = _41188_ & _41876_ /*27687*/;
assign _41880_ = _41188_ ^ _41876_ /*27690*/;
assign _41881_ = _41872_ & _41880_ /*27688*/;
assign _41636_ = _41872_ ^ _41880_ /*27689*/;
assign _41878_ = _41879_ | _41881_ /*27686*/;
assign _41883_ = ~Q[17] /*27685*/;
assign _41882_ = _41883_ & D[36] /*27684*/;
assign _41885_ = _41189_ & _41882_ /*27679*/;
assign _41886_ = _41189_ ^ _41882_ /*27682*/;
assign _41887_ = _41878_ & _41886_ /*27680*/;
assign _41637_ = _41878_ ^ _41886_ /*27681*/;
assign _41884_ = _41885_ | _41887_ /*27678*/;
assign _41889_ = ~Q[17] /*27677*/;
assign _41888_ = _41889_ & D[37] /*27676*/;
assign _41891_ = _41190_ & _41888_ /*27671*/;
assign _41892_ = _41190_ ^ _41888_ /*27674*/;
assign _41893_ = _41884_ & _41892_ /*27672*/;
assign _41638_ = _41884_ ^ _41892_ /*27673*/;
assign _41890_ = _41891_ | _41893_ /*27670*/;
assign _41895_ = ~Q[17] /*27669*/;
assign _41894_ = _41895_ & D[38] /*27668*/;
assign _41897_ = _41191_ & _41894_ /*27663*/;
assign _41898_ = _41191_ ^ _41894_ /*27666*/;
assign _41899_ = _41890_ & _41898_ /*27664*/;
assign _41639_ = _41890_ ^ _41898_ /*27665*/;
assign _41896_ = _41897_ | _41899_ /*27662*/;
assign _41901_ = ~Q[17] /*27661*/;
assign _41900_ = _41901_ & D[39] /*27660*/;
assign _41903_ = _41192_ & _41900_ /*27655*/;
assign _41904_ = _41192_ ^ _41900_ /*27658*/;
assign _41905_ = _41896_ & _41904_ /*27656*/;
assign _41640_ = _41896_ ^ _41904_ /*27657*/;
assign _41902_ = _41903_ | _41905_ /*27654*/;
assign _41907_ = ~Q[17] /*27653*/;
assign _41906_ = _41907_ & D[40] /*27652*/;
assign _41909_ = _41193_ & _41906_ /*27647*/;
assign _41910_ = _41193_ ^ _41906_ /*27650*/;
assign _41911_ = _41902_ & _41910_ /*27648*/;
assign _41641_ = _41902_ ^ _41910_ /*27649*/;
assign _41908_ = _41909_ | _41911_ /*27646*/;
assign _41913_ = ~Q[17] /*27645*/;
assign _41912_ = _41913_ & D[41] /*27644*/;
assign _41915_ = _41194_ & _41912_ /*27639*/;
assign _41916_ = _41194_ ^ _41912_ /*27642*/;
assign _41917_ = _41908_ & _41916_ /*27640*/;
assign _41642_ = _41908_ ^ _41916_ /*27641*/;
assign _41914_ = _41915_ | _41917_ /*27638*/;
assign _41919_ = ~Q[17] /*27637*/;
assign _41918_ = _41919_ & D[42] /*27636*/;
assign _41921_ = _41195_ & _41918_ /*27631*/;
assign _41922_ = _41195_ ^ _41918_ /*27634*/;
assign _41923_ = _41914_ & _41922_ /*27632*/;
assign _41643_ = _41914_ ^ _41922_ /*27633*/;
assign _41920_ = _41921_ | _41923_ /*27630*/;
assign _41925_ = ~Q[17] /*27629*/;
assign _41924_ = _41925_ & D[43] /*27628*/;
assign _41927_ = _41196_ & _41924_ /*27623*/;
assign _41928_ = _41196_ ^ _41924_ /*27626*/;
assign _41929_ = _41920_ & _41928_ /*27624*/;
assign _41644_ = _41920_ ^ _41928_ /*27625*/;
assign _41926_ = _41927_ | _41929_ /*27622*/;
assign _41931_ = ~Q[17] /*27621*/;
assign _41930_ = _41931_ & D[44] /*27620*/;
assign _41933_ = _41197_ & _41930_ /*27615*/;
assign _41934_ = _41197_ ^ _41930_ /*27618*/;
assign _41935_ = _41926_ & _41934_ /*27616*/;
assign _41645_ = _41926_ ^ _41934_ /*27617*/;
assign _41932_ = _41933_ | _41935_ /*27614*/;
assign _41937_ = ~Q[17] /*27613*/;
assign _41936_ = _41937_ & D[45] /*27612*/;
assign _41939_ = _41198_ & _41936_ /*27607*/;
assign _41940_ = _41198_ ^ _41936_ /*27610*/;
assign _41941_ = _41932_ & _41940_ /*27608*/;
assign _41646_ = _41932_ ^ _41940_ /*27609*/;
assign _41938_ = _41939_ | _41941_ /*27606*/;
assign _41943_ = ~Q[17] /*27605*/;
assign _41942_ = _41943_ & D[46] /*27604*/;
assign _41945_ = _41199_ & _41942_ /*27599*/;
assign _41946_ = _41199_ ^ _41942_ /*27602*/;
assign _41947_ = _41938_ & _41946_ /*27600*/;
assign _41647_ = _41938_ ^ _41946_ /*27601*/;
assign _41944_ = _41945_ | _41947_ /*27598*/;
assign _41949_ = ~Q[17] /*27597*/;
assign _41948_ = _41949_ & D[47] /*27596*/;
assign _41951_ = _41200_ & _41948_ /*27591*/;
assign _41952_ = _41200_ ^ _41948_ /*27594*/;
assign _41953_ = _41944_ & _41952_ /*27592*/;
assign _41648_ = _41944_ ^ _41952_ /*27593*/;
assign _41950_ = _41951_ | _41953_ /*27590*/;
assign _41955_ = ~Q[17] /*27589*/;
assign _41954_ = _41955_ & D[48] /*27588*/;
assign _41957_ = _41201_ & _41954_ /*27583*/;
assign _41958_ = _41201_ ^ _41954_ /*27586*/;
assign _41959_ = _41950_ & _41958_ /*27584*/;
assign _41649_ = _41950_ ^ _41958_ /*27585*/;
assign _41956_ = _41957_ | _41959_ /*27582*/;
assign _41961_ = ~Q[17] /*27581*/;
assign _41960_ = _41961_ & D[49] /*27580*/;
assign _41963_ = _41202_ & _41960_ /*27575*/;
assign _41964_ = _41202_ ^ _41960_ /*27578*/;
assign _41965_ = _41956_ & _41964_ /*27576*/;
assign _41650_ = _41956_ ^ _41964_ /*27577*/;
assign _41962_ = _41963_ | _41965_ /*27574*/;
assign _41967_ = ~Q[17] /*27573*/;
assign _41966_ = _41967_ & D[50] /*27572*/;
assign _41969_ = _41203_ & _41966_ /*27567*/;
assign _41970_ = _41203_ ^ _41966_ /*27570*/;
assign _41971_ = _41962_ & _41970_ /*27568*/;
assign _41651_ = _41962_ ^ _41970_ /*27569*/;
assign _41968_ = _41969_ | _41971_ /*27566*/;
assign _41973_ = ~Q[17] /*27565*/;
assign _41972_ = _41973_ & D[51] /*27564*/;
assign _41975_ = _41204_ & _41972_ /*27559*/;
assign _41976_ = _41204_ ^ _41972_ /*27562*/;
assign _41977_ = _41968_ & _41976_ /*27560*/;
assign _41652_ = _41968_ ^ _41976_ /*27561*/;
assign _41974_ = _41975_ | _41977_ /*27558*/;
assign _41979_ = ~Q[17] /*27557*/;
assign _41978_ = _41979_ & D[52] /*27556*/;
assign _41981_ = _41205_ & _41978_ /*27551*/;
assign _41982_ = _41205_ ^ _41978_ /*27554*/;
assign _41983_ = _41974_ & _41982_ /*27552*/;
assign _41653_ = _41974_ ^ _41982_ /*27553*/;
assign _41980_ = _41981_ | _41983_ /*27550*/;
assign _41985_ = ~Q[17] /*27549*/;
assign _41984_ = _41985_ & D[53] /*27548*/;
assign _41987_ = _41206_ & _41984_ /*27543*/;
assign _41988_ = _41206_ ^ _41984_ /*27546*/;
assign _41989_ = _41980_ & _41988_ /*27544*/;
assign _41654_ = _41980_ ^ _41988_ /*27545*/;
assign _41986_ = _41987_ | _41989_ /*27542*/;
assign _41991_ = ~Q[17] /*27541*/;
assign _41990_ = _41991_ & D[54] /*27540*/;
assign _41993_ = _41207_ & _41990_ /*27535*/;
assign _41994_ = _41207_ ^ _41990_ /*27538*/;
assign _41995_ = _41986_ & _41994_ /*27536*/;
assign _41655_ = _41986_ ^ _41994_ /*27537*/;
assign _41992_ = _41993_ | _41995_ /*27534*/;
assign _41997_ = ~Q[17] /*27533*/;
assign _41996_ = _41997_ & D[55] /*27532*/;
assign _41999_ = _41208_ & _41996_ /*27527*/;
assign _42000_ = _41208_ ^ _41996_ /*27530*/;
assign _42001_ = _41992_ & _42000_ /*27528*/;
assign _41656_ = _41992_ ^ _42000_ /*27529*/;
assign _41998_ = _41999_ | _42001_ /*27526*/;
assign _42003_ = ~Q[17] /*27525*/;
assign _42002_ = _42003_ & D[56] /*27524*/;
assign _42005_ = _41209_ & _42002_ /*27519*/;
assign _42006_ = _41209_ ^ _42002_ /*27522*/;
assign _42007_ = _41998_ & _42006_ /*27520*/;
assign _41657_ = _41998_ ^ _42006_ /*27521*/;
assign _42004_ = _42005_ | _42007_ /*27518*/;
assign _42009_ = ~Q[17] /*27517*/;
assign _42008_ = _42009_ & D[57] /*27516*/;
assign _42011_ = _41210_ & _42008_ /*27511*/;
assign _42012_ = _41210_ ^ _42008_ /*27514*/;
assign _42013_ = _42004_ & _42012_ /*27512*/;
assign _41658_ = _42004_ ^ _42012_ /*27513*/;
assign _42010_ = _42011_ | _42013_ /*27510*/;
assign _42015_ = ~Q[17] /*27509*/;
assign _42014_ = _42015_ & D[58] /*27508*/;
assign _42017_ = _41211_ & _42014_ /*27503*/;
assign _42018_ = _41211_ ^ _42014_ /*27506*/;
assign _42019_ = _42010_ & _42018_ /*27504*/;
assign _41659_ = _42010_ ^ _42018_ /*27505*/;
assign _42016_ = _42017_ | _42019_ /*27502*/;
assign _42021_ = ~Q[17] /*27501*/;
assign _42020_ = _42021_ & D[59] /*27500*/;
assign _42023_ = _41212_ & _42020_ /*27495*/;
assign _42024_ = _41212_ ^ _42020_ /*27498*/;
assign _42025_ = _42016_ & _42024_ /*27496*/;
assign _41660_ = _42016_ ^ _42024_ /*27497*/;
assign _42022_ = _42023_ | _42025_ /*27494*/;
assign _42027_ = ~Q[17] /*27493*/;
assign _42026_ = _42027_ & D[60] /*27492*/;
assign _42029_ = _41213_ & _42026_ /*27487*/;
assign _42030_ = _41213_ ^ _42026_ /*27490*/;
assign _42031_ = _42022_ & _42030_ /*27488*/;
assign _41661_ = _42022_ ^ _42030_ /*27489*/;
assign _42028_ = _42029_ | _42031_ /*27486*/;
assign _42033_ = ~Q[17] /*27485*/;
assign _42032_ = _42033_ & D[61] /*27484*/;
assign _42035_ = _41214_ & _42032_ /*27479*/;
assign _42036_ = _41214_ ^ _42032_ /*27482*/;
assign _42037_ = _42028_ & _42036_ /*27480*/;
assign _41662_ = _42028_ ^ _42036_ /*27481*/;
assign _42034_ = _42035_ | _42037_ /*27478*/;
assign _42039_ = ~Q[17] /*27477*/;
assign _42038_ = _42039_ & D[62] /*27476*/;
assign _42041_ = _41215_ & _42038_ /*27471*/;
assign _42042_ = _41215_ ^ _42038_ /*27474*/;
assign _42043_ = _42034_ & _42042_ /*27472*/;
assign _41663_ = _42034_ ^ _42042_ /*27473*/;
assign _42040_ = _42041_ | _42043_ /*27470*/;
assign _42045_ = ~Q[17] /*27469*/;
assign _42044_ = _42045_ & zeroWire /*27468*/;
assign _42046_ = _41216_ ^ _42044_ /*27466*/;
assign _41664_ = _42046_ ^ _42040_ /*27465*/;
assign _42117_ = ~D[0] /*27211*/;
assign _42114_ = R_0[16] & _42117_ /*27207*/;
assign _42115_ = R_0[16] ^ _42117_ /*27210*/;
assign _42116_ = oneWire & _42115_ /*27208*/;
assign _42049_ = oneWire ^ _42115_ /*27209*/;
assign _42113_ = _42114_ | _42116_ /*27206*/;
assign _42122_ = ~D[1] /*27205*/;
assign _42119_ = _41601_ & _42122_ /*27201*/;
assign _42120_ = _41601_ ^ _42122_ /*27204*/;
assign _42121_ = _42113_ & _42120_ /*27202*/;
assign _42050_ = _42113_ ^ _42120_ /*27203*/;
assign _42118_ = _42119_ | _42121_ /*27200*/;
assign _42127_ = ~D[2] /*27199*/;
assign _42124_ = _41602_ & _42127_ /*27195*/;
assign _42125_ = _41602_ ^ _42127_ /*27198*/;
assign _42126_ = _42118_ & _42125_ /*27196*/;
assign _42051_ = _42118_ ^ _42125_ /*27197*/;
assign _42123_ = _42124_ | _42126_ /*27194*/;
assign _42132_ = ~D[3] /*27193*/;
assign _42129_ = _41603_ & _42132_ /*27189*/;
assign _42130_ = _41603_ ^ _42132_ /*27192*/;
assign _42131_ = _42123_ & _42130_ /*27190*/;
assign _42052_ = _42123_ ^ _42130_ /*27191*/;
assign _42128_ = _42129_ | _42131_ /*27188*/;
assign _42137_ = ~D[4] /*27187*/;
assign _42134_ = _41604_ & _42137_ /*27183*/;
assign _42135_ = _41604_ ^ _42137_ /*27186*/;
assign _42136_ = _42128_ & _42135_ /*27184*/;
assign _42053_ = _42128_ ^ _42135_ /*27185*/;
assign _42133_ = _42134_ | _42136_ /*27182*/;
assign _42142_ = ~D[5] /*27181*/;
assign _42139_ = _41605_ & _42142_ /*27177*/;
assign _42140_ = _41605_ ^ _42142_ /*27180*/;
assign _42141_ = _42133_ & _42140_ /*27178*/;
assign _42054_ = _42133_ ^ _42140_ /*27179*/;
assign _42138_ = _42139_ | _42141_ /*27176*/;
assign _42147_ = ~D[6] /*27175*/;
assign _42144_ = _41606_ & _42147_ /*27171*/;
assign _42145_ = _41606_ ^ _42147_ /*27174*/;
assign _42146_ = _42138_ & _42145_ /*27172*/;
assign _42055_ = _42138_ ^ _42145_ /*27173*/;
assign _42143_ = _42144_ | _42146_ /*27170*/;
assign _42152_ = ~D[7] /*27169*/;
assign _42149_ = _41607_ & _42152_ /*27165*/;
assign _42150_ = _41607_ ^ _42152_ /*27168*/;
assign _42151_ = _42143_ & _42150_ /*27166*/;
assign _42056_ = _42143_ ^ _42150_ /*27167*/;
assign _42148_ = _42149_ | _42151_ /*27164*/;
assign _42157_ = ~D[8] /*27163*/;
assign _42154_ = _41608_ & _42157_ /*27159*/;
assign _42155_ = _41608_ ^ _42157_ /*27162*/;
assign _42156_ = _42148_ & _42155_ /*27160*/;
assign _42057_ = _42148_ ^ _42155_ /*27161*/;
assign _42153_ = _42154_ | _42156_ /*27158*/;
assign _42162_ = ~D[9] /*27157*/;
assign _42159_ = _41609_ & _42162_ /*27153*/;
assign _42160_ = _41609_ ^ _42162_ /*27156*/;
assign _42161_ = _42153_ & _42160_ /*27154*/;
assign _42058_ = _42153_ ^ _42160_ /*27155*/;
assign _42158_ = _42159_ | _42161_ /*27152*/;
assign _42167_ = ~D[10] /*27151*/;
assign _42164_ = _41610_ & _42167_ /*27147*/;
assign _42165_ = _41610_ ^ _42167_ /*27150*/;
assign _42166_ = _42158_ & _42165_ /*27148*/;
assign _42059_ = _42158_ ^ _42165_ /*27149*/;
assign _42163_ = _42164_ | _42166_ /*27146*/;
assign _42172_ = ~D[11] /*27145*/;
assign _42169_ = _41611_ & _42172_ /*27141*/;
assign _42170_ = _41611_ ^ _42172_ /*27144*/;
assign _42171_ = _42163_ & _42170_ /*27142*/;
assign _42060_ = _42163_ ^ _42170_ /*27143*/;
assign _42168_ = _42169_ | _42171_ /*27140*/;
assign _42177_ = ~D[12] /*27139*/;
assign _42174_ = _41612_ & _42177_ /*27135*/;
assign _42175_ = _41612_ ^ _42177_ /*27138*/;
assign _42176_ = _42168_ & _42175_ /*27136*/;
assign _42061_ = _42168_ ^ _42175_ /*27137*/;
assign _42173_ = _42174_ | _42176_ /*27134*/;
assign _42182_ = ~D[13] /*27133*/;
assign _42179_ = _41613_ & _42182_ /*27129*/;
assign _42180_ = _41613_ ^ _42182_ /*27132*/;
assign _42181_ = _42173_ & _42180_ /*27130*/;
assign _42062_ = _42173_ ^ _42180_ /*27131*/;
assign _42178_ = _42179_ | _42181_ /*27128*/;
assign _42187_ = ~D[14] /*27127*/;
assign _42184_ = _41614_ & _42187_ /*27123*/;
assign _42185_ = _41614_ ^ _42187_ /*27126*/;
assign _42186_ = _42178_ & _42185_ /*27124*/;
assign _42063_ = _42178_ ^ _42185_ /*27125*/;
assign _42183_ = _42184_ | _42186_ /*27122*/;
assign _42192_ = ~D[15] /*27121*/;
assign _42189_ = _41615_ & _42192_ /*27117*/;
assign _42190_ = _41615_ ^ _42192_ /*27120*/;
assign _42191_ = _42183_ & _42190_ /*27118*/;
assign _42064_ = _42183_ ^ _42190_ /*27119*/;
assign _42188_ = _42189_ | _42191_ /*27116*/;
assign _42197_ = ~D[16] /*27115*/;
assign _42194_ = _41616_ & _42197_ /*27111*/;
assign _42195_ = _41616_ ^ _42197_ /*27114*/;
assign _42196_ = _42188_ & _42195_ /*27112*/;
assign _42065_ = _42188_ ^ _42195_ /*27113*/;
assign _42193_ = _42194_ | _42196_ /*27110*/;
assign _42202_ = ~D[17] /*27109*/;
assign _42199_ = _41617_ & _42202_ /*27105*/;
assign _42200_ = _41617_ ^ _42202_ /*27108*/;
assign _42201_ = _42193_ & _42200_ /*27106*/;
assign _42066_ = _42193_ ^ _42200_ /*27107*/;
assign _42198_ = _42199_ | _42201_ /*27104*/;
assign _42207_ = ~D[18] /*27103*/;
assign _42204_ = _41618_ & _42207_ /*27099*/;
assign _42205_ = _41618_ ^ _42207_ /*27102*/;
assign _42206_ = _42198_ & _42205_ /*27100*/;
assign _42067_ = _42198_ ^ _42205_ /*27101*/;
assign _42203_ = _42204_ | _42206_ /*27098*/;
assign _42212_ = ~D[19] /*27097*/;
assign _42209_ = _41619_ & _42212_ /*27093*/;
assign _42210_ = _41619_ ^ _42212_ /*27096*/;
assign _42211_ = _42203_ & _42210_ /*27094*/;
assign _42068_ = _42203_ ^ _42210_ /*27095*/;
assign _42208_ = _42209_ | _42211_ /*27092*/;
assign _42217_ = ~D[20] /*27091*/;
assign _42214_ = _41620_ & _42217_ /*27087*/;
assign _42215_ = _41620_ ^ _42217_ /*27090*/;
assign _42216_ = _42208_ & _42215_ /*27088*/;
assign _42069_ = _42208_ ^ _42215_ /*27089*/;
assign _42213_ = _42214_ | _42216_ /*27086*/;
assign _42222_ = ~D[21] /*27085*/;
assign _42219_ = _41621_ & _42222_ /*27081*/;
assign _42220_ = _41621_ ^ _42222_ /*27084*/;
assign _42221_ = _42213_ & _42220_ /*27082*/;
assign _42070_ = _42213_ ^ _42220_ /*27083*/;
assign _42218_ = _42219_ | _42221_ /*27080*/;
assign _42227_ = ~D[22] /*27079*/;
assign _42224_ = _41622_ & _42227_ /*27075*/;
assign _42225_ = _41622_ ^ _42227_ /*27078*/;
assign _42226_ = _42218_ & _42225_ /*27076*/;
assign _42071_ = _42218_ ^ _42225_ /*27077*/;
assign _42223_ = _42224_ | _42226_ /*27074*/;
assign _42232_ = ~D[23] /*27073*/;
assign _42229_ = _41623_ & _42232_ /*27069*/;
assign _42230_ = _41623_ ^ _42232_ /*27072*/;
assign _42231_ = _42223_ & _42230_ /*27070*/;
assign _42072_ = _42223_ ^ _42230_ /*27071*/;
assign _42228_ = _42229_ | _42231_ /*27068*/;
assign _42237_ = ~D[24] /*27067*/;
assign _42234_ = _41624_ & _42237_ /*27063*/;
assign _42235_ = _41624_ ^ _42237_ /*27066*/;
assign _42236_ = _42228_ & _42235_ /*27064*/;
assign _42073_ = _42228_ ^ _42235_ /*27065*/;
assign _42233_ = _42234_ | _42236_ /*27062*/;
assign _42242_ = ~D[25] /*27061*/;
assign _42239_ = _41625_ & _42242_ /*27057*/;
assign _42240_ = _41625_ ^ _42242_ /*27060*/;
assign _42241_ = _42233_ & _42240_ /*27058*/;
assign _42074_ = _42233_ ^ _42240_ /*27059*/;
assign _42238_ = _42239_ | _42241_ /*27056*/;
assign _42247_ = ~D[26] /*27055*/;
assign _42244_ = _41626_ & _42247_ /*27051*/;
assign _42245_ = _41626_ ^ _42247_ /*27054*/;
assign _42246_ = _42238_ & _42245_ /*27052*/;
assign _42075_ = _42238_ ^ _42245_ /*27053*/;
assign _42243_ = _42244_ | _42246_ /*27050*/;
assign _42252_ = ~D[27] /*27049*/;
assign _42249_ = _41627_ & _42252_ /*27045*/;
assign _42250_ = _41627_ ^ _42252_ /*27048*/;
assign _42251_ = _42243_ & _42250_ /*27046*/;
assign _42076_ = _42243_ ^ _42250_ /*27047*/;
assign _42248_ = _42249_ | _42251_ /*27044*/;
assign _42257_ = ~D[28] /*27043*/;
assign _42254_ = _41628_ & _42257_ /*27039*/;
assign _42255_ = _41628_ ^ _42257_ /*27042*/;
assign _42256_ = _42248_ & _42255_ /*27040*/;
assign _42077_ = _42248_ ^ _42255_ /*27041*/;
assign _42253_ = _42254_ | _42256_ /*27038*/;
assign _42262_ = ~D[29] /*27037*/;
assign _42259_ = _41629_ & _42262_ /*27033*/;
assign _42260_ = _41629_ ^ _42262_ /*27036*/;
assign _42261_ = _42253_ & _42260_ /*27034*/;
assign _42078_ = _42253_ ^ _42260_ /*27035*/;
assign _42258_ = _42259_ | _42261_ /*27032*/;
assign _42267_ = ~D[30] /*27031*/;
assign _42264_ = _41630_ & _42267_ /*27027*/;
assign _42265_ = _41630_ ^ _42267_ /*27030*/;
assign _42266_ = _42258_ & _42265_ /*27028*/;
assign _42079_ = _42258_ ^ _42265_ /*27029*/;
assign _42263_ = _42264_ | _42266_ /*27026*/;
assign _42272_ = ~D[31] /*27025*/;
assign _42269_ = _41631_ & _42272_ /*27021*/;
assign _42270_ = _41631_ ^ _42272_ /*27024*/;
assign _42271_ = _42263_ & _42270_ /*27022*/;
assign _42080_ = _42263_ ^ _42270_ /*27023*/;
assign _42268_ = _42269_ | _42271_ /*27020*/;
assign _42277_ = ~D[32] /*27019*/;
assign _42274_ = _41632_ & _42277_ /*27015*/;
assign _42275_ = _41632_ ^ _42277_ /*27018*/;
assign _42276_ = _42268_ & _42275_ /*27016*/;
assign _42081_ = _42268_ ^ _42275_ /*27017*/;
assign _42273_ = _42274_ | _42276_ /*27014*/;
assign _42282_ = ~D[33] /*27013*/;
assign _42279_ = _41633_ & _42282_ /*27009*/;
assign _42280_ = _41633_ ^ _42282_ /*27012*/;
assign _42281_ = _42273_ & _42280_ /*27010*/;
assign _42082_ = _42273_ ^ _42280_ /*27011*/;
assign _42278_ = _42279_ | _42281_ /*27008*/;
assign _42287_ = ~D[34] /*27007*/;
assign _42284_ = _41634_ & _42287_ /*27003*/;
assign _42285_ = _41634_ ^ _42287_ /*27006*/;
assign _42286_ = _42278_ & _42285_ /*27004*/;
assign _42083_ = _42278_ ^ _42285_ /*27005*/;
assign _42283_ = _42284_ | _42286_ /*27002*/;
assign _42292_ = ~D[35] /*27001*/;
assign _42289_ = _41635_ & _42292_ /*26997*/;
assign _42290_ = _41635_ ^ _42292_ /*27000*/;
assign _42291_ = _42283_ & _42290_ /*26998*/;
assign _42084_ = _42283_ ^ _42290_ /*26999*/;
assign _42288_ = _42289_ | _42291_ /*26996*/;
assign _42297_ = ~D[36] /*26995*/;
assign _42294_ = _41636_ & _42297_ /*26991*/;
assign _42295_ = _41636_ ^ _42297_ /*26994*/;
assign _42296_ = _42288_ & _42295_ /*26992*/;
assign _42085_ = _42288_ ^ _42295_ /*26993*/;
assign _42293_ = _42294_ | _42296_ /*26990*/;
assign _42302_ = ~D[37] /*26989*/;
assign _42299_ = _41637_ & _42302_ /*26985*/;
assign _42300_ = _41637_ ^ _42302_ /*26988*/;
assign _42301_ = _42293_ & _42300_ /*26986*/;
assign _42086_ = _42293_ ^ _42300_ /*26987*/;
assign _42298_ = _42299_ | _42301_ /*26984*/;
assign _42307_ = ~D[38] /*26983*/;
assign _42304_ = _41638_ & _42307_ /*26979*/;
assign _42305_ = _41638_ ^ _42307_ /*26982*/;
assign _42306_ = _42298_ & _42305_ /*26980*/;
assign _42087_ = _42298_ ^ _42305_ /*26981*/;
assign _42303_ = _42304_ | _42306_ /*26978*/;
assign _42312_ = ~D[39] /*26977*/;
assign _42309_ = _41639_ & _42312_ /*26973*/;
assign _42310_ = _41639_ ^ _42312_ /*26976*/;
assign _42311_ = _42303_ & _42310_ /*26974*/;
assign _42088_ = _42303_ ^ _42310_ /*26975*/;
assign _42308_ = _42309_ | _42311_ /*26972*/;
assign _42317_ = ~D[40] /*26971*/;
assign _42314_ = _41640_ & _42317_ /*26967*/;
assign _42315_ = _41640_ ^ _42317_ /*26970*/;
assign _42316_ = _42308_ & _42315_ /*26968*/;
assign _42089_ = _42308_ ^ _42315_ /*26969*/;
assign _42313_ = _42314_ | _42316_ /*26966*/;
assign _42322_ = ~D[41] /*26965*/;
assign _42319_ = _41641_ & _42322_ /*26961*/;
assign _42320_ = _41641_ ^ _42322_ /*26964*/;
assign _42321_ = _42313_ & _42320_ /*26962*/;
assign _42090_ = _42313_ ^ _42320_ /*26963*/;
assign _42318_ = _42319_ | _42321_ /*26960*/;
assign _42327_ = ~D[42] /*26959*/;
assign _42324_ = _41642_ & _42327_ /*26955*/;
assign _42325_ = _41642_ ^ _42327_ /*26958*/;
assign _42326_ = _42318_ & _42325_ /*26956*/;
assign _42091_ = _42318_ ^ _42325_ /*26957*/;
assign _42323_ = _42324_ | _42326_ /*26954*/;
assign _42332_ = ~D[43] /*26953*/;
assign _42329_ = _41643_ & _42332_ /*26949*/;
assign _42330_ = _41643_ ^ _42332_ /*26952*/;
assign _42331_ = _42323_ & _42330_ /*26950*/;
assign _42092_ = _42323_ ^ _42330_ /*26951*/;
assign _42328_ = _42329_ | _42331_ /*26948*/;
assign _42337_ = ~D[44] /*26947*/;
assign _42334_ = _41644_ & _42337_ /*26943*/;
assign _42335_ = _41644_ ^ _42337_ /*26946*/;
assign _42336_ = _42328_ & _42335_ /*26944*/;
assign _42093_ = _42328_ ^ _42335_ /*26945*/;
assign _42333_ = _42334_ | _42336_ /*26942*/;
assign _42342_ = ~D[45] /*26941*/;
assign _42339_ = _41645_ & _42342_ /*26937*/;
assign _42340_ = _41645_ ^ _42342_ /*26940*/;
assign _42341_ = _42333_ & _42340_ /*26938*/;
assign _42094_ = _42333_ ^ _42340_ /*26939*/;
assign _42338_ = _42339_ | _42341_ /*26936*/;
assign _42347_ = ~D[46] /*26935*/;
assign _42344_ = _41646_ & _42347_ /*26931*/;
assign _42345_ = _41646_ ^ _42347_ /*26934*/;
assign _42346_ = _42338_ & _42345_ /*26932*/;
assign _42095_ = _42338_ ^ _42345_ /*26933*/;
assign _42343_ = _42344_ | _42346_ /*26930*/;
assign _42352_ = ~D[47] /*26929*/;
assign _42349_ = _41647_ & _42352_ /*26925*/;
assign _42350_ = _41647_ ^ _42352_ /*26928*/;
assign _42351_ = _42343_ & _42350_ /*26926*/;
assign _42096_ = _42343_ ^ _42350_ /*26927*/;
assign _42348_ = _42349_ | _42351_ /*26924*/;
assign _42357_ = ~D[48] /*26923*/;
assign _42354_ = _41648_ & _42357_ /*26919*/;
assign _42355_ = _41648_ ^ _42357_ /*26922*/;
assign _42356_ = _42348_ & _42355_ /*26920*/;
assign _42097_ = _42348_ ^ _42355_ /*26921*/;
assign _42353_ = _42354_ | _42356_ /*26918*/;
assign _42362_ = ~D[49] /*26917*/;
assign _42359_ = _41649_ & _42362_ /*26913*/;
assign _42360_ = _41649_ ^ _42362_ /*26916*/;
assign _42361_ = _42353_ & _42360_ /*26914*/;
assign _42098_ = _42353_ ^ _42360_ /*26915*/;
assign _42358_ = _42359_ | _42361_ /*26912*/;
assign _42367_ = ~D[50] /*26911*/;
assign _42364_ = _41650_ & _42367_ /*26907*/;
assign _42365_ = _41650_ ^ _42367_ /*26910*/;
assign _42366_ = _42358_ & _42365_ /*26908*/;
assign _42099_ = _42358_ ^ _42365_ /*26909*/;
assign _42363_ = _42364_ | _42366_ /*26906*/;
assign _42372_ = ~D[51] /*26905*/;
assign _42369_ = _41651_ & _42372_ /*26901*/;
assign _42370_ = _41651_ ^ _42372_ /*26904*/;
assign _42371_ = _42363_ & _42370_ /*26902*/;
assign _42100_ = _42363_ ^ _42370_ /*26903*/;
assign _42368_ = _42369_ | _42371_ /*26900*/;
assign _42377_ = ~D[52] /*26899*/;
assign _42374_ = _41652_ & _42377_ /*26895*/;
assign _42375_ = _41652_ ^ _42377_ /*26898*/;
assign _42376_ = _42368_ & _42375_ /*26896*/;
assign _42101_ = _42368_ ^ _42375_ /*26897*/;
assign _42373_ = _42374_ | _42376_ /*26894*/;
assign _42382_ = ~D[53] /*26893*/;
assign _42379_ = _41653_ & _42382_ /*26889*/;
assign _42380_ = _41653_ ^ _42382_ /*26892*/;
assign _42381_ = _42373_ & _42380_ /*26890*/;
assign _42102_ = _42373_ ^ _42380_ /*26891*/;
assign _42378_ = _42379_ | _42381_ /*26888*/;
assign _42387_ = ~D[54] /*26887*/;
assign _42384_ = _41654_ & _42387_ /*26883*/;
assign _42385_ = _41654_ ^ _42387_ /*26886*/;
assign _42386_ = _42378_ & _42385_ /*26884*/;
assign _42103_ = _42378_ ^ _42385_ /*26885*/;
assign _42383_ = _42384_ | _42386_ /*26882*/;
assign _42392_ = ~D[55] /*26881*/;
assign _42389_ = _41655_ & _42392_ /*26877*/;
assign _42390_ = _41655_ ^ _42392_ /*26880*/;
assign _42391_ = _42383_ & _42390_ /*26878*/;
assign _42104_ = _42383_ ^ _42390_ /*26879*/;
assign _42388_ = _42389_ | _42391_ /*26876*/;
assign _42397_ = ~D[56] /*26875*/;
assign _42394_ = _41656_ & _42397_ /*26871*/;
assign _42395_ = _41656_ ^ _42397_ /*26874*/;
assign _42396_ = _42388_ & _42395_ /*26872*/;
assign _42105_ = _42388_ ^ _42395_ /*26873*/;
assign _42393_ = _42394_ | _42396_ /*26870*/;
assign _42402_ = ~D[57] /*26869*/;
assign _42399_ = _41657_ & _42402_ /*26865*/;
assign _42400_ = _41657_ ^ _42402_ /*26868*/;
assign _42401_ = _42393_ & _42400_ /*26866*/;
assign _42106_ = _42393_ ^ _42400_ /*26867*/;
assign _42398_ = _42399_ | _42401_ /*26864*/;
assign _42407_ = ~D[58] /*26863*/;
assign _42404_ = _41658_ & _42407_ /*26859*/;
assign _42405_ = _41658_ ^ _42407_ /*26862*/;
assign _42406_ = _42398_ & _42405_ /*26860*/;
assign _42107_ = _42398_ ^ _42405_ /*26861*/;
assign _42403_ = _42404_ | _42406_ /*26858*/;
assign _42412_ = ~D[59] /*26857*/;
assign _42409_ = _41659_ & _42412_ /*26853*/;
assign _42410_ = _41659_ ^ _42412_ /*26856*/;
assign _42411_ = _42403_ & _42410_ /*26854*/;
assign _42108_ = _42403_ ^ _42410_ /*26855*/;
assign _42408_ = _42409_ | _42411_ /*26852*/;
assign _42417_ = ~D[60] /*26851*/;
assign _42414_ = _41660_ & _42417_ /*26847*/;
assign _42415_ = _41660_ ^ _42417_ /*26850*/;
assign _42416_ = _42408_ & _42415_ /*26848*/;
assign _42109_ = _42408_ ^ _42415_ /*26849*/;
assign _42413_ = _42414_ | _42416_ /*26846*/;
assign _42422_ = ~D[61] /*26845*/;
assign _42419_ = _41661_ & _42422_ /*26841*/;
assign _42420_ = _41661_ ^ _42422_ /*26844*/;
assign _42421_ = _42413_ & _42420_ /*26842*/;
assign _42110_ = _42413_ ^ _42420_ /*26843*/;
assign _42418_ = _42419_ | _42421_ /*26840*/;
assign _42427_ = ~D[62] /*26839*/;
assign _42424_ = _41662_ & _42427_ /*26835*/;
assign _42425_ = _41662_ ^ _42427_ /*26838*/;
assign _42426_ = _42418_ & _42425_ /*26836*/;
assign _42111_ = _42418_ ^ _42425_ /*26837*/;
assign _42423_ = _42424_ | _42426_ /*26834*/;
assign _42428_ = _41663_ & oneWire /*26829*/;
assign _42429_ = _41663_ ^ oneWire /*26832*/;
assign _42430_ = _42423_ & _42429_ /*26830*/;
assign _42112_ = _42423_ ^ _42429_ /*26831*/;
assign Q[16] = _42428_ | _42430_ /*26828*/;
assign _42563_ = ~Q[16] /*26443*/;
assign _42562_ = _42563_ & D[0] /*26442*/;
assign _42565_ = _42049_ & _42562_ /*26437*/;
assign _42566_ = _42049_ ^ _42562_ /*26440*/;
assign _42567_ = zeroWire & _42566_ /*26438*/;
assign _42497_ = zeroWire ^ _42566_ /*26439*/;
assign _42564_ = _42565_ | _42567_ /*26436*/;
assign _42569_ = ~Q[16] /*26435*/;
assign _42568_ = _42569_ & D[1] /*26434*/;
assign _42571_ = _42050_ & _42568_ /*26429*/;
assign _42572_ = _42050_ ^ _42568_ /*26432*/;
assign _42573_ = _42564_ & _42572_ /*26430*/;
assign _42498_ = _42564_ ^ _42572_ /*26431*/;
assign _42570_ = _42571_ | _42573_ /*26428*/;
assign _42575_ = ~Q[16] /*26427*/;
assign _42574_ = _42575_ & D[2] /*26426*/;
assign _42577_ = _42051_ & _42574_ /*26421*/;
assign _42578_ = _42051_ ^ _42574_ /*26424*/;
assign _42579_ = _42570_ & _42578_ /*26422*/;
assign _42499_ = _42570_ ^ _42578_ /*26423*/;
assign _42576_ = _42577_ | _42579_ /*26420*/;
assign _42581_ = ~Q[16] /*26419*/;
assign _42580_ = _42581_ & D[3] /*26418*/;
assign _42583_ = _42052_ & _42580_ /*26413*/;
assign _42584_ = _42052_ ^ _42580_ /*26416*/;
assign _42585_ = _42576_ & _42584_ /*26414*/;
assign _42500_ = _42576_ ^ _42584_ /*26415*/;
assign _42582_ = _42583_ | _42585_ /*26412*/;
assign _42587_ = ~Q[16] /*26411*/;
assign _42586_ = _42587_ & D[4] /*26410*/;
assign _42589_ = _42053_ & _42586_ /*26405*/;
assign _42590_ = _42053_ ^ _42586_ /*26408*/;
assign _42591_ = _42582_ & _42590_ /*26406*/;
assign _42501_ = _42582_ ^ _42590_ /*26407*/;
assign _42588_ = _42589_ | _42591_ /*26404*/;
assign _42593_ = ~Q[16] /*26403*/;
assign _42592_ = _42593_ & D[5] /*26402*/;
assign _42595_ = _42054_ & _42592_ /*26397*/;
assign _42596_ = _42054_ ^ _42592_ /*26400*/;
assign _42597_ = _42588_ & _42596_ /*26398*/;
assign _42502_ = _42588_ ^ _42596_ /*26399*/;
assign _42594_ = _42595_ | _42597_ /*26396*/;
assign _42599_ = ~Q[16] /*26395*/;
assign _42598_ = _42599_ & D[6] /*26394*/;
assign _42601_ = _42055_ & _42598_ /*26389*/;
assign _42602_ = _42055_ ^ _42598_ /*26392*/;
assign _42603_ = _42594_ & _42602_ /*26390*/;
assign _42503_ = _42594_ ^ _42602_ /*26391*/;
assign _42600_ = _42601_ | _42603_ /*26388*/;
assign _42605_ = ~Q[16] /*26387*/;
assign _42604_ = _42605_ & D[7] /*26386*/;
assign _42607_ = _42056_ & _42604_ /*26381*/;
assign _42608_ = _42056_ ^ _42604_ /*26384*/;
assign _42609_ = _42600_ & _42608_ /*26382*/;
assign _42504_ = _42600_ ^ _42608_ /*26383*/;
assign _42606_ = _42607_ | _42609_ /*26380*/;
assign _42611_ = ~Q[16] /*26379*/;
assign _42610_ = _42611_ & D[8] /*26378*/;
assign _42613_ = _42057_ & _42610_ /*26373*/;
assign _42614_ = _42057_ ^ _42610_ /*26376*/;
assign _42615_ = _42606_ & _42614_ /*26374*/;
assign _42505_ = _42606_ ^ _42614_ /*26375*/;
assign _42612_ = _42613_ | _42615_ /*26372*/;
assign _42617_ = ~Q[16] /*26371*/;
assign _42616_ = _42617_ & D[9] /*26370*/;
assign _42619_ = _42058_ & _42616_ /*26365*/;
assign _42620_ = _42058_ ^ _42616_ /*26368*/;
assign _42621_ = _42612_ & _42620_ /*26366*/;
assign _42506_ = _42612_ ^ _42620_ /*26367*/;
assign _42618_ = _42619_ | _42621_ /*26364*/;
assign _42623_ = ~Q[16] /*26363*/;
assign _42622_ = _42623_ & D[10] /*26362*/;
assign _42625_ = _42059_ & _42622_ /*26357*/;
assign _42626_ = _42059_ ^ _42622_ /*26360*/;
assign _42627_ = _42618_ & _42626_ /*26358*/;
assign _42507_ = _42618_ ^ _42626_ /*26359*/;
assign _42624_ = _42625_ | _42627_ /*26356*/;
assign _42629_ = ~Q[16] /*26355*/;
assign _42628_ = _42629_ & D[11] /*26354*/;
assign _42631_ = _42060_ & _42628_ /*26349*/;
assign _42632_ = _42060_ ^ _42628_ /*26352*/;
assign _42633_ = _42624_ & _42632_ /*26350*/;
assign _42508_ = _42624_ ^ _42632_ /*26351*/;
assign _42630_ = _42631_ | _42633_ /*26348*/;
assign _42635_ = ~Q[16] /*26347*/;
assign _42634_ = _42635_ & D[12] /*26346*/;
assign _42637_ = _42061_ & _42634_ /*26341*/;
assign _42638_ = _42061_ ^ _42634_ /*26344*/;
assign _42639_ = _42630_ & _42638_ /*26342*/;
assign _42509_ = _42630_ ^ _42638_ /*26343*/;
assign _42636_ = _42637_ | _42639_ /*26340*/;
assign _42641_ = ~Q[16] /*26339*/;
assign _42640_ = _42641_ & D[13] /*26338*/;
assign _42643_ = _42062_ & _42640_ /*26333*/;
assign _42644_ = _42062_ ^ _42640_ /*26336*/;
assign _42645_ = _42636_ & _42644_ /*26334*/;
assign _42510_ = _42636_ ^ _42644_ /*26335*/;
assign _42642_ = _42643_ | _42645_ /*26332*/;
assign _42647_ = ~Q[16] /*26331*/;
assign _42646_ = _42647_ & D[14] /*26330*/;
assign _42649_ = _42063_ & _42646_ /*26325*/;
assign _42650_ = _42063_ ^ _42646_ /*26328*/;
assign _42651_ = _42642_ & _42650_ /*26326*/;
assign _42511_ = _42642_ ^ _42650_ /*26327*/;
assign _42648_ = _42649_ | _42651_ /*26324*/;
assign _42653_ = ~Q[16] /*26323*/;
assign _42652_ = _42653_ & D[15] /*26322*/;
assign _42655_ = _42064_ & _42652_ /*26317*/;
assign _42656_ = _42064_ ^ _42652_ /*26320*/;
assign _42657_ = _42648_ & _42656_ /*26318*/;
assign _42512_ = _42648_ ^ _42656_ /*26319*/;
assign _42654_ = _42655_ | _42657_ /*26316*/;
assign _42659_ = ~Q[16] /*26315*/;
assign _42658_ = _42659_ & D[16] /*26314*/;
assign _42661_ = _42065_ & _42658_ /*26309*/;
assign _42662_ = _42065_ ^ _42658_ /*26312*/;
assign _42663_ = _42654_ & _42662_ /*26310*/;
assign _42513_ = _42654_ ^ _42662_ /*26311*/;
assign _42660_ = _42661_ | _42663_ /*26308*/;
assign _42665_ = ~Q[16] /*26307*/;
assign _42664_ = _42665_ & D[17] /*26306*/;
assign _42667_ = _42066_ & _42664_ /*26301*/;
assign _42668_ = _42066_ ^ _42664_ /*26304*/;
assign _42669_ = _42660_ & _42668_ /*26302*/;
assign _42514_ = _42660_ ^ _42668_ /*26303*/;
assign _42666_ = _42667_ | _42669_ /*26300*/;
assign _42671_ = ~Q[16] /*26299*/;
assign _42670_ = _42671_ & D[18] /*26298*/;
assign _42673_ = _42067_ & _42670_ /*26293*/;
assign _42674_ = _42067_ ^ _42670_ /*26296*/;
assign _42675_ = _42666_ & _42674_ /*26294*/;
assign _42515_ = _42666_ ^ _42674_ /*26295*/;
assign _42672_ = _42673_ | _42675_ /*26292*/;
assign _42677_ = ~Q[16] /*26291*/;
assign _42676_ = _42677_ & D[19] /*26290*/;
assign _42679_ = _42068_ & _42676_ /*26285*/;
assign _42680_ = _42068_ ^ _42676_ /*26288*/;
assign _42681_ = _42672_ & _42680_ /*26286*/;
assign _42516_ = _42672_ ^ _42680_ /*26287*/;
assign _42678_ = _42679_ | _42681_ /*26284*/;
assign _42683_ = ~Q[16] /*26283*/;
assign _42682_ = _42683_ & D[20] /*26282*/;
assign _42685_ = _42069_ & _42682_ /*26277*/;
assign _42686_ = _42069_ ^ _42682_ /*26280*/;
assign _42687_ = _42678_ & _42686_ /*26278*/;
assign _42517_ = _42678_ ^ _42686_ /*26279*/;
assign _42684_ = _42685_ | _42687_ /*26276*/;
assign _42689_ = ~Q[16] /*26275*/;
assign _42688_ = _42689_ & D[21] /*26274*/;
assign _42691_ = _42070_ & _42688_ /*26269*/;
assign _42692_ = _42070_ ^ _42688_ /*26272*/;
assign _42693_ = _42684_ & _42692_ /*26270*/;
assign _42518_ = _42684_ ^ _42692_ /*26271*/;
assign _42690_ = _42691_ | _42693_ /*26268*/;
assign _42695_ = ~Q[16] /*26267*/;
assign _42694_ = _42695_ & D[22] /*26266*/;
assign _42697_ = _42071_ & _42694_ /*26261*/;
assign _42698_ = _42071_ ^ _42694_ /*26264*/;
assign _42699_ = _42690_ & _42698_ /*26262*/;
assign _42519_ = _42690_ ^ _42698_ /*26263*/;
assign _42696_ = _42697_ | _42699_ /*26260*/;
assign _42701_ = ~Q[16] /*26259*/;
assign _42700_ = _42701_ & D[23] /*26258*/;
assign _42703_ = _42072_ & _42700_ /*26253*/;
assign _42704_ = _42072_ ^ _42700_ /*26256*/;
assign _42705_ = _42696_ & _42704_ /*26254*/;
assign _42520_ = _42696_ ^ _42704_ /*26255*/;
assign _42702_ = _42703_ | _42705_ /*26252*/;
assign _42707_ = ~Q[16] /*26251*/;
assign _42706_ = _42707_ & D[24] /*26250*/;
assign _42709_ = _42073_ & _42706_ /*26245*/;
assign _42710_ = _42073_ ^ _42706_ /*26248*/;
assign _42711_ = _42702_ & _42710_ /*26246*/;
assign _42521_ = _42702_ ^ _42710_ /*26247*/;
assign _42708_ = _42709_ | _42711_ /*26244*/;
assign _42713_ = ~Q[16] /*26243*/;
assign _42712_ = _42713_ & D[25] /*26242*/;
assign _42715_ = _42074_ & _42712_ /*26237*/;
assign _42716_ = _42074_ ^ _42712_ /*26240*/;
assign _42717_ = _42708_ & _42716_ /*26238*/;
assign _42522_ = _42708_ ^ _42716_ /*26239*/;
assign _42714_ = _42715_ | _42717_ /*26236*/;
assign _42719_ = ~Q[16] /*26235*/;
assign _42718_ = _42719_ & D[26] /*26234*/;
assign _42721_ = _42075_ & _42718_ /*26229*/;
assign _42722_ = _42075_ ^ _42718_ /*26232*/;
assign _42723_ = _42714_ & _42722_ /*26230*/;
assign _42523_ = _42714_ ^ _42722_ /*26231*/;
assign _42720_ = _42721_ | _42723_ /*26228*/;
assign _42725_ = ~Q[16] /*26227*/;
assign _42724_ = _42725_ & D[27] /*26226*/;
assign _42727_ = _42076_ & _42724_ /*26221*/;
assign _42728_ = _42076_ ^ _42724_ /*26224*/;
assign _42729_ = _42720_ & _42728_ /*26222*/;
assign _42524_ = _42720_ ^ _42728_ /*26223*/;
assign _42726_ = _42727_ | _42729_ /*26220*/;
assign _42731_ = ~Q[16] /*26219*/;
assign _42730_ = _42731_ & D[28] /*26218*/;
assign _42733_ = _42077_ & _42730_ /*26213*/;
assign _42734_ = _42077_ ^ _42730_ /*26216*/;
assign _42735_ = _42726_ & _42734_ /*26214*/;
assign _42525_ = _42726_ ^ _42734_ /*26215*/;
assign _42732_ = _42733_ | _42735_ /*26212*/;
assign _42737_ = ~Q[16] /*26211*/;
assign _42736_ = _42737_ & D[29] /*26210*/;
assign _42739_ = _42078_ & _42736_ /*26205*/;
assign _42740_ = _42078_ ^ _42736_ /*26208*/;
assign _42741_ = _42732_ & _42740_ /*26206*/;
assign _42526_ = _42732_ ^ _42740_ /*26207*/;
assign _42738_ = _42739_ | _42741_ /*26204*/;
assign _42743_ = ~Q[16] /*26203*/;
assign _42742_ = _42743_ & D[30] /*26202*/;
assign _42745_ = _42079_ & _42742_ /*26197*/;
assign _42746_ = _42079_ ^ _42742_ /*26200*/;
assign _42747_ = _42738_ & _42746_ /*26198*/;
assign _42527_ = _42738_ ^ _42746_ /*26199*/;
assign _42744_ = _42745_ | _42747_ /*26196*/;
assign _42749_ = ~Q[16] /*26195*/;
assign _42748_ = _42749_ & D[31] /*26194*/;
assign _42751_ = _42080_ & _42748_ /*26189*/;
assign _42752_ = _42080_ ^ _42748_ /*26192*/;
assign _42753_ = _42744_ & _42752_ /*26190*/;
assign _42528_ = _42744_ ^ _42752_ /*26191*/;
assign _42750_ = _42751_ | _42753_ /*26188*/;
assign _42755_ = ~Q[16] /*26187*/;
assign _42754_ = _42755_ & D[32] /*26186*/;
assign _42757_ = _42081_ & _42754_ /*26181*/;
assign _42758_ = _42081_ ^ _42754_ /*26184*/;
assign _42759_ = _42750_ & _42758_ /*26182*/;
assign _42529_ = _42750_ ^ _42758_ /*26183*/;
assign _42756_ = _42757_ | _42759_ /*26180*/;
assign _42761_ = ~Q[16] /*26179*/;
assign _42760_ = _42761_ & D[33] /*26178*/;
assign _42763_ = _42082_ & _42760_ /*26173*/;
assign _42764_ = _42082_ ^ _42760_ /*26176*/;
assign _42765_ = _42756_ & _42764_ /*26174*/;
assign _42530_ = _42756_ ^ _42764_ /*26175*/;
assign _42762_ = _42763_ | _42765_ /*26172*/;
assign _42767_ = ~Q[16] /*26171*/;
assign _42766_ = _42767_ & D[34] /*26170*/;
assign _42769_ = _42083_ & _42766_ /*26165*/;
assign _42770_ = _42083_ ^ _42766_ /*26168*/;
assign _42771_ = _42762_ & _42770_ /*26166*/;
assign _42531_ = _42762_ ^ _42770_ /*26167*/;
assign _42768_ = _42769_ | _42771_ /*26164*/;
assign _42773_ = ~Q[16] /*26163*/;
assign _42772_ = _42773_ & D[35] /*26162*/;
assign _42775_ = _42084_ & _42772_ /*26157*/;
assign _42776_ = _42084_ ^ _42772_ /*26160*/;
assign _42777_ = _42768_ & _42776_ /*26158*/;
assign _42532_ = _42768_ ^ _42776_ /*26159*/;
assign _42774_ = _42775_ | _42777_ /*26156*/;
assign _42779_ = ~Q[16] /*26155*/;
assign _42778_ = _42779_ & D[36] /*26154*/;
assign _42781_ = _42085_ & _42778_ /*26149*/;
assign _42782_ = _42085_ ^ _42778_ /*26152*/;
assign _42783_ = _42774_ & _42782_ /*26150*/;
assign _42533_ = _42774_ ^ _42782_ /*26151*/;
assign _42780_ = _42781_ | _42783_ /*26148*/;
assign _42785_ = ~Q[16] /*26147*/;
assign _42784_ = _42785_ & D[37] /*26146*/;
assign _42787_ = _42086_ & _42784_ /*26141*/;
assign _42788_ = _42086_ ^ _42784_ /*26144*/;
assign _42789_ = _42780_ & _42788_ /*26142*/;
assign _42534_ = _42780_ ^ _42788_ /*26143*/;
assign _42786_ = _42787_ | _42789_ /*26140*/;
assign _42791_ = ~Q[16] /*26139*/;
assign _42790_ = _42791_ & D[38] /*26138*/;
assign _42793_ = _42087_ & _42790_ /*26133*/;
assign _42794_ = _42087_ ^ _42790_ /*26136*/;
assign _42795_ = _42786_ & _42794_ /*26134*/;
assign _42535_ = _42786_ ^ _42794_ /*26135*/;
assign _42792_ = _42793_ | _42795_ /*26132*/;
assign _42797_ = ~Q[16] /*26131*/;
assign _42796_ = _42797_ & D[39] /*26130*/;
assign _42799_ = _42088_ & _42796_ /*26125*/;
assign _42800_ = _42088_ ^ _42796_ /*26128*/;
assign _42801_ = _42792_ & _42800_ /*26126*/;
assign _42536_ = _42792_ ^ _42800_ /*26127*/;
assign _42798_ = _42799_ | _42801_ /*26124*/;
assign _42803_ = ~Q[16] /*26123*/;
assign _42802_ = _42803_ & D[40] /*26122*/;
assign _42805_ = _42089_ & _42802_ /*26117*/;
assign _42806_ = _42089_ ^ _42802_ /*26120*/;
assign _42807_ = _42798_ & _42806_ /*26118*/;
assign _42537_ = _42798_ ^ _42806_ /*26119*/;
assign _42804_ = _42805_ | _42807_ /*26116*/;
assign _42809_ = ~Q[16] /*26115*/;
assign _42808_ = _42809_ & D[41] /*26114*/;
assign _42811_ = _42090_ & _42808_ /*26109*/;
assign _42812_ = _42090_ ^ _42808_ /*26112*/;
assign _42813_ = _42804_ & _42812_ /*26110*/;
assign _42538_ = _42804_ ^ _42812_ /*26111*/;
assign _42810_ = _42811_ | _42813_ /*26108*/;
assign _42815_ = ~Q[16] /*26107*/;
assign _42814_ = _42815_ & D[42] /*26106*/;
assign _42817_ = _42091_ & _42814_ /*26101*/;
assign _42818_ = _42091_ ^ _42814_ /*26104*/;
assign _42819_ = _42810_ & _42818_ /*26102*/;
assign _42539_ = _42810_ ^ _42818_ /*26103*/;
assign _42816_ = _42817_ | _42819_ /*26100*/;
assign _42821_ = ~Q[16] /*26099*/;
assign _42820_ = _42821_ & D[43] /*26098*/;
assign _42823_ = _42092_ & _42820_ /*26093*/;
assign _42824_ = _42092_ ^ _42820_ /*26096*/;
assign _42825_ = _42816_ & _42824_ /*26094*/;
assign _42540_ = _42816_ ^ _42824_ /*26095*/;
assign _42822_ = _42823_ | _42825_ /*26092*/;
assign _42827_ = ~Q[16] /*26091*/;
assign _42826_ = _42827_ & D[44] /*26090*/;
assign _42829_ = _42093_ & _42826_ /*26085*/;
assign _42830_ = _42093_ ^ _42826_ /*26088*/;
assign _42831_ = _42822_ & _42830_ /*26086*/;
assign _42541_ = _42822_ ^ _42830_ /*26087*/;
assign _42828_ = _42829_ | _42831_ /*26084*/;
assign _42833_ = ~Q[16] /*26083*/;
assign _42832_ = _42833_ & D[45] /*26082*/;
assign _42835_ = _42094_ & _42832_ /*26077*/;
assign _42836_ = _42094_ ^ _42832_ /*26080*/;
assign _42837_ = _42828_ & _42836_ /*26078*/;
assign _42542_ = _42828_ ^ _42836_ /*26079*/;
assign _42834_ = _42835_ | _42837_ /*26076*/;
assign _42839_ = ~Q[16] /*26075*/;
assign _42838_ = _42839_ & D[46] /*26074*/;
assign _42841_ = _42095_ & _42838_ /*26069*/;
assign _42842_ = _42095_ ^ _42838_ /*26072*/;
assign _42843_ = _42834_ & _42842_ /*26070*/;
assign _42543_ = _42834_ ^ _42842_ /*26071*/;
assign _42840_ = _42841_ | _42843_ /*26068*/;
assign _42845_ = ~Q[16] /*26067*/;
assign _42844_ = _42845_ & D[47] /*26066*/;
assign _42847_ = _42096_ & _42844_ /*26061*/;
assign _42848_ = _42096_ ^ _42844_ /*26064*/;
assign _42849_ = _42840_ & _42848_ /*26062*/;
assign _42544_ = _42840_ ^ _42848_ /*26063*/;
assign _42846_ = _42847_ | _42849_ /*26060*/;
assign _42851_ = ~Q[16] /*26059*/;
assign _42850_ = _42851_ & D[48] /*26058*/;
assign _42853_ = _42097_ & _42850_ /*26053*/;
assign _42854_ = _42097_ ^ _42850_ /*26056*/;
assign _42855_ = _42846_ & _42854_ /*26054*/;
assign _42545_ = _42846_ ^ _42854_ /*26055*/;
assign _42852_ = _42853_ | _42855_ /*26052*/;
assign _42857_ = ~Q[16] /*26051*/;
assign _42856_ = _42857_ & D[49] /*26050*/;
assign _42859_ = _42098_ & _42856_ /*26045*/;
assign _42860_ = _42098_ ^ _42856_ /*26048*/;
assign _42861_ = _42852_ & _42860_ /*26046*/;
assign _42546_ = _42852_ ^ _42860_ /*26047*/;
assign _42858_ = _42859_ | _42861_ /*26044*/;
assign _42863_ = ~Q[16] /*26043*/;
assign _42862_ = _42863_ & D[50] /*26042*/;
assign _42865_ = _42099_ & _42862_ /*26037*/;
assign _42866_ = _42099_ ^ _42862_ /*26040*/;
assign _42867_ = _42858_ & _42866_ /*26038*/;
assign _42547_ = _42858_ ^ _42866_ /*26039*/;
assign _42864_ = _42865_ | _42867_ /*26036*/;
assign _42869_ = ~Q[16] /*26035*/;
assign _42868_ = _42869_ & D[51] /*26034*/;
assign _42871_ = _42100_ & _42868_ /*26029*/;
assign _42872_ = _42100_ ^ _42868_ /*26032*/;
assign _42873_ = _42864_ & _42872_ /*26030*/;
assign _42548_ = _42864_ ^ _42872_ /*26031*/;
assign _42870_ = _42871_ | _42873_ /*26028*/;
assign _42875_ = ~Q[16] /*26027*/;
assign _42874_ = _42875_ & D[52] /*26026*/;
assign _42877_ = _42101_ & _42874_ /*26021*/;
assign _42878_ = _42101_ ^ _42874_ /*26024*/;
assign _42879_ = _42870_ & _42878_ /*26022*/;
assign _42549_ = _42870_ ^ _42878_ /*26023*/;
assign _42876_ = _42877_ | _42879_ /*26020*/;
assign _42881_ = ~Q[16] /*26019*/;
assign _42880_ = _42881_ & D[53] /*26018*/;
assign _42883_ = _42102_ & _42880_ /*26013*/;
assign _42884_ = _42102_ ^ _42880_ /*26016*/;
assign _42885_ = _42876_ & _42884_ /*26014*/;
assign _42550_ = _42876_ ^ _42884_ /*26015*/;
assign _42882_ = _42883_ | _42885_ /*26012*/;
assign _42887_ = ~Q[16] /*26011*/;
assign _42886_ = _42887_ & D[54] /*26010*/;
assign _42889_ = _42103_ & _42886_ /*26005*/;
assign _42890_ = _42103_ ^ _42886_ /*26008*/;
assign _42891_ = _42882_ & _42890_ /*26006*/;
assign _42551_ = _42882_ ^ _42890_ /*26007*/;
assign _42888_ = _42889_ | _42891_ /*26004*/;
assign _42893_ = ~Q[16] /*26003*/;
assign _42892_ = _42893_ & D[55] /*26002*/;
assign _42895_ = _42104_ & _42892_ /*25997*/;
assign _42896_ = _42104_ ^ _42892_ /*26000*/;
assign _42897_ = _42888_ & _42896_ /*25998*/;
assign _42552_ = _42888_ ^ _42896_ /*25999*/;
assign _42894_ = _42895_ | _42897_ /*25996*/;
assign _42899_ = ~Q[16] /*25995*/;
assign _42898_ = _42899_ & D[56] /*25994*/;
assign _42901_ = _42105_ & _42898_ /*25989*/;
assign _42902_ = _42105_ ^ _42898_ /*25992*/;
assign _42903_ = _42894_ & _42902_ /*25990*/;
assign _42553_ = _42894_ ^ _42902_ /*25991*/;
assign _42900_ = _42901_ | _42903_ /*25988*/;
assign _42905_ = ~Q[16] /*25987*/;
assign _42904_ = _42905_ & D[57] /*25986*/;
assign _42907_ = _42106_ & _42904_ /*25981*/;
assign _42908_ = _42106_ ^ _42904_ /*25984*/;
assign _42909_ = _42900_ & _42908_ /*25982*/;
assign _42554_ = _42900_ ^ _42908_ /*25983*/;
assign _42906_ = _42907_ | _42909_ /*25980*/;
assign _42911_ = ~Q[16] /*25979*/;
assign _42910_ = _42911_ & D[58] /*25978*/;
assign _42913_ = _42107_ & _42910_ /*25973*/;
assign _42914_ = _42107_ ^ _42910_ /*25976*/;
assign _42915_ = _42906_ & _42914_ /*25974*/;
assign _42555_ = _42906_ ^ _42914_ /*25975*/;
assign _42912_ = _42913_ | _42915_ /*25972*/;
assign _42917_ = ~Q[16] /*25971*/;
assign _42916_ = _42917_ & D[59] /*25970*/;
assign _42919_ = _42108_ & _42916_ /*25965*/;
assign _42920_ = _42108_ ^ _42916_ /*25968*/;
assign _42921_ = _42912_ & _42920_ /*25966*/;
assign _42556_ = _42912_ ^ _42920_ /*25967*/;
assign _42918_ = _42919_ | _42921_ /*25964*/;
assign _42923_ = ~Q[16] /*25963*/;
assign _42922_ = _42923_ & D[60] /*25962*/;
assign _42925_ = _42109_ & _42922_ /*25957*/;
assign _42926_ = _42109_ ^ _42922_ /*25960*/;
assign _42927_ = _42918_ & _42926_ /*25958*/;
assign _42557_ = _42918_ ^ _42926_ /*25959*/;
assign _42924_ = _42925_ | _42927_ /*25956*/;
assign _42929_ = ~Q[16] /*25955*/;
assign _42928_ = _42929_ & D[61] /*25954*/;
assign _42931_ = _42110_ & _42928_ /*25949*/;
assign _42932_ = _42110_ ^ _42928_ /*25952*/;
assign _42933_ = _42924_ & _42932_ /*25950*/;
assign _42558_ = _42924_ ^ _42932_ /*25951*/;
assign _42930_ = _42931_ | _42933_ /*25948*/;
assign _42935_ = ~Q[16] /*25947*/;
assign _42934_ = _42935_ & D[62] /*25946*/;
assign _42937_ = _42111_ & _42934_ /*25941*/;
assign _42938_ = _42111_ ^ _42934_ /*25944*/;
assign _42939_ = _42930_ & _42938_ /*25942*/;
assign _42559_ = _42930_ ^ _42938_ /*25943*/;
assign _42936_ = _42937_ | _42939_ /*25940*/;
assign _42941_ = ~Q[16] /*25939*/;
assign _42940_ = _42941_ & zeroWire /*25938*/;
assign _42942_ = _42112_ ^ _42940_ /*25936*/;
assign _42560_ = _42942_ ^ _42936_ /*25935*/;
assign _43013_ = ~D[0] /*25681*/;
assign _43010_ = R_0[15] & _43013_ /*25677*/;
assign _43011_ = R_0[15] ^ _43013_ /*25680*/;
assign _43012_ = oneWire & _43011_ /*25678*/;
assign _42945_ = oneWire ^ _43011_ /*25679*/;
assign _43009_ = _43010_ | _43012_ /*25676*/;
assign _43018_ = ~D[1] /*25675*/;
assign _43015_ = _42497_ & _43018_ /*25671*/;
assign _43016_ = _42497_ ^ _43018_ /*25674*/;
assign _43017_ = _43009_ & _43016_ /*25672*/;
assign _42946_ = _43009_ ^ _43016_ /*25673*/;
assign _43014_ = _43015_ | _43017_ /*25670*/;
assign _43023_ = ~D[2] /*25669*/;
assign _43020_ = _42498_ & _43023_ /*25665*/;
assign _43021_ = _42498_ ^ _43023_ /*25668*/;
assign _43022_ = _43014_ & _43021_ /*25666*/;
assign _42947_ = _43014_ ^ _43021_ /*25667*/;
assign _43019_ = _43020_ | _43022_ /*25664*/;
assign _43028_ = ~D[3] /*25663*/;
assign _43025_ = _42499_ & _43028_ /*25659*/;
assign _43026_ = _42499_ ^ _43028_ /*25662*/;
assign _43027_ = _43019_ & _43026_ /*25660*/;
assign _42948_ = _43019_ ^ _43026_ /*25661*/;
assign _43024_ = _43025_ | _43027_ /*25658*/;
assign _43033_ = ~D[4] /*25657*/;
assign _43030_ = _42500_ & _43033_ /*25653*/;
assign _43031_ = _42500_ ^ _43033_ /*25656*/;
assign _43032_ = _43024_ & _43031_ /*25654*/;
assign _42949_ = _43024_ ^ _43031_ /*25655*/;
assign _43029_ = _43030_ | _43032_ /*25652*/;
assign _43038_ = ~D[5] /*25651*/;
assign _43035_ = _42501_ & _43038_ /*25647*/;
assign _43036_ = _42501_ ^ _43038_ /*25650*/;
assign _43037_ = _43029_ & _43036_ /*25648*/;
assign _42950_ = _43029_ ^ _43036_ /*25649*/;
assign _43034_ = _43035_ | _43037_ /*25646*/;
assign _43043_ = ~D[6] /*25645*/;
assign _43040_ = _42502_ & _43043_ /*25641*/;
assign _43041_ = _42502_ ^ _43043_ /*25644*/;
assign _43042_ = _43034_ & _43041_ /*25642*/;
assign _42951_ = _43034_ ^ _43041_ /*25643*/;
assign _43039_ = _43040_ | _43042_ /*25640*/;
assign _43048_ = ~D[7] /*25639*/;
assign _43045_ = _42503_ & _43048_ /*25635*/;
assign _43046_ = _42503_ ^ _43048_ /*25638*/;
assign _43047_ = _43039_ & _43046_ /*25636*/;
assign _42952_ = _43039_ ^ _43046_ /*25637*/;
assign _43044_ = _43045_ | _43047_ /*25634*/;
assign _43053_ = ~D[8] /*25633*/;
assign _43050_ = _42504_ & _43053_ /*25629*/;
assign _43051_ = _42504_ ^ _43053_ /*25632*/;
assign _43052_ = _43044_ & _43051_ /*25630*/;
assign _42953_ = _43044_ ^ _43051_ /*25631*/;
assign _43049_ = _43050_ | _43052_ /*25628*/;
assign _43058_ = ~D[9] /*25627*/;
assign _43055_ = _42505_ & _43058_ /*25623*/;
assign _43056_ = _42505_ ^ _43058_ /*25626*/;
assign _43057_ = _43049_ & _43056_ /*25624*/;
assign _42954_ = _43049_ ^ _43056_ /*25625*/;
assign _43054_ = _43055_ | _43057_ /*25622*/;
assign _43063_ = ~D[10] /*25621*/;
assign _43060_ = _42506_ & _43063_ /*25617*/;
assign _43061_ = _42506_ ^ _43063_ /*25620*/;
assign _43062_ = _43054_ & _43061_ /*25618*/;
assign _42955_ = _43054_ ^ _43061_ /*25619*/;
assign _43059_ = _43060_ | _43062_ /*25616*/;
assign _43068_ = ~D[11] /*25615*/;
assign _43065_ = _42507_ & _43068_ /*25611*/;
assign _43066_ = _42507_ ^ _43068_ /*25614*/;
assign _43067_ = _43059_ & _43066_ /*25612*/;
assign _42956_ = _43059_ ^ _43066_ /*25613*/;
assign _43064_ = _43065_ | _43067_ /*25610*/;
assign _43073_ = ~D[12] /*25609*/;
assign _43070_ = _42508_ & _43073_ /*25605*/;
assign _43071_ = _42508_ ^ _43073_ /*25608*/;
assign _43072_ = _43064_ & _43071_ /*25606*/;
assign _42957_ = _43064_ ^ _43071_ /*25607*/;
assign _43069_ = _43070_ | _43072_ /*25604*/;
assign _43078_ = ~D[13] /*25603*/;
assign _43075_ = _42509_ & _43078_ /*25599*/;
assign _43076_ = _42509_ ^ _43078_ /*25602*/;
assign _43077_ = _43069_ & _43076_ /*25600*/;
assign _42958_ = _43069_ ^ _43076_ /*25601*/;
assign _43074_ = _43075_ | _43077_ /*25598*/;
assign _43083_ = ~D[14] /*25597*/;
assign _43080_ = _42510_ & _43083_ /*25593*/;
assign _43081_ = _42510_ ^ _43083_ /*25596*/;
assign _43082_ = _43074_ & _43081_ /*25594*/;
assign _42959_ = _43074_ ^ _43081_ /*25595*/;
assign _43079_ = _43080_ | _43082_ /*25592*/;
assign _43088_ = ~D[15] /*25591*/;
assign _43085_ = _42511_ & _43088_ /*25587*/;
assign _43086_ = _42511_ ^ _43088_ /*25590*/;
assign _43087_ = _43079_ & _43086_ /*25588*/;
assign _42960_ = _43079_ ^ _43086_ /*25589*/;
assign _43084_ = _43085_ | _43087_ /*25586*/;
assign _43093_ = ~D[16] /*25585*/;
assign _43090_ = _42512_ & _43093_ /*25581*/;
assign _43091_ = _42512_ ^ _43093_ /*25584*/;
assign _43092_ = _43084_ & _43091_ /*25582*/;
assign _42961_ = _43084_ ^ _43091_ /*25583*/;
assign _43089_ = _43090_ | _43092_ /*25580*/;
assign _43098_ = ~D[17] /*25579*/;
assign _43095_ = _42513_ & _43098_ /*25575*/;
assign _43096_ = _42513_ ^ _43098_ /*25578*/;
assign _43097_ = _43089_ & _43096_ /*25576*/;
assign _42962_ = _43089_ ^ _43096_ /*25577*/;
assign _43094_ = _43095_ | _43097_ /*25574*/;
assign _43103_ = ~D[18] /*25573*/;
assign _43100_ = _42514_ & _43103_ /*25569*/;
assign _43101_ = _42514_ ^ _43103_ /*25572*/;
assign _43102_ = _43094_ & _43101_ /*25570*/;
assign _42963_ = _43094_ ^ _43101_ /*25571*/;
assign _43099_ = _43100_ | _43102_ /*25568*/;
assign _43108_ = ~D[19] /*25567*/;
assign _43105_ = _42515_ & _43108_ /*25563*/;
assign _43106_ = _42515_ ^ _43108_ /*25566*/;
assign _43107_ = _43099_ & _43106_ /*25564*/;
assign _42964_ = _43099_ ^ _43106_ /*25565*/;
assign _43104_ = _43105_ | _43107_ /*25562*/;
assign _43113_ = ~D[20] /*25561*/;
assign _43110_ = _42516_ & _43113_ /*25557*/;
assign _43111_ = _42516_ ^ _43113_ /*25560*/;
assign _43112_ = _43104_ & _43111_ /*25558*/;
assign _42965_ = _43104_ ^ _43111_ /*25559*/;
assign _43109_ = _43110_ | _43112_ /*25556*/;
assign _43118_ = ~D[21] /*25555*/;
assign _43115_ = _42517_ & _43118_ /*25551*/;
assign _43116_ = _42517_ ^ _43118_ /*25554*/;
assign _43117_ = _43109_ & _43116_ /*25552*/;
assign _42966_ = _43109_ ^ _43116_ /*25553*/;
assign _43114_ = _43115_ | _43117_ /*25550*/;
assign _43123_ = ~D[22] /*25549*/;
assign _43120_ = _42518_ & _43123_ /*25545*/;
assign _43121_ = _42518_ ^ _43123_ /*25548*/;
assign _43122_ = _43114_ & _43121_ /*25546*/;
assign _42967_ = _43114_ ^ _43121_ /*25547*/;
assign _43119_ = _43120_ | _43122_ /*25544*/;
assign _43128_ = ~D[23] /*25543*/;
assign _43125_ = _42519_ & _43128_ /*25539*/;
assign _43126_ = _42519_ ^ _43128_ /*25542*/;
assign _43127_ = _43119_ & _43126_ /*25540*/;
assign _42968_ = _43119_ ^ _43126_ /*25541*/;
assign _43124_ = _43125_ | _43127_ /*25538*/;
assign _43133_ = ~D[24] /*25537*/;
assign _43130_ = _42520_ & _43133_ /*25533*/;
assign _43131_ = _42520_ ^ _43133_ /*25536*/;
assign _43132_ = _43124_ & _43131_ /*25534*/;
assign _42969_ = _43124_ ^ _43131_ /*25535*/;
assign _43129_ = _43130_ | _43132_ /*25532*/;
assign _43138_ = ~D[25] /*25531*/;
assign _43135_ = _42521_ & _43138_ /*25527*/;
assign _43136_ = _42521_ ^ _43138_ /*25530*/;
assign _43137_ = _43129_ & _43136_ /*25528*/;
assign _42970_ = _43129_ ^ _43136_ /*25529*/;
assign _43134_ = _43135_ | _43137_ /*25526*/;
assign _43143_ = ~D[26] /*25525*/;
assign _43140_ = _42522_ & _43143_ /*25521*/;
assign _43141_ = _42522_ ^ _43143_ /*25524*/;
assign _43142_ = _43134_ & _43141_ /*25522*/;
assign _42971_ = _43134_ ^ _43141_ /*25523*/;
assign _43139_ = _43140_ | _43142_ /*25520*/;
assign _43148_ = ~D[27] /*25519*/;
assign _43145_ = _42523_ & _43148_ /*25515*/;
assign _43146_ = _42523_ ^ _43148_ /*25518*/;
assign _43147_ = _43139_ & _43146_ /*25516*/;
assign _42972_ = _43139_ ^ _43146_ /*25517*/;
assign _43144_ = _43145_ | _43147_ /*25514*/;
assign _43153_ = ~D[28] /*25513*/;
assign _43150_ = _42524_ & _43153_ /*25509*/;
assign _43151_ = _42524_ ^ _43153_ /*25512*/;
assign _43152_ = _43144_ & _43151_ /*25510*/;
assign _42973_ = _43144_ ^ _43151_ /*25511*/;
assign _43149_ = _43150_ | _43152_ /*25508*/;
assign _43158_ = ~D[29] /*25507*/;
assign _43155_ = _42525_ & _43158_ /*25503*/;
assign _43156_ = _42525_ ^ _43158_ /*25506*/;
assign _43157_ = _43149_ & _43156_ /*25504*/;
assign _42974_ = _43149_ ^ _43156_ /*25505*/;
assign _43154_ = _43155_ | _43157_ /*25502*/;
assign _43163_ = ~D[30] /*25501*/;
assign _43160_ = _42526_ & _43163_ /*25497*/;
assign _43161_ = _42526_ ^ _43163_ /*25500*/;
assign _43162_ = _43154_ & _43161_ /*25498*/;
assign _42975_ = _43154_ ^ _43161_ /*25499*/;
assign _43159_ = _43160_ | _43162_ /*25496*/;
assign _43168_ = ~D[31] /*25495*/;
assign _43165_ = _42527_ & _43168_ /*25491*/;
assign _43166_ = _42527_ ^ _43168_ /*25494*/;
assign _43167_ = _43159_ & _43166_ /*25492*/;
assign _42976_ = _43159_ ^ _43166_ /*25493*/;
assign _43164_ = _43165_ | _43167_ /*25490*/;
assign _43173_ = ~D[32] /*25489*/;
assign _43170_ = _42528_ & _43173_ /*25485*/;
assign _43171_ = _42528_ ^ _43173_ /*25488*/;
assign _43172_ = _43164_ & _43171_ /*25486*/;
assign _42977_ = _43164_ ^ _43171_ /*25487*/;
assign _43169_ = _43170_ | _43172_ /*25484*/;
assign _43178_ = ~D[33] /*25483*/;
assign _43175_ = _42529_ & _43178_ /*25479*/;
assign _43176_ = _42529_ ^ _43178_ /*25482*/;
assign _43177_ = _43169_ & _43176_ /*25480*/;
assign _42978_ = _43169_ ^ _43176_ /*25481*/;
assign _43174_ = _43175_ | _43177_ /*25478*/;
assign _43183_ = ~D[34] /*25477*/;
assign _43180_ = _42530_ & _43183_ /*25473*/;
assign _43181_ = _42530_ ^ _43183_ /*25476*/;
assign _43182_ = _43174_ & _43181_ /*25474*/;
assign _42979_ = _43174_ ^ _43181_ /*25475*/;
assign _43179_ = _43180_ | _43182_ /*25472*/;
assign _43188_ = ~D[35] /*25471*/;
assign _43185_ = _42531_ & _43188_ /*25467*/;
assign _43186_ = _42531_ ^ _43188_ /*25470*/;
assign _43187_ = _43179_ & _43186_ /*25468*/;
assign _42980_ = _43179_ ^ _43186_ /*25469*/;
assign _43184_ = _43185_ | _43187_ /*25466*/;
assign _43193_ = ~D[36] /*25465*/;
assign _43190_ = _42532_ & _43193_ /*25461*/;
assign _43191_ = _42532_ ^ _43193_ /*25464*/;
assign _43192_ = _43184_ & _43191_ /*25462*/;
assign _42981_ = _43184_ ^ _43191_ /*25463*/;
assign _43189_ = _43190_ | _43192_ /*25460*/;
assign _43198_ = ~D[37] /*25459*/;
assign _43195_ = _42533_ & _43198_ /*25455*/;
assign _43196_ = _42533_ ^ _43198_ /*25458*/;
assign _43197_ = _43189_ & _43196_ /*25456*/;
assign _42982_ = _43189_ ^ _43196_ /*25457*/;
assign _43194_ = _43195_ | _43197_ /*25454*/;
assign _43203_ = ~D[38] /*25453*/;
assign _43200_ = _42534_ & _43203_ /*25449*/;
assign _43201_ = _42534_ ^ _43203_ /*25452*/;
assign _43202_ = _43194_ & _43201_ /*25450*/;
assign _42983_ = _43194_ ^ _43201_ /*25451*/;
assign _43199_ = _43200_ | _43202_ /*25448*/;
assign _43208_ = ~D[39] /*25447*/;
assign _43205_ = _42535_ & _43208_ /*25443*/;
assign _43206_ = _42535_ ^ _43208_ /*25446*/;
assign _43207_ = _43199_ & _43206_ /*25444*/;
assign _42984_ = _43199_ ^ _43206_ /*25445*/;
assign _43204_ = _43205_ | _43207_ /*25442*/;
assign _43213_ = ~D[40] /*25441*/;
assign _43210_ = _42536_ & _43213_ /*25437*/;
assign _43211_ = _42536_ ^ _43213_ /*25440*/;
assign _43212_ = _43204_ & _43211_ /*25438*/;
assign _42985_ = _43204_ ^ _43211_ /*25439*/;
assign _43209_ = _43210_ | _43212_ /*25436*/;
assign _43218_ = ~D[41] /*25435*/;
assign _43215_ = _42537_ & _43218_ /*25431*/;
assign _43216_ = _42537_ ^ _43218_ /*25434*/;
assign _43217_ = _43209_ & _43216_ /*25432*/;
assign _42986_ = _43209_ ^ _43216_ /*25433*/;
assign _43214_ = _43215_ | _43217_ /*25430*/;
assign _43223_ = ~D[42] /*25429*/;
assign _43220_ = _42538_ & _43223_ /*25425*/;
assign _43221_ = _42538_ ^ _43223_ /*25428*/;
assign _43222_ = _43214_ & _43221_ /*25426*/;
assign _42987_ = _43214_ ^ _43221_ /*25427*/;
assign _43219_ = _43220_ | _43222_ /*25424*/;
assign _43228_ = ~D[43] /*25423*/;
assign _43225_ = _42539_ & _43228_ /*25419*/;
assign _43226_ = _42539_ ^ _43228_ /*25422*/;
assign _43227_ = _43219_ & _43226_ /*25420*/;
assign _42988_ = _43219_ ^ _43226_ /*25421*/;
assign _43224_ = _43225_ | _43227_ /*25418*/;
assign _43233_ = ~D[44] /*25417*/;
assign _43230_ = _42540_ & _43233_ /*25413*/;
assign _43231_ = _42540_ ^ _43233_ /*25416*/;
assign _43232_ = _43224_ & _43231_ /*25414*/;
assign _42989_ = _43224_ ^ _43231_ /*25415*/;
assign _43229_ = _43230_ | _43232_ /*25412*/;
assign _43238_ = ~D[45] /*25411*/;
assign _43235_ = _42541_ & _43238_ /*25407*/;
assign _43236_ = _42541_ ^ _43238_ /*25410*/;
assign _43237_ = _43229_ & _43236_ /*25408*/;
assign _42990_ = _43229_ ^ _43236_ /*25409*/;
assign _43234_ = _43235_ | _43237_ /*25406*/;
assign _43243_ = ~D[46] /*25405*/;
assign _43240_ = _42542_ & _43243_ /*25401*/;
assign _43241_ = _42542_ ^ _43243_ /*25404*/;
assign _43242_ = _43234_ & _43241_ /*25402*/;
assign _42991_ = _43234_ ^ _43241_ /*25403*/;
assign _43239_ = _43240_ | _43242_ /*25400*/;
assign _43248_ = ~D[47] /*25399*/;
assign _43245_ = _42543_ & _43248_ /*25395*/;
assign _43246_ = _42543_ ^ _43248_ /*25398*/;
assign _43247_ = _43239_ & _43246_ /*25396*/;
assign _42992_ = _43239_ ^ _43246_ /*25397*/;
assign _43244_ = _43245_ | _43247_ /*25394*/;
assign _43253_ = ~D[48] /*25393*/;
assign _43250_ = _42544_ & _43253_ /*25389*/;
assign _43251_ = _42544_ ^ _43253_ /*25392*/;
assign _43252_ = _43244_ & _43251_ /*25390*/;
assign _42993_ = _43244_ ^ _43251_ /*25391*/;
assign _43249_ = _43250_ | _43252_ /*25388*/;
assign _43258_ = ~D[49] /*25387*/;
assign _43255_ = _42545_ & _43258_ /*25383*/;
assign _43256_ = _42545_ ^ _43258_ /*25386*/;
assign _43257_ = _43249_ & _43256_ /*25384*/;
assign _42994_ = _43249_ ^ _43256_ /*25385*/;
assign _43254_ = _43255_ | _43257_ /*25382*/;
assign _43263_ = ~D[50] /*25381*/;
assign _43260_ = _42546_ & _43263_ /*25377*/;
assign _43261_ = _42546_ ^ _43263_ /*25380*/;
assign _43262_ = _43254_ & _43261_ /*25378*/;
assign _42995_ = _43254_ ^ _43261_ /*25379*/;
assign _43259_ = _43260_ | _43262_ /*25376*/;
assign _43268_ = ~D[51] /*25375*/;
assign _43265_ = _42547_ & _43268_ /*25371*/;
assign _43266_ = _42547_ ^ _43268_ /*25374*/;
assign _43267_ = _43259_ & _43266_ /*25372*/;
assign _42996_ = _43259_ ^ _43266_ /*25373*/;
assign _43264_ = _43265_ | _43267_ /*25370*/;
assign _43273_ = ~D[52] /*25369*/;
assign _43270_ = _42548_ & _43273_ /*25365*/;
assign _43271_ = _42548_ ^ _43273_ /*25368*/;
assign _43272_ = _43264_ & _43271_ /*25366*/;
assign _42997_ = _43264_ ^ _43271_ /*25367*/;
assign _43269_ = _43270_ | _43272_ /*25364*/;
assign _43278_ = ~D[53] /*25363*/;
assign _43275_ = _42549_ & _43278_ /*25359*/;
assign _43276_ = _42549_ ^ _43278_ /*25362*/;
assign _43277_ = _43269_ & _43276_ /*25360*/;
assign _42998_ = _43269_ ^ _43276_ /*25361*/;
assign _43274_ = _43275_ | _43277_ /*25358*/;
assign _43283_ = ~D[54] /*25357*/;
assign _43280_ = _42550_ & _43283_ /*25353*/;
assign _43281_ = _42550_ ^ _43283_ /*25356*/;
assign _43282_ = _43274_ & _43281_ /*25354*/;
assign _42999_ = _43274_ ^ _43281_ /*25355*/;
assign _43279_ = _43280_ | _43282_ /*25352*/;
assign _43288_ = ~D[55] /*25351*/;
assign _43285_ = _42551_ & _43288_ /*25347*/;
assign _43286_ = _42551_ ^ _43288_ /*25350*/;
assign _43287_ = _43279_ & _43286_ /*25348*/;
assign _43000_ = _43279_ ^ _43286_ /*25349*/;
assign _43284_ = _43285_ | _43287_ /*25346*/;
assign _43293_ = ~D[56] /*25345*/;
assign _43290_ = _42552_ & _43293_ /*25341*/;
assign _43291_ = _42552_ ^ _43293_ /*25344*/;
assign _43292_ = _43284_ & _43291_ /*25342*/;
assign _43001_ = _43284_ ^ _43291_ /*25343*/;
assign _43289_ = _43290_ | _43292_ /*25340*/;
assign _43298_ = ~D[57] /*25339*/;
assign _43295_ = _42553_ & _43298_ /*25335*/;
assign _43296_ = _42553_ ^ _43298_ /*25338*/;
assign _43297_ = _43289_ & _43296_ /*25336*/;
assign _43002_ = _43289_ ^ _43296_ /*25337*/;
assign _43294_ = _43295_ | _43297_ /*25334*/;
assign _43303_ = ~D[58] /*25333*/;
assign _43300_ = _42554_ & _43303_ /*25329*/;
assign _43301_ = _42554_ ^ _43303_ /*25332*/;
assign _43302_ = _43294_ & _43301_ /*25330*/;
assign _43003_ = _43294_ ^ _43301_ /*25331*/;
assign _43299_ = _43300_ | _43302_ /*25328*/;
assign _43308_ = ~D[59] /*25327*/;
assign _43305_ = _42555_ & _43308_ /*25323*/;
assign _43306_ = _42555_ ^ _43308_ /*25326*/;
assign _43307_ = _43299_ & _43306_ /*25324*/;
assign _43004_ = _43299_ ^ _43306_ /*25325*/;
assign _43304_ = _43305_ | _43307_ /*25322*/;
assign _43313_ = ~D[60] /*25321*/;
assign _43310_ = _42556_ & _43313_ /*25317*/;
assign _43311_ = _42556_ ^ _43313_ /*25320*/;
assign _43312_ = _43304_ & _43311_ /*25318*/;
assign _43005_ = _43304_ ^ _43311_ /*25319*/;
assign _43309_ = _43310_ | _43312_ /*25316*/;
assign _43318_ = ~D[61] /*25315*/;
assign _43315_ = _42557_ & _43318_ /*25311*/;
assign _43316_ = _42557_ ^ _43318_ /*25314*/;
assign _43317_ = _43309_ & _43316_ /*25312*/;
assign _43006_ = _43309_ ^ _43316_ /*25313*/;
assign _43314_ = _43315_ | _43317_ /*25310*/;
assign _43323_ = ~D[62] /*25309*/;
assign _43320_ = _42558_ & _43323_ /*25305*/;
assign _43321_ = _42558_ ^ _43323_ /*25308*/;
assign _43322_ = _43314_ & _43321_ /*25306*/;
assign _43007_ = _43314_ ^ _43321_ /*25307*/;
assign _43319_ = _43320_ | _43322_ /*25304*/;
assign _43324_ = _42559_ & oneWire /*25299*/;
assign _43325_ = _42559_ ^ oneWire /*25302*/;
assign _43326_ = _43319_ & _43325_ /*25300*/;
assign _43008_ = _43319_ ^ _43325_ /*25301*/;
assign Q[15] = _43324_ | _43326_ /*25298*/;
assign _43459_ = ~Q[15] /*24913*/;
assign _43458_ = _43459_ & D[0] /*24912*/;
assign _43461_ = _42945_ & _43458_ /*24907*/;
assign _43462_ = _42945_ ^ _43458_ /*24910*/;
assign _43463_ = zeroWire & _43462_ /*24908*/;
assign _43393_ = zeroWire ^ _43462_ /*24909*/;
assign _43460_ = _43461_ | _43463_ /*24906*/;
assign _43465_ = ~Q[15] /*24905*/;
assign _43464_ = _43465_ & D[1] /*24904*/;
assign _43467_ = _42946_ & _43464_ /*24899*/;
assign _43468_ = _42946_ ^ _43464_ /*24902*/;
assign _43469_ = _43460_ & _43468_ /*24900*/;
assign _43394_ = _43460_ ^ _43468_ /*24901*/;
assign _43466_ = _43467_ | _43469_ /*24898*/;
assign _43471_ = ~Q[15] /*24897*/;
assign _43470_ = _43471_ & D[2] /*24896*/;
assign _43473_ = _42947_ & _43470_ /*24891*/;
assign _43474_ = _42947_ ^ _43470_ /*24894*/;
assign _43475_ = _43466_ & _43474_ /*24892*/;
assign _43395_ = _43466_ ^ _43474_ /*24893*/;
assign _43472_ = _43473_ | _43475_ /*24890*/;
assign _43477_ = ~Q[15] /*24889*/;
assign _43476_ = _43477_ & D[3] /*24888*/;
assign _43479_ = _42948_ & _43476_ /*24883*/;
assign _43480_ = _42948_ ^ _43476_ /*24886*/;
assign _43481_ = _43472_ & _43480_ /*24884*/;
assign _43396_ = _43472_ ^ _43480_ /*24885*/;
assign _43478_ = _43479_ | _43481_ /*24882*/;
assign _43483_ = ~Q[15] /*24881*/;
assign _43482_ = _43483_ & D[4] /*24880*/;
assign _43485_ = _42949_ & _43482_ /*24875*/;
assign _43486_ = _42949_ ^ _43482_ /*24878*/;
assign _43487_ = _43478_ & _43486_ /*24876*/;
assign _43397_ = _43478_ ^ _43486_ /*24877*/;
assign _43484_ = _43485_ | _43487_ /*24874*/;
assign _43489_ = ~Q[15] /*24873*/;
assign _43488_ = _43489_ & D[5] /*24872*/;
assign _43491_ = _42950_ & _43488_ /*24867*/;
assign _43492_ = _42950_ ^ _43488_ /*24870*/;
assign _43493_ = _43484_ & _43492_ /*24868*/;
assign _43398_ = _43484_ ^ _43492_ /*24869*/;
assign _43490_ = _43491_ | _43493_ /*24866*/;
assign _43495_ = ~Q[15] /*24865*/;
assign _43494_ = _43495_ & D[6] /*24864*/;
assign _43497_ = _42951_ & _43494_ /*24859*/;
assign _43498_ = _42951_ ^ _43494_ /*24862*/;
assign _43499_ = _43490_ & _43498_ /*24860*/;
assign _43399_ = _43490_ ^ _43498_ /*24861*/;
assign _43496_ = _43497_ | _43499_ /*24858*/;
assign _43501_ = ~Q[15] /*24857*/;
assign _43500_ = _43501_ & D[7] /*24856*/;
assign _43503_ = _42952_ & _43500_ /*24851*/;
assign _43504_ = _42952_ ^ _43500_ /*24854*/;
assign _43505_ = _43496_ & _43504_ /*24852*/;
assign _43400_ = _43496_ ^ _43504_ /*24853*/;
assign _43502_ = _43503_ | _43505_ /*24850*/;
assign _43507_ = ~Q[15] /*24849*/;
assign _43506_ = _43507_ & D[8] /*24848*/;
assign _43509_ = _42953_ & _43506_ /*24843*/;
assign _43510_ = _42953_ ^ _43506_ /*24846*/;
assign _43511_ = _43502_ & _43510_ /*24844*/;
assign _43401_ = _43502_ ^ _43510_ /*24845*/;
assign _43508_ = _43509_ | _43511_ /*24842*/;
assign _43513_ = ~Q[15] /*24841*/;
assign _43512_ = _43513_ & D[9] /*24840*/;
assign _43515_ = _42954_ & _43512_ /*24835*/;
assign _43516_ = _42954_ ^ _43512_ /*24838*/;
assign _43517_ = _43508_ & _43516_ /*24836*/;
assign _43402_ = _43508_ ^ _43516_ /*24837*/;
assign _43514_ = _43515_ | _43517_ /*24834*/;
assign _43519_ = ~Q[15] /*24833*/;
assign _43518_ = _43519_ & D[10] /*24832*/;
assign _43521_ = _42955_ & _43518_ /*24827*/;
assign _43522_ = _42955_ ^ _43518_ /*24830*/;
assign _43523_ = _43514_ & _43522_ /*24828*/;
assign _43403_ = _43514_ ^ _43522_ /*24829*/;
assign _43520_ = _43521_ | _43523_ /*24826*/;
assign _43525_ = ~Q[15] /*24825*/;
assign _43524_ = _43525_ & D[11] /*24824*/;
assign _43527_ = _42956_ & _43524_ /*24819*/;
assign _43528_ = _42956_ ^ _43524_ /*24822*/;
assign _43529_ = _43520_ & _43528_ /*24820*/;
assign _43404_ = _43520_ ^ _43528_ /*24821*/;
assign _43526_ = _43527_ | _43529_ /*24818*/;
assign _43531_ = ~Q[15] /*24817*/;
assign _43530_ = _43531_ & D[12] /*24816*/;
assign _43533_ = _42957_ & _43530_ /*24811*/;
assign _43534_ = _42957_ ^ _43530_ /*24814*/;
assign _43535_ = _43526_ & _43534_ /*24812*/;
assign _43405_ = _43526_ ^ _43534_ /*24813*/;
assign _43532_ = _43533_ | _43535_ /*24810*/;
assign _43537_ = ~Q[15] /*24809*/;
assign _43536_ = _43537_ & D[13] /*24808*/;
assign _43539_ = _42958_ & _43536_ /*24803*/;
assign _43540_ = _42958_ ^ _43536_ /*24806*/;
assign _43541_ = _43532_ & _43540_ /*24804*/;
assign _43406_ = _43532_ ^ _43540_ /*24805*/;
assign _43538_ = _43539_ | _43541_ /*24802*/;
assign _43543_ = ~Q[15] /*24801*/;
assign _43542_ = _43543_ & D[14] /*24800*/;
assign _43545_ = _42959_ & _43542_ /*24795*/;
assign _43546_ = _42959_ ^ _43542_ /*24798*/;
assign _43547_ = _43538_ & _43546_ /*24796*/;
assign _43407_ = _43538_ ^ _43546_ /*24797*/;
assign _43544_ = _43545_ | _43547_ /*24794*/;
assign _43549_ = ~Q[15] /*24793*/;
assign _43548_ = _43549_ & D[15] /*24792*/;
assign _43551_ = _42960_ & _43548_ /*24787*/;
assign _43552_ = _42960_ ^ _43548_ /*24790*/;
assign _43553_ = _43544_ & _43552_ /*24788*/;
assign _43408_ = _43544_ ^ _43552_ /*24789*/;
assign _43550_ = _43551_ | _43553_ /*24786*/;
assign _43555_ = ~Q[15] /*24785*/;
assign _43554_ = _43555_ & D[16] /*24784*/;
assign _43557_ = _42961_ & _43554_ /*24779*/;
assign _43558_ = _42961_ ^ _43554_ /*24782*/;
assign _43559_ = _43550_ & _43558_ /*24780*/;
assign _43409_ = _43550_ ^ _43558_ /*24781*/;
assign _43556_ = _43557_ | _43559_ /*24778*/;
assign _43561_ = ~Q[15] /*24777*/;
assign _43560_ = _43561_ & D[17] /*24776*/;
assign _43563_ = _42962_ & _43560_ /*24771*/;
assign _43564_ = _42962_ ^ _43560_ /*24774*/;
assign _43565_ = _43556_ & _43564_ /*24772*/;
assign _43410_ = _43556_ ^ _43564_ /*24773*/;
assign _43562_ = _43563_ | _43565_ /*24770*/;
assign _43567_ = ~Q[15] /*24769*/;
assign _43566_ = _43567_ & D[18] /*24768*/;
assign _43569_ = _42963_ & _43566_ /*24763*/;
assign _43570_ = _42963_ ^ _43566_ /*24766*/;
assign _43571_ = _43562_ & _43570_ /*24764*/;
assign _43411_ = _43562_ ^ _43570_ /*24765*/;
assign _43568_ = _43569_ | _43571_ /*24762*/;
assign _43573_ = ~Q[15] /*24761*/;
assign _43572_ = _43573_ & D[19] /*24760*/;
assign _43575_ = _42964_ & _43572_ /*24755*/;
assign _43576_ = _42964_ ^ _43572_ /*24758*/;
assign _43577_ = _43568_ & _43576_ /*24756*/;
assign _43412_ = _43568_ ^ _43576_ /*24757*/;
assign _43574_ = _43575_ | _43577_ /*24754*/;
assign _43579_ = ~Q[15] /*24753*/;
assign _43578_ = _43579_ & D[20] /*24752*/;
assign _43581_ = _42965_ & _43578_ /*24747*/;
assign _43582_ = _42965_ ^ _43578_ /*24750*/;
assign _43583_ = _43574_ & _43582_ /*24748*/;
assign _43413_ = _43574_ ^ _43582_ /*24749*/;
assign _43580_ = _43581_ | _43583_ /*24746*/;
assign _43585_ = ~Q[15] /*24745*/;
assign _43584_ = _43585_ & D[21] /*24744*/;
assign _43587_ = _42966_ & _43584_ /*24739*/;
assign _43588_ = _42966_ ^ _43584_ /*24742*/;
assign _43589_ = _43580_ & _43588_ /*24740*/;
assign _43414_ = _43580_ ^ _43588_ /*24741*/;
assign _43586_ = _43587_ | _43589_ /*24738*/;
assign _43591_ = ~Q[15] /*24737*/;
assign _43590_ = _43591_ & D[22] /*24736*/;
assign _43593_ = _42967_ & _43590_ /*24731*/;
assign _43594_ = _42967_ ^ _43590_ /*24734*/;
assign _43595_ = _43586_ & _43594_ /*24732*/;
assign _43415_ = _43586_ ^ _43594_ /*24733*/;
assign _43592_ = _43593_ | _43595_ /*24730*/;
assign _43597_ = ~Q[15] /*24729*/;
assign _43596_ = _43597_ & D[23] /*24728*/;
assign _43599_ = _42968_ & _43596_ /*24723*/;
assign _43600_ = _42968_ ^ _43596_ /*24726*/;
assign _43601_ = _43592_ & _43600_ /*24724*/;
assign _43416_ = _43592_ ^ _43600_ /*24725*/;
assign _43598_ = _43599_ | _43601_ /*24722*/;
assign _43603_ = ~Q[15] /*24721*/;
assign _43602_ = _43603_ & D[24] /*24720*/;
assign _43605_ = _42969_ & _43602_ /*24715*/;
assign _43606_ = _42969_ ^ _43602_ /*24718*/;
assign _43607_ = _43598_ & _43606_ /*24716*/;
assign _43417_ = _43598_ ^ _43606_ /*24717*/;
assign _43604_ = _43605_ | _43607_ /*24714*/;
assign _43609_ = ~Q[15] /*24713*/;
assign _43608_ = _43609_ & D[25] /*24712*/;
assign _43611_ = _42970_ & _43608_ /*24707*/;
assign _43612_ = _42970_ ^ _43608_ /*24710*/;
assign _43613_ = _43604_ & _43612_ /*24708*/;
assign _43418_ = _43604_ ^ _43612_ /*24709*/;
assign _43610_ = _43611_ | _43613_ /*24706*/;
assign _43615_ = ~Q[15] /*24705*/;
assign _43614_ = _43615_ & D[26] /*24704*/;
assign _43617_ = _42971_ & _43614_ /*24699*/;
assign _43618_ = _42971_ ^ _43614_ /*24702*/;
assign _43619_ = _43610_ & _43618_ /*24700*/;
assign _43419_ = _43610_ ^ _43618_ /*24701*/;
assign _43616_ = _43617_ | _43619_ /*24698*/;
assign _43621_ = ~Q[15] /*24697*/;
assign _43620_ = _43621_ & D[27] /*24696*/;
assign _43623_ = _42972_ & _43620_ /*24691*/;
assign _43624_ = _42972_ ^ _43620_ /*24694*/;
assign _43625_ = _43616_ & _43624_ /*24692*/;
assign _43420_ = _43616_ ^ _43624_ /*24693*/;
assign _43622_ = _43623_ | _43625_ /*24690*/;
assign _43627_ = ~Q[15] /*24689*/;
assign _43626_ = _43627_ & D[28] /*24688*/;
assign _43629_ = _42973_ & _43626_ /*24683*/;
assign _43630_ = _42973_ ^ _43626_ /*24686*/;
assign _43631_ = _43622_ & _43630_ /*24684*/;
assign _43421_ = _43622_ ^ _43630_ /*24685*/;
assign _43628_ = _43629_ | _43631_ /*24682*/;
assign _43633_ = ~Q[15] /*24681*/;
assign _43632_ = _43633_ & D[29] /*24680*/;
assign _43635_ = _42974_ & _43632_ /*24675*/;
assign _43636_ = _42974_ ^ _43632_ /*24678*/;
assign _43637_ = _43628_ & _43636_ /*24676*/;
assign _43422_ = _43628_ ^ _43636_ /*24677*/;
assign _43634_ = _43635_ | _43637_ /*24674*/;
assign _43639_ = ~Q[15] /*24673*/;
assign _43638_ = _43639_ & D[30] /*24672*/;
assign _43641_ = _42975_ & _43638_ /*24667*/;
assign _43642_ = _42975_ ^ _43638_ /*24670*/;
assign _43643_ = _43634_ & _43642_ /*24668*/;
assign _43423_ = _43634_ ^ _43642_ /*24669*/;
assign _43640_ = _43641_ | _43643_ /*24666*/;
assign _43645_ = ~Q[15] /*24665*/;
assign _43644_ = _43645_ & D[31] /*24664*/;
assign _43647_ = _42976_ & _43644_ /*24659*/;
assign _43648_ = _42976_ ^ _43644_ /*24662*/;
assign _43649_ = _43640_ & _43648_ /*24660*/;
assign _43424_ = _43640_ ^ _43648_ /*24661*/;
assign _43646_ = _43647_ | _43649_ /*24658*/;
assign _43651_ = ~Q[15] /*24657*/;
assign _43650_ = _43651_ & D[32] /*24656*/;
assign _43653_ = _42977_ & _43650_ /*24651*/;
assign _43654_ = _42977_ ^ _43650_ /*24654*/;
assign _43655_ = _43646_ & _43654_ /*24652*/;
assign _43425_ = _43646_ ^ _43654_ /*24653*/;
assign _43652_ = _43653_ | _43655_ /*24650*/;
assign _43657_ = ~Q[15] /*24649*/;
assign _43656_ = _43657_ & D[33] /*24648*/;
assign _43659_ = _42978_ & _43656_ /*24643*/;
assign _43660_ = _42978_ ^ _43656_ /*24646*/;
assign _43661_ = _43652_ & _43660_ /*24644*/;
assign _43426_ = _43652_ ^ _43660_ /*24645*/;
assign _43658_ = _43659_ | _43661_ /*24642*/;
assign _43663_ = ~Q[15] /*24641*/;
assign _43662_ = _43663_ & D[34] /*24640*/;
assign _43665_ = _42979_ & _43662_ /*24635*/;
assign _43666_ = _42979_ ^ _43662_ /*24638*/;
assign _43667_ = _43658_ & _43666_ /*24636*/;
assign _43427_ = _43658_ ^ _43666_ /*24637*/;
assign _43664_ = _43665_ | _43667_ /*24634*/;
assign _43669_ = ~Q[15] /*24633*/;
assign _43668_ = _43669_ & D[35] /*24632*/;
assign _43671_ = _42980_ & _43668_ /*24627*/;
assign _43672_ = _42980_ ^ _43668_ /*24630*/;
assign _43673_ = _43664_ & _43672_ /*24628*/;
assign _43428_ = _43664_ ^ _43672_ /*24629*/;
assign _43670_ = _43671_ | _43673_ /*24626*/;
assign _43675_ = ~Q[15] /*24625*/;
assign _43674_ = _43675_ & D[36] /*24624*/;
assign _43677_ = _42981_ & _43674_ /*24619*/;
assign _43678_ = _42981_ ^ _43674_ /*24622*/;
assign _43679_ = _43670_ & _43678_ /*24620*/;
assign _43429_ = _43670_ ^ _43678_ /*24621*/;
assign _43676_ = _43677_ | _43679_ /*24618*/;
assign _43681_ = ~Q[15] /*24617*/;
assign _43680_ = _43681_ & D[37] /*24616*/;
assign _43683_ = _42982_ & _43680_ /*24611*/;
assign _43684_ = _42982_ ^ _43680_ /*24614*/;
assign _43685_ = _43676_ & _43684_ /*24612*/;
assign _43430_ = _43676_ ^ _43684_ /*24613*/;
assign _43682_ = _43683_ | _43685_ /*24610*/;
assign _43687_ = ~Q[15] /*24609*/;
assign _43686_ = _43687_ & D[38] /*24608*/;
assign _43689_ = _42983_ & _43686_ /*24603*/;
assign _43690_ = _42983_ ^ _43686_ /*24606*/;
assign _43691_ = _43682_ & _43690_ /*24604*/;
assign _43431_ = _43682_ ^ _43690_ /*24605*/;
assign _43688_ = _43689_ | _43691_ /*24602*/;
assign _43693_ = ~Q[15] /*24601*/;
assign _43692_ = _43693_ & D[39] /*24600*/;
assign _43695_ = _42984_ & _43692_ /*24595*/;
assign _43696_ = _42984_ ^ _43692_ /*24598*/;
assign _43697_ = _43688_ & _43696_ /*24596*/;
assign _43432_ = _43688_ ^ _43696_ /*24597*/;
assign _43694_ = _43695_ | _43697_ /*24594*/;
assign _43699_ = ~Q[15] /*24593*/;
assign _43698_ = _43699_ & D[40] /*24592*/;
assign _43701_ = _42985_ & _43698_ /*24587*/;
assign _43702_ = _42985_ ^ _43698_ /*24590*/;
assign _43703_ = _43694_ & _43702_ /*24588*/;
assign _43433_ = _43694_ ^ _43702_ /*24589*/;
assign _43700_ = _43701_ | _43703_ /*24586*/;
assign _43705_ = ~Q[15] /*24585*/;
assign _43704_ = _43705_ & D[41] /*24584*/;
assign _43707_ = _42986_ & _43704_ /*24579*/;
assign _43708_ = _42986_ ^ _43704_ /*24582*/;
assign _43709_ = _43700_ & _43708_ /*24580*/;
assign _43434_ = _43700_ ^ _43708_ /*24581*/;
assign _43706_ = _43707_ | _43709_ /*24578*/;
assign _43711_ = ~Q[15] /*24577*/;
assign _43710_ = _43711_ & D[42] /*24576*/;
assign _43713_ = _42987_ & _43710_ /*24571*/;
assign _43714_ = _42987_ ^ _43710_ /*24574*/;
assign _43715_ = _43706_ & _43714_ /*24572*/;
assign _43435_ = _43706_ ^ _43714_ /*24573*/;
assign _43712_ = _43713_ | _43715_ /*24570*/;
assign _43717_ = ~Q[15] /*24569*/;
assign _43716_ = _43717_ & D[43] /*24568*/;
assign _43719_ = _42988_ & _43716_ /*24563*/;
assign _43720_ = _42988_ ^ _43716_ /*24566*/;
assign _43721_ = _43712_ & _43720_ /*24564*/;
assign _43436_ = _43712_ ^ _43720_ /*24565*/;
assign _43718_ = _43719_ | _43721_ /*24562*/;
assign _43723_ = ~Q[15] /*24561*/;
assign _43722_ = _43723_ & D[44] /*24560*/;
assign _43725_ = _42989_ & _43722_ /*24555*/;
assign _43726_ = _42989_ ^ _43722_ /*24558*/;
assign _43727_ = _43718_ & _43726_ /*24556*/;
assign _43437_ = _43718_ ^ _43726_ /*24557*/;
assign _43724_ = _43725_ | _43727_ /*24554*/;
assign _43729_ = ~Q[15] /*24553*/;
assign _43728_ = _43729_ & D[45] /*24552*/;
assign _43731_ = _42990_ & _43728_ /*24547*/;
assign _43732_ = _42990_ ^ _43728_ /*24550*/;
assign _43733_ = _43724_ & _43732_ /*24548*/;
assign _43438_ = _43724_ ^ _43732_ /*24549*/;
assign _43730_ = _43731_ | _43733_ /*24546*/;
assign _43735_ = ~Q[15] /*24545*/;
assign _43734_ = _43735_ & D[46] /*24544*/;
assign _43737_ = _42991_ & _43734_ /*24539*/;
assign _43738_ = _42991_ ^ _43734_ /*24542*/;
assign _43739_ = _43730_ & _43738_ /*24540*/;
assign _43439_ = _43730_ ^ _43738_ /*24541*/;
assign _43736_ = _43737_ | _43739_ /*24538*/;
assign _43741_ = ~Q[15] /*24537*/;
assign _43740_ = _43741_ & D[47] /*24536*/;
assign _43743_ = _42992_ & _43740_ /*24531*/;
assign _43744_ = _42992_ ^ _43740_ /*24534*/;
assign _43745_ = _43736_ & _43744_ /*24532*/;
assign _43440_ = _43736_ ^ _43744_ /*24533*/;
assign _43742_ = _43743_ | _43745_ /*24530*/;
assign _43747_ = ~Q[15] /*24529*/;
assign _43746_ = _43747_ & D[48] /*24528*/;
assign _43749_ = _42993_ & _43746_ /*24523*/;
assign _43750_ = _42993_ ^ _43746_ /*24526*/;
assign _43751_ = _43742_ & _43750_ /*24524*/;
assign _43441_ = _43742_ ^ _43750_ /*24525*/;
assign _43748_ = _43749_ | _43751_ /*24522*/;
assign _43753_ = ~Q[15] /*24521*/;
assign _43752_ = _43753_ & D[49] /*24520*/;
assign _43755_ = _42994_ & _43752_ /*24515*/;
assign _43756_ = _42994_ ^ _43752_ /*24518*/;
assign _43757_ = _43748_ & _43756_ /*24516*/;
assign _43442_ = _43748_ ^ _43756_ /*24517*/;
assign _43754_ = _43755_ | _43757_ /*24514*/;
assign _43759_ = ~Q[15] /*24513*/;
assign _43758_ = _43759_ & D[50] /*24512*/;
assign _43761_ = _42995_ & _43758_ /*24507*/;
assign _43762_ = _42995_ ^ _43758_ /*24510*/;
assign _43763_ = _43754_ & _43762_ /*24508*/;
assign _43443_ = _43754_ ^ _43762_ /*24509*/;
assign _43760_ = _43761_ | _43763_ /*24506*/;
assign _43765_ = ~Q[15] /*24505*/;
assign _43764_ = _43765_ & D[51] /*24504*/;
assign _43767_ = _42996_ & _43764_ /*24499*/;
assign _43768_ = _42996_ ^ _43764_ /*24502*/;
assign _43769_ = _43760_ & _43768_ /*24500*/;
assign _43444_ = _43760_ ^ _43768_ /*24501*/;
assign _43766_ = _43767_ | _43769_ /*24498*/;
assign _43771_ = ~Q[15] /*24497*/;
assign _43770_ = _43771_ & D[52] /*24496*/;
assign _43773_ = _42997_ & _43770_ /*24491*/;
assign _43774_ = _42997_ ^ _43770_ /*24494*/;
assign _43775_ = _43766_ & _43774_ /*24492*/;
assign _43445_ = _43766_ ^ _43774_ /*24493*/;
assign _43772_ = _43773_ | _43775_ /*24490*/;
assign _43777_ = ~Q[15] /*24489*/;
assign _43776_ = _43777_ & D[53] /*24488*/;
assign _43779_ = _42998_ & _43776_ /*24483*/;
assign _43780_ = _42998_ ^ _43776_ /*24486*/;
assign _43781_ = _43772_ & _43780_ /*24484*/;
assign _43446_ = _43772_ ^ _43780_ /*24485*/;
assign _43778_ = _43779_ | _43781_ /*24482*/;
assign _43783_ = ~Q[15] /*24481*/;
assign _43782_ = _43783_ & D[54] /*24480*/;
assign _43785_ = _42999_ & _43782_ /*24475*/;
assign _43786_ = _42999_ ^ _43782_ /*24478*/;
assign _43787_ = _43778_ & _43786_ /*24476*/;
assign _43447_ = _43778_ ^ _43786_ /*24477*/;
assign _43784_ = _43785_ | _43787_ /*24474*/;
assign _43789_ = ~Q[15] /*24473*/;
assign _43788_ = _43789_ & D[55] /*24472*/;
assign _43791_ = _43000_ & _43788_ /*24467*/;
assign _43792_ = _43000_ ^ _43788_ /*24470*/;
assign _43793_ = _43784_ & _43792_ /*24468*/;
assign _43448_ = _43784_ ^ _43792_ /*24469*/;
assign _43790_ = _43791_ | _43793_ /*24466*/;
assign _43795_ = ~Q[15] /*24465*/;
assign _43794_ = _43795_ & D[56] /*24464*/;
assign _43797_ = _43001_ & _43794_ /*24459*/;
assign _43798_ = _43001_ ^ _43794_ /*24462*/;
assign _43799_ = _43790_ & _43798_ /*24460*/;
assign _43449_ = _43790_ ^ _43798_ /*24461*/;
assign _43796_ = _43797_ | _43799_ /*24458*/;
assign _43801_ = ~Q[15] /*24457*/;
assign _43800_ = _43801_ & D[57] /*24456*/;
assign _43803_ = _43002_ & _43800_ /*24451*/;
assign _43804_ = _43002_ ^ _43800_ /*24454*/;
assign _43805_ = _43796_ & _43804_ /*24452*/;
assign _43450_ = _43796_ ^ _43804_ /*24453*/;
assign _43802_ = _43803_ | _43805_ /*24450*/;
assign _43807_ = ~Q[15] /*24449*/;
assign _43806_ = _43807_ & D[58] /*24448*/;
assign _43809_ = _43003_ & _43806_ /*24443*/;
assign _43810_ = _43003_ ^ _43806_ /*24446*/;
assign _43811_ = _43802_ & _43810_ /*24444*/;
assign _43451_ = _43802_ ^ _43810_ /*24445*/;
assign _43808_ = _43809_ | _43811_ /*24442*/;
assign _43813_ = ~Q[15] /*24441*/;
assign _43812_ = _43813_ & D[59] /*24440*/;
assign _43815_ = _43004_ & _43812_ /*24435*/;
assign _43816_ = _43004_ ^ _43812_ /*24438*/;
assign _43817_ = _43808_ & _43816_ /*24436*/;
assign _43452_ = _43808_ ^ _43816_ /*24437*/;
assign _43814_ = _43815_ | _43817_ /*24434*/;
assign _43819_ = ~Q[15] /*24433*/;
assign _43818_ = _43819_ & D[60] /*24432*/;
assign _43821_ = _43005_ & _43818_ /*24427*/;
assign _43822_ = _43005_ ^ _43818_ /*24430*/;
assign _43823_ = _43814_ & _43822_ /*24428*/;
assign _43453_ = _43814_ ^ _43822_ /*24429*/;
assign _43820_ = _43821_ | _43823_ /*24426*/;
assign _43825_ = ~Q[15] /*24425*/;
assign _43824_ = _43825_ & D[61] /*24424*/;
assign _43827_ = _43006_ & _43824_ /*24419*/;
assign _43828_ = _43006_ ^ _43824_ /*24422*/;
assign _43829_ = _43820_ & _43828_ /*24420*/;
assign _43454_ = _43820_ ^ _43828_ /*24421*/;
assign _43826_ = _43827_ | _43829_ /*24418*/;
assign _43831_ = ~Q[15] /*24417*/;
assign _43830_ = _43831_ & D[62] /*24416*/;
assign _43833_ = _43007_ & _43830_ /*24411*/;
assign _43834_ = _43007_ ^ _43830_ /*24414*/;
assign _43835_ = _43826_ & _43834_ /*24412*/;
assign _43455_ = _43826_ ^ _43834_ /*24413*/;
assign _43832_ = _43833_ | _43835_ /*24410*/;
assign _43837_ = ~Q[15] /*24409*/;
assign _43836_ = _43837_ & zeroWire /*24408*/;
assign _43838_ = _43008_ ^ _43836_ /*24406*/;
assign _43456_ = _43838_ ^ _43832_ /*24405*/;
assign _43909_ = ~D[0] /*24151*/;
assign _43906_ = R_0[14] & _43909_ /*24147*/;
assign _43907_ = R_0[14] ^ _43909_ /*24150*/;
assign _43908_ = oneWire & _43907_ /*24148*/;
assign _43841_ = oneWire ^ _43907_ /*24149*/;
assign _43905_ = _43906_ | _43908_ /*24146*/;
assign _43914_ = ~D[1] /*24145*/;
assign _43911_ = _43393_ & _43914_ /*24141*/;
assign _43912_ = _43393_ ^ _43914_ /*24144*/;
assign _43913_ = _43905_ & _43912_ /*24142*/;
assign _43842_ = _43905_ ^ _43912_ /*24143*/;
assign _43910_ = _43911_ | _43913_ /*24140*/;
assign _43919_ = ~D[2] /*24139*/;
assign _43916_ = _43394_ & _43919_ /*24135*/;
assign _43917_ = _43394_ ^ _43919_ /*24138*/;
assign _43918_ = _43910_ & _43917_ /*24136*/;
assign _43843_ = _43910_ ^ _43917_ /*24137*/;
assign _43915_ = _43916_ | _43918_ /*24134*/;
assign _43924_ = ~D[3] /*24133*/;
assign _43921_ = _43395_ & _43924_ /*24129*/;
assign _43922_ = _43395_ ^ _43924_ /*24132*/;
assign _43923_ = _43915_ & _43922_ /*24130*/;
assign _43844_ = _43915_ ^ _43922_ /*24131*/;
assign _43920_ = _43921_ | _43923_ /*24128*/;
assign _43929_ = ~D[4] /*24127*/;
assign _43926_ = _43396_ & _43929_ /*24123*/;
assign _43927_ = _43396_ ^ _43929_ /*24126*/;
assign _43928_ = _43920_ & _43927_ /*24124*/;
assign _43845_ = _43920_ ^ _43927_ /*24125*/;
assign _43925_ = _43926_ | _43928_ /*24122*/;
assign _43934_ = ~D[5] /*24121*/;
assign _43931_ = _43397_ & _43934_ /*24117*/;
assign _43932_ = _43397_ ^ _43934_ /*24120*/;
assign _43933_ = _43925_ & _43932_ /*24118*/;
assign _43846_ = _43925_ ^ _43932_ /*24119*/;
assign _43930_ = _43931_ | _43933_ /*24116*/;
assign _43939_ = ~D[6] /*24115*/;
assign _43936_ = _43398_ & _43939_ /*24111*/;
assign _43937_ = _43398_ ^ _43939_ /*24114*/;
assign _43938_ = _43930_ & _43937_ /*24112*/;
assign _43847_ = _43930_ ^ _43937_ /*24113*/;
assign _43935_ = _43936_ | _43938_ /*24110*/;
assign _43944_ = ~D[7] /*24109*/;
assign _43941_ = _43399_ & _43944_ /*24105*/;
assign _43942_ = _43399_ ^ _43944_ /*24108*/;
assign _43943_ = _43935_ & _43942_ /*24106*/;
assign _43848_ = _43935_ ^ _43942_ /*24107*/;
assign _43940_ = _43941_ | _43943_ /*24104*/;
assign _43949_ = ~D[8] /*24103*/;
assign _43946_ = _43400_ & _43949_ /*24099*/;
assign _43947_ = _43400_ ^ _43949_ /*24102*/;
assign _43948_ = _43940_ & _43947_ /*24100*/;
assign _43849_ = _43940_ ^ _43947_ /*24101*/;
assign _43945_ = _43946_ | _43948_ /*24098*/;
assign _43954_ = ~D[9] /*24097*/;
assign _43951_ = _43401_ & _43954_ /*24093*/;
assign _43952_ = _43401_ ^ _43954_ /*24096*/;
assign _43953_ = _43945_ & _43952_ /*24094*/;
assign _43850_ = _43945_ ^ _43952_ /*24095*/;
assign _43950_ = _43951_ | _43953_ /*24092*/;
assign _43959_ = ~D[10] /*24091*/;
assign _43956_ = _43402_ & _43959_ /*24087*/;
assign _43957_ = _43402_ ^ _43959_ /*24090*/;
assign _43958_ = _43950_ & _43957_ /*24088*/;
assign _43851_ = _43950_ ^ _43957_ /*24089*/;
assign _43955_ = _43956_ | _43958_ /*24086*/;
assign _43964_ = ~D[11] /*24085*/;
assign _43961_ = _43403_ & _43964_ /*24081*/;
assign _43962_ = _43403_ ^ _43964_ /*24084*/;
assign _43963_ = _43955_ & _43962_ /*24082*/;
assign _43852_ = _43955_ ^ _43962_ /*24083*/;
assign _43960_ = _43961_ | _43963_ /*24080*/;
assign _43969_ = ~D[12] /*24079*/;
assign _43966_ = _43404_ & _43969_ /*24075*/;
assign _43967_ = _43404_ ^ _43969_ /*24078*/;
assign _43968_ = _43960_ & _43967_ /*24076*/;
assign _43853_ = _43960_ ^ _43967_ /*24077*/;
assign _43965_ = _43966_ | _43968_ /*24074*/;
assign _43974_ = ~D[13] /*24073*/;
assign _43971_ = _43405_ & _43974_ /*24069*/;
assign _43972_ = _43405_ ^ _43974_ /*24072*/;
assign _43973_ = _43965_ & _43972_ /*24070*/;
assign _43854_ = _43965_ ^ _43972_ /*24071*/;
assign _43970_ = _43971_ | _43973_ /*24068*/;
assign _43979_ = ~D[14] /*24067*/;
assign _43976_ = _43406_ & _43979_ /*24063*/;
assign _43977_ = _43406_ ^ _43979_ /*24066*/;
assign _43978_ = _43970_ & _43977_ /*24064*/;
assign _43855_ = _43970_ ^ _43977_ /*24065*/;
assign _43975_ = _43976_ | _43978_ /*24062*/;
assign _43984_ = ~D[15] /*24061*/;
assign _43981_ = _43407_ & _43984_ /*24057*/;
assign _43982_ = _43407_ ^ _43984_ /*24060*/;
assign _43983_ = _43975_ & _43982_ /*24058*/;
assign _43856_ = _43975_ ^ _43982_ /*24059*/;
assign _43980_ = _43981_ | _43983_ /*24056*/;
assign _43989_ = ~D[16] /*24055*/;
assign _43986_ = _43408_ & _43989_ /*24051*/;
assign _43987_ = _43408_ ^ _43989_ /*24054*/;
assign _43988_ = _43980_ & _43987_ /*24052*/;
assign _43857_ = _43980_ ^ _43987_ /*24053*/;
assign _43985_ = _43986_ | _43988_ /*24050*/;
assign _43994_ = ~D[17] /*24049*/;
assign _43991_ = _43409_ & _43994_ /*24045*/;
assign _43992_ = _43409_ ^ _43994_ /*24048*/;
assign _43993_ = _43985_ & _43992_ /*24046*/;
assign _43858_ = _43985_ ^ _43992_ /*24047*/;
assign _43990_ = _43991_ | _43993_ /*24044*/;
assign _43999_ = ~D[18] /*24043*/;
assign _43996_ = _43410_ & _43999_ /*24039*/;
assign _43997_ = _43410_ ^ _43999_ /*24042*/;
assign _43998_ = _43990_ & _43997_ /*24040*/;
assign _43859_ = _43990_ ^ _43997_ /*24041*/;
assign _43995_ = _43996_ | _43998_ /*24038*/;
assign _44004_ = ~D[19] /*24037*/;
assign _44001_ = _43411_ & _44004_ /*24033*/;
assign _44002_ = _43411_ ^ _44004_ /*24036*/;
assign _44003_ = _43995_ & _44002_ /*24034*/;
assign _43860_ = _43995_ ^ _44002_ /*24035*/;
assign _44000_ = _44001_ | _44003_ /*24032*/;
assign _44009_ = ~D[20] /*24031*/;
assign _44006_ = _43412_ & _44009_ /*24027*/;
assign _44007_ = _43412_ ^ _44009_ /*24030*/;
assign _44008_ = _44000_ & _44007_ /*24028*/;
assign _43861_ = _44000_ ^ _44007_ /*24029*/;
assign _44005_ = _44006_ | _44008_ /*24026*/;
assign _44014_ = ~D[21] /*24025*/;
assign _44011_ = _43413_ & _44014_ /*24021*/;
assign _44012_ = _43413_ ^ _44014_ /*24024*/;
assign _44013_ = _44005_ & _44012_ /*24022*/;
assign _43862_ = _44005_ ^ _44012_ /*24023*/;
assign _44010_ = _44011_ | _44013_ /*24020*/;
assign _44019_ = ~D[22] /*24019*/;
assign _44016_ = _43414_ & _44019_ /*24015*/;
assign _44017_ = _43414_ ^ _44019_ /*24018*/;
assign _44018_ = _44010_ & _44017_ /*24016*/;
assign _43863_ = _44010_ ^ _44017_ /*24017*/;
assign _44015_ = _44016_ | _44018_ /*24014*/;
assign _44024_ = ~D[23] /*24013*/;
assign _44021_ = _43415_ & _44024_ /*24009*/;
assign _44022_ = _43415_ ^ _44024_ /*24012*/;
assign _44023_ = _44015_ & _44022_ /*24010*/;
assign _43864_ = _44015_ ^ _44022_ /*24011*/;
assign _44020_ = _44021_ | _44023_ /*24008*/;
assign _44029_ = ~D[24] /*24007*/;
assign _44026_ = _43416_ & _44029_ /*24003*/;
assign _44027_ = _43416_ ^ _44029_ /*24006*/;
assign _44028_ = _44020_ & _44027_ /*24004*/;
assign _43865_ = _44020_ ^ _44027_ /*24005*/;
assign _44025_ = _44026_ | _44028_ /*24002*/;
assign _44034_ = ~D[25] /*24001*/;
assign _44031_ = _43417_ & _44034_ /*23997*/;
assign _44032_ = _43417_ ^ _44034_ /*24000*/;
assign _44033_ = _44025_ & _44032_ /*23998*/;
assign _43866_ = _44025_ ^ _44032_ /*23999*/;
assign _44030_ = _44031_ | _44033_ /*23996*/;
assign _44039_ = ~D[26] /*23995*/;
assign _44036_ = _43418_ & _44039_ /*23991*/;
assign _44037_ = _43418_ ^ _44039_ /*23994*/;
assign _44038_ = _44030_ & _44037_ /*23992*/;
assign _43867_ = _44030_ ^ _44037_ /*23993*/;
assign _44035_ = _44036_ | _44038_ /*23990*/;
assign _44044_ = ~D[27] /*23989*/;
assign _44041_ = _43419_ & _44044_ /*23985*/;
assign _44042_ = _43419_ ^ _44044_ /*23988*/;
assign _44043_ = _44035_ & _44042_ /*23986*/;
assign _43868_ = _44035_ ^ _44042_ /*23987*/;
assign _44040_ = _44041_ | _44043_ /*23984*/;
assign _44049_ = ~D[28] /*23983*/;
assign _44046_ = _43420_ & _44049_ /*23979*/;
assign _44047_ = _43420_ ^ _44049_ /*23982*/;
assign _44048_ = _44040_ & _44047_ /*23980*/;
assign _43869_ = _44040_ ^ _44047_ /*23981*/;
assign _44045_ = _44046_ | _44048_ /*23978*/;
assign _44054_ = ~D[29] /*23977*/;
assign _44051_ = _43421_ & _44054_ /*23973*/;
assign _44052_ = _43421_ ^ _44054_ /*23976*/;
assign _44053_ = _44045_ & _44052_ /*23974*/;
assign _43870_ = _44045_ ^ _44052_ /*23975*/;
assign _44050_ = _44051_ | _44053_ /*23972*/;
assign _44059_ = ~D[30] /*23971*/;
assign _44056_ = _43422_ & _44059_ /*23967*/;
assign _44057_ = _43422_ ^ _44059_ /*23970*/;
assign _44058_ = _44050_ & _44057_ /*23968*/;
assign _43871_ = _44050_ ^ _44057_ /*23969*/;
assign _44055_ = _44056_ | _44058_ /*23966*/;
assign _44064_ = ~D[31] /*23965*/;
assign _44061_ = _43423_ & _44064_ /*23961*/;
assign _44062_ = _43423_ ^ _44064_ /*23964*/;
assign _44063_ = _44055_ & _44062_ /*23962*/;
assign _43872_ = _44055_ ^ _44062_ /*23963*/;
assign _44060_ = _44061_ | _44063_ /*23960*/;
assign _44069_ = ~D[32] /*23959*/;
assign _44066_ = _43424_ & _44069_ /*23955*/;
assign _44067_ = _43424_ ^ _44069_ /*23958*/;
assign _44068_ = _44060_ & _44067_ /*23956*/;
assign _43873_ = _44060_ ^ _44067_ /*23957*/;
assign _44065_ = _44066_ | _44068_ /*23954*/;
assign _44074_ = ~D[33] /*23953*/;
assign _44071_ = _43425_ & _44074_ /*23949*/;
assign _44072_ = _43425_ ^ _44074_ /*23952*/;
assign _44073_ = _44065_ & _44072_ /*23950*/;
assign _43874_ = _44065_ ^ _44072_ /*23951*/;
assign _44070_ = _44071_ | _44073_ /*23948*/;
assign _44079_ = ~D[34] /*23947*/;
assign _44076_ = _43426_ & _44079_ /*23943*/;
assign _44077_ = _43426_ ^ _44079_ /*23946*/;
assign _44078_ = _44070_ & _44077_ /*23944*/;
assign _43875_ = _44070_ ^ _44077_ /*23945*/;
assign _44075_ = _44076_ | _44078_ /*23942*/;
assign _44084_ = ~D[35] /*23941*/;
assign _44081_ = _43427_ & _44084_ /*23937*/;
assign _44082_ = _43427_ ^ _44084_ /*23940*/;
assign _44083_ = _44075_ & _44082_ /*23938*/;
assign _43876_ = _44075_ ^ _44082_ /*23939*/;
assign _44080_ = _44081_ | _44083_ /*23936*/;
assign _44089_ = ~D[36] /*23935*/;
assign _44086_ = _43428_ & _44089_ /*23931*/;
assign _44087_ = _43428_ ^ _44089_ /*23934*/;
assign _44088_ = _44080_ & _44087_ /*23932*/;
assign _43877_ = _44080_ ^ _44087_ /*23933*/;
assign _44085_ = _44086_ | _44088_ /*23930*/;
assign _44094_ = ~D[37] /*23929*/;
assign _44091_ = _43429_ & _44094_ /*23925*/;
assign _44092_ = _43429_ ^ _44094_ /*23928*/;
assign _44093_ = _44085_ & _44092_ /*23926*/;
assign _43878_ = _44085_ ^ _44092_ /*23927*/;
assign _44090_ = _44091_ | _44093_ /*23924*/;
assign _44099_ = ~D[38] /*23923*/;
assign _44096_ = _43430_ & _44099_ /*23919*/;
assign _44097_ = _43430_ ^ _44099_ /*23922*/;
assign _44098_ = _44090_ & _44097_ /*23920*/;
assign _43879_ = _44090_ ^ _44097_ /*23921*/;
assign _44095_ = _44096_ | _44098_ /*23918*/;
assign _44104_ = ~D[39] /*23917*/;
assign _44101_ = _43431_ & _44104_ /*23913*/;
assign _44102_ = _43431_ ^ _44104_ /*23916*/;
assign _44103_ = _44095_ & _44102_ /*23914*/;
assign _43880_ = _44095_ ^ _44102_ /*23915*/;
assign _44100_ = _44101_ | _44103_ /*23912*/;
assign _44109_ = ~D[40] /*23911*/;
assign _44106_ = _43432_ & _44109_ /*23907*/;
assign _44107_ = _43432_ ^ _44109_ /*23910*/;
assign _44108_ = _44100_ & _44107_ /*23908*/;
assign _43881_ = _44100_ ^ _44107_ /*23909*/;
assign _44105_ = _44106_ | _44108_ /*23906*/;
assign _44114_ = ~D[41] /*23905*/;
assign _44111_ = _43433_ & _44114_ /*23901*/;
assign _44112_ = _43433_ ^ _44114_ /*23904*/;
assign _44113_ = _44105_ & _44112_ /*23902*/;
assign _43882_ = _44105_ ^ _44112_ /*23903*/;
assign _44110_ = _44111_ | _44113_ /*23900*/;
assign _44119_ = ~D[42] /*23899*/;
assign _44116_ = _43434_ & _44119_ /*23895*/;
assign _44117_ = _43434_ ^ _44119_ /*23898*/;
assign _44118_ = _44110_ & _44117_ /*23896*/;
assign _43883_ = _44110_ ^ _44117_ /*23897*/;
assign _44115_ = _44116_ | _44118_ /*23894*/;
assign _44124_ = ~D[43] /*23893*/;
assign _44121_ = _43435_ & _44124_ /*23889*/;
assign _44122_ = _43435_ ^ _44124_ /*23892*/;
assign _44123_ = _44115_ & _44122_ /*23890*/;
assign _43884_ = _44115_ ^ _44122_ /*23891*/;
assign _44120_ = _44121_ | _44123_ /*23888*/;
assign _44129_ = ~D[44] /*23887*/;
assign _44126_ = _43436_ & _44129_ /*23883*/;
assign _44127_ = _43436_ ^ _44129_ /*23886*/;
assign _44128_ = _44120_ & _44127_ /*23884*/;
assign _43885_ = _44120_ ^ _44127_ /*23885*/;
assign _44125_ = _44126_ | _44128_ /*23882*/;
assign _44134_ = ~D[45] /*23881*/;
assign _44131_ = _43437_ & _44134_ /*23877*/;
assign _44132_ = _43437_ ^ _44134_ /*23880*/;
assign _44133_ = _44125_ & _44132_ /*23878*/;
assign _43886_ = _44125_ ^ _44132_ /*23879*/;
assign _44130_ = _44131_ | _44133_ /*23876*/;
assign _44139_ = ~D[46] /*23875*/;
assign _44136_ = _43438_ & _44139_ /*23871*/;
assign _44137_ = _43438_ ^ _44139_ /*23874*/;
assign _44138_ = _44130_ & _44137_ /*23872*/;
assign _43887_ = _44130_ ^ _44137_ /*23873*/;
assign _44135_ = _44136_ | _44138_ /*23870*/;
assign _44144_ = ~D[47] /*23869*/;
assign _44141_ = _43439_ & _44144_ /*23865*/;
assign _44142_ = _43439_ ^ _44144_ /*23868*/;
assign _44143_ = _44135_ & _44142_ /*23866*/;
assign _43888_ = _44135_ ^ _44142_ /*23867*/;
assign _44140_ = _44141_ | _44143_ /*23864*/;
assign _44149_ = ~D[48] /*23863*/;
assign _44146_ = _43440_ & _44149_ /*23859*/;
assign _44147_ = _43440_ ^ _44149_ /*23862*/;
assign _44148_ = _44140_ & _44147_ /*23860*/;
assign _43889_ = _44140_ ^ _44147_ /*23861*/;
assign _44145_ = _44146_ | _44148_ /*23858*/;
assign _44154_ = ~D[49] /*23857*/;
assign _44151_ = _43441_ & _44154_ /*23853*/;
assign _44152_ = _43441_ ^ _44154_ /*23856*/;
assign _44153_ = _44145_ & _44152_ /*23854*/;
assign _43890_ = _44145_ ^ _44152_ /*23855*/;
assign _44150_ = _44151_ | _44153_ /*23852*/;
assign _44159_ = ~D[50] /*23851*/;
assign _44156_ = _43442_ & _44159_ /*23847*/;
assign _44157_ = _43442_ ^ _44159_ /*23850*/;
assign _44158_ = _44150_ & _44157_ /*23848*/;
assign _43891_ = _44150_ ^ _44157_ /*23849*/;
assign _44155_ = _44156_ | _44158_ /*23846*/;
assign _44164_ = ~D[51] /*23845*/;
assign _44161_ = _43443_ & _44164_ /*23841*/;
assign _44162_ = _43443_ ^ _44164_ /*23844*/;
assign _44163_ = _44155_ & _44162_ /*23842*/;
assign _43892_ = _44155_ ^ _44162_ /*23843*/;
assign _44160_ = _44161_ | _44163_ /*23840*/;
assign _44169_ = ~D[52] /*23839*/;
assign _44166_ = _43444_ & _44169_ /*23835*/;
assign _44167_ = _43444_ ^ _44169_ /*23838*/;
assign _44168_ = _44160_ & _44167_ /*23836*/;
assign _43893_ = _44160_ ^ _44167_ /*23837*/;
assign _44165_ = _44166_ | _44168_ /*23834*/;
assign _44174_ = ~D[53] /*23833*/;
assign _44171_ = _43445_ & _44174_ /*23829*/;
assign _44172_ = _43445_ ^ _44174_ /*23832*/;
assign _44173_ = _44165_ & _44172_ /*23830*/;
assign _43894_ = _44165_ ^ _44172_ /*23831*/;
assign _44170_ = _44171_ | _44173_ /*23828*/;
assign _44179_ = ~D[54] /*23827*/;
assign _44176_ = _43446_ & _44179_ /*23823*/;
assign _44177_ = _43446_ ^ _44179_ /*23826*/;
assign _44178_ = _44170_ & _44177_ /*23824*/;
assign _43895_ = _44170_ ^ _44177_ /*23825*/;
assign _44175_ = _44176_ | _44178_ /*23822*/;
assign _44184_ = ~D[55] /*23821*/;
assign _44181_ = _43447_ & _44184_ /*23817*/;
assign _44182_ = _43447_ ^ _44184_ /*23820*/;
assign _44183_ = _44175_ & _44182_ /*23818*/;
assign _43896_ = _44175_ ^ _44182_ /*23819*/;
assign _44180_ = _44181_ | _44183_ /*23816*/;
assign _44189_ = ~D[56] /*23815*/;
assign _44186_ = _43448_ & _44189_ /*23811*/;
assign _44187_ = _43448_ ^ _44189_ /*23814*/;
assign _44188_ = _44180_ & _44187_ /*23812*/;
assign _43897_ = _44180_ ^ _44187_ /*23813*/;
assign _44185_ = _44186_ | _44188_ /*23810*/;
assign _44194_ = ~D[57] /*23809*/;
assign _44191_ = _43449_ & _44194_ /*23805*/;
assign _44192_ = _43449_ ^ _44194_ /*23808*/;
assign _44193_ = _44185_ & _44192_ /*23806*/;
assign _43898_ = _44185_ ^ _44192_ /*23807*/;
assign _44190_ = _44191_ | _44193_ /*23804*/;
assign _44199_ = ~D[58] /*23803*/;
assign _44196_ = _43450_ & _44199_ /*23799*/;
assign _44197_ = _43450_ ^ _44199_ /*23802*/;
assign _44198_ = _44190_ & _44197_ /*23800*/;
assign _43899_ = _44190_ ^ _44197_ /*23801*/;
assign _44195_ = _44196_ | _44198_ /*23798*/;
assign _44204_ = ~D[59] /*23797*/;
assign _44201_ = _43451_ & _44204_ /*23793*/;
assign _44202_ = _43451_ ^ _44204_ /*23796*/;
assign _44203_ = _44195_ & _44202_ /*23794*/;
assign _43900_ = _44195_ ^ _44202_ /*23795*/;
assign _44200_ = _44201_ | _44203_ /*23792*/;
assign _44209_ = ~D[60] /*23791*/;
assign _44206_ = _43452_ & _44209_ /*23787*/;
assign _44207_ = _43452_ ^ _44209_ /*23790*/;
assign _44208_ = _44200_ & _44207_ /*23788*/;
assign _43901_ = _44200_ ^ _44207_ /*23789*/;
assign _44205_ = _44206_ | _44208_ /*23786*/;
assign _44214_ = ~D[61] /*23785*/;
assign _44211_ = _43453_ & _44214_ /*23781*/;
assign _44212_ = _43453_ ^ _44214_ /*23784*/;
assign _44213_ = _44205_ & _44212_ /*23782*/;
assign _43902_ = _44205_ ^ _44212_ /*23783*/;
assign _44210_ = _44211_ | _44213_ /*23780*/;
assign _44219_ = ~D[62] /*23779*/;
assign _44216_ = _43454_ & _44219_ /*23775*/;
assign _44217_ = _43454_ ^ _44219_ /*23778*/;
assign _44218_ = _44210_ & _44217_ /*23776*/;
assign _43903_ = _44210_ ^ _44217_ /*23777*/;
assign _44215_ = _44216_ | _44218_ /*23774*/;
assign _44220_ = _43455_ & oneWire /*23769*/;
assign _44221_ = _43455_ ^ oneWire /*23772*/;
assign _44222_ = _44215_ & _44221_ /*23770*/;
assign _43904_ = _44215_ ^ _44221_ /*23771*/;
assign Q[14] = _44220_ | _44222_ /*23768*/;
assign _44355_ = ~Q[14] /*23383*/;
assign _44354_ = _44355_ & D[0] /*23382*/;
assign _44357_ = _43841_ & _44354_ /*23377*/;
assign _44358_ = _43841_ ^ _44354_ /*23380*/;
assign _44359_ = zeroWire & _44358_ /*23378*/;
assign _44289_ = zeroWire ^ _44358_ /*23379*/;
assign _44356_ = _44357_ | _44359_ /*23376*/;
assign _44361_ = ~Q[14] /*23375*/;
assign _44360_ = _44361_ & D[1] /*23374*/;
assign _44363_ = _43842_ & _44360_ /*23369*/;
assign _44364_ = _43842_ ^ _44360_ /*23372*/;
assign _44365_ = _44356_ & _44364_ /*23370*/;
assign _44290_ = _44356_ ^ _44364_ /*23371*/;
assign _44362_ = _44363_ | _44365_ /*23368*/;
assign _44367_ = ~Q[14] /*23367*/;
assign _44366_ = _44367_ & D[2] /*23366*/;
assign _44369_ = _43843_ & _44366_ /*23361*/;
assign _44370_ = _43843_ ^ _44366_ /*23364*/;
assign _44371_ = _44362_ & _44370_ /*23362*/;
assign _44291_ = _44362_ ^ _44370_ /*23363*/;
assign _44368_ = _44369_ | _44371_ /*23360*/;
assign _44373_ = ~Q[14] /*23359*/;
assign _44372_ = _44373_ & D[3] /*23358*/;
assign _44375_ = _43844_ & _44372_ /*23353*/;
assign _44376_ = _43844_ ^ _44372_ /*23356*/;
assign _44377_ = _44368_ & _44376_ /*23354*/;
assign _44292_ = _44368_ ^ _44376_ /*23355*/;
assign _44374_ = _44375_ | _44377_ /*23352*/;
assign _44379_ = ~Q[14] /*23351*/;
assign _44378_ = _44379_ & D[4] /*23350*/;
assign _44381_ = _43845_ & _44378_ /*23345*/;
assign _44382_ = _43845_ ^ _44378_ /*23348*/;
assign _44383_ = _44374_ & _44382_ /*23346*/;
assign _44293_ = _44374_ ^ _44382_ /*23347*/;
assign _44380_ = _44381_ | _44383_ /*23344*/;
assign _44385_ = ~Q[14] /*23343*/;
assign _44384_ = _44385_ & D[5] /*23342*/;
assign _44387_ = _43846_ & _44384_ /*23337*/;
assign _44388_ = _43846_ ^ _44384_ /*23340*/;
assign _44389_ = _44380_ & _44388_ /*23338*/;
assign _44294_ = _44380_ ^ _44388_ /*23339*/;
assign _44386_ = _44387_ | _44389_ /*23336*/;
assign _44391_ = ~Q[14] /*23335*/;
assign _44390_ = _44391_ & D[6] /*23334*/;
assign _44393_ = _43847_ & _44390_ /*23329*/;
assign _44394_ = _43847_ ^ _44390_ /*23332*/;
assign _44395_ = _44386_ & _44394_ /*23330*/;
assign _44295_ = _44386_ ^ _44394_ /*23331*/;
assign _44392_ = _44393_ | _44395_ /*23328*/;
assign _44397_ = ~Q[14] /*23327*/;
assign _44396_ = _44397_ & D[7] /*23326*/;
assign _44399_ = _43848_ & _44396_ /*23321*/;
assign _44400_ = _43848_ ^ _44396_ /*23324*/;
assign _44401_ = _44392_ & _44400_ /*23322*/;
assign _44296_ = _44392_ ^ _44400_ /*23323*/;
assign _44398_ = _44399_ | _44401_ /*23320*/;
assign _44403_ = ~Q[14] /*23319*/;
assign _44402_ = _44403_ & D[8] /*23318*/;
assign _44405_ = _43849_ & _44402_ /*23313*/;
assign _44406_ = _43849_ ^ _44402_ /*23316*/;
assign _44407_ = _44398_ & _44406_ /*23314*/;
assign _44297_ = _44398_ ^ _44406_ /*23315*/;
assign _44404_ = _44405_ | _44407_ /*23312*/;
assign _44409_ = ~Q[14] /*23311*/;
assign _44408_ = _44409_ & D[9] /*23310*/;
assign _44411_ = _43850_ & _44408_ /*23305*/;
assign _44412_ = _43850_ ^ _44408_ /*23308*/;
assign _44413_ = _44404_ & _44412_ /*23306*/;
assign _44298_ = _44404_ ^ _44412_ /*23307*/;
assign _44410_ = _44411_ | _44413_ /*23304*/;
assign _44415_ = ~Q[14] /*23303*/;
assign _44414_ = _44415_ & D[10] /*23302*/;
assign _44417_ = _43851_ & _44414_ /*23297*/;
assign _44418_ = _43851_ ^ _44414_ /*23300*/;
assign _44419_ = _44410_ & _44418_ /*23298*/;
assign _44299_ = _44410_ ^ _44418_ /*23299*/;
assign _44416_ = _44417_ | _44419_ /*23296*/;
assign _44421_ = ~Q[14] /*23295*/;
assign _44420_ = _44421_ & D[11] /*23294*/;
assign _44423_ = _43852_ & _44420_ /*23289*/;
assign _44424_ = _43852_ ^ _44420_ /*23292*/;
assign _44425_ = _44416_ & _44424_ /*23290*/;
assign _44300_ = _44416_ ^ _44424_ /*23291*/;
assign _44422_ = _44423_ | _44425_ /*23288*/;
assign _44427_ = ~Q[14] /*23287*/;
assign _44426_ = _44427_ & D[12] /*23286*/;
assign _44429_ = _43853_ & _44426_ /*23281*/;
assign _44430_ = _43853_ ^ _44426_ /*23284*/;
assign _44431_ = _44422_ & _44430_ /*23282*/;
assign _44301_ = _44422_ ^ _44430_ /*23283*/;
assign _44428_ = _44429_ | _44431_ /*23280*/;
assign _44433_ = ~Q[14] /*23279*/;
assign _44432_ = _44433_ & D[13] /*23278*/;
assign _44435_ = _43854_ & _44432_ /*23273*/;
assign _44436_ = _43854_ ^ _44432_ /*23276*/;
assign _44437_ = _44428_ & _44436_ /*23274*/;
assign _44302_ = _44428_ ^ _44436_ /*23275*/;
assign _44434_ = _44435_ | _44437_ /*23272*/;
assign _44439_ = ~Q[14] /*23271*/;
assign _44438_ = _44439_ & D[14] /*23270*/;
assign _44441_ = _43855_ & _44438_ /*23265*/;
assign _44442_ = _43855_ ^ _44438_ /*23268*/;
assign _44443_ = _44434_ & _44442_ /*23266*/;
assign _44303_ = _44434_ ^ _44442_ /*23267*/;
assign _44440_ = _44441_ | _44443_ /*23264*/;
assign _44445_ = ~Q[14] /*23263*/;
assign _44444_ = _44445_ & D[15] /*23262*/;
assign _44447_ = _43856_ & _44444_ /*23257*/;
assign _44448_ = _43856_ ^ _44444_ /*23260*/;
assign _44449_ = _44440_ & _44448_ /*23258*/;
assign _44304_ = _44440_ ^ _44448_ /*23259*/;
assign _44446_ = _44447_ | _44449_ /*23256*/;
assign _44451_ = ~Q[14] /*23255*/;
assign _44450_ = _44451_ & D[16] /*23254*/;
assign _44453_ = _43857_ & _44450_ /*23249*/;
assign _44454_ = _43857_ ^ _44450_ /*23252*/;
assign _44455_ = _44446_ & _44454_ /*23250*/;
assign _44305_ = _44446_ ^ _44454_ /*23251*/;
assign _44452_ = _44453_ | _44455_ /*23248*/;
assign _44457_ = ~Q[14] /*23247*/;
assign _44456_ = _44457_ & D[17] /*23246*/;
assign _44459_ = _43858_ & _44456_ /*23241*/;
assign _44460_ = _43858_ ^ _44456_ /*23244*/;
assign _44461_ = _44452_ & _44460_ /*23242*/;
assign _44306_ = _44452_ ^ _44460_ /*23243*/;
assign _44458_ = _44459_ | _44461_ /*23240*/;
assign _44463_ = ~Q[14] /*23239*/;
assign _44462_ = _44463_ & D[18] /*23238*/;
assign _44465_ = _43859_ & _44462_ /*23233*/;
assign _44466_ = _43859_ ^ _44462_ /*23236*/;
assign _44467_ = _44458_ & _44466_ /*23234*/;
assign _44307_ = _44458_ ^ _44466_ /*23235*/;
assign _44464_ = _44465_ | _44467_ /*23232*/;
assign _44469_ = ~Q[14] /*23231*/;
assign _44468_ = _44469_ & D[19] /*23230*/;
assign _44471_ = _43860_ & _44468_ /*23225*/;
assign _44472_ = _43860_ ^ _44468_ /*23228*/;
assign _44473_ = _44464_ & _44472_ /*23226*/;
assign _44308_ = _44464_ ^ _44472_ /*23227*/;
assign _44470_ = _44471_ | _44473_ /*23224*/;
assign _44475_ = ~Q[14] /*23223*/;
assign _44474_ = _44475_ & D[20] /*23222*/;
assign _44477_ = _43861_ & _44474_ /*23217*/;
assign _44478_ = _43861_ ^ _44474_ /*23220*/;
assign _44479_ = _44470_ & _44478_ /*23218*/;
assign _44309_ = _44470_ ^ _44478_ /*23219*/;
assign _44476_ = _44477_ | _44479_ /*23216*/;
assign _44481_ = ~Q[14] /*23215*/;
assign _44480_ = _44481_ & D[21] /*23214*/;
assign _44483_ = _43862_ & _44480_ /*23209*/;
assign _44484_ = _43862_ ^ _44480_ /*23212*/;
assign _44485_ = _44476_ & _44484_ /*23210*/;
assign _44310_ = _44476_ ^ _44484_ /*23211*/;
assign _44482_ = _44483_ | _44485_ /*23208*/;
assign _44487_ = ~Q[14] /*23207*/;
assign _44486_ = _44487_ & D[22] /*23206*/;
assign _44489_ = _43863_ & _44486_ /*23201*/;
assign _44490_ = _43863_ ^ _44486_ /*23204*/;
assign _44491_ = _44482_ & _44490_ /*23202*/;
assign _44311_ = _44482_ ^ _44490_ /*23203*/;
assign _44488_ = _44489_ | _44491_ /*23200*/;
assign _44493_ = ~Q[14] /*23199*/;
assign _44492_ = _44493_ & D[23] /*23198*/;
assign _44495_ = _43864_ & _44492_ /*23193*/;
assign _44496_ = _43864_ ^ _44492_ /*23196*/;
assign _44497_ = _44488_ & _44496_ /*23194*/;
assign _44312_ = _44488_ ^ _44496_ /*23195*/;
assign _44494_ = _44495_ | _44497_ /*23192*/;
assign _44499_ = ~Q[14] /*23191*/;
assign _44498_ = _44499_ & D[24] /*23190*/;
assign _44501_ = _43865_ & _44498_ /*23185*/;
assign _44502_ = _43865_ ^ _44498_ /*23188*/;
assign _44503_ = _44494_ & _44502_ /*23186*/;
assign _44313_ = _44494_ ^ _44502_ /*23187*/;
assign _44500_ = _44501_ | _44503_ /*23184*/;
assign _44505_ = ~Q[14] /*23183*/;
assign _44504_ = _44505_ & D[25] /*23182*/;
assign _44507_ = _43866_ & _44504_ /*23177*/;
assign _44508_ = _43866_ ^ _44504_ /*23180*/;
assign _44509_ = _44500_ & _44508_ /*23178*/;
assign _44314_ = _44500_ ^ _44508_ /*23179*/;
assign _44506_ = _44507_ | _44509_ /*23176*/;
assign _44511_ = ~Q[14] /*23175*/;
assign _44510_ = _44511_ & D[26] /*23174*/;
assign _44513_ = _43867_ & _44510_ /*23169*/;
assign _44514_ = _43867_ ^ _44510_ /*23172*/;
assign _44515_ = _44506_ & _44514_ /*23170*/;
assign _44315_ = _44506_ ^ _44514_ /*23171*/;
assign _44512_ = _44513_ | _44515_ /*23168*/;
assign _44517_ = ~Q[14] /*23167*/;
assign _44516_ = _44517_ & D[27] /*23166*/;
assign _44519_ = _43868_ & _44516_ /*23161*/;
assign _44520_ = _43868_ ^ _44516_ /*23164*/;
assign _44521_ = _44512_ & _44520_ /*23162*/;
assign _44316_ = _44512_ ^ _44520_ /*23163*/;
assign _44518_ = _44519_ | _44521_ /*23160*/;
assign _44523_ = ~Q[14] /*23159*/;
assign _44522_ = _44523_ & D[28] /*23158*/;
assign _44525_ = _43869_ & _44522_ /*23153*/;
assign _44526_ = _43869_ ^ _44522_ /*23156*/;
assign _44527_ = _44518_ & _44526_ /*23154*/;
assign _44317_ = _44518_ ^ _44526_ /*23155*/;
assign _44524_ = _44525_ | _44527_ /*23152*/;
assign _44529_ = ~Q[14] /*23151*/;
assign _44528_ = _44529_ & D[29] /*23150*/;
assign _44531_ = _43870_ & _44528_ /*23145*/;
assign _44532_ = _43870_ ^ _44528_ /*23148*/;
assign _44533_ = _44524_ & _44532_ /*23146*/;
assign _44318_ = _44524_ ^ _44532_ /*23147*/;
assign _44530_ = _44531_ | _44533_ /*23144*/;
assign _44535_ = ~Q[14] /*23143*/;
assign _44534_ = _44535_ & D[30] /*23142*/;
assign _44537_ = _43871_ & _44534_ /*23137*/;
assign _44538_ = _43871_ ^ _44534_ /*23140*/;
assign _44539_ = _44530_ & _44538_ /*23138*/;
assign _44319_ = _44530_ ^ _44538_ /*23139*/;
assign _44536_ = _44537_ | _44539_ /*23136*/;
assign _44541_ = ~Q[14] /*23135*/;
assign _44540_ = _44541_ & D[31] /*23134*/;
assign _44543_ = _43872_ & _44540_ /*23129*/;
assign _44544_ = _43872_ ^ _44540_ /*23132*/;
assign _44545_ = _44536_ & _44544_ /*23130*/;
assign _44320_ = _44536_ ^ _44544_ /*23131*/;
assign _44542_ = _44543_ | _44545_ /*23128*/;
assign _44547_ = ~Q[14] /*23127*/;
assign _44546_ = _44547_ & D[32] /*23126*/;
assign _44549_ = _43873_ & _44546_ /*23121*/;
assign _44550_ = _43873_ ^ _44546_ /*23124*/;
assign _44551_ = _44542_ & _44550_ /*23122*/;
assign _44321_ = _44542_ ^ _44550_ /*23123*/;
assign _44548_ = _44549_ | _44551_ /*23120*/;
assign _44553_ = ~Q[14] /*23119*/;
assign _44552_ = _44553_ & D[33] /*23118*/;
assign _44555_ = _43874_ & _44552_ /*23113*/;
assign _44556_ = _43874_ ^ _44552_ /*23116*/;
assign _44557_ = _44548_ & _44556_ /*23114*/;
assign _44322_ = _44548_ ^ _44556_ /*23115*/;
assign _44554_ = _44555_ | _44557_ /*23112*/;
assign _44559_ = ~Q[14] /*23111*/;
assign _44558_ = _44559_ & D[34] /*23110*/;
assign _44561_ = _43875_ & _44558_ /*23105*/;
assign _44562_ = _43875_ ^ _44558_ /*23108*/;
assign _44563_ = _44554_ & _44562_ /*23106*/;
assign _44323_ = _44554_ ^ _44562_ /*23107*/;
assign _44560_ = _44561_ | _44563_ /*23104*/;
assign _44565_ = ~Q[14] /*23103*/;
assign _44564_ = _44565_ & D[35] /*23102*/;
assign _44567_ = _43876_ & _44564_ /*23097*/;
assign _44568_ = _43876_ ^ _44564_ /*23100*/;
assign _44569_ = _44560_ & _44568_ /*23098*/;
assign _44324_ = _44560_ ^ _44568_ /*23099*/;
assign _44566_ = _44567_ | _44569_ /*23096*/;
assign _44571_ = ~Q[14] /*23095*/;
assign _44570_ = _44571_ & D[36] /*23094*/;
assign _44573_ = _43877_ & _44570_ /*23089*/;
assign _44574_ = _43877_ ^ _44570_ /*23092*/;
assign _44575_ = _44566_ & _44574_ /*23090*/;
assign _44325_ = _44566_ ^ _44574_ /*23091*/;
assign _44572_ = _44573_ | _44575_ /*23088*/;
assign _44577_ = ~Q[14] /*23087*/;
assign _44576_ = _44577_ & D[37] /*23086*/;
assign _44579_ = _43878_ & _44576_ /*23081*/;
assign _44580_ = _43878_ ^ _44576_ /*23084*/;
assign _44581_ = _44572_ & _44580_ /*23082*/;
assign _44326_ = _44572_ ^ _44580_ /*23083*/;
assign _44578_ = _44579_ | _44581_ /*23080*/;
assign _44583_ = ~Q[14] /*23079*/;
assign _44582_ = _44583_ & D[38] /*23078*/;
assign _44585_ = _43879_ & _44582_ /*23073*/;
assign _44586_ = _43879_ ^ _44582_ /*23076*/;
assign _44587_ = _44578_ & _44586_ /*23074*/;
assign _44327_ = _44578_ ^ _44586_ /*23075*/;
assign _44584_ = _44585_ | _44587_ /*23072*/;
assign _44589_ = ~Q[14] /*23071*/;
assign _44588_ = _44589_ & D[39] /*23070*/;
assign _44591_ = _43880_ & _44588_ /*23065*/;
assign _44592_ = _43880_ ^ _44588_ /*23068*/;
assign _44593_ = _44584_ & _44592_ /*23066*/;
assign _44328_ = _44584_ ^ _44592_ /*23067*/;
assign _44590_ = _44591_ | _44593_ /*23064*/;
assign _44595_ = ~Q[14] /*23063*/;
assign _44594_ = _44595_ & D[40] /*23062*/;
assign _44597_ = _43881_ & _44594_ /*23057*/;
assign _44598_ = _43881_ ^ _44594_ /*23060*/;
assign _44599_ = _44590_ & _44598_ /*23058*/;
assign _44329_ = _44590_ ^ _44598_ /*23059*/;
assign _44596_ = _44597_ | _44599_ /*23056*/;
assign _44601_ = ~Q[14] /*23055*/;
assign _44600_ = _44601_ & D[41] /*23054*/;
assign _44603_ = _43882_ & _44600_ /*23049*/;
assign _44604_ = _43882_ ^ _44600_ /*23052*/;
assign _44605_ = _44596_ & _44604_ /*23050*/;
assign _44330_ = _44596_ ^ _44604_ /*23051*/;
assign _44602_ = _44603_ | _44605_ /*23048*/;
assign _44607_ = ~Q[14] /*23047*/;
assign _44606_ = _44607_ & D[42] /*23046*/;
assign _44609_ = _43883_ & _44606_ /*23041*/;
assign _44610_ = _43883_ ^ _44606_ /*23044*/;
assign _44611_ = _44602_ & _44610_ /*23042*/;
assign _44331_ = _44602_ ^ _44610_ /*23043*/;
assign _44608_ = _44609_ | _44611_ /*23040*/;
assign _44613_ = ~Q[14] /*23039*/;
assign _44612_ = _44613_ & D[43] /*23038*/;
assign _44615_ = _43884_ & _44612_ /*23033*/;
assign _44616_ = _43884_ ^ _44612_ /*23036*/;
assign _44617_ = _44608_ & _44616_ /*23034*/;
assign _44332_ = _44608_ ^ _44616_ /*23035*/;
assign _44614_ = _44615_ | _44617_ /*23032*/;
assign _44619_ = ~Q[14] /*23031*/;
assign _44618_ = _44619_ & D[44] /*23030*/;
assign _44621_ = _43885_ & _44618_ /*23025*/;
assign _44622_ = _43885_ ^ _44618_ /*23028*/;
assign _44623_ = _44614_ & _44622_ /*23026*/;
assign _44333_ = _44614_ ^ _44622_ /*23027*/;
assign _44620_ = _44621_ | _44623_ /*23024*/;
assign _44625_ = ~Q[14] /*23023*/;
assign _44624_ = _44625_ & D[45] /*23022*/;
assign _44627_ = _43886_ & _44624_ /*23017*/;
assign _44628_ = _43886_ ^ _44624_ /*23020*/;
assign _44629_ = _44620_ & _44628_ /*23018*/;
assign _44334_ = _44620_ ^ _44628_ /*23019*/;
assign _44626_ = _44627_ | _44629_ /*23016*/;
assign _44631_ = ~Q[14] /*23015*/;
assign _44630_ = _44631_ & D[46] /*23014*/;
assign _44633_ = _43887_ & _44630_ /*23009*/;
assign _44634_ = _43887_ ^ _44630_ /*23012*/;
assign _44635_ = _44626_ & _44634_ /*23010*/;
assign _44335_ = _44626_ ^ _44634_ /*23011*/;
assign _44632_ = _44633_ | _44635_ /*23008*/;
assign _44637_ = ~Q[14] /*23007*/;
assign _44636_ = _44637_ & D[47] /*23006*/;
assign _44639_ = _43888_ & _44636_ /*23001*/;
assign _44640_ = _43888_ ^ _44636_ /*23004*/;
assign _44641_ = _44632_ & _44640_ /*23002*/;
assign _44336_ = _44632_ ^ _44640_ /*23003*/;
assign _44638_ = _44639_ | _44641_ /*23000*/;
assign _44643_ = ~Q[14] /*22999*/;
assign _44642_ = _44643_ & D[48] /*22998*/;
assign _44645_ = _43889_ & _44642_ /*22993*/;
assign _44646_ = _43889_ ^ _44642_ /*22996*/;
assign _44647_ = _44638_ & _44646_ /*22994*/;
assign _44337_ = _44638_ ^ _44646_ /*22995*/;
assign _44644_ = _44645_ | _44647_ /*22992*/;
assign _44649_ = ~Q[14] /*22991*/;
assign _44648_ = _44649_ & D[49] /*22990*/;
assign _44651_ = _43890_ & _44648_ /*22985*/;
assign _44652_ = _43890_ ^ _44648_ /*22988*/;
assign _44653_ = _44644_ & _44652_ /*22986*/;
assign _44338_ = _44644_ ^ _44652_ /*22987*/;
assign _44650_ = _44651_ | _44653_ /*22984*/;
assign _44655_ = ~Q[14] /*22983*/;
assign _44654_ = _44655_ & D[50] /*22982*/;
assign _44657_ = _43891_ & _44654_ /*22977*/;
assign _44658_ = _43891_ ^ _44654_ /*22980*/;
assign _44659_ = _44650_ & _44658_ /*22978*/;
assign _44339_ = _44650_ ^ _44658_ /*22979*/;
assign _44656_ = _44657_ | _44659_ /*22976*/;
assign _44661_ = ~Q[14] /*22975*/;
assign _44660_ = _44661_ & D[51] /*22974*/;
assign _44663_ = _43892_ & _44660_ /*22969*/;
assign _44664_ = _43892_ ^ _44660_ /*22972*/;
assign _44665_ = _44656_ & _44664_ /*22970*/;
assign _44340_ = _44656_ ^ _44664_ /*22971*/;
assign _44662_ = _44663_ | _44665_ /*22968*/;
assign _44667_ = ~Q[14] /*22967*/;
assign _44666_ = _44667_ & D[52] /*22966*/;
assign _44669_ = _43893_ & _44666_ /*22961*/;
assign _44670_ = _43893_ ^ _44666_ /*22964*/;
assign _44671_ = _44662_ & _44670_ /*22962*/;
assign _44341_ = _44662_ ^ _44670_ /*22963*/;
assign _44668_ = _44669_ | _44671_ /*22960*/;
assign _44673_ = ~Q[14] /*22959*/;
assign _44672_ = _44673_ & D[53] /*22958*/;
assign _44675_ = _43894_ & _44672_ /*22953*/;
assign _44676_ = _43894_ ^ _44672_ /*22956*/;
assign _44677_ = _44668_ & _44676_ /*22954*/;
assign _44342_ = _44668_ ^ _44676_ /*22955*/;
assign _44674_ = _44675_ | _44677_ /*22952*/;
assign _44679_ = ~Q[14] /*22951*/;
assign _44678_ = _44679_ & D[54] /*22950*/;
assign _44681_ = _43895_ & _44678_ /*22945*/;
assign _44682_ = _43895_ ^ _44678_ /*22948*/;
assign _44683_ = _44674_ & _44682_ /*22946*/;
assign _44343_ = _44674_ ^ _44682_ /*22947*/;
assign _44680_ = _44681_ | _44683_ /*22944*/;
assign _44685_ = ~Q[14] /*22943*/;
assign _44684_ = _44685_ & D[55] /*22942*/;
assign _44687_ = _43896_ & _44684_ /*22937*/;
assign _44688_ = _43896_ ^ _44684_ /*22940*/;
assign _44689_ = _44680_ & _44688_ /*22938*/;
assign _44344_ = _44680_ ^ _44688_ /*22939*/;
assign _44686_ = _44687_ | _44689_ /*22936*/;
assign _44691_ = ~Q[14] /*22935*/;
assign _44690_ = _44691_ & D[56] /*22934*/;
assign _44693_ = _43897_ & _44690_ /*22929*/;
assign _44694_ = _43897_ ^ _44690_ /*22932*/;
assign _44695_ = _44686_ & _44694_ /*22930*/;
assign _44345_ = _44686_ ^ _44694_ /*22931*/;
assign _44692_ = _44693_ | _44695_ /*22928*/;
assign _44697_ = ~Q[14] /*22927*/;
assign _44696_ = _44697_ & D[57] /*22926*/;
assign _44699_ = _43898_ & _44696_ /*22921*/;
assign _44700_ = _43898_ ^ _44696_ /*22924*/;
assign _44701_ = _44692_ & _44700_ /*22922*/;
assign _44346_ = _44692_ ^ _44700_ /*22923*/;
assign _44698_ = _44699_ | _44701_ /*22920*/;
assign _44703_ = ~Q[14] /*22919*/;
assign _44702_ = _44703_ & D[58] /*22918*/;
assign _44705_ = _43899_ & _44702_ /*22913*/;
assign _44706_ = _43899_ ^ _44702_ /*22916*/;
assign _44707_ = _44698_ & _44706_ /*22914*/;
assign _44347_ = _44698_ ^ _44706_ /*22915*/;
assign _44704_ = _44705_ | _44707_ /*22912*/;
assign _44709_ = ~Q[14] /*22911*/;
assign _44708_ = _44709_ & D[59] /*22910*/;
assign _44711_ = _43900_ & _44708_ /*22905*/;
assign _44712_ = _43900_ ^ _44708_ /*22908*/;
assign _44713_ = _44704_ & _44712_ /*22906*/;
assign _44348_ = _44704_ ^ _44712_ /*22907*/;
assign _44710_ = _44711_ | _44713_ /*22904*/;
assign _44715_ = ~Q[14] /*22903*/;
assign _44714_ = _44715_ & D[60] /*22902*/;
assign _44717_ = _43901_ & _44714_ /*22897*/;
assign _44718_ = _43901_ ^ _44714_ /*22900*/;
assign _44719_ = _44710_ & _44718_ /*22898*/;
assign _44349_ = _44710_ ^ _44718_ /*22899*/;
assign _44716_ = _44717_ | _44719_ /*22896*/;
assign _44721_ = ~Q[14] /*22895*/;
assign _44720_ = _44721_ & D[61] /*22894*/;
assign _44723_ = _43902_ & _44720_ /*22889*/;
assign _44724_ = _43902_ ^ _44720_ /*22892*/;
assign _44725_ = _44716_ & _44724_ /*22890*/;
assign _44350_ = _44716_ ^ _44724_ /*22891*/;
assign _44722_ = _44723_ | _44725_ /*22888*/;
assign _44727_ = ~Q[14] /*22887*/;
assign _44726_ = _44727_ & D[62] /*22886*/;
assign _44729_ = _43903_ & _44726_ /*22881*/;
assign _44730_ = _43903_ ^ _44726_ /*22884*/;
assign _44731_ = _44722_ & _44730_ /*22882*/;
assign _44351_ = _44722_ ^ _44730_ /*22883*/;
assign _44728_ = _44729_ | _44731_ /*22880*/;
assign _44733_ = ~Q[14] /*22879*/;
assign _44732_ = _44733_ & zeroWire /*22878*/;
assign _44734_ = _43904_ ^ _44732_ /*22876*/;
assign _44352_ = _44734_ ^ _44728_ /*22875*/;
assign _44805_ = ~D[0] /*22621*/;
assign _44802_ = R_0[13] & _44805_ /*22617*/;
assign _44803_ = R_0[13] ^ _44805_ /*22620*/;
assign _44804_ = oneWire & _44803_ /*22618*/;
assign _44737_ = oneWire ^ _44803_ /*22619*/;
assign _44801_ = _44802_ | _44804_ /*22616*/;
assign _44810_ = ~D[1] /*22615*/;
assign _44807_ = _44289_ & _44810_ /*22611*/;
assign _44808_ = _44289_ ^ _44810_ /*22614*/;
assign _44809_ = _44801_ & _44808_ /*22612*/;
assign _44738_ = _44801_ ^ _44808_ /*22613*/;
assign _44806_ = _44807_ | _44809_ /*22610*/;
assign _44815_ = ~D[2] /*22609*/;
assign _44812_ = _44290_ & _44815_ /*22605*/;
assign _44813_ = _44290_ ^ _44815_ /*22608*/;
assign _44814_ = _44806_ & _44813_ /*22606*/;
assign _44739_ = _44806_ ^ _44813_ /*22607*/;
assign _44811_ = _44812_ | _44814_ /*22604*/;
assign _44820_ = ~D[3] /*22603*/;
assign _44817_ = _44291_ & _44820_ /*22599*/;
assign _44818_ = _44291_ ^ _44820_ /*22602*/;
assign _44819_ = _44811_ & _44818_ /*22600*/;
assign _44740_ = _44811_ ^ _44818_ /*22601*/;
assign _44816_ = _44817_ | _44819_ /*22598*/;
assign _44825_ = ~D[4] /*22597*/;
assign _44822_ = _44292_ & _44825_ /*22593*/;
assign _44823_ = _44292_ ^ _44825_ /*22596*/;
assign _44824_ = _44816_ & _44823_ /*22594*/;
assign _44741_ = _44816_ ^ _44823_ /*22595*/;
assign _44821_ = _44822_ | _44824_ /*22592*/;
assign _44830_ = ~D[5] /*22591*/;
assign _44827_ = _44293_ & _44830_ /*22587*/;
assign _44828_ = _44293_ ^ _44830_ /*22590*/;
assign _44829_ = _44821_ & _44828_ /*22588*/;
assign _44742_ = _44821_ ^ _44828_ /*22589*/;
assign _44826_ = _44827_ | _44829_ /*22586*/;
assign _44835_ = ~D[6] /*22585*/;
assign _44832_ = _44294_ & _44835_ /*22581*/;
assign _44833_ = _44294_ ^ _44835_ /*22584*/;
assign _44834_ = _44826_ & _44833_ /*22582*/;
assign _44743_ = _44826_ ^ _44833_ /*22583*/;
assign _44831_ = _44832_ | _44834_ /*22580*/;
assign _44840_ = ~D[7] /*22579*/;
assign _44837_ = _44295_ & _44840_ /*22575*/;
assign _44838_ = _44295_ ^ _44840_ /*22578*/;
assign _44839_ = _44831_ & _44838_ /*22576*/;
assign _44744_ = _44831_ ^ _44838_ /*22577*/;
assign _44836_ = _44837_ | _44839_ /*22574*/;
assign _44845_ = ~D[8] /*22573*/;
assign _44842_ = _44296_ & _44845_ /*22569*/;
assign _44843_ = _44296_ ^ _44845_ /*22572*/;
assign _44844_ = _44836_ & _44843_ /*22570*/;
assign _44745_ = _44836_ ^ _44843_ /*22571*/;
assign _44841_ = _44842_ | _44844_ /*22568*/;
assign _44850_ = ~D[9] /*22567*/;
assign _44847_ = _44297_ & _44850_ /*22563*/;
assign _44848_ = _44297_ ^ _44850_ /*22566*/;
assign _44849_ = _44841_ & _44848_ /*22564*/;
assign _44746_ = _44841_ ^ _44848_ /*22565*/;
assign _44846_ = _44847_ | _44849_ /*22562*/;
assign _44855_ = ~D[10] /*22561*/;
assign _44852_ = _44298_ & _44855_ /*22557*/;
assign _44853_ = _44298_ ^ _44855_ /*22560*/;
assign _44854_ = _44846_ & _44853_ /*22558*/;
assign _44747_ = _44846_ ^ _44853_ /*22559*/;
assign _44851_ = _44852_ | _44854_ /*22556*/;
assign _44860_ = ~D[11] /*22555*/;
assign _44857_ = _44299_ & _44860_ /*22551*/;
assign _44858_ = _44299_ ^ _44860_ /*22554*/;
assign _44859_ = _44851_ & _44858_ /*22552*/;
assign _44748_ = _44851_ ^ _44858_ /*22553*/;
assign _44856_ = _44857_ | _44859_ /*22550*/;
assign _44865_ = ~D[12] /*22549*/;
assign _44862_ = _44300_ & _44865_ /*22545*/;
assign _44863_ = _44300_ ^ _44865_ /*22548*/;
assign _44864_ = _44856_ & _44863_ /*22546*/;
assign _44749_ = _44856_ ^ _44863_ /*22547*/;
assign _44861_ = _44862_ | _44864_ /*22544*/;
assign _44870_ = ~D[13] /*22543*/;
assign _44867_ = _44301_ & _44870_ /*22539*/;
assign _44868_ = _44301_ ^ _44870_ /*22542*/;
assign _44869_ = _44861_ & _44868_ /*22540*/;
assign _44750_ = _44861_ ^ _44868_ /*22541*/;
assign _44866_ = _44867_ | _44869_ /*22538*/;
assign _44875_ = ~D[14] /*22537*/;
assign _44872_ = _44302_ & _44875_ /*22533*/;
assign _44873_ = _44302_ ^ _44875_ /*22536*/;
assign _44874_ = _44866_ & _44873_ /*22534*/;
assign _44751_ = _44866_ ^ _44873_ /*22535*/;
assign _44871_ = _44872_ | _44874_ /*22532*/;
assign _44880_ = ~D[15] /*22531*/;
assign _44877_ = _44303_ & _44880_ /*22527*/;
assign _44878_ = _44303_ ^ _44880_ /*22530*/;
assign _44879_ = _44871_ & _44878_ /*22528*/;
assign _44752_ = _44871_ ^ _44878_ /*22529*/;
assign _44876_ = _44877_ | _44879_ /*22526*/;
assign _44885_ = ~D[16] /*22525*/;
assign _44882_ = _44304_ & _44885_ /*22521*/;
assign _44883_ = _44304_ ^ _44885_ /*22524*/;
assign _44884_ = _44876_ & _44883_ /*22522*/;
assign _44753_ = _44876_ ^ _44883_ /*22523*/;
assign _44881_ = _44882_ | _44884_ /*22520*/;
assign _44890_ = ~D[17] /*22519*/;
assign _44887_ = _44305_ & _44890_ /*22515*/;
assign _44888_ = _44305_ ^ _44890_ /*22518*/;
assign _44889_ = _44881_ & _44888_ /*22516*/;
assign _44754_ = _44881_ ^ _44888_ /*22517*/;
assign _44886_ = _44887_ | _44889_ /*22514*/;
assign _44895_ = ~D[18] /*22513*/;
assign _44892_ = _44306_ & _44895_ /*22509*/;
assign _44893_ = _44306_ ^ _44895_ /*22512*/;
assign _44894_ = _44886_ & _44893_ /*22510*/;
assign _44755_ = _44886_ ^ _44893_ /*22511*/;
assign _44891_ = _44892_ | _44894_ /*22508*/;
assign _44900_ = ~D[19] /*22507*/;
assign _44897_ = _44307_ & _44900_ /*22503*/;
assign _44898_ = _44307_ ^ _44900_ /*22506*/;
assign _44899_ = _44891_ & _44898_ /*22504*/;
assign _44756_ = _44891_ ^ _44898_ /*22505*/;
assign _44896_ = _44897_ | _44899_ /*22502*/;
assign _44905_ = ~D[20] /*22501*/;
assign _44902_ = _44308_ & _44905_ /*22497*/;
assign _44903_ = _44308_ ^ _44905_ /*22500*/;
assign _44904_ = _44896_ & _44903_ /*22498*/;
assign _44757_ = _44896_ ^ _44903_ /*22499*/;
assign _44901_ = _44902_ | _44904_ /*22496*/;
assign _44910_ = ~D[21] /*22495*/;
assign _44907_ = _44309_ & _44910_ /*22491*/;
assign _44908_ = _44309_ ^ _44910_ /*22494*/;
assign _44909_ = _44901_ & _44908_ /*22492*/;
assign _44758_ = _44901_ ^ _44908_ /*22493*/;
assign _44906_ = _44907_ | _44909_ /*22490*/;
assign _44915_ = ~D[22] /*22489*/;
assign _44912_ = _44310_ & _44915_ /*22485*/;
assign _44913_ = _44310_ ^ _44915_ /*22488*/;
assign _44914_ = _44906_ & _44913_ /*22486*/;
assign _44759_ = _44906_ ^ _44913_ /*22487*/;
assign _44911_ = _44912_ | _44914_ /*22484*/;
assign _44920_ = ~D[23] /*22483*/;
assign _44917_ = _44311_ & _44920_ /*22479*/;
assign _44918_ = _44311_ ^ _44920_ /*22482*/;
assign _44919_ = _44911_ & _44918_ /*22480*/;
assign _44760_ = _44911_ ^ _44918_ /*22481*/;
assign _44916_ = _44917_ | _44919_ /*22478*/;
assign _44925_ = ~D[24] /*22477*/;
assign _44922_ = _44312_ & _44925_ /*22473*/;
assign _44923_ = _44312_ ^ _44925_ /*22476*/;
assign _44924_ = _44916_ & _44923_ /*22474*/;
assign _44761_ = _44916_ ^ _44923_ /*22475*/;
assign _44921_ = _44922_ | _44924_ /*22472*/;
assign _44930_ = ~D[25] /*22471*/;
assign _44927_ = _44313_ & _44930_ /*22467*/;
assign _44928_ = _44313_ ^ _44930_ /*22470*/;
assign _44929_ = _44921_ & _44928_ /*22468*/;
assign _44762_ = _44921_ ^ _44928_ /*22469*/;
assign _44926_ = _44927_ | _44929_ /*22466*/;
assign _44935_ = ~D[26] /*22465*/;
assign _44932_ = _44314_ & _44935_ /*22461*/;
assign _44933_ = _44314_ ^ _44935_ /*22464*/;
assign _44934_ = _44926_ & _44933_ /*22462*/;
assign _44763_ = _44926_ ^ _44933_ /*22463*/;
assign _44931_ = _44932_ | _44934_ /*22460*/;
assign _44940_ = ~D[27] /*22459*/;
assign _44937_ = _44315_ & _44940_ /*22455*/;
assign _44938_ = _44315_ ^ _44940_ /*22458*/;
assign _44939_ = _44931_ & _44938_ /*22456*/;
assign _44764_ = _44931_ ^ _44938_ /*22457*/;
assign _44936_ = _44937_ | _44939_ /*22454*/;
assign _44945_ = ~D[28] /*22453*/;
assign _44942_ = _44316_ & _44945_ /*22449*/;
assign _44943_ = _44316_ ^ _44945_ /*22452*/;
assign _44944_ = _44936_ & _44943_ /*22450*/;
assign _44765_ = _44936_ ^ _44943_ /*22451*/;
assign _44941_ = _44942_ | _44944_ /*22448*/;
assign _44950_ = ~D[29] /*22447*/;
assign _44947_ = _44317_ & _44950_ /*22443*/;
assign _44948_ = _44317_ ^ _44950_ /*22446*/;
assign _44949_ = _44941_ & _44948_ /*22444*/;
assign _44766_ = _44941_ ^ _44948_ /*22445*/;
assign _44946_ = _44947_ | _44949_ /*22442*/;
assign _44955_ = ~D[30] /*22441*/;
assign _44952_ = _44318_ & _44955_ /*22437*/;
assign _44953_ = _44318_ ^ _44955_ /*22440*/;
assign _44954_ = _44946_ & _44953_ /*22438*/;
assign _44767_ = _44946_ ^ _44953_ /*22439*/;
assign _44951_ = _44952_ | _44954_ /*22436*/;
assign _44960_ = ~D[31] /*22435*/;
assign _44957_ = _44319_ & _44960_ /*22431*/;
assign _44958_ = _44319_ ^ _44960_ /*22434*/;
assign _44959_ = _44951_ & _44958_ /*22432*/;
assign _44768_ = _44951_ ^ _44958_ /*22433*/;
assign _44956_ = _44957_ | _44959_ /*22430*/;
assign _44965_ = ~D[32] /*22429*/;
assign _44962_ = _44320_ & _44965_ /*22425*/;
assign _44963_ = _44320_ ^ _44965_ /*22428*/;
assign _44964_ = _44956_ & _44963_ /*22426*/;
assign _44769_ = _44956_ ^ _44963_ /*22427*/;
assign _44961_ = _44962_ | _44964_ /*22424*/;
assign _44970_ = ~D[33] /*22423*/;
assign _44967_ = _44321_ & _44970_ /*22419*/;
assign _44968_ = _44321_ ^ _44970_ /*22422*/;
assign _44969_ = _44961_ & _44968_ /*22420*/;
assign _44770_ = _44961_ ^ _44968_ /*22421*/;
assign _44966_ = _44967_ | _44969_ /*22418*/;
assign _44975_ = ~D[34] /*22417*/;
assign _44972_ = _44322_ & _44975_ /*22413*/;
assign _44973_ = _44322_ ^ _44975_ /*22416*/;
assign _44974_ = _44966_ & _44973_ /*22414*/;
assign _44771_ = _44966_ ^ _44973_ /*22415*/;
assign _44971_ = _44972_ | _44974_ /*22412*/;
assign _44980_ = ~D[35] /*22411*/;
assign _44977_ = _44323_ & _44980_ /*22407*/;
assign _44978_ = _44323_ ^ _44980_ /*22410*/;
assign _44979_ = _44971_ & _44978_ /*22408*/;
assign _44772_ = _44971_ ^ _44978_ /*22409*/;
assign _44976_ = _44977_ | _44979_ /*22406*/;
assign _44985_ = ~D[36] /*22405*/;
assign _44982_ = _44324_ & _44985_ /*22401*/;
assign _44983_ = _44324_ ^ _44985_ /*22404*/;
assign _44984_ = _44976_ & _44983_ /*22402*/;
assign _44773_ = _44976_ ^ _44983_ /*22403*/;
assign _44981_ = _44982_ | _44984_ /*22400*/;
assign _44990_ = ~D[37] /*22399*/;
assign _44987_ = _44325_ & _44990_ /*22395*/;
assign _44988_ = _44325_ ^ _44990_ /*22398*/;
assign _44989_ = _44981_ & _44988_ /*22396*/;
assign _44774_ = _44981_ ^ _44988_ /*22397*/;
assign _44986_ = _44987_ | _44989_ /*22394*/;
assign _44995_ = ~D[38] /*22393*/;
assign _44992_ = _44326_ & _44995_ /*22389*/;
assign _44993_ = _44326_ ^ _44995_ /*22392*/;
assign _44994_ = _44986_ & _44993_ /*22390*/;
assign _44775_ = _44986_ ^ _44993_ /*22391*/;
assign _44991_ = _44992_ | _44994_ /*22388*/;
assign _45000_ = ~D[39] /*22387*/;
assign _44997_ = _44327_ & _45000_ /*22383*/;
assign _44998_ = _44327_ ^ _45000_ /*22386*/;
assign _44999_ = _44991_ & _44998_ /*22384*/;
assign _44776_ = _44991_ ^ _44998_ /*22385*/;
assign _44996_ = _44997_ | _44999_ /*22382*/;
assign _45005_ = ~D[40] /*22381*/;
assign _45002_ = _44328_ & _45005_ /*22377*/;
assign _45003_ = _44328_ ^ _45005_ /*22380*/;
assign _45004_ = _44996_ & _45003_ /*22378*/;
assign _44777_ = _44996_ ^ _45003_ /*22379*/;
assign _45001_ = _45002_ | _45004_ /*22376*/;
assign _45010_ = ~D[41] /*22375*/;
assign _45007_ = _44329_ & _45010_ /*22371*/;
assign _45008_ = _44329_ ^ _45010_ /*22374*/;
assign _45009_ = _45001_ & _45008_ /*22372*/;
assign _44778_ = _45001_ ^ _45008_ /*22373*/;
assign _45006_ = _45007_ | _45009_ /*22370*/;
assign _45015_ = ~D[42] /*22369*/;
assign _45012_ = _44330_ & _45015_ /*22365*/;
assign _45013_ = _44330_ ^ _45015_ /*22368*/;
assign _45014_ = _45006_ & _45013_ /*22366*/;
assign _44779_ = _45006_ ^ _45013_ /*22367*/;
assign _45011_ = _45012_ | _45014_ /*22364*/;
assign _45020_ = ~D[43] /*22363*/;
assign _45017_ = _44331_ & _45020_ /*22359*/;
assign _45018_ = _44331_ ^ _45020_ /*22362*/;
assign _45019_ = _45011_ & _45018_ /*22360*/;
assign _44780_ = _45011_ ^ _45018_ /*22361*/;
assign _45016_ = _45017_ | _45019_ /*22358*/;
assign _45025_ = ~D[44] /*22357*/;
assign _45022_ = _44332_ & _45025_ /*22353*/;
assign _45023_ = _44332_ ^ _45025_ /*22356*/;
assign _45024_ = _45016_ & _45023_ /*22354*/;
assign _44781_ = _45016_ ^ _45023_ /*22355*/;
assign _45021_ = _45022_ | _45024_ /*22352*/;
assign _45030_ = ~D[45] /*22351*/;
assign _45027_ = _44333_ & _45030_ /*22347*/;
assign _45028_ = _44333_ ^ _45030_ /*22350*/;
assign _45029_ = _45021_ & _45028_ /*22348*/;
assign _44782_ = _45021_ ^ _45028_ /*22349*/;
assign _45026_ = _45027_ | _45029_ /*22346*/;
assign _45035_ = ~D[46] /*22345*/;
assign _45032_ = _44334_ & _45035_ /*22341*/;
assign _45033_ = _44334_ ^ _45035_ /*22344*/;
assign _45034_ = _45026_ & _45033_ /*22342*/;
assign _44783_ = _45026_ ^ _45033_ /*22343*/;
assign _45031_ = _45032_ | _45034_ /*22340*/;
assign _45040_ = ~D[47] /*22339*/;
assign _45037_ = _44335_ & _45040_ /*22335*/;
assign _45038_ = _44335_ ^ _45040_ /*22338*/;
assign _45039_ = _45031_ & _45038_ /*22336*/;
assign _44784_ = _45031_ ^ _45038_ /*22337*/;
assign _45036_ = _45037_ | _45039_ /*22334*/;
assign _45045_ = ~D[48] /*22333*/;
assign _45042_ = _44336_ & _45045_ /*22329*/;
assign _45043_ = _44336_ ^ _45045_ /*22332*/;
assign _45044_ = _45036_ & _45043_ /*22330*/;
assign _44785_ = _45036_ ^ _45043_ /*22331*/;
assign _45041_ = _45042_ | _45044_ /*22328*/;
assign _45050_ = ~D[49] /*22327*/;
assign _45047_ = _44337_ & _45050_ /*22323*/;
assign _45048_ = _44337_ ^ _45050_ /*22326*/;
assign _45049_ = _45041_ & _45048_ /*22324*/;
assign _44786_ = _45041_ ^ _45048_ /*22325*/;
assign _45046_ = _45047_ | _45049_ /*22322*/;
assign _45055_ = ~D[50] /*22321*/;
assign _45052_ = _44338_ & _45055_ /*22317*/;
assign _45053_ = _44338_ ^ _45055_ /*22320*/;
assign _45054_ = _45046_ & _45053_ /*22318*/;
assign _44787_ = _45046_ ^ _45053_ /*22319*/;
assign _45051_ = _45052_ | _45054_ /*22316*/;
assign _45060_ = ~D[51] /*22315*/;
assign _45057_ = _44339_ & _45060_ /*22311*/;
assign _45058_ = _44339_ ^ _45060_ /*22314*/;
assign _45059_ = _45051_ & _45058_ /*22312*/;
assign _44788_ = _45051_ ^ _45058_ /*22313*/;
assign _45056_ = _45057_ | _45059_ /*22310*/;
assign _45065_ = ~D[52] /*22309*/;
assign _45062_ = _44340_ & _45065_ /*22305*/;
assign _45063_ = _44340_ ^ _45065_ /*22308*/;
assign _45064_ = _45056_ & _45063_ /*22306*/;
assign _44789_ = _45056_ ^ _45063_ /*22307*/;
assign _45061_ = _45062_ | _45064_ /*22304*/;
assign _45070_ = ~D[53] /*22303*/;
assign _45067_ = _44341_ & _45070_ /*22299*/;
assign _45068_ = _44341_ ^ _45070_ /*22302*/;
assign _45069_ = _45061_ & _45068_ /*22300*/;
assign _44790_ = _45061_ ^ _45068_ /*22301*/;
assign _45066_ = _45067_ | _45069_ /*22298*/;
assign _45075_ = ~D[54] /*22297*/;
assign _45072_ = _44342_ & _45075_ /*22293*/;
assign _45073_ = _44342_ ^ _45075_ /*22296*/;
assign _45074_ = _45066_ & _45073_ /*22294*/;
assign _44791_ = _45066_ ^ _45073_ /*22295*/;
assign _45071_ = _45072_ | _45074_ /*22292*/;
assign _45080_ = ~D[55] /*22291*/;
assign _45077_ = _44343_ & _45080_ /*22287*/;
assign _45078_ = _44343_ ^ _45080_ /*22290*/;
assign _45079_ = _45071_ & _45078_ /*22288*/;
assign _44792_ = _45071_ ^ _45078_ /*22289*/;
assign _45076_ = _45077_ | _45079_ /*22286*/;
assign _45085_ = ~D[56] /*22285*/;
assign _45082_ = _44344_ & _45085_ /*22281*/;
assign _45083_ = _44344_ ^ _45085_ /*22284*/;
assign _45084_ = _45076_ & _45083_ /*22282*/;
assign _44793_ = _45076_ ^ _45083_ /*22283*/;
assign _45081_ = _45082_ | _45084_ /*22280*/;
assign _45090_ = ~D[57] /*22279*/;
assign _45087_ = _44345_ & _45090_ /*22275*/;
assign _45088_ = _44345_ ^ _45090_ /*22278*/;
assign _45089_ = _45081_ & _45088_ /*22276*/;
assign _44794_ = _45081_ ^ _45088_ /*22277*/;
assign _45086_ = _45087_ | _45089_ /*22274*/;
assign _45095_ = ~D[58] /*22273*/;
assign _45092_ = _44346_ & _45095_ /*22269*/;
assign _45093_ = _44346_ ^ _45095_ /*22272*/;
assign _45094_ = _45086_ & _45093_ /*22270*/;
assign _44795_ = _45086_ ^ _45093_ /*22271*/;
assign _45091_ = _45092_ | _45094_ /*22268*/;
assign _45100_ = ~D[59] /*22267*/;
assign _45097_ = _44347_ & _45100_ /*22263*/;
assign _45098_ = _44347_ ^ _45100_ /*22266*/;
assign _45099_ = _45091_ & _45098_ /*22264*/;
assign _44796_ = _45091_ ^ _45098_ /*22265*/;
assign _45096_ = _45097_ | _45099_ /*22262*/;
assign _45105_ = ~D[60] /*22261*/;
assign _45102_ = _44348_ & _45105_ /*22257*/;
assign _45103_ = _44348_ ^ _45105_ /*22260*/;
assign _45104_ = _45096_ & _45103_ /*22258*/;
assign _44797_ = _45096_ ^ _45103_ /*22259*/;
assign _45101_ = _45102_ | _45104_ /*22256*/;
assign _45110_ = ~D[61] /*22255*/;
assign _45107_ = _44349_ & _45110_ /*22251*/;
assign _45108_ = _44349_ ^ _45110_ /*22254*/;
assign _45109_ = _45101_ & _45108_ /*22252*/;
assign _44798_ = _45101_ ^ _45108_ /*22253*/;
assign _45106_ = _45107_ | _45109_ /*22250*/;
assign _45115_ = ~D[62] /*22249*/;
assign _45112_ = _44350_ & _45115_ /*22245*/;
assign _45113_ = _44350_ ^ _45115_ /*22248*/;
assign _45114_ = _45106_ & _45113_ /*22246*/;
assign _44799_ = _45106_ ^ _45113_ /*22247*/;
assign _45111_ = _45112_ | _45114_ /*22244*/;
assign _45116_ = _44351_ & oneWire /*22239*/;
assign _45117_ = _44351_ ^ oneWire /*22242*/;
assign _45118_ = _45111_ & _45117_ /*22240*/;
assign _44800_ = _45111_ ^ _45117_ /*22241*/;
assign Q[13] = _45116_ | _45118_ /*22238*/;
assign _45251_ = ~Q[13] /*21853*/;
assign _45250_ = _45251_ & D[0] /*21852*/;
assign _45253_ = _44737_ & _45250_ /*21847*/;
assign _45254_ = _44737_ ^ _45250_ /*21850*/;
assign _45255_ = zeroWire & _45254_ /*21848*/;
assign _45185_ = zeroWire ^ _45254_ /*21849*/;
assign _45252_ = _45253_ | _45255_ /*21846*/;
assign _45257_ = ~Q[13] /*21845*/;
assign _45256_ = _45257_ & D[1] /*21844*/;
assign _45259_ = _44738_ & _45256_ /*21839*/;
assign _45260_ = _44738_ ^ _45256_ /*21842*/;
assign _45261_ = _45252_ & _45260_ /*21840*/;
assign _45186_ = _45252_ ^ _45260_ /*21841*/;
assign _45258_ = _45259_ | _45261_ /*21838*/;
assign _45263_ = ~Q[13] /*21837*/;
assign _45262_ = _45263_ & D[2] /*21836*/;
assign _45265_ = _44739_ & _45262_ /*21831*/;
assign _45266_ = _44739_ ^ _45262_ /*21834*/;
assign _45267_ = _45258_ & _45266_ /*21832*/;
assign _45187_ = _45258_ ^ _45266_ /*21833*/;
assign _45264_ = _45265_ | _45267_ /*21830*/;
assign _45269_ = ~Q[13] /*21829*/;
assign _45268_ = _45269_ & D[3] /*21828*/;
assign _45271_ = _44740_ & _45268_ /*21823*/;
assign _45272_ = _44740_ ^ _45268_ /*21826*/;
assign _45273_ = _45264_ & _45272_ /*21824*/;
assign _45188_ = _45264_ ^ _45272_ /*21825*/;
assign _45270_ = _45271_ | _45273_ /*21822*/;
assign _45275_ = ~Q[13] /*21821*/;
assign _45274_ = _45275_ & D[4] /*21820*/;
assign _45277_ = _44741_ & _45274_ /*21815*/;
assign _45278_ = _44741_ ^ _45274_ /*21818*/;
assign _45279_ = _45270_ & _45278_ /*21816*/;
assign _45189_ = _45270_ ^ _45278_ /*21817*/;
assign _45276_ = _45277_ | _45279_ /*21814*/;
assign _45281_ = ~Q[13] /*21813*/;
assign _45280_ = _45281_ & D[5] /*21812*/;
assign _45283_ = _44742_ & _45280_ /*21807*/;
assign _45284_ = _44742_ ^ _45280_ /*21810*/;
assign _45285_ = _45276_ & _45284_ /*21808*/;
assign _45190_ = _45276_ ^ _45284_ /*21809*/;
assign _45282_ = _45283_ | _45285_ /*21806*/;
assign _45287_ = ~Q[13] /*21805*/;
assign _45286_ = _45287_ & D[6] /*21804*/;
assign _45289_ = _44743_ & _45286_ /*21799*/;
assign _45290_ = _44743_ ^ _45286_ /*21802*/;
assign _45291_ = _45282_ & _45290_ /*21800*/;
assign _45191_ = _45282_ ^ _45290_ /*21801*/;
assign _45288_ = _45289_ | _45291_ /*21798*/;
assign _45293_ = ~Q[13] /*21797*/;
assign _45292_ = _45293_ & D[7] /*21796*/;
assign _45295_ = _44744_ & _45292_ /*21791*/;
assign _45296_ = _44744_ ^ _45292_ /*21794*/;
assign _45297_ = _45288_ & _45296_ /*21792*/;
assign _45192_ = _45288_ ^ _45296_ /*21793*/;
assign _45294_ = _45295_ | _45297_ /*21790*/;
assign _45299_ = ~Q[13] /*21789*/;
assign _45298_ = _45299_ & D[8] /*21788*/;
assign _45301_ = _44745_ & _45298_ /*21783*/;
assign _45302_ = _44745_ ^ _45298_ /*21786*/;
assign _45303_ = _45294_ & _45302_ /*21784*/;
assign _45193_ = _45294_ ^ _45302_ /*21785*/;
assign _45300_ = _45301_ | _45303_ /*21782*/;
assign _45305_ = ~Q[13] /*21781*/;
assign _45304_ = _45305_ & D[9] /*21780*/;
assign _45307_ = _44746_ & _45304_ /*21775*/;
assign _45308_ = _44746_ ^ _45304_ /*21778*/;
assign _45309_ = _45300_ & _45308_ /*21776*/;
assign _45194_ = _45300_ ^ _45308_ /*21777*/;
assign _45306_ = _45307_ | _45309_ /*21774*/;
assign _45311_ = ~Q[13] /*21773*/;
assign _45310_ = _45311_ & D[10] /*21772*/;
assign _45313_ = _44747_ & _45310_ /*21767*/;
assign _45314_ = _44747_ ^ _45310_ /*21770*/;
assign _45315_ = _45306_ & _45314_ /*21768*/;
assign _45195_ = _45306_ ^ _45314_ /*21769*/;
assign _45312_ = _45313_ | _45315_ /*21766*/;
assign _45317_ = ~Q[13] /*21765*/;
assign _45316_ = _45317_ & D[11] /*21764*/;
assign _45319_ = _44748_ & _45316_ /*21759*/;
assign _45320_ = _44748_ ^ _45316_ /*21762*/;
assign _45321_ = _45312_ & _45320_ /*21760*/;
assign _45196_ = _45312_ ^ _45320_ /*21761*/;
assign _45318_ = _45319_ | _45321_ /*21758*/;
assign _45323_ = ~Q[13] /*21757*/;
assign _45322_ = _45323_ & D[12] /*21756*/;
assign _45325_ = _44749_ & _45322_ /*21751*/;
assign _45326_ = _44749_ ^ _45322_ /*21754*/;
assign _45327_ = _45318_ & _45326_ /*21752*/;
assign _45197_ = _45318_ ^ _45326_ /*21753*/;
assign _45324_ = _45325_ | _45327_ /*21750*/;
assign _45329_ = ~Q[13] /*21749*/;
assign _45328_ = _45329_ & D[13] /*21748*/;
assign _45331_ = _44750_ & _45328_ /*21743*/;
assign _45332_ = _44750_ ^ _45328_ /*21746*/;
assign _45333_ = _45324_ & _45332_ /*21744*/;
assign _45198_ = _45324_ ^ _45332_ /*21745*/;
assign _45330_ = _45331_ | _45333_ /*21742*/;
assign _45335_ = ~Q[13] /*21741*/;
assign _45334_ = _45335_ & D[14] /*21740*/;
assign _45337_ = _44751_ & _45334_ /*21735*/;
assign _45338_ = _44751_ ^ _45334_ /*21738*/;
assign _45339_ = _45330_ & _45338_ /*21736*/;
assign _45199_ = _45330_ ^ _45338_ /*21737*/;
assign _45336_ = _45337_ | _45339_ /*21734*/;
assign _45341_ = ~Q[13] /*21733*/;
assign _45340_ = _45341_ & D[15] /*21732*/;
assign _45343_ = _44752_ & _45340_ /*21727*/;
assign _45344_ = _44752_ ^ _45340_ /*21730*/;
assign _45345_ = _45336_ & _45344_ /*21728*/;
assign _45200_ = _45336_ ^ _45344_ /*21729*/;
assign _45342_ = _45343_ | _45345_ /*21726*/;
assign _45347_ = ~Q[13] /*21725*/;
assign _45346_ = _45347_ & D[16] /*21724*/;
assign _45349_ = _44753_ & _45346_ /*21719*/;
assign _45350_ = _44753_ ^ _45346_ /*21722*/;
assign _45351_ = _45342_ & _45350_ /*21720*/;
assign _45201_ = _45342_ ^ _45350_ /*21721*/;
assign _45348_ = _45349_ | _45351_ /*21718*/;
assign _45353_ = ~Q[13] /*21717*/;
assign _45352_ = _45353_ & D[17] /*21716*/;
assign _45355_ = _44754_ & _45352_ /*21711*/;
assign _45356_ = _44754_ ^ _45352_ /*21714*/;
assign _45357_ = _45348_ & _45356_ /*21712*/;
assign _45202_ = _45348_ ^ _45356_ /*21713*/;
assign _45354_ = _45355_ | _45357_ /*21710*/;
assign _45359_ = ~Q[13] /*21709*/;
assign _45358_ = _45359_ & D[18] /*21708*/;
assign _45361_ = _44755_ & _45358_ /*21703*/;
assign _45362_ = _44755_ ^ _45358_ /*21706*/;
assign _45363_ = _45354_ & _45362_ /*21704*/;
assign _45203_ = _45354_ ^ _45362_ /*21705*/;
assign _45360_ = _45361_ | _45363_ /*21702*/;
assign _45365_ = ~Q[13] /*21701*/;
assign _45364_ = _45365_ & D[19] /*21700*/;
assign _45367_ = _44756_ & _45364_ /*21695*/;
assign _45368_ = _44756_ ^ _45364_ /*21698*/;
assign _45369_ = _45360_ & _45368_ /*21696*/;
assign _45204_ = _45360_ ^ _45368_ /*21697*/;
assign _45366_ = _45367_ | _45369_ /*21694*/;
assign _45371_ = ~Q[13] /*21693*/;
assign _45370_ = _45371_ & D[20] /*21692*/;
assign _45373_ = _44757_ & _45370_ /*21687*/;
assign _45374_ = _44757_ ^ _45370_ /*21690*/;
assign _45375_ = _45366_ & _45374_ /*21688*/;
assign _45205_ = _45366_ ^ _45374_ /*21689*/;
assign _45372_ = _45373_ | _45375_ /*21686*/;
assign _45377_ = ~Q[13] /*21685*/;
assign _45376_ = _45377_ & D[21] /*21684*/;
assign _45379_ = _44758_ & _45376_ /*21679*/;
assign _45380_ = _44758_ ^ _45376_ /*21682*/;
assign _45381_ = _45372_ & _45380_ /*21680*/;
assign _45206_ = _45372_ ^ _45380_ /*21681*/;
assign _45378_ = _45379_ | _45381_ /*21678*/;
assign _45383_ = ~Q[13] /*21677*/;
assign _45382_ = _45383_ & D[22] /*21676*/;
assign _45385_ = _44759_ & _45382_ /*21671*/;
assign _45386_ = _44759_ ^ _45382_ /*21674*/;
assign _45387_ = _45378_ & _45386_ /*21672*/;
assign _45207_ = _45378_ ^ _45386_ /*21673*/;
assign _45384_ = _45385_ | _45387_ /*21670*/;
assign _45389_ = ~Q[13] /*21669*/;
assign _45388_ = _45389_ & D[23] /*21668*/;
assign _45391_ = _44760_ & _45388_ /*21663*/;
assign _45392_ = _44760_ ^ _45388_ /*21666*/;
assign _45393_ = _45384_ & _45392_ /*21664*/;
assign _45208_ = _45384_ ^ _45392_ /*21665*/;
assign _45390_ = _45391_ | _45393_ /*21662*/;
assign _45395_ = ~Q[13] /*21661*/;
assign _45394_ = _45395_ & D[24] /*21660*/;
assign _45397_ = _44761_ & _45394_ /*21655*/;
assign _45398_ = _44761_ ^ _45394_ /*21658*/;
assign _45399_ = _45390_ & _45398_ /*21656*/;
assign _45209_ = _45390_ ^ _45398_ /*21657*/;
assign _45396_ = _45397_ | _45399_ /*21654*/;
assign _45401_ = ~Q[13] /*21653*/;
assign _45400_ = _45401_ & D[25] /*21652*/;
assign _45403_ = _44762_ & _45400_ /*21647*/;
assign _45404_ = _44762_ ^ _45400_ /*21650*/;
assign _45405_ = _45396_ & _45404_ /*21648*/;
assign _45210_ = _45396_ ^ _45404_ /*21649*/;
assign _45402_ = _45403_ | _45405_ /*21646*/;
assign _45407_ = ~Q[13] /*21645*/;
assign _45406_ = _45407_ & D[26] /*21644*/;
assign _45409_ = _44763_ & _45406_ /*21639*/;
assign _45410_ = _44763_ ^ _45406_ /*21642*/;
assign _45411_ = _45402_ & _45410_ /*21640*/;
assign _45211_ = _45402_ ^ _45410_ /*21641*/;
assign _45408_ = _45409_ | _45411_ /*21638*/;
assign _45413_ = ~Q[13] /*21637*/;
assign _45412_ = _45413_ & D[27] /*21636*/;
assign _45415_ = _44764_ & _45412_ /*21631*/;
assign _45416_ = _44764_ ^ _45412_ /*21634*/;
assign _45417_ = _45408_ & _45416_ /*21632*/;
assign _45212_ = _45408_ ^ _45416_ /*21633*/;
assign _45414_ = _45415_ | _45417_ /*21630*/;
assign _45419_ = ~Q[13] /*21629*/;
assign _45418_ = _45419_ & D[28] /*21628*/;
assign _45421_ = _44765_ & _45418_ /*21623*/;
assign _45422_ = _44765_ ^ _45418_ /*21626*/;
assign _45423_ = _45414_ & _45422_ /*21624*/;
assign _45213_ = _45414_ ^ _45422_ /*21625*/;
assign _45420_ = _45421_ | _45423_ /*21622*/;
assign _45425_ = ~Q[13] /*21621*/;
assign _45424_ = _45425_ & D[29] /*21620*/;
assign _45427_ = _44766_ & _45424_ /*21615*/;
assign _45428_ = _44766_ ^ _45424_ /*21618*/;
assign _45429_ = _45420_ & _45428_ /*21616*/;
assign _45214_ = _45420_ ^ _45428_ /*21617*/;
assign _45426_ = _45427_ | _45429_ /*21614*/;
assign _45431_ = ~Q[13] /*21613*/;
assign _45430_ = _45431_ & D[30] /*21612*/;
assign _45433_ = _44767_ & _45430_ /*21607*/;
assign _45434_ = _44767_ ^ _45430_ /*21610*/;
assign _45435_ = _45426_ & _45434_ /*21608*/;
assign _45215_ = _45426_ ^ _45434_ /*21609*/;
assign _45432_ = _45433_ | _45435_ /*21606*/;
assign _45437_ = ~Q[13] /*21605*/;
assign _45436_ = _45437_ & D[31] /*21604*/;
assign _45439_ = _44768_ & _45436_ /*21599*/;
assign _45440_ = _44768_ ^ _45436_ /*21602*/;
assign _45441_ = _45432_ & _45440_ /*21600*/;
assign _45216_ = _45432_ ^ _45440_ /*21601*/;
assign _45438_ = _45439_ | _45441_ /*21598*/;
assign _45443_ = ~Q[13] /*21597*/;
assign _45442_ = _45443_ & D[32] /*21596*/;
assign _45445_ = _44769_ & _45442_ /*21591*/;
assign _45446_ = _44769_ ^ _45442_ /*21594*/;
assign _45447_ = _45438_ & _45446_ /*21592*/;
assign _45217_ = _45438_ ^ _45446_ /*21593*/;
assign _45444_ = _45445_ | _45447_ /*21590*/;
assign _45449_ = ~Q[13] /*21589*/;
assign _45448_ = _45449_ & D[33] /*21588*/;
assign _45451_ = _44770_ & _45448_ /*21583*/;
assign _45452_ = _44770_ ^ _45448_ /*21586*/;
assign _45453_ = _45444_ & _45452_ /*21584*/;
assign _45218_ = _45444_ ^ _45452_ /*21585*/;
assign _45450_ = _45451_ | _45453_ /*21582*/;
assign _45455_ = ~Q[13] /*21581*/;
assign _45454_ = _45455_ & D[34] /*21580*/;
assign _45457_ = _44771_ & _45454_ /*21575*/;
assign _45458_ = _44771_ ^ _45454_ /*21578*/;
assign _45459_ = _45450_ & _45458_ /*21576*/;
assign _45219_ = _45450_ ^ _45458_ /*21577*/;
assign _45456_ = _45457_ | _45459_ /*21574*/;
assign _45461_ = ~Q[13] /*21573*/;
assign _45460_ = _45461_ & D[35] /*21572*/;
assign _45463_ = _44772_ & _45460_ /*21567*/;
assign _45464_ = _44772_ ^ _45460_ /*21570*/;
assign _45465_ = _45456_ & _45464_ /*21568*/;
assign _45220_ = _45456_ ^ _45464_ /*21569*/;
assign _45462_ = _45463_ | _45465_ /*21566*/;
assign _45467_ = ~Q[13] /*21565*/;
assign _45466_ = _45467_ & D[36] /*21564*/;
assign _45469_ = _44773_ & _45466_ /*21559*/;
assign _45470_ = _44773_ ^ _45466_ /*21562*/;
assign _45471_ = _45462_ & _45470_ /*21560*/;
assign _45221_ = _45462_ ^ _45470_ /*21561*/;
assign _45468_ = _45469_ | _45471_ /*21558*/;
assign _45473_ = ~Q[13] /*21557*/;
assign _45472_ = _45473_ & D[37] /*21556*/;
assign _45475_ = _44774_ & _45472_ /*21551*/;
assign _45476_ = _44774_ ^ _45472_ /*21554*/;
assign _45477_ = _45468_ & _45476_ /*21552*/;
assign _45222_ = _45468_ ^ _45476_ /*21553*/;
assign _45474_ = _45475_ | _45477_ /*21550*/;
assign _45479_ = ~Q[13] /*21549*/;
assign _45478_ = _45479_ & D[38] /*21548*/;
assign _45481_ = _44775_ & _45478_ /*21543*/;
assign _45482_ = _44775_ ^ _45478_ /*21546*/;
assign _45483_ = _45474_ & _45482_ /*21544*/;
assign _45223_ = _45474_ ^ _45482_ /*21545*/;
assign _45480_ = _45481_ | _45483_ /*21542*/;
assign _45485_ = ~Q[13] /*21541*/;
assign _45484_ = _45485_ & D[39] /*21540*/;
assign _45487_ = _44776_ & _45484_ /*21535*/;
assign _45488_ = _44776_ ^ _45484_ /*21538*/;
assign _45489_ = _45480_ & _45488_ /*21536*/;
assign _45224_ = _45480_ ^ _45488_ /*21537*/;
assign _45486_ = _45487_ | _45489_ /*21534*/;
assign _45491_ = ~Q[13] /*21533*/;
assign _45490_ = _45491_ & D[40] /*21532*/;
assign _45493_ = _44777_ & _45490_ /*21527*/;
assign _45494_ = _44777_ ^ _45490_ /*21530*/;
assign _45495_ = _45486_ & _45494_ /*21528*/;
assign _45225_ = _45486_ ^ _45494_ /*21529*/;
assign _45492_ = _45493_ | _45495_ /*21526*/;
assign _45497_ = ~Q[13] /*21525*/;
assign _45496_ = _45497_ & D[41] /*21524*/;
assign _45499_ = _44778_ & _45496_ /*21519*/;
assign _45500_ = _44778_ ^ _45496_ /*21522*/;
assign _45501_ = _45492_ & _45500_ /*21520*/;
assign _45226_ = _45492_ ^ _45500_ /*21521*/;
assign _45498_ = _45499_ | _45501_ /*21518*/;
assign _45503_ = ~Q[13] /*21517*/;
assign _45502_ = _45503_ & D[42] /*21516*/;
assign _45505_ = _44779_ & _45502_ /*21511*/;
assign _45506_ = _44779_ ^ _45502_ /*21514*/;
assign _45507_ = _45498_ & _45506_ /*21512*/;
assign _45227_ = _45498_ ^ _45506_ /*21513*/;
assign _45504_ = _45505_ | _45507_ /*21510*/;
assign _45509_ = ~Q[13] /*21509*/;
assign _45508_ = _45509_ & D[43] /*21508*/;
assign _45511_ = _44780_ & _45508_ /*21503*/;
assign _45512_ = _44780_ ^ _45508_ /*21506*/;
assign _45513_ = _45504_ & _45512_ /*21504*/;
assign _45228_ = _45504_ ^ _45512_ /*21505*/;
assign _45510_ = _45511_ | _45513_ /*21502*/;
assign _45515_ = ~Q[13] /*21501*/;
assign _45514_ = _45515_ & D[44] /*21500*/;
assign _45517_ = _44781_ & _45514_ /*21495*/;
assign _45518_ = _44781_ ^ _45514_ /*21498*/;
assign _45519_ = _45510_ & _45518_ /*21496*/;
assign _45229_ = _45510_ ^ _45518_ /*21497*/;
assign _45516_ = _45517_ | _45519_ /*21494*/;
assign _45521_ = ~Q[13] /*21493*/;
assign _45520_ = _45521_ & D[45] /*21492*/;
assign _45523_ = _44782_ & _45520_ /*21487*/;
assign _45524_ = _44782_ ^ _45520_ /*21490*/;
assign _45525_ = _45516_ & _45524_ /*21488*/;
assign _45230_ = _45516_ ^ _45524_ /*21489*/;
assign _45522_ = _45523_ | _45525_ /*21486*/;
assign _45527_ = ~Q[13] /*21485*/;
assign _45526_ = _45527_ & D[46] /*21484*/;
assign _45529_ = _44783_ & _45526_ /*21479*/;
assign _45530_ = _44783_ ^ _45526_ /*21482*/;
assign _45531_ = _45522_ & _45530_ /*21480*/;
assign _45231_ = _45522_ ^ _45530_ /*21481*/;
assign _45528_ = _45529_ | _45531_ /*21478*/;
assign _45533_ = ~Q[13] /*21477*/;
assign _45532_ = _45533_ & D[47] /*21476*/;
assign _45535_ = _44784_ & _45532_ /*21471*/;
assign _45536_ = _44784_ ^ _45532_ /*21474*/;
assign _45537_ = _45528_ & _45536_ /*21472*/;
assign _45232_ = _45528_ ^ _45536_ /*21473*/;
assign _45534_ = _45535_ | _45537_ /*21470*/;
assign _45539_ = ~Q[13] /*21469*/;
assign _45538_ = _45539_ & D[48] /*21468*/;
assign _45541_ = _44785_ & _45538_ /*21463*/;
assign _45542_ = _44785_ ^ _45538_ /*21466*/;
assign _45543_ = _45534_ & _45542_ /*21464*/;
assign _45233_ = _45534_ ^ _45542_ /*21465*/;
assign _45540_ = _45541_ | _45543_ /*21462*/;
assign _45545_ = ~Q[13] /*21461*/;
assign _45544_ = _45545_ & D[49] /*21460*/;
assign _45547_ = _44786_ & _45544_ /*21455*/;
assign _45548_ = _44786_ ^ _45544_ /*21458*/;
assign _45549_ = _45540_ & _45548_ /*21456*/;
assign _45234_ = _45540_ ^ _45548_ /*21457*/;
assign _45546_ = _45547_ | _45549_ /*21454*/;
assign _45551_ = ~Q[13] /*21453*/;
assign _45550_ = _45551_ & D[50] /*21452*/;
assign _45553_ = _44787_ & _45550_ /*21447*/;
assign _45554_ = _44787_ ^ _45550_ /*21450*/;
assign _45555_ = _45546_ & _45554_ /*21448*/;
assign _45235_ = _45546_ ^ _45554_ /*21449*/;
assign _45552_ = _45553_ | _45555_ /*21446*/;
assign _45557_ = ~Q[13] /*21445*/;
assign _45556_ = _45557_ & D[51] /*21444*/;
assign _45559_ = _44788_ & _45556_ /*21439*/;
assign _45560_ = _44788_ ^ _45556_ /*21442*/;
assign _45561_ = _45552_ & _45560_ /*21440*/;
assign _45236_ = _45552_ ^ _45560_ /*21441*/;
assign _45558_ = _45559_ | _45561_ /*21438*/;
assign _45563_ = ~Q[13] /*21437*/;
assign _45562_ = _45563_ & D[52] /*21436*/;
assign _45565_ = _44789_ & _45562_ /*21431*/;
assign _45566_ = _44789_ ^ _45562_ /*21434*/;
assign _45567_ = _45558_ & _45566_ /*21432*/;
assign _45237_ = _45558_ ^ _45566_ /*21433*/;
assign _45564_ = _45565_ | _45567_ /*21430*/;
assign _45569_ = ~Q[13] /*21429*/;
assign _45568_ = _45569_ & D[53] /*21428*/;
assign _45571_ = _44790_ & _45568_ /*21423*/;
assign _45572_ = _44790_ ^ _45568_ /*21426*/;
assign _45573_ = _45564_ & _45572_ /*21424*/;
assign _45238_ = _45564_ ^ _45572_ /*21425*/;
assign _45570_ = _45571_ | _45573_ /*21422*/;
assign _45575_ = ~Q[13] /*21421*/;
assign _45574_ = _45575_ & D[54] /*21420*/;
assign _45577_ = _44791_ & _45574_ /*21415*/;
assign _45578_ = _44791_ ^ _45574_ /*21418*/;
assign _45579_ = _45570_ & _45578_ /*21416*/;
assign _45239_ = _45570_ ^ _45578_ /*21417*/;
assign _45576_ = _45577_ | _45579_ /*21414*/;
assign _45581_ = ~Q[13] /*21413*/;
assign _45580_ = _45581_ & D[55] /*21412*/;
assign _45583_ = _44792_ & _45580_ /*21407*/;
assign _45584_ = _44792_ ^ _45580_ /*21410*/;
assign _45585_ = _45576_ & _45584_ /*21408*/;
assign _45240_ = _45576_ ^ _45584_ /*21409*/;
assign _45582_ = _45583_ | _45585_ /*21406*/;
assign _45587_ = ~Q[13] /*21405*/;
assign _45586_ = _45587_ & D[56] /*21404*/;
assign _45589_ = _44793_ & _45586_ /*21399*/;
assign _45590_ = _44793_ ^ _45586_ /*21402*/;
assign _45591_ = _45582_ & _45590_ /*21400*/;
assign _45241_ = _45582_ ^ _45590_ /*21401*/;
assign _45588_ = _45589_ | _45591_ /*21398*/;
assign _45593_ = ~Q[13] /*21397*/;
assign _45592_ = _45593_ & D[57] /*21396*/;
assign _45595_ = _44794_ & _45592_ /*21391*/;
assign _45596_ = _44794_ ^ _45592_ /*21394*/;
assign _45597_ = _45588_ & _45596_ /*21392*/;
assign _45242_ = _45588_ ^ _45596_ /*21393*/;
assign _45594_ = _45595_ | _45597_ /*21390*/;
assign _45599_ = ~Q[13] /*21389*/;
assign _45598_ = _45599_ & D[58] /*21388*/;
assign _45601_ = _44795_ & _45598_ /*21383*/;
assign _45602_ = _44795_ ^ _45598_ /*21386*/;
assign _45603_ = _45594_ & _45602_ /*21384*/;
assign _45243_ = _45594_ ^ _45602_ /*21385*/;
assign _45600_ = _45601_ | _45603_ /*21382*/;
assign _45605_ = ~Q[13] /*21381*/;
assign _45604_ = _45605_ & D[59] /*21380*/;
assign _45607_ = _44796_ & _45604_ /*21375*/;
assign _45608_ = _44796_ ^ _45604_ /*21378*/;
assign _45609_ = _45600_ & _45608_ /*21376*/;
assign _45244_ = _45600_ ^ _45608_ /*21377*/;
assign _45606_ = _45607_ | _45609_ /*21374*/;
assign _45611_ = ~Q[13] /*21373*/;
assign _45610_ = _45611_ & D[60] /*21372*/;
assign _45613_ = _44797_ & _45610_ /*21367*/;
assign _45614_ = _44797_ ^ _45610_ /*21370*/;
assign _45615_ = _45606_ & _45614_ /*21368*/;
assign _45245_ = _45606_ ^ _45614_ /*21369*/;
assign _45612_ = _45613_ | _45615_ /*21366*/;
assign _45617_ = ~Q[13] /*21365*/;
assign _45616_ = _45617_ & D[61] /*21364*/;
assign _45619_ = _44798_ & _45616_ /*21359*/;
assign _45620_ = _44798_ ^ _45616_ /*21362*/;
assign _45621_ = _45612_ & _45620_ /*21360*/;
assign _45246_ = _45612_ ^ _45620_ /*21361*/;
assign _45618_ = _45619_ | _45621_ /*21358*/;
assign _45623_ = ~Q[13] /*21357*/;
assign _45622_ = _45623_ & D[62] /*21356*/;
assign _45625_ = _44799_ & _45622_ /*21351*/;
assign _45626_ = _44799_ ^ _45622_ /*21354*/;
assign _45627_ = _45618_ & _45626_ /*21352*/;
assign _45247_ = _45618_ ^ _45626_ /*21353*/;
assign _45624_ = _45625_ | _45627_ /*21350*/;
assign _45629_ = ~Q[13] /*21349*/;
assign _45628_ = _45629_ & zeroWire /*21348*/;
assign _45630_ = _44800_ ^ _45628_ /*21346*/;
assign _45248_ = _45630_ ^ _45624_ /*21345*/;
assign _45701_ = ~D[0] /*21091*/;
assign _45698_ = R_0[12] & _45701_ /*21087*/;
assign _45699_ = R_0[12] ^ _45701_ /*21090*/;
assign _45700_ = oneWire & _45699_ /*21088*/;
assign _45633_ = oneWire ^ _45699_ /*21089*/;
assign _45697_ = _45698_ | _45700_ /*21086*/;
assign _45706_ = ~D[1] /*21085*/;
assign _45703_ = _45185_ & _45706_ /*21081*/;
assign _45704_ = _45185_ ^ _45706_ /*21084*/;
assign _45705_ = _45697_ & _45704_ /*21082*/;
assign _45634_ = _45697_ ^ _45704_ /*21083*/;
assign _45702_ = _45703_ | _45705_ /*21080*/;
assign _45711_ = ~D[2] /*21079*/;
assign _45708_ = _45186_ & _45711_ /*21075*/;
assign _45709_ = _45186_ ^ _45711_ /*21078*/;
assign _45710_ = _45702_ & _45709_ /*21076*/;
assign _45635_ = _45702_ ^ _45709_ /*21077*/;
assign _45707_ = _45708_ | _45710_ /*21074*/;
assign _45716_ = ~D[3] /*21073*/;
assign _45713_ = _45187_ & _45716_ /*21069*/;
assign _45714_ = _45187_ ^ _45716_ /*21072*/;
assign _45715_ = _45707_ & _45714_ /*21070*/;
assign _45636_ = _45707_ ^ _45714_ /*21071*/;
assign _45712_ = _45713_ | _45715_ /*21068*/;
assign _45721_ = ~D[4] /*21067*/;
assign _45718_ = _45188_ & _45721_ /*21063*/;
assign _45719_ = _45188_ ^ _45721_ /*21066*/;
assign _45720_ = _45712_ & _45719_ /*21064*/;
assign _45637_ = _45712_ ^ _45719_ /*21065*/;
assign _45717_ = _45718_ | _45720_ /*21062*/;
assign _45726_ = ~D[5] /*21061*/;
assign _45723_ = _45189_ & _45726_ /*21057*/;
assign _45724_ = _45189_ ^ _45726_ /*21060*/;
assign _45725_ = _45717_ & _45724_ /*21058*/;
assign _45638_ = _45717_ ^ _45724_ /*21059*/;
assign _45722_ = _45723_ | _45725_ /*21056*/;
assign _45731_ = ~D[6] /*21055*/;
assign _45728_ = _45190_ & _45731_ /*21051*/;
assign _45729_ = _45190_ ^ _45731_ /*21054*/;
assign _45730_ = _45722_ & _45729_ /*21052*/;
assign _45639_ = _45722_ ^ _45729_ /*21053*/;
assign _45727_ = _45728_ | _45730_ /*21050*/;
assign _45736_ = ~D[7] /*21049*/;
assign _45733_ = _45191_ & _45736_ /*21045*/;
assign _45734_ = _45191_ ^ _45736_ /*21048*/;
assign _45735_ = _45727_ & _45734_ /*21046*/;
assign _45640_ = _45727_ ^ _45734_ /*21047*/;
assign _45732_ = _45733_ | _45735_ /*21044*/;
assign _45741_ = ~D[8] /*21043*/;
assign _45738_ = _45192_ & _45741_ /*21039*/;
assign _45739_ = _45192_ ^ _45741_ /*21042*/;
assign _45740_ = _45732_ & _45739_ /*21040*/;
assign _45641_ = _45732_ ^ _45739_ /*21041*/;
assign _45737_ = _45738_ | _45740_ /*21038*/;
assign _45746_ = ~D[9] /*21037*/;
assign _45743_ = _45193_ & _45746_ /*21033*/;
assign _45744_ = _45193_ ^ _45746_ /*21036*/;
assign _45745_ = _45737_ & _45744_ /*21034*/;
assign _45642_ = _45737_ ^ _45744_ /*21035*/;
assign _45742_ = _45743_ | _45745_ /*21032*/;
assign _45751_ = ~D[10] /*21031*/;
assign _45748_ = _45194_ & _45751_ /*21027*/;
assign _45749_ = _45194_ ^ _45751_ /*21030*/;
assign _45750_ = _45742_ & _45749_ /*21028*/;
assign _45643_ = _45742_ ^ _45749_ /*21029*/;
assign _45747_ = _45748_ | _45750_ /*21026*/;
assign _45756_ = ~D[11] /*21025*/;
assign _45753_ = _45195_ & _45756_ /*21021*/;
assign _45754_ = _45195_ ^ _45756_ /*21024*/;
assign _45755_ = _45747_ & _45754_ /*21022*/;
assign _45644_ = _45747_ ^ _45754_ /*21023*/;
assign _45752_ = _45753_ | _45755_ /*21020*/;
assign _45761_ = ~D[12] /*21019*/;
assign _45758_ = _45196_ & _45761_ /*21015*/;
assign _45759_ = _45196_ ^ _45761_ /*21018*/;
assign _45760_ = _45752_ & _45759_ /*21016*/;
assign _45645_ = _45752_ ^ _45759_ /*21017*/;
assign _45757_ = _45758_ | _45760_ /*21014*/;
assign _45766_ = ~D[13] /*21013*/;
assign _45763_ = _45197_ & _45766_ /*21009*/;
assign _45764_ = _45197_ ^ _45766_ /*21012*/;
assign _45765_ = _45757_ & _45764_ /*21010*/;
assign _45646_ = _45757_ ^ _45764_ /*21011*/;
assign _45762_ = _45763_ | _45765_ /*21008*/;
assign _45771_ = ~D[14] /*21007*/;
assign _45768_ = _45198_ & _45771_ /*21003*/;
assign _45769_ = _45198_ ^ _45771_ /*21006*/;
assign _45770_ = _45762_ & _45769_ /*21004*/;
assign _45647_ = _45762_ ^ _45769_ /*21005*/;
assign _45767_ = _45768_ | _45770_ /*21002*/;
assign _45776_ = ~D[15] /*21001*/;
assign _45773_ = _45199_ & _45776_ /*20997*/;
assign _45774_ = _45199_ ^ _45776_ /*21000*/;
assign _45775_ = _45767_ & _45774_ /*20998*/;
assign _45648_ = _45767_ ^ _45774_ /*20999*/;
assign _45772_ = _45773_ | _45775_ /*20996*/;
assign _45781_ = ~D[16] /*20995*/;
assign _45778_ = _45200_ & _45781_ /*20991*/;
assign _45779_ = _45200_ ^ _45781_ /*20994*/;
assign _45780_ = _45772_ & _45779_ /*20992*/;
assign _45649_ = _45772_ ^ _45779_ /*20993*/;
assign _45777_ = _45778_ | _45780_ /*20990*/;
assign _45786_ = ~D[17] /*20989*/;
assign _45783_ = _45201_ & _45786_ /*20985*/;
assign _45784_ = _45201_ ^ _45786_ /*20988*/;
assign _45785_ = _45777_ & _45784_ /*20986*/;
assign _45650_ = _45777_ ^ _45784_ /*20987*/;
assign _45782_ = _45783_ | _45785_ /*20984*/;
assign _45791_ = ~D[18] /*20983*/;
assign _45788_ = _45202_ & _45791_ /*20979*/;
assign _45789_ = _45202_ ^ _45791_ /*20982*/;
assign _45790_ = _45782_ & _45789_ /*20980*/;
assign _45651_ = _45782_ ^ _45789_ /*20981*/;
assign _45787_ = _45788_ | _45790_ /*20978*/;
assign _45796_ = ~D[19] /*20977*/;
assign _45793_ = _45203_ & _45796_ /*20973*/;
assign _45794_ = _45203_ ^ _45796_ /*20976*/;
assign _45795_ = _45787_ & _45794_ /*20974*/;
assign _45652_ = _45787_ ^ _45794_ /*20975*/;
assign _45792_ = _45793_ | _45795_ /*20972*/;
assign _45801_ = ~D[20] /*20971*/;
assign _45798_ = _45204_ & _45801_ /*20967*/;
assign _45799_ = _45204_ ^ _45801_ /*20970*/;
assign _45800_ = _45792_ & _45799_ /*20968*/;
assign _45653_ = _45792_ ^ _45799_ /*20969*/;
assign _45797_ = _45798_ | _45800_ /*20966*/;
assign _45806_ = ~D[21] /*20965*/;
assign _45803_ = _45205_ & _45806_ /*20961*/;
assign _45804_ = _45205_ ^ _45806_ /*20964*/;
assign _45805_ = _45797_ & _45804_ /*20962*/;
assign _45654_ = _45797_ ^ _45804_ /*20963*/;
assign _45802_ = _45803_ | _45805_ /*20960*/;
assign _45811_ = ~D[22] /*20959*/;
assign _45808_ = _45206_ & _45811_ /*20955*/;
assign _45809_ = _45206_ ^ _45811_ /*20958*/;
assign _45810_ = _45802_ & _45809_ /*20956*/;
assign _45655_ = _45802_ ^ _45809_ /*20957*/;
assign _45807_ = _45808_ | _45810_ /*20954*/;
assign _45816_ = ~D[23] /*20953*/;
assign _45813_ = _45207_ & _45816_ /*20949*/;
assign _45814_ = _45207_ ^ _45816_ /*20952*/;
assign _45815_ = _45807_ & _45814_ /*20950*/;
assign _45656_ = _45807_ ^ _45814_ /*20951*/;
assign _45812_ = _45813_ | _45815_ /*20948*/;
assign _45821_ = ~D[24] /*20947*/;
assign _45818_ = _45208_ & _45821_ /*20943*/;
assign _45819_ = _45208_ ^ _45821_ /*20946*/;
assign _45820_ = _45812_ & _45819_ /*20944*/;
assign _45657_ = _45812_ ^ _45819_ /*20945*/;
assign _45817_ = _45818_ | _45820_ /*20942*/;
assign _45826_ = ~D[25] /*20941*/;
assign _45823_ = _45209_ & _45826_ /*20937*/;
assign _45824_ = _45209_ ^ _45826_ /*20940*/;
assign _45825_ = _45817_ & _45824_ /*20938*/;
assign _45658_ = _45817_ ^ _45824_ /*20939*/;
assign _45822_ = _45823_ | _45825_ /*20936*/;
assign _45831_ = ~D[26] /*20935*/;
assign _45828_ = _45210_ & _45831_ /*20931*/;
assign _45829_ = _45210_ ^ _45831_ /*20934*/;
assign _45830_ = _45822_ & _45829_ /*20932*/;
assign _45659_ = _45822_ ^ _45829_ /*20933*/;
assign _45827_ = _45828_ | _45830_ /*20930*/;
assign _45836_ = ~D[27] /*20929*/;
assign _45833_ = _45211_ & _45836_ /*20925*/;
assign _45834_ = _45211_ ^ _45836_ /*20928*/;
assign _45835_ = _45827_ & _45834_ /*20926*/;
assign _45660_ = _45827_ ^ _45834_ /*20927*/;
assign _45832_ = _45833_ | _45835_ /*20924*/;
assign _45841_ = ~D[28] /*20923*/;
assign _45838_ = _45212_ & _45841_ /*20919*/;
assign _45839_ = _45212_ ^ _45841_ /*20922*/;
assign _45840_ = _45832_ & _45839_ /*20920*/;
assign _45661_ = _45832_ ^ _45839_ /*20921*/;
assign _45837_ = _45838_ | _45840_ /*20918*/;
assign _45846_ = ~D[29] /*20917*/;
assign _45843_ = _45213_ & _45846_ /*20913*/;
assign _45844_ = _45213_ ^ _45846_ /*20916*/;
assign _45845_ = _45837_ & _45844_ /*20914*/;
assign _45662_ = _45837_ ^ _45844_ /*20915*/;
assign _45842_ = _45843_ | _45845_ /*20912*/;
assign _45851_ = ~D[30] /*20911*/;
assign _45848_ = _45214_ & _45851_ /*20907*/;
assign _45849_ = _45214_ ^ _45851_ /*20910*/;
assign _45850_ = _45842_ & _45849_ /*20908*/;
assign _45663_ = _45842_ ^ _45849_ /*20909*/;
assign _45847_ = _45848_ | _45850_ /*20906*/;
assign _45856_ = ~D[31] /*20905*/;
assign _45853_ = _45215_ & _45856_ /*20901*/;
assign _45854_ = _45215_ ^ _45856_ /*20904*/;
assign _45855_ = _45847_ & _45854_ /*20902*/;
assign _45664_ = _45847_ ^ _45854_ /*20903*/;
assign _45852_ = _45853_ | _45855_ /*20900*/;
assign _45861_ = ~D[32] /*20899*/;
assign _45858_ = _45216_ & _45861_ /*20895*/;
assign _45859_ = _45216_ ^ _45861_ /*20898*/;
assign _45860_ = _45852_ & _45859_ /*20896*/;
assign _45665_ = _45852_ ^ _45859_ /*20897*/;
assign _45857_ = _45858_ | _45860_ /*20894*/;
assign _45866_ = ~D[33] /*20893*/;
assign _45863_ = _45217_ & _45866_ /*20889*/;
assign _45864_ = _45217_ ^ _45866_ /*20892*/;
assign _45865_ = _45857_ & _45864_ /*20890*/;
assign _45666_ = _45857_ ^ _45864_ /*20891*/;
assign _45862_ = _45863_ | _45865_ /*20888*/;
assign _45871_ = ~D[34] /*20887*/;
assign _45868_ = _45218_ & _45871_ /*20883*/;
assign _45869_ = _45218_ ^ _45871_ /*20886*/;
assign _45870_ = _45862_ & _45869_ /*20884*/;
assign _45667_ = _45862_ ^ _45869_ /*20885*/;
assign _45867_ = _45868_ | _45870_ /*20882*/;
assign _45876_ = ~D[35] /*20881*/;
assign _45873_ = _45219_ & _45876_ /*20877*/;
assign _45874_ = _45219_ ^ _45876_ /*20880*/;
assign _45875_ = _45867_ & _45874_ /*20878*/;
assign _45668_ = _45867_ ^ _45874_ /*20879*/;
assign _45872_ = _45873_ | _45875_ /*20876*/;
assign _45881_ = ~D[36] /*20875*/;
assign _45878_ = _45220_ & _45881_ /*20871*/;
assign _45879_ = _45220_ ^ _45881_ /*20874*/;
assign _45880_ = _45872_ & _45879_ /*20872*/;
assign _45669_ = _45872_ ^ _45879_ /*20873*/;
assign _45877_ = _45878_ | _45880_ /*20870*/;
assign _45886_ = ~D[37] /*20869*/;
assign _45883_ = _45221_ & _45886_ /*20865*/;
assign _45884_ = _45221_ ^ _45886_ /*20868*/;
assign _45885_ = _45877_ & _45884_ /*20866*/;
assign _45670_ = _45877_ ^ _45884_ /*20867*/;
assign _45882_ = _45883_ | _45885_ /*20864*/;
assign _45891_ = ~D[38] /*20863*/;
assign _45888_ = _45222_ & _45891_ /*20859*/;
assign _45889_ = _45222_ ^ _45891_ /*20862*/;
assign _45890_ = _45882_ & _45889_ /*20860*/;
assign _45671_ = _45882_ ^ _45889_ /*20861*/;
assign _45887_ = _45888_ | _45890_ /*20858*/;
assign _45896_ = ~D[39] /*20857*/;
assign _45893_ = _45223_ & _45896_ /*20853*/;
assign _45894_ = _45223_ ^ _45896_ /*20856*/;
assign _45895_ = _45887_ & _45894_ /*20854*/;
assign _45672_ = _45887_ ^ _45894_ /*20855*/;
assign _45892_ = _45893_ | _45895_ /*20852*/;
assign _45901_ = ~D[40] /*20851*/;
assign _45898_ = _45224_ & _45901_ /*20847*/;
assign _45899_ = _45224_ ^ _45901_ /*20850*/;
assign _45900_ = _45892_ & _45899_ /*20848*/;
assign _45673_ = _45892_ ^ _45899_ /*20849*/;
assign _45897_ = _45898_ | _45900_ /*20846*/;
assign _45906_ = ~D[41] /*20845*/;
assign _45903_ = _45225_ & _45906_ /*20841*/;
assign _45904_ = _45225_ ^ _45906_ /*20844*/;
assign _45905_ = _45897_ & _45904_ /*20842*/;
assign _45674_ = _45897_ ^ _45904_ /*20843*/;
assign _45902_ = _45903_ | _45905_ /*20840*/;
assign _45911_ = ~D[42] /*20839*/;
assign _45908_ = _45226_ & _45911_ /*20835*/;
assign _45909_ = _45226_ ^ _45911_ /*20838*/;
assign _45910_ = _45902_ & _45909_ /*20836*/;
assign _45675_ = _45902_ ^ _45909_ /*20837*/;
assign _45907_ = _45908_ | _45910_ /*20834*/;
assign _45916_ = ~D[43] /*20833*/;
assign _45913_ = _45227_ & _45916_ /*20829*/;
assign _45914_ = _45227_ ^ _45916_ /*20832*/;
assign _45915_ = _45907_ & _45914_ /*20830*/;
assign _45676_ = _45907_ ^ _45914_ /*20831*/;
assign _45912_ = _45913_ | _45915_ /*20828*/;
assign _45921_ = ~D[44] /*20827*/;
assign _45918_ = _45228_ & _45921_ /*20823*/;
assign _45919_ = _45228_ ^ _45921_ /*20826*/;
assign _45920_ = _45912_ & _45919_ /*20824*/;
assign _45677_ = _45912_ ^ _45919_ /*20825*/;
assign _45917_ = _45918_ | _45920_ /*20822*/;
assign _45926_ = ~D[45] /*20821*/;
assign _45923_ = _45229_ & _45926_ /*20817*/;
assign _45924_ = _45229_ ^ _45926_ /*20820*/;
assign _45925_ = _45917_ & _45924_ /*20818*/;
assign _45678_ = _45917_ ^ _45924_ /*20819*/;
assign _45922_ = _45923_ | _45925_ /*20816*/;
assign _45931_ = ~D[46] /*20815*/;
assign _45928_ = _45230_ & _45931_ /*20811*/;
assign _45929_ = _45230_ ^ _45931_ /*20814*/;
assign _45930_ = _45922_ & _45929_ /*20812*/;
assign _45679_ = _45922_ ^ _45929_ /*20813*/;
assign _45927_ = _45928_ | _45930_ /*20810*/;
assign _45936_ = ~D[47] /*20809*/;
assign _45933_ = _45231_ & _45936_ /*20805*/;
assign _45934_ = _45231_ ^ _45936_ /*20808*/;
assign _45935_ = _45927_ & _45934_ /*20806*/;
assign _45680_ = _45927_ ^ _45934_ /*20807*/;
assign _45932_ = _45933_ | _45935_ /*20804*/;
assign _45941_ = ~D[48] /*20803*/;
assign _45938_ = _45232_ & _45941_ /*20799*/;
assign _45939_ = _45232_ ^ _45941_ /*20802*/;
assign _45940_ = _45932_ & _45939_ /*20800*/;
assign _45681_ = _45932_ ^ _45939_ /*20801*/;
assign _45937_ = _45938_ | _45940_ /*20798*/;
assign _45946_ = ~D[49] /*20797*/;
assign _45943_ = _45233_ & _45946_ /*20793*/;
assign _45944_ = _45233_ ^ _45946_ /*20796*/;
assign _45945_ = _45937_ & _45944_ /*20794*/;
assign _45682_ = _45937_ ^ _45944_ /*20795*/;
assign _45942_ = _45943_ | _45945_ /*20792*/;
assign _45951_ = ~D[50] /*20791*/;
assign _45948_ = _45234_ & _45951_ /*20787*/;
assign _45949_ = _45234_ ^ _45951_ /*20790*/;
assign _45950_ = _45942_ & _45949_ /*20788*/;
assign _45683_ = _45942_ ^ _45949_ /*20789*/;
assign _45947_ = _45948_ | _45950_ /*20786*/;
assign _45956_ = ~D[51] /*20785*/;
assign _45953_ = _45235_ & _45956_ /*20781*/;
assign _45954_ = _45235_ ^ _45956_ /*20784*/;
assign _45955_ = _45947_ & _45954_ /*20782*/;
assign _45684_ = _45947_ ^ _45954_ /*20783*/;
assign _45952_ = _45953_ | _45955_ /*20780*/;
assign _45961_ = ~D[52] /*20779*/;
assign _45958_ = _45236_ & _45961_ /*20775*/;
assign _45959_ = _45236_ ^ _45961_ /*20778*/;
assign _45960_ = _45952_ & _45959_ /*20776*/;
assign _45685_ = _45952_ ^ _45959_ /*20777*/;
assign _45957_ = _45958_ | _45960_ /*20774*/;
assign _45966_ = ~D[53] /*20773*/;
assign _45963_ = _45237_ & _45966_ /*20769*/;
assign _45964_ = _45237_ ^ _45966_ /*20772*/;
assign _45965_ = _45957_ & _45964_ /*20770*/;
assign _45686_ = _45957_ ^ _45964_ /*20771*/;
assign _45962_ = _45963_ | _45965_ /*20768*/;
assign _45971_ = ~D[54] /*20767*/;
assign _45968_ = _45238_ & _45971_ /*20763*/;
assign _45969_ = _45238_ ^ _45971_ /*20766*/;
assign _45970_ = _45962_ & _45969_ /*20764*/;
assign _45687_ = _45962_ ^ _45969_ /*20765*/;
assign _45967_ = _45968_ | _45970_ /*20762*/;
assign _45976_ = ~D[55] /*20761*/;
assign _45973_ = _45239_ & _45976_ /*20757*/;
assign _45974_ = _45239_ ^ _45976_ /*20760*/;
assign _45975_ = _45967_ & _45974_ /*20758*/;
assign _45688_ = _45967_ ^ _45974_ /*20759*/;
assign _45972_ = _45973_ | _45975_ /*20756*/;
assign _45981_ = ~D[56] /*20755*/;
assign _45978_ = _45240_ & _45981_ /*20751*/;
assign _45979_ = _45240_ ^ _45981_ /*20754*/;
assign _45980_ = _45972_ & _45979_ /*20752*/;
assign _45689_ = _45972_ ^ _45979_ /*20753*/;
assign _45977_ = _45978_ | _45980_ /*20750*/;
assign _45986_ = ~D[57] /*20749*/;
assign _45983_ = _45241_ & _45986_ /*20745*/;
assign _45984_ = _45241_ ^ _45986_ /*20748*/;
assign _45985_ = _45977_ & _45984_ /*20746*/;
assign _45690_ = _45977_ ^ _45984_ /*20747*/;
assign _45982_ = _45983_ | _45985_ /*20744*/;
assign _45991_ = ~D[58] /*20743*/;
assign _45988_ = _45242_ & _45991_ /*20739*/;
assign _45989_ = _45242_ ^ _45991_ /*20742*/;
assign _45990_ = _45982_ & _45989_ /*20740*/;
assign _45691_ = _45982_ ^ _45989_ /*20741*/;
assign _45987_ = _45988_ | _45990_ /*20738*/;
assign _45996_ = ~D[59] /*20737*/;
assign _45993_ = _45243_ & _45996_ /*20733*/;
assign _45994_ = _45243_ ^ _45996_ /*20736*/;
assign _45995_ = _45987_ & _45994_ /*20734*/;
assign _45692_ = _45987_ ^ _45994_ /*20735*/;
assign _45992_ = _45993_ | _45995_ /*20732*/;
assign _46001_ = ~D[60] /*20731*/;
assign _45998_ = _45244_ & _46001_ /*20727*/;
assign _45999_ = _45244_ ^ _46001_ /*20730*/;
assign _46000_ = _45992_ & _45999_ /*20728*/;
assign _45693_ = _45992_ ^ _45999_ /*20729*/;
assign _45997_ = _45998_ | _46000_ /*20726*/;
assign _46006_ = ~D[61] /*20725*/;
assign _46003_ = _45245_ & _46006_ /*20721*/;
assign _46004_ = _45245_ ^ _46006_ /*20724*/;
assign _46005_ = _45997_ & _46004_ /*20722*/;
assign _45694_ = _45997_ ^ _46004_ /*20723*/;
assign _46002_ = _46003_ | _46005_ /*20720*/;
assign _46011_ = ~D[62] /*20719*/;
assign _46008_ = _45246_ & _46011_ /*20715*/;
assign _46009_ = _45246_ ^ _46011_ /*20718*/;
assign _46010_ = _46002_ & _46009_ /*20716*/;
assign _45695_ = _46002_ ^ _46009_ /*20717*/;
assign _46007_ = _46008_ | _46010_ /*20714*/;
assign _46012_ = _45247_ & oneWire /*20709*/;
assign _46013_ = _45247_ ^ oneWire /*20712*/;
assign _46014_ = _46007_ & _46013_ /*20710*/;
assign _45696_ = _46007_ ^ _46013_ /*20711*/;
assign Q[12] = _46012_ | _46014_ /*20708*/;
assign _46147_ = ~Q[12] /*20323*/;
assign _46146_ = _46147_ & D[0] /*20322*/;
assign _46149_ = _45633_ & _46146_ /*20317*/;
assign _46150_ = _45633_ ^ _46146_ /*20320*/;
assign _46151_ = zeroWire & _46150_ /*20318*/;
assign _46081_ = zeroWire ^ _46150_ /*20319*/;
assign _46148_ = _46149_ | _46151_ /*20316*/;
assign _46153_ = ~Q[12] /*20315*/;
assign _46152_ = _46153_ & D[1] /*20314*/;
assign _46155_ = _45634_ & _46152_ /*20309*/;
assign _46156_ = _45634_ ^ _46152_ /*20312*/;
assign _46157_ = _46148_ & _46156_ /*20310*/;
assign _46082_ = _46148_ ^ _46156_ /*20311*/;
assign _46154_ = _46155_ | _46157_ /*20308*/;
assign _46159_ = ~Q[12] /*20307*/;
assign _46158_ = _46159_ & D[2] /*20306*/;
assign _46161_ = _45635_ & _46158_ /*20301*/;
assign _46162_ = _45635_ ^ _46158_ /*20304*/;
assign _46163_ = _46154_ & _46162_ /*20302*/;
assign _46083_ = _46154_ ^ _46162_ /*20303*/;
assign _46160_ = _46161_ | _46163_ /*20300*/;
assign _46165_ = ~Q[12] /*20299*/;
assign _46164_ = _46165_ & D[3] /*20298*/;
assign _46167_ = _45636_ & _46164_ /*20293*/;
assign _46168_ = _45636_ ^ _46164_ /*20296*/;
assign _46169_ = _46160_ & _46168_ /*20294*/;
assign _46084_ = _46160_ ^ _46168_ /*20295*/;
assign _46166_ = _46167_ | _46169_ /*20292*/;
assign _46171_ = ~Q[12] /*20291*/;
assign _46170_ = _46171_ & D[4] /*20290*/;
assign _46173_ = _45637_ & _46170_ /*20285*/;
assign _46174_ = _45637_ ^ _46170_ /*20288*/;
assign _46175_ = _46166_ & _46174_ /*20286*/;
assign _46085_ = _46166_ ^ _46174_ /*20287*/;
assign _46172_ = _46173_ | _46175_ /*20284*/;
assign _46177_ = ~Q[12] /*20283*/;
assign _46176_ = _46177_ & D[5] /*20282*/;
assign _46179_ = _45638_ & _46176_ /*20277*/;
assign _46180_ = _45638_ ^ _46176_ /*20280*/;
assign _46181_ = _46172_ & _46180_ /*20278*/;
assign _46086_ = _46172_ ^ _46180_ /*20279*/;
assign _46178_ = _46179_ | _46181_ /*20276*/;
assign _46183_ = ~Q[12] /*20275*/;
assign _46182_ = _46183_ & D[6] /*20274*/;
assign _46185_ = _45639_ & _46182_ /*20269*/;
assign _46186_ = _45639_ ^ _46182_ /*20272*/;
assign _46187_ = _46178_ & _46186_ /*20270*/;
assign _46087_ = _46178_ ^ _46186_ /*20271*/;
assign _46184_ = _46185_ | _46187_ /*20268*/;
assign _46189_ = ~Q[12] /*20267*/;
assign _46188_ = _46189_ & D[7] /*20266*/;
assign _46191_ = _45640_ & _46188_ /*20261*/;
assign _46192_ = _45640_ ^ _46188_ /*20264*/;
assign _46193_ = _46184_ & _46192_ /*20262*/;
assign _46088_ = _46184_ ^ _46192_ /*20263*/;
assign _46190_ = _46191_ | _46193_ /*20260*/;
assign _46195_ = ~Q[12] /*20259*/;
assign _46194_ = _46195_ & D[8] /*20258*/;
assign _46197_ = _45641_ & _46194_ /*20253*/;
assign _46198_ = _45641_ ^ _46194_ /*20256*/;
assign _46199_ = _46190_ & _46198_ /*20254*/;
assign _46089_ = _46190_ ^ _46198_ /*20255*/;
assign _46196_ = _46197_ | _46199_ /*20252*/;
assign _46201_ = ~Q[12] /*20251*/;
assign _46200_ = _46201_ & D[9] /*20250*/;
assign _46203_ = _45642_ & _46200_ /*20245*/;
assign _46204_ = _45642_ ^ _46200_ /*20248*/;
assign _46205_ = _46196_ & _46204_ /*20246*/;
assign _46090_ = _46196_ ^ _46204_ /*20247*/;
assign _46202_ = _46203_ | _46205_ /*20244*/;
assign _46207_ = ~Q[12] /*20243*/;
assign _46206_ = _46207_ & D[10] /*20242*/;
assign _46209_ = _45643_ & _46206_ /*20237*/;
assign _46210_ = _45643_ ^ _46206_ /*20240*/;
assign _46211_ = _46202_ & _46210_ /*20238*/;
assign _46091_ = _46202_ ^ _46210_ /*20239*/;
assign _46208_ = _46209_ | _46211_ /*20236*/;
assign _46213_ = ~Q[12] /*20235*/;
assign _46212_ = _46213_ & D[11] /*20234*/;
assign _46215_ = _45644_ & _46212_ /*20229*/;
assign _46216_ = _45644_ ^ _46212_ /*20232*/;
assign _46217_ = _46208_ & _46216_ /*20230*/;
assign _46092_ = _46208_ ^ _46216_ /*20231*/;
assign _46214_ = _46215_ | _46217_ /*20228*/;
assign _46219_ = ~Q[12] /*20227*/;
assign _46218_ = _46219_ & D[12] /*20226*/;
assign _46221_ = _45645_ & _46218_ /*20221*/;
assign _46222_ = _45645_ ^ _46218_ /*20224*/;
assign _46223_ = _46214_ & _46222_ /*20222*/;
assign _46093_ = _46214_ ^ _46222_ /*20223*/;
assign _46220_ = _46221_ | _46223_ /*20220*/;
assign _46225_ = ~Q[12] /*20219*/;
assign _46224_ = _46225_ & D[13] /*20218*/;
assign _46227_ = _45646_ & _46224_ /*20213*/;
assign _46228_ = _45646_ ^ _46224_ /*20216*/;
assign _46229_ = _46220_ & _46228_ /*20214*/;
assign _46094_ = _46220_ ^ _46228_ /*20215*/;
assign _46226_ = _46227_ | _46229_ /*20212*/;
assign _46231_ = ~Q[12] /*20211*/;
assign _46230_ = _46231_ & D[14] /*20210*/;
assign _46233_ = _45647_ & _46230_ /*20205*/;
assign _46234_ = _45647_ ^ _46230_ /*20208*/;
assign _46235_ = _46226_ & _46234_ /*20206*/;
assign _46095_ = _46226_ ^ _46234_ /*20207*/;
assign _46232_ = _46233_ | _46235_ /*20204*/;
assign _46237_ = ~Q[12] /*20203*/;
assign _46236_ = _46237_ & D[15] /*20202*/;
assign _46239_ = _45648_ & _46236_ /*20197*/;
assign _46240_ = _45648_ ^ _46236_ /*20200*/;
assign _46241_ = _46232_ & _46240_ /*20198*/;
assign _46096_ = _46232_ ^ _46240_ /*20199*/;
assign _46238_ = _46239_ | _46241_ /*20196*/;
assign _46243_ = ~Q[12] /*20195*/;
assign _46242_ = _46243_ & D[16] /*20194*/;
assign _46245_ = _45649_ & _46242_ /*20189*/;
assign _46246_ = _45649_ ^ _46242_ /*20192*/;
assign _46247_ = _46238_ & _46246_ /*20190*/;
assign _46097_ = _46238_ ^ _46246_ /*20191*/;
assign _46244_ = _46245_ | _46247_ /*20188*/;
assign _46249_ = ~Q[12] /*20187*/;
assign _46248_ = _46249_ & D[17] /*20186*/;
assign _46251_ = _45650_ & _46248_ /*20181*/;
assign _46252_ = _45650_ ^ _46248_ /*20184*/;
assign _46253_ = _46244_ & _46252_ /*20182*/;
assign _46098_ = _46244_ ^ _46252_ /*20183*/;
assign _46250_ = _46251_ | _46253_ /*20180*/;
assign _46255_ = ~Q[12] /*20179*/;
assign _46254_ = _46255_ & D[18] /*20178*/;
assign _46257_ = _45651_ & _46254_ /*20173*/;
assign _46258_ = _45651_ ^ _46254_ /*20176*/;
assign _46259_ = _46250_ & _46258_ /*20174*/;
assign _46099_ = _46250_ ^ _46258_ /*20175*/;
assign _46256_ = _46257_ | _46259_ /*20172*/;
assign _46261_ = ~Q[12] /*20171*/;
assign _46260_ = _46261_ & D[19] /*20170*/;
assign _46263_ = _45652_ & _46260_ /*20165*/;
assign _46264_ = _45652_ ^ _46260_ /*20168*/;
assign _46265_ = _46256_ & _46264_ /*20166*/;
assign _46100_ = _46256_ ^ _46264_ /*20167*/;
assign _46262_ = _46263_ | _46265_ /*20164*/;
assign _46267_ = ~Q[12] /*20163*/;
assign _46266_ = _46267_ & D[20] /*20162*/;
assign _46269_ = _45653_ & _46266_ /*20157*/;
assign _46270_ = _45653_ ^ _46266_ /*20160*/;
assign _46271_ = _46262_ & _46270_ /*20158*/;
assign _46101_ = _46262_ ^ _46270_ /*20159*/;
assign _46268_ = _46269_ | _46271_ /*20156*/;
assign _46273_ = ~Q[12] /*20155*/;
assign _46272_ = _46273_ & D[21] /*20154*/;
assign _46275_ = _45654_ & _46272_ /*20149*/;
assign _46276_ = _45654_ ^ _46272_ /*20152*/;
assign _46277_ = _46268_ & _46276_ /*20150*/;
assign _46102_ = _46268_ ^ _46276_ /*20151*/;
assign _46274_ = _46275_ | _46277_ /*20148*/;
assign _46279_ = ~Q[12] /*20147*/;
assign _46278_ = _46279_ & D[22] /*20146*/;
assign _46281_ = _45655_ & _46278_ /*20141*/;
assign _46282_ = _45655_ ^ _46278_ /*20144*/;
assign _46283_ = _46274_ & _46282_ /*20142*/;
assign _46103_ = _46274_ ^ _46282_ /*20143*/;
assign _46280_ = _46281_ | _46283_ /*20140*/;
assign _46285_ = ~Q[12] /*20139*/;
assign _46284_ = _46285_ & D[23] /*20138*/;
assign _46287_ = _45656_ & _46284_ /*20133*/;
assign _46288_ = _45656_ ^ _46284_ /*20136*/;
assign _46289_ = _46280_ & _46288_ /*20134*/;
assign _46104_ = _46280_ ^ _46288_ /*20135*/;
assign _46286_ = _46287_ | _46289_ /*20132*/;
assign _46291_ = ~Q[12] /*20131*/;
assign _46290_ = _46291_ & D[24] /*20130*/;
assign _46293_ = _45657_ & _46290_ /*20125*/;
assign _46294_ = _45657_ ^ _46290_ /*20128*/;
assign _46295_ = _46286_ & _46294_ /*20126*/;
assign _46105_ = _46286_ ^ _46294_ /*20127*/;
assign _46292_ = _46293_ | _46295_ /*20124*/;
assign _46297_ = ~Q[12] /*20123*/;
assign _46296_ = _46297_ & D[25] /*20122*/;
assign _46299_ = _45658_ & _46296_ /*20117*/;
assign _46300_ = _45658_ ^ _46296_ /*20120*/;
assign _46301_ = _46292_ & _46300_ /*20118*/;
assign _46106_ = _46292_ ^ _46300_ /*20119*/;
assign _46298_ = _46299_ | _46301_ /*20116*/;
assign _46303_ = ~Q[12] /*20115*/;
assign _46302_ = _46303_ & D[26] /*20114*/;
assign _46305_ = _45659_ & _46302_ /*20109*/;
assign _46306_ = _45659_ ^ _46302_ /*20112*/;
assign _46307_ = _46298_ & _46306_ /*20110*/;
assign _46107_ = _46298_ ^ _46306_ /*20111*/;
assign _46304_ = _46305_ | _46307_ /*20108*/;
assign _46309_ = ~Q[12] /*20107*/;
assign _46308_ = _46309_ & D[27] /*20106*/;
assign _46311_ = _45660_ & _46308_ /*20101*/;
assign _46312_ = _45660_ ^ _46308_ /*20104*/;
assign _46313_ = _46304_ & _46312_ /*20102*/;
assign _46108_ = _46304_ ^ _46312_ /*20103*/;
assign _46310_ = _46311_ | _46313_ /*20100*/;
assign _46315_ = ~Q[12] /*20099*/;
assign _46314_ = _46315_ & D[28] /*20098*/;
assign _46317_ = _45661_ & _46314_ /*20093*/;
assign _46318_ = _45661_ ^ _46314_ /*20096*/;
assign _46319_ = _46310_ & _46318_ /*20094*/;
assign _46109_ = _46310_ ^ _46318_ /*20095*/;
assign _46316_ = _46317_ | _46319_ /*20092*/;
assign _46321_ = ~Q[12] /*20091*/;
assign _46320_ = _46321_ & D[29] /*20090*/;
assign _46323_ = _45662_ & _46320_ /*20085*/;
assign _46324_ = _45662_ ^ _46320_ /*20088*/;
assign _46325_ = _46316_ & _46324_ /*20086*/;
assign _46110_ = _46316_ ^ _46324_ /*20087*/;
assign _46322_ = _46323_ | _46325_ /*20084*/;
assign _46327_ = ~Q[12] /*20083*/;
assign _46326_ = _46327_ & D[30] /*20082*/;
assign _46329_ = _45663_ & _46326_ /*20077*/;
assign _46330_ = _45663_ ^ _46326_ /*20080*/;
assign _46331_ = _46322_ & _46330_ /*20078*/;
assign _46111_ = _46322_ ^ _46330_ /*20079*/;
assign _46328_ = _46329_ | _46331_ /*20076*/;
assign _46333_ = ~Q[12] /*20075*/;
assign _46332_ = _46333_ & D[31] /*20074*/;
assign _46335_ = _45664_ & _46332_ /*20069*/;
assign _46336_ = _45664_ ^ _46332_ /*20072*/;
assign _46337_ = _46328_ & _46336_ /*20070*/;
assign _46112_ = _46328_ ^ _46336_ /*20071*/;
assign _46334_ = _46335_ | _46337_ /*20068*/;
assign _46339_ = ~Q[12] /*20067*/;
assign _46338_ = _46339_ & D[32] /*20066*/;
assign _46341_ = _45665_ & _46338_ /*20061*/;
assign _46342_ = _45665_ ^ _46338_ /*20064*/;
assign _46343_ = _46334_ & _46342_ /*20062*/;
assign _46113_ = _46334_ ^ _46342_ /*20063*/;
assign _46340_ = _46341_ | _46343_ /*20060*/;
assign _46345_ = ~Q[12] /*20059*/;
assign _46344_ = _46345_ & D[33] /*20058*/;
assign _46347_ = _45666_ & _46344_ /*20053*/;
assign _46348_ = _45666_ ^ _46344_ /*20056*/;
assign _46349_ = _46340_ & _46348_ /*20054*/;
assign _46114_ = _46340_ ^ _46348_ /*20055*/;
assign _46346_ = _46347_ | _46349_ /*20052*/;
assign _46351_ = ~Q[12] /*20051*/;
assign _46350_ = _46351_ & D[34] /*20050*/;
assign _46353_ = _45667_ & _46350_ /*20045*/;
assign _46354_ = _45667_ ^ _46350_ /*20048*/;
assign _46355_ = _46346_ & _46354_ /*20046*/;
assign _46115_ = _46346_ ^ _46354_ /*20047*/;
assign _46352_ = _46353_ | _46355_ /*20044*/;
assign _46357_ = ~Q[12] /*20043*/;
assign _46356_ = _46357_ & D[35] /*20042*/;
assign _46359_ = _45668_ & _46356_ /*20037*/;
assign _46360_ = _45668_ ^ _46356_ /*20040*/;
assign _46361_ = _46352_ & _46360_ /*20038*/;
assign _46116_ = _46352_ ^ _46360_ /*20039*/;
assign _46358_ = _46359_ | _46361_ /*20036*/;
assign _46363_ = ~Q[12] /*20035*/;
assign _46362_ = _46363_ & D[36] /*20034*/;
assign _46365_ = _45669_ & _46362_ /*20029*/;
assign _46366_ = _45669_ ^ _46362_ /*20032*/;
assign _46367_ = _46358_ & _46366_ /*20030*/;
assign _46117_ = _46358_ ^ _46366_ /*20031*/;
assign _46364_ = _46365_ | _46367_ /*20028*/;
assign _46369_ = ~Q[12] /*20027*/;
assign _46368_ = _46369_ & D[37] /*20026*/;
assign _46371_ = _45670_ & _46368_ /*20021*/;
assign _46372_ = _45670_ ^ _46368_ /*20024*/;
assign _46373_ = _46364_ & _46372_ /*20022*/;
assign _46118_ = _46364_ ^ _46372_ /*20023*/;
assign _46370_ = _46371_ | _46373_ /*20020*/;
assign _46375_ = ~Q[12] /*20019*/;
assign _46374_ = _46375_ & D[38] /*20018*/;
assign _46377_ = _45671_ & _46374_ /*20013*/;
assign _46378_ = _45671_ ^ _46374_ /*20016*/;
assign _46379_ = _46370_ & _46378_ /*20014*/;
assign _46119_ = _46370_ ^ _46378_ /*20015*/;
assign _46376_ = _46377_ | _46379_ /*20012*/;
assign _46381_ = ~Q[12] /*20011*/;
assign _46380_ = _46381_ & D[39] /*20010*/;
assign _46383_ = _45672_ & _46380_ /*20005*/;
assign _46384_ = _45672_ ^ _46380_ /*20008*/;
assign _46385_ = _46376_ & _46384_ /*20006*/;
assign _46120_ = _46376_ ^ _46384_ /*20007*/;
assign _46382_ = _46383_ | _46385_ /*20004*/;
assign _46387_ = ~Q[12] /*20003*/;
assign _46386_ = _46387_ & D[40] /*20002*/;
assign _46389_ = _45673_ & _46386_ /*19997*/;
assign _46390_ = _45673_ ^ _46386_ /*20000*/;
assign _46391_ = _46382_ & _46390_ /*19998*/;
assign _46121_ = _46382_ ^ _46390_ /*19999*/;
assign _46388_ = _46389_ | _46391_ /*19996*/;
assign _46393_ = ~Q[12] /*19995*/;
assign _46392_ = _46393_ & D[41] /*19994*/;
assign _46395_ = _45674_ & _46392_ /*19989*/;
assign _46396_ = _45674_ ^ _46392_ /*19992*/;
assign _46397_ = _46388_ & _46396_ /*19990*/;
assign _46122_ = _46388_ ^ _46396_ /*19991*/;
assign _46394_ = _46395_ | _46397_ /*19988*/;
assign _46399_ = ~Q[12] /*19987*/;
assign _46398_ = _46399_ & D[42] /*19986*/;
assign _46401_ = _45675_ & _46398_ /*19981*/;
assign _46402_ = _45675_ ^ _46398_ /*19984*/;
assign _46403_ = _46394_ & _46402_ /*19982*/;
assign _46123_ = _46394_ ^ _46402_ /*19983*/;
assign _46400_ = _46401_ | _46403_ /*19980*/;
assign _46405_ = ~Q[12] /*19979*/;
assign _46404_ = _46405_ & D[43] /*19978*/;
assign _46407_ = _45676_ & _46404_ /*19973*/;
assign _46408_ = _45676_ ^ _46404_ /*19976*/;
assign _46409_ = _46400_ & _46408_ /*19974*/;
assign _46124_ = _46400_ ^ _46408_ /*19975*/;
assign _46406_ = _46407_ | _46409_ /*19972*/;
assign _46411_ = ~Q[12] /*19971*/;
assign _46410_ = _46411_ & D[44] /*19970*/;
assign _46413_ = _45677_ & _46410_ /*19965*/;
assign _46414_ = _45677_ ^ _46410_ /*19968*/;
assign _46415_ = _46406_ & _46414_ /*19966*/;
assign _46125_ = _46406_ ^ _46414_ /*19967*/;
assign _46412_ = _46413_ | _46415_ /*19964*/;
assign _46417_ = ~Q[12] /*19963*/;
assign _46416_ = _46417_ & D[45] /*19962*/;
assign _46419_ = _45678_ & _46416_ /*19957*/;
assign _46420_ = _45678_ ^ _46416_ /*19960*/;
assign _46421_ = _46412_ & _46420_ /*19958*/;
assign _46126_ = _46412_ ^ _46420_ /*19959*/;
assign _46418_ = _46419_ | _46421_ /*19956*/;
assign _46423_ = ~Q[12] /*19955*/;
assign _46422_ = _46423_ & D[46] /*19954*/;
assign _46425_ = _45679_ & _46422_ /*19949*/;
assign _46426_ = _45679_ ^ _46422_ /*19952*/;
assign _46427_ = _46418_ & _46426_ /*19950*/;
assign _46127_ = _46418_ ^ _46426_ /*19951*/;
assign _46424_ = _46425_ | _46427_ /*19948*/;
assign _46429_ = ~Q[12] /*19947*/;
assign _46428_ = _46429_ & D[47] /*19946*/;
assign _46431_ = _45680_ & _46428_ /*19941*/;
assign _46432_ = _45680_ ^ _46428_ /*19944*/;
assign _46433_ = _46424_ & _46432_ /*19942*/;
assign _46128_ = _46424_ ^ _46432_ /*19943*/;
assign _46430_ = _46431_ | _46433_ /*19940*/;
assign _46435_ = ~Q[12] /*19939*/;
assign _46434_ = _46435_ & D[48] /*19938*/;
assign _46437_ = _45681_ & _46434_ /*19933*/;
assign _46438_ = _45681_ ^ _46434_ /*19936*/;
assign _46439_ = _46430_ & _46438_ /*19934*/;
assign _46129_ = _46430_ ^ _46438_ /*19935*/;
assign _46436_ = _46437_ | _46439_ /*19932*/;
assign _46441_ = ~Q[12] /*19931*/;
assign _46440_ = _46441_ & D[49] /*19930*/;
assign _46443_ = _45682_ & _46440_ /*19925*/;
assign _46444_ = _45682_ ^ _46440_ /*19928*/;
assign _46445_ = _46436_ & _46444_ /*19926*/;
assign _46130_ = _46436_ ^ _46444_ /*19927*/;
assign _46442_ = _46443_ | _46445_ /*19924*/;
assign _46447_ = ~Q[12] /*19923*/;
assign _46446_ = _46447_ & D[50] /*19922*/;
assign _46449_ = _45683_ & _46446_ /*19917*/;
assign _46450_ = _45683_ ^ _46446_ /*19920*/;
assign _46451_ = _46442_ & _46450_ /*19918*/;
assign _46131_ = _46442_ ^ _46450_ /*19919*/;
assign _46448_ = _46449_ | _46451_ /*19916*/;
assign _46453_ = ~Q[12] /*19915*/;
assign _46452_ = _46453_ & D[51] /*19914*/;
assign _46455_ = _45684_ & _46452_ /*19909*/;
assign _46456_ = _45684_ ^ _46452_ /*19912*/;
assign _46457_ = _46448_ & _46456_ /*19910*/;
assign _46132_ = _46448_ ^ _46456_ /*19911*/;
assign _46454_ = _46455_ | _46457_ /*19908*/;
assign _46459_ = ~Q[12] /*19907*/;
assign _46458_ = _46459_ & D[52] /*19906*/;
assign _46461_ = _45685_ & _46458_ /*19901*/;
assign _46462_ = _45685_ ^ _46458_ /*19904*/;
assign _46463_ = _46454_ & _46462_ /*19902*/;
assign _46133_ = _46454_ ^ _46462_ /*19903*/;
assign _46460_ = _46461_ | _46463_ /*19900*/;
assign _46465_ = ~Q[12] /*19899*/;
assign _46464_ = _46465_ & D[53] /*19898*/;
assign _46467_ = _45686_ & _46464_ /*19893*/;
assign _46468_ = _45686_ ^ _46464_ /*19896*/;
assign _46469_ = _46460_ & _46468_ /*19894*/;
assign _46134_ = _46460_ ^ _46468_ /*19895*/;
assign _46466_ = _46467_ | _46469_ /*19892*/;
assign _46471_ = ~Q[12] /*19891*/;
assign _46470_ = _46471_ & D[54] /*19890*/;
assign _46473_ = _45687_ & _46470_ /*19885*/;
assign _46474_ = _45687_ ^ _46470_ /*19888*/;
assign _46475_ = _46466_ & _46474_ /*19886*/;
assign _46135_ = _46466_ ^ _46474_ /*19887*/;
assign _46472_ = _46473_ | _46475_ /*19884*/;
assign _46477_ = ~Q[12] /*19883*/;
assign _46476_ = _46477_ & D[55] /*19882*/;
assign _46479_ = _45688_ & _46476_ /*19877*/;
assign _46480_ = _45688_ ^ _46476_ /*19880*/;
assign _46481_ = _46472_ & _46480_ /*19878*/;
assign _46136_ = _46472_ ^ _46480_ /*19879*/;
assign _46478_ = _46479_ | _46481_ /*19876*/;
assign _46483_ = ~Q[12] /*19875*/;
assign _46482_ = _46483_ & D[56] /*19874*/;
assign _46485_ = _45689_ & _46482_ /*19869*/;
assign _46486_ = _45689_ ^ _46482_ /*19872*/;
assign _46487_ = _46478_ & _46486_ /*19870*/;
assign _46137_ = _46478_ ^ _46486_ /*19871*/;
assign _46484_ = _46485_ | _46487_ /*19868*/;
assign _46489_ = ~Q[12] /*19867*/;
assign _46488_ = _46489_ & D[57] /*19866*/;
assign _46491_ = _45690_ & _46488_ /*19861*/;
assign _46492_ = _45690_ ^ _46488_ /*19864*/;
assign _46493_ = _46484_ & _46492_ /*19862*/;
assign _46138_ = _46484_ ^ _46492_ /*19863*/;
assign _46490_ = _46491_ | _46493_ /*19860*/;
assign _46495_ = ~Q[12] /*19859*/;
assign _46494_ = _46495_ & D[58] /*19858*/;
assign _46497_ = _45691_ & _46494_ /*19853*/;
assign _46498_ = _45691_ ^ _46494_ /*19856*/;
assign _46499_ = _46490_ & _46498_ /*19854*/;
assign _46139_ = _46490_ ^ _46498_ /*19855*/;
assign _46496_ = _46497_ | _46499_ /*19852*/;
assign _46501_ = ~Q[12] /*19851*/;
assign _46500_ = _46501_ & D[59] /*19850*/;
assign _46503_ = _45692_ & _46500_ /*19845*/;
assign _46504_ = _45692_ ^ _46500_ /*19848*/;
assign _46505_ = _46496_ & _46504_ /*19846*/;
assign _46140_ = _46496_ ^ _46504_ /*19847*/;
assign _46502_ = _46503_ | _46505_ /*19844*/;
assign _46507_ = ~Q[12] /*19843*/;
assign _46506_ = _46507_ & D[60] /*19842*/;
assign _46509_ = _45693_ & _46506_ /*19837*/;
assign _46510_ = _45693_ ^ _46506_ /*19840*/;
assign _46511_ = _46502_ & _46510_ /*19838*/;
assign _46141_ = _46502_ ^ _46510_ /*19839*/;
assign _46508_ = _46509_ | _46511_ /*19836*/;
assign _46513_ = ~Q[12] /*19835*/;
assign _46512_ = _46513_ & D[61] /*19834*/;
assign _46515_ = _45694_ & _46512_ /*19829*/;
assign _46516_ = _45694_ ^ _46512_ /*19832*/;
assign _46517_ = _46508_ & _46516_ /*19830*/;
assign _46142_ = _46508_ ^ _46516_ /*19831*/;
assign _46514_ = _46515_ | _46517_ /*19828*/;
assign _46519_ = ~Q[12] /*19827*/;
assign _46518_ = _46519_ & D[62] /*19826*/;
assign _46521_ = _45695_ & _46518_ /*19821*/;
assign _46522_ = _45695_ ^ _46518_ /*19824*/;
assign _46523_ = _46514_ & _46522_ /*19822*/;
assign _46143_ = _46514_ ^ _46522_ /*19823*/;
assign _46520_ = _46521_ | _46523_ /*19820*/;
assign _46525_ = ~Q[12] /*19819*/;
assign _46524_ = _46525_ & zeroWire /*19818*/;
assign _46526_ = _45696_ ^ _46524_ /*19816*/;
assign _46144_ = _46526_ ^ _46520_ /*19815*/;
assign _46597_ = ~D[0] /*19561*/;
assign _46594_ = R_0[11] & _46597_ /*19557*/;
assign _46595_ = R_0[11] ^ _46597_ /*19560*/;
assign _46596_ = oneWire & _46595_ /*19558*/;
assign _46529_ = oneWire ^ _46595_ /*19559*/;
assign _46593_ = _46594_ | _46596_ /*19556*/;
assign _46602_ = ~D[1] /*19555*/;
assign _46599_ = _46081_ & _46602_ /*19551*/;
assign _46600_ = _46081_ ^ _46602_ /*19554*/;
assign _46601_ = _46593_ & _46600_ /*19552*/;
assign _46530_ = _46593_ ^ _46600_ /*19553*/;
assign _46598_ = _46599_ | _46601_ /*19550*/;
assign _46607_ = ~D[2] /*19549*/;
assign _46604_ = _46082_ & _46607_ /*19545*/;
assign _46605_ = _46082_ ^ _46607_ /*19548*/;
assign _46606_ = _46598_ & _46605_ /*19546*/;
assign _46531_ = _46598_ ^ _46605_ /*19547*/;
assign _46603_ = _46604_ | _46606_ /*19544*/;
assign _46612_ = ~D[3] /*19543*/;
assign _46609_ = _46083_ & _46612_ /*19539*/;
assign _46610_ = _46083_ ^ _46612_ /*19542*/;
assign _46611_ = _46603_ & _46610_ /*19540*/;
assign _46532_ = _46603_ ^ _46610_ /*19541*/;
assign _46608_ = _46609_ | _46611_ /*19538*/;
assign _46617_ = ~D[4] /*19537*/;
assign _46614_ = _46084_ & _46617_ /*19533*/;
assign _46615_ = _46084_ ^ _46617_ /*19536*/;
assign _46616_ = _46608_ & _46615_ /*19534*/;
assign _46533_ = _46608_ ^ _46615_ /*19535*/;
assign _46613_ = _46614_ | _46616_ /*19532*/;
assign _46622_ = ~D[5] /*19531*/;
assign _46619_ = _46085_ & _46622_ /*19527*/;
assign _46620_ = _46085_ ^ _46622_ /*19530*/;
assign _46621_ = _46613_ & _46620_ /*19528*/;
assign _46534_ = _46613_ ^ _46620_ /*19529*/;
assign _46618_ = _46619_ | _46621_ /*19526*/;
assign _46627_ = ~D[6] /*19525*/;
assign _46624_ = _46086_ & _46627_ /*19521*/;
assign _46625_ = _46086_ ^ _46627_ /*19524*/;
assign _46626_ = _46618_ & _46625_ /*19522*/;
assign _46535_ = _46618_ ^ _46625_ /*19523*/;
assign _46623_ = _46624_ | _46626_ /*19520*/;
assign _46632_ = ~D[7] /*19519*/;
assign _46629_ = _46087_ & _46632_ /*19515*/;
assign _46630_ = _46087_ ^ _46632_ /*19518*/;
assign _46631_ = _46623_ & _46630_ /*19516*/;
assign _46536_ = _46623_ ^ _46630_ /*19517*/;
assign _46628_ = _46629_ | _46631_ /*19514*/;
assign _46637_ = ~D[8] /*19513*/;
assign _46634_ = _46088_ & _46637_ /*19509*/;
assign _46635_ = _46088_ ^ _46637_ /*19512*/;
assign _46636_ = _46628_ & _46635_ /*19510*/;
assign _46537_ = _46628_ ^ _46635_ /*19511*/;
assign _46633_ = _46634_ | _46636_ /*19508*/;
assign _46642_ = ~D[9] /*19507*/;
assign _46639_ = _46089_ & _46642_ /*19503*/;
assign _46640_ = _46089_ ^ _46642_ /*19506*/;
assign _46641_ = _46633_ & _46640_ /*19504*/;
assign _46538_ = _46633_ ^ _46640_ /*19505*/;
assign _46638_ = _46639_ | _46641_ /*19502*/;
assign _46647_ = ~D[10] /*19501*/;
assign _46644_ = _46090_ & _46647_ /*19497*/;
assign _46645_ = _46090_ ^ _46647_ /*19500*/;
assign _46646_ = _46638_ & _46645_ /*19498*/;
assign _46539_ = _46638_ ^ _46645_ /*19499*/;
assign _46643_ = _46644_ | _46646_ /*19496*/;
assign _46652_ = ~D[11] /*19495*/;
assign _46649_ = _46091_ & _46652_ /*19491*/;
assign _46650_ = _46091_ ^ _46652_ /*19494*/;
assign _46651_ = _46643_ & _46650_ /*19492*/;
assign _46540_ = _46643_ ^ _46650_ /*19493*/;
assign _46648_ = _46649_ | _46651_ /*19490*/;
assign _46657_ = ~D[12] /*19489*/;
assign _46654_ = _46092_ & _46657_ /*19485*/;
assign _46655_ = _46092_ ^ _46657_ /*19488*/;
assign _46656_ = _46648_ & _46655_ /*19486*/;
assign _46541_ = _46648_ ^ _46655_ /*19487*/;
assign _46653_ = _46654_ | _46656_ /*19484*/;
assign _46662_ = ~D[13] /*19483*/;
assign _46659_ = _46093_ & _46662_ /*19479*/;
assign _46660_ = _46093_ ^ _46662_ /*19482*/;
assign _46661_ = _46653_ & _46660_ /*19480*/;
assign _46542_ = _46653_ ^ _46660_ /*19481*/;
assign _46658_ = _46659_ | _46661_ /*19478*/;
assign _46667_ = ~D[14] /*19477*/;
assign _46664_ = _46094_ & _46667_ /*19473*/;
assign _46665_ = _46094_ ^ _46667_ /*19476*/;
assign _46666_ = _46658_ & _46665_ /*19474*/;
assign _46543_ = _46658_ ^ _46665_ /*19475*/;
assign _46663_ = _46664_ | _46666_ /*19472*/;
assign _46672_ = ~D[15] /*19471*/;
assign _46669_ = _46095_ & _46672_ /*19467*/;
assign _46670_ = _46095_ ^ _46672_ /*19470*/;
assign _46671_ = _46663_ & _46670_ /*19468*/;
assign _46544_ = _46663_ ^ _46670_ /*19469*/;
assign _46668_ = _46669_ | _46671_ /*19466*/;
assign _46677_ = ~D[16] /*19465*/;
assign _46674_ = _46096_ & _46677_ /*19461*/;
assign _46675_ = _46096_ ^ _46677_ /*19464*/;
assign _46676_ = _46668_ & _46675_ /*19462*/;
assign _46545_ = _46668_ ^ _46675_ /*19463*/;
assign _46673_ = _46674_ | _46676_ /*19460*/;
assign _46682_ = ~D[17] /*19459*/;
assign _46679_ = _46097_ & _46682_ /*19455*/;
assign _46680_ = _46097_ ^ _46682_ /*19458*/;
assign _46681_ = _46673_ & _46680_ /*19456*/;
assign _46546_ = _46673_ ^ _46680_ /*19457*/;
assign _46678_ = _46679_ | _46681_ /*19454*/;
assign _46687_ = ~D[18] /*19453*/;
assign _46684_ = _46098_ & _46687_ /*19449*/;
assign _46685_ = _46098_ ^ _46687_ /*19452*/;
assign _46686_ = _46678_ & _46685_ /*19450*/;
assign _46547_ = _46678_ ^ _46685_ /*19451*/;
assign _46683_ = _46684_ | _46686_ /*19448*/;
assign _46692_ = ~D[19] /*19447*/;
assign _46689_ = _46099_ & _46692_ /*19443*/;
assign _46690_ = _46099_ ^ _46692_ /*19446*/;
assign _46691_ = _46683_ & _46690_ /*19444*/;
assign _46548_ = _46683_ ^ _46690_ /*19445*/;
assign _46688_ = _46689_ | _46691_ /*19442*/;
assign _46697_ = ~D[20] /*19441*/;
assign _46694_ = _46100_ & _46697_ /*19437*/;
assign _46695_ = _46100_ ^ _46697_ /*19440*/;
assign _46696_ = _46688_ & _46695_ /*19438*/;
assign _46549_ = _46688_ ^ _46695_ /*19439*/;
assign _46693_ = _46694_ | _46696_ /*19436*/;
assign _46702_ = ~D[21] /*19435*/;
assign _46699_ = _46101_ & _46702_ /*19431*/;
assign _46700_ = _46101_ ^ _46702_ /*19434*/;
assign _46701_ = _46693_ & _46700_ /*19432*/;
assign _46550_ = _46693_ ^ _46700_ /*19433*/;
assign _46698_ = _46699_ | _46701_ /*19430*/;
assign _46707_ = ~D[22] /*19429*/;
assign _46704_ = _46102_ & _46707_ /*19425*/;
assign _46705_ = _46102_ ^ _46707_ /*19428*/;
assign _46706_ = _46698_ & _46705_ /*19426*/;
assign _46551_ = _46698_ ^ _46705_ /*19427*/;
assign _46703_ = _46704_ | _46706_ /*19424*/;
assign _46712_ = ~D[23] /*19423*/;
assign _46709_ = _46103_ & _46712_ /*19419*/;
assign _46710_ = _46103_ ^ _46712_ /*19422*/;
assign _46711_ = _46703_ & _46710_ /*19420*/;
assign _46552_ = _46703_ ^ _46710_ /*19421*/;
assign _46708_ = _46709_ | _46711_ /*19418*/;
assign _46717_ = ~D[24] /*19417*/;
assign _46714_ = _46104_ & _46717_ /*19413*/;
assign _46715_ = _46104_ ^ _46717_ /*19416*/;
assign _46716_ = _46708_ & _46715_ /*19414*/;
assign _46553_ = _46708_ ^ _46715_ /*19415*/;
assign _46713_ = _46714_ | _46716_ /*19412*/;
assign _46722_ = ~D[25] /*19411*/;
assign _46719_ = _46105_ & _46722_ /*19407*/;
assign _46720_ = _46105_ ^ _46722_ /*19410*/;
assign _46721_ = _46713_ & _46720_ /*19408*/;
assign _46554_ = _46713_ ^ _46720_ /*19409*/;
assign _46718_ = _46719_ | _46721_ /*19406*/;
assign _46727_ = ~D[26] /*19405*/;
assign _46724_ = _46106_ & _46727_ /*19401*/;
assign _46725_ = _46106_ ^ _46727_ /*19404*/;
assign _46726_ = _46718_ & _46725_ /*19402*/;
assign _46555_ = _46718_ ^ _46725_ /*19403*/;
assign _46723_ = _46724_ | _46726_ /*19400*/;
assign _46732_ = ~D[27] /*19399*/;
assign _46729_ = _46107_ & _46732_ /*19395*/;
assign _46730_ = _46107_ ^ _46732_ /*19398*/;
assign _46731_ = _46723_ & _46730_ /*19396*/;
assign _46556_ = _46723_ ^ _46730_ /*19397*/;
assign _46728_ = _46729_ | _46731_ /*19394*/;
assign _46737_ = ~D[28] /*19393*/;
assign _46734_ = _46108_ & _46737_ /*19389*/;
assign _46735_ = _46108_ ^ _46737_ /*19392*/;
assign _46736_ = _46728_ & _46735_ /*19390*/;
assign _46557_ = _46728_ ^ _46735_ /*19391*/;
assign _46733_ = _46734_ | _46736_ /*19388*/;
assign _46742_ = ~D[29] /*19387*/;
assign _46739_ = _46109_ & _46742_ /*19383*/;
assign _46740_ = _46109_ ^ _46742_ /*19386*/;
assign _46741_ = _46733_ & _46740_ /*19384*/;
assign _46558_ = _46733_ ^ _46740_ /*19385*/;
assign _46738_ = _46739_ | _46741_ /*19382*/;
assign _46747_ = ~D[30] /*19381*/;
assign _46744_ = _46110_ & _46747_ /*19377*/;
assign _46745_ = _46110_ ^ _46747_ /*19380*/;
assign _46746_ = _46738_ & _46745_ /*19378*/;
assign _46559_ = _46738_ ^ _46745_ /*19379*/;
assign _46743_ = _46744_ | _46746_ /*19376*/;
assign _46752_ = ~D[31] /*19375*/;
assign _46749_ = _46111_ & _46752_ /*19371*/;
assign _46750_ = _46111_ ^ _46752_ /*19374*/;
assign _46751_ = _46743_ & _46750_ /*19372*/;
assign _46560_ = _46743_ ^ _46750_ /*19373*/;
assign _46748_ = _46749_ | _46751_ /*19370*/;
assign _46757_ = ~D[32] /*19369*/;
assign _46754_ = _46112_ & _46757_ /*19365*/;
assign _46755_ = _46112_ ^ _46757_ /*19368*/;
assign _46756_ = _46748_ & _46755_ /*19366*/;
assign _46561_ = _46748_ ^ _46755_ /*19367*/;
assign _46753_ = _46754_ | _46756_ /*19364*/;
assign _46762_ = ~D[33] /*19363*/;
assign _46759_ = _46113_ & _46762_ /*19359*/;
assign _46760_ = _46113_ ^ _46762_ /*19362*/;
assign _46761_ = _46753_ & _46760_ /*19360*/;
assign _46562_ = _46753_ ^ _46760_ /*19361*/;
assign _46758_ = _46759_ | _46761_ /*19358*/;
assign _46767_ = ~D[34] /*19357*/;
assign _46764_ = _46114_ & _46767_ /*19353*/;
assign _46765_ = _46114_ ^ _46767_ /*19356*/;
assign _46766_ = _46758_ & _46765_ /*19354*/;
assign _46563_ = _46758_ ^ _46765_ /*19355*/;
assign _46763_ = _46764_ | _46766_ /*19352*/;
assign _46772_ = ~D[35] /*19351*/;
assign _46769_ = _46115_ & _46772_ /*19347*/;
assign _46770_ = _46115_ ^ _46772_ /*19350*/;
assign _46771_ = _46763_ & _46770_ /*19348*/;
assign _46564_ = _46763_ ^ _46770_ /*19349*/;
assign _46768_ = _46769_ | _46771_ /*19346*/;
assign _46777_ = ~D[36] /*19345*/;
assign _46774_ = _46116_ & _46777_ /*19341*/;
assign _46775_ = _46116_ ^ _46777_ /*19344*/;
assign _46776_ = _46768_ & _46775_ /*19342*/;
assign _46565_ = _46768_ ^ _46775_ /*19343*/;
assign _46773_ = _46774_ | _46776_ /*19340*/;
assign _46782_ = ~D[37] /*19339*/;
assign _46779_ = _46117_ & _46782_ /*19335*/;
assign _46780_ = _46117_ ^ _46782_ /*19338*/;
assign _46781_ = _46773_ & _46780_ /*19336*/;
assign _46566_ = _46773_ ^ _46780_ /*19337*/;
assign _46778_ = _46779_ | _46781_ /*19334*/;
assign _46787_ = ~D[38] /*19333*/;
assign _46784_ = _46118_ & _46787_ /*19329*/;
assign _46785_ = _46118_ ^ _46787_ /*19332*/;
assign _46786_ = _46778_ & _46785_ /*19330*/;
assign _46567_ = _46778_ ^ _46785_ /*19331*/;
assign _46783_ = _46784_ | _46786_ /*19328*/;
assign _46792_ = ~D[39] /*19327*/;
assign _46789_ = _46119_ & _46792_ /*19323*/;
assign _46790_ = _46119_ ^ _46792_ /*19326*/;
assign _46791_ = _46783_ & _46790_ /*19324*/;
assign _46568_ = _46783_ ^ _46790_ /*19325*/;
assign _46788_ = _46789_ | _46791_ /*19322*/;
assign _46797_ = ~D[40] /*19321*/;
assign _46794_ = _46120_ & _46797_ /*19317*/;
assign _46795_ = _46120_ ^ _46797_ /*19320*/;
assign _46796_ = _46788_ & _46795_ /*19318*/;
assign _46569_ = _46788_ ^ _46795_ /*19319*/;
assign _46793_ = _46794_ | _46796_ /*19316*/;
assign _46802_ = ~D[41] /*19315*/;
assign _46799_ = _46121_ & _46802_ /*19311*/;
assign _46800_ = _46121_ ^ _46802_ /*19314*/;
assign _46801_ = _46793_ & _46800_ /*19312*/;
assign _46570_ = _46793_ ^ _46800_ /*19313*/;
assign _46798_ = _46799_ | _46801_ /*19310*/;
assign _46807_ = ~D[42] /*19309*/;
assign _46804_ = _46122_ & _46807_ /*19305*/;
assign _46805_ = _46122_ ^ _46807_ /*19308*/;
assign _46806_ = _46798_ & _46805_ /*19306*/;
assign _46571_ = _46798_ ^ _46805_ /*19307*/;
assign _46803_ = _46804_ | _46806_ /*19304*/;
assign _46812_ = ~D[43] /*19303*/;
assign _46809_ = _46123_ & _46812_ /*19299*/;
assign _46810_ = _46123_ ^ _46812_ /*19302*/;
assign _46811_ = _46803_ & _46810_ /*19300*/;
assign _46572_ = _46803_ ^ _46810_ /*19301*/;
assign _46808_ = _46809_ | _46811_ /*19298*/;
assign _46817_ = ~D[44] /*19297*/;
assign _46814_ = _46124_ & _46817_ /*19293*/;
assign _46815_ = _46124_ ^ _46817_ /*19296*/;
assign _46816_ = _46808_ & _46815_ /*19294*/;
assign _46573_ = _46808_ ^ _46815_ /*19295*/;
assign _46813_ = _46814_ | _46816_ /*19292*/;
assign _46822_ = ~D[45] /*19291*/;
assign _46819_ = _46125_ & _46822_ /*19287*/;
assign _46820_ = _46125_ ^ _46822_ /*19290*/;
assign _46821_ = _46813_ & _46820_ /*19288*/;
assign _46574_ = _46813_ ^ _46820_ /*19289*/;
assign _46818_ = _46819_ | _46821_ /*19286*/;
assign _46827_ = ~D[46] /*19285*/;
assign _46824_ = _46126_ & _46827_ /*19281*/;
assign _46825_ = _46126_ ^ _46827_ /*19284*/;
assign _46826_ = _46818_ & _46825_ /*19282*/;
assign _46575_ = _46818_ ^ _46825_ /*19283*/;
assign _46823_ = _46824_ | _46826_ /*19280*/;
assign _46832_ = ~D[47] /*19279*/;
assign _46829_ = _46127_ & _46832_ /*19275*/;
assign _46830_ = _46127_ ^ _46832_ /*19278*/;
assign _46831_ = _46823_ & _46830_ /*19276*/;
assign _46576_ = _46823_ ^ _46830_ /*19277*/;
assign _46828_ = _46829_ | _46831_ /*19274*/;
assign _46837_ = ~D[48] /*19273*/;
assign _46834_ = _46128_ & _46837_ /*19269*/;
assign _46835_ = _46128_ ^ _46837_ /*19272*/;
assign _46836_ = _46828_ & _46835_ /*19270*/;
assign _46577_ = _46828_ ^ _46835_ /*19271*/;
assign _46833_ = _46834_ | _46836_ /*19268*/;
assign _46842_ = ~D[49] /*19267*/;
assign _46839_ = _46129_ & _46842_ /*19263*/;
assign _46840_ = _46129_ ^ _46842_ /*19266*/;
assign _46841_ = _46833_ & _46840_ /*19264*/;
assign _46578_ = _46833_ ^ _46840_ /*19265*/;
assign _46838_ = _46839_ | _46841_ /*19262*/;
assign _46847_ = ~D[50] /*19261*/;
assign _46844_ = _46130_ & _46847_ /*19257*/;
assign _46845_ = _46130_ ^ _46847_ /*19260*/;
assign _46846_ = _46838_ & _46845_ /*19258*/;
assign _46579_ = _46838_ ^ _46845_ /*19259*/;
assign _46843_ = _46844_ | _46846_ /*19256*/;
assign _46852_ = ~D[51] /*19255*/;
assign _46849_ = _46131_ & _46852_ /*19251*/;
assign _46850_ = _46131_ ^ _46852_ /*19254*/;
assign _46851_ = _46843_ & _46850_ /*19252*/;
assign _46580_ = _46843_ ^ _46850_ /*19253*/;
assign _46848_ = _46849_ | _46851_ /*19250*/;
assign _46857_ = ~D[52] /*19249*/;
assign _46854_ = _46132_ & _46857_ /*19245*/;
assign _46855_ = _46132_ ^ _46857_ /*19248*/;
assign _46856_ = _46848_ & _46855_ /*19246*/;
assign _46581_ = _46848_ ^ _46855_ /*19247*/;
assign _46853_ = _46854_ | _46856_ /*19244*/;
assign _46862_ = ~D[53] /*19243*/;
assign _46859_ = _46133_ & _46862_ /*19239*/;
assign _46860_ = _46133_ ^ _46862_ /*19242*/;
assign _46861_ = _46853_ & _46860_ /*19240*/;
assign _46582_ = _46853_ ^ _46860_ /*19241*/;
assign _46858_ = _46859_ | _46861_ /*19238*/;
assign _46867_ = ~D[54] /*19237*/;
assign _46864_ = _46134_ & _46867_ /*19233*/;
assign _46865_ = _46134_ ^ _46867_ /*19236*/;
assign _46866_ = _46858_ & _46865_ /*19234*/;
assign _46583_ = _46858_ ^ _46865_ /*19235*/;
assign _46863_ = _46864_ | _46866_ /*19232*/;
assign _46872_ = ~D[55] /*19231*/;
assign _46869_ = _46135_ & _46872_ /*19227*/;
assign _46870_ = _46135_ ^ _46872_ /*19230*/;
assign _46871_ = _46863_ & _46870_ /*19228*/;
assign _46584_ = _46863_ ^ _46870_ /*19229*/;
assign _46868_ = _46869_ | _46871_ /*19226*/;
assign _46877_ = ~D[56] /*19225*/;
assign _46874_ = _46136_ & _46877_ /*19221*/;
assign _46875_ = _46136_ ^ _46877_ /*19224*/;
assign _46876_ = _46868_ & _46875_ /*19222*/;
assign _46585_ = _46868_ ^ _46875_ /*19223*/;
assign _46873_ = _46874_ | _46876_ /*19220*/;
assign _46882_ = ~D[57] /*19219*/;
assign _46879_ = _46137_ & _46882_ /*19215*/;
assign _46880_ = _46137_ ^ _46882_ /*19218*/;
assign _46881_ = _46873_ & _46880_ /*19216*/;
assign _46586_ = _46873_ ^ _46880_ /*19217*/;
assign _46878_ = _46879_ | _46881_ /*19214*/;
assign _46887_ = ~D[58] /*19213*/;
assign _46884_ = _46138_ & _46887_ /*19209*/;
assign _46885_ = _46138_ ^ _46887_ /*19212*/;
assign _46886_ = _46878_ & _46885_ /*19210*/;
assign _46587_ = _46878_ ^ _46885_ /*19211*/;
assign _46883_ = _46884_ | _46886_ /*19208*/;
assign _46892_ = ~D[59] /*19207*/;
assign _46889_ = _46139_ & _46892_ /*19203*/;
assign _46890_ = _46139_ ^ _46892_ /*19206*/;
assign _46891_ = _46883_ & _46890_ /*19204*/;
assign _46588_ = _46883_ ^ _46890_ /*19205*/;
assign _46888_ = _46889_ | _46891_ /*19202*/;
assign _46897_ = ~D[60] /*19201*/;
assign _46894_ = _46140_ & _46897_ /*19197*/;
assign _46895_ = _46140_ ^ _46897_ /*19200*/;
assign _46896_ = _46888_ & _46895_ /*19198*/;
assign _46589_ = _46888_ ^ _46895_ /*19199*/;
assign _46893_ = _46894_ | _46896_ /*19196*/;
assign _46902_ = ~D[61] /*19195*/;
assign _46899_ = _46141_ & _46902_ /*19191*/;
assign _46900_ = _46141_ ^ _46902_ /*19194*/;
assign _46901_ = _46893_ & _46900_ /*19192*/;
assign _46590_ = _46893_ ^ _46900_ /*19193*/;
assign _46898_ = _46899_ | _46901_ /*19190*/;
assign _46907_ = ~D[62] /*19189*/;
assign _46904_ = _46142_ & _46907_ /*19185*/;
assign _46905_ = _46142_ ^ _46907_ /*19188*/;
assign _46906_ = _46898_ & _46905_ /*19186*/;
assign _46591_ = _46898_ ^ _46905_ /*19187*/;
assign _46903_ = _46904_ | _46906_ /*19184*/;
assign _46908_ = _46143_ & oneWire /*19179*/;
assign _46909_ = _46143_ ^ oneWire /*19182*/;
assign _46910_ = _46903_ & _46909_ /*19180*/;
assign _46592_ = _46903_ ^ _46909_ /*19181*/;
assign Q[11] = _46908_ | _46910_ /*19178*/;
assign _47043_ = ~Q[11] /*18793*/;
assign _47042_ = _47043_ & D[0] /*18792*/;
assign _47045_ = _46529_ & _47042_ /*18787*/;
assign _47046_ = _46529_ ^ _47042_ /*18790*/;
assign _47047_ = zeroWire & _47046_ /*18788*/;
assign _46977_ = zeroWire ^ _47046_ /*18789*/;
assign _47044_ = _47045_ | _47047_ /*18786*/;
assign _47049_ = ~Q[11] /*18785*/;
assign _47048_ = _47049_ & D[1] /*18784*/;
assign _47051_ = _46530_ & _47048_ /*18779*/;
assign _47052_ = _46530_ ^ _47048_ /*18782*/;
assign _47053_ = _47044_ & _47052_ /*18780*/;
assign _46978_ = _47044_ ^ _47052_ /*18781*/;
assign _47050_ = _47051_ | _47053_ /*18778*/;
assign _47055_ = ~Q[11] /*18777*/;
assign _47054_ = _47055_ & D[2] /*18776*/;
assign _47057_ = _46531_ & _47054_ /*18771*/;
assign _47058_ = _46531_ ^ _47054_ /*18774*/;
assign _47059_ = _47050_ & _47058_ /*18772*/;
assign _46979_ = _47050_ ^ _47058_ /*18773*/;
assign _47056_ = _47057_ | _47059_ /*18770*/;
assign _47061_ = ~Q[11] /*18769*/;
assign _47060_ = _47061_ & D[3] /*18768*/;
assign _47063_ = _46532_ & _47060_ /*18763*/;
assign _47064_ = _46532_ ^ _47060_ /*18766*/;
assign _47065_ = _47056_ & _47064_ /*18764*/;
assign _46980_ = _47056_ ^ _47064_ /*18765*/;
assign _47062_ = _47063_ | _47065_ /*18762*/;
assign _47067_ = ~Q[11] /*18761*/;
assign _47066_ = _47067_ & D[4] /*18760*/;
assign _47069_ = _46533_ & _47066_ /*18755*/;
assign _47070_ = _46533_ ^ _47066_ /*18758*/;
assign _47071_ = _47062_ & _47070_ /*18756*/;
assign _46981_ = _47062_ ^ _47070_ /*18757*/;
assign _47068_ = _47069_ | _47071_ /*18754*/;
assign _47073_ = ~Q[11] /*18753*/;
assign _47072_ = _47073_ & D[5] /*18752*/;
assign _47075_ = _46534_ & _47072_ /*18747*/;
assign _47076_ = _46534_ ^ _47072_ /*18750*/;
assign _47077_ = _47068_ & _47076_ /*18748*/;
assign _46982_ = _47068_ ^ _47076_ /*18749*/;
assign _47074_ = _47075_ | _47077_ /*18746*/;
assign _47079_ = ~Q[11] /*18745*/;
assign _47078_ = _47079_ & D[6] /*18744*/;
assign _47081_ = _46535_ & _47078_ /*18739*/;
assign _47082_ = _46535_ ^ _47078_ /*18742*/;
assign _47083_ = _47074_ & _47082_ /*18740*/;
assign _46983_ = _47074_ ^ _47082_ /*18741*/;
assign _47080_ = _47081_ | _47083_ /*18738*/;
assign _47085_ = ~Q[11] /*18737*/;
assign _47084_ = _47085_ & D[7] /*18736*/;
assign _47087_ = _46536_ & _47084_ /*18731*/;
assign _47088_ = _46536_ ^ _47084_ /*18734*/;
assign _47089_ = _47080_ & _47088_ /*18732*/;
assign _46984_ = _47080_ ^ _47088_ /*18733*/;
assign _47086_ = _47087_ | _47089_ /*18730*/;
assign _47091_ = ~Q[11] /*18729*/;
assign _47090_ = _47091_ & D[8] /*18728*/;
assign _47093_ = _46537_ & _47090_ /*18723*/;
assign _47094_ = _46537_ ^ _47090_ /*18726*/;
assign _47095_ = _47086_ & _47094_ /*18724*/;
assign _46985_ = _47086_ ^ _47094_ /*18725*/;
assign _47092_ = _47093_ | _47095_ /*18722*/;
assign _47097_ = ~Q[11] /*18721*/;
assign _47096_ = _47097_ & D[9] /*18720*/;
assign _47099_ = _46538_ & _47096_ /*18715*/;
assign _47100_ = _46538_ ^ _47096_ /*18718*/;
assign _47101_ = _47092_ & _47100_ /*18716*/;
assign _46986_ = _47092_ ^ _47100_ /*18717*/;
assign _47098_ = _47099_ | _47101_ /*18714*/;
assign _47103_ = ~Q[11] /*18713*/;
assign _47102_ = _47103_ & D[10] /*18712*/;
assign _47105_ = _46539_ & _47102_ /*18707*/;
assign _47106_ = _46539_ ^ _47102_ /*18710*/;
assign _47107_ = _47098_ & _47106_ /*18708*/;
assign _46987_ = _47098_ ^ _47106_ /*18709*/;
assign _47104_ = _47105_ | _47107_ /*18706*/;
assign _47109_ = ~Q[11] /*18705*/;
assign _47108_ = _47109_ & D[11] /*18704*/;
assign _47111_ = _46540_ & _47108_ /*18699*/;
assign _47112_ = _46540_ ^ _47108_ /*18702*/;
assign _47113_ = _47104_ & _47112_ /*18700*/;
assign _46988_ = _47104_ ^ _47112_ /*18701*/;
assign _47110_ = _47111_ | _47113_ /*18698*/;
assign _47115_ = ~Q[11] /*18697*/;
assign _47114_ = _47115_ & D[12] /*18696*/;
assign _47117_ = _46541_ & _47114_ /*18691*/;
assign _47118_ = _46541_ ^ _47114_ /*18694*/;
assign _47119_ = _47110_ & _47118_ /*18692*/;
assign _46989_ = _47110_ ^ _47118_ /*18693*/;
assign _47116_ = _47117_ | _47119_ /*18690*/;
assign _47121_ = ~Q[11] /*18689*/;
assign _47120_ = _47121_ & D[13] /*18688*/;
assign _47123_ = _46542_ & _47120_ /*18683*/;
assign _47124_ = _46542_ ^ _47120_ /*18686*/;
assign _47125_ = _47116_ & _47124_ /*18684*/;
assign _46990_ = _47116_ ^ _47124_ /*18685*/;
assign _47122_ = _47123_ | _47125_ /*18682*/;
assign _47127_ = ~Q[11] /*18681*/;
assign _47126_ = _47127_ & D[14] /*18680*/;
assign _47129_ = _46543_ & _47126_ /*18675*/;
assign _47130_ = _46543_ ^ _47126_ /*18678*/;
assign _47131_ = _47122_ & _47130_ /*18676*/;
assign _46991_ = _47122_ ^ _47130_ /*18677*/;
assign _47128_ = _47129_ | _47131_ /*18674*/;
assign _47133_ = ~Q[11] /*18673*/;
assign _47132_ = _47133_ & D[15] /*18672*/;
assign _47135_ = _46544_ & _47132_ /*18667*/;
assign _47136_ = _46544_ ^ _47132_ /*18670*/;
assign _47137_ = _47128_ & _47136_ /*18668*/;
assign _46992_ = _47128_ ^ _47136_ /*18669*/;
assign _47134_ = _47135_ | _47137_ /*18666*/;
assign _47139_ = ~Q[11] /*18665*/;
assign _47138_ = _47139_ & D[16] /*18664*/;
assign _47141_ = _46545_ & _47138_ /*18659*/;
assign _47142_ = _46545_ ^ _47138_ /*18662*/;
assign _47143_ = _47134_ & _47142_ /*18660*/;
assign _46993_ = _47134_ ^ _47142_ /*18661*/;
assign _47140_ = _47141_ | _47143_ /*18658*/;
assign _47145_ = ~Q[11] /*18657*/;
assign _47144_ = _47145_ & D[17] /*18656*/;
assign _47147_ = _46546_ & _47144_ /*18651*/;
assign _47148_ = _46546_ ^ _47144_ /*18654*/;
assign _47149_ = _47140_ & _47148_ /*18652*/;
assign _46994_ = _47140_ ^ _47148_ /*18653*/;
assign _47146_ = _47147_ | _47149_ /*18650*/;
assign _47151_ = ~Q[11] /*18649*/;
assign _47150_ = _47151_ & D[18] /*18648*/;
assign _47153_ = _46547_ & _47150_ /*18643*/;
assign _47154_ = _46547_ ^ _47150_ /*18646*/;
assign _47155_ = _47146_ & _47154_ /*18644*/;
assign _46995_ = _47146_ ^ _47154_ /*18645*/;
assign _47152_ = _47153_ | _47155_ /*18642*/;
assign _47157_ = ~Q[11] /*18641*/;
assign _47156_ = _47157_ & D[19] /*18640*/;
assign _47159_ = _46548_ & _47156_ /*18635*/;
assign _47160_ = _46548_ ^ _47156_ /*18638*/;
assign _47161_ = _47152_ & _47160_ /*18636*/;
assign _46996_ = _47152_ ^ _47160_ /*18637*/;
assign _47158_ = _47159_ | _47161_ /*18634*/;
assign _47163_ = ~Q[11] /*18633*/;
assign _47162_ = _47163_ & D[20] /*18632*/;
assign _47165_ = _46549_ & _47162_ /*18627*/;
assign _47166_ = _46549_ ^ _47162_ /*18630*/;
assign _47167_ = _47158_ & _47166_ /*18628*/;
assign _46997_ = _47158_ ^ _47166_ /*18629*/;
assign _47164_ = _47165_ | _47167_ /*18626*/;
assign _47169_ = ~Q[11] /*18625*/;
assign _47168_ = _47169_ & D[21] /*18624*/;
assign _47171_ = _46550_ & _47168_ /*18619*/;
assign _47172_ = _46550_ ^ _47168_ /*18622*/;
assign _47173_ = _47164_ & _47172_ /*18620*/;
assign _46998_ = _47164_ ^ _47172_ /*18621*/;
assign _47170_ = _47171_ | _47173_ /*18618*/;
assign _47175_ = ~Q[11] /*18617*/;
assign _47174_ = _47175_ & D[22] /*18616*/;
assign _47177_ = _46551_ & _47174_ /*18611*/;
assign _47178_ = _46551_ ^ _47174_ /*18614*/;
assign _47179_ = _47170_ & _47178_ /*18612*/;
assign _46999_ = _47170_ ^ _47178_ /*18613*/;
assign _47176_ = _47177_ | _47179_ /*18610*/;
assign _47181_ = ~Q[11] /*18609*/;
assign _47180_ = _47181_ & D[23] /*18608*/;
assign _47183_ = _46552_ & _47180_ /*18603*/;
assign _47184_ = _46552_ ^ _47180_ /*18606*/;
assign _47185_ = _47176_ & _47184_ /*18604*/;
assign _47000_ = _47176_ ^ _47184_ /*18605*/;
assign _47182_ = _47183_ | _47185_ /*18602*/;
assign _47187_ = ~Q[11] /*18601*/;
assign _47186_ = _47187_ & D[24] /*18600*/;
assign _47189_ = _46553_ & _47186_ /*18595*/;
assign _47190_ = _46553_ ^ _47186_ /*18598*/;
assign _47191_ = _47182_ & _47190_ /*18596*/;
assign _47001_ = _47182_ ^ _47190_ /*18597*/;
assign _47188_ = _47189_ | _47191_ /*18594*/;
assign _47193_ = ~Q[11] /*18593*/;
assign _47192_ = _47193_ & D[25] /*18592*/;
assign _47195_ = _46554_ & _47192_ /*18587*/;
assign _47196_ = _46554_ ^ _47192_ /*18590*/;
assign _47197_ = _47188_ & _47196_ /*18588*/;
assign _47002_ = _47188_ ^ _47196_ /*18589*/;
assign _47194_ = _47195_ | _47197_ /*18586*/;
assign _47199_ = ~Q[11] /*18585*/;
assign _47198_ = _47199_ & D[26] /*18584*/;
assign _47201_ = _46555_ & _47198_ /*18579*/;
assign _47202_ = _46555_ ^ _47198_ /*18582*/;
assign _47203_ = _47194_ & _47202_ /*18580*/;
assign _47003_ = _47194_ ^ _47202_ /*18581*/;
assign _47200_ = _47201_ | _47203_ /*18578*/;
assign _47205_ = ~Q[11] /*18577*/;
assign _47204_ = _47205_ & D[27] /*18576*/;
assign _47207_ = _46556_ & _47204_ /*18571*/;
assign _47208_ = _46556_ ^ _47204_ /*18574*/;
assign _47209_ = _47200_ & _47208_ /*18572*/;
assign _47004_ = _47200_ ^ _47208_ /*18573*/;
assign _47206_ = _47207_ | _47209_ /*18570*/;
assign _47211_ = ~Q[11] /*18569*/;
assign _47210_ = _47211_ & D[28] /*18568*/;
assign _47213_ = _46557_ & _47210_ /*18563*/;
assign _47214_ = _46557_ ^ _47210_ /*18566*/;
assign _47215_ = _47206_ & _47214_ /*18564*/;
assign _47005_ = _47206_ ^ _47214_ /*18565*/;
assign _47212_ = _47213_ | _47215_ /*18562*/;
assign _47217_ = ~Q[11] /*18561*/;
assign _47216_ = _47217_ & D[29] /*18560*/;
assign _47219_ = _46558_ & _47216_ /*18555*/;
assign _47220_ = _46558_ ^ _47216_ /*18558*/;
assign _47221_ = _47212_ & _47220_ /*18556*/;
assign _47006_ = _47212_ ^ _47220_ /*18557*/;
assign _47218_ = _47219_ | _47221_ /*18554*/;
assign _47223_ = ~Q[11] /*18553*/;
assign _47222_ = _47223_ & D[30] /*18552*/;
assign _47225_ = _46559_ & _47222_ /*18547*/;
assign _47226_ = _46559_ ^ _47222_ /*18550*/;
assign _47227_ = _47218_ & _47226_ /*18548*/;
assign _47007_ = _47218_ ^ _47226_ /*18549*/;
assign _47224_ = _47225_ | _47227_ /*18546*/;
assign _47229_ = ~Q[11] /*18545*/;
assign _47228_ = _47229_ & D[31] /*18544*/;
assign _47231_ = _46560_ & _47228_ /*18539*/;
assign _47232_ = _46560_ ^ _47228_ /*18542*/;
assign _47233_ = _47224_ & _47232_ /*18540*/;
assign _47008_ = _47224_ ^ _47232_ /*18541*/;
assign _47230_ = _47231_ | _47233_ /*18538*/;
assign _47235_ = ~Q[11] /*18537*/;
assign _47234_ = _47235_ & D[32] /*18536*/;
assign _47237_ = _46561_ & _47234_ /*18531*/;
assign _47238_ = _46561_ ^ _47234_ /*18534*/;
assign _47239_ = _47230_ & _47238_ /*18532*/;
assign _47009_ = _47230_ ^ _47238_ /*18533*/;
assign _47236_ = _47237_ | _47239_ /*18530*/;
assign _47241_ = ~Q[11] /*18529*/;
assign _47240_ = _47241_ & D[33] /*18528*/;
assign _47243_ = _46562_ & _47240_ /*18523*/;
assign _47244_ = _46562_ ^ _47240_ /*18526*/;
assign _47245_ = _47236_ & _47244_ /*18524*/;
assign _47010_ = _47236_ ^ _47244_ /*18525*/;
assign _47242_ = _47243_ | _47245_ /*18522*/;
assign _47247_ = ~Q[11] /*18521*/;
assign _47246_ = _47247_ & D[34] /*18520*/;
assign _47249_ = _46563_ & _47246_ /*18515*/;
assign _47250_ = _46563_ ^ _47246_ /*18518*/;
assign _47251_ = _47242_ & _47250_ /*18516*/;
assign _47011_ = _47242_ ^ _47250_ /*18517*/;
assign _47248_ = _47249_ | _47251_ /*18514*/;
assign _47253_ = ~Q[11] /*18513*/;
assign _47252_ = _47253_ & D[35] /*18512*/;
assign _47255_ = _46564_ & _47252_ /*18507*/;
assign _47256_ = _46564_ ^ _47252_ /*18510*/;
assign _47257_ = _47248_ & _47256_ /*18508*/;
assign _47012_ = _47248_ ^ _47256_ /*18509*/;
assign _47254_ = _47255_ | _47257_ /*18506*/;
assign _47259_ = ~Q[11] /*18505*/;
assign _47258_ = _47259_ & D[36] /*18504*/;
assign _47261_ = _46565_ & _47258_ /*18499*/;
assign _47262_ = _46565_ ^ _47258_ /*18502*/;
assign _47263_ = _47254_ & _47262_ /*18500*/;
assign _47013_ = _47254_ ^ _47262_ /*18501*/;
assign _47260_ = _47261_ | _47263_ /*18498*/;
assign _47265_ = ~Q[11] /*18497*/;
assign _47264_ = _47265_ & D[37] /*18496*/;
assign _47267_ = _46566_ & _47264_ /*18491*/;
assign _47268_ = _46566_ ^ _47264_ /*18494*/;
assign _47269_ = _47260_ & _47268_ /*18492*/;
assign _47014_ = _47260_ ^ _47268_ /*18493*/;
assign _47266_ = _47267_ | _47269_ /*18490*/;
assign _47271_ = ~Q[11] /*18489*/;
assign _47270_ = _47271_ & D[38] /*18488*/;
assign _47273_ = _46567_ & _47270_ /*18483*/;
assign _47274_ = _46567_ ^ _47270_ /*18486*/;
assign _47275_ = _47266_ & _47274_ /*18484*/;
assign _47015_ = _47266_ ^ _47274_ /*18485*/;
assign _47272_ = _47273_ | _47275_ /*18482*/;
assign _47277_ = ~Q[11] /*18481*/;
assign _47276_ = _47277_ & D[39] /*18480*/;
assign _47279_ = _46568_ & _47276_ /*18475*/;
assign _47280_ = _46568_ ^ _47276_ /*18478*/;
assign _47281_ = _47272_ & _47280_ /*18476*/;
assign _47016_ = _47272_ ^ _47280_ /*18477*/;
assign _47278_ = _47279_ | _47281_ /*18474*/;
assign _47283_ = ~Q[11] /*18473*/;
assign _47282_ = _47283_ & D[40] /*18472*/;
assign _47285_ = _46569_ & _47282_ /*18467*/;
assign _47286_ = _46569_ ^ _47282_ /*18470*/;
assign _47287_ = _47278_ & _47286_ /*18468*/;
assign _47017_ = _47278_ ^ _47286_ /*18469*/;
assign _47284_ = _47285_ | _47287_ /*18466*/;
assign _47289_ = ~Q[11] /*18465*/;
assign _47288_ = _47289_ & D[41] /*18464*/;
assign _47291_ = _46570_ & _47288_ /*18459*/;
assign _47292_ = _46570_ ^ _47288_ /*18462*/;
assign _47293_ = _47284_ & _47292_ /*18460*/;
assign _47018_ = _47284_ ^ _47292_ /*18461*/;
assign _47290_ = _47291_ | _47293_ /*18458*/;
assign _47295_ = ~Q[11] /*18457*/;
assign _47294_ = _47295_ & D[42] /*18456*/;
assign _47297_ = _46571_ & _47294_ /*18451*/;
assign _47298_ = _46571_ ^ _47294_ /*18454*/;
assign _47299_ = _47290_ & _47298_ /*18452*/;
assign _47019_ = _47290_ ^ _47298_ /*18453*/;
assign _47296_ = _47297_ | _47299_ /*18450*/;
assign _47301_ = ~Q[11] /*18449*/;
assign _47300_ = _47301_ & D[43] /*18448*/;
assign _47303_ = _46572_ & _47300_ /*18443*/;
assign _47304_ = _46572_ ^ _47300_ /*18446*/;
assign _47305_ = _47296_ & _47304_ /*18444*/;
assign _47020_ = _47296_ ^ _47304_ /*18445*/;
assign _47302_ = _47303_ | _47305_ /*18442*/;
assign _47307_ = ~Q[11] /*18441*/;
assign _47306_ = _47307_ & D[44] /*18440*/;
assign _47309_ = _46573_ & _47306_ /*18435*/;
assign _47310_ = _46573_ ^ _47306_ /*18438*/;
assign _47311_ = _47302_ & _47310_ /*18436*/;
assign _47021_ = _47302_ ^ _47310_ /*18437*/;
assign _47308_ = _47309_ | _47311_ /*18434*/;
assign _47313_ = ~Q[11] /*18433*/;
assign _47312_ = _47313_ & D[45] /*18432*/;
assign _47315_ = _46574_ & _47312_ /*18427*/;
assign _47316_ = _46574_ ^ _47312_ /*18430*/;
assign _47317_ = _47308_ & _47316_ /*18428*/;
assign _47022_ = _47308_ ^ _47316_ /*18429*/;
assign _47314_ = _47315_ | _47317_ /*18426*/;
assign _47319_ = ~Q[11] /*18425*/;
assign _47318_ = _47319_ & D[46] /*18424*/;
assign _47321_ = _46575_ & _47318_ /*18419*/;
assign _47322_ = _46575_ ^ _47318_ /*18422*/;
assign _47323_ = _47314_ & _47322_ /*18420*/;
assign _47023_ = _47314_ ^ _47322_ /*18421*/;
assign _47320_ = _47321_ | _47323_ /*18418*/;
assign _47325_ = ~Q[11] /*18417*/;
assign _47324_ = _47325_ & D[47] /*18416*/;
assign _47327_ = _46576_ & _47324_ /*18411*/;
assign _47328_ = _46576_ ^ _47324_ /*18414*/;
assign _47329_ = _47320_ & _47328_ /*18412*/;
assign _47024_ = _47320_ ^ _47328_ /*18413*/;
assign _47326_ = _47327_ | _47329_ /*18410*/;
assign _47331_ = ~Q[11] /*18409*/;
assign _47330_ = _47331_ & D[48] /*18408*/;
assign _47333_ = _46577_ & _47330_ /*18403*/;
assign _47334_ = _46577_ ^ _47330_ /*18406*/;
assign _47335_ = _47326_ & _47334_ /*18404*/;
assign _47025_ = _47326_ ^ _47334_ /*18405*/;
assign _47332_ = _47333_ | _47335_ /*18402*/;
assign _47337_ = ~Q[11] /*18401*/;
assign _47336_ = _47337_ & D[49] /*18400*/;
assign _47339_ = _46578_ & _47336_ /*18395*/;
assign _47340_ = _46578_ ^ _47336_ /*18398*/;
assign _47341_ = _47332_ & _47340_ /*18396*/;
assign _47026_ = _47332_ ^ _47340_ /*18397*/;
assign _47338_ = _47339_ | _47341_ /*18394*/;
assign _47343_ = ~Q[11] /*18393*/;
assign _47342_ = _47343_ & D[50] /*18392*/;
assign _47345_ = _46579_ & _47342_ /*18387*/;
assign _47346_ = _46579_ ^ _47342_ /*18390*/;
assign _47347_ = _47338_ & _47346_ /*18388*/;
assign _47027_ = _47338_ ^ _47346_ /*18389*/;
assign _47344_ = _47345_ | _47347_ /*18386*/;
assign _47349_ = ~Q[11] /*18385*/;
assign _47348_ = _47349_ & D[51] /*18384*/;
assign _47351_ = _46580_ & _47348_ /*18379*/;
assign _47352_ = _46580_ ^ _47348_ /*18382*/;
assign _47353_ = _47344_ & _47352_ /*18380*/;
assign _47028_ = _47344_ ^ _47352_ /*18381*/;
assign _47350_ = _47351_ | _47353_ /*18378*/;
assign _47355_ = ~Q[11] /*18377*/;
assign _47354_ = _47355_ & D[52] /*18376*/;
assign _47357_ = _46581_ & _47354_ /*18371*/;
assign _47358_ = _46581_ ^ _47354_ /*18374*/;
assign _47359_ = _47350_ & _47358_ /*18372*/;
assign _47029_ = _47350_ ^ _47358_ /*18373*/;
assign _47356_ = _47357_ | _47359_ /*18370*/;
assign _47361_ = ~Q[11] /*18369*/;
assign _47360_ = _47361_ & D[53] /*18368*/;
assign _47363_ = _46582_ & _47360_ /*18363*/;
assign _47364_ = _46582_ ^ _47360_ /*18366*/;
assign _47365_ = _47356_ & _47364_ /*18364*/;
assign _47030_ = _47356_ ^ _47364_ /*18365*/;
assign _47362_ = _47363_ | _47365_ /*18362*/;
assign _47367_ = ~Q[11] /*18361*/;
assign _47366_ = _47367_ & D[54] /*18360*/;
assign _47369_ = _46583_ & _47366_ /*18355*/;
assign _47370_ = _46583_ ^ _47366_ /*18358*/;
assign _47371_ = _47362_ & _47370_ /*18356*/;
assign _47031_ = _47362_ ^ _47370_ /*18357*/;
assign _47368_ = _47369_ | _47371_ /*18354*/;
assign _47373_ = ~Q[11] /*18353*/;
assign _47372_ = _47373_ & D[55] /*18352*/;
assign _47375_ = _46584_ & _47372_ /*18347*/;
assign _47376_ = _46584_ ^ _47372_ /*18350*/;
assign _47377_ = _47368_ & _47376_ /*18348*/;
assign _47032_ = _47368_ ^ _47376_ /*18349*/;
assign _47374_ = _47375_ | _47377_ /*18346*/;
assign _47379_ = ~Q[11] /*18345*/;
assign _47378_ = _47379_ & D[56] /*18344*/;
assign _47381_ = _46585_ & _47378_ /*18339*/;
assign _47382_ = _46585_ ^ _47378_ /*18342*/;
assign _47383_ = _47374_ & _47382_ /*18340*/;
assign _47033_ = _47374_ ^ _47382_ /*18341*/;
assign _47380_ = _47381_ | _47383_ /*18338*/;
assign _47385_ = ~Q[11] /*18337*/;
assign _47384_ = _47385_ & D[57] /*18336*/;
assign _47387_ = _46586_ & _47384_ /*18331*/;
assign _47388_ = _46586_ ^ _47384_ /*18334*/;
assign _47389_ = _47380_ & _47388_ /*18332*/;
assign _47034_ = _47380_ ^ _47388_ /*18333*/;
assign _47386_ = _47387_ | _47389_ /*18330*/;
assign _47391_ = ~Q[11] /*18329*/;
assign _47390_ = _47391_ & D[58] /*18328*/;
assign _47393_ = _46587_ & _47390_ /*18323*/;
assign _47394_ = _46587_ ^ _47390_ /*18326*/;
assign _47395_ = _47386_ & _47394_ /*18324*/;
assign _47035_ = _47386_ ^ _47394_ /*18325*/;
assign _47392_ = _47393_ | _47395_ /*18322*/;
assign _47397_ = ~Q[11] /*18321*/;
assign _47396_ = _47397_ & D[59] /*18320*/;
assign _47399_ = _46588_ & _47396_ /*18315*/;
assign _47400_ = _46588_ ^ _47396_ /*18318*/;
assign _47401_ = _47392_ & _47400_ /*18316*/;
assign _47036_ = _47392_ ^ _47400_ /*18317*/;
assign _47398_ = _47399_ | _47401_ /*18314*/;
assign _47403_ = ~Q[11] /*18313*/;
assign _47402_ = _47403_ & D[60] /*18312*/;
assign _47405_ = _46589_ & _47402_ /*18307*/;
assign _47406_ = _46589_ ^ _47402_ /*18310*/;
assign _47407_ = _47398_ & _47406_ /*18308*/;
assign _47037_ = _47398_ ^ _47406_ /*18309*/;
assign _47404_ = _47405_ | _47407_ /*18306*/;
assign _47409_ = ~Q[11] /*18305*/;
assign _47408_ = _47409_ & D[61] /*18304*/;
assign _47411_ = _46590_ & _47408_ /*18299*/;
assign _47412_ = _46590_ ^ _47408_ /*18302*/;
assign _47413_ = _47404_ & _47412_ /*18300*/;
assign _47038_ = _47404_ ^ _47412_ /*18301*/;
assign _47410_ = _47411_ | _47413_ /*18298*/;
assign _47415_ = ~Q[11] /*18297*/;
assign _47414_ = _47415_ & D[62] /*18296*/;
assign _47417_ = _46591_ & _47414_ /*18291*/;
assign _47418_ = _46591_ ^ _47414_ /*18294*/;
assign _47419_ = _47410_ & _47418_ /*18292*/;
assign _47039_ = _47410_ ^ _47418_ /*18293*/;
assign _47416_ = _47417_ | _47419_ /*18290*/;
assign _47421_ = ~Q[11] /*18289*/;
assign _47420_ = _47421_ & zeroWire /*18288*/;
assign _47422_ = _46592_ ^ _47420_ /*18286*/;
assign _47040_ = _47422_ ^ _47416_ /*18285*/;
assign _47493_ = ~D[0] /*18031*/;
assign _47490_ = R_0[10] & _47493_ /*18027*/;
assign _47491_ = R_0[10] ^ _47493_ /*18030*/;
assign _47492_ = oneWire & _47491_ /*18028*/;
assign _47425_ = oneWire ^ _47491_ /*18029*/;
assign _47489_ = _47490_ | _47492_ /*18026*/;
assign _47498_ = ~D[1] /*18025*/;
assign _47495_ = _46977_ & _47498_ /*18021*/;
assign _47496_ = _46977_ ^ _47498_ /*18024*/;
assign _47497_ = _47489_ & _47496_ /*18022*/;
assign _47426_ = _47489_ ^ _47496_ /*18023*/;
assign _47494_ = _47495_ | _47497_ /*18020*/;
assign _47503_ = ~D[2] /*18019*/;
assign _47500_ = _46978_ & _47503_ /*18015*/;
assign _47501_ = _46978_ ^ _47503_ /*18018*/;
assign _47502_ = _47494_ & _47501_ /*18016*/;
assign _47427_ = _47494_ ^ _47501_ /*18017*/;
assign _47499_ = _47500_ | _47502_ /*18014*/;
assign _47508_ = ~D[3] /*18013*/;
assign _47505_ = _46979_ & _47508_ /*18009*/;
assign _47506_ = _46979_ ^ _47508_ /*18012*/;
assign _47507_ = _47499_ & _47506_ /*18010*/;
assign _47428_ = _47499_ ^ _47506_ /*18011*/;
assign _47504_ = _47505_ | _47507_ /*18008*/;
assign _47513_ = ~D[4] /*18007*/;
assign _47510_ = _46980_ & _47513_ /*18003*/;
assign _47511_ = _46980_ ^ _47513_ /*18006*/;
assign _47512_ = _47504_ & _47511_ /*18004*/;
assign _47429_ = _47504_ ^ _47511_ /*18005*/;
assign _47509_ = _47510_ | _47512_ /*18002*/;
assign _47518_ = ~D[5] /*18001*/;
assign _47515_ = _46981_ & _47518_ /*17997*/;
assign _47516_ = _46981_ ^ _47518_ /*18000*/;
assign _47517_ = _47509_ & _47516_ /*17998*/;
assign _47430_ = _47509_ ^ _47516_ /*17999*/;
assign _47514_ = _47515_ | _47517_ /*17996*/;
assign _47523_ = ~D[6] /*17995*/;
assign _47520_ = _46982_ & _47523_ /*17991*/;
assign _47521_ = _46982_ ^ _47523_ /*17994*/;
assign _47522_ = _47514_ & _47521_ /*17992*/;
assign _47431_ = _47514_ ^ _47521_ /*17993*/;
assign _47519_ = _47520_ | _47522_ /*17990*/;
assign _47528_ = ~D[7] /*17989*/;
assign _47525_ = _46983_ & _47528_ /*17985*/;
assign _47526_ = _46983_ ^ _47528_ /*17988*/;
assign _47527_ = _47519_ & _47526_ /*17986*/;
assign _47432_ = _47519_ ^ _47526_ /*17987*/;
assign _47524_ = _47525_ | _47527_ /*17984*/;
assign _47533_ = ~D[8] /*17983*/;
assign _47530_ = _46984_ & _47533_ /*17979*/;
assign _47531_ = _46984_ ^ _47533_ /*17982*/;
assign _47532_ = _47524_ & _47531_ /*17980*/;
assign _47433_ = _47524_ ^ _47531_ /*17981*/;
assign _47529_ = _47530_ | _47532_ /*17978*/;
assign _47538_ = ~D[9] /*17977*/;
assign _47535_ = _46985_ & _47538_ /*17973*/;
assign _47536_ = _46985_ ^ _47538_ /*17976*/;
assign _47537_ = _47529_ & _47536_ /*17974*/;
assign _47434_ = _47529_ ^ _47536_ /*17975*/;
assign _47534_ = _47535_ | _47537_ /*17972*/;
assign _47543_ = ~D[10] /*17971*/;
assign _47540_ = _46986_ & _47543_ /*17967*/;
assign _47541_ = _46986_ ^ _47543_ /*17970*/;
assign _47542_ = _47534_ & _47541_ /*17968*/;
assign _47435_ = _47534_ ^ _47541_ /*17969*/;
assign _47539_ = _47540_ | _47542_ /*17966*/;
assign _47548_ = ~D[11] /*17965*/;
assign _47545_ = _46987_ & _47548_ /*17961*/;
assign _47546_ = _46987_ ^ _47548_ /*17964*/;
assign _47547_ = _47539_ & _47546_ /*17962*/;
assign _47436_ = _47539_ ^ _47546_ /*17963*/;
assign _47544_ = _47545_ | _47547_ /*17960*/;
assign _47553_ = ~D[12] /*17959*/;
assign _47550_ = _46988_ & _47553_ /*17955*/;
assign _47551_ = _46988_ ^ _47553_ /*17958*/;
assign _47552_ = _47544_ & _47551_ /*17956*/;
assign _47437_ = _47544_ ^ _47551_ /*17957*/;
assign _47549_ = _47550_ | _47552_ /*17954*/;
assign _47558_ = ~D[13] /*17953*/;
assign _47555_ = _46989_ & _47558_ /*17949*/;
assign _47556_ = _46989_ ^ _47558_ /*17952*/;
assign _47557_ = _47549_ & _47556_ /*17950*/;
assign _47438_ = _47549_ ^ _47556_ /*17951*/;
assign _47554_ = _47555_ | _47557_ /*17948*/;
assign _47563_ = ~D[14] /*17947*/;
assign _47560_ = _46990_ & _47563_ /*17943*/;
assign _47561_ = _46990_ ^ _47563_ /*17946*/;
assign _47562_ = _47554_ & _47561_ /*17944*/;
assign _47439_ = _47554_ ^ _47561_ /*17945*/;
assign _47559_ = _47560_ | _47562_ /*17942*/;
assign _47568_ = ~D[15] /*17941*/;
assign _47565_ = _46991_ & _47568_ /*17937*/;
assign _47566_ = _46991_ ^ _47568_ /*17940*/;
assign _47567_ = _47559_ & _47566_ /*17938*/;
assign _47440_ = _47559_ ^ _47566_ /*17939*/;
assign _47564_ = _47565_ | _47567_ /*17936*/;
assign _47573_ = ~D[16] /*17935*/;
assign _47570_ = _46992_ & _47573_ /*17931*/;
assign _47571_ = _46992_ ^ _47573_ /*17934*/;
assign _47572_ = _47564_ & _47571_ /*17932*/;
assign _47441_ = _47564_ ^ _47571_ /*17933*/;
assign _47569_ = _47570_ | _47572_ /*17930*/;
assign _47578_ = ~D[17] /*17929*/;
assign _47575_ = _46993_ & _47578_ /*17925*/;
assign _47576_ = _46993_ ^ _47578_ /*17928*/;
assign _47577_ = _47569_ & _47576_ /*17926*/;
assign _47442_ = _47569_ ^ _47576_ /*17927*/;
assign _47574_ = _47575_ | _47577_ /*17924*/;
assign _47583_ = ~D[18] /*17923*/;
assign _47580_ = _46994_ & _47583_ /*17919*/;
assign _47581_ = _46994_ ^ _47583_ /*17922*/;
assign _47582_ = _47574_ & _47581_ /*17920*/;
assign _47443_ = _47574_ ^ _47581_ /*17921*/;
assign _47579_ = _47580_ | _47582_ /*17918*/;
assign _47588_ = ~D[19] /*17917*/;
assign _47585_ = _46995_ & _47588_ /*17913*/;
assign _47586_ = _46995_ ^ _47588_ /*17916*/;
assign _47587_ = _47579_ & _47586_ /*17914*/;
assign _47444_ = _47579_ ^ _47586_ /*17915*/;
assign _47584_ = _47585_ | _47587_ /*17912*/;
assign _47593_ = ~D[20] /*17911*/;
assign _47590_ = _46996_ & _47593_ /*17907*/;
assign _47591_ = _46996_ ^ _47593_ /*17910*/;
assign _47592_ = _47584_ & _47591_ /*17908*/;
assign _47445_ = _47584_ ^ _47591_ /*17909*/;
assign _47589_ = _47590_ | _47592_ /*17906*/;
assign _47598_ = ~D[21] /*17905*/;
assign _47595_ = _46997_ & _47598_ /*17901*/;
assign _47596_ = _46997_ ^ _47598_ /*17904*/;
assign _47597_ = _47589_ & _47596_ /*17902*/;
assign _47446_ = _47589_ ^ _47596_ /*17903*/;
assign _47594_ = _47595_ | _47597_ /*17900*/;
assign _47603_ = ~D[22] /*17899*/;
assign _47600_ = _46998_ & _47603_ /*17895*/;
assign _47601_ = _46998_ ^ _47603_ /*17898*/;
assign _47602_ = _47594_ & _47601_ /*17896*/;
assign _47447_ = _47594_ ^ _47601_ /*17897*/;
assign _47599_ = _47600_ | _47602_ /*17894*/;
assign _47608_ = ~D[23] /*17893*/;
assign _47605_ = _46999_ & _47608_ /*17889*/;
assign _47606_ = _46999_ ^ _47608_ /*17892*/;
assign _47607_ = _47599_ & _47606_ /*17890*/;
assign _47448_ = _47599_ ^ _47606_ /*17891*/;
assign _47604_ = _47605_ | _47607_ /*17888*/;
assign _47613_ = ~D[24] /*17887*/;
assign _47610_ = _47000_ & _47613_ /*17883*/;
assign _47611_ = _47000_ ^ _47613_ /*17886*/;
assign _47612_ = _47604_ & _47611_ /*17884*/;
assign _47449_ = _47604_ ^ _47611_ /*17885*/;
assign _47609_ = _47610_ | _47612_ /*17882*/;
assign _47618_ = ~D[25] /*17881*/;
assign _47615_ = _47001_ & _47618_ /*17877*/;
assign _47616_ = _47001_ ^ _47618_ /*17880*/;
assign _47617_ = _47609_ & _47616_ /*17878*/;
assign _47450_ = _47609_ ^ _47616_ /*17879*/;
assign _47614_ = _47615_ | _47617_ /*17876*/;
assign _47623_ = ~D[26] /*17875*/;
assign _47620_ = _47002_ & _47623_ /*17871*/;
assign _47621_ = _47002_ ^ _47623_ /*17874*/;
assign _47622_ = _47614_ & _47621_ /*17872*/;
assign _47451_ = _47614_ ^ _47621_ /*17873*/;
assign _47619_ = _47620_ | _47622_ /*17870*/;
assign _47628_ = ~D[27] /*17869*/;
assign _47625_ = _47003_ & _47628_ /*17865*/;
assign _47626_ = _47003_ ^ _47628_ /*17868*/;
assign _47627_ = _47619_ & _47626_ /*17866*/;
assign _47452_ = _47619_ ^ _47626_ /*17867*/;
assign _47624_ = _47625_ | _47627_ /*17864*/;
assign _47633_ = ~D[28] /*17863*/;
assign _47630_ = _47004_ & _47633_ /*17859*/;
assign _47631_ = _47004_ ^ _47633_ /*17862*/;
assign _47632_ = _47624_ & _47631_ /*17860*/;
assign _47453_ = _47624_ ^ _47631_ /*17861*/;
assign _47629_ = _47630_ | _47632_ /*17858*/;
assign _47638_ = ~D[29] /*17857*/;
assign _47635_ = _47005_ & _47638_ /*17853*/;
assign _47636_ = _47005_ ^ _47638_ /*17856*/;
assign _47637_ = _47629_ & _47636_ /*17854*/;
assign _47454_ = _47629_ ^ _47636_ /*17855*/;
assign _47634_ = _47635_ | _47637_ /*17852*/;
assign _47643_ = ~D[30] /*17851*/;
assign _47640_ = _47006_ & _47643_ /*17847*/;
assign _47641_ = _47006_ ^ _47643_ /*17850*/;
assign _47642_ = _47634_ & _47641_ /*17848*/;
assign _47455_ = _47634_ ^ _47641_ /*17849*/;
assign _47639_ = _47640_ | _47642_ /*17846*/;
assign _47648_ = ~D[31] /*17845*/;
assign _47645_ = _47007_ & _47648_ /*17841*/;
assign _47646_ = _47007_ ^ _47648_ /*17844*/;
assign _47647_ = _47639_ & _47646_ /*17842*/;
assign _47456_ = _47639_ ^ _47646_ /*17843*/;
assign _47644_ = _47645_ | _47647_ /*17840*/;
assign _47653_ = ~D[32] /*17839*/;
assign _47650_ = _47008_ & _47653_ /*17835*/;
assign _47651_ = _47008_ ^ _47653_ /*17838*/;
assign _47652_ = _47644_ & _47651_ /*17836*/;
assign _47457_ = _47644_ ^ _47651_ /*17837*/;
assign _47649_ = _47650_ | _47652_ /*17834*/;
assign _47658_ = ~D[33] /*17833*/;
assign _47655_ = _47009_ & _47658_ /*17829*/;
assign _47656_ = _47009_ ^ _47658_ /*17832*/;
assign _47657_ = _47649_ & _47656_ /*17830*/;
assign _47458_ = _47649_ ^ _47656_ /*17831*/;
assign _47654_ = _47655_ | _47657_ /*17828*/;
assign _47663_ = ~D[34] /*17827*/;
assign _47660_ = _47010_ & _47663_ /*17823*/;
assign _47661_ = _47010_ ^ _47663_ /*17826*/;
assign _47662_ = _47654_ & _47661_ /*17824*/;
assign _47459_ = _47654_ ^ _47661_ /*17825*/;
assign _47659_ = _47660_ | _47662_ /*17822*/;
assign _47668_ = ~D[35] /*17821*/;
assign _47665_ = _47011_ & _47668_ /*17817*/;
assign _47666_ = _47011_ ^ _47668_ /*17820*/;
assign _47667_ = _47659_ & _47666_ /*17818*/;
assign _47460_ = _47659_ ^ _47666_ /*17819*/;
assign _47664_ = _47665_ | _47667_ /*17816*/;
assign _47673_ = ~D[36] /*17815*/;
assign _47670_ = _47012_ & _47673_ /*17811*/;
assign _47671_ = _47012_ ^ _47673_ /*17814*/;
assign _47672_ = _47664_ & _47671_ /*17812*/;
assign _47461_ = _47664_ ^ _47671_ /*17813*/;
assign _47669_ = _47670_ | _47672_ /*17810*/;
assign _47678_ = ~D[37] /*17809*/;
assign _47675_ = _47013_ & _47678_ /*17805*/;
assign _47676_ = _47013_ ^ _47678_ /*17808*/;
assign _47677_ = _47669_ & _47676_ /*17806*/;
assign _47462_ = _47669_ ^ _47676_ /*17807*/;
assign _47674_ = _47675_ | _47677_ /*17804*/;
assign _47683_ = ~D[38] /*17803*/;
assign _47680_ = _47014_ & _47683_ /*17799*/;
assign _47681_ = _47014_ ^ _47683_ /*17802*/;
assign _47682_ = _47674_ & _47681_ /*17800*/;
assign _47463_ = _47674_ ^ _47681_ /*17801*/;
assign _47679_ = _47680_ | _47682_ /*17798*/;
assign _47688_ = ~D[39] /*17797*/;
assign _47685_ = _47015_ & _47688_ /*17793*/;
assign _47686_ = _47015_ ^ _47688_ /*17796*/;
assign _47687_ = _47679_ & _47686_ /*17794*/;
assign _47464_ = _47679_ ^ _47686_ /*17795*/;
assign _47684_ = _47685_ | _47687_ /*17792*/;
assign _47693_ = ~D[40] /*17791*/;
assign _47690_ = _47016_ & _47693_ /*17787*/;
assign _47691_ = _47016_ ^ _47693_ /*17790*/;
assign _47692_ = _47684_ & _47691_ /*17788*/;
assign _47465_ = _47684_ ^ _47691_ /*17789*/;
assign _47689_ = _47690_ | _47692_ /*17786*/;
assign _47698_ = ~D[41] /*17785*/;
assign _47695_ = _47017_ & _47698_ /*17781*/;
assign _47696_ = _47017_ ^ _47698_ /*17784*/;
assign _47697_ = _47689_ & _47696_ /*17782*/;
assign _47466_ = _47689_ ^ _47696_ /*17783*/;
assign _47694_ = _47695_ | _47697_ /*17780*/;
assign _47703_ = ~D[42] /*17779*/;
assign _47700_ = _47018_ & _47703_ /*17775*/;
assign _47701_ = _47018_ ^ _47703_ /*17778*/;
assign _47702_ = _47694_ & _47701_ /*17776*/;
assign _47467_ = _47694_ ^ _47701_ /*17777*/;
assign _47699_ = _47700_ | _47702_ /*17774*/;
assign _47708_ = ~D[43] /*17773*/;
assign _47705_ = _47019_ & _47708_ /*17769*/;
assign _47706_ = _47019_ ^ _47708_ /*17772*/;
assign _47707_ = _47699_ & _47706_ /*17770*/;
assign _47468_ = _47699_ ^ _47706_ /*17771*/;
assign _47704_ = _47705_ | _47707_ /*17768*/;
assign _47713_ = ~D[44] /*17767*/;
assign _47710_ = _47020_ & _47713_ /*17763*/;
assign _47711_ = _47020_ ^ _47713_ /*17766*/;
assign _47712_ = _47704_ & _47711_ /*17764*/;
assign _47469_ = _47704_ ^ _47711_ /*17765*/;
assign _47709_ = _47710_ | _47712_ /*17762*/;
assign _47718_ = ~D[45] /*17761*/;
assign _47715_ = _47021_ & _47718_ /*17757*/;
assign _47716_ = _47021_ ^ _47718_ /*17760*/;
assign _47717_ = _47709_ & _47716_ /*17758*/;
assign _47470_ = _47709_ ^ _47716_ /*17759*/;
assign _47714_ = _47715_ | _47717_ /*17756*/;
assign _47723_ = ~D[46] /*17755*/;
assign _47720_ = _47022_ & _47723_ /*17751*/;
assign _47721_ = _47022_ ^ _47723_ /*17754*/;
assign _47722_ = _47714_ & _47721_ /*17752*/;
assign _47471_ = _47714_ ^ _47721_ /*17753*/;
assign _47719_ = _47720_ | _47722_ /*17750*/;
assign _47728_ = ~D[47] /*17749*/;
assign _47725_ = _47023_ & _47728_ /*17745*/;
assign _47726_ = _47023_ ^ _47728_ /*17748*/;
assign _47727_ = _47719_ & _47726_ /*17746*/;
assign _47472_ = _47719_ ^ _47726_ /*17747*/;
assign _47724_ = _47725_ | _47727_ /*17744*/;
assign _47733_ = ~D[48] /*17743*/;
assign _47730_ = _47024_ & _47733_ /*17739*/;
assign _47731_ = _47024_ ^ _47733_ /*17742*/;
assign _47732_ = _47724_ & _47731_ /*17740*/;
assign _47473_ = _47724_ ^ _47731_ /*17741*/;
assign _47729_ = _47730_ | _47732_ /*17738*/;
assign _47738_ = ~D[49] /*17737*/;
assign _47735_ = _47025_ & _47738_ /*17733*/;
assign _47736_ = _47025_ ^ _47738_ /*17736*/;
assign _47737_ = _47729_ & _47736_ /*17734*/;
assign _47474_ = _47729_ ^ _47736_ /*17735*/;
assign _47734_ = _47735_ | _47737_ /*17732*/;
assign _47743_ = ~D[50] /*17731*/;
assign _47740_ = _47026_ & _47743_ /*17727*/;
assign _47741_ = _47026_ ^ _47743_ /*17730*/;
assign _47742_ = _47734_ & _47741_ /*17728*/;
assign _47475_ = _47734_ ^ _47741_ /*17729*/;
assign _47739_ = _47740_ | _47742_ /*17726*/;
assign _47748_ = ~D[51] /*17725*/;
assign _47745_ = _47027_ & _47748_ /*17721*/;
assign _47746_ = _47027_ ^ _47748_ /*17724*/;
assign _47747_ = _47739_ & _47746_ /*17722*/;
assign _47476_ = _47739_ ^ _47746_ /*17723*/;
assign _47744_ = _47745_ | _47747_ /*17720*/;
assign _47753_ = ~D[52] /*17719*/;
assign _47750_ = _47028_ & _47753_ /*17715*/;
assign _47751_ = _47028_ ^ _47753_ /*17718*/;
assign _47752_ = _47744_ & _47751_ /*17716*/;
assign _47477_ = _47744_ ^ _47751_ /*17717*/;
assign _47749_ = _47750_ | _47752_ /*17714*/;
assign _47758_ = ~D[53] /*17713*/;
assign _47755_ = _47029_ & _47758_ /*17709*/;
assign _47756_ = _47029_ ^ _47758_ /*17712*/;
assign _47757_ = _47749_ & _47756_ /*17710*/;
assign _47478_ = _47749_ ^ _47756_ /*17711*/;
assign _47754_ = _47755_ | _47757_ /*17708*/;
assign _47763_ = ~D[54] /*17707*/;
assign _47760_ = _47030_ & _47763_ /*17703*/;
assign _47761_ = _47030_ ^ _47763_ /*17706*/;
assign _47762_ = _47754_ & _47761_ /*17704*/;
assign _47479_ = _47754_ ^ _47761_ /*17705*/;
assign _47759_ = _47760_ | _47762_ /*17702*/;
assign _47768_ = ~D[55] /*17701*/;
assign _47765_ = _47031_ & _47768_ /*17697*/;
assign _47766_ = _47031_ ^ _47768_ /*17700*/;
assign _47767_ = _47759_ & _47766_ /*17698*/;
assign _47480_ = _47759_ ^ _47766_ /*17699*/;
assign _47764_ = _47765_ | _47767_ /*17696*/;
assign _47773_ = ~D[56] /*17695*/;
assign _47770_ = _47032_ & _47773_ /*17691*/;
assign _47771_ = _47032_ ^ _47773_ /*17694*/;
assign _47772_ = _47764_ & _47771_ /*17692*/;
assign _47481_ = _47764_ ^ _47771_ /*17693*/;
assign _47769_ = _47770_ | _47772_ /*17690*/;
assign _47778_ = ~D[57] /*17689*/;
assign _47775_ = _47033_ & _47778_ /*17685*/;
assign _47776_ = _47033_ ^ _47778_ /*17688*/;
assign _47777_ = _47769_ & _47776_ /*17686*/;
assign _47482_ = _47769_ ^ _47776_ /*17687*/;
assign _47774_ = _47775_ | _47777_ /*17684*/;
assign _47783_ = ~D[58] /*17683*/;
assign _47780_ = _47034_ & _47783_ /*17679*/;
assign _47781_ = _47034_ ^ _47783_ /*17682*/;
assign _47782_ = _47774_ & _47781_ /*17680*/;
assign _47483_ = _47774_ ^ _47781_ /*17681*/;
assign _47779_ = _47780_ | _47782_ /*17678*/;
assign _47788_ = ~D[59] /*17677*/;
assign _47785_ = _47035_ & _47788_ /*17673*/;
assign _47786_ = _47035_ ^ _47788_ /*17676*/;
assign _47787_ = _47779_ & _47786_ /*17674*/;
assign _47484_ = _47779_ ^ _47786_ /*17675*/;
assign _47784_ = _47785_ | _47787_ /*17672*/;
assign _47793_ = ~D[60] /*17671*/;
assign _47790_ = _47036_ & _47793_ /*17667*/;
assign _47791_ = _47036_ ^ _47793_ /*17670*/;
assign _47792_ = _47784_ & _47791_ /*17668*/;
assign _47485_ = _47784_ ^ _47791_ /*17669*/;
assign _47789_ = _47790_ | _47792_ /*17666*/;
assign _47798_ = ~D[61] /*17665*/;
assign _47795_ = _47037_ & _47798_ /*17661*/;
assign _47796_ = _47037_ ^ _47798_ /*17664*/;
assign _47797_ = _47789_ & _47796_ /*17662*/;
assign _47486_ = _47789_ ^ _47796_ /*17663*/;
assign _47794_ = _47795_ | _47797_ /*17660*/;
assign _47803_ = ~D[62] /*17659*/;
assign _47800_ = _47038_ & _47803_ /*17655*/;
assign _47801_ = _47038_ ^ _47803_ /*17658*/;
assign _47802_ = _47794_ & _47801_ /*17656*/;
assign _47487_ = _47794_ ^ _47801_ /*17657*/;
assign _47799_ = _47800_ | _47802_ /*17654*/;
assign _47804_ = _47039_ & oneWire /*17649*/;
assign _47805_ = _47039_ ^ oneWire /*17652*/;
assign _47806_ = _47799_ & _47805_ /*17650*/;
assign _47488_ = _47799_ ^ _47805_ /*17651*/;
assign Q[10] = _47804_ | _47806_ /*17648*/;
assign _47939_ = ~Q[10] /*17263*/;
assign _47938_ = _47939_ & D[0] /*17262*/;
assign _47941_ = _47425_ & _47938_ /*17257*/;
assign _47942_ = _47425_ ^ _47938_ /*17260*/;
assign _47943_ = zeroWire & _47942_ /*17258*/;
assign _47873_ = zeroWire ^ _47942_ /*17259*/;
assign _47940_ = _47941_ | _47943_ /*17256*/;
assign _47945_ = ~Q[10] /*17255*/;
assign _47944_ = _47945_ & D[1] /*17254*/;
assign _47947_ = _47426_ & _47944_ /*17249*/;
assign _47948_ = _47426_ ^ _47944_ /*17252*/;
assign _47949_ = _47940_ & _47948_ /*17250*/;
assign _47874_ = _47940_ ^ _47948_ /*17251*/;
assign _47946_ = _47947_ | _47949_ /*17248*/;
assign _47951_ = ~Q[10] /*17247*/;
assign _47950_ = _47951_ & D[2] /*17246*/;
assign _47953_ = _47427_ & _47950_ /*17241*/;
assign _47954_ = _47427_ ^ _47950_ /*17244*/;
assign _47955_ = _47946_ & _47954_ /*17242*/;
assign _47875_ = _47946_ ^ _47954_ /*17243*/;
assign _47952_ = _47953_ | _47955_ /*17240*/;
assign _47957_ = ~Q[10] /*17239*/;
assign _47956_ = _47957_ & D[3] /*17238*/;
assign _47959_ = _47428_ & _47956_ /*17233*/;
assign _47960_ = _47428_ ^ _47956_ /*17236*/;
assign _47961_ = _47952_ & _47960_ /*17234*/;
assign _47876_ = _47952_ ^ _47960_ /*17235*/;
assign _47958_ = _47959_ | _47961_ /*17232*/;
assign _47963_ = ~Q[10] /*17231*/;
assign _47962_ = _47963_ & D[4] /*17230*/;
assign _47965_ = _47429_ & _47962_ /*17225*/;
assign _47966_ = _47429_ ^ _47962_ /*17228*/;
assign _47967_ = _47958_ & _47966_ /*17226*/;
assign _47877_ = _47958_ ^ _47966_ /*17227*/;
assign _47964_ = _47965_ | _47967_ /*17224*/;
assign _47969_ = ~Q[10] /*17223*/;
assign _47968_ = _47969_ & D[5] /*17222*/;
assign _47971_ = _47430_ & _47968_ /*17217*/;
assign _47972_ = _47430_ ^ _47968_ /*17220*/;
assign _47973_ = _47964_ & _47972_ /*17218*/;
assign _47878_ = _47964_ ^ _47972_ /*17219*/;
assign _47970_ = _47971_ | _47973_ /*17216*/;
assign _47975_ = ~Q[10] /*17215*/;
assign _47974_ = _47975_ & D[6] /*17214*/;
assign _47977_ = _47431_ & _47974_ /*17209*/;
assign _47978_ = _47431_ ^ _47974_ /*17212*/;
assign _47979_ = _47970_ & _47978_ /*17210*/;
assign _47879_ = _47970_ ^ _47978_ /*17211*/;
assign _47976_ = _47977_ | _47979_ /*17208*/;
assign _47981_ = ~Q[10] /*17207*/;
assign _47980_ = _47981_ & D[7] /*17206*/;
assign _47983_ = _47432_ & _47980_ /*17201*/;
assign _47984_ = _47432_ ^ _47980_ /*17204*/;
assign _47985_ = _47976_ & _47984_ /*17202*/;
assign _47880_ = _47976_ ^ _47984_ /*17203*/;
assign _47982_ = _47983_ | _47985_ /*17200*/;
assign _47987_ = ~Q[10] /*17199*/;
assign _47986_ = _47987_ & D[8] /*17198*/;
assign _47989_ = _47433_ & _47986_ /*17193*/;
assign _47990_ = _47433_ ^ _47986_ /*17196*/;
assign _47991_ = _47982_ & _47990_ /*17194*/;
assign _47881_ = _47982_ ^ _47990_ /*17195*/;
assign _47988_ = _47989_ | _47991_ /*17192*/;
assign _47993_ = ~Q[10] /*17191*/;
assign _47992_ = _47993_ & D[9] /*17190*/;
assign _47995_ = _47434_ & _47992_ /*17185*/;
assign _47996_ = _47434_ ^ _47992_ /*17188*/;
assign _47997_ = _47988_ & _47996_ /*17186*/;
assign _47882_ = _47988_ ^ _47996_ /*17187*/;
assign _47994_ = _47995_ | _47997_ /*17184*/;
assign _47999_ = ~Q[10] /*17183*/;
assign _47998_ = _47999_ & D[10] /*17182*/;
assign _48001_ = _47435_ & _47998_ /*17177*/;
assign _48002_ = _47435_ ^ _47998_ /*17180*/;
assign _48003_ = _47994_ & _48002_ /*17178*/;
assign _47883_ = _47994_ ^ _48002_ /*17179*/;
assign _48000_ = _48001_ | _48003_ /*17176*/;
assign _48005_ = ~Q[10] /*17175*/;
assign _48004_ = _48005_ & D[11] /*17174*/;
assign _48007_ = _47436_ & _48004_ /*17169*/;
assign _48008_ = _47436_ ^ _48004_ /*17172*/;
assign _48009_ = _48000_ & _48008_ /*17170*/;
assign _47884_ = _48000_ ^ _48008_ /*17171*/;
assign _48006_ = _48007_ | _48009_ /*17168*/;
assign _48011_ = ~Q[10] /*17167*/;
assign _48010_ = _48011_ & D[12] /*17166*/;
assign _48013_ = _47437_ & _48010_ /*17161*/;
assign _48014_ = _47437_ ^ _48010_ /*17164*/;
assign _48015_ = _48006_ & _48014_ /*17162*/;
assign _47885_ = _48006_ ^ _48014_ /*17163*/;
assign _48012_ = _48013_ | _48015_ /*17160*/;
assign _48017_ = ~Q[10] /*17159*/;
assign _48016_ = _48017_ & D[13] /*17158*/;
assign _48019_ = _47438_ & _48016_ /*17153*/;
assign _48020_ = _47438_ ^ _48016_ /*17156*/;
assign _48021_ = _48012_ & _48020_ /*17154*/;
assign _47886_ = _48012_ ^ _48020_ /*17155*/;
assign _48018_ = _48019_ | _48021_ /*17152*/;
assign _48023_ = ~Q[10] /*17151*/;
assign _48022_ = _48023_ & D[14] /*17150*/;
assign _48025_ = _47439_ & _48022_ /*17145*/;
assign _48026_ = _47439_ ^ _48022_ /*17148*/;
assign _48027_ = _48018_ & _48026_ /*17146*/;
assign _47887_ = _48018_ ^ _48026_ /*17147*/;
assign _48024_ = _48025_ | _48027_ /*17144*/;
assign _48029_ = ~Q[10] /*17143*/;
assign _48028_ = _48029_ & D[15] /*17142*/;
assign _48031_ = _47440_ & _48028_ /*17137*/;
assign _48032_ = _47440_ ^ _48028_ /*17140*/;
assign _48033_ = _48024_ & _48032_ /*17138*/;
assign _47888_ = _48024_ ^ _48032_ /*17139*/;
assign _48030_ = _48031_ | _48033_ /*17136*/;
assign _48035_ = ~Q[10] /*17135*/;
assign _48034_ = _48035_ & D[16] /*17134*/;
assign _48037_ = _47441_ & _48034_ /*17129*/;
assign _48038_ = _47441_ ^ _48034_ /*17132*/;
assign _48039_ = _48030_ & _48038_ /*17130*/;
assign _47889_ = _48030_ ^ _48038_ /*17131*/;
assign _48036_ = _48037_ | _48039_ /*17128*/;
assign _48041_ = ~Q[10] /*17127*/;
assign _48040_ = _48041_ & D[17] /*17126*/;
assign _48043_ = _47442_ & _48040_ /*17121*/;
assign _48044_ = _47442_ ^ _48040_ /*17124*/;
assign _48045_ = _48036_ & _48044_ /*17122*/;
assign _47890_ = _48036_ ^ _48044_ /*17123*/;
assign _48042_ = _48043_ | _48045_ /*17120*/;
assign _48047_ = ~Q[10] /*17119*/;
assign _48046_ = _48047_ & D[18] /*17118*/;
assign _48049_ = _47443_ & _48046_ /*17113*/;
assign _48050_ = _47443_ ^ _48046_ /*17116*/;
assign _48051_ = _48042_ & _48050_ /*17114*/;
assign _47891_ = _48042_ ^ _48050_ /*17115*/;
assign _48048_ = _48049_ | _48051_ /*17112*/;
assign _48053_ = ~Q[10] /*17111*/;
assign _48052_ = _48053_ & D[19] /*17110*/;
assign _48055_ = _47444_ & _48052_ /*17105*/;
assign _48056_ = _47444_ ^ _48052_ /*17108*/;
assign _48057_ = _48048_ & _48056_ /*17106*/;
assign _47892_ = _48048_ ^ _48056_ /*17107*/;
assign _48054_ = _48055_ | _48057_ /*17104*/;
assign _48059_ = ~Q[10] /*17103*/;
assign _48058_ = _48059_ & D[20] /*17102*/;
assign _48061_ = _47445_ & _48058_ /*17097*/;
assign _48062_ = _47445_ ^ _48058_ /*17100*/;
assign _48063_ = _48054_ & _48062_ /*17098*/;
assign _47893_ = _48054_ ^ _48062_ /*17099*/;
assign _48060_ = _48061_ | _48063_ /*17096*/;
assign _48065_ = ~Q[10] /*17095*/;
assign _48064_ = _48065_ & D[21] /*17094*/;
assign _48067_ = _47446_ & _48064_ /*17089*/;
assign _48068_ = _47446_ ^ _48064_ /*17092*/;
assign _48069_ = _48060_ & _48068_ /*17090*/;
assign _47894_ = _48060_ ^ _48068_ /*17091*/;
assign _48066_ = _48067_ | _48069_ /*17088*/;
assign _48071_ = ~Q[10] /*17087*/;
assign _48070_ = _48071_ & D[22] /*17086*/;
assign _48073_ = _47447_ & _48070_ /*17081*/;
assign _48074_ = _47447_ ^ _48070_ /*17084*/;
assign _48075_ = _48066_ & _48074_ /*17082*/;
assign _47895_ = _48066_ ^ _48074_ /*17083*/;
assign _48072_ = _48073_ | _48075_ /*17080*/;
assign _48077_ = ~Q[10] /*17079*/;
assign _48076_ = _48077_ & D[23] /*17078*/;
assign _48079_ = _47448_ & _48076_ /*17073*/;
assign _48080_ = _47448_ ^ _48076_ /*17076*/;
assign _48081_ = _48072_ & _48080_ /*17074*/;
assign _47896_ = _48072_ ^ _48080_ /*17075*/;
assign _48078_ = _48079_ | _48081_ /*17072*/;
assign _48083_ = ~Q[10] /*17071*/;
assign _48082_ = _48083_ & D[24] /*17070*/;
assign _48085_ = _47449_ & _48082_ /*17065*/;
assign _48086_ = _47449_ ^ _48082_ /*17068*/;
assign _48087_ = _48078_ & _48086_ /*17066*/;
assign _47897_ = _48078_ ^ _48086_ /*17067*/;
assign _48084_ = _48085_ | _48087_ /*17064*/;
assign _48089_ = ~Q[10] /*17063*/;
assign _48088_ = _48089_ & D[25] /*17062*/;
assign _48091_ = _47450_ & _48088_ /*17057*/;
assign _48092_ = _47450_ ^ _48088_ /*17060*/;
assign _48093_ = _48084_ & _48092_ /*17058*/;
assign _47898_ = _48084_ ^ _48092_ /*17059*/;
assign _48090_ = _48091_ | _48093_ /*17056*/;
assign _48095_ = ~Q[10] /*17055*/;
assign _48094_ = _48095_ & D[26] /*17054*/;
assign _48097_ = _47451_ & _48094_ /*17049*/;
assign _48098_ = _47451_ ^ _48094_ /*17052*/;
assign _48099_ = _48090_ & _48098_ /*17050*/;
assign _47899_ = _48090_ ^ _48098_ /*17051*/;
assign _48096_ = _48097_ | _48099_ /*17048*/;
assign _48101_ = ~Q[10] /*17047*/;
assign _48100_ = _48101_ & D[27] /*17046*/;
assign _48103_ = _47452_ & _48100_ /*17041*/;
assign _48104_ = _47452_ ^ _48100_ /*17044*/;
assign _48105_ = _48096_ & _48104_ /*17042*/;
assign _47900_ = _48096_ ^ _48104_ /*17043*/;
assign _48102_ = _48103_ | _48105_ /*17040*/;
assign _48107_ = ~Q[10] /*17039*/;
assign _48106_ = _48107_ & D[28] /*17038*/;
assign _48109_ = _47453_ & _48106_ /*17033*/;
assign _48110_ = _47453_ ^ _48106_ /*17036*/;
assign _48111_ = _48102_ & _48110_ /*17034*/;
assign _47901_ = _48102_ ^ _48110_ /*17035*/;
assign _48108_ = _48109_ | _48111_ /*17032*/;
assign _48113_ = ~Q[10] /*17031*/;
assign _48112_ = _48113_ & D[29] /*17030*/;
assign _48115_ = _47454_ & _48112_ /*17025*/;
assign _48116_ = _47454_ ^ _48112_ /*17028*/;
assign _48117_ = _48108_ & _48116_ /*17026*/;
assign _47902_ = _48108_ ^ _48116_ /*17027*/;
assign _48114_ = _48115_ | _48117_ /*17024*/;
assign _48119_ = ~Q[10] /*17023*/;
assign _48118_ = _48119_ & D[30] /*17022*/;
assign _48121_ = _47455_ & _48118_ /*17017*/;
assign _48122_ = _47455_ ^ _48118_ /*17020*/;
assign _48123_ = _48114_ & _48122_ /*17018*/;
assign _47903_ = _48114_ ^ _48122_ /*17019*/;
assign _48120_ = _48121_ | _48123_ /*17016*/;
assign _48125_ = ~Q[10] /*17015*/;
assign _48124_ = _48125_ & D[31] /*17014*/;
assign _48127_ = _47456_ & _48124_ /*17009*/;
assign _48128_ = _47456_ ^ _48124_ /*17012*/;
assign _48129_ = _48120_ & _48128_ /*17010*/;
assign _47904_ = _48120_ ^ _48128_ /*17011*/;
assign _48126_ = _48127_ | _48129_ /*17008*/;
assign _48131_ = ~Q[10] /*17007*/;
assign _48130_ = _48131_ & D[32] /*17006*/;
assign _48133_ = _47457_ & _48130_ /*17001*/;
assign _48134_ = _47457_ ^ _48130_ /*17004*/;
assign _48135_ = _48126_ & _48134_ /*17002*/;
assign _47905_ = _48126_ ^ _48134_ /*17003*/;
assign _48132_ = _48133_ | _48135_ /*17000*/;
assign _48137_ = ~Q[10] /*16999*/;
assign _48136_ = _48137_ & D[33] /*16998*/;
assign _48139_ = _47458_ & _48136_ /*16993*/;
assign _48140_ = _47458_ ^ _48136_ /*16996*/;
assign _48141_ = _48132_ & _48140_ /*16994*/;
assign _47906_ = _48132_ ^ _48140_ /*16995*/;
assign _48138_ = _48139_ | _48141_ /*16992*/;
assign _48143_ = ~Q[10] /*16991*/;
assign _48142_ = _48143_ & D[34] /*16990*/;
assign _48145_ = _47459_ & _48142_ /*16985*/;
assign _48146_ = _47459_ ^ _48142_ /*16988*/;
assign _48147_ = _48138_ & _48146_ /*16986*/;
assign _47907_ = _48138_ ^ _48146_ /*16987*/;
assign _48144_ = _48145_ | _48147_ /*16984*/;
assign _48149_ = ~Q[10] /*16983*/;
assign _48148_ = _48149_ & D[35] /*16982*/;
assign _48151_ = _47460_ & _48148_ /*16977*/;
assign _48152_ = _47460_ ^ _48148_ /*16980*/;
assign _48153_ = _48144_ & _48152_ /*16978*/;
assign _47908_ = _48144_ ^ _48152_ /*16979*/;
assign _48150_ = _48151_ | _48153_ /*16976*/;
assign _48155_ = ~Q[10] /*16975*/;
assign _48154_ = _48155_ & D[36] /*16974*/;
assign _48157_ = _47461_ & _48154_ /*16969*/;
assign _48158_ = _47461_ ^ _48154_ /*16972*/;
assign _48159_ = _48150_ & _48158_ /*16970*/;
assign _47909_ = _48150_ ^ _48158_ /*16971*/;
assign _48156_ = _48157_ | _48159_ /*16968*/;
assign _48161_ = ~Q[10] /*16967*/;
assign _48160_ = _48161_ & D[37] /*16966*/;
assign _48163_ = _47462_ & _48160_ /*16961*/;
assign _48164_ = _47462_ ^ _48160_ /*16964*/;
assign _48165_ = _48156_ & _48164_ /*16962*/;
assign _47910_ = _48156_ ^ _48164_ /*16963*/;
assign _48162_ = _48163_ | _48165_ /*16960*/;
assign _48167_ = ~Q[10] /*16959*/;
assign _48166_ = _48167_ & D[38] /*16958*/;
assign _48169_ = _47463_ & _48166_ /*16953*/;
assign _48170_ = _47463_ ^ _48166_ /*16956*/;
assign _48171_ = _48162_ & _48170_ /*16954*/;
assign _47911_ = _48162_ ^ _48170_ /*16955*/;
assign _48168_ = _48169_ | _48171_ /*16952*/;
assign _48173_ = ~Q[10] /*16951*/;
assign _48172_ = _48173_ & D[39] /*16950*/;
assign _48175_ = _47464_ & _48172_ /*16945*/;
assign _48176_ = _47464_ ^ _48172_ /*16948*/;
assign _48177_ = _48168_ & _48176_ /*16946*/;
assign _47912_ = _48168_ ^ _48176_ /*16947*/;
assign _48174_ = _48175_ | _48177_ /*16944*/;
assign _48179_ = ~Q[10] /*16943*/;
assign _48178_ = _48179_ & D[40] /*16942*/;
assign _48181_ = _47465_ & _48178_ /*16937*/;
assign _48182_ = _47465_ ^ _48178_ /*16940*/;
assign _48183_ = _48174_ & _48182_ /*16938*/;
assign _47913_ = _48174_ ^ _48182_ /*16939*/;
assign _48180_ = _48181_ | _48183_ /*16936*/;
assign _48185_ = ~Q[10] /*16935*/;
assign _48184_ = _48185_ & D[41] /*16934*/;
assign _48187_ = _47466_ & _48184_ /*16929*/;
assign _48188_ = _47466_ ^ _48184_ /*16932*/;
assign _48189_ = _48180_ & _48188_ /*16930*/;
assign _47914_ = _48180_ ^ _48188_ /*16931*/;
assign _48186_ = _48187_ | _48189_ /*16928*/;
assign _48191_ = ~Q[10] /*16927*/;
assign _48190_ = _48191_ & D[42] /*16926*/;
assign _48193_ = _47467_ & _48190_ /*16921*/;
assign _48194_ = _47467_ ^ _48190_ /*16924*/;
assign _48195_ = _48186_ & _48194_ /*16922*/;
assign _47915_ = _48186_ ^ _48194_ /*16923*/;
assign _48192_ = _48193_ | _48195_ /*16920*/;
assign _48197_ = ~Q[10] /*16919*/;
assign _48196_ = _48197_ & D[43] /*16918*/;
assign _48199_ = _47468_ & _48196_ /*16913*/;
assign _48200_ = _47468_ ^ _48196_ /*16916*/;
assign _48201_ = _48192_ & _48200_ /*16914*/;
assign _47916_ = _48192_ ^ _48200_ /*16915*/;
assign _48198_ = _48199_ | _48201_ /*16912*/;
assign _48203_ = ~Q[10] /*16911*/;
assign _48202_ = _48203_ & D[44] /*16910*/;
assign _48205_ = _47469_ & _48202_ /*16905*/;
assign _48206_ = _47469_ ^ _48202_ /*16908*/;
assign _48207_ = _48198_ & _48206_ /*16906*/;
assign _47917_ = _48198_ ^ _48206_ /*16907*/;
assign _48204_ = _48205_ | _48207_ /*16904*/;
assign _48209_ = ~Q[10] /*16903*/;
assign _48208_ = _48209_ & D[45] /*16902*/;
assign _48211_ = _47470_ & _48208_ /*16897*/;
assign _48212_ = _47470_ ^ _48208_ /*16900*/;
assign _48213_ = _48204_ & _48212_ /*16898*/;
assign _47918_ = _48204_ ^ _48212_ /*16899*/;
assign _48210_ = _48211_ | _48213_ /*16896*/;
assign _48215_ = ~Q[10] /*16895*/;
assign _48214_ = _48215_ & D[46] /*16894*/;
assign _48217_ = _47471_ & _48214_ /*16889*/;
assign _48218_ = _47471_ ^ _48214_ /*16892*/;
assign _48219_ = _48210_ & _48218_ /*16890*/;
assign _47919_ = _48210_ ^ _48218_ /*16891*/;
assign _48216_ = _48217_ | _48219_ /*16888*/;
assign _48221_ = ~Q[10] /*16887*/;
assign _48220_ = _48221_ & D[47] /*16886*/;
assign _48223_ = _47472_ & _48220_ /*16881*/;
assign _48224_ = _47472_ ^ _48220_ /*16884*/;
assign _48225_ = _48216_ & _48224_ /*16882*/;
assign _47920_ = _48216_ ^ _48224_ /*16883*/;
assign _48222_ = _48223_ | _48225_ /*16880*/;
assign _48227_ = ~Q[10] /*16879*/;
assign _48226_ = _48227_ & D[48] /*16878*/;
assign _48229_ = _47473_ & _48226_ /*16873*/;
assign _48230_ = _47473_ ^ _48226_ /*16876*/;
assign _48231_ = _48222_ & _48230_ /*16874*/;
assign _47921_ = _48222_ ^ _48230_ /*16875*/;
assign _48228_ = _48229_ | _48231_ /*16872*/;
assign _48233_ = ~Q[10] /*16871*/;
assign _48232_ = _48233_ & D[49] /*16870*/;
assign _48235_ = _47474_ & _48232_ /*16865*/;
assign _48236_ = _47474_ ^ _48232_ /*16868*/;
assign _48237_ = _48228_ & _48236_ /*16866*/;
assign _47922_ = _48228_ ^ _48236_ /*16867*/;
assign _48234_ = _48235_ | _48237_ /*16864*/;
assign _48239_ = ~Q[10] /*16863*/;
assign _48238_ = _48239_ & D[50] /*16862*/;
assign _48241_ = _47475_ & _48238_ /*16857*/;
assign _48242_ = _47475_ ^ _48238_ /*16860*/;
assign _48243_ = _48234_ & _48242_ /*16858*/;
assign _47923_ = _48234_ ^ _48242_ /*16859*/;
assign _48240_ = _48241_ | _48243_ /*16856*/;
assign _48245_ = ~Q[10] /*16855*/;
assign _48244_ = _48245_ & D[51] /*16854*/;
assign _48247_ = _47476_ & _48244_ /*16849*/;
assign _48248_ = _47476_ ^ _48244_ /*16852*/;
assign _48249_ = _48240_ & _48248_ /*16850*/;
assign _47924_ = _48240_ ^ _48248_ /*16851*/;
assign _48246_ = _48247_ | _48249_ /*16848*/;
assign _48251_ = ~Q[10] /*16847*/;
assign _48250_ = _48251_ & D[52] /*16846*/;
assign _48253_ = _47477_ & _48250_ /*16841*/;
assign _48254_ = _47477_ ^ _48250_ /*16844*/;
assign _48255_ = _48246_ & _48254_ /*16842*/;
assign _47925_ = _48246_ ^ _48254_ /*16843*/;
assign _48252_ = _48253_ | _48255_ /*16840*/;
assign _48257_ = ~Q[10] /*16839*/;
assign _48256_ = _48257_ & D[53] /*16838*/;
assign _48259_ = _47478_ & _48256_ /*16833*/;
assign _48260_ = _47478_ ^ _48256_ /*16836*/;
assign _48261_ = _48252_ & _48260_ /*16834*/;
assign _47926_ = _48252_ ^ _48260_ /*16835*/;
assign _48258_ = _48259_ | _48261_ /*16832*/;
assign _48263_ = ~Q[10] /*16831*/;
assign _48262_ = _48263_ & D[54] /*16830*/;
assign _48265_ = _47479_ & _48262_ /*16825*/;
assign _48266_ = _47479_ ^ _48262_ /*16828*/;
assign _48267_ = _48258_ & _48266_ /*16826*/;
assign _47927_ = _48258_ ^ _48266_ /*16827*/;
assign _48264_ = _48265_ | _48267_ /*16824*/;
assign _48269_ = ~Q[10] /*16823*/;
assign _48268_ = _48269_ & D[55] /*16822*/;
assign _48271_ = _47480_ & _48268_ /*16817*/;
assign _48272_ = _47480_ ^ _48268_ /*16820*/;
assign _48273_ = _48264_ & _48272_ /*16818*/;
assign _47928_ = _48264_ ^ _48272_ /*16819*/;
assign _48270_ = _48271_ | _48273_ /*16816*/;
assign _48275_ = ~Q[10] /*16815*/;
assign _48274_ = _48275_ & D[56] /*16814*/;
assign _48277_ = _47481_ & _48274_ /*16809*/;
assign _48278_ = _47481_ ^ _48274_ /*16812*/;
assign _48279_ = _48270_ & _48278_ /*16810*/;
assign _47929_ = _48270_ ^ _48278_ /*16811*/;
assign _48276_ = _48277_ | _48279_ /*16808*/;
assign _48281_ = ~Q[10] /*16807*/;
assign _48280_ = _48281_ & D[57] /*16806*/;
assign _48283_ = _47482_ & _48280_ /*16801*/;
assign _48284_ = _47482_ ^ _48280_ /*16804*/;
assign _48285_ = _48276_ & _48284_ /*16802*/;
assign _47930_ = _48276_ ^ _48284_ /*16803*/;
assign _48282_ = _48283_ | _48285_ /*16800*/;
assign _48287_ = ~Q[10] /*16799*/;
assign _48286_ = _48287_ & D[58] /*16798*/;
assign _48289_ = _47483_ & _48286_ /*16793*/;
assign _48290_ = _47483_ ^ _48286_ /*16796*/;
assign _48291_ = _48282_ & _48290_ /*16794*/;
assign _47931_ = _48282_ ^ _48290_ /*16795*/;
assign _48288_ = _48289_ | _48291_ /*16792*/;
assign _48293_ = ~Q[10] /*16791*/;
assign _48292_ = _48293_ & D[59] /*16790*/;
assign _48295_ = _47484_ & _48292_ /*16785*/;
assign _48296_ = _47484_ ^ _48292_ /*16788*/;
assign _48297_ = _48288_ & _48296_ /*16786*/;
assign _47932_ = _48288_ ^ _48296_ /*16787*/;
assign _48294_ = _48295_ | _48297_ /*16784*/;
assign _48299_ = ~Q[10] /*16783*/;
assign _48298_ = _48299_ & D[60] /*16782*/;
assign _48301_ = _47485_ & _48298_ /*16777*/;
assign _48302_ = _47485_ ^ _48298_ /*16780*/;
assign _48303_ = _48294_ & _48302_ /*16778*/;
assign _47933_ = _48294_ ^ _48302_ /*16779*/;
assign _48300_ = _48301_ | _48303_ /*16776*/;
assign _48305_ = ~Q[10] /*16775*/;
assign _48304_ = _48305_ & D[61] /*16774*/;
assign _48307_ = _47486_ & _48304_ /*16769*/;
assign _48308_ = _47486_ ^ _48304_ /*16772*/;
assign _48309_ = _48300_ & _48308_ /*16770*/;
assign _47934_ = _48300_ ^ _48308_ /*16771*/;
assign _48306_ = _48307_ | _48309_ /*16768*/;
assign _48311_ = ~Q[10] /*16767*/;
assign _48310_ = _48311_ & D[62] /*16766*/;
assign _48313_ = _47487_ & _48310_ /*16761*/;
assign _48314_ = _47487_ ^ _48310_ /*16764*/;
assign _48315_ = _48306_ & _48314_ /*16762*/;
assign _47935_ = _48306_ ^ _48314_ /*16763*/;
assign _48312_ = _48313_ | _48315_ /*16760*/;
assign _48317_ = ~Q[10] /*16759*/;
assign _48316_ = _48317_ & zeroWire /*16758*/;
assign _48318_ = _47488_ ^ _48316_ /*16756*/;
assign _47936_ = _48318_ ^ _48312_ /*16755*/;
assign _48389_ = ~D[0] /*16501*/;
assign _48386_ = R_0[9] & _48389_ /*16497*/;
assign _48387_ = R_0[9] ^ _48389_ /*16500*/;
assign _48388_ = oneWire & _48387_ /*16498*/;
assign _48321_ = oneWire ^ _48387_ /*16499*/;
assign _48385_ = _48386_ | _48388_ /*16496*/;
assign _48394_ = ~D[1] /*16495*/;
assign _48391_ = _47873_ & _48394_ /*16491*/;
assign _48392_ = _47873_ ^ _48394_ /*16494*/;
assign _48393_ = _48385_ & _48392_ /*16492*/;
assign _48322_ = _48385_ ^ _48392_ /*16493*/;
assign _48390_ = _48391_ | _48393_ /*16490*/;
assign _48399_ = ~D[2] /*16489*/;
assign _48396_ = _47874_ & _48399_ /*16485*/;
assign _48397_ = _47874_ ^ _48399_ /*16488*/;
assign _48398_ = _48390_ & _48397_ /*16486*/;
assign _48323_ = _48390_ ^ _48397_ /*16487*/;
assign _48395_ = _48396_ | _48398_ /*16484*/;
assign _48404_ = ~D[3] /*16483*/;
assign _48401_ = _47875_ & _48404_ /*16479*/;
assign _48402_ = _47875_ ^ _48404_ /*16482*/;
assign _48403_ = _48395_ & _48402_ /*16480*/;
assign _48324_ = _48395_ ^ _48402_ /*16481*/;
assign _48400_ = _48401_ | _48403_ /*16478*/;
assign _48409_ = ~D[4] /*16477*/;
assign _48406_ = _47876_ & _48409_ /*16473*/;
assign _48407_ = _47876_ ^ _48409_ /*16476*/;
assign _48408_ = _48400_ & _48407_ /*16474*/;
assign _48325_ = _48400_ ^ _48407_ /*16475*/;
assign _48405_ = _48406_ | _48408_ /*16472*/;
assign _48414_ = ~D[5] /*16471*/;
assign _48411_ = _47877_ & _48414_ /*16467*/;
assign _48412_ = _47877_ ^ _48414_ /*16470*/;
assign _48413_ = _48405_ & _48412_ /*16468*/;
assign _48326_ = _48405_ ^ _48412_ /*16469*/;
assign _48410_ = _48411_ | _48413_ /*16466*/;
assign _48419_ = ~D[6] /*16465*/;
assign _48416_ = _47878_ & _48419_ /*16461*/;
assign _48417_ = _47878_ ^ _48419_ /*16464*/;
assign _48418_ = _48410_ & _48417_ /*16462*/;
assign _48327_ = _48410_ ^ _48417_ /*16463*/;
assign _48415_ = _48416_ | _48418_ /*16460*/;
assign _48424_ = ~D[7] /*16459*/;
assign _48421_ = _47879_ & _48424_ /*16455*/;
assign _48422_ = _47879_ ^ _48424_ /*16458*/;
assign _48423_ = _48415_ & _48422_ /*16456*/;
assign _48328_ = _48415_ ^ _48422_ /*16457*/;
assign _48420_ = _48421_ | _48423_ /*16454*/;
assign _48429_ = ~D[8] /*16453*/;
assign _48426_ = _47880_ & _48429_ /*16449*/;
assign _48427_ = _47880_ ^ _48429_ /*16452*/;
assign _48428_ = _48420_ & _48427_ /*16450*/;
assign _48329_ = _48420_ ^ _48427_ /*16451*/;
assign _48425_ = _48426_ | _48428_ /*16448*/;
assign _48434_ = ~D[9] /*16447*/;
assign _48431_ = _47881_ & _48434_ /*16443*/;
assign _48432_ = _47881_ ^ _48434_ /*16446*/;
assign _48433_ = _48425_ & _48432_ /*16444*/;
assign _48330_ = _48425_ ^ _48432_ /*16445*/;
assign _48430_ = _48431_ | _48433_ /*16442*/;
assign _48439_ = ~D[10] /*16441*/;
assign _48436_ = _47882_ & _48439_ /*16437*/;
assign _48437_ = _47882_ ^ _48439_ /*16440*/;
assign _48438_ = _48430_ & _48437_ /*16438*/;
assign _48331_ = _48430_ ^ _48437_ /*16439*/;
assign _48435_ = _48436_ | _48438_ /*16436*/;
assign _48444_ = ~D[11] /*16435*/;
assign _48441_ = _47883_ & _48444_ /*16431*/;
assign _48442_ = _47883_ ^ _48444_ /*16434*/;
assign _48443_ = _48435_ & _48442_ /*16432*/;
assign _48332_ = _48435_ ^ _48442_ /*16433*/;
assign _48440_ = _48441_ | _48443_ /*16430*/;
assign _48449_ = ~D[12] /*16429*/;
assign _48446_ = _47884_ & _48449_ /*16425*/;
assign _48447_ = _47884_ ^ _48449_ /*16428*/;
assign _48448_ = _48440_ & _48447_ /*16426*/;
assign _48333_ = _48440_ ^ _48447_ /*16427*/;
assign _48445_ = _48446_ | _48448_ /*16424*/;
assign _48454_ = ~D[13] /*16423*/;
assign _48451_ = _47885_ & _48454_ /*16419*/;
assign _48452_ = _47885_ ^ _48454_ /*16422*/;
assign _48453_ = _48445_ & _48452_ /*16420*/;
assign _48334_ = _48445_ ^ _48452_ /*16421*/;
assign _48450_ = _48451_ | _48453_ /*16418*/;
assign _48459_ = ~D[14] /*16417*/;
assign _48456_ = _47886_ & _48459_ /*16413*/;
assign _48457_ = _47886_ ^ _48459_ /*16416*/;
assign _48458_ = _48450_ & _48457_ /*16414*/;
assign _48335_ = _48450_ ^ _48457_ /*16415*/;
assign _48455_ = _48456_ | _48458_ /*16412*/;
assign _48464_ = ~D[15] /*16411*/;
assign _48461_ = _47887_ & _48464_ /*16407*/;
assign _48462_ = _47887_ ^ _48464_ /*16410*/;
assign _48463_ = _48455_ & _48462_ /*16408*/;
assign _48336_ = _48455_ ^ _48462_ /*16409*/;
assign _48460_ = _48461_ | _48463_ /*16406*/;
assign _48469_ = ~D[16] /*16405*/;
assign _48466_ = _47888_ & _48469_ /*16401*/;
assign _48467_ = _47888_ ^ _48469_ /*16404*/;
assign _48468_ = _48460_ & _48467_ /*16402*/;
assign _48337_ = _48460_ ^ _48467_ /*16403*/;
assign _48465_ = _48466_ | _48468_ /*16400*/;
assign _48474_ = ~D[17] /*16399*/;
assign _48471_ = _47889_ & _48474_ /*16395*/;
assign _48472_ = _47889_ ^ _48474_ /*16398*/;
assign _48473_ = _48465_ & _48472_ /*16396*/;
assign _48338_ = _48465_ ^ _48472_ /*16397*/;
assign _48470_ = _48471_ | _48473_ /*16394*/;
assign _48479_ = ~D[18] /*16393*/;
assign _48476_ = _47890_ & _48479_ /*16389*/;
assign _48477_ = _47890_ ^ _48479_ /*16392*/;
assign _48478_ = _48470_ & _48477_ /*16390*/;
assign _48339_ = _48470_ ^ _48477_ /*16391*/;
assign _48475_ = _48476_ | _48478_ /*16388*/;
assign _48484_ = ~D[19] /*16387*/;
assign _48481_ = _47891_ & _48484_ /*16383*/;
assign _48482_ = _47891_ ^ _48484_ /*16386*/;
assign _48483_ = _48475_ & _48482_ /*16384*/;
assign _48340_ = _48475_ ^ _48482_ /*16385*/;
assign _48480_ = _48481_ | _48483_ /*16382*/;
assign _48489_ = ~D[20] /*16381*/;
assign _48486_ = _47892_ & _48489_ /*16377*/;
assign _48487_ = _47892_ ^ _48489_ /*16380*/;
assign _48488_ = _48480_ & _48487_ /*16378*/;
assign _48341_ = _48480_ ^ _48487_ /*16379*/;
assign _48485_ = _48486_ | _48488_ /*16376*/;
assign _48494_ = ~D[21] /*16375*/;
assign _48491_ = _47893_ & _48494_ /*16371*/;
assign _48492_ = _47893_ ^ _48494_ /*16374*/;
assign _48493_ = _48485_ & _48492_ /*16372*/;
assign _48342_ = _48485_ ^ _48492_ /*16373*/;
assign _48490_ = _48491_ | _48493_ /*16370*/;
assign _48499_ = ~D[22] /*16369*/;
assign _48496_ = _47894_ & _48499_ /*16365*/;
assign _48497_ = _47894_ ^ _48499_ /*16368*/;
assign _48498_ = _48490_ & _48497_ /*16366*/;
assign _48343_ = _48490_ ^ _48497_ /*16367*/;
assign _48495_ = _48496_ | _48498_ /*16364*/;
assign _48504_ = ~D[23] /*16363*/;
assign _48501_ = _47895_ & _48504_ /*16359*/;
assign _48502_ = _47895_ ^ _48504_ /*16362*/;
assign _48503_ = _48495_ & _48502_ /*16360*/;
assign _48344_ = _48495_ ^ _48502_ /*16361*/;
assign _48500_ = _48501_ | _48503_ /*16358*/;
assign _48509_ = ~D[24] /*16357*/;
assign _48506_ = _47896_ & _48509_ /*16353*/;
assign _48507_ = _47896_ ^ _48509_ /*16356*/;
assign _48508_ = _48500_ & _48507_ /*16354*/;
assign _48345_ = _48500_ ^ _48507_ /*16355*/;
assign _48505_ = _48506_ | _48508_ /*16352*/;
assign _48514_ = ~D[25] /*16351*/;
assign _48511_ = _47897_ & _48514_ /*16347*/;
assign _48512_ = _47897_ ^ _48514_ /*16350*/;
assign _48513_ = _48505_ & _48512_ /*16348*/;
assign _48346_ = _48505_ ^ _48512_ /*16349*/;
assign _48510_ = _48511_ | _48513_ /*16346*/;
assign _48519_ = ~D[26] /*16345*/;
assign _48516_ = _47898_ & _48519_ /*16341*/;
assign _48517_ = _47898_ ^ _48519_ /*16344*/;
assign _48518_ = _48510_ & _48517_ /*16342*/;
assign _48347_ = _48510_ ^ _48517_ /*16343*/;
assign _48515_ = _48516_ | _48518_ /*16340*/;
assign _48524_ = ~D[27] /*16339*/;
assign _48521_ = _47899_ & _48524_ /*16335*/;
assign _48522_ = _47899_ ^ _48524_ /*16338*/;
assign _48523_ = _48515_ & _48522_ /*16336*/;
assign _48348_ = _48515_ ^ _48522_ /*16337*/;
assign _48520_ = _48521_ | _48523_ /*16334*/;
assign _48529_ = ~D[28] /*16333*/;
assign _48526_ = _47900_ & _48529_ /*16329*/;
assign _48527_ = _47900_ ^ _48529_ /*16332*/;
assign _48528_ = _48520_ & _48527_ /*16330*/;
assign _48349_ = _48520_ ^ _48527_ /*16331*/;
assign _48525_ = _48526_ | _48528_ /*16328*/;
assign _48534_ = ~D[29] /*16327*/;
assign _48531_ = _47901_ & _48534_ /*16323*/;
assign _48532_ = _47901_ ^ _48534_ /*16326*/;
assign _48533_ = _48525_ & _48532_ /*16324*/;
assign _48350_ = _48525_ ^ _48532_ /*16325*/;
assign _48530_ = _48531_ | _48533_ /*16322*/;
assign _48539_ = ~D[30] /*16321*/;
assign _48536_ = _47902_ & _48539_ /*16317*/;
assign _48537_ = _47902_ ^ _48539_ /*16320*/;
assign _48538_ = _48530_ & _48537_ /*16318*/;
assign _48351_ = _48530_ ^ _48537_ /*16319*/;
assign _48535_ = _48536_ | _48538_ /*16316*/;
assign _48544_ = ~D[31] /*16315*/;
assign _48541_ = _47903_ & _48544_ /*16311*/;
assign _48542_ = _47903_ ^ _48544_ /*16314*/;
assign _48543_ = _48535_ & _48542_ /*16312*/;
assign _48352_ = _48535_ ^ _48542_ /*16313*/;
assign _48540_ = _48541_ | _48543_ /*16310*/;
assign _48549_ = ~D[32] /*16309*/;
assign _48546_ = _47904_ & _48549_ /*16305*/;
assign _48547_ = _47904_ ^ _48549_ /*16308*/;
assign _48548_ = _48540_ & _48547_ /*16306*/;
assign _48353_ = _48540_ ^ _48547_ /*16307*/;
assign _48545_ = _48546_ | _48548_ /*16304*/;
assign _48554_ = ~D[33] /*16303*/;
assign _48551_ = _47905_ & _48554_ /*16299*/;
assign _48552_ = _47905_ ^ _48554_ /*16302*/;
assign _48553_ = _48545_ & _48552_ /*16300*/;
assign _48354_ = _48545_ ^ _48552_ /*16301*/;
assign _48550_ = _48551_ | _48553_ /*16298*/;
assign _48559_ = ~D[34] /*16297*/;
assign _48556_ = _47906_ & _48559_ /*16293*/;
assign _48557_ = _47906_ ^ _48559_ /*16296*/;
assign _48558_ = _48550_ & _48557_ /*16294*/;
assign _48355_ = _48550_ ^ _48557_ /*16295*/;
assign _48555_ = _48556_ | _48558_ /*16292*/;
assign _48564_ = ~D[35] /*16291*/;
assign _48561_ = _47907_ & _48564_ /*16287*/;
assign _48562_ = _47907_ ^ _48564_ /*16290*/;
assign _48563_ = _48555_ & _48562_ /*16288*/;
assign _48356_ = _48555_ ^ _48562_ /*16289*/;
assign _48560_ = _48561_ | _48563_ /*16286*/;
assign _48569_ = ~D[36] /*16285*/;
assign _48566_ = _47908_ & _48569_ /*16281*/;
assign _48567_ = _47908_ ^ _48569_ /*16284*/;
assign _48568_ = _48560_ & _48567_ /*16282*/;
assign _48357_ = _48560_ ^ _48567_ /*16283*/;
assign _48565_ = _48566_ | _48568_ /*16280*/;
assign _48574_ = ~D[37] /*16279*/;
assign _48571_ = _47909_ & _48574_ /*16275*/;
assign _48572_ = _47909_ ^ _48574_ /*16278*/;
assign _48573_ = _48565_ & _48572_ /*16276*/;
assign _48358_ = _48565_ ^ _48572_ /*16277*/;
assign _48570_ = _48571_ | _48573_ /*16274*/;
assign _48579_ = ~D[38] /*16273*/;
assign _48576_ = _47910_ & _48579_ /*16269*/;
assign _48577_ = _47910_ ^ _48579_ /*16272*/;
assign _48578_ = _48570_ & _48577_ /*16270*/;
assign _48359_ = _48570_ ^ _48577_ /*16271*/;
assign _48575_ = _48576_ | _48578_ /*16268*/;
assign _48584_ = ~D[39] /*16267*/;
assign _48581_ = _47911_ & _48584_ /*16263*/;
assign _48582_ = _47911_ ^ _48584_ /*16266*/;
assign _48583_ = _48575_ & _48582_ /*16264*/;
assign _48360_ = _48575_ ^ _48582_ /*16265*/;
assign _48580_ = _48581_ | _48583_ /*16262*/;
assign _48589_ = ~D[40] /*16261*/;
assign _48586_ = _47912_ & _48589_ /*16257*/;
assign _48587_ = _47912_ ^ _48589_ /*16260*/;
assign _48588_ = _48580_ & _48587_ /*16258*/;
assign _48361_ = _48580_ ^ _48587_ /*16259*/;
assign _48585_ = _48586_ | _48588_ /*16256*/;
assign _48594_ = ~D[41] /*16255*/;
assign _48591_ = _47913_ & _48594_ /*16251*/;
assign _48592_ = _47913_ ^ _48594_ /*16254*/;
assign _48593_ = _48585_ & _48592_ /*16252*/;
assign _48362_ = _48585_ ^ _48592_ /*16253*/;
assign _48590_ = _48591_ | _48593_ /*16250*/;
assign _48599_ = ~D[42] /*16249*/;
assign _48596_ = _47914_ & _48599_ /*16245*/;
assign _48597_ = _47914_ ^ _48599_ /*16248*/;
assign _48598_ = _48590_ & _48597_ /*16246*/;
assign _48363_ = _48590_ ^ _48597_ /*16247*/;
assign _48595_ = _48596_ | _48598_ /*16244*/;
assign _48604_ = ~D[43] /*16243*/;
assign _48601_ = _47915_ & _48604_ /*16239*/;
assign _48602_ = _47915_ ^ _48604_ /*16242*/;
assign _48603_ = _48595_ & _48602_ /*16240*/;
assign _48364_ = _48595_ ^ _48602_ /*16241*/;
assign _48600_ = _48601_ | _48603_ /*16238*/;
assign _48609_ = ~D[44] /*16237*/;
assign _48606_ = _47916_ & _48609_ /*16233*/;
assign _48607_ = _47916_ ^ _48609_ /*16236*/;
assign _48608_ = _48600_ & _48607_ /*16234*/;
assign _48365_ = _48600_ ^ _48607_ /*16235*/;
assign _48605_ = _48606_ | _48608_ /*16232*/;
assign _48614_ = ~D[45] /*16231*/;
assign _48611_ = _47917_ & _48614_ /*16227*/;
assign _48612_ = _47917_ ^ _48614_ /*16230*/;
assign _48613_ = _48605_ & _48612_ /*16228*/;
assign _48366_ = _48605_ ^ _48612_ /*16229*/;
assign _48610_ = _48611_ | _48613_ /*16226*/;
assign _48619_ = ~D[46] /*16225*/;
assign _48616_ = _47918_ & _48619_ /*16221*/;
assign _48617_ = _47918_ ^ _48619_ /*16224*/;
assign _48618_ = _48610_ & _48617_ /*16222*/;
assign _48367_ = _48610_ ^ _48617_ /*16223*/;
assign _48615_ = _48616_ | _48618_ /*16220*/;
assign _48624_ = ~D[47] /*16219*/;
assign _48621_ = _47919_ & _48624_ /*16215*/;
assign _48622_ = _47919_ ^ _48624_ /*16218*/;
assign _48623_ = _48615_ & _48622_ /*16216*/;
assign _48368_ = _48615_ ^ _48622_ /*16217*/;
assign _48620_ = _48621_ | _48623_ /*16214*/;
assign _48629_ = ~D[48] /*16213*/;
assign _48626_ = _47920_ & _48629_ /*16209*/;
assign _48627_ = _47920_ ^ _48629_ /*16212*/;
assign _48628_ = _48620_ & _48627_ /*16210*/;
assign _48369_ = _48620_ ^ _48627_ /*16211*/;
assign _48625_ = _48626_ | _48628_ /*16208*/;
assign _48634_ = ~D[49] /*16207*/;
assign _48631_ = _47921_ & _48634_ /*16203*/;
assign _48632_ = _47921_ ^ _48634_ /*16206*/;
assign _48633_ = _48625_ & _48632_ /*16204*/;
assign _48370_ = _48625_ ^ _48632_ /*16205*/;
assign _48630_ = _48631_ | _48633_ /*16202*/;
assign _48639_ = ~D[50] /*16201*/;
assign _48636_ = _47922_ & _48639_ /*16197*/;
assign _48637_ = _47922_ ^ _48639_ /*16200*/;
assign _48638_ = _48630_ & _48637_ /*16198*/;
assign _48371_ = _48630_ ^ _48637_ /*16199*/;
assign _48635_ = _48636_ | _48638_ /*16196*/;
assign _48644_ = ~D[51] /*16195*/;
assign _48641_ = _47923_ & _48644_ /*16191*/;
assign _48642_ = _47923_ ^ _48644_ /*16194*/;
assign _48643_ = _48635_ & _48642_ /*16192*/;
assign _48372_ = _48635_ ^ _48642_ /*16193*/;
assign _48640_ = _48641_ | _48643_ /*16190*/;
assign _48649_ = ~D[52] /*16189*/;
assign _48646_ = _47924_ & _48649_ /*16185*/;
assign _48647_ = _47924_ ^ _48649_ /*16188*/;
assign _48648_ = _48640_ & _48647_ /*16186*/;
assign _48373_ = _48640_ ^ _48647_ /*16187*/;
assign _48645_ = _48646_ | _48648_ /*16184*/;
assign _48654_ = ~D[53] /*16183*/;
assign _48651_ = _47925_ & _48654_ /*16179*/;
assign _48652_ = _47925_ ^ _48654_ /*16182*/;
assign _48653_ = _48645_ & _48652_ /*16180*/;
assign _48374_ = _48645_ ^ _48652_ /*16181*/;
assign _48650_ = _48651_ | _48653_ /*16178*/;
assign _48659_ = ~D[54] /*16177*/;
assign _48656_ = _47926_ & _48659_ /*16173*/;
assign _48657_ = _47926_ ^ _48659_ /*16176*/;
assign _48658_ = _48650_ & _48657_ /*16174*/;
assign _48375_ = _48650_ ^ _48657_ /*16175*/;
assign _48655_ = _48656_ | _48658_ /*16172*/;
assign _48664_ = ~D[55] /*16171*/;
assign _48661_ = _47927_ & _48664_ /*16167*/;
assign _48662_ = _47927_ ^ _48664_ /*16170*/;
assign _48663_ = _48655_ & _48662_ /*16168*/;
assign _48376_ = _48655_ ^ _48662_ /*16169*/;
assign _48660_ = _48661_ | _48663_ /*16166*/;
assign _48669_ = ~D[56] /*16165*/;
assign _48666_ = _47928_ & _48669_ /*16161*/;
assign _48667_ = _47928_ ^ _48669_ /*16164*/;
assign _48668_ = _48660_ & _48667_ /*16162*/;
assign _48377_ = _48660_ ^ _48667_ /*16163*/;
assign _48665_ = _48666_ | _48668_ /*16160*/;
assign _48674_ = ~D[57] /*16159*/;
assign _48671_ = _47929_ & _48674_ /*16155*/;
assign _48672_ = _47929_ ^ _48674_ /*16158*/;
assign _48673_ = _48665_ & _48672_ /*16156*/;
assign _48378_ = _48665_ ^ _48672_ /*16157*/;
assign _48670_ = _48671_ | _48673_ /*16154*/;
assign _48679_ = ~D[58] /*16153*/;
assign _48676_ = _47930_ & _48679_ /*16149*/;
assign _48677_ = _47930_ ^ _48679_ /*16152*/;
assign _48678_ = _48670_ & _48677_ /*16150*/;
assign _48379_ = _48670_ ^ _48677_ /*16151*/;
assign _48675_ = _48676_ | _48678_ /*16148*/;
assign _48684_ = ~D[59] /*16147*/;
assign _48681_ = _47931_ & _48684_ /*16143*/;
assign _48682_ = _47931_ ^ _48684_ /*16146*/;
assign _48683_ = _48675_ & _48682_ /*16144*/;
assign _48380_ = _48675_ ^ _48682_ /*16145*/;
assign _48680_ = _48681_ | _48683_ /*16142*/;
assign _48689_ = ~D[60] /*16141*/;
assign _48686_ = _47932_ & _48689_ /*16137*/;
assign _48687_ = _47932_ ^ _48689_ /*16140*/;
assign _48688_ = _48680_ & _48687_ /*16138*/;
assign _48381_ = _48680_ ^ _48687_ /*16139*/;
assign _48685_ = _48686_ | _48688_ /*16136*/;
assign _48694_ = ~D[61] /*16135*/;
assign _48691_ = _47933_ & _48694_ /*16131*/;
assign _48692_ = _47933_ ^ _48694_ /*16134*/;
assign _48693_ = _48685_ & _48692_ /*16132*/;
assign _48382_ = _48685_ ^ _48692_ /*16133*/;
assign _48690_ = _48691_ | _48693_ /*16130*/;
assign _48699_ = ~D[62] /*16129*/;
assign _48696_ = _47934_ & _48699_ /*16125*/;
assign _48697_ = _47934_ ^ _48699_ /*16128*/;
assign _48698_ = _48690_ & _48697_ /*16126*/;
assign _48383_ = _48690_ ^ _48697_ /*16127*/;
assign _48695_ = _48696_ | _48698_ /*16124*/;
assign _48700_ = _47935_ & oneWire /*16119*/;
assign _48701_ = _47935_ ^ oneWire /*16122*/;
assign _48702_ = _48695_ & _48701_ /*16120*/;
assign _48384_ = _48695_ ^ _48701_ /*16121*/;
assign Q[9] = _48700_ | _48702_ /*16118*/;
assign _48835_ = ~Q[9] /*15733*/;
assign _48834_ = _48835_ & D[0] /*15732*/;
assign _48837_ = _48321_ & _48834_ /*15727*/;
assign _48838_ = _48321_ ^ _48834_ /*15730*/;
assign _48839_ = zeroWire & _48838_ /*15728*/;
assign _48769_ = zeroWire ^ _48838_ /*15729*/;
assign _48836_ = _48837_ | _48839_ /*15726*/;
assign _48841_ = ~Q[9] /*15725*/;
assign _48840_ = _48841_ & D[1] /*15724*/;
assign _48843_ = _48322_ & _48840_ /*15719*/;
assign _48844_ = _48322_ ^ _48840_ /*15722*/;
assign _48845_ = _48836_ & _48844_ /*15720*/;
assign _48770_ = _48836_ ^ _48844_ /*15721*/;
assign _48842_ = _48843_ | _48845_ /*15718*/;
assign _48847_ = ~Q[9] /*15717*/;
assign _48846_ = _48847_ & D[2] /*15716*/;
assign _48849_ = _48323_ & _48846_ /*15711*/;
assign _48850_ = _48323_ ^ _48846_ /*15714*/;
assign _48851_ = _48842_ & _48850_ /*15712*/;
assign _48771_ = _48842_ ^ _48850_ /*15713*/;
assign _48848_ = _48849_ | _48851_ /*15710*/;
assign _48853_ = ~Q[9] /*15709*/;
assign _48852_ = _48853_ & D[3] /*15708*/;
assign _48855_ = _48324_ & _48852_ /*15703*/;
assign _48856_ = _48324_ ^ _48852_ /*15706*/;
assign _48857_ = _48848_ & _48856_ /*15704*/;
assign _48772_ = _48848_ ^ _48856_ /*15705*/;
assign _48854_ = _48855_ | _48857_ /*15702*/;
assign _48859_ = ~Q[9] /*15701*/;
assign _48858_ = _48859_ & D[4] /*15700*/;
assign _48861_ = _48325_ & _48858_ /*15695*/;
assign _48862_ = _48325_ ^ _48858_ /*15698*/;
assign _48863_ = _48854_ & _48862_ /*15696*/;
assign _48773_ = _48854_ ^ _48862_ /*15697*/;
assign _48860_ = _48861_ | _48863_ /*15694*/;
assign _48865_ = ~Q[9] /*15693*/;
assign _48864_ = _48865_ & D[5] /*15692*/;
assign _48867_ = _48326_ & _48864_ /*15687*/;
assign _48868_ = _48326_ ^ _48864_ /*15690*/;
assign _48869_ = _48860_ & _48868_ /*15688*/;
assign _48774_ = _48860_ ^ _48868_ /*15689*/;
assign _48866_ = _48867_ | _48869_ /*15686*/;
assign _48871_ = ~Q[9] /*15685*/;
assign _48870_ = _48871_ & D[6] /*15684*/;
assign _48873_ = _48327_ & _48870_ /*15679*/;
assign _48874_ = _48327_ ^ _48870_ /*15682*/;
assign _48875_ = _48866_ & _48874_ /*15680*/;
assign _48775_ = _48866_ ^ _48874_ /*15681*/;
assign _48872_ = _48873_ | _48875_ /*15678*/;
assign _48877_ = ~Q[9] /*15677*/;
assign _48876_ = _48877_ & D[7] /*15676*/;
assign _48879_ = _48328_ & _48876_ /*15671*/;
assign _48880_ = _48328_ ^ _48876_ /*15674*/;
assign _48881_ = _48872_ & _48880_ /*15672*/;
assign _48776_ = _48872_ ^ _48880_ /*15673*/;
assign _48878_ = _48879_ | _48881_ /*15670*/;
assign _48883_ = ~Q[9] /*15669*/;
assign _48882_ = _48883_ & D[8] /*15668*/;
assign _48885_ = _48329_ & _48882_ /*15663*/;
assign _48886_ = _48329_ ^ _48882_ /*15666*/;
assign _48887_ = _48878_ & _48886_ /*15664*/;
assign _48777_ = _48878_ ^ _48886_ /*15665*/;
assign _48884_ = _48885_ | _48887_ /*15662*/;
assign _48889_ = ~Q[9] /*15661*/;
assign _48888_ = _48889_ & D[9] /*15660*/;
assign _48891_ = _48330_ & _48888_ /*15655*/;
assign _48892_ = _48330_ ^ _48888_ /*15658*/;
assign _48893_ = _48884_ & _48892_ /*15656*/;
assign _48778_ = _48884_ ^ _48892_ /*15657*/;
assign _48890_ = _48891_ | _48893_ /*15654*/;
assign _48895_ = ~Q[9] /*15653*/;
assign _48894_ = _48895_ & D[10] /*15652*/;
assign _48897_ = _48331_ & _48894_ /*15647*/;
assign _48898_ = _48331_ ^ _48894_ /*15650*/;
assign _48899_ = _48890_ & _48898_ /*15648*/;
assign _48779_ = _48890_ ^ _48898_ /*15649*/;
assign _48896_ = _48897_ | _48899_ /*15646*/;
assign _48901_ = ~Q[9] /*15645*/;
assign _48900_ = _48901_ & D[11] /*15644*/;
assign _48903_ = _48332_ & _48900_ /*15639*/;
assign _48904_ = _48332_ ^ _48900_ /*15642*/;
assign _48905_ = _48896_ & _48904_ /*15640*/;
assign _48780_ = _48896_ ^ _48904_ /*15641*/;
assign _48902_ = _48903_ | _48905_ /*15638*/;
assign _48907_ = ~Q[9] /*15637*/;
assign _48906_ = _48907_ & D[12] /*15636*/;
assign _48909_ = _48333_ & _48906_ /*15631*/;
assign _48910_ = _48333_ ^ _48906_ /*15634*/;
assign _48911_ = _48902_ & _48910_ /*15632*/;
assign _48781_ = _48902_ ^ _48910_ /*15633*/;
assign _48908_ = _48909_ | _48911_ /*15630*/;
assign _48913_ = ~Q[9] /*15629*/;
assign _48912_ = _48913_ & D[13] /*15628*/;
assign _48915_ = _48334_ & _48912_ /*15623*/;
assign _48916_ = _48334_ ^ _48912_ /*15626*/;
assign _48917_ = _48908_ & _48916_ /*15624*/;
assign _48782_ = _48908_ ^ _48916_ /*15625*/;
assign _48914_ = _48915_ | _48917_ /*15622*/;
assign _48919_ = ~Q[9] /*15621*/;
assign _48918_ = _48919_ & D[14] /*15620*/;
assign _48921_ = _48335_ & _48918_ /*15615*/;
assign _48922_ = _48335_ ^ _48918_ /*15618*/;
assign _48923_ = _48914_ & _48922_ /*15616*/;
assign _48783_ = _48914_ ^ _48922_ /*15617*/;
assign _48920_ = _48921_ | _48923_ /*15614*/;
assign _48925_ = ~Q[9] /*15613*/;
assign _48924_ = _48925_ & D[15] /*15612*/;
assign _48927_ = _48336_ & _48924_ /*15607*/;
assign _48928_ = _48336_ ^ _48924_ /*15610*/;
assign _48929_ = _48920_ & _48928_ /*15608*/;
assign _48784_ = _48920_ ^ _48928_ /*15609*/;
assign _48926_ = _48927_ | _48929_ /*15606*/;
assign _48931_ = ~Q[9] /*15605*/;
assign _48930_ = _48931_ & D[16] /*15604*/;
assign _48933_ = _48337_ & _48930_ /*15599*/;
assign _48934_ = _48337_ ^ _48930_ /*15602*/;
assign _48935_ = _48926_ & _48934_ /*15600*/;
assign _48785_ = _48926_ ^ _48934_ /*15601*/;
assign _48932_ = _48933_ | _48935_ /*15598*/;
assign _48937_ = ~Q[9] /*15597*/;
assign _48936_ = _48937_ & D[17] /*15596*/;
assign _48939_ = _48338_ & _48936_ /*15591*/;
assign _48940_ = _48338_ ^ _48936_ /*15594*/;
assign _48941_ = _48932_ & _48940_ /*15592*/;
assign _48786_ = _48932_ ^ _48940_ /*15593*/;
assign _48938_ = _48939_ | _48941_ /*15590*/;
assign _48943_ = ~Q[9] /*15589*/;
assign _48942_ = _48943_ & D[18] /*15588*/;
assign _48945_ = _48339_ & _48942_ /*15583*/;
assign _48946_ = _48339_ ^ _48942_ /*15586*/;
assign _48947_ = _48938_ & _48946_ /*15584*/;
assign _48787_ = _48938_ ^ _48946_ /*15585*/;
assign _48944_ = _48945_ | _48947_ /*15582*/;
assign _48949_ = ~Q[9] /*15581*/;
assign _48948_ = _48949_ & D[19] /*15580*/;
assign _48951_ = _48340_ & _48948_ /*15575*/;
assign _48952_ = _48340_ ^ _48948_ /*15578*/;
assign _48953_ = _48944_ & _48952_ /*15576*/;
assign _48788_ = _48944_ ^ _48952_ /*15577*/;
assign _48950_ = _48951_ | _48953_ /*15574*/;
assign _48955_ = ~Q[9] /*15573*/;
assign _48954_ = _48955_ & D[20] /*15572*/;
assign _48957_ = _48341_ & _48954_ /*15567*/;
assign _48958_ = _48341_ ^ _48954_ /*15570*/;
assign _48959_ = _48950_ & _48958_ /*15568*/;
assign _48789_ = _48950_ ^ _48958_ /*15569*/;
assign _48956_ = _48957_ | _48959_ /*15566*/;
assign _48961_ = ~Q[9] /*15565*/;
assign _48960_ = _48961_ & D[21] /*15564*/;
assign _48963_ = _48342_ & _48960_ /*15559*/;
assign _48964_ = _48342_ ^ _48960_ /*15562*/;
assign _48965_ = _48956_ & _48964_ /*15560*/;
assign _48790_ = _48956_ ^ _48964_ /*15561*/;
assign _48962_ = _48963_ | _48965_ /*15558*/;
assign _48967_ = ~Q[9] /*15557*/;
assign _48966_ = _48967_ & D[22] /*15556*/;
assign _48969_ = _48343_ & _48966_ /*15551*/;
assign _48970_ = _48343_ ^ _48966_ /*15554*/;
assign _48971_ = _48962_ & _48970_ /*15552*/;
assign _48791_ = _48962_ ^ _48970_ /*15553*/;
assign _48968_ = _48969_ | _48971_ /*15550*/;
assign _48973_ = ~Q[9] /*15549*/;
assign _48972_ = _48973_ & D[23] /*15548*/;
assign _48975_ = _48344_ & _48972_ /*15543*/;
assign _48976_ = _48344_ ^ _48972_ /*15546*/;
assign _48977_ = _48968_ & _48976_ /*15544*/;
assign _48792_ = _48968_ ^ _48976_ /*15545*/;
assign _48974_ = _48975_ | _48977_ /*15542*/;
assign _48979_ = ~Q[9] /*15541*/;
assign _48978_ = _48979_ & D[24] /*15540*/;
assign _48981_ = _48345_ & _48978_ /*15535*/;
assign _48982_ = _48345_ ^ _48978_ /*15538*/;
assign _48983_ = _48974_ & _48982_ /*15536*/;
assign _48793_ = _48974_ ^ _48982_ /*15537*/;
assign _48980_ = _48981_ | _48983_ /*15534*/;
assign _48985_ = ~Q[9] /*15533*/;
assign _48984_ = _48985_ & D[25] /*15532*/;
assign _48987_ = _48346_ & _48984_ /*15527*/;
assign _48988_ = _48346_ ^ _48984_ /*15530*/;
assign _48989_ = _48980_ & _48988_ /*15528*/;
assign _48794_ = _48980_ ^ _48988_ /*15529*/;
assign _48986_ = _48987_ | _48989_ /*15526*/;
assign _48991_ = ~Q[9] /*15525*/;
assign _48990_ = _48991_ & D[26] /*15524*/;
assign _48993_ = _48347_ & _48990_ /*15519*/;
assign _48994_ = _48347_ ^ _48990_ /*15522*/;
assign _48995_ = _48986_ & _48994_ /*15520*/;
assign _48795_ = _48986_ ^ _48994_ /*15521*/;
assign _48992_ = _48993_ | _48995_ /*15518*/;
assign _48997_ = ~Q[9] /*15517*/;
assign _48996_ = _48997_ & D[27] /*15516*/;
assign _48999_ = _48348_ & _48996_ /*15511*/;
assign _49000_ = _48348_ ^ _48996_ /*15514*/;
assign _49001_ = _48992_ & _49000_ /*15512*/;
assign _48796_ = _48992_ ^ _49000_ /*15513*/;
assign _48998_ = _48999_ | _49001_ /*15510*/;
assign _49003_ = ~Q[9] /*15509*/;
assign _49002_ = _49003_ & D[28] /*15508*/;
assign _49005_ = _48349_ & _49002_ /*15503*/;
assign _49006_ = _48349_ ^ _49002_ /*15506*/;
assign _49007_ = _48998_ & _49006_ /*15504*/;
assign _48797_ = _48998_ ^ _49006_ /*15505*/;
assign _49004_ = _49005_ | _49007_ /*15502*/;
assign _49009_ = ~Q[9] /*15501*/;
assign _49008_ = _49009_ & D[29] /*15500*/;
assign _49011_ = _48350_ & _49008_ /*15495*/;
assign _49012_ = _48350_ ^ _49008_ /*15498*/;
assign _49013_ = _49004_ & _49012_ /*15496*/;
assign _48798_ = _49004_ ^ _49012_ /*15497*/;
assign _49010_ = _49011_ | _49013_ /*15494*/;
assign _49015_ = ~Q[9] /*15493*/;
assign _49014_ = _49015_ & D[30] /*15492*/;
assign _49017_ = _48351_ & _49014_ /*15487*/;
assign _49018_ = _48351_ ^ _49014_ /*15490*/;
assign _49019_ = _49010_ & _49018_ /*15488*/;
assign _48799_ = _49010_ ^ _49018_ /*15489*/;
assign _49016_ = _49017_ | _49019_ /*15486*/;
assign _49021_ = ~Q[9] /*15485*/;
assign _49020_ = _49021_ & D[31] /*15484*/;
assign _49023_ = _48352_ & _49020_ /*15479*/;
assign _49024_ = _48352_ ^ _49020_ /*15482*/;
assign _49025_ = _49016_ & _49024_ /*15480*/;
assign _48800_ = _49016_ ^ _49024_ /*15481*/;
assign _49022_ = _49023_ | _49025_ /*15478*/;
assign _49027_ = ~Q[9] /*15477*/;
assign _49026_ = _49027_ & D[32] /*15476*/;
assign _49029_ = _48353_ & _49026_ /*15471*/;
assign _49030_ = _48353_ ^ _49026_ /*15474*/;
assign _49031_ = _49022_ & _49030_ /*15472*/;
assign _48801_ = _49022_ ^ _49030_ /*15473*/;
assign _49028_ = _49029_ | _49031_ /*15470*/;
assign _49033_ = ~Q[9] /*15469*/;
assign _49032_ = _49033_ & D[33] /*15468*/;
assign _49035_ = _48354_ & _49032_ /*15463*/;
assign _49036_ = _48354_ ^ _49032_ /*15466*/;
assign _49037_ = _49028_ & _49036_ /*15464*/;
assign _48802_ = _49028_ ^ _49036_ /*15465*/;
assign _49034_ = _49035_ | _49037_ /*15462*/;
assign _49039_ = ~Q[9] /*15461*/;
assign _49038_ = _49039_ & D[34] /*15460*/;
assign _49041_ = _48355_ & _49038_ /*15455*/;
assign _49042_ = _48355_ ^ _49038_ /*15458*/;
assign _49043_ = _49034_ & _49042_ /*15456*/;
assign _48803_ = _49034_ ^ _49042_ /*15457*/;
assign _49040_ = _49041_ | _49043_ /*15454*/;
assign _49045_ = ~Q[9] /*15453*/;
assign _49044_ = _49045_ & D[35] /*15452*/;
assign _49047_ = _48356_ & _49044_ /*15447*/;
assign _49048_ = _48356_ ^ _49044_ /*15450*/;
assign _49049_ = _49040_ & _49048_ /*15448*/;
assign _48804_ = _49040_ ^ _49048_ /*15449*/;
assign _49046_ = _49047_ | _49049_ /*15446*/;
assign _49051_ = ~Q[9] /*15445*/;
assign _49050_ = _49051_ & D[36] /*15444*/;
assign _49053_ = _48357_ & _49050_ /*15439*/;
assign _49054_ = _48357_ ^ _49050_ /*15442*/;
assign _49055_ = _49046_ & _49054_ /*15440*/;
assign _48805_ = _49046_ ^ _49054_ /*15441*/;
assign _49052_ = _49053_ | _49055_ /*15438*/;
assign _49057_ = ~Q[9] /*15437*/;
assign _49056_ = _49057_ & D[37] /*15436*/;
assign _49059_ = _48358_ & _49056_ /*15431*/;
assign _49060_ = _48358_ ^ _49056_ /*15434*/;
assign _49061_ = _49052_ & _49060_ /*15432*/;
assign _48806_ = _49052_ ^ _49060_ /*15433*/;
assign _49058_ = _49059_ | _49061_ /*15430*/;
assign _49063_ = ~Q[9] /*15429*/;
assign _49062_ = _49063_ & D[38] /*15428*/;
assign _49065_ = _48359_ & _49062_ /*15423*/;
assign _49066_ = _48359_ ^ _49062_ /*15426*/;
assign _49067_ = _49058_ & _49066_ /*15424*/;
assign _48807_ = _49058_ ^ _49066_ /*15425*/;
assign _49064_ = _49065_ | _49067_ /*15422*/;
assign _49069_ = ~Q[9] /*15421*/;
assign _49068_ = _49069_ & D[39] /*15420*/;
assign _49071_ = _48360_ & _49068_ /*15415*/;
assign _49072_ = _48360_ ^ _49068_ /*15418*/;
assign _49073_ = _49064_ & _49072_ /*15416*/;
assign _48808_ = _49064_ ^ _49072_ /*15417*/;
assign _49070_ = _49071_ | _49073_ /*15414*/;
assign _49075_ = ~Q[9] /*15413*/;
assign _49074_ = _49075_ & D[40] /*15412*/;
assign _49077_ = _48361_ & _49074_ /*15407*/;
assign _49078_ = _48361_ ^ _49074_ /*15410*/;
assign _49079_ = _49070_ & _49078_ /*15408*/;
assign _48809_ = _49070_ ^ _49078_ /*15409*/;
assign _49076_ = _49077_ | _49079_ /*15406*/;
assign _49081_ = ~Q[9] /*15405*/;
assign _49080_ = _49081_ & D[41] /*15404*/;
assign _49083_ = _48362_ & _49080_ /*15399*/;
assign _49084_ = _48362_ ^ _49080_ /*15402*/;
assign _49085_ = _49076_ & _49084_ /*15400*/;
assign _48810_ = _49076_ ^ _49084_ /*15401*/;
assign _49082_ = _49083_ | _49085_ /*15398*/;
assign _49087_ = ~Q[9] /*15397*/;
assign _49086_ = _49087_ & D[42] /*15396*/;
assign _49089_ = _48363_ & _49086_ /*15391*/;
assign _49090_ = _48363_ ^ _49086_ /*15394*/;
assign _49091_ = _49082_ & _49090_ /*15392*/;
assign _48811_ = _49082_ ^ _49090_ /*15393*/;
assign _49088_ = _49089_ | _49091_ /*15390*/;
assign _49093_ = ~Q[9] /*15389*/;
assign _49092_ = _49093_ & D[43] /*15388*/;
assign _49095_ = _48364_ & _49092_ /*15383*/;
assign _49096_ = _48364_ ^ _49092_ /*15386*/;
assign _49097_ = _49088_ & _49096_ /*15384*/;
assign _48812_ = _49088_ ^ _49096_ /*15385*/;
assign _49094_ = _49095_ | _49097_ /*15382*/;
assign _49099_ = ~Q[9] /*15381*/;
assign _49098_ = _49099_ & D[44] /*15380*/;
assign _49101_ = _48365_ & _49098_ /*15375*/;
assign _49102_ = _48365_ ^ _49098_ /*15378*/;
assign _49103_ = _49094_ & _49102_ /*15376*/;
assign _48813_ = _49094_ ^ _49102_ /*15377*/;
assign _49100_ = _49101_ | _49103_ /*15374*/;
assign _49105_ = ~Q[9] /*15373*/;
assign _49104_ = _49105_ & D[45] /*15372*/;
assign _49107_ = _48366_ & _49104_ /*15367*/;
assign _49108_ = _48366_ ^ _49104_ /*15370*/;
assign _49109_ = _49100_ & _49108_ /*15368*/;
assign _48814_ = _49100_ ^ _49108_ /*15369*/;
assign _49106_ = _49107_ | _49109_ /*15366*/;
assign _49111_ = ~Q[9] /*15365*/;
assign _49110_ = _49111_ & D[46] /*15364*/;
assign _49113_ = _48367_ & _49110_ /*15359*/;
assign _49114_ = _48367_ ^ _49110_ /*15362*/;
assign _49115_ = _49106_ & _49114_ /*15360*/;
assign _48815_ = _49106_ ^ _49114_ /*15361*/;
assign _49112_ = _49113_ | _49115_ /*15358*/;
assign _49117_ = ~Q[9] /*15357*/;
assign _49116_ = _49117_ & D[47] /*15356*/;
assign _49119_ = _48368_ & _49116_ /*15351*/;
assign _49120_ = _48368_ ^ _49116_ /*15354*/;
assign _49121_ = _49112_ & _49120_ /*15352*/;
assign _48816_ = _49112_ ^ _49120_ /*15353*/;
assign _49118_ = _49119_ | _49121_ /*15350*/;
assign _49123_ = ~Q[9] /*15349*/;
assign _49122_ = _49123_ & D[48] /*15348*/;
assign _49125_ = _48369_ & _49122_ /*15343*/;
assign _49126_ = _48369_ ^ _49122_ /*15346*/;
assign _49127_ = _49118_ & _49126_ /*15344*/;
assign _48817_ = _49118_ ^ _49126_ /*15345*/;
assign _49124_ = _49125_ | _49127_ /*15342*/;
assign _49129_ = ~Q[9] /*15341*/;
assign _49128_ = _49129_ & D[49] /*15340*/;
assign _49131_ = _48370_ & _49128_ /*15335*/;
assign _49132_ = _48370_ ^ _49128_ /*15338*/;
assign _49133_ = _49124_ & _49132_ /*15336*/;
assign _48818_ = _49124_ ^ _49132_ /*15337*/;
assign _49130_ = _49131_ | _49133_ /*15334*/;
assign _49135_ = ~Q[9] /*15333*/;
assign _49134_ = _49135_ & D[50] /*15332*/;
assign _49137_ = _48371_ & _49134_ /*15327*/;
assign _49138_ = _48371_ ^ _49134_ /*15330*/;
assign _49139_ = _49130_ & _49138_ /*15328*/;
assign _48819_ = _49130_ ^ _49138_ /*15329*/;
assign _49136_ = _49137_ | _49139_ /*15326*/;
assign _49141_ = ~Q[9] /*15325*/;
assign _49140_ = _49141_ & D[51] /*15324*/;
assign _49143_ = _48372_ & _49140_ /*15319*/;
assign _49144_ = _48372_ ^ _49140_ /*15322*/;
assign _49145_ = _49136_ & _49144_ /*15320*/;
assign _48820_ = _49136_ ^ _49144_ /*15321*/;
assign _49142_ = _49143_ | _49145_ /*15318*/;
assign _49147_ = ~Q[9] /*15317*/;
assign _49146_ = _49147_ & D[52] /*15316*/;
assign _49149_ = _48373_ & _49146_ /*15311*/;
assign _49150_ = _48373_ ^ _49146_ /*15314*/;
assign _49151_ = _49142_ & _49150_ /*15312*/;
assign _48821_ = _49142_ ^ _49150_ /*15313*/;
assign _49148_ = _49149_ | _49151_ /*15310*/;
assign _49153_ = ~Q[9] /*15309*/;
assign _49152_ = _49153_ & D[53] /*15308*/;
assign _49155_ = _48374_ & _49152_ /*15303*/;
assign _49156_ = _48374_ ^ _49152_ /*15306*/;
assign _49157_ = _49148_ & _49156_ /*15304*/;
assign _48822_ = _49148_ ^ _49156_ /*15305*/;
assign _49154_ = _49155_ | _49157_ /*15302*/;
assign _49159_ = ~Q[9] /*15301*/;
assign _49158_ = _49159_ & D[54] /*15300*/;
assign _49161_ = _48375_ & _49158_ /*15295*/;
assign _49162_ = _48375_ ^ _49158_ /*15298*/;
assign _49163_ = _49154_ & _49162_ /*15296*/;
assign _48823_ = _49154_ ^ _49162_ /*15297*/;
assign _49160_ = _49161_ | _49163_ /*15294*/;
assign _49165_ = ~Q[9] /*15293*/;
assign _49164_ = _49165_ & D[55] /*15292*/;
assign _49167_ = _48376_ & _49164_ /*15287*/;
assign _49168_ = _48376_ ^ _49164_ /*15290*/;
assign _49169_ = _49160_ & _49168_ /*15288*/;
assign _48824_ = _49160_ ^ _49168_ /*15289*/;
assign _49166_ = _49167_ | _49169_ /*15286*/;
assign _49171_ = ~Q[9] /*15285*/;
assign _49170_ = _49171_ & D[56] /*15284*/;
assign _49173_ = _48377_ & _49170_ /*15279*/;
assign _49174_ = _48377_ ^ _49170_ /*15282*/;
assign _49175_ = _49166_ & _49174_ /*15280*/;
assign _48825_ = _49166_ ^ _49174_ /*15281*/;
assign _49172_ = _49173_ | _49175_ /*15278*/;
assign _49177_ = ~Q[9] /*15277*/;
assign _49176_ = _49177_ & D[57] /*15276*/;
assign _49179_ = _48378_ & _49176_ /*15271*/;
assign _49180_ = _48378_ ^ _49176_ /*15274*/;
assign _49181_ = _49172_ & _49180_ /*15272*/;
assign _48826_ = _49172_ ^ _49180_ /*15273*/;
assign _49178_ = _49179_ | _49181_ /*15270*/;
assign _49183_ = ~Q[9] /*15269*/;
assign _49182_ = _49183_ & D[58] /*15268*/;
assign _49185_ = _48379_ & _49182_ /*15263*/;
assign _49186_ = _48379_ ^ _49182_ /*15266*/;
assign _49187_ = _49178_ & _49186_ /*15264*/;
assign _48827_ = _49178_ ^ _49186_ /*15265*/;
assign _49184_ = _49185_ | _49187_ /*15262*/;
assign _49189_ = ~Q[9] /*15261*/;
assign _49188_ = _49189_ & D[59] /*15260*/;
assign _49191_ = _48380_ & _49188_ /*15255*/;
assign _49192_ = _48380_ ^ _49188_ /*15258*/;
assign _49193_ = _49184_ & _49192_ /*15256*/;
assign _48828_ = _49184_ ^ _49192_ /*15257*/;
assign _49190_ = _49191_ | _49193_ /*15254*/;
assign _49195_ = ~Q[9] /*15253*/;
assign _49194_ = _49195_ & D[60] /*15252*/;
assign _49197_ = _48381_ & _49194_ /*15247*/;
assign _49198_ = _48381_ ^ _49194_ /*15250*/;
assign _49199_ = _49190_ & _49198_ /*15248*/;
assign _48829_ = _49190_ ^ _49198_ /*15249*/;
assign _49196_ = _49197_ | _49199_ /*15246*/;
assign _49201_ = ~Q[9] /*15245*/;
assign _49200_ = _49201_ & D[61] /*15244*/;
assign _49203_ = _48382_ & _49200_ /*15239*/;
assign _49204_ = _48382_ ^ _49200_ /*15242*/;
assign _49205_ = _49196_ & _49204_ /*15240*/;
assign _48830_ = _49196_ ^ _49204_ /*15241*/;
assign _49202_ = _49203_ | _49205_ /*15238*/;
assign _49207_ = ~Q[9] /*15237*/;
assign _49206_ = _49207_ & D[62] /*15236*/;
assign _49209_ = _48383_ & _49206_ /*15231*/;
assign _49210_ = _48383_ ^ _49206_ /*15234*/;
assign _49211_ = _49202_ & _49210_ /*15232*/;
assign _48831_ = _49202_ ^ _49210_ /*15233*/;
assign _49208_ = _49209_ | _49211_ /*15230*/;
assign _49213_ = ~Q[9] /*15229*/;
assign _49212_ = _49213_ & zeroWire /*15228*/;
assign _49214_ = _48384_ ^ _49212_ /*15226*/;
assign _48832_ = _49214_ ^ _49208_ /*15225*/;
assign _49285_ = ~D[0] /*14971*/;
assign _49282_ = R_0[8] & _49285_ /*14967*/;
assign _49283_ = R_0[8] ^ _49285_ /*14970*/;
assign _49284_ = oneWire & _49283_ /*14968*/;
assign _49217_ = oneWire ^ _49283_ /*14969*/;
assign _49281_ = _49282_ | _49284_ /*14966*/;
assign _49290_ = ~D[1] /*14965*/;
assign _49287_ = _48769_ & _49290_ /*14961*/;
assign _49288_ = _48769_ ^ _49290_ /*14964*/;
assign _49289_ = _49281_ & _49288_ /*14962*/;
assign _49218_ = _49281_ ^ _49288_ /*14963*/;
assign _49286_ = _49287_ | _49289_ /*14960*/;
assign _49295_ = ~D[2] /*14959*/;
assign _49292_ = _48770_ & _49295_ /*14955*/;
assign _49293_ = _48770_ ^ _49295_ /*14958*/;
assign _49294_ = _49286_ & _49293_ /*14956*/;
assign _49219_ = _49286_ ^ _49293_ /*14957*/;
assign _49291_ = _49292_ | _49294_ /*14954*/;
assign _49300_ = ~D[3] /*14953*/;
assign _49297_ = _48771_ & _49300_ /*14949*/;
assign _49298_ = _48771_ ^ _49300_ /*14952*/;
assign _49299_ = _49291_ & _49298_ /*14950*/;
assign _49220_ = _49291_ ^ _49298_ /*14951*/;
assign _49296_ = _49297_ | _49299_ /*14948*/;
assign _49305_ = ~D[4] /*14947*/;
assign _49302_ = _48772_ & _49305_ /*14943*/;
assign _49303_ = _48772_ ^ _49305_ /*14946*/;
assign _49304_ = _49296_ & _49303_ /*14944*/;
assign _49221_ = _49296_ ^ _49303_ /*14945*/;
assign _49301_ = _49302_ | _49304_ /*14942*/;
assign _49310_ = ~D[5] /*14941*/;
assign _49307_ = _48773_ & _49310_ /*14937*/;
assign _49308_ = _48773_ ^ _49310_ /*14940*/;
assign _49309_ = _49301_ & _49308_ /*14938*/;
assign _49222_ = _49301_ ^ _49308_ /*14939*/;
assign _49306_ = _49307_ | _49309_ /*14936*/;
assign _49315_ = ~D[6] /*14935*/;
assign _49312_ = _48774_ & _49315_ /*14931*/;
assign _49313_ = _48774_ ^ _49315_ /*14934*/;
assign _49314_ = _49306_ & _49313_ /*14932*/;
assign _49223_ = _49306_ ^ _49313_ /*14933*/;
assign _49311_ = _49312_ | _49314_ /*14930*/;
assign _49320_ = ~D[7] /*14929*/;
assign _49317_ = _48775_ & _49320_ /*14925*/;
assign _49318_ = _48775_ ^ _49320_ /*14928*/;
assign _49319_ = _49311_ & _49318_ /*14926*/;
assign _49224_ = _49311_ ^ _49318_ /*14927*/;
assign _49316_ = _49317_ | _49319_ /*14924*/;
assign _49325_ = ~D[8] /*14923*/;
assign _49322_ = _48776_ & _49325_ /*14919*/;
assign _49323_ = _48776_ ^ _49325_ /*14922*/;
assign _49324_ = _49316_ & _49323_ /*14920*/;
assign _49225_ = _49316_ ^ _49323_ /*14921*/;
assign _49321_ = _49322_ | _49324_ /*14918*/;
assign _49330_ = ~D[9] /*14917*/;
assign _49327_ = _48777_ & _49330_ /*14913*/;
assign _49328_ = _48777_ ^ _49330_ /*14916*/;
assign _49329_ = _49321_ & _49328_ /*14914*/;
assign _49226_ = _49321_ ^ _49328_ /*14915*/;
assign _49326_ = _49327_ | _49329_ /*14912*/;
assign _49335_ = ~D[10] /*14911*/;
assign _49332_ = _48778_ & _49335_ /*14907*/;
assign _49333_ = _48778_ ^ _49335_ /*14910*/;
assign _49334_ = _49326_ & _49333_ /*14908*/;
assign _49227_ = _49326_ ^ _49333_ /*14909*/;
assign _49331_ = _49332_ | _49334_ /*14906*/;
assign _49340_ = ~D[11] /*14905*/;
assign _49337_ = _48779_ & _49340_ /*14901*/;
assign _49338_ = _48779_ ^ _49340_ /*14904*/;
assign _49339_ = _49331_ & _49338_ /*14902*/;
assign _49228_ = _49331_ ^ _49338_ /*14903*/;
assign _49336_ = _49337_ | _49339_ /*14900*/;
assign _49345_ = ~D[12] /*14899*/;
assign _49342_ = _48780_ & _49345_ /*14895*/;
assign _49343_ = _48780_ ^ _49345_ /*14898*/;
assign _49344_ = _49336_ & _49343_ /*14896*/;
assign _49229_ = _49336_ ^ _49343_ /*14897*/;
assign _49341_ = _49342_ | _49344_ /*14894*/;
assign _49350_ = ~D[13] /*14893*/;
assign _49347_ = _48781_ & _49350_ /*14889*/;
assign _49348_ = _48781_ ^ _49350_ /*14892*/;
assign _49349_ = _49341_ & _49348_ /*14890*/;
assign _49230_ = _49341_ ^ _49348_ /*14891*/;
assign _49346_ = _49347_ | _49349_ /*14888*/;
assign _49355_ = ~D[14] /*14887*/;
assign _49352_ = _48782_ & _49355_ /*14883*/;
assign _49353_ = _48782_ ^ _49355_ /*14886*/;
assign _49354_ = _49346_ & _49353_ /*14884*/;
assign _49231_ = _49346_ ^ _49353_ /*14885*/;
assign _49351_ = _49352_ | _49354_ /*14882*/;
assign _49360_ = ~D[15] /*14881*/;
assign _49357_ = _48783_ & _49360_ /*14877*/;
assign _49358_ = _48783_ ^ _49360_ /*14880*/;
assign _49359_ = _49351_ & _49358_ /*14878*/;
assign _49232_ = _49351_ ^ _49358_ /*14879*/;
assign _49356_ = _49357_ | _49359_ /*14876*/;
assign _49365_ = ~D[16] /*14875*/;
assign _49362_ = _48784_ & _49365_ /*14871*/;
assign _49363_ = _48784_ ^ _49365_ /*14874*/;
assign _49364_ = _49356_ & _49363_ /*14872*/;
assign _49233_ = _49356_ ^ _49363_ /*14873*/;
assign _49361_ = _49362_ | _49364_ /*14870*/;
assign _49370_ = ~D[17] /*14869*/;
assign _49367_ = _48785_ & _49370_ /*14865*/;
assign _49368_ = _48785_ ^ _49370_ /*14868*/;
assign _49369_ = _49361_ & _49368_ /*14866*/;
assign _49234_ = _49361_ ^ _49368_ /*14867*/;
assign _49366_ = _49367_ | _49369_ /*14864*/;
assign _49375_ = ~D[18] /*14863*/;
assign _49372_ = _48786_ & _49375_ /*14859*/;
assign _49373_ = _48786_ ^ _49375_ /*14862*/;
assign _49374_ = _49366_ & _49373_ /*14860*/;
assign _49235_ = _49366_ ^ _49373_ /*14861*/;
assign _49371_ = _49372_ | _49374_ /*14858*/;
assign _49380_ = ~D[19] /*14857*/;
assign _49377_ = _48787_ & _49380_ /*14853*/;
assign _49378_ = _48787_ ^ _49380_ /*14856*/;
assign _49379_ = _49371_ & _49378_ /*14854*/;
assign _49236_ = _49371_ ^ _49378_ /*14855*/;
assign _49376_ = _49377_ | _49379_ /*14852*/;
assign _49385_ = ~D[20] /*14851*/;
assign _49382_ = _48788_ & _49385_ /*14847*/;
assign _49383_ = _48788_ ^ _49385_ /*14850*/;
assign _49384_ = _49376_ & _49383_ /*14848*/;
assign _49237_ = _49376_ ^ _49383_ /*14849*/;
assign _49381_ = _49382_ | _49384_ /*14846*/;
assign _49390_ = ~D[21] /*14845*/;
assign _49387_ = _48789_ & _49390_ /*14841*/;
assign _49388_ = _48789_ ^ _49390_ /*14844*/;
assign _49389_ = _49381_ & _49388_ /*14842*/;
assign _49238_ = _49381_ ^ _49388_ /*14843*/;
assign _49386_ = _49387_ | _49389_ /*14840*/;
assign _49395_ = ~D[22] /*14839*/;
assign _49392_ = _48790_ & _49395_ /*14835*/;
assign _49393_ = _48790_ ^ _49395_ /*14838*/;
assign _49394_ = _49386_ & _49393_ /*14836*/;
assign _49239_ = _49386_ ^ _49393_ /*14837*/;
assign _49391_ = _49392_ | _49394_ /*14834*/;
assign _49400_ = ~D[23] /*14833*/;
assign _49397_ = _48791_ & _49400_ /*14829*/;
assign _49398_ = _48791_ ^ _49400_ /*14832*/;
assign _49399_ = _49391_ & _49398_ /*14830*/;
assign _49240_ = _49391_ ^ _49398_ /*14831*/;
assign _49396_ = _49397_ | _49399_ /*14828*/;
assign _49405_ = ~D[24] /*14827*/;
assign _49402_ = _48792_ & _49405_ /*14823*/;
assign _49403_ = _48792_ ^ _49405_ /*14826*/;
assign _49404_ = _49396_ & _49403_ /*14824*/;
assign _49241_ = _49396_ ^ _49403_ /*14825*/;
assign _49401_ = _49402_ | _49404_ /*14822*/;
assign _49410_ = ~D[25] /*14821*/;
assign _49407_ = _48793_ & _49410_ /*14817*/;
assign _49408_ = _48793_ ^ _49410_ /*14820*/;
assign _49409_ = _49401_ & _49408_ /*14818*/;
assign _49242_ = _49401_ ^ _49408_ /*14819*/;
assign _49406_ = _49407_ | _49409_ /*14816*/;
assign _49415_ = ~D[26] /*14815*/;
assign _49412_ = _48794_ & _49415_ /*14811*/;
assign _49413_ = _48794_ ^ _49415_ /*14814*/;
assign _49414_ = _49406_ & _49413_ /*14812*/;
assign _49243_ = _49406_ ^ _49413_ /*14813*/;
assign _49411_ = _49412_ | _49414_ /*14810*/;
assign _49420_ = ~D[27] /*14809*/;
assign _49417_ = _48795_ & _49420_ /*14805*/;
assign _49418_ = _48795_ ^ _49420_ /*14808*/;
assign _49419_ = _49411_ & _49418_ /*14806*/;
assign _49244_ = _49411_ ^ _49418_ /*14807*/;
assign _49416_ = _49417_ | _49419_ /*14804*/;
assign _49425_ = ~D[28] /*14803*/;
assign _49422_ = _48796_ & _49425_ /*14799*/;
assign _49423_ = _48796_ ^ _49425_ /*14802*/;
assign _49424_ = _49416_ & _49423_ /*14800*/;
assign _49245_ = _49416_ ^ _49423_ /*14801*/;
assign _49421_ = _49422_ | _49424_ /*14798*/;
assign _49430_ = ~D[29] /*14797*/;
assign _49427_ = _48797_ & _49430_ /*14793*/;
assign _49428_ = _48797_ ^ _49430_ /*14796*/;
assign _49429_ = _49421_ & _49428_ /*14794*/;
assign _49246_ = _49421_ ^ _49428_ /*14795*/;
assign _49426_ = _49427_ | _49429_ /*14792*/;
assign _49435_ = ~D[30] /*14791*/;
assign _49432_ = _48798_ & _49435_ /*14787*/;
assign _49433_ = _48798_ ^ _49435_ /*14790*/;
assign _49434_ = _49426_ & _49433_ /*14788*/;
assign _49247_ = _49426_ ^ _49433_ /*14789*/;
assign _49431_ = _49432_ | _49434_ /*14786*/;
assign _49440_ = ~D[31] /*14785*/;
assign _49437_ = _48799_ & _49440_ /*14781*/;
assign _49438_ = _48799_ ^ _49440_ /*14784*/;
assign _49439_ = _49431_ & _49438_ /*14782*/;
assign _49248_ = _49431_ ^ _49438_ /*14783*/;
assign _49436_ = _49437_ | _49439_ /*14780*/;
assign _49445_ = ~D[32] /*14779*/;
assign _49442_ = _48800_ & _49445_ /*14775*/;
assign _49443_ = _48800_ ^ _49445_ /*14778*/;
assign _49444_ = _49436_ & _49443_ /*14776*/;
assign _49249_ = _49436_ ^ _49443_ /*14777*/;
assign _49441_ = _49442_ | _49444_ /*14774*/;
assign _49450_ = ~D[33] /*14773*/;
assign _49447_ = _48801_ & _49450_ /*14769*/;
assign _49448_ = _48801_ ^ _49450_ /*14772*/;
assign _49449_ = _49441_ & _49448_ /*14770*/;
assign _49250_ = _49441_ ^ _49448_ /*14771*/;
assign _49446_ = _49447_ | _49449_ /*14768*/;
assign _49455_ = ~D[34] /*14767*/;
assign _49452_ = _48802_ & _49455_ /*14763*/;
assign _49453_ = _48802_ ^ _49455_ /*14766*/;
assign _49454_ = _49446_ & _49453_ /*14764*/;
assign _49251_ = _49446_ ^ _49453_ /*14765*/;
assign _49451_ = _49452_ | _49454_ /*14762*/;
assign _49460_ = ~D[35] /*14761*/;
assign _49457_ = _48803_ & _49460_ /*14757*/;
assign _49458_ = _48803_ ^ _49460_ /*14760*/;
assign _49459_ = _49451_ & _49458_ /*14758*/;
assign _49252_ = _49451_ ^ _49458_ /*14759*/;
assign _49456_ = _49457_ | _49459_ /*14756*/;
assign _49465_ = ~D[36] /*14755*/;
assign _49462_ = _48804_ & _49465_ /*14751*/;
assign _49463_ = _48804_ ^ _49465_ /*14754*/;
assign _49464_ = _49456_ & _49463_ /*14752*/;
assign _49253_ = _49456_ ^ _49463_ /*14753*/;
assign _49461_ = _49462_ | _49464_ /*14750*/;
assign _49470_ = ~D[37] /*14749*/;
assign _49467_ = _48805_ & _49470_ /*14745*/;
assign _49468_ = _48805_ ^ _49470_ /*14748*/;
assign _49469_ = _49461_ & _49468_ /*14746*/;
assign _49254_ = _49461_ ^ _49468_ /*14747*/;
assign _49466_ = _49467_ | _49469_ /*14744*/;
assign _49475_ = ~D[38] /*14743*/;
assign _49472_ = _48806_ & _49475_ /*14739*/;
assign _49473_ = _48806_ ^ _49475_ /*14742*/;
assign _49474_ = _49466_ & _49473_ /*14740*/;
assign _49255_ = _49466_ ^ _49473_ /*14741*/;
assign _49471_ = _49472_ | _49474_ /*14738*/;
assign _49480_ = ~D[39] /*14737*/;
assign _49477_ = _48807_ & _49480_ /*14733*/;
assign _49478_ = _48807_ ^ _49480_ /*14736*/;
assign _49479_ = _49471_ & _49478_ /*14734*/;
assign _49256_ = _49471_ ^ _49478_ /*14735*/;
assign _49476_ = _49477_ | _49479_ /*14732*/;
assign _49485_ = ~D[40] /*14731*/;
assign _49482_ = _48808_ & _49485_ /*14727*/;
assign _49483_ = _48808_ ^ _49485_ /*14730*/;
assign _49484_ = _49476_ & _49483_ /*14728*/;
assign _49257_ = _49476_ ^ _49483_ /*14729*/;
assign _49481_ = _49482_ | _49484_ /*14726*/;
assign _49490_ = ~D[41] /*14725*/;
assign _49487_ = _48809_ & _49490_ /*14721*/;
assign _49488_ = _48809_ ^ _49490_ /*14724*/;
assign _49489_ = _49481_ & _49488_ /*14722*/;
assign _49258_ = _49481_ ^ _49488_ /*14723*/;
assign _49486_ = _49487_ | _49489_ /*14720*/;
assign _49495_ = ~D[42] /*14719*/;
assign _49492_ = _48810_ & _49495_ /*14715*/;
assign _49493_ = _48810_ ^ _49495_ /*14718*/;
assign _49494_ = _49486_ & _49493_ /*14716*/;
assign _49259_ = _49486_ ^ _49493_ /*14717*/;
assign _49491_ = _49492_ | _49494_ /*14714*/;
assign _49500_ = ~D[43] /*14713*/;
assign _49497_ = _48811_ & _49500_ /*14709*/;
assign _49498_ = _48811_ ^ _49500_ /*14712*/;
assign _49499_ = _49491_ & _49498_ /*14710*/;
assign _49260_ = _49491_ ^ _49498_ /*14711*/;
assign _49496_ = _49497_ | _49499_ /*14708*/;
assign _49505_ = ~D[44] /*14707*/;
assign _49502_ = _48812_ & _49505_ /*14703*/;
assign _49503_ = _48812_ ^ _49505_ /*14706*/;
assign _49504_ = _49496_ & _49503_ /*14704*/;
assign _49261_ = _49496_ ^ _49503_ /*14705*/;
assign _49501_ = _49502_ | _49504_ /*14702*/;
assign _49510_ = ~D[45] /*14701*/;
assign _49507_ = _48813_ & _49510_ /*14697*/;
assign _49508_ = _48813_ ^ _49510_ /*14700*/;
assign _49509_ = _49501_ & _49508_ /*14698*/;
assign _49262_ = _49501_ ^ _49508_ /*14699*/;
assign _49506_ = _49507_ | _49509_ /*14696*/;
assign _49515_ = ~D[46] /*14695*/;
assign _49512_ = _48814_ & _49515_ /*14691*/;
assign _49513_ = _48814_ ^ _49515_ /*14694*/;
assign _49514_ = _49506_ & _49513_ /*14692*/;
assign _49263_ = _49506_ ^ _49513_ /*14693*/;
assign _49511_ = _49512_ | _49514_ /*14690*/;
assign _49520_ = ~D[47] /*14689*/;
assign _49517_ = _48815_ & _49520_ /*14685*/;
assign _49518_ = _48815_ ^ _49520_ /*14688*/;
assign _49519_ = _49511_ & _49518_ /*14686*/;
assign _49264_ = _49511_ ^ _49518_ /*14687*/;
assign _49516_ = _49517_ | _49519_ /*14684*/;
assign _49525_ = ~D[48] /*14683*/;
assign _49522_ = _48816_ & _49525_ /*14679*/;
assign _49523_ = _48816_ ^ _49525_ /*14682*/;
assign _49524_ = _49516_ & _49523_ /*14680*/;
assign _49265_ = _49516_ ^ _49523_ /*14681*/;
assign _49521_ = _49522_ | _49524_ /*14678*/;
assign _49530_ = ~D[49] /*14677*/;
assign _49527_ = _48817_ & _49530_ /*14673*/;
assign _49528_ = _48817_ ^ _49530_ /*14676*/;
assign _49529_ = _49521_ & _49528_ /*14674*/;
assign _49266_ = _49521_ ^ _49528_ /*14675*/;
assign _49526_ = _49527_ | _49529_ /*14672*/;
assign _49535_ = ~D[50] /*14671*/;
assign _49532_ = _48818_ & _49535_ /*14667*/;
assign _49533_ = _48818_ ^ _49535_ /*14670*/;
assign _49534_ = _49526_ & _49533_ /*14668*/;
assign _49267_ = _49526_ ^ _49533_ /*14669*/;
assign _49531_ = _49532_ | _49534_ /*14666*/;
assign _49540_ = ~D[51] /*14665*/;
assign _49537_ = _48819_ & _49540_ /*14661*/;
assign _49538_ = _48819_ ^ _49540_ /*14664*/;
assign _49539_ = _49531_ & _49538_ /*14662*/;
assign _49268_ = _49531_ ^ _49538_ /*14663*/;
assign _49536_ = _49537_ | _49539_ /*14660*/;
assign _49545_ = ~D[52] /*14659*/;
assign _49542_ = _48820_ & _49545_ /*14655*/;
assign _49543_ = _48820_ ^ _49545_ /*14658*/;
assign _49544_ = _49536_ & _49543_ /*14656*/;
assign _49269_ = _49536_ ^ _49543_ /*14657*/;
assign _49541_ = _49542_ | _49544_ /*14654*/;
assign _49550_ = ~D[53] /*14653*/;
assign _49547_ = _48821_ & _49550_ /*14649*/;
assign _49548_ = _48821_ ^ _49550_ /*14652*/;
assign _49549_ = _49541_ & _49548_ /*14650*/;
assign _49270_ = _49541_ ^ _49548_ /*14651*/;
assign _49546_ = _49547_ | _49549_ /*14648*/;
assign _49555_ = ~D[54] /*14647*/;
assign _49552_ = _48822_ & _49555_ /*14643*/;
assign _49553_ = _48822_ ^ _49555_ /*14646*/;
assign _49554_ = _49546_ & _49553_ /*14644*/;
assign _49271_ = _49546_ ^ _49553_ /*14645*/;
assign _49551_ = _49552_ | _49554_ /*14642*/;
assign _49560_ = ~D[55] /*14641*/;
assign _49557_ = _48823_ & _49560_ /*14637*/;
assign _49558_ = _48823_ ^ _49560_ /*14640*/;
assign _49559_ = _49551_ & _49558_ /*14638*/;
assign _49272_ = _49551_ ^ _49558_ /*14639*/;
assign _49556_ = _49557_ | _49559_ /*14636*/;
assign _49565_ = ~D[56] /*14635*/;
assign _49562_ = _48824_ & _49565_ /*14631*/;
assign _49563_ = _48824_ ^ _49565_ /*14634*/;
assign _49564_ = _49556_ & _49563_ /*14632*/;
assign _49273_ = _49556_ ^ _49563_ /*14633*/;
assign _49561_ = _49562_ | _49564_ /*14630*/;
assign _49570_ = ~D[57] /*14629*/;
assign _49567_ = _48825_ & _49570_ /*14625*/;
assign _49568_ = _48825_ ^ _49570_ /*14628*/;
assign _49569_ = _49561_ & _49568_ /*14626*/;
assign _49274_ = _49561_ ^ _49568_ /*14627*/;
assign _49566_ = _49567_ | _49569_ /*14624*/;
assign _49575_ = ~D[58] /*14623*/;
assign _49572_ = _48826_ & _49575_ /*14619*/;
assign _49573_ = _48826_ ^ _49575_ /*14622*/;
assign _49574_ = _49566_ & _49573_ /*14620*/;
assign _49275_ = _49566_ ^ _49573_ /*14621*/;
assign _49571_ = _49572_ | _49574_ /*14618*/;
assign _49580_ = ~D[59] /*14617*/;
assign _49577_ = _48827_ & _49580_ /*14613*/;
assign _49578_ = _48827_ ^ _49580_ /*14616*/;
assign _49579_ = _49571_ & _49578_ /*14614*/;
assign _49276_ = _49571_ ^ _49578_ /*14615*/;
assign _49576_ = _49577_ | _49579_ /*14612*/;
assign _49585_ = ~D[60] /*14611*/;
assign _49582_ = _48828_ & _49585_ /*14607*/;
assign _49583_ = _48828_ ^ _49585_ /*14610*/;
assign _49584_ = _49576_ & _49583_ /*14608*/;
assign _49277_ = _49576_ ^ _49583_ /*14609*/;
assign _49581_ = _49582_ | _49584_ /*14606*/;
assign _49590_ = ~D[61] /*14605*/;
assign _49587_ = _48829_ & _49590_ /*14601*/;
assign _49588_ = _48829_ ^ _49590_ /*14604*/;
assign _49589_ = _49581_ & _49588_ /*14602*/;
assign _49278_ = _49581_ ^ _49588_ /*14603*/;
assign _49586_ = _49587_ | _49589_ /*14600*/;
assign _49595_ = ~D[62] /*14599*/;
assign _49592_ = _48830_ & _49595_ /*14595*/;
assign _49593_ = _48830_ ^ _49595_ /*14598*/;
assign _49594_ = _49586_ & _49593_ /*14596*/;
assign _49279_ = _49586_ ^ _49593_ /*14597*/;
assign _49591_ = _49592_ | _49594_ /*14594*/;
assign _49596_ = _48831_ & oneWire /*14589*/;
assign _49597_ = _48831_ ^ oneWire /*14592*/;
assign _49598_ = _49591_ & _49597_ /*14590*/;
assign _49280_ = _49591_ ^ _49597_ /*14591*/;
assign Q[8] = _49596_ | _49598_ /*14588*/;
assign _49731_ = ~Q[8] /*14203*/;
assign _49730_ = _49731_ & D[0] /*14202*/;
assign _49733_ = _49217_ & _49730_ /*14197*/;
assign _49734_ = _49217_ ^ _49730_ /*14200*/;
assign _49735_ = zeroWire & _49734_ /*14198*/;
assign _49665_ = zeroWire ^ _49734_ /*14199*/;
assign _49732_ = _49733_ | _49735_ /*14196*/;
assign _49737_ = ~Q[8] /*14195*/;
assign _49736_ = _49737_ & D[1] /*14194*/;
assign _49739_ = _49218_ & _49736_ /*14189*/;
assign _49740_ = _49218_ ^ _49736_ /*14192*/;
assign _49741_ = _49732_ & _49740_ /*14190*/;
assign _49666_ = _49732_ ^ _49740_ /*14191*/;
assign _49738_ = _49739_ | _49741_ /*14188*/;
assign _49743_ = ~Q[8] /*14187*/;
assign _49742_ = _49743_ & D[2] /*14186*/;
assign _49745_ = _49219_ & _49742_ /*14181*/;
assign _49746_ = _49219_ ^ _49742_ /*14184*/;
assign _49747_ = _49738_ & _49746_ /*14182*/;
assign _49667_ = _49738_ ^ _49746_ /*14183*/;
assign _49744_ = _49745_ | _49747_ /*14180*/;
assign _49749_ = ~Q[8] /*14179*/;
assign _49748_ = _49749_ & D[3] /*14178*/;
assign _49751_ = _49220_ & _49748_ /*14173*/;
assign _49752_ = _49220_ ^ _49748_ /*14176*/;
assign _49753_ = _49744_ & _49752_ /*14174*/;
assign _49668_ = _49744_ ^ _49752_ /*14175*/;
assign _49750_ = _49751_ | _49753_ /*14172*/;
assign _49755_ = ~Q[8] /*14171*/;
assign _49754_ = _49755_ & D[4] /*14170*/;
assign _49757_ = _49221_ & _49754_ /*14165*/;
assign _49758_ = _49221_ ^ _49754_ /*14168*/;
assign _49759_ = _49750_ & _49758_ /*14166*/;
assign _49669_ = _49750_ ^ _49758_ /*14167*/;
assign _49756_ = _49757_ | _49759_ /*14164*/;
assign _49761_ = ~Q[8] /*14163*/;
assign _49760_ = _49761_ & D[5] /*14162*/;
assign _49763_ = _49222_ & _49760_ /*14157*/;
assign _49764_ = _49222_ ^ _49760_ /*14160*/;
assign _49765_ = _49756_ & _49764_ /*14158*/;
assign _49670_ = _49756_ ^ _49764_ /*14159*/;
assign _49762_ = _49763_ | _49765_ /*14156*/;
assign _49767_ = ~Q[8] /*14155*/;
assign _49766_ = _49767_ & D[6] /*14154*/;
assign _49769_ = _49223_ & _49766_ /*14149*/;
assign _49770_ = _49223_ ^ _49766_ /*14152*/;
assign _49771_ = _49762_ & _49770_ /*14150*/;
assign _49671_ = _49762_ ^ _49770_ /*14151*/;
assign _49768_ = _49769_ | _49771_ /*14148*/;
assign _49773_ = ~Q[8] /*14147*/;
assign _49772_ = _49773_ & D[7] /*14146*/;
assign _49775_ = _49224_ & _49772_ /*14141*/;
assign _49776_ = _49224_ ^ _49772_ /*14144*/;
assign _49777_ = _49768_ & _49776_ /*14142*/;
assign _49672_ = _49768_ ^ _49776_ /*14143*/;
assign _49774_ = _49775_ | _49777_ /*14140*/;
assign _49779_ = ~Q[8] /*14139*/;
assign _49778_ = _49779_ & D[8] /*14138*/;
assign _49781_ = _49225_ & _49778_ /*14133*/;
assign _49782_ = _49225_ ^ _49778_ /*14136*/;
assign _49783_ = _49774_ & _49782_ /*14134*/;
assign _49673_ = _49774_ ^ _49782_ /*14135*/;
assign _49780_ = _49781_ | _49783_ /*14132*/;
assign _49785_ = ~Q[8] /*14131*/;
assign _49784_ = _49785_ & D[9] /*14130*/;
assign _49787_ = _49226_ & _49784_ /*14125*/;
assign _49788_ = _49226_ ^ _49784_ /*14128*/;
assign _49789_ = _49780_ & _49788_ /*14126*/;
assign _49674_ = _49780_ ^ _49788_ /*14127*/;
assign _49786_ = _49787_ | _49789_ /*14124*/;
assign _49791_ = ~Q[8] /*14123*/;
assign _49790_ = _49791_ & D[10] /*14122*/;
assign _49793_ = _49227_ & _49790_ /*14117*/;
assign _49794_ = _49227_ ^ _49790_ /*14120*/;
assign _49795_ = _49786_ & _49794_ /*14118*/;
assign _49675_ = _49786_ ^ _49794_ /*14119*/;
assign _49792_ = _49793_ | _49795_ /*14116*/;
assign _49797_ = ~Q[8] /*14115*/;
assign _49796_ = _49797_ & D[11] /*14114*/;
assign _49799_ = _49228_ & _49796_ /*14109*/;
assign _49800_ = _49228_ ^ _49796_ /*14112*/;
assign _49801_ = _49792_ & _49800_ /*14110*/;
assign _49676_ = _49792_ ^ _49800_ /*14111*/;
assign _49798_ = _49799_ | _49801_ /*14108*/;
assign _49803_ = ~Q[8] /*14107*/;
assign _49802_ = _49803_ & D[12] /*14106*/;
assign _49805_ = _49229_ & _49802_ /*14101*/;
assign _49806_ = _49229_ ^ _49802_ /*14104*/;
assign _49807_ = _49798_ & _49806_ /*14102*/;
assign _49677_ = _49798_ ^ _49806_ /*14103*/;
assign _49804_ = _49805_ | _49807_ /*14100*/;
assign _49809_ = ~Q[8] /*14099*/;
assign _49808_ = _49809_ & D[13] /*14098*/;
assign _49811_ = _49230_ & _49808_ /*14093*/;
assign _49812_ = _49230_ ^ _49808_ /*14096*/;
assign _49813_ = _49804_ & _49812_ /*14094*/;
assign _49678_ = _49804_ ^ _49812_ /*14095*/;
assign _49810_ = _49811_ | _49813_ /*14092*/;
assign _49815_ = ~Q[8] /*14091*/;
assign _49814_ = _49815_ & D[14] /*14090*/;
assign _49817_ = _49231_ & _49814_ /*14085*/;
assign _49818_ = _49231_ ^ _49814_ /*14088*/;
assign _49819_ = _49810_ & _49818_ /*14086*/;
assign _49679_ = _49810_ ^ _49818_ /*14087*/;
assign _49816_ = _49817_ | _49819_ /*14084*/;
assign _49821_ = ~Q[8] /*14083*/;
assign _49820_ = _49821_ & D[15] /*14082*/;
assign _49823_ = _49232_ & _49820_ /*14077*/;
assign _49824_ = _49232_ ^ _49820_ /*14080*/;
assign _49825_ = _49816_ & _49824_ /*14078*/;
assign _49680_ = _49816_ ^ _49824_ /*14079*/;
assign _49822_ = _49823_ | _49825_ /*14076*/;
assign _49827_ = ~Q[8] /*14075*/;
assign _49826_ = _49827_ & D[16] /*14074*/;
assign _49829_ = _49233_ & _49826_ /*14069*/;
assign _49830_ = _49233_ ^ _49826_ /*14072*/;
assign _49831_ = _49822_ & _49830_ /*14070*/;
assign _49681_ = _49822_ ^ _49830_ /*14071*/;
assign _49828_ = _49829_ | _49831_ /*14068*/;
assign _49833_ = ~Q[8] /*14067*/;
assign _49832_ = _49833_ & D[17] /*14066*/;
assign _49835_ = _49234_ & _49832_ /*14061*/;
assign _49836_ = _49234_ ^ _49832_ /*14064*/;
assign _49837_ = _49828_ & _49836_ /*14062*/;
assign _49682_ = _49828_ ^ _49836_ /*14063*/;
assign _49834_ = _49835_ | _49837_ /*14060*/;
assign _49839_ = ~Q[8] /*14059*/;
assign _49838_ = _49839_ & D[18] /*14058*/;
assign _49841_ = _49235_ & _49838_ /*14053*/;
assign _49842_ = _49235_ ^ _49838_ /*14056*/;
assign _49843_ = _49834_ & _49842_ /*14054*/;
assign _49683_ = _49834_ ^ _49842_ /*14055*/;
assign _49840_ = _49841_ | _49843_ /*14052*/;
assign _49845_ = ~Q[8] /*14051*/;
assign _49844_ = _49845_ & D[19] /*14050*/;
assign _49847_ = _49236_ & _49844_ /*14045*/;
assign _49848_ = _49236_ ^ _49844_ /*14048*/;
assign _49849_ = _49840_ & _49848_ /*14046*/;
assign _49684_ = _49840_ ^ _49848_ /*14047*/;
assign _49846_ = _49847_ | _49849_ /*14044*/;
assign _49851_ = ~Q[8] /*14043*/;
assign _49850_ = _49851_ & D[20] /*14042*/;
assign _49853_ = _49237_ & _49850_ /*14037*/;
assign _49854_ = _49237_ ^ _49850_ /*14040*/;
assign _49855_ = _49846_ & _49854_ /*14038*/;
assign _49685_ = _49846_ ^ _49854_ /*14039*/;
assign _49852_ = _49853_ | _49855_ /*14036*/;
assign _49857_ = ~Q[8] /*14035*/;
assign _49856_ = _49857_ & D[21] /*14034*/;
assign _49859_ = _49238_ & _49856_ /*14029*/;
assign _49860_ = _49238_ ^ _49856_ /*14032*/;
assign _49861_ = _49852_ & _49860_ /*14030*/;
assign _49686_ = _49852_ ^ _49860_ /*14031*/;
assign _49858_ = _49859_ | _49861_ /*14028*/;
assign _49863_ = ~Q[8] /*14027*/;
assign _49862_ = _49863_ & D[22] /*14026*/;
assign _49865_ = _49239_ & _49862_ /*14021*/;
assign _49866_ = _49239_ ^ _49862_ /*14024*/;
assign _49867_ = _49858_ & _49866_ /*14022*/;
assign _49687_ = _49858_ ^ _49866_ /*14023*/;
assign _49864_ = _49865_ | _49867_ /*14020*/;
assign _49869_ = ~Q[8] /*14019*/;
assign _49868_ = _49869_ & D[23] /*14018*/;
assign _49871_ = _49240_ & _49868_ /*14013*/;
assign _49872_ = _49240_ ^ _49868_ /*14016*/;
assign _49873_ = _49864_ & _49872_ /*14014*/;
assign _49688_ = _49864_ ^ _49872_ /*14015*/;
assign _49870_ = _49871_ | _49873_ /*14012*/;
assign _49875_ = ~Q[8] /*14011*/;
assign _49874_ = _49875_ & D[24] /*14010*/;
assign _49877_ = _49241_ & _49874_ /*14005*/;
assign _49878_ = _49241_ ^ _49874_ /*14008*/;
assign _49879_ = _49870_ & _49878_ /*14006*/;
assign _49689_ = _49870_ ^ _49878_ /*14007*/;
assign _49876_ = _49877_ | _49879_ /*14004*/;
assign _49881_ = ~Q[8] /*14003*/;
assign _49880_ = _49881_ & D[25] /*14002*/;
assign _49883_ = _49242_ & _49880_ /*13997*/;
assign _49884_ = _49242_ ^ _49880_ /*14000*/;
assign _49885_ = _49876_ & _49884_ /*13998*/;
assign _49690_ = _49876_ ^ _49884_ /*13999*/;
assign _49882_ = _49883_ | _49885_ /*13996*/;
assign _49887_ = ~Q[8] /*13995*/;
assign _49886_ = _49887_ & D[26] /*13994*/;
assign _49889_ = _49243_ & _49886_ /*13989*/;
assign _49890_ = _49243_ ^ _49886_ /*13992*/;
assign _49891_ = _49882_ & _49890_ /*13990*/;
assign _49691_ = _49882_ ^ _49890_ /*13991*/;
assign _49888_ = _49889_ | _49891_ /*13988*/;
assign _49893_ = ~Q[8] /*13987*/;
assign _49892_ = _49893_ & D[27] /*13986*/;
assign _49895_ = _49244_ & _49892_ /*13981*/;
assign _49896_ = _49244_ ^ _49892_ /*13984*/;
assign _49897_ = _49888_ & _49896_ /*13982*/;
assign _49692_ = _49888_ ^ _49896_ /*13983*/;
assign _49894_ = _49895_ | _49897_ /*13980*/;
assign _49899_ = ~Q[8] /*13979*/;
assign _49898_ = _49899_ & D[28] /*13978*/;
assign _49901_ = _49245_ & _49898_ /*13973*/;
assign _49902_ = _49245_ ^ _49898_ /*13976*/;
assign _49903_ = _49894_ & _49902_ /*13974*/;
assign _49693_ = _49894_ ^ _49902_ /*13975*/;
assign _49900_ = _49901_ | _49903_ /*13972*/;
assign _49905_ = ~Q[8] /*13971*/;
assign _49904_ = _49905_ & D[29] /*13970*/;
assign _49907_ = _49246_ & _49904_ /*13965*/;
assign _49908_ = _49246_ ^ _49904_ /*13968*/;
assign _49909_ = _49900_ & _49908_ /*13966*/;
assign _49694_ = _49900_ ^ _49908_ /*13967*/;
assign _49906_ = _49907_ | _49909_ /*13964*/;
assign _49911_ = ~Q[8] /*13963*/;
assign _49910_ = _49911_ & D[30] /*13962*/;
assign _49913_ = _49247_ & _49910_ /*13957*/;
assign _49914_ = _49247_ ^ _49910_ /*13960*/;
assign _49915_ = _49906_ & _49914_ /*13958*/;
assign _49695_ = _49906_ ^ _49914_ /*13959*/;
assign _49912_ = _49913_ | _49915_ /*13956*/;
assign _49917_ = ~Q[8] /*13955*/;
assign _49916_ = _49917_ & D[31] /*13954*/;
assign _49919_ = _49248_ & _49916_ /*13949*/;
assign _49920_ = _49248_ ^ _49916_ /*13952*/;
assign _49921_ = _49912_ & _49920_ /*13950*/;
assign _49696_ = _49912_ ^ _49920_ /*13951*/;
assign _49918_ = _49919_ | _49921_ /*13948*/;
assign _49923_ = ~Q[8] /*13947*/;
assign _49922_ = _49923_ & D[32] /*13946*/;
assign _49925_ = _49249_ & _49922_ /*13941*/;
assign _49926_ = _49249_ ^ _49922_ /*13944*/;
assign _49927_ = _49918_ & _49926_ /*13942*/;
assign _49697_ = _49918_ ^ _49926_ /*13943*/;
assign _49924_ = _49925_ | _49927_ /*13940*/;
assign _49929_ = ~Q[8] /*13939*/;
assign _49928_ = _49929_ & D[33] /*13938*/;
assign _49931_ = _49250_ & _49928_ /*13933*/;
assign _49932_ = _49250_ ^ _49928_ /*13936*/;
assign _49933_ = _49924_ & _49932_ /*13934*/;
assign _49698_ = _49924_ ^ _49932_ /*13935*/;
assign _49930_ = _49931_ | _49933_ /*13932*/;
assign _49935_ = ~Q[8] /*13931*/;
assign _49934_ = _49935_ & D[34] /*13930*/;
assign _49937_ = _49251_ & _49934_ /*13925*/;
assign _49938_ = _49251_ ^ _49934_ /*13928*/;
assign _49939_ = _49930_ & _49938_ /*13926*/;
assign _49699_ = _49930_ ^ _49938_ /*13927*/;
assign _49936_ = _49937_ | _49939_ /*13924*/;
assign _49941_ = ~Q[8] /*13923*/;
assign _49940_ = _49941_ & D[35] /*13922*/;
assign _49943_ = _49252_ & _49940_ /*13917*/;
assign _49944_ = _49252_ ^ _49940_ /*13920*/;
assign _49945_ = _49936_ & _49944_ /*13918*/;
assign _49700_ = _49936_ ^ _49944_ /*13919*/;
assign _49942_ = _49943_ | _49945_ /*13916*/;
assign _49947_ = ~Q[8] /*13915*/;
assign _49946_ = _49947_ & D[36] /*13914*/;
assign _49949_ = _49253_ & _49946_ /*13909*/;
assign _49950_ = _49253_ ^ _49946_ /*13912*/;
assign _49951_ = _49942_ & _49950_ /*13910*/;
assign _49701_ = _49942_ ^ _49950_ /*13911*/;
assign _49948_ = _49949_ | _49951_ /*13908*/;
assign _49953_ = ~Q[8] /*13907*/;
assign _49952_ = _49953_ & D[37] /*13906*/;
assign _49955_ = _49254_ & _49952_ /*13901*/;
assign _49956_ = _49254_ ^ _49952_ /*13904*/;
assign _49957_ = _49948_ & _49956_ /*13902*/;
assign _49702_ = _49948_ ^ _49956_ /*13903*/;
assign _49954_ = _49955_ | _49957_ /*13900*/;
assign _49959_ = ~Q[8] /*13899*/;
assign _49958_ = _49959_ & D[38] /*13898*/;
assign _49961_ = _49255_ & _49958_ /*13893*/;
assign _49962_ = _49255_ ^ _49958_ /*13896*/;
assign _49963_ = _49954_ & _49962_ /*13894*/;
assign _49703_ = _49954_ ^ _49962_ /*13895*/;
assign _49960_ = _49961_ | _49963_ /*13892*/;
assign _49965_ = ~Q[8] /*13891*/;
assign _49964_ = _49965_ & D[39] /*13890*/;
assign _49967_ = _49256_ & _49964_ /*13885*/;
assign _49968_ = _49256_ ^ _49964_ /*13888*/;
assign _49969_ = _49960_ & _49968_ /*13886*/;
assign _49704_ = _49960_ ^ _49968_ /*13887*/;
assign _49966_ = _49967_ | _49969_ /*13884*/;
assign _49971_ = ~Q[8] /*13883*/;
assign _49970_ = _49971_ & D[40] /*13882*/;
assign _49973_ = _49257_ & _49970_ /*13877*/;
assign _49974_ = _49257_ ^ _49970_ /*13880*/;
assign _49975_ = _49966_ & _49974_ /*13878*/;
assign _49705_ = _49966_ ^ _49974_ /*13879*/;
assign _49972_ = _49973_ | _49975_ /*13876*/;
assign _49977_ = ~Q[8] /*13875*/;
assign _49976_ = _49977_ & D[41] /*13874*/;
assign _49979_ = _49258_ & _49976_ /*13869*/;
assign _49980_ = _49258_ ^ _49976_ /*13872*/;
assign _49981_ = _49972_ & _49980_ /*13870*/;
assign _49706_ = _49972_ ^ _49980_ /*13871*/;
assign _49978_ = _49979_ | _49981_ /*13868*/;
assign _49983_ = ~Q[8] /*13867*/;
assign _49982_ = _49983_ & D[42] /*13866*/;
assign _49985_ = _49259_ & _49982_ /*13861*/;
assign _49986_ = _49259_ ^ _49982_ /*13864*/;
assign _49987_ = _49978_ & _49986_ /*13862*/;
assign _49707_ = _49978_ ^ _49986_ /*13863*/;
assign _49984_ = _49985_ | _49987_ /*13860*/;
assign _49989_ = ~Q[8] /*13859*/;
assign _49988_ = _49989_ & D[43] /*13858*/;
assign _49991_ = _49260_ & _49988_ /*13853*/;
assign _49992_ = _49260_ ^ _49988_ /*13856*/;
assign _49993_ = _49984_ & _49992_ /*13854*/;
assign _49708_ = _49984_ ^ _49992_ /*13855*/;
assign _49990_ = _49991_ | _49993_ /*13852*/;
assign _49995_ = ~Q[8] /*13851*/;
assign _49994_ = _49995_ & D[44] /*13850*/;
assign _49997_ = _49261_ & _49994_ /*13845*/;
assign _49998_ = _49261_ ^ _49994_ /*13848*/;
assign _49999_ = _49990_ & _49998_ /*13846*/;
assign _49709_ = _49990_ ^ _49998_ /*13847*/;
assign _49996_ = _49997_ | _49999_ /*13844*/;
assign _50001_ = ~Q[8] /*13843*/;
assign _50000_ = _50001_ & D[45] /*13842*/;
assign _50003_ = _49262_ & _50000_ /*13837*/;
assign _50004_ = _49262_ ^ _50000_ /*13840*/;
assign _50005_ = _49996_ & _50004_ /*13838*/;
assign _49710_ = _49996_ ^ _50004_ /*13839*/;
assign _50002_ = _50003_ | _50005_ /*13836*/;
assign _50007_ = ~Q[8] /*13835*/;
assign _50006_ = _50007_ & D[46] /*13834*/;
assign _50009_ = _49263_ & _50006_ /*13829*/;
assign _50010_ = _49263_ ^ _50006_ /*13832*/;
assign _50011_ = _50002_ & _50010_ /*13830*/;
assign _49711_ = _50002_ ^ _50010_ /*13831*/;
assign _50008_ = _50009_ | _50011_ /*13828*/;
assign _50013_ = ~Q[8] /*13827*/;
assign _50012_ = _50013_ & D[47] /*13826*/;
assign _50015_ = _49264_ & _50012_ /*13821*/;
assign _50016_ = _49264_ ^ _50012_ /*13824*/;
assign _50017_ = _50008_ & _50016_ /*13822*/;
assign _49712_ = _50008_ ^ _50016_ /*13823*/;
assign _50014_ = _50015_ | _50017_ /*13820*/;
assign _50019_ = ~Q[8] /*13819*/;
assign _50018_ = _50019_ & D[48] /*13818*/;
assign _50021_ = _49265_ & _50018_ /*13813*/;
assign _50022_ = _49265_ ^ _50018_ /*13816*/;
assign _50023_ = _50014_ & _50022_ /*13814*/;
assign _49713_ = _50014_ ^ _50022_ /*13815*/;
assign _50020_ = _50021_ | _50023_ /*13812*/;
assign _50025_ = ~Q[8] /*13811*/;
assign _50024_ = _50025_ & D[49] /*13810*/;
assign _50027_ = _49266_ & _50024_ /*13805*/;
assign _50028_ = _49266_ ^ _50024_ /*13808*/;
assign _50029_ = _50020_ & _50028_ /*13806*/;
assign _49714_ = _50020_ ^ _50028_ /*13807*/;
assign _50026_ = _50027_ | _50029_ /*13804*/;
assign _50031_ = ~Q[8] /*13803*/;
assign _50030_ = _50031_ & D[50] /*13802*/;
assign _50033_ = _49267_ & _50030_ /*13797*/;
assign _50034_ = _49267_ ^ _50030_ /*13800*/;
assign _50035_ = _50026_ & _50034_ /*13798*/;
assign _49715_ = _50026_ ^ _50034_ /*13799*/;
assign _50032_ = _50033_ | _50035_ /*13796*/;
assign _50037_ = ~Q[8] /*13795*/;
assign _50036_ = _50037_ & D[51] /*13794*/;
assign _50039_ = _49268_ & _50036_ /*13789*/;
assign _50040_ = _49268_ ^ _50036_ /*13792*/;
assign _50041_ = _50032_ & _50040_ /*13790*/;
assign _49716_ = _50032_ ^ _50040_ /*13791*/;
assign _50038_ = _50039_ | _50041_ /*13788*/;
assign _50043_ = ~Q[8] /*13787*/;
assign _50042_ = _50043_ & D[52] /*13786*/;
assign _50045_ = _49269_ & _50042_ /*13781*/;
assign _50046_ = _49269_ ^ _50042_ /*13784*/;
assign _50047_ = _50038_ & _50046_ /*13782*/;
assign _49717_ = _50038_ ^ _50046_ /*13783*/;
assign _50044_ = _50045_ | _50047_ /*13780*/;
assign _50049_ = ~Q[8] /*13779*/;
assign _50048_ = _50049_ & D[53] /*13778*/;
assign _50051_ = _49270_ & _50048_ /*13773*/;
assign _50052_ = _49270_ ^ _50048_ /*13776*/;
assign _50053_ = _50044_ & _50052_ /*13774*/;
assign _49718_ = _50044_ ^ _50052_ /*13775*/;
assign _50050_ = _50051_ | _50053_ /*13772*/;
assign _50055_ = ~Q[8] /*13771*/;
assign _50054_ = _50055_ & D[54] /*13770*/;
assign _50057_ = _49271_ & _50054_ /*13765*/;
assign _50058_ = _49271_ ^ _50054_ /*13768*/;
assign _50059_ = _50050_ & _50058_ /*13766*/;
assign _49719_ = _50050_ ^ _50058_ /*13767*/;
assign _50056_ = _50057_ | _50059_ /*13764*/;
assign _50061_ = ~Q[8] /*13763*/;
assign _50060_ = _50061_ & D[55] /*13762*/;
assign _50063_ = _49272_ & _50060_ /*13757*/;
assign _50064_ = _49272_ ^ _50060_ /*13760*/;
assign _50065_ = _50056_ & _50064_ /*13758*/;
assign _49720_ = _50056_ ^ _50064_ /*13759*/;
assign _50062_ = _50063_ | _50065_ /*13756*/;
assign _50067_ = ~Q[8] /*13755*/;
assign _50066_ = _50067_ & D[56] /*13754*/;
assign _50069_ = _49273_ & _50066_ /*13749*/;
assign _50070_ = _49273_ ^ _50066_ /*13752*/;
assign _50071_ = _50062_ & _50070_ /*13750*/;
assign _49721_ = _50062_ ^ _50070_ /*13751*/;
assign _50068_ = _50069_ | _50071_ /*13748*/;
assign _50073_ = ~Q[8] /*13747*/;
assign _50072_ = _50073_ & D[57] /*13746*/;
assign _50075_ = _49274_ & _50072_ /*13741*/;
assign _50076_ = _49274_ ^ _50072_ /*13744*/;
assign _50077_ = _50068_ & _50076_ /*13742*/;
assign _49722_ = _50068_ ^ _50076_ /*13743*/;
assign _50074_ = _50075_ | _50077_ /*13740*/;
assign _50079_ = ~Q[8] /*13739*/;
assign _50078_ = _50079_ & D[58] /*13738*/;
assign _50081_ = _49275_ & _50078_ /*13733*/;
assign _50082_ = _49275_ ^ _50078_ /*13736*/;
assign _50083_ = _50074_ & _50082_ /*13734*/;
assign _49723_ = _50074_ ^ _50082_ /*13735*/;
assign _50080_ = _50081_ | _50083_ /*13732*/;
assign _50085_ = ~Q[8] /*13731*/;
assign _50084_ = _50085_ & D[59] /*13730*/;
assign _50087_ = _49276_ & _50084_ /*13725*/;
assign _50088_ = _49276_ ^ _50084_ /*13728*/;
assign _50089_ = _50080_ & _50088_ /*13726*/;
assign _49724_ = _50080_ ^ _50088_ /*13727*/;
assign _50086_ = _50087_ | _50089_ /*13724*/;
assign _50091_ = ~Q[8] /*13723*/;
assign _50090_ = _50091_ & D[60] /*13722*/;
assign _50093_ = _49277_ & _50090_ /*13717*/;
assign _50094_ = _49277_ ^ _50090_ /*13720*/;
assign _50095_ = _50086_ & _50094_ /*13718*/;
assign _49725_ = _50086_ ^ _50094_ /*13719*/;
assign _50092_ = _50093_ | _50095_ /*13716*/;
assign _50097_ = ~Q[8] /*13715*/;
assign _50096_ = _50097_ & D[61] /*13714*/;
assign _50099_ = _49278_ & _50096_ /*13709*/;
assign _50100_ = _49278_ ^ _50096_ /*13712*/;
assign _50101_ = _50092_ & _50100_ /*13710*/;
assign _49726_ = _50092_ ^ _50100_ /*13711*/;
assign _50098_ = _50099_ | _50101_ /*13708*/;
assign _50103_ = ~Q[8] /*13707*/;
assign _50102_ = _50103_ & D[62] /*13706*/;
assign _50105_ = _49279_ & _50102_ /*13701*/;
assign _50106_ = _49279_ ^ _50102_ /*13704*/;
assign _50107_ = _50098_ & _50106_ /*13702*/;
assign _49727_ = _50098_ ^ _50106_ /*13703*/;
assign _50104_ = _50105_ | _50107_ /*13700*/;
assign _50109_ = ~Q[8] /*13699*/;
assign _50108_ = _50109_ & zeroWire /*13698*/;
assign _50110_ = _49280_ ^ _50108_ /*13696*/;
assign _49728_ = _50110_ ^ _50104_ /*13695*/;
assign _50181_ = ~D[0] /*13441*/;
assign _50178_ = R_0[7] & _50181_ /*13437*/;
assign _50179_ = R_0[7] ^ _50181_ /*13440*/;
assign _50180_ = oneWire & _50179_ /*13438*/;
assign _50113_ = oneWire ^ _50179_ /*13439*/;
assign _50177_ = _50178_ | _50180_ /*13436*/;
assign _50186_ = ~D[1] /*13435*/;
assign _50183_ = _49665_ & _50186_ /*13431*/;
assign _50184_ = _49665_ ^ _50186_ /*13434*/;
assign _50185_ = _50177_ & _50184_ /*13432*/;
assign _50114_ = _50177_ ^ _50184_ /*13433*/;
assign _50182_ = _50183_ | _50185_ /*13430*/;
assign _50191_ = ~D[2] /*13429*/;
assign _50188_ = _49666_ & _50191_ /*13425*/;
assign _50189_ = _49666_ ^ _50191_ /*13428*/;
assign _50190_ = _50182_ & _50189_ /*13426*/;
assign _50115_ = _50182_ ^ _50189_ /*13427*/;
assign _50187_ = _50188_ | _50190_ /*13424*/;
assign _50196_ = ~D[3] /*13423*/;
assign _50193_ = _49667_ & _50196_ /*13419*/;
assign _50194_ = _49667_ ^ _50196_ /*13422*/;
assign _50195_ = _50187_ & _50194_ /*13420*/;
assign _50116_ = _50187_ ^ _50194_ /*13421*/;
assign _50192_ = _50193_ | _50195_ /*13418*/;
assign _50201_ = ~D[4] /*13417*/;
assign _50198_ = _49668_ & _50201_ /*13413*/;
assign _50199_ = _49668_ ^ _50201_ /*13416*/;
assign _50200_ = _50192_ & _50199_ /*13414*/;
assign _50117_ = _50192_ ^ _50199_ /*13415*/;
assign _50197_ = _50198_ | _50200_ /*13412*/;
assign _50206_ = ~D[5] /*13411*/;
assign _50203_ = _49669_ & _50206_ /*13407*/;
assign _50204_ = _49669_ ^ _50206_ /*13410*/;
assign _50205_ = _50197_ & _50204_ /*13408*/;
assign _50118_ = _50197_ ^ _50204_ /*13409*/;
assign _50202_ = _50203_ | _50205_ /*13406*/;
assign _50211_ = ~D[6] /*13405*/;
assign _50208_ = _49670_ & _50211_ /*13401*/;
assign _50209_ = _49670_ ^ _50211_ /*13404*/;
assign _50210_ = _50202_ & _50209_ /*13402*/;
assign _50119_ = _50202_ ^ _50209_ /*13403*/;
assign _50207_ = _50208_ | _50210_ /*13400*/;
assign _50216_ = ~D[7] /*13399*/;
assign _50213_ = _49671_ & _50216_ /*13395*/;
assign _50214_ = _49671_ ^ _50216_ /*13398*/;
assign _50215_ = _50207_ & _50214_ /*13396*/;
assign _50120_ = _50207_ ^ _50214_ /*13397*/;
assign _50212_ = _50213_ | _50215_ /*13394*/;
assign _50221_ = ~D[8] /*13393*/;
assign _50218_ = _49672_ & _50221_ /*13389*/;
assign _50219_ = _49672_ ^ _50221_ /*13392*/;
assign _50220_ = _50212_ & _50219_ /*13390*/;
assign _50121_ = _50212_ ^ _50219_ /*13391*/;
assign _50217_ = _50218_ | _50220_ /*13388*/;
assign _50226_ = ~D[9] /*13387*/;
assign _50223_ = _49673_ & _50226_ /*13383*/;
assign _50224_ = _49673_ ^ _50226_ /*13386*/;
assign _50225_ = _50217_ & _50224_ /*13384*/;
assign _50122_ = _50217_ ^ _50224_ /*13385*/;
assign _50222_ = _50223_ | _50225_ /*13382*/;
assign _50231_ = ~D[10] /*13381*/;
assign _50228_ = _49674_ & _50231_ /*13377*/;
assign _50229_ = _49674_ ^ _50231_ /*13380*/;
assign _50230_ = _50222_ & _50229_ /*13378*/;
assign _50123_ = _50222_ ^ _50229_ /*13379*/;
assign _50227_ = _50228_ | _50230_ /*13376*/;
assign _50236_ = ~D[11] /*13375*/;
assign _50233_ = _49675_ & _50236_ /*13371*/;
assign _50234_ = _49675_ ^ _50236_ /*13374*/;
assign _50235_ = _50227_ & _50234_ /*13372*/;
assign _50124_ = _50227_ ^ _50234_ /*13373*/;
assign _50232_ = _50233_ | _50235_ /*13370*/;
assign _50241_ = ~D[12] /*13369*/;
assign _50238_ = _49676_ & _50241_ /*13365*/;
assign _50239_ = _49676_ ^ _50241_ /*13368*/;
assign _50240_ = _50232_ & _50239_ /*13366*/;
assign _50125_ = _50232_ ^ _50239_ /*13367*/;
assign _50237_ = _50238_ | _50240_ /*13364*/;
assign _50246_ = ~D[13] /*13363*/;
assign _50243_ = _49677_ & _50246_ /*13359*/;
assign _50244_ = _49677_ ^ _50246_ /*13362*/;
assign _50245_ = _50237_ & _50244_ /*13360*/;
assign _50126_ = _50237_ ^ _50244_ /*13361*/;
assign _50242_ = _50243_ | _50245_ /*13358*/;
assign _50251_ = ~D[14] /*13357*/;
assign _50248_ = _49678_ & _50251_ /*13353*/;
assign _50249_ = _49678_ ^ _50251_ /*13356*/;
assign _50250_ = _50242_ & _50249_ /*13354*/;
assign _50127_ = _50242_ ^ _50249_ /*13355*/;
assign _50247_ = _50248_ | _50250_ /*13352*/;
assign _50256_ = ~D[15] /*13351*/;
assign _50253_ = _49679_ & _50256_ /*13347*/;
assign _50254_ = _49679_ ^ _50256_ /*13350*/;
assign _50255_ = _50247_ & _50254_ /*13348*/;
assign _50128_ = _50247_ ^ _50254_ /*13349*/;
assign _50252_ = _50253_ | _50255_ /*13346*/;
assign _50261_ = ~D[16] /*13345*/;
assign _50258_ = _49680_ & _50261_ /*13341*/;
assign _50259_ = _49680_ ^ _50261_ /*13344*/;
assign _50260_ = _50252_ & _50259_ /*13342*/;
assign _50129_ = _50252_ ^ _50259_ /*13343*/;
assign _50257_ = _50258_ | _50260_ /*13340*/;
assign _50266_ = ~D[17] /*13339*/;
assign _50263_ = _49681_ & _50266_ /*13335*/;
assign _50264_ = _49681_ ^ _50266_ /*13338*/;
assign _50265_ = _50257_ & _50264_ /*13336*/;
assign _50130_ = _50257_ ^ _50264_ /*13337*/;
assign _50262_ = _50263_ | _50265_ /*13334*/;
assign _50271_ = ~D[18] /*13333*/;
assign _50268_ = _49682_ & _50271_ /*13329*/;
assign _50269_ = _49682_ ^ _50271_ /*13332*/;
assign _50270_ = _50262_ & _50269_ /*13330*/;
assign _50131_ = _50262_ ^ _50269_ /*13331*/;
assign _50267_ = _50268_ | _50270_ /*13328*/;
assign _50276_ = ~D[19] /*13327*/;
assign _50273_ = _49683_ & _50276_ /*13323*/;
assign _50274_ = _49683_ ^ _50276_ /*13326*/;
assign _50275_ = _50267_ & _50274_ /*13324*/;
assign _50132_ = _50267_ ^ _50274_ /*13325*/;
assign _50272_ = _50273_ | _50275_ /*13322*/;
assign _50281_ = ~D[20] /*13321*/;
assign _50278_ = _49684_ & _50281_ /*13317*/;
assign _50279_ = _49684_ ^ _50281_ /*13320*/;
assign _50280_ = _50272_ & _50279_ /*13318*/;
assign _50133_ = _50272_ ^ _50279_ /*13319*/;
assign _50277_ = _50278_ | _50280_ /*13316*/;
assign _50286_ = ~D[21] /*13315*/;
assign _50283_ = _49685_ & _50286_ /*13311*/;
assign _50284_ = _49685_ ^ _50286_ /*13314*/;
assign _50285_ = _50277_ & _50284_ /*13312*/;
assign _50134_ = _50277_ ^ _50284_ /*13313*/;
assign _50282_ = _50283_ | _50285_ /*13310*/;
assign _50291_ = ~D[22] /*13309*/;
assign _50288_ = _49686_ & _50291_ /*13305*/;
assign _50289_ = _49686_ ^ _50291_ /*13308*/;
assign _50290_ = _50282_ & _50289_ /*13306*/;
assign _50135_ = _50282_ ^ _50289_ /*13307*/;
assign _50287_ = _50288_ | _50290_ /*13304*/;
assign _50296_ = ~D[23] /*13303*/;
assign _50293_ = _49687_ & _50296_ /*13299*/;
assign _50294_ = _49687_ ^ _50296_ /*13302*/;
assign _50295_ = _50287_ & _50294_ /*13300*/;
assign _50136_ = _50287_ ^ _50294_ /*13301*/;
assign _50292_ = _50293_ | _50295_ /*13298*/;
assign _50301_ = ~D[24] /*13297*/;
assign _50298_ = _49688_ & _50301_ /*13293*/;
assign _50299_ = _49688_ ^ _50301_ /*13296*/;
assign _50300_ = _50292_ & _50299_ /*13294*/;
assign _50137_ = _50292_ ^ _50299_ /*13295*/;
assign _50297_ = _50298_ | _50300_ /*13292*/;
assign _50306_ = ~D[25] /*13291*/;
assign _50303_ = _49689_ & _50306_ /*13287*/;
assign _50304_ = _49689_ ^ _50306_ /*13290*/;
assign _50305_ = _50297_ & _50304_ /*13288*/;
assign _50138_ = _50297_ ^ _50304_ /*13289*/;
assign _50302_ = _50303_ | _50305_ /*13286*/;
assign _50311_ = ~D[26] /*13285*/;
assign _50308_ = _49690_ & _50311_ /*13281*/;
assign _50309_ = _49690_ ^ _50311_ /*13284*/;
assign _50310_ = _50302_ & _50309_ /*13282*/;
assign _50139_ = _50302_ ^ _50309_ /*13283*/;
assign _50307_ = _50308_ | _50310_ /*13280*/;
assign _50316_ = ~D[27] /*13279*/;
assign _50313_ = _49691_ & _50316_ /*13275*/;
assign _50314_ = _49691_ ^ _50316_ /*13278*/;
assign _50315_ = _50307_ & _50314_ /*13276*/;
assign _50140_ = _50307_ ^ _50314_ /*13277*/;
assign _50312_ = _50313_ | _50315_ /*13274*/;
assign _50321_ = ~D[28] /*13273*/;
assign _50318_ = _49692_ & _50321_ /*13269*/;
assign _50319_ = _49692_ ^ _50321_ /*13272*/;
assign _50320_ = _50312_ & _50319_ /*13270*/;
assign _50141_ = _50312_ ^ _50319_ /*13271*/;
assign _50317_ = _50318_ | _50320_ /*13268*/;
assign _50326_ = ~D[29] /*13267*/;
assign _50323_ = _49693_ & _50326_ /*13263*/;
assign _50324_ = _49693_ ^ _50326_ /*13266*/;
assign _50325_ = _50317_ & _50324_ /*13264*/;
assign _50142_ = _50317_ ^ _50324_ /*13265*/;
assign _50322_ = _50323_ | _50325_ /*13262*/;
assign _50331_ = ~D[30] /*13261*/;
assign _50328_ = _49694_ & _50331_ /*13257*/;
assign _50329_ = _49694_ ^ _50331_ /*13260*/;
assign _50330_ = _50322_ & _50329_ /*13258*/;
assign _50143_ = _50322_ ^ _50329_ /*13259*/;
assign _50327_ = _50328_ | _50330_ /*13256*/;
assign _50336_ = ~D[31] /*13255*/;
assign _50333_ = _49695_ & _50336_ /*13251*/;
assign _50334_ = _49695_ ^ _50336_ /*13254*/;
assign _50335_ = _50327_ & _50334_ /*13252*/;
assign _50144_ = _50327_ ^ _50334_ /*13253*/;
assign _50332_ = _50333_ | _50335_ /*13250*/;
assign _50341_ = ~D[32] /*13249*/;
assign _50338_ = _49696_ & _50341_ /*13245*/;
assign _50339_ = _49696_ ^ _50341_ /*13248*/;
assign _50340_ = _50332_ & _50339_ /*13246*/;
assign _50145_ = _50332_ ^ _50339_ /*13247*/;
assign _50337_ = _50338_ | _50340_ /*13244*/;
assign _50346_ = ~D[33] /*13243*/;
assign _50343_ = _49697_ & _50346_ /*13239*/;
assign _50344_ = _49697_ ^ _50346_ /*13242*/;
assign _50345_ = _50337_ & _50344_ /*13240*/;
assign _50146_ = _50337_ ^ _50344_ /*13241*/;
assign _50342_ = _50343_ | _50345_ /*13238*/;
assign _50351_ = ~D[34] /*13237*/;
assign _50348_ = _49698_ & _50351_ /*13233*/;
assign _50349_ = _49698_ ^ _50351_ /*13236*/;
assign _50350_ = _50342_ & _50349_ /*13234*/;
assign _50147_ = _50342_ ^ _50349_ /*13235*/;
assign _50347_ = _50348_ | _50350_ /*13232*/;
assign _50356_ = ~D[35] /*13231*/;
assign _50353_ = _49699_ & _50356_ /*13227*/;
assign _50354_ = _49699_ ^ _50356_ /*13230*/;
assign _50355_ = _50347_ & _50354_ /*13228*/;
assign _50148_ = _50347_ ^ _50354_ /*13229*/;
assign _50352_ = _50353_ | _50355_ /*13226*/;
assign _50361_ = ~D[36] /*13225*/;
assign _50358_ = _49700_ & _50361_ /*13221*/;
assign _50359_ = _49700_ ^ _50361_ /*13224*/;
assign _50360_ = _50352_ & _50359_ /*13222*/;
assign _50149_ = _50352_ ^ _50359_ /*13223*/;
assign _50357_ = _50358_ | _50360_ /*13220*/;
assign _50366_ = ~D[37] /*13219*/;
assign _50363_ = _49701_ & _50366_ /*13215*/;
assign _50364_ = _49701_ ^ _50366_ /*13218*/;
assign _50365_ = _50357_ & _50364_ /*13216*/;
assign _50150_ = _50357_ ^ _50364_ /*13217*/;
assign _50362_ = _50363_ | _50365_ /*13214*/;
assign _50371_ = ~D[38] /*13213*/;
assign _50368_ = _49702_ & _50371_ /*13209*/;
assign _50369_ = _49702_ ^ _50371_ /*13212*/;
assign _50370_ = _50362_ & _50369_ /*13210*/;
assign _50151_ = _50362_ ^ _50369_ /*13211*/;
assign _50367_ = _50368_ | _50370_ /*13208*/;
assign _50376_ = ~D[39] /*13207*/;
assign _50373_ = _49703_ & _50376_ /*13203*/;
assign _50374_ = _49703_ ^ _50376_ /*13206*/;
assign _50375_ = _50367_ & _50374_ /*13204*/;
assign _50152_ = _50367_ ^ _50374_ /*13205*/;
assign _50372_ = _50373_ | _50375_ /*13202*/;
assign _50381_ = ~D[40] /*13201*/;
assign _50378_ = _49704_ & _50381_ /*13197*/;
assign _50379_ = _49704_ ^ _50381_ /*13200*/;
assign _50380_ = _50372_ & _50379_ /*13198*/;
assign _50153_ = _50372_ ^ _50379_ /*13199*/;
assign _50377_ = _50378_ | _50380_ /*13196*/;
assign _50386_ = ~D[41] /*13195*/;
assign _50383_ = _49705_ & _50386_ /*13191*/;
assign _50384_ = _49705_ ^ _50386_ /*13194*/;
assign _50385_ = _50377_ & _50384_ /*13192*/;
assign _50154_ = _50377_ ^ _50384_ /*13193*/;
assign _50382_ = _50383_ | _50385_ /*13190*/;
assign _50391_ = ~D[42] /*13189*/;
assign _50388_ = _49706_ & _50391_ /*13185*/;
assign _50389_ = _49706_ ^ _50391_ /*13188*/;
assign _50390_ = _50382_ & _50389_ /*13186*/;
assign _50155_ = _50382_ ^ _50389_ /*13187*/;
assign _50387_ = _50388_ | _50390_ /*13184*/;
assign _50396_ = ~D[43] /*13183*/;
assign _50393_ = _49707_ & _50396_ /*13179*/;
assign _50394_ = _49707_ ^ _50396_ /*13182*/;
assign _50395_ = _50387_ & _50394_ /*13180*/;
assign _50156_ = _50387_ ^ _50394_ /*13181*/;
assign _50392_ = _50393_ | _50395_ /*13178*/;
assign _50401_ = ~D[44] /*13177*/;
assign _50398_ = _49708_ & _50401_ /*13173*/;
assign _50399_ = _49708_ ^ _50401_ /*13176*/;
assign _50400_ = _50392_ & _50399_ /*13174*/;
assign _50157_ = _50392_ ^ _50399_ /*13175*/;
assign _50397_ = _50398_ | _50400_ /*13172*/;
assign _50406_ = ~D[45] /*13171*/;
assign _50403_ = _49709_ & _50406_ /*13167*/;
assign _50404_ = _49709_ ^ _50406_ /*13170*/;
assign _50405_ = _50397_ & _50404_ /*13168*/;
assign _50158_ = _50397_ ^ _50404_ /*13169*/;
assign _50402_ = _50403_ | _50405_ /*13166*/;
assign _50411_ = ~D[46] /*13165*/;
assign _50408_ = _49710_ & _50411_ /*13161*/;
assign _50409_ = _49710_ ^ _50411_ /*13164*/;
assign _50410_ = _50402_ & _50409_ /*13162*/;
assign _50159_ = _50402_ ^ _50409_ /*13163*/;
assign _50407_ = _50408_ | _50410_ /*13160*/;
assign _50416_ = ~D[47] /*13159*/;
assign _50413_ = _49711_ & _50416_ /*13155*/;
assign _50414_ = _49711_ ^ _50416_ /*13158*/;
assign _50415_ = _50407_ & _50414_ /*13156*/;
assign _50160_ = _50407_ ^ _50414_ /*13157*/;
assign _50412_ = _50413_ | _50415_ /*13154*/;
assign _50421_ = ~D[48] /*13153*/;
assign _50418_ = _49712_ & _50421_ /*13149*/;
assign _50419_ = _49712_ ^ _50421_ /*13152*/;
assign _50420_ = _50412_ & _50419_ /*13150*/;
assign _50161_ = _50412_ ^ _50419_ /*13151*/;
assign _50417_ = _50418_ | _50420_ /*13148*/;
assign _50426_ = ~D[49] /*13147*/;
assign _50423_ = _49713_ & _50426_ /*13143*/;
assign _50424_ = _49713_ ^ _50426_ /*13146*/;
assign _50425_ = _50417_ & _50424_ /*13144*/;
assign _50162_ = _50417_ ^ _50424_ /*13145*/;
assign _50422_ = _50423_ | _50425_ /*13142*/;
assign _50431_ = ~D[50] /*13141*/;
assign _50428_ = _49714_ & _50431_ /*13137*/;
assign _50429_ = _49714_ ^ _50431_ /*13140*/;
assign _50430_ = _50422_ & _50429_ /*13138*/;
assign _50163_ = _50422_ ^ _50429_ /*13139*/;
assign _50427_ = _50428_ | _50430_ /*13136*/;
assign _50436_ = ~D[51] /*13135*/;
assign _50433_ = _49715_ & _50436_ /*13131*/;
assign _50434_ = _49715_ ^ _50436_ /*13134*/;
assign _50435_ = _50427_ & _50434_ /*13132*/;
assign _50164_ = _50427_ ^ _50434_ /*13133*/;
assign _50432_ = _50433_ | _50435_ /*13130*/;
assign _50441_ = ~D[52] /*13129*/;
assign _50438_ = _49716_ & _50441_ /*13125*/;
assign _50439_ = _49716_ ^ _50441_ /*13128*/;
assign _50440_ = _50432_ & _50439_ /*13126*/;
assign _50165_ = _50432_ ^ _50439_ /*13127*/;
assign _50437_ = _50438_ | _50440_ /*13124*/;
assign _50446_ = ~D[53] /*13123*/;
assign _50443_ = _49717_ & _50446_ /*13119*/;
assign _50444_ = _49717_ ^ _50446_ /*13122*/;
assign _50445_ = _50437_ & _50444_ /*13120*/;
assign _50166_ = _50437_ ^ _50444_ /*13121*/;
assign _50442_ = _50443_ | _50445_ /*13118*/;
assign _50451_ = ~D[54] /*13117*/;
assign _50448_ = _49718_ & _50451_ /*13113*/;
assign _50449_ = _49718_ ^ _50451_ /*13116*/;
assign _50450_ = _50442_ & _50449_ /*13114*/;
assign _50167_ = _50442_ ^ _50449_ /*13115*/;
assign _50447_ = _50448_ | _50450_ /*13112*/;
assign _50456_ = ~D[55] /*13111*/;
assign _50453_ = _49719_ & _50456_ /*13107*/;
assign _50454_ = _49719_ ^ _50456_ /*13110*/;
assign _50455_ = _50447_ & _50454_ /*13108*/;
assign _50168_ = _50447_ ^ _50454_ /*13109*/;
assign _50452_ = _50453_ | _50455_ /*13106*/;
assign _50461_ = ~D[56] /*13105*/;
assign _50458_ = _49720_ & _50461_ /*13101*/;
assign _50459_ = _49720_ ^ _50461_ /*13104*/;
assign _50460_ = _50452_ & _50459_ /*13102*/;
assign _50169_ = _50452_ ^ _50459_ /*13103*/;
assign _50457_ = _50458_ | _50460_ /*13100*/;
assign _50466_ = ~D[57] /*13099*/;
assign _50463_ = _49721_ & _50466_ /*13095*/;
assign _50464_ = _49721_ ^ _50466_ /*13098*/;
assign _50465_ = _50457_ & _50464_ /*13096*/;
assign _50170_ = _50457_ ^ _50464_ /*13097*/;
assign _50462_ = _50463_ | _50465_ /*13094*/;
assign _50471_ = ~D[58] /*13093*/;
assign _50468_ = _49722_ & _50471_ /*13089*/;
assign _50469_ = _49722_ ^ _50471_ /*13092*/;
assign _50470_ = _50462_ & _50469_ /*13090*/;
assign _50171_ = _50462_ ^ _50469_ /*13091*/;
assign _50467_ = _50468_ | _50470_ /*13088*/;
assign _50476_ = ~D[59] /*13087*/;
assign _50473_ = _49723_ & _50476_ /*13083*/;
assign _50474_ = _49723_ ^ _50476_ /*13086*/;
assign _50475_ = _50467_ & _50474_ /*13084*/;
assign _50172_ = _50467_ ^ _50474_ /*13085*/;
assign _50472_ = _50473_ | _50475_ /*13082*/;
assign _50481_ = ~D[60] /*13081*/;
assign _50478_ = _49724_ & _50481_ /*13077*/;
assign _50479_ = _49724_ ^ _50481_ /*13080*/;
assign _50480_ = _50472_ & _50479_ /*13078*/;
assign _50173_ = _50472_ ^ _50479_ /*13079*/;
assign _50477_ = _50478_ | _50480_ /*13076*/;
assign _50486_ = ~D[61] /*13075*/;
assign _50483_ = _49725_ & _50486_ /*13071*/;
assign _50484_ = _49725_ ^ _50486_ /*13074*/;
assign _50485_ = _50477_ & _50484_ /*13072*/;
assign _50174_ = _50477_ ^ _50484_ /*13073*/;
assign _50482_ = _50483_ | _50485_ /*13070*/;
assign _50491_ = ~D[62] /*13069*/;
assign _50488_ = _49726_ & _50491_ /*13065*/;
assign _50489_ = _49726_ ^ _50491_ /*13068*/;
assign _50490_ = _50482_ & _50489_ /*13066*/;
assign _50175_ = _50482_ ^ _50489_ /*13067*/;
assign _50487_ = _50488_ | _50490_ /*13064*/;
assign _50492_ = _49727_ & oneWire /*13059*/;
assign _50493_ = _49727_ ^ oneWire /*13062*/;
assign _50494_ = _50487_ & _50493_ /*13060*/;
assign _50176_ = _50487_ ^ _50493_ /*13061*/;
assign Q[7] = _50492_ | _50494_ /*13058*/;
assign _50627_ = ~Q[7] /*12673*/;
assign _50626_ = _50627_ & D[0] /*12672*/;
assign _50629_ = _50113_ & _50626_ /*12667*/;
assign _50630_ = _50113_ ^ _50626_ /*12670*/;
assign _50631_ = zeroWire & _50630_ /*12668*/;
assign _50561_ = zeroWire ^ _50630_ /*12669*/;
assign _50628_ = _50629_ | _50631_ /*12666*/;
assign _50633_ = ~Q[7] /*12665*/;
assign _50632_ = _50633_ & D[1] /*12664*/;
assign _50635_ = _50114_ & _50632_ /*12659*/;
assign _50636_ = _50114_ ^ _50632_ /*12662*/;
assign _50637_ = _50628_ & _50636_ /*12660*/;
assign _50562_ = _50628_ ^ _50636_ /*12661*/;
assign _50634_ = _50635_ | _50637_ /*12658*/;
assign _50639_ = ~Q[7] /*12657*/;
assign _50638_ = _50639_ & D[2] /*12656*/;
assign _50641_ = _50115_ & _50638_ /*12651*/;
assign _50642_ = _50115_ ^ _50638_ /*12654*/;
assign _50643_ = _50634_ & _50642_ /*12652*/;
assign _50563_ = _50634_ ^ _50642_ /*12653*/;
assign _50640_ = _50641_ | _50643_ /*12650*/;
assign _50645_ = ~Q[7] /*12649*/;
assign _50644_ = _50645_ & D[3] /*12648*/;
assign _50647_ = _50116_ & _50644_ /*12643*/;
assign _50648_ = _50116_ ^ _50644_ /*12646*/;
assign _50649_ = _50640_ & _50648_ /*12644*/;
assign _50564_ = _50640_ ^ _50648_ /*12645*/;
assign _50646_ = _50647_ | _50649_ /*12642*/;
assign _50651_ = ~Q[7] /*12641*/;
assign _50650_ = _50651_ & D[4] /*12640*/;
assign _50653_ = _50117_ & _50650_ /*12635*/;
assign _50654_ = _50117_ ^ _50650_ /*12638*/;
assign _50655_ = _50646_ & _50654_ /*12636*/;
assign _50565_ = _50646_ ^ _50654_ /*12637*/;
assign _50652_ = _50653_ | _50655_ /*12634*/;
assign _50657_ = ~Q[7] /*12633*/;
assign _50656_ = _50657_ & D[5] /*12632*/;
assign _50659_ = _50118_ & _50656_ /*12627*/;
assign _50660_ = _50118_ ^ _50656_ /*12630*/;
assign _50661_ = _50652_ & _50660_ /*12628*/;
assign _50566_ = _50652_ ^ _50660_ /*12629*/;
assign _50658_ = _50659_ | _50661_ /*12626*/;
assign _50663_ = ~Q[7] /*12625*/;
assign _50662_ = _50663_ & D[6] /*12624*/;
assign _50665_ = _50119_ & _50662_ /*12619*/;
assign _50666_ = _50119_ ^ _50662_ /*12622*/;
assign _50667_ = _50658_ & _50666_ /*12620*/;
assign _50567_ = _50658_ ^ _50666_ /*12621*/;
assign _50664_ = _50665_ | _50667_ /*12618*/;
assign _50669_ = ~Q[7] /*12617*/;
assign _50668_ = _50669_ & D[7] /*12616*/;
assign _50671_ = _50120_ & _50668_ /*12611*/;
assign _50672_ = _50120_ ^ _50668_ /*12614*/;
assign _50673_ = _50664_ & _50672_ /*12612*/;
assign _50568_ = _50664_ ^ _50672_ /*12613*/;
assign _50670_ = _50671_ | _50673_ /*12610*/;
assign _50675_ = ~Q[7] /*12609*/;
assign _50674_ = _50675_ & D[8] /*12608*/;
assign _50677_ = _50121_ & _50674_ /*12603*/;
assign _50678_ = _50121_ ^ _50674_ /*12606*/;
assign _50679_ = _50670_ & _50678_ /*12604*/;
assign _50569_ = _50670_ ^ _50678_ /*12605*/;
assign _50676_ = _50677_ | _50679_ /*12602*/;
assign _50681_ = ~Q[7] /*12601*/;
assign _50680_ = _50681_ & D[9] /*12600*/;
assign _50683_ = _50122_ & _50680_ /*12595*/;
assign _50684_ = _50122_ ^ _50680_ /*12598*/;
assign _50685_ = _50676_ & _50684_ /*12596*/;
assign _50570_ = _50676_ ^ _50684_ /*12597*/;
assign _50682_ = _50683_ | _50685_ /*12594*/;
assign _50687_ = ~Q[7] /*12593*/;
assign _50686_ = _50687_ & D[10] /*12592*/;
assign _50689_ = _50123_ & _50686_ /*12587*/;
assign _50690_ = _50123_ ^ _50686_ /*12590*/;
assign _50691_ = _50682_ & _50690_ /*12588*/;
assign _50571_ = _50682_ ^ _50690_ /*12589*/;
assign _50688_ = _50689_ | _50691_ /*12586*/;
assign _50693_ = ~Q[7] /*12585*/;
assign _50692_ = _50693_ & D[11] /*12584*/;
assign _50695_ = _50124_ & _50692_ /*12579*/;
assign _50696_ = _50124_ ^ _50692_ /*12582*/;
assign _50697_ = _50688_ & _50696_ /*12580*/;
assign _50572_ = _50688_ ^ _50696_ /*12581*/;
assign _50694_ = _50695_ | _50697_ /*12578*/;
assign _50699_ = ~Q[7] /*12577*/;
assign _50698_ = _50699_ & D[12] /*12576*/;
assign _50701_ = _50125_ & _50698_ /*12571*/;
assign _50702_ = _50125_ ^ _50698_ /*12574*/;
assign _50703_ = _50694_ & _50702_ /*12572*/;
assign _50573_ = _50694_ ^ _50702_ /*12573*/;
assign _50700_ = _50701_ | _50703_ /*12570*/;
assign _50705_ = ~Q[7] /*12569*/;
assign _50704_ = _50705_ & D[13] /*12568*/;
assign _50707_ = _50126_ & _50704_ /*12563*/;
assign _50708_ = _50126_ ^ _50704_ /*12566*/;
assign _50709_ = _50700_ & _50708_ /*12564*/;
assign _50574_ = _50700_ ^ _50708_ /*12565*/;
assign _50706_ = _50707_ | _50709_ /*12562*/;
assign _50711_ = ~Q[7] /*12561*/;
assign _50710_ = _50711_ & D[14] /*12560*/;
assign _50713_ = _50127_ & _50710_ /*12555*/;
assign _50714_ = _50127_ ^ _50710_ /*12558*/;
assign _50715_ = _50706_ & _50714_ /*12556*/;
assign _50575_ = _50706_ ^ _50714_ /*12557*/;
assign _50712_ = _50713_ | _50715_ /*12554*/;
assign _50717_ = ~Q[7] /*12553*/;
assign _50716_ = _50717_ & D[15] /*12552*/;
assign _50719_ = _50128_ & _50716_ /*12547*/;
assign _50720_ = _50128_ ^ _50716_ /*12550*/;
assign _50721_ = _50712_ & _50720_ /*12548*/;
assign _50576_ = _50712_ ^ _50720_ /*12549*/;
assign _50718_ = _50719_ | _50721_ /*12546*/;
assign _50723_ = ~Q[7] /*12545*/;
assign _50722_ = _50723_ & D[16] /*12544*/;
assign _50725_ = _50129_ & _50722_ /*12539*/;
assign _50726_ = _50129_ ^ _50722_ /*12542*/;
assign _50727_ = _50718_ & _50726_ /*12540*/;
assign _50577_ = _50718_ ^ _50726_ /*12541*/;
assign _50724_ = _50725_ | _50727_ /*12538*/;
assign _50729_ = ~Q[7] /*12537*/;
assign _50728_ = _50729_ & D[17] /*12536*/;
assign _50731_ = _50130_ & _50728_ /*12531*/;
assign _50732_ = _50130_ ^ _50728_ /*12534*/;
assign _50733_ = _50724_ & _50732_ /*12532*/;
assign _50578_ = _50724_ ^ _50732_ /*12533*/;
assign _50730_ = _50731_ | _50733_ /*12530*/;
assign _50735_ = ~Q[7] /*12529*/;
assign _50734_ = _50735_ & D[18] /*12528*/;
assign _50737_ = _50131_ & _50734_ /*12523*/;
assign _50738_ = _50131_ ^ _50734_ /*12526*/;
assign _50739_ = _50730_ & _50738_ /*12524*/;
assign _50579_ = _50730_ ^ _50738_ /*12525*/;
assign _50736_ = _50737_ | _50739_ /*12522*/;
assign _50741_ = ~Q[7] /*12521*/;
assign _50740_ = _50741_ & D[19] /*12520*/;
assign _50743_ = _50132_ & _50740_ /*12515*/;
assign _50744_ = _50132_ ^ _50740_ /*12518*/;
assign _50745_ = _50736_ & _50744_ /*12516*/;
assign _50580_ = _50736_ ^ _50744_ /*12517*/;
assign _50742_ = _50743_ | _50745_ /*12514*/;
assign _50747_ = ~Q[7] /*12513*/;
assign _50746_ = _50747_ & D[20] /*12512*/;
assign _50749_ = _50133_ & _50746_ /*12507*/;
assign _50750_ = _50133_ ^ _50746_ /*12510*/;
assign _50751_ = _50742_ & _50750_ /*12508*/;
assign _50581_ = _50742_ ^ _50750_ /*12509*/;
assign _50748_ = _50749_ | _50751_ /*12506*/;
assign _50753_ = ~Q[7] /*12505*/;
assign _50752_ = _50753_ & D[21] /*12504*/;
assign _50755_ = _50134_ & _50752_ /*12499*/;
assign _50756_ = _50134_ ^ _50752_ /*12502*/;
assign _50757_ = _50748_ & _50756_ /*12500*/;
assign _50582_ = _50748_ ^ _50756_ /*12501*/;
assign _50754_ = _50755_ | _50757_ /*12498*/;
assign _50759_ = ~Q[7] /*12497*/;
assign _50758_ = _50759_ & D[22] /*12496*/;
assign _50761_ = _50135_ & _50758_ /*12491*/;
assign _50762_ = _50135_ ^ _50758_ /*12494*/;
assign _50763_ = _50754_ & _50762_ /*12492*/;
assign _50583_ = _50754_ ^ _50762_ /*12493*/;
assign _50760_ = _50761_ | _50763_ /*12490*/;
assign _50765_ = ~Q[7] /*12489*/;
assign _50764_ = _50765_ & D[23] /*12488*/;
assign _50767_ = _50136_ & _50764_ /*12483*/;
assign _50768_ = _50136_ ^ _50764_ /*12486*/;
assign _50769_ = _50760_ & _50768_ /*12484*/;
assign _50584_ = _50760_ ^ _50768_ /*12485*/;
assign _50766_ = _50767_ | _50769_ /*12482*/;
assign _50771_ = ~Q[7] /*12481*/;
assign _50770_ = _50771_ & D[24] /*12480*/;
assign _50773_ = _50137_ & _50770_ /*12475*/;
assign _50774_ = _50137_ ^ _50770_ /*12478*/;
assign _50775_ = _50766_ & _50774_ /*12476*/;
assign _50585_ = _50766_ ^ _50774_ /*12477*/;
assign _50772_ = _50773_ | _50775_ /*12474*/;
assign _50777_ = ~Q[7] /*12473*/;
assign _50776_ = _50777_ & D[25] /*12472*/;
assign _50779_ = _50138_ & _50776_ /*12467*/;
assign _50780_ = _50138_ ^ _50776_ /*12470*/;
assign _50781_ = _50772_ & _50780_ /*12468*/;
assign _50586_ = _50772_ ^ _50780_ /*12469*/;
assign _50778_ = _50779_ | _50781_ /*12466*/;
assign _50783_ = ~Q[7] /*12465*/;
assign _50782_ = _50783_ & D[26] /*12464*/;
assign _50785_ = _50139_ & _50782_ /*12459*/;
assign _50786_ = _50139_ ^ _50782_ /*12462*/;
assign _50787_ = _50778_ & _50786_ /*12460*/;
assign _50587_ = _50778_ ^ _50786_ /*12461*/;
assign _50784_ = _50785_ | _50787_ /*12458*/;
assign _50789_ = ~Q[7] /*12457*/;
assign _50788_ = _50789_ & D[27] /*12456*/;
assign _50791_ = _50140_ & _50788_ /*12451*/;
assign _50792_ = _50140_ ^ _50788_ /*12454*/;
assign _50793_ = _50784_ & _50792_ /*12452*/;
assign _50588_ = _50784_ ^ _50792_ /*12453*/;
assign _50790_ = _50791_ | _50793_ /*12450*/;
assign _50795_ = ~Q[7] /*12449*/;
assign _50794_ = _50795_ & D[28] /*12448*/;
assign _50797_ = _50141_ & _50794_ /*12443*/;
assign _50798_ = _50141_ ^ _50794_ /*12446*/;
assign _50799_ = _50790_ & _50798_ /*12444*/;
assign _50589_ = _50790_ ^ _50798_ /*12445*/;
assign _50796_ = _50797_ | _50799_ /*12442*/;
assign _50801_ = ~Q[7] /*12441*/;
assign _50800_ = _50801_ & D[29] /*12440*/;
assign _50803_ = _50142_ & _50800_ /*12435*/;
assign _50804_ = _50142_ ^ _50800_ /*12438*/;
assign _50805_ = _50796_ & _50804_ /*12436*/;
assign _50590_ = _50796_ ^ _50804_ /*12437*/;
assign _50802_ = _50803_ | _50805_ /*12434*/;
assign _50807_ = ~Q[7] /*12433*/;
assign _50806_ = _50807_ & D[30] /*12432*/;
assign _50809_ = _50143_ & _50806_ /*12427*/;
assign _50810_ = _50143_ ^ _50806_ /*12430*/;
assign _50811_ = _50802_ & _50810_ /*12428*/;
assign _50591_ = _50802_ ^ _50810_ /*12429*/;
assign _50808_ = _50809_ | _50811_ /*12426*/;
assign _50813_ = ~Q[7] /*12425*/;
assign _50812_ = _50813_ & D[31] /*12424*/;
assign _50815_ = _50144_ & _50812_ /*12419*/;
assign _50816_ = _50144_ ^ _50812_ /*12422*/;
assign _50817_ = _50808_ & _50816_ /*12420*/;
assign _50592_ = _50808_ ^ _50816_ /*12421*/;
assign _50814_ = _50815_ | _50817_ /*12418*/;
assign _50819_ = ~Q[7] /*12417*/;
assign _50818_ = _50819_ & D[32] /*12416*/;
assign _50821_ = _50145_ & _50818_ /*12411*/;
assign _50822_ = _50145_ ^ _50818_ /*12414*/;
assign _50823_ = _50814_ & _50822_ /*12412*/;
assign _50593_ = _50814_ ^ _50822_ /*12413*/;
assign _50820_ = _50821_ | _50823_ /*12410*/;
assign _50825_ = ~Q[7] /*12409*/;
assign _50824_ = _50825_ & D[33] /*12408*/;
assign _50827_ = _50146_ & _50824_ /*12403*/;
assign _50828_ = _50146_ ^ _50824_ /*12406*/;
assign _50829_ = _50820_ & _50828_ /*12404*/;
assign _50594_ = _50820_ ^ _50828_ /*12405*/;
assign _50826_ = _50827_ | _50829_ /*12402*/;
assign _50831_ = ~Q[7] /*12401*/;
assign _50830_ = _50831_ & D[34] /*12400*/;
assign _50833_ = _50147_ & _50830_ /*12395*/;
assign _50834_ = _50147_ ^ _50830_ /*12398*/;
assign _50835_ = _50826_ & _50834_ /*12396*/;
assign _50595_ = _50826_ ^ _50834_ /*12397*/;
assign _50832_ = _50833_ | _50835_ /*12394*/;
assign _50837_ = ~Q[7] /*12393*/;
assign _50836_ = _50837_ & D[35] /*12392*/;
assign _50839_ = _50148_ & _50836_ /*12387*/;
assign _50840_ = _50148_ ^ _50836_ /*12390*/;
assign _50841_ = _50832_ & _50840_ /*12388*/;
assign _50596_ = _50832_ ^ _50840_ /*12389*/;
assign _50838_ = _50839_ | _50841_ /*12386*/;
assign _50843_ = ~Q[7] /*12385*/;
assign _50842_ = _50843_ & D[36] /*12384*/;
assign _50845_ = _50149_ & _50842_ /*12379*/;
assign _50846_ = _50149_ ^ _50842_ /*12382*/;
assign _50847_ = _50838_ & _50846_ /*12380*/;
assign _50597_ = _50838_ ^ _50846_ /*12381*/;
assign _50844_ = _50845_ | _50847_ /*12378*/;
assign _50849_ = ~Q[7] /*12377*/;
assign _50848_ = _50849_ & D[37] /*12376*/;
assign _50851_ = _50150_ & _50848_ /*12371*/;
assign _50852_ = _50150_ ^ _50848_ /*12374*/;
assign _50853_ = _50844_ & _50852_ /*12372*/;
assign _50598_ = _50844_ ^ _50852_ /*12373*/;
assign _50850_ = _50851_ | _50853_ /*12370*/;
assign _50855_ = ~Q[7] /*12369*/;
assign _50854_ = _50855_ & D[38] /*12368*/;
assign _50857_ = _50151_ & _50854_ /*12363*/;
assign _50858_ = _50151_ ^ _50854_ /*12366*/;
assign _50859_ = _50850_ & _50858_ /*12364*/;
assign _50599_ = _50850_ ^ _50858_ /*12365*/;
assign _50856_ = _50857_ | _50859_ /*12362*/;
assign _50861_ = ~Q[7] /*12361*/;
assign _50860_ = _50861_ & D[39] /*12360*/;
assign _50863_ = _50152_ & _50860_ /*12355*/;
assign _50864_ = _50152_ ^ _50860_ /*12358*/;
assign _50865_ = _50856_ & _50864_ /*12356*/;
assign _50600_ = _50856_ ^ _50864_ /*12357*/;
assign _50862_ = _50863_ | _50865_ /*12354*/;
assign _50867_ = ~Q[7] /*12353*/;
assign _50866_ = _50867_ & D[40] /*12352*/;
assign _50869_ = _50153_ & _50866_ /*12347*/;
assign _50870_ = _50153_ ^ _50866_ /*12350*/;
assign _50871_ = _50862_ & _50870_ /*12348*/;
assign _50601_ = _50862_ ^ _50870_ /*12349*/;
assign _50868_ = _50869_ | _50871_ /*12346*/;
assign _50873_ = ~Q[7] /*12345*/;
assign _50872_ = _50873_ & D[41] /*12344*/;
assign _50875_ = _50154_ & _50872_ /*12339*/;
assign _50876_ = _50154_ ^ _50872_ /*12342*/;
assign _50877_ = _50868_ & _50876_ /*12340*/;
assign _50602_ = _50868_ ^ _50876_ /*12341*/;
assign _50874_ = _50875_ | _50877_ /*12338*/;
assign _50879_ = ~Q[7] /*12337*/;
assign _50878_ = _50879_ & D[42] /*12336*/;
assign _50881_ = _50155_ & _50878_ /*12331*/;
assign _50882_ = _50155_ ^ _50878_ /*12334*/;
assign _50883_ = _50874_ & _50882_ /*12332*/;
assign _50603_ = _50874_ ^ _50882_ /*12333*/;
assign _50880_ = _50881_ | _50883_ /*12330*/;
assign _50885_ = ~Q[7] /*12329*/;
assign _50884_ = _50885_ & D[43] /*12328*/;
assign _50887_ = _50156_ & _50884_ /*12323*/;
assign _50888_ = _50156_ ^ _50884_ /*12326*/;
assign _50889_ = _50880_ & _50888_ /*12324*/;
assign _50604_ = _50880_ ^ _50888_ /*12325*/;
assign _50886_ = _50887_ | _50889_ /*12322*/;
assign _50891_ = ~Q[7] /*12321*/;
assign _50890_ = _50891_ & D[44] /*12320*/;
assign _50893_ = _50157_ & _50890_ /*12315*/;
assign _50894_ = _50157_ ^ _50890_ /*12318*/;
assign _50895_ = _50886_ & _50894_ /*12316*/;
assign _50605_ = _50886_ ^ _50894_ /*12317*/;
assign _50892_ = _50893_ | _50895_ /*12314*/;
assign _50897_ = ~Q[7] /*12313*/;
assign _50896_ = _50897_ & D[45] /*12312*/;
assign _50899_ = _50158_ & _50896_ /*12307*/;
assign _50900_ = _50158_ ^ _50896_ /*12310*/;
assign _50901_ = _50892_ & _50900_ /*12308*/;
assign _50606_ = _50892_ ^ _50900_ /*12309*/;
assign _50898_ = _50899_ | _50901_ /*12306*/;
assign _50903_ = ~Q[7] /*12305*/;
assign _50902_ = _50903_ & D[46] /*12304*/;
assign _50905_ = _50159_ & _50902_ /*12299*/;
assign _50906_ = _50159_ ^ _50902_ /*12302*/;
assign _50907_ = _50898_ & _50906_ /*12300*/;
assign _50607_ = _50898_ ^ _50906_ /*12301*/;
assign _50904_ = _50905_ | _50907_ /*12298*/;
assign _50909_ = ~Q[7] /*12297*/;
assign _50908_ = _50909_ & D[47] /*12296*/;
assign _50911_ = _50160_ & _50908_ /*12291*/;
assign _50912_ = _50160_ ^ _50908_ /*12294*/;
assign _50913_ = _50904_ & _50912_ /*12292*/;
assign _50608_ = _50904_ ^ _50912_ /*12293*/;
assign _50910_ = _50911_ | _50913_ /*12290*/;
assign _50915_ = ~Q[7] /*12289*/;
assign _50914_ = _50915_ & D[48] /*12288*/;
assign _50917_ = _50161_ & _50914_ /*12283*/;
assign _50918_ = _50161_ ^ _50914_ /*12286*/;
assign _50919_ = _50910_ & _50918_ /*12284*/;
assign _50609_ = _50910_ ^ _50918_ /*12285*/;
assign _50916_ = _50917_ | _50919_ /*12282*/;
assign _50921_ = ~Q[7] /*12281*/;
assign _50920_ = _50921_ & D[49] /*12280*/;
assign _50923_ = _50162_ & _50920_ /*12275*/;
assign _50924_ = _50162_ ^ _50920_ /*12278*/;
assign _50925_ = _50916_ & _50924_ /*12276*/;
assign _50610_ = _50916_ ^ _50924_ /*12277*/;
assign _50922_ = _50923_ | _50925_ /*12274*/;
assign _50927_ = ~Q[7] /*12273*/;
assign _50926_ = _50927_ & D[50] /*12272*/;
assign _50929_ = _50163_ & _50926_ /*12267*/;
assign _50930_ = _50163_ ^ _50926_ /*12270*/;
assign _50931_ = _50922_ & _50930_ /*12268*/;
assign _50611_ = _50922_ ^ _50930_ /*12269*/;
assign _50928_ = _50929_ | _50931_ /*12266*/;
assign _50933_ = ~Q[7] /*12265*/;
assign _50932_ = _50933_ & D[51] /*12264*/;
assign _50935_ = _50164_ & _50932_ /*12259*/;
assign _50936_ = _50164_ ^ _50932_ /*12262*/;
assign _50937_ = _50928_ & _50936_ /*12260*/;
assign _50612_ = _50928_ ^ _50936_ /*12261*/;
assign _50934_ = _50935_ | _50937_ /*12258*/;
assign _50939_ = ~Q[7] /*12257*/;
assign _50938_ = _50939_ & D[52] /*12256*/;
assign _50941_ = _50165_ & _50938_ /*12251*/;
assign _50942_ = _50165_ ^ _50938_ /*12254*/;
assign _50943_ = _50934_ & _50942_ /*12252*/;
assign _50613_ = _50934_ ^ _50942_ /*12253*/;
assign _50940_ = _50941_ | _50943_ /*12250*/;
assign _50945_ = ~Q[7] /*12249*/;
assign _50944_ = _50945_ & D[53] /*12248*/;
assign _50947_ = _50166_ & _50944_ /*12243*/;
assign _50948_ = _50166_ ^ _50944_ /*12246*/;
assign _50949_ = _50940_ & _50948_ /*12244*/;
assign _50614_ = _50940_ ^ _50948_ /*12245*/;
assign _50946_ = _50947_ | _50949_ /*12242*/;
assign _50951_ = ~Q[7] /*12241*/;
assign _50950_ = _50951_ & D[54] /*12240*/;
assign _50953_ = _50167_ & _50950_ /*12235*/;
assign _50954_ = _50167_ ^ _50950_ /*12238*/;
assign _50955_ = _50946_ & _50954_ /*12236*/;
assign _50615_ = _50946_ ^ _50954_ /*12237*/;
assign _50952_ = _50953_ | _50955_ /*12234*/;
assign _50957_ = ~Q[7] /*12233*/;
assign _50956_ = _50957_ & D[55] /*12232*/;
assign _50959_ = _50168_ & _50956_ /*12227*/;
assign _50960_ = _50168_ ^ _50956_ /*12230*/;
assign _50961_ = _50952_ & _50960_ /*12228*/;
assign _50616_ = _50952_ ^ _50960_ /*12229*/;
assign _50958_ = _50959_ | _50961_ /*12226*/;
assign _50963_ = ~Q[7] /*12225*/;
assign _50962_ = _50963_ & D[56] /*12224*/;
assign _50965_ = _50169_ & _50962_ /*12219*/;
assign _50966_ = _50169_ ^ _50962_ /*12222*/;
assign _50967_ = _50958_ & _50966_ /*12220*/;
assign _50617_ = _50958_ ^ _50966_ /*12221*/;
assign _50964_ = _50965_ | _50967_ /*12218*/;
assign _50969_ = ~Q[7] /*12217*/;
assign _50968_ = _50969_ & D[57] /*12216*/;
assign _50971_ = _50170_ & _50968_ /*12211*/;
assign _50972_ = _50170_ ^ _50968_ /*12214*/;
assign _50973_ = _50964_ & _50972_ /*12212*/;
assign _50618_ = _50964_ ^ _50972_ /*12213*/;
assign _50970_ = _50971_ | _50973_ /*12210*/;
assign _50975_ = ~Q[7] /*12209*/;
assign _50974_ = _50975_ & D[58] /*12208*/;
assign _50977_ = _50171_ & _50974_ /*12203*/;
assign _50978_ = _50171_ ^ _50974_ /*12206*/;
assign _50979_ = _50970_ & _50978_ /*12204*/;
assign _50619_ = _50970_ ^ _50978_ /*12205*/;
assign _50976_ = _50977_ | _50979_ /*12202*/;
assign _50981_ = ~Q[7] /*12201*/;
assign _50980_ = _50981_ & D[59] /*12200*/;
assign _50983_ = _50172_ & _50980_ /*12195*/;
assign _50984_ = _50172_ ^ _50980_ /*12198*/;
assign _50985_ = _50976_ & _50984_ /*12196*/;
assign _50620_ = _50976_ ^ _50984_ /*12197*/;
assign _50982_ = _50983_ | _50985_ /*12194*/;
assign _50987_ = ~Q[7] /*12193*/;
assign _50986_ = _50987_ & D[60] /*12192*/;
assign _50989_ = _50173_ & _50986_ /*12187*/;
assign _50990_ = _50173_ ^ _50986_ /*12190*/;
assign _50991_ = _50982_ & _50990_ /*12188*/;
assign _50621_ = _50982_ ^ _50990_ /*12189*/;
assign _50988_ = _50989_ | _50991_ /*12186*/;
assign _50993_ = ~Q[7] /*12185*/;
assign _50992_ = _50993_ & D[61] /*12184*/;
assign _50995_ = _50174_ & _50992_ /*12179*/;
assign _50996_ = _50174_ ^ _50992_ /*12182*/;
assign _50997_ = _50988_ & _50996_ /*12180*/;
assign _50622_ = _50988_ ^ _50996_ /*12181*/;
assign _50994_ = _50995_ | _50997_ /*12178*/;
assign _50999_ = ~Q[7] /*12177*/;
assign _50998_ = _50999_ & D[62] /*12176*/;
assign _51001_ = _50175_ & _50998_ /*12171*/;
assign _51002_ = _50175_ ^ _50998_ /*12174*/;
assign _51003_ = _50994_ & _51002_ /*12172*/;
assign _50623_ = _50994_ ^ _51002_ /*12173*/;
assign _51000_ = _51001_ | _51003_ /*12170*/;
assign _51005_ = ~Q[7] /*12169*/;
assign _51004_ = _51005_ & zeroWire /*12168*/;
assign _51006_ = _50176_ ^ _51004_ /*12166*/;
assign _50624_ = _51006_ ^ _51000_ /*12165*/;
assign _51077_ = ~D[0] /*11911*/;
assign _51074_ = R_0[6] & _51077_ /*11907*/;
assign _51075_ = R_0[6] ^ _51077_ /*11910*/;
assign _51076_ = oneWire & _51075_ /*11908*/;
assign _51009_ = oneWire ^ _51075_ /*11909*/;
assign _51073_ = _51074_ | _51076_ /*11906*/;
assign _51082_ = ~D[1] /*11905*/;
assign _51079_ = _50561_ & _51082_ /*11901*/;
assign _51080_ = _50561_ ^ _51082_ /*11904*/;
assign _51081_ = _51073_ & _51080_ /*11902*/;
assign _51010_ = _51073_ ^ _51080_ /*11903*/;
assign _51078_ = _51079_ | _51081_ /*11900*/;
assign _51087_ = ~D[2] /*11899*/;
assign _51084_ = _50562_ & _51087_ /*11895*/;
assign _51085_ = _50562_ ^ _51087_ /*11898*/;
assign _51086_ = _51078_ & _51085_ /*11896*/;
assign _51011_ = _51078_ ^ _51085_ /*11897*/;
assign _51083_ = _51084_ | _51086_ /*11894*/;
assign _51092_ = ~D[3] /*11893*/;
assign _51089_ = _50563_ & _51092_ /*11889*/;
assign _51090_ = _50563_ ^ _51092_ /*11892*/;
assign _51091_ = _51083_ & _51090_ /*11890*/;
assign _51012_ = _51083_ ^ _51090_ /*11891*/;
assign _51088_ = _51089_ | _51091_ /*11888*/;
assign _51097_ = ~D[4] /*11887*/;
assign _51094_ = _50564_ & _51097_ /*11883*/;
assign _51095_ = _50564_ ^ _51097_ /*11886*/;
assign _51096_ = _51088_ & _51095_ /*11884*/;
assign _51013_ = _51088_ ^ _51095_ /*11885*/;
assign _51093_ = _51094_ | _51096_ /*11882*/;
assign _51102_ = ~D[5] /*11881*/;
assign _51099_ = _50565_ & _51102_ /*11877*/;
assign _51100_ = _50565_ ^ _51102_ /*11880*/;
assign _51101_ = _51093_ & _51100_ /*11878*/;
assign _51014_ = _51093_ ^ _51100_ /*11879*/;
assign _51098_ = _51099_ | _51101_ /*11876*/;
assign _51107_ = ~D[6] /*11875*/;
assign _51104_ = _50566_ & _51107_ /*11871*/;
assign _51105_ = _50566_ ^ _51107_ /*11874*/;
assign _51106_ = _51098_ & _51105_ /*11872*/;
assign _51015_ = _51098_ ^ _51105_ /*11873*/;
assign _51103_ = _51104_ | _51106_ /*11870*/;
assign _51112_ = ~D[7] /*11869*/;
assign _51109_ = _50567_ & _51112_ /*11865*/;
assign _51110_ = _50567_ ^ _51112_ /*11868*/;
assign _51111_ = _51103_ & _51110_ /*11866*/;
assign _51016_ = _51103_ ^ _51110_ /*11867*/;
assign _51108_ = _51109_ | _51111_ /*11864*/;
assign _51117_ = ~D[8] /*11863*/;
assign _51114_ = _50568_ & _51117_ /*11859*/;
assign _51115_ = _50568_ ^ _51117_ /*11862*/;
assign _51116_ = _51108_ & _51115_ /*11860*/;
assign _51017_ = _51108_ ^ _51115_ /*11861*/;
assign _51113_ = _51114_ | _51116_ /*11858*/;
assign _51122_ = ~D[9] /*11857*/;
assign _51119_ = _50569_ & _51122_ /*11853*/;
assign _51120_ = _50569_ ^ _51122_ /*11856*/;
assign _51121_ = _51113_ & _51120_ /*11854*/;
assign _51018_ = _51113_ ^ _51120_ /*11855*/;
assign _51118_ = _51119_ | _51121_ /*11852*/;
assign _51127_ = ~D[10] /*11851*/;
assign _51124_ = _50570_ & _51127_ /*11847*/;
assign _51125_ = _50570_ ^ _51127_ /*11850*/;
assign _51126_ = _51118_ & _51125_ /*11848*/;
assign _51019_ = _51118_ ^ _51125_ /*11849*/;
assign _51123_ = _51124_ | _51126_ /*11846*/;
assign _51132_ = ~D[11] /*11845*/;
assign _51129_ = _50571_ & _51132_ /*11841*/;
assign _51130_ = _50571_ ^ _51132_ /*11844*/;
assign _51131_ = _51123_ & _51130_ /*11842*/;
assign _51020_ = _51123_ ^ _51130_ /*11843*/;
assign _51128_ = _51129_ | _51131_ /*11840*/;
assign _51137_ = ~D[12] /*11839*/;
assign _51134_ = _50572_ & _51137_ /*11835*/;
assign _51135_ = _50572_ ^ _51137_ /*11838*/;
assign _51136_ = _51128_ & _51135_ /*11836*/;
assign _51021_ = _51128_ ^ _51135_ /*11837*/;
assign _51133_ = _51134_ | _51136_ /*11834*/;
assign _51142_ = ~D[13] /*11833*/;
assign _51139_ = _50573_ & _51142_ /*11829*/;
assign _51140_ = _50573_ ^ _51142_ /*11832*/;
assign _51141_ = _51133_ & _51140_ /*11830*/;
assign _51022_ = _51133_ ^ _51140_ /*11831*/;
assign _51138_ = _51139_ | _51141_ /*11828*/;
assign _51147_ = ~D[14] /*11827*/;
assign _51144_ = _50574_ & _51147_ /*11823*/;
assign _51145_ = _50574_ ^ _51147_ /*11826*/;
assign _51146_ = _51138_ & _51145_ /*11824*/;
assign _51023_ = _51138_ ^ _51145_ /*11825*/;
assign _51143_ = _51144_ | _51146_ /*11822*/;
assign _51152_ = ~D[15] /*11821*/;
assign _51149_ = _50575_ & _51152_ /*11817*/;
assign _51150_ = _50575_ ^ _51152_ /*11820*/;
assign _51151_ = _51143_ & _51150_ /*11818*/;
assign _51024_ = _51143_ ^ _51150_ /*11819*/;
assign _51148_ = _51149_ | _51151_ /*11816*/;
assign _51157_ = ~D[16] /*11815*/;
assign _51154_ = _50576_ & _51157_ /*11811*/;
assign _51155_ = _50576_ ^ _51157_ /*11814*/;
assign _51156_ = _51148_ & _51155_ /*11812*/;
assign _51025_ = _51148_ ^ _51155_ /*11813*/;
assign _51153_ = _51154_ | _51156_ /*11810*/;
assign _51162_ = ~D[17] /*11809*/;
assign _51159_ = _50577_ & _51162_ /*11805*/;
assign _51160_ = _50577_ ^ _51162_ /*11808*/;
assign _51161_ = _51153_ & _51160_ /*11806*/;
assign _51026_ = _51153_ ^ _51160_ /*11807*/;
assign _51158_ = _51159_ | _51161_ /*11804*/;
assign _51167_ = ~D[18] /*11803*/;
assign _51164_ = _50578_ & _51167_ /*11799*/;
assign _51165_ = _50578_ ^ _51167_ /*11802*/;
assign _51166_ = _51158_ & _51165_ /*11800*/;
assign _51027_ = _51158_ ^ _51165_ /*11801*/;
assign _51163_ = _51164_ | _51166_ /*11798*/;
assign _51172_ = ~D[19] /*11797*/;
assign _51169_ = _50579_ & _51172_ /*11793*/;
assign _51170_ = _50579_ ^ _51172_ /*11796*/;
assign _51171_ = _51163_ & _51170_ /*11794*/;
assign _51028_ = _51163_ ^ _51170_ /*11795*/;
assign _51168_ = _51169_ | _51171_ /*11792*/;
assign _51177_ = ~D[20] /*11791*/;
assign _51174_ = _50580_ & _51177_ /*11787*/;
assign _51175_ = _50580_ ^ _51177_ /*11790*/;
assign _51176_ = _51168_ & _51175_ /*11788*/;
assign _51029_ = _51168_ ^ _51175_ /*11789*/;
assign _51173_ = _51174_ | _51176_ /*11786*/;
assign _51182_ = ~D[21] /*11785*/;
assign _51179_ = _50581_ & _51182_ /*11781*/;
assign _51180_ = _50581_ ^ _51182_ /*11784*/;
assign _51181_ = _51173_ & _51180_ /*11782*/;
assign _51030_ = _51173_ ^ _51180_ /*11783*/;
assign _51178_ = _51179_ | _51181_ /*11780*/;
assign _51187_ = ~D[22] /*11779*/;
assign _51184_ = _50582_ & _51187_ /*11775*/;
assign _51185_ = _50582_ ^ _51187_ /*11778*/;
assign _51186_ = _51178_ & _51185_ /*11776*/;
assign _51031_ = _51178_ ^ _51185_ /*11777*/;
assign _51183_ = _51184_ | _51186_ /*11774*/;
assign _51192_ = ~D[23] /*11773*/;
assign _51189_ = _50583_ & _51192_ /*11769*/;
assign _51190_ = _50583_ ^ _51192_ /*11772*/;
assign _51191_ = _51183_ & _51190_ /*11770*/;
assign _51032_ = _51183_ ^ _51190_ /*11771*/;
assign _51188_ = _51189_ | _51191_ /*11768*/;
assign _51197_ = ~D[24] /*11767*/;
assign _51194_ = _50584_ & _51197_ /*11763*/;
assign _51195_ = _50584_ ^ _51197_ /*11766*/;
assign _51196_ = _51188_ & _51195_ /*11764*/;
assign _51033_ = _51188_ ^ _51195_ /*11765*/;
assign _51193_ = _51194_ | _51196_ /*11762*/;
assign _51202_ = ~D[25] /*11761*/;
assign _51199_ = _50585_ & _51202_ /*11757*/;
assign _51200_ = _50585_ ^ _51202_ /*11760*/;
assign _51201_ = _51193_ & _51200_ /*11758*/;
assign _51034_ = _51193_ ^ _51200_ /*11759*/;
assign _51198_ = _51199_ | _51201_ /*11756*/;
assign _51207_ = ~D[26] /*11755*/;
assign _51204_ = _50586_ & _51207_ /*11751*/;
assign _51205_ = _50586_ ^ _51207_ /*11754*/;
assign _51206_ = _51198_ & _51205_ /*11752*/;
assign _51035_ = _51198_ ^ _51205_ /*11753*/;
assign _51203_ = _51204_ | _51206_ /*11750*/;
assign _51212_ = ~D[27] /*11749*/;
assign _51209_ = _50587_ & _51212_ /*11745*/;
assign _51210_ = _50587_ ^ _51212_ /*11748*/;
assign _51211_ = _51203_ & _51210_ /*11746*/;
assign _51036_ = _51203_ ^ _51210_ /*11747*/;
assign _51208_ = _51209_ | _51211_ /*11744*/;
assign _51217_ = ~D[28] /*11743*/;
assign _51214_ = _50588_ & _51217_ /*11739*/;
assign _51215_ = _50588_ ^ _51217_ /*11742*/;
assign _51216_ = _51208_ & _51215_ /*11740*/;
assign _51037_ = _51208_ ^ _51215_ /*11741*/;
assign _51213_ = _51214_ | _51216_ /*11738*/;
assign _51222_ = ~D[29] /*11737*/;
assign _51219_ = _50589_ & _51222_ /*11733*/;
assign _51220_ = _50589_ ^ _51222_ /*11736*/;
assign _51221_ = _51213_ & _51220_ /*11734*/;
assign _51038_ = _51213_ ^ _51220_ /*11735*/;
assign _51218_ = _51219_ | _51221_ /*11732*/;
assign _51227_ = ~D[30] /*11731*/;
assign _51224_ = _50590_ & _51227_ /*11727*/;
assign _51225_ = _50590_ ^ _51227_ /*11730*/;
assign _51226_ = _51218_ & _51225_ /*11728*/;
assign _51039_ = _51218_ ^ _51225_ /*11729*/;
assign _51223_ = _51224_ | _51226_ /*11726*/;
assign _51232_ = ~D[31] /*11725*/;
assign _51229_ = _50591_ & _51232_ /*11721*/;
assign _51230_ = _50591_ ^ _51232_ /*11724*/;
assign _51231_ = _51223_ & _51230_ /*11722*/;
assign _51040_ = _51223_ ^ _51230_ /*11723*/;
assign _51228_ = _51229_ | _51231_ /*11720*/;
assign _51237_ = ~D[32] /*11719*/;
assign _51234_ = _50592_ & _51237_ /*11715*/;
assign _51235_ = _50592_ ^ _51237_ /*11718*/;
assign _51236_ = _51228_ & _51235_ /*11716*/;
assign _51041_ = _51228_ ^ _51235_ /*11717*/;
assign _51233_ = _51234_ | _51236_ /*11714*/;
assign _51242_ = ~D[33] /*11713*/;
assign _51239_ = _50593_ & _51242_ /*11709*/;
assign _51240_ = _50593_ ^ _51242_ /*11712*/;
assign _51241_ = _51233_ & _51240_ /*11710*/;
assign _51042_ = _51233_ ^ _51240_ /*11711*/;
assign _51238_ = _51239_ | _51241_ /*11708*/;
assign _51247_ = ~D[34] /*11707*/;
assign _51244_ = _50594_ & _51247_ /*11703*/;
assign _51245_ = _50594_ ^ _51247_ /*11706*/;
assign _51246_ = _51238_ & _51245_ /*11704*/;
assign _51043_ = _51238_ ^ _51245_ /*11705*/;
assign _51243_ = _51244_ | _51246_ /*11702*/;
assign _51252_ = ~D[35] /*11701*/;
assign _51249_ = _50595_ & _51252_ /*11697*/;
assign _51250_ = _50595_ ^ _51252_ /*11700*/;
assign _51251_ = _51243_ & _51250_ /*11698*/;
assign _51044_ = _51243_ ^ _51250_ /*11699*/;
assign _51248_ = _51249_ | _51251_ /*11696*/;
assign _51257_ = ~D[36] /*11695*/;
assign _51254_ = _50596_ & _51257_ /*11691*/;
assign _51255_ = _50596_ ^ _51257_ /*11694*/;
assign _51256_ = _51248_ & _51255_ /*11692*/;
assign _51045_ = _51248_ ^ _51255_ /*11693*/;
assign _51253_ = _51254_ | _51256_ /*11690*/;
assign _51262_ = ~D[37] /*11689*/;
assign _51259_ = _50597_ & _51262_ /*11685*/;
assign _51260_ = _50597_ ^ _51262_ /*11688*/;
assign _51261_ = _51253_ & _51260_ /*11686*/;
assign _51046_ = _51253_ ^ _51260_ /*11687*/;
assign _51258_ = _51259_ | _51261_ /*11684*/;
assign _51267_ = ~D[38] /*11683*/;
assign _51264_ = _50598_ & _51267_ /*11679*/;
assign _51265_ = _50598_ ^ _51267_ /*11682*/;
assign _51266_ = _51258_ & _51265_ /*11680*/;
assign _51047_ = _51258_ ^ _51265_ /*11681*/;
assign _51263_ = _51264_ | _51266_ /*11678*/;
assign _51272_ = ~D[39] /*11677*/;
assign _51269_ = _50599_ & _51272_ /*11673*/;
assign _51270_ = _50599_ ^ _51272_ /*11676*/;
assign _51271_ = _51263_ & _51270_ /*11674*/;
assign _51048_ = _51263_ ^ _51270_ /*11675*/;
assign _51268_ = _51269_ | _51271_ /*11672*/;
assign _51277_ = ~D[40] /*11671*/;
assign _51274_ = _50600_ & _51277_ /*11667*/;
assign _51275_ = _50600_ ^ _51277_ /*11670*/;
assign _51276_ = _51268_ & _51275_ /*11668*/;
assign _51049_ = _51268_ ^ _51275_ /*11669*/;
assign _51273_ = _51274_ | _51276_ /*11666*/;
assign _51282_ = ~D[41] /*11665*/;
assign _51279_ = _50601_ & _51282_ /*11661*/;
assign _51280_ = _50601_ ^ _51282_ /*11664*/;
assign _51281_ = _51273_ & _51280_ /*11662*/;
assign _51050_ = _51273_ ^ _51280_ /*11663*/;
assign _51278_ = _51279_ | _51281_ /*11660*/;
assign _51287_ = ~D[42] /*11659*/;
assign _51284_ = _50602_ & _51287_ /*11655*/;
assign _51285_ = _50602_ ^ _51287_ /*11658*/;
assign _51286_ = _51278_ & _51285_ /*11656*/;
assign _51051_ = _51278_ ^ _51285_ /*11657*/;
assign _51283_ = _51284_ | _51286_ /*11654*/;
assign _51292_ = ~D[43] /*11653*/;
assign _51289_ = _50603_ & _51292_ /*11649*/;
assign _51290_ = _50603_ ^ _51292_ /*11652*/;
assign _51291_ = _51283_ & _51290_ /*11650*/;
assign _51052_ = _51283_ ^ _51290_ /*11651*/;
assign _51288_ = _51289_ | _51291_ /*11648*/;
assign _51297_ = ~D[44] /*11647*/;
assign _51294_ = _50604_ & _51297_ /*11643*/;
assign _51295_ = _50604_ ^ _51297_ /*11646*/;
assign _51296_ = _51288_ & _51295_ /*11644*/;
assign _51053_ = _51288_ ^ _51295_ /*11645*/;
assign _51293_ = _51294_ | _51296_ /*11642*/;
assign _51302_ = ~D[45] /*11641*/;
assign _51299_ = _50605_ & _51302_ /*11637*/;
assign _51300_ = _50605_ ^ _51302_ /*11640*/;
assign _51301_ = _51293_ & _51300_ /*11638*/;
assign _51054_ = _51293_ ^ _51300_ /*11639*/;
assign _51298_ = _51299_ | _51301_ /*11636*/;
assign _51307_ = ~D[46] /*11635*/;
assign _51304_ = _50606_ & _51307_ /*11631*/;
assign _51305_ = _50606_ ^ _51307_ /*11634*/;
assign _51306_ = _51298_ & _51305_ /*11632*/;
assign _51055_ = _51298_ ^ _51305_ /*11633*/;
assign _51303_ = _51304_ | _51306_ /*11630*/;
assign _51312_ = ~D[47] /*11629*/;
assign _51309_ = _50607_ & _51312_ /*11625*/;
assign _51310_ = _50607_ ^ _51312_ /*11628*/;
assign _51311_ = _51303_ & _51310_ /*11626*/;
assign _51056_ = _51303_ ^ _51310_ /*11627*/;
assign _51308_ = _51309_ | _51311_ /*11624*/;
assign _51317_ = ~D[48] /*11623*/;
assign _51314_ = _50608_ & _51317_ /*11619*/;
assign _51315_ = _50608_ ^ _51317_ /*11622*/;
assign _51316_ = _51308_ & _51315_ /*11620*/;
assign _51057_ = _51308_ ^ _51315_ /*11621*/;
assign _51313_ = _51314_ | _51316_ /*11618*/;
assign _51322_ = ~D[49] /*11617*/;
assign _51319_ = _50609_ & _51322_ /*11613*/;
assign _51320_ = _50609_ ^ _51322_ /*11616*/;
assign _51321_ = _51313_ & _51320_ /*11614*/;
assign _51058_ = _51313_ ^ _51320_ /*11615*/;
assign _51318_ = _51319_ | _51321_ /*11612*/;
assign _51327_ = ~D[50] /*11611*/;
assign _51324_ = _50610_ & _51327_ /*11607*/;
assign _51325_ = _50610_ ^ _51327_ /*11610*/;
assign _51326_ = _51318_ & _51325_ /*11608*/;
assign _51059_ = _51318_ ^ _51325_ /*11609*/;
assign _51323_ = _51324_ | _51326_ /*11606*/;
assign _51332_ = ~D[51] /*11605*/;
assign _51329_ = _50611_ & _51332_ /*11601*/;
assign _51330_ = _50611_ ^ _51332_ /*11604*/;
assign _51331_ = _51323_ & _51330_ /*11602*/;
assign _51060_ = _51323_ ^ _51330_ /*11603*/;
assign _51328_ = _51329_ | _51331_ /*11600*/;
assign _51337_ = ~D[52] /*11599*/;
assign _51334_ = _50612_ & _51337_ /*11595*/;
assign _51335_ = _50612_ ^ _51337_ /*11598*/;
assign _51336_ = _51328_ & _51335_ /*11596*/;
assign _51061_ = _51328_ ^ _51335_ /*11597*/;
assign _51333_ = _51334_ | _51336_ /*11594*/;
assign _51342_ = ~D[53] /*11593*/;
assign _51339_ = _50613_ & _51342_ /*11589*/;
assign _51340_ = _50613_ ^ _51342_ /*11592*/;
assign _51341_ = _51333_ & _51340_ /*11590*/;
assign _51062_ = _51333_ ^ _51340_ /*11591*/;
assign _51338_ = _51339_ | _51341_ /*11588*/;
assign _51347_ = ~D[54] /*11587*/;
assign _51344_ = _50614_ & _51347_ /*11583*/;
assign _51345_ = _50614_ ^ _51347_ /*11586*/;
assign _51346_ = _51338_ & _51345_ /*11584*/;
assign _51063_ = _51338_ ^ _51345_ /*11585*/;
assign _51343_ = _51344_ | _51346_ /*11582*/;
assign _51352_ = ~D[55] /*11581*/;
assign _51349_ = _50615_ & _51352_ /*11577*/;
assign _51350_ = _50615_ ^ _51352_ /*11580*/;
assign _51351_ = _51343_ & _51350_ /*11578*/;
assign _51064_ = _51343_ ^ _51350_ /*11579*/;
assign _51348_ = _51349_ | _51351_ /*11576*/;
assign _51357_ = ~D[56] /*11575*/;
assign _51354_ = _50616_ & _51357_ /*11571*/;
assign _51355_ = _50616_ ^ _51357_ /*11574*/;
assign _51356_ = _51348_ & _51355_ /*11572*/;
assign _51065_ = _51348_ ^ _51355_ /*11573*/;
assign _51353_ = _51354_ | _51356_ /*11570*/;
assign _51362_ = ~D[57] /*11569*/;
assign _51359_ = _50617_ & _51362_ /*11565*/;
assign _51360_ = _50617_ ^ _51362_ /*11568*/;
assign _51361_ = _51353_ & _51360_ /*11566*/;
assign _51066_ = _51353_ ^ _51360_ /*11567*/;
assign _51358_ = _51359_ | _51361_ /*11564*/;
assign _51367_ = ~D[58] /*11563*/;
assign _51364_ = _50618_ & _51367_ /*11559*/;
assign _51365_ = _50618_ ^ _51367_ /*11562*/;
assign _51366_ = _51358_ & _51365_ /*11560*/;
assign _51067_ = _51358_ ^ _51365_ /*11561*/;
assign _51363_ = _51364_ | _51366_ /*11558*/;
assign _51372_ = ~D[59] /*11557*/;
assign _51369_ = _50619_ & _51372_ /*11553*/;
assign _51370_ = _50619_ ^ _51372_ /*11556*/;
assign _51371_ = _51363_ & _51370_ /*11554*/;
assign _51068_ = _51363_ ^ _51370_ /*11555*/;
assign _51368_ = _51369_ | _51371_ /*11552*/;
assign _51377_ = ~D[60] /*11551*/;
assign _51374_ = _50620_ & _51377_ /*11547*/;
assign _51375_ = _50620_ ^ _51377_ /*11550*/;
assign _51376_ = _51368_ & _51375_ /*11548*/;
assign _51069_ = _51368_ ^ _51375_ /*11549*/;
assign _51373_ = _51374_ | _51376_ /*11546*/;
assign _51382_ = ~D[61] /*11545*/;
assign _51379_ = _50621_ & _51382_ /*11541*/;
assign _51380_ = _50621_ ^ _51382_ /*11544*/;
assign _51381_ = _51373_ & _51380_ /*11542*/;
assign _51070_ = _51373_ ^ _51380_ /*11543*/;
assign _51378_ = _51379_ | _51381_ /*11540*/;
assign _51387_ = ~D[62] /*11539*/;
assign _51384_ = _50622_ & _51387_ /*11535*/;
assign _51385_ = _50622_ ^ _51387_ /*11538*/;
assign _51386_ = _51378_ & _51385_ /*11536*/;
assign _51071_ = _51378_ ^ _51385_ /*11537*/;
assign _51383_ = _51384_ | _51386_ /*11534*/;
assign _51388_ = _50623_ & oneWire /*11529*/;
assign _51389_ = _50623_ ^ oneWire /*11532*/;
assign _51390_ = _51383_ & _51389_ /*11530*/;
assign _51072_ = _51383_ ^ _51389_ /*11531*/;
assign Q[6] = _51388_ | _51390_ /*11528*/;
assign _51523_ = ~Q[6] /*11143*/;
assign _51522_ = _51523_ & D[0] /*11142*/;
assign _51525_ = _51009_ & _51522_ /*11137*/;
assign _51526_ = _51009_ ^ _51522_ /*11140*/;
assign _51527_ = zeroWire & _51526_ /*11138*/;
assign _51457_ = zeroWire ^ _51526_ /*11139*/;
assign _51524_ = _51525_ | _51527_ /*11136*/;
assign _51529_ = ~Q[6] /*11135*/;
assign _51528_ = _51529_ & D[1] /*11134*/;
assign _51531_ = _51010_ & _51528_ /*11129*/;
assign _51532_ = _51010_ ^ _51528_ /*11132*/;
assign _51533_ = _51524_ & _51532_ /*11130*/;
assign _51458_ = _51524_ ^ _51532_ /*11131*/;
assign _51530_ = _51531_ | _51533_ /*11128*/;
assign _51535_ = ~Q[6] /*11127*/;
assign _51534_ = _51535_ & D[2] /*11126*/;
assign _51537_ = _51011_ & _51534_ /*11121*/;
assign _51538_ = _51011_ ^ _51534_ /*11124*/;
assign _51539_ = _51530_ & _51538_ /*11122*/;
assign _51459_ = _51530_ ^ _51538_ /*11123*/;
assign _51536_ = _51537_ | _51539_ /*11120*/;
assign _51541_ = ~Q[6] /*11119*/;
assign _51540_ = _51541_ & D[3] /*11118*/;
assign _51543_ = _51012_ & _51540_ /*11113*/;
assign _51544_ = _51012_ ^ _51540_ /*11116*/;
assign _51545_ = _51536_ & _51544_ /*11114*/;
assign _51460_ = _51536_ ^ _51544_ /*11115*/;
assign _51542_ = _51543_ | _51545_ /*11112*/;
assign _51547_ = ~Q[6] /*11111*/;
assign _51546_ = _51547_ & D[4] /*11110*/;
assign _51549_ = _51013_ & _51546_ /*11105*/;
assign _51550_ = _51013_ ^ _51546_ /*11108*/;
assign _51551_ = _51542_ & _51550_ /*11106*/;
assign _51461_ = _51542_ ^ _51550_ /*11107*/;
assign _51548_ = _51549_ | _51551_ /*11104*/;
assign _51553_ = ~Q[6] /*11103*/;
assign _51552_ = _51553_ & D[5] /*11102*/;
assign _51555_ = _51014_ & _51552_ /*11097*/;
assign _51556_ = _51014_ ^ _51552_ /*11100*/;
assign _51557_ = _51548_ & _51556_ /*11098*/;
assign _51462_ = _51548_ ^ _51556_ /*11099*/;
assign _51554_ = _51555_ | _51557_ /*11096*/;
assign _51559_ = ~Q[6] /*11095*/;
assign _51558_ = _51559_ & D[6] /*11094*/;
assign _51561_ = _51015_ & _51558_ /*11089*/;
assign _51562_ = _51015_ ^ _51558_ /*11092*/;
assign _51563_ = _51554_ & _51562_ /*11090*/;
assign _51463_ = _51554_ ^ _51562_ /*11091*/;
assign _51560_ = _51561_ | _51563_ /*11088*/;
assign _51565_ = ~Q[6] /*11087*/;
assign _51564_ = _51565_ & D[7] /*11086*/;
assign _51567_ = _51016_ & _51564_ /*11081*/;
assign _51568_ = _51016_ ^ _51564_ /*11084*/;
assign _51569_ = _51560_ & _51568_ /*11082*/;
assign _51464_ = _51560_ ^ _51568_ /*11083*/;
assign _51566_ = _51567_ | _51569_ /*11080*/;
assign _51571_ = ~Q[6] /*11079*/;
assign _51570_ = _51571_ & D[8] /*11078*/;
assign _51573_ = _51017_ & _51570_ /*11073*/;
assign _51574_ = _51017_ ^ _51570_ /*11076*/;
assign _51575_ = _51566_ & _51574_ /*11074*/;
assign _51465_ = _51566_ ^ _51574_ /*11075*/;
assign _51572_ = _51573_ | _51575_ /*11072*/;
assign _51577_ = ~Q[6] /*11071*/;
assign _51576_ = _51577_ & D[9] /*11070*/;
assign _51579_ = _51018_ & _51576_ /*11065*/;
assign _51580_ = _51018_ ^ _51576_ /*11068*/;
assign _51581_ = _51572_ & _51580_ /*11066*/;
assign _51466_ = _51572_ ^ _51580_ /*11067*/;
assign _51578_ = _51579_ | _51581_ /*11064*/;
assign _51583_ = ~Q[6] /*11063*/;
assign _51582_ = _51583_ & D[10] /*11062*/;
assign _51585_ = _51019_ & _51582_ /*11057*/;
assign _51586_ = _51019_ ^ _51582_ /*11060*/;
assign _51587_ = _51578_ & _51586_ /*11058*/;
assign _51467_ = _51578_ ^ _51586_ /*11059*/;
assign _51584_ = _51585_ | _51587_ /*11056*/;
assign _51589_ = ~Q[6] /*11055*/;
assign _51588_ = _51589_ & D[11] /*11054*/;
assign _51591_ = _51020_ & _51588_ /*11049*/;
assign _51592_ = _51020_ ^ _51588_ /*11052*/;
assign _51593_ = _51584_ & _51592_ /*11050*/;
assign _51468_ = _51584_ ^ _51592_ /*11051*/;
assign _51590_ = _51591_ | _51593_ /*11048*/;
assign _51595_ = ~Q[6] /*11047*/;
assign _51594_ = _51595_ & D[12] /*11046*/;
assign _51597_ = _51021_ & _51594_ /*11041*/;
assign _51598_ = _51021_ ^ _51594_ /*11044*/;
assign _51599_ = _51590_ & _51598_ /*11042*/;
assign _51469_ = _51590_ ^ _51598_ /*11043*/;
assign _51596_ = _51597_ | _51599_ /*11040*/;
assign _51601_ = ~Q[6] /*11039*/;
assign _51600_ = _51601_ & D[13] /*11038*/;
assign _51603_ = _51022_ & _51600_ /*11033*/;
assign _51604_ = _51022_ ^ _51600_ /*11036*/;
assign _51605_ = _51596_ & _51604_ /*11034*/;
assign _51470_ = _51596_ ^ _51604_ /*11035*/;
assign _51602_ = _51603_ | _51605_ /*11032*/;
assign _51607_ = ~Q[6] /*11031*/;
assign _51606_ = _51607_ & D[14] /*11030*/;
assign _51609_ = _51023_ & _51606_ /*11025*/;
assign _51610_ = _51023_ ^ _51606_ /*11028*/;
assign _51611_ = _51602_ & _51610_ /*11026*/;
assign _51471_ = _51602_ ^ _51610_ /*11027*/;
assign _51608_ = _51609_ | _51611_ /*11024*/;
assign _51613_ = ~Q[6] /*11023*/;
assign _51612_ = _51613_ & D[15] /*11022*/;
assign _51615_ = _51024_ & _51612_ /*11017*/;
assign _51616_ = _51024_ ^ _51612_ /*11020*/;
assign _51617_ = _51608_ & _51616_ /*11018*/;
assign _51472_ = _51608_ ^ _51616_ /*11019*/;
assign _51614_ = _51615_ | _51617_ /*11016*/;
assign _51619_ = ~Q[6] /*11015*/;
assign _51618_ = _51619_ & D[16] /*11014*/;
assign _51621_ = _51025_ & _51618_ /*11009*/;
assign _51622_ = _51025_ ^ _51618_ /*11012*/;
assign _51623_ = _51614_ & _51622_ /*11010*/;
assign _51473_ = _51614_ ^ _51622_ /*11011*/;
assign _51620_ = _51621_ | _51623_ /*11008*/;
assign _51625_ = ~Q[6] /*11007*/;
assign _51624_ = _51625_ & D[17] /*11006*/;
assign _51627_ = _51026_ & _51624_ /*11001*/;
assign _51628_ = _51026_ ^ _51624_ /*11004*/;
assign _51629_ = _51620_ & _51628_ /*11002*/;
assign _51474_ = _51620_ ^ _51628_ /*11003*/;
assign _51626_ = _51627_ | _51629_ /*11000*/;
assign _51631_ = ~Q[6] /*10999*/;
assign _51630_ = _51631_ & D[18] /*10998*/;
assign _51633_ = _51027_ & _51630_ /*10993*/;
assign _51634_ = _51027_ ^ _51630_ /*10996*/;
assign _51635_ = _51626_ & _51634_ /*10994*/;
assign _51475_ = _51626_ ^ _51634_ /*10995*/;
assign _51632_ = _51633_ | _51635_ /*10992*/;
assign _51637_ = ~Q[6] /*10991*/;
assign _51636_ = _51637_ & D[19] /*10990*/;
assign _51639_ = _51028_ & _51636_ /*10985*/;
assign _51640_ = _51028_ ^ _51636_ /*10988*/;
assign _51641_ = _51632_ & _51640_ /*10986*/;
assign _51476_ = _51632_ ^ _51640_ /*10987*/;
assign _51638_ = _51639_ | _51641_ /*10984*/;
assign _51643_ = ~Q[6] /*10983*/;
assign _51642_ = _51643_ & D[20] /*10982*/;
assign _51645_ = _51029_ & _51642_ /*10977*/;
assign _51646_ = _51029_ ^ _51642_ /*10980*/;
assign _51647_ = _51638_ & _51646_ /*10978*/;
assign _51477_ = _51638_ ^ _51646_ /*10979*/;
assign _51644_ = _51645_ | _51647_ /*10976*/;
assign _51649_ = ~Q[6] /*10975*/;
assign _51648_ = _51649_ & D[21] /*10974*/;
assign _51651_ = _51030_ & _51648_ /*10969*/;
assign _51652_ = _51030_ ^ _51648_ /*10972*/;
assign _51653_ = _51644_ & _51652_ /*10970*/;
assign _51478_ = _51644_ ^ _51652_ /*10971*/;
assign _51650_ = _51651_ | _51653_ /*10968*/;
assign _51655_ = ~Q[6] /*10967*/;
assign _51654_ = _51655_ & D[22] /*10966*/;
assign _51657_ = _51031_ & _51654_ /*10961*/;
assign _51658_ = _51031_ ^ _51654_ /*10964*/;
assign _51659_ = _51650_ & _51658_ /*10962*/;
assign _51479_ = _51650_ ^ _51658_ /*10963*/;
assign _51656_ = _51657_ | _51659_ /*10960*/;
assign _51661_ = ~Q[6] /*10959*/;
assign _51660_ = _51661_ & D[23] /*10958*/;
assign _51663_ = _51032_ & _51660_ /*10953*/;
assign _51664_ = _51032_ ^ _51660_ /*10956*/;
assign _51665_ = _51656_ & _51664_ /*10954*/;
assign _51480_ = _51656_ ^ _51664_ /*10955*/;
assign _51662_ = _51663_ | _51665_ /*10952*/;
assign _51667_ = ~Q[6] /*10951*/;
assign _51666_ = _51667_ & D[24] /*10950*/;
assign _51669_ = _51033_ & _51666_ /*10945*/;
assign _51670_ = _51033_ ^ _51666_ /*10948*/;
assign _51671_ = _51662_ & _51670_ /*10946*/;
assign _51481_ = _51662_ ^ _51670_ /*10947*/;
assign _51668_ = _51669_ | _51671_ /*10944*/;
assign _51673_ = ~Q[6] /*10943*/;
assign _51672_ = _51673_ & D[25] /*10942*/;
assign _51675_ = _51034_ & _51672_ /*10937*/;
assign _51676_ = _51034_ ^ _51672_ /*10940*/;
assign _51677_ = _51668_ & _51676_ /*10938*/;
assign _51482_ = _51668_ ^ _51676_ /*10939*/;
assign _51674_ = _51675_ | _51677_ /*10936*/;
assign _51679_ = ~Q[6] /*10935*/;
assign _51678_ = _51679_ & D[26] /*10934*/;
assign _51681_ = _51035_ & _51678_ /*10929*/;
assign _51682_ = _51035_ ^ _51678_ /*10932*/;
assign _51683_ = _51674_ & _51682_ /*10930*/;
assign _51483_ = _51674_ ^ _51682_ /*10931*/;
assign _51680_ = _51681_ | _51683_ /*10928*/;
assign _51685_ = ~Q[6] /*10927*/;
assign _51684_ = _51685_ & D[27] /*10926*/;
assign _51687_ = _51036_ & _51684_ /*10921*/;
assign _51688_ = _51036_ ^ _51684_ /*10924*/;
assign _51689_ = _51680_ & _51688_ /*10922*/;
assign _51484_ = _51680_ ^ _51688_ /*10923*/;
assign _51686_ = _51687_ | _51689_ /*10920*/;
assign _51691_ = ~Q[6] /*10919*/;
assign _51690_ = _51691_ & D[28] /*10918*/;
assign _51693_ = _51037_ & _51690_ /*10913*/;
assign _51694_ = _51037_ ^ _51690_ /*10916*/;
assign _51695_ = _51686_ & _51694_ /*10914*/;
assign _51485_ = _51686_ ^ _51694_ /*10915*/;
assign _51692_ = _51693_ | _51695_ /*10912*/;
assign _51697_ = ~Q[6] /*10911*/;
assign _51696_ = _51697_ & D[29] /*10910*/;
assign _51699_ = _51038_ & _51696_ /*10905*/;
assign _51700_ = _51038_ ^ _51696_ /*10908*/;
assign _51701_ = _51692_ & _51700_ /*10906*/;
assign _51486_ = _51692_ ^ _51700_ /*10907*/;
assign _51698_ = _51699_ | _51701_ /*10904*/;
assign _51703_ = ~Q[6] /*10903*/;
assign _51702_ = _51703_ & D[30] /*10902*/;
assign _51705_ = _51039_ & _51702_ /*10897*/;
assign _51706_ = _51039_ ^ _51702_ /*10900*/;
assign _51707_ = _51698_ & _51706_ /*10898*/;
assign _51487_ = _51698_ ^ _51706_ /*10899*/;
assign _51704_ = _51705_ | _51707_ /*10896*/;
assign _51709_ = ~Q[6] /*10895*/;
assign _51708_ = _51709_ & D[31] /*10894*/;
assign _51711_ = _51040_ & _51708_ /*10889*/;
assign _51712_ = _51040_ ^ _51708_ /*10892*/;
assign _51713_ = _51704_ & _51712_ /*10890*/;
assign _51488_ = _51704_ ^ _51712_ /*10891*/;
assign _51710_ = _51711_ | _51713_ /*10888*/;
assign _51715_ = ~Q[6] /*10887*/;
assign _51714_ = _51715_ & D[32] /*10886*/;
assign _51717_ = _51041_ & _51714_ /*10881*/;
assign _51718_ = _51041_ ^ _51714_ /*10884*/;
assign _51719_ = _51710_ & _51718_ /*10882*/;
assign _51489_ = _51710_ ^ _51718_ /*10883*/;
assign _51716_ = _51717_ | _51719_ /*10880*/;
assign _51721_ = ~Q[6] /*10879*/;
assign _51720_ = _51721_ & D[33] /*10878*/;
assign _51723_ = _51042_ & _51720_ /*10873*/;
assign _51724_ = _51042_ ^ _51720_ /*10876*/;
assign _51725_ = _51716_ & _51724_ /*10874*/;
assign _51490_ = _51716_ ^ _51724_ /*10875*/;
assign _51722_ = _51723_ | _51725_ /*10872*/;
assign _51727_ = ~Q[6] /*10871*/;
assign _51726_ = _51727_ & D[34] /*10870*/;
assign _51729_ = _51043_ & _51726_ /*10865*/;
assign _51730_ = _51043_ ^ _51726_ /*10868*/;
assign _51731_ = _51722_ & _51730_ /*10866*/;
assign _51491_ = _51722_ ^ _51730_ /*10867*/;
assign _51728_ = _51729_ | _51731_ /*10864*/;
assign _51733_ = ~Q[6] /*10863*/;
assign _51732_ = _51733_ & D[35] /*10862*/;
assign _51735_ = _51044_ & _51732_ /*10857*/;
assign _51736_ = _51044_ ^ _51732_ /*10860*/;
assign _51737_ = _51728_ & _51736_ /*10858*/;
assign _51492_ = _51728_ ^ _51736_ /*10859*/;
assign _51734_ = _51735_ | _51737_ /*10856*/;
assign _51739_ = ~Q[6] /*10855*/;
assign _51738_ = _51739_ & D[36] /*10854*/;
assign _51741_ = _51045_ & _51738_ /*10849*/;
assign _51742_ = _51045_ ^ _51738_ /*10852*/;
assign _51743_ = _51734_ & _51742_ /*10850*/;
assign _51493_ = _51734_ ^ _51742_ /*10851*/;
assign _51740_ = _51741_ | _51743_ /*10848*/;
assign _51745_ = ~Q[6] /*10847*/;
assign _51744_ = _51745_ & D[37] /*10846*/;
assign _51747_ = _51046_ & _51744_ /*10841*/;
assign _51748_ = _51046_ ^ _51744_ /*10844*/;
assign _51749_ = _51740_ & _51748_ /*10842*/;
assign _51494_ = _51740_ ^ _51748_ /*10843*/;
assign _51746_ = _51747_ | _51749_ /*10840*/;
assign _51751_ = ~Q[6] /*10839*/;
assign _51750_ = _51751_ & D[38] /*10838*/;
assign _51753_ = _51047_ & _51750_ /*10833*/;
assign _51754_ = _51047_ ^ _51750_ /*10836*/;
assign _51755_ = _51746_ & _51754_ /*10834*/;
assign _51495_ = _51746_ ^ _51754_ /*10835*/;
assign _51752_ = _51753_ | _51755_ /*10832*/;
assign _51757_ = ~Q[6] /*10831*/;
assign _51756_ = _51757_ & D[39] /*10830*/;
assign _51759_ = _51048_ & _51756_ /*10825*/;
assign _51760_ = _51048_ ^ _51756_ /*10828*/;
assign _51761_ = _51752_ & _51760_ /*10826*/;
assign _51496_ = _51752_ ^ _51760_ /*10827*/;
assign _51758_ = _51759_ | _51761_ /*10824*/;
assign _51763_ = ~Q[6] /*10823*/;
assign _51762_ = _51763_ & D[40] /*10822*/;
assign _51765_ = _51049_ & _51762_ /*10817*/;
assign _51766_ = _51049_ ^ _51762_ /*10820*/;
assign _51767_ = _51758_ & _51766_ /*10818*/;
assign _51497_ = _51758_ ^ _51766_ /*10819*/;
assign _51764_ = _51765_ | _51767_ /*10816*/;
assign _51769_ = ~Q[6] /*10815*/;
assign _51768_ = _51769_ & D[41] /*10814*/;
assign _51771_ = _51050_ & _51768_ /*10809*/;
assign _51772_ = _51050_ ^ _51768_ /*10812*/;
assign _51773_ = _51764_ & _51772_ /*10810*/;
assign _51498_ = _51764_ ^ _51772_ /*10811*/;
assign _51770_ = _51771_ | _51773_ /*10808*/;
assign _51775_ = ~Q[6] /*10807*/;
assign _51774_ = _51775_ & D[42] /*10806*/;
assign _51777_ = _51051_ & _51774_ /*10801*/;
assign _51778_ = _51051_ ^ _51774_ /*10804*/;
assign _51779_ = _51770_ & _51778_ /*10802*/;
assign _51499_ = _51770_ ^ _51778_ /*10803*/;
assign _51776_ = _51777_ | _51779_ /*10800*/;
assign _51781_ = ~Q[6] /*10799*/;
assign _51780_ = _51781_ & D[43] /*10798*/;
assign _51783_ = _51052_ & _51780_ /*10793*/;
assign _51784_ = _51052_ ^ _51780_ /*10796*/;
assign _51785_ = _51776_ & _51784_ /*10794*/;
assign _51500_ = _51776_ ^ _51784_ /*10795*/;
assign _51782_ = _51783_ | _51785_ /*10792*/;
assign _51787_ = ~Q[6] /*10791*/;
assign _51786_ = _51787_ & D[44] /*10790*/;
assign _51789_ = _51053_ & _51786_ /*10785*/;
assign _51790_ = _51053_ ^ _51786_ /*10788*/;
assign _51791_ = _51782_ & _51790_ /*10786*/;
assign _51501_ = _51782_ ^ _51790_ /*10787*/;
assign _51788_ = _51789_ | _51791_ /*10784*/;
assign _51793_ = ~Q[6] /*10783*/;
assign _51792_ = _51793_ & D[45] /*10782*/;
assign _51795_ = _51054_ & _51792_ /*10777*/;
assign _51796_ = _51054_ ^ _51792_ /*10780*/;
assign _51797_ = _51788_ & _51796_ /*10778*/;
assign _51502_ = _51788_ ^ _51796_ /*10779*/;
assign _51794_ = _51795_ | _51797_ /*10776*/;
assign _51799_ = ~Q[6] /*10775*/;
assign _51798_ = _51799_ & D[46] /*10774*/;
assign _51801_ = _51055_ & _51798_ /*10769*/;
assign _51802_ = _51055_ ^ _51798_ /*10772*/;
assign _51803_ = _51794_ & _51802_ /*10770*/;
assign _51503_ = _51794_ ^ _51802_ /*10771*/;
assign _51800_ = _51801_ | _51803_ /*10768*/;
assign _51805_ = ~Q[6] /*10767*/;
assign _51804_ = _51805_ & D[47] /*10766*/;
assign _51807_ = _51056_ & _51804_ /*10761*/;
assign _51808_ = _51056_ ^ _51804_ /*10764*/;
assign _51809_ = _51800_ & _51808_ /*10762*/;
assign _51504_ = _51800_ ^ _51808_ /*10763*/;
assign _51806_ = _51807_ | _51809_ /*10760*/;
assign _51811_ = ~Q[6] /*10759*/;
assign _51810_ = _51811_ & D[48] /*10758*/;
assign _51813_ = _51057_ & _51810_ /*10753*/;
assign _51814_ = _51057_ ^ _51810_ /*10756*/;
assign _51815_ = _51806_ & _51814_ /*10754*/;
assign _51505_ = _51806_ ^ _51814_ /*10755*/;
assign _51812_ = _51813_ | _51815_ /*10752*/;
assign _51817_ = ~Q[6] /*10751*/;
assign _51816_ = _51817_ & D[49] /*10750*/;
assign _51819_ = _51058_ & _51816_ /*10745*/;
assign _51820_ = _51058_ ^ _51816_ /*10748*/;
assign _51821_ = _51812_ & _51820_ /*10746*/;
assign _51506_ = _51812_ ^ _51820_ /*10747*/;
assign _51818_ = _51819_ | _51821_ /*10744*/;
assign _51823_ = ~Q[6] /*10743*/;
assign _51822_ = _51823_ & D[50] /*10742*/;
assign _51825_ = _51059_ & _51822_ /*10737*/;
assign _51826_ = _51059_ ^ _51822_ /*10740*/;
assign _51827_ = _51818_ & _51826_ /*10738*/;
assign _51507_ = _51818_ ^ _51826_ /*10739*/;
assign _51824_ = _51825_ | _51827_ /*10736*/;
assign _51829_ = ~Q[6] /*10735*/;
assign _51828_ = _51829_ & D[51] /*10734*/;
assign _51831_ = _51060_ & _51828_ /*10729*/;
assign _51832_ = _51060_ ^ _51828_ /*10732*/;
assign _51833_ = _51824_ & _51832_ /*10730*/;
assign _51508_ = _51824_ ^ _51832_ /*10731*/;
assign _51830_ = _51831_ | _51833_ /*10728*/;
assign _51835_ = ~Q[6] /*10727*/;
assign _51834_ = _51835_ & D[52] /*10726*/;
assign _51837_ = _51061_ & _51834_ /*10721*/;
assign _51838_ = _51061_ ^ _51834_ /*10724*/;
assign _51839_ = _51830_ & _51838_ /*10722*/;
assign _51509_ = _51830_ ^ _51838_ /*10723*/;
assign _51836_ = _51837_ | _51839_ /*10720*/;
assign _51841_ = ~Q[6] /*10719*/;
assign _51840_ = _51841_ & D[53] /*10718*/;
assign _51843_ = _51062_ & _51840_ /*10713*/;
assign _51844_ = _51062_ ^ _51840_ /*10716*/;
assign _51845_ = _51836_ & _51844_ /*10714*/;
assign _51510_ = _51836_ ^ _51844_ /*10715*/;
assign _51842_ = _51843_ | _51845_ /*10712*/;
assign _51847_ = ~Q[6] /*10711*/;
assign _51846_ = _51847_ & D[54] /*10710*/;
assign _51849_ = _51063_ & _51846_ /*10705*/;
assign _51850_ = _51063_ ^ _51846_ /*10708*/;
assign _51851_ = _51842_ & _51850_ /*10706*/;
assign _51511_ = _51842_ ^ _51850_ /*10707*/;
assign _51848_ = _51849_ | _51851_ /*10704*/;
assign _51853_ = ~Q[6] /*10703*/;
assign _51852_ = _51853_ & D[55] /*10702*/;
assign _51855_ = _51064_ & _51852_ /*10697*/;
assign _51856_ = _51064_ ^ _51852_ /*10700*/;
assign _51857_ = _51848_ & _51856_ /*10698*/;
assign _51512_ = _51848_ ^ _51856_ /*10699*/;
assign _51854_ = _51855_ | _51857_ /*10696*/;
assign _51859_ = ~Q[6] /*10695*/;
assign _51858_ = _51859_ & D[56] /*10694*/;
assign _51861_ = _51065_ & _51858_ /*10689*/;
assign _51862_ = _51065_ ^ _51858_ /*10692*/;
assign _51863_ = _51854_ & _51862_ /*10690*/;
assign _51513_ = _51854_ ^ _51862_ /*10691*/;
assign _51860_ = _51861_ | _51863_ /*10688*/;
assign _51865_ = ~Q[6] /*10687*/;
assign _51864_ = _51865_ & D[57] /*10686*/;
assign _51867_ = _51066_ & _51864_ /*10681*/;
assign _51868_ = _51066_ ^ _51864_ /*10684*/;
assign _51869_ = _51860_ & _51868_ /*10682*/;
assign _51514_ = _51860_ ^ _51868_ /*10683*/;
assign _51866_ = _51867_ | _51869_ /*10680*/;
assign _51871_ = ~Q[6] /*10679*/;
assign _51870_ = _51871_ & D[58] /*10678*/;
assign _51873_ = _51067_ & _51870_ /*10673*/;
assign _51874_ = _51067_ ^ _51870_ /*10676*/;
assign _51875_ = _51866_ & _51874_ /*10674*/;
assign _51515_ = _51866_ ^ _51874_ /*10675*/;
assign _51872_ = _51873_ | _51875_ /*10672*/;
assign _51877_ = ~Q[6] /*10671*/;
assign _51876_ = _51877_ & D[59] /*10670*/;
assign _51879_ = _51068_ & _51876_ /*10665*/;
assign _51880_ = _51068_ ^ _51876_ /*10668*/;
assign _51881_ = _51872_ & _51880_ /*10666*/;
assign _51516_ = _51872_ ^ _51880_ /*10667*/;
assign _51878_ = _51879_ | _51881_ /*10664*/;
assign _51883_ = ~Q[6] /*10663*/;
assign _51882_ = _51883_ & D[60] /*10662*/;
assign _51885_ = _51069_ & _51882_ /*10657*/;
assign _51886_ = _51069_ ^ _51882_ /*10660*/;
assign _51887_ = _51878_ & _51886_ /*10658*/;
assign _51517_ = _51878_ ^ _51886_ /*10659*/;
assign _51884_ = _51885_ | _51887_ /*10656*/;
assign _51889_ = ~Q[6] /*10655*/;
assign _51888_ = _51889_ & D[61] /*10654*/;
assign _51891_ = _51070_ & _51888_ /*10649*/;
assign _51892_ = _51070_ ^ _51888_ /*10652*/;
assign _51893_ = _51884_ & _51892_ /*10650*/;
assign _51518_ = _51884_ ^ _51892_ /*10651*/;
assign _51890_ = _51891_ | _51893_ /*10648*/;
assign _51895_ = ~Q[6] /*10647*/;
assign _51894_ = _51895_ & D[62] /*10646*/;
assign _51897_ = _51071_ & _51894_ /*10641*/;
assign _51898_ = _51071_ ^ _51894_ /*10644*/;
assign _51899_ = _51890_ & _51898_ /*10642*/;
assign _51519_ = _51890_ ^ _51898_ /*10643*/;
assign _51896_ = _51897_ | _51899_ /*10640*/;
assign _51901_ = ~Q[6] /*10639*/;
assign _51900_ = _51901_ & zeroWire /*10638*/;
assign _51902_ = _51072_ ^ _51900_ /*10636*/;
assign _51520_ = _51902_ ^ _51896_ /*10635*/;
assign _51973_ = ~D[0] /*10381*/;
assign _51970_ = R_0[5] & _51973_ /*10377*/;
assign _51971_ = R_0[5] ^ _51973_ /*10380*/;
assign _51972_ = oneWire & _51971_ /*10378*/;
assign _51905_ = oneWire ^ _51971_ /*10379*/;
assign _51969_ = _51970_ | _51972_ /*10376*/;
assign _51978_ = ~D[1] /*10375*/;
assign _51975_ = _51457_ & _51978_ /*10371*/;
assign _51976_ = _51457_ ^ _51978_ /*10374*/;
assign _51977_ = _51969_ & _51976_ /*10372*/;
assign _51906_ = _51969_ ^ _51976_ /*10373*/;
assign _51974_ = _51975_ | _51977_ /*10370*/;
assign _51983_ = ~D[2] /*10369*/;
assign _51980_ = _51458_ & _51983_ /*10365*/;
assign _51981_ = _51458_ ^ _51983_ /*10368*/;
assign _51982_ = _51974_ & _51981_ /*10366*/;
assign _51907_ = _51974_ ^ _51981_ /*10367*/;
assign _51979_ = _51980_ | _51982_ /*10364*/;
assign _51988_ = ~D[3] /*10363*/;
assign _51985_ = _51459_ & _51988_ /*10359*/;
assign _51986_ = _51459_ ^ _51988_ /*10362*/;
assign _51987_ = _51979_ & _51986_ /*10360*/;
assign _51908_ = _51979_ ^ _51986_ /*10361*/;
assign _51984_ = _51985_ | _51987_ /*10358*/;
assign _51993_ = ~D[4] /*10357*/;
assign _51990_ = _51460_ & _51993_ /*10353*/;
assign _51991_ = _51460_ ^ _51993_ /*10356*/;
assign _51992_ = _51984_ & _51991_ /*10354*/;
assign _51909_ = _51984_ ^ _51991_ /*10355*/;
assign _51989_ = _51990_ | _51992_ /*10352*/;
assign _51998_ = ~D[5] /*10351*/;
assign _51995_ = _51461_ & _51998_ /*10347*/;
assign _51996_ = _51461_ ^ _51998_ /*10350*/;
assign _51997_ = _51989_ & _51996_ /*10348*/;
assign _51910_ = _51989_ ^ _51996_ /*10349*/;
assign _51994_ = _51995_ | _51997_ /*10346*/;
assign _52003_ = ~D[6] /*10345*/;
assign _52000_ = _51462_ & _52003_ /*10341*/;
assign _52001_ = _51462_ ^ _52003_ /*10344*/;
assign _52002_ = _51994_ & _52001_ /*10342*/;
assign _51911_ = _51994_ ^ _52001_ /*10343*/;
assign _51999_ = _52000_ | _52002_ /*10340*/;
assign _52008_ = ~D[7] /*10339*/;
assign _52005_ = _51463_ & _52008_ /*10335*/;
assign _52006_ = _51463_ ^ _52008_ /*10338*/;
assign _52007_ = _51999_ & _52006_ /*10336*/;
assign _51912_ = _51999_ ^ _52006_ /*10337*/;
assign _52004_ = _52005_ | _52007_ /*10334*/;
assign _52013_ = ~D[8] /*10333*/;
assign _52010_ = _51464_ & _52013_ /*10329*/;
assign _52011_ = _51464_ ^ _52013_ /*10332*/;
assign _52012_ = _52004_ & _52011_ /*10330*/;
assign _51913_ = _52004_ ^ _52011_ /*10331*/;
assign _52009_ = _52010_ | _52012_ /*10328*/;
assign _52018_ = ~D[9] /*10327*/;
assign _52015_ = _51465_ & _52018_ /*10323*/;
assign _52016_ = _51465_ ^ _52018_ /*10326*/;
assign _52017_ = _52009_ & _52016_ /*10324*/;
assign _51914_ = _52009_ ^ _52016_ /*10325*/;
assign _52014_ = _52015_ | _52017_ /*10322*/;
assign _52023_ = ~D[10] /*10321*/;
assign _52020_ = _51466_ & _52023_ /*10317*/;
assign _52021_ = _51466_ ^ _52023_ /*10320*/;
assign _52022_ = _52014_ & _52021_ /*10318*/;
assign _51915_ = _52014_ ^ _52021_ /*10319*/;
assign _52019_ = _52020_ | _52022_ /*10316*/;
assign _52028_ = ~D[11] /*10315*/;
assign _52025_ = _51467_ & _52028_ /*10311*/;
assign _52026_ = _51467_ ^ _52028_ /*10314*/;
assign _52027_ = _52019_ & _52026_ /*10312*/;
assign _51916_ = _52019_ ^ _52026_ /*10313*/;
assign _52024_ = _52025_ | _52027_ /*10310*/;
assign _52033_ = ~D[12] /*10309*/;
assign _52030_ = _51468_ & _52033_ /*10305*/;
assign _52031_ = _51468_ ^ _52033_ /*10308*/;
assign _52032_ = _52024_ & _52031_ /*10306*/;
assign _51917_ = _52024_ ^ _52031_ /*10307*/;
assign _52029_ = _52030_ | _52032_ /*10304*/;
assign _52038_ = ~D[13] /*10303*/;
assign _52035_ = _51469_ & _52038_ /*10299*/;
assign _52036_ = _51469_ ^ _52038_ /*10302*/;
assign _52037_ = _52029_ & _52036_ /*10300*/;
assign _51918_ = _52029_ ^ _52036_ /*10301*/;
assign _52034_ = _52035_ | _52037_ /*10298*/;
assign _52043_ = ~D[14] /*10297*/;
assign _52040_ = _51470_ & _52043_ /*10293*/;
assign _52041_ = _51470_ ^ _52043_ /*10296*/;
assign _52042_ = _52034_ & _52041_ /*10294*/;
assign _51919_ = _52034_ ^ _52041_ /*10295*/;
assign _52039_ = _52040_ | _52042_ /*10292*/;
assign _52048_ = ~D[15] /*10291*/;
assign _52045_ = _51471_ & _52048_ /*10287*/;
assign _52046_ = _51471_ ^ _52048_ /*10290*/;
assign _52047_ = _52039_ & _52046_ /*10288*/;
assign _51920_ = _52039_ ^ _52046_ /*10289*/;
assign _52044_ = _52045_ | _52047_ /*10286*/;
assign _52053_ = ~D[16] /*10285*/;
assign _52050_ = _51472_ & _52053_ /*10281*/;
assign _52051_ = _51472_ ^ _52053_ /*10284*/;
assign _52052_ = _52044_ & _52051_ /*10282*/;
assign _51921_ = _52044_ ^ _52051_ /*10283*/;
assign _52049_ = _52050_ | _52052_ /*10280*/;
assign _52058_ = ~D[17] /*10279*/;
assign _52055_ = _51473_ & _52058_ /*10275*/;
assign _52056_ = _51473_ ^ _52058_ /*10278*/;
assign _52057_ = _52049_ & _52056_ /*10276*/;
assign _51922_ = _52049_ ^ _52056_ /*10277*/;
assign _52054_ = _52055_ | _52057_ /*10274*/;
assign _52063_ = ~D[18] /*10273*/;
assign _52060_ = _51474_ & _52063_ /*10269*/;
assign _52061_ = _51474_ ^ _52063_ /*10272*/;
assign _52062_ = _52054_ & _52061_ /*10270*/;
assign _51923_ = _52054_ ^ _52061_ /*10271*/;
assign _52059_ = _52060_ | _52062_ /*10268*/;
assign _52068_ = ~D[19] /*10267*/;
assign _52065_ = _51475_ & _52068_ /*10263*/;
assign _52066_ = _51475_ ^ _52068_ /*10266*/;
assign _52067_ = _52059_ & _52066_ /*10264*/;
assign _51924_ = _52059_ ^ _52066_ /*10265*/;
assign _52064_ = _52065_ | _52067_ /*10262*/;
assign _52073_ = ~D[20] /*10261*/;
assign _52070_ = _51476_ & _52073_ /*10257*/;
assign _52071_ = _51476_ ^ _52073_ /*10260*/;
assign _52072_ = _52064_ & _52071_ /*10258*/;
assign _51925_ = _52064_ ^ _52071_ /*10259*/;
assign _52069_ = _52070_ | _52072_ /*10256*/;
assign _52078_ = ~D[21] /*10255*/;
assign _52075_ = _51477_ & _52078_ /*10251*/;
assign _52076_ = _51477_ ^ _52078_ /*10254*/;
assign _52077_ = _52069_ & _52076_ /*10252*/;
assign _51926_ = _52069_ ^ _52076_ /*10253*/;
assign _52074_ = _52075_ | _52077_ /*10250*/;
assign _52083_ = ~D[22] /*10249*/;
assign _52080_ = _51478_ & _52083_ /*10245*/;
assign _52081_ = _51478_ ^ _52083_ /*10248*/;
assign _52082_ = _52074_ & _52081_ /*10246*/;
assign _51927_ = _52074_ ^ _52081_ /*10247*/;
assign _52079_ = _52080_ | _52082_ /*10244*/;
assign _52088_ = ~D[23] /*10243*/;
assign _52085_ = _51479_ & _52088_ /*10239*/;
assign _52086_ = _51479_ ^ _52088_ /*10242*/;
assign _52087_ = _52079_ & _52086_ /*10240*/;
assign _51928_ = _52079_ ^ _52086_ /*10241*/;
assign _52084_ = _52085_ | _52087_ /*10238*/;
assign _52093_ = ~D[24] /*10237*/;
assign _52090_ = _51480_ & _52093_ /*10233*/;
assign _52091_ = _51480_ ^ _52093_ /*10236*/;
assign _52092_ = _52084_ & _52091_ /*10234*/;
assign _51929_ = _52084_ ^ _52091_ /*10235*/;
assign _52089_ = _52090_ | _52092_ /*10232*/;
assign _52098_ = ~D[25] /*10231*/;
assign _52095_ = _51481_ & _52098_ /*10227*/;
assign _52096_ = _51481_ ^ _52098_ /*10230*/;
assign _52097_ = _52089_ & _52096_ /*10228*/;
assign _51930_ = _52089_ ^ _52096_ /*10229*/;
assign _52094_ = _52095_ | _52097_ /*10226*/;
assign _52103_ = ~D[26] /*10225*/;
assign _52100_ = _51482_ & _52103_ /*10221*/;
assign _52101_ = _51482_ ^ _52103_ /*10224*/;
assign _52102_ = _52094_ & _52101_ /*10222*/;
assign _51931_ = _52094_ ^ _52101_ /*10223*/;
assign _52099_ = _52100_ | _52102_ /*10220*/;
assign _52108_ = ~D[27] /*10219*/;
assign _52105_ = _51483_ & _52108_ /*10215*/;
assign _52106_ = _51483_ ^ _52108_ /*10218*/;
assign _52107_ = _52099_ & _52106_ /*10216*/;
assign _51932_ = _52099_ ^ _52106_ /*10217*/;
assign _52104_ = _52105_ | _52107_ /*10214*/;
assign _52113_ = ~D[28] /*10213*/;
assign _52110_ = _51484_ & _52113_ /*10209*/;
assign _52111_ = _51484_ ^ _52113_ /*10212*/;
assign _52112_ = _52104_ & _52111_ /*10210*/;
assign _51933_ = _52104_ ^ _52111_ /*10211*/;
assign _52109_ = _52110_ | _52112_ /*10208*/;
assign _52118_ = ~D[29] /*10207*/;
assign _52115_ = _51485_ & _52118_ /*10203*/;
assign _52116_ = _51485_ ^ _52118_ /*10206*/;
assign _52117_ = _52109_ & _52116_ /*10204*/;
assign _51934_ = _52109_ ^ _52116_ /*10205*/;
assign _52114_ = _52115_ | _52117_ /*10202*/;
assign _52123_ = ~D[30] /*10201*/;
assign _52120_ = _51486_ & _52123_ /*10197*/;
assign _52121_ = _51486_ ^ _52123_ /*10200*/;
assign _52122_ = _52114_ & _52121_ /*10198*/;
assign _51935_ = _52114_ ^ _52121_ /*10199*/;
assign _52119_ = _52120_ | _52122_ /*10196*/;
assign _52128_ = ~D[31] /*10195*/;
assign _52125_ = _51487_ & _52128_ /*10191*/;
assign _52126_ = _51487_ ^ _52128_ /*10194*/;
assign _52127_ = _52119_ & _52126_ /*10192*/;
assign _51936_ = _52119_ ^ _52126_ /*10193*/;
assign _52124_ = _52125_ | _52127_ /*10190*/;
assign _52133_ = ~D[32] /*10189*/;
assign _52130_ = _51488_ & _52133_ /*10185*/;
assign _52131_ = _51488_ ^ _52133_ /*10188*/;
assign _52132_ = _52124_ & _52131_ /*10186*/;
assign _51937_ = _52124_ ^ _52131_ /*10187*/;
assign _52129_ = _52130_ | _52132_ /*10184*/;
assign _52138_ = ~D[33] /*10183*/;
assign _52135_ = _51489_ & _52138_ /*10179*/;
assign _52136_ = _51489_ ^ _52138_ /*10182*/;
assign _52137_ = _52129_ & _52136_ /*10180*/;
assign _51938_ = _52129_ ^ _52136_ /*10181*/;
assign _52134_ = _52135_ | _52137_ /*10178*/;
assign _52143_ = ~D[34] /*10177*/;
assign _52140_ = _51490_ & _52143_ /*10173*/;
assign _52141_ = _51490_ ^ _52143_ /*10176*/;
assign _52142_ = _52134_ & _52141_ /*10174*/;
assign _51939_ = _52134_ ^ _52141_ /*10175*/;
assign _52139_ = _52140_ | _52142_ /*10172*/;
assign _52148_ = ~D[35] /*10171*/;
assign _52145_ = _51491_ & _52148_ /*10167*/;
assign _52146_ = _51491_ ^ _52148_ /*10170*/;
assign _52147_ = _52139_ & _52146_ /*10168*/;
assign _51940_ = _52139_ ^ _52146_ /*10169*/;
assign _52144_ = _52145_ | _52147_ /*10166*/;
assign _52153_ = ~D[36] /*10165*/;
assign _52150_ = _51492_ & _52153_ /*10161*/;
assign _52151_ = _51492_ ^ _52153_ /*10164*/;
assign _52152_ = _52144_ & _52151_ /*10162*/;
assign _51941_ = _52144_ ^ _52151_ /*10163*/;
assign _52149_ = _52150_ | _52152_ /*10160*/;
assign _52158_ = ~D[37] /*10159*/;
assign _52155_ = _51493_ & _52158_ /*10155*/;
assign _52156_ = _51493_ ^ _52158_ /*10158*/;
assign _52157_ = _52149_ & _52156_ /*10156*/;
assign _51942_ = _52149_ ^ _52156_ /*10157*/;
assign _52154_ = _52155_ | _52157_ /*10154*/;
assign _52163_ = ~D[38] /*10153*/;
assign _52160_ = _51494_ & _52163_ /*10149*/;
assign _52161_ = _51494_ ^ _52163_ /*10152*/;
assign _52162_ = _52154_ & _52161_ /*10150*/;
assign _51943_ = _52154_ ^ _52161_ /*10151*/;
assign _52159_ = _52160_ | _52162_ /*10148*/;
assign _52168_ = ~D[39] /*10147*/;
assign _52165_ = _51495_ & _52168_ /*10143*/;
assign _52166_ = _51495_ ^ _52168_ /*10146*/;
assign _52167_ = _52159_ & _52166_ /*10144*/;
assign _51944_ = _52159_ ^ _52166_ /*10145*/;
assign _52164_ = _52165_ | _52167_ /*10142*/;
assign _52173_ = ~D[40] /*10141*/;
assign _52170_ = _51496_ & _52173_ /*10137*/;
assign _52171_ = _51496_ ^ _52173_ /*10140*/;
assign _52172_ = _52164_ & _52171_ /*10138*/;
assign _51945_ = _52164_ ^ _52171_ /*10139*/;
assign _52169_ = _52170_ | _52172_ /*10136*/;
assign _52178_ = ~D[41] /*10135*/;
assign _52175_ = _51497_ & _52178_ /*10131*/;
assign _52176_ = _51497_ ^ _52178_ /*10134*/;
assign _52177_ = _52169_ & _52176_ /*10132*/;
assign _51946_ = _52169_ ^ _52176_ /*10133*/;
assign _52174_ = _52175_ | _52177_ /*10130*/;
assign _52183_ = ~D[42] /*10129*/;
assign _52180_ = _51498_ & _52183_ /*10125*/;
assign _52181_ = _51498_ ^ _52183_ /*10128*/;
assign _52182_ = _52174_ & _52181_ /*10126*/;
assign _51947_ = _52174_ ^ _52181_ /*10127*/;
assign _52179_ = _52180_ | _52182_ /*10124*/;
assign _52188_ = ~D[43] /*10123*/;
assign _52185_ = _51499_ & _52188_ /*10119*/;
assign _52186_ = _51499_ ^ _52188_ /*10122*/;
assign _52187_ = _52179_ & _52186_ /*10120*/;
assign _51948_ = _52179_ ^ _52186_ /*10121*/;
assign _52184_ = _52185_ | _52187_ /*10118*/;
assign _52193_ = ~D[44] /*10117*/;
assign _52190_ = _51500_ & _52193_ /*10113*/;
assign _52191_ = _51500_ ^ _52193_ /*10116*/;
assign _52192_ = _52184_ & _52191_ /*10114*/;
assign _51949_ = _52184_ ^ _52191_ /*10115*/;
assign _52189_ = _52190_ | _52192_ /*10112*/;
assign _52198_ = ~D[45] /*10111*/;
assign _52195_ = _51501_ & _52198_ /*10107*/;
assign _52196_ = _51501_ ^ _52198_ /*10110*/;
assign _52197_ = _52189_ & _52196_ /*10108*/;
assign _51950_ = _52189_ ^ _52196_ /*10109*/;
assign _52194_ = _52195_ | _52197_ /*10106*/;
assign _52203_ = ~D[46] /*10105*/;
assign _52200_ = _51502_ & _52203_ /*10101*/;
assign _52201_ = _51502_ ^ _52203_ /*10104*/;
assign _52202_ = _52194_ & _52201_ /*10102*/;
assign _51951_ = _52194_ ^ _52201_ /*10103*/;
assign _52199_ = _52200_ | _52202_ /*10100*/;
assign _52208_ = ~D[47] /*10099*/;
assign _52205_ = _51503_ & _52208_ /*10095*/;
assign _52206_ = _51503_ ^ _52208_ /*10098*/;
assign _52207_ = _52199_ & _52206_ /*10096*/;
assign _51952_ = _52199_ ^ _52206_ /*10097*/;
assign _52204_ = _52205_ | _52207_ /*10094*/;
assign _52213_ = ~D[48] /*10093*/;
assign _52210_ = _51504_ & _52213_ /*10089*/;
assign _52211_ = _51504_ ^ _52213_ /*10092*/;
assign _52212_ = _52204_ & _52211_ /*10090*/;
assign _51953_ = _52204_ ^ _52211_ /*10091*/;
assign _52209_ = _52210_ | _52212_ /*10088*/;
assign _52218_ = ~D[49] /*10087*/;
assign _52215_ = _51505_ & _52218_ /*10083*/;
assign _52216_ = _51505_ ^ _52218_ /*10086*/;
assign _52217_ = _52209_ & _52216_ /*10084*/;
assign _51954_ = _52209_ ^ _52216_ /*10085*/;
assign _52214_ = _52215_ | _52217_ /*10082*/;
assign _52223_ = ~D[50] /*10081*/;
assign _52220_ = _51506_ & _52223_ /*10077*/;
assign _52221_ = _51506_ ^ _52223_ /*10080*/;
assign _52222_ = _52214_ & _52221_ /*10078*/;
assign _51955_ = _52214_ ^ _52221_ /*10079*/;
assign _52219_ = _52220_ | _52222_ /*10076*/;
assign _52228_ = ~D[51] /*10075*/;
assign _52225_ = _51507_ & _52228_ /*10071*/;
assign _52226_ = _51507_ ^ _52228_ /*10074*/;
assign _52227_ = _52219_ & _52226_ /*10072*/;
assign _51956_ = _52219_ ^ _52226_ /*10073*/;
assign _52224_ = _52225_ | _52227_ /*10070*/;
assign _52233_ = ~D[52] /*10069*/;
assign _52230_ = _51508_ & _52233_ /*10065*/;
assign _52231_ = _51508_ ^ _52233_ /*10068*/;
assign _52232_ = _52224_ & _52231_ /*10066*/;
assign _51957_ = _52224_ ^ _52231_ /*10067*/;
assign _52229_ = _52230_ | _52232_ /*10064*/;
assign _52238_ = ~D[53] /*10063*/;
assign _52235_ = _51509_ & _52238_ /*10059*/;
assign _52236_ = _51509_ ^ _52238_ /*10062*/;
assign _52237_ = _52229_ & _52236_ /*10060*/;
assign _51958_ = _52229_ ^ _52236_ /*10061*/;
assign _52234_ = _52235_ | _52237_ /*10058*/;
assign _52243_ = ~D[54] /*10057*/;
assign _52240_ = _51510_ & _52243_ /*10053*/;
assign _52241_ = _51510_ ^ _52243_ /*10056*/;
assign _52242_ = _52234_ & _52241_ /*10054*/;
assign _51959_ = _52234_ ^ _52241_ /*10055*/;
assign _52239_ = _52240_ | _52242_ /*10052*/;
assign _52248_ = ~D[55] /*10051*/;
assign _52245_ = _51511_ & _52248_ /*10047*/;
assign _52246_ = _51511_ ^ _52248_ /*10050*/;
assign _52247_ = _52239_ & _52246_ /*10048*/;
assign _51960_ = _52239_ ^ _52246_ /*10049*/;
assign _52244_ = _52245_ | _52247_ /*10046*/;
assign _52253_ = ~D[56] /*10045*/;
assign _52250_ = _51512_ & _52253_ /*10041*/;
assign _52251_ = _51512_ ^ _52253_ /*10044*/;
assign _52252_ = _52244_ & _52251_ /*10042*/;
assign _51961_ = _52244_ ^ _52251_ /*10043*/;
assign _52249_ = _52250_ | _52252_ /*10040*/;
assign _52258_ = ~D[57] /*10039*/;
assign _52255_ = _51513_ & _52258_ /*10035*/;
assign _52256_ = _51513_ ^ _52258_ /*10038*/;
assign _52257_ = _52249_ & _52256_ /*10036*/;
assign _51962_ = _52249_ ^ _52256_ /*10037*/;
assign _52254_ = _52255_ | _52257_ /*10034*/;
assign _52263_ = ~D[58] /*10033*/;
assign _52260_ = _51514_ & _52263_ /*10029*/;
assign _52261_ = _51514_ ^ _52263_ /*10032*/;
assign _52262_ = _52254_ & _52261_ /*10030*/;
assign _51963_ = _52254_ ^ _52261_ /*10031*/;
assign _52259_ = _52260_ | _52262_ /*10028*/;
assign _52268_ = ~D[59] /*10027*/;
assign _52265_ = _51515_ & _52268_ /*10023*/;
assign _52266_ = _51515_ ^ _52268_ /*10026*/;
assign _52267_ = _52259_ & _52266_ /*10024*/;
assign _51964_ = _52259_ ^ _52266_ /*10025*/;
assign _52264_ = _52265_ | _52267_ /*10022*/;
assign _52273_ = ~D[60] /*10021*/;
assign _52270_ = _51516_ & _52273_ /*10017*/;
assign _52271_ = _51516_ ^ _52273_ /*10020*/;
assign _52272_ = _52264_ & _52271_ /*10018*/;
assign _51965_ = _52264_ ^ _52271_ /*10019*/;
assign _52269_ = _52270_ | _52272_ /*10016*/;
assign _52278_ = ~D[61] /*10015*/;
assign _52275_ = _51517_ & _52278_ /*10011*/;
assign _52276_ = _51517_ ^ _52278_ /*10014*/;
assign _52277_ = _52269_ & _52276_ /*10012*/;
assign _51966_ = _52269_ ^ _52276_ /*10013*/;
assign _52274_ = _52275_ | _52277_ /*10010*/;
assign _52283_ = ~D[62] /*10009*/;
assign _52280_ = _51518_ & _52283_ /*10005*/;
assign _52281_ = _51518_ ^ _52283_ /*10008*/;
assign _52282_ = _52274_ & _52281_ /*10006*/;
assign _51967_ = _52274_ ^ _52281_ /*10007*/;
assign _52279_ = _52280_ | _52282_ /*10004*/;
assign _52284_ = _51519_ & oneWire /*9999*/;
assign _52285_ = _51519_ ^ oneWire /*10002*/;
assign _52286_ = _52279_ & _52285_ /*10000*/;
assign _51968_ = _52279_ ^ _52285_ /*10001*/;
assign Q[5] = _52284_ | _52286_ /*9998*/;
assign _52419_ = ~Q[5] /*9613*/;
assign _52418_ = _52419_ & D[0] /*9612*/;
assign _52421_ = _51905_ & _52418_ /*9607*/;
assign _52422_ = _51905_ ^ _52418_ /*9610*/;
assign _52423_ = zeroWire & _52422_ /*9608*/;
assign _52353_ = zeroWire ^ _52422_ /*9609*/;
assign _52420_ = _52421_ | _52423_ /*9606*/;
assign _52425_ = ~Q[5] /*9605*/;
assign _52424_ = _52425_ & D[1] /*9604*/;
assign _52427_ = _51906_ & _52424_ /*9599*/;
assign _52428_ = _51906_ ^ _52424_ /*9602*/;
assign _52429_ = _52420_ & _52428_ /*9600*/;
assign _52354_ = _52420_ ^ _52428_ /*9601*/;
assign _52426_ = _52427_ | _52429_ /*9598*/;
assign _52431_ = ~Q[5] /*9597*/;
assign _52430_ = _52431_ & D[2] /*9596*/;
assign _52433_ = _51907_ & _52430_ /*9591*/;
assign _52434_ = _51907_ ^ _52430_ /*9594*/;
assign _52435_ = _52426_ & _52434_ /*9592*/;
assign _52355_ = _52426_ ^ _52434_ /*9593*/;
assign _52432_ = _52433_ | _52435_ /*9590*/;
assign _52437_ = ~Q[5] /*9589*/;
assign _52436_ = _52437_ & D[3] /*9588*/;
assign _52439_ = _51908_ & _52436_ /*9583*/;
assign _52440_ = _51908_ ^ _52436_ /*9586*/;
assign _52441_ = _52432_ & _52440_ /*9584*/;
assign _52356_ = _52432_ ^ _52440_ /*9585*/;
assign _52438_ = _52439_ | _52441_ /*9582*/;
assign _52443_ = ~Q[5] /*9581*/;
assign _52442_ = _52443_ & D[4] /*9580*/;
assign _52445_ = _51909_ & _52442_ /*9575*/;
assign _52446_ = _51909_ ^ _52442_ /*9578*/;
assign _52447_ = _52438_ & _52446_ /*9576*/;
assign _52357_ = _52438_ ^ _52446_ /*9577*/;
assign _52444_ = _52445_ | _52447_ /*9574*/;
assign _52449_ = ~Q[5] /*9573*/;
assign _52448_ = _52449_ & D[5] /*9572*/;
assign _52451_ = _51910_ & _52448_ /*9567*/;
assign _52452_ = _51910_ ^ _52448_ /*9570*/;
assign _52453_ = _52444_ & _52452_ /*9568*/;
assign _52358_ = _52444_ ^ _52452_ /*9569*/;
assign _52450_ = _52451_ | _52453_ /*9566*/;
assign _52455_ = ~Q[5] /*9565*/;
assign _52454_ = _52455_ & D[6] /*9564*/;
assign _52457_ = _51911_ & _52454_ /*9559*/;
assign _52458_ = _51911_ ^ _52454_ /*9562*/;
assign _52459_ = _52450_ & _52458_ /*9560*/;
assign _52359_ = _52450_ ^ _52458_ /*9561*/;
assign _52456_ = _52457_ | _52459_ /*9558*/;
assign _52461_ = ~Q[5] /*9557*/;
assign _52460_ = _52461_ & D[7] /*9556*/;
assign _52463_ = _51912_ & _52460_ /*9551*/;
assign _52464_ = _51912_ ^ _52460_ /*9554*/;
assign _52465_ = _52456_ & _52464_ /*9552*/;
assign _52360_ = _52456_ ^ _52464_ /*9553*/;
assign _52462_ = _52463_ | _52465_ /*9550*/;
assign _52467_ = ~Q[5] /*9549*/;
assign _52466_ = _52467_ & D[8] /*9548*/;
assign _52469_ = _51913_ & _52466_ /*9543*/;
assign _52470_ = _51913_ ^ _52466_ /*9546*/;
assign _52471_ = _52462_ & _52470_ /*9544*/;
assign _52361_ = _52462_ ^ _52470_ /*9545*/;
assign _52468_ = _52469_ | _52471_ /*9542*/;
assign _52473_ = ~Q[5] /*9541*/;
assign _52472_ = _52473_ & D[9] /*9540*/;
assign _52475_ = _51914_ & _52472_ /*9535*/;
assign _52476_ = _51914_ ^ _52472_ /*9538*/;
assign _52477_ = _52468_ & _52476_ /*9536*/;
assign _52362_ = _52468_ ^ _52476_ /*9537*/;
assign _52474_ = _52475_ | _52477_ /*9534*/;
assign _52479_ = ~Q[5] /*9533*/;
assign _52478_ = _52479_ & D[10] /*9532*/;
assign _52481_ = _51915_ & _52478_ /*9527*/;
assign _52482_ = _51915_ ^ _52478_ /*9530*/;
assign _52483_ = _52474_ & _52482_ /*9528*/;
assign _52363_ = _52474_ ^ _52482_ /*9529*/;
assign _52480_ = _52481_ | _52483_ /*9526*/;
assign _52485_ = ~Q[5] /*9525*/;
assign _52484_ = _52485_ & D[11] /*9524*/;
assign _52487_ = _51916_ & _52484_ /*9519*/;
assign _52488_ = _51916_ ^ _52484_ /*9522*/;
assign _52489_ = _52480_ & _52488_ /*9520*/;
assign _52364_ = _52480_ ^ _52488_ /*9521*/;
assign _52486_ = _52487_ | _52489_ /*9518*/;
assign _52491_ = ~Q[5] /*9517*/;
assign _52490_ = _52491_ & D[12] /*9516*/;
assign _52493_ = _51917_ & _52490_ /*9511*/;
assign _52494_ = _51917_ ^ _52490_ /*9514*/;
assign _52495_ = _52486_ & _52494_ /*9512*/;
assign _52365_ = _52486_ ^ _52494_ /*9513*/;
assign _52492_ = _52493_ | _52495_ /*9510*/;
assign _52497_ = ~Q[5] /*9509*/;
assign _52496_ = _52497_ & D[13] /*9508*/;
assign _52499_ = _51918_ & _52496_ /*9503*/;
assign _52500_ = _51918_ ^ _52496_ /*9506*/;
assign _52501_ = _52492_ & _52500_ /*9504*/;
assign _52366_ = _52492_ ^ _52500_ /*9505*/;
assign _52498_ = _52499_ | _52501_ /*9502*/;
assign _52503_ = ~Q[5] /*9501*/;
assign _52502_ = _52503_ & D[14] /*9500*/;
assign _52505_ = _51919_ & _52502_ /*9495*/;
assign _52506_ = _51919_ ^ _52502_ /*9498*/;
assign _52507_ = _52498_ & _52506_ /*9496*/;
assign _52367_ = _52498_ ^ _52506_ /*9497*/;
assign _52504_ = _52505_ | _52507_ /*9494*/;
assign _52509_ = ~Q[5] /*9493*/;
assign _52508_ = _52509_ & D[15] /*9492*/;
assign _52511_ = _51920_ & _52508_ /*9487*/;
assign _52512_ = _51920_ ^ _52508_ /*9490*/;
assign _52513_ = _52504_ & _52512_ /*9488*/;
assign _52368_ = _52504_ ^ _52512_ /*9489*/;
assign _52510_ = _52511_ | _52513_ /*9486*/;
assign _52515_ = ~Q[5] /*9485*/;
assign _52514_ = _52515_ & D[16] /*9484*/;
assign _52517_ = _51921_ & _52514_ /*9479*/;
assign _52518_ = _51921_ ^ _52514_ /*9482*/;
assign _52519_ = _52510_ & _52518_ /*9480*/;
assign _52369_ = _52510_ ^ _52518_ /*9481*/;
assign _52516_ = _52517_ | _52519_ /*9478*/;
assign _52521_ = ~Q[5] /*9477*/;
assign _52520_ = _52521_ & D[17] /*9476*/;
assign _52523_ = _51922_ & _52520_ /*9471*/;
assign _52524_ = _51922_ ^ _52520_ /*9474*/;
assign _52525_ = _52516_ & _52524_ /*9472*/;
assign _52370_ = _52516_ ^ _52524_ /*9473*/;
assign _52522_ = _52523_ | _52525_ /*9470*/;
assign _52527_ = ~Q[5] /*9469*/;
assign _52526_ = _52527_ & D[18] /*9468*/;
assign _52529_ = _51923_ & _52526_ /*9463*/;
assign _52530_ = _51923_ ^ _52526_ /*9466*/;
assign _52531_ = _52522_ & _52530_ /*9464*/;
assign _52371_ = _52522_ ^ _52530_ /*9465*/;
assign _52528_ = _52529_ | _52531_ /*9462*/;
assign _52533_ = ~Q[5] /*9461*/;
assign _52532_ = _52533_ & D[19] /*9460*/;
assign _52535_ = _51924_ & _52532_ /*9455*/;
assign _52536_ = _51924_ ^ _52532_ /*9458*/;
assign _52537_ = _52528_ & _52536_ /*9456*/;
assign _52372_ = _52528_ ^ _52536_ /*9457*/;
assign _52534_ = _52535_ | _52537_ /*9454*/;
assign _52539_ = ~Q[5] /*9453*/;
assign _52538_ = _52539_ & D[20] /*9452*/;
assign _52541_ = _51925_ & _52538_ /*9447*/;
assign _52542_ = _51925_ ^ _52538_ /*9450*/;
assign _52543_ = _52534_ & _52542_ /*9448*/;
assign _52373_ = _52534_ ^ _52542_ /*9449*/;
assign _52540_ = _52541_ | _52543_ /*9446*/;
assign _52545_ = ~Q[5] /*9445*/;
assign _52544_ = _52545_ & D[21] /*9444*/;
assign _52547_ = _51926_ & _52544_ /*9439*/;
assign _52548_ = _51926_ ^ _52544_ /*9442*/;
assign _52549_ = _52540_ & _52548_ /*9440*/;
assign _52374_ = _52540_ ^ _52548_ /*9441*/;
assign _52546_ = _52547_ | _52549_ /*9438*/;
assign _52551_ = ~Q[5] /*9437*/;
assign _52550_ = _52551_ & D[22] /*9436*/;
assign _52553_ = _51927_ & _52550_ /*9431*/;
assign _52554_ = _51927_ ^ _52550_ /*9434*/;
assign _52555_ = _52546_ & _52554_ /*9432*/;
assign _52375_ = _52546_ ^ _52554_ /*9433*/;
assign _52552_ = _52553_ | _52555_ /*9430*/;
assign _52557_ = ~Q[5] /*9429*/;
assign _52556_ = _52557_ & D[23] /*9428*/;
assign _52559_ = _51928_ & _52556_ /*9423*/;
assign _52560_ = _51928_ ^ _52556_ /*9426*/;
assign _52561_ = _52552_ & _52560_ /*9424*/;
assign _52376_ = _52552_ ^ _52560_ /*9425*/;
assign _52558_ = _52559_ | _52561_ /*9422*/;
assign _52563_ = ~Q[5] /*9421*/;
assign _52562_ = _52563_ & D[24] /*9420*/;
assign _52565_ = _51929_ & _52562_ /*9415*/;
assign _52566_ = _51929_ ^ _52562_ /*9418*/;
assign _52567_ = _52558_ & _52566_ /*9416*/;
assign _52377_ = _52558_ ^ _52566_ /*9417*/;
assign _52564_ = _52565_ | _52567_ /*9414*/;
assign _52569_ = ~Q[5] /*9413*/;
assign _52568_ = _52569_ & D[25] /*9412*/;
assign _52571_ = _51930_ & _52568_ /*9407*/;
assign _52572_ = _51930_ ^ _52568_ /*9410*/;
assign _52573_ = _52564_ & _52572_ /*9408*/;
assign _52378_ = _52564_ ^ _52572_ /*9409*/;
assign _52570_ = _52571_ | _52573_ /*9406*/;
assign _52575_ = ~Q[5] /*9405*/;
assign _52574_ = _52575_ & D[26] /*9404*/;
assign _52577_ = _51931_ & _52574_ /*9399*/;
assign _52578_ = _51931_ ^ _52574_ /*9402*/;
assign _52579_ = _52570_ & _52578_ /*9400*/;
assign _52379_ = _52570_ ^ _52578_ /*9401*/;
assign _52576_ = _52577_ | _52579_ /*9398*/;
assign _52581_ = ~Q[5] /*9397*/;
assign _52580_ = _52581_ & D[27] /*9396*/;
assign _52583_ = _51932_ & _52580_ /*9391*/;
assign _52584_ = _51932_ ^ _52580_ /*9394*/;
assign _52585_ = _52576_ & _52584_ /*9392*/;
assign _52380_ = _52576_ ^ _52584_ /*9393*/;
assign _52582_ = _52583_ | _52585_ /*9390*/;
assign _52587_ = ~Q[5] /*9389*/;
assign _52586_ = _52587_ & D[28] /*9388*/;
assign _52589_ = _51933_ & _52586_ /*9383*/;
assign _52590_ = _51933_ ^ _52586_ /*9386*/;
assign _52591_ = _52582_ & _52590_ /*9384*/;
assign _52381_ = _52582_ ^ _52590_ /*9385*/;
assign _52588_ = _52589_ | _52591_ /*9382*/;
assign _52593_ = ~Q[5] /*9381*/;
assign _52592_ = _52593_ & D[29] /*9380*/;
assign _52595_ = _51934_ & _52592_ /*9375*/;
assign _52596_ = _51934_ ^ _52592_ /*9378*/;
assign _52597_ = _52588_ & _52596_ /*9376*/;
assign _52382_ = _52588_ ^ _52596_ /*9377*/;
assign _52594_ = _52595_ | _52597_ /*9374*/;
assign _52599_ = ~Q[5] /*9373*/;
assign _52598_ = _52599_ & D[30] /*9372*/;
assign _52601_ = _51935_ & _52598_ /*9367*/;
assign _52602_ = _51935_ ^ _52598_ /*9370*/;
assign _52603_ = _52594_ & _52602_ /*9368*/;
assign _52383_ = _52594_ ^ _52602_ /*9369*/;
assign _52600_ = _52601_ | _52603_ /*9366*/;
assign _52605_ = ~Q[5] /*9365*/;
assign _52604_ = _52605_ & D[31] /*9364*/;
assign _52607_ = _51936_ & _52604_ /*9359*/;
assign _52608_ = _51936_ ^ _52604_ /*9362*/;
assign _52609_ = _52600_ & _52608_ /*9360*/;
assign _52384_ = _52600_ ^ _52608_ /*9361*/;
assign _52606_ = _52607_ | _52609_ /*9358*/;
assign _52611_ = ~Q[5] /*9357*/;
assign _52610_ = _52611_ & D[32] /*9356*/;
assign _52613_ = _51937_ & _52610_ /*9351*/;
assign _52614_ = _51937_ ^ _52610_ /*9354*/;
assign _52615_ = _52606_ & _52614_ /*9352*/;
assign _52385_ = _52606_ ^ _52614_ /*9353*/;
assign _52612_ = _52613_ | _52615_ /*9350*/;
assign _52617_ = ~Q[5] /*9349*/;
assign _52616_ = _52617_ & D[33] /*9348*/;
assign _52619_ = _51938_ & _52616_ /*9343*/;
assign _52620_ = _51938_ ^ _52616_ /*9346*/;
assign _52621_ = _52612_ & _52620_ /*9344*/;
assign _52386_ = _52612_ ^ _52620_ /*9345*/;
assign _52618_ = _52619_ | _52621_ /*9342*/;
assign _52623_ = ~Q[5] /*9341*/;
assign _52622_ = _52623_ & D[34] /*9340*/;
assign _52625_ = _51939_ & _52622_ /*9335*/;
assign _52626_ = _51939_ ^ _52622_ /*9338*/;
assign _52627_ = _52618_ & _52626_ /*9336*/;
assign _52387_ = _52618_ ^ _52626_ /*9337*/;
assign _52624_ = _52625_ | _52627_ /*9334*/;
assign _52629_ = ~Q[5] /*9333*/;
assign _52628_ = _52629_ & D[35] /*9332*/;
assign _52631_ = _51940_ & _52628_ /*9327*/;
assign _52632_ = _51940_ ^ _52628_ /*9330*/;
assign _52633_ = _52624_ & _52632_ /*9328*/;
assign _52388_ = _52624_ ^ _52632_ /*9329*/;
assign _52630_ = _52631_ | _52633_ /*9326*/;
assign _52635_ = ~Q[5] /*9325*/;
assign _52634_ = _52635_ & D[36] /*9324*/;
assign _52637_ = _51941_ & _52634_ /*9319*/;
assign _52638_ = _51941_ ^ _52634_ /*9322*/;
assign _52639_ = _52630_ & _52638_ /*9320*/;
assign _52389_ = _52630_ ^ _52638_ /*9321*/;
assign _52636_ = _52637_ | _52639_ /*9318*/;
assign _52641_ = ~Q[5] /*9317*/;
assign _52640_ = _52641_ & D[37] /*9316*/;
assign _52643_ = _51942_ & _52640_ /*9311*/;
assign _52644_ = _51942_ ^ _52640_ /*9314*/;
assign _52645_ = _52636_ & _52644_ /*9312*/;
assign _52390_ = _52636_ ^ _52644_ /*9313*/;
assign _52642_ = _52643_ | _52645_ /*9310*/;
assign _52647_ = ~Q[5] /*9309*/;
assign _52646_ = _52647_ & D[38] /*9308*/;
assign _52649_ = _51943_ & _52646_ /*9303*/;
assign _52650_ = _51943_ ^ _52646_ /*9306*/;
assign _52651_ = _52642_ & _52650_ /*9304*/;
assign _52391_ = _52642_ ^ _52650_ /*9305*/;
assign _52648_ = _52649_ | _52651_ /*9302*/;
assign _52653_ = ~Q[5] /*9301*/;
assign _52652_ = _52653_ & D[39] /*9300*/;
assign _52655_ = _51944_ & _52652_ /*9295*/;
assign _52656_ = _51944_ ^ _52652_ /*9298*/;
assign _52657_ = _52648_ & _52656_ /*9296*/;
assign _52392_ = _52648_ ^ _52656_ /*9297*/;
assign _52654_ = _52655_ | _52657_ /*9294*/;
assign _52659_ = ~Q[5] /*9293*/;
assign _52658_ = _52659_ & D[40] /*9292*/;
assign _52661_ = _51945_ & _52658_ /*9287*/;
assign _52662_ = _51945_ ^ _52658_ /*9290*/;
assign _52663_ = _52654_ & _52662_ /*9288*/;
assign _52393_ = _52654_ ^ _52662_ /*9289*/;
assign _52660_ = _52661_ | _52663_ /*9286*/;
assign _52665_ = ~Q[5] /*9285*/;
assign _52664_ = _52665_ & D[41] /*9284*/;
assign _52667_ = _51946_ & _52664_ /*9279*/;
assign _52668_ = _51946_ ^ _52664_ /*9282*/;
assign _52669_ = _52660_ & _52668_ /*9280*/;
assign _52394_ = _52660_ ^ _52668_ /*9281*/;
assign _52666_ = _52667_ | _52669_ /*9278*/;
assign _52671_ = ~Q[5] /*9277*/;
assign _52670_ = _52671_ & D[42] /*9276*/;
assign _52673_ = _51947_ & _52670_ /*9271*/;
assign _52674_ = _51947_ ^ _52670_ /*9274*/;
assign _52675_ = _52666_ & _52674_ /*9272*/;
assign _52395_ = _52666_ ^ _52674_ /*9273*/;
assign _52672_ = _52673_ | _52675_ /*9270*/;
assign _52677_ = ~Q[5] /*9269*/;
assign _52676_ = _52677_ & D[43] /*9268*/;
assign _52679_ = _51948_ & _52676_ /*9263*/;
assign _52680_ = _51948_ ^ _52676_ /*9266*/;
assign _52681_ = _52672_ & _52680_ /*9264*/;
assign _52396_ = _52672_ ^ _52680_ /*9265*/;
assign _52678_ = _52679_ | _52681_ /*9262*/;
assign _52683_ = ~Q[5] /*9261*/;
assign _52682_ = _52683_ & D[44] /*9260*/;
assign _52685_ = _51949_ & _52682_ /*9255*/;
assign _52686_ = _51949_ ^ _52682_ /*9258*/;
assign _52687_ = _52678_ & _52686_ /*9256*/;
assign _52397_ = _52678_ ^ _52686_ /*9257*/;
assign _52684_ = _52685_ | _52687_ /*9254*/;
assign _52689_ = ~Q[5] /*9253*/;
assign _52688_ = _52689_ & D[45] /*9252*/;
assign _52691_ = _51950_ & _52688_ /*9247*/;
assign _52692_ = _51950_ ^ _52688_ /*9250*/;
assign _52693_ = _52684_ & _52692_ /*9248*/;
assign _52398_ = _52684_ ^ _52692_ /*9249*/;
assign _52690_ = _52691_ | _52693_ /*9246*/;
assign _52695_ = ~Q[5] /*9245*/;
assign _52694_ = _52695_ & D[46] /*9244*/;
assign _52697_ = _51951_ & _52694_ /*9239*/;
assign _52698_ = _51951_ ^ _52694_ /*9242*/;
assign _52699_ = _52690_ & _52698_ /*9240*/;
assign _52399_ = _52690_ ^ _52698_ /*9241*/;
assign _52696_ = _52697_ | _52699_ /*9238*/;
assign _52701_ = ~Q[5] /*9237*/;
assign _52700_ = _52701_ & D[47] /*9236*/;
assign _52703_ = _51952_ & _52700_ /*9231*/;
assign _52704_ = _51952_ ^ _52700_ /*9234*/;
assign _52705_ = _52696_ & _52704_ /*9232*/;
assign _52400_ = _52696_ ^ _52704_ /*9233*/;
assign _52702_ = _52703_ | _52705_ /*9230*/;
assign _52707_ = ~Q[5] /*9229*/;
assign _52706_ = _52707_ & D[48] /*9228*/;
assign _52709_ = _51953_ & _52706_ /*9223*/;
assign _52710_ = _51953_ ^ _52706_ /*9226*/;
assign _52711_ = _52702_ & _52710_ /*9224*/;
assign _52401_ = _52702_ ^ _52710_ /*9225*/;
assign _52708_ = _52709_ | _52711_ /*9222*/;
assign _52713_ = ~Q[5] /*9221*/;
assign _52712_ = _52713_ & D[49] /*9220*/;
assign _52715_ = _51954_ & _52712_ /*9215*/;
assign _52716_ = _51954_ ^ _52712_ /*9218*/;
assign _52717_ = _52708_ & _52716_ /*9216*/;
assign _52402_ = _52708_ ^ _52716_ /*9217*/;
assign _52714_ = _52715_ | _52717_ /*9214*/;
assign _52719_ = ~Q[5] /*9213*/;
assign _52718_ = _52719_ & D[50] /*9212*/;
assign _52721_ = _51955_ & _52718_ /*9207*/;
assign _52722_ = _51955_ ^ _52718_ /*9210*/;
assign _52723_ = _52714_ & _52722_ /*9208*/;
assign _52403_ = _52714_ ^ _52722_ /*9209*/;
assign _52720_ = _52721_ | _52723_ /*9206*/;
assign _52725_ = ~Q[5] /*9205*/;
assign _52724_ = _52725_ & D[51] /*9204*/;
assign _52727_ = _51956_ & _52724_ /*9199*/;
assign _52728_ = _51956_ ^ _52724_ /*9202*/;
assign _52729_ = _52720_ & _52728_ /*9200*/;
assign _52404_ = _52720_ ^ _52728_ /*9201*/;
assign _52726_ = _52727_ | _52729_ /*9198*/;
assign _52731_ = ~Q[5] /*9197*/;
assign _52730_ = _52731_ & D[52] /*9196*/;
assign _52733_ = _51957_ & _52730_ /*9191*/;
assign _52734_ = _51957_ ^ _52730_ /*9194*/;
assign _52735_ = _52726_ & _52734_ /*9192*/;
assign _52405_ = _52726_ ^ _52734_ /*9193*/;
assign _52732_ = _52733_ | _52735_ /*9190*/;
assign _52737_ = ~Q[5] /*9189*/;
assign _52736_ = _52737_ & D[53] /*9188*/;
assign _52739_ = _51958_ & _52736_ /*9183*/;
assign _52740_ = _51958_ ^ _52736_ /*9186*/;
assign _52741_ = _52732_ & _52740_ /*9184*/;
assign _52406_ = _52732_ ^ _52740_ /*9185*/;
assign _52738_ = _52739_ | _52741_ /*9182*/;
assign _52743_ = ~Q[5] /*9181*/;
assign _52742_ = _52743_ & D[54] /*9180*/;
assign _52745_ = _51959_ & _52742_ /*9175*/;
assign _52746_ = _51959_ ^ _52742_ /*9178*/;
assign _52747_ = _52738_ & _52746_ /*9176*/;
assign _52407_ = _52738_ ^ _52746_ /*9177*/;
assign _52744_ = _52745_ | _52747_ /*9174*/;
assign _52749_ = ~Q[5] /*9173*/;
assign _52748_ = _52749_ & D[55] /*9172*/;
assign _52751_ = _51960_ & _52748_ /*9167*/;
assign _52752_ = _51960_ ^ _52748_ /*9170*/;
assign _52753_ = _52744_ & _52752_ /*9168*/;
assign _52408_ = _52744_ ^ _52752_ /*9169*/;
assign _52750_ = _52751_ | _52753_ /*9166*/;
assign _52755_ = ~Q[5] /*9165*/;
assign _52754_ = _52755_ & D[56] /*9164*/;
assign _52757_ = _51961_ & _52754_ /*9159*/;
assign _52758_ = _51961_ ^ _52754_ /*9162*/;
assign _52759_ = _52750_ & _52758_ /*9160*/;
assign _52409_ = _52750_ ^ _52758_ /*9161*/;
assign _52756_ = _52757_ | _52759_ /*9158*/;
assign _52761_ = ~Q[5] /*9157*/;
assign _52760_ = _52761_ & D[57] /*9156*/;
assign _52763_ = _51962_ & _52760_ /*9151*/;
assign _52764_ = _51962_ ^ _52760_ /*9154*/;
assign _52765_ = _52756_ & _52764_ /*9152*/;
assign _52410_ = _52756_ ^ _52764_ /*9153*/;
assign _52762_ = _52763_ | _52765_ /*9150*/;
assign _52767_ = ~Q[5] /*9149*/;
assign _52766_ = _52767_ & D[58] /*9148*/;
assign _52769_ = _51963_ & _52766_ /*9143*/;
assign _52770_ = _51963_ ^ _52766_ /*9146*/;
assign _52771_ = _52762_ & _52770_ /*9144*/;
assign _52411_ = _52762_ ^ _52770_ /*9145*/;
assign _52768_ = _52769_ | _52771_ /*9142*/;
assign _52773_ = ~Q[5] /*9141*/;
assign _52772_ = _52773_ & D[59] /*9140*/;
assign _52775_ = _51964_ & _52772_ /*9135*/;
assign _52776_ = _51964_ ^ _52772_ /*9138*/;
assign _52777_ = _52768_ & _52776_ /*9136*/;
assign _52412_ = _52768_ ^ _52776_ /*9137*/;
assign _52774_ = _52775_ | _52777_ /*9134*/;
assign _52779_ = ~Q[5] /*9133*/;
assign _52778_ = _52779_ & D[60] /*9132*/;
assign _52781_ = _51965_ & _52778_ /*9127*/;
assign _52782_ = _51965_ ^ _52778_ /*9130*/;
assign _52783_ = _52774_ & _52782_ /*9128*/;
assign _52413_ = _52774_ ^ _52782_ /*9129*/;
assign _52780_ = _52781_ | _52783_ /*9126*/;
assign _52785_ = ~Q[5] /*9125*/;
assign _52784_ = _52785_ & D[61] /*9124*/;
assign _52787_ = _51966_ & _52784_ /*9119*/;
assign _52788_ = _51966_ ^ _52784_ /*9122*/;
assign _52789_ = _52780_ & _52788_ /*9120*/;
assign _52414_ = _52780_ ^ _52788_ /*9121*/;
assign _52786_ = _52787_ | _52789_ /*9118*/;
assign _52791_ = ~Q[5] /*9117*/;
assign _52790_ = _52791_ & D[62] /*9116*/;
assign _52793_ = _51967_ & _52790_ /*9111*/;
assign _52794_ = _51967_ ^ _52790_ /*9114*/;
assign _52795_ = _52786_ & _52794_ /*9112*/;
assign _52415_ = _52786_ ^ _52794_ /*9113*/;
assign _52792_ = _52793_ | _52795_ /*9110*/;
assign _52797_ = ~Q[5] /*9109*/;
assign _52796_ = _52797_ & zeroWire /*9108*/;
assign _52798_ = _51968_ ^ _52796_ /*9106*/;
assign _52416_ = _52798_ ^ _52792_ /*9105*/;
assign _52869_ = ~D[0] /*8851*/;
assign _52866_ = R_0[4] & _52869_ /*8847*/;
assign _52867_ = R_0[4] ^ _52869_ /*8850*/;
assign _52868_ = oneWire & _52867_ /*8848*/;
assign _52801_ = oneWire ^ _52867_ /*8849*/;
assign _52865_ = _52866_ | _52868_ /*8846*/;
assign _52874_ = ~D[1] /*8845*/;
assign _52871_ = _52353_ & _52874_ /*8841*/;
assign _52872_ = _52353_ ^ _52874_ /*8844*/;
assign _52873_ = _52865_ & _52872_ /*8842*/;
assign _52802_ = _52865_ ^ _52872_ /*8843*/;
assign _52870_ = _52871_ | _52873_ /*8840*/;
assign _52879_ = ~D[2] /*8839*/;
assign _52876_ = _52354_ & _52879_ /*8835*/;
assign _52877_ = _52354_ ^ _52879_ /*8838*/;
assign _52878_ = _52870_ & _52877_ /*8836*/;
assign _52803_ = _52870_ ^ _52877_ /*8837*/;
assign _52875_ = _52876_ | _52878_ /*8834*/;
assign _52884_ = ~D[3] /*8833*/;
assign _52881_ = _52355_ & _52884_ /*8829*/;
assign _52882_ = _52355_ ^ _52884_ /*8832*/;
assign _52883_ = _52875_ & _52882_ /*8830*/;
assign _52804_ = _52875_ ^ _52882_ /*8831*/;
assign _52880_ = _52881_ | _52883_ /*8828*/;
assign _52889_ = ~D[4] /*8827*/;
assign _52886_ = _52356_ & _52889_ /*8823*/;
assign _52887_ = _52356_ ^ _52889_ /*8826*/;
assign _52888_ = _52880_ & _52887_ /*8824*/;
assign _52805_ = _52880_ ^ _52887_ /*8825*/;
assign _52885_ = _52886_ | _52888_ /*8822*/;
assign _52894_ = ~D[5] /*8821*/;
assign _52891_ = _52357_ & _52894_ /*8817*/;
assign _52892_ = _52357_ ^ _52894_ /*8820*/;
assign _52893_ = _52885_ & _52892_ /*8818*/;
assign _52806_ = _52885_ ^ _52892_ /*8819*/;
assign _52890_ = _52891_ | _52893_ /*8816*/;
assign _52899_ = ~D[6] /*8815*/;
assign _52896_ = _52358_ & _52899_ /*8811*/;
assign _52897_ = _52358_ ^ _52899_ /*8814*/;
assign _52898_ = _52890_ & _52897_ /*8812*/;
assign _52807_ = _52890_ ^ _52897_ /*8813*/;
assign _52895_ = _52896_ | _52898_ /*8810*/;
assign _52904_ = ~D[7] /*8809*/;
assign _52901_ = _52359_ & _52904_ /*8805*/;
assign _52902_ = _52359_ ^ _52904_ /*8808*/;
assign _52903_ = _52895_ & _52902_ /*8806*/;
assign _52808_ = _52895_ ^ _52902_ /*8807*/;
assign _52900_ = _52901_ | _52903_ /*8804*/;
assign _52909_ = ~D[8] /*8803*/;
assign _52906_ = _52360_ & _52909_ /*8799*/;
assign _52907_ = _52360_ ^ _52909_ /*8802*/;
assign _52908_ = _52900_ & _52907_ /*8800*/;
assign _52809_ = _52900_ ^ _52907_ /*8801*/;
assign _52905_ = _52906_ | _52908_ /*8798*/;
assign _52914_ = ~D[9] /*8797*/;
assign _52911_ = _52361_ & _52914_ /*8793*/;
assign _52912_ = _52361_ ^ _52914_ /*8796*/;
assign _52913_ = _52905_ & _52912_ /*8794*/;
assign _52810_ = _52905_ ^ _52912_ /*8795*/;
assign _52910_ = _52911_ | _52913_ /*8792*/;
assign _52919_ = ~D[10] /*8791*/;
assign _52916_ = _52362_ & _52919_ /*8787*/;
assign _52917_ = _52362_ ^ _52919_ /*8790*/;
assign _52918_ = _52910_ & _52917_ /*8788*/;
assign _52811_ = _52910_ ^ _52917_ /*8789*/;
assign _52915_ = _52916_ | _52918_ /*8786*/;
assign _52924_ = ~D[11] /*8785*/;
assign _52921_ = _52363_ & _52924_ /*8781*/;
assign _52922_ = _52363_ ^ _52924_ /*8784*/;
assign _52923_ = _52915_ & _52922_ /*8782*/;
assign _52812_ = _52915_ ^ _52922_ /*8783*/;
assign _52920_ = _52921_ | _52923_ /*8780*/;
assign _52929_ = ~D[12] /*8779*/;
assign _52926_ = _52364_ & _52929_ /*8775*/;
assign _52927_ = _52364_ ^ _52929_ /*8778*/;
assign _52928_ = _52920_ & _52927_ /*8776*/;
assign _52813_ = _52920_ ^ _52927_ /*8777*/;
assign _52925_ = _52926_ | _52928_ /*8774*/;
assign _52934_ = ~D[13] /*8773*/;
assign _52931_ = _52365_ & _52934_ /*8769*/;
assign _52932_ = _52365_ ^ _52934_ /*8772*/;
assign _52933_ = _52925_ & _52932_ /*8770*/;
assign _52814_ = _52925_ ^ _52932_ /*8771*/;
assign _52930_ = _52931_ | _52933_ /*8768*/;
assign _52939_ = ~D[14] /*8767*/;
assign _52936_ = _52366_ & _52939_ /*8763*/;
assign _52937_ = _52366_ ^ _52939_ /*8766*/;
assign _52938_ = _52930_ & _52937_ /*8764*/;
assign _52815_ = _52930_ ^ _52937_ /*8765*/;
assign _52935_ = _52936_ | _52938_ /*8762*/;
assign _52944_ = ~D[15] /*8761*/;
assign _52941_ = _52367_ & _52944_ /*8757*/;
assign _52942_ = _52367_ ^ _52944_ /*8760*/;
assign _52943_ = _52935_ & _52942_ /*8758*/;
assign _52816_ = _52935_ ^ _52942_ /*8759*/;
assign _52940_ = _52941_ | _52943_ /*8756*/;
assign _52949_ = ~D[16] /*8755*/;
assign _52946_ = _52368_ & _52949_ /*8751*/;
assign _52947_ = _52368_ ^ _52949_ /*8754*/;
assign _52948_ = _52940_ & _52947_ /*8752*/;
assign _52817_ = _52940_ ^ _52947_ /*8753*/;
assign _52945_ = _52946_ | _52948_ /*8750*/;
assign _52954_ = ~D[17] /*8749*/;
assign _52951_ = _52369_ & _52954_ /*8745*/;
assign _52952_ = _52369_ ^ _52954_ /*8748*/;
assign _52953_ = _52945_ & _52952_ /*8746*/;
assign _52818_ = _52945_ ^ _52952_ /*8747*/;
assign _52950_ = _52951_ | _52953_ /*8744*/;
assign _52959_ = ~D[18] /*8743*/;
assign _52956_ = _52370_ & _52959_ /*8739*/;
assign _52957_ = _52370_ ^ _52959_ /*8742*/;
assign _52958_ = _52950_ & _52957_ /*8740*/;
assign _52819_ = _52950_ ^ _52957_ /*8741*/;
assign _52955_ = _52956_ | _52958_ /*8738*/;
assign _52964_ = ~D[19] /*8737*/;
assign _52961_ = _52371_ & _52964_ /*8733*/;
assign _52962_ = _52371_ ^ _52964_ /*8736*/;
assign _52963_ = _52955_ & _52962_ /*8734*/;
assign _52820_ = _52955_ ^ _52962_ /*8735*/;
assign _52960_ = _52961_ | _52963_ /*8732*/;
assign _52969_ = ~D[20] /*8731*/;
assign _52966_ = _52372_ & _52969_ /*8727*/;
assign _52967_ = _52372_ ^ _52969_ /*8730*/;
assign _52968_ = _52960_ & _52967_ /*8728*/;
assign _52821_ = _52960_ ^ _52967_ /*8729*/;
assign _52965_ = _52966_ | _52968_ /*8726*/;
assign _52974_ = ~D[21] /*8725*/;
assign _52971_ = _52373_ & _52974_ /*8721*/;
assign _52972_ = _52373_ ^ _52974_ /*8724*/;
assign _52973_ = _52965_ & _52972_ /*8722*/;
assign _52822_ = _52965_ ^ _52972_ /*8723*/;
assign _52970_ = _52971_ | _52973_ /*8720*/;
assign _52979_ = ~D[22] /*8719*/;
assign _52976_ = _52374_ & _52979_ /*8715*/;
assign _52977_ = _52374_ ^ _52979_ /*8718*/;
assign _52978_ = _52970_ & _52977_ /*8716*/;
assign _52823_ = _52970_ ^ _52977_ /*8717*/;
assign _52975_ = _52976_ | _52978_ /*8714*/;
assign _52984_ = ~D[23] /*8713*/;
assign _52981_ = _52375_ & _52984_ /*8709*/;
assign _52982_ = _52375_ ^ _52984_ /*8712*/;
assign _52983_ = _52975_ & _52982_ /*8710*/;
assign _52824_ = _52975_ ^ _52982_ /*8711*/;
assign _52980_ = _52981_ | _52983_ /*8708*/;
assign _52989_ = ~D[24] /*8707*/;
assign _52986_ = _52376_ & _52989_ /*8703*/;
assign _52987_ = _52376_ ^ _52989_ /*8706*/;
assign _52988_ = _52980_ & _52987_ /*8704*/;
assign _52825_ = _52980_ ^ _52987_ /*8705*/;
assign _52985_ = _52986_ | _52988_ /*8702*/;
assign _52994_ = ~D[25] /*8701*/;
assign _52991_ = _52377_ & _52994_ /*8697*/;
assign _52992_ = _52377_ ^ _52994_ /*8700*/;
assign _52993_ = _52985_ & _52992_ /*8698*/;
assign _52826_ = _52985_ ^ _52992_ /*8699*/;
assign _52990_ = _52991_ | _52993_ /*8696*/;
assign _52999_ = ~D[26] /*8695*/;
assign _52996_ = _52378_ & _52999_ /*8691*/;
assign _52997_ = _52378_ ^ _52999_ /*8694*/;
assign _52998_ = _52990_ & _52997_ /*8692*/;
assign _52827_ = _52990_ ^ _52997_ /*8693*/;
assign _52995_ = _52996_ | _52998_ /*8690*/;
assign _53004_ = ~D[27] /*8689*/;
assign _53001_ = _52379_ & _53004_ /*8685*/;
assign _53002_ = _52379_ ^ _53004_ /*8688*/;
assign _53003_ = _52995_ & _53002_ /*8686*/;
assign _52828_ = _52995_ ^ _53002_ /*8687*/;
assign _53000_ = _53001_ | _53003_ /*8684*/;
assign _53009_ = ~D[28] /*8683*/;
assign _53006_ = _52380_ & _53009_ /*8679*/;
assign _53007_ = _52380_ ^ _53009_ /*8682*/;
assign _53008_ = _53000_ & _53007_ /*8680*/;
assign _52829_ = _53000_ ^ _53007_ /*8681*/;
assign _53005_ = _53006_ | _53008_ /*8678*/;
assign _53014_ = ~D[29] /*8677*/;
assign _53011_ = _52381_ & _53014_ /*8673*/;
assign _53012_ = _52381_ ^ _53014_ /*8676*/;
assign _53013_ = _53005_ & _53012_ /*8674*/;
assign _52830_ = _53005_ ^ _53012_ /*8675*/;
assign _53010_ = _53011_ | _53013_ /*8672*/;
assign _53019_ = ~D[30] /*8671*/;
assign _53016_ = _52382_ & _53019_ /*8667*/;
assign _53017_ = _52382_ ^ _53019_ /*8670*/;
assign _53018_ = _53010_ & _53017_ /*8668*/;
assign _52831_ = _53010_ ^ _53017_ /*8669*/;
assign _53015_ = _53016_ | _53018_ /*8666*/;
assign _53024_ = ~D[31] /*8665*/;
assign _53021_ = _52383_ & _53024_ /*8661*/;
assign _53022_ = _52383_ ^ _53024_ /*8664*/;
assign _53023_ = _53015_ & _53022_ /*8662*/;
assign _52832_ = _53015_ ^ _53022_ /*8663*/;
assign _53020_ = _53021_ | _53023_ /*8660*/;
assign _53029_ = ~D[32] /*8659*/;
assign _53026_ = _52384_ & _53029_ /*8655*/;
assign _53027_ = _52384_ ^ _53029_ /*8658*/;
assign _53028_ = _53020_ & _53027_ /*8656*/;
assign _52833_ = _53020_ ^ _53027_ /*8657*/;
assign _53025_ = _53026_ | _53028_ /*8654*/;
assign _53034_ = ~D[33] /*8653*/;
assign _53031_ = _52385_ & _53034_ /*8649*/;
assign _53032_ = _52385_ ^ _53034_ /*8652*/;
assign _53033_ = _53025_ & _53032_ /*8650*/;
assign _52834_ = _53025_ ^ _53032_ /*8651*/;
assign _53030_ = _53031_ | _53033_ /*8648*/;
assign _53039_ = ~D[34] /*8647*/;
assign _53036_ = _52386_ & _53039_ /*8643*/;
assign _53037_ = _52386_ ^ _53039_ /*8646*/;
assign _53038_ = _53030_ & _53037_ /*8644*/;
assign _52835_ = _53030_ ^ _53037_ /*8645*/;
assign _53035_ = _53036_ | _53038_ /*8642*/;
assign _53044_ = ~D[35] /*8641*/;
assign _53041_ = _52387_ & _53044_ /*8637*/;
assign _53042_ = _52387_ ^ _53044_ /*8640*/;
assign _53043_ = _53035_ & _53042_ /*8638*/;
assign _52836_ = _53035_ ^ _53042_ /*8639*/;
assign _53040_ = _53041_ | _53043_ /*8636*/;
assign _53049_ = ~D[36] /*8635*/;
assign _53046_ = _52388_ & _53049_ /*8631*/;
assign _53047_ = _52388_ ^ _53049_ /*8634*/;
assign _53048_ = _53040_ & _53047_ /*8632*/;
assign _52837_ = _53040_ ^ _53047_ /*8633*/;
assign _53045_ = _53046_ | _53048_ /*8630*/;
assign _53054_ = ~D[37] /*8629*/;
assign _53051_ = _52389_ & _53054_ /*8625*/;
assign _53052_ = _52389_ ^ _53054_ /*8628*/;
assign _53053_ = _53045_ & _53052_ /*8626*/;
assign _52838_ = _53045_ ^ _53052_ /*8627*/;
assign _53050_ = _53051_ | _53053_ /*8624*/;
assign _53059_ = ~D[38] /*8623*/;
assign _53056_ = _52390_ & _53059_ /*8619*/;
assign _53057_ = _52390_ ^ _53059_ /*8622*/;
assign _53058_ = _53050_ & _53057_ /*8620*/;
assign _52839_ = _53050_ ^ _53057_ /*8621*/;
assign _53055_ = _53056_ | _53058_ /*8618*/;
assign _53064_ = ~D[39] /*8617*/;
assign _53061_ = _52391_ & _53064_ /*8613*/;
assign _53062_ = _52391_ ^ _53064_ /*8616*/;
assign _53063_ = _53055_ & _53062_ /*8614*/;
assign _52840_ = _53055_ ^ _53062_ /*8615*/;
assign _53060_ = _53061_ | _53063_ /*8612*/;
assign _53069_ = ~D[40] /*8611*/;
assign _53066_ = _52392_ & _53069_ /*8607*/;
assign _53067_ = _52392_ ^ _53069_ /*8610*/;
assign _53068_ = _53060_ & _53067_ /*8608*/;
assign _52841_ = _53060_ ^ _53067_ /*8609*/;
assign _53065_ = _53066_ | _53068_ /*8606*/;
assign _53074_ = ~D[41] /*8605*/;
assign _53071_ = _52393_ & _53074_ /*8601*/;
assign _53072_ = _52393_ ^ _53074_ /*8604*/;
assign _53073_ = _53065_ & _53072_ /*8602*/;
assign _52842_ = _53065_ ^ _53072_ /*8603*/;
assign _53070_ = _53071_ | _53073_ /*8600*/;
assign _53079_ = ~D[42] /*8599*/;
assign _53076_ = _52394_ & _53079_ /*8595*/;
assign _53077_ = _52394_ ^ _53079_ /*8598*/;
assign _53078_ = _53070_ & _53077_ /*8596*/;
assign _52843_ = _53070_ ^ _53077_ /*8597*/;
assign _53075_ = _53076_ | _53078_ /*8594*/;
assign _53084_ = ~D[43] /*8593*/;
assign _53081_ = _52395_ & _53084_ /*8589*/;
assign _53082_ = _52395_ ^ _53084_ /*8592*/;
assign _53083_ = _53075_ & _53082_ /*8590*/;
assign _52844_ = _53075_ ^ _53082_ /*8591*/;
assign _53080_ = _53081_ | _53083_ /*8588*/;
assign _53089_ = ~D[44] /*8587*/;
assign _53086_ = _52396_ & _53089_ /*8583*/;
assign _53087_ = _52396_ ^ _53089_ /*8586*/;
assign _53088_ = _53080_ & _53087_ /*8584*/;
assign _52845_ = _53080_ ^ _53087_ /*8585*/;
assign _53085_ = _53086_ | _53088_ /*8582*/;
assign _53094_ = ~D[45] /*8581*/;
assign _53091_ = _52397_ & _53094_ /*8577*/;
assign _53092_ = _52397_ ^ _53094_ /*8580*/;
assign _53093_ = _53085_ & _53092_ /*8578*/;
assign _52846_ = _53085_ ^ _53092_ /*8579*/;
assign _53090_ = _53091_ | _53093_ /*8576*/;
assign _53099_ = ~D[46] /*8575*/;
assign _53096_ = _52398_ & _53099_ /*8571*/;
assign _53097_ = _52398_ ^ _53099_ /*8574*/;
assign _53098_ = _53090_ & _53097_ /*8572*/;
assign _52847_ = _53090_ ^ _53097_ /*8573*/;
assign _53095_ = _53096_ | _53098_ /*8570*/;
assign _53104_ = ~D[47] /*8569*/;
assign _53101_ = _52399_ & _53104_ /*8565*/;
assign _53102_ = _52399_ ^ _53104_ /*8568*/;
assign _53103_ = _53095_ & _53102_ /*8566*/;
assign _52848_ = _53095_ ^ _53102_ /*8567*/;
assign _53100_ = _53101_ | _53103_ /*8564*/;
assign _53109_ = ~D[48] /*8563*/;
assign _53106_ = _52400_ & _53109_ /*8559*/;
assign _53107_ = _52400_ ^ _53109_ /*8562*/;
assign _53108_ = _53100_ & _53107_ /*8560*/;
assign _52849_ = _53100_ ^ _53107_ /*8561*/;
assign _53105_ = _53106_ | _53108_ /*8558*/;
assign _53114_ = ~D[49] /*8557*/;
assign _53111_ = _52401_ & _53114_ /*8553*/;
assign _53112_ = _52401_ ^ _53114_ /*8556*/;
assign _53113_ = _53105_ & _53112_ /*8554*/;
assign _52850_ = _53105_ ^ _53112_ /*8555*/;
assign _53110_ = _53111_ | _53113_ /*8552*/;
assign _53119_ = ~D[50] /*8551*/;
assign _53116_ = _52402_ & _53119_ /*8547*/;
assign _53117_ = _52402_ ^ _53119_ /*8550*/;
assign _53118_ = _53110_ & _53117_ /*8548*/;
assign _52851_ = _53110_ ^ _53117_ /*8549*/;
assign _53115_ = _53116_ | _53118_ /*8546*/;
assign _53124_ = ~D[51] /*8545*/;
assign _53121_ = _52403_ & _53124_ /*8541*/;
assign _53122_ = _52403_ ^ _53124_ /*8544*/;
assign _53123_ = _53115_ & _53122_ /*8542*/;
assign _52852_ = _53115_ ^ _53122_ /*8543*/;
assign _53120_ = _53121_ | _53123_ /*8540*/;
assign _53129_ = ~D[52] /*8539*/;
assign _53126_ = _52404_ & _53129_ /*8535*/;
assign _53127_ = _52404_ ^ _53129_ /*8538*/;
assign _53128_ = _53120_ & _53127_ /*8536*/;
assign _52853_ = _53120_ ^ _53127_ /*8537*/;
assign _53125_ = _53126_ | _53128_ /*8534*/;
assign _53134_ = ~D[53] /*8533*/;
assign _53131_ = _52405_ & _53134_ /*8529*/;
assign _53132_ = _52405_ ^ _53134_ /*8532*/;
assign _53133_ = _53125_ & _53132_ /*8530*/;
assign _52854_ = _53125_ ^ _53132_ /*8531*/;
assign _53130_ = _53131_ | _53133_ /*8528*/;
assign _53139_ = ~D[54] /*8527*/;
assign _53136_ = _52406_ & _53139_ /*8523*/;
assign _53137_ = _52406_ ^ _53139_ /*8526*/;
assign _53138_ = _53130_ & _53137_ /*8524*/;
assign _52855_ = _53130_ ^ _53137_ /*8525*/;
assign _53135_ = _53136_ | _53138_ /*8522*/;
assign _53144_ = ~D[55] /*8521*/;
assign _53141_ = _52407_ & _53144_ /*8517*/;
assign _53142_ = _52407_ ^ _53144_ /*8520*/;
assign _53143_ = _53135_ & _53142_ /*8518*/;
assign _52856_ = _53135_ ^ _53142_ /*8519*/;
assign _53140_ = _53141_ | _53143_ /*8516*/;
assign _53149_ = ~D[56] /*8515*/;
assign _53146_ = _52408_ & _53149_ /*8511*/;
assign _53147_ = _52408_ ^ _53149_ /*8514*/;
assign _53148_ = _53140_ & _53147_ /*8512*/;
assign _52857_ = _53140_ ^ _53147_ /*8513*/;
assign _53145_ = _53146_ | _53148_ /*8510*/;
assign _53154_ = ~D[57] /*8509*/;
assign _53151_ = _52409_ & _53154_ /*8505*/;
assign _53152_ = _52409_ ^ _53154_ /*8508*/;
assign _53153_ = _53145_ & _53152_ /*8506*/;
assign _52858_ = _53145_ ^ _53152_ /*8507*/;
assign _53150_ = _53151_ | _53153_ /*8504*/;
assign _53159_ = ~D[58] /*8503*/;
assign _53156_ = _52410_ & _53159_ /*8499*/;
assign _53157_ = _52410_ ^ _53159_ /*8502*/;
assign _53158_ = _53150_ & _53157_ /*8500*/;
assign _52859_ = _53150_ ^ _53157_ /*8501*/;
assign _53155_ = _53156_ | _53158_ /*8498*/;
assign _53164_ = ~D[59] /*8497*/;
assign _53161_ = _52411_ & _53164_ /*8493*/;
assign _53162_ = _52411_ ^ _53164_ /*8496*/;
assign _53163_ = _53155_ & _53162_ /*8494*/;
assign _52860_ = _53155_ ^ _53162_ /*8495*/;
assign _53160_ = _53161_ | _53163_ /*8492*/;
assign _53169_ = ~D[60] /*8491*/;
assign _53166_ = _52412_ & _53169_ /*8487*/;
assign _53167_ = _52412_ ^ _53169_ /*8490*/;
assign _53168_ = _53160_ & _53167_ /*8488*/;
assign _52861_ = _53160_ ^ _53167_ /*8489*/;
assign _53165_ = _53166_ | _53168_ /*8486*/;
assign _53174_ = ~D[61] /*8485*/;
assign _53171_ = _52413_ & _53174_ /*8481*/;
assign _53172_ = _52413_ ^ _53174_ /*8484*/;
assign _53173_ = _53165_ & _53172_ /*8482*/;
assign _52862_ = _53165_ ^ _53172_ /*8483*/;
assign _53170_ = _53171_ | _53173_ /*8480*/;
assign _53179_ = ~D[62] /*8479*/;
assign _53176_ = _52414_ & _53179_ /*8475*/;
assign _53177_ = _52414_ ^ _53179_ /*8478*/;
assign _53178_ = _53170_ & _53177_ /*8476*/;
assign _52863_ = _53170_ ^ _53177_ /*8477*/;
assign _53175_ = _53176_ | _53178_ /*8474*/;
assign _53180_ = _52415_ & oneWire /*8469*/;
assign _53181_ = _52415_ ^ oneWire /*8472*/;
assign _53182_ = _53175_ & _53181_ /*8470*/;
assign _52864_ = _53175_ ^ _53181_ /*8471*/;
assign Q[4] = _53180_ | _53182_ /*8468*/;
assign _53315_ = ~Q[4] /*8083*/;
assign _53314_ = _53315_ & D[0] /*8082*/;
assign _53317_ = _52801_ & _53314_ /*8077*/;
assign _53318_ = _52801_ ^ _53314_ /*8080*/;
assign _53319_ = zeroWire & _53318_ /*8078*/;
assign _53249_ = zeroWire ^ _53318_ /*8079*/;
assign _53316_ = _53317_ | _53319_ /*8076*/;
assign _53321_ = ~Q[4] /*8075*/;
assign _53320_ = _53321_ & D[1] /*8074*/;
assign _53323_ = _52802_ & _53320_ /*8069*/;
assign _53324_ = _52802_ ^ _53320_ /*8072*/;
assign _53325_ = _53316_ & _53324_ /*8070*/;
assign _53250_ = _53316_ ^ _53324_ /*8071*/;
assign _53322_ = _53323_ | _53325_ /*8068*/;
assign _53327_ = ~Q[4] /*8067*/;
assign _53326_ = _53327_ & D[2] /*8066*/;
assign _53329_ = _52803_ & _53326_ /*8061*/;
assign _53330_ = _52803_ ^ _53326_ /*8064*/;
assign _53331_ = _53322_ & _53330_ /*8062*/;
assign _53251_ = _53322_ ^ _53330_ /*8063*/;
assign _53328_ = _53329_ | _53331_ /*8060*/;
assign _53333_ = ~Q[4] /*8059*/;
assign _53332_ = _53333_ & D[3] /*8058*/;
assign _53335_ = _52804_ & _53332_ /*8053*/;
assign _53336_ = _52804_ ^ _53332_ /*8056*/;
assign _53337_ = _53328_ & _53336_ /*8054*/;
assign _53252_ = _53328_ ^ _53336_ /*8055*/;
assign _53334_ = _53335_ | _53337_ /*8052*/;
assign _53339_ = ~Q[4] /*8051*/;
assign _53338_ = _53339_ & D[4] /*8050*/;
assign _53341_ = _52805_ & _53338_ /*8045*/;
assign _53342_ = _52805_ ^ _53338_ /*8048*/;
assign _53343_ = _53334_ & _53342_ /*8046*/;
assign _53253_ = _53334_ ^ _53342_ /*8047*/;
assign _53340_ = _53341_ | _53343_ /*8044*/;
assign _53345_ = ~Q[4] /*8043*/;
assign _53344_ = _53345_ & D[5] /*8042*/;
assign _53347_ = _52806_ & _53344_ /*8037*/;
assign _53348_ = _52806_ ^ _53344_ /*8040*/;
assign _53349_ = _53340_ & _53348_ /*8038*/;
assign _53254_ = _53340_ ^ _53348_ /*8039*/;
assign _53346_ = _53347_ | _53349_ /*8036*/;
assign _53351_ = ~Q[4] /*8035*/;
assign _53350_ = _53351_ & D[6] /*8034*/;
assign _53353_ = _52807_ & _53350_ /*8029*/;
assign _53354_ = _52807_ ^ _53350_ /*8032*/;
assign _53355_ = _53346_ & _53354_ /*8030*/;
assign _53255_ = _53346_ ^ _53354_ /*8031*/;
assign _53352_ = _53353_ | _53355_ /*8028*/;
assign _53357_ = ~Q[4] /*8027*/;
assign _53356_ = _53357_ & D[7] /*8026*/;
assign _53359_ = _52808_ & _53356_ /*8021*/;
assign _53360_ = _52808_ ^ _53356_ /*8024*/;
assign _53361_ = _53352_ & _53360_ /*8022*/;
assign _53256_ = _53352_ ^ _53360_ /*8023*/;
assign _53358_ = _53359_ | _53361_ /*8020*/;
assign _53363_ = ~Q[4] /*8019*/;
assign _53362_ = _53363_ & D[8] /*8018*/;
assign _53365_ = _52809_ & _53362_ /*8013*/;
assign _53366_ = _52809_ ^ _53362_ /*8016*/;
assign _53367_ = _53358_ & _53366_ /*8014*/;
assign _53257_ = _53358_ ^ _53366_ /*8015*/;
assign _53364_ = _53365_ | _53367_ /*8012*/;
assign _53369_ = ~Q[4] /*8011*/;
assign _53368_ = _53369_ & D[9] /*8010*/;
assign _53371_ = _52810_ & _53368_ /*8005*/;
assign _53372_ = _52810_ ^ _53368_ /*8008*/;
assign _53373_ = _53364_ & _53372_ /*8006*/;
assign _53258_ = _53364_ ^ _53372_ /*8007*/;
assign _53370_ = _53371_ | _53373_ /*8004*/;
assign _53375_ = ~Q[4] /*8003*/;
assign _53374_ = _53375_ & D[10] /*8002*/;
assign _53377_ = _52811_ & _53374_ /*7997*/;
assign _53378_ = _52811_ ^ _53374_ /*8000*/;
assign _53379_ = _53370_ & _53378_ /*7998*/;
assign _53259_ = _53370_ ^ _53378_ /*7999*/;
assign _53376_ = _53377_ | _53379_ /*7996*/;
assign _53381_ = ~Q[4] /*7995*/;
assign _53380_ = _53381_ & D[11] /*7994*/;
assign _53383_ = _52812_ & _53380_ /*7989*/;
assign _53384_ = _52812_ ^ _53380_ /*7992*/;
assign _53385_ = _53376_ & _53384_ /*7990*/;
assign _53260_ = _53376_ ^ _53384_ /*7991*/;
assign _53382_ = _53383_ | _53385_ /*7988*/;
assign _53387_ = ~Q[4] /*7987*/;
assign _53386_ = _53387_ & D[12] /*7986*/;
assign _53389_ = _52813_ & _53386_ /*7981*/;
assign _53390_ = _52813_ ^ _53386_ /*7984*/;
assign _53391_ = _53382_ & _53390_ /*7982*/;
assign _53261_ = _53382_ ^ _53390_ /*7983*/;
assign _53388_ = _53389_ | _53391_ /*7980*/;
assign _53393_ = ~Q[4] /*7979*/;
assign _53392_ = _53393_ & D[13] /*7978*/;
assign _53395_ = _52814_ & _53392_ /*7973*/;
assign _53396_ = _52814_ ^ _53392_ /*7976*/;
assign _53397_ = _53388_ & _53396_ /*7974*/;
assign _53262_ = _53388_ ^ _53396_ /*7975*/;
assign _53394_ = _53395_ | _53397_ /*7972*/;
assign _53399_ = ~Q[4] /*7971*/;
assign _53398_ = _53399_ & D[14] /*7970*/;
assign _53401_ = _52815_ & _53398_ /*7965*/;
assign _53402_ = _52815_ ^ _53398_ /*7968*/;
assign _53403_ = _53394_ & _53402_ /*7966*/;
assign _53263_ = _53394_ ^ _53402_ /*7967*/;
assign _53400_ = _53401_ | _53403_ /*7964*/;
assign _53405_ = ~Q[4] /*7963*/;
assign _53404_ = _53405_ & D[15] /*7962*/;
assign _53407_ = _52816_ & _53404_ /*7957*/;
assign _53408_ = _52816_ ^ _53404_ /*7960*/;
assign _53409_ = _53400_ & _53408_ /*7958*/;
assign _53264_ = _53400_ ^ _53408_ /*7959*/;
assign _53406_ = _53407_ | _53409_ /*7956*/;
assign _53411_ = ~Q[4] /*7955*/;
assign _53410_ = _53411_ & D[16] /*7954*/;
assign _53413_ = _52817_ & _53410_ /*7949*/;
assign _53414_ = _52817_ ^ _53410_ /*7952*/;
assign _53415_ = _53406_ & _53414_ /*7950*/;
assign _53265_ = _53406_ ^ _53414_ /*7951*/;
assign _53412_ = _53413_ | _53415_ /*7948*/;
assign _53417_ = ~Q[4] /*7947*/;
assign _53416_ = _53417_ & D[17] /*7946*/;
assign _53419_ = _52818_ & _53416_ /*7941*/;
assign _53420_ = _52818_ ^ _53416_ /*7944*/;
assign _53421_ = _53412_ & _53420_ /*7942*/;
assign _53266_ = _53412_ ^ _53420_ /*7943*/;
assign _53418_ = _53419_ | _53421_ /*7940*/;
assign _53423_ = ~Q[4] /*7939*/;
assign _53422_ = _53423_ & D[18] /*7938*/;
assign _53425_ = _52819_ & _53422_ /*7933*/;
assign _53426_ = _52819_ ^ _53422_ /*7936*/;
assign _53427_ = _53418_ & _53426_ /*7934*/;
assign _53267_ = _53418_ ^ _53426_ /*7935*/;
assign _53424_ = _53425_ | _53427_ /*7932*/;
assign _53429_ = ~Q[4] /*7931*/;
assign _53428_ = _53429_ & D[19] /*7930*/;
assign _53431_ = _52820_ & _53428_ /*7925*/;
assign _53432_ = _52820_ ^ _53428_ /*7928*/;
assign _53433_ = _53424_ & _53432_ /*7926*/;
assign _53268_ = _53424_ ^ _53432_ /*7927*/;
assign _53430_ = _53431_ | _53433_ /*7924*/;
assign _53435_ = ~Q[4] /*7923*/;
assign _53434_ = _53435_ & D[20] /*7922*/;
assign _53437_ = _52821_ & _53434_ /*7917*/;
assign _53438_ = _52821_ ^ _53434_ /*7920*/;
assign _53439_ = _53430_ & _53438_ /*7918*/;
assign _53269_ = _53430_ ^ _53438_ /*7919*/;
assign _53436_ = _53437_ | _53439_ /*7916*/;
assign _53441_ = ~Q[4] /*7915*/;
assign _53440_ = _53441_ & D[21] /*7914*/;
assign _53443_ = _52822_ & _53440_ /*7909*/;
assign _53444_ = _52822_ ^ _53440_ /*7912*/;
assign _53445_ = _53436_ & _53444_ /*7910*/;
assign _53270_ = _53436_ ^ _53444_ /*7911*/;
assign _53442_ = _53443_ | _53445_ /*7908*/;
assign _53447_ = ~Q[4] /*7907*/;
assign _53446_ = _53447_ & D[22] /*7906*/;
assign _53449_ = _52823_ & _53446_ /*7901*/;
assign _53450_ = _52823_ ^ _53446_ /*7904*/;
assign _53451_ = _53442_ & _53450_ /*7902*/;
assign _53271_ = _53442_ ^ _53450_ /*7903*/;
assign _53448_ = _53449_ | _53451_ /*7900*/;
assign _53453_ = ~Q[4] /*7899*/;
assign _53452_ = _53453_ & D[23] /*7898*/;
assign _53455_ = _52824_ & _53452_ /*7893*/;
assign _53456_ = _52824_ ^ _53452_ /*7896*/;
assign _53457_ = _53448_ & _53456_ /*7894*/;
assign _53272_ = _53448_ ^ _53456_ /*7895*/;
assign _53454_ = _53455_ | _53457_ /*7892*/;
assign _53459_ = ~Q[4] /*7891*/;
assign _53458_ = _53459_ & D[24] /*7890*/;
assign _53461_ = _52825_ & _53458_ /*7885*/;
assign _53462_ = _52825_ ^ _53458_ /*7888*/;
assign _53463_ = _53454_ & _53462_ /*7886*/;
assign _53273_ = _53454_ ^ _53462_ /*7887*/;
assign _53460_ = _53461_ | _53463_ /*7884*/;
assign _53465_ = ~Q[4] /*7883*/;
assign _53464_ = _53465_ & D[25] /*7882*/;
assign _53467_ = _52826_ & _53464_ /*7877*/;
assign _53468_ = _52826_ ^ _53464_ /*7880*/;
assign _53469_ = _53460_ & _53468_ /*7878*/;
assign _53274_ = _53460_ ^ _53468_ /*7879*/;
assign _53466_ = _53467_ | _53469_ /*7876*/;
assign _53471_ = ~Q[4] /*7875*/;
assign _53470_ = _53471_ & D[26] /*7874*/;
assign _53473_ = _52827_ & _53470_ /*7869*/;
assign _53474_ = _52827_ ^ _53470_ /*7872*/;
assign _53475_ = _53466_ & _53474_ /*7870*/;
assign _53275_ = _53466_ ^ _53474_ /*7871*/;
assign _53472_ = _53473_ | _53475_ /*7868*/;
assign _53477_ = ~Q[4] /*7867*/;
assign _53476_ = _53477_ & D[27] /*7866*/;
assign _53479_ = _52828_ & _53476_ /*7861*/;
assign _53480_ = _52828_ ^ _53476_ /*7864*/;
assign _53481_ = _53472_ & _53480_ /*7862*/;
assign _53276_ = _53472_ ^ _53480_ /*7863*/;
assign _53478_ = _53479_ | _53481_ /*7860*/;
assign _53483_ = ~Q[4] /*7859*/;
assign _53482_ = _53483_ & D[28] /*7858*/;
assign _53485_ = _52829_ & _53482_ /*7853*/;
assign _53486_ = _52829_ ^ _53482_ /*7856*/;
assign _53487_ = _53478_ & _53486_ /*7854*/;
assign _53277_ = _53478_ ^ _53486_ /*7855*/;
assign _53484_ = _53485_ | _53487_ /*7852*/;
assign _53489_ = ~Q[4] /*7851*/;
assign _53488_ = _53489_ & D[29] /*7850*/;
assign _53491_ = _52830_ & _53488_ /*7845*/;
assign _53492_ = _52830_ ^ _53488_ /*7848*/;
assign _53493_ = _53484_ & _53492_ /*7846*/;
assign _53278_ = _53484_ ^ _53492_ /*7847*/;
assign _53490_ = _53491_ | _53493_ /*7844*/;
assign _53495_ = ~Q[4] /*7843*/;
assign _53494_ = _53495_ & D[30] /*7842*/;
assign _53497_ = _52831_ & _53494_ /*7837*/;
assign _53498_ = _52831_ ^ _53494_ /*7840*/;
assign _53499_ = _53490_ & _53498_ /*7838*/;
assign _53279_ = _53490_ ^ _53498_ /*7839*/;
assign _53496_ = _53497_ | _53499_ /*7836*/;
assign _53501_ = ~Q[4] /*7835*/;
assign _53500_ = _53501_ & D[31] /*7834*/;
assign _53503_ = _52832_ & _53500_ /*7829*/;
assign _53504_ = _52832_ ^ _53500_ /*7832*/;
assign _53505_ = _53496_ & _53504_ /*7830*/;
assign _53280_ = _53496_ ^ _53504_ /*7831*/;
assign _53502_ = _53503_ | _53505_ /*7828*/;
assign _53507_ = ~Q[4] /*7827*/;
assign _53506_ = _53507_ & D[32] /*7826*/;
assign _53509_ = _52833_ & _53506_ /*7821*/;
assign _53510_ = _52833_ ^ _53506_ /*7824*/;
assign _53511_ = _53502_ & _53510_ /*7822*/;
assign _53281_ = _53502_ ^ _53510_ /*7823*/;
assign _53508_ = _53509_ | _53511_ /*7820*/;
assign _53513_ = ~Q[4] /*7819*/;
assign _53512_ = _53513_ & D[33] /*7818*/;
assign _53515_ = _52834_ & _53512_ /*7813*/;
assign _53516_ = _52834_ ^ _53512_ /*7816*/;
assign _53517_ = _53508_ & _53516_ /*7814*/;
assign _53282_ = _53508_ ^ _53516_ /*7815*/;
assign _53514_ = _53515_ | _53517_ /*7812*/;
assign _53519_ = ~Q[4] /*7811*/;
assign _53518_ = _53519_ & D[34] /*7810*/;
assign _53521_ = _52835_ & _53518_ /*7805*/;
assign _53522_ = _52835_ ^ _53518_ /*7808*/;
assign _53523_ = _53514_ & _53522_ /*7806*/;
assign _53283_ = _53514_ ^ _53522_ /*7807*/;
assign _53520_ = _53521_ | _53523_ /*7804*/;
assign _53525_ = ~Q[4] /*7803*/;
assign _53524_ = _53525_ & D[35] /*7802*/;
assign _53527_ = _52836_ & _53524_ /*7797*/;
assign _53528_ = _52836_ ^ _53524_ /*7800*/;
assign _53529_ = _53520_ & _53528_ /*7798*/;
assign _53284_ = _53520_ ^ _53528_ /*7799*/;
assign _53526_ = _53527_ | _53529_ /*7796*/;
assign _53531_ = ~Q[4] /*7795*/;
assign _53530_ = _53531_ & D[36] /*7794*/;
assign _53533_ = _52837_ & _53530_ /*7789*/;
assign _53534_ = _52837_ ^ _53530_ /*7792*/;
assign _53535_ = _53526_ & _53534_ /*7790*/;
assign _53285_ = _53526_ ^ _53534_ /*7791*/;
assign _53532_ = _53533_ | _53535_ /*7788*/;
assign _53537_ = ~Q[4] /*7787*/;
assign _53536_ = _53537_ & D[37] /*7786*/;
assign _53539_ = _52838_ & _53536_ /*7781*/;
assign _53540_ = _52838_ ^ _53536_ /*7784*/;
assign _53541_ = _53532_ & _53540_ /*7782*/;
assign _53286_ = _53532_ ^ _53540_ /*7783*/;
assign _53538_ = _53539_ | _53541_ /*7780*/;
assign _53543_ = ~Q[4] /*7779*/;
assign _53542_ = _53543_ & D[38] /*7778*/;
assign _53545_ = _52839_ & _53542_ /*7773*/;
assign _53546_ = _52839_ ^ _53542_ /*7776*/;
assign _53547_ = _53538_ & _53546_ /*7774*/;
assign _53287_ = _53538_ ^ _53546_ /*7775*/;
assign _53544_ = _53545_ | _53547_ /*7772*/;
assign _53549_ = ~Q[4] /*7771*/;
assign _53548_ = _53549_ & D[39] /*7770*/;
assign _53551_ = _52840_ & _53548_ /*7765*/;
assign _53552_ = _52840_ ^ _53548_ /*7768*/;
assign _53553_ = _53544_ & _53552_ /*7766*/;
assign _53288_ = _53544_ ^ _53552_ /*7767*/;
assign _53550_ = _53551_ | _53553_ /*7764*/;
assign _53555_ = ~Q[4] /*7763*/;
assign _53554_ = _53555_ & D[40] /*7762*/;
assign _53557_ = _52841_ & _53554_ /*7757*/;
assign _53558_ = _52841_ ^ _53554_ /*7760*/;
assign _53559_ = _53550_ & _53558_ /*7758*/;
assign _53289_ = _53550_ ^ _53558_ /*7759*/;
assign _53556_ = _53557_ | _53559_ /*7756*/;
assign _53561_ = ~Q[4] /*7755*/;
assign _53560_ = _53561_ & D[41] /*7754*/;
assign _53563_ = _52842_ & _53560_ /*7749*/;
assign _53564_ = _52842_ ^ _53560_ /*7752*/;
assign _53565_ = _53556_ & _53564_ /*7750*/;
assign _53290_ = _53556_ ^ _53564_ /*7751*/;
assign _53562_ = _53563_ | _53565_ /*7748*/;
assign _53567_ = ~Q[4] /*7747*/;
assign _53566_ = _53567_ & D[42] /*7746*/;
assign _53569_ = _52843_ & _53566_ /*7741*/;
assign _53570_ = _52843_ ^ _53566_ /*7744*/;
assign _53571_ = _53562_ & _53570_ /*7742*/;
assign _53291_ = _53562_ ^ _53570_ /*7743*/;
assign _53568_ = _53569_ | _53571_ /*7740*/;
assign _53573_ = ~Q[4] /*7739*/;
assign _53572_ = _53573_ & D[43] /*7738*/;
assign _53575_ = _52844_ & _53572_ /*7733*/;
assign _53576_ = _52844_ ^ _53572_ /*7736*/;
assign _53577_ = _53568_ & _53576_ /*7734*/;
assign _53292_ = _53568_ ^ _53576_ /*7735*/;
assign _53574_ = _53575_ | _53577_ /*7732*/;
assign _53579_ = ~Q[4] /*7731*/;
assign _53578_ = _53579_ & D[44] /*7730*/;
assign _53581_ = _52845_ & _53578_ /*7725*/;
assign _53582_ = _52845_ ^ _53578_ /*7728*/;
assign _53583_ = _53574_ & _53582_ /*7726*/;
assign _53293_ = _53574_ ^ _53582_ /*7727*/;
assign _53580_ = _53581_ | _53583_ /*7724*/;
assign _53585_ = ~Q[4] /*7723*/;
assign _53584_ = _53585_ & D[45] /*7722*/;
assign _53587_ = _52846_ & _53584_ /*7717*/;
assign _53588_ = _52846_ ^ _53584_ /*7720*/;
assign _53589_ = _53580_ & _53588_ /*7718*/;
assign _53294_ = _53580_ ^ _53588_ /*7719*/;
assign _53586_ = _53587_ | _53589_ /*7716*/;
assign _53591_ = ~Q[4] /*7715*/;
assign _53590_ = _53591_ & D[46] /*7714*/;
assign _53593_ = _52847_ & _53590_ /*7709*/;
assign _53594_ = _52847_ ^ _53590_ /*7712*/;
assign _53595_ = _53586_ & _53594_ /*7710*/;
assign _53295_ = _53586_ ^ _53594_ /*7711*/;
assign _53592_ = _53593_ | _53595_ /*7708*/;
assign _53597_ = ~Q[4] /*7707*/;
assign _53596_ = _53597_ & D[47] /*7706*/;
assign _53599_ = _52848_ & _53596_ /*7701*/;
assign _53600_ = _52848_ ^ _53596_ /*7704*/;
assign _53601_ = _53592_ & _53600_ /*7702*/;
assign _53296_ = _53592_ ^ _53600_ /*7703*/;
assign _53598_ = _53599_ | _53601_ /*7700*/;
assign _53603_ = ~Q[4] /*7699*/;
assign _53602_ = _53603_ & D[48] /*7698*/;
assign _53605_ = _52849_ & _53602_ /*7693*/;
assign _53606_ = _52849_ ^ _53602_ /*7696*/;
assign _53607_ = _53598_ & _53606_ /*7694*/;
assign _53297_ = _53598_ ^ _53606_ /*7695*/;
assign _53604_ = _53605_ | _53607_ /*7692*/;
assign _53609_ = ~Q[4] /*7691*/;
assign _53608_ = _53609_ & D[49] /*7690*/;
assign _53611_ = _52850_ & _53608_ /*7685*/;
assign _53612_ = _52850_ ^ _53608_ /*7688*/;
assign _53613_ = _53604_ & _53612_ /*7686*/;
assign _53298_ = _53604_ ^ _53612_ /*7687*/;
assign _53610_ = _53611_ | _53613_ /*7684*/;
assign _53615_ = ~Q[4] /*7683*/;
assign _53614_ = _53615_ & D[50] /*7682*/;
assign _53617_ = _52851_ & _53614_ /*7677*/;
assign _53618_ = _52851_ ^ _53614_ /*7680*/;
assign _53619_ = _53610_ & _53618_ /*7678*/;
assign _53299_ = _53610_ ^ _53618_ /*7679*/;
assign _53616_ = _53617_ | _53619_ /*7676*/;
assign _53621_ = ~Q[4] /*7675*/;
assign _53620_ = _53621_ & D[51] /*7674*/;
assign _53623_ = _52852_ & _53620_ /*7669*/;
assign _53624_ = _52852_ ^ _53620_ /*7672*/;
assign _53625_ = _53616_ & _53624_ /*7670*/;
assign _53300_ = _53616_ ^ _53624_ /*7671*/;
assign _53622_ = _53623_ | _53625_ /*7668*/;
assign _53627_ = ~Q[4] /*7667*/;
assign _53626_ = _53627_ & D[52] /*7666*/;
assign _53629_ = _52853_ & _53626_ /*7661*/;
assign _53630_ = _52853_ ^ _53626_ /*7664*/;
assign _53631_ = _53622_ & _53630_ /*7662*/;
assign _53301_ = _53622_ ^ _53630_ /*7663*/;
assign _53628_ = _53629_ | _53631_ /*7660*/;
assign _53633_ = ~Q[4] /*7659*/;
assign _53632_ = _53633_ & D[53] /*7658*/;
assign _53635_ = _52854_ & _53632_ /*7653*/;
assign _53636_ = _52854_ ^ _53632_ /*7656*/;
assign _53637_ = _53628_ & _53636_ /*7654*/;
assign _53302_ = _53628_ ^ _53636_ /*7655*/;
assign _53634_ = _53635_ | _53637_ /*7652*/;
assign _53639_ = ~Q[4] /*7651*/;
assign _53638_ = _53639_ & D[54] /*7650*/;
assign _53641_ = _52855_ & _53638_ /*7645*/;
assign _53642_ = _52855_ ^ _53638_ /*7648*/;
assign _53643_ = _53634_ & _53642_ /*7646*/;
assign _53303_ = _53634_ ^ _53642_ /*7647*/;
assign _53640_ = _53641_ | _53643_ /*7644*/;
assign _53645_ = ~Q[4] /*7643*/;
assign _53644_ = _53645_ & D[55] /*7642*/;
assign _53647_ = _52856_ & _53644_ /*7637*/;
assign _53648_ = _52856_ ^ _53644_ /*7640*/;
assign _53649_ = _53640_ & _53648_ /*7638*/;
assign _53304_ = _53640_ ^ _53648_ /*7639*/;
assign _53646_ = _53647_ | _53649_ /*7636*/;
assign _53651_ = ~Q[4] /*7635*/;
assign _53650_ = _53651_ & D[56] /*7634*/;
assign _53653_ = _52857_ & _53650_ /*7629*/;
assign _53654_ = _52857_ ^ _53650_ /*7632*/;
assign _53655_ = _53646_ & _53654_ /*7630*/;
assign _53305_ = _53646_ ^ _53654_ /*7631*/;
assign _53652_ = _53653_ | _53655_ /*7628*/;
assign _53657_ = ~Q[4] /*7627*/;
assign _53656_ = _53657_ & D[57] /*7626*/;
assign _53659_ = _52858_ & _53656_ /*7621*/;
assign _53660_ = _52858_ ^ _53656_ /*7624*/;
assign _53661_ = _53652_ & _53660_ /*7622*/;
assign _53306_ = _53652_ ^ _53660_ /*7623*/;
assign _53658_ = _53659_ | _53661_ /*7620*/;
assign _53663_ = ~Q[4] /*7619*/;
assign _53662_ = _53663_ & D[58] /*7618*/;
assign _53665_ = _52859_ & _53662_ /*7613*/;
assign _53666_ = _52859_ ^ _53662_ /*7616*/;
assign _53667_ = _53658_ & _53666_ /*7614*/;
assign _53307_ = _53658_ ^ _53666_ /*7615*/;
assign _53664_ = _53665_ | _53667_ /*7612*/;
assign _53669_ = ~Q[4] /*7611*/;
assign _53668_ = _53669_ & D[59] /*7610*/;
assign _53671_ = _52860_ & _53668_ /*7605*/;
assign _53672_ = _52860_ ^ _53668_ /*7608*/;
assign _53673_ = _53664_ & _53672_ /*7606*/;
assign _53308_ = _53664_ ^ _53672_ /*7607*/;
assign _53670_ = _53671_ | _53673_ /*7604*/;
assign _53675_ = ~Q[4] /*7603*/;
assign _53674_ = _53675_ & D[60] /*7602*/;
assign _53677_ = _52861_ & _53674_ /*7597*/;
assign _53678_ = _52861_ ^ _53674_ /*7600*/;
assign _53679_ = _53670_ & _53678_ /*7598*/;
assign _53309_ = _53670_ ^ _53678_ /*7599*/;
assign _53676_ = _53677_ | _53679_ /*7596*/;
assign _53681_ = ~Q[4] /*7595*/;
assign _53680_ = _53681_ & D[61] /*7594*/;
assign _53683_ = _52862_ & _53680_ /*7589*/;
assign _53684_ = _52862_ ^ _53680_ /*7592*/;
assign _53685_ = _53676_ & _53684_ /*7590*/;
assign _53310_ = _53676_ ^ _53684_ /*7591*/;
assign _53682_ = _53683_ | _53685_ /*7588*/;
assign _53687_ = ~Q[4] /*7587*/;
assign _53686_ = _53687_ & D[62] /*7586*/;
assign _53689_ = _52863_ & _53686_ /*7581*/;
assign _53690_ = _52863_ ^ _53686_ /*7584*/;
assign _53691_ = _53682_ & _53690_ /*7582*/;
assign _53311_ = _53682_ ^ _53690_ /*7583*/;
assign _53688_ = _53689_ | _53691_ /*7580*/;
assign _53693_ = ~Q[4] /*7579*/;
assign _53692_ = _53693_ & zeroWire /*7578*/;
assign _53694_ = _52864_ ^ _53692_ /*7576*/;
assign _53312_ = _53694_ ^ _53688_ /*7575*/;
assign _53765_ = ~D[0] /*7321*/;
assign _53762_ = R_0[3] & _53765_ /*7317*/;
assign _53763_ = R_0[3] ^ _53765_ /*7320*/;
assign _53764_ = oneWire & _53763_ /*7318*/;
assign _53697_ = oneWire ^ _53763_ /*7319*/;
assign _53761_ = _53762_ | _53764_ /*7316*/;
assign _53770_ = ~D[1] /*7315*/;
assign _53767_ = _53249_ & _53770_ /*7311*/;
assign _53768_ = _53249_ ^ _53770_ /*7314*/;
assign _53769_ = _53761_ & _53768_ /*7312*/;
assign _53698_ = _53761_ ^ _53768_ /*7313*/;
assign _53766_ = _53767_ | _53769_ /*7310*/;
assign _53775_ = ~D[2] /*7309*/;
assign _53772_ = _53250_ & _53775_ /*7305*/;
assign _53773_ = _53250_ ^ _53775_ /*7308*/;
assign _53774_ = _53766_ & _53773_ /*7306*/;
assign _53699_ = _53766_ ^ _53773_ /*7307*/;
assign _53771_ = _53772_ | _53774_ /*7304*/;
assign _53780_ = ~D[3] /*7303*/;
assign _53777_ = _53251_ & _53780_ /*7299*/;
assign _53778_ = _53251_ ^ _53780_ /*7302*/;
assign _53779_ = _53771_ & _53778_ /*7300*/;
assign _53700_ = _53771_ ^ _53778_ /*7301*/;
assign _53776_ = _53777_ | _53779_ /*7298*/;
assign _53785_ = ~D[4] /*7297*/;
assign _53782_ = _53252_ & _53785_ /*7293*/;
assign _53783_ = _53252_ ^ _53785_ /*7296*/;
assign _53784_ = _53776_ & _53783_ /*7294*/;
assign _53701_ = _53776_ ^ _53783_ /*7295*/;
assign _53781_ = _53782_ | _53784_ /*7292*/;
assign _53790_ = ~D[5] /*7291*/;
assign _53787_ = _53253_ & _53790_ /*7287*/;
assign _53788_ = _53253_ ^ _53790_ /*7290*/;
assign _53789_ = _53781_ & _53788_ /*7288*/;
assign _53702_ = _53781_ ^ _53788_ /*7289*/;
assign _53786_ = _53787_ | _53789_ /*7286*/;
assign _53795_ = ~D[6] /*7285*/;
assign _53792_ = _53254_ & _53795_ /*7281*/;
assign _53793_ = _53254_ ^ _53795_ /*7284*/;
assign _53794_ = _53786_ & _53793_ /*7282*/;
assign _53703_ = _53786_ ^ _53793_ /*7283*/;
assign _53791_ = _53792_ | _53794_ /*7280*/;
assign _53800_ = ~D[7] /*7279*/;
assign _53797_ = _53255_ & _53800_ /*7275*/;
assign _53798_ = _53255_ ^ _53800_ /*7278*/;
assign _53799_ = _53791_ & _53798_ /*7276*/;
assign _53704_ = _53791_ ^ _53798_ /*7277*/;
assign _53796_ = _53797_ | _53799_ /*7274*/;
assign _53805_ = ~D[8] /*7273*/;
assign _53802_ = _53256_ & _53805_ /*7269*/;
assign _53803_ = _53256_ ^ _53805_ /*7272*/;
assign _53804_ = _53796_ & _53803_ /*7270*/;
assign _53705_ = _53796_ ^ _53803_ /*7271*/;
assign _53801_ = _53802_ | _53804_ /*7268*/;
assign _53810_ = ~D[9] /*7267*/;
assign _53807_ = _53257_ & _53810_ /*7263*/;
assign _53808_ = _53257_ ^ _53810_ /*7266*/;
assign _53809_ = _53801_ & _53808_ /*7264*/;
assign _53706_ = _53801_ ^ _53808_ /*7265*/;
assign _53806_ = _53807_ | _53809_ /*7262*/;
assign _53815_ = ~D[10] /*7261*/;
assign _53812_ = _53258_ & _53815_ /*7257*/;
assign _53813_ = _53258_ ^ _53815_ /*7260*/;
assign _53814_ = _53806_ & _53813_ /*7258*/;
assign _53707_ = _53806_ ^ _53813_ /*7259*/;
assign _53811_ = _53812_ | _53814_ /*7256*/;
assign _53820_ = ~D[11] /*7255*/;
assign _53817_ = _53259_ & _53820_ /*7251*/;
assign _53818_ = _53259_ ^ _53820_ /*7254*/;
assign _53819_ = _53811_ & _53818_ /*7252*/;
assign _53708_ = _53811_ ^ _53818_ /*7253*/;
assign _53816_ = _53817_ | _53819_ /*7250*/;
assign _53825_ = ~D[12] /*7249*/;
assign _53822_ = _53260_ & _53825_ /*7245*/;
assign _53823_ = _53260_ ^ _53825_ /*7248*/;
assign _53824_ = _53816_ & _53823_ /*7246*/;
assign _53709_ = _53816_ ^ _53823_ /*7247*/;
assign _53821_ = _53822_ | _53824_ /*7244*/;
assign _53830_ = ~D[13] /*7243*/;
assign _53827_ = _53261_ & _53830_ /*7239*/;
assign _53828_ = _53261_ ^ _53830_ /*7242*/;
assign _53829_ = _53821_ & _53828_ /*7240*/;
assign _53710_ = _53821_ ^ _53828_ /*7241*/;
assign _53826_ = _53827_ | _53829_ /*7238*/;
assign _53835_ = ~D[14] /*7237*/;
assign _53832_ = _53262_ & _53835_ /*7233*/;
assign _53833_ = _53262_ ^ _53835_ /*7236*/;
assign _53834_ = _53826_ & _53833_ /*7234*/;
assign _53711_ = _53826_ ^ _53833_ /*7235*/;
assign _53831_ = _53832_ | _53834_ /*7232*/;
assign _53840_ = ~D[15] /*7231*/;
assign _53837_ = _53263_ & _53840_ /*7227*/;
assign _53838_ = _53263_ ^ _53840_ /*7230*/;
assign _53839_ = _53831_ & _53838_ /*7228*/;
assign _53712_ = _53831_ ^ _53838_ /*7229*/;
assign _53836_ = _53837_ | _53839_ /*7226*/;
assign _53845_ = ~D[16] /*7225*/;
assign _53842_ = _53264_ & _53845_ /*7221*/;
assign _53843_ = _53264_ ^ _53845_ /*7224*/;
assign _53844_ = _53836_ & _53843_ /*7222*/;
assign _53713_ = _53836_ ^ _53843_ /*7223*/;
assign _53841_ = _53842_ | _53844_ /*7220*/;
assign _53850_ = ~D[17] /*7219*/;
assign _53847_ = _53265_ & _53850_ /*7215*/;
assign _53848_ = _53265_ ^ _53850_ /*7218*/;
assign _53849_ = _53841_ & _53848_ /*7216*/;
assign _53714_ = _53841_ ^ _53848_ /*7217*/;
assign _53846_ = _53847_ | _53849_ /*7214*/;
assign _53855_ = ~D[18] /*7213*/;
assign _53852_ = _53266_ & _53855_ /*7209*/;
assign _53853_ = _53266_ ^ _53855_ /*7212*/;
assign _53854_ = _53846_ & _53853_ /*7210*/;
assign _53715_ = _53846_ ^ _53853_ /*7211*/;
assign _53851_ = _53852_ | _53854_ /*7208*/;
assign _53860_ = ~D[19] /*7207*/;
assign _53857_ = _53267_ & _53860_ /*7203*/;
assign _53858_ = _53267_ ^ _53860_ /*7206*/;
assign _53859_ = _53851_ & _53858_ /*7204*/;
assign _53716_ = _53851_ ^ _53858_ /*7205*/;
assign _53856_ = _53857_ | _53859_ /*7202*/;
assign _53865_ = ~D[20] /*7201*/;
assign _53862_ = _53268_ & _53865_ /*7197*/;
assign _53863_ = _53268_ ^ _53865_ /*7200*/;
assign _53864_ = _53856_ & _53863_ /*7198*/;
assign _53717_ = _53856_ ^ _53863_ /*7199*/;
assign _53861_ = _53862_ | _53864_ /*7196*/;
assign _53870_ = ~D[21] /*7195*/;
assign _53867_ = _53269_ & _53870_ /*7191*/;
assign _53868_ = _53269_ ^ _53870_ /*7194*/;
assign _53869_ = _53861_ & _53868_ /*7192*/;
assign _53718_ = _53861_ ^ _53868_ /*7193*/;
assign _53866_ = _53867_ | _53869_ /*7190*/;
assign _53875_ = ~D[22] /*7189*/;
assign _53872_ = _53270_ & _53875_ /*7185*/;
assign _53873_ = _53270_ ^ _53875_ /*7188*/;
assign _53874_ = _53866_ & _53873_ /*7186*/;
assign _53719_ = _53866_ ^ _53873_ /*7187*/;
assign _53871_ = _53872_ | _53874_ /*7184*/;
assign _53880_ = ~D[23] /*7183*/;
assign _53877_ = _53271_ & _53880_ /*7179*/;
assign _53878_ = _53271_ ^ _53880_ /*7182*/;
assign _53879_ = _53871_ & _53878_ /*7180*/;
assign _53720_ = _53871_ ^ _53878_ /*7181*/;
assign _53876_ = _53877_ | _53879_ /*7178*/;
assign _53885_ = ~D[24] /*7177*/;
assign _53882_ = _53272_ & _53885_ /*7173*/;
assign _53883_ = _53272_ ^ _53885_ /*7176*/;
assign _53884_ = _53876_ & _53883_ /*7174*/;
assign _53721_ = _53876_ ^ _53883_ /*7175*/;
assign _53881_ = _53882_ | _53884_ /*7172*/;
assign _53890_ = ~D[25] /*7171*/;
assign _53887_ = _53273_ & _53890_ /*7167*/;
assign _53888_ = _53273_ ^ _53890_ /*7170*/;
assign _53889_ = _53881_ & _53888_ /*7168*/;
assign _53722_ = _53881_ ^ _53888_ /*7169*/;
assign _53886_ = _53887_ | _53889_ /*7166*/;
assign _53895_ = ~D[26] /*7165*/;
assign _53892_ = _53274_ & _53895_ /*7161*/;
assign _53893_ = _53274_ ^ _53895_ /*7164*/;
assign _53894_ = _53886_ & _53893_ /*7162*/;
assign _53723_ = _53886_ ^ _53893_ /*7163*/;
assign _53891_ = _53892_ | _53894_ /*7160*/;
assign _53900_ = ~D[27] /*7159*/;
assign _53897_ = _53275_ & _53900_ /*7155*/;
assign _53898_ = _53275_ ^ _53900_ /*7158*/;
assign _53899_ = _53891_ & _53898_ /*7156*/;
assign _53724_ = _53891_ ^ _53898_ /*7157*/;
assign _53896_ = _53897_ | _53899_ /*7154*/;
assign _53905_ = ~D[28] /*7153*/;
assign _53902_ = _53276_ & _53905_ /*7149*/;
assign _53903_ = _53276_ ^ _53905_ /*7152*/;
assign _53904_ = _53896_ & _53903_ /*7150*/;
assign _53725_ = _53896_ ^ _53903_ /*7151*/;
assign _53901_ = _53902_ | _53904_ /*7148*/;
assign _53910_ = ~D[29] /*7147*/;
assign _53907_ = _53277_ & _53910_ /*7143*/;
assign _53908_ = _53277_ ^ _53910_ /*7146*/;
assign _53909_ = _53901_ & _53908_ /*7144*/;
assign _53726_ = _53901_ ^ _53908_ /*7145*/;
assign _53906_ = _53907_ | _53909_ /*7142*/;
assign _53915_ = ~D[30] /*7141*/;
assign _53912_ = _53278_ & _53915_ /*7137*/;
assign _53913_ = _53278_ ^ _53915_ /*7140*/;
assign _53914_ = _53906_ & _53913_ /*7138*/;
assign _53727_ = _53906_ ^ _53913_ /*7139*/;
assign _53911_ = _53912_ | _53914_ /*7136*/;
assign _53920_ = ~D[31] /*7135*/;
assign _53917_ = _53279_ & _53920_ /*7131*/;
assign _53918_ = _53279_ ^ _53920_ /*7134*/;
assign _53919_ = _53911_ & _53918_ /*7132*/;
assign _53728_ = _53911_ ^ _53918_ /*7133*/;
assign _53916_ = _53917_ | _53919_ /*7130*/;
assign _53925_ = ~D[32] /*7129*/;
assign _53922_ = _53280_ & _53925_ /*7125*/;
assign _53923_ = _53280_ ^ _53925_ /*7128*/;
assign _53924_ = _53916_ & _53923_ /*7126*/;
assign _53729_ = _53916_ ^ _53923_ /*7127*/;
assign _53921_ = _53922_ | _53924_ /*7124*/;
assign _53930_ = ~D[33] /*7123*/;
assign _53927_ = _53281_ & _53930_ /*7119*/;
assign _53928_ = _53281_ ^ _53930_ /*7122*/;
assign _53929_ = _53921_ & _53928_ /*7120*/;
assign _53730_ = _53921_ ^ _53928_ /*7121*/;
assign _53926_ = _53927_ | _53929_ /*7118*/;
assign _53935_ = ~D[34] /*7117*/;
assign _53932_ = _53282_ & _53935_ /*7113*/;
assign _53933_ = _53282_ ^ _53935_ /*7116*/;
assign _53934_ = _53926_ & _53933_ /*7114*/;
assign _53731_ = _53926_ ^ _53933_ /*7115*/;
assign _53931_ = _53932_ | _53934_ /*7112*/;
assign _53940_ = ~D[35] /*7111*/;
assign _53937_ = _53283_ & _53940_ /*7107*/;
assign _53938_ = _53283_ ^ _53940_ /*7110*/;
assign _53939_ = _53931_ & _53938_ /*7108*/;
assign _53732_ = _53931_ ^ _53938_ /*7109*/;
assign _53936_ = _53937_ | _53939_ /*7106*/;
assign _53945_ = ~D[36] /*7105*/;
assign _53942_ = _53284_ & _53945_ /*7101*/;
assign _53943_ = _53284_ ^ _53945_ /*7104*/;
assign _53944_ = _53936_ & _53943_ /*7102*/;
assign _53733_ = _53936_ ^ _53943_ /*7103*/;
assign _53941_ = _53942_ | _53944_ /*7100*/;
assign _53950_ = ~D[37] /*7099*/;
assign _53947_ = _53285_ & _53950_ /*7095*/;
assign _53948_ = _53285_ ^ _53950_ /*7098*/;
assign _53949_ = _53941_ & _53948_ /*7096*/;
assign _53734_ = _53941_ ^ _53948_ /*7097*/;
assign _53946_ = _53947_ | _53949_ /*7094*/;
assign _53955_ = ~D[38] /*7093*/;
assign _53952_ = _53286_ & _53955_ /*7089*/;
assign _53953_ = _53286_ ^ _53955_ /*7092*/;
assign _53954_ = _53946_ & _53953_ /*7090*/;
assign _53735_ = _53946_ ^ _53953_ /*7091*/;
assign _53951_ = _53952_ | _53954_ /*7088*/;
assign _53960_ = ~D[39] /*7087*/;
assign _53957_ = _53287_ & _53960_ /*7083*/;
assign _53958_ = _53287_ ^ _53960_ /*7086*/;
assign _53959_ = _53951_ & _53958_ /*7084*/;
assign _53736_ = _53951_ ^ _53958_ /*7085*/;
assign _53956_ = _53957_ | _53959_ /*7082*/;
assign _53965_ = ~D[40] /*7081*/;
assign _53962_ = _53288_ & _53965_ /*7077*/;
assign _53963_ = _53288_ ^ _53965_ /*7080*/;
assign _53964_ = _53956_ & _53963_ /*7078*/;
assign _53737_ = _53956_ ^ _53963_ /*7079*/;
assign _53961_ = _53962_ | _53964_ /*7076*/;
assign _53970_ = ~D[41] /*7075*/;
assign _53967_ = _53289_ & _53970_ /*7071*/;
assign _53968_ = _53289_ ^ _53970_ /*7074*/;
assign _53969_ = _53961_ & _53968_ /*7072*/;
assign _53738_ = _53961_ ^ _53968_ /*7073*/;
assign _53966_ = _53967_ | _53969_ /*7070*/;
assign _53975_ = ~D[42] /*7069*/;
assign _53972_ = _53290_ & _53975_ /*7065*/;
assign _53973_ = _53290_ ^ _53975_ /*7068*/;
assign _53974_ = _53966_ & _53973_ /*7066*/;
assign _53739_ = _53966_ ^ _53973_ /*7067*/;
assign _53971_ = _53972_ | _53974_ /*7064*/;
assign _53980_ = ~D[43] /*7063*/;
assign _53977_ = _53291_ & _53980_ /*7059*/;
assign _53978_ = _53291_ ^ _53980_ /*7062*/;
assign _53979_ = _53971_ & _53978_ /*7060*/;
assign _53740_ = _53971_ ^ _53978_ /*7061*/;
assign _53976_ = _53977_ | _53979_ /*7058*/;
assign _53985_ = ~D[44] /*7057*/;
assign _53982_ = _53292_ & _53985_ /*7053*/;
assign _53983_ = _53292_ ^ _53985_ /*7056*/;
assign _53984_ = _53976_ & _53983_ /*7054*/;
assign _53741_ = _53976_ ^ _53983_ /*7055*/;
assign _53981_ = _53982_ | _53984_ /*7052*/;
assign _53990_ = ~D[45] /*7051*/;
assign _53987_ = _53293_ & _53990_ /*7047*/;
assign _53988_ = _53293_ ^ _53990_ /*7050*/;
assign _53989_ = _53981_ & _53988_ /*7048*/;
assign _53742_ = _53981_ ^ _53988_ /*7049*/;
assign _53986_ = _53987_ | _53989_ /*7046*/;
assign _53995_ = ~D[46] /*7045*/;
assign _53992_ = _53294_ & _53995_ /*7041*/;
assign _53993_ = _53294_ ^ _53995_ /*7044*/;
assign _53994_ = _53986_ & _53993_ /*7042*/;
assign _53743_ = _53986_ ^ _53993_ /*7043*/;
assign _53991_ = _53992_ | _53994_ /*7040*/;
assign _54000_ = ~D[47] /*7039*/;
assign _53997_ = _53295_ & _54000_ /*7035*/;
assign _53998_ = _53295_ ^ _54000_ /*7038*/;
assign _53999_ = _53991_ & _53998_ /*7036*/;
assign _53744_ = _53991_ ^ _53998_ /*7037*/;
assign _53996_ = _53997_ | _53999_ /*7034*/;
assign _54005_ = ~D[48] /*7033*/;
assign _54002_ = _53296_ & _54005_ /*7029*/;
assign _54003_ = _53296_ ^ _54005_ /*7032*/;
assign _54004_ = _53996_ & _54003_ /*7030*/;
assign _53745_ = _53996_ ^ _54003_ /*7031*/;
assign _54001_ = _54002_ | _54004_ /*7028*/;
assign _54010_ = ~D[49] /*7027*/;
assign _54007_ = _53297_ & _54010_ /*7023*/;
assign _54008_ = _53297_ ^ _54010_ /*7026*/;
assign _54009_ = _54001_ & _54008_ /*7024*/;
assign _53746_ = _54001_ ^ _54008_ /*7025*/;
assign _54006_ = _54007_ | _54009_ /*7022*/;
assign _54015_ = ~D[50] /*7021*/;
assign _54012_ = _53298_ & _54015_ /*7017*/;
assign _54013_ = _53298_ ^ _54015_ /*7020*/;
assign _54014_ = _54006_ & _54013_ /*7018*/;
assign _53747_ = _54006_ ^ _54013_ /*7019*/;
assign _54011_ = _54012_ | _54014_ /*7016*/;
assign _54020_ = ~D[51] /*7015*/;
assign _54017_ = _53299_ & _54020_ /*7011*/;
assign _54018_ = _53299_ ^ _54020_ /*7014*/;
assign _54019_ = _54011_ & _54018_ /*7012*/;
assign _53748_ = _54011_ ^ _54018_ /*7013*/;
assign _54016_ = _54017_ | _54019_ /*7010*/;
assign _54025_ = ~D[52] /*7009*/;
assign _54022_ = _53300_ & _54025_ /*7005*/;
assign _54023_ = _53300_ ^ _54025_ /*7008*/;
assign _54024_ = _54016_ & _54023_ /*7006*/;
assign _53749_ = _54016_ ^ _54023_ /*7007*/;
assign _54021_ = _54022_ | _54024_ /*7004*/;
assign _54030_ = ~D[53] /*7003*/;
assign _54027_ = _53301_ & _54030_ /*6999*/;
assign _54028_ = _53301_ ^ _54030_ /*7002*/;
assign _54029_ = _54021_ & _54028_ /*7000*/;
assign _53750_ = _54021_ ^ _54028_ /*7001*/;
assign _54026_ = _54027_ | _54029_ /*6998*/;
assign _54035_ = ~D[54] /*6997*/;
assign _54032_ = _53302_ & _54035_ /*6993*/;
assign _54033_ = _53302_ ^ _54035_ /*6996*/;
assign _54034_ = _54026_ & _54033_ /*6994*/;
assign _53751_ = _54026_ ^ _54033_ /*6995*/;
assign _54031_ = _54032_ | _54034_ /*6992*/;
assign _54040_ = ~D[55] /*6991*/;
assign _54037_ = _53303_ & _54040_ /*6987*/;
assign _54038_ = _53303_ ^ _54040_ /*6990*/;
assign _54039_ = _54031_ & _54038_ /*6988*/;
assign _53752_ = _54031_ ^ _54038_ /*6989*/;
assign _54036_ = _54037_ | _54039_ /*6986*/;
assign _54045_ = ~D[56] /*6985*/;
assign _54042_ = _53304_ & _54045_ /*6981*/;
assign _54043_ = _53304_ ^ _54045_ /*6984*/;
assign _54044_ = _54036_ & _54043_ /*6982*/;
assign _53753_ = _54036_ ^ _54043_ /*6983*/;
assign _54041_ = _54042_ | _54044_ /*6980*/;
assign _54050_ = ~D[57] /*6979*/;
assign _54047_ = _53305_ & _54050_ /*6975*/;
assign _54048_ = _53305_ ^ _54050_ /*6978*/;
assign _54049_ = _54041_ & _54048_ /*6976*/;
assign _53754_ = _54041_ ^ _54048_ /*6977*/;
assign _54046_ = _54047_ | _54049_ /*6974*/;
assign _54055_ = ~D[58] /*6973*/;
assign _54052_ = _53306_ & _54055_ /*6969*/;
assign _54053_ = _53306_ ^ _54055_ /*6972*/;
assign _54054_ = _54046_ & _54053_ /*6970*/;
assign _53755_ = _54046_ ^ _54053_ /*6971*/;
assign _54051_ = _54052_ | _54054_ /*6968*/;
assign _54060_ = ~D[59] /*6967*/;
assign _54057_ = _53307_ & _54060_ /*6963*/;
assign _54058_ = _53307_ ^ _54060_ /*6966*/;
assign _54059_ = _54051_ & _54058_ /*6964*/;
assign _53756_ = _54051_ ^ _54058_ /*6965*/;
assign _54056_ = _54057_ | _54059_ /*6962*/;
assign _54065_ = ~D[60] /*6961*/;
assign _54062_ = _53308_ & _54065_ /*6957*/;
assign _54063_ = _53308_ ^ _54065_ /*6960*/;
assign _54064_ = _54056_ & _54063_ /*6958*/;
assign _53757_ = _54056_ ^ _54063_ /*6959*/;
assign _54061_ = _54062_ | _54064_ /*6956*/;
assign _54070_ = ~D[61] /*6955*/;
assign _54067_ = _53309_ & _54070_ /*6951*/;
assign _54068_ = _53309_ ^ _54070_ /*6954*/;
assign _54069_ = _54061_ & _54068_ /*6952*/;
assign _53758_ = _54061_ ^ _54068_ /*6953*/;
assign _54066_ = _54067_ | _54069_ /*6950*/;
assign _54075_ = ~D[62] /*6949*/;
assign _54072_ = _53310_ & _54075_ /*6945*/;
assign _54073_ = _53310_ ^ _54075_ /*6948*/;
assign _54074_ = _54066_ & _54073_ /*6946*/;
assign _53759_ = _54066_ ^ _54073_ /*6947*/;
assign _54071_ = _54072_ | _54074_ /*6944*/;
assign _54076_ = _53311_ & oneWire /*6939*/;
assign _54077_ = _53311_ ^ oneWire /*6942*/;
assign _54078_ = _54071_ & _54077_ /*6940*/;
assign _53760_ = _54071_ ^ _54077_ /*6941*/;
assign Q[3] = _54076_ | _54078_ /*6938*/;
assign _54211_ = ~Q[3] /*6553*/;
assign _54210_ = _54211_ & D[0] /*6552*/;
assign _54213_ = _53697_ & _54210_ /*6547*/;
assign _54214_ = _53697_ ^ _54210_ /*6550*/;
assign _54215_ = zeroWire & _54214_ /*6548*/;
assign _54145_ = zeroWire ^ _54214_ /*6549*/;
assign _54212_ = _54213_ | _54215_ /*6546*/;
assign _54217_ = ~Q[3] /*6545*/;
assign _54216_ = _54217_ & D[1] /*6544*/;
assign _54219_ = _53698_ & _54216_ /*6539*/;
assign _54220_ = _53698_ ^ _54216_ /*6542*/;
assign _54221_ = _54212_ & _54220_ /*6540*/;
assign _54146_ = _54212_ ^ _54220_ /*6541*/;
assign _54218_ = _54219_ | _54221_ /*6538*/;
assign _54223_ = ~Q[3] /*6537*/;
assign _54222_ = _54223_ & D[2] /*6536*/;
assign _54225_ = _53699_ & _54222_ /*6531*/;
assign _54226_ = _53699_ ^ _54222_ /*6534*/;
assign _54227_ = _54218_ & _54226_ /*6532*/;
assign _54147_ = _54218_ ^ _54226_ /*6533*/;
assign _54224_ = _54225_ | _54227_ /*6530*/;
assign _54229_ = ~Q[3] /*6529*/;
assign _54228_ = _54229_ & D[3] /*6528*/;
assign _54231_ = _53700_ & _54228_ /*6523*/;
assign _54232_ = _53700_ ^ _54228_ /*6526*/;
assign _54233_ = _54224_ & _54232_ /*6524*/;
assign _54148_ = _54224_ ^ _54232_ /*6525*/;
assign _54230_ = _54231_ | _54233_ /*6522*/;
assign _54235_ = ~Q[3] /*6521*/;
assign _54234_ = _54235_ & D[4] /*6520*/;
assign _54237_ = _53701_ & _54234_ /*6515*/;
assign _54238_ = _53701_ ^ _54234_ /*6518*/;
assign _54239_ = _54230_ & _54238_ /*6516*/;
assign _54149_ = _54230_ ^ _54238_ /*6517*/;
assign _54236_ = _54237_ | _54239_ /*6514*/;
assign _54241_ = ~Q[3] /*6513*/;
assign _54240_ = _54241_ & D[5] /*6512*/;
assign _54243_ = _53702_ & _54240_ /*6507*/;
assign _54244_ = _53702_ ^ _54240_ /*6510*/;
assign _54245_ = _54236_ & _54244_ /*6508*/;
assign _54150_ = _54236_ ^ _54244_ /*6509*/;
assign _54242_ = _54243_ | _54245_ /*6506*/;
assign _54247_ = ~Q[3] /*6505*/;
assign _54246_ = _54247_ & D[6] /*6504*/;
assign _54249_ = _53703_ & _54246_ /*6499*/;
assign _54250_ = _53703_ ^ _54246_ /*6502*/;
assign _54251_ = _54242_ & _54250_ /*6500*/;
assign _54151_ = _54242_ ^ _54250_ /*6501*/;
assign _54248_ = _54249_ | _54251_ /*6498*/;
assign _54253_ = ~Q[3] /*6497*/;
assign _54252_ = _54253_ & D[7] /*6496*/;
assign _54255_ = _53704_ & _54252_ /*6491*/;
assign _54256_ = _53704_ ^ _54252_ /*6494*/;
assign _54257_ = _54248_ & _54256_ /*6492*/;
assign _54152_ = _54248_ ^ _54256_ /*6493*/;
assign _54254_ = _54255_ | _54257_ /*6490*/;
assign _54259_ = ~Q[3] /*6489*/;
assign _54258_ = _54259_ & D[8] /*6488*/;
assign _54261_ = _53705_ & _54258_ /*6483*/;
assign _54262_ = _53705_ ^ _54258_ /*6486*/;
assign _54263_ = _54254_ & _54262_ /*6484*/;
assign _54153_ = _54254_ ^ _54262_ /*6485*/;
assign _54260_ = _54261_ | _54263_ /*6482*/;
assign _54265_ = ~Q[3] /*6481*/;
assign _54264_ = _54265_ & D[9] /*6480*/;
assign _54267_ = _53706_ & _54264_ /*6475*/;
assign _54268_ = _53706_ ^ _54264_ /*6478*/;
assign _54269_ = _54260_ & _54268_ /*6476*/;
assign _54154_ = _54260_ ^ _54268_ /*6477*/;
assign _54266_ = _54267_ | _54269_ /*6474*/;
assign _54271_ = ~Q[3] /*6473*/;
assign _54270_ = _54271_ & D[10] /*6472*/;
assign _54273_ = _53707_ & _54270_ /*6467*/;
assign _54274_ = _53707_ ^ _54270_ /*6470*/;
assign _54275_ = _54266_ & _54274_ /*6468*/;
assign _54155_ = _54266_ ^ _54274_ /*6469*/;
assign _54272_ = _54273_ | _54275_ /*6466*/;
assign _54277_ = ~Q[3] /*6465*/;
assign _54276_ = _54277_ & D[11] /*6464*/;
assign _54279_ = _53708_ & _54276_ /*6459*/;
assign _54280_ = _53708_ ^ _54276_ /*6462*/;
assign _54281_ = _54272_ & _54280_ /*6460*/;
assign _54156_ = _54272_ ^ _54280_ /*6461*/;
assign _54278_ = _54279_ | _54281_ /*6458*/;
assign _54283_ = ~Q[3] /*6457*/;
assign _54282_ = _54283_ & D[12] /*6456*/;
assign _54285_ = _53709_ & _54282_ /*6451*/;
assign _54286_ = _53709_ ^ _54282_ /*6454*/;
assign _54287_ = _54278_ & _54286_ /*6452*/;
assign _54157_ = _54278_ ^ _54286_ /*6453*/;
assign _54284_ = _54285_ | _54287_ /*6450*/;
assign _54289_ = ~Q[3] /*6449*/;
assign _54288_ = _54289_ & D[13] /*6448*/;
assign _54291_ = _53710_ & _54288_ /*6443*/;
assign _54292_ = _53710_ ^ _54288_ /*6446*/;
assign _54293_ = _54284_ & _54292_ /*6444*/;
assign _54158_ = _54284_ ^ _54292_ /*6445*/;
assign _54290_ = _54291_ | _54293_ /*6442*/;
assign _54295_ = ~Q[3] /*6441*/;
assign _54294_ = _54295_ & D[14] /*6440*/;
assign _54297_ = _53711_ & _54294_ /*6435*/;
assign _54298_ = _53711_ ^ _54294_ /*6438*/;
assign _54299_ = _54290_ & _54298_ /*6436*/;
assign _54159_ = _54290_ ^ _54298_ /*6437*/;
assign _54296_ = _54297_ | _54299_ /*6434*/;
assign _54301_ = ~Q[3] /*6433*/;
assign _54300_ = _54301_ & D[15] /*6432*/;
assign _54303_ = _53712_ & _54300_ /*6427*/;
assign _54304_ = _53712_ ^ _54300_ /*6430*/;
assign _54305_ = _54296_ & _54304_ /*6428*/;
assign _54160_ = _54296_ ^ _54304_ /*6429*/;
assign _54302_ = _54303_ | _54305_ /*6426*/;
assign _54307_ = ~Q[3] /*6425*/;
assign _54306_ = _54307_ & D[16] /*6424*/;
assign _54309_ = _53713_ & _54306_ /*6419*/;
assign _54310_ = _53713_ ^ _54306_ /*6422*/;
assign _54311_ = _54302_ & _54310_ /*6420*/;
assign _54161_ = _54302_ ^ _54310_ /*6421*/;
assign _54308_ = _54309_ | _54311_ /*6418*/;
assign _54313_ = ~Q[3] /*6417*/;
assign _54312_ = _54313_ & D[17] /*6416*/;
assign _54315_ = _53714_ & _54312_ /*6411*/;
assign _54316_ = _53714_ ^ _54312_ /*6414*/;
assign _54317_ = _54308_ & _54316_ /*6412*/;
assign _54162_ = _54308_ ^ _54316_ /*6413*/;
assign _54314_ = _54315_ | _54317_ /*6410*/;
assign _54319_ = ~Q[3] /*6409*/;
assign _54318_ = _54319_ & D[18] /*6408*/;
assign _54321_ = _53715_ & _54318_ /*6403*/;
assign _54322_ = _53715_ ^ _54318_ /*6406*/;
assign _54323_ = _54314_ & _54322_ /*6404*/;
assign _54163_ = _54314_ ^ _54322_ /*6405*/;
assign _54320_ = _54321_ | _54323_ /*6402*/;
assign _54325_ = ~Q[3] /*6401*/;
assign _54324_ = _54325_ & D[19] /*6400*/;
assign _54327_ = _53716_ & _54324_ /*6395*/;
assign _54328_ = _53716_ ^ _54324_ /*6398*/;
assign _54329_ = _54320_ & _54328_ /*6396*/;
assign _54164_ = _54320_ ^ _54328_ /*6397*/;
assign _54326_ = _54327_ | _54329_ /*6394*/;
assign _54331_ = ~Q[3] /*6393*/;
assign _54330_ = _54331_ & D[20] /*6392*/;
assign _54333_ = _53717_ & _54330_ /*6387*/;
assign _54334_ = _53717_ ^ _54330_ /*6390*/;
assign _54335_ = _54326_ & _54334_ /*6388*/;
assign _54165_ = _54326_ ^ _54334_ /*6389*/;
assign _54332_ = _54333_ | _54335_ /*6386*/;
assign _54337_ = ~Q[3] /*6385*/;
assign _54336_ = _54337_ & D[21] /*6384*/;
assign _54339_ = _53718_ & _54336_ /*6379*/;
assign _54340_ = _53718_ ^ _54336_ /*6382*/;
assign _54341_ = _54332_ & _54340_ /*6380*/;
assign _54166_ = _54332_ ^ _54340_ /*6381*/;
assign _54338_ = _54339_ | _54341_ /*6378*/;
assign _54343_ = ~Q[3] /*6377*/;
assign _54342_ = _54343_ & D[22] /*6376*/;
assign _54345_ = _53719_ & _54342_ /*6371*/;
assign _54346_ = _53719_ ^ _54342_ /*6374*/;
assign _54347_ = _54338_ & _54346_ /*6372*/;
assign _54167_ = _54338_ ^ _54346_ /*6373*/;
assign _54344_ = _54345_ | _54347_ /*6370*/;
assign _54349_ = ~Q[3] /*6369*/;
assign _54348_ = _54349_ & D[23] /*6368*/;
assign _54351_ = _53720_ & _54348_ /*6363*/;
assign _54352_ = _53720_ ^ _54348_ /*6366*/;
assign _54353_ = _54344_ & _54352_ /*6364*/;
assign _54168_ = _54344_ ^ _54352_ /*6365*/;
assign _54350_ = _54351_ | _54353_ /*6362*/;
assign _54355_ = ~Q[3] /*6361*/;
assign _54354_ = _54355_ & D[24] /*6360*/;
assign _54357_ = _53721_ & _54354_ /*6355*/;
assign _54358_ = _53721_ ^ _54354_ /*6358*/;
assign _54359_ = _54350_ & _54358_ /*6356*/;
assign _54169_ = _54350_ ^ _54358_ /*6357*/;
assign _54356_ = _54357_ | _54359_ /*6354*/;
assign _54361_ = ~Q[3] /*6353*/;
assign _54360_ = _54361_ & D[25] /*6352*/;
assign _54363_ = _53722_ & _54360_ /*6347*/;
assign _54364_ = _53722_ ^ _54360_ /*6350*/;
assign _54365_ = _54356_ & _54364_ /*6348*/;
assign _54170_ = _54356_ ^ _54364_ /*6349*/;
assign _54362_ = _54363_ | _54365_ /*6346*/;
assign _54367_ = ~Q[3] /*6345*/;
assign _54366_ = _54367_ & D[26] /*6344*/;
assign _54369_ = _53723_ & _54366_ /*6339*/;
assign _54370_ = _53723_ ^ _54366_ /*6342*/;
assign _54371_ = _54362_ & _54370_ /*6340*/;
assign _54171_ = _54362_ ^ _54370_ /*6341*/;
assign _54368_ = _54369_ | _54371_ /*6338*/;
assign _54373_ = ~Q[3] /*6337*/;
assign _54372_ = _54373_ & D[27] /*6336*/;
assign _54375_ = _53724_ & _54372_ /*6331*/;
assign _54376_ = _53724_ ^ _54372_ /*6334*/;
assign _54377_ = _54368_ & _54376_ /*6332*/;
assign _54172_ = _54368_ ^ _54376_ /*6333*/;
assign _54374_ = _54375_ | _54377_ /*6330*/;
assign _54379_ = ~Q[3] /*6329*/;
assign _54378_ = _54379_ & D[28] /*6328*/;
assign _54381_ = _53725_ & _54378_ /*6323*/;
assign _54382_ = _53725_ ^ _54378_ /*6326*/;
assign _54383_ = _54374_ & _54382_ /*6324*/;
assign _54173_ = _54374_ ^ _54382_ /*6325*/;
assign _54380_ = _54381_ | _54383_ /*6322*/;
assign _54385_ = ~Q[3] /*6321*/;
assign _54384_ = _54385_ & D[29] /*6320*/;
assign _54387_ = _53726_ & _54384_ /*6315*/;
assign _54388_ = _53726_ ^ _54384_ /*6318*/;
assign _54389_ = _54380_ & _54388_ /*6316*/;
assign _54174_ = _54380_ ^ _54388_ /*6317*/;
assign _54386_ = _54387_ | _54389_ /*6314*/;
assign _54391_ = ~Q[3] /*6313*/;
assign _54390_ = _54391_ & D[30] /*6312*/;
assign _54393_ = _53727_ & _54390_ /*6307*/;
assign _54394_ = _53727_ ^ _54390_ /*6310*/;
assign _54395_ = _54386_ & _54394_ /*6308*/;
assign _54175_ = _54386_ ^ _54394_ /*6309*/;
assign _54392_ = _54393_ | _54395_ /*6306*/;
assign _54397_ = ~Q[3] /*6305*/;
assign _54396_ = _54397_ & D[31] /*6304*/;
assign _54399_ = _53728_ & _54396_ /*6299*/;
assign _54400_ = _53728_ ^ _54396_ /*6302*/;
assign _54401_ = _54392_ & _54400_ /*6300*/;
assign _54176_ = _54392_ ^ _54400_ /*6301*/;
assign _54398_ = _54399_ | _54401_ /*6298*/;
assign _54403_ = ~Q[3] /*6297*/;
assign _54402_ = _54403_ & D[32] /*6296*/;
assign _54405_ = _53729_ & _54402_ /*6291*/;
assign _54406_ = _53729_ ^ _54402_ /*6294*/;
assign _54407_ = _54398_ & _54406_ /*6292*/;
assign _54177_ = _54398_ ^ _54406_ /*6293*/;
assign _54404_ = _54405_ | _54407_ /*6290*/;
assign _54409_ = ~Q[3] /*6289*/;
assign _54408_ = _54409_ & D[33] /*6288*/;
assign _54411_ = _53730_ & _54408_ /*6283*/;
assign _54412_ = _53730_ ^ _54408_ /*6286*/;
assign _54413_ = _54404_ & _54412_ /*6284*/;
assign _54178_ = _54404_ ^ _54412_ /*6285*/;
assign _54410_ = _54411_ | _54413_ /*6282*/;
assign _54415_ = ~Q[3] /*6281*/;
assign _54414_ = _54415_ & D[34] /*6280*/;
assign _54417_ = _53731_ & _54414_ /*6275*/;
assign _54418_ = _53731_ ^ _54414_ /*6278*/;
assign _54419_ = _54410_ & _54418_ /*6276*/;
assign _54179_ = _54410_ ^ _54418_ /*6277*/;
assign _54416_ = _54417_ | _54419_ /*6274*/;
assign _54421_ = ~Q[3] /*6273*/;
assign _54420_ = _54421_ & D[35] /*6272*/;
assign _54423_ = _53732_ & _54420_ /*6267*/;
assign _54424_ = _53732_ ^ _54420_ /*6270*/;
assign _54425_ = _54416_ & _54424_ /*6268*/;
assign _54180_ = _54416_ ^ _54424_ /*6269*/;
assign _54422_ = _54423_ | _54425_ /*6266*/;
assign _54427_ = ~Q[3] /*6265*/;
assign _54426_ = _54427_ & D[36] /*6264*/;
assign _54429_ = _53733_ & _54426_ /*6259*/;
assign _54430_ = _53733_ ^ _54426_ /*6262*/;
assign _54431_ = _54422_ & _54430_ /*6260*/;
assign _54181_ = _54422_ ^ _54430_ /*6261*/;
assign _54428_ = _54429_ | _54431_ /*6258*/;
assign _54433_ = ~Q[3] /*6257*/;
assign _54432_ = _54433_ & D[37] /*6256*/;
assign _54435_ = _53734_ & _54432_ /*6251*/;
assign _54436_ = _53734_ ^ _54432_ /*6254*/;
assign _54437_ = _54428_ & _54436_ /*6252*/;
assign _54182_ = _54428_ ^ _54436_ /*6253*/;
assign _54434_ = _54435_ | _54437_ /*6250*/;
assign _54439_ = ~Q[3] /*6249*/;
assign _54438_ = _54439_ & D[38] /*6248*/;
assign _54441_ = _53735_ & _54438_ /*6243*/;
assign _54442_ = _53735_ ^ _54438_ /*6246*/;
assign _54443_ = _54434_ & _54442_ /*6244*/;
assign _54183_ = _54434_ ^ _54442_ /*6245*/;
assign _54440_ = _54441_ | _54443_ /*6242*/;
assign _54445_ = ~Q[3] /*6241*/;
assign _54444_ = _54445_ & D[39] /*6240*/;
assign _54447_ = _53736_ & _54444_ /*6235*/;
assign _54448_ = _53736_ ^ _54444_ /*6238*/;
assign _54449_ = _54440_ & _54448_ /*6236*/;
assign _54184_ = _54440_ ^ _54448_ /*6237*/;
assign _54446_ = _54447_ | _54449_ /*6234*/;
assign _54451_ = ~Q[3] /*6233*/;
assign _54450_ = _54451_ & D[40] /*6232*/;
assign _54453_ = _53737_ & _54450_ /*6227*/;
assign _54454_ = _53737_ ^ _54450_ /*6230*/;
assign _54455_ = _54446_ & _54454_ /*6228*/;
assign _54185_ = _54446_ ^ _54454_ /*6229*/;
assign _54452_ = _54453_ | _54455_ /*6226*/;
assign _54457_ = ~Q[3] /*6225*/;
assign _54456_ = _54457_ & D[41] /*6224*/;
assign _54459_ = _53738_ & _54456_ /*6219*/;
assign _54460_ = _53738_ ^ _54456_ /*6222*/;
assign _54461_ = _54452_ & _54460_ /*6220*/;
assign _54186_ = _54452_ ^ _54460_ /*6221*/;
assign _54458_ = _54459_ | _54461_ /*6218*/;
assign _54463_ = ~Q[3] /*6217*/;
assign _54462_ = _54463_ & D[42] /*6216*/;
assign _54465_ = _53739_ & _54462_ /*6211*/;
assign _54466_ = _53739_ ^ _54462_ /*6214*/;
assign _54467_ = _54458_ & _54466_ /*6212*/;
assign _54187_ = _54458_ ^ _54466_ /*6213*/;
assign _54464_ = _54465_ | _54467_ /*6210*/;
assign _54469_ = ~Q[3] /*6209*/;
assign _54468_ = _54469_ & D[43] /*6208*/;
assign _54471_ = _53740_ & _54468_ /*6203*/;
assign _54472_ = _53740_ ^ _54468_ /*6206*/;
assign _54473_ = _54464_ & _54472_ /*6204*/;
assign _54188_ = _54464_ ^ _54472_ /*6205*/;
assign _54470_ = _54471_ | _54473_ /*6202*/;
assign _54475_ = ~Q[3] /*6201*/;
assign _54474_ = _54475_ & D[44] /*6200*/;
assign _54477_ = _53741_ & _54474_ /*6195*/;
assign _54478_ = _53741_ ^ _54474_ /*6198*/;
assign _54479_ = _54470_ & _54478_ /*6196*/;
assign _54189_ = _54470_ ^ _54478_ /*6197*/;
assign _54476_ = _54477_ | _54479_ /*6194*/;
assign _54481_ = ~Q[3] /*6193*/;
assign _54480_ = _54481_ & D[45] /*6192*/;
assign _54483_ = _53742_ & _54480_ /*6187*/;
assign _54484_ = _53742_ ^ _54480_ /*6190*/;
assign _54485_ = _54476_ & _54484_ /*6188*/;
assign _54190_ = _54476_ ^ _54484_ /*6189*/;
assign _54482_ = _54483_ | _54485_ /*6186*/;
assign _54487_ = ~Q[3] /*6185*/;
assign _54486_ = _54487_ & D[46] /*6184*/;
assign _54489_ = _53743_ & _54486_ /*6179*/;
assign _54490_ = _53743_ ^ _54486_ /*6182*/;
assign _54491_ = _54482_ & _54490_ /*6180*/;
assign _54191_ = _54482_ ^ _54490_ /*6181*/;
assign _54488_ = _54489_ | _54491_ /*6178*/;
assign _54493_ = ~Q[3] /*6177*/;
assign _54492_ = _54493_ & D[47] /*6176*/;
assign _54495_ = _53744_ & _54492_ /*6171*/;
assign _54496_ = _53744_ ^ _54492_ /*6174*/;
assign _54497_ = _54488_ & _54496_ /*6172*/;
assign _54192_ = _54488_ ^ _54496_ /*6173*/;
assign _54494_ = _54495_ | _54497_ /*6170*/;
assign _54499_ = ~Q[3] /*6169*/;
assign _54498_ = _54499_ & D[48] /*6168*/;
assign _54501_ = _53745_ & _54498_ /*6163*/;
assign _54502_ = _53745_ ^ _54498_ /*6166*/;
assign _54503_ = _54494_ & _54502_ /*6164*/;
assign _54193_ = _54494_ ^ _54502_ /*6165*/;
assign _54500_ = _54501_ | _54503_ /*6162*/;
assign _54505_ = ~Q[3] /*6161*/;
assign _54504_ = _54505_ & D[49] /*6160*/;
assign _54507_ = _53746_ & _54504_ /*6155*/;
assign _54508_ = _53746_ ^ _54504_ /*6158*/;
assign _54509_ = _54500_ & _54508_ /*6156*/;
assign _54194_ = _54500_ ^ _54508_ /*6157*/;
assign _54506_ = _54507_ | _54509_ /*6154*/;
assign _54511_ = ~Q[3] /*6153*/;
assign _54510_ = _54511_ & D[50] /*6152*/;
assign _54513_ = _53747_ & _54510_ /*6147*/;
assign _54514_ = _53747_ ^ _54510_ /*6150*/;
assign _54515_ = _54506_ & _54514_ /*6148*/;
assign _54195_ = _54506_ ^ _54514_ /*6149*/;
assign _54512_ = _54513_ | _54515_ /*6146*/;
assign _54517_ = ~Q[3] /*6145*/;
assign _54516_ = _54517_ & D[51] /*6144*/;
assign _54519_ = _53748_ & _54516_ /*6139*/;
assign _54520_ = _53748_ ^ _54516_ /*6142*/;
assign _54521_ = _54512_ & _54520_ /*6140*/;
assign _54196_ = _54512_ ^ _54520_ /*6141*/;
assign _54518_ = _54519_ | _54521_ /*6138*/;
assign _54523_ = ~Q[3] /*6137*/;
assign _54522_ = _54523_ & D[52] /*6136*/;
assign _54525_ = _53749_ & _54522_ /*6131*/;
assign _54526_ = _53749_ ^ _54522_ /*6134*/;
assign _54527_ = _54518_ & _54526_ /*6132*/;
assign _54197_ = _54518_ ^ _54526_ /*6133*/;
assign _54524_ = _54525_ | _54527_ /*6130*/;
assign _54529_ = ~Q[3] /*6129*/;
assign _54528_ = _54529_ & D[53] /*6128*/;
assign _54531_ = _53750_ & _54528_ /*6123*/;
assign _54532_ = _53750_ ^ _54528_ /*6126*/;
assign _54533_ = _54524_ & _54532_ /*6124*/;
assign _54198_ = _54524_ ^ _54532_ /*6125*/;
assign _54530_ = _54531_ | _54533_ /*6122*/;
assign _54535_ = ~Q[3] /*6121*/;
assign _54534_ = _54535_ & D[54] /*6120*/;
assign _54537_ = _53751_ & _54534_ /*6115*/;
assign _54538_ = _53751_ ^ _54534_ /*6118*/;
assign _54539_ = _54530_ & _54538_ /*6116*/;
assign _54199_ = _54530_ ^ _54538_ /*6117*/;
assign _54536_ = _54537_ | _54539_ /*6114*/;
assign _54541_ = ~Q[3] /*6113*/;
assign _54540_ = _54541_ & D[55] /*6112*/;
assign _54543_ = _53752_ & _54540_ /*6107*/;
assign _54544_ = _53752_ ^ _54540_ /*6110*/;
assign _54545_ = _54536_ & _54544_ /*6108*/;
assign _54200_ = _54536_ ^ _54544_ /*6109*/;
assign _54542_ = _54543_ | _54545_ /*6106*/;
assign _54547_ = ~Q[3] /*6105*/;
assign _54546_ = _54547_ & D[56] /*6104*/;
assign _54549_ = _53753_ & _54546_ /*6099*/;
assign _54550_ = _53753_ ^ _54546_ /*6102*/;
assign _54551_ = _54542_ & _54550_ /*6100*/;
assign _54201_ = _54542_ ^ _54550_ /*6101*/;
assign _54548_ = _54549_ | _54551_ /*6098*/;
assign _54553_ = ~Q[3] /*6097*/;
assign _54552_ = _54553_ & D[57] /*6096*/;
assign _54555_ = _53754_ & _54552_ /*6091*/;
assign _54556_ = _53754_ ^ _54552_ /*6094*/;
assign _54557_ = _54548_ & _54556_ /*6092*/;
assign _54202_ = _54548_ ^ _54556_ /*6093*/;
assign _54554_ = _54555_ | _54557_ /*6090*/;
assign _54559_ = ~Q[3] /*6089*/;
assign _54558_ = _54559_ & D[58] /*6088*/;
assign _54561_ = _53755_ & _54558_ /*6083*/;
assign _54562_ = _53755_ ^ _54558_ /*6086*/;
assign _54563_ = _54554_ & _54562_ /*6084*/;
assign _54203_ = _54554_ ^ _54562_ /*6085*/;
assign _54560_ = _54561_ | _54563_ /*6082*/;
assign _54565_ = ~Q[3] /*6081*/;
assign _54564_ = _54565_ & D[59] /*6080*/;
assign _54567_ = _53756_ & _54564_ /*6075*/;
assign _54568_ = _53756_ ^ _54564_ /*6078*/;
assign _54569_ = _54560_ & _54568_ /*6076*/;
assign _54204_ = _54560_ ^ _54568_ /*6077*/;
assign _54566_ = _54567_ | _54569_ /*6074*/;
assign _54571_ = ~Q[3] /*6073*/;
assign _54570_ = _54571_ & D[60] /*6072*/;
assign _54573_ = _53757_ & _54570_ /*6067*/;
assign _54574_ = _53757_ ^ _54570_ /*6070*/;
assign _54575_ = _54566_ & _54574_ /*6068*/;
assign _54205_ = _54566_ ^ _54574_ /*6069*/;
assign _54572_ = _54573_ | _54575_ /*6066*/;
assign _54577_ = ~Q[3] /*6065*/;
assign _54576_ = _54577_ & D[61] /*6064*/;
assign _54579_ = _53758_ & _54576_ /*6059*/;
assign _54580_ = _53758_ ^ _54576_ /*6062*/;
assign _54581_ = _54572_ & _54580_ /*6060*/;
assign _54206_ = _54572_ ^ _54580_ /*6061*/;
assign _54578_ = _54579_ | _54581_ /*6058*/;
assign _54583_ = ~Q[3] /*6057*/;
assign _54582_ = _54583_ & D[62] /*6056*/;
assign _54585_ = _53759_ & _54582_ /*6051*/;
assign _54586_ = _53759_ ^ _54582_ /*6054*/;
assign _54587_ = _54578_ & _54586_ /*6052*/;
assign _54207_ = _54578_ ^ _54586_ /*6053*/;
assign _54584_ = _54585_ | _54587_ /*6050*/;
assign _54589_ = ~Q[3] /*6049*/;
assign _54588_ = _54589_ & zeroWire /*6048*/;
assign _54590_ = _53760_ ^ _54588_ /*6046*/;
assign _54208_ = _54590_ ^ _54584_ /*6045*/;
assign _54661_ = ~D[0] /*5791*/;
assign _54658_ = R_0[2] & _54661_ /*5787*/;
assign _54659_ = R_0[2] ^ _54661_ /*5790*/;
assign _54660_ = oneWire & _54659_ /*5788*/;
assign _54593_ = oneWire ^ _54659_ /*5789*/;
assign _54657_ = _54658_ | _54660_ /*5786*/;
assign _54666_ = ~D[1] /*5785*/;
assign _54663_ = _54145_ & _54666_ /*5781*/;
assign _54664_ = _54145_ ^ _54666_ /*5784*/;
assign _54665_ = _54657_ & _54664_ /*5782*/;
assign _54594_ = _54657_ ^ _54664_ /*5783*/;
assign _54662_ = _54663_ | _54665_ /*5780*/;
assign _54671_ = ~D[2] /*5779*/;
assign _54668_ = _54146_ & _54671_ /*5775*/;
assign _54669_ = _54146_ ^ _54671_ /*5778*/;
assign _54670_ = _54662_ & _54669_ /*5776*/;
assign _54595_ = _54662_ ^ _54669_ /*5777*/;
assign _54667_ = _54668_ | _54670_ /*5774*/;
assign _54676_ = ~D[3] /*5773*/;
assign _54673_ = _54147_ & _54676_ /*5769*/;
assign _54674_ = _54147_ ^ _54676_ /*5772*/;
assign _54675_ = _54667_ & _54674_ /*5770*/;
assign _54596_ = _54667_ ^ _54674_ /*5771*/;
assign _54672_ = _54673_ | _54675_ /*5768*/;
assign _54681_ = ~D[4] /*5767*/;
assign _54678_ = _54148_ & _54681_ /*5763*/;
assign _54679_ = _54148_ ^ _54681_ /*5766*/;
assign _54680_ = _54672_ & _54679_ /*5764*/;
assign _54597_ = _54672_ ^ _54679_ /*5765*/;
assign _54677_ = _54678_ | _54680_ /*5762*/;
assign _54686_ = ~D[5] /*5761*/;
assign _54683_ = _54149_ & _54686_ /*5757*/;
assign _54684_ = _54149_ ^ _54686_ /*5760*/;
assign _54685_ = _54677_ & _54684_ /*5758*/;
assign _54598_ = _54677_ ^ _54684_ /*5759*/;
assign _54682_ = _54683_ | _54685_ /*5756*/;
assign _54691_ = ~D[6] /*5755*/;
assign _54688_ = _54150_ & _54691_ /*5751*/;
assign _54689_ = _54150_ ^ _54691_ /*5754*/;
assign _54690_ = _54682_ & _54689_ /*5752*/;
assign _54599_ = _54682_ ^ _54689_ /*5753*/;
assign _54687_ = _54688_ | _54690_ /*5750*/;
assign _54696_ = ~D[7] /*5749*/;
assign _54693_ = _54151_ & _54696_ /*5745*/;
assign _54694_ = _54151_ ^ _54696_ /*5748*/;
assign _54695_ = _54687_ & _54694_ /*5746*/;
assign _54600_ = _54687_ ^ _54694_ /*5747*/;
assign _54692_ = _54693_ | _54695_ /*5744*/;
assign _54701_ = ~D[8] /*5743*/;
assign _54698_ = _54152_ & _54701_ /*5739*/;
assign _54699_ = _54152_ ^ _54701_ /*5742*/;
assign _54700_ = _54692_ & _54699_ /*5740*/;
assign _54601_ = _54692_ ^ _54699_ /*5741*/;
assign _54697_ = _54698_ | _54700_ /*5738*/;
assign _54706_ = ~D[9] /*5737*/;
assign _54703_ = _54153_ & _54706_ /*5733*/;
assign _54704_ = _54153_ ^ _54706_ /*5736*/;
assign _54705_ = _54697_ & _54704_ /*5734*/;
assign _54602_ = _54697_ ^ _54704_ /*5735*/;
assign _54702_ = _54703_ | _54705_ /*5732*/;
assign _54711_ = ~D[10] /*5731*/;
assign _54708_ = _54154_ & _54711_ /*5727*/;
assign _54709_ = _54154_ ^ _54711_ /*5730*/;
assign _54710_ = _54702_ & _54709_ /*5728*/;
assign _54603_ = _54702_ ^ _54709_ /*5729*/;
assign _54707_ = _54708_ | _54710_ /*5726*/;
assign _54716_ = ~D[11] /*5725*/;
assign _54713_ = _54155_ & _54716_ /*5721*/;
assign _54714_ = _54155_ ^ _54716_ /*5724*/;
assign _54715_ = _54707_ & _54714_ /*5722*/;
assign _54604_ = _54707_ ^ _54714_ /*5723*/;
assign _54712_ = _54713_ | _54715_ /*5720*/;
assign _54721_ = ~D[12] /*5719*/;
assign _54718_ = _54156_ & _54721_ /*5715*/;
assign _54719_ = _54156_ ^ _54721_ /*5718*/;
assign _54720_ = _54712_ & _54719_ /*5716*/;
assign _54605_ = _54712_ ^ _54719_ /*5717*/;
assign _54717_ = _54718_ | _54720_ /*5714*/;
assign _54726_ = ~D[13] /*5713*/;
assign _54723_ = _54157_ & _54726_ /*5709*/;
assign _54724_ = _54157_ ^ _54726_ /*5712*/;
assign _54725_ = _54717_ & _54724_ /*5710*/;
assign _54606_ = _54717_ ^ _54724_ /*5711*/;
assign _54722_ = _54723_ | _54725_ /*5708*/;
assign _54731_ = ~D[14] /*5707*/;
assign _54728_ = _54158_ & _54731_ /*5703*/;
assign _54729_ = _54158_ ^ _54731_ /*5706*/;
assign _54730_ = _54722_ & _54729_ /*5704*/;
assign _54607_ = _54722_ ^ _54729_ /*5705*/;
assign _54727_ = _54728_ | _54730_ /*5702*/;
assign _54736_ = ~D[15] /*5701*/;
assign _54733_ = _54159_ & _54736_ /*5697*/;
assign _54734_ = _54159_ ^ _54736_ /*5700*/;
assign _54735_ = _54727_ & _54734_ /*5698*/;
assign _54608_ = _54727_ ^ _54734_ /*5699*/;
assign _54732_ = _54733_ | _54735_ /*5696*/;
assign _54741_ = ~D[16] /*5695*/;
assign _54738_ = _54160_ & _54741_ /*5691*/;
assign _54739_ = _54160_ ^ _54741_ /*5694*/;
assign _54740_ = _54732_ & _54739_ /*5692*/;
assign _54609_ = _54732_ ^ _54739_ /*5693*/;
assign _54737_ = _54738_ | _54740_ /*5690*/;
assign _54746_ = ~D[17] /*5689*/;
assign _54743_ = _54161_ & _54746_ /*5685*/;
assign _54744_ = _54161_ ^ _54746_ /*5688*/;
assign _54745_ = _54737_ & _54744_ /*5686*/;
assign _54610_ = _54737_ ^ _54744_ /*5687*/;
assign _54742_ = _54743_ | _54745_ /*5684*/;
assign _54751_ = ~D[18] /*5683*/;
assign _54748_ = _54162_ & _54751_ /*5679*/;
assign _54749_ = _54162_ ^ _54751_ /*5682*/;
assign _54750_ = _54742_ & _54749_ /*5680*/;
assign _54611_ = _54742_ ^ _54749_ /*5681*/;
assign _54747_ = _54748_ | _54750_ /*5678*/;
assign _54756_ = ~D[19] /*5677*/;
assign _54753_ = _54163_ & _54756_ /*5673*/;
assign _54754_ = _54163_ ^ _54756_ /*5676*/;
assign _54755_ = _54747_ & _54754_ /*5674*/;
assign _54612_ = _54747_ ^ _54754_ /*5675*/;
assign _54752_ = _54753_ | _54755_ /*5672*/;
assign _54761_ = ~D[20] /*5671*/;
assign _54758_ = _54164_ & _54761_ /*5667*/;
assign _54759_ = _54164_ ^ _54761_ /*5670*/;
assign _54760_ = _54752_ & _54759_ /*5668*/;
assign _54613_ = _54752_ ^ _54759_ /*5669*/;
assign _54757_ = _54758_ | _54760_ /*5666*/;
assign _54766_ = ~D[21] /*5665*/;
assign _54763_ = _54165_ & _54766_ /*5661*/;
assign _54764_ = _54165_ ^ _54766_ /*5664*/;
assign _54765_ = _54757_ & _54764_ /*5662*/;
assign _54614_ = _54757_ ^ _54764_ /*5663*/;
assign _54762_ = _54763_ | _54765_ /*5660*/;
assign _54771_ = ~D[22] /*5659*/;
assign _54768_ = _54166_ & _54771_ /*5655*/;
assign _54769_ = _54166_ ^ _54771_ /*5658*/;
assign _54770_ = _54762_ & _54769_ /*5656*/;
assign _54615_ = _54762_ ^ _54769_ /*5657*/;
assign _54767_ = _54768_ | _54770_ /*5654*/;
assign _54776_ = ~D[23] /*5653*/;
assign _54773_ = _54167_ & _54776_ /*5649*/;
assign _54774_ = _54167_ ^ _54776_ /*5652*/;
assign _54775_ = _54767_ & _54774_ /*5650*/;
assign _54616_ = _54767_ ^ _54774_ /*5651*/;
assign _54772_ = _54773_ | _54775_ /*5648*/;
assign _54781_ = ~D[24] /*5647*/;
assign _54778_ = _54168_ & _54781_ /*5643*/;
assign _54779_ = _54168_ ^ _54781_ /*5646*/;
assign _54780_ = _54772_ & _54779_ /*5644*/;
assign _54617_ = _54772_ ^ _54779_ /*5645*/;
assign _54777_ = _54778_ | _54780_ /*5642*/;
assign _54786_ = ~D[25] /*5641*/;
assign _54783_ = _54169_ & _54786_ /*5637*/;
assign _54784_ = _54169_ ^ _54786_ /*5640*/;
assign _54785_ = _54777_ & _54784_ /*5638*/;
assign _54618_ = _54777_ ^ _54784_ /*5639*/;
assign _54782_ = _54783_ | _54785_ /*5636*/;
assign _54791_ = ~D[26] /*5635*/;
assign _54788_ = _54170_ & _54791_ /*5631*/;
assign _54789_ = _54170_ ^ _54791_ /*5634*/;
assign _54790_ = _54782_ & _54789_ /*5632*/;
assign _54619_ = _54782_ ^ _54789_ /*5633*/;
assign _54787_ = _54788_ | _54790_ /*5630*/;
assign _54796_ = ~D[27] /*5629*/;
assign _54793_ = _54171_ & _54796_ /*5625*/;
assign _54794_ = _54171_ ^ _54796_ /*5628*/;
assign _54795_ = _54787_ & _54794_ /*5626*/;
assign _54620_ = _54787_ ^ _54794_ /*5627*/;
assign _54792_ = _54793_ | _54795_ /*5624*/;
assign _54801_ = ~D[28] /*5623*/;
assign _54798_ = _54172_ & _54801_ /*5619*/;
assign _54799_ = _54172_ ^ _54801_ /*5622*/;
assign _54800_ = _54792_ & _54799_ /*5620*/;
assign _54621_ = _54792_ ^ _54799_ /*5621*/;
assign _54797_ = _54798_ | _54800_ /*5618*/;
assign _54806_ = ~D[29] /*5617*/;
assign _54803_ = _54173_ & _54806_ /*5613*/;
assign _54804_ = _54173_ ^ _54806_ /*5616*/;
assign _54805_ = _54797_ & _54804_ /*5614*/;
assign _54622_ = _54797_ ^ _54804_ /*5615*/;
assign _54802_ = _54803_ | _54805_ /*5612*/;
assign _54811_ = ~D[30] /*5611*/;
assign _54808_ = _54174_ & _54811_ /*5607*/;
assign _54809_ = _54174_ ^ _54811_ /*5610*/;
assign _54810_ = _54802_ & _54809_ /*5608*/;
assign _54623_ = _54802_ ^ _54809_ /*5609*/;
assign _54807_ = _54808_ | _54810_ /*5606*/;
assign _54816_ = ~D[31] /*5605*/;
assign _54813_ = _54175_ & _54816_ /*5601*/;
assign _54814_ = _54175_ ^ _54816_ /*5604*/;
assign _54815_ = _54807_ & _54814_ /*5602*/;
assign _54624_ = _54807_ ^ _54814_ /*5603*/;
assign _54812_ = _54813_ | _54815_ /*5600*/;
assign _54821_ = ~D[32] /*5599*/;
assign _54818_ = _54176_ & _54821_ /*5595*/;
assign _54819_ = _54176_ ^ _54821_ /*5598*/;
assign _54820_ = _54812_ & _54819_ /*5596*/;
assign _54625_ = _54812_ ^ _54819_ /*5597*/;
assign _54817_ = _54818_ | _54820_ /*5594*/;
assign _54826_ = ~D[33] /*5593*/;
assign _54823_ = _54177_ & _54826_ /*5589*/;
assign _54824_ = _54177_ ^ _54826_ /*5592*/;
assign _54825_ = _54817_ & _54824_ /*5590*/;
assign _54626_ = _54817_ ^ _54824_ /*5591*/;
assign _54822_ = _54823_ | _54825_ /*5588*/;
assign _54831_ = ~D[34] /*5587*/;
assign _54828_ = _54178_ & _54831_ /*5583*/;
assign _54829_ = _54178_ ^ _54831_ /*5586*/;
assign _54830_ = _54822_ & _54829_ /*5584*/;
assign _54627_ = _54822_ ^ _54829_ /*5585*/;
assign _54827_ = _54828_ | _54830_ /*5582*/;
assign _54836_ = ~D[35] /*5581*/;
assign _54833_ = _54179_ & _54836_ /*5577*/;
assign _54834_ = _54179_ ^ _54836_ /*5580*/;
assign _54835_ = _54827_ & _54834_ /*5578*/;
assign _54628_ = _54827_ ^ _54834_ /*5579*/;
assign _54832_ = _54833_ | _54835_ /*5576*/;
assign _54841_ = ~D[36] /*5575*/;
assign _54838_ = _54180_ & _54841_ /*5571*/;
assign _54839_ = _54180_ ^ _54841_ /*5574*/;
assign _54840_ = _54832_ & _54839_ /*5572*/;
assign _54629_ = _54832_ ^ _54839_ /*5573*/;
assign _54837_ = _54838_ | _54840_ /*5570*/;
assign _54846_ = ~D[37] /*5569*/;
assign _54843_ = _54181_ & _54846_ /*5565*/;
assign _54844_ = _54181_ ^ _54846_ /*5568*/;
assign _54845_ = _54837_ & _54844_ /*5566*/;
assign _54630_ = _54837_ ^ _54844_ /*5567*/;
assign _54842_ = _54843_ | _54845_ /*5564*/;
assign _54851_ = ~D[38] /*5563*/;
assign _54848_ = _54182_ & _54851_ /*5559*/;
assign _54849_ = _54182_ ^ _54851_ /*5562*/;
assign _54850_ = _54842_ & _54849_ /*5560*/;
assign _54631_ = _54842_ ^ _54849_ /*5561*/;
assign _54847_ = _54848_ | _54850_ /*5558*/;
assign _54856_ = ~D[39] /*5557*/;
assign _54853_ = _54183_ & _54856_ /*5553*/;
assign _54854_ = _54183_ ^ _54856_ /*5556*/;
assign _54855_ = _54847_ & _54854_ /*5554*/;
assign _54632_ = _54847_ ^ _54854_ /*5555*/;
assign _54852_ = _54853_ | _54855_ /*5552*/;
assign _54861_ = ~D[40] /*5551*/;
assign _54858_ = _54184_ & _54861_ /*5547*/;
assign _54859_ = _54184_ ^ _54861_ /*5550*/;
assign _54860_ = _54852_ & _54859_ /*5548*/;
assign _54633_ = _54852_ ^ _54859_ /*5549*/;
assign _54857_ = _54858_ | _54860_ /*5546*/;
assign _54866_ = ~D[41] /*5545*/;
assign _54863_ = _54185_ & _54866_ /*5541*/;
assign _54864_ = _54185_ ^ _54866_ /*5544*/;
assign _54865_ = _54857_ & _54864_ /*5542*/;
assign _54634_ = _54857_ ^ _54864_ /*5543*/;
assign _54862_ = _54863_ | _54865_ /*5540*/;
assign _54871_ = ~D[42] /*5539*/;
assign _54868_ = _54186_ & _54871_ /*5535*/;
assign _54869_ = _54186_ ^ _54871_ /*5538*/;
assign _54870_ = _54862_ & _54869_ /*5536*/;
assign _54635_ = _54862_ ^ _54869_ /*5537*/;
assign _54867_ = _54868_ | _54870_ /*5534*/;
assign _54876_ = ~D[43] /*5533*/;
assign _54873_ = _54187_ & _54876_ /*5529*/;
assign _54874_ = _54187_ ^ _54876_ /*5532*/;
assign _54875_ = _54867_ & _54874_ /*5530*/;
assign _54636_ = _54867_ ^ _54874_ /*5531*/;
assign _54872_ = _54873_ | _54875_ /*5528*/;
assign _54881_ = ~D[44] /*5527*/;
assign _54878_ = _54188_ & _54881_ /*5523*/;
assign _54879_ = _54188_ ^ _54881_ /*5526*/;
assign _54880_ = _54872_ & _54879_ /*5524*/;
assign _54637_ = _54872_ ^ _54879_ /*5525*/;
assign _54877_ = _54878_ | _54880_ /*5522*/;
assign _54886_ = ~D[45] /*5521*/;
assign _54883_ = _54189_ & _54886_ /*5517*/;
assign _54884_ = _54189_ ^ _54886_ /*5520*/;
assign _54885_ = _54877_ & _54884_ /*5518*/;
assign _54638_ = _54877_ ^ _54884_ /*5519*/;
assign _54882_ = _54883_ | _54885_ /*5516*/;
assign _54891_ = ~D[46] /*5515*/;
assign _54888_ = _54190_ & _54891_ /*5511*/;
assign _54889_ = _54190_ ^ _54891_ /*5514*/;
assign _54890_ = _54882_ & _54889_ /*5512*/;
assign _54639_ = _54882_ ^ _54889_ /*5513*/;
assign _54887_ = _54888_ | _54890_ /*5510*/;
assign _54896_ = ~D[47] /*5509*/;
assign _54893_ = _54191_ & _54896_ /*5505*/;
assign _54894_ = _54191_ ^ _54896_ /*5508*/;
assign _54895_ = _54887_ & _54894_ /*5506*/;
assign _54640_ = _54887_ ^ _54894_ /*5507*/;
assign _54892_ = _54893_ | _54895_ /*5504*/;
assign _54901_ = ~D[48] /*5503*/;
assign _54898_ = _54192_ & _54901_ /*5499*/;
assign _54899_ = _54192_ ^ _54901_ /*5502*/;
assign _54900_ = _54892_ & _54899_ /*5500*/;
assign _54641_ = _54892_ ^ _54899_ /*5501*/;
assign _54897_ = _54898_ | _54900_ /*5498*/;
assign _54906_ = ~D[49] /*5497*/;
assign _54903_ = _54193_ & _54906_ /*5493*/;
assign _54904_ = _54193_ ^ _54906_ /*5496*/;
assign _54905_ = _54897_ & _54904_ /*5494*/;
assign _54642_ = _54897_ ^ _54904_ /*5495*/;
assign _54902_ = _54903_ | _54905_ /*5492*/;
assign _54911_ = ~D[50] /*5491*/;
assign _54908_ = _54194_ & _54911_ /*5487*/;
assign _54909_ = _54194_ ^ _54911_ /*5490*/;
assign _54910_ = _54902_ & _54909_ /*5488*/;
assign _54643_ = _54902_ ^ _54909_ /*5489*/;
assign _54907_ = _54908_ | _54910_ /*5486*/;
assign _54916_ = ~D[51] /*5485*/;
assign _54913_ = _54195_ & _54916_ /*5481*/;
assign _54914_ = _54195_ ^ _54916_ /*5484*/;
assign _54915_ = _54907_ & _54914_ /*5482*/;
assign _54644_ = _54907_ ^ _54914_ /*5483*/;
assign _54912_ = _54913_ | _54915_ /*5480*/;
assign _54921_ = ~D[52] /*5479*/;
assign _54918_ = _54196_ & _54921_ /*5475*/;
assign _54919_ = _54196_ ^ _54921_ /*5478*/;
assign _54920_ = _54912_ & _54919_ /*5476*/;
assign _54645_ = _54912_ ^ _54919_ /*5477*/;
assign _54917_ = _54918_ | _54920_ /*5474*/;
assign _54926_ = ~D[53] /*5473*/;
assign _54923_ = _54197_ & _54926_ /*5469*/;
assign _54924_ = _54197_ ^ _54926_ /*5472*/;
assign _54925_ = _54917_ & _54924_ /*5470*/;
assign _54646_ = _54917_ ^ _54924_ /*5471*/;
assign _54922_ = _54923_ | _54925_ /*5468*/;
assign _54931_ = ~D[54] /*5467*/;
assign _54928_ = _54198_ & _54931_ /*5463*/;
assign _54929_ = _54198_ ^ _54931_ /*5466*/;
assign _54930_ = _54922_ & _54929_ /*5464*/;
assign _54647_ = _54922_ ^ _54929_ /*5465*/;
assign _54927_ = _54928_ | _54930_ /*5462*/;
assign _54936_ = ~D[55] /*5461*/;
assign _54933_ = _54199_ & _54936_ /*5457*/;
assign _54934_ = _54199_ ^ _54936_ /*5460*/;
assign _54935_ = _54927_ & _54934_ /*5458*/;
assign _54648_ = _54927_ ^ _54934_ /*5459*/;
assign _54932_ = _54933_ | _54935_ /*5456*/;
assign _54941_ = ~D[56] /*5455*/;
assign _54938_ = _54200_ & _54941_ /*5451*/;
assign _54939_ = _54200_ ^ _54941_ /*5454*/;
assign _54940_ = _54932_ & _54939_ /*5452*/;
assign _54649_ = _54932_ ^ _54939_ /*5453*/;
assign _54937_ = _54938_ | _54940_ /*5450*/;
assign _54946_ = ~D[57] /*5449*/;
assign _54943_ = _54201_ & _54946_ /*5445*/;
assign _54944_ = _54201_ ^ _54946_ /*5448*/;
assign _54945_ = _54937_ & _54944_ /*5446*/;
assign _54650_ = _54937_ ^ _54944_ /*5447*/;
assign _54942_ = _54943_ | _54945_ /*5444*/;
assign _54951_ = ~D[58] /*5443*/;
assign _54948_ = _54202_ & _54951_ /*5439*/;
assign _54949_ = _54202_ ^ _54951_ /*5442*/;
assign _54950_ = _54942_ & _54949_ /*5440*/;
assign _54651_ = _54942_ ^ _54949_ /*5441*/;
assign _54947_ = _54948_ | _54950_ /*5438*/;
assign _54956_ = ~D[59] /*5437*/;
assign _54953_ = _54203_ & _54956_ /*5433*/;
assign _54954_ = _54203_ ^ _54956_ /*5436*/;
assign _54955_ = _54947_ & _54954_ /*5434*/;
assign _54652_ = _54947_ ^ _54954_ /*5435*/;
assign _54952_ = _54953_ | _54955_ /*5432*/;
assign _54961_ = ~D[60] /*5431*/;
assign _54958_ = _54204_ & _54961_ /*5427*/;
assign _54959_ = _54204_ ^ _54961_ /*5430*/;
assign _54960_ = _54952_ & _54959_ /*5428*/;
assign _54653_ = _54952_ ^ _54959_ /*5429*/;
assign _54957_ = _54958_ | _54960_ /*5426*/;
assign _54966_ = ~D[61] /*5425*/;
assign _54963_ = _54205_ & _54966_ /*5421*/;
assign _54964_ = _54205_ ^ _54966_ /*5424*/;
assign _54965_ = _54957_ & _54964_ /*5422*/;
assign _54654_ = _54957_ ^ _54964_ /*5423*/;
assign _54962_ = _54963_ | _54965_ /*5420*/;
assign _54971_ = ~D[62] /*5419*/;
assign _54968_ = _54206_ & _54971_ /*5415*/;
assign _54969_ = _54206_ ^ _54971_ /*5418*/;
assign _54970_ = _54962_ & _54969_ /*5416*/;
assign _54655_ = _54962_ ^ _54969_ /*5417*/;
assign _54967_ = _54968_ | _54970_ /*5414*/;
assign _54972_ = _54207_ & oneWire /*5409*/;
assign _54973_ = _54207_ ^ oneWire /*5412*/;
assign _54974_ = _54967_ & _54973_ /*5410*/;
assign _54656_ = _54967_ ^ _54973_ /*5411*/;
assign Q[2] = _54972_ | _54974_ /*5408*/;
assign _55107_ = ~Q[2] /*5023*/;
assign _55106_ = _55107_ & D[0] /*5022*/;
assign _55109_ = _54593_ & _55106_ /*5017*/;
assign _55110_ = _54593_ ^ _55106_ /*5020*/;
assign _55111_ = zeroWire & _55110_ /*5018*/;
assign _55041_ = zeroWire ^ _55110_ /*5019*/;
assign _55108_ = _55109_ | _55111_ /*5016*/;
assign _55113_ = ~Q[2] /*5015*/;
assign _55112_ = _55113_ & D[1] /*5014*/;
assign _55115_ = _54594_ & _55112_ /*5009*/;
assign _55116_ = _54594_ ^ _55112_ /*5012*/;
assign _55117_ = _55108_ & _55116_ /*5010*/;
assign _55042_ = _55108_ ^ _55116_ /*5011*/;
assign _55114_ = _55115_ | _55117_ /*5008*/;
assign _55119_ = ~Q[2] /*5007*/;
assign _55118_ = _55119_ & D[2] /*5006*/;
assign _55121_ = _54595_ & _55118_ /*5001*/;
assign _55122_ = _54595_ ^ _55118_ /*5004*/;
assign _55123_ = _55114_ & _55122_ /*5002*/;
assign _55043_ = _55114_ ^ _55122_ /*5003*/;
assign _55120_ = _55121_ | _55123_ /*5000*/;
assign _55125_ = ~Q[2] /*4999*/;
assign _55124_ = _55125_ & D[3] /*4998*/;
assign _55127_ = _54596_ & _55124_ /*4993*/;
assign _55128_ = _54596_ ^ _55124_ /*4996*/;
assign _55129_ = _55120_ & _55128_ /*4994*/;
assign _55044_ = _55120_ ^ _55128_ /*4995*/;
assign _55126_ = _55127_ | _55129_ /*4992*/;
assign _55131_ = ~Q[2] /*4991*/;
assign _55130_ = _55131_ & D[4] /*4990*/;
assign _55133_ = _54597_ & _55130_ /*4985*/;
assign _55134_ = _54597_ ^ _55130_ /*4988*/;
assign _55135_ = _55126_ & _55134_ /*4986*/;
assign _55045_ = _55126_ ^ _55134_ /*4987*/;
assign _55132_ = _55133_ | _55135_ /*4984*/;
assign _55137_ = ~Q[2] /*4983*/;
assign _55136_ = _55137_ & D[5] /*4982*/;
assign _55139_ = _54598_ & _55136_ /*4977*/;
assign _55140_ = _54598_ ^ _55136_ /*4980*/;
assign _55141_ = _55132_ & _55140_ /*4978*/;
assign _55046_ = _55132_ ^ _55140_ /*4979*/;
assign _55138_ = _55139_ | _55141_ /*4976*/;
assign _55143_ = ~Q[2] /*4975*/;
assign _55142_ = _55143_ & D[6] /*4974*/;
assign _55145_ = _54599_ & _55142_ /*4969*/;
assign _55146_ = _54599_ ^ _55142_ /*4972*/;
assign _55147_ = _55138_ & _55146_ /*4970*/;
assign _55047_ = _55138_ ^ _55146_ /*4971*/;
assign _55144_ = _55145_ | _55147_ /*4968*/;
assign _55149_ = ~Q[2] /*4967*/;
assign _55148_ = _55149_ & D[7] /*4966*/;
assign _55151_ = _54600_ & _55148_ /*4961*/;
assign _55152_ = _54600_ ^ _55148_ /*4964*/;
assign _55153_ = _55144_ & _55152_ /*4962*/;
assign _55048_ = _55144_ ^ _55152_ /*4963*/;
assign _55150_ = _55151_ | _55153_ /*4960*/;
assign _55155_ = ~Q[2] /*4959*/;
assign _55154_ = _55155_ & D[8] /*4958*/;
assign _55157_ = _54601_ & _55154_ /*4953*/;
assign _55158_ = _54601_ ^ _55154_ /*4956*/;
assign _55159_ = _55150_ & _55158_ /*4954*/;
assign _55049_ = _55150_ ^ _55158_ /*4955*/;
assign _55156_ = _55157_ | _55159_ /*4952*/;
assign _55161_ = ~Q[2] /*4951*/;
assign _55160_ = _55161_ & D[9] /*4950*/;
assign _55163_ = _54602_ & _55160_ /*4945*/;
assign _55164_ = _54602_ ^ _55160_ /*4948*/;
assign _55165_ = _55156_ & _55164_ /*4946*/;
assign _55050_ = _55156_ ^ _55164_ /*4947*/;
assign _55162_ = _55163_ | _55165_ /*4944*/;
assign _55167_ = ~Q[2] /*4943*/;
assign _55166_ = _55167_ & D[10] /*4942*/;
assign _55169_ = _54603_ & _55166_ /*4937*/;
assign _55170_ = _54603_ ^ _55166_ /*4940*/;
assign _55171_ = _55162_ & _55170_ /*4938*/;
assign _55051_ = _55162_ ^ _55170_ /*4939*/;
assign _55168_ = _55169_ | _55171_ /*4936*/;
assign _55173_ = ~Q[2] /*4935*/;
assign _55172_ = _55173_ & D[11] /*4934*/;
assign _55175_ = _54604_ & _55172_ /*4929*/;
assign _55176_ = _54604_ ^ _55172_ /*4932*/;
assign _55177_ = _55168_ & _55176_ /*4930*/;
assign _55052_ = _55168_ ^ _55176_ /*4931*/;
assign _55174_ = _55175_ | _55177_ /*4928*/;
assign _55179_ = ~Q[2] /*4927*/;
assign _55178_ = _55179_ & D[12] /*4926*/;
assign _55181_ = _54605_ & _55178_ /*4921*/;
assign _55182_ = _54605_ ^ _55178_ /*4924*/;
assign _55183_ = _55174_ & _55182_ /*4922*/;
assign _55053_ = _55174_ ^ _55182_ /*4923*/;
assign _55180_ = _55181_ | _55183_ /*4920*/;
assign _55185_ = ~Q[2] /*4919*/;
assign _55184_ = _55185_ & D[13] /*4918*/;
assign _55187_ = _54606_ & _55184_ /*4913*/;
assign _55188_ = _54606_ ^ _55184_ /*4916*/;
assign _55189_ = _55180_ & _55188_ /*4914*/;
assign _55054_ = _55180_ ^ _55188_ /*4915*/;
assign _55186_ = _55187_ | _55189_ /*4912*/;
assign _55191_ = ~Q[2] /*4911*/;
assign _55190_ = _55191_ & D[14] /*4910*/;
assign _55193_ = _54607_ & _55190_ /*4905*/;
assign _55194_ = _54607_ ^ _55190_ /*4908*/;
assign _55195_ = _55186_ & _55194_ /*4906*/;
assign _55055_ = _55186_ ^ _55194_ /*4907*/;
assign _55192_ = _55193_ | _55195_ /*4904*/;
assign _55197_ = ~Q[2] /*4903*/;
assign _55196_ = _55197_ & D[15] /*4902*/;
assign _55199_ = _54608_ & _55196_ /*4897*/;
assign _55200_ = _54608_ ^ _55196_ /*4900*/;
assign _55201_ = _55192_ & _55200_ /*4898*/;
assign _55056_ = _55192_ ^ _55200_ /*4899*/;
assign _55198_ = _55199_ | _55201_ /*4896*/;
assign _55203_ = ~Q[2] /*4895*/;
assign _55202_ = _55203_ & D[16] /*4894*/;
assign _55205_ = _54609_ & _55202_ /*4889*/;
assign _55206_ = _54609_ ^ _55202_ /*4892*/;
assign _55207_ = _55198_ & _55206_ /*4890*/;
assign _55057_ = _55198_ ^ _55206_ /*4891*/;
assign _55204_ = _55205_ | _55207_ /*4888*/;
assign _55209_ = ~Q[2] /*4887*/;
assign _55208_ = _55209_ & D[17] /*4886*/;
assign _55211_ = _54610_ & _55208_ /*4881*/;
assign _55212_ = _54610_ ^ _55208_ /*4884*/;
assign _55213_ = _55204_ & _55212_ /*4882*/;
assign _55058_ = _55204_ ^ _55212_ /*4883*/;
assign _55210_ = _55211_ | _55213_ /*4880*/;
assign _55215_ = ~Q[2] /*4879*/;
assign _55214_ = _55215_ & D[18] /*4878*/;
assign _55217_ = _54611_ & _55214_ /*4873*/;
assign _55218_ = _54611_ ^ _55214_ /*4876*/;
assign _55219_ = _55210_ & _55218_ /*4874*/;
assign _55059_ = _55210_ ^ _55218_ /*4875*/;
assign _55216_ = _55217_ | _55219_ /*4872*/;
assign _55221_ = ~Q[2] /*4871*/;
assign _55220_ = _55221_ & D[19] /*4870*/;
assign _55223_ = _54612_ & _55220_ /*4865*/;
assign _55224_ = _54612_ ^ _55220_ /*4868*/;
assign _55225_ = _55216_ & _55224_ /*4866*/;
assign _55060_ = _55216_ ^ _55224_ /*4867*/;
assign _55222_ = _55223_ | _55225_ /*4864*/;
assign _55227_ = ~Q[2] /*4863*/;
assign _55226_ = _55227_ & D[20] /*4862*/;
assign _55229_ = _54613_ & _55226_ /*4857*/;
assign _55230_ = _54613_ ^ _55226_ /*4860*/;
assign _55231_ = _55222_ & _55230_ /*4858*/;
assign _55061_ = _55222_ ^ _55230_ /*4859*/;
assign _55228_ = _55229_ | _55231_ /*4856*/;
assign _55233_ = ~Q[2] /*4855*/;
assign _55232_ = _55233_ & D[21] /*4854*/;
assign _55235_ = _54614_ & _55232_ /*4849*/;
assign _55236_ = _54614_ ^ _55232_ /*4852*/;
assign _55237_ = _55228_ & _55236_ /*4850*/;
assign _55062_ = _55228_ ^ _55236_ /*4851*/;
assign _55234_ = _55235_ | _55237_ /*4848*/;
assign _55239_ = ~Q[2] /*4847*/;
assign _55238_ = _55239_ & D[22] /*4846*/;
assign _55241_ = _54615_ & _55238_ /*4841*/;
assign _55242_ = _54615_ ^ _55238_ /*4844*/;
assign _55243_ = _55234_ & _55242_ /*4842*/;
assign _55063_ = _55234_ ^ _55242_ /*4843*/;
assign _55240_ = _55241_ | _55243_ /*4840*/;
assign _55245_ = ~Q[2] /*4839*/;
assign _55244_ = _55245_ & D[23] /*4838*/;
assign _55247_ = _54616_ & _55244_ /*4833*/;
assign _55248_ = _54616_ ^ _55244_ /*4836*/;
assign _55249_ = _55240_ & _55248_ /*4834*/;
assign _55064_ = _55240_ ^ _55248_ /*4835*/;
assign _55246_ = _55247_ | _55249_ /*4832*/;
assign _55251_ = ~Q[2] /*4831*/;
assign _55250_ = _55251_ & D[24] /*4830*/;
assign _55253_ = _54617_ & _55250_ /*4825*/;
assign _55254_ = _54617_ ^ _55250_ /*4828*/;
assign _55255_ = _55246_ & _55254_ /*4826*/;
assign _55065_ = _55246_ ^ _55254_ /*4827*/;
assign _55252_ = _55253_ | _55255_ /*4824*/;
assign _55257_ = ~Q[2] /*4823*/;
assign _55256_ = _55257_ & D[25] /*4822*/;
assign _55259_ = _54618_ & _55256_ /*4817*/;
assign _55260_ = _54618_ ^ _55256_ /*4820*/;
assign _55261_ = _55252_ & _55260_ /*4818*/;
assign _55066_ = _55252_ ^ _55260_ /*4819*/;
assign _55258_ = _55259_ | _55261_ /*4816*/;
assign _55263_ = ~Q[2] /*4815*/;
assign _55262_ = _55263_ & D[26] /*4814*/;
assign _55265_ = _54619_ & _55262_ /*4809*/;
assign _55266_ = _54619_ ^ _55262_ /*4812*/;
assign _55267_ = _55258_ & _55266_ /*4810*/;
assign _55067_ = _55258_ ^ _55266_ /*4811*/;
assign _55264_ = _55265_ | _55267_ /*4808*/;
assign _55269_ = ~Q[2] /*4807*/;
assign _55268_ = _55269_ & D[27] /*4806*/;
assign _55271_ = _54620_ & _55268_ /*4801*/;
assign _55272_ = _54620_ ^ _55268_ /*4804*/;
assign _55273_ = _55264_ & _55272_ /*4802*/;
assign _55068_ = _55264_ ^ _55272_ /*4803*/;
assign _55270_ = _55271_ | _55273_ /*4800*/;
assign _55275_ = ~Q[2] /*4799*/;
assign _55274_ = _55275_ & D[28] /*4798*/;
assign _55277_ = _54621_ & _55274_ /*4793*/;
assign _55278_ = _54621_ ^ _55274_ /*4796*/;
assign _55279_ = _55270_ & _55278_ /*4794*/;
assign _55069_ = _55270_ ^ _55278_ /*4795*/;
assign _55276_ = _55277_ | _55279_ /*4792*/;
assign _55281_ = ~Q[2] /*4791*/;
assign _55280_ = _55281_ & D[29] /*4790*/;
assign _55283_ = _54622_ & _55280_ /*4785*/;
assign _55284_ = _54622_ ^ _55280_ /*4788*/;
assign _55285_ = _55276_ & _55284_ /*4786*/;
assign _55070_ = _55276_ ^ _55284_ /*4787*/;
assign _55282_ = _55283_ | _55285_ /*4784*/;
assign _55287_ = ~Q[2] /*4783*/;
assign _55286_ = _55287_ & D[30] /*4782*/;
assign _55289_ = _54623_ & _55286_ /*4777*/;
assign _55290_ = _54623_ ^ _55286_ /*4780*/;
assign _55291_ = _55282_ & _55290_ /*4778*/;
assign _55071_ = _55282_ ^ _55290_ /*4779*/;
assign _55288_ = _55289_ | _55291_ /*4776*/;
assign _55293_ = ~Q[2] /*4775*/;
assign _55292_ = _55293_ & D[31] /*4774*/;
assign _55295_ = _54624_ & _55292_ /*4769*/;
assign _55296_ = _54624_ ^ _55292_ /*4772*/;
assign _55297_ = _55288_ & _55296_ /*4770*/;
assign _55072_ = _55288_ ^ _55296_ /*4771*/;
assign _55294_ = _55295_ | _55297_ /*4768*/;
assign _55299_ = ~Q[2] /*4767*/;
assign _55298_ = _55299_ & D[32] /*4766*/;
assign _55301_ = _54625_ & _55298_ /*4761*/;
assign _55302_ = _54625_ ^ _55298_ /*4764*/;
assign _55303_ = _55294_ & _55302_ /*4762*/;
assign _55073_ = _55294_ ^ _55302_ /*4763*/;
assign _55300_ = _55301_ | _55303_ /*4760*/;
assign _55305_ = ~Q[2] /*4759*/;
assign _55304_ = _55305_ & D[33] /*4758*/;
assign _55307_ = _54626_ & _55304_ /*4753*/;
assign _55308_ = _54626_ ^ _55304_ /*4756*/;
assign _55309_ = _55300_ & _55308_ /*4754*/;
assign _55074_ = _55300_ ^ _55308_ /*4755*/;
assign _55306_ = _55307_ | _55309_ /*4752*/;
assign _55311_ = ~Q[2] /*4751*/;
assign _55310_ = _55311_ & D[34] /*4750*/;
assign _55313_ = _54627_ & _55310_ /*4745*/;
assign _55314_ = _54627_ ^ _55310_ /*4748*/;
assign _55315_ = _55306_ & _55314_ /*4746*/;
assign _55075_ = _55306_ ^ _55314_ /*4747*/;
assign _55312_ = _55313_ | _55315_ /*4744*/;
assign _55317_ = ~Q[2] /*4743*/;
assign _55316_ = _55317_ & D[35] /*4742*/;
assign _55319_ = _54628_ & _55316_ /*4737*/;
assign _55320_ = _54628_ ^ _55316_ /*4740*/;
assign _55321_ = _55312_ & _55320_ /*4738*/;
assign _55076_ = _55312_ ^ _55320_ /*4739*/;
assign _55318_ = _55319_ | _55321_ /*4736*/;
assign _55323_ = ~Q[2] /*4735*/;
assign _55322_ = _55323_ & D[36] /*4734*/;
assign _55325_ = _54629_ & _55322_ /*4729*/;
assign _55326_ = _54629_ ^ _55322_ /*4732*/;
assign _55327_ = _55318_ & _55326_ /*4730*/;
assign _55077_ = _55318_ ^ _55326_ /*4731*/;
assign _55324_ = _55325_ | _55327_ /*4728*/;
assign _55329_ = ~Q[2] /*4727*/;
assign _55328_ = _55329_ & D[37] /*4726*/;
assign _55331_ = _54630_ & _55328_ /*4721*/;
assign _55332_ = _54630_ ^ _55328_ /*4724*/;
assign _55333_ = _55324_ & _55332_ /*4722*/;
assign _55078_ = _55324_ ^ _55332_ /*4723*/;
assign _55330_ = _55331_ | _55333_ /*4720*/;
assign _55335_ = ~Q[2] /*4719*/;
assign _55334_ = _55335_ & D[38] /*4718*/;
assign _55337_ = _54631_ & _55334_ /*4713*/;
assign _55338_ = _54631_ ^ _55334_ /*4716*/;
assign _55339_ = _55330_ & _55338_ /*4714*/;
assign _55079_ = _55330_ ^ _55338_ /*4715*/;
assign _55336_ = _55337_ | _55339_ /*4712*/;
assign _55341_ = ~Q[2] /*4711*/;
assign _55340_ = _55341_ & D[39] /*4710*/;
assign _55343_ = _54632_ & _55340_ /*4705*/;
assign _55344_ = _54632_ ^ _55340_ /*4708*/;
assign _55345_ = _55336_ & _55344_ /*4706*/;
assign _55080_ = _55336_ ^ _55344_ /*4707*/;
assign _55342_ = _55343_ | _55345_ /*4704*/;
assign _55347_ = ~Q[2] /*4703*/;
assign _55346_ = _55347_ & D[40] /*4702*/;
assign _55349_ = _54633_ & _55346_ /*4697*/;
assign _55350_ = _54633_ ^ _55346_ /*4700*/;
assign _55351_ = _55342_ & _55350_ /*4698*/;
assign _55081_ = _55342_ ^ _55350_ /*4699*/;
assign _55348_ = _55349_ | _55351_ /*4696*/;
assign _55353_ = ~Q[2] /*4695*/;
assign _55352_ = _55353_ & D[41] /*4694*/;
assign _55355_ = _54634_ & _55352_ /*4689*/;
assign _55356_ = _54634_ ^ _55352_ /*4692*/;
assign _55357_ = _55348_ & _55356_ /*4690*/;
assign _55082_ = _55348_ ^ _55356_ /*4691*/;
assign _55354_ = _55355_ | _55357_ /*4688*/;
assign _55359_ = ~Q[2] /*4687*/;
assign _55358_ = _55359_ & D[42] /*4686*/;
assign _55361_ = _54635_ & _55358_ /*4681*/;
assign _55362_ = _54635_ ^ _55358_ /*4684*/;
assign _55363_ = _55354_ & _55362_ /*4682*/;
assign _55083_ = _55354_ ^ _55362_ /*4683*/;
assign _55360_ = _55361_ | _55363_ /*4680*/;
assign _55365_ = ~Q[2] /*4679*/;
assign _55364_ = _55365_ & D[43] /*4678*/;
assign _55367_ = _54636_ & _55364_ /*4673*/;
assign _55368_ = _54636_ ^ _55364_ /*4676*/;
assign _55369_ = _55360_ & _55368_ /*4674*/;
assign _55084_ = _55360_ ^ _55368_ /*4675*/;
assign _55366_ = _55367_ | _55369_ /*4672*/;
assign _55371_ = ~Q[2] /*4671*/;
assign _55370_ = _55371_ & D[44] /*4670*/;
assign _55373_ = _54637_ & _55370_ /*4665*/;
assign _55374_ = _54637_ ^ _55370_ /*4668*/;
assign _55375_ = _55366_ & _55374_ /*4666*/;
assign _55085_ = _55366_ ^ _55374_ /*4667*/;
assign _55372_ = _55373_ | _55375_ /*4664*/;
assign _55377_ = ~Q[2] /*4663*/;
assign _55376_ = _55377_ & D[45] /*4662*/;
assign _55379_ = _54638_ & _55376_ /*4657*/;
assign _55380_ = _54638_ ^ _55376_ /*4660*/;
assign _55381_ = _55372_ & _55380_ /*4658*/;
assign _55086_ = _55372_ ^ _55380_ /*4659*/;
assign _55378_ = _55379_ | _55381_ /*4656*/;
assign _55383_ = ~Q[2] /*4655*/;
assign _55382_ = _55383_ & D[46] /*4654*/;
assign _55385_ = _54639_ & _55382_ /*4649*/;
assign _55386_ = _54639_ ^ _55382_ /*4652*/;
assign _55387_ = _55378_ & _55386_ /*4650*/;
assign _55087_ = _55378_ ^ _55386_ /*4651*/;
assign _55384_ = _55385_ | _55387_ /*4648*/;
assign _55389_ = ~Q[2] /*4647*/;
assign _55388_ = _55389_ & D[47] /*4646*/;
assign _55391_ = _54640_ & _55388_ /*4641*/;
assign _55392_ = _54640_ ^ _55388_ /*4644*/;
assign _55393_ = _55384_ & _55392_ /*4642*/;
assign _55088_ = _55384_ ^ _55392_ /*4643*/;
assign _55390_ = _55391_ | _55393_ /*4640*/;
assign _55395_ = ~Q[2] /*4639*/;
assign _55394_ = _55395_ & D[48] /*4638*/;
assign _55397_ = _54641_ & _55394_ /*4633*/;
assign _55398_ = _54641_ ^ _55394_ /*4636*/;
assign _55399_ = _55390_ & _55398_ /*4634*/;
assign _55089_ = _55390_ ^ _55398_ /*4635*/;
assign _55396_ = _55397_ | _55399_ /*4632*/;
assign _55401_ = ~Q[2] /*4631*/;
assign _55400_ = _55401_ & D[49] /*4630*/;
assign _55403_ = _54642_ & _55400_ /*4625*/;
assign _55404_ = _54642_ ^ _55400_ /*4628*/;
assign _55405_ = _55396_ & _55404_ /*4626*/;
assign _55090_ = _55396_ ^ _55404_ /*4627*/;
assign _55402_ = _55403_ | _55405_ /*4624*/;
assign _55407_ = ~Q[2] /*4623*/;
assign _55406_ = _55407_ & D[50] /*4622*/;
assign _55409_ = _54643_ & _55406_ /*4617*/;
assign _55410_ = _54643_ ^ _55406_ /*4620*/;
assign _55411_ = _55402_ & _55410_ /*4618*/;
assign _55091_ = _55402_ ^ _55410_ /*4619*/;
assign _55408_ = _55409_ | _55411_ /*4616*/;
assign _55413_ = ~Q[2] /*4615*/;
assign _55412_ = _55413_ & D[51] /*4614*/;
assign _55415_ = _54644_ & _55412_ /*4609*/;
assign _55416_ = _54644_ ^ _55412_ /*4612*/;
assign _55417_ = _55408_ & _55416_ /*4610*/;
assign _55092_ = _55408_ ^ _55416_ /*4611*/;
assign _55414_ = _55415_ | _55417_ /*4608*/;
assign _55419_ = ~Q[2] /*4607*/;
assign _55418_ = _55419_ & D[52] /*4606*/;
assign _55421_ = _54645_ & _55418_ /*4601*/;
assign _55422_ = _54645_ ^ _55418_ /*4604*/;
assign _55423_ = _55414_ & _55422_ /*4602*/;
assign _55093_ = _55414_ ^ _55422_ /*4603*/;
assign _55420_ = _55421_ | _55423_ /*4600*/;
assign _55425_ = ~Q[2] /*4599*/;
assign _55424_ = _55425_ & D[53] /*4598*/;
assign _55427_ = _54646_ & _55424_ /*4593*/;
assign _55428_ = _54646_ ^ _55424_ /*4596*/;
assign _55429_ = _55420_ & _55428_ /*4594*/;
assign _55094_ = _55420_ ^ _55428_ /*4595*/;
assign _55426_ = _55427_ | _55429_ /*4592*/;
assign _55431_ = ~Q[2] /*4591*/;
assign _55430_ = _55431_ & D[54] /*4590*/;
assign _55433_ = _54647_ & _55430_ /*4585*/;
assign _55434_ = _54647_ ^ _55430_ /*4588*/;
assign _55435_ = _55426_ & _55434_ /*4586*/;
assign _55095_ = _55426_ ^ _55434_ /*4587*/;
assign _55432_ = _55433_ | _55435_ /*4584*/;
assign _55437_ = ~Q[2] /*4583*/;
assign _55436_ = _55437_ & D[55] /*4582*/;
assign _55439_ = _54648_ & _55436_ /*4577*/;
assign _55440_ = _54648_ ^ _55436_ /*4580*/;
assign _55441_ = _55432_ & _55440_ /*4578*/;
assign _55096_ = _55432_ ^ _55440_ /*4579*/;
assign _55438_ = _55439_ | _55441_ /*4576*/;
assign _55443_ = ~Q[2] /*4575*/;
assign _55442_ = _55443_ & D[56] /*4574*/;
assign _55445_ = _54649_ & _55442_ /*4569*/;
assign _55446_ = _54649_ ^ _55442_ /*4572*/;
assign _55447_ = _55438_ & _55446_ /*4570*/;
assign _55097_ = _55438_ ^ _55446_ /*4571*/;
assign _55444_ = _55445_ | _55447_ /*4568*/;
assign _55449_ = ~Q[2] /*4567*/;
assign _55448_ = _55449_ & D[57] /*4566*/;
assign _55451_ = _54650_ & _55448_ /*4561*/;
assign _55452_ = _54650_ ^ _55448_ /*4564*/;
assign _55453_ = _55444_ & _55452_ /*4562*/;
assign _55098_ = _55444_ ^ _55452_ /*4563*/;
assign _55450_ = _55451_ | _55453_ /*4560*/;
assign _55455_ = ~Q[2] /*4559*/;
assign _55454_ = _55455_ & D[58] /*4558*/;
assign _55457_ = _54651_ & _55454_ /*4553*/;
assign _55458_ = _54651_ ^ _55454_ /*4556*/;
assign _55459_ = _55450_ & _55458_ /*4554*/;
assign _55099_ = _55450_ ^ _55458_ /*4555*/;
assign _55456_ = _55457_ | _55459_ /*4552*/;
assign _55461_ = ~Q[2] /*4551*/;
assign _55460_ = _55461_ & D[59] /*4550*/;
assign _55463_ = _54652_ & _55460_ /*4545*/;
assign _55464_ = _54652_ ^ _55460_ /*4548*/;
assign _55465_ = _55456_ & _55464_ /*4546*/;
assign _55100_ = _55456_ ^ _55464_ /*4547*/;
assign _55462_ = _55463_ | _55465_ /*4544*/;
assign _55467_ = ~Q[2] /*4543*/;
assign _55466_ = _55467_ & D[60] /*4542*/;
assign _55469_ = _54653_ & _55466_ /*4537*/;
assign _55470_ = _54653_ ^ _55466_ /*4540*/;
assign _55471_ = _55462_ & _55470_ /*4538*/;
assign _55101_ = _55462_ ^ _55470_ /*4539*/;
assign _55468_ = _55469_ | _55471_ /*4536*/;
assign _55473_ = ~Q[2] /*4535*/;
assign _55472_ = _55473_ & D[61] /*4534*/;
assign _55475_ = _54654_ & _55472_ /*4529*/;
assign _55476_ = _54654_ ^ _55472_ /*4532*/;
assign _55477_ = _55468_ & _55476_ /*4530*/;
assign _55102_ = _55468_ ^ _55476_ /*4531*/;
assign _55474_ = _55475_ | _55477_ /*4528*/;
assign _55479_ = ~Q[2] /*4527*/;
assign _55478_ = _55479_ & D[62] /*4526*/;
assign _55481_ = _54655_ & _55478_ /*4521*/;
assign _55482_ = _54655_ ^ _55478_ /*4524*/;
assign _55483_ = _55474_ & _55482_ /*4522*/;
assign _55103_ = _55474_ ^ _55482_ /*4523*/;
assign _55480_ = _55481_ | _55483_ /*4520*/;
assign _55485_ = ~Q[2] /*4519*/;
assign _55484_ = _55485_ & zeroWire /*4518*/;
assign _55486_ = _54656_ ^ _55484_ /*4516*/;
assign _55104_ = _55486_ ^ _55480_ /*4515*/;
assign _55557_ = ~D[0] /*4261*/;
assign _55554_ = R_0[1] & _55557_ /*4257*/;
assign _55555_ = R_0[1] ^ _55557_ /*4260*/;
assign _55556_ = oneWire & _55555_ /*4258*/;
assign _55489_ = oneWire ^ _55555_ /*4259*/;
assign _55553_ = _55554_ | _55556_ /*4256*/;
assign _55562_ = ~D[1] /*4255*/;
assign _55559_ = _55041_ & _55562_ /*4251*/;
assign _55560_ = _55041_ ^ _55562_ /*4254*/;
assign _55561_ = _55553_ & _55560_ /*4252*/;
assign _55490_ = _55553_ ^ _55560_ /*4253*/;
assign _55558_ = _55559_ | _55561_ /*4250*/;
assign _55567_ = ~D[2] /*4249*/;
assign _55564_ = _55042_ & _55567_ /*4245*/;
assign _55565_ = _55042_ ^ _55567_ /*4248*/;
assign _55566_ = _55558_ & _55565_ /*4246*/;
assign _55491_ = _55558_ ^ _55565_ /*4247*/;
assign _55563_ = _55564_ | _55566_ /*4244*/;
assign _55572_ = ~D[3] /*4243*/;
assign _55569_ = _55043_ & _55572_ /*4239*/;
assign _55570_ = _55043_ ^ _55572_ /*4242*/;
assign _55571_ = _55563_ & _55570_ /*4240*/;
assign _55492_ = _55563_ ^ _55570_ /*4241*/;
assign _55568_ = _55569_ | _55571_ /*4238*/;
assign _55577_ = ~D[4] /*4237*/;
assign _55574_ = _55044_ & _55577_ /*4233*/;
assign _55575_ = _55044_ ^ _55577_ /*4236*/;
assign _55576_ = _55568_ & _55575_ /*4234*/;
assign _55493_ = _55568_ ^ _55575_ /*4235*/;
assign _55573_ = _55574_ | _55576_ /*4232*/;
assign _55582_ = ~D[5] /*4231*/;
assign _55579_ = _55045_ & _55582_ /*4227*/;
assign _55580_ = _55045_ ^ _55582_ /*4230*/;
assign _55581_ = _55573_ & _55580_ /*4228*/;
assign _55494_ = _55573_ ^ _55580_ /*4229*/;
assign _55578_ = _55579_ | _55581_ /*4226*/;
assign _55587_ = ~D[6] /*4225*/;
assign _55584_ = _55046_ & _55587_ /*4221*/;
assign _55585_ = _55046_ ^ _55587_ /*4224*/;
assign _55586_ = _55578_ & _55585_ /*4222*/;
assign _55495_ = _55578_ ^ _55585_ /*4223*/;
assign _55583_ = _55584_ | _55586_ /*4220*/;
assign _55592_ = ~D[7] /*4219*/;
assign _55589_ = _55047_ & _55592_ /*4215*/;
assign _55590_ = _55047_ ^ _55592_ /*4218*/;
assign _55591_ = _55583_ & _55590_ /*4216*/;
assign _55496_ = _55583_ ^ _55590_ /*4217*/;
assign _55588_ = _55589_ | _55591_ /*4214*/;
assign _55597_ = ~D[8] /*4213*/;
assign _55594_ = _55048_ & _55597_ /*4209*/;
assign _55595_ = _55048_ ^ _55597_ /*4212*/;
assign _55596_ = _55588_ & _55595_ /*4210*/;
assign _55497_ = _55588_ ^ _55595_ /*4211*/;
assign _55593_ = _55594_ | _55596_ /*4208*/;
assign _55602_ = ~D[9] /*4207*/;
assign _55599_ = _55049_ & _55602_ /*4203*/;
assign _55600_ = _55049_ ^ _55602_ /*4206*/;
assign _55601_ = _55593_ & _55600_ /*4204*/;
assign _55498_ = _55593_ ^ _55600_ /*4205*/;
assign _55598_ = _55599_ | _55601_ /*4202*/;
assign _55607_ = ~D[10] /*4201*/;
assign _55604_ = _55050_ & _55607_ /*4197*/;
assign _55605_ = _55050_ ^ _55607_ /*4200*/;
assign _55606_ = _55598_ & _55605_ /*4198*/;
assign _55499_ = _55598_ ^ _55605_ /*4199*/;
assign _55603_ = _55604_ | _55606_ /*4196*/;
assign _55612_ = ~D[11] /*4195*/;
assign _55609_ = _55051_ & _55612_ /*4191*/;
assign _55610_ = _55051_ ^ _55612_ /*4194*/;
assign _55611_ = _55603_ & _55610_ /*4192*/;
assign _55500_ = _55603_ ^ _55610_ /*4193*/;
assign _55608_ = _55609_ | _55611_ /*4190*/;
assign _55617_ = ~D[12] /*4189*/;
assign _55614_ = _55052_ & _55617_ /*4185*/;
assign _55615_ = _55052_ ^ _55617_ /*4188*/;
assign _55616_ = _55608_ & _55615_ /*4186*/;
assign _55501_ = _55608_ ^ _55615_ /*4187*/;
assign _55613_ = _55614_ | _55616_ /*4184*/;
assign _55622_ = ~D[13] /*4183*/;
assign _55619_ = _55053_ & _55622_ /*4179*/;
assign _55620_ = _55053_ ^ _55622_ /*4182*/;
assign _55621_ = _55613_ & _55620_ /*4180*/;
assign _55502_ = _55613_ ^ _55620_ /*4181*/;
assign _55618_ = _55619_ | _55621_ /*4178*/;
assign _55627_ = ~D[14] /*4177*/;
assign _55624_ = _55054_ & _55627_ /*4173*/;
assign _55625_ = _55054_ ^ _55627_ /*4176*/;
assign _55626_ = _55618_ & _55625_ /*4174*/;
assign _55503_ = _55618_ ^ _55625_ /*4175*/;
assign _55623_ = _55624_ | _55626_ /*4172*/;
assign _55632_ = ~D[15] /*4171*/;
assign _55629_ = _55055_ & _55632_ /*4167*/;
assign _55630_ = _55055_ ^ _55632_ /*4170*/;
assign _55631_ = _55623_ & _55630_ /*4168*/;
assign _55504_ = _55623_ ^ _55630_ /*4169*/;
assign _55628_ = _55629_ | _55631_ /*4166*/;
assign _55637_ = ~D[16] /*4165*/;
assign _55634_ = _55056_ & _55637_ /*4161*/;
assign _55635_ = _55056_ ^ _55637_ /*4164*/;
assign _55636_ = _55628_ & _55635_ /*4162*/;
assign _55505_ = _55628_ ^ _55635_ /*4163*/;
assign _55633_ = _55634_ | _55636_ /*4160*/;
assign _55642_ = ~D[17] /*4159*/;
assign _55639_ = _55057_ & _55642_ /*4155*/;
assign _55640_ = _55057_ ^ _55642_ /*4158*/;
assign _55641_ = _55633_ & _55640_ /*4156*/;
assign _55506_ = _55633_ ^ _55640_ /*4157*/;
assign _55638_ = _55639_ | _55641_ /*4154*/;
assign _55647_ = ~D[18] /*4153*/;
assign _55644_ = _55058_ & _55647_ /*4149*/;
assign _55645_ = _55058_ ^ _55647_ /*4152*/;
assign _55646_ = _55638_ & _55645_ /*4150*/;
assign _55507_ = _55638_ ^ _55645_ /*4151*/;
assign _55643_ = _55644_ | _55646_ /*4148*/;
assign _55652_ = ~D[19] /*4147*/;
assign _55649_ = _55059_ & _55652_ /*4143*/;
assign _55650_ = _55059_ ^ _55652_ /*4146*/;
assign _55651_ = _55643_ & _55650_ /*4144*/;
assign _55508_ = _55643_ ^ _55650_ /*4145*/;
assign _55648_ = _55649_ | _55651_ /*4142*/;
assign _55657_ = ~D[20] /*4141*/;
assign _55654_ = _55060_ & _55657_ /*4137*/;
assign _55655_ = _55060_ ^ _55657_ /*4140*/;
assign _55656_ = _55648_ & _55655_ /*4138*/;
assign _55509_ = _55648_ ^ _55655_ /*4139*/;
assign _55653_ = _55654_ | _55656_ /*4136*/;
assign _55662_ = ~D[21] /*4135*/;
assign _55659_ = _55061_ & _55662_ /*4131*/;
assign _55660_ = _55061_ ^ _55662_ /*4134*/;
assign _55661_ = _55653_ & _55660_ /*4132*/;
assign _55510_ = _55653_ ^ _55660_ /*4133*/;
assign _55658_ = _55659_ | _55661_ /*4130*/;
assign _55667_ = ~D[22] /*4129*/;
assign _55664_ = _55062_ & _55667_ /*4125*/;
assign _55665_ = _55062_ ^ _55667_ /*4128*/;
assign _55666_ = _55658_ & _55665_ /*4126*/;
assign _55511_ = _55658_ ^ _55665_ /*4127*/;
assign _55663_ = _55664_ | _55666_ /*4124*/;
assign _55672_ = ~D[23] /*4123*/;
assign _55669_ = _55063_ & _55672_ /*4119*/;
assign _55670_ = _55063_ ^ _55672_ /*4122*/;
assign _55671_ = _55663_ & _55670_ /*4120*/;
assign _55512_ = _55663_ ^ _55670_ /*4121*/;
assign _55668_ = _55669_ | _55671_ /*4118*/;
assign _55677_ = ~D[24] /*4117*/;
assign _55674_ = _55064_ & _55677_ /*4113*/;
assign _55675_ = _55064_ ^ _55677_ /*4116*/;
assign _55676_ = _55668_ & _55675_ /*4114*/;
assign _55513_ = _55668_ ^ _55675_ /*4115*/;
assign _55673_ = _55674_ | _55676_ /*4112*/;
assign _55682_ = ~D[25] /*4111*/;
assign _55679_ = _55065_ & _55682_ /*4107*/;
assign _55680_ = _55065_ ^ _55682_ /*4110*/;
assign _55681_ = _55673_ & _55680_ /*4108*/;
assign _55514_ = _55673_ ^ _55680_ /*4109*/;
assign _55678_ = _55679_ | _55681_ /*4106*/;
assign _55687_ = ~D[26] /*4105*/;
assign _55684_ = _55066_ & _55687_ /*4101*/;
assign _55685_ = _55066_ ^ _55687_ /*4104*/;
assign _55686_ = _55678_ & _55685_ /*4102*/;
assign _55515_ = _55678_ ^ _55685_ /*4103*/;
assign _55683_ = _55684_ | _55686_ /*4100*/;
assign _55692_ = ~D[27] /*4099*/;
assign _55689_ = _55067_ & _55692_ /*4095*/;
assign _55690_ = _55067_ ^ _55692_ /*4098*/;
assign _55691_ = _55683_ & _55690_ /*4096*/;
assign _55516_ = _55683_ ^ _55690_ /*4097*/;
assign _55688_ = _55689_ | _55691_ /*4094*/;
assign _55697_ = ~D[28] /*4093*/;
assign _55694_ = _55068_ & _55697_ /*4089*/;
assign _55695_ = _55068_ ^ _55697_ /*4092*/;
assign _55696_ = _55688_ & _55695_ /*4090*/;
assign _55517_ = _55688_ ^ _55695_ /*4091*/;
assign _55693_ = _55694_ | _55696_ /*4088*/;
assign _55702_ = ~D[29] /*4087*/;
assign _55699_ = _55069_ & _55702_ /*4083*/;
assign _55700_ = _55069_ ^ _55702_ /*4086*/;
assign _55701_ = _55693_ & _55700_ /*4084*/;
assign _55518_ = _55693_ ^ _55700_ /*4085*/;
assign _55698_ = _55699_ | _55701_ /*4082*/;
assign _55707_ = ~D[30] /*4081*/;
assign _55704_ = _55070_ & _55707_ /*4077*/;
assign _55705_ = _55070_ ^ _55707_ /*4080*/;
assign _55706_ = _55698_ & _55705_ /*4078*/;
assign _55519_ = _55698_ ^ _55705_ /*4079*/;
assign _55703_ = _55704_ | _55706_ /*4076*/;
assign _55712_ = ~D[31] /*4075*/;
assign _55709_ = _55071_ & _55712_ /*4071*/;
assign _55710_ = _55071_ ^ _55712_ /*4074*/;
assign _55711_ = _55703_ & _55710_ /*4072*/;
assign _55520_ = _55703_ ^ _55710_ /*4073*/;
assign _55708_ = _55709_ | _55711_ /*4070*/;
assign _55717_ = ~D[32] /*4069*/;
assign _55714_ = _55072_ & _55717_ /*4065*/;
assign _55715_ = _55072_ ^ _55717_ /*4068*/;
assign _55716_ = _55708_ & _55715_ /*4066*/;
assign _55521_ = _55708_ ^ _55715_ /*4067*/;
assign _55713_ = _55714_ | _55716_ /*4064*/;
assign _55722_ = ~D[33] /*4063*/;
assign _55719_ = _55073_ & _55722_ /*4059*/;
assign _55720_ = _55073_ ^ _55722_ /*4062*/;
assign _55721_ = _55713_ & _55720_ /*4060*/;
assign _55522_ = _55713_ ^ _55720_ /*4061*/;
assign _55718_ = _55719_ | _55721_ /*4058*/;
assign _55727_ = ~D[34] /*4057*/;
assign _55724_ = _55074_ & _55727_ /*4053*/;
assign _55725_ = _55074_ ^ _55727_ /*4056*/;
assign _55726_ = _55718_ & _55725_ /*4054*/;
assign _55523_ = _55718_ ^ _55725_ /*4055*/;
assign _55723_ = _55724_ | _55726_ /*4052*/;
assign _55732_ = ~D[35] /*4051*/;
assign _55729_ = _55075_ & _55732_ /*4047*/;
assign _55730_ = _55075_ ^ _55732_ /*4050*/;
assign _55731_ = _55723_ & _55730_ /*4048*/;
assign _55524_ = _55723_ ^ _55730_ /*4049*/;
assign _55728_ = _55729_ | _55731_ /*4046*/;
assign _55737_ = ~D[36] /*4045*/;
assign _55734_ = _55076_ & _55737_ /*4041*/;
assign _55735_ = _55076_ ^ _55737_ /*4044*/;
assign _55736_ = _55728_ & _55735_ /*4042*/;
assign _55525_ = _55728_ ^ _55735_ /*4043*/;
assign _55733_ = _55734_ | _55736_ /*4040*/;
assign _55742_ = ~D[37] /*4039*/;
assign _55739_ = _55077_ & _55742_ /*4035*/;
assign _55740_ = _55077_ ^ _55742_ /*4038*/;
assign _55741_ = _55733_ & _55740_ /*4036*/;
assign _55526_ = _55733_ ^ _55740_ /*4037*/;
assign _55738_ = _55739_ | _55741_ /*4034*/;
assign _55747_ = ~D[38] /*4033*/;
assign _55744_ = _55078_ & _55747_ /*4029*/;
assign _55745_ = _55078_ ^ _55747_ /*4032*/;
assign _55746_ = _55738_ & _55745_ /*4030*/;
assign _55527_ = _55738_ ^ _55745_ /*4031*/;
assign _55743_ = _55744_ | _55746_ /*4028*/;
assign _55752_ = ~D[39] /*4027*/;
assign _55749_ = _55079_ & _55752_ /*4023*/;
assign _55750_ = _55079_ ^ _55752_ /*4026*/;
assign _55751_ = _55743_ & _55750_ /*4024*/;
assign _55528_ = _55743_ ^ _55750_ /*4025*/;
assign _55748_ = _55749_ | _55751_ /*4022*/;
assign _55757_ = ~D[40] /*4021*/;
assign _55754_ = _55080_ & _55757_ /*4017*/;
assign _55755_ = _55080_ ^ _55757_ /*4020*/;
assign _55756_ = _55748_ & _55755_ /*4018*/;
assign _55529_ = _55748_ ^ _55755_ /*4019*/;
assign _55753_ = _55754_ | _55756_ /*4016*/;
assign _55762_ = ~D[41] /*4015*/;
assign _55759_ = _55081_ & _55762_ /*4011*/;
assign _55760_ = _55081_ ^ _55762_ /*4014*/;
assign _55761_ = _55753_ & _55760_ /*4012*/;
assign _55530_ = _55753_ ^ _55760_ /*4013*/;
assign _55758_ = _55759_ | _55761_ /*4010*/;
assign _55767_ = ~D[42] /*4009*/;
assign _55764_ = _55082_ & _55767_ /*4005*/;
assign _55765_ = _55082_ ^ _55767_ /*4008*/;
assign _55766_ = _55758_ & _55765_ /*4006*/;
assign _55531_ = _55758_ ^ _55765_ /*4007*/;
assign _55763_ = _55764_ | _55766_ /*4004*/;
assign _55772_ = ~D[43] /*4003*/;
assign _55769_ = _55083_ & _55772_ /*3999*/;
assign _55770_ = _55083_ ^ _55772_ /*4002*/;
assign _55771_ = _55763_ & _55770_ /*4000*/;
assign _55532_ = _55763_ ^ _55770_ /*4001*/;
assign _55768_ = _55769_ | _55771_ /*3998*/;
assign _55777_ = ~D[44] /*3997*/;
assign _55774_ = _55084_ & _55777_ /*3993*/;
assign _55775_ = _55084_ ^ _55777_ /*3996*/;
assign _55776_ = _55768_ & _55775_ /*3994*/;
assign _55533_ = _55768_ ^ _55775_ /*3995*/;
assign _55773_ = _55774_ | _55776_ /*3992*/;
assign _55782_ = ~D[45] /*3991*/;
assign _55779_ = _55085_ & _55782_ /*3987*/;
assign _55780_ = _55085_ ^ _55782_ /*3990*/;
assign _55781_ = _55773_ & _55780_ /*3988*/;
assign _55534_ = _55773_ ^ _55780_ /*3989*/;
assign _55778_ = _55779_ | _55781_ /*3986*/;
assign _55787_ = ~D[46] /*3985*/;
assign _55784_ = _55086_ & _55787_ /*3981*/;
assign _55785_ = _55086_ ^ _55787_ /*3984*/;
assign _55786_ = _55778_ & _55785_ /*3982*/;
assign _55535_ = _55778_ ^ _55785_ /*3983*/;
assign _55783_ = _55784_ | _55786_ /*3980*/;
assign _55792_ = ~D[47] /*3979*/;
assign _55789_ = _55087_ & _55792_ /*3975*/;
assign _55790_ = _55087_ ^ _55792_ /*3978*/;
assign _55791_ = _55783_ & _55790_ /*3976*/;
assign _55536_ = _55783_ ^ _55790_ /*3977*/;
assign _55788_ = _55789_ | _55791_ /*3974*/;
assign _55797_ = ~D[48] /*3973*/;
assign _55794_ = _55088_ & _55797_ /*3969*/;
assign _55795_ = _55088_ ^ _55797_ /*3972*/;
assign _55796_ = _55788_ & _55795_ /*3970*/;
assign _55537_ = _55788_ ^ _55795_ /*3971*/;
assign _55793_ = _55794_ | _55796_ /*3968*/;
assign _55802_ = ~D[49] /*3967*/;
assign _55799_ = _55089_ & _55802_ /*3963*/;
assign _55800_ = _55089_ ^ _55802_ /*3966*/;
assign _55801_ = _55793_ & _55800_ /*3964*/;
assign _55538_ = _55793_ ^ _55800_ /*3965*/;
assign _55798_ = _55799_ | _55801_ /*3962*/;
assign _55807_ = ~D[50] /*3961*/;
assign _55804_ = _55090_ & _55807_ /*3957*/;
assign _55805_ = _55090_ ^ _55807_ /*3960*/;
assign _55806_ = _55798_ & _55805_ /*3958*/;
assign _55539_ = _55798_ ^ _55805_ /*3959*/;
assign _55803_ = _55804_ | _55806_ /*3956*/;
assign _55812_ = ~D[51] /*3955*/;
assign _55809_ = _55091_ & _55812_ /*3951*/;
assign _55810_ = _55091_ ^ _55812_ /*3954*/;
assign _55811_ = _55803_ & _55810_ /*3952*/;
assign _55540_ = _55803_ ^ _55810_ /*3953*/;
assign _55808_ = _55809_ | _55811_ /*3950*/;
assign _55817_ = ~D[52] /*3949*/;
assign _55814_ = _55092_ & _55817_ /*3945*/;
assign _55815_ = _55092_ ^ _55817_ /*3948*/;
assign _55816_ = _55808_ & _55815_ /*3946*/;
assign _55541_ = _55808_ ^ _55815_ /*3947*/;
assign _55813_ = _55814_ | _55816_ /*3944*/;
assign _55822_ = ~D[53] /*3943*/;
assign _55819_ = _55093_ & _55822_ /*3939*/;
assign _55820_ = _55093_ ^ _55822_ /*3942*/;
assign _55821_ = _55813_ & _55820_ /*3940*/;
assign _55542_ = _55813_ ^ _55820_ /*3941*/;
assign _55818_ = _55819_ | _55821_ /*3938*/;
assign _55827_ = ~D[54] /*3937*/;
assign _55824_ = _55094_ & _55827_ /*3933*/;
assign _55825_ = _55094_ ^ _55827_ /*3936*/;
assign _55826_ = _55818_ & _55825_ /*3934*/;
assign _55543_ = _55818_ ^ _55825_ /*3935*/;
assign _55823_ = _55824_ | _55826_ /*3932*/;
assign _55832_ = ~D[55] /*3931*/;
assign _55829_ = _55095_ & _55832_ /*3927*/;
assign _55830_ = _55095_ ^ _55832_ /*3930*/;
assign _55831_ = _55823_ & _55830_ /*3928*/;
assign _55544_ = _55823_ ^ _55830_ /*3929*/;
assign _55828_ = _55829_ | _55831_ /*3926*/;
assign _55837_ = ~D[56] /*3925*/;
assign _55834_ = _55096_ & _55837_ /*3921*/;
assign _55835_ = _55096_ ^ _55837_ /*3924*/;
assign _55836_ = _55828_ & _55835_ /*3922*/;
assign _55545_ = _55828_ ^ _55835_ /*3923*/;
assign _55833_ = _55834_ | _55836_ /*3920*/;
assign _55842_ = ~D[57] /*3919*/;
assign _55839_ = _55097_ & _55842_ /*3915*/;
assign _55840_ = _55097_ ^ _55842_ /*3918*/;
assign _55841_ = _55833_ & _55840_ /*3916*/;
assign _55546_ = _55833_ ^ _55840_ /*3917*/;
assign _55838_ = _55839_ | _55841_ /*3914*/;
assign _55847_ = ~D[58] /*3913*/;
assign _55844_ = _55098_ & _55847_ /*3909*/;
assign _55845_ = _55098_ ^ _55847_ /*3912*/;
assign _55846_ = _55838_ & _55845_ /*3910*/;
assign _55547_ = _55838_ ^ _55845_ /*3911*/;
assign _55843_ = _55844_ | _55846_ /*3908*/;
assign _55852_ = ~D[59] /*3907*/;
assign _55849_ = _55099_ & _55852_ /*3903*/;
assign _55850_ = _55099_ ^ _55852_ /*3906*/;
assign _55851_ = _55843_ & _55850_ /*3904*/;
assign _55548_ = _55843_ ^ _55850_ /*3905*/;
assign _55848_ = _55849_ | _55851_ /*3902*/;
assign _55857_ = ~D[60] /*3901*/;
assign _55854_ = _55100_ & _55857_ /*3897*/;
assign _55855_ = _55100_ ^ _55857_ /*3900*/;
assign _55856_ = _55848_ & _55855_ /*3898*/;
assign _55549_ = _55848_ ^ _55855_ /*3899*/;
assign _55853_ = _55854_ | _55856_ /*3896*/;
assign _55862_ = ~D[61] /*3895*/;
assign _55859_ = _55101_ & _55862_ /*3891*/;
assign _55860_ = _55101_ ^ _55862_ /*3894*/;
assign _55861_ = _55853_ & _55860_ /*3892*/;
assign _55550_ = _55853_ ^ _55860_ /*3893*/;
assign _55858_ = _55859_ | _55861_ /*3890*/;
assign _55867_ = ~D[62] /*3889*/;
assign _55864_ = _55102_ & _55867_ /*3885*/;
assign _55865_ = _55102_ ^ _55867_ /*3888*/;
assign _55866_ = _55858_ & _55865_ /*3886*/;
assign _55551_ = _55858_ ^ _55865_ /*3887*/;
assign _55863_ = _55864_ | _55866_ /*3884*/;
assign _55868_ = _55103_ & oneWire /*3879*/;
assign _55869_ = _55103_ ^ oneWire /*3882*/;
assign _55870_ = _55863_ & _55869_ /*3880*/;
assign _55552_ = _55863_ ^ _55869_ /*3881*/;
assign Q[1] = _55868_ | _55870_ /*3878*/;
assign _56003_ = ~Q[1] /*3493*/;
assign _56002_ = _56003_ & D[0] /*3492*/;
assign _56005_ = _55489_ & _56002_ /*3487*/;
assign _56006_ = _55489_ ^ _56002_ /*3490*/;
assign _56007_ = zeroWire & _56006_ /*3488*/;
assign _55937_ = zeroWire ^ _56006_ /*3489*/;
assign _56004_ = _56005_ | _56007_ /*3486*/;
assign _56009_ = ~Q[1] /*3485*/;
assign _56008_ = _56009_ & D[1] /*3484*/;
assign _56011_ = _55490_ & _56008_ /*3479*/;
assign _56012_ = _55490_ ^ _56008_ /*3482*/;
assign _56013_ = _56004_ & _56012_ /*3480*/;
assign _55938_ = _56004_ ^ _56012_ /*3481*/;
assign _56010_ = _56011_ | _56013_ /*3478*/;
assign _56015_ = ~Q[1] /*3477*/;
assign _56014_ = _56015_ & D[2] /*3476*/;
assign _56017_ = _55491_ & _56014_ /*3471*/;
assign _56018_ = _55491_ ^ _56014_ /*3474*/;
assign _56019_ = _56010_ & _56018_ /*3472*/;
assign _55939_ = _56010_ ^ _56018_ /*3473*/;
assign _56016_ = _56017_ | _56019_ /*3470*/;
assign _56021_ = ~Q[1] /*3469*/;
assign _56020_ = _56021_ & D[3] /*3468*/;
assign _56023_ = _55492_ & _56020_ /*3463*/;
assign _56024_ = _55492_ ^ _56020_ /*3466*/;
assign _56025_ = _56016_ & _56024_ /*3464*/;
assign _55940_ = _56016_ ^ _56024_ /*3465*/;
assign _56022_ = _56023_ | _56025_ /*3462*/;
assign _56027_ = ~Q[1] /*3461*/;
assign _56026_ = _56027_ & D[4] /*3460*/;
assign _56029_ = _55493_ & _56026_ /*3455*/;
assign _56030_ = _55493_ ^ _56026_ /*3458*/;
assign _56031_ = _56022_ & _56030_ /*3456*/;
assign _55941_ = _56022_ ^ _56030_ /*3457*/;
assign _56028_ = _56029_ | _56031_ /*3454*/;
assign _56033_ = ~Q[1] /*3453*/;
assign _56032_ = _56033_ & D[5] /*3452*/;
assign _56035_ = _55494_ & _56032_ /*3447*/;
assign _56036_ = _55494_ ^ _56032_ /*3450*/;
assign _56037_ = _56028_ & _56036_ /*3448*/;
assign _55942_ = _56028_ ^ _56036_ /*3449*/;
assign _56034_ = _56035_ | _56037_ /*3446*/;
assign _56039_ = ~Q[1] /*3445*/;
assign _56038_ = _56039_ & D[6] /*3444*/;
assign _56041_ = _55495_ & _56038_ /*3439*/;
assign _56042_ = _55495_ ^ _56038_ /*3442*/;
assign _56043_ = _56034_ & _56042_ /*3440*/;
assign _55943_ = _56034_ ^ _56042_ /*3441*/;
assign _56040_ = _56041_ | _56043_ /*3438*/;
assign _56045_ = ~Q[1] /*3437*/;
assign _56044_ = _56045_ & D[7] /*3436*/;
assign _56047_ = _55496_ & _56044_ /*3431*/;
assign _56048_ = _55496_ ^ _56044_ /*3434*/;
assign _56049_ = _56040_ & _56048_ /*3432*/;
assign _55944_ = _56040_ ^ _56048_ /*3433*/;
assign _56046_ = _56047_ | _56049_ /*3430*/;
assign _56051_ = ~Q[1] /*3429*/;
assign _56050_ = _56051_ & D[8] /*3428*/;
assign _56053_ = _55497_ & _56050_ /*3423*/;
assign _56054_ = _55497_ ^ _56050_ /*3426*/;
assign _56055_ = _56046_ & _56054_ /*3424*/;
assign _55945_ = _56046_ ^ _56054_ /*3425*/;
assign _56052_ = _56053_ | _56055_ /*3422*/;
assign _56057_ = ~Q[1] /*3421*/;
assign _56056_ = _56057_ & D[9] /*3420*/;
assign _56059_ = _55498_ & _56056_ /*3415*/;
assign _56060_ = _55498_ ^ _56056_ /*3418*/;
assign _56061_ = _56052_ & _56060_ /*3416*/;
assign _55946_ = _56052_ ^ _56060_ /*3417*/;
assign _56058_ = _56059_ | _56061_ /*3414*/;
assign _56063_ = ~Q[1] /*3413*/;
assign _56062_ = _56063_ & D[10] /*3412*/;
assign _56065_ = _55499_ & _56062_ /*3407*/;
assign _56066_ = _55499_ ^ _56062_ /*3410*/;
assign _56067_ = _56058_ & _56066_ /*3408*/;
assign _55947_ = _56058_ ^ _56066_ /*3409*/;
assign _56064_ = _56065_ | _56067_ /*3406*/;
assign _56069_ = ~Q[1] /*3405*/;
assign _56068_ = _56069_ & D[11] /*3404*/;
assign _56071_ = _55500_ & _56068_ /*3399*/;
assign _56072_ = _55500_ ^ _56068_ /*3402*/;
assign _56073_ = _56064_ & _56072_ /*3400*/;
assign _55948_ = _56064_ ^ _56072_ /*3401*/;
assign _56070_ = _56071_ | _56073_ /*3398*/;
assign _56075_ = ~Q[1] /*3397*/;
assign _56074_ = _56075_ & D[12] /*3396*/;
assign _56077_ = _55501_ & _56074_ /*3391*/;
assign _56078_ = _55501_ ^ _56074_ /*3394*/;
assign _56079_ = _56070_ & _56078_ /*3392*/;
assign _55949_ = _56070_ ^ _56078_ /*3393*/;
assign _56076_ = _56077_ | _56079_ /*3390*/;
assign _56081_ = ~Q[1] /*3389*/;
assign _56080_ = _56081_ & D[13] /*3388*/;
assign _56083_ = _55502_ & _56080_ /*3383*/;
assign _56084_ = _55502_ ^ _56080_ /*3386*/;
assign _56085_ = _56076_ & _56084_ /*3384*/;
assign _55950_ = _56076_ ^ _56084_ /*3385*/;
assign _56082_ = _56083_ | _56085_ /*3382*/;
assign _56087_ = ~Q[1] /*3381*/;
assign _56086_ = _56087_ & D[14] /*3380*/;
assign _56089_ = _55503_ & _56086_ /*3375*/;
assign _56090_ = _55503_ ^ _56086_ /*3378*/;
assign _56091_ = _56082_ & _56090_ /*3376*/;
assign _55951_ = _56082_ ^ _56090_ /*3377*/;
assign _56088_ = _56089_ | _56091_ /*3374*/;
assign _56093_ = ~Q[1] /*3373*/;
assign _56092_ = _56093_ & D[15] /*3372*/;
assign _56095_ = _55504_ & _56092_ /*3367*/;
assign _56096_ = _55504_ ^ _56092_ /*3370*/;
assign _56097_ = _56088_ & _56096_ /*3368*/;
assign _55952_ = _56088_ ^ _56096_ /*3369*/;
assign _56094_ = _56095_ | _56097_ /*3366*/;
assign _56099_ = ~Q[1] /*3365*/;
assign _56098_ = _56099_ & D[16] /*3364*/;
assign _56101_ = _55505_ & _56098_ /*3359*/;
assign _56102_ = _55505_ ^ _56098_ /*3362*/;
assign _56103_ = _56094_ & _56102_ /*3360*/;
assign _55953_ = _56094_ ^ _56102_ /*3361*/;
assign _56100_ = _56101_ | _56103_ /*3358*/;
assign _56105_ = ~Q[1] /*3357*/;
assign _56104_ = _56105_ & D[17] /*3356*/;
assign _56107_ = _55506_ & _56104_ /*3351*/;
assign _56108_ = _55506_ ^ _56104_ /*3354*/;
assign _56109_ = _56100_ & _56108_ /*3352*/;
assign _55954_ = _56100_ ^ _56108_ /*3353*/;
assign _56106_ = _56107_ | _56109_ /*3350*/;
assign _56111_ = ~Q[1] /*3349*/;
assign _56110_ = _56111_ & D[18] /*3348*/;
assign _56113_ = _55507_ & _56110_ /*3343*/;
assign _56114_ = _55507_ ^ _56110_ /*3346*/;
assign _56115_ = _56106_ & _56114_ /*3344*/;
assign _55955_ = _56106_ ^ _56114_ /*3345*/;
assign _56112_ = _56113_ | _56115_ /*3342*/;
assign _56117_ = ~Q[1] /*3341*/;
assign _56116_ = _56117_ & D[19] /*3340*/;
assign _56119_ = _55508_ & _56116_ /*3335*/;
assign _56120_ = _55508_ ^ _56116_ /*3338*/;
assign _56121_ = _56112_ & _56120_ /*3336*/;
assign _55956_ = _56112_ ^ _56120_ /*3337*/;
assign _56118_ = _56119_ | _56121_ /*3334*/;
assign _56123_ = ~Q[1] /*3333*/;
assign _56122_ = _56123_ & D[20] /*3332*/;
assign _56125_ = _55509_ & _56122_ /*3327*/;
assign _56126_ = _55509_ ^ _56122_ /*3330*/;
assign _56127_ = _56118_ & _56126_ /*3328*/;
assign _55957_ = _56118_ ^ _56126_ /*3329*/;
assign _56124_ = _56125_ | _56127_ /*3326*/;
assign _56129_ = ~Q[1] /*3325*/;
assign _56128_ = _56129_ & D[21] /*3324*/;
assign _56131_ = _55510_ & _56128_ /*3319*/;
assign _56132_ = _55510_ ^ _56128_ /*3322*/;
assign _56133_ = _56124_ & _56132_ /*3320*/;
assign _55958_ = _56124_ ^ _56132_ /*3321*/;
assign _56130_ = _56131_ | _56133_ /*3318*/;
assign _56135_ = ~Q[1] /*3317*/;
assign _56134_ = _56135_ & D[22] /*3316*/;
assign _56137_ = _55511_ & _56134_ /*3311*/;
assign _56138_ = _55511_ ^ _56134_ /*3314*/;
assign _56139_ = _56130_ & _56138_ /*3312*/;
assign _55959_ = _56130_ ^ _56138_ /*3313*/;
assign _56136_ = _56137_ | _56139_ /*3310*/;
assign _56141_ = ~Q[1] /*3309*/;
assign _56140_ = _56141_ & D[23] /*3308*/;
assign _56143_ = _55512_ & _56140_ /*3303*/;
assign _56144_ = _55512_ ^ _56140_ /*3306*/;
assign _56145_ = _56136_ & _56144_ /*3304*/;
assign _55960_ = _56136_ ^ _56144_ /*3305*/;
assign _56142_ = _56143_ | _56145_ /*3302*/;
assign _56147_ = ~Q[1] /*3301*/;
assign _56146_ = _56147_ & D[24] /*3300*/;
assign _56149_ = _55513_ & _56146_ /*3295*/;
assign _56150_ = _55513_ ^ _56146_ /*3298*/;
assign _56151_ = _56142_ & _56150_ /*3296*/;
assign _55961_ = _56142_ ^ _56150_ /*3297*/;
assign _56148_ = _56149_ | _56151_ /*3294*/;
assign _56153_ = ~Q[1] /*3293*/;
assign _56152_ = _56153_ & D[25] /*3292*/;
assign _56155_ = _55514_ & _56152_ /*3287*/;
assign _56156_ = _55514_ ^ _56152_ /*3290*/;
assign _56157_ = _56148_ & _56156_ /*3288*/;
assign _55962_ = _56148_ ^ _56156_ /*3289*/;
assign _56154_ = _56155_ | _56157_ /*3286*/;
assign _56159_ = ~Q[1] /*3285*/;
assign _56158_ = _56159_ & D[26] /*3284*/;
assign _56161_ = _55515_ & _56158_ /*3279*/;
assign _56162_ = _55515_ ^ _56158_ /*3282*/;
assign _56163_ = _56154_ & _56162_ /*3280*/;
assign _55963_ = _56154_ ^ _56162_ /*3281*/;
assign _56160_ = _56161_ | _56163_ /*3278*/;
assign _56165_ = ~Q[1] /*3277*/;
assign _56164_ = _56165_ & D[27] /*3276*/;
assign _56167_ = _55516_ & _56164_ /*3271*/;
assign _56168_ = _55516_ ^ _56164_ /*3274*/;
assign _56169_ = _56160_ & _56168_ /*3272*/;
assign _55964_ = _56160_ ^ _56168_ /*3273*/;
assign _56166_ = _56167_ | _56169_ /*3270*/;
assign _56171_ = ~Q[1] /*3269*/;
assign _56170_ = _56171_ & D[28] /*3268*/;
assign _56173_ = _55517_ & _56170_ /*3263*/;
assign _56174_ = _55517_ ^ _56170_ /*3266*/;
assign _56175_ = _56166_ & _56174_ /*3264*/;
assign _55965_ = _56166_ ^ _56174_ /*3265*/;
assign _56172_ = _56173_ | _56175_ /*3262*/;
assign _56177_ = ~Q[1] /*3261*/;
assign _56176_ = _56177_ & D[29] /*3260*/;
assign _56179_ = _55518_ & _56176_ /*3255*/;
assign _56180_ = _55518_ ^ _56176_ /*3258*/;
assign _56181_ = _56172_ & _56180_ /*3256*/;
assign _55966_ = _56172_ ^ _56180_ /*3257*/;
assign _56178_ = _56179_ | _56181_ /*3254*/;
assign _56183_ = ~Q[1] /*3253*/;
assign _56182_ = _56183_ & D[30] /*3252*/;
assign _56185_ = _55519_ & _56182_ /*3247*/;
assign _56186_ = _55519_ ^ _56182_ /*3250*/;
assign _56187_ = _56178_ & _56186_ /*3248*/;
assign _55967_ = _56178_ ^ _56186_ /*3249*/;
assign _56184_ = _56185_ | _56187_ /*3246*/;
assign _56189_ = ~Q[1] /*3245*/;
assign _56188_ = _56189_ & D[31] /*3244*/;
assign _56191_ = _55520_ & _56188_ /*3239*/;
assign _56192_ = _55520_ ^ _56188_ /*3242*/;
assign _56193_ = _56184_ & _56192_ /*3240*/;
assign _55968_ = _56184_ ^ _56192_ /*3241*/;
assign _56190_ = _56191_ | _56193_ /*3238*/;
assign _56195_ = ~Q[1] /*3237*/;
assign _56194_ = _56195_ & D[32] /*3236*/;
assign _56197_ = _55521_ & _56194_ /*3231*/;
assign _56198_ = _55521_ ^ _56194_ /*3234*/;
assign _56199_ = _56190_ & _56198_ /*3232*/;
assign _55969_ = _56190_ ^ _56198_ /*3233*/;
assign _56196_ = _56197_ | _56199_ /*3230*/;
assign _56201_ = ~Q[1] /*3229*/;
assign _56200_ = _56201_ & D[33] /*3228*/;
assign _56203_ = _55522_ & _56200_ /*3223*/;
assign _56204_ = _55522_ ^ _56200_ /*3226*/;
assign _56205_ = _56196_ & _56204_ /*3224*/;
assign _55970_ = _56196_ ^ _56204_ /*3225*/;
assign _56202_ = _56203_ | _56205_ /*3222*/;
assign _56207_ = ~Q[1] /*3221*/;
assign _56206_ = _56207_ & D[34] /*3220*/;
assign _56209_ = _55523_ & _56206_ /*3215*/;
assign _56210_ = _55523_ ^ _56206_ /*3218*/;
assign _56211_ = _56202_ & _56210_ /*3216*/;
assign _55971_ = _56202_ ^ _56210_ /*3217*/;
assign _56208_ = _56209_ | _56211_ /*3214*/;
assign _56213_ = ~Q[1] /*3213*/;
assign _56212_ = _56213_ & D[35] /*3212*/;
assign _56215_ = _55524_ & _56212_ /*3207*/;
assign _56216_ = _55524_ ^ _56212_ /*3210*/;
assign _56217_ = _56208_ & _56216_ /*3208*/;
assign _55972_ = _56208_ ^ _56216_ /*3209*/;
assign _56214_ = _56215_ | _56217_ /*3206*/;
assign _56219_ = ~Q[1] /*3205*/;
assign _56218_ = _56219_ & D[36] /*3204*/;
assign _56221_ = _55525_ & _56218_ /*3199*/;
assign _56222_ = _55525_ ^ _56218_ /*3202*/;
assign _56223_ = _56214_ & _56222_ /*3200*/;
assign _55973_ = _56214_ ^ _56222_ /*3201*/;
assign _56220_ = _56221_ | _56223_ /*3198*/;
assign _56225_ = ~Q[1] /*3197*/;
assign _56224_ = _56225_ & D[37] /*3196*/;
assign _56227_ = _55526_ & _56224_ /*3191*/;
assign _56228_ = _55526_ ^ _56224_ /*3194*/;
assign _56229_ = _56220_ & _56228_ /*3192*/;
assign _55974_ = _56220_ ^ _56228_ /*3193*/;
assign _56226_ = _56227_ | _56229_ /*3190*/;
assign _56231_ = ~Q[1] /*3189*/;
assign _56230_ = _56231_ & D[38] /*3188*/;
assign _56233_ = _55527_ & _56230_ /*3183*/;
assign _56234_ = _55527_ ^ _56230_ /*3186*/;
assign _56235_ = _56226_ & _56234_ /*3184*/;
assign _55975_ = _56226_ ^ _56234_ /*3185*/;
assign _56232_ = _56233_ | _56235_ /*3182*/;
assign _56237_ = ~Q[1] /*3181*/;
assign _56236_ = _56237_ & D[39] /*3180*/;
assign _56239_ = _55528_ & _56236_ /*3175*/;
assign _56240_ = _55528_ ^ _56236_ /*3178*/;
assign _56241_ = _56232_ & _56240_ /*3176*/;
assign _55976_ = _56232_ ^ _56240_ /*3177*/;
assign _56238_ = _56239_ | _56241_ /*3174*/;
assign _56243_ = ~Q[1] /*3173*/;
assign _56242_ = _56243_ & D[40] /*3172*/;
assign _56245_ = _55529_ & _56242_ /*3167*/;
assign _56246_ = _55529_ ^ _56242_ /*3170*/;
assign _56247_ = _56238_ & _56246_ /*3168*/;
assign _55977_ = _56238_ ^ _56246_ /*3169*/;
assign _56244_ = _56245_ | _56247_ /*3166*/;
assign _56249_ = ~Q[1] /*3165*/;
assign _56248_ = _56249_ & D[41] /*3164*/;
assign _56251_ = _55530_ & _56248_ /*3159*/;
assign _56252_ = _55530_ ^ _56248_ /*3162*/;
assign _56253_ = _56244_ & _56252_ /*3160*/;
assign _55978_ = _56244_ ^ _56252_ /*3161*/;
assign _56250_ = _56251_ | _56253_ /*3158*/;
assign _56255_ = ~Q[1] /*3157*/;
assign _56254_ = _56255_ & D[42] /*3156*/;
assign _56257_ = _55531_ & _56254_ /*3151*/;
assign _56258_ = _55531_ ^ _56254_ /*3154*/;
assign _56259_ = _56250_ & _56258_ /*3152*/;
assign _55979_ = _56250_ ^ _56258_ /*3153*/;
assign _56256_ = _56257_ | _56259_ /*3150*/;
assign _56261_ = ~Q[1] /*3149*/;
assign _56260_ = _56261_ & D[43] /*3148*/;
assign _56263_ = _55532_ & _56260_ /*3143*/;
assign _56264_ = _55532_ ^ _56260_ /*3146*/;
assign _56265_ = _56256_ & _56264_ /*3144*/;
assign _55980_ = _56256_ ^ _56264_ /*3145*/;
assign _56262_ = _56263_ | _56265_ /*3142*/;
assign _56267_ = ~Q[1] /*3141*/;
assign _56266_ = _56267_ & D[44] /*3140*/;
assign _56269_ = _55533_ & _56266_ /*3135*/;
assign _56270_ = _55533_ ^ _56266_ /*3138*/;
assign _56271_ = _56262_ & _56270_ /*3136*/;
assign _55981_ = _56262_ ^ _56270_ /*3137*/;
assign _56268_ = _56269_ | _56271_ /*3134*/;
assign _56273_ = ~Q[1] /*3133*/;
assign _56272_ = _56273_ & D[45] /*3132*/;
assign _56275_ = _55534_ & _56272_ /*3127*/;
assign _56276_ = _55534_ ^ _56272_ /*3130*/;
assign _56277_ = _56268_ & _56276_ /*3128*/;
assign _55982_ = _56268_ ^ _56276_ /*3129*/;
assign _56274_ = _56275_ | _56277_ /*3126*/;
assign _56279_ = ~Q[1] /*3125*/;
assign _56278_ = _56279_ & D[46] /*3124*/;
assign _56281_ = _55535_ & _56278_ /*3119*/;
assign _56282_ = _55535_ ^ _56278_ /*3122*/;
assign _56283_ = _56274_ & _56282_ /*3120*/;
assign _55983_ = _56274_ ^ _56282_ /*3121*/;
assign _56280_ = _56281_ | _56283_ /*3118*/;
assign _56285_ = ~Q[1] /*3117*/;
assign _56284_ = _56285_ & D[47] /*3116*/;
assign _56287_ = _55536_ & _56284_ /*3111*/;
assign _56288_ = _55536_ ^ _56284_ /*3114*/;
assign _56289_ = _56280_ & _56288_ /*3112*/;
assign _55984_ = _56280_ ^ _56288_ /*3113*/;
assign _56286_ = _56287_ | _56289_ /*3110*/;
assign _56291_ = ~Q[1] /*3109*/;
assign _56290_ = _56291_ & D[48] /*3108*/;
assign _56293_ = _55537_ & _56290_ /*3103*/;
assign _56294_ = _55537_ ^ _56290_ /*3106*/;
assign _56295_ = _56286_ & _56294_ /*3104*/;
assign _55985_ = _56286_ ^ _56294_ /*3105*/;
assign _56292_ = _56293_ | _56295_ /*3102*/;
assign _56297_ = ~Q[1] /*3101*/;
assign _56296_ = _56297_ & D[49] /*3100*/;
assign _56299_ = _55538_ & _56296_ /*3095*/;
assign _56300_ = _55538_ ^ _56296_ /*3098*/;
assign _56301_ = _56292_ & _56300_ /*3096*/;
assign _55986_ = _56292_ ^ _56300_ /*3097*/;
assign _56298_ = _56299_ | _56301_ /*3094*/;
assign _56303_ = ~Q[1] /*3093*/;
assign _56302_ = _56303_ & D[50] /*3092*/;
assign _56305_ = _55539_ & _56302_ /*3087*/;
assign _56306_ = _55539_ ^ _56302_ /*3090*/;
assign _56307_ = _56298_ & _56306_ /*3088*/;
assign _55987_ = _56298_ ^ _56306_ /*3089*/;
assign _56304_ = _56305_ | _56307_ /*3086*/;
assign _56309_ = ~Q[1] /*3085*/;
assign _56308_ = _56309_ & D[51] /*3084*/;
assign _56311_ = _55540_ & _56308_ /*3079*/;
assign _56312_ = _55540_ ^ _56308_ /*3082*/;
assign _56313_ = _56304_ & _56312_ /*3080*/;
assign _55988_ = _56304_ ^ _56312_ /*3081*/;
assign _56310_ = _56311_ | _56313_ /*3078*/;
assign _56315_ = ~Q[1] /*3077*/;
assign _56314_ = _56315_ & D[52] /*3076*/;
assign _56317_ = _55541_ & _56314_ /*3071*/;
assign _56318_ = _55541_ ^ _56314_ /*3074*/;
assign _56319_ = _56310_ & _56318_ /*3072*/;
assign _55989_ = _56310_ ^ _56318_ /*3073*/;
assign _56316_ = _56317_ | _56319_ /*3070*/;
assign _56321_ = ~Q[1] /*3069*/;
assign _56320_ = _56321_ & D[53] /*3068*/;
assign _56323_ = _55542_ & _56320_ /*3063*/;
assign _56324_ = _55542_ ^ _56320_ /*3066*/;
assign _56325_ = _56316_ & _56324_ /*3064*/;
assign _55990_ = _56316_ ^ _56324_ /*3065*/;
assign _56322_ = _56323_ | _56325_ /*3062*/;
assign _56327_ = ~Q[1] /*3061*/;
assign _56326_ = _56327_ & D[54] /*3060*/;
assign _56329_ = _55543_ & _56326_ /*3055*/;
assign _56330_ = _55543_ ^ _56326_ /*3058*/;
assign _56331_ = _56322_ & _56330_ /*3056*/;
assign _55991_ = _56322_ ^ _56330_ /*3057*/;
assign _56328_ = _56329_ | _56331_ /*3054*/;
assign _56333_ = ~Q[1] /*3053*/;
assign _56332_ = _56333_ & D[55] /*3052*/;
assign _56335_ = _55544_ & _56332_ /*3047*/;
assign _56336_ = _55544_ ^ _56332_ /*3050*/;
assign _56337_ = _56328_ & _56336_ /*3048*/;
assign _55992_ = _56328_ ^ _56336_ /*3049*/;
assign _56334_ = _56335_ | _56337_ /*3046*/;
assign _56339_ = ~Q[1] /*3045*/;
assign _56338_ = _56339_ & D[56] /*3044*/;
assign _56341_ = _55545_ & _56338_ /*3039*/;
assign _56342_ = _55545_ ^ _56338_ /*3042*/;
assign _56343_ = _56334_ & _56342_ /*3040*/;
assign _55993_ = _56334_ ^ _56342_ /*3041*/;
assign _56340_ = _56341_ | _56343_ /*3038*/;
assign _56345_ = ~Q[1] /*3037*/;
assign _56344_ = _56345_ & D[57] /*3036*/;
assign _56347_ = _55546_ & _56344_ /*3031*/;
assign _56348_ = _55546_ ^ _56344_ /*3034*/;
assign _56349_ = _56340_ & _56348_ /*3032*/;
assign _55994_ = _56340_ ^ _56348_ /*3033*/;
assign _56346_ = _56347_ | _56349_ /*3030*/;
assign _56351_ = ~Q[1] /*3029*/;
assign _56350_ = _56351_ & D[58] /*3028*/;
assign _56353_ = _55547_ & _56350_ /*3023*/;
assign _56354_ = _55547_ ^ _56350_ /*3026*/;
assign _56355_ = _56346_ & _56354_ /*3024*/;
assign _55995_ = _56346_ ^ _56354_ /*3025*/;
assign _56352_ = _56353_ | _56355_ /*3022*/;
assign _56357_ = ~Q[1] /*3021*/;
assign _56356_ = _56357_ & D[59] /*3020*/;
assign _56359_ = _55548_ & _56356_ /*3015*/;
assign _56360_ = _55548_ ^ _56356_ /*3018*/;
assign _56361_ = _56352_ & _56360_ /*3016*/;
assign _55996_ = _56352_ ^ _56360_ /*3017*/;
assign _56358_ = _56359_ | _56361_ /*3014*/;
assign _56363_ = ~Q[1] /*3013*/;
assign _56362_ = _56363_ & D[60] /*3012*/;
assign _56365_ = _55549_ & _56362_ /*3007*/;
assign _56366_ = _55549_ ^ _56362_ /*3010*/;
assign _56367_ = _56358_ & _56366_ /*3008*/;
assign _55997_ = _56358_ ^ _56366_ /*3009*/;
assign _56364_ = _56365_ | _56367_ /*3006*/;
assign _56369_ = ~Q[1] /*3005*/;
assign _56368_ = _56369_ & D[61] /*3004*/;
assign _56371_ = _55550_ & _56368_ /*2999*/;
assign _56372_ = _55550_ ^ _56368_ /*3002*/;
assign _56373_ = _56364_ & _56372_ /*3000*/;
assign _55998_ = _56364_ ^ _56372_ /*3001*/;
assign _56370_ = _56371_ | _56373_ /*2998*/;
assign _56375_ = ~Q[1] /*2997*/;
assign _56374_ = _56375_ & D[62] /*2996*/;
assign _56377_ = _55551_ & _56374_ /*2991*/;
assign _56378_ = _55551_ ^ _56374_ /*2994*/;
assign _56379_ = _56370_ & _56378_ /*2992*/;
assign _55999_ = _56370_ ^ _56378_ /*2993*/;
assign _56376_ = _56377_ | _56379_ /*2990*/;
assign _56381_ = ~Q[1] /*2989*/;
assign _56380_ = _56381_ & zeroWire /*2988*/;
assign _56382_ = _55552_ ^ _56380_ /*2986*/;
assign _56000_ = _56382_ ^ _56376_ /*2985*/;
assign _56453_ = ~D[0] /*2731*/;
assign _56450_ = R_0[0] & _56453_ /*2727*/;
assign _56451_ = R_0[0] ^ _56453_ /*2730*/;
assign _56452_ = oneWire & _56451_ /*2728*/;
assign _56385_ = oneWire ^ _56451_ /*2729*/;
assign _56449_ = _56450_ | _56452_ /*2726*/;
assign _56458_ = ~D[1] /*2725*/;
assign _56455_ = _55937_ & _56458_ /*2721*/;
assign _56456_ = _55937_ ^ _56458_ /*2724*/;
assign _56457_ = _56449_ & _56456_ /*2722*/;
assign _56386_ = _56449_ ^ _56456_ /*2723*/;
assign _56454_ = _56455_ | _56457_ /*2720*/;
assign _56463_ = ~D[2] /*2719*/;
assign _56460_ = _55938_ & _56463_ /*2715*/;
assign _56461_ = _55938_ ^ _56463_ /*2718*/;
assign _56462_ = _56454_ & _56461_ /*2716*/;
assign _56387_ = _56454_ ^ _56461_ /*2717*/;
assign _56459_ = _56460_ | _56462_ /*2714*/;
assign _56468_ = ~D[3] /*2713*/;
assign _56465_ = _55939_ & _56468_ /*2709*/;
assign _56466_ = _55939_ ^ _56468_ /*2712*/;
assign _56467_ = _56459_ & _56466_ /*2710*/;
assign _56388_ = _56459_ ^ _56466_ /*2711*/;
assign _56464_ = _56465_ | _56467_ /*2708*/;
assign _56473_ = ~D[4] /*2707*/;
assign _56470_ = _55940_ & _56473_ /*2703*/;
assign _56471_ = _55940_ ^ _56473_ /*2706*/;
assign _56472_ = _56464_ & _56471_ /*2704*/;
assign _56389_ = _56464_ ^ _56471_ /*2705*/;
assign _56469_ = _56470_ | _56472_ /*2702*/;
assign _56478_ = ~D[5] /*2701*/;
assign _56475_ = _55941_ & _56478_ /*2697*/;
assign _56476_ = _55941_ ^ _56478_ /*2700*/;
assign _56477_ = _56469_ & _56476_ /*2698*/;
assign _56390_ = _56469_ ^ _56476_ /*2699*/;
assign _56474_ = _56475_ | _56477_ /*2696*/;
assign _56483_ = ~D[6] /*2695*/;
assign _56480_ = _55942_ & _56483_ /*2691*/;
assign _56481_ = _55942_ ^ _56483_ /*2694*/;
assign _56482_ = _56474_ & _56481_ /*2692*/;
assign _56391_ = _56474_ ^ _56481_ /*2693*/;
assign _56479_ = _56480_ | _56482_ /*2690*/;
assign _56488_ = ~D[7] /*2689*/;
assign _56485_ = _55943_ & _56488_ /*2685*/;
assign _56486_ = _55943_ ^ _56488_ /*2688*/;
assign _56487_ = _56479_ & _56486_ /*2686*/;
assign _56392_ = _56479_ ^ _56486_ /*2687*/;
assign _56484_ = _56485_ | _56487_ /*2684*/;
assign _56493_ = ~D[8] /*2683*/;
assign _56490_ = _55944_ & _56493_ /*2679*/;
assign _56491_ = _55944_ ^ _56493_ /*2682*/;
assign _56492_ = _56484_ & _56491_ /*2680*/;
assign _56393_ = _56484_ ^ _56491_ /*2681*/;
assign _56489_ = _56490_ | _56492_ /*2678*/;
assign _56498_ = ~D[9] /*2677*/;
assign _56495_ = _55945_ & _56498_ /*2673*/;
assign _56496_ = _55945_ ^ _56498_ /*2676*/;
assign _56497_ = _56489_ & _56496_ /*2674*/;
assign _56394_ = _56489_ ^ _56496_ /*2675*/;
assign _56494_ = _56495_ | _56497_ /*2672*/;
assign _56503_ = ~D[10] /*2671*/;
assign _56500_ = _55946_ & _56503_ /*2667*/;
assign _56501_ = _55946_ ^ _56503_ /*2670*/;
assign _56502_ = _56494_ & _56501_ /*2668*/;
assign _56395_ = _56494_ ^ _56501_ /*2669*/;
assign _56499_ = _56500_ | _56502_ /*2666*/;
assign _56508_ = ~D[11] /*2665*/;
assign _56505_ = _55947_ & _56508_ /*2661*/;
assign _56506_ = _55947_ ^ _56508_ /*2664*/;
assign _56507_ = _56499_ & _56506_ /*2662*/;
assign _56396_ = _56499_ ^ _56506_ /*2663*/;
assign _56504_ = _56505_ | _56507_ /*2660*/;
assign _56513_ = ~D[12] /*2659*/;
assign _56510_ = _55948_ & _56513_ /*2655*/;
assign _56511_ = _55948_ ^ _56513_ /*2658*/;
assign _56512_ = _56504_ & _56511_ /*2656*/;
assign _56397_ = _56504_ ^ _56511_ /*2657*/;
assign _56509_ = _56510_ | _56512_ /*2654*/;
assign _56518_ = ~D[13] /*2653*/;
assign _56515_ = _55949_ & _56518_ /*2649*/;
assign _56516_ = _55949_ ^ _56518_ /*2652*/;
assign _56517_ = _56509_ & _56516_ /*2650*/;
assign _56398_ = _56509_ ^ _56516_ /*2651*/;
assign _56514_ = _56515_ | _56517_ /*2648*/;
assign _56523_ = ~D[14] /*2647*/;
assign _56520_ = _55950_ & _56523_ /*2643*/;
assign _56521_ = _55950_ ^ _56523_ /*2646*/;
assign _56522_ = _56514_ & _56521_ /*2644*/;
assign _56399_ = _56514_ ^ _56521_ /*2645*/;
assign _56519_ = _56520_ | _56522_ /*2642*/;
assign _56528_ = ~D[15] /*2641*/;
assign _56525_ = _55951_ & _56528_ /*2637*/;
assign _56526_ = _55951_ ^ _56528_ /*2640*/;
assign _56527_ = _56519_ & _56526_ /*2638*/;
assign _56400_ = _56519_ ^ _56526_ /*2639*/;
assign _56524_ = _56525_ | _56527_ /*2636*/;
assign _56533_ = ~D[16] /*2635*/;
assign _56530_ = _55952_ & _56533_ /*2631*/;
assign _56531_ = _55952_ ^ _56533_ /*2634*/;
assign _56532_ = _56524_ & _56531_ /*2632*/;
assign _56401_ = _56524_ ^ _56531_ /*2633*/;
assign _56529_ = _56530_ | _56532_ /*2630*/;
assign _56538_ = ~D[17] /*2629*/;
assign _56535_ = _55953_ & _56538_ /*2625*/;
assign _56536_ = _55953_ ^ _56538_ /*2628*/;
assign _56537_ = _56529_ & _56536_ /*2626*/;
assign _56402_ = _56529_ ^ _56536_ /*2627*/;
assign _56534_ = _56535_ | _56537_ /*2624*/;
assign _56543_ = ~D[18] /*2623*/;
assign _56540_ = _55954_ & _56543_ /*2619*/;
assign _56541_ = _55954_ ^ _56543_ /*2622*/;
assign _56542_ = _56534_ & _56541_ /*2620*/;
assign _56403_ = _56534_ ^ _56541_ /*2621*/;
assign _56539_ = _56540_ | _56542_ /*2618*/;
assign _56548_ = ~D[19] /*2617*/;
assign _56545_ = _55955_ & _56548_ /*2613*/;
assign _56546_ = _55955_ ^ _56548_ /*2616*/;
assign _56547_ = _56539_ & _56546_ /*2614*/;
assign _56404_ = _56539_ ^ _56546_ /*2615*/;
assign _56544_ = _56545_ | _56547_ /*2612*/;
assign _56553_ = ~D[20] /*2611*/;
assign _56550_ = _55956_ & _56553_ /*2607*/;
assign _56551_ = _55956_ ^ _56553_ /*2610*/;
assign _56552_ = _56544_ & _56551_ /*2608*/;
assign _56405_ = _56544_ ^ _56551_ /*2609*/;
assign _56549_ = _56550_ | _56552_ /*2606*/;
assign _56558_ = ~D[21] /*2605*/;
assign _56555_ = _55957_ & _56558_ /*2601*/;
assign _56556_ = _55957_ ^ _56558_ /*2604*/;
assign _56557_ = _56549_ & _56556_ /*2602*/;
assign _56406_ = _56549_ ^ _56556_ /*2603*/;
assign _56554_ = _56555_ | _56557_ /*2600*/;
assign _56563_ = ~D[22] /*2599*/;
assign _56560_ = _55958_ & _56563_ /*2595*/;
assign _56561_ = _55958_ ^ _56563_ /*2598*/;
assign _56562_ = _56554_ & _56561_ /*2596*/;
assign _56407_ = _56554_ ^ _56561_ /*2597*/;
assign _56559_ = _56560_ | _56562_ /*2594*/;
assign _56568_ = ~D[23] /*2593*/;
assign _56565_ = _55959_ & _56568_ /*2589*/;
assign _56566_ = _55959_ ^ _56568_ /*2592*/;
assign _56567_ = _56559_ & _56566_ /*2590*/;
assign _56408_ = _56559_ ^ _56566_ /*2591*/;
assign _56564_ = _56565_ | _56567_ /*2588*/;
assign _56573_ = ~D[24] /*2587*/;
assign _56570_ = _55960_ & _56573_ /*2583*/;
assign _56571_ = _55960_ ^ _56573_ /*2586*/;
assign _56572_ = _56564_ & _56571_ /*2584*/;
assign _56409_ = _56564_ ^ _56571_ /*2585*/;
assign _56569_ = _56570_ | _56572_ /*2582*/;
assign _56578_ = ~D[25] /*2581*/;
assign _56575_ = _55961_ & _56578_ /*2577*/;
assign _56576_ = _55961_ ^ _56578_ /*2580*/;
assign _56577_ = _56569_ & _56576_ /*2578*/;
assign _56410_ = _56569_ ^ _56576_ /*2579*/;
assign _56574_ = _56575_ | _56577_ /*2576*/;
assign _56583_ = ~D[26] /*2575*/;
assign _56580_ = _55962_ & _56583_ /*2571*/;
assign _56581_ = _55962_ ^ _56583_ /*2574*/;
assign _56582_ = _56574_ & _56581_ /*2572*/;
assign _56411_ = _56574_ ^ _56581_ /*2573*/;
assign _56579_ = _56580_ | _56582_ /*2570*/;
assign _56588_ = ~D[27] /*2569*/;
assign _56585_ = _55963_ & _56588_ /*2565*/;
assign _56586_ = _55963_ ^ _56588_ /*2568*/;
assign _56587_ = _56579_ & _56586_ /*2566*/;
assign _56412_ = _56579_ ^ _56586_ /*2567*/;
assign _56584_ = _56585_ | _56587_ /*2564*/;
assign _56593_ = ~D[28] /*2563*/;
assign _56590_ = _55964_ & _56593_ /*2559*/;
assign _56591_ = _55964_ ^ _56593_ /*2562*/;
assign _56592_ = _56584_ & _56591_ /*2560*/;
assign _56413_ = _56584_ ^ _56591_ /*2561*/;
assign _56589_ = _56590_ | _56592_ /*2558*/;
assign _56598_ = ~D[29] /*2557*/;
assign _56595_ = _55965_ & _56598_ /*2553*/;
assign _56596_ = _55965_ ^ _56598_ /*2556*/;
assign _56597_ = _56589_ & _56596_ /*2554*/;
assign _56414_ = _56589_ ^ _56596_ /*2555*/;
assign _56594_ = _56595_ | _56597_ /*2552*/;
assign _56603_ = ~D[30] /*2551*/;
assign _56600_ = _55966_ & _56603_ /*2547*/;
assign _56601_ = _55966_ ^ _56603_ /*2550*/;
assign _56602_ = _56594_ & _56601_ /*2548*/;
assign _56415_ = _56594_ ^ _56601_ /*2549*/;
assign _56599_ = _56600_ | _56602_ /*2546*/;
assign _56608_ = ~D[31] /*2545*/;
assign _56605_ = _55967_ & _56608_ /*2541*/;
assign _56606_ = _55967_ ^ _56608_ /*2544*/;
assign _56607_ = _56599_ & _56606_ /*2542*/;
assign _56416_ = _56599_ ^ _56606_ /*2543*/;
assign _56604_ = _56605_ | _56607_ /*2540*/;
assign _56613_ = ~D[32] /*2539*/;
assign _56610_ = _55968_ & _56613_ /*2535*/;
assign _56611_ = _55968_ ^ _56613_ /*2538*/;
assign _56612_ = _56604_ & _56611_ /*2536*/;
assign _56417_ = _56604_ ^ _56611_ /*2537*/;
assign _56609_ = _56610_ | _56612_ /*2534*/;
assign _56618_ = ~D[33] /*2533*/;
assign _56615_ = _55969_ & _56618_ /*2529*/;
assign _56616_ = _55969_ ^ _56618_ /*2532*/;
assign _56617_ = _56609_ & _56616_ /*2530*/;
assign _56418_ = _56609_ ^ _56616_ /*2531*/;
assign _56614_ = _56615_ | _56617_ /*2528*/;
assign _56623_ = ~D[34] /*2527*/;
assign _56620_ = _55970_ & _56623_ /*2523*/;
assign _56621_ = _55970_ ^ _56623_ /*2526*/;
assign _56622_ = _56614_ & _56621_ /*2524*/;
assign _56419_ = _56614_ ^ _56621_ /*2525*/;
assign _56619_ = _56620_ | _56622_ /*2522*/;
assign _56628_ = ~D[35] /*2521*/;
assign _56625_ = _55971_ & _56628_ /*2517*/;
assign _56626_ = _55971_ ^ _56628_ /*2520*/;
assign _56627_ = _56619_ & _56626_ /*2518*/;
assign _56420_ = _56619_ ^ _56626_ /*2519*/;
assign _56624_ = _56625_ | _56627_ /*2516*/;
assign _56633_ = ~D[36] /*2515*/;
assign _56630_ = _55972_ & _56633_ /*2511*/;
assign _56631_ = _55972_ ^ _56633_ /*2514*/;
assign _56632_ = _56624_ & _56631_ /*2512*/;
assign _56421_ = _56624_ ^ _56631_ /*2513*/;
assign _56629_ = _56630_ | _56632_ /*2510*/;
assign _56638_ = ~D[37] /*2509*/;
assign _56635_ = _55973_ & _56638_ /*2505*/;
assign _56636_ = _55973_ ^ _56638_ /*2508*/;
assign _56637_ = _56629_ & _56636_ /*2506*/;
assign _56422_ = _56629_ ^ _56636_ /*2507*/;
assign _56634_ = _56635_ | _56637_ /*2504*/;
assign _56643_ = ~D[38] /*2503*/;
assign _56640_ = _55974_ & _56643_ /*2499*/;
assign _56641_ = _55974_ ^ _56643_ /*2502*/;
assign _56642_ = _56634_ & _56641_ /*2500*/;
assign _56423_ = _56634_ ^ _56641_ /*2501*/;
assign _56639_ = _56640_ | _56642_ /*2498*/;
assign _56648_ = ~D[39] /*2497*/;
assign _56645_ = _55975_ & _56648_ /*2493*/;
assign _56646_ = _55975_ ^ _56648_ /*2496*/;
assign _56647_ = _56639_ & _56646_ /*2494*/;
assign _56424_ = _56639_ ^ _56646_ /*2495*/;
assign _56644_ = _56645_ | _56647_ /*2492*/;
assign _56653_ = ~D[40] /*2491*/;
assign _56650_ = _55976_ & _56653_ /*2487*/;
assign _56651_ = _55976_ ^ _56653_ /*2490*/;
assign _56652_ = _56644_ & _56651_ /*2488*/;
assign _56425_ = _56644_ ^ _56651_ /*2489*/;
assign _56649_ = _56650_ | _56652_ /*2486*/;
assign _56658_ = ~D[41] /*2485*/;
assign _56655_ = _55977_ & _56658_ /*2481*/;
assign _56656_ = _55977_ ^ _56658_ /*2484*/;
assign _56657_ = _56649_ & _56656_ /*2482*/;
assign _56426_ = _56649_ ^ _56656_ /*2483*/;
assign _56654_ = _56655_ | _56657_ /*2480*/;
assign _56663_ = ~D[42] /*2479*/;
assign _56660_ = _55978_ & _56663_ /*2475*/;
assign _56661_ = _55978_ ^ _56663_ /*2478*/;
assign _56662_ = _56654_ & _56661_ /*2476*/;
assign _56427_ = _56654_ ^ _56661_ /*2477*/;
assign _56659_ = _56660_ | _56662_ /*2474*/;
assign _56668_ = ~D[43] /*2473*/;
assign _56665_ = _55979_ & _56668_ /*2469*/;
assign _56666_ = _55979_ ^ _56668_ /*2472*/;
assign _56667_ = _56659_ & _56666_ /*2470*/;
assign _56428_ = _56659_ ^ _56666_ /*2471*/;
assign _56664_ = _56665_ | _56667_ /*2468*/;
assign _56673_ = ~D[44] /*2467*/;
assign _56670_ = _55980_ & _56673_ /*2463*/;
assign _56671_ = _55980_ ^ _56673_ /*2466*/;
assign _56672_ = _56664_ & _56671_ /*2464*/;
assign _56429_ = _56664_ ^ _56671_ /*2465*/;
assign _56669_ = _56670_ | _56672_ /*2462*/;
assign _56678_ = ~D[45] /*2461*/;
assign _56675_ = _55981_ & _56678_ /*2457*/;
assign _56676_ = _55981_ ^ _56678_ /*2460*/;
assign _56677_ = _56669_ & _56676_ /*2458*/;
assign _56430_ = _56669_ ^ _56676_ /*2459*/;
assign _56674_ = _56675_ | _56677_ /*2456*/;
assign _56683_ = ~D[46] /*2455*/;
assign _56680_ = _55982_ & _56683_ /*2451*/;
assign _56681_ = _55982_ ^ _56683_ /*2454*/;
assign _56682_ = _56674_ & _56681_ /*2452*/;
assign _56431_ = _56674_ ^ _56681_ /*2453*/;
assign _56679_ = _56680_ | _56682_ /*2450*/;
assign _56688_ = ~D[47] /*2449*/;
assign _56685_ = _55983_ & _56688_ /*2445*/;
assign _56686_ = _55983_ ^ _56688_ /*2448*/;
assign _56687_ = _56679_ & _56686_ /*2446*/;
assign _56432_ = _56679_ ^ _56686_ /*2447*/;
assign _56684_ = _56685_ | _56687_ /*2444*/;
assign _56693_ = ~D[48] /*2443*/;
assign _56690_ = _55984_ & _56693_ /*2439*/;
assign _56691_ = _55984_ ^ _56693_ /*2442*/;
assign _56692_ = _56684_ & _56691_ /*2440*/;
assign _56433_ = _56684_ ^ _56691_ /*2441*/;
assign _56689_ = _56690_ | _56692_ /*2438*/;
assign _56698_ = ~D[49] /*2437*/;
assign _56695_ = _55985_ & _56698_ /*2433*/;
assign _56696_ = _55985_ ^ _56698_ /*2436*/;
assign _56697_ = _56689_ & _56696_ /*2434*/;
assign _56434_ = _56689_ ^ _56696_ /*2435*/;
assign _56694_ = _56695_ | _56697_ /*2432*/;
assign _56703_ = ~D[50] /*2431*/;
assign _56700_ = _55986_ & _56703_ /*2427*/;
assign _56701_ = _55986_ ^ _56703_ /*2430*/;
assign _56702_ = _56694_ & _56701_ /*2428*/;
assign _56435_ = _56694_ ^ _56701_ /*2429*/;
assign _56699_ = _56700_ | _56702_ /*2426*/;
assign _56708_ = ~D[51] /*2425*/;
assign _56705_ = _55987_ & _56708_ /*2421*/;
assign _56706_ = _55987_ ^ _56708_ /*2424*/;
assign _56707_ = _56699_ & _56706_ /*2422*/;
assign _56436_ = _56699_ ^ _56706_ /*2423*/;
assign _56704_ = _56705_ | _56707_ /*2420*/;
assign _56713_ = ~D[52] /*2419*/;
assign _56710_ = _55988_ & _56713_ /*2415*/;
assign _56711_ = _55988_ ^ _56713_ /*2418*/;
assign _56712_ = _56704_ & _56711_ /*2416*/;
assign _56437_ = _56704_ ^ _56711_ /*2417*/;
assign _56709_ = _56710_ | _56712_ /*2414*/;
assign _56718_ = ~D[53] /*2413*/;
assign _56715_ = _55989_ & _56718_ /*2409*/;
assign _56716_ = _55989_ ^ _56718_ /*2412*/;
assign _56717_ = _56709_ & _56716_ /*2410*/;
assign _56438_ = _56709_ ^ _56716_ /*2411*/;
assign _56714_ = _56715_ | _56717_ /*2408*/;
assign _56723_ = ~D[54] /*2407*/;
assign _56720_ = _55990_ & _56723_ /*2403*/;
assign _56721_ = _55990_ ^ _56723_ /*2406*/;
assign _56722_ = _56714_ & _56721_ /*2404*/;
assign _56439_ = _56714_ ^ _56721_ /*2405*/;
assign _56719_ = _56720_ | _56722_ /*2402*/;
assign _56728_ = ~D[55] /*2401*/;
assign _56725_ = _55991_ & _56728_ /*2397*/;
assign _56726_ = _55991_ ^ _56728_ /*2400*/;
assign _56727_ = _56719_ & _56726_ /*2398*/;
assign _56440_ = _56719_ ^ _56726_ /*2399*/;
assign _56724_ = _56725_ | _56727_ /*2396*/;
assign _56733_ = ~D[56] /*2395*/;
assign _56730_ = _55992_ & _56733_ /*2391*/;
assign _56731_ = _55992_ ^ _56733_ /*2394*/;
assign _56732_ = _56724_ & _56731_ /*2392*/;
assign _56441_ = _56724_ ^ _56731_ /*2393*/;
assign _56729_ = _56730_ | _56732_ /*2390*/;
assign _56738_ = ~D[57] /*2389*/;
assign _56735_ = _55993_ & _56738_ /*2385*/;
assign _56736_ = _55993_ ^ _56738_ /*2388*/;
assign _56737_ = _56729_ & _56736_ /*2386*/;
assign _56442_ = _56729_ ^ _56736_ /*2387*/;
assign _56734_ = _56735_ | _56737_ /*2384*/;
assign _56743_ = ~D[58] /*2383*/;
assign _56740_ = _55994_ & _56743_ /*2379*/;
assign _56741_ = _55994_ ^ _56743_ /*2382*/;
assign _56742_ = _56734_ & _56741_ /*2380*/;
assign _56443_ = _56734_ ^ _56741_ /*2381*/;
assign _56739_ = _56740_ | _56742_ /*2378*/;
assign _56748_ = ~D[59] /*2377*/;
assign _56745_ = _55995_ & _56748_ /*2373*/;
assign _56746_ = _55995_ ^ _56748_ /*2376*/;
assign _56747_ = _56739_ & _56746_ /*2374*/;
assign _56444_ = _56739_ ^ _56746_ /*2375*/;
assign _56744_ = _56745_ | _56747_ /*2372*/;
assign _56753_ = ~D[60] /*2371*/;
assign _56750_ = _55996_ & _56753_ /*2367*/;
assign _56751_ = _55996_ ^ _56753_ /*2370*/;
assign _56752_ = _56744_ & _56751_ /*2368*/;
assign _56445_ = _56744_ ^ _56751_ /*2369*/;
assign _56749_ = _56750_ | _56752_ /*2366*/;
assign _56758_ = ~D[61] /*2365*/;
assign _56755_ = _55997_ & _56758_ /*2361*/;
assign _56756_ = _55997_ ^ _56758_ /*2364*/;
assign _56757_ = _56749_ & _56756_ /*2362*/;
assign _56446_ = _56749_ ^ _56756_ /*2363*/;
assign _56754_ = _56755_ | _56757_ /*2360*/;
assign _56763_ = ~D[62] /*2359*/;
assign _56760_ = _55998_ & _56763_ /*2355*/;
assign _56761_ = _55998_ ^ _56763_ /*2358*/;
assign _56762_ = _56754_ & _56761_ /*2356*/;
assign _56447_ = _56754_ ^ _56761_ /*2357*/;
assign _56759_ = _56760_ | _56762_ /*2354*/;
assign _56764_ = _55999_ & oneWire /*2349*/;
assign _56765_ = _55999_ ^ oneWire /*2352*/;
assign _56766_ = _56759_ & _56765_ /*2350*/;
assign _56448_ = _56759_ ^ _56765_ /*2351*/;
assign Q[0] = _56764_ | _56766_ /*2348*/;
assign _56899_ = ~Q[0] /*1963*/;
assign _56898_ = _56899_ & D[0] /*1962*/;
assign _56901_ = _56385_ & _56898_ /*1957*/;
assign _56902_ = _56385_ ^ _56898_ /*1960*/;
assign _56903_ = zeroWire & _56902_ /*1958*/;
assign R_n1[0] = zeroWire ^ _56902_ /*1959*/;
assign _56900_ = _56901_ | _56903_ /*1956*/;
assign _56905_ = ~Q[0] /*1955*/;
assign _56904_ = _56905_ & D[1] /*1954*/;
assign _56907_ = _56386_ & _56904_ /*1949*/;
assign _56908_ = _56386_ ^ _56904_ /*1952*/;
assign _56909_ = _56900_ & _56908_ /*1950*/;
assign R_n1[1] = _56900_ ^ _56908_ /*1951*/;
assign _56906_ = _56907_ | _56909_ /*1948*/;
assign _56911_ = ~Q[0] /*1947*/;
assign _56910_ = _56911_ & D[2] /*1946*/;
assign _56913_ = _56387_ & _56910_ /*1941*/;
assign _56914_ = _56387_ ^ _56910_ /*1944*/;
assign _56915_ = _56906_ & _56914_ /*1942*/;
assign R_n1[2] = _56906_ ^ _56914_ /*1943*/;
assign _56912_ = _56913_ | _56915_ /*1940*/;
assign _56917_ = ~Q[0] /*1939*/;
assign _56916_ = _56917_ & D[3] /*1938*/;
assign _56919_ = _56388_ & _56916_ /*1933*/;
assign _56920_ = _56388_ ^ _56916_ /*1936*/;
assign _56921_ = _56912_ & _56920_ /*1934*/;
assign R_n1[3] = _56912_ ^ _56920_ /*1935*/;
assign _56918_ = _56919_ | _56921_ /*1932*/;
assign _56923_ = ~Q[0] /*1931*/;
assign _56922_ = _56923_ & D[4] /*1930*/;
assign _56925_ = _56389_ & _56922_ /*1925*/;
assign _56926_ = _56389_ ^ _56922_ /*1928*/;
assign _56927_ = _56918_ & _56926_ /*1926*/;
assign R_n1[4] = _56918_ ^ _56926_ /*1927*/;
assign _56924_ = _56925_ | _56927_ /*1924*/;
assign _56929_ = ~Q[0] /*1923*/;
assign _56928_ = _56929_ & D[5] /*1922*/;
assign _56931_ = _56390_ & _56928_ /*1917*/;
assign _56932_ = _56390_ ^ _56928_ /*1920*/;
assign _56933_ = _56924_ & _56932_ /*1918*/;
assign R_n1[5] = _56924_ ^ _56932_ /*1919*/;
assign _56930_ = _56931_ | _56933_ /*1916*/;
assign _56935_ = ~Q[0] /*1915*/;
assign _56934_ = _56935_ & D[6] /*1914*/;
assign _56937_ = _56391_ & _56934_ /*1909*/;
assign _56938_ = _56391_ ^ _56934_ /*1912*/;
assign _56939_ = _56930_ & _56938_ /*1910*/;
assign R_n1[6] = _56930_ ^ _56938_ /*1911*/;
assign _56936_ = _56937_ | _56939_ /*1908*/;
assign _56941_ = ~Q[0] /*1907*/;
assign _56940_ = _56941_ & D[7] /*1906*/;
assign _56943_ = _56392_ & _56940_ /*1901*/;
assign _56944_ = _56392_ ^ _56940_ /*1904*/;
assign _56945_ = _56936_ & _56944_ /*1902*/;
assign R_n1[7] = _56936_ ^ _56944_ /*1903*/;
assign _56942_ = _56943_ | _56945_ /*1900*/;
assign _56947_ = ~Q[0] /*1899*/;
assign _56946_ = _56947_ & D[8] /*1898*/;
assign _56949_ = _56393_ & _56946_ /*1893*/;
assign _56950_ = _56393_ ^ _56946_ /*1896*/;
assign _56951_ = _56942_ & _56950_ /*1894*/;
assign R_n1[8] = _56942_ ^ _56950_ /*1895*/;
assign _56948_ = _56949_ | _56951_ /*1892*/;
assign _56953_ = ~Q[0] /*1891*/;
assign _56952_ = _56953_ & D[9] /*1890*/;
assign _56955_ = _56394_ & _56952_ /*1885*/;
assign _56956_ = _56394_ ^ _56952_ /*1888*/;
assign _56957_ = _56948_ & _56956_ /*1886*/;
assign R_n1[9] = _56948_ ^ _56956_ /*1887*/;
assign _56954_ = _56955_ | _56957_ /*1884*/;
assign _56959_ = ~Q[0] /*1883*/;
assign _56958_ = _56959_ & D[10] /*1882*/;
assign _56961_ = _56395_ & _56958_ /*1877*/;
assign _56962_ = _56395_ ^ _56958_ /*1880*/;
assign _56963_ = _56954_ & _56962_ /*1878*/;
assign R_n1[10] = _56954_ ^ _56962_ /*1879*/;
assign _56960_ = _56961_ | _56963_ /*1876*/;
assign _56965_ = ~Q[0] /*1875*/;
assign _56964_ = _56965_ & D[11] /*1874*/;
assign _56967_ = _56396_ & _56964_ /*1869*/;
assign _56968_ = _56396_ ^ _56964_ /*1872*/;
assign _56969_ = _56960_ & _56968_ /*1870*/;
assign R_n1[11] = _56960_ ^ _56968_ /*1871*/;
assign _56966_ = _56967_ | _56969_ /*1868*/;
assign _56971_ = ~Q[0] /*1867*/;
assign _56970_ = _56971_ & D[12] /*1866*/;
assign _56973_ = _56397_ & _56970_ /*1861*/;
assign _56974_ = _56397_ ^ _56970_ /*1864*/;
assign _56975_ = _56966_ & _56974_ /*1862*/;
assign R_n1[12] = _56966_ ^ _56974_ /*1863*/;
assign _56972_ = _56973_ | _56975_ /*1860*/;
assign _56977_ = ~Q[0] /*1859*/;
assign _56976_ = _56977_ & D[13] /*1858*/;
assign _56979_ = _56398_ & _56976_ /*1853*/;
assign _56980_ = _56398_ ^ _56976_ /*1856*/;
assign _56981_ = _56972_ & _56980_ /*1854*/;
assign R_n1[13] = _56972_ ^ _56980_ /*1855*/;
assign _56978_ = _56979_ | _56981_ /*1852*/;
assign _56983_ = ~Q[0] /*1851*/;
assign _56982_ = _56983_ & D[14] /*1850*/;
assign _56985_ = _56399_ & _56982_ /*1845*/;
assign _56986_ = _56399_ ^ _56982_ /*1848*/;
assign _56987_ = _56978_ & _56986_ /*1846*/;
assign R_n1[14] = _56978_ ^ _56986_ /*1847*/;
assign _56984_ = _56985_ | _56987_ /*1844*/;
assign _56989_ = ~Q[0] /*1843*/;
assign _56988_ = _56989_ & D[15] /*1842*/;
assign _56991_ = _56400_ & _56988_ /*1837*/;
assign _56992_ = _56400_ ^ _56988_ /*1840*/;
assign _56993_ = _56984_ & _56992_ /*1838*/;
assign R_n1[15] = _56984_ ^ _56992_ /*1839*/;
assign _56990_ = _56991_ | _56993_ /*1836*/;
assign _56995_ = ~Q[0] /*1835*/;
assign _56994_ = _56995_ & D[16] /*1834*/;
assign _56997_ = _56401_ & _56994_ /*1829*/;
assign _56998_ = _56401_ ^ _56994_ /*1832*/;
assign _56999_ = _56990_ & _56998_ /*1830*/;
assign R_n1[16] = _56990_ ^ _56998_ /*1831*/;
assign _56996_ = _56997_ | _56999_ /*1828*/;
assign _57001_ = ~Q[0] /*1827*/;
assign _57000_ = _57001_ & D[17] /*1826*/;
assign _57003_ = _56402_ & _57000_ /*1821*/;
assign _57004_ = _56402_ ^ _57000_ /*1824*/;
assign _57005_ = _56996_ & _57004_ /*1822*/;
assign R_n1[17] = _56996_ ^ _57004_ /*1823*/;
assign _57002_ = _57003_ | _57005_ /*1820*/;
assign _57007_ = ~Q[0] /*1819*/;
assign _57006_ = _57007_ & D[18] /*1818*/;
assign _57009_ = _56403_ & _57006_ /*1813*/;
assign _57010_ = _56403_ ^ _57006_ /*1816*/;
assign _57011_ = _57002_ & _57010_ /*1814*/;
assign R_n1[18] = _57002_ ^ _57010_ /*1815*/;
assign _57008_ = _57009_ | _57011_ /*1812*/;
assign _57013_ = ~Q[0] /*1811*/;
assign _57012_ = _57013_ & D[19] /*1810*/;
assign _57015_ = _56404_ & _57012_ /*1805*/;
assign _57016_ = _56404_ ^ _57012_ /*1808*/;
assign _57017_ = _57008_ & _57016_ /*1806*/;
assign R_n1[19] = _57008_ ^ _57016_ /*1807*/;
assign _57014_ = _57015_ | _57017_ /*1804*/;
assign _57019_ = ~Q[0] /*1803*/;
assign _57018_ = _57019_ & D[20] /*1802*/;
assign _57021_ = _56405_ & _57018_ /*1797*/;
assign _57022_ = _56405_ ^ _57018_ /*1800*/;
assign _57023_ = _57014_ & _57022_ /*1798*/;
assign R_n1[20] = _57014_ ^ _57022_ /*1799*/;
assign _57020_ = _57021_ | _57023_ /*1796*/;
assign _57025_ = ~Q[0] /*1795*/;
assign _57024_ = _57025_ & D[21] /*1794*/;
assign _57027_ = _56406_ & _57024_ /*1789*/;
assign _57028_ = _56406_ ^ _57024_ /*1792*/;
assign _57029_ = _57020_ & _57028_ /*1790*/;
assign R_n1[21] = _57020_ ^ _57028_ /*1791*/;
assign _57026_ = _57027_ | _57029_ /*1788*/;
assign _57031_ = ~Q[0] /*1787*/;
assign _57030_ = _57031_ & D[22] /*1786*/;
assign _57033_ = _56407_ & _57030_ /*1781*/;
assign _57034_ = _56407_ ^ _57030_ /*1784*/;
assign _57035_ = _57026_ & _57034_ /*1782*/;
assign R_n1[22] = _57026_ ^ _57034_ /*1783*/;
assign _57032_ = _57033_ | _57035_ /*1780*/;
assign _57037_ = ~Q[0] /*1779*/;
assign _57036_ = _57037_ & D[23] /*1778*/;
assign _57039_ = _56408_ & _57036_ /*1773*/;
assign _57040_ = _56408_ ^ _57036_ /*1776*/;
assign _57041_ = _57032_ & _57040_ /*1774*/;
assign R_n1[23] = _57032_ ^ _57040_ /*1775*/;
assign _57038_ = _57039_ | _57041_ /*1772*/;
assign _57043_ = ~Q[0] /*1771*/;
assign _57042_ = _57043_ & D[24] /*1770*/;
assign _57045_ = _56409_ & _57042_ /*1765*/;
assign _57046_ = _56409_ ^ _57042_ /*1768*/;
assign _57047_ = _57038_ & _57046_ /*1766*/;
assign R_n1[24] = _57038_ ^ _57046_ /*1767*/;
assign _57044_ = _57045_ | _57047_ /*1764*/;
assign _57049_ = ~Q[0] /*1763*/;
assign _57048_ = _57049_ & D[25] /*1762*/;
assign _57051_ = _56410_ & _57048_ /*1757*/;
assign _57052_ = _56410_ ^ _57048_ /*1760*/;
assign _57053_ = _57044_ & _57052_ /*1758*/;
assign R_n1[25] = _57044_ ^ _57052_ /*1759*/;
assign _57050_ = _57051_ | _57053_ /*1756*/;
assign _57055_ = ~Q[0] /*1755*/;
assign _57054_ = _57055_ & D[26] /*1754*/;
assign _57057_ = _56411_ & _57054_ /*1749*/;
assign _57058_ = _56411_ ^ _57054_ /*1752*/;
assign _57059_ = _57050_ & _57058_ /*1750*/;
assign R_n1[26] = _57050_ ^ _57058_ /*1751*/;
assign _57056_ = _57057_ | _57059_ /*1748*/;
assign _57061_ = ~Q[0] /*1747*/;
assign _57060_ = _57061_ & D[27] /*1746*/;
assign _57063_ = _56412_ & _57060_ /*1741*/;
assign _57064_ = _56412_ ^ _57060_ /*1744*/;
assign _57065_ = _57056_ & _57064_ /*1742*/;
assign R_n1[27] = _57056_ ^ _57064_ /*1743*/;
assign _57062_ = _57063_ | _57065_ /*1740*/;
assign _57067_ = ~Q[0] /*1739*/;
assign _57066_ = _57067_ & D[28] /*1738*/;
assign _57069_ = _56413_ & _57066_ /*1733*/;
assign _57070_ = _56413_ ^ _57066_ /*1736*/;
assign _57071_ = _57062_ & _57070_ /*1734*/;
assign R_n1[28] = _57062_ ^ _57070_ /*1735*/;
assign _57068_ = _57069_ | _57071_ /*1732*/;
assign _57073_ = ~Q[0] /*1731*/;
assign _57072_ = _57073_ & D[29] /*1730*/;
assign _57075_ = _56414_ & _57072_ /*1725*/;
assign _57076_ = _56414_ ^ _57072_ /*1728*/;
assign _57077_ = _57068_ & _57076_ /*1726*/;
assign R_n1[29] = _57068_ ^ _57076_ /*1727*/;
assign _57074_ = _57075_ | _57077_ /*1724*/;
assign _57079_ = ~Q[0] /*1723*/;
assign _57078_ = _57079_ & D[30] /*1722*/;
assign _57081_ = _56415_ & _57078_ /*1717*/;
assign _57082_ = _56415_ ^ _57078_ /*1720*/;
assign _57083_ = _57074_ & _57082_ /*1718*/;
assign R_n1[30] = _57074_ ^ _57082_ /*1719*/;
assign _57080_ = _57081_ | _57083_ /*1716*/;
assign _57085_ = ~Q[0] /*1715*/;
assign _57084_ = _57085_ & D[31] /*1714*/;
assign _57087_ = _56416_ & _57084_ /*1709*/;
assign _57088_ = _56416_ ^ _57084_ /*1712*/;
assign _57089_ = _57080_ & _57088_ /*1710*/;
assign R_n1[31] = _57080_ ^ _57088_ /*1711*/;
assign _57086_ = _57087_ | _57089_ /*1708*/;
assign _57091_ = ~Q[0] /*1707*/;
assign _57090_ = _57091_ & D[32] /*1706*/;
assign _57093_ = _56417_ & _57090_ /*1701*/;
assign _57094_ = _56417_ ^ _57090_ /*1704*/;
assign _57095_ = _57086_ & _57094_ /*1702*/;
assign R_n1[32] = _57086_ ^ _57094_ /*1703*/;
assign _57092_ = _57093_ | _57095_ /*1700*/;
assign _57097_ = ~Q[0] /*1699*/;
assign _57096_ = _57097_ & D[33] /*1698*/;
assign _57099_ = _56418_ & _57096_ /*1693*/;
assign _57100_ = _56418_ ^ _57096_ /*1696*/;
assign _57101_ = _57092_ & _57100_ /*1694*/;
assign R_n1[33] = _57092_ ^ _57100_ /*1695*/;
assign _57098_ = _57099_ | _57101_ /*1692*/;
assign _57103_ = ~Q[0] /*1691*/;
assign _57102_ = _57103_ & D[34] /*1690*/;
assign _57105_ = _56419_ & _57102_ /*1685*/;
assign _57106_ = _56419_ ^ _57102_ /*1688*/;
assign _57107_ = _57098_ & _57106_ /*1686*/;
assign R_n1[34] = _57098_ ^ _57106_ /*1687*/;
assign _57104_ = _57105_ | _57107_ /*1684*/;
assign _57109_ = ~Q[0] /*1683*/;
assign _57108_ = _57109_ & D[35] /*1682*/;
assign _57111_ = _56420_ & _57108_ /*1677*/;
assign _57112_ = _56420_ ^ _57108_ /*1680*/;
assign _57113_ = _57104_ & _57112_ /*1678*/;
assign R_n1[35] = _57104_ ^ _57112_ /*1679*/;
assign _57110_ = _57111_ | _57113_ /*1676*/;
assign _57115_ = ~Q[0] /*1675*/;
assign _57114_ = _57115_ & D[36] /*1674*/;
assign _57117_ = _56421_ & _57114_ /*1669*/;
assign _57118_ = _56421_ ^ _57114_ /*1672*/;
assign _57119_ = _57110_ & _57118_ /*1670*/;
assign R_n1[36] = _57110_ ^ _57118_ /*1671*/;
assign _57116_ = _57117_ | _57119_ /*1668*/;
assign _57121_ = ~Q[0] /*1667*/;
assign _57120_ = _57121_ & D[37] /*1666*/;
assign _57123_ = _56422_ & _57120_ /*1661*/;
assign _57124_ = _56422_ ^ _57120_ /*1664*/;
assign _57125_ = _57116_ & _57124_ /*1662*/;
assign R_n1[37] = _57116_ ^ _57124_ /*1663*/;
assign _57122_ = _57123_ | _57125_ /*1660*/;
assign _57127_ = ~Q[0] /*1659*/;
assign _57126_ = _57127_ & D[38] /*1658*/;
assign _57129_ = _56423_ & _57126_ /*1653*/;
assign _57130_ = _56423_ ^ _57126_ /*1656*/;
assign _57131_ = _57122_ & _57130_ /*1654*/;
assign R_n1[38] = _57122_ ^ _57130_ /*1655*/;
assign _57128_ = _57129_ | _57131_ /*1652*/;
assign _57133_ = ~Q[0] /*1651*/;
assign _57132_ = _57133_ & D[39] /*1650*/;
assign _57135_ = _56424_ & _57132_ /*1645*/;
assign _57136_ = _56424_ ^ _57132_ /*1648*/;
assign _57137_ = _57128_ & _57136_ /*1646*/;
assign R_n1[39] = _57128_ ^ _57136_ /*1647*/;
assign _57134_ = _57135_ | _57137_ /*1644*/;
assign _57139_ = ~Q[0] /*1643*/;
assign _57138_ = _57139_ & D[40] /*1642*/;
assign _57141_ = _56425_ & _57138_ /*1637*/;
assign _57142_ = _56425_ ^ _57138_ /*1640*/;
assign _57143_ = _57134_ & _57142_ /*1638*/;
assign R_n1[40] = _57134_ ^ _57142_ /*1639*/;
assign _57140_ = _57141_ | _57143_ /*1636*/;
assign _57145_ = ~Q[0] /*1635*/;
assign _57144_ = _57145_ & D[41] /*1634*/;
assign _57147_ = _56426_ & _57144_ /*1629*/;
assign _57148_ = _56426_ ^ _57144_ /*1632*/;
assign _57149_ = _57140_ & _57148_ /*1630*/;
assign R_n1[41] = _57140_ ^ _57148_ /*1631*/;
assign _57146_ = _57147_ | _57149_ /*1628*/;
assign _57151_ = ~Q[0] /*1627*/;
assign _57150_ = _57151_ & D[42] /*1626*/;
assign _57153_ = _56427_ & _57150_ /*1621*/;
assign _57154_ = _56427_ ^ _57150_ /*1624*/;
assign _57155_ = _57146_ & _57154_ /*1622*/;
assign R_n1[42] = _57146_ ^ _57154_ /*1623*/;
assign _57152_ = _57153_ | _57155_ /*1620*/;
assign _57157_ = ~Q[0] /*1619*/;
assign _57156_ = _57157_ & D[43] /*1618*/;
assign _57159_ = _56428_ & _57156_ /*1613*/;
assign _57160_ = _56428_ ^ _57156_ /*1616*/;
assign _57161_ = _57152_ & _57160_ /*1614*/;
assign R_n1[43] = _57152_ ^ _57160_ /*1615*/;
assign _57158_ = _57159_ | _57161_ /*1612*/;
assign _57163_ = ~Q[0] /*1611*/;
assign _57162_ = _57163_ & D[44] /*1610*/;
assign _57165_ = _56429_ & _57162_ /*1605*/;
assign _57166_ = _56429_ ^ _57162_ /*1608*/;
assign _57167_ = _57158_ & _57166_ /*1606*/;
assign R_n1[44] = _57158_ ^ _57166_ /*1607*/;
assign _57164_ = _57165_ | _57167_ /*1604*/;
assign _57169_ = ~Q[0] /*1603*/;
assign _57168_ = _57169_ & D[45] /*1602*/;
assign _57171_ = _56430_ & _57168_ /*1597*/;
assign _57172_ = _56430_ ^ _57168_ /*1600*/;
assign _57173_ = _57164_ & _57172_ /*1598*/;
assign R_n1[45] = _57164_ ^ _57172_ /*1599*/;
assign _57170_ = _57171_ | _57173_ /*1596*/;
assign _57175_ = ~Q[0] /*1595*/;
assign _57174_ = _57175_ & D[46] /*1594*/;
assign _57177_ = _56431_ & _57174_ /*1589*/;
assign _57178_ = _56431_ ^ _57174_ /*1592*/;
assign _57179_ = _57170_ & _57178_ /*1590*/;
assign R_n1[46] = _57170_ ^ _57178_ /*1591*/;
assign _57176_ = _57177_ | _57179_ /*1588*/;
assign _57181_ = ~Q[0] /*1587*/;
assign _57180_ = _57181_ & D[47] /*1586*/;
assign _57183_ = _56432_ & _57180_ /*1581*/;
assign _57184_ = _56432_ ^ _57180_ /*1584*/;
assign _57185_ = _57176_ & _57184_ /*1582*/;
assign R_n1[47] = _57176_ ^ _57184_ /*1583*/;
assign _57182_ = _57183_ | _57185_ /*1580*/;
assign _57187_ = ~Q[0] /*1579*/;
assign _57186_ = _57187_ & D[48] /*1578*/;
assign _57189_ = _56433_ & _57186_ /*1573*/;
assign _57190_ = _56433_ ^ _57186_ /*1576*/;
assign _57191_ = _57182_ & _57190_ /*1574*/;
assign R_n1[48] = _57182_ ^ _57190_ /*1575*/;
assign _57188_ = _57189_ | _57191_ /*1572*/;
assign _57193_ = ~Q[0] /*1571*/;
assign _57192_ = _57193_ & D[49] /*1570*/;
assign _57195_ = _56434_ & _57192_ /*1565*/;
assign _57196_ = _56434_ ^ _57192_ /*1568*/;
assign _57197_ = _57188_ & _57196_ /*1566*/;
assign R_n1[49] = _57188_ ^ _57196_ /*1567*/;
assign _57194_ = _57195_ | _57197_ /*1564*/;
assign _57199_ = ~Q[0] /*1563*/;
assign _57198_ = _57199_ & D[50] /*1562*/;
assign _57201_ = _56435_ & _57198_ /*1557*/;
assign _57202_ = _56435_ ^ _57198_ /*1560*/;
assign _57203_ = _57194_ & _57202_ /*1558*/;
assign R_n1[50] = _57194_ ^ _57202_ /*1559*/;
assign _57200_ = _57201_ | _57203_ /*1556*/;
assign _57205_ = ~Q[0] /*1555*/;
assign _57204_ = _57205_ & D[51] /*1554*/;
assign _57207_ = _56436_ & _57204_ /*1549*/;
assign _57208_ = _56436_ ^ _57204_ /*1552*/;
assign _57209_ = _57200_ & _57208_ /*1550*/;
assign R_n1[51] = _57200_ ^ _57208_ /*1551*/;
assign _57206_ = _57207_ | _57209_ /*1548*/;
assign _57211_ = ~Q[0] /*1547*/;
assign _57210_ = _57211_ & D[52] /*1546*/;
assign _57213_ = _56437_ & _57210_ /*1541*/;
assign _57214_ = _56437_ ^ _57210_ /*1544*/;
assign _57215_ = _57206_ & _57214_ /*1542*/;
assign R_n1[52] = _57206_ ^ _57214_ /*1543*/;
assign _57212_ = _57213_ | _57215_ /*1540*/;
assign _57217_ = ~Q[0] /*1539*/;
assign _57216_ = _57217_ & D[53] /*1538*/;
assign _57219_ = _56438_ & _57216_ /*1533*/;
assign _57220_ = _56438_ ^ _57216_ /*1536*/;
assign _57221_ = _57212_ & _57220_ /*1534*/;
assign R_n1[53] = _57212_ ^ _57220_ /*1535*/;
assign _57218_ = _57219_ | _57221_ /*1532*/;
assign _57223_ = ~Q[0] /*1531*/;
assign _57222_ = _57223_ & D[54] /*1530*/;
assign _57225_ = _56439_ & _57222_ /*1525*/;
assign _57226_ = _56439_ ^ _57222_ /*1528*/;
assign _57227_ = _57218_ & _57226_ /*1526*/;
assign R_n1[54] = _57218_ ^ _57226_ /*1527*/;
assign _57224_ = _57225_ | _57227_ /*1524*/;
assign _57229_ = ~Q[0] /*1523*/;
assign _57228_ = _57229_ & D[55] /*1522*/;
assign _57231_ = _56440_ & _57228_ /*1517*/;
assign _57232_ = _56440_ ^ _57228_ /*1520*/;
assign _57233_ = _57224_ & _57232_ /*1518*/;
assign R_n1[55] = _57224_ ^ _57232_ /*1519*/;
assign _57230_ = _57231_ | _57233_ /*1516*/;
assign _57235_ = ~Q[0] /*1515*/;
assign _57234_ = _57235_ & D[56] /*1514*/;
assign _57237_ = _56441_ & _57234_ /*1509*/;
assign _57238_ = _56441_ ^ _57234_ /*1512*/;
assign _57239_ = _57230_ & _57238_ /*1510*/;
assign R_n1[56] = _57230_ ^ _57238_ /*1511*/;
assign _57236_ = _57237_ | _57239_ /*1508*/;
assign _57241_ = ~Q[0] /*1507*/;
assign _57240_ = _57241_ & D[57] /*1506*/;
assign _57243_ = _56442_ & _57240_ /*1501*/;
assign _57244_ = _56442_ ^ _57240_ /*1504*/;
assign _57245_ = _57236_ & _57244_ /*1502*/;
assign R_n1[57] = _57236_ ^ _57244_ /*1503*/;
assign _57242_ = _57243_ | _57245_ /*1500*/;
assign _57247_ = ~Q[0] /*1499*/;
assign _57246_ = _57247_ & D[58] /*1498*/;
assign _57249_ = _56443_ & _57246_ /*1493*/;
assign _57250_ = _56443_ ^ _57246_ /*1496*/;
assign _57251_ = _57242_ & _57250_ /*1494*/;
assign R_n1[58] = _57242_ ^ _57250_ /*1495*/;
assign _57248_ = _57249_ | _57251_ /*1492*/;
assign _57253_ = ~Q[0] /*1491*/;
assign _57252_ = _57253_ & D[59] /*1490*/;
assign _57255_ = _56444_ & _57252_ /*1485*/;
assign _57256_ = _56444_ ^ _57252_ /*1488*/;
assign _57257_ = _57248_ & _57256_ /*1486*/;
assign R_n1[59] = _57248_ ^ _57256_ /*1487*/;
assign _57254_ = _57255_ | _57257_ /*1484*/;
assign _57259_ = ~Q[0] /*1483*/;
assign _57258_ = _57259_ & D[60] /*1482*/;
assign _57261_ = _56445_ & _57258_ /*1477*/;
assign _57262_ = _56445_ ^ _57258_ /*1480*/;
assign _57263_ = _57254_ & _57262_ /*1478*/;
assign R_n1[60] = _57254_ ^ _57262_ /*1479*/;
assign _57260_ = _57261_ | _57263_ /*1476*/;
assign _57265_ = ~Q[0] /*1475*/;
assign _57264_ = _57265_ & D[61] /*1474*/;
assign _57267_ = _56446_ & _57264_ /*1469*/;
assign _57268_ = _56446_ ^ _57264_ /*1472*/;
assign _57269_ = _57260_ & _57268_ /*1470*/;
assign R_n1[61] = _57260_ ^ _57268_ /*1471*/;
assign _57266_ = _57267_ | _57269_ /*1468*/;
assign _57271_ = ~Q[0] /*1467*/;
assign _57270_ = _57271_ & D[62] /*1466*/;
assign _57273_ = _56447_ & _57270_ /*1461*/;
assign _57274_ = _56447_ ^ _57270_ /*1464*/;
assign _57275_ = _57266_ & _57274_ /*1462*/;
assign R_n1[62] = _57266_ ^ _57274_ /*1463*/;
assign _57272_ = _57273_ | _57275_ /*1460*/;
endmodule
