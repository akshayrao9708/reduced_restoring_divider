module divider(q, rout, rin, div);
  wire _0_;
  wire _1_;
  wire _2_;
  wire _3_;
  wire _4_;
  wire _5_;
  wire _6_;
  wire _7_;
  wire _8_;
  wire _9_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  wire _38_;
  wire _39_;
  wire _40_;
  wire _41_;
  wire _42_;
  wire _43_;
  wire _44_;
  wire _45_;
  wire _46_;
  wire _47_;
  wire _48_;
  wire _49_;
  wire _50_;
  wire _51_;
  wire _52_;
  wire _53_;
  wire _54_;
  wire _55_;
  wire _56_;
  wire _57_;
  wire _58_;
  wire _59_;
  wire _60_;
  wire _61_;
  wire _62_;
  wire _63_;
  wire _64_;
  wire _65_;
  wire _66_;
  wire _67_;
  wire _68_;
  wire _69_;
  wire _70_;
  wire _71_;
  wire _72_;
  wire _73_;
  wire _74_;
  wire _75_;
  wire _76_;
  wire _77_;
  wire _78_;
  wire _79_;
  wire _80_;
  wire _81_;
  wire _82_;
  wire _83_;
  wire _84_;
  wire _85_;
  wire _86_;
  wire _87_;
  wire _88_;
  wire _89_;
  wire _90_;
  wire _91_;
  wire _92_;
  wire _93_;
  wire _94_;
  wire _95_;
  wire _96_;
  wire _97_;
  wire _98_;
  wire _99_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire _304_;
  wire _305_;
  wire _306_;
  wire _307_;
  wire _308_;
  wire _309_;
  wire _310_;
  wire _311_;
  wire _312_;
  wire _313_;
  wire _314_;
  wire _315_;
  wire _316_;
  wire _317_;
  wire _318_;
  wire _319_;
  wire _320_;
  wire _321_;
  wire _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire _326_;
  wire _327_;
  wire _328_;
  wire _329_;
  wire _330_;
  wire _331_;
  wire _332_;
  wire _333_;
  wire _334_;
  wire _335_;
  wire _336_;
  wire _337_;
  wire _338_;
  wire _339_;
  wire _340_;
  wire _341_;
  wire _342_;
  wire _343_;
  wire _344_;
  wire _345_;
  wire _346_;
  wire _347_;
  wire _348_;
  wire _349_;
  wire _350_;
  wire _351_;
  wire _352_;
  wire _353_;
  wire _354_;
  wire _355_;
  wire _356_;
  wire _357_;
  wire _358_;
  wire _359_;
  wire _360_;
  wire _361_;
  wire _362_;
  wire _363_;
  wire _364_;
  wire _365_;
  wire _366_;
  wire _367_;
  wire _368_;
  wire _369_;
  wire _370_;
  wire _371_;
  wire _372_;
  wire _373_;
  wire _374_;
  wire _375_;
  wire _376_;
  wire _377_;
  wire _378_;
  wire _379_;
  wire _380_;
  wire _381_;
  wire _382_;
  wire _383_;
  wire _384_;
  wire _385_;
  wire _386_;
  wire _387_;
  wire _388_;
  wire _389_;
  wire _390_;
  wire _391_;
  wire _392_;
  wire _393_;
  wire _394_;
  wire _395_;
  wire _396_;
  wire _397_;
  wire _398_;
  wire _399_;
  wire _400_;
  wire _401_;
  wire _402_;
  wire _403_;
  wire _404_;
  wire _405_;
  wire _406_;
  wire _407_;
  wire _408_;
  wire _409_;
  wire _410_;
  wire _411_;
  wire _412_;
  wire _413_;
  wire _414_;
  wire _415_;
  wire _416_;
  wire _417_;
  wire _418_;
  wire _419_;
  wire _420_;
  wire _421_;
  wire _422_;
  wire _423_;
  wire _424_;
  wire _425_;
  wire _426_;
  wire _427_;
  wire _428_;
  wire _429_;
  wire _430_;
  wire _431_;
  wire _432_;
  wire _433_;
  wire _434_;
  wire _435_;
  wire _436_;
  wire _437_;
  wire _438_;
  wire _439_;
  wire _440_;
  wire _441_;
  wire _442_;
  wire _443_;
  wire _444_;
  wire _445_;
  wire _446_;
  wire _447_;
  wire _448_;
  wire _449_;
  wire _450_;
  wire _451_;
  wire _452_;
  wire _453_;
  wire _454_;
  wire _455_;
  wire _456_;
  wire _457_;
  wire _458_;
  wire _459_;
  wire _460_;
  wire _461_;
  wire _462_;
  wire _463_;
  wire _464_;
  wire _465_;
  wire _466_;
  wire _467_;
  wire _468_;
  wire _469_;
  wire _470_;
  wire _471_;
  wire _472_;
  wire _473_;
  wire _474_;
  wire _475_;
  wire _476_;
  wire _477_;
  wire _478_;
  wire _479_;
  wire _480_;
  wire _481_;
  wire _482_;
  wire _483_;
  wire _484_;
  wire _485_;
  wire _486_;
  wire _487_;
  wire _488_;
  wire _489_;
  wire _490_;
  wire _491_;
  wire _492_;
  wire _493_;
  wire _494_;
  wire _495_;
  wire _496_;
  wire _497_;
  wire _498_;
  wire _499_;
  wire _500_;
  wire _501_;
  wire _502_;
  wire _503_;
  wire _504_;
  wire _505_;
  wire _506_;
  wire _507_;
  wire _508_;
  wire _509_;
  wire _510_;
  wire _511_;
  wire _512_;
  wire _513_;
  wire _514_;
  wire _515_;
  wire _516_;
  wire _517_;
  wire _518_;
  wire _519_;
  wire _520_;
  wire _521_;
  wire _522_;
  wire _523_;
  wire _524_;
  wire _525_;
  wire _526_;
  wire _527_;
  wire _528_;
  wire _529_;
  wire _530_;
  wire _531_;
  wire _532_;
  wire _533_;
  wire _534_;
  wire _535_;
  wire _536_;
  wire _537_;
  wire _538_;
  wire _539_;
  wire _540_;
  wire _541_;
  wire _542_;
  wire _543_;
  wire _544_;
  wire _545_;
  wire _546_;
  wire _547_;
  wire _548_;
  wire _549_;
  wire _550_;
  wire _551_;
  wire _552_;
  wire _553_;
  wire _554_;
  wire _555_;
  wire _556_;
  wire _557_;
  wire _558_;
  wire _559_;
  wire _560_;
  wire _561_;
  wire _562_;
  wire _563_;
  wire _564_;
  wire _565_;
  wire _566_;
  wire _567_;
  wire _568_;
  wire _569_;
  wire _570_;
  wire _571_;
  wire _572_;
  wire _573_;
  wire _574_;
  wire _575_;
  wire _576_;
  wire _577_;
  wire _578_;
  wire _579_;
  wire _580_;
  wire _581_;
  wire _582_;
  wire _583_;
  wire _584_;
  wire _585_;
  wire _586_;
  wire _587_;
  wire _588_;
  wire _589_;
  wire _590_;
  wire _591_;
  wire _592_;
  wire _593_;
  wire _594_;
  wire _595_;
  wire _596_;
  wire _597_;
  wire _598_;
  wire _599_;
  wire _600_;
  wire _601_;
  wire _602_;
  wire _603_;
  wire _604_;
  wire _605_;
  wire _606_;
  wire _607_;
  wire _608_;
  wire _609_;
  wire _610_;
  wire _611_;
  wire _612_;
  wire _613_;
  wire _614_;
  wire _615_;
  wire _616_;
  wire _617_;
  wire _618_;
  wire _619_;
  wire _620_;
  wire _621_;
  wire _622_;
  wire _623_;
  wire _624_;
  wire _625_;
  wire _626_;
  wire _627_;
  wire _628_;
  wire _629_;
  wire _630_;
  wire _631_;
  wire _632_;
  wire _633_;
  wire _634_;
  wire _635_;
  wire _636_;
  wire _637_;
  wire _638_;
  wire _639_;
  wire _640_;
  wire _641_;
  wire _642_;
  wire _643_;
  wire _644_;
  wire _645_;
  wire _646_;
  wire _647_;
  wire _648_;
  wire _649_;
  wire _650_;
  wire _651_;
  wire _652_;
  wire _653_;
  wire _654_;
  wire _655_;
  wire _656_;
  wire _657_;
  wire _658_;
  wire _659_;
  wire _660_;
  wire _661_;
  wire _662_;
  wire _663_;
  wire _664_;
  wire _665_;
  wire _666_;
  wire _667_;
  wire _668_;
  wire _669_;
  wire _670_;
  wire _671_;
  wire _672_;
  wire _673_;
  wire _674_;
  wire _675_;
  wire _676_;
  wire _677_;
  wire _678_;
  wire _679_;
  wire _680_;
  wire _681_;
  wire _682_;
  wire _683_;
  wire _684_;
  wire _685_;
  wire _686_;
  wire _687_;
  wire _688_;
  wire _689_;
  wire _690_;
  wire _691_;
  wire _692_;
  wire _693_;
  wire _694_;
  wire _695_;
  wire _696_;
  wire _697_;
  wire _698_;
  wire _699_;
  wire _700_;
  wire _701_;
  wire _702_;
  wire _703_;
  wire _704_;
  wire _705_;
  wire _706_;
  wire _707_;
  wire _708_;
  wire _709_;
  wire _710_;
  wire _711_;
  wire _712_;
  wire _713_;
  wire _714_;
  wire _715_;
  wire _716_;
  wire _717_;
  wire _718_;
  wire _719_;
  wire _720_;
  wire _721_;
  wire _722_;
  wire _723_;
  wire _724_;
  wire _725_;
  wire _726_;
  wire _727_;
  wire _728_;
  wire _729_;
  wire _730_;
  wire _731_;
  wire _732_;
  wire _733_;
  wire _734_;
  wire _735_;
  wire _736_;
  wire _737_;
  wire _738_;
  wire _739_;
  wire _740_;
  wire _741_;
  wire _742_;
  wire _743_;
  wire _744_;
  wire _745_;
  wire _746_;
  wire _747_;
  wire _748_;
  wire _749_;
  wire _750_;
  wire _751_;
  wire _752_;
  wire _753_;
  wire _754_;
  wire _755_;
  wire _756_;
  wire _757_;
  wire _758_;
  wire _759_;
  wire _760_;
  wire _761_;
  wire _762_;
  wire _763_;
  wire _764_;
  wire _765_;
  wire _766_;
  wire _767_;
  wire _768_;
  wire _769_;
  wire _770_;
  wire _771_;
  wire _772_;
  wire _773_;
  wire _774_;
  wire _775_;
  wire _776_;
  wire _777_;
  wire _778_;
  wire _779_;
  wire _780_;
  wire _781_;
  wire _782_;
  wire _783_;
  wire _784_;
  wire _785_;
  wire _786_;
  wire _787_;
  wire _788_;
  wire _789_;
  wire _790_;
  wire _791_;
  wire _792_;
  wire _793_;
  wire _794_;
  wire _795_;
  wire _796_;
  wire _797_;
  wire _798_;
  wire _799_;
  wire _800_;
  wire _801_;
  wire _802_;
  wire _803_;
  wire _804_;
  wire _805_;
  wire _806_;
  wire _807_;
  wire _808_;
  wire _809_;
  wire _810_;
  wire _811_;
  wire _812_;
  wire _813_;
  wire _814_;
  wire _815_;
  wire _816_;
  wire _817_;
  wire _818_;
  wire _819_;
  wire _820_;
  wire _821_;
  wire _822_;
  wire _823_;
  wire _824_;
  wire _825_;
  wire _826_;
  wire _827_;
  wire _828_;
  wire _829_;
  wire _830_;
  wire _831_;
  wire _832_;
  wire _833_;
  wire _834_;
  wire _835_;
  wire _836_;
  wire _837_;
  wire _838_;
  wire _839_;
  wire _840_;
  wire _841_;
  wire _842_;
  wire _843_;
  wire _844_;
  wire _845_;
  wire _846_;
  wire _847_;
  wire _848_;
  wire _849_;
  wire _850_;
  wire _851_;
  wire _852_;
  wire _853_;
  wire _854_;
  wire _855_;
  wire _856_;
  wire _857_;
  wire _858_;
  wire _859_;
  wire _860_;
  wire _861_;
  wire _862_;
  wire _863_;
  wire _864_;
  wire _865_;
  wire _866_;
  wire _867_;
  wire _868_;
  wire _869_;
  wire _870_;
  wire _871_;
  wire _872_;
  wire _873_;
  wire _874_;
  wire _875_;
  wire _876_;
  wire _877_;
  wire _878_;
  wire _879_;
  wire _880_;
  wire _881_;
  wire _882_;
  wire _883_;
  wire _884_;
  wire _885_;
  wire _886_;
  wire _887_;
  wire _888_;
  wire _889_;
  wire _890_;
  wire _891_;
  wire _892_;
  wire _893_;
  wire _894_;
  wire _895_;
  wire _896_;
  wire _897_;
  wire _898_;
  wire _899_;
  wire _900_;
  wire _901_;
  wire _902_;
  wire _903_;
  wire _904_;
  wire _905_;
  wire _906_;
  wire _907_;
  wire _908_;
  wire _909_;
  wire _910_;
  wire _911_;
  wire _912_;
  wire _913_;
  wire _914_;
  wire _915_;
  wire _916_;
  wire _917_;
  wire _918_;
  wire _919_;
  wire _920_;
  wire _921_;
  wire _922_;
  wire _923_;
  wire _924_;
  wire _925_;
  wire _926_;
  wire _927_;
  wire _928_;
  wire _929_;
  wire _930_;
  wire _931_;
  wire _932_;
  wire _933_;
  wire _934_;
  wire _935_;
  wire _936_;
  wire _937_;
  wire _938_;
  wire _939_;
  wire _940_;
  wire _941_;
  wire _942_;
  wire _943_;
  wire _944_;
  wire _945_;
  wire _946_;
  wire _947_;
  wire _948_;
  wire _949_;
  wire _950_;
  wire _951_;
  wire _952_;
  wire _953_;
  wire _954_;
  wire _955_;
  wire _956_;
  wire _957_;
  wire _958_;
  wire _959_;
  wire _960_;
  wire _961_;
  wire _962_;
  wire _963_;
  wire _964_;
  wire _965_;
  wire _966_;
  wire _967_;
  wire _968_;
  wire _969_;
  wire _970_;
  wire _971_;
  wire _972_;
  wire _973_;
  wire _974_;
  wire _975_;
  wire _976_;
  wire _977_;
  wire _978_;
  wire _979_;
  wire _980_;
  wire _981_;
  wire _982_;
  wire _983_;
  wire _984_;
  wire _985_;
  wire _986_;
  wire _987_;
  wire _988_;
  wire _989_;
  wire _990_;
  wire _991_;
  wire _992_;
  wire _993_;
  wire _994_;
  wire _995_;
  wire _996_;
  wire _997_;
  wire _998_;
  wire _999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire [22:0] r_0;
  wire [22:0] r_1;
  wire [11:0] m_1;
  wire [11:0] sum_1;
  wire [11:0] inv_1;
  wire [21:0] r_2;
  wire [11:0] m_2;
  wire [11:0] sum_2;
  wire [11:0] inv_2;
  wire [20:0] r_3;
  wire [11:0] m_3;
  wire [11:0] sum_3;
  wire [11:0] inv_3;
  wire [19:0] r_4;
  wire [11:0] m_4;
  wire [11:0] sum_4;
  wire [11:0] inv_4;
  wire [18:0] r_5;
  wire [11:0] m_5;
  wire [11:0] sum_5;
  wire [11:0] inv_5;
  wire [17:0] r_6;
  wire [11:0] m_6;
  wire [11:0] sum_6;
  wire [11:0] inv_6;
  wire [16:0] r_7;
  wire [11:0] m_7;
  wire [11:0] sum_7;
  wire [11:0] inv_7;
  wire [15:0] r_8;
  wire [11:0] m_8;
  wire [11:0] sum_8;
  wire [11:0] inv_8;
  wire [14:0] r_9;
  wire [11:0] m_9;
  wire [11:0] sum_9;
  wire [11:0] inv_9;
  wire [13:0] r_10;
  wire [11:0] m_10;
  wire [11:0] sum_10;
  wire [11:0] inv_10;
  wire [12:0] r_11;
  wire [11:0] m_11;
  wire [11:0] sum_11;
  wire [11:0] inv_11;
  wire [11:0] r_12;
  wire [11:0] m_12;
  wire [11:0] sum_12;
  wire [11:0] inv_12;
  wire zeroWire;
  wire oneWire;
  input [21:0] rin;
  input [10:0] div;
  output [11:0] q;
  output [11:0] rout;
  assign zeroWire = 1'b0 /*0*/;
  assign oneWire = 1'b1 /*0*/;
  assign r_0[0] = rin[0] /*3155*/;
  assign r_0[1] = rin[1] /*3154*/;
  assign r_0[2] = rin[2] /*3153*/;
  assign r_0[3] = rin[3] /*3152*/;
  assign r_0[4] = rin[4] /*3151*/;
  assign r_0[5] = rin[5] /*3150*/;
  assign r_0[6] = rin[6] /*3149*/;
  assign r_0[7] = rin[7] /*3148*/;
  assign r_0[8] = rin[8] /*3147*/;
  assign r_0[9] = rin[9] /*3146*/;
  assign r_0[10] = rin[10] /*3145*/;
  assign r_0[11] = rin[11] /*3144*/;
  assign r_0[12] = rin[12] /*3143*/;
  assign r_0[13] = rin[13] /*3142*/;
  assign r_0[14] = rin[14] /*3141*/;
  assign r_0[15] = rin[15] /*3140*/;
  assign r_0[16] = rin[16] /*3139*/;
  assign r_0[17] = rin[17] /*3138*/;
  assign r_0[18] = rin[18] /*3137*/;
  assign r_0[19] = rin[19] /*3136*/;
  assign r_0[20] = rin[20] /*3135*/;
  assign r_0[21] = rin[21] /*3134*/;
  assign r_0[22] = zeroWire /*3133*/;
  assign inv_1[0] = ~div[0] /*3132*/;
  assign inv_1[1] = ~div[1] /*3131*/;
  assign inv_1[2] = ~div[2] /*3130*/;
  assign inv_1[3] = ~div[3] /*3129*/;
  assign inv_1[4] = ~div[4] /*3128*/;
  assign inv_1[5] = ~div[5] /*3127*/;
  assign inv_1[6] = ~div[6] /*3126*/;
  assign inv_1[7] = ~div[7] /*3125*/;
  assign inv_1[8] = ~div[8] /*3124*/;
  assign inv_1[9] = ~div[9] /*3123*/;
  assign inv_1[10] = ~div[10] /*3122*/;
assign inv_1[11] = oneWire /*3121*/;
  assign _0_ = inv_1[0] ^ r_0[11] /*3119*/;
  assign sum_1[0] = _0_ ^ oneWire /*3118*/;
  assign _1_ = _0_ & oneWire /*3117*/;
  assign _2_ = inv_1[0] & r_0[11] /*3116*/;
  assign _3_ = _1_ | _2_ /*3115*/;
  assign _4_ = inv_1[1] ^ r_0[12] /*3114*/;
  assign sum_1[1] = _4_ ^ _3_ /*3113*/;
  assign _5_ = _4_ & _3_ /*3112*/;
  assign _6_ = inv_1[1] & r_0[12] /*3111*/;
  assign _7_ = _5_ | _6_ /*3110*/;
  assign _8_ = inv_1[2] ^ r_0[13] /*3108*/;
  assign sum_1[2] = _8_ ^ _7_ /*3107*/;
  assign _9_ = _8_ & _7_ /*3106*/;
  assign _10_ = inv_1[2] & r_0[13] /*3105*/;
  assign _11_ = _9_ | _10_ /*3104*/;
  assign _12_ = inv_1[3] ^ r_0[14] /*3102*/;
  assign sum_1[3] = _12_ ^ _11_ /*3101*/;
  assign _13_ = _12_ & _11_ /*3100*/;
  assign _14_ = inv_1[3] & r_0[14] /*3099*/;
  assign _15_ = _13_ | _14_ /*3098*/;
  assign _16_ = inv_1[4] ^ r_0[15] /*3096*/;
  assign sum_1[4] = _16_ ^ _15_ /*3095*/;
  assign _17_ = _16_ & _15_ /*3094*/;
  assign _18_ = inv_1[4] & r_0[15] /*3093*/;
  assign _19_ = _17_ | _18_ /*3092*/;
  assign _20_ = inv_1[5] ^ r_0[16] /*3090*/;
  assign sum_1[5] = _20_ ^ _19_ /*3089*/;
  assign _21_ = _20_ & _19_ /*3088*/;
  assign _22_ = inv_1[5] & r_0[16] /*3087*/;
  assign _23_ = _21_ | _22_ /*3086*/;
  assign _24_ = inv_1[6] ^ r_0[17] /*3084*/;
  assign sum_1[6] = _24_ ^ _23_ /*3083*/;
  assign _25_ = _24_ & _23_ /*3082*/;
  assign _26_ = inv_1[6] & r_0[17] /*3081*/;
  assign _27_ = _25_ | _26_ /*3080*/;
  assign _28_ = inv_1[7] ^ r_0[18] /*3078*/;
  assign sum_1[7] = _28_ ^ _27_ /*3077*/;
  assign _29_ = _28_ & _27_ /*3076*/;
  assign _30_ = inv_1[7] & r_0[18] /*3075*/;
  assign _31_ = _29_ | _30_ /*3074*/;
  assign _32_ = inv_1[8] ^ r_0[19] /*3072*/;
  assign sum_1[8] = _32_ ^ _31_ /*3071*/;
  assign _33_ = _32_ & _31_ /*3070*/;
  assign _34_ = inv_1[8] & r_0[19] /*3069*/;
  assign _35_ = _33_ | _34_ /*3068*/;
  assign _36_ = inv_1[9] ^ r_0[20] /*3066*/;
  assign sum_1[9] = _36_ ^ _35_ /*3065*/;
  assign _37_ = _36_ & _35_ /*3064*/;
  assign _38_ = inv_1[9] & r_0[20] /*3063*/;
  assign _39_ = _37_ | _38_ /*3062*/;
  assign _40_ = inv_1[10] ^ r_0[21] /*3060*/;
  assign sum_1[10] = _40_ ^ _39_ /*3059*/;
  assign _41_ = _40_ & _39_ /*3058*/;
  assign _42_ = inv_1[10] & r_0[21] /*3057*/;
  assign _43_ = _41_ | _42_ /*3056*/;
  assign _44_ = inv_1[11] ^ r_0[22] /*3054*/;
  assign sum_1[11] = _44_ ^ _43_ /*3053*/;
  assign _45_ = _44_ & _43_ /*3052*/;
  assign _46_ = inv_1[11] & r_0[22] /*3051*/;
  assign _47_ = _45_ | _46_ /*3050*/;
  assign q[11] = ~sum_1[11] /*3057*/;
  assign m_1[0] = r_0[11] /*3056*/;
  assign m_1[1] = r_0[12] /*3055*/;
  assign m_1[2] = r_0[13] /*3054*/;
  assign m_1[3] = r_0[14] /*3053*/;
  assign m_1[4] = r_0[15] /*3052*/;
  assign m_1[5] = r_0[16] /*3051*/;
  assign m_1[6] = r_0[17] /*3050*/;
  assign m_1[7] = r_0[18] /*3049*/;
  assign m_1[8] = r_0[19] /*3048*/;
  assign m_1[9] = r_0[20] /*3047*/;
  assign m_1[10] = r_0[21] /*3046*/;
  assign m_1[11] = r_0[22] /*3045*/;
  assign _48_ = ~q[11] /*3043*/;
  assign _49_ = sum_1[0] & q[11] /*3042*/;
  assign _50_ = m_1[0] & _48_ /*3041*/;
  assign r_1[11] = _50_ | _49_ /*3040*/;
  assign _51_ = ~q[11] /*3039*/;
  assign _52_ = sum_1[1] & q[11] /*3038*/;
  assign _53_ = m_1[1] & _51_ /*3037*/;
  assign r_1[12] = _53_ | _52_ /*3036*/;
  assign _54_ = ~q[11] /*3035*/;
  assign _55_ = sum_1[2] & q[11] /*3034*/;
  assign _56_ = m_1[2] & _54_ /*3033*/;
  assign r_1[13] = _56_ | _55_ /*3032*/;
  assign _57_ = ~q[11] /*3031*/;
  assign _58_ = sum_1[3] & q[11] /*3030*/;
  assign _59_ = m_1[3] & _57_ /*3029*/;
  assign r_1[14] = _59_ | _58_ /*3028*/;
  assign _60_ = ~q[11] /*3027*/;
  assign _61_ = sum_1[4] & q[11] /*3026*/;
  assign _62_ = m_1[4] & _60_ /*3025*/;
  assign r_1[15] = _62_ | _61_ /*3024*/;
  assign _63_ = ~q[11] /*3023*/;
  assign _64_ = sum_1[5] & q[11] /*3022*/;
  assign _65_ = m_1[5] & _63_ /*3021*/;
  assign r_1[16] = _65_ | _64_ /*3020*/;
  assign _66_ = ~q[11] /*3019*/;
  assign _67_ = sum_1[6] & q[11] /*3018*/;
  assign _68_ = m_1[6] & _66_ /*3017*/;
  assign r_1[17] = _68_ | _67_ /*3016*/;
  assign _69_ = ~q[11] /*3015*/;
  assign _70_ = sum_1[7] & q[11] /*3014*/;
  assign _71_ = m_1[7] & _69_ /*3013*/;
  assign r_1[18] = _71_ | _70_ /*3012*/;
  assign _72_ = ~q[11] /*3011*/;
  assign _73_ = sum_1[8] & q[11] /*3010*/;
  assign _74_ = m_1[8] & _72_ /*3009*/;
  assign r_1[19] = _74_ | _73_ /*3008*/;
  assign _75_ = ~q[11] /*3007*/;
  assign _76_ = sum_1[9] & q[11] /*3006*/;
  assign _77_ = m_1[9] & _75_ /*3005*/;
  assign r_1[20] = _77_ | _76_ /*3004*/;
  assign _78_ = ~q[11] /*3003*/;
  assign _79_ = sum_1[10] & q[11] /*3002*/;
  assign _80_ = m_1[10] & _78_ /*3001*/;
  assign r_1[21] = _80_ | _79_ /*3000*/;
  assign _81_ = ~q[11] /*2999*/;
  assign _82_ = sum_1[11] & q[11] /*2998*/;
  assign _83_ = m_1[11] & _81_ /*2997*/;
  assign r_1[22] = _83_ | _82_ /*2996*/;
assign r_1[0]= r_0[0] /*2995*/;
assign r_1[1]= r_0[1] /*2994*/;
assign r_1[2]= r_0[2] /*2993*/;
assign r_1[3]= r_0[3] /*2992*/;
assign r_1[4]= r_0[4] /*2991*/;
assign r_1[5]= r_0[5] /*2990*/;
assign r_1[6]= r_0[6] /*2989*/;
assign r_1[7]= r_0[7] /*2988*/;
assign r_1[8]= r_0[8] /*2987*/;
assign r_1[9]= r_0[9] /*2986*/;
assign r_1[10]= r_0[10] /*2985*/;
  assign inv_2[0] = ~div[0] /*2964*/;
  assign inv_2[1] = ~div[1] /*2963*/;
  assign inv_2[2] = ~div[2] /*2962*/;
  assign inv_2[3] = ~div[3] /*2961*/;
  assign inv_2[4] = ~div[4] /*2960*/;
  assign inv_2[5] = ~div[5] /*2959*/;
  assign inv_2[6] = ~div[6] /*2958*/;
  assign inv_2[7] = ~div[7] /*2957*/;
  assign inv_2[8] = ~div[8] /*2956*/;
  assign inv_2[9] = ~div[9] /*2955*/;
  assign inv_2[10] = ~div[10] /*2954*/;
assign inv_2[11] = oneWire /*2953*/;
  assign _84_ = inv_2[0] ^ r_1[10] /*2951*/;
  assign sum_2[0] = _84_ ^ oneWire /*2950*/;
  assign _85_ = _84_ & oneWire /*2949*/;
  assign _86_ = inv_2[0] & r_1[10] /*2948*/;
  assign _87_ = _85_ | _86_ /*2947*/;
  assign _88_ = inv_2[1] ^ r_1[11] /*2946*/;
  assign sum_2[1] = _88_ ^ _87_ /*2945*/;
  assign _89_ = _88_ & _87_ /*2944*/;
  assign _90_ = inv_2[1] & r_1[11] /*2943*/;
  assign _91_ = _89_ | _90_ /*2942*/;
  assign _92_ = inv_2[2] ^ r_1[12] /*2940*/;
  assign sum_2[2] = _92_ ^ _91_ /*2939*/;
  assign _93_ = _92_ & _91_ /*2938*/;
  assign _94_ = inv_2[2] & r_1[12] /*2937*/;
  assign _95_ = _93_ | _94_ /*2936*/;
  assign _96_ = inv_2[3] ^ r_1[13] /*2934*/;
  assign sum_2[3] = _96_ ^ _95_ /*2933*/;
  assign _97_ = _96_ & _95_ /*2932*/;
  assign _98_ = inv_2[3] & r_1[13] /*2931*/;
  assign _99_ = _97_ | _98_ /*2930*/;
  assign _100_ = inv_2[4] ^ r_1[14] /*2928*/;
  assign sum_2[4] = _100_ ^ _99_ /*2927*/;
  assign _101_ = _100_ & _99_ /*2926*/;
  assign _102_ = inv_2[4] & r_1[14] /*2925*/;
  assign _103_ = _101_ | _102_ /*2924*/;
  assign _104_ = inv_2[5] ^ r_1[15] /*2922*/;
  assign sum_2[5] = _104_ ^ _103_ /*2921*/;
  assign _105_ = _104_ & _103_ /*2920*/;
  assign _106_ = inv_2[5] & r_1[15] /*2919*/;
  assign _107_ = _105_ | _106_ /*2918*/;
  assign _108_ = inv_2[6] ^ r_1[16] /*2916*/;
  assign sum_2[6] = _108_ ^ _107_ /*2915*/;
  assign _109_ = _108_ & _107_ /*2914*/;
  assign _110_ = inv_2[6] & r_1[16] /*2913*/;
  assign _111_ = _109_ | _110_ /*2912*/;
  assign _112_ = inv_2[7] ^ r_1[17] /*2910*/;
  assign sum_2[7] = _112_ ^ _111_ /*2909*/;
  assign _113_ = _112_ & _111_ /*2908*/;
  assign _114_ = inv_2[7] & r_1[17] /*2907*/;
  assign _115_ = _113_ | _114_ /*2906*/;
  assign _116_ = inv_2[8] ^ r_1[18] /*2904*/;
  assign sum_2[8] = _116_ ^ _115_ /*2903*/;
  assign _117_ = _116_ & _115_ /*2902*/;
  assign _118_ = inv_2[8] & r_1[18] /*2901*/;
  assign _119_ = _117_ | _118_ /*2900*/;
  assign _120_ = inv_2[9] ^ r_1[19] /*2898*/;
  assign sum_2[9] = _120_ ^ _119_ /*2897*/;
  assign _121_ = _120_ & _119_ /*2896*/;
  assign _122_ = inv_2[9] & r_1[19] /*2895*/;
  assign _123_ = _121_ | _122_ /*2894*/;
  assign _124_ = inv_2[10] ^ r_1[20] /*2892*/;
  assign sum_2[10] = _124_ ^ _123_ /*2891*/;
  assign _125_ = _124_ & _123_ /*2890*/;
  assign _126_ = inv_2[10] & r_1[20] /*2889*/;
  assign _127_ = _125_ | _126_ /*2888*/;
  assign _128_ = inv_2[11] ^ r_1[21] /*2886*/;
  assign sum_2[11] = _128_ ^ _127_ /*2885*/;
  assign _129_ = _128_ & _127_ /*2884*/;
  assign _130_ = inv_2[11] & r_1[21] /*2883*/;
  assign _131_ = _129_ | _130_ /*2882*/;
  assign q[10] = ~sum_2[11] /*2889*/;
  assign m_2[0] = r_1[10] /*2888*/;
  assign m_2[1] = r_1[11] /*2887*/;
  assign m_2[2] = r_1[12] /*2886*/;
  assign m_2[3] = r_1[13] /*2885*/;
  assign m_2[4] = r_1[14] /*2884*/;
  assign m_2[5] = r_1[15] /*2883*/;
  assign m_2[6] = r_1[16] /*2882*/;
  assign m_2[7] = r_1[17] /*2881*/;
  assign m_2[8] = r_1[18] /*2880*/;
  assign m_2[9] = r_1[19] /*2879*/;
  assign m_2[10] = r_1[20] /*2878*/;
  assign m_2[11] = r_1[21] /*2877*/;
  assign _132_ = ~q[10] /*2875*/;
  assign _133_ = sum_2[0] & q[10] /*2874*/;
  assign _134_ = m_2[0] & _132_ /*2873*/;
  assign r_2[10] = _134_ | _133_ /*2872*/;
  assign _135_ = ~q[10] /*2871*/;
  assign _136_ = sum_2[1] & q[10] /*2870*/;
  assign _137_ = m_2[1] & _135_ /*2869*/;
  assign r_2[11] = _137_ | _136_ /*2868*/;
  assign _138_ = ~q[10] /*2867*/;
  assign _139_ = sum_2[2] & q[10] /*2866*/;
  assign _140_ = m_2[2] & _138_ /*2865*/;
  assign r_2[12] = _140_ | _139_ /*2864*/;
  assign _141_ = ~q[10] /*2863*/;
  assign _142_ = sum_2[3] & q[10] /*2862*/;
  assign _143_ = m_2[3] & _141_ /*2861*/;
  assign r_2[13] = _143_ | _142_ /*2860*/;
  assign _144_ = ~q[10] /*2859*/;
  assign _145_ = sum_2[4] & q[10] /*2858*/;
  assign _146_ = m_2[4] & _144_ /*2857*/;
  assign r_2[14] = _146_ | _145_ /*2856*/;
  assign _147_ = ~q[10] /*2855*/;
  assign _148_ = sum_2[5] & q[10] /*2854*/;
  assign _149_ = m_2[5] & _147_ /*2853*/;
  assign r_2[15] = _149_ | _148_ /*2852*/;
  assign _150_ = ~q[10] /*2851*/;
  assign _151_ = sum_2[6] & q[10] /*2850*/;
  assign _152_ = m_2[6] & _150_ /*2849*/;
  assign r_2[16] = _152_ | _151_ /*2848*/;
  assign _153_ = ~q[10] /*2847*/;
  assign _154_ = sum_2[7] & q[10] /*2846*/;
  assign _155_ = m_2[7] & _153_ /*2845*/;
  assign r_2[17] = _155_ | _154_ /*2844*/;
  assign _156_ = ~q[10] /*2843*/;
  assign _157_ = sum_2[8] & q[10] /*2842*/;
  assign _158_ = m_2[8] & _156_ /*2841*/;
  assign r_2[18] = _158_ | _157_ /*2840*/;
  assign _159_ = ~q[10] /*2839*/;
  assign _160_ = sum_2[9] & q[10] /*2838*/;
  assign _161_ = m_2[9] & _159_ /*2837*/;
  assign r_2[19] = _161_ | _160_ /*2836*/;
  assign _162_ = ~q[10] /*2835*/;
  assign _163_ = sum_2[10] & q[10] /*2834*/;
  assign _164_ = m_2[10] & _162_ /*2833*/;
  assign r_2[20] = _164_ | _163_ /*2832*/;
  assign _165_ = ~q[10] /*2831*/;
  assign _166_ = sum_2[11] & q[10] /*2830*/;
  assign _167_ = m_2[11] & _165_ /*2829*/;
  assign r_2[21] = _167_ | _166_ /*2828*/;
assign r_2[0]= r_1[0] /*2827*/;
assign r_2[1]= r_1[1] /*2826*/;
assign r_2[2]= r_1[2] /*2825*/;
assign r_2[3]= r_1[3] /*2824*/;
assign r_2[4]= r_1[4] /*2823*/;
assign r_2[5]= r_1[5] /*2822*/;
assign r_2[6]= r_1[6] /*2821*/;
assign r_2[7]= r_1[7] /*2820*/;
assign r_2[8]= r_1[8] /*2819*/;
assign r_2[9]= r_1[9] /*2818*/;
  assign inv_3[0] = ~div[0] /*2796*/;
  assign inv_3[1] = ~div[1] /*2795*/;
  assign inv_3[2] = ~div[2] /*2794*/;
  assign inv_3[3] = ~div[3] /*2793*/;
  assign inv_3[4] = ~div[4] /*2792*/;
  assign inv_3[5] = ~div[5] /*2791*/;
  assign inv_3[6] = ~div[6] /*2790*/;
  assign inv_3[7] = ~div[7] /*2789*/;
  assign inv_3[8] = ~div[8] /*2788*/;
  assign inv_3[9] = ~div[9] /*2787*/;
  assign inv_3[10] = ~div[10] /*2786*/;
assign inv_3[11] = oneWire /*2785*/;
  assign _168_ = inv_3[0] ^ r_2[9] /*2783*/;
  assign sum_3[0] = _168_ ^ oneWire /*2782*/;
  assign _169_ = _168_ & oneWire /*2781*/;
  assign _170_ = inv_3[0] & r_2[9] /*2780*/;
  assign _171_ = _169_ | _170_ /*2779*/;
  assign _172_ = inv_3[1] ^ r_2[10] /*2778*/;
  assign sum_3[1] = _172_ ^ _171_ /*2777*/;
  assign _173_ = _172_ & _171_ /*2776*/;
  assign _174_ = inv_3[1] & r_2[10] /*2775*/;
  assign _175_ = _173_ | _174_ /*2774*/;
  assign _176_ = inv_3[2] ^ r_2[11] /*2772*/;
  assign sum_3[2] = _176_ ^ _175_ /*2771*/;
  assign _177_ = _176_ & _175_ /*2770*/;
  assign _178_ = inv_3[2] & r_2[11] /*2769*/;
  assign _179_ = _177_ | _178_ /*2768*/;
  assign _180_ = inv_3[3] ^ r_2[12] /*2766*/;
  assign sum_3[3] = _180_ ^ _179_ /*2765*/;
  assign _181_ = _180_ & _179_ /*2764*/;
  assign _182_ = inv_3[3] & r_2[12] /*2763*/;
  assign _183_ = _181_ | _182_ /*2762*/;
  assign _184_ = inv_3[4] ^ r_2[13] /*2760*/;
  assign sum_3[4] = _184_ ^ _183_ /*2759*/;
  assign _185_ = _184_ & _183_ /*2758*/;
  assign _186_ = inv_3[4] & r_2[13] /*2757*/;
  assign _187_ = _185_ | _186_ /*2756*/;
  assign _188_ = inv_3[5] ^ r_2[14] /*2754*/;
  assign sum_3[5] = _188_ ^ _187_ /*2753*/;
  assign _189_ = _188_ & _187_ /*2752*/;
  assign _190_ = inv_3[5] & r_2[14] /*2751*/;
  assign _191_ = _189_ | _190_ /*2750*/;
  assign _192_ = inv_3[6] ^ r_2[15] /*2748*/;
  assign sum_3[6] = _192_ ^ _191_ /*2747*/;
  assign _193_ = _192_ & _191_ /*2746*/;
  assign _194_ = inv_3[6] & r_2[15] /*2745*/;
  assign _195_ = _193_ | _194_ /*2744*/;
  assign _196_ = inv_3[7] ^ r_2[16] /*2742*/;
  assign sum_3[7] = _196_ ^ _195_ /*2741*/;
  assign _197_ = _196_ & _195_ /*2740*/;
  assign _198_ = inv_3[7] & r_2[16] /*2739*/;
  assign _199_ = _197_ | _198_ /*2738*/;
  assign _200_ = inv_3[8] ^ r_2[17] /*2736*/;
  assign sum_3[8] = _200_ ^ _199_ /*2735*/;
  assign _201_ = _200_ & _199_ /*2734*/;
  assign _202_ = inv_3[8] & r_2[17] /*2733*/;
  assign _203_ = _201_ | _202_ /*2732*/;
  assign _204_ = inv_3[9] ^ r_2[18] /*2730*/;
  assign sum_3[9] = _204_ ^ _203_ /*2729*/;
  assign _205_ = _204_ & _203_ /*2728*/;
  assign _206_ = inv_3[9] & r_2[18] /*2727*/;
  assign _207_ = _205_ | _206_ /*2726*/;
  assign _208_ = inv_3[10] ^ r_2[19] /*2724*/;
  assign sum_3[10] = _208_ ^ _207_ /*2723*/;
  assign _209_ = _208_ & _207_ /*2722*/;
  assign _210_ = inv_3[10] & r_2[19] /*2721*/;
  assign _211_ = _209_ | _210_ /*2720*/;
  assign _212_ = inv_3[11] ^ r_2[20] /*2718*/;
  assign sum_3[11] = _212_ ^ _211_ /*2717*/;
  assign _213_ = _212_ & _211_ /*2716*/;
  assign _214_ = inv_3[11] & r_2[20] /*2715*/;
  assign _215_ = _213_ | _214_ /*2714*/;
  assign q[9] = ~sum_3[11] /*2721*/;
  assign m_3[0] = r_2[9] /*2720*/;
  assign m_3[1] = r_2[10] /*2719*/;
  assign m_3[2] = r_2[11] /*2718*/;
  assign m_3[3] = r_2[12] /*2717*/;
  assign m_3[4] = r_2[13] /*2716*/;
  assign m_3[5] = r_2[14] /*2715*/;
  assign m_3[6] = r_2[15] /*2714*/;
  assign m_3[7] = r_2[16] /*2713*/;
  assign m_3[8] = r_2[17] /*2712*/;
  assign m_3[9] = r_2[18] /*2711*/;
  assign m_3[10] = r_2[19] /*2710*/;
  assign m_3[11] = r_2[20] /*2709*/;
  assign _216_ = ~q[9] /*2707*/;
  assign _217_ = sum_3[0] & q[9] /*2706*/;
  assign _218_ = m_3[0] & _216_ /*2705*/;
  assign r_3[9] = _218_ | _217_ /*2704*/;
  assign _219_ = ~q[9] /*2703*/;
  assign _220_ = sum_3[1] & q[9] /*2702*/;
  assign _221_ = m_3[1] & _219_ /*2701*/;
  assign r_3[10] = _221_ | _220_ /*2700*/;
  assign _222_ = ~q[9] /*2699*/;
  assign _223_ = sum_3[2] & q[9] /*2698*/;
  assign _224_ = m_3[2] & _222_ /*2697*/;
  assign r_3[11] = _224_ | _223_ /*2696*/;
  assign _225_ = ~q[9] /*2695*/;
  assign _226_ = sum_3[3] & q[9] /*2694*/;
  assign _227_ = m_3[3] & _225_ /*2693*/;
  assign r_3[12] = _227_ | _226_ /*2692*/;
  assign _228_ = ~q[9] /*2691*/;
  assign _229_ = sum_3[4] & q[9] /*2690*/;
  assign _230_ = m_3[4] & _228_ /*2689*/;
  assign r_3[13] = _230_ | _229_ /*2688*/;
  assign _231_ = ~q[9] /*2687*/;
  assign _232_ = sum_3[5] & q[9] /*2686*/;
  assign _233_ = m_3[5] & _231_ /*2685*/;
  assign r_3[14] = _233_ | _232_ /*2684*/;
  assign _234_ = ~q[9] /*2683*/;
  assign _235_ = sum_3[6] & q[9] /*2682*/;
  assign _236_ = m_3[6] & _234_ /*2681*/;
  assign r_3[15] = _236_ | _235_ /*2680*/;
  assign _237_ = ~q[9] /*2679*/;
  assign _238_ = sum_3[7] & q[9] /*2678*/;
  assign _239_ = m_3[7] & _237_ /*2677*/;
  assign r_3[16] = _239_ | _238_ /*2676*/;
  assign _240_ = ~q[9] /*2675*/;
  assign _241_ = sum_3[8] & q[9] /*2674*/;
  assign _242_ = m_3[8] & _240_ /*2673*/;
  assign r_3[17] = _242_ | _241_ /*2672*/;
  assign _243_ = ~q[9] /*2671*/;
  assign _244_ = sum_3[9] & q[9] /*2670*/;
  assign _245_ = m_3[9] & _243_ /*2669*/;
  assign r_3[18] = _245_ | _244_ /*2668*/;
  assign _246_ = ~q[9] /*2667*/;
  assign _247_ = sum_3[10] & q[9] /*2666*/;
  assign _248_ = m_3[10] & _246_ /*2665*/;
  assign r_3[19] = _248_ | _247_ /*2664*/;
  assign _249_ = ~q[9] /*2663*/;
  assign _250_ = sum_3[11] & q[9] /*2662*/;
  assign _251_ = m_3[11] & _249_ /*2661*/;
  assign r_3[20] = _251_ | _250_ /*2660*/;
assign r_3[0]= r_2[0] /*2659*/;
assign r_3[1]= r_2[1] /*2658*/;
assign r_3[2]= r_2[2] /*2657*/;
assign r_3[3]= r_2[3] /*2656*/;
assign r_3[4]= r_2[4] /*2655*/;
assign r_3[5]= r_2[5] /*2654*/;
assign r_3[6]= r_2[6] /*2653*/;
assign r_3[7]= r_2[7] /*2652*/;
assign r_3[8]= r_2[8] /*2651*/;
  assign inv_4[0] = ~div[0] /*2628*/;
  assign inv_4[1] = ~div[1] /*2627*/;
  assign inv_4[2] = ~div[2] /*2626*/;
  assign inv_4[3] = ~div[3] /*2625*/;
  assign inv_4[4] = ~div[4] /*2624*/;
  assign inv_4[5] = ~div[5] /*2623*/;
  assign inv_4[6] = ~div[6] /*2622*/;
  assign inv_4[7] = ~div[7] /*2621*/;
  assign inv_4[8] = ~div[8] /*2620*/;
  assign inv_4[9] = ~div[9] /*2619*/;
  assign inv_4[10] = ~div[10] /*2618*/;
assign inv_4[11] = oneWire /*2617*/;
  assign _252_ = inv_4[0] ^ r_3[8] /*2615*/;
  assign sum_4[0] = _252_ ^ oneWire /*2614*/;
  assign _253_ = _252_ & oneWire /*2613*/;
  assign _254_ = inv_4[0] & r_3[8] /*2612*/;
  assign _255_ = _253_ | _254_ /*2611*/;
  assign _256_ = inv_4[1] ^ r_3[9] /*2610*/;
  assign sum_4[1] = _256_ ^ _255_ /*2609*/;
  assign _257_ = _256_ & _255_ /*2608*/;
  assign _258_ = inv_4[1] & r_3[9] /*2607*/;
  assign _259_ = _257_ | _258_ /*2606*/;
  assign _260_ = inv_4[2] ^ r_3[10] /*2604*/;
  assign sum_4[2] = _260_ ^ _259_ /*2603*/;
  assign _261_ = _260_ & _259_ /*2602*/;
  assign _262_ = inv_4[2] & r_3[10] /*2601*/;
  assign _263_ = _261_ | _262_ /*2600*/;
  assign _264_ = inv_4[3] ^ r_3[11] /*2598*/;
  assign sum_4[3] = _264_ ^ _263_ /*2597*/;
  assign _265_ = _264_ & _263_ /*2596*/;
  assign _266_ = inv_4[3] & r_3[11] /*2595*/;
  assign _267_ = _265_ | _266_ /*2594*/;
  assign _268_ = inv_4[4] ^ r_3[12] /*2592*/;
  assign sum_4[4] = _268_ ^ _267_ /*2591*/;
  assign _269_ = _268_ & _267_ /*2590*/;
  assign _270_ = inv_4[4] & r_3[12] /*2589*/;
  assign _271_ = _269_ | _270_ /*2588*/;
  assign _272_ = inv_4[5] ^ r_3[13] /*2586*/;
  assign sum_4[5] = _272_ ^ _271_ /*2585*/;
  assign _273_ = _272_ & _271_ /*2584*/;
  assign _274_ = inv_4[5] & r_3[13] /*2583*/;
  assign _275_ = _273_ | _274_ /*2582*/;
  assign _276_ = inv_4[6] ^ r_3[14] /*2580*/;
  assign sum_4[6] = _276_ ^ _275_ /*2579*/;
  assign _277_ = _276_ & _275_ /*2578*/;
  assign _278_ = inv_4[6] & r_3[14] /*2577*/;
  assign _279_ = _277_ | _278_ /*2576*/;
  assign _280_ = inv_4[7] ^ r_3[15] /*2574*/;
  assign sum_4[7] = _280_ ^ _279_ /*2573*/;
  assign _281_ = _280_ & _279_ /*2572*/;
  assign _282_ = inv_4[7] & r_3[15] /*2571*/;
  assign _283_ = _281_ | _282_ /*2570*/;
  assign _284_ = inv_4[8] ^ r_3[16] /*2568*/;
  assign sum_4[8] = _284_ ^ _283_ /*2567*/;
  assign _285_ = _284_ & _283_ /*2566*/;
  assign _286_ = inv_4[8] & r_3[16] /*2565*/;
  assign _287_ = _285_ | _286_ /*2564*/;
  assign _288_ = inv_4[9] ^ r_3[17] /*2562*/;
  assign sum_4[9] = _288_ ^ _287_ /*2561*/;
  assign _289_ = _288_ & _287_ /*2560*/;
  assign _290_ = inv_4[9] & r_3[17] /*2559*/;
  assign _291_ = _289_ | _290_ /*2558*/;
  assign _292_ = inv_4[10] ^ r_3[18] /*2556*/;
  assign sum_4[10] = _292_ ^ _291_ /*2555*/;
  assign _293_ = _292_ & _291_ /*2554*/;
  assign _294_ = inv_4[10] & r_3[18] /*2553*/;
  assign _295_ = _293_ | _294_ /*2552*/;
  assign _296_ = inv_4[11] ^ r_3[19] /*2550*/;
  assign sum_4[11] = _296_ ^ _295_ /*2549*/;
  assign _297_ = _296_ & _295_ /*2548*/;
  assign _298_ = inv_4[11] & r_3[19] /*2547*/;
  assign _299_ = _297_ | _298_ /*2546*/;
  assign q[8] = ~sum_4[11] /*2553*/;
  assign m_4[0] = r_3[8] /*2552*/;
  assign m_4[1] = r_3[9] /*2551*/;
  assign m_4[2] = r_3[10] /*2550*/;
  assign m_4[3] = r_3[11] /*2549*/;
  assign m_4[4] = r_3[12] /*2548*/;
  assign m_4[5] = r_3[13] /*2547*/;
  assign m_4[6] = r_3[14] /*2546*/;
  assign m_4[7] = r_3[15] /*2545*/;
  assign m_4[8] = r_3[16] /*2544*/;
  assign m_4[9] = r_3[17] /*2543*/;
  assign m_4[10] = r_3[18] /*2542*/;
  assign m_4[11] = r_3[19] /*2541*/;
  assign _300_ = ~q[8] /*2539*/;
  assign _301_ = sum_4[0] & q[8] /*2538*/;
  assign _302_ = m_4[0] & _300_ /*2537*/;
  assign r_4[8] = _302_ | _301_ /*2536*/;
  assign _303_ = ~q[8] /*2535*/;
  assign _304_ = sum_4[1] & q[8] /*2534*/;
  assign _305_ = m_4[1] & _303_ /*2533*/;
  assign r_4[9] = _305_ | _304_ /*2532*/;
  assign _306_ = ~q[8] /*2531*/;
  assign _307_ = sum_4[2] & q[8] /*2530*/;
  assign _308_ = m_4[2] & _306_ /*2529*/;
  assign r_4[10] = _308_ | _307_ /*2528*/;
  assign _309_ = ~q[8] /*2527*/;
  assign _310_ = sum_4[3] & q[8] /*2526*/;
  assign _311_ = m_4[3] & _309_ /*2525*/;
  assign r_4[11] = _311_ | _310_ /*2524*/;
  assign _312_ = ~q[8] /*2523*/;
  assign _313_ = sum_4[4] & q[8] /*2522*/;
  assign _314_ = m_4[4] & _312_ /*2521*/;
  assign r_4[12] = _314_ | _313_ /*2520*/;
  assign _315_ = ~q[8] /*2519*/;
  assign _316_ = sum_4[5] & q[8] /*2518*/;
  assign _317_ = m_4[5] & _315_ /*2517*/;
  assign r_4[13] = _317_ | _316_ /*2516*/;
  assign _318_ = ~q[8] /*2515*/;
  assign _319_ = sum_4[6] & q[8] /*2514*/;
  assign _320_ = m_4[6] & _318_ /*2513*/;
  assign r_4[14] = _320_ | _319_ /*2512*/;
  assign _321_ = ~q[8] /*2511*/;
  assign _322_ = sum_4[7] & q[8] /*2510*/;
  assign _323_ = m_4[7] & _321_ /*2509*/;
  assign r_4[15] = _323_ | _322_ /*2508*/;
  assign _324_ = ~q[8] /*2507*/;
  assign _325_ = sum_4[8] & q[8] /*2506*/;
  assign _326_ = m_4[8] & _324_ /*2505*/;
  assign r_4[16] = _326_ | _325_ /*2504*/;
  assign _327_ = ~q[8] /*2503*/;
  assign _328_ = sum_4[9] & q[8] /*2502*/;
  assign _329_ = m_4[9] & _327_ /*2501*/;
  assign r_4[17] = _329_ | _328_ /*2500*/;
  assign _330_ = ~q[8] /*2499*/;
  assign _331_ = sum_4[10] & q[8] /*2498*/;
  assign _332_ = m_4[10] & _330_ /*2497*/;
  assign r_4[18] = _332_ | _331_ /*2496*/;
  assign _333_ = ~q[8] /*2495*/;
  assign _334_ = sum_4[11] & q[8] /*2494*/;
  assign _335_ = m_4[11] & _333_ /*2493*/;
  assign r_4[19] = _335_ | _334_ /*2492*/;
assign r_4[0]= r_3[0] /*2491*/;
assign r_4[1]= r_3[1] /*2490*/;
assign r_4[2]= r_3[2] /*2489*/;
assign r_4[3]= r_3[3] /*2488*/;
assign r_4[4]= r_3[4] /*2487*/;
assign r_4[5]= r_3[5] /*2486*/;
assign r_4[6]= r_3[6] /*2485*/;
assign r_4[7]= r_3[7] /*2484*/;
  assign inv_5[0] = ~div[0] /*2460*/;
  assign inv_5[1] = ~div[1] /*2459*/;
  assign inv_5[2] = ~div[2] /*2458*/;
  assign inv_5[3] = ~div[3] /*2457*/;
  assign inv_5[4] = ~div[4] /*2456*/;
  assign inv_5[5] = ~div[5] /*2455*/;
  assign inv_5[6] = ~div[6] /*2454*/;
  assign inv_5[7] = ~div[7] /*2453*/;
  assign inv_5[8] = ~div[8] /*2452*/;
  assign inv_5[9] = ~div[9] /*2451*/;
  assign inv_5[10] = ~div[10] /*2450*/;
assign inv_5[11] = oneWire /*2449*/;
  assign _336_ = inv_5[0] ^ r_4[7] /*2447*/;
  assign sum_5[0] = _336_ ^ oneWire /*2446*/;
  assign _337_ = _336_ & oneWire /*2445*/;
  assign _338_ = inv_5[0] & r_4[7] /*2444*/;
  assign _339_ = _337_ | _338_ /*2443*/;
  assign _340_ = inv_5[1] ^ r_4[8] /*2442*/;
  assign sum_5[1] = _340_ ^ _339_ /*2441*/;
  assign _341_ = _340_ & _339_ /*2440*/;
  assign _342_ = inv_5[1] & r_4[8] /*2439*/;
  assign _343_ = _341_ | _342_ /*2438*/;
  assign _344_ = inv_5[2] ^ r_4[9] /*2436*/;
  assign sum_5[2] = _344_ ^ _343_ /*2435*/;
  assign _345_ = _344_ & _343_ /*2434*/;
  assign _346_ = inv_5[2] & r_4[9] /*2433*/;
  assign _347_ = _345_ | _346_ /*2432*/;
  assign _348_ = inv_5[3] ^ r_4[10] /*2430*/;
  assign sum_5[3] = _348_ ^ _347_ /*2429*/;
  assign _349_ = _348_ & _347_ /*2428*/;
  assign _350_ = inv_5[3] & r_4[10] /*2427*/;
  assign _351_ = _349_ | _350_ /*2426*/;
  assign _352_ = inv_5[4] ^ r_4[11] /*2424*/;
  assign sum_5[4] = _352_ ^ _351_ /*2423*/;
  assign _353_ = _352_ & _351_ /*2422*/;
  assign _354_ = inv_5[4] & r_4[11] /*2421*/;
  assign _355_ = _353_ | _354_ /*2420*/;
  assign _356_ = inv_5[5] ^ r_4[12] /*2418*/;
  assign sum_5[5] = _356_ ^ _355_ /*2417*/;
  assign _357_ = _356_ & _355_ /*2416*/;
  assign _358_ = inv_5[5] & r_4[12] /*2415*/;
  assign _359_ = _357_ | _358_ /*2414*/;
  assign _360_ = inv_5[6] ^ r_4[13] /*2412*/;
  assign sum_5[6] = _360_ ^ _359_ /*2411*/;
  assign _361_ = _360_ & _359_ /*2410*/;
  assign _362_ = inv_5[6] & r_4[13] /*2409*/;
  assign _363_ = _361_ | _362_ /*2408*/;
  assign _364_ = inv_5[7] ^ r_4[14] /*2406*/;
  assign sum_5[7] = _364_ ^ _363_ /*2405*/;
  assign _365_ = _364_ & _363_ /*2404*/;
  assign _366_ = inv_5[7] & r_4[14] /*2403*/;
  assign _367_ = _365_ | _366_ /*2402*/;
  assign _368_ = inv_5[8] ^ r_4[15] /*2400*/;
  assign sum_5[8] = _368_ ^ _367_ /*2399*/;
  assign _369_ = _368_ & _367_ /*2398*/;
  assign _370_ = inv_5[8] & r_4[15] /*2397*/;
  assign _371_ = _369_ | _370_ /*2396*/;
  assign _372_ = inv_5[9] ^ r_4[16] /*2394*/;
  assign sum_5[9] = _372_ ^ _371_ /*2393*/;
  assign _373_ = _372_ & _371_ /*2392*/;
  assign _374_ = inv_5[9] & r_4[16] /*2391*/;
  assign _375_ = _373_ | _374_ /*2390*/;
  assign _376_ = inv_5[10] ^ r_4[17] /*2388*/;
  assign sum_5[10] = _376_ ^ _375_ /*2387*/;
  assign _377_ = _376_ & _375_ /*2386*/;
  assign _378_ = inv_5[10] & r_4[17] /*2385*/;
  assign _379_ = _377_ | _378_ /*2384*/;
  assign _380_ = inv_5[11] ^ r_4[18] /*2382*/;
  assign sum_5[11] = _380_ ^ _379_ /*2381*/;
  assign _381_ = _380_ & _379_ /*2380*/;
  assign _382_ = inv_5[11] & r_4[18] /*2379*/;
  assign _383_ = _381_ | _382_ /*2378*/;
  assign q[7] = ~sum_5[11] /*2385*/;
  assign m_5[0] = r_4[7] /*2384*/;
  assign m_5[1] = r_4[8] /*2383*/;
  assign m_5[2] = r_4[9] /*2382*/;
  assign m_5[3] = r_4[10] /*2381*/;
  assign m_5[4] = r_4[11] /*2380*/;
  assign m_5[5] = r_4[12] /*2379*/;
  assign m_5[6] = r_4[13] /*2378*/;
  assign m_5[7] = r_4[14] /*2377*/;
  assign m_5[8] = r_4[15] /*2376*/;
  assign m_5[9] = r_4[16] /*2375*/;
  assign m_5[10] = r_4[17] /*2374*/;
  assign m_5[11] = r_4[18] /*2373*/;
  assign _384_ = ~q[7] /*2371*/;
  assign _385_ = sum_5[0] & q[7] /*2370*/;
  assign _386_ = m_5[0] & _384_ /*2369*/;
  assign r_5[7] = _386_ | _385_ /*2368*/;
  assign _387_ = ~q[7] /*2367*/;
  assign _388_ = sum_5[1] & q[7] /*2366*/;
  assign _389_ = m_5[1] & _387_ /*2365*/;
  assign r_5[8] = _389_ | _388_ /*2364*/;
  assign _390_ = ~q[7] /*2363*/;
  assign _391_ = sum_5[2] & q[7] /*2362*/;
  assign _392_ = m_5[2] & _390_ /*2361*/;
  assign r_5[9] = _392_ | _391_ /*2360*/;
  assign _393_ = ~q[7] /*2359*/;
  assign _394_ = sum_5[3] & q[7] /*2358*/;
  assign _395_ = m_5[3] & _393_ /*2357*/;
  assign r_5[10] = _395_ | _394_ /*2356*/;
  assign _396_ = ~q[7] /*2355*/;
  assign _397_ = sum_5[4] & q[7] /*2354*/;
  assign _398_ = m_5[4] & _396_ /*2353*/;
  assign r_5[11] = _398_ | _397_ /*2352*/;
  assign _399_ = ~q[7] /*2351*/;
  assign _400_ = sum_5[5] & q[7] /*2350*/;
  assign _401_ = m_5[5] & _399_ /*2349*/;
  assign r_5[12] = _401_ | _400_ /*2348*/;
  assign _402_ = ~q[7] /*2347*/;
  assign _403_ = sum_5[6] & q[7] /*2346*/;
  assign _404_ = m_5[6] & _402_ /*2345*/;
  assign r_5[13] = _404_ | _403_ /*2344*/;
  assign _405_ = ~q[7] /*2343*/;
  assign _406_ = sum_5[7] & q[7] /*2342*/;
  assign _407_ = m_5[7] & _405_ /*2341*/;
  assign r_5[14] = _407_ | _406_ /*2340*/;
  assign _408_ = ~q[7] /*2339*/;
  assign _409_ = sum_5[8] & q[7] /*2338*/;
  assign _410_ = m_5[8] & _408_ /*2337*/;
  assign r_5[15] = _410_ | _409_ /*2336*/;
  assign _411_ = ~q[7] /*2335*/;
  assign _412_ = sum_5[9] & q[7] /*2334*/;
  assign _413_ = m_5[9] & _411_ /*2333*/;
  assign r_5[16] = _413_ | _412_ /*2332*/;
  assign _414_ = ~q[7] /*2331*/;
  assign _415_ = sum_5[10] & q[7] /*2330*/;
  assign _416_ = m_5[10] & _414_ /*2329*/;
  assign r_5[17] = _416_ | _415_ /*2328*/;
  assign _417_ = ~q[7] /*2327*/;
  assign _418_ = sum_5[11] & q[7] /*2326*/;
  assign _419_ = m_5[11] & _417_ /*2325*/;
  assign r_5[18] = _419_ | _418_ /*2324*/;
assign r_5[0]= r_4[0] /*2323*/;
assign r_5[1]= r_4[1] /*2322*/;
assign r_5[2]= r_4[2] /*2321*/;
assign r_5[3]= r_4[3] /*2320*/;
assign r_5[4]= r_4[4] /*2319*/;
assign r_5[5]= r_4[5] /*2318*/;
assign r_5[6]= r_4[6] /*2317*/;
  assign inv_6[0] = ~div[0] /*2292*/;
  assign inv_6[1] = ~div[1] /*2291*/;
  assign inv_6[2] = ~div[2] /*2290*/;
  assign inv_6[3] = ~div[3] /*2289*/;
  assign inv_6[4] = ~div[4] /*2288*/;
  assign inv_6[5] = ~div[5] /*2287*/;
  assign inv_6[6] = ~div[6] /*2286*/;
  assign inv_6[7] = ~div[7] /*2285*/;
  assign inv_6[8] = ~div[8] /*2284*/;
  assign inv_6[9] = ~div[9] /*2283*/;
  assign inv_6[10] = ~div[10] /*2282*/;
assign inv_6[11] = oneWire /*2281*/;
  assign _420_ = inv_6[0] ^ r_5[6] /*2279*/;
  assign sum_6[0] = _420_ ^ oneWire /*2278*/;
  assign _421_ = _420_ & oneWire /*2277*/;
  assign _422_ = inv_6[0] & r_5[6] /*2276*/;
  assign _423_ = _421_ | _422_ /*2275*/;
  assign _424_ = inv_6[1] ^ r_5[7] /*2274*/;
  assign sum_6[1] = _424_ ^ _423_ /*2273*/;
  assign _425_ = _424_ & _423_ /*2272*/;
  assign _426_ = inv_6[1] & r_5[7] /*2271*/;
  assign _427_ = _425_ | _426_ /*2270*/;
  assign _428_ = inv_6[2] ^ r_5[8] /*2268*/;
  assign sum_6[2] = _428_ ^ _427_ /*2267*/;
  assign _429_ = _428_ & _427_ /*2266*/;
  assign _430_ = inv_6[2] & r_5[8] /*2265*/;
  assign _431_ = _429_ | _430_ /*2264*/;
  assign _432_ = inv_6[3] ^ r_5[9] /*2262*/;
  assign sum_6[3] = _432_ ^ _431_ /*2261*/;
  assign _433_ = _432_ & _431_ /*2260*/;
  assign _434_ = inv_6[3] & r_5[9] /*2259*/;
  assign _435_ = _433_ | _434_ /*2258*/;
  assign _436_ = inv_6[4] ^ r_5[10] /*2256*/;
  assign sum_6[4] = _436_ ^ _435_ /*2255*/;
  assign _437_ = _436_ & _435_ /*2254*/;
  assign _438_ = inv_6[4] & r_5[10] /*2253*/;
  assign _439_ = _437_ | _438_ /*2252*/;
  assign _440_ = inv_6[5] ^ r_5[11] /*2250*/;
  assign sum_6[5] = _440_ ^ _439_ /*2249*/;
  assign _441_ = _440_ & _439_ /*2248*/;
  assign _442_ = inv_6[5] & r_5[11] /*2247*/;
  assign _443_ = _441_ | _442_ /*2246*/;
  assign _444_ = inv_6[6] ^ r_5[12] /*2244*/;
  assign sum_6[6] = _444_ ^ _443_ /*2243*/;
  assign _445_ = _444_ & _443_ /*2242*/;
  assign _446_ = inv_6[6] & r_5[12] /*2241*/;
  assign _447_ = _445_ | _446_ /*2240*/;
  assign _448_ = inv_6[7] ^ r_5[13] /*2238*/;
  assign sum_6[7] = _448_ ^ _447_ /*2237*/;
  assign _449_ = _448_ & _447_ /*2236*/;
  assign _450_ = inv_6[7] & r_5[13] /*2235*/;
  assign _451_ = _449_ | _450_ /*2234*/;
  assign _452_ = inv_6[8] ^ r_5[14] /*2232*/;
  assign sum_6[8] = _452_ ^ _451_ /*2231*/;
  assign _453_ = _452_ & _451_ /*2230*/;
  assign _454_ = inv_6[8] & r_5[14] /*2229*/;
  assign _455_ = _453_ | _454_ /*2228*/;
  assign _456_ = inv_6[9] ^ r_5[15] /*2226*/;
  assign sum_6[9] = _456_ ^ _455_ /*2225*/;
  assign _457_ = _456_ & _455_ /*2224*/;
  assign _458_ = inv_6[9] & r_5[15] /*2223*/;
  assign _459_ = _457_ | _458_ /*2222*/;
  assign _460_ = inv_6[10] ^ r_5[16] /*2220*/;
  assign sum_6[10] = _460_ ^ _459_ /*2219*/;
  assign _461_ = _460_ & _459_ /*2218*/;
  assign _462_ = inv_6[10] & r_5[16] /*2217*/;
  assign _463_ = _461_ | _462_ /*2216*/;
  assign _464_ = inv_6[11] ^ r_5[17] /*2214*/;
  assign sum_6[11] = _464_ ^ _463_ /*2213*/;
  assign _465_ = _464_ & _463_ /*2212*/;
  assign _466_ = inv_6[11] & r_5[17] /*2211*/;
  assign _467_ = _465_ | _466_ /*2210*/;
  assign q[6] = ~sum_6[11] /*2217*/;
  assign m_6[0] = r_5[6] /*2216*/;
  assign m_6[1] = r_5[7] /*2215*/;
  assign m_6[2] = r_5[8] /*2214*/;
  assign m_6[3] = r_5[9] /*2213*/;
  assign m_6[4] = r_5[10] /*2212*/;
  assign m_6[5] = r_5[11] /*2211*/;
  assign m_6[6] = r_5[12] /*2210*/;
  assign m_6[7] = r_5[13] /*2209*/;
  assign m_6[8] = r_5[14] /*2208*/;
  assign m_6[9] = r_5[15] /*2207*/;
  assign m_6[10] = r_5[16] /*2206*/;
  assign m_6[11] = r_5[17] /*2205*/;
  assign _468_ = ~q[6] /*2203*/;
  assign _469_ = sum_6[0] & q[6] /*2202*/;
  assign _470_ = m_6[0] & _468_ /*2201*/;
  assign r_6[6] = _470_ | _469_ /*2200*/;
  assign _471_ = ~q[6] /*2199*/;
  assign _472_ = sum_6[1] & q[6] /*2198*/;
  assign _473_ = m_6[1] & _471_ /*2197*/;
  assign r_6[7] = _473_ | _472_ /*2196*/;
  assign _474_ = ~q[6] /*2195*/;
  assign _475_ = sum_6[2] & q[6] /*2194*/;
  assign _476_ = m_6[2] & _474_ /*2193*/;
  assign r_6[8] = _476_ | _475_ /*2192*/;
  assign _477_ = ~q[6] /*2191*/;
  assign _478_ = sum_6[3] & q[6] /*2190*/;
  assign _479_ = m_6[3] & _477_ /*2189*/;
  assign r_6[9] = _479_ | _478_ /*2188*/;
  assign _480_ = ~q[6] /*2187*/;
  assign _481_ = sum_6[4] & q[6] /*2186*/;
  assign _482_ = m_6[4] & _480_ /*2185*/;
  assign r_6[10] = _482_ | _481_ /*2184*/;
  assign _483_ = ~q[6] /*2183*/;
  assign _484_ = sum_6[5] & q[6] /*2182*/;
  assign _485_ = m_6[5] & _483_ /*2181*/;
  assign r_6[11] = _485_ | _484_ /*2180*/;
  assign _486_ = ~q[6] /*2179*/;
  assign _487_ = sum_6[6] & q[6] /*2178*/;
  assign _488_ = m_6[6] & _486_ /*2177*/;
  assign r_6[12] = _488_ | _487_ /*2176*/;
  assign _489_ = ~q[6] /*2175*/;
  assign _490_ = sum_6[7] & q[6] /*2174*/;
  assign _491_ = m_6[7] & _489_ /*2173*/;
  assign r_6[13] = _491_ | _490_ /*2172*/;
  assign _492_ = ~q[6] /*2171*/;
  assign _493_ = sum_6[8] & q[6] /*2170*/;
  assign _494_ = m_6[8] & _492_ /*2169*/;
  assign r_6[14] = _494_ | _493_ /*2168*/;
  assign _495_ = ~q[6] /*2167*/;
  assign _496_ = sum_6[9] & q[6] /*2166*/;
  assign _497_ = m_6[9] & _495_ /*2165*/;
  assign r_6[15] = _497_ | _496_ /*2164*/;
  assign _498_ = ~q[6] /*2163*/;
  assign _499_ = sum_6[10] & q[6] /*2162*/;
  assign _500_ = m_6[10] & _498_ /*2161*/;
  assign r_6[16] = _500_ | _499_ /*2160*/;
  assign _501_ = ~q[6] /*2159*/;
  assign _502_ = sum_6[11] & q[6] /*2158*/;
  assign _503_ = m_6[11] & _501_ /*2157*/;
  assign r_6[17] = _503_ | _502_ /*2156*/;
assign r_6[0]= r_5[0] /*2155*/;
assign r_6[1]= r_5[1] /*2154*/;
assign r_6[2]= r_5[2] /*2153*/;
assign r_6[3]= r_5[3] /*2152*/;
assign r_6[4]= r_5[4] /*2151*/;
assign r_6[5]= r_5[5] /*2150*/;
  assign inv_7[0] = ~div[0] /*2124*/;
  assign inv_7[1] = ~div[1] /*2123*/;
  assign inv_7[2] = ~div[2] /*2122*/;
  assign inv_7[3] = ~div[3] /*2121*/;
  assign inv_7[4] = ~div[4] /*2120*/;
  assign inv_7[5] = ~div[5] /*2119*/;
  assign inv_7[6] = ~div[6] /*2118*/;
  assign inv_7[7] = ~div[7] /*2117*/;
  assign inv_7[8] = ~div[8] /*2116*/;
  assign inv_7[9] = ~div[9] /*2115*/;
  assign inv_7[10] = ~div[10] /*2114*/;
assign inv_7[11] = oneWire /*2113*/;
  assign _504_ = inv_7[0] ^ r_6[5] /*2111*/;
  assign sum_7[0] = _504_ ^ oneWire /*2110*/;
  assign _505_ = _504_ & oneWire /*2109*/;
  assign _506_ = inv_7[0] & r_6[5] /*2108*/;
  assign _507_ = _505_ | _506_ /*2107*/;
  assign _508_ = inv_7[1] ^ r_6[6] /*2106*/;
  assign sum_7[1] = _508_ ^ _507_ /*2105*/;
  assign _509_ = _508_ & _507_ /*2104*/;
  assign _510_ = inv_7[1] & r_6[6] /*2103*/;
  assign _511_ = _509_ | _510_ /*2102*/;
  assign _512_ = inv_7[2] ^ r_6[7] /*2100*/;
  assign sum_7[2] = _512_ ^ _511_ /*2099*/;
  assign _513_ = _512_ & _511_ /*2098*/;
  assign _514_ = inv_7[2] & r_6[7] /*2097*/;
  assign _515_ = _513_ | _514_ /*2096*/;
  assign _516_ = inv_7[3] ^ r_6[8] /*2094*/;
  assign sum_7[3] = _516_ ^ _515_ /*2093*/;
  assign _517_ = _516_ & _515_ /*2092*/;
  assign _518_ = inv_7[3] & r_6[8] /*2091*/;
  assign _519_ = _517_ | _518_ /*2090*/;
  assign _520_ = inv_7[4] ^ r_6[9] /*2088*/;
  assign sum_7[4] = _520_ ^ _519_ /*2087*/;
  assign _521_ = _520_ & _519_ /*2086*/;
  assign _522_ = inv_7[4] & r_6[9] /*2085*/;
  assign _523_ = _521_ | _522_ /*2084*/;
  assign _524_ = inv_7[5] ^ r_6[10] /*2082*/;
  assign sum_7[5] = _524_ ^ _523_ /*2081*/;
  assign _525_ = _524_ & _523_ /*2080*/;
  assign _526_ = inv_7[5] & r_6[10] /*2079*/;
  assign _527_ = _525_ | _526_ /*2078*/;
  assign _528_ = inv_7[6] ^ r_6[11] /*2076*/;
  assign sum_7[6] = _528_ ^ _527_ /*2075*/;
  assign _529_ = _528_ & _527_ /*2074*/;
  assign _530_ = inv_7[6] & r_6[11] /*2073*/;
  assign _531_ = _529_ | _530_ /*2072*/;
  assign _532_ = inv_7[7] ^ r_6[12] /*2070*/;
  assign sum_7[7] = _532_ ^ _531_ /*2069*/;
  assign _533_ = _532_ & _531_ /*2068*/;
  assign _534_ = inv_7[7] & r_6[12] /*2067*/;
  assign _535_ = _533_ | _534_ /*2066*/;
  assign _536_ = inv_7[8] ^ r_6[13] /*2064*/;
  assign sum_7[8] = _536_ ^ _535_ /*2063*/;
  assign _537_ = _536_ & _535_ /*2062*/;
  assign _538_ = inv_7[8] & r_6[13] /*2061*/;
  assign _539_ = _537_ | _538_ /*2060*/;
  assign _540_ = inv_7[9] ^ r_6[14] /*2058*/;
  assign sum_7[9] = _540_ ^ _539_ /*2057*/;
  assign _541_ = _540_ & _539_ /*2056*/;
  assign _542_ = inv_7[9] & r_6[14] /*2055*/;
  assign _543_ = _541_ | _542_ /*2054*/;
  assign _544_ = inv_7[10] ^ r_6[15] /*2052*/;
  assign sum_7[10] = _544_ ^ _543_ /*2051*/;
  assign _545_ = _544_ & _543_ /*2050*/;
  assign _546_ = inv_7[10] & r_6[15] /*2049*/;
  assign _547_ = _545_ | _546_ /*2048*/;
  assign _548_ = inv_7[11] ^ r_6[16] /*2046*/;
  assign sum_7[11] = _548_ ^ _547_ /*2045*/;
  assign _549_ = _548_ & _547_ /*2044*/;
  assign _550_ = inv_7[11] & r_6[16] /*2043*/;
  assign _551_ = _549_ | _550_ /*2042*/;
  assign q[5] = ~sum_7[11] /*2049*/;
  assign m_7[0] = r_6[5] /*2048*/;
  assign m_7[1] = r_6[6] /*2047*/;
  assign m_7[2] = r_6[7] /*2046*/;
  assign m_7[3] = r_6[8] /*2045*/;
  assign m_7[4] = r_6[9] /*2044*/;
  assign m_7[5] = r_6[10] /*2043*/;
  assign m_7[6] = r_6[11] /*2042*/;
  assign m_7[7] = r_6[12] /*2041*/;
  assign m_7[8] = r_6[13] /*2040*/;
  assign m_7[9] = r_6[14] /*2039*/;
  assign m_7[10] = r_6[15] /*2038*/;
  assign m_7[11] = r_6[16] /*2037*/;
  assign _552_ = ~q[5] /*2035*/;
  assign _553_ = sum_7[0] & q[5] /*2034*/;
  assign _554_ = m_7[0] & _552_ /*2033*/;
  assign r_7[5] = _554_ | _553_ /*2032*/;
  assign _555_ = ~q[5] /*2031*/;
  assign _556_ = sum_7[1] & q[5] /*2030*/;
  assign _557_ = m_7[1] & _555_ /*2029*/;
  assign r_7[6] = _557_ | _556_ /*2028*/;
  assign _558_ = ~q[5] /*2027*/;
  assign _559_ = sum_7[2] & q[5] /*2026*/;
  assign _560_ = m_7[2] & _558_ /*2025*/;
  assign r_7[7] = _560_ | _559_ /*2024*/;
  assign _561_ = ~q[5] /*2023*/;
  assign _562_ = sum_7[3] & q[5] /*2022*/;
  assign _563_ = m_7[3] & _561_ /*2021*/;
  assign r_7[8] = _563_ | _562_ /*2020*/;
  assign _564_ = ~q[5] /*2019*/;
  assign _565_ = sum_7[4] & q[5] /*2018*/;
  assign _566_ = m_7[4] & _564_ /*2017*/;
  assign r_7[9] = _566_ | _565_ /*2016*/;
  assign _567_ = ~q[5] /*2015*/;
  assign _568_ = sum_7[5] & q[5] /*2014*/;
  assign _569_ = m_7[5] & _567_ /*2013*/;
  assign r_7[10] = _569_ | _568_ /*2012*/;
  assign _570_ = ~q[5] /*2011*/;
  assign _571_ = sum_7[6] & q[5] /*2010*/;
  assign _572_ = m_7[6] & _570_ /*2009*/;
  assign r_7[11] = _572_ | _571_ /*2008*/;
  assign _573_ = ~q[5] /*2007*/;
  assign _574_ = sum_7[7] & q[5] /*2006*/;
  assign _575_ = m_7[7] & _573_ /*2005*/;
  assign r_7[12] = _575_ | _574_ /*2004*/;
  assign _576_ = ~q[5] /*2003*/;
  assign _577_ = sum_7[8] & q[5] /*2002*/;
  assign _578_ = m_7[8] & _576_ /*2001*/;
  assign r_7[13] = _578_ | _577_ /*2000*/;
  assign _579_ = ~q[5] /*1999*/;
  assign _580_ = sum_7[9] & q[5] /*1998*/;
  assign _581_ = m_7[9] & _579_ /*1997*/;
  assign r_7[14] = _581_ | _580_ /*1996*/;
  assign _582_ = ~q[5] /*1995*/;
  assign _583_ = sum_7[10] & q[5] /*1994*/;
  assign _584_ = m_7[10] & _582_ /*1993*/;
  assign r_7[15] = _584_ | _583_ /*1992*/;
  assign _585_ = ~q[5] /*1991*/;
  assign _586_ = sum_7[11] & q[5] /*1990*/;
  assign _587_ = m_7[11] & _585_ /*1989*/;
  assign r_7[16] = _587_ | _586_ /*1988*/;
assign r_7[0]= r_6[0] /*1987*/;
assign r_7[1]= r_6[1] /*1986*/;
assign r_7[2]= r_6[2] /*1985*/;
assign r_7[3]= r_6[3] /*1984*/;
assign r_7[4]= r_6[4] /*1983*/;
  assign inv_8[0] = ~div[0] /*1956*/;
  assign inv_8[1] = ~div[1] /*1955*/;
  assign inv_8[2] = ~div[2] /*1954*/;
  assign inv_8[3] = ~div[3] /*1953*/;
  assign inv_8[4] = ~div[4] /*1952*/;
  assign inv_8[5] = ~div[5] /*1951*/;
  assign inv_8[6] = ~div[6] /*1950*/;
  assign inv_8[7] = ~div[7] /*1949*/;
  assign inv_8[8] = ~div[8] /*1948*/;
  assign inv_8[9] = ~div[9] /*1947*/;
  assign inv_8[10] = ~div[10] /*1946*/;
assign inv_8[11] = oneWire /*1945*/;
  assign _588_ = inv_8[0] ^ r_7[4] /*1943*/;
  assign sum_8[0] = _588_ ^ oneWire /*1942*/;
  assign _589_ = _588_ & oneWire /*1941*/;
  assign _590_ = inv_8[0] & r_7[4] /*1940*/;
  assign _591_ = _589_ | _590_ /*1939*/;
  assign _592_ = inv_8[1] ^ r_7[5] /*1938*/;
  assign sum_8[1] = _592_ ^ _591_ /*1937*/;
  assign _593_ = _592_ & _591_ /*1936*/;
  assign _594_ = inv_8[1] & r_7[5] /*1935*/;
  assign _595_ = _593_ | _594_ /*1934*/;
  assign _596_ = inv_8[2] ^ r_7[6] /*1932*/;
  assign sum_8[2] = _596_ ^ _595_ /*1931*/;
  assign _597_ = _596_ & _595_ /*1930*/;
  assign _598_ = inv_8[2] & r_7[6] /*1929*/;
  assign _599_ = _597_ | _598_ /*1928*/;
  assign _600_ = inv_8[3] ^ r_7[7] /*1926*/;
  assign sum_8[3] = _600_ ^ _599_ /*1925*/;
  assign _601_ = _600_ & _599_ /*1924*/;
  assign _602_ = inv_8[3] & r_7[7] /*1923*/;
  assign _603_ = _601_ | _602_ /*1922*/;
  assign _604_ = inv_8[4] ^ r_7[8] /*1920*/;
  assign sum_8[4] = _604_ ^ _603_ /*1919*/;
  assign _605_ = _604_ & _603_ /*1918*/;
  assign _606_ = inv_8[4] & r_7[8] /*1917*/;
  assign _607_ = _605_ | _606_ /*1916*/;
  assign _608_ = inv_8[5] ^ r_7[9] /*1914*/;
  assign sum_8[5] = _608_ ^ _607_ /*1913*/;
  assign _609_ = _608_ & _607_ /*1912*/;
  assign _610_ = inv_8[5] & r_7[9] /*1911*/;
  assign _611_ = _609_ | _610_ /*1910*/;
  assign _612_ = inv_8[6] ^ r_7[10] /*1908*/;
  assign sum_8[6] = _612_ ^ _611_ /*1907*/;
  assign _613_ = _612_ & _611_ /*1906*/;
  assign _614_ = inv_8[6] & r_7[10] /*1905*/;
  assign _615_ = _613_ | _614_ /*1904*/;
  assign _616_ = inv_8[7] ^ r_7[11] /*1902*/;
  assign sum_8[7] = _616_ ^ _615_ /*1901*/;
  assign _617_ = _616_ & _615_ /*1900*/;
  assign _618_ = inv_8[7] & r_7[11] /*1899*/;
  assign _619_ = _617_ | _618_ /*1898*/;
  assign _620_ = inv_8[8] ^ r_7[12] /*1896*/;
  assign sum_8[8] = _620_ ^ _619_ /*1895*/;
  assign _621_ = _620_ & _619_ /*1894*/;
  assign _622_ = inv_8[8] & r_7[12] /*1893*/;
  assign _623_ = _621_ | _622_ /*1892*/;
  assign _624_ = inv_8[9] ^ r_7[13] /*1890*/;
  assign sum_8[9] = _624_ ^ _623_ /*1889*/;
  assign _625_ = _624_ & _623_ /*1888*/;
  assign _626_ = inv_8[9] & r_7[13] /*1887*/;
  assign _627_ = _625_ | _626_ /*1886*/;
  assign _628_ = inv_8[10] ^ r_7[14] /*1884*/;
  assign sum_8[10] = _628_ ^ _627_ /*1883*/;
  assign _629_ = _628_ & _627_ /*1882*/;
  assign _630_ = inv_8[10] & r_7[14] /*1881*/;
  assign _631_ = _629_ | _630_ /*1880*/;
  assign _632_ = inv_8[11] ^ r_7[15] /*1878*/;
  assign sum_8[11] = _632_ ^ _631_ /*1877*/;
  assign _633_ = _632_ & _631_ /*1876*/;
  assign _634_ = inv_8[11] & r_7[15] /*1875*/;
  assign _635_ = _633_ | _634_ /*1874*/;
  assign q[4] = ~sum_8[11] /*1881*/;
  assign m_8[0] = r_7[4] /*1880*/;
  assign m_8[1] = r_7[5] /*1879*/;
  assign m_8[2] = r_7[6] /*1878*/;
  assign m_8[3] = r_7[7] /*1877*/;
  assign m_8[4] = r_7[8] /*1876*/;
  assign m_8[5] = r_7[9] /*1875*/;
  assign m_8[6] = r_7[10] /*1874*/;
  assign m_8[7] = r_7[11] /*1873*/;
  assign m_8[8] = r_7[12] /*1872*/;
  assign m_8[9] = r_7[13] /*1871*/;
  assign m_8[10] = r_7[14] /*1870*/;
  assign m_8[11] = r_7[15] /*1869*/;
  assign _636_ = ~q[4] /*1867*/;
  assign _637_ = sum_8[0] & q[4] /*1866*/;
  assign _638_ = m_8[0] & _636_ /*1865*/;
  assign r_8[4] = _638_ | _637_ /*1864*/;
  assign _639_ = ~q[4] /*1863*/;
  assign _640_ = sum_8[1] & q[4] /*1862*/;
  assign _641_ = m_8[1] & _639_ /*1861*/;
  assign r_8[5] = _641_ | _640_ /*1860*/;
  assign _642_ = ~q[4] /*1859*/;
  assign _643_ = sum_8[2] & q[4] /*1858*/;
  assign _644_ = m_8[2] & _642_ /*1857*/;
  assign r_8[6] = _644_ | _643_ /*1856*/;
  assign _645_ = ~q[4] /*1855*/;
  assign _646_ = sum_8[3] & q[4] /*1854*/;
  assign _647_ = m_8[3] & _645_ /*1853*/;
  assign r_8[7] = _647_ | _646_ /*1852*/;
  assign _648_ = ~q[4] /*1851*/;
  assign _649_ = sum_8[4] & q[4] /*1850*/;
  assign _650_ = m_8[4] & _648_ /*1849*/;
  assign r_8[8] = _650_ | _649_ /*1848*/;
  assign _651_ = ~q[4] /*1847*/;
  assign _652_ = sum_8[5] & q[4] /*1846*/;
  assign _653_ = m_8[5] & _651_ /*1845*/;
  assign r_8[9] = _653_ | _652_ /*1844*/;
  assign _654_ = ~q[4] /*1843*/;
  assign _655_ = sum_8[6] & q[4] /*1842*/;
  assign _656_ = m_8[6] & _654_ /*1841*/;
  assign r_8[10] = _656_ | _655_ /*1840*/;
  assign _657_ = ~q[4] /*1839*/;
  assign _658_ = sum_8[7] & q[4] /*1838*/;
  assign _659_ = m_8[7] & _657_ /*1837*/;
  assign r_8[11] = _659_ | _658_ /*1836*/;
  assign _660_ = ~q[4] /*1835*/;
  assign _661_ = sum_8[8] & q[4] /*1834*/;
  assign _662_ = m_8[8] & _660_ /*1833*/;
  assign r_8[12] = _662_ | _661_ /*1832*/;
  assign _663_ = ~q[4] /*1831*/;
  assign _664_ = sum_8[9] & q[4] /*1830*/;
  assign _665_ = m_8[9] & _663_ /*1829*/;
  assign r_8[13] = _665_ | _664_ /*1828*/;
  assign _666_ = ~q[4] /*1827*/;
  assign _667_ = sum_8[10] & q[4] /*1826*/;
  assign _668_ = m_8[10] & _666_ /*1825*/;
  assign r_8[14] = _668_ | _667_ /*1824*/;
  assign _669_ = ~q[4] /*1823*/;
  assign _670_ = sum_8[11] & q[4] /*1822*/;
  assign _671_ = m_8[11] & _669_ /*1821*/;
  assign r_8[15] = _671_ | _670_ /*1820*/;
assign r_8[0]= r_7[0] /*1819*/;
assign r_8[1]= r_7[1] /*1818*/;
assign r_8[2]= r_7[2] /*1817*/;
assign r_8[3]= r_7[3] /*1816*/;
  assign inv_9[0] = ~div[0] /*1788*/;
  assign inv_9[1] = ~div[1] /*1787*/;
  assign inv_9[2] = ~div[2] /*1786*/;
  assign inv_9[3] = ~div[3] /*1785*/;
  assign inv_9[4] = ~div[4] /*1784*/;
  assign inv_9[5] = ~div[5] /*1783*/;
  assign inv_9[6] = ~div[6] /*1782*/;
  assign inv_9[7] = ~div[7] /*1781*/;
  assign inv_9[8] = ~div[8] /*1780*/;
  assign inv_9[9] = ~div[9] /*1779*/;
  assign inv_9[10] = ~div[10] /*1778*/;
assign inv_9[11] = oneWire /*1777*/;
  assign _672_ = inv_9[0] ^ r_8[3] /*1775*/;
  assign sum_9[0] = _672_ ^ oneWire /*1774*/;
  assign _673_ = _672_ & oneWire /*1773*/;
  assign _674_ = inv_9[0] & r_8[3] /*1772*/;
  assign _675_ = _673_ | _674_ /*1771*/;
  assign _676_ = inv_9[1] ^ r_8[4] /*1770*/;
  assign sum_9[1] = _676_ ^ _675_ /*1769*/;
  assign _677_ = _676_ & _675_ /*1768*/;
  assign _678_ = inv_9[1] & r_8[4] /*1767*/;
  assign _679_ = _677_ | _678_ /*1766*/;
  assign _680_ = inv_9[2] ^ r_8[5] /*1764*/;
  assign sum_9[2] = _680_ ^ _679_ /*1763*/;
  assign _681_ = _680_ & _679_ /*1762*/;
  assign _682_ = inv_9[2] & r_8[5] /*1761*/;
  assign _683_ = _681_ | _682_ /*1760*/;
  assign _684_ = inv_9[3] ^ r_8[6] /*1758*/;
  assign sum_9[3] = _684_ ^ _683_ /*1757*/;
  assign _685_ = _684_ & _683_ /*1756*/;
  assign _686_ = inv_9[3] & r_8[6] /*1755*/;
  assign _687_ = _685_ | _686_ /*1754*/;
  assign _688_ = inv_9[4] ^ r_8[7] /*1752*/;
  assign sum_9[4] = _688_ ^ _687_ /*1751*/;
  assign _689_ = _688_ & _687_ /*1750*/;
  assign _690_ = inv_9[4] & r_8[7] /*1749*/;
  assign _691_ = _689_ | _690_ /*1748*/;
  assign _692_ = inv_9[5] ^ r_8[8] /*1746*/;
  assign sum_9[5] = _692_ ^ _691_ /*1745*/;
  assign _693_ = _692_ & _691_ /*1744*/;
  assign _694_ = inv_9[5] & r_8[8] /*1743*/;
  assign _695_ = _693_ | _694_ /*1742*/;
  assign _696_ = inv_9[6] ^ r_8[9] /*1740*/;
  assign sum_9[6] = _696_ ^ _695_ /*1739*/;
  assign _697_ = _696_ & _695_ /*1738*/;
  assign _698_ = inv_9[6] & r_8[9] /*1737*/;
  assign _699_ = _697_ | _698_ /*1736*/;
  assign _700_ = inv_9[7] ^ r_8[10] /*1734*/;
  assign sum_9[7] = _700_ ^ _699_ /*1733*/;
  assign _701_ = _700_ & _699_ /*1732*/;
  assign _702_ = inv_9[7] & r_8[10] /*1731*/;
  assign _703_ = _701_ | _702_ /*1730*/;
  assign _704_ = inv_9[8] ^ r_8[11] /*1728*/;
  assign sum_9[8] = _704_ ^ _703_ /*1727*/;
  assign _705_ = _704_ & _703_ /*1726*/;
  assign _706_ = inv_9[8] & r_8[11] /*1725*/;
  assign _707_ = _705_ | _706_ /*1724*/;
  assign _708_ = inv_9[9] ^ r_8[12] /*1722*/;
  assign sum_9[9] = _708_ ^ _707_ /*1721*/;
  assign _709_ = _708_ & _707_ /*1720*/;
  assign _710_ = inv_9[9] & r_8[12] /*1719*/;
  assign _711_ = _709_ | _710_ /*1718*/;
  assign _712_ = inv_9[10] ^ r_8[13] /*1716*/;
  assign sum_9[10] = _712_ ^ _711_ /*1715*/;
  assign _713_ = _712_ & _711_ /*1714*/;
  assign _714_ = inv_9[10] & r_8[13] /*1713*/;
  assign _715_ = _713_ | _714_ /*1712*/;
  assign _716_ = inv_9[11] ^ r_8[14] /*1710*/;
  assign sum_9[11] = _716_ ^ _715_ /*1709*/;
  assign _717_ = _716_ & _715_ /*1708*/;
  assign _718_ = inv_9[11] & r_8[14] /*1707*/;
  assign _719_ = _717_ | _718_ /*1706*/;
  assign q[3] = ~sum_9[11] /*1713*/;
  assign m_9[0] = r_8[3] /*1712*/;
  assign m_9[1] = r_8[4] /*1711*/;
  assign m_9[2] = r_8[5] /*1710*/;
  assign m_9[3] = r_8[6] /*1709*/;
  assign m_9[4] = r_8[7] /*1708*/;
  assign m_9[5] = r_8[8] /*1707*/;
  assign m_9[6] = r_8[9] /*1706*/;
  assign m_9[7] = r_8[10] /*1705*/;
  assign m_9[8] = r_8[11] /*1704*/;
  assign m_9[9] = r_8[12] /*1703*/;
  assign m_9[10] = r_8[13] /*1702*/;
  assign m_9[11] = r_8[14] /*1701*/;
  assign _720_ = ~q[3] /*1699*/;
  assign _721_ = sum_9[0] & q[3] /*1698*/;
  assign _722_ = m_9[0] & _720_ /*1697*/;
  assign r_9[3] = _722_ | _721_ /*1696*/;
  assign _723_ = ~q[3] /*1695*/;
  assign _724_ = sum_9[1] & q[3] /*1694*/;
  assign _725_ = m_9[1] & _723_ /*1693*/;
  assign r_9[4] = _725_ | _724_ /*1692*/;
  assign _726_ = ~q[3] /*1691*/;
  assign _727_ = sum_9[2] & q[3] /*1690*/;
  assign _728_ = m_9[2] & _726_ /*1689*/;
  assign r_9[5] = _728_ | _727_ /*1688*/;
  assign _729_ = ~q[3] /*1687*/;
  assign _730_ = sum_9[3] & q[3] /*1686*/;
  assign _731_ = m_9[3] & _729_ /*1685*/;
  assign r_9[6] = _731_ | _730_ /*1684*/;
  assign _732_ = ~q[3] /*1683*/;
  assign _733_ = sum_9[4] & q[3] /*1682*/;
  assign _734_ = m_9[4] & _732_ /*1681*/;
  assign r_9[7] = _734_ | _733_ /*1680*/;
  assign _735_ = ~q[3] /*1679*/;
  assign _736_ = sum_9[5] & q[3] /*1678*/;
  assign _737_ = m_9[5] & _735_ /*1677*/;
  assign r_9[8] = _737_ | _736_ /*1676*/;
  assign _738_ = ~q[3] /*1675*/;
  assign _739_ = sum_9[6] & q[3] /*1674*/;
  assign _740_ = m_9[6] & _738_ /*1673*/;
  assign r_9[9] = _740_ | _739_ /*1672*/;
  assign _741_ = ~q[3] /*1671*/;
  assign _742_ = sum_9[7] & q[3] /*1670*/;
  assign _743_ = m_9[7] & _741_ /*1669*/;
  assign r_9[10] = _743_ | _742_ /*1668*/;
  assign _744_ = ~q[3] /*1667*/;
  assign _745_ = sum_9[8] & q[3] /*1666*/;
  assign _746_ = m_9[8] & _744_ /*1665*/;
  assign r_9[11] = _746_ | _745_ /*1664*/;
  assign _747_ = ~q[3] /*1663*/;
  assign _748_ = sum_9[9] & q[3] /*1662*/;
  assign _749_ = m_9[9] & _747_ /*1661*/;
  assign r_9[12] = _749_ | _748_ /*1660*/;
  assign _750_ = ~q[3] /*1659*/;
  assign _751_ = sum_9[10] & q[3] /*1658*/;
  assign _752_ = m_9[10] & _750_ /*1657*/;
  assign r_9[13] = _752_ | _751_ /*1656*/;
  assign _753_ = ~q[3] /*1655*/;
  assign _754_ = sum_9[11] & q[3] /*1654*/;
  assign _755_ = m_9[11] & _753_ /*1653*/;
  assign r_9[14] = _755_ | _754_ /*1652*/;
assign r_9[0]= r_8[0] /*1651*/;
assign r_9[1]= r_8[1] /*1650*/;
assign r_9[2]= r_8[2] /*1649*/;
  assign inv_10[0] = ~div[0] /*1620*/;
  assign inv_10[1] = ~div[1] /*1619*/;
  assign inv_10[2] = ~div[2] /*1618*/;
  assign inv_10[3] = ~div[3] /*1617*/;
  assign inv_10[4] = ~div[4] /*1616*/;
  assign inv_10[5] = ~div[5] /*1615*/;
  assign inv_10[6] = ~div[6] /*1614*/;
  assign inv_10[7] = ~div[7] /*1613*/;
  assign inv_10[8] = ~div[8] /*1612*/;
  assign inv_10[9] = ~div[9] /*1611*/;
  assign inv_10[10] = ~div[10] /*1610*/;
assign inv_10[11] = oneWire /*1609*/;
  assign _756_ = inv_10[0] ^ r_9[2] /*1607*/;
  assign sum_10[0] = _756_ ^ oneWire /*1606*/;
  assign _757_ = _756_ & oneWire /*1605*/;
  assign _758_ = inv_10[0] & r_9[2] /*1604*/;
  assign _759_ = _757_ | _758_ /*1603*/;
  assign _760_ = inv_10[1] ^ r_9[3] /*1602*/;
  assign sum_10[1] = _760_ ^ _759_ /*1601*/;
  assign _761_ = _760_ & _759_ /*1600*/;
  assign _762_ = inv_10[1] & r_9[3] /*1599*/;
  assign _763_ = _761_ | _762_ /*1598*/;
  assign _764_ = inv_10[2] ^ r_9[4] /*1596*/;
  assign sum_10[2] = _764_ ^ _763_ /*1595*/;
  assign _765_ = _764_ & _763_ /*1594*/;
  assign _766_ = inv_10[2] & r_9[4] /*1593*/;
  assign _767_ = _765_ | _766_ /*1592*/;
  assign _768_ = inv_10[3] ^ r_9[5] /*1590*/;
  assign sum_10[3] = _768_ ^ _767_ /*1589*/;
  assign _769_ = _768_ & _767_ /*1588*/;
  assign _770_ = inv_10[3] & r_9[5] /*1587*/;
  assign _771_ = _769_ | _770_ /*1586*/;
  assign _772_ = inv_10[4] ^ r_9[6] /*1584*/;
  assign sum_10[4] = _772_ ^ _771_ /*1583*/;
  assign _773_ = _772_ & _771_ /*1582*/;
  assign _774_ = inv_10[4] & r_9[6] /*1581*/;
  assign _775_ = _773_ | _774_ /*1580*/;
  assign _776_ = inv_10[5] ^ r_9[7] /*1578*/;
  assign sum_10[5] = _776_ ^ _775_ /*1577*/;
  assign _777_ = _776_ & _775_ /*1576*/;
  assign _778_ = inv_10[5] & r_9[7] /*1575*/;
  assign _779_ = _777_ | _778_ /*1574*/;
  assign _780_ = inv_10[6] ^ r_9[8] /*1572*/;
  assign sum_10[6] = _780_ ^ _779_ /*1571*/;
  assign _781_ = _780_ & _779_ /*1570*/;
  assign _782_ = inv_10[6] & r_9[8] /*1569*/;
  assign _783_ = _781_ | _782_ /*1568*/;
  assign _784_ = inv_10[7] ^ r_9[9] /*1566*/;
  assign sum_10[7] = _784_ ^ _783_ /*1565*/;
  assign _785_ = _784_ & _783_ /*1564*/;
  assign _786_ = inv_10[7] & r_9[9] /*1563*/;
  assign _787_ = _785_ | _786_ /*1562*/;
  assign _788_ = inv_10[8] ^ r_9[10] /*1560*/;
  assign sum_10[8] = _788_ ^ _787_ /*1559*/;
  assign _789_ = _788_ & _787_ /*1558*/;
  assign _790_ = inv_10[8] & r_9[10] /*1557*/;
  assign _791_ = _789_ | _790_ /*1556*/;
  assign _792_ = inv_10[9] ^ r_9[11] /*1554*/;
  assign sum_10[9] = _792_ ^ _791_ /*1553*/;
  assign _793_ = _792_ & _791_ /*1552*/;
  assign _794_ = inv_10[9] & r_9[11] /*1551*/;
  assign _795_ = _793_ | _794_ /*1550*/;
  assign _796_ = inv_10[10] ^ r_9[12] /*1548*/;
  assign sum_10[10] = _796_ ^ _795_ /*1547*/;
  assign _797_ = _796_ & _795_ /*1546*/;
  assign _798_ = inv_10[10] & r_9[12] /*1545*/;
  assign _799_ = _797_ | _798_ /*1544*/;
  assign _800_ = inv_10[11] ^ r_9[13] /*1542*/;
  assign sum_10[11] = _800_ ^ _799_ /*1541*/;
  assign _801_ = _800_ & _799_ /*1540*/;
  assign _802_ = inv_10[11] & r_9[13] /*1539*/;
  assign _803_ = _801_ | _802_ /*1538*/;
  assign q[2] = ~sum_10[11] /*1545*/;
  assign m_10[0] = r_9[2] /*1544*/;
  assign m_10[1] = r_9[3] /*1543*/;
  assign m_10[2] = r_9[4] /*1542*/;
  assign m_10[3] = r_9[5] /*1541*/;
  assign m_10[4] = r_9[6] /*1540*/;
  assign m_10[5] = r_9[7] /*1539*/;
  assign m_10[6] = r_9[8] /*1538*/;
  assign m_10[7] = r_9[9] /*1537*/;
  assign m_10[8] = r_9[10] /*1536*/;
  assign m_10[9] = r_9[11] /*1535*/;
  assign m_10[10] = r_9[12] /*1534*/;
  assign m_10[11] = r_9[13] /*1533*/;
  assign _804_ = ~q[2] /*1531*/;
  assign _805_ = sum_10[0] & q[2] /*1530*/;
  assign _806_ = m_10[0] & _804_ /*1529*/;
  assign r_10[2] = _806_ | _805_ /*1528*/;
  assign _807_ = ~q[2] /*1527*/;
  assign _808_ = sum_10[1] & q[2] /*1526*/;
  assign _809_ = m_10[1] & _807_ /*1525*/;
  assign r_10[3] = _809_ | _808_ /*1524*/;
  assign _810_ = ~q[2] /*1523*/;
  assign _811_ = sum_10[2] & q[2] /*1522*/;
  assign _812_ = m_10[2] & _810_ /*1521*/;
  assign r_10[4] = _812_ | _811_ /*1520*/;
  assign _813_ = ~q[2] /*1519*/;
  assign _814_ = sum_10[3] & q[2] /*1518*/;
  assign _815_ = m_10[3] & _813_ /*1517*/;
  assign r_10[5] = _815_ | _814_ /*1516*/;
  assign _816_ = ~q[2] /*1515*/;
  assign _817_ = sum_10[4] & q[2] /*1514*/;
  assign _818_ = m_10[4] & _816_ /*1513*/;
  assign r_10[6] = _818_ | _817_ /*1512*/;
  assign _819_ = ~q[2] /*1511*/;
  assign _820_ = sum_10[5] & q[2] /*1510*/;
  assign _821_ = m_10[5] & _819_ /*1509*/;
  assign r_10[7] = _821_ | _820_ /*1508*/;
  assign _822_ = ~q[2] /*1507*/;
  assign _823_ = sum_10[6] & q[2] /*1506*/;
  assign _824_ = m_10[6] & _822_ /*1505*/;
  assign r_10[8] = _824_ | _823_ /*1504*/;
  assign _825_ = ~q[2] /*1503*/;
  assign _826_ = sum_10[7] & q[2] /*1502*/;
  assign _827_ = m_10[7] & _825_ /*1501*/;
  assign r_10[9] = _827_ | _826_ /*1500*/;
  assign _828_ = ~q[2] /*1499*/;
  assign _829_ = sum_10[8] & q[2] /*1498*/;
  assign _830_ = m_10[8] & _828_ /*1497*/;
  assign r_10[10] = _830_ | _829_ /*1496*/;
  assign _831_ = ~q[2] /*1495*/;
  assign _832_ = sum_10[9] & q[2] /*1494*/;
  assign _833_ = m_10[9] & _831_ /*1493*/;
  assign r_10[11] = _833_ | _832_ /*1492*/;
  assign _834_ = ~q[2] /*1491*/;
  assign _835_ = sum_10[10] & q[2] /*1490*/;
  assign _836_ = m_10[10] & _834_ /*1489*/;
  assign r_10[12] = _836_ | _835_ /*1488*/;
  assign _837_ = ~q[2] /*1487*/;
  assign _838_ = sum_10[11] & q[2] /*1486*/;
  assign _839_ = m_10[11] & _837_ /*1485*/;
  assign r_10[13] = _839_ | _838_ /*1484*/;
assign r_10[0]= r_9[0] /*1483*/;
assign r_10[1]= r_9[1] /*1482*/;
  assign inv_11[0] = ~div[0] /*1452*/;
  assign inv_11[1] = ~div[1] /*1451*/;
  assign inv_11[2] = ~div[2] /*1450*/;
  assign inv_11[3] = ~div[3] /*1449*/;
  assign inv_11[4] = ~div[4] /*1448*/;
  assign inv_11[5] = ~div[5] /*1447*/;
  assign inv_11[6] = ~div[6] /*1446*/;
  assign inv_11[7] = ~div[7] /*1445*/;
  assign inv_11[8] = ~div[8] /*1444*/;
  assign inv_11[9] = ~div[9] /*1443*/;
  assign inv_11[10] = ~div[10] /*1442*/;
assign inv_11[11] = oneWire /*1441*/;
  assign _840_ = inv_11[0] ^ r_10[1] /*1439*/;
  assign sum_11[0] = _840_ ^ oneWire /*1438*/;
  assign _841_ = _840_ & oneWire /*1437*/;
  assign _842_ = inv_11[0] & r_10[1] /*1436*/;
  assign _843_ = _841_ | _842_ /*1435*/;
  assign _844_ = inv_11[1] ^ r_10[2] /*1434*/;
  assign sum_11[1] = _844_ ^ _843_ /*1433*/;
  assign _845_ = _844_ & _843_ /*1432*/;
  assign _846_ = inv_11[1] & r_10[2] /*1431*/;
  assign _847_ = _845_ | _846_ /*1430*/;
  assign _848_ = inv_11[2] ^ r_10[3] /*1428*/;
  assign sum_11[2] = _848_ ^ _847_ /*1427*/;
  assign _849_ = _848_ & _847_ /*1426*/;
  assign _850_ = inv_11[2] & r_10[3] /*1425*/;
  assign _851_ = _849_ | _850_ /*1424*/;
  assign _852_ = inv_11[3] ^ r_10[4] /*1422*/;
  assign sum_11[3] = _852_ ^ _851_ /*1421*/;
  assign _853_ = _852_ & _851_ /*1420*/;
  assign _854_ = inv_11[3] & r_10[4] /*1419*/;
  assign _855_ = _853_ | _854_ /*1418*/;
  assign _856_ = inv_11[4] ^ r_10[5] /*1416*/;
  assign sum_11[4] = _856_ ^ _855_ /*1415*/;
  assign _857_ = _856_ & _855_ /*1414*/;
  assign _858_ = inv_11[4] & r_10[5] /*1413*/;
  assign _859_ = _857_ | _858_ /*1412*/;
  assign _860_ = inv_11[5] ^ r_10[6] /*1410*/;
  assign sum_11[5] = _860_ ^ _859_ /*1409*/;
  assign _861_ = _860_ & _859_ /*1408*/;
  assign _862_ = inv_11[5] & r_10[6] /*1407*/;
  assign _863_ = _861_ | _862_ /*1406*/;
  assign _864_ = inv_11[6] ^ r_10[7] /*1404*/;
  assign sum_11[6] = _864_ ^ _863_ /*1403*/;
  assign _865_ = _864_ & _863_ /*1402*/;
  assign _866_ = inv_11[6] & r_10[7] /*1401*/;
  assign _867_ = _865_ | _866_ /*1400*/;
  assign _868_ = inv_11[7] ^ r_10[8] /*1398*/;
  assign sum_11[7] = _868_ ^ _867_ /*1397*/;
  assign _869_ = _868_ & _867_ /*1396*/;
  assign _870_ = inv_11[7] & r_10[8] /*1395*/;
  assign _871_ = _869_ | _870_ /*1394*/;
  assign _872_ = inv_11[8] ^ r_10[9] /*1392*/;
  assign sum_11[8] = _872_ ^ _871_ /*1391*/;
  assign _873_ = _872_ & _871_ /*1390*/;
  assign _874_ = inv_11[8] & r_10[9] /*1389*/;
  assign _875_ = _873_ | _874_ /*1388*/;
  assign _876_ = inv_11[9] ^ r_10[10] /*1386*/;
  assign sum_11[9] = _876_ ^ _875_ /*1385*/;
  assign _877_ = _876_ & _875_ /*1384*/;
  assign _878_ = inv_11[9] & r_10[10] /*1383*/;
  assign _879_ = _877_ | _878_ /*1382*/;
  assign _880_ = inv_11[10] ^ r_10[11] /*1380*/;
  assign sum_11[10] = _880_ ^ _879_ /*1379*/;
  assign _881_ = _880_ & _879_ /*1378*/;
  assign _882_ = inv_11[10] & r_10[11] /*1377*/;
  assign _883_ = _881_ | _882_ /*1376*/;
  assign _884_ = inv_11[11] ^ r_10[12] /*1374*/;
  assign sum_11[11] = _884_ ^ _883_ /*1373*/;
  assign _885_ = _884_ & _883_ /*1372*/;
  assign _886_ = inv_11[11] & r_10[12] /*1371*/;
  assign _887_ = _885_ | _886_ /*1370*/;
  assign q[1] = ~sum_11[11] /*1377*/;
  assign m_11[0] = r_10[1] /*1376*/;
  assign m_11[1] = r_10[2] /*1375*/;
  assign m_11[2] = r_10[3] /*1374*/;
  assign m_11[3] = r_10[4] /*1373*/;
  assign m_11[4] = r_10[5] /*1372*/;
  assign m_11[5] = r_10[6] /*1371*/;
  assign m_11[6] = r_10[7] /*1370*/;
  assign m_11[7] = r_10[8] /*1369*/;
  assign m_11[8] = r_10[9] /*1368*/;
  assign m_11[9] = r_10[10] /*1367*/;
  assign m_11[10] = r_10[11] /*1366*/;
  assign m_11[11] = r_10[12] /*1365*/;
  assign _888_ = ~q[1] /*1363*/;
  assign _889_ = sum_11[0] & q[1] /*1362*/;
  assign _890_ = m_11[0] & _888_ /*1361*/;
  assign r_11[1] = _890_ | _889_ /*1360*/;
  assign _891_ = ~q[1] /*1359*/;
  assign _892_ = sum_11[1] & q[1] /*1358*/;
  assign _893_ = m_11[1] & _891_ /*1357*/;
  assign r_11[2] = _893_ | _892_ /*1356*/;
  assign _894_ = ~q[1] /*1355*/;
  assign _895_ = sum_11[2] & q[1] /*1354*/;
  assign _896_ = m_11[2] & _894_ /*1353*/;
  assign r_11[3] = _896_ | _895_ /*1352*/;
  assign _897_ = ~q[1] /*1351*/;
  assign _898_ = sum_11[3] & q[1] /*1350*/;
  assign _899_ = m_11[3] & _897_ /*1349*/;
  assign r_11[4] = _899_ | _898_ /*1348*/;
  assign _900_ = ~q[1] /*1347*/;
  assign _901_ = sum_11[4] & q[1] /*1346*/;
  assign _902_ = m_11[4] & _900_ /*1345*/;
  assign r_11[5] = _902_ | _901_ /*1344*/;
  assign _903_ = ~q[1] /*1343*/;
  assign _904_ = sum_11[5] & q[1] /*1342*/;
  assign _905_ = m_11[5] & _903_ /*1341*/;
  assign r_11[6] = _905_ | _904_ /*1340*/;
  assign _906_ = ~q[1] /*1339*/;
  assign _907_ = sum_11[6] & q[1] /*1338*/;
  assign _908_ = m_11[6] & _906_ /*1337*/;
  assign r_11[7] = _908_ | _907_ /*1336*/;
  assign _909_ = ~q[1] /*1335*/;
  assign _910_ = sum_11[7] & q[1] /*1334*/;
  assign _911_ = m_11[7] & _909_ /*1333*/;
  assign r_11[8] = _911_ | _910_ /*1332*/;
  assign _912_ = ~q[1] /*1331*/;
  assign _913_ = sum_11[8] & q[1] /*1330*/;
  assign _914_ = m_11[8] & _912_ /*1329*/;
  assign r_11[9] = _914_ | _913_ /*1328*/;
  assign _915_ = ~q[1] /*1327*/;
  assign _916_ = sum_11[9] & q[1] /*1326*/;
  assign _917_ = m_11[9] & _915_ /*1325*/;
  assign r_11[10] = _917_ | _916_ /*1324*/;
  assign _918_ = ~q[1] /*1323*/;
  assign _919_ = sum_11[10] & q[1] /*1322*/;
  assign _920_ = m_11[10] & _918_ /*1321*/;
  assign r_11[11] = _920_ | _919_ /*1320*/;
  assign _921_ = ~q[1] /*1319*/;
  assign _922_ = sum_11[11] & q[1] /*1318*/;
  assign _923_ = m_11[11] & _921_ /*1317*/;
  assign r_11[12] = _923_ | _922_ /*1316*/;
assign r_11[0]= r_10[0] /*1315*/;
  assign inv_12[0] = ~div[0] /*1284*/;
  assign inv_12[1] = ~div[1] /*1283*/;
  assign inv_12[2] = ~div[2] /*1282*/;
  assign inv_12[3] = ~div[3] /*1281*/;
  assign inv_12[4] = ~div[4] /*1280*/;
  assign inv_12[5] = ~div[5] /*1279*/;
  assign inv_12[6] = ~div[6] /*1278*/;
  assign inv_12[7] = ~div[7] /*1277*/;
  assign inv_12[8] = ~div[8] /*1276*/;
  assign inv_12[9] = ~div[9] /*1275*/;
  assign inv_12[10] = ~div[10] /*1274*/;
assign inv_12[11] = oneWire /*1273*/;
  assign _924_ = inv_12[0] ^ r_11[0] /*1271*/;
  assign sum_12[0] = _924_ ^ oneWire /*1270*/;
  assign _925_ = _924_ & oneWire /*1269*/;
  assign _926_ = inv_12[0] & r_11[0] /*1268*/;
  assign _927_ = _925_ | _926_ /*1267*/;
  assign _928_ = inv_12[1] ^ r_11[1] /*1266*/;
  assign sum_12[1] = _928_ ^ _927_ /*1265*/;
  assign _929_ = _928_ & _927_ /*1264*/;
  assign _930_ = inv_12[1] & r_11[1] /*1263*/;
  assign _931_ = _929_ | _930_ /*1262*/;
  assign _932_ = inv_12[2] ^ r_11[2] /*1260*/;
  assign sum_12[2] = _932_ ^ _931_ /*1259*/;
  assign _933_ = _932_ & _931_ /*1258*/;
  assign _934_ = inv_12[2] & r_11[2] /*1257*/;
  assign _935_ = _933_ | _934_ /*1256*/;
  assign _936_ = inv_12[3] ^ r_11[3] /*1254*/;
  assign sum_12[3] = _936_ ^ _935_ /*1253*/;
  assign _937_ = _936_ & _935_ /*1252*/;
  assign _938_ = inv_12[3] & r_11[3] /*1251*/;
  assign _939_ = _937_ | _938_ /*1250*/;
  assign _940_ = inv_12[4] ^ r_11[4] /*1248*/;
  assign sum_12[4] = _940_ ^ _939_ /*1247*/;
  assign _941_ = _940_ & _939_ /*1246*/;
  assign _942_ = inv_12[4] & r_11[4] /*1245*/;
  assign _943_ = _941_ | _942_ /*1244*/;
  assign _944_ = inv_12[5] ^ r_11[5] /*1242*/;
  assign sum_12[5] = _944_ ^ _943_ /*1241*/;
  assign _945_ = _944_ & _943_ /*1240*/;
  assign _946_ = inv_12[5] & r_11[5] /*1239*/;
  assign _947_ = _945_ | _946_ /*1238*/;
  assign _948_ = inv_12[6] ^ r_11[6] /*1236*/;
  assign sum_12[6] = _948_ ^ _947_ /*1235*/;
  assign _949_ = _948_ & _947_ /*1234*/;
  assign _950_ = inv_12[6] & r_11[6] /*1233*/;
  assign _951_ = _949_ | _950_ /*1232*/;
  assign _952_ = inv_12[7] ^ r_11[7] /*1230*/;
  assign sum_12[7] = _952_ ^ _951_ /*1229*/;
  assign _953_ = _952_ & _951_ /*1228*/;
  assign _954_ = inv_12[7] & r_11[7] /*1227*/;
  assign _955_ = _953_ | _954_ /*1226*/;
  assign _956_ = inv_12[8] ^ r_11[8] /*1224*/;
  assign sum_12[8] = _956_ ^ _955_ /*1223*/;
  assign _957_ = _956_ & _955_ /*1222*/;
  assign _958_ = inv_12[8] & r_11[8] /*1221*/;
  assign _959_ = _957_ | _958_ /*1220*/;
  assign _960_ = inv_12[9] ^ r_11[9] /*1218*/;
  assign sum_12[9] = _960_ ^ _959_ /*1217*/;
  assign _961_ = _960_ & _959_ /*1216*/;
  assign _962_ = inv_12[9] & r_11[9] /*1215*/;
  assign _963_ = _961_ | _962_ /*1214*/;
  assign _964_ = inv_12[10] ^ r_11[10] /*1212*/;
  assign sum_12[10] = _964_ ^ _963_ /*1211*/;
  assign _965_ = _964_ & _963_ /*1210*/;
  assign _966_ = inv_12[10] & r_11[10] /*1209*/;
  assign _967_ = _965_ | _966_ /*1208*/;
  assign _968_ = inv_12[11] ^ r_11[11] /*1206*/;
  assign sum_12[11] = _968_ ^ _967_ /*1205*/;
  assign _969_ = _968_ & _967_ /*1204*/;
  assign _970_ = inv_12[11] & r_11[11] /*1203*/;
  assign _971_ = _969_ | _970_ /*1202*/;
  assign q[0] = ~sum_12[11] /*1209*/;
  assign m_12[0] = r_11[0] /*1208*/;
  assign m_12[1] = r_11[1] /*1207*/;
  assign m_12[2] = r_11[2] /*1206*/;
  assign m_12[3] = r_11[3] /*1205*/;
  assign m_12[4] = r_11[4] /*1204*/;
  assign m_12[5] = r_11[5] /*1203*/;
  assign m_12[6] = r_11[6] /*1202*/;
  assign m_12[7] = r_11[7] /*1201*/;
  assign m_12[8] = r_11[8] /*1200*/;
  assign m_12[9] = r_11[9] /*1199*/;
  assign m_12[10] = r_11[10] /*1198*/;
  assign m_12[11] = r_11[11] /*1197*/;
  assign _972_ = ~q[0] /*1195*/;
  assign _973_ = sum_12[0] & q[0] /*1194*/;
  assign _974_ = m_12[0] & _972_ /*1193*/;
  assign r_12[0] = _974_ | _973_ /*1192*/;
  assign _975_ = ~q[0] /*1191*/;
  assign _976_ = sum_12[1] & q[0] /*1190*/;
  assign _977_ = m_12[1] & _975_ /*1189*/;
  assign r_12[1] = _977_ | _976_ /*1188*/;
  assign _978_ = ~q[0] /*1187*/;
  assign _979_ = sum_12[2] & q[0] /*1186*/;
  assign _980_ = m_12[2] & _978_ /*1185*/;
  assign r_12[2] = _980_ | _979_ /*1184*/;
  assign _981_ = ~q[0] /*1183*/;
  assign _982_ = sum_12[3] & q[0] /*1182*/;
  assign _983_ = m_12[3] & _981_ /*1181*/;
  assign r_12[3] = _983_ | _982_ /*1180*/;
  assign _984_ = ~q[0] /*1179*/;
  assign _985_ = sum_12[4] & q[0] /*1178*/;
  assign _986_ = m_12[4] & _984_ /*1177*/;
  assign r_12[4] = _986_ | _985_ /*1176*/;
  assign _987_ = ~q[0] /*1175*/;
  assign _988_ = sum_12[5] & q[0] /*1174*/;
  assign _989_ = m_12[5] & _987_ /*1173*/;
  assign r_12[5] = _989_ | _988_ /*1172*/;
  assign _990_ = ~q[0] /*1171*/;
  assign _991_ = sum_12[6] & q[0] /*1170*/;
  assign _992_ = m_12[6] & _990_ /*1169*/;
  assign r_12[6] = _992_ | _991_ /*1168*/;
  assign _993_ = ~q[0] /*1167*/;
  assign _994_ = sum_12[7] & q[0] /*1166*/;
  assign _995_ = m_12[7] & _993_ /*1165*/;
  assign r_12[7] = _995_ | _994_ /*1164*/;
  assign _996_ = ~q[0] /*1163*/;
  assign _997_ = sum_12[8] & q[0] /*1162*/;
  assign _998_ = m_12[8] & _996_ /*1161*/;
  assign r_12[8] = _998_ | _997_ /*1160*/;
  assign _999_ = ~q[0] /*1159*/;
  assign _1000_ = sum_12[9] & q[0] /*1158*/;
  assign _1001_ = m_12[9] & _999_ /*1157*/;
  assign r_12[9] = _1001_ | _1000_ /*1156*/;
  assign _1002_ = ~q[0] /*1155*/;
  assign _1003_ = sum_12[10] & q[0] /*1154*/;
  assign _1004_ = m_12[10] & _1002_ /*1153*/;
  assign r_12[10] = _1004_ | _1003_ /*1152*/;
  assign _1005_ = ~q[0] /*1151*/;
  assign _1006_ = sum_12[11] & q[0] /*1150*/;
  assign _1007_ = m_12[11] & _1005_ /*1149*/;
  assign r_12[11] = _1007_ | _1006_ /*1148*/;
  assign rout[0] = r_12[0] /*0*/;
  assign rout[1] = r_12[1] /*1*/;
  assign rout[2] = r_12[2] /*2*/;
  assign rout[3] = r_12[3] /*3*/;
  assign rout[4] = r_12[4] /*4*/;
  assign rout[5] = r_12[5] /*5*/;
  assign rout[6] = r_12[6] /*6*/;
  assign rout[7] = r_12[7] /*7*/;
  assign rout[8] = r_12[8] /*8*/;
  assign rout[9] = r_12[9] /*9*/;
  assign rout[10] = r_12[10] /*10*/;
  assign rout[11] = r_12[11] /*11*/;
endmodule