module divider(q, rout, rin, div);
  wire _0_;
  wire _1_;
  wire _2_;
  wire _3_;
  wire _4_;
  wire _5_;
  wire _6_;
  wire _7_;
  wire _8_;
  wire _9_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  wire _38_;
  wire _39_;
  wire _40_;
  wire _41_;
  wire _42_;
  wire _43_;
  wire _44_;
  wire _45_;
  wire _46_;
  wire _47_;
  wire _48_;
  wire _49_;
  wire _50_;
  wire _51_;
  wire _52_;
  wire _53_;
  wire _54_;
  wire _55_;
  wire _56_;
  wire _57_;
  wire _58_;
  wire _59_;
  wire _60_;
  wire _61_;
  wire _62_;
  wire _63_;
  wire _64_;
  wire _65_;
  wire _66_;
  wire _67_;
  wire _68_;
  wire _69_;
  wire _70_;
  wire _71_;
  wire _72_;
  wire _73_;
  wire _74_;
  wire _75_;
  wire _76_;
  wire _77_;
  wire _78_;
  wire _79_;
  wire _80_;
  wire _81_;
  wire _82_;
  wire _83_;
  wire _84_;
  wire _85_;
  wire _86_;
  wire _87_;
  wire _88_;
  wire _89_;
  wire _90_;
  wire _91_;
  wire _92_;
  wire _93_;
  wire _94_;
  wire _95_;
  wire _96_;
  wire _97_;
  wire _98_;
  wire _99_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire _304_;
  wire _305_;
  wire _306_;
  wire _307_;
  wire _308_;
  wire _309_;
  wire _310_;
  wire _311_;
  wire _312_;
  wire _313_;
  wire _314_;
  wire _315_;
  wire _316_;
  wire _317_;
  wire _318_;
  wire _319_;
  wire _320_;
  wire _321_;
  wire _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire _326_;
  wire _327_;
  wire _328_;
  wire _329_;
  wire _330_;
  wire _331_;
  wire _332_;
  wire _333_;
  wire _334_;
  wire _335_;
  wire _336_;
  wire _337_;
  wire _338_;
  wire _339_;
  wire _340_;
  wire _341_;
  wire _342_;
  wire _343_;
  wire _344_;
  wire _345_;
  wire _346_;
  wire _347_;
  wire _348_;
  wire _349_;
  wire _350_;
  wire _351_;
  wire _352_;
  wire _353_;
  wire _354_;
  wire _355_;
  wire _356_;
  wire _357_;
  wire _358_;
  wire _359_;
  wire _360_;
  wire _361_;
  wire _362_;
  wire _363_;
  wire _364_;
  wire _365_;
  wire _366_;
  wire _367_;
  wire _368_;
  wire _369_;
  wire _370_;
  wire _371_;
  wire _372_;
  wire _373_;
  wire _374_;
  wire _375_;
  wire _376_;
  wire _377_;
  wire _378_;
  wire _379_;
  wire _380_;
  wire _381_;
  wire _382_;
  wire _383_;
  wire _384_;
  wire _385_;
  wire _386_;
  wire _387_;
  wire _388_;
  wire _389_;
  wire _390_;
  wire _391_;
  wire _392_;
  wire _393_;
  wire _394_;
  wire _395_;
  wire _396_;
  wire _397_;
  wire _398_;
  wire _399_;
  wire _400_;
  wire _401_;
  wire _402_;
  wire _403_;
  wire _404_;
  wire _405_;
  wire _406_;
  wire _407_;
  wire _408_;
  wire _409_;
  wire _410_;
  wire _411_;
  wire _412_;
  wire _413_;
  wire _414_;
  wire _415_;
  wire _416_;
  wire _417_;
  wire _418_;
  wire _419_;
  wire _420_;
  wire _421_;
  wire _422_;
  wire _423_;
  wire _424_;
  wire _425_;
  wire _426_;
  wire _427_;
  wire _428_;
  wire _429_;
  wire _430_;
  wire _431_;
  wire _432_;
  wire _433_;
  wire _434_;
  wire _435_;
  wire _436_;
  wire _437_;
  wire _438_;
  wire _439_;
  wire _440_;
  wire _441_;
  wire _442_;
  wire _443_;
  wire _444_;
  wire _445_;
  wire _446_;
  wire _447_;
  wire _448_;
  wire _449_;
  wire _450_;
  wire _451_;
  wire _452_;
  wire _453_;
  wire _454_;
  wire _455_;
  wire _456_;
  wire _457_;
  wire _458_;
  wire _459_;
  wire _460_;
  wire _461_;
  wire _462_;
  wire _463_;
  wire _464_;
  wire _465_;
  wire _466_;
  wire _467_;
  wire _468_;
  wire _469_;
  wire _470_;
  wire _471_;
  wire _472_;
  wire _473_;
  wire _474_;
  wire _475_;
  wire _476_;
  wire _477_;
  wire _478_;
  wire _479_;
  wire _480_;
  wire _481_;
  wire _482_;
  wire _483_;
  wire _484_;
  wire _485_;
  wire _486_;
  wire _487_;
  wire _488_;
  wire _489_;
  wire _490_;
  wire _491_;
  wire _492_;
  wire _493_;
  wire _494_;
  wire _495_;
  wire _496_;
  wire _497_;
  wire _498_;
  wire _499_;
  wire _500_;
  wire _501_;
  wire _502_;
  wire _503_;
  wire _504_;
  wire _505_;
  wire _506_;
  wire _507_;
  wire _508_;
  wire _509_;
  wire _510_;
  wire _511_;
  wire _512_;
  wire _513_;
  wire _514_;
  wire _515_;
  wire _516_;
  wire _517_;
  wire _518_;
  wire _519_;
  wire _520_;
  wire _521_;
  wire _522_;
  wire _523_;
  wire _524_;
  wire _525_;
  wire _526_;
  wire _527_;
  wire _528_;
  wire _529_;
  wire _530_;
  wire _531_;
  wire _532_;
  wire _533_;
  wire _534_;
  wire _535_;
  wire _536_;
  wire _537_;
  wire _538_;
  wire _539_;
  wire _540_;
  wire _541_;
  wire _542_;
  wire _543_;
  wire _544_;
  wire _545_;
  wire _546_;
  wire _547_;
  wire _548_;
  wire _549_;
  wire _550_;
  wire _551_;
  wire _552_;
  wire _553_;
  wire _554_;
  wire _555_;
  wire _556_;
  wire _557_;
  wire _558_;
  wire _559_;
  wire _560_;
  wire _561_;
  wire _562_;
  wire _563_;
  wire _564_;
  wire _565_;
  wire _566_;
  wire _567_;
  wire _568_;
  wire _569_;
  wire _570_;
  wire _571_;
  wire _572_;
  wire _573_;
  wire _574_;
  wire _575_;
  wire _576_;
  wire _577_;
  wire _578_;
  wire _579_;
  wire _580_;
  wire _581_;
  wire _582_;
  wire _583_;
  wire _584_;
  wire _585_;
  wire _586_;
  wire _587_;
  wire _588_;
  wire _589_;
  wire _590_;
  wire _591_;
  wire _592_;
  wire _593_;
  wire _594_;
  wire _595_;
  wire _596_;
  wire _597_;
  wire _598_;
  wire _599_;
  wire _600_;
  wire _601_;
  wire _602_;
  wire _603_;
  wire _604_;
  wire _605_;
  wire _606_;
  wire _607_;
  wire _608_;
  wire _609_;
  wire _610_;
  wire _611_;
  wire _612_;
  wire _613_;
  wire _614_;
  wire _615_;
  wire _616_;
  wire _617_;
  wire _618_;
  wire _619_;
  wire _620_;
  wire _621_;
  wire _622_;
  wire _623_;
  wire _624_;
  wire _625_;
  wire _626_;
  wire _627_;
  wire _628_;
  wire _629_;
  wire _630_;
  wire _631_;
  wire _632_;
  wire _633_;
  wire _634_;
  wire _635_;
  wire _636_;
  wire _637_;
  wire _638_;
  wire _639_;
  wire _640_;
  wire _641_;
  wire _642_;
  wire _643_;
  wire _644_;
  wire _645_;
  wire _646_;
  wire _647_;
  wire _648_;
  wire _649_;
  wire _650_;
  wire _651_;
  wire _652_;
  wire _653_;
  wire _654_;
  wire _655_;
  wire _656_;
  wire _657_;
  wire _658_;
  wire _659_;
  wire _660_;
  wire _661_;
  wire _662_;
  wire _663_;
  wire _664_;
  wire _665_;
  wire _666_;
  wire _667_;
  wire _668_;
  wire _669_;
  wire _670_;
  wire _671_;
  wire _672_;
  wire _673_;
  wire _674_;
  wire _675_;
  wire _676_;
  wire _677_;
  wire _678_;
  wire _679_;
  wire _680_;
  wire _681_;
  wire _682_;
  wire _683_;
  wire _684_;
  wire _685_;
  wire _686_;
  wire _687_;
  wire _688_;
  wire _689_;
  wire _690_;
  wire _691_;
  wire _692_;
  wire _693_;
  wire _694_;
  wire _695_;
  wire _696_;
  wire _697_;
  wire _698_;
  wire _699_;
  wire _700_;
  wire _701_;
  wire _702_;
  wire _703_;
  wire _704_;
  wire _705_;
  wire _706_;
  wire _707_;
  wire _708_;
  wire _709_;
  wire _710_;
  wire _711_;
  wire _712_;
  wire _713_;
  wire _714_;
  wire _715_;
  wire _716_;
  wire _717_;
  wire _718_;
  wire _719_;
  wire _720_;
  wire _721_;
  wire _722_;
  wire _723_;
  wire _724_;
  wire _725_;
  wire _726_;
  wire _727_;
  wire _728_;
  wire _729_;
  wire _730_;
  wire _731_;
  wire _732_;
  wire _733_;
  wire _734_;
  wire _735_;
  wire _736_;
  wire _737_;
  wire _738_;
  wire _739_;
  wire _740_;
  wire _741_;
  wire _742_;
  wire _743_;
  wire _744_;
  wire _745_;
  wire _746_;
  wire _747_;
  wire _748_;
  wire _749_;
  wire _750_;
  wire _751_;
  wire _752_;
  wire _753_;
  wire _754_;
  wire _755_;
  wire _756_;
  wire _757_;
  wire _758_;
  wire _759_;
  wire _760_;
  wire _761_;
  wire _762_;
  wire _763_;
  wire _764_;
  wire _765_;
  wire _766_;
  wire _767_;
  wire _768_;
  wire _769_;
  wire _770_;
  wire _771_;
  wire _772_;
  wire _773_;
  wire _774_;
  wire _775_;
  wire _776_;
  wire _777_;
  wire _778_;
  wire _779_;
  wire _780_;
  wire _781_;
  wire _782_;
  wire _783_;
  wire _784_;
  wire _785_;
  wire _786_;
  wire _787_;
  wire _788_;
  wire _789_;
  wire _790_;
  wire _791_;
  wire _792_;
  wire _793_;
  wire _794_;
  wire _795_;
  wire _796_;
  wire _797_;
  wire _798_;
  wire _799_;
  wire _800_;
  wire _801_;
  wire _802_;
  wire _803_;
  wire _804_;
  wire _805_;
  wire _806_;
  wire _807_;
  wire _808_;
  wire _809_;
  wire _810_;
  wire _811_;
  wire _812_;
  wire _813_;
  wire _814_;
  wire _815_;
  wire _816_;
  wire _817_;
  wire _818_;
  wire _819_;
  wire _820_;
  wire _821_;
  wire _822_;
  wire _823_;
  wire _824_;
  wire _825_;
  wire _826_;
  wire _827_;
  wire _828_;
  wire _829_;
  wire _830_;
  wire _831_;
  wire _832_;
  wire _833_;
  wire _834_;
  wire _835_;
  wire _836_;
  wire _837_;
  wire _838_;
  wire _839_;
  wire _840_;
  wire _841_;
  wire _842_;
  wire _843_;
  wire _844_;
  wire _845_;
  wire _846_;
  wire _847_;
  wire _848_;
  wire _849_;
  wire _850_;
  wire _851_;
  wire _852_;
  wire _853_;
  wire _854_;
  wire _855_;
  wire _856_;
  wire _857_;
  wire _858_;
  wire _859_;
  wire _860_;
  wire _861_;
  wire _862_;
  wire _863_;
  wire _864_;
  wire _865_;
  wire _866_;
  wire _867_;
  wire _868_;
  wire _869_;
  wire _870_;
  wire _871_;
  wire _872_;
  wire _873_;
  wire _874_;
  wire _875_;
  wire _876_;
  wire _877_;
  wire _878_;
  wire _879_;
  wire _880_;
  wire _881_;
  wire _882_;
  wire _883_;
  wire _884_;
  wire _885_;
  wire _886_;
  wire _887_;
  wire _888_;
  wire _889_;
  wire _890_;
  wire _891_;
  wire _892_;
  wire _893_;
  wire _894_;
  wire _895_;
  wire _896_;
  wire _897_;
  wire _898_;
  wire _899_;
  wire _900_;
  wire _901_;
  wire _902_;
  wire _903_;
  wire _904_;
  wire _905_;
  wire _906_;
  wire _907_;
  wire _908_;
  wire _909_;
  wire _910_;
  wire _911_;
  wire _912_;
  wire _913_;
  wire _914_;
  wire _915_;
  wire _916_;
  wire _917_;
  wire _918_;
  wire _919_;
  wire _920_;
  wire _921_;
  wire _922_;
  wire _923_;
  wire _924_;
  wire _925_;
  wire _926_;
  wire _927_;
  wire _928_;
  wire _929_;
  wire _930_;
  wire _931_;
  wire _932_;
  wire _933_;
  wire _934_;
  wire _935_;
  wire _936_;
  wire _937_;
  wire _938_;
  wire _939_;
  wire _940_;
  wire _941_;
  wire _942_;
  wire _943_;
  wire _944_;
  wire _945_;
  wire _946_;
  wire _947_;
  wire _948_;
  wire _949_;
  wire _950_;
  wire _951_;
  wire _952_;
  wire _953_;
  wire _954_;
  wire _955_;
  wire _956_;
  wire _957_;
  wire _958_;
  wire _959_;
  wire _960_;
  wire _961_;
  wire _962_;
  wire _963_;
  wire _964_;
  wire _965_;
  wire _966_;
  wire _967_;
  wire _968_;
  wire _969_;
  wire _970_;
  wire _971_;
  wire _972_;
  wire _973_;
  wire _974_;
  wire _975_;
  wire _976_;
  wire _977_;
  wire _978_;
  wire _979_;
  wire _980_;
  wire _981_;
  wire _982_;
  wire _983_;
  wire _984_;
  wire _985_;
  wire _986_;
  wire _987_;
  wire _988_;
  wire _989_;
  wire _990_;
  wire _991_;
  wire _992_;
  wire _993_;
  wire _994_;
  wire _995_;
  wire _996_;
  wire _997_;
  wire _998_;
  wire _999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire [14:0] r_0;
  wire [15:0] r_1;
  wire [15:0] m_1;
  wire [15:0] sum_1;
  wire [14:0] inv_1;
  wire [16:0] r_2;
  wire [16:0] m_2;
  wire [16:0] sum_2;
  wire [15:0] inv_2;
  wire [17:0] r_3;
  wire [17:0] m_3;
  wire [17:0] sum_3;
  wire [16:0] inv_3;
  wire [18:0] r_4;
  wire [18:0] m_4;
  wire [18:0] sum_4;
  wire [17:0] inv_4;
  wire [19:0] r_5;
  wire [19:0] m_5;
  wire [19:0] sum_5;
  wire [18:0] inv_5;
  wire [20:0] r_6;
  wire [20:0] m_6;
  wire [20:0] sum_6;
  wire [19:0] inv_6;
  wire [21:0] r_7;
  wire [21:0] m_7;
  wire [21:0] sum_7;
  wire [20:0] inv_7;
  wire [22:0] r_8;
  wire [22:0] m_8;
  wire [22:0] sum_8;
  wire [21:0] inv_8;
  wire zeroWire;
  wire oneWire;
  input [13:0] rin;
  input [6:0] div;
  output [7:0] q;
  output [22:0] rout;
  assign zeroWire = 1'b0 /*0*/;
  assign oneWire = 1'b1 /*0*/;
  assign r_0[0] = rin[0] /*2408*/;
  assign r_0[1] = rin[1] /*2407*/;
  assign r_0[2] = rin[2] /*2406*/;
  assign r_0[3] = rin[3] /*2405*/;
  assign r_0[4] = rin[4] /*2404*/;
  assign r_0[5] = rin[5] /*2403*/;
  assign r_0[6] = rin[6] /*2402*/;
  assign r_0[7] = rin[7] /*2401*/;
  assign r_0[8] = rin[8] /*2400*/;
  assign r_0[9] = rin[9] /*2399*/;
  assign r_0[10] = rin[10] /*2398*/;
  assign r_0[11] = rin[11] /*2397*/;
  assign r_0[12] = rin[12] /*2396*/;
  assign r_0[13] = rin[13] /*2395*/;
  assign r_0[14] = zeroWire /*2394*/;
  assign inv_1[0] = oneWire /*2080*/;
  assign inv_1[1] = oneWire /*2074*/;
  assign inv_1[2] = oneWire /*2068*/;
  assign inv_1[3] = oneWire /*2062*/;
  assign inv_1[4] = oneWire /*2056*/;
  assign inv_1[5] = oneWire /*2050*/;
  assign inv_1[6] = oneWire /*2044*/;
  assign inv_1[7] = ~div[0] /*2038*/;
  assign inv_1[8] = ~div[1] /*2032*/;
  assign inv_1[9] = ~div[2] /*2026*/;
  assign inv_1[10] = ~div[3] /*2020*/;
  assign inv_1[11] = ~div[4] /*2014*/;
  assign inv_1[12] = ~div[5] /*2008*/;
  assign inv_1[13] = ~div[6] /*2002*/;
  assign inv_1[14] = oneWire /*1996*/;
  assign _0_ = inv_1[0] ^ r_0[0] /*2079*/;
  assign sum_1[0] = _0_ ^ oneWire /*2078*/;
  assign _1_ = _0_ & oneWire /*2077*/;
  assign _2_ = inv_1[0] & r_0[0] /*2076*/;
  assign _3_ = _1_ | _2_ /*2075*/;
  assign _4_ = inv_1[1] ^ r_0[1] /*2073*/;
  assign sum_1[1] = _4_ ^ _3_ /*2072*/;
  assign _5_ = _4_ & _3_ /*2071*/;
  assign _6_ = inv_1[1] & r_0[1] /*2070*/;
  assign _7_ = _5_ | _6_ /*2069*/;
  assign _8_ = inv_1[2] ^ r_0[2] /*2067*/;
  assign sum_1[2] = _8_ ^ _7_ /*2066*/;
  assign _9_ = _8_ & _7_ /*2065*/;
  assign _10_ = inv_1[2] & r_0[2] /*2064*/;
  assign _11_ = _9_ | _10_ /*2063*/;
  assign _12_ = inv_1[3] ^ r_0[3] /*2061*/;
  assign sum_1[3] = _12_ ^ _11_ /*2060*/;
  assign _13_ = _12_ & _11_ /*2059*/;
  assign _14_ = inv_1[3] & r_0[3] /*2058*/;
  assign _15_ = _13_ | _14_ /*2057*/;
  assign _16_ = inv_1[4] ^ r_0[4] /*2055*/;
  assign sum_1[4] = _16_ ^ _15_ /*2054*/;
  assign _17_ = _16_ & _15_ /*2053*/;
  assign _18_ = inv_1[4] & r_0[4] /*2052*/;
  assign _19_ = _17_ | _18_ /*2051*/;
  assign _20_ = inv_1[5] ^ r_0[5] /*2049*/;
  assign sum_1[5] = _20_ ^ _19_ /*2048*/;
  assign _21_ = _20_ & _19_ /*2047*/;
  assign _22_ = inv_1[5] & r_0[5] /*2046*/;
  assign _23_ = _21_ | _22_ /*2045*/;
  assign _24_ = inv_1[6] ^ r_0[6] /*2043*/;
  assign sum_1[6] = _24_ ^ _23_ /*2042*/;
  assign _25_ = _24_ & _23_ /*2041*/;
  assign _26_ = inv_1[6] & r_0[6] /*2040*/;
  assign _27_ = _25_ | _26_ /*2039*/;
  assign _28_ = inv_1[7] ^ r_0[7] /*2037*/;
  assign sum_1[7] = _28_ ^ _27_ /*2036*/;
  assign _29_ = _28_ & _27_ /*2035*/;
  assign _30_ = inv_1[7] & r_0[7] /*2034*/;
  assign _31_ = _29_ | _30_ /*2033*/;
  assign _32_ = inv_1[8] ^ r_0[8] /*2031*/;
  assign sum_1[8] = _32_ ^ _31_ /*2030*/;
  assign _33_ = _32_ & _31_ /*2029*/;
  assign _34_ = inv_1[8] & r_0[8] /*2028*/;
  assign _35_ = _33_ | _34_ /*2027*/;
  assign _36_ = inv_1[9] ^ r_0[9] /*2025*/;
  assign sum_1[9] = _36_ ^ _35_ /*2024*/;
  assign _37_ = _36_ & _35_ /*2023*/;
  assign _38_ = inv_1[9] & r_0[9] /*2022*/;
  assign _39_ = _37_ | _38_ /*2021*/;
  assign _40_ = inv_1[10] ^ r_0[10] /*2019*/;
  assign sum_1[10] = _40_ ^ _39_ /*2018*/;
  assign _41_ = _40_ & _39_ /*2017*/;
  assign _42_ = inv_1[10] & r_0[10] /*2016*/;
  assign _43_ = _41_ | _42_ /*2015*/;
  assign _44_ = inv_1[11] ^ r_0[11] /*2013*/;
  assign sum_1[11] = _44_ ^ _43_ /*2012*/;
  assign _45_ = _44_ & _43_ /*2011*/;
  assign _46_ = inv_1[11] & r_0[11] /*2010*/;
  assign _47_ = _45_ | _46_ /*2009*/;
  assign _48_ = inv_1[12] ^ r_0[12] /*2007*/;
  assign sum_1[12] = _48_ ^ _47_ /*2006*/;
  assign _49_ = _48_ & _47_ /*2005*/;
  assign _50_ = inv_1[12] & r_0[12] /*2004*/;
  assign _51_ = _49_ | _50_ /*2003*/;
  assign _52_ = inv_1[13] ^ r_0[13] /*2001*/;
  assign sum_1[13] = _52_ ^ _51_ /*2000*/;
  assign _53_ = _52_ & _51_ /*1999*/;
  assign _54_ = inv_1[13] & r_0[13] /*1998*/;
  assign _55_ = _53_ | _54_ /*1997*/;
  assign _56_ = inv_1[14] ^ r_0[14] /*1995*/;
  assign sum_1[14] = _56_ ^ _55_ /*1994*/;
  assign _57_ = _56_ & _55_ /*1993*/;
  assign _58_ = inv_1[14] & r_0[14] /*1992*/;
  assign _59_ = _57_ | _58_ /*1991*/;
  assign _60_ = _59_ ^ _55_ /*1990*/;
  assign _61_ = ~_60_ /*1989*/;
  assign _62_ = sum_1[14] & _61_ /*1988*/;
  assign _63_ = _60_ & _59_ /*1987*/;
  assign sum_1[15] = _63_ | _62_ /*1986*/;
  assign q[7] = ~sum_1[15] /*1985*/;
  assign m_1[0] = r_0[0] /*1984*/;
  assign m_1[1] = r_0[1] /*1983*/;
  assign m_1[2] = r_0[2] /*1982*/;
  assign m_1[3] = r_0[3] /*1981*/;
  assign m_1[4] = r_0[4] /*1980*/;
  assign m_1[5] = r_0[5] /*1979*/;
  assign m_1[6] = r_0[6] /*1978*/;
  assign m_1[7] = r_0[7] /*1977*/;
  assign m_1[8] = r_0[8] /*1976*/;
  assign m_1[9] = r_0[9] /*1975*/;
  assign m_1[10] = r_0[10] /*1974*/;
  assign m_1[11] = r_0[11] /*1973*/;
  assign m_1[12] = r_0[12] /*1972*/;
  assign m_1[13] = r_0[13] /*1971*/;
  assign m_1[14] = r_0[14] /*1970*/;
  assign m_1[15] = r_0[14] /*1969*/;
  assign _65_ = ~q[7] /*1968*/;
  assign _66_ = sum_1[0] & q[7] /*1967*/;
  assign _67_ = m_1[0] & _65_ /*1966*/;
  assign r_1[0] = _67_ | _66_ /*1965*/;
  assign _68_ = sum_1[1] & q[7] /*1964*/;
  assign _69_ = m_1[1] & _65_ /*1963*/;
  assign r_1[1] = _69_ | _68_ /*1962*/;
  assign _70_ = sum_1[2] & q[7] /*1961*/;
  assign _71_ = m_1[2] & _65_ /*1960*/;
  assign r_1[2] = _71_ | _70_ /*1959*/;
  assign _72_ = sum_1[3] & q[7] /*1958*/;
  assign _73_ = m_1[3] & _65_ /*1957*/;
  assign r_1[3] = _73_ | _72_ /*1956*/;
  assign _74_ = sum_1[4] & q[7] /*1955*/;
  assign _75_ = m_1[4] & _65_ /*1954*/;
  assign r_1[4] = _75_ | _74_ /*1953*/;
  assign _76_ = sum_1[5] & q[7] /*1952*/;
  assign _77_ = m_1[5] & _65_ /*1951*/;
  assign r_1[5] = _77_ | _76_ /*1950*/;
  assign _78_ = sum_1[6] & q[7] /*1949*/;
  assign _79_ = m_1[6] & _65_ /*1948*/;
  assign r_1[6] = _79_ | _78_ /*1947*/;
  assign _80_ = sum_1[7] & q[7] /*1946*/;
  assign _81_ = m_1[7] & _65_ /*1945*/;
  assign r_1[7] = _81_ | _80_ /*1944*/;
  assign _82_ = sum_1[8] & q[7] /*1943*/;
  assign _83_ = m_1[8] & _65_ /*1942*/;
  assign r_1[8] = _83_ | _82_ /*1941*/;
  assign _84_ = sum_1[9] & q[7] /*1940*/;
  assign _85_ = m_1[9] & _65_ /*1939*/;
  assign r_1[9] = _85_ | _84_ /*1938*/;
  assign _86_ = sum_1[10] & q[7] /*1937*/;
  assign _87_ = m_1[10] & _65_ /*1936*/;
  assign r_1[10] = _87_ | _86_ /*1935*/;
  assign _88_ = sum_1[11] & q[7] /*1934*/;
  assign _89_ = m_1[11] & _65_ /*1933*/;
  assign r_1[11] = _89_ | _88_ /*1932*/;
  assign _90_ = sum_1[12] & q[7] /*1931*/;
  assign _91_ = m_1[12] & _65_ /*1930*/;
  assign r_1[12] = _91_ | _90_ /*1929*/;
  assign _92_ = sum_1[13] & q[7] /*1928*/;
  assign _93_ = m_1[13] & _65_ /*1927*/;
  assign r_1[13] = _93_ | _92_ /*1926*/;
  assign _94_ = sum_1[14] & q[7] /*1925*/;
  assign _95_ = m_1[14] & _65_ /*1924*/;
  assign r_1[14] = _95_ | _94_ /*1923*/;
  assign _96_ = sum_1[15] & q[7] /*1922*/;
  assign _97_ = m_1[15] & _65_ /*1921*/;
  assign r_1[15] = _97_ | _96_ /*1920*/;
  assign inv_2[0] = oneWire /*1819*/;
  assign inv_2[1] = oneWire /*1813*/;
  assign inv_2[2] = oneWire /*1807*/;
  assign inv_2[3] = oneWire /*1801*/;
  assign inv_2[4] = oneWire /*1795*/;
  assign inv_2[5] = oneWire /*1789*/;
  assign inv_2[6] = ~div[0] /*1783*/;
  assign inv_2[7] = ~div[1] /*1777*/;
  assign inv_2[8] = ~div[2] /*1771*/;
  assign inv_2[9] = ~div[3] /*1765*/;
  assign inv_2[10] = ~div[4] /*1759*/;
  assign inv_2[11] = ~div[5] /*1753*/;
  assign inv_2[12] = ~div[6] /*1747*/;
  assign inv_2[13] = oneWire /*1741*/;
  assign inv_2[14] = oneWire /*1735*/;
  assign inv_2[15] = oneWire /*1729*/;
  assign _98_ = inv_2[0] ^ r_1[0] /*1818*/;
  assign sum_2[0] = _98_ ^ oneWire /*1817*/;
  assign _99_ = _98_ & oneWire /*1816*/;
  assign _100_ = inv_2[0] & r_1[0] /*1815*/;
  assign _101_ = _99_ | _100_ /*1814*/;
  assign _102_ = inv_2[1] ^ r_1[1] /*1812*/;
  assign sum_2[1] = _102_ ^ _101_ /*1811*/;
  assign _103_ = _102_ & _101_ /*1810*/;
  assign _104_ = inv_2[1] & r_1[1] /*1809*/;
  assign _105_ = _103_ | _104_ /*1808*/;
  assign _106_ = inv_2[2] ^ r_1[2] /*1806*/;
  assign sum_2[2] = _106_ ^ _105_ /*1805*/;
  assign _107_ = _106_ & _105_ /*1804*/;
  assign _108_ = inv_2[2] & r_1[2] /*1803*/;
  assign _109_ = _107_ | _108_ /*1802*/;
  assign _110_ = inv_2[3] ^ r_1[3] /*1800*/;
  assign sum_2[3] = _110_ ^ _109_ /*1799*/;
  assign _111_ = _110_ & _109_ /*1798*/;
  assign _112_ = inv_2[3] & r_1[3] /*1797*/;
  assign _113_ = _111_ | _112_ /*1796*/;
  assign _114_ = inv_2[4] ^ r_1[4] /*1794*/;
  assign sum_2[4] = _114_ ^ _113_ /*1793*/;
  assign _115_ = _114_ & _113_ /*1792*/;
  assign _116_ = inv_2[4] & r_1[4] /*1791*/;
  assign _117_ = _115_ | _116_ /*1790*/;
  assign _118_ = inv_2[5] ^ r_1[5] /*1788*/;
  assign sum_2[5] = _118_ ^ _117_ /*1787*/;
  assign _119_ = _118_ & _117_ /*1786*/;
  assign _120_ = inv_2[5] & r_1[5] /*1785*/;
  assign _121_ = _119_ | _120_ /*1784*/;
  assign _122_ = inv_2[6] ^ r_1[6] /*1782*/;
  assign sum_2[6] = _122_ ^ _121_ /*1781*/;
  assign _123_ = _122_ & _121_ /*1780*/;
  assign _124_ = inv_2[6] & r_1[6] /*1779*/;
  assign _125_ = _123_ | _124_ /*1778*/;
  assign _126_ = inv_2[7] ^ r_1[7] /*1776*/;
  assign sum_2[7] = _126_ ^ _125_ /*1775*/;
  assign _127_ = _126_ & _125_ /*1774*/;
  assign _128_ = inv_2[7] & r_1[7] /*1773*/;
  assign _129_ = _127_ | _128_ /*1772*/;
  assign _130_ = inv_2[8] ^ r_1[8] /*1770*/;
  assign sum_2[8] = _130_ ^ _129_ /*1769*/;
  assign _131_ = _130_ & _129_ /*1768*/;
  assign _132_ = inv_2[8] & r_1[8] /*1767*/;
  assign _133_ = _131_ | _132_ /*1766*/;
  assign _134_ = inv_2[9] ^ r_1[9] /*1764*/;
  assign sum_2[9] = _134_ ^ _133_ /*1763*/;
  assign _135_ = _134_ & _133_ /*1762*/;
  assign _136_ = inv_2[9] & r_1[9] /*1761*/;
  assign _137_ = _135_ | _136_ /*1760*/;
  assign _138_ = inv_2[10] ^ r_1[10] /*1758*/;
  assign sum_2[10] = _138_ ^ _137_ /*1757*/;
  assign _139_ = _138_ & _137_ /*1756*/;
  assign _140_ = inv_2[10] & r_1[10] /*1755*/;
  assign _141_ = _139_ | _140_ /*1754*/;
  assign _142_ = inv_2[11] ^ r_1[11] /*1752*/;
  assign sum_2[11] = _142_ ^ _141_ /*1751*/;
  assign _143_ = _142_ & _141_ /*1750*/;
  assign _144_ = inv_2[11] & r_1[11] /*1749*/;
  assign _145_ = _143_ | _144_ /*1748*/;
  assign _146_ = inv_2[12] ^ r_1[12] /*1746*/;
  assign sum_2[12] = _146_ ^ _145_ /*1745*/;
  assign _147_ = _146_ & _145_ /*1744*/;
  assign _148_ = inv_2[12] & r_1[12] /*1743*/;
  assign _149_ = _147_ | _148_ /*1742*/;
  assign _150_ = inv_2[13] ^ r_1[13] /*1740*/;
  assign sum_2[13] = _150_ ^ _149_ /*1739*/;
  assign _151_ = _150_ & _149_ /*1738*/;
  assign _152_ = inv_2[13] & r_1[13] /*1737*/;
  assign _153_ = _151_ | _152_ /*1736*/;
  assign _154_ = inv_2[14] ^ r_1[14] /*1734*/;
  assign sum_2[14] = _154_ ^ _153_ /*1733*/;
  assign _155_ = _154_ & _153_ /*1732*/;
  assign _156_ = inv_2[14] & r_1[14] /*1731*/;
  assign _157_ = _155_ | _156_ /*1730*/;
  assign _158_ = inv_2[15] ^ r_1[15] /*1728*/;
  assign sum_2[15] = _158_ ^ _157_ /*1727*/;
  assign _159_ = _158_ & _157_ /*1726*/;
  assign _160_ = inv_2[15] & r_1[15] /*1725*/;
  assign _161_ = _159_ | _160_ /*1724*/;
  assign _162_ = _161_ ^ _157_ /*1723*/;
  assign _163_ = ~_162_ /*1722*/;
  assign _164_ = sum_2[15] & _163_ /*1721*/;
  assign _165_ = _162_ & _161_ /*1720*/;
  assign sum_2[16] = _165_ | _164_ /*1719*/;
  assign q[6] = ~sum_2[16] /*1718*/;
  assign m_2[0] = r_1[0] /*1717*/;
  assign m_2[1] = r_1[1] /*1716*/;
  assign m_2[2] = r_1[2] /*1715*/;
  assign m_2[3] = r_1[3] /*1714*/;
  assign m_2[4] = r_1[4] /*1713*/;
  assign m_2[5] = r_1[5] /*1712*/;
  assign m_2[6] = r_1[6] /*1711*/;
  assign m_2[7] = r_1[7] /*1710*/;
  assign m_2[8] = r_1[8] /*1709*/;
  assign m_2[9] = r_1[9] /*1708*/;
  assign m_2[10] = r_1[10] /*1707*/;
  assign m_2[11] = r_1[11] /*1706*/;
  assign m_2[12] = r_1[12] /*1705*/;
  assign m_2[13] = r_1[13] /*1704*/;
  assign m_2[14] = r_1[14] /*1703*/;
  assign m_2[15] = r_1[15] /*1702*/;
  assign m_2[16] = r_1[15] /*1701*/;
  assign _167_ = ~q[6] /*1700*/;
  assign _168_ = sum_2[0] & q[6] /*1699*/;
  assign _169_ = m_2[0] & _167_ /*1698*/;
  assign r_2[0] = _169_ | _168_ /*1697*/;
  assign _170_ = sum_2[1] & q[6] /*1696*/;
  assign _171_ = m_2[1] & _167_ /*1695*/;
  assign r_2[1] = _171_ | _170_ /*1694*/;
  assign _172_ = sum_2[2] & q[6] /*1693*/;
  assign _173_ = m_2[2] & _167_ /*1692*/;
  assign r_2[2] = _173_ | _172_ /*1691*/;
  assign _174_ = sum_2[3] & q[6] /*1690*/;
  assign _175_ = m_2[3] & _167_ /*1689*/;
  assign r_2[3] = _175_ | _174_ /*1688*/;
  assign _176_ = sum_2[4] & q[6] /*1687*/;
  assign _177_ = m_2[4] & _167_ /*1686*/;
  assign r_2[4] = _177_ | _176_ /*1685*/;
  assign _178_ = sum_2[5] & q[6] /*1684*/;
  assign _179_ = m_2[5] & _167_ /*1683*/;
  assign r_2[5] = _179_ | _178_ /*1682*/;
  assign _180_ = sum_2[6] & q[6] /*1681*/;
  assign _181_ = m_2[6] & _167_ /*1680*/;
  assign r_2[6] = _181_ | _180_ /*1679*/;
  assign _182_ = sum_2[7] & q[6] /*1678*/;
  assign _183_ = m_2[7] & _167_ /*1677*/;
  assign r_2[7] = _183_ | _182_ /*1676*/;
  assign _184_ = sum_2[8] & q[6] /*1675*/;
  assign _185_ = m_2[8] & _167_ /*1674*/;
  assign r_2[8] = _185_ | _184_ /*1673*/;
  assign _186_ = sum_2[9] & q[6] /*1672*/;
  assign _187_ = m_2[9] & _167_ /*1671*/;
  assign r_2[9] = _187_ | _186_ /*1670*/;
  assign _188_ = sum_2[10] & q[6] /*1669*/;
  assign _189_ = m_2[10] & _167_ /*1668*/;
  assign r_2[10] = _189_ | _188_ /*1667*/;
  assign _190_ = sum_2[11] & q[6] /*1666*/;
  assign _191_ = m_2[11] & _167_ /*1665*/;
  assign r_2[11] = _191_ | _190_ /*1664*/;
  assign _192_ = sum_2[12] & q[6] /*1663*/;
  assign _193_ = m_2[12] & _167_ /*1662*/;
  assign r_2[12] = _193_ | _192_ /*1661*/;
  assign _194_ = sum_2[13] & q[6] /*1660*/;
  assign _195_ = m_2[13] & _167_ /*1659*/;
  assign r_2[13] = _195_ | _194_ /*1658*/;
  assign _196_ = sum_2[14] & q[6] /*1657*/;
  assign _197_ = m_2[14] & _167_ /*1656*/;
  assign r_2[14] = _197_ | _196_ /*1655*/;
  assign _198_ = sum_2[15] & q[6] /*1654*/;
  assign _199_ = m_2[15] & _167_ /*1653*/;
  assign r_2[15] = _199_ | _198_ /*1652*/;
  assign _200_ = sum_2[16] & q[6] /*1651*/;
  assign _201_ = m_2[16] & _167_ /*1650*/;
  assign r_2[16] = _201_ | _200_ /*1649*/;
  assign inv_3[0] = oneWire /*1558*/;
  assign inv_3[1] = oneWire /*1552*/;
  assign inv_3[2] = oneWire /*1546*/;
  assign inv_3[3] = oneWire /*1540*/;
  assign inv_3[4] = oneWire /*1534*/;
  assign inv_3[5] = ~div[0] /*1528*/;
  assign inv_3[6] = ~div[1] /*1522*/;
  assign inv_3[7] = ~div[2] /*1516*/;
  assign inv_3[8] = ~div[3] /*1510*/;
  assign inv_3[9] = ~div[4] /*1504*/;
  assign inv_3[10] = ~div[5] /*1498*/;
  assign inv_3[11] = ~div[6] /*1492*/;
  assign inv_3[12] = oneWire /*1486*/;
  assign inv_3[13] = oneWire /*1480*/;
  assign inv_3[14] = oneWire /*1474*/;
  assign inv_3[15] = oneWire /*1468*/;
  assign inv_3[16] = oneWire /*1462*/;
  assign _202_ = inv_3[0] ^ r_2[0] /*1557*/;
  assign sum_3[0] = _202_ ^ oneWire /*1556*/;
  assign _203_ = _202_ & oneWire /*1555*/;
  assign _204_ = inv_3[0] & r_2[0] /*1554*/;
  assign _205_ = _203_ | _204_ /*1553*/;
  assign _206_ = inv_3[1] ^ r_2[1] /*1551*/;
  assign sum_3[1] = _206_ ^ _205_ /*1550*/;
  assign _207_ = _206_ & _205_ /*1549*/;
  assign _208_ = inv_3[1] & r_2[1] /*1548*/;
  assign _209_ = _207_ | _208_ /*1547*/;
  assign _210_ = inv_3[2] ^ r_2[2] /*1545*/;
  assign sum_3[2] = _210_ ^ _209_ /*1544*/;
  assign _211_ = _210_ & _209_ /*1543*/;
  assign _212_ = inv_3[2] & r_2[2] /*1542*/;
  assign _213_ = _211_ | _212_ /*1541*/;
  assign _214_ = inv_3[3] ^ r_2[3] /*1539*/;
  assign sum_3[3] = _214_ ^ _213_ /*1538*/;
  assign _215_ = _214_ & _213_ /*1537*/;
  assign _216_ = inv_3[3] & r_2[3] /*1536*/;
  assign _217_ = _215_ | _216_ /*1535*/;
  assign _218_ = inv_3[4] ^ r_2[4] /*1533*/;
  assign sum_3[4] = _218_ ^ _217_ /*1532*/;
  assign _219_ = _218_ & _217_ /*1531*/;
  assign _220_ = inv_3[4] & r_2[4] /*1530*/;
  assign _221_ = _219_ | _220_ /*1529*/;
  assign _222_ = inv_3[5] ^ r_2[5] /*1527*/;
  assign sum_3[5] = _222_ ^ _221_ /*1526*/;
  assign _223_ = _222_ & _221_ /*1525*/;
  assign _224_ = inv_3[5] & r_2[5] /*1524*/;
  assign _225_ = _223_ | _224_ /*1523*/;
  assign _226_ = inv_3[6] ^ r_2[6] /*1521*/;
  assign sum_3[6] = _226_ ^ _225_ /*1520*/;
  assign _227_ = _226_ & _225_ /*1519*/;
  assign _228_ = inv_3[6] & r_2[6] /*1518*/;
  assign _229_ = _227_ | _228_ /*1517*/;
  assign _230_ = inv_3[7] ^ r_2[7] /*1515*/;
  assign sum_3[7] = _230_ ^ _229_ /*1514*/;
  assign _231_ = _230_ & _229_ /*1513*/;
  assign _232_ = inv_3[7] & r_2[7] /*1512*/;
  assign _233_ = _231_ | _232_ /*1511*/;
  assign _234_ = inv_3[8] ^ r_2[8] /*1509*/;
  assign sum_3[8] = _234_ ^ _233_ /*1508*/;
  assign _235_ = _234_ & _233_ /*1507*/;
  assign _236_ = inv_3[8] & r_2[8] /*1506*/;
  assign _237_ = _235_ | _236_ /*1505*/;
  assign _238_ = inv_3[9] ^ r_2[9] /*1503*/;
  assign sum_3[9] = _238_ ^ _237_ /*1502*/;
  assign _239_ = _238_ & _237_ /*1501*/;
  assign _240_ = inv_3[9] & r_2[9] /*1500*/;
  assign _241_ = _239_ | _240_ /*1499*/;
  assign _242_ = inv_3[10] ^ r_2[10] /*1497*/;
  assign sum_3[10] = _242_ ^ _241_ /*1496*/;
  assign _243_ = _242_ & _241_ /*1495*/;
  assign _244_ = inv_3[10] & r_2[10] /*1494*/;
  assign _245_ = _243_ | _244_ /*1493*/;
  assign _246_ = inv_3[11] ^ r_2[11] /*1491*/;
  assign sum_3[11] = _246_ ^ _245_ /*1490*/;
  assign _247_ = _246_ & _245_ /*1489*/;
  assign _248_ = inv_3[11] & r_2[11] /*1488*/;
  assign _249_ = _247_ | _248_ /*1487*/;
  assign _250_ = inv_3[12] ^ r_2[12] /*1485*/;
  assign sum_3[12] = _250_ ^ _249_ /*1484*/;
  assign _251_ = _250_ & _249_ /*1483*/;
  assign _252_ = inv_3[12] & r_2[12] /*1482*/;
  assign _253_ = _251_ | _252_ /*1481*/;
  assign _254_ = inv_3[13] ^ r_2[13] /*1479*/;
  assign sum_3[13] = _254_ ^ _253_ /*1478*/;
  assign _255_ = _254_ & _253_ /*1477*/;
  assign _256_ = inv_3[13] & r_2[13] /*1476*/;
  assign _257_ = _255_ | _256_ /*1475*/;
  assign _258_ = inv_3[14] ^ r_2[14] /*1473*/;
  assign sum_3[14] = _258_ ^ _257_ /*1472*/;
  assign _259_ = _258_ & _257_ /*1471*/;
  assign _260_ = inv_3[14] & r_2[14] /*1470*/;
  assign _261_ = _259_ | _260_ /*1469*/;
  assign _262_ = inv_3[15] ^ r_2[15] /*1467*/;
  assign sum_3[15] = _262_ ^ _261_ /*1466*/;
  assign _263_ = _262_ & _261_ /*1465*/;
  assign _264_ = inv_3[15] & r_2[15] /*1464*/;
  assign _265_ = _263_ | _264_ /*1463*/;
  assign _266_ = inv_3[16] ^ r_2[16] /*1461*/;
  assign sum_3[16] = _266_ ^ _265_ /*1460*/;
  assign _267_ = _266_ & _265_ /*1459*/;
  assign _268_ = inv_3[16] & r_2[16] /*1458*/;
  assign _269_ = _267_ | _268_ /*1457*/;
  assign _270_ = _269_ ^ _265_ /*1456*/;
  assign _271_ = ~_270_ /*1455*/;
  assign _272_ = sum_3[16] & _271_ /*1454*/;
  assign _273_ = _270_ & _269_ /*1453*/;
  assign sum_3[17] = _273_ | _272_ /*1452*/;
  assign q[5] = ~sum_3[17] /*1451*/;
  assign m_3[0] = r_2[0] /*1450*/;
  assign m_3[1] = r_2[1] /*1449*/;
  assign m_3[2] = r_2[2] /*1448*/;
  assign m_3[3] = r_2[3] /*1447*/;
  assign m_3[4] = r_2[4] /*1446*/;
  assign m_3[5] = r_2[5] /*1445*/;
  assign m_3[6] = r_2[6] /*1444*/;
  assign m_3[7] = r_2[7] /*1443*/;
  assign m_3[8] = r_2[8] /*1442*/;
  assign m_3[9] = r_2[9] /*1441*/;
  assign m_3[10] = r_2[10] /*1440*/;
  assign m_3[11] = r_2[11] /*1439*/;
  assign m_3[12] = r_2[12] /*1438*/;
  assign m_3[13] = r_2[13] /*1437*/;
  assign m_3[14] = r_2[14] /*1436*/;
  assign m_3[15] = r_2[15] /*1435*/;
  assign m_3[16] = r_2[16] /*1434*/;
  assign m_3[17] = r_2[16] /*1433*/;
  assign _275_ = ~q[5] /*1432*/;
  assign _276_ = sum_3[0] & q[5] /*1431*/;
  assign _277_ = m_3[0] & _275_ /*1430*/;
  assign r_3[0] = _277_ | _276_ /*1429*/;
  assign _278_ = sum_3[1] & q[5] /*1428*/;
  assign _279_ = m_3[1] & _275_ /*1427*/;
  assign r_3[1] = _279_ | _278_ /*1426*/;
  assign _280_ = sum_3[2] & q[5] /*1425*/;
  assign _281_ = m_3[2] & _275_ /*1424*/;
  assign r_3[2] = _281_ | _280_ /*1423*/;
  assign _282_ = sum_3[3] & q[5] /*1422*/;
  assign _283_ = m_3[3] & _275_ /*1421*/;
  assign r_3[3] = _283_ | _282_ /*1420*/;
  assign _284_ = sum_3[4] & q[5] /*1419*/;
  assign _285_ = m_3[4] & _275_ /*1418*/;
  assign r_3[4] = _285_ | _284_ /*1417*/;
  assign _286_ = sum_3[5] & q[5] /*1416*/;
  assign _287_ = m_3[5] & _275_ /*1415*/;
  assign r_3[5] = _287_ | _286_ /*1414*/;
  assign _288_ = sum_3[6] & q[5] /*1413*/;
  assign _289_ = m_3[6] & _275_ /*1412*/;
  assign r_3[6] = _289_ | _288_ /*1411*/;
  assign _290_ = sum_3[7] & q[5] /*1410*/;
  assign _291_ = m_3[7] & _275_ /*1409*/;
  assign r_3[7] = _291_ | _290_ /*1408*/;
  assign _292_ = sum_3[8] & q[5] /*1407*/;
  assign _293_ = m_3[8] & _275_ /*1406*/;
  assign r_3[8] = _293_ | _292_ /*1405*/;
  assign _294_ = sum_3[9] & q[5] /*1404*/;
  assign _295_ = m_3[9] & _275_ /*1403*/;
  assign r_3[9] = _295_ | _294_ /*1402*/;
  assign _296_ = sum_3[10] & q[5] /*1401*/;
  assign _297_ = m_3[10] & _275_ /*1400*/;
  assign r_3[10] = _297_ | _296_ /*1399*/;
  assign _298_ = sum_3[11] & q[5] /*1398*/;
  assign _299_ = m_3[11] & _275_ /*1397*/;
  assign r_3[11] = _299_ | _298_ /*1396*/;
  assign _300_ = sum_3[12] & q[5] /*1395*/;
  assign _301_ = m_3[12] & _275_ /*1394*/;
  assign r_3[12] = _301_ | _300_ /*1393*/;
  assign _302_ = sum_3[13] & q[5] /*1392*/;
  assign _303_ = m_3[13] & _275_ /*1391*/;
  assign r_3[13] = _303_ | _302_ /*1390*/;
  assign _304_ = sum_3[14] & q[5] /*1389*/;
  assign _305_ = m_3[14] & _275_ /*1388*/;
  assign r_3[14] = _305_ | _304_ /*1387*/;
  assign _306_ = sum_3[15] & q[5] /*1386*/;
  assign _307_ = m_3[15] & _275_ /*1385*/;
  assign r_3[15] = _307_ | _306_ /*1384*/;
  assign _308_ = sum_3[16] & q[5] /*1383*/;
  assign _309_ = m_3[16] & _275_ /*1382*/;
  assign r_3[16] = _309_ | _308_ /*1381*/;
  assign _310_ = sum_3[17] & q[5] /*1380*/;
  assign _311_ = m_3[17] & _275_ /*1379*/;
  assign r_3[17] = _311_ | _310_ /*1378*/;
  assign inv_4[0] = oneWire /*1297*/;
  assign inv_4[1] = oneWire /*1291*/;
  assign inv_4[2] = oneWire /*1285*/;
  assign inv_4[3] = oneWire /*1279*/;
  assign inv_4[4] = ~div[0] /*1273*/;
  assign inv_4[5] = ~div[1] /*1267*/;
  assign inv_4[6] = ~div[2] /*1261*/;
  assign inv_4[7] = ~div[3] /*1255*/;
  assign inv_4[8] = ~div[4] /*1249*/;
  assign inv_4[9] = ~div[5] /*1243*/;
  assign inv_4[10] = ~div[6] /*1237*/;
  assign inv_4[11] = oneWire /*1231*/;
  assign inv_4[12] = oneWire /*1225*/;
  assign inv_4[13] = oneWire /*1219*/;
  assign inv_4[14] = oneWire /*1213*/;
  assign inv_4[15] = oneWire /*1207*/;
  assign inv_4[16] = oneWire /*1201*/;
  assign inv_4[17] = oneWire /*1195*/;
  assign _312_ = inv_4[0] ^ r_3[0] /*1296*/;
  assign sum_4[0] = _312_ ^ oneWire /*1295*/;
  assign _313_ = _312_ & oneWire /*1294*/;
  assign _314_ = inv_4[0] & r_3[0] /*1293*/;
  assign _315_ = _313_ | _314_ /*1292*/;
  assign _316_ = inv_4[1] ^ r_3[1] /*1290*/;
  assign sum_4[1] = _316_ ^ _315_ /*1289*/;
  assign _317_ = _316_ & _315_ /*1288*/;
  assign _318_ = inv_4[1] & r_3[1] /*1287*/;
  assign _319_ = _317_ | _318_ /*1286*/;
  assign _320_ = inv_4[2] ^ r_3[2] /*1284*/;
  assign sum_4[2] = _320_ ^ _319_ /*1283*/;
  assign _321_ = _320_ & _319_ /*1282*/;
  assign _322_ = inv_4[2] & r_3[2] /*1281*/;
  assign _323_ = _321_ | _322_ /*1280*/;
  assign _324_ = inv_4[3] ^ r_3[3] /*1278*/;
  assign sum_4[3] = _324_ ^ _323_ /*1277*/;
  assign _325_ = _324_ & _323_ /*1276*/;
  assign _326_ = inv_4[3] & r_3[3] /*1275*/;
  assign _327_ = _325_ | _326_ /*1274*/;
  assign _328_ = inv_4[4] ^ r_3[4] /*1272*/;
  assign sum_4[4] = _328_ ^ _327_ /*1271*/;
  assign _329_ = _328_ & _327_ /*1270*/;
  assign _330_ = inv_4[4] & r_3[4] /*1269*/;
  assign _331_ = _329_ | _330_ /*1268*/;
  assign _332_ = inv_4[5] ^ r_3[5] /*1266*/;
  assign sum_4[5] = _332_ ^ _331_ /*1265*/;
  assign _333_ = _332_ & _331_ /*1264*/;
  assign _334_ = inv_4[5] & r_3[5] /*1263*/;
  assign _335_ = _333_ | _334_ /*1262*/;
  assign _336_ = inv_4[6] ^ r_3[6] /*1260*/;
  assign sum_4[6] = _336_ ^ _335_ /*1259*/;
  assign _337_ = _336_ & _335_ /*1258*/;
  assign _338_ = inv_4[6] & r_3[6] /*1257*/;
  assign _339_ = _337_ | _338_ /*1256*/;
  assign _340_ = inv_4[7] ^ r_3[7] /*1254*/;
  assign sum_4[7] = _340_ ^ _339_ /*1253*/;
  assign _341_ = _340_ & _339_ /*1252*/;
  assign _342_ = inv_4[7] & r_3[7] /*1251*/;
  assign _343_ = _341_ | _342_ /*1250*/;
  assign _344_ = inv_4[8] ^ r_3[8] /*1248*/;
  assign sum_4[8] = _344_ ^ _343_ /*1247*/;
  assign _345_ = _344_ & _343_ /*1246*/;
  assign _346_ = inv_4[8] & r_3[8] /*1245*/;
  assign _347_ = _345_ | _346_ /*1244*/;
  assign _348_ = inv_4[9] ^ r_3[9] /*1242*/;
  assign sum_4[9] = _348_ ^ _347_ /*1241*/;
  assign _349_ = _348_ & _347_ /*1240*/;
  assign _350_ = inv_4[9] & r_3[9] /*1239*/;
  assign _351_ = _349_ | _350_ /*1238*/;
  assign _352_ = inv_4[10] ^ r_3[10] /*1236*/;
  assign sum_4[10] = _352_ ^ _351_ /*1235*/;
  assign _353_ = _352_ & _351_ /*1234*/;
  assign _354_ = inv_4[10] & r_3[10] /*1233*/;
  assign _355_ = _353_ | _354_ /*1232*/;
  assign _356_ = inv_4[11] ^ r_3[11] /*1230*/;
  assign sum_4[11] = _356_ ^ _355_ /*1229*/;
  assign _357_ = _356_ & _355_ /*1228*/;
  assign _358_ = inv_4[11] & r_3[11] /*1227*/;
  assign _359_ = _357_ | _358_ /*1226*/;
  assign _360_ = inv_4[12] ^ r_3[12] /*1224*/;
  assign sum_4[12] = _360_ ^ _359_ /*1223*/;
  assign _361_ = _360_ & _359_ /*1222*/;
  assign _362_ = inv_4[12] & r_3[12] /*1221*/;
  assign _363_ = _361_ | _362_ /*1220*/;
  assign _364_ = inv_4[13] ^ r_3[13] /*1218*/;
  assign sum_4[13] = _364_ ^ _363_ /*1217*/;
  assign _365_ = _364_ & _363_ /*1216*/;
  assign _366_ = inv_4[13] & r_3[13] /*1215*/;
  assign _367_ = _365_ | _366_ /*1214*/;
  assign _368_ = inv_4[14] ^ r_3[14] /*1212*/;
  assign sum_4[14] = _368_ ^ _367_ /*1211*/;
  assign _369_ = _368_ & _367_ /*1210*/;
  assign _370_ = inv_4[14] & r_3[14] /*1209*/;
  assign _371_ = _369_ | _370_ /*1208*/;
  assign _372_ = inv_4[15] ^ r_3[15] /*1206*/;
  assign sum_4[15] = _372_ ^ _371_ /*1205*/;
  assign _373_ = _372_ & _371_ /*1204*/;
  assign _374_ = inv_4[15] & r_3[15] /*1203*/;
  assign _375_ = _373_ | _374_ /*1202*/;
  assign _376_ = inv_4[16] ^ r_3[16] /*1200*/;
  assign sum_4[16] = _376_ ^ _375_ /*1199*/;
  assign _377_ = _376_ & _375_ /*1198*/;
  assign _378_ = inv_4[16] & r_3[16] /*1197*/;
  assign _379_ = _377_ | _378_ /*1196*/;
  assign _380_ = inv_4[17] ^ r_3[17] /*1194*/;
  assign sum_4[17] = _380_ ^ _379_ /*1193*/;
  assign _381_ = _380_ & _379_ /*1192*/;
  assign _382_ = inv_4[17] & r_3[17] /*1191*/;
  assign _383_ = _381_ | _382_ /*1190*/;
  assign _384_ = _383_ ^ _379_ /*1189*/;
  assign _385_ = ~_384_ /*1188*/;
  assign _386_ = sum_4[17] & _385_ /*1187*/;
  assign _387_ = _384_ & _383_ /*1186*/;
  assign sum_4[18] = _387_ | _386_ /*1185*/;
  assign q[4] = ~sum_4[18] /*1184*/;
  assign m_4[0] = r_3[0] /*1183*/;
  assign m_4[1] = r_3[1] /*1182*/;
  assign m_4[2] = r_3[2] /*1181*/;
  assign m_4[3] = r_3[3] /*1180*/;
  assign m_4[4] = r_3[4] /*1179*/;
  assign m_4[5] = r_3[5] /*1178*/;
  assign m_4[6] = r_3[6] /*1177*/;
  assign m_4[7] = r_3[7] /*1176*/;
  assign m_4[8] = r_3[8] /*1175*/;
  assign m_4[9] = r_3[9] /*1174*/;
  assign m_4[10] = r_3[10] /*1173*/;
  assign m_4[11] = r_3[11] /*1172*/;
  assign m_4[12] = r_3[12] /*1171*/;
  assign m_4[13] = r_3[13] /*1170*/;
  assign m_4[14] = r_3[14] /*1169*/;
  assign m_4[15] = r_3[15] /*1168*/;
  assign m_4[16] = r_3[16] /*1167*/;
  assign m_4[17] = r_3[17] /*1166*/;
  assign m_4[18] = r_3[17] /*1165*/;
  assign _389_ = ~q[4] /*1164*/;
  assign _390_ = sum_4[0] & q[4] /*1163*/;
  assign _391_ = m_4[0] & _389_ /*1162*/;
  assign r_4[0] = _391_ | _390_ /*1161*/;
  assign _392_ = sum_4[1] & q[4] /*1160*/;
  assign _393_ = m_4[1] & _389_ /*1159*/;
  assign r_4[1] = _393_ | _392_ /*1158*/;
  assign _394_ = sum_4[2] & q[4] /*1157*/;
  assign _395_ = m_4[2] & _389_ /*1156*/;
  assign r_4[2] = _395_ | _394_ /*1155*/;
  assign _396_ = sum_4[3] & q[4] /*1154*/;
  assign _397_ = m_4[3] & _389_ /*1153*/;
  assign r_4[3] = _397_ | _396_ /*1152*/;
  assign _398_ = sum_4[4] & q[4] /*1151*/;
  assign _399_ = m_4[4] & _389_ /*1150*/;
  assign r_4[4] = _399_ | _398_ /*1149*/;
  assign _400_ = sum_4[5] & q[4] /*1148*/;
  assign _401_ = m_4[5] & _389_ /*1147*/;
  assign r_4[5] = _401_ | _400_ /*1146*/;
  assign _402_ = sum_4[6] & q[4] /*1145*/;
  assign _403_ = m_4[6] & _389_ /*1144*/;
  assign r_4[6] = _403_ | _402_ /*1143*/;
  assign _404_ = sum_4[7] & q[4] /*1142*/;
  assign _405_ = m_4[7] & _389_ /*1141*/;
  assign r_4[7] = _405_ | _404_ /*1140*/;
  assign _406_ = sum_4[8] & q[4] /*1139*/;
  assign _407_ = m_4[8] & _389_ /*1138*/;
  assign r_4[8] = _407_ | _406_ /*1137*/;
  assign _408_ = sum_4[9] & q[4] /*1136*/;
  assign _409_ = m_4[9] & _389_ /*1135*/;
  assign r_4[9] = _409_ | _408_ /*1134*/;
  assign _410_ = sum_4[10] & q[4] /*1133*/;
  assign _411_ = m_4[10] & _389_ /*1132*/;
  assign r_4[10] = _411_ | _410_ /*1131*/;
  assign _412_ = sum_4[11] & q[4] /*1130*/;
  assign _413_ = m_4[11] & _389_ /*1129*/;
  assign r_4[11] = _413_ | _412_ /*1128*/;
  assign _414_ = sum_4[12] & q[4] /*1127*/;
  assign _415_ = m_4[12] & _389_ /*1126*/;
  assign r_4[12] = _415_ | _414_ /*1125*/;
  assign _416_ = sum_4[13] & q[4] /*1124*/;
  assign _417_ = m_4[13] & _389_ /*1123*/;
  assign r_4[13] = _417_ | _416_ /*1122*/;
  assign _418_ = sum_4[14] & q[4] /*1121*/;
  assign _419_ = m_4[14] & _389_ /*1120*/;
  assign r_4[14] = _419_ | _418_ /*1119*/;
  assign _420_ = sum_4[15] & q[4] /*1118*/;
  assign _421_ = m_4[15] & _389_ /*1117*/;
  assign r_4[15] = _421_ | _420_ /*1116*/;
  assign _422_ = sum_4[16] & q[4] /*1115*/;
  assign _423_ = m_4[16] & _389_ /*1114*/;
  assign r_4[16] = _423_ | _422_ /*1113*/;
  assign _424_ = sum_4[17] & q[4] /*1112*/;
  assign _425_ = m_4[17] & _389_ /*1111*/;
  assign r_4[17] = _425_ | _424_ /*1110*/;
  assign _426_ = sum_4[18] & q[4] /*1109*/;
  assign _427_ = m_4[18] & _389_ /*1108*/;
  assign r_4[18] = _427_ | _426_ /*1107*/;
  assign inv_5[0] = oneWire /*1036*/;
  assign inv_5[1] = oneWire /*1030*/;
  assign inv_5[2] = oneWire /*1024*/;
  assign inv_5[3] = ~div[0] /*1018*/;
  assign inv_5[4] = ~div[1] /*1012*/;
  assign inv_5[5] = ~div[2] /*1006*/;
  assign inv_5[6] = ~div[3] /*1000*/;
  assign inv_5[7] = ~div[4] /*994*/;
  assign inv_5[8] = ~div[5] /*988*/;
  assign inv_5[9] = ~div[6] /*982*/;
  assign inv_5[10] = oneWire /*976*/;
  assign inv_5[11] = oneWire /*970*/;
  assign inv_5[12] = oneWire /*964*/;
  assign inv_5[13] = oneWire /*958*/;
  assign inv_5[14] = oneWire /*952*/;
  assign inv_5[15] = oneWire /*946*/;
  assign inv_5[16] = oneWire /*940*/;
  assign inv_5[17] = oneWire /*934*/;
  assign inv_5[18] = oneWire /*928*/;
  assign _428_ = inv_5[0] ^ r_4[0] /*1035*/;
  assign sum_5[0] = _428_ ^ oneWire /*1034*/;
  assign _429_ = _428_ & oneWire /*1033*/;
  assign _430_ = inv_5[0] & r_4[0] /*1032*/;
  assign _431_ = _429_ | _430_ /*1031*/;
  assign _432_ = inv_5[1] ^ r_4[1] /*1029*/;
  assign sum_5[1] = _432_ ^ _431_ /*1028*/;
  assign _433_ = _432_ & _431_ /*1027*/;
  assign _434_ = inv_5[1] & r_4[1] /*1026*/;
  assign _435_ = _433_ | _434_ /*1025*/;
  assign _436_ = inv_5[2] ^ r_4[2] /*1023*/;
  assign sum_5[2] = _436_ ^ _435_ /*1022*/;
  assign _437_ = _436_ & _435_ /*1021*/;
  assign _438_ = inv_5[2] & r_4[2] /*1020*/;
  assign _439_ = _437_ | _438_ /*1019*/;
  assign _440_ = inv_5[3] ^ r_4[3] /*1017*/;
  assign sum_5[3] = _440_ ^ _439_ /*1016*/;
  assign _441_ = _440_ & _439_ /*1015*/;
  assign _442_ = inv_5[3] & r_4[3] /*1014*/;
  assign _443_ = _441_ | _442_ /*1013*/;
  assign _444_ = inv_5[4] ^ r_4[4] /*1011*/;
  assign sum_5[4] = _444_ ^ _443_ /*1010*/;
  assign _445_ = _444_ & _443_ /*1009*/;
  assign _446_ = inv_5[4] & r_4[4] /*1008*/;
  assign _447_ = _445_ | _446_ /*1007*/;
  assign _448_ = inv_5[5] ^ r_4[5] /*1005*/;
  assign sum_5[5] = _448_ ^ _447_ /*1004*/;
  assign _449_ = _448_ & _447_ /*1003*/;
  assign _450_ = inv_5[5] & r_4[5] /*1002*/;
  assign _451_ = _449_ | _450_ /*1001*/;
  assign _452_ = inv_5[6] ^ r_4[6] /*999*/;
  assign sum_5[6] = _452_ ^ _451_ /*998*/;
  assign _453_ = _452_ & _451_ /*997*/;
  assign _454_ = inv_5[6] & r_4[6] /*996*/;
  assign _455_ = _453_ | _454_ /*995*/;
  assign _456_ = inv_5[7] ^ r_4[7] /*993*/;
  assign sum_5[7] = _456_ ^ _455_ /*992*/;
  assign _457_ = _456_ & _455_ /*991*/;
  assign _458_ = inv_5[7] & r_4[7] /*990*/;
  assign _459_ = _457_ | _458_ /*989*/;
  assign _460_ = inv_5[8] ^ r_4[8] /*987*/;
  assign sum_5[8] = _460_ ^ _459_ /*986*/;
  assign _461_ = _460_ & _459_ /*985*/;
  assign _462_ = inv_5[8] & r_4[8] /*984*/;
  assign _463_ = _461_ | _462_ /*983*/;
  assign _464_ = inv_5[9] ^ r_4[9] /*981*/;
  assign sum_5[9] = _464_ ^ _463_ /*980*/;
  assign _465_ = _464_ & _463_ /*979*/;
  assign _466_ = inv_5[9] & r_4[9] /*978*/;
  assign _467_ = _465_ | _466_ /*977*/;
  assign _468_ = inv_5[10] ^ r_4[10] /*975*/;
  assign sum_5[10] = _468_ ^ _467_ /*974*/;
  assign _469_ = _468_ & _467_ /*973*/;
  assign _470_ = inv_5[10] & r_4[10] /*972*/;
  assign _471_ = _469_ | _470_ /*971*/;
  assign _472_ = inv_5[11] ^ r_4[11] /*969*/;
  assign sum_5[11] = _472_ ^ _471_ /*968*/;
  assign _473_ = _472_ & _471_ /*967*/;
  assign _474_ = inv_5[11] & r_4[11] /*966*/;
  assign _475_ = _473_ | _474_ /*965*/;
  assign _476_ = inv_5[12] ^ r_4[12] /*963*/;
  assign sum_5[12] = _476_ ^ _475_ /*962*/;
  assign _477_ = _476_ & _475_ /*961*/;
  assign _478_ = inv_5[12] & r_4[12] /*960*/;
  assign _479_ = _477_ | _478_ /*959*/;
  assign _480_ = inv_5[13] ^ r_4[13] /*957*/;
  assign sum_5[13] = _480_ ^ _479_ /*956*/;
  assign _481_ = _480_ & _479_ /*955*/;
  assign _482_ = inv_5[13] & r_4[13] /*954*/;
  assign _483_ = _481_ | _482_ /*953*/;
  assign _484_ = inv_5[14] ^ r_4[14] /*951*/;
  assign sum_5[14] = _484_ ^ _483_ /*950*/;
  assign _485_ = _484_ & _483_ /*949*/;
  assign _486_ = inv_5[14] & r_4[14] /*948*/;
  assign _487_ = _485_ | _486_ /*947*/;
  assign _488_ = inv_5[15] ^ r_4[15] /*945*/;
  assign sum_5[15] = _488_ ^ _487_ /*944*/;
  assign _489_ = _488_ & _487_ /*943*/;
  assign _490_ = inv_5[15] & r_4[15] /*942*/;
  assign _491_ = _489_ | _490_ /*941*/;
  assign _492_ = inv_5[16] ^ r_4[16] /*939*/;
  assign sum_5[16] = _492_ ^ _491_ /*938*/;
  assign _493_ = _492_ & _491_ /*937*/;
  assign _494_ = inv_5[16] & r_4[16] /*936*/;
  assign _495_ = _493_ | _494_ /*935*/;
  assign _496_ = inv_5[17] ^ r_4[17] /*933*/;
  assign sum_5[17] = _496_ ^ _495_ /*932*/;
  assign _497_ = _496_ & _495_ /*931*/;
  assign _498_ = inv_5[17] & r_4[17] /*930*/;
  assign _499_ = _497_ | _498_ /*929*/;
  assign _500_ = inv_5[18] ^ r_4[18] /*927*/;
  assign sum_5[18] = _500_ ^ _499_ /*926*/;
  assign _501_ = _500_ & _499_ /*925*/;
  assign _502_ = inv_5[18] & r_4[18] /*924*/;
  assign _503_ = _501_ | _502_ /*923*/;
  assign _504_ = _503_ ^ _499_ /*922*/;
  assign _505_ = ~_504_ /*921*/;
  assign _506_ = sum_5[18] & _505_ /*920*/;
  assign _507_ = _504_ & _503_ /*919*/;
  assign sum_5[19] = _507_ | _506_ /*918*/;
  assign q[3] = ~sum_5[19] /*917*/;
  assign m_5[0] = r_4[0] /*916*/;
  assign m_5[1] = r_4[1] /*915*/;
  assign m_5[2] = r_4[2] /*914*/;
  assign m_5[3] = r_4[3] /*913*/;
  assign m_5[4] = r_4[4] /*912*/;
  assign m_5[5] = r_4[5] /*911*/;
  assign m_5[6] = r_4[6] /*910*/;
  assign m_5[7] = r_4[7] /*909*/;
  assign m_5[8] = r_4[8] /*908*/;
  assign m_5[9] = r_4[9] /*907*/;
  assign m_5[10] = r_4[10] /*906*/;
  assign m_5[11] = r_4[11] /*905*/;
  assign m_5[12] = r_4[12] /*904*/;
  assign m_5[13] = r_4[13] /*903*/;
  assign m_5[14] = r_4[14] /*902*/;
  assign m_5[15] = r_4[15] /*901*/;
  assign m_5[16] = r_4[16] /*900*/;
  assign m_5[17] = r_4[17] /*899*/;
  assign m_5[18] = r_4[18] /*898*/;
  assign m_5[19] = r_4[18] /*897*/;
  assign _509_ = ~q[3] /*896*/;
  assign _510_ = sum_5[0] & q[3] /*895*/;
  assign _511_ = m_5[0] & _509_ /*894*/;
  assign r_5[0] = _511_ | _510_ /*893*/;
  assign _512_ = sum_5[1] & q[3] /*892*/;
  assign _513_ = m_5[1] & _509_ /*891*/;
  assign r_5[1] = _513_ | _512_ /*890*/;
  assign _514_ = sum_5[2] & q[3] /*889*/;
  assign _515_ = m_5[2] & _509_ /*888*/;
  assign r_5[2] = _515_ | _514_ /*887*/;
  assign _516_ = sum_5[3] & q[3] /*886*/;
  assign _517_ = m_5[3] & _509_ /*885*/;
  assign r_5[3] = _517_ | _516_ /*884*/;
  assign _518_ = sum_5[4] & q[3] /*883*/;
  assign _519_ = m_5[4] & _509_ /*882*/;
  assign r_5[4] = _519_ | _518_ /*881*/;
  assign _520_ = sum_5[5] & q[3] /*880*/;
  assign _521_ = m_5[5] & _509_ /*879*/;
  assign r_5[5] = _521_ | _520_ /*878*/;
  assign _522_ = sum_5[6] & q[3] /*877*/;
  assign _523_ = m_5[6] & _509_ /*876*/;
  assign r_5[6] = _523_ | _522_ /*875*/;
  assign _524_ = sum_5[7] & q[3] /*874*/;
  assign _525_ = m_5[7] & _509_ /*873*/;
  assign r_5[7] = _525_ | _524_ /*872*/;
  assign _526_ = sum_5[8] & q[3] /*871*/;
  assign _527_ = m_5[8] & _509_ /*870*/;
  assign r_5[8] = _527_ | _526_ /*869*/;
  assign _528_ = sum_5[9] & q[3] /*868*/;
  assign _529_ = m_5[9] & _509_ /*867*/;
  assign r_5[9] = _529_ | _528_ /*866*/;
  assign _530_ = sum_5[10] & q[3] /*865*/;
  assign _531_ = m_5[10] & _509_ /*864*/;
  assign r_5[10] = _531_ | _530_ /*863*/;
  assign _532_ = sum_5[11] & q[3] /*862*/;
  assign _533_ = m_5[11] & _509_ /*861*/;
  assign r_5[11] = _533_ | _532_ /*860*/;
  assign _534_ = sum_5[12] & q[3] /*859*/;
  assign _535_ = m_5[12] & _509_ /*858*/;
  assign r_5[12] = _535_ | _534_ /*857*/;
  assign _536_ = sum_5[13] & q[3] /*856*/;
  assign _537_ = m_5[13] & _509_ /*855*/;
  assign r_5[13] = _537_ | _536_ /*854*/;
  assign _538_ = sum_5[14] & q[3] /*853*/;
  assign _539_ = m_5[14] & _509_ /*852*/;
  assign r_5[14] = _539_ | _538_ /*851*/;
  assign _540_ = sum_5[15] & q[3] /*850*/;
  assign _541_ = m_5[15] & _509_ /*849*/;
  assign r_5[15] = _541_ | _540_ /*848*/;
  assign _542_ = sum_5[16] & q[3] /*847*/;
  assign _543_ = m_5[16] & _509_ /*846*/;
  assign r_5[16] = _543_ | _542_ /*845*/;
  assign _544_ = sum_5[17] & q[3] /*844*/;
  assign _545_ = m_5[17] & _509_ /*843*/;
  assign r_5[17] = _545_ | _544_ /*842*/;
  assign _546_ = sum_5[18] & q[3] /*841*/;
  assign _547_ = m_5[18] & _509_ /*840*/;
  assign r_5[18] = _547_ | _546_ /*839*/;
  assign _548_ = sum_5[19] & q[3] /*838*/;
  assign _549_ = m_5[19] & _509_ /*837*/;
  assign r_5[19] = _549_ | _548_ /*836*/;
  assign inv_6[0] = oneWire /*775*/;
  assign inv_6[1] = oneWire /*769*/;
  assign inv_6[2] = ~div[0] /*763*/;
  assign inv_6[3] = ~div[1] /*757*/;
  assign inv_6[4] = ~div[2] /*751*/;
  assign inv_6[5] = ~div[3] /*745*/;
  assign inv_6[6] = ~div[4] /*739*/;
  assign inv_6[7] = ~div[5] /*733*/;
  assign inv_6[8] = ~div[6] /*727*/;
  assign inv_6[9] = oneWire /*721*/;
  assign inv_6[10] = oneWire /*715*/;
  assign inv_6[11] = oneWire /*709*/;
  assign inv_6[12] = oneWire /*703*/;
  assign inv_6[13] = oneWire /*697*/;
  assign inv_6[14] = oneWire /*691*/;
  assign inv_6[15] = oneWire /*685*/;
  assign inv_6[16] = oneWire /*679*/;
  assign inv_6[17] = oneWire /*673*/;
  assign inv_6[18] = oneWire /*667*/;
  assign inv_6[19] = oneWire /*661*/;
  assign _550_ = inv_6[0] ^ r_5[0] /*774*/;
  assign sum_6[0] = _550_ ^ oneWire /*773*/;
  assign _551_ = _550_ & oneWire /*772*/;
  assign _552_ = inv_6[0] & r_5[0] /*771*/;
  assign _553_ = _551_ | _552_ /*770*/;
  assign _554_ = inv_6[1] ^ r_5[1] /*768*/;
  assign sum_6[1] = _554_ ^ _553_ /*767*/;
  assign _555_ = _554_ & _553_ /*766*/;
  assign _556_ = inv_6[1] & r_5[1] /*765*/;
  assign _557_ = _555_ | _556_ /*764*/;
  assign _558_ = inv_6[2] ^ r_5[2] /*762*/;
  assign sum_6[2] = _558_ ^ _557_ /*761*/;
  assign _559_ = _558_ & _557_ /*760*/;
  assign _560_ = inv_6[2] & r_5[2] /*759*/;
  assign _561_ = _559_ | _560_ /*758*/;
  assign _562_ = inv_6[3] ^ r_5[3] /*756*/;
  assign sum_6[3] = _562_ ^ _561_ /*755*/;
  assign _563_ = _562_ & _561_ /*754*/;
  assign _564_ = inv_6[3] & r_5[3] /*753*/;
  assign _565_ = _563_ | _564_ /*752*/;
  assign _566_ = inv_6[4] ^ r_5[4] /*750*/;
  assign sum_6[4] = _566_ ^ _565_ /*749*/;
  assign _567_ = _566_ & _565_ /*748*/;
  assign _568_ = inv_6[4] & r_5[4] /*747*/;
  assign _569_ = _567_ | _568_ /*746*/;
  assign _570_ = inv_6[5] ^ r_5[5] /*744*/;
  assign sum_6[5] = _570_ ^ _569_ /*743*/;
  assign _571_ = _570_ & _569_ /*742*/;
  assign _572_ = inv_6[5] & r_5[5] /*741*/;
  assign _573_ = _571_ | _572_ /*740*/;
  assign _574_ = inv_6[6] ^ r_5[6] /*738*/;
  assign sum_6[6] = _574_ ^ _573_ /*737*/;
  assign _575_ = _574_ & _573_ /*736*/;
  assign _576_ = inv_6[6] & r_5[6] /*735*/;
  assign _577_ = _575_ | _576_ /*734*/;
  assign _578_ = inv_6[7] ^ r_5[7] /*732*/;
  assign sum_6[7] = _578_ ^ _577_ /*731*/;
  assign _579_ = _578_ & _577_ /*730*/;
  assign _580_ = inv_6[7] & r_5[7] /*729*/;
  assign _581_ = _579_ | _580_ /*728*/;
  assign _582_ = inv_6[8] ^ r_5[8] /*726*/;
  assign sum_6[8] = _582_ ^ _581_ /*725*/;
  assign _583_ = _582_ & _581_ /*724*/;
  assign _584_ = inv_6[8] & r_5[8] /*723*/;
  assign _585_ = _583_ | _584_ /*722*/;
  assign _586_ = inv_6[9] ^ r_5[9] /*720*/;
  assign sum_6[9] = _586_ ^ _585_ /*719*/;
  assign _587_ = _586_ & _585_ /*718*/;
  assign _588_ = inv_6[9] & r_5[9] /*717*/;
  assign _589_ = _587_ | _588_ /*716*/;
  assign _590_ = inv_6[10] ^ r_5[10] /*714*/;
  assign sum_6[10] = _590_ ^ _589_ /*713*/;
  assign _591_ = _590_ & _589_ /*712*/;
  assign _592_ = inv_6[10] & r_5[10] /*711*/;
  assign _593_ = _591_ | _592_ /*710*/;
  assign _594_ = inv_6[11] ^ r_5[11] /*708*/;
  assign sum_6[11] = _594_ ^ _593_ /*707*/;
  assign _595_ = _594_ & _593_ /*706*/;
  assign _596_ = inv_6[11] & r_5[11] /*705*/;
  assign _597_ = _595_ | _596_ /*704*/;
  assign _598_ = inv_6[12] ^ r_5[12] /*702*/;
  assign sum_6[12] = _598_ ^ _597_ /*701*/;
  assign _599_ = _598_ & _597_ /*700*/;
  assign _600_ = inv_6[12] & r_5[12] /*699*/;
  assign _601_ = _599_ | _600_ /*698*/;
  assign _602_ = inv_6[13] ^ r_5[13] /*696*/;
  assign sum_6[13] = _602_ ^ _601_ /*695*/;
  assign _603_ = _602_ & _601_ /*694*/;
  assign _604_ = inv_6[13] & r_5[13] /*693*/;
  assign _605_ = _603_ | _604_ /*692*/;
  assign _606_ = inv_6[14] ^ r_5[14] /*690*/;
  assign sum_6[14] = _606_ ^ _605_ /*689*/;
  assign _607_ = _606_ & _605_ /*688*/;
  assign _608_ = inv_6[14] & r_5[14] /*687*/;
  assign _609_ = _607_ | _608_ /*686*/;
  assign _610_ = inv_6[15] ^ r_5[15] /*684*/;
  assign sum_6[15] = _610_ ^ _609_ /*683*/;
  assign _611_ = _610_ & _609_ /*682*/;
  assign _612_ = inv_6[15] & r_5[15] /*681*/;
  assign _613_ = _611_ | _612_ /*680*/;
  assign _614_ = inv_6[16] ^ r_5[16] /*678*/;
  assign sum_6[16] = _614_ ^ _613_ /*677*/;
  assign _615_ = _614_ & _613_ /*676*/;
  assign _616_ = inv_6[16] & r_5[16] /*675*/;
  assign _617_ = _615_ | _616_ /*674*/;
  assign _618_ = inv_6[17] ^ r_5[17] /*672*/;
  assign sum_6[17] = _618_ ^ _617_ /*671*/;
  assign _619_ = _618_ & _617_ /*670*/;
  assign _620_ = inv_6[17] & r_5[17] /*669*/;
  assign _621_ = _619_ | _620_ /*668*/;
  assign _622_ = inv_6[18] ^ r_5[18] /*666*/;
  assign sum_6[18] = _622_ ^ _621_ /*665*/;
  assign _623_ = _622_ & _621_ /*664*/;
  assign _624_ = inv_6[18] & r_5[18] /*663*/;
  assign _625_ = _623_ | _624_ /*662*/;
  assign _626_ = inv_6[19] ^ r_5[19] /*660*/;
  assign sum_6[19] = _626_ ^ _625_ /*659*/;
  assign _627_ = _626_ & _625_ /*658*/;
  assign _628_ = inv_6[19] & r_5[19] /*657*/;
  assign _629_ = _627_ | _628_ /*656*/;
  assign _630_ = _629_ ^ _625_ /*655*/;
  assign _631_ = ~_630_ /*654*/;
  assign _632_ = sum_6[19] & _631_ /*653*/;
  assign _633_ = _630_ & _629_ /*652*/;
  assign sum_6[20] = _633_ | _632_ /*651*/;
  assign q[2] = ~sum_6[20] /*650*/;
  assign m_6[0] = r_5[0] /*649*/;
  assign m_6[1] = r_5[1] /*648*/;
  assign m_6[2] = r_5[2] /*647*/;
  assign m_6[3] = r_5[3] /*646*/;
  assign m_6[4] = r_5[4] /*645*/;
  assign m_6[5] = r_5[5] /*644*/;
  assign m_6[6] = r_5[6] /*643*/;
  assign m_6[7] = r_5[7] /*642*/;
  assign m_6[8] = r_5[8] /*641*/;
  assign m_6[9] = r_5[9] /*640*/;
  assign m_6[10] = r_5[10] /*639*/;
  assign m_6[11] = r_5[11] /*638*/;
  assign m_6[12] = r_5[12] /*637*/;
  assign m_6[13] = r_5[13] /*636*/;
  assign m_6[14] = r_5[14] /*635*/;
  assign m_6[15] = r_5[15] /*634*/;
  assign m_6[16] = r_5[16] /*633*/;
  assign m_6[17] = r_5[17] /*632*/;
  assign m_6[18] = r_5[18] /*631*/;
  assign m_6[19] = r_5[19] /*630*/;
  assign m_6[20] = r_5[19] /*629*/;
  assign _635_ = ~q[2] /*628*/;
  assign _636_ = sum_6[0] & q[2] /*627*/;
  assign _637_ = m_6[0] & _635_ /*626*/;
  assign r_6[0] = _637_ | _636_ /*625*/;
  assign _638_ = sum_6[1] & q[2] /*624*/;
  assign _639_ = m_6[1] & _635_ /*623*/;
  assign r_6[1] = _639_ | _638_ /*622*/;
  assign _640_ = sum_6[2] & q[2] /*621*/;
  assign _641_ = m_6[2] & _635_ /*620*/;
  assign r_6[2] = _641_ | _640_ /*619*/;
  assign _642_ = sum_6[3] & q[2] /*618*/;
  assign _643_ = m_6[3] & _635_ /*617*/;
  assign r_6[3] = _643_ | _642_ /*616*/;
  assign _644_ = sum_6[4] & q[2] /*615*/;
  assign _645_ = m_6[4] & _635_ /*614*/;
  assign r_6[4] = _645_ | _644_ /*613*/;
  assign _646_ = sum_6[5] & q[2] /*612*/;
  assign _647_ = m_6[5] & _635_ /*611*/;
  assign r_6[5] = _647_ | _646_ /*610*/;
  assign _648_ = sum_6[6] & q[2] /*609*/;
  assign _649_ = m_6[6] & _635_ /*608*/;
  assign r_6[6] = _649_ | _648_ /*607*/;
  assign _650_ = sum_6[7] & q[2] /*606*/;
  assign _651_ = m_6[7] & _635_ /*605*/;
  assign r_6[7] = _651_ | _650_ /*604*/;
  assign _652_ = sum_6[8] & q[2] /*603*/;
  assign _653_ = m_6[8] & _635_ /*602*/;
  assign r_6[8] = _653_ | _652_ /*601*/;
  assign _654_ = sum_6[9] & q[2] /*600*/;
  assign _655_ = m_6[9] & _635_ /*599*/;
  assign r_6[9] = _655_ | _654_ /*598*/;
  assign _656_ = sum_6[10] & q[2] /*597*/;
  assign _657_ = m_6[10] & _635_ /*596*/;
  assign r_6[10] = _657_ | _656_ /*595*/;
  assign _658_ = sum_6[11] & q[2] /*594*/;
  assign _659_ = m_6[11] & _635_ /*593*/;
  assign r_6[11] = _659_ | _658_ /*592*/;
  assign _660_ = sum_6[12] & q[2] /*591*/;
  assign _661_ = m_6[12] & _635_ /*590*/;
  assign r_6[12] = _661_ | _660_ /*589*/;
  assign _662_ = sum_6[13] & q[2] /*588*/;
  assign _663_ = m_6[13] & _635_ /*587*/;
  assign r_6[13] = _663_ | _662_ /*586*/;
  assign _664_ = sum_6[14] & q[2] /*585*/;
  assign _665_ = m_6[14] & _635_ /*584*/;
  assign r_6[14] = _665_ | _664_ /*583*/;
  assign _666_ = sum_6[15] & q[2] /*582*/;
  assign _667_ = m_6[15] & _635_ /*581*/;
  assign r_6[15] = _667_ | _666_ /*580*/;
  assign _668_ = sum_6[16] & q[2] /*579*/;
  assign _669_ = m_6[16] & _635_ /*578*/;
  assign r_6[16] = _669_ | _668_ /*577*/;
  assign _670_ = sum_6[17] & q[2] /*576*/;
  assign _671_ = m_6[17] & _635_ /*575*/;
  assign r_6[17] = _671_ | _670_ /*574*/;
  assign _672_ = sum_6[18] & q[2] /*573*/;
  assign _673_ = m_6[18] & _635_ /*572*/;
  assign r_6[18] = _673_ | _672_ /*571*/;
  assign _674_ = sum_6[19] & q[2] /*570*/;
  assign _675_ = m_6[19] & _635_ /*569*/;
  assign r_6[19] = _675_ | _674_ /*568*/;
  assign _676_ = sum_6[20] & q[2] /*567*/;
  assign _677_ = m_6[20] & _635_ /*566*/;
  assign r_6[20] = _677_ | _676_ /*565*/;
  assign inv_7[0] = oneWire /*514*/;
  assign inv_7[1] = ~div[0] /*508*/;
  assign inv_7[2] = ~div[1] /*502*/;
  assign inv_7[3] = ~div[2] /*496*/;
  assign inv_7[4] = ~div[3] /*490*/;
  assign inv_7[5] = ~div[4] /*484*/;
  assign inv_7[6] = ~div[5] /*478*/;
  assign inv_7[7] = ~div[6] /*472*/;
  assign inv_7[8] = oneWire /*466*/;
  assign inv_7[9] = oneWire /*460*/;
  assign inv_7[10] = oneWire /*454*/;
  assign inv_7[11] = oneWire /*448*/;
  assign inv_7[12] = oneWire /*442*/;
  assign inv_7[13] = oneWire /*436*/;
  assign inv_7[14] = oneWire /*430*/;
  assign inv_7[15] = oneWire /*424*/;
  assign inv_7[16] = oneWire /*418*/;
  assign inv_7[17] = oneWire /*412*/;
  assign inv_7[18] = oneWire /*406*/;
  assign inv_7[19] = oneWire /*400*/;
  assign inv_7[20] = oneWire /*394*/;
  assign _678_ = inv_7[0] ^ r_6[0] /*513*/;
  assign sum_7[0] = _678_ ^ oneWire /*512*/;
  assign _679_ = _678_ & oneWire /*511*/;
  assign _680_ = inv_7[0] & r_6[0] /*510*/;
  assign _681_ = _679_ | _680_ /*509*/;
  assign _682_ = inv_7[1] ^ r_6[1] /*507*/;
  assign sum_7[1] = _682_ ^ _681_ /*506*/;
  assign _683_ = _682_ & _681_ /*505*/;
  assign _684_ = inv_7[1] & r_6[1] /*504*/;
  assign _685_ = _683_ | _684_ /*503*/;
  assign _686_ = inv_7[2] ^ r_6[2] /*501*/;
  assign sum_7[2] = _686_ ^ _685_ /*500*/;
  assign _687_ = _686_ & _685_ /*499*/;
  assign _688_ = inv_7[2] & r_6[2] /*498*/;
  assign _689_ = _687_ | _688_ /*497*/;
  assign _690_ = inv_7[3] ^ r_6[3] /*495*/;
  assign sum_7[3] = _690_ ^ _689_ /*494*/;
  assign _691_ = _690_ & _689_ /*493*/;
  assign _692_ = inv_7[3] & r_6[3] /*492*/;
  assign _693_ = _691_ | _692_ /*491*/;
  assign _694_ = inv_7[4] ^ r_6[4] /*489*/;
  assign sum_7[4] = _694_ ^ _693_ /*488*/;
  assign _695_ = _694_ & _693_ /*487*/;
  assign _696_ = inv_7[4] & r_6[4] /*486*/;
  assign _697_ = _695_ | _696_ /*485*/;
  assign _698_ = inv_7[5] ^ r_6[5] /*483*/;
  assign sum_7[5] = _698_ ^ _697_ /*482*/;
  assign _699_ = _698_ & _697_ /*481*/;
  assign _700_ = inv_7[5] & r_6[5] /*480*/;
  assign _701_ = _699_ | _700_ /*479*/;
  assign _702_ = inv_7[6] ^ r_6[6] /*477*/;
  assign sum_7[6] = _702_ ^ _701_ /*476*/;
  assign _703_ = _702_ & _701_ /*475*/;
  assign _704_ = inv_7[6] & r_6[6] /*474*/;
  assign _705_ = _703_ | _704_ /*473*/;
  assign _706_ = inv_7[7] ^ r_6[7] /*471*/;
  assign sum_7[7] = _706_ ^ _705_ /*470*/;
  assign _707_ = _706_ & _705_ /*469*/;
  assign _708_ = inv_7[7] & r_6[7] /*468*/;
  assign _709_ = _707_ | _708_ /*467*/;
  assign _710_ = inv_7[8] ^ r_6[8] /*465*/;
  assign sum_7[8] = _710_ ^ _709_ /*464*/;
  assign _711_ = _710_ & _709_ /*463*/;
  assign _712_ = inv_7[8] & r_6[8] /*462*/;
  assign _713_ = _711_ | _712_ /*461*/;
  assign _714_ = inv_7[9] ^ r_6[9] /*459*/;
  assign sum_7[9] = _714_ ^ _713_ /*458*/;
  assign _715_ = _714_ & _713_ /*457*/;
  assign _716_ = inv_7[9] & r_6[9] /*456*/;
  assign _717_ = _715_ | _716_ /*455*/;
  assign _718_ = inv_7[10] ^ r_6[10] /*453*/;
  assign sum_7[10] = _718_ ^ _717_ /*452*/;
  assign _719_ = _718_ & _717_ /*451*/;
  assign _720_ = inv_7[10] & r_6[10] /*450*/;
  assign _721_ = _719_ | _720_ /*449*/;
  assign _722_ = inv_7[11] ^ r_6[11] /*447*/;
  assign sum_7[11] = _722_ ^ _721_ /*446*/;
  assign _723_ = _722_ & _721_ /*445*/;
  assign _724_ = inv_7[11] & r_6[11] /*444*/;
  assign _725_ = _723_ | _724_ /*443*/;
  assign _726_ = inv_7[12] ^ r_6[12] /*441*/;
  assign sum_7[12] = _726_ ^ _725_ /*440*/;
  assign _727_ = _726_ & _725_ /*439*/;
  assign _728_ = inv_7[12] & r_6[12] /*438*/;
  assign _729_ = _727_ | _728_ /*437*/;
  assign _730_ = inv_7[13] ^ r_6[13] /*435*/;
  assign sum_7[13] = _730_ ^ _729_ /*434*/;
  assign _731_ = _730_ & _729_ /*433*/;
  assign _732_ = inv_7[13] & r_6[13] /*432*/;
  assign _733_ = _731_ | _732_ /*431*/;
  assign _734_ = inv_7[14] ^ r_6[14] /*429*/;
  assign sum_7[14] = _734_ ^ _733_ /*428*/;
  assign _735_ = _734_ & _733_ /*427*/;
  assign _736_ = inv_7[14] & r_6[14] /*426*/;
  assign _737_ = _735_ | _736_ /*425*/;
  assign _738_ = inv_7[15] ^ r_6[15] /*423*/;
  assign sum_7[15] = _738_ ^ _737_ /*422*/;
  assign _739_ = _738_ & _737_ /*421*/;
  assign _740_ = inv_7[15] & r_6[15] /*420*/;
  assign _741_ = _739_ | _740_ /*419*/;
  assign _742_ = inv_7[16] ^ r_6[16] /*417*/;
  assign sum_7[16] = _742_ ^ _741_ /*416*/;
  assign _743_ = _742_ & _741_ /*415*/;
  assign _744_ = inv_7[16] & r_6[16] /*414*/;
  assign _745_ = _743_ | _744_ /*413*/;
  assign _746_ = inv_7[17] ^ r_6[17] /*411*/;
  assign sum_7[17] = _746_ ^ _745_ /*410*/;
  assign _747_ = _746_ & _745_ /*409*/;
  assign _748_ = inv_7[17] & r_6[17] /*408*/;
  assign _749_ = _747_ | _748_ /*407*/;
  assign _750_ = inv_7[18] ^ r_6[18] /*405*/;
  assign sum_7[18] = _750_ ^ _749_ /*404*/;
  assign _751_ = _750_ & _749_ /*403*/;
  assign _752_ = inv_7[18] & r_6[18] /*402*/;
  assign _753_ = _751_ | _752_ /*401*/;
  assign _754_ = inv_7[19] ^ r_6[19] /*399*/;
  assign sum_7[19] = _754_ ^ _753_ /*398*/;
  assign _755_ = _754_ & _753_ /*397*/;
  assign _756_ = inv_7[19] & r_6[19] /*396*/;
  assign _757_ = _755_ | _756_ /*395*/;
  assign _758_ = inv_7[20] ^ r_6[20] /*393*/;
  assign sum_7[20] = _758_ ^ _757_ /*392*/;
  assign _759_ = _758_ & _757_ /*391*/;
  assign _760_ = inv_7[20] & r_6[20] /*390*/;
  assign _761_ = _759_ | _760_ /*389*/;
  assign _762_ = _761_ ^ _757_ /*388*/;
  assign _763_ = ~_762_ /*387*/;
  assign _764_ = sum_7[20] & _763_ /*386*/;
  assign _765_ = _762_ & _761_ /*385*/;
  assign sum_7[21] = _765_ | _764_ /*384*/;
  assign q[1] = ~sum_7[21] /*383*/;
  assign m_7[0] = r_6[0] /*382*/;
  assign m_7[1] = r_6[1] /*381*/;
  assign m_7[2] = r_6[2] /*380*/;
  assign m_7[3] = r_6[3] /*379*/;
  assign m_7[4] = r_6[4] /*378*/;
  assign m_7[5] = r_6[5] /*377*/;
  assign m_7[6] = r_6[6] /*376*/;
  assign m_7[7] = r_6[7] /*375*/;
  assign m_7[8] = r_6[8] /*374*/;
  assign m_7[9] = r_6[9] /*373*/;
  assign m_7[10] = r_6[10] /*372*/;
  assign m_7[11] = r_6[11] /*371*/;
  assign m_7[12] = r_6[12] /*370*/;
  assign m_7[13] = r_6[13] /*369*/;
  assign m_7[14] = r_6[14] /*368*/;
  assign m_7[15] = r_6[15] /*367*/;
  assign m_7[16] = r_6[16] /*366*/;
  assign m_7[17] = r_6[17] /*365*/;
  assign m_7[18] = r_6[18] /*364*/;
  assign m_7[19] = r_6[19] /*363*/;
  assign m_7[20] = r_6[20] /*362*/;
  assign m_7[21] = r_6[20] /*361*/;
  assign _767_ = ~q[1] /*360*/;
  assign _768_ = sum_7[0] & q[1] /*359*/;
  assign _769_ = m_7[0] & _767_ /*358*/;
  assign r_7[0] = _769_ | _768_ /*357*/;
  assign _770_ = sum_7[1] & q[1] /*356*/;
  assign _771_ = m_7[1] & _767_ /*355*/;
  assign r_7[1] = _771_ | _770_ /*354*/;
  assign _772_ = sum_7[2] & q[1] /*353*/;
  assign _773_ = m_7[2] & _767_ /*352*/;
  assign r_7[2] = _773_ | _772_ /*351*/;
  assign _774_ = sum_7[3] & q[1] /*350*/;
  assign _775_ = m_7[3] & _767_ /*349*/;
  assign r_7[3] = _775_ | _774_ /*348*/;
  assign _776_ = sum_7[4] & q[1] /*347*/;
  assign _777_ = m_7[4] & _767_ /*346*/;
  assign r_7[4] = _777_ | _776_ /*345*/;
  assign _778_ = sum_7[5] & q[1] /*344*/;
  assign _779_ = m_7[5] & _767_ /*343*/;
  assign r_7[5] = _779_ | _778_ /*342*/;
  assign _780_ = sum_7[6] & q[1] /*341*/;
  assign _781_ = m_7[6] & _767_ /*340*/;
  assign r_7[6] = _781_ | _780_ /*339*/;
  assign _782_ = sum_7[7] & q[1] /*338*/;
  assign _783_ = m_7[7] & _767_ /*337*/;
  assign r_7[7] = _783_ | _782_ /*336*/;
  assign _784_ = sum_7[8] & q[1] /*335*/;
  assign _785_ = m_7[8] & _767_ /*334*/;
  assign r_7[8] = _785_ | _784_ /*333*/;
  assign _786_ = sum_7[9] & q[1] /*332*/;
  assign _787_ = m_7[9] & _767_ /*331*/;
  assign r_7[9] = _787_ | _786_ /*330*/;
  assign _788_ = sum_7[10] & q[1] /*329*/;
  assign _789_ = m_7[10] & _767_ /*328*/;
  assign r_7[10] = _789_ | _788_ /*327*/;
  assign _790_ = sum_7[11] & q[1] /*326*/;
  assign _791_ = m_7[11] & _767_ /*325*/;
  assign r_7[11] = _791_ | _790_ /*324*/;
  assign _792_ = sum_7[12] & q[1] /*323*/;
  assign _793_ = m_7[12] & _767_ /*322*/;
  assign r_7[12] = _793_ | _792_ /*321*/;
  assign _794_ = sum_7[13] & q[1] /*320*/;
  assign _795_ = m_7[13] & _767_ /*319*/;
  assign r_7[13] = _795_ | _794_ /*318*/;
  assign _796_ = sum_7[14] & q[1] /*317*/;
  assign _797_ = m_7[14] & _767_ /*316*/;
  assign r_7[14] = _797_ | _796_ /*315*/;
  assign _798_ = sum_7[15] & q[1] /*314*/;
  assign _799_ = m_7[15] & _767_ /*313*/;
  assign r_7[15] = _799_ | _798_ /*312*/;
  assign _800_ = sum_7[16] & q[1] /*311*/;
  assign _801_ = m_7[16] & _767_ /*310*/;
  assign r_7[16] = _801_ | _800_ /*309*/;
  assign _802_ = sum_7[17] & q[1] /*308*/;
  assign _803_ = m_7[17] & _767_ /*307*/;
  assign r_7[17] = _803_ | _802_ /*306*/;
  assign _804_ = sum_7[18] & q[1] /*305*/;
  assign _805_ = m_7[18] & _767_ /*304*/;
  assign r_7[18] = _805_ | _804_ /*303*/;
  assign _806_ = sum_7[19] & q[1] /*302*/;
  assign _807_ = m_7[19] & _767_ /*301*/;
  assign r_7[19] = _807_ | _806_ /*300*/;
  assign _808_ = sum_7[20] & q[1] /*299*/;
  assign _809_ = m_7[20] & _767_ /*298*/;
  assign r_7[20] = _809_ | _808_ /*297*/;
  assign _810_ = sum_7[21] & q[1] /*296*/;
  assign _811_ = m_7[21] & _767_ /*295*/;
  assign r_7[21] = _811_ | _810_ /*294*/;
  assign inv_8[0] = ~div[0] /*253*/;
  assign inv_8[1] = ~div[1] /*247*/;
  assign inv_8[2] = ~div[2] /*241*/;
  assign inv_8[3] = ~div[3] /*235*/;
  assign inv_8[4] = ~div[4] /*229*/;
  assign inv_8[5] = ~div[5] /*223*/;
  assign inv_8[6] = ~div[6] /*217*/;
  assign inv_8[7] = oneWire /*211*/;
  assign inv_8[8] = oneWire /*205*/;
  assign inv_8[9] = oneWire /*199*/;
  assign inv_8[10] = oneWire /*193*/;
  assign inv_8[11] = oneWire /*187*/;
  assign inv_8[12] = oneWire /*181*/;
  assign inv_8[13] = oneWire /*175*/;
  assign inv_8[14] = oneWire /*169*/;
  assign inv_8[15] = oneWire /*163*/;
  assign inv_8[16] = oneWire /*157*/;
  assign inv_8[17] = oneWire /*151*/;
  assign inv_8[18] = oneWire /*145*/;
  assign inv_8[19] = oneWire /*139*/;
  assign inv_8[20] = oneWire /*133*/;
  assign inv_8[21] = oneWire /*127*/;
  assign _812_ = inv_8[0] ^ r_7[0] /*252*/;
  assign sum_8[0] = _812_ ^ oneWire /*251*/;
  assign _813_ = _812_ & oneWire /*250*/;
  assign _814_ = inv_8[0] & r_7[0] /*249*/;
  assign _815_ = _813_ | _814_ /*248*/;
  assign _816_ = inv_8[1] ^ r_7[1] /*246*/;
  assign sum_8[1] = _816_ ^ _815_ /*245*/;
  assign _817_ = _816_ & _815_ /*244*/;
  assign _818_ = inv_8[1] & r_7[1] /*243*/;
  assign _819_ = _817_ | _818_ /*242*/;
  assign _820_ = inv_8[2] ^ r_7[2] /*240*/;
  assign sum_8[2] = _820_ ^ _819_ /*239*/;
  assign _821_ = _820_ & _819_ /*238*/;
  assign _822_ = inv_8[2] & r_7[2] /*237*/;
  assign _823_ = _821_ | _822_ /*236*/;
  assign _824_ = inv_8[3] ^ r_7[3] /*234*/;
  assign sum_8[3] = _824_ ^ _823_ /*233*/;
  assign _825_ = _824_ & _823_ /*232*/;
  assign _826_ = inv_8[3] & r_7[3] /*231*/;
  assign _827_ = _825_ | _826_ /*230*/;
  assign _828_ = inv_8[4] ^ r_7[4] /*228*/;
  assign sum_8[4] = _828_ ^ _827_ /*227*/;
  assign _829_ = _828_ & _827_ /*226*/;
  assign _830_ = inv_8[4] & r_7[4] /*225*/;
  assign _831_ = _829_ | _830_ /*224*/;
  assign _832_ = inv_8[5] ^ r_7[5] /*222*/;
  assign sum_8[5] = _832_ ^ _831_ /*221*/;
  assign _833_ = _832_ & _831_ /*220*/;
  assign _834_ = inv_8[5] & r_7[5] /*219*/;
  assign _835_ = _833_ | _834_ /*218*/;
  assign _836_ = inv_8[6] ^ r_7[6] /*216*/;
  assign sum_8[6] = _836_ ^ _835_ /*215*/;
  assign _837_ = _836_ & _835_ /*214*/;
  assign _838_ = inv_8[6] & r_7[6] /*213*/;
  assign _839_ = _837_ | _838_ /*212*/;
  assign _840_ = inv_8[7] ^ r_7[7] /*210*/;
  assign sum_8[7] = _840_ ^ _839_ /*209*/;
  assign _841_ = _840_ & _839_ /*208*/;
  assign _842_ = inv_8[7] & r_7[7] /*207*/;
  assign _843_ = _841_ | _842_ /*206*/;
  assign _844_ = inv_8[8] ^ r_7[8] /*204*/;
  assign sum_8[8] = _844_ ^ _843_ /*203*/;
  assign _845_ = _844_ & _843_ /*202*/;
  assign _846_ = inv_8[8] & r_7[8] /*201*/;
  assign _847_ = _845_ | _846_ /*200*/;
  assign _848_ = inv_8[9] ^ r_7[9] /*198*/;
  assign sum_8[9] = _848_ ^ _847_ /*197*/;
  assign _849_ = _848_ & _847_ /*196*/;
  assign _850_ = inv_8[9] & r_7[9] /*195*/;
  assign _851_ = _849_ | _850_ /*194*/;
  assign _852_ = inv_8[10] ^ r_7[10] /*192*/;
  assign sum_8[10] = _852_ ^ _851_ /*191*/;
  assign _853_ = _852_ & _851_ /*190*/;
  assign _854_ = inv_8[10] & r_7[10] /*189*/;
  assign _855_ = _853_ | _854_ /*188*/;
  assign _856_ = inv_8[11] ^ r_7[11] /*186*/;
  assign sum_8[11] = _856_ ^ _855_ /*185*/;
  assign _857_ = _856_ & _855_ /*184*/;
  assign _858_ = inv_8[11] & r_7[11] /*183*/;
  assign _859_ = _857_ | _858_ /*182*/;
  assign _860_ = inv_8[12] ^ r_7[12] /*180*/;
  assign sum_8[12] = _860_ ^ _859_ /*179*/;
  assign _861_ = _860_ & _859_ /*178*/;
  assign _862_ = inv_8[12] & r_7[12] /*177*/;
  assign _863_ = _861_ | _862_ /*176*/;
  assign _864_ = inv_8[13] ^ r_7[13] /*174*/;
  assign sum_8[13] = _864_ ^ _863_ /*173*/;
  assign _865_ = _864_ & _863_ /*172*/;
  assign _866_ = inv_8[13] & r_7[13] /*171*/;
  assign _867_ = _865_ | _866_ /*170*/;
  assign _868_ = inv_8[14] ^ r_7[14] /*168*/;
  assign sum_8[14] = _868_ ^ _867_ /*167*/;
  assign _869_ = _868_ & _867_ /*166*/;
  assign _870_ = inv_8[14] & r_7[14] /*165*/;
  assign _871_ = _869_ | _870_ /*164*/;
  assign _872_ = inv_8[15] ^ r_7[15] /*162*/;
  assign sum_8[15] = _872_ ^ _871_ /*161*/;
  assign _873_ = _872_ & _871_ /*160*/;
  assign _874_ = inv_8[15] & r_7[15] /*159*/;
  assign _875_ = _873_ | _874_ /*158*/;
  assign _876_ = inv_8[16] ^ r_7[16] /*156*/;
  assign sum_8[16] = _876_ ^ _875_ /*155*/;
  assign _877_ = _876_ & _875_ /*154*/;
  assign _878_ = inv_8[16] & r_7[16] /*153*/;
  assign _879_ = _877_ | _878_ /*152*/;
  assign _880_ = inv_8[17] ^ r_7[17] /*150*/;
  assign sum_8[17] = _880_ ^ _879_ /*149*/;
  assign _881_ = _880_ & _879_ /*148*/;
  assign _882_ = inv_8[17] & r_7[17] /*147*/;
  assign _883_ = _881_ | _882_ /*146*/;
  assign _884_ = inv_8[18] ^ r_7[18] /*144*/;
  assign sum_8[18] = _884_ ^ _883_ /*143*/;
  assign _885_ = _884_ & _883_ /*142*/;
  assign _886_ = inv_8[18] & r_7[18] /*141*/;
  assign _887_ = _885_ | _886_ /*140*/;
  assign _888_ = inv_8[19] ^ r_7[19] /*138*/;
  assign sum_8[19] = _888_ ^ _887_ /*137*/;
  assign _889_ = _888_ & _887_ /*136*/;
  assign _890_ = inv_8[19] & r_7[19] /*135*/;
  assign _891_ = _889_ | _890_ /*134*/;
  assign _892_ = inv_8[20] ^ r_7[20] /*132*/;
  assign sum_8[20] = _892_ ^ _891_ /*131*/;
  assign _893_ = _892_ & _891_ /*130*/;
  assign _894_ = inv_8[20] & r_7[20] /*129*/;
  assign _895_ = _893_ | _894_ /*128*/;
  assign _896_ = inv_8[21] ^ r_7[21] /*126*/;
  assign sum_8[21] = _896_ ^ _895_ /*125*/;
  assign _897_ = _896_ & _895_ /*124*/;
  assign _898_ = inv_8[21] & r_7[21] /*123*/;
  assign _899_ = _897_ | _898_ /*122*/;
  assign _900_ = _899_ ^ _895_ /*121*/;
  assign _901_ = ~_900_ /*120*/;
  assign _902_ = sum_8[21] & _901_ /*119*/;
  assign _903_ = _900_ & _899_ /*118*/;
  assign sum_8[22] = _903_ | _902_ /*117*/;
  assign q[0] = ~sum_8[22] /*116*/;
  assign m_8[0] = r_7[0] /*115*/;
  assign m_8[1] = r_7[1] /*114*/;
  assign m_8[2] = r_7[2] /*113*/;
  assign m_8[3] = r_7[3] /*112*/;
  assign m_8[4] = r_7[4] /*111*/;
  assign m_8[5] = r_7[5] /*110*/;
  assign m_8[6] = r_7[6] /*109*/;
  assign m_8[7] = r_7[7] /*108*/;
  assign m_8[8] = r_7[8] /*107*/;
  assign m_8[9] = r_7[9] /*106*/;
  assign m_8[10] = r_7[10] /*105*/;
  assign m_8[11] = r_7[11] /*104*/;
  assign m_8[12] = r_7[12] /*103*/;
  assign m_8[13] = r_7[13] /*102*/;
  assign m_8[14] = r_7[14] /*101*/;
  assign m_8[15] = r_7[15] /*100*/;
  assign m_8[16] = r_7[16] /*99*/;
  assign m_8[17] = r_7[17] /*98*/;
  assign m_8[18] = r_7[18] /*97*/;
  assign m_8[19] = r_7[19] /*96*/;
  assign m_8[20] = r_7[20] /*95*/;
  assign m_8[21] = r_7[21] /*94*/;
  assign m_8[22] = r_7[21] /*93*/;
  assign _905_ = ~q[0] /*92*/;
  assign _906_ = sum_8[0] & q[0] /*91*/;
  assign _907_ = m_8[0] & _905_ /*90*/;
  assign r_8[0] = _907_ | _906_ /*89*/;
  assign _908_ = sum_8[1] & q[0] /*88*/;
  assign _909_ = m_8[1] & _905_ /*87*/;
  assign r_8[1] = _909_ | _908_ /*86*/;
  assign _910_ = sum_8[2] & q[0] /*85*/;
  assign _911_ = m_8[2] & _905_ /*84*/;
  assign r_8[2] = _911_ | _910_ /*83*/;
  assign _912_ = sum_8[3] & q[0] /*82*/;
  assign _913_ = m_8[3] & _905_ /*81*/;
  assign r_8[3] = _913_ | _912_ /*80*/;
  assign _914_ = sum_8[4] & q[0] /*79*/;
  assign _915_ = m_8[4] & _905_ /*78*/;
  assign r_8[4] = _915_ | _914_ /*77*/;
  assign _916_ = sum_8[5] & q[0] /*76*/;
  assign _917_ = m_8[5] & _905_ /*75*/;
  assign r_8[5] = _917_ | _916_ /*74*/;
  assign _918_ = sum_8[6] & q[0] /*73*/;
  assign _919_ = m_8[6] & _905_ /*72*/;
  assign r_8[6] = _919_ | _918_ /*71*/;
  assign _920_ = sum_8[7] & q[0] /*70*/;
  assign _921_ = m_8[7] & _905_ /*69*/;
  assign r_8[7] = _921_ | _920_ /*68*/;
  assign _922_ = sum_8[8] & q[0] /*67*/;
  assign _923_ = m_8[8] & _905_ /*66*/;
  assign r_8[8] = _923_ | _922_ /*65*/;
  assign _924_ = sum_8[9] & q[0] /*64*/;
  assign _925_ = m_8[9] & _905_ /*63*/;
  assign r_8[9] = _925_ | _924_ /*62*/;
  assign _926_ = sum_8[10] & q[0] /*61*/;
  assign _927_ = m_8[10] & _905_ /*60*/;
  assign r_8[10] = _927_ | _926_ /*59*/;
  assign _928_ = sum_8[11] & q[0] /*58*/;
  assign _929_ = m_8[11] & _905_ /*57*/;
  assign r_8[11] = _929_ | _928_ /*56*/;
  assign _930_ = sum_8[12] & q[0] /*55*/;
  assign _931_ = m_8[12] & _905_ /*54*/;
  assign r_8[12] = _931_ | _930_ /*53*/;
  assign _932_ = sum_8[13] & q[0] /*52*/;
  assign _933_ = m_8[13] & _905_ /*51*/;
  assign r_8[13] = _933_ | _932_ /*50*/;
  assign _934_ = sum_8[14] & q[0] /*49*/;
  assign _935_ = m_8[14] & _905_ /*48*/;
  assign r_8[14] = _935_ | _934_ /*47*/;
  assign _936_ = sum_8[15] & q[0] /*46*/;
  assign _937_ = m_8[15] & _905_ /*45*/;
  assign r_8[15] = _937_ | _936_ /*44*/;
  assign _938_ = sum_8[16] & q[0] /*43*/;
  assign _939_ = m_8[16] & _905_ /*42*/;
  assign r_8[16] = _939_ | _938_ /*41*/;
  assign _940_ = sum_8[17] & q[0] /*40*/;
  assign _941_ = m_8[17] & _905_ /*39*/;
  assign r_8[17] = _941_ | _940_ /*38*/;
  assign _942_ = sum_8[18] & q[0] /*37*/;
  assign _943_ = m_8[18] & _905_ /*36*/;
  assign r_8[18] = _943_ | _942_ /*35*/;
  assign _944_ = sum_8[19] & q[0] /*34*/;
  assign _945_ = m_8[19] & _905_ /*33*/;
  assign r_8[19] = _945_ | _944_ /*32*/;
  assign _946_ = sum_8[20] & q[0] /*31*/;
  assign _947_ = m_8[20] & _905_ /*30*/;
  assign r_8[20] = _947_ | _946_ /*29*/;
  assign _948_ = sum_8[21] & q[0] /*28*/;
  assign _949_ = m_8[21] & _905_ /*27*/;
  assign r_8[21] = _949_ | _948_ /*26*/;
  assign _950_ = sum_8[22] & q[0] /*25*/;
  assign _951_ = m_8[22] & _905_ /*24*/;
  assign r_8[22] = _951_ | _950_ /*23*/;
  assign rout[0] = r_8[0] /*0*/;
  assign rout[1] = r_8[1] /*1*/;
  assign rout[2] = r_8[2] /*2*/;
  assign rout[3] = r_8[3] /*3*/;
  assign rout[4] = r_8[4] /*4*/;
  assign rout[5] = r_8[5] /*5*/;
  assign rout[6] = r_8[6] /*6*/;
  assign rout[7] = r_8[7] /*7*/;
  assign rout[8] = r_8[8] /*8*/;
  assign rout[9] = r_8[9] /*9*/;
  assign rout[10] = r_8[10] /*10*/;
  assign rout[11] = r_8[11] /*11*/;
  assign rout[12] = r_8[12] /*12*/;
  assign rout[13] = r_8[13] /*13*/;
  assign rout[14] = r_8[14] /*14*/;
  assign rout[15] = r_8[15] /*15*/;
  assign rout[16] = r_8[16] /*16*/;
  assign rout[17] = r_8[17] /*17*/;
  assign rout[18] = r_8[18] /*18*/;
  assign rout[19] = r_8[19] /*19*/;
  assign rout[20] = r_8[20] /*20*/;
  assign rout[21] = r_8[21] /*21*/;
  assign rout[22] = r_8[22] /*22*/;
endmodule