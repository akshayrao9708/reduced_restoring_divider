module divider(q, rout, rin, div);
  wire _0_;
  wire _1_;
  wire _2_;
  wire _3_;
  wire _4_;
  wire _5_;
  wire _6_;
  wire _7_;
  wire _8_;
  wire _9_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  wire _38_;
  wire _39_;
  wire _40_;
  wire _41_;
  wire _42_;
  wire _43_;
  wire _44_;
  wire _45_;
  wire _46_;
  wire _47_;
  wire _48_;
  wire _49_;
  wire _50_;
  wire _51_;
  wire _52_;
  wire _53_;
  wire _54_;
  wire _55_;
  wire _56_;
  wire _57_;
  wire _58_;
  wire _59_;
  wire _60_;
  wire _61_;
  wire _62_;
  wire _63_;
  wire _64_;
  wire _65_;
  wire _66_;
  wire _67_;
  wire _68_;
  wire _69_;
  wire _70_;
  wire _71_;
  wire _72_;
  wire _73_;
  wire _74_;
  wire _75_;
  wire _76_;
  wire _77_;
  wire _78_;
  wire _79_;
  wire _80_;
  wire _81_;
  wire _82_;
  wire _83_;
  wire _84_;
  wire _85_;
  wire _86_;
  wire _87_;
  wire _88_;
  wire _89_;
  wire _90_;
  wire _91_;
  wire _92_;
  wire _93_;
  wire _94_;
  wire _95_;
  wire _96_;
  wire _97_;
  wire _98_;
  wire _99_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire _304_;
  wire _305_;
  wire _306_;
  wire _307_;
  wire _308_;
  wire _309_;
  wire _310_;
  wire _311_;
  wire _312_;
  wire _313_;
  wire _314_;
  wire _315_;
  wire _316_;
  wire _317_;
  wire _318_;
  wire _319_;
  wire _320_;
  wire _321_;
  wire _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire _326_;
  wire _327_;
  wire _328_;
  wire _329_;
  wire _330_;
  wire _331_;
  wire _332_;
  wire _333_;
  wire _334_;
  wire _335_;
  wire _336_;
  wire _337_;
  wire _338_;
  wire _339_;
  wire _340_;
  wire _341_;
  wire _342_;
  wire _343_;
  wire _344_;
  wire _345_;
  wire _346_;
  wire _347_;
  wire _348_;
  wire _349_;
  wire _350_;
  wire _351_;
  wire _352_;
  wire _353_;
  wire _354_;
  wire _355_;
  wire _356_;
  wire _357_;
  wire _358_;
  wire _359_;
  wire _360_;
  wire _361_;
  wire _362_;
  wire _363_;
  wire _364_;
  wire _365_;
  wire _366_;
  wire _367_;
  wire _368_;
  wire _369_;
  wire _370_;
  wire _371_;
  wire _372_;
  wire _373_;
  wire _374_;
  wire _375_;
  wire _376_;
  wire _377_;
  wire _378_;
  wire _379_;
  wire _380_;
  wire _381_;
  wire _382_;
  wire _383_;
  wire _384_;
  wire _385_;
  wire _386_;
  wire _387_;
  wire _388_;
  wire _389_;
  wire _390_;
  wire _391_;
  wire _392_;
  wire _393_;
  wire _394_;
  wire _395_;
  wire _396_;
  wire _397_;
  wire _398_;
  wire _399_;
  wire _400_;
  wire _401_;
  wire _402_;
  wire _403_;
  wire _404_;
  wire _405_;
  wire _406_;
  wire _407_;
  wire _408_;
  wire _409_;
  wire _410_;
  wire _411_;
  wire _412_;
  wire _413_;
  wire _414_;
  wire _415_;
  wire _416_;
  wire _417_;
  wire _418_;
  wire _419_;
  wire _420_;
  wire _421_;
  wire _422_;
  wire _423_;
  wire _424_;
  wire _425_;
  wire _426_;
  wire _427_;
  wire _428_;
  wire _429_;
  wire _430_;
  wire _431_;
  wire _432_;
  wire _433_;
  wire _434_;
  wire _435_;
  wire _436_;
  wire _437_;
  wire _438_;
  wire _439_;
  wire _440_;
  wire _441_;
  wire _442_;
  wire _443_;
  wire _444_;
  wire _445_;
  wire _446_;
  wire _447_;
  wire _448_;
  wire _449_;
  wire _450_;
  wire _451_;
  wire _452_;
  wire _453_;
  wire _454_;
  wire _455_;
  wire _456_;
  wire _457_;
  wire _458_;
  wire _459_;
  wire _460_;
  wire _461_;
  wire _462_;
  wire _463_;
  wire _464_;
  wire _465_;
  wire _466_;
  wire _467_;
  wire _468_;
  wire _469_;
  wire _470_;
  wire _471_;
  wire _472_;
  wire _473_;
  wire _474_;
  wire _475_;
  wire _476_;
  wire _477_;
  wire _478_;
  wire _479_;
  wire _480_;
  wire _481_;
  wire _482_;
  wire _483_;
  wire _484_;
  wire _485_;
  wire _486_;
  wire _487_;
  wire _488_;
  wire _489_;
  wire _490_;
  wire _491_;
  wire _492_;
  wire _493_;
  wire _494_;
  wire _495_;
  wire _496_;
  wire _497_;
  wire _498_;
  wire _499_;
  wire _500_;
  wire _501_;
  wire _502_;
  wire _503_;
  wire _504_;
  wire _505_;
  wire _506_;
  wire _507_;
  wire _508_;
  wire _509_;
  wire _510_;
  wire _511_;
  wire _512_;
  wire _513_;
  wire _514_;
  wire _515_;
  wire _516_;
  wire _517_;
  wire _518_;
  wire _519_;
  wire _520_;
  wire _521_;
  wire _522_;
  wire _523_;
  wire _524_;
  wire _525_;
  wire _526_;
  wire _527_;
  wire _528_;
  wire _529_;
  wire _530_;
  wire _531_;
  wire _532_;
  wire _533_;
  wire _534_;
  wire _535_;
  wire _536_;
  wire _537_;
  wire _538_;
  wire _539_;
  wire _540_;
  wire _541_;
  wire _542_;
  wire _543_;
  wire _544_;
  wire _545_;
  wire _546_;
  wire _547_;
  wire _548_;
  wire _549_;
  wire _550_;
  wire _551_;
  wire _552_;
  wire _553_;
  wire _554_;
  wire _555_;
  wire _556_;
  wire _557_;
  wire _558_;
  wire _559_;
  wire _560_;
  wire _561_;
  wire _562_;
  wire _563_;
  wire _564_;
  wire _565_;
  wire _566_;
  wire _567_;
  wire _568_;
  wire _569_;
  wire _570_;
  wire _571_;
  wire _572_;
  wire _573_;
  wire _574_;
  wire _575_;
  wire _576_;
  wire _577_;
  wire _578_;
  wire _579_;
  wire _580_;
  wire _581_;
  wire _582_;
  wire _583_;
  wire _584_;
  wire _585_;
  wire _586_;
  wire _587_;
  wire _588_;
  wire _589_;
  wire _590_;
  wire _591_;
  wire _592_;
  wire _593_;
  wire _594_;
  wire _595_;
  wire _596_;
  wire _597_;
  wire _598_;
  wire _599_;
  wire _600_;
  wire _601_;
  wire _602_;
  wire _603_;
  wire _604_;
  wire _605_;
  wire _606_;
  wire _607_;
  wire _608_;
  wire _609_;
  wire _610_;
  wire _611_;
  wire _612_;
  wire _613_;
  wire _614_;
  wire _615_;
  wire _616_;
  wire _617_;
  wire _618_;
  wire _619_;
  wire _620_;
  wire _621_;
  wire _622_;
  wire _623_;
  wire _624_;
  wire _625_;
  wire _626_;
  wire _627_;
  wire _628_;
  wire _629_;
  wire _630_;
  wire _631_;
  wire _632_;
  wire _633_;
  wire _634_;
  wire _635_;
  wire _636_;
  wire _637_;
  wire _638_;
  wire _639_;
  wire _640_;
  wire _641_;
  wire _642_;
  wire _643_;
  wire _644_;
  wire _645_;
  wire _646_;
  wire _647_;
  wire _648_;
  wire _649_;
  wire _650_;
  wire _651_;
  wire _652_;
  wire _653_;
  wire _654_;
  wire _655_;
  wire _656_;
  wire _657_;
  wire _658_;
  wire _659_;
  wire _660_;
  wire _661_;
  wire _662_;
  wire _663_;
  wire _664_;
  wire _665_;
  wire _666_;
  wire _667_;
  wire _668_;
  wire _669_;
  wire _670_;
  wire _671_;
  wire _672_;
  wire _673_;
  wire _674_;
  wire _675_;
  wire _676_;
  wire _677_;
  wire _678_;
  wire _679_;
  wire _680_;
  wire _681_;
  wire _682_;
  wire _683_;
  wire _684_;
  wire _685_;
  wire _686_;
  wire _687_;
  wire _688_;
  wire _689_;
  wire _690_;
  wire _691_;
  wire _692_;
  wire _693_;
  wire _694_;
  wire _695_;
  wire _696_;
  wire _697_;
  wire _698_;
  wire _699_;
  wire _700_;
  wire _701_;
  wire _702_;
  wire _703_;
  wire _704_;
  wire _705_;
  wire _706_;
  wire _707_;
  wire _708_;
  wire _709_;
  wire _710_;
  wire _711_;
  wire _712_;
  wire _713_;
  wire _714_;
  wire _715_;
  wire _716_;
  wire _717_;
  wire _718_;
  wire _719_;
  wire _720_;
  wire _721_;
  wire _722_;
  wire _723_;
  wire _724_;
  wire _725_;
  wire _726_;
  wire _727_;
  wire _728_;
  wire _729_;
  wire _730_;
  wire _731_;
  wire _732_;
  wire _733_;
  wire _734_;
  wire _735_;
  wire _736_;
  wire _737_;
  wire _738_;
  wire _739_;
  wire _740_;
  wire _741_;
  wire _742_;
  wire _743_;
  wire _744_;
  wire _745_;
  wire _746_;
  wire _747_;
  wire _748_;
  wire _749_;
  wire _750_;
  wire _751_;
  wire _752_;
  wire _753_;
  wire _754_;
  wire _755_;
  wire _756_;
  wire _757_;
  wire _758_;
  wire _759_;
  wire _760_;
  wire _761_;
  wire _762_;
  wire _763_;
  wire _764_;
  wire _765_;
  wire _766_;
  wire _767_;
  wire _768_;
  wire _769_;
  wire _770_;
  wire _771_;
  wire _772_;
  wire _773_;
  wire _774_;
  wire _775_;
  wire _776_;
  wire _777_;
  wire _778_;
  wire _779_;
  wire _780_;
  wire _781_;
  wire _782_;
  wire _783_;
  wire _784_;
  wire _785_;
  wire _786_;
  wire _787_;
  wire _788_;
  wire _789_;
  wire _790_;
  wire _791_;
  wire _792_;
  wire _793_;
  wire _794_;
  wire _795_;
  wire _796_;
  wire _797_;
  wire _798_;
  wire _799_;
  wire _800_;
  wire _801_;
  wire _802_;
  wire _803_;
  wire _804_;
  wire _805_;
  wire _806_;
  wire _807_;
  wire _808_;
  wire _809_;
  wire _810_;
  wire _811_;
  wire _812_;
  wire _813_;
  wire _814_;
  wire _815_;
  wire _816_;
  wire _817_;
  wire _818_;
  wire _819_;
  wire _820_;
  wire _821_;
  wire _822_;
  wire _823_;
  wire _824_;
  wire _825_;
  wire _826_;
  wire _827_;
  wire _828_;
  wire _829_;
  wire _830_;
  wire _831_;
  wire _832_;
  wire _833_;
  wire _834_;
  wire _835_;
  wire _836_;
  wire _837_;
  wire _838_;
  wire _839_;
  wire _840_;
  wire _841_;
  wire _842_;
  wire _843_;
  wire _844_;
  wire _845_;
  wire _846_;
  wire _847_;
  wire _848_;
  wire _849_;
  wire _850_;
  wire _851_;
  wire _852_;
  wire _853_;
  wire _854_;
  wire _855_;
  wire _856_;
  wire _857_;
  wire _858_;
  wire _859_;
  wire _860_;
  wire _861_;
  wire _862_;
  wire _863_;
  wire _864_;
  wire _865_;
  wire _866_;
  wire _867_;
  wire _868_;
  wire _869_;
  wire _870_;
  wire _871_;
  wire _872_;
  wire _873_;
  wire _874_;
  wire _875_;
  wire _876_;
  wire _877_;
  wire _878_;
  wire _879_;
  wire _880_;
  wire _881_;
  wire _882_;
  wire _883_;
  wire _884_;
  wire _885_;
  wire _886_;
  wire _887_;
  wire _888_;
  wire _889_;
  wire _890_;
  wire _891_;
  wire _892_;
  wire _893_;
  wire _894_;
  wire _895_;
  wire _896_;
  wire _897_;
  wire _898_;
  wire _899_;
  wire _900_;
  wire _901_;
  wire _902_;
  wire _903_;
  wire _904_;
  wire _905_;
  wire _906_;
  wire _907_;
  wire _908_;
  wire _909_;
  wire _910_;
  wire _911_;
  wire _912_;
  wire _913_;
  wire _914_;
  wire _915_;
  wire _916_;
  wire _917_;
  wire _918_;
  wire _919_;
  wire _920_;
  wire _921_;
  wire _922_;
  wire _923_;
  wire _924_;
  wire _925_;
  wire _926_;
  wire _927_;
  wire _928_;
  wire _929_;
  wire _930_;
  wire _931_;
  wire _932_;
  wire _933_;
  wire _934_;
  wire _935_;
  wire _936_;
  wire _937_;
  wire _938_;
  wire _939_;
  wire _940_;
  wire _941_;
  wire _942_;
  wire _943_;
  wire _944_;
  wire _945_;
  wire _946_;
  wire _947_;
  wire _948_;
  wire _949_;
  wire _950_;
  wire _951_;
  wire _952_;
  wire _953_;
  wire _954_;
  wire _955_;
  wire _956_;
  wire _957_;
  wire _958_;
  wire _959_;
  wire _960_;
  wire _961_;
  wire _962_;
  wire _963_;
  wire _964_;
  wire _965_;
  wire _966_;
  wire _967_;
  wire _968_;
  wire _969_;
  wire _970_;
  wire _971_;
  wire _972_;
  wire _973_;
  wire _974_;
  wire _975_;
  wire _976_;
  wire _977_;
  wire _978_;
  wire _979_;
  wire _980_;
  wire _981_;
  wire _982_;
  wire _983_;
  wire _984_;
  wire _985_;
  wire _986_;
  wire _987_;
  wire _988_;
  wire _989_;
  wire _990_;
  wire _991_;
  wire _992_;
  wire _993_;
  wire _994_;
  wire _995_;
  wire _996_;
  wire _997_;
  wire _998_;
  wire _999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire _1601_;
  wire _1602_;
  wire _1603_;
  wire _1604_;
  wire _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire _1611_;
  wire _1612_;
  wire _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire _1629_;
  wire _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire _1720_;
  wire _1721_;
  wire _1722_;
  wire _1723_;
  wire _1724_;
  wire _1725_;
  wire _1726_;
  wire _1727_;
  wire _1728_;
  wire _1729_;
  wire _1730_;
  wire _1731_;
  wire _1732_;
  wire _1733_;
  wire _1734_;
  wire _1735_;
  wire _1736_;
  wire _1737_;
  wire _1738_;
  wire _1739_;
  wire _1740_;
  wire _1741_;
  wire _1742_;
  wire _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire _1751_;
  wire _1752_;
  wire _1753_;
  wire _1754_;
  wire _1755_;
  wire _1756_;
  wire _1757_;
  wire _1758_;
  wire _1759_;
  wire _1760_;
  wire _1761_;
  wire _1762_;
  wire _1763_;
  wire _1764_;
  wire _1765_;
  wire _1766_;
  wire _1767_;
  wire _1768_;
  wire _1769_;
  wire _1770_;
  wire _1771_;
  wire _1772_;
  wire _1773_;
  wire _1774_;
  wire _1775_;
  wire _1776_;
  wire _1777_;
  wire _1778_;
  wire _1779_;
  wire _1780_;
  wire _1781_;
  wire _1782_;
  wire _1783_;
  wire _1784_;
  wire _1785_;
  wire _1786_;
  wire _1787_;
  wire _1788_;
  wire _1789_;
  wire _1790_;
  wire _1791_;
  wire _1792_;
  wire _1793_;
  wire _1794_;
  wire _1795_;
  wire _1796_;
  wire _1797_;
  wire _1798_;
  wire _1799_;
  wire _1800_;
  wire _1801_;
  wire _1802_;
  wire _1803_;
  wire _1804_;
  wire _1805_;
  wire _1806_;
  wire _1807_;
  wire _1808_;
  wire _1809_;
  wire _1810_;
  wire _1811_;
  wire _1812_;
  wire _1813_;
  wire _1814_;
  wire _1815_;
  wire _1816_;
  wire _1817_;
  wire _1818_;
  wire _1819_;
  wire _1820_;
  wire _1821_;
  wire _1822_;
  wire _1823_;
  wire _1824_;
  wire _1825_;
  wire _1826_;
  wire _1827_;
  wire _1828_;
  wire _1829_;
  wire _1830_;
  wire _1831_;
  wire _1832_;
  wire _1833_;
  wire _1834_;
  wire _1835_;
  wire _1836_;
  wire _1837_;
  wire _1838_;
  wire _1839_;
  wire _1840_;
  wire _1841_;
  wire _1842_;
  wire _1843_;
  wire _1844_;
  wire _1845_;
  wire _1846_;
  wire _1847_;
  wire _1848_;
  wire _1849_;
  wire _1850_;
  wire _1851_;
  wire _1852_;
  wire _1853_;
  wire _1854_;
  wire _1855_;
  wire _1856_;
  wire _1857_;
  wire _1858_;
  wire _1859_;
  wire _1860_;
  wire _1861_;
  wire _1862_;
  wire _1863_;
  wire _1864_;
  wire _1865_;
  wire _1866_;
  wire _1867_;
  wire _1868_;
  wire _1869_;
  wire _1870_;
  wire _1871_;
  wire _1872_;
  wire _1873_;
  wire _1874_;
  wire _1875_;
  wire _1876_;
  wire _1877_;
  wire _1878_;
  wire _1879_;
  wire _1880_;
  wire _1881_;
  wire _1882_;
  wire _1883_;
  wire _1884_;
  wire _1885_;
  wire _1886_;
  wire _1887_;
  wire _1888_;
  wire _1889_;
  wire _1890_;
  wire _1891_;
  wire _1892_;
  wire _1893_;
  wire _1894_;
  wire _1895_;
  wire _1896_;
  wire _1897_;
  wire _1898_;
  wire _1899_;
  wire _1900_;
  wire _1901_;
  wire _1902_;
  wire _1903_;
  wire _1904_;
  wire _1905_;
  wire _1906_;
  wire _1907_;
  wire _1908_;
  wire _1909_;
  wire _1910_;
  wire _1911_;
  wire _1912_;
  wire _1913_;
  wire _1914_;
  wire _1915_;
  wire _1916_;
  wire _1917_;
  wire _1918_;
  wire _1919_;
  wire _1920_;
  wire _1921_;
  wire _1922_;
  wire _1923_;
  wire _1924_;
  wire _1925_;
  wire _1926_;
  wire _1927_;
  wire _1928_;
  wire _1929_;
  wire _1930_;
  wire _1931_;
  wire _1932_;
  wire _1933_;
  wire _1934_;
  wire _1935_;
  wire _1936_;
  wire _1937_;
  wire _1938_;
  wire _1939_;
  wire _1940_;
  wire _1941_;
  wire _1942_;
  wire _1943_;
  wire _1944_;
  wire _1945_;
  wire _1946_;
  wire _1947_;
  wire _1948_;
  wire _1949_;
  wire _1950_;
  wire _1951_;
  wire _1952_;
  wire _1953_;
  wire _1954_;
  wire _1955_;
  wire _1956_;
  wire _1957_;
  wire _1958_;
  wire _1959_;
  wire _1960_;
  wire _1961_;
  wire _1962_;
  wire _1963_;
  wire _1964_;
  wire _1965_;
  wire _1966_;
  wire _1967_;
  wire _1968_;
  wire _1969_;
  wire _1970_;
  wire _1971_;
  wire _1972_;
  wire _1973_;
  wire _1974_;
  wire _1975_;
  wire _1976_;
  wire _1977_;
  wire _1978_;
  wire _1979_;
  wire _1980_;
  wire _1981_;
  wire _1982_;
  wire _1983_;
  wire _1984_;
  wire _1985_;
  wire _1986_;
  wire _1987_;
  wire _1988_;
  wire _1989_;
  wire _1990_;
  wire _1991_;
  wire _1992_;
  wire _1993_;
  wire _1994_;
  wire _1995_;
  wire _1996_;
  wire _1997_;
  wire _1998_;
  wire _1999_;
  wire _2000_;
  wire _2001_;
  wire _2002_;
  wire _2003_;
  wire _2004_;
  wire _2005_;
  wire _2006_;
  wire _2007_;
  wire _2008_;
  wire _2009_;
  wire _2010_;
  wire _2011_;
  wire _2012_;
  wire _2013_;
  wire _2014_;
  wire _2015_;
  wire _2016_;
  wire _2017_;
  wire _2018_;
  wire _2019_;
  wire _2020_;
  wire _2021_;
  wire _2022_;
  wire _2023_;
  wire _2024_;
  wire _2025_;
  wire _2026_;
  wire _2027_;
  wire _2028_;
  wire _2029_;
  wire _2030_;
  wire _2031_;
  wire _2032_;
  wire _2033_;
  wire _2034_;
  wire _2035_;
  wire _2036_;
  wire _2037_;
  wire _2038_;
  wire _2039_;
  wire _2040_;
  wire _2041_;
  wire _2042_;
  wire _2043_;
  wire _2044_;
  wire _2045_;
  wire _2046_;
  wire _2047_;
  wire _2048_;
  wire _2049_;
  wire _2050_;
  wire _2051_;
  wire _2052_;
  wire _2053_;
  wire _2054_;
  wire _2055_;
  wire _2056_;
  wire _2057_;
  wire _2058_;
  wire _2059_;
  wire _2060_;
  wire _2061_;
  wire _2062_;
  wire _2063_;
  wire _2064_;
  wire _2065_;
  wire _2066_;
  wire _2067_;
  wire _2068_;
  wire _2069_;
  wire _2070_;
  wire _2071_;
  wire _2072_;
  wire _2073_;
  wire _2074_;
  wire _2075_;
  wire _2076_;
  wire _2077_;
  wire _2078_;
  wire _2079_;
  wire _2080_;
  wire _2081_;
  wire _2082_;
  wire _2083_;
  wire _2084_;
  wire _2085_;
  wire _2086_;
  wire _2087_;
  wire _2088_;
  wire _2089_;
  wire _2090_;
  wire _2091_;
  wire _2092_;
  wire _2093_;
  wire _2094_;
  wire _2095_;
  wire _2096_;
  wire _2097_;
  wire _2098_;
  wire _2099_;
  wire _2100_;
  wire _2101_;
  wire _2102_;
  wire _2103_;
  wire _2104_;
  wire _2105_;
  wire _2106_;
  wire _2107_;
  wire _2108_;
  wire _2109_;
  wire _2110_;
  wire _2111_;
  wire _2112_;
  wire _2113_;
  wire _2114_;
  wire _2115_;
  wire _2116_;
  wire _2117_;
  wire _2118_;
  wire _2119_;
  wire _2120_;
  wire _2121_;
  wire _2122_;
  wire _2123_;
  wire _2124_;
  wire _2125_;
  wire _2126_;
  wire _2127_;
  wire _2128_;
  wire _2129_;
  wire _2130_;
  wire _2131_;
  wire _2132_;
  wire _2133_;
  wire _2134_;
  wire _2135_;
  wire _2136_;
  wire _2137_;
  wire _2138_;
  wire _2139_;
  wire _2140_;
  wire _2141_;
  wire _2142_;
  wire _2143_;
  wire _2144_;
  wire _2145_;
  wire _2146_;
  wire _2147_;
  wire _2148_;
  wire _2149_;
  wire _2150_;
  wire _2151_;
  wire _2152_;
  wire _2153_;
  wire _2154_;
  wire _2155_;
  wire _2156_;
  wire _2157_;
  wire _2158_;
  wire _2159_;
  wire _2160_;
  wire _2161_;
  wire _2162_;
  wire _2163_;
  wire _2164_;
  wire _2165_;
  wire _2166_;
  wire _2167_;
  wire _2168_;
  wire _2169_;
  wire _2170_;
  wire _2171_;
  wire _2172_;
  wire _2173_;
  wire _2174_;
  wire _2175_;
  wire _2176_;
  wire _2177_;
  wire _2178_;
  wire _2179_;
  wire _2180_;
  wire _2181_;
  wire _2182_;
  wire _2183_;
  wire _2184_;
  wire _2185_;
  wire _2186_;
  wire _2187_;
  wire _2188_;
  wire _2189_;
  wire _2190_;
  wire _2191_;
  wire _2192_;
  wire _2193_;
  wire _2194_;
  wire _2195_;
  wire _2196_;
  wire _2197_;
  wire _2198_;
  wire _2199_;
  wire _2200_;
  wire _2201_;
  wire _2202_;
  wire _2203_;
  wire _2204_;
  wire _2205_;
  wire _2206_;
  wire _2207_;
  wire _2208_;
  wire _2209_;
  wire _2210_;
  wire _2211_;
  wire _2212_;
  wire _2213_;
  wire _2214_;
  wire _2215_;
  wire _2216_;
  wire _2217_;
  wire _2218_;
  wire _2219_;
  wire _2220_;
  wire _2221_;
  wire _2222_;
  wire _2223_;
  wire _2224_;
  wire _2225_;
  wire _2226_;
  wire _2227_;
  wire _2228_;
  wire _2229_;
  wire _2230_;
  wire _2231_;
  wire _2232_;
  wire _2233_;
  wire _2234_;
  wire _2235_;
  wire _2236_;
  wire _2237_;
  wire _2238_;
  wire _2239_;
  wire _2240_;
  wire _2241_;
  wire _2242_;
  wire _2243_;
  wire _2244_;
  wire _2245_;
  wire _2246_;
  wire _2247_;
  wire _2248_;
  wire _2249_;
  wire _2250_;
  wire _2251_;
  wire _2252_;
  wire _2253_;
  wire _2254_;
  wire _2255_;
  wire _2256_;
  wire _2257_;
  wire _2258_;
  wire _2259_;
  wire _2260_;
  wire _2261_;
  wire _2262_;
  wire _2263_;
  wire _2264_;
  wire _2265_;
  wire _2266_;
  wire _2267_;
  wire _2268_;
  wire _2269_;
  wire _2270_;
  wire _2271_;
  wire _2272_;
  wire _2273_;
  wire _2274_;
  wire _2275_;
  wire _2276_;
  wire _2277_;
  wire _2278_;
  wire _2279_;
  wire _2280_;
  wire _2281_;
  wire _2282_;
  wire _2283_;
  wire _2284_;
  wire _2285_;
  wire _2286_;
  wire _2287_;
  wire _2288_;
  wire _2289_;
  wire _2290_;
  wire _2291_;
  wire _2292_;
  wire _2293_;
  wire _2294_;
  wire _2295_;
  wire _2296_;
  wire _2297_;
  wire _2298_;
  wire _2299_;
  wire _2300_;
  wire _2301_;
  wire _2302_;
  wire _2303_;
  wire _2304_;
  wire _2305_;
  wire _2306_;
  wire _2307_;
  wire _2308_;
  wire _2309_;
  wire _2310_;
  wire _2311_;
  wire _2312_;
  wire _2313_;
  wire _2314_;
  wire _2315_;
  wire _2316_;
  wire _2317_;
  wire _2318_;
  wire _2319_;
  wire _2320_;
  wire _2321_;
  wire _2322_;
  wire _2323_;
  wire _2324_;
  wire _2325_;
  wire _2326_;
  wire _2327_;
  wire _2328_;
  wire _2329_;
  wire _2330_;
  wire _2331_;
  wire _2332_;
  wire _2333_;
  wire _2334_;
  wire _2335_;
  wire _2336_;
  wire _2337_;
  wire _2338_;
  wire _2339_;
  wire _2340_;
  wire _2341_;
  wire _2342_;
  wire _2343_;
  wire _2344_;
  wire _2345_;
  wire _2346_;
  wire _2347_;
  wire _2348_;
  wire _2349_;
  wire _2350_;
  wire _2351_;
  wire _2352_;
  wire _2353_;
  wire _2354_;
  wire _2355_;
  wire _2356_;
  wire _2357_;
  wire _2358_;
  wire _2359_;
  wire _2360_;
  wire _2361_;
  wire _2362_;
  wire _2363_;
  wire _2364_;
  wire _2365_;
  wire _2366_;
  wire _2367_;
  wire _2368_;
  wire _2369_;
  wire _2370_;
  wire _2371_;
  wire _2372_;
  wire _2373_;
  wire _2374_;
  wire _2375_;
  wire _2376_;
  wire _2377_;
  wire _2378_;
  wire _2379_;
  wire _2380_;
  wire _2381_;
  wire _2382_;
  wire _2383_;
  wire _2384_;
  wire _2385_;
  wire _2386_;
  wire _2387_;
  wire _2388_;
  wire _2389_;
  wire _2390_;
  wire _2391_;
  wire _2392_;
  wire _2393_;
  wire _2394_;
  wire _2395_;
  wire _2396_;
  wire _2397_;
  wire _2398_;
  wire _2399_;
  wire _2400_;
  wire _2401_;
  wire _2402_;
  wire _2403_;
  wire _2404_;
  wire _2405_;
  wire _2406_;
  wire _2407_;
  wire _2408_;
  wire _2409_;
  wire _2410_;
  wire _2411_;
  wire _2412_;
  wire _2413_;
  wire _2414_;
  wire _2415_;
  wire _2416_;
  wire _2417_;
  wire _2418_;
  wire _2419_;
  wire _2420_;
  wire _2421_;
  wire _2422_;
  wire _2423_;
  wire _2424_;
  wire _2425_;
  wire _2426_;
  wire _2427_;
  wire _2428_;
  wire _2429_;
  wire _2430_;
  wire _2431_;
  wire _2432_;
  wire _2433_;
  wire _2434_;
  wire _2435_;
  wire _2436_;
  wire _2437_;
  wire _2438_;
  wire _2439_;
  wire _2440_;
  wire _2441_;
  wire _2442_;
  wire _2443_;
  wire _2444_;
  wire _2445_;
  wire _2446_;
  wire _2447_;
  wire _2448_;
  wire _2449_;
  wire _2450_;
  wire _2451_;
  wire _2452_;
  wire _2453_;
  wire _2454_;
  wire _2455_;
  wire _2456_;
  wire _2457_;
  wire _2458_;
  wire _2459_;
  wire _2460_;
  wire _2461_;
  wire _2462_;
  wire _2463_;
  wire _2464_;
  wire _2465_;
  wire _2466_;
  wire _2467_;
  wire _2468_;
  wire _2469_;
  wire _2470_;
  wire _2471_;
  wire _2472_;
  wire _2473_;
  wire _2474_;
  wire _2475_;
  wire _2476_;
  wire _2477_;
  wire _2478_;
  wire _2479_;
  wire _2480_;
  wire _2481_;
  wire _2482_;
  wire _2483_;
  wire _2484_;
  wire _2485_;
  wire _2486_;
  wire _2487_;
  wire _2488_;
  wire _2489_;
  wire _2490_;
  wire _2491_;
  wire _2492_;
  wire _2493_;
  wire _2494_;
  wire _2495_;
  wire _2496_;
  wire _2497_;
  wire _2498_;
  wire _2499_;
  wire _2500_;
  wire _2501_;
  wire _2502_;
  wire _2503_;
  wire _2504_;
  wire _2505_;
  wire _2506_;
  wire _2507_;
  wire _2508_;
  wire _2509_;
  wire _2510_;
  wire _2511_;
  wire _2512_;
  wire _2513_;
  wire _2514_;
  wire _2515_;
  wire _2516_;
  wire _2517_;
  wire _2518_;
  wire _2519_;
  wire _2520_;
  wire _2521_;
  wire _2522_;
  wire _2523_;
  wire _2524_;
  wire _2525_;
  wire _2526_;
  wire _2527_;
  wire _2528_;
  wire _2529_;
  wire _2530_;
  wire _2531_;
  wire _2532_;
  wire _2533_;
  wire _2534_;
  wire _2535_;
  wire _2536_;
  wire _2537_;
  wire _2538_;
  wire _2539_;
  wire _2540_;
  wire _2541_;
  wire _2542_;
  wire _2543_;
  wire _2544_;
  wire _2545_;
  wire _2546_;
  wire _2547_;
  wire _2548_;
  wire _2549_;
  wire _2550_;
  wire _2551_;
  wire _2552_;
  wire _2553_;
  wire _2554_;
  wire _2555_;
  wire _2556_;
  wire _2557_;
  wire _2558_;
  wire _2559_;
  wire _2560_;
  wire _2561_;
  wire _2562_;
  wire _2563_;
  wire _2564_;
  wire _2565_;
  wire _2566_;
  wire _2567_;
  wire _2568_;
  wire _2569_;
  wire _2570_;
  wire _2571_;
  wire _2572_;
  wire _2573_;
  wire _2574_;
  wire _2575_;
  wire _2576_;
  wire _2577_;
  wire _2578_;
  wire _2579_;
  wire _2580_;
  wire _2581_;
  wire _2582_;
  wire _2583_;
  wire _2584_;
  wire _2585_;
  wire _2586_;
  wire _2587_;
  wire _2588_;
  wire _2589_;
  wire _2590_;
  wire _2591_;
  wire _2592_;
  wire _2593_;
  wire _2594_;
  wire _2595_;
  wire _2596_;
  wire _2597_;
  wire _2598_;
  wire _2599_;
  wire _2600_;
  wire _2601_;
  wire _2602_;
  wire _2603_;
  wire _2604_;
  wire _2605_;
  wire _2606_;
  wire _2607_;
  wire _2608_;
  wire _2609_;
  wire _2610_;
  wire _2611_;
  wire _2612_;
  wire _2613_;
  wire _2614_;
  wire _2615_;
  wire _2616_;
  wire _2617_;
  wire _2618_;
  wire _2619_;
  wire _2620_;
  wire _2621_;
  wire _2622_;
  wire _2623_;
  wire _2624_;
  wire _2625_;
  wire _2626_;
  wire _2627_;
  wire _2628_;
  wire _2629_;
  wire _2630_;
  wire _2631_;
  wire _2632_;
  wire _2633_;
  wire _2634_;
  wire _2635_;
  wire _2636_;
  wire _2637_;
  wire _2638_;
  wire _2639_;
  wire _2640_;
  wire _2641_;
  wire _2642_;
  wire _2643_;
  wire _2644_;
  wire _2645_;
  wire _2646_;
  wire _2647_;
  wire _2648_;
  wire _2649_;
  wire _2650_;
  wire _2651_;
  wire _2652_;
  wire _2653_;
  wire _2654_;
  wire _2655_;
  wire _2656_;
  wire _2657_;
  wire _2658_;
  wire _2659_;
  wire _2660_;
  wire _2661_;
  wire _2662_;
  wire _2663_;
  wire _2664_;
  wire _2665_;
  wire _2666_;
  wire _2667_;
  wire _2668_;
  wire _2669_;
  wire _2670_;
  wire _2671_;
  wire _2672_;
  wire _2673_;
  wire _2674_;
  wire _2675_;
  wire _2676_;
  wire _2677_;
  wire _2678_;
  wire _2679_;
  wire _2680_;
  wire _2681_;
  wire _2682_;
  wire _2683_;
  wire _2684_;
  wire _2685_;
  wire _2686_;
  wire _2687_;
  wire _2688_;
  wire _2689_;
  wire _2690_;
  wire _2691_;
  wire _2692_;
  wire _2693_;
  wire _2694_;
  wire _2695_;
  wire _2696_;
  wire _2697_;
  wire _2698_;
  wire _2699_;
  wire _2700_;
  wire _2701_;
  wire _2702_;
  wire _2703_;
  wire _2704_;
  wire _2705_;
  wire _2706_;
  wire _2707_;
  wire _2708_;
  wire _2709_;
  wire _2710_;
  wire _2711_;
  wire _2712_;
  wire _2713_;
  wire _2714_;
  wire _2715_;
  wire _2716_;
  wire _2717_;
  wire _2718_;
  wire _2719_;
  wire _2720_;
  wire _2721_;
  wire _2722_;
  wire _2723_;
  wire _2724_;
  wire _2725_;
  wire _2726_;
  wire _2727_;
  wire _2728_;
  wire _2729_;
  wire _2730_;
  wire _2731_;
  wire _2732_;
  wire _2733_;
  wire _2734_;
  wire _2735_;
  wire _2736_;
  wire _2737_;
  wire _2738_;
  wire _2739_;
  wire _2740_;
  wire _2741_;
  wire _2742_;
  wire _2743_;
  wire _2744_;
  wire _2745_;
  wire _2746_;
  wire _2747_;
  wire _2748_;
  wire _2749_;
  wire _2750_;
  wire _2751_;
  wire _2752_;
  wire _2753_;
  wire _2754_;
  wire _2755_;
  wire _2756_;
  wire _2757_;
  wire _2758_;
  wire _2759_;
  wire _2760_;
  wire _2761_;
  wire _2762_;
  wire _2763_;
  wire _2764_;
  wire _2765_;
  wire _2766_;
  wire _2767_;
  wire _2768_;
  wire _2769_;
  wire _2770_;
  wire _2771_;
  wire _2772_;
  wire _2773_;
  wire _2774_;
  wire _2775_;
  wire _2776_;
  wire _2777_;
  wire _2778_;
  wire _2779_;
  wire _2780_;
  wire _2781_;
  wire _2782_;
  wire _2783_;
  wire _2784_;
  wire _2785_;
  wire _2786_;
  wire _2787_;
  wire _2788_;
  wire _2789_;
  wire _2790_;
  wire _2791_;
  wire _2792_;
  wire _2793_;
  wire _2794_;
  wire _2795_;
  wire _2796_;
  wire _2797_;
  wire _2798_;
  wire _2799_;
  wire _2800_;
  wire _2801_;
  wire _2802_;
  wire _2803_;
  wire _2804_;
  wire _2805_;
  wire _2806_;
  wire _2807_;
  wire _2808_;
  wire _2809_;
  wire _2810_;
  wire _2811_;
  wire _2812_;
  wire _2813_;
  wire _2814_;
  wire _2815_;
  wire _2816_;
  wire _2817_;
  wire _2818_;
  wire _2819_;
  wire _2820_;
  wire _2821_;
  wire _2822_;
  wire _2823_;
  wire _2824_;
  wire _2825_;
  wire _2826_;
  wire _2827_;
  wire _2828_;
  wire _2829_;
  wire _2830_;
  wire _2831_;
  wire _2832_;
  wire _2833_;
  wire _2834_;
  wire _2835_;
  wire _2836_;
  wire _2837_;
  wire _2838_;
  wire _2839_;
  wire _2840_;
  wire _2841_;
  wire _2842_;
  wire _2843_;
  wire _2844_;
  wire _2845_;
  wire _2846_;
  wire _2847_;
  wire _2848_;
  wire _2849_;
  wire _2850_;
  wire _2851_;
  wire _2852_;
  wire _2853_;
  wire _2854_;
  wire _2855_;
  wire _2856_;
  wire _2857_;
  wire _2858_;
  wire _2859_;
  wire _2860_;
  wire _2861_;
  wire _2862_;
  wire _2863_;
  wire _2864_;
  wire _2865_;
  wire _2866_;
  wire _2867_;
  wire _2868_;
  wire _2869_;
  wire _2870_;
  wire _2871_;
  wire _2872_;
  wire _2873_;
  wire _2874_;
  wire _2875_;
  wire _2876_;
  wire _2877_;
  wire _2878_;
  wire _2879_;
  wire _2880_;
  wire _2881_;
  wire _2882_;
  wire _2883_;
  wire _2884_;
  wire _2885_;
  wire _2886_;
  wire _2887_;
  wire _2888_;
  wire _2889_;
  wire _2890_;
  wire _2891_;
  wire _2892_;
  wire _2893_;
  wire _2894_;
  wire _2895_;
  wire _2896_;
  wire _2897_;
  wire _2898_;
  wire _2899_;
  wire _2900_;
  wire _2901_;
  wire _2902_;
  wire _2903_;
  wire _2904_;
  wire _2905_;
  wire _2906_;
  wire _2907_;
  wire _2908_;
  wire _2909_;
  wire _2910_;
  wire _2911_;
  wire _2912_;
  wire _2913_;
  wire _2914_;
  wire _2915_;
  wire _2916_;
  wire _2917_;
  wire _2918_;
  wire _2919_;
  wire _2920_;
  wire _2921_;
  wire _2922_;
  wire _2923_;
  wire _2924_;
  wire _2925_;
  wire _2926_;
  wire _2927_;
  wire _2928_;
  wire _2929_;
  wire _2930_;
  wire _2931_;
  wire _2932_;
  wire _2933_;
  wire _2934_;
  wire _2935_;
  wire _2936_;
  wire _2937_;
  wire _2938_;
  wire _2939_;
  wire _2940_;
  wire _2941_;
  wire _2942_;
  wire _2943_;
  wire _2944_;
  wire _2945_;
  wire _2946_;
  wire _2947_;
  wire _2948_;
  wire _2949_;
  wire _2950_;
  wire _2951_;
  wire _2952_;
  wire _2953_;
  wire _2954_;
  wire _2955_;
  wire _2956_;
  wire _2957_;
  wire _2958_;
  wire _2959_;
  wire _2960_;
  wire _2961_;
  wire _2962_;
  wire _2963_;
  wire _2964_;
  wire _2965_;
  wire _2966_;
  wire _2967_;
  wire _2968_;
  wire _2969_;
  wire _2970_;
  wire _2971_;
  wire _2972_;
  wire _2973_;
  wire _2974_;
  wire _2975_;
  wire _2976_;
  wire _2977_;
  wire _2978_;
  wire _2979_;
  wire _2980_;
  wire _2981_;
  wire _2982_;
  wire _2983_;
  wire _2984_;
  wire _2985_;
  wire _2986_;
  wire _2987_;
  wire _2988_;
  wire _2989_;
  wire _2990_;
  wire _2991_;
  wire _2992_;
  wire _2993_;
  wire _2994_;
  wire _2995_;
  wire _2996_;
  wire _2997_;
  wire _2998_;
  wire _2999_;
  wire _3000_;
  wire _3001_;
  wire _3002_;
  wire _3003_;
  wire _3004_;
  wire _3005_;
  wire _3006_;
  wire _3007_;
  wire _3008_;
  wire _3009_;
  wire _3010_;
  wire _3011_;
  wire _3012_;
  wire _3013_;
  wire _3014_;
  wire _3015_;
  wire _3016_;
  wire _3017_;
  wire _3018_;
  wire _3019_;
  wire _3020_;
  wire _3021_;
  wire _3022_;
  wire _3023_;
  wire _3024_;
  wire _3025_;
  wire _3026_;
  wire _3027_;
  wire _3028_;
  wire _3029_;
  wire _3030_;
  wire _3031_;
  wire _3032_;
  wire _3033_;
  wire _3034_;
  wire _3035_;
  wire _3036_;
  wire _3037_;
  wire _3038_;
  wire _3039_;
  wire _3040_;
  wire _3041_;
  wire _3042_;
  wire _3043_;
  wire _3044_;
  wire _3045_;
  wire _3046_;
  wire _3047_;
  wire _3048_;
  wire _3049_;
  wire _3050_;
  wire _3051_;
  wire _3052_;
  wire _3053_;
  wire _3054_;
  wire _3055_;
  wire _3056_;
  wire _3057_;
  wire _3058_;
  wire _3059_;
  wire _3060_;
  wire _3061_;
  wire _3062_;
  wire _3063_;
  wire _3064_;
  wire _3065_;
  wire _3066_;
  wire _3067_;
  wire _3068_;
  wire _3069_;
  wire _3070_;
  wire _3071_;
  wire _3072_;
  wire _3073_;
  wire _3074_;
  wire _3075_;
  wire _3076_;
  wire _3077_;
  wire _3078_;
  wire _3079_;
  wire _3080_;
  wire _3081_;
  wire _3082_;
  wire _3083_;
  wire _3084_;
  wire _3085_;
  wire _3086_;
  wire _3087_;
  wire _3088_;
  wire _3089_;
  wire _3090_;
  wire _3091_;
  wire _3092_;
  wire _3093_;
  wire _3094_;
  wire _3095_;
  wire _3096_;
  wire _3097_;
  wire _3098_;
  wire _3099_;
  wire _3100_;
  wire _3101_;
  wire _3102_;
  wire _3103_;
  wire _3104_;
  wire _3105_;
  wire _3106_;
  wire _3107_;
  wire _3108_;
  wire _3109_;
  wire _3110_;
  wire _3111_;
  wire _3112_;
  wire _3113_;
  wire _3114_;
  wire _3115_;
  wire _3116_;
  wire _3117_;
  wire _3118_;
  wire _3119_;
  wire _3120_;
  wire _3121_;
  wire _3122_;
  wire _3123_;
  wire _3124_;
  wire _3125_;
  wire _3126_;
  wire _3127_;
  wire _3128_;
  wire _3129_;
  wire _3130_;
  wire _3131_;
  wire _3132_;
  wire _3133_;
  wire _3134_;
  wire _3135_;
  wire _3136_;
  wire _3137_;
  wire _3138_;
  wire _3139_;
  wire _3140_;
  wire _3141_;
  wire _3142_;
  wire _3143_;
  wire _3144_;
  wire _3145_;
  wire _3146_;
  wire _3147_;
  wire _3148_;
  wire _3149_;
  wire _3150_;
  wire _3151_;
  wire _3152_;
  wire _3153_;
  wire _3154_;
  wire _3155_;
  wire _3156_;
  wire _3157_;
  wire _3158_;
  wire _3159_;
  wire _3160_;
  wire _3161_;
  wire _3162_;
  wire _3163_;
  wire _3164_;
  wire _3165_;
  wire _3166_;
  wire _3167_;
  wire _3168_;
  wire _3169_;
  wire _3170_;
  wire _3171_;
  wire _3172_;
  wire _3173_;
  wire _3174_;
  wire _3175_;
  wire _3176_;
  wire _3177_;
  wire _3178_;
  wire _3179_;
  wire _3180_;
  wire _3181_;
  wire _3182_;
  wire _3183_;
  wire _3184_;
  wire _3185_;
  wire _3186_;
  wire _3187_;
  wire _3188_;
  wire _3189_;
  wire _3190_;
  wire _3191_;
  wire _3192_;
  wire _3193_;
  wire _3194_;
  wire _3195_;
  wire _3196_;
  wire _3197_;
  wire _3198_;
  wire _3199_;
  wire _3200_;
  wire _3201_;
  wire _3202_;
  wire _3203_;
  wire _3204_;
  wire _3205_;
  wire _3206_;
  wire _3207_;
  wire _3208_;
  wire _3209_;
  wire _3210_;
  wire _3211_;
  wire _3212_;
  wire _3213_;
  wire _3214_;
  wire _3215_;
  wire _3216_;
  wire _3217_;
  wire _3218_;
  wire _3219_;
  wire _3220_;
  wire _3221_;
  wire _3222_;
  wire _3223_;
  wire _3224_;
  wire _3225_;
  wire _3226_;
  wire _3227_;
  wire _3228_;
  wire _3229_;
  wire _3230_;
  wire _3231_;
  wire _3232_;
  wire _3233_;
  wire _3234_;
  wire _3235_;
  wire _3236_;
  wire _3237_;
  wire _3238_;
  wire _3239_;
  wire _3240_;
  wire _3241_;
  wire _3242_;
  wire _3243_;
  wire _3244_;
  wire _3245_;
  wire _3246_;
  wire _3247_;
  wire _3248_;
  wire _3249_;
  wire _3250_;
  wire _3251_;
  wire _3252_;
  wire _3253_;
  wire _3254_;
  wire _3255_;
  wire _3256_;
  wire _3257_;
  wire _3258_;
  wire _3259_;
  wire _3260_;
  wire _3261_;
  wire _3262_;
  wire _3263_;
  wire _3264_;
  wire _3265_;
  wire _3266_;
  wire _3267_;
  wire _3268_;
  wire _3269_;
  wire _3270_;
  wire _3271_;
  wire _3272_;
  wire _3273_;
  wire _3274_;
  wire _3275_;
  wire _3276_;
  wire _3277_;
  wire _3278_;
  wire _3279_;
  wire _3280_;
  wire _3281_;
  wire _3282_;
  wire _3283_;
  wire _3284_;
  wire _3285_;
  wire _3286_;
  wire _3287_;
  wire _3288_;
  wire _3289_;
  wire _3290_;
  wire _3291_;
  wire _3292_;
  wire _3293_;
  wire _3294_;
  wire _3295_;
  wire _3296_;
  wire _3297_;
  wire _3298_;
  wire _3299_;
  wire _3300_;
  wire _3301_;
  wire _3302_;
  wire _3303_;
  wire _3304_;
  wire _3305_;
  wire _3306_;
  wire _3307_;
  wire _3308_;
  wire _3309_;
  wire _3310_;
  wire _3311_;
  wire _3312_;
  wire _3313_;
  wire _3314_;
  wire _3315_;
  wire _3316_;
  wire _3317_;
  wire _3318_;
  wire _3319_;
  wire _3320_;
  wire _3321_;
  wire _3322_;
  wire _3323_;
  wire _3324_;
  wire _3325_;
  wire _3326_;
  wire _3327_;
  wire _3328_;
  wire _3329_;
  wire _3330_;
  wire _3331_;
  wire _3332_;
  wire _3333_;
  wire _3334_;
  wire _3335_;
  wire _3336_;
  wire _3337_;
  wire _3338_;
  wire _3339_;
  wire _3340_;
  wire _3341_;
  wire _3342_;
  wire _3343_;
  wire _3344_;
  wire _3345_;
  wire _3346_;
  wire _3347_;
  wire _3348_;
  wire _3349_;
  wire _3350_;
  wire _3351_;
  wire _3352_;
  wire _3353_;
  wire _3354_;
  wire _3355_;
  wire _3356_;
  wire _3357_;
  wire _3358_;
  wire _3359_;
  wire _3360_;
  wire _3361_;
  wire _3362_;
  wire _3363_;
  wire _3364_;
  wire _3365_;
  wire _3366_;
  wire _3367_;
  wire _3368_;
  wire _3369_;
  wire _3370_;
  wire _3371_;
  wire _3372_;
  wire _3373_;
  wire _3374_;
  wire _3375_;
  wire _3376_;
  wire _3377_;
  wire _3378_;
  wire _3379_;
  wire _3380_;
  wire _3381_;
  wire _3382_;
  wire _3383_;
  wire _3384_;
  wire _3385_;
  wire _3386_;
  wire _3387_;
  wire _3388_;
  wire _3389_;
  wire _3390_;
  wire _3391_;
  wire _3392_;
  wire _3393_;
  wire _3394_;
  wire _3395_;
  wire _3396_;
  wire _3397_;
  wire _3398_;
  wire _3399_;
  wire _3400_;
  wire _3401_;
  wire _3402_;
  wire _3403_;
  wire _3404_;
  wire _3405_;
  wire _3406_;
  wire _3407_;
  wire _3408_;
  wire _3409_;
  wire _3410_;
  wire _3411_;
  wire _3412_;
  wire _3413_;
  wire _3414_;
  wire _3415_;
  wire _3416_;
  wire _3417_;
  wire _3418_;
  wire _3419_;
  wire _3420_;
  wire _3421_;
  wire _3422_;
  wire _3423_;
  wire _3424_;
  wire _3425_;
  wire _3426_;
  wire _3427_;
  wire _3428_;
  wire _3429_;
  wire _3430_;
  wire _3431_;
  wire _3432_;
  wire _3433_;
  wire _3434_;
  wire _3435_;
  wire _3436_;
  wire _3437_;
  wire _3438_;
  wire _3439_;
  wire _3440_;
  wire _3441_;
  wire _3442_;
  wire _3443_;
  wire _3444_;
  wire _3445_;
  wire _3446_;
  wire _3447_;
  wire _3448_;
  wire _3449_;
  wire _3450_;
  wire _3451_;
  wire _3452_;
  wire _3453_;
  wire _3454_;
  wire _3455_;
  wire _3456_;
  wire _3457_;
  wire _3458_;
  wire _3459_;
  wire _3460_;
  wire _3461_;
  wire _3462_;
  wire _3463_;
  wire _3464_;
  wire _3465_;
  wire _3466_;
  wire _3467_;
  wire _3468_;
  wire _3469_;
  wire _3470_;
  wire _3471_;
  wire _3472_;
  wire _3473_;
  wire _3474_;
  wire _3475_;
  wire _3476_;
  wire _3477_;
  wire _3478_;
  wire _3479_;
  wire _3480_;
  wire _3481_;
  wire _3482_;
  wire _3483_;
  wire _3484_;
  wire _3485_;
  wire _3486_;
  wire _3487_;
  wire _3488_;
  wire _3489_;
  wire _3490_;
  wire _3491_;
  wire _3492_;
  wire _3493_;
  wire _3494_;
  wire _3495_;
  wire _3496_;
  wire _3497_;
  wire _3498_;
  wire _3499_;
  wire _3500_;
  wire _3501_;
  wire _3502_;
  wire _3503_;
  wire _3504_;
  wire _3505_;
  wire _3506_;
  wire _3507_;
  wire _3508_;
  wire _3509_;
  wire _3510_;
  wire _3511_;
  wire _3512_;
  wire _3513_;
  wire _3514_;
  wire _3515_;
  wire _3516_;
  wire _3517_;
  wire _3518_;
  wire _3519_;
  wire _3520_;
  wire _3521_;
  wire _3522_;
  wire _3523_;
  wire _3524_;
  wire _3525_;
  wire _3526_;
  wire _3527_;
  wire _3528_;
  wire _3529_;
  wire _3530_;
  wire _3531_;
  wire _3532_;
  wire _3533_;
  wire _3534_;
  wire _3535_;
  wire _3536_;
  wire _3537_;
  wire _3538_;
  wire _3539_;
  wire _3540_;
  wire _3541_;
  wire _3542_;
  wire _3543_;
  wire _3544_;
  wire _3545_;
  wire _3546_;
  wire _3547_;
  wire _3548_;
  wire _3549_;
  wire _3550_;
  wire _3551_;
  wire _3552_;
  wire _3553_;
  wire _3554_;
  wire _3555_;
  wire _3556_;
  wire _3557_;
  wire _3558_;
  wire _3559_;
  wire _3560_;
  wire _3561_;
  wire _3562_;
  wire _3563_;
  wire _3564_;
  wire _3565_;
  wire _3566_;
  wire _3567_;
  wire _3568_;
  wire _3569_;
  wire _3570_;
  wire _3571_;
  wire _3572_;
  wire _3573_;
  wire _3574_;
  wire _3575_;
  wire _3576_;
  wire _3577_;
  wire _3578_;
  wire _3579_;
  wire _3580_;
  wire _3581_;
  wire _3582_;
  wire _3583_;
  wire _3584_;
  wire _3585_;
  wire _3586_;
  wire _3587_;
  wire _3588_;
  wire _3589_;
  wire _3590_;
  wire _3591_;
  wire _3592_;
  wire _3593_;
  wire _3594_;
  wire _3595_;
  wire _3596_;
  wire _3597_;
  wire _3598_;
  wire _3599_;
  wire _3600_;
  wire _3601_;
  wire _3602_;
  wire _3603_;
  wire _3604_;
  wire _3605_;
  wire _3606_;
  wire _3607_;
  wire _3608_;
  wire _3609_;
  wire _3610_;
  wire _3611_;
  wire _3612_;
  wire _3613_;
  wire _3614_;
  wire _3615_;
  wire _3616_;
  wire _3617_;
  wire _3618_;
  wire _3619_;
  wire _3620_;
  wire _3621_;
  wire _3622_;
  wire _3623_;
  wire _3624_;
  wire _3625_;
  wire _3626_;
  wire _3627_;
  wire _3628_;
  wire _3629_;
  wire _3630_;
  wire _3631_;
  wire _3632_;
  wire _3633_;
  wire _3634_;
  wire _3635_;
  wire _3636_;
  wire _3637_;
  wire _3638_;
  wire _3639_;
  wire _3640_;
  wire _3641_;
  wire _3642_;
  wire _3643_;
  wire _3644_;
  wire _3645_;
  wire _3646_;
  wire _3647_;
  wire _3648_;
  wire _3649_;
  wire _3650_;
  wire _3651_;
  wire _3652_;
  wire _3653_;
  wire _3654_;
  wire _3655_;
  wire _3656_;
  wire _3657_;
  wire _3658_;
  wire _3659_;
  wire _3660_;
  wire _3661_;
  wire _3662_;
  wire _3663_;
  wire _3664_;
  wire _3665_;
  wire _3666_;
  wire _3667_;
  wire _3668_;
  wire _3669_;
  wire _3670_;
  wire _3671_;
  wire _3672_;
  wire _3673_;
  wire _3674_;
  wire _3675_;
  wire _3676_;
  wire _3677_;
  wire _3678_;
  wire _3679_;
  wire _3680_;
  wire _3681_;
  wire _3682_;
  wire _3683_;
  wire _3684_;
  wire _3685_;
  wire _3686_;
  wire _3687_;
  wire _3688_;
  wire _3689_;
  wire _3690_;
  wire _3691_;
  wire _3692_;
  wire _3693_;
  wire _3694_;
  wire _3695_;
  wire _3696_;
  wire _3697_;
  wire _3698_;
  wire _3699_;
  wire _3700_;
  wire _3701_;
  wire _3702_;
  wire _3703_;
  wire _3704_;
  wire _3705_;
  wire _3706_;
  wire _3707_;
  wire _3708_;
  wire _3709_;
  wire _3710_;
  wire _3711_;
  wire _3712_;
  wire _3713_;
  wire _3714_;
  wire _3715_;
  wire _3716_;
  wire _3717_;
  wire _3718_;
  wire _3719_;
  wire _3720_;
  wire _3721_;
  wire _3722_;
  wire _3723_;
  wire _3724_;
  wire _3725_;
  wire _3726_;
  wire _3727_;
  wire _3728_;
  wire _3729_;
  wire _3730_;
  wire _3731_;
  wire _3732_;
  wire _3733_;
  wire _3734_;
  wire _3735_;
  wire _3736_;
  wire _3737_;
  wire _3738_;
  wire _3739_;
  wire _3740_;
  wire _3741_;
  wire _3742_;
  wire _3743_;
  wire _3744_;
  wire _3745_;
  wire _3746_;
  wire _3747_;
  wire _3748_;
  wire _3749_;
  wire _3750_;
  wire _3751_;
  wire _3752_;
  wire _3753_;
  wire _3754_;
  wire _3755_;
  wire _3756_;
  wire _3757_;
  wire _3758_;
  wire _3759_;
  wire _3760_;
  wire _3761_;
  wire _3762_;
  wire _3763_;
  wire _3764_;
  wire _3765_;
  wire _3766_;
  wire _3767_;
  wire _3768_;
  wire _3769_;
  wire _3770_;
  wire _3771_;
  wire _3772_;
  wire _3773_;
  wire _3774_;
  wire _3775_;
  wire _3776_;
  wire _3777_;
  wire _3778_;
  wire _3779_;
  wire _3780_;
  wire _3781_;
  wire _3782_;
  wire _3783_;
  wire _3784_;
  wire _3785_;
  wire _3786_;
  wire _3787_;
  wire _3788_;
  wire _3789_;
  wire _3790_;
  wire _3791_;
  wire _3792_;
  wire _3793_;
  wire _3794_;
  wire _3795_;
  wire _3796_;
  wire _3797_;
  wire _3798_;
  wire _3799_;
  wire _3800_;
  wire _3801_;
  wire _3802_;
  wire _3803_;
  wire _3804_;
  wire _3805_;
  wire _3806_;
  wire _3807_;
  wire _3808_;
  wire _3809_;
  wire _3810_;
  wire _3811_;
  wire _3812_;
  wire _3813_;
  wire _3814_;
  wire _3815_;
  wire _3816_;
  wire _3817_;
  wire _3818_;
  wire _3819_;
  wire _3820_;
  wire _3821_;
  wire _3822_;
  wire _3823_;
  wire _3824_;
  wire _3825_;
  wire _3826_;
  wire _3827_;
  wire _3828_;
  wire _3829_;
  wire _3830_;
  wire _3831_;
  wire _3832_;
  wire _3833_;
  wire _3834_;
  wire _3835_;
  wire _3836_;
  wire _3837_;
  wire _3838_;
  wire _3839_;
  wire _3840_;
  wire _3841_;
  wire _3842_;
  wire _3843_;
  wire _3844_;
  wire _3845_;
  wire _3846_;
  wire _3847_;
  wire _3848_;
  wire _3849_;
  wire _3850_;
  wire _3851_;
  wire _3852_;
  wire _3853_;
  wire _3854_;
  wire _3855_;
  wire _3856_;
  wire _3857_;
  wire _3858_;
  wire _3859_;
  wire _3860_;
  wire _3861_;
  wire _3862_;
  wire _3863_;
  wire _3864_;
  wire _3865_;
  wire _3866_;
  wire _3867_;
  wire _3868_;
  wire _3869_;
  wire _3870_;
  wire _3871_;
  wire _3872_;
  wire _3873_;
  wire _3874_;
  wire _3875_;
  wire _3876_;
  wire _3877_;
  wire _3878_;
  wire _3879_;
  wire _3880_;
  wire _3881_;
  wire _3882_;
  wire _3883_;
  wire _3884_;
  wire _3885_;
  wire _3886_;
  wire _3887_;
  wire _3888_;
  wire _3889_;
  wire _3890_;
  wire _3891_;
  wire _3892_;
  wire _3893_;
  wire _3894_;
  wire _3895_;
  wire _3896_;
  wire _3897_;
  wire _3898_;
  wire _3899_;
  wire _3900_;
  wire _3901_;
  wire _3902_;
  wire _3903_;
  wire _3904_;
  wire _3905_;
  wire _3906_;
  wire _3907_;
  wire _3908_;
  wire _3909_;
  wire _3910_;
  wire _3911_;
  wire _3912_;
  wire _3913_;
  wire _3914_;
  wire _3915_;
  wire _3916_;
  wire _3917_;
  wire _3918_;
  wire _3919_;
  wire _3920_;
  wire _3921_;
  wire _3922_;
  wire _3923_;
  wire _3924_;
  wire _3925_;
  wire _3926_;
  wire _3927_;
  wire _3928_;
  wire _3929_;
  wire _3930_;
  wire _3931_;
  wire _3932_;
  wire _3933_;
  wire _3934_;
  wire _3935_;
  wire _3936_;
  wire _3937_;
  wire _3938_;
  wire _3939_;
  wire _3940_;
  wire _3941_;
  wire _3942_;
  wire _3943_;
  wire _3944_;
  wire _3945_;
  wire _3946_;
  wire _3947_;
  wire _3948_;
  wire _3949_;
  wire _3950_;
  wire _3951_;
  wire _3952_;
  wire _3953_;
  wire _3954_;
  wire _3955_;
  wire _3956_;
  wire _3957_;
  wire _3958_;
  wire _3959_;
  wire _3960_;
  wire _3961_;
  wire _3962_;
  wire _3963_;
  wire _3964_;
  wire _3965_;
  wire _3966_;
  wire _3967_;
  wire _3968_;
  wire _3969_;
  wire _3970_;
  wire _3971_;
  wire _3972_;
  wire _3973_;
  wire _3974_;
  wire _3975_;
  wire _3976_;
  wire _3977_;
  wire _3978_;
  wire _3979_;
  wire _3980_;
  wire _3981_;
  wire _3982_;
  wire _3983_;
  wire _3984_;
  wire _3985_;
  wire _3986_;
  wire _3987_;
  wire _3988_;
  wire _3989_;
  wire _3990_;
  wire _3991_;
  wire _3992_;
  wire _3993_;
  wire _3994_;
  wire _3995_;
  wire _3996_;
  wire _3997_;
  wire _3998_;
  wire _3999_;
  wire _4000_;
  wire _4001_;
  wire _4002_;
  wire _4003_;
  wire _4004_;
  wire _4005_;
  wire _4006_;
  wire _4007_;
  wire _4008_;
  wire _4009_;
  wire _4010_;
  wire _4011_;
  wire _4012_;
  wire _4013_;
  wire _4014_;
  wire _4015_;
  wire _4016_;
  wire _4017_;
  wire _4018_;
  wire _4019_;
  wire _4020_;
  wire _4021_;
  wire _4022_;
  wire _4023_;
  wire _4024_;
  wire _4025_;
  wire _4026_;
  wire _4027_;
  wire _4028_;
  wire _4029_;
  wire _4030_;
  wire _4031_;
  wire _4032_;
  wire _4033_;
  wire _4034_;
  wire _4035_;
  wire _4036_;
  wire _4037_;
  wire _4038_;
  wire _4039_;
  wire _4040_;
  wire _4041_;
  wire _4042_;
  wire _4043_;
  wire _4044_;
  wire _4045_;
  wire _4046_;
  wire _4047_;
  wire _4048_;
  wire _4049_;
  wire _4050_;
  wire _4051_;
  wire _4052_;
  wire _4053_;
  wire _4054_;
  wire _4055_;
  wire _4056_;
  wire _4057_;
  wire _4058_;
  wire _4059_;
  wire _4060_;
  wire _4061_;
  wire _4062_;
  wire _4063_;
  wire _4064_;
  wire _4065_;
  wire _4066_;
  wire _4067_;
  wire _4068_;
  wire _4069_;
  wire _4070_;
  wire _4071_;
  wire _4072_;
  wire _4073_;
  wire _4074_;
  wire _4075_;
  wire _4076_;
  wire _4077_;
  wire _4078_;
  wire _4079_;
  wire _4080_;
  wire _4081_;
  wire _4082_;
  wire _4083_;
  wire _4084_;
  wire _4085_;
  wire _4086_;
  wire _4087_;
  wire _4088_;
  wire _4089_;
  wire _4090_;
  wire _4091_;
  wire _4092_;
  wire _4093_;
  wire _4094_;
  wire _4095_;
  wire _4096_;
  wire _4097_;
  wire _4098_;
  wire _4099_;
  wire _4100_;
  wire _4101_;
  wire _4102_;
  wire _4103_;
  wire _4104_;
  wire _4105_;
  wire _4106_;
  wire _4107_;
  wire _4108_;
  wire _4109_;
  wire _4110_;
  wire _4111_;
  wire _4112_;
  wire _4113_;
  wire _4114_;
  wire _4115_;
  wire _4116_;
  wire _4117_;
  wire _4118_;
  wire _4119_;
  wire _4120_;
  wire _4121_;
  wire _4122_;
  wire _4123_;
  wire _4124_;
  wire _4125_;
  wire _4126_;
  wire _4127_;
  wire _4128_;
  wire _4129_;
  wire _4130_;
  wire _4131_;
  wire _4132_;
  wire _4133_;
  wire _4134_;
  wire _4135_;
  wire _4136_;
  wire _4137_;
  wire _4138_;
  wire _4139_;
  wire _4140_;
  wire _4141_;
  wire _4142_;
  wire _4143_;
  wire _4144_;
  wire _4145_;
  wire _4146_;
  wire _4147_;
  wire _4148_;
  wire _4149_;
  wire _4150_;
  wire _4151_;
  wire _4152_;
  wire _4153_;
  wire _4154_;
  wire _4155_;
  wire _4156_;
  wire _4157_;
  wire _4158_;
  wire _4159_;
  wire _4160_;
  wire _4161_;
  wire _4162_;
  wire _4163_;
  wire _4164_;
  wire _4165_;
  wire _4166_;
  wire _4167_;
  wire _4168_;
  wire _4169_;
  wire _4170_;
  wire _4171_;
  wire _4172_;
  wire _4173_;
  wire _4174_;
  wire _4175_;
  wire _4176_;
  wire _4177_;
  wire _4178_;
  wire _4179_;
  wire _4180_;
  wire _4181_;
  wire _4182_;
  wire _4183_;
  wire _4184_;
  wire _4185_;
  wire _4186_;
  wire _4187_;
  wire _4188_;
  wire _4189_;
  wire _4190_;
  wire _4191_;
  wire _4192_;
  wire _4193_;
  wire _4194_;
  wire _4195_;
  wire _4196_;
  wire _4197_;
  wire _4198_;
  wire _4199_;
  wire _4200_;
  wire _4201_;
  wire _4202_;
  wire _4203_;
  wire _4204_;
  wire _4205_;
  wire _4206_;
  wire _4207_;
  wire _4208_;
  wire _4209_;
  wire _4210_;
  wire _4211_;
  wire _4212_;
  wire _4213_;
  wire _4214_;
  wire _4215_;
  wire _4216_;
  wire _4217_;
  wire _4218_;
  wire _4219_;
  wire _4220_;
  wire _4221_;
  wire _4222_;
  wire _4223_;
  wire _4224_;
  wire _4225_;
  wire _4226_;
  wire _4227_;
  wire _4228_;
  wire _4229_;
  wire _4230_;
  wire _4231_;
  wire _4232_;
  wire _4233_;
  wire _4234_;
  wire _4235_;
  wire _4236_;
  wire _4237_;
  wire _4238_;
  wire _4239_;
  wire _4240_;
  wire _4241_;
  wire _4242_;
  wire _4243_;
  wire _4244_;
  wire _4245_;
  wire _4246_;
  wire _4247_;
  wire _4248_;
  wire _4249_;
  wire _4250_;
  wire _4251_;
  wire _4252_;
  wire _4253_;
  wire _4254_;
  wire _4255_;
  wire _4256_;
  wire _4257_;
  wire _4258_;
  wire _4259_;
  wire _4260_;
  wire _4261_;
  wire _4262_;
  wire _4263_;
  wire _4264_;
  wire _4265_;
  wire _4266_;
  wire _4267_;
  wire _4268_;
  wire _4269_;
  wire _4270_;
  wire _4271_;
  wire _4272_;
  wire _4273_;
  wire _4274_;
  wire _4275_;
  wire _4276_;
  wire _4277_;
  wire _4278_;
  wire _4279_;
  wire _4280_;
  wire _4281_;
  wire _4282_;
  wire _4283_;
  wire _4284_;
  wire _4285_;
  wire _4286_;
  wire _4287_;
  wire _4288_;
  wire _4289_;
  wire _4290_;
  wire _4291_;
  wire _4292_;
  wire _4293_;
  wire _4294_;
  wire _4295_;
  wire _4296_;
  wire _4297_;
  wire _4298_;
  wire _4299_;
  wire _4300_;
  wire _4301_;
  wire _4302_;
  wire _4303_;
  wire _4304_;
  wire _4305_;
  wire _4306_;
  wire _4307_;
  wire _4308_;
  wire _4309_;
  wire _4310_;
  wire _4311_;
  wire _4312_;
  wire _4313_;
  wire _4314_;
  wire _4315_;
  wire _4316_;
  wire _4317_;
  wire _4318_;
  wire _4319_;
  wire _4320_;
  wire _4321_;
  wire _4322_;
  wire _4323_;
  wire _4324_;
  wire _4325_;
  wire _4326_;
  wire _4327_;
  wire _4328_;
  wire _4329_;
  wire _4330_;
  wire _4331_;
  wire _4332_;
  wire _4333_;
  wire _4334_;
  wire _4335_;
  wire _4336_;
  wire _4337_;
  wire _4338_;
  wire _4339_;
  wire _4340_;
  wire _4341_;
  wire _4342_;
  wire _4343_;
  wire _4344_;
  wire _4345_;
  wire _4346_;
  wire _4347_;
  wire _4348_;
  wire _4349_;
  wire _4350_;
  wire _4351_;
  wire _4352_;
  wire _4353_;
  wire _4354_;
  wire _4355_;
  wire _4356_;
  wire _4357_;
  wire _4358_;
  wire _4359_;
  wire _4360_;
  wire _4361_;
  wire _4362_;
  wire _4363_;
  wire _4364_;
  wire _4365_;
  wire _4366_;
  wire _4367_;
  wire _4368_;
  wire _4369_;
  wire _4370_;
  wire _4371_;
  wire _4372_;
  wire _4373_;
  wire _4374_;
  wire _4375_;
  wire _4376_;
  wire _4377_;
  wire _4378_;
  wire _4379_;
  wire _4380_;
  wire _4381_;
  wire _4382_;
  wire _4383_;
  wire _4384_;
  wire _4385_;
  wire _4386_;
  wire _4387_;
  wire _4388_;
  wire _4389_;
  wire _4390_;
  wire _4391_;
  wire _4392_;
  wire _4393_;
  wire _4394_;
  wire _4395_;
  wire _4396_;
  wire _4397_;
  wire _4398_;
  wire _4399_;
  wire _4400_;
  wire _4401_;
  wire _4402_;
  wire _4403_;
  wire _4404_;
  wire _4405_;
  wire _4406_;
  wire _4407_;
  wire _4408_;
  wire _4409_;
  wire _4410_;
  wire _4411_;
  wire _4412_;
  wire _4413_;
  wire _4414_;
  wire _4415_;
  wire _4416_;
  wire _4417_;
  wire _4418_;
  wire _4419_;
  wire _4420_;
  wire _4421_;
  wire _4422_;
  wire _4423_;
  wire _4424_;
  wire _4425_;
  wire _4426_;
  wire _4427_;
  wire _4428_;
  wire _4429_;
  wire _4430_;
  wire _4431_;
  wire _4432_;
  wire _4433_;
  wire _4434_;
  wire _4435_;
  wire _4436_;
  wire _4437_;
  wire _4438_;
  wire _4439_;
  wire _4440_;
  wire _4441_;
  wire _4442_;
  wire _4443_;
  wire _4444_;
  wire _4445_;
  wire _4446_;
  wire _4447_;
  wire _4448_;
  wire _4449_;
  wire _4450_;
  wire _4451_;
  wire _4452_;
  wire _4453_;
  wire _4454_;
  wire _4455_;
  wire _4456_;
  wire _4457_;
  wire _4458_;
  wire _4459_;
  wire _4460_;
  wire _4461_;
  wire _4462_;
  wire _4463_;
  wire _4464_;
  wire _4465_;
  wire _4466_;
  wire _4467_;
  wire _4468_;
  wire _4469_;
  wire _4470_;
  wire _4471_;
  wire _4472_;
  wire _4473_;
  wire _4474_;
  wire _4475_;
  wire _4476_;
  wire _4477_;
  wire _4478_;
  wire _4479_;
  wire _4480_;
  wire _4481_;
  wire _4482_;
  wire _4483_;
  wire _4484_;
  wire _4485_;
  wire _4486_;
  wire _4487_;
  wire _4488_;
  wire _4489_;
  wire _4490_;
  wire _4491_;
  wire _4492_;
  wire _4493_;
  wire _4494_;
  wire _4495_;
  wire _4496_;
  wire _4497_;
  wire _4498_;
  wire _4499_;
  wire _4500_;
  wire _4501_;
  wire _4502_;
  wire _4503_;
  wire _4504_;
  wire _4505_;
  wire _4506_;
  wire _4507_;
  wire _4508_;
  wire _4509_;
  wire _4510_;
  wire _4511_;
  wire _4512_;
  wire _4513_;
  wire _4514_;
  wire _4515_;
  wire _4516_;
  wire _4517_;
  wire _4518_;
  wire _4519_;
  wire _4520_;
  wire _4521_;
  wire _4522_;
  wire _4523_;
  wire _4524_;
  wire _4525_;
  wire _4526_;
  wire _4527_;
  wire _4528_;
  wire _4529_;
  wire _4530_;
  wire _4531_;
  wire _4532_;
  wire _4533_;
  wire _4534_;
  wire _4535_;
  wire _4536_;
  wire _4537_;
  wire _4538_;
  wire _4539_;
  wire _4540_;
  wire _4541_;
  wire _4542_;
  wire _4543_;
  wire _4544_;
  wire _4545_;
  wire _4546_;
  wire _4547_;
  wire _4548_;
  wire _4549_;
  wire _4550_;
  wire _4551_;
  wire _4552_;
  wire _4553_;
  wire _4554_;
  wire _4555_;
  wire _4556_;
  wire _4557_;
  wire _4558_;
  wire _4559_;
  wire _4560_;
  wire _4561_;
  wire _4562_;
  wire _4563_;
  wire _4564_;
  wire _4565_;
  wire _4566_;
  wire _4567_;
  wire _4568_;
  wire _4569_;
  wire _4570_;
  wire _4571_;
  wire _4572_;
  wire _4573_;
  wire _4574_;
  wire _4575_;
  wire _4576_;
  wire _4577_;
  wire _4578_;
  wire _4579_;
  wire _4580_;
  wire _4581_;
  wire _4582_;
  wire _4583_;
  wire _4584_;
  wire _4585_;
  wire _4586_;
  wire _4587_;
  wire _4588_;
  wire _4589_;
  wire _4590_;
  wire _4591_;
  wire _4592_;
  wire _4593_;
  wire _4594_;
  wire _4595_;
  wire _4596_;
  wire _4597_;
  wire _4598_;
  wire _4599_;
  wire _4600_;
  wire _4601_;
  wire _4602_;
  wire _4603_;
  wire _4604_;
  wire _4605_;
  wire _4606_;
  wire _4607_;
  wire _4608_;
  wire _4609_;
  wire _4610_;
  wire _4611_;
  wire _4612_;
  wire _4613_;
  wire _4614_;
  wire _4615_;
  wire _4616_;
  wire _4617_;
  wire _4618_;
  wire _4619_;
  wire _4620_;
  wire _4621_;
  wire _4622_;
  wire _4623_;
  wire _4624_;
  wire _4625_;
  wire _4626_;
  wire _4627_;
  wire _4628_;
  wire _4629_;
  wire _4630_;
  wire _4631_;
  wire _4632_;
  wire _4633_;
  wire _4634_;
  wire _4635_;
  wire _4636_;
  wire _4637_;
  wire _4638_;
  wire _4639_;
  wire _4640_;
  wire _4641_;
  wire _4642_;
  wire _4643_;
  wire _4644_;
  wire _4645_;
  wire _4646_;
  wire _4647_;
  wire _4648_;
  wire _4649_;
  wire _4650_;
  wire _4651_;
  wire _4652_;
  wire _4653_;
  wire _4654_;
  wire _4655_;
  wire _4656_;
  wire _4657_;
  wire _4658_;
  wire _4659_;
  wire _4660_;
  wire _4661_;
  wire _4662_;
  wire _4663_;
  wire _4664_;
  wire _4665_;
  wire _4666_;
  wire _4667_;
  wire _4668_;
  wire _4669_;
  wire _4670_;
  wire _4671_;
  wire _4672_;
  wire _4673_;
  wire _4674_;
  wire _4675_;
  wire _4676_;
  wire _4677_;
  wire _4678_;
  wire _4679_;
  wire _4680_;
  wire _4681_;
  wire _4682_;
  wire _4683_;
  wire _4684_;
  wire _4685_;
  wire _4686_;
  wire _4687_;
  wire _4688_;
  wire _4689_;
  wire _4690_;
  wire _4691_;
  wire _4692_;
  wire _4693_;
  wire _4694_;
  wire _4695_;
  wire _4696_;
  wire _4697_;
  wire _4698_;
  wire _4699_;
  wire _4700_;
  wire _4701_;
  wire _4702_;
  wire _4703_;
  wire _4704_;
  wire _4705_;
  wire _4706_;
  wire _4707_;
  wire _4708_;
  wire _4709_;
  wire _4710_;
  wire _4711_;
  wire _4712_;
  wire _4713_;
  wire _4714_;
  wire _4715_;
  wire _4716_;
  wire _4717_;
  wire _4718_;
  wire _4719_;
  wire _4720_;
  wire _4721_;
  wire _4722_;
  wire _4723_;
  wire _4724_;
  wire _4725_;
  wire _4726_;
  wire _4727_;
  wire _4728_;
  wire _4729_;
  wire _4730_;
  wire _4731_;
  wire _4732_;
  wire _4733_;
  wire _4734_;
  wire _4735_;
  wire _4736_;
  wire _4737_;
  wire _4738_;
  wire _4739_;
  wire _4740_;
  wire _4741_;
  wire _4742_;
  wire _4743_;
  wire _4744_;
  wire _4745_;
  wire _4746_;
  wire _4747_;
  wire _4748_;
  wire _4749_;
  wire _4750_;
  wire _4751_;
  wire _4752_;
  wire _4753_;
  wire _4754_;
  wire _4755_;
  wire _4756_;
  wire _4757_;
  wire _4758_;
  wire _4759_;
  wire _4760_;
  wire _4761_;
  wire _4762_;
  wire _4763_;
  wire _4764_;
  wire _4765_;
  wire _4766_;
  wire _4767_;
  wire _4768_;
  wire _4769_;
  wire _4770_;
  wire _4771_;
  wire _4772_;
  wire _4773_;
  wire _4774_;
  wire _4775_;
  wire _4776_;
  wire _4777_;
  wire _4778_;
  wire _4779_;
  wire _4780_;
  wire _4781_;
  wire _4782_;
  wire _4783_;
  wire _4784_;
  wire _4785_;
  wire _4786_;
  wire _4787_;
  wire _4788_;
  wire _4789_;
  wire _4790_;
  wire _4791_;
  wire _4792_;
  wire _4793_;
  wire _4794_;
  wire _4795_;
  wire _4796_;
  wire _4797_;
  wire _4798_;
  wire _4799_;
  wire _4800_;
  wire _4801_;
  wire _4802_;
  wire _4803_;
  wire _4804_;
  wire _4805_;
  wire _4806_;
  wire _4807_;
  wire _4808_;
  wire _4809_;
  wire _4810_;
  wire _4811_;
  wire _4812_;
  wire _4813_;
  wire _4814_;
  wire _4815_;
  wire _4816_;
  wire _4817_;
  wire _4818_;
  wire _4819_;
  wire _4820_;
  wire _4821_;
  wire _4822_;
  wire _4823_;
  wire _4824_;
  wire _4825_;
  wire _4826_;
  wire _4827_;
  wire _4828_;
  wire _4829_;
  wire _4830_;
  wire _4831_;
  wire _4832_;
  wire _4833_;
  wire _4834_;
  wire _4835_;
  wire _4836_;
  wire _4837_;
  wire _4838_;
  wire _4839_;
  wire _4840_;
  wire _4841_;
  wire _4842_;
  wire _4843_;
  wire _4844_;
  wire _4845_;
  wire _4846_;
  wire _4847_;
  wire _4848_;
  wire _4849_;
  wire _4850_;
  wire _4851_;
  wire _4852_;
  wire _4853_;
  wire _4854_;
  wire _4855_;
  wire _4856_;
  wire _4857_;
  wire _4858_;
  wire _4859_;
  wire _4860_;
  wire _4861_;
  wire _4862_;
  wire _4863_;
  wire _4864_;
  wire _4865_;
  wire _4866_;
  wire _4867_;
  wire _4868_;
  wire _4869_;
  wire _4870_;
  wire _4871_;
  wire _4872_;
  wire _4873_;
  wire _4874_;
  wire _4875_;
  wire _4876_;
  wire _4877_;
  wire _4878_;
  wire _4879_;
  wire _4880_;
  wire _4881_;
  wire _4882_;
  wire _4883_;
  wire _4884_;
  wire _4885_;
  wire _4886_;
  wire _4887_;
  wire _4888_;
  wire _4889_;
  wire _4890_;
  wire _4891_;
  wire _4892_;
  wire _4893_;
  wire _4894_;
  wire _4895_;
  wire _4896_;
  wire _4897_;
  wire _4898_;
  wire _4899_;
  wire _4900_;
  wire _4901_;
  wire _4902_;
  wire _4903_;
  wire _4904_;
  wire _4905_;
  wire _4906_;
  wire _4907_;
  wire _4908_;
  wire _4909_;
  wire _4910_;
  wire _4911_;
  wire _4912_;
  wire _4913_;
  wire _4914_;
  wire _4915_;
  wire _4916_;
  wire _4917_;
  wire _4918_;
  wire _4919_;
  wire _4920_;
  wire _4921_;
  wire _4922_;
  wire _4923_;
  wire _4924_;
  wire _4925_;
  wire _4926_;
  wire _4927_;
  wire _4928_;
  wire _4929_;
  wire _4930_;
  wire _4931_;
  wire _4932_;
  wire _4933_;
  wire _4934_;
  wire _4935_;
  wire _4936_;
  wire _4937_;
  wire _4938_;
  wire _4939_;
  wire _4940_;
  wire _4941_;
  wire _4942_;
  wire _4943_;
  wire _4944_;
  wire _4945_;
  wire _4946_;
  wire _4947_;
  wire _4948_;
  wire _4949_;
  wire _4950_;
  wire _4951_;
  wire _4952_;
  wire _4953_;
  wire _4954_;
  wire _4955_;
  wire _4956_;
  wire _4957_;
  wire _4958_;
  wire _4959_;
  wire _4960_;
  wire _4961_;
  wire _4962_;
  wire _4963_;
  wire _4964_;
  wire _4965_;
  wire _4966_;
  wire _4967_;
  wire _4968_;
  wire _4969_;
  wire _4970_;
  wire _4971_;
  wire _4972_;
  wire _4973_;
  wire _4974_;
  wire _4975_;
  wire _4976_;
  wire _4977_;
  wire _4978_;
  wire _4979_;
  wire _4980_;
  wire _4981_;
  wire _4982_;
  wire _4983_;
  wire _4984_;
  wire _4985_;
  wire _4986_;
  wire _4987_;
  wire _4988_;
  wire _4989_;
  wire _4990_;
  wire _4991_;
  wire _4992_;
  wire _4993_;
  wire _4994_;
  wire _4995_;
  wire _4996_;
  wire _4997_;
  wire _4998_;
  wire _4999_;
  wire _5000_;
  wire _5001_;
  wire _5002_;
  wire _5003_;
  wire _5004_;
  wire _5005_;
  wire _5006_;
  wire _5007_;
  wire _5008_;
  wire _5009_;
  wire _5010_;
  wire _5011_;
  wire _5012_;
  wire _5013_;
  wire _5014_;
  wire _5015_;
  wire _5016_;
  wire _5017_;
  wire _5018_;
  wire _5019_;
  wire _5020_;
  wire _5021_;
  wire _5022_;
  wire _5023_;
  wire _5024_;
  wire _5025_;
  wire _5026_;
  wire _5027_;
  wire _5028_;
  wire _5029_;
  wire _5030_;
  wire _5031_;
  wire _5032_;
  wire _5033_;
  wire _5034_;
  wire _5035_;
  wire _5036_;
  wire _5037_;
  wire _5038_;
  wire _5039_;
  wire _5040_;
  wire _5041_;
  wire _5042_;
  wire _5043_;
  wire _5044_;
  wire _5045_;
  wire _5046_;
  wire _5047_;
  wire _5048_;
  wire _5049_;
  wire _5050_;
  wire _5051_;
  wire _5052_;
  wire _5053_;
  wire _5054_;
  wire _5055_;
  wire _5056_;
  wire _5057_;
  wire _5058_;
  wire _5059_;
  wire _5060_;
  wire _5061_;
  wire _5062_;
  wire _5063_;
  wire _5064_;
  wire _5065_;
  wire _5066_;
  wire _5067_;
  wire _5068_;
  wire _5069_;
  wire _5070_;
  wire _5071_;
  wire _5072_;
  wire _5073_;
  wire _5074_;
  wire _5075_;
  wire _5076_;
  wire _5077_;
  wire _5078_;
  wire _5079_;
  wire _5080_;
  wire _5081_;
  wire _5082_;
  wire _5083_;
  wire _5084_;
  wire _5085_;
  wire _5086_;
  wire _5087_;
  wire _5088_;
  wire _5089_;
  wire _5090_;
  wire _5091_;
  wire _5092_;
  wire _5093_;
  wire _5094_;
  wire _5095_;
  wire _5096_;
  wire _5097_;
  wire _5098_;
  wire _5099_;
  wire _5100_;
  wire _5101_;
  wire _5102_;
  wire _5103_;
  wire _5104_;
  wire _5105_;
  wire _5106_;
  wire _5107_;
  wire _5108_;
  wire _5109_;
  wire _5110_;
  wire _5111_;
  wire _5112_;
  wire _5113_;
  wire _5114_;
  wire _5115_;
  wire _5116_;
  wire _5117_;
  wire _5118_;
  wire _5119_;
  wire _5120_;
  wire _5121_;
  wire _5122_;
  wire _5123_;
  wire _5124_;
  wire _5125_;
  wire _5126_;
  wire _5127_;
  wire _5128_;
  wire _5129_;
  wire _5130_;
  wire _5131_;
  wire _5132_;
  wire _5133_;
  wire _5134_;
  wire _5135_;
  wire _5136_;
  wire _5137_;
  wire _5138_;
  wire _5139_;
  wire _5140_;
  wire _5141_;
  wire _5142_;
  wire _5143_;
  wire _5144_;
  wire _5145_;
  wire _5146_;
  wire _5147_;
  wire _5148_;
  wire _5149_;
  wire _5150_;
  wire _5151_;
  wire _5152_;
  wire _5153_;
  wire _5154_;
  wire _5155_;
  wire _5156_;
  wire _5157_;
  wire _5158_;
  wire _5159_;
  wire _5160_;
  wire _5161_;
  wire _5162_;
  wire _5163_;
  wire _5164_;
  wire _5165_;
  wire _5166_;
  wire _5167_;
  wire _5168_;
  wire _5169_;
  wire _5170_;
  wire _5171_;
  wire _5172_;
  wire _5173_;
  wire _5174_;
  wire _5175_;
  wire _5176_;
  wire _5177_;
  wire _5178_;
  wire _5179_;
  wire _5180_;
  wire _5181_;
  wire _5182_;
  wire _5183_;
  wire _5184_;
  wire _5185_;
  wire _5186_;
  wire _5187_;
  wire _5188_;
  wire _5189_;
  wire _5190_;
  wire _5191_;
  wire _5192_;
  wire _5193_;
  wire _5194_;
  wire _5195_;
  wire _5196_;
  wire _5197_;
  wire _5198_;
  wire _5199_;
  wire _5200_;
  wire _5201_;
  wire _5202_;
  wire _5203_;
  wire _5204_;
  wire _5205_;
  wire _5206_;
  wire _5207_;
  wire _5208_;
  wire _5209_;
  wire _5210_;
  wire _5211_;
  wire _5212_;
  wire _5213_;
  wire _5214_;
  wire _5215_;
  wire _5216_;
  wire _5217_;
  wire _5218_;
  wire _5219_;
  wire _5220_;
  wire _5221_;
  wire _5222_;
  wire _5223_;
  wire _5224_;
  wire _5225_;
  wire _5226_;
  wire _5227_;
  wire _5228_;
  wire _5229_;
  wire _5230_;
  wire _5231_;
  wire _5232_;
  wire _5233_;
  wire _5234_;
  wire _5235_;
  wire _5236_;
  wire _5237_;
  wire _5238_;
  wire _5239_;
  wire _5240_;
  wire _5241_;
  wire _5242_;
  wire _5243_;
  wire _5244_;
  wire _5245_;
  wire _5246_;
  wire _5247_;
  wire _5248_;
  wire _5249_;
  wire _5250_;
  wire _5251_;
  wire _5252_;
  wire _5253_;
  wire _5254_;
  wire _5255_;
  wire _5256_;
  wire _5257_;
  wire _5258_;
  wire _5259_;
  wire _5260_;
  wire _5261_;
  wire _5262_;
  wire _5263_;
  wire _5264_;
  wire _5265_;
  wire _5266_;
  wire _5267_;
  wire _5268_;
  wire _5269_;
  wire _5270_;
  wire _5271_;
  wire _5272_;
  wire _5273_;
  wire _5274_;
  wire _5275_;
  wire _5276_;
  wire _5277_;
  wire _5278_;
  wire _5279_;
  wire _5280_;
  wire _5281_;
  wire _5282_;
  wire _5283_;
  wire _5284_;
  wire _5285_;
  wire _5286_;
  wire _5287_;
  wire _5288_;
  wire _5289_;
  wire _5290_;
  wire _5291_;
  wire _5292_;
  wire _5293_;
  wire _5294_;
  wire _5295_;
  wire _5296_;
  wire _5297_;
  wire _5298_;
  wire _5299_;
  wire _5300_;
  wire _5301_;
  wire _5302_;
  wire _5303_;
  wire _5304_;
  wire _5305_;
  wire _5306_;
  wire _5307_;
  wire _5308_;
  wire _5309_;
  wire _5310_;
  wire _5311_;
  wire _5312_;
  wire _5313_;
  wire _5314_;
  wire _5315_;
  wire _5316_;
  wire _5317_;
  wire _5318_;
  wire _5319_;
  wire _5320_;
  wire _5321_;
  wire _5322_;
  wire _5323_;
  wire _5324_;
  wire _5325_;
  wire _5326_;
  wire _5327_;
  wire _5328_;
  wire _5329_;
  wire _5330_;
  wire _5331_;
  wire _5332_;
  wire _5333_;
  wire _5334_;
  wire _5335_;
  wire _5336_;
  wire _5337_;
  wire _5338_;
  wire _5339_;
  wire _5340_;
  wire _5341_;
  wire _5342_;
  wire _5343_;
  wire _5344_;
  wire _5345_;
  wire _5346_;
  wire _5347_;
  wire _5348_;
  wire _5349_;
  wire _5350_;
  wire _5351_;
  wire _5352_;
  wire _5353_;
  wire _5354_;
  wire _5355_;
  wire _5356_;
  wire _5357_;
  wire _5358_;
  wire _5359_;
  wire _5360_;
  wire _5361_;
  wire _5362_;
  wire _5363_;
  wire _5364_;
  wire _5365_;
  wire _5366_;
  wire _5367_;
  wire _5368_;
  wire _5369_;
  wire _5370_;
  wire _5371_;
  wire _5372_;
  wire _5373_;
  wire _5374_;
  wire _5375_;
  wire _5376_;
  wire _5377_;
  wire _5378_;
  wire _5379_;
  wire _5380_;
  wire _5381_;
  wire _5382_;
  wire _5383_;
  wire _5384_;
  wire _5385_;
  wire _5386_;
  wire _5387_;
  wire _5388_;
  wire _5389_;
  wire _5390_;
  wire _5391_;
  wire _5392_;
  wire _5393_;
  wire _5394_;
  wire _5395_;
  wire _5396_;
  wire _5397_;
  wire _5398_;
  wire _5399_;
  wire _5400_;
  wire _5401_;
  wire _5402_;
  wire _5403_;
  wire _5404_;
  wire _5405_;
  wire _5406_;
  wire _5407_;
  wire _5408_;
  wire _5409_;
  wire _5410_;
  wire _5411_;
  wire _5412_;
  wire _5413_;
  wire _5414_;
  wire _5415_;
  wire _5416_;
  wire _5417_;
  wire _5418_;
  wire _5419_;
  wire _5420_;
  wire _5421_;
  wire _5422_;
  wire _5423_;
  wire _5424_;
  wire _5425_;
  wire _5426_;
  wire _5427_;
  wire _5428_;
  wire _5429_;
  wire _5430_;
  wire _5431_;
  wire _5432_;
  wire _5433_;
  wire _5434_;
  wire _5435_;
  wire _5436_;
  wire _5437_;
  wire _5438_;
  wire _5439_;
  wire _5440_;
  wire _5441_;
  wire _5442_;
  wire _5443_;
  wire _5444_;
  wire _5445_;
  wire _5446_;
  wire _5447_;
  wire _5448_;
  wire _5449_;
  wire _5450_;
  wire _5451_;
  wire _5452_;
  wire _5453_;
  wire _5454_;
  wire _5455_;
  wire _5456_;
  wire _5457_;
  wire _5458_;
  wire _5459_;
  wire _5460_;
  wire _5461_;
  wire _5462_;
  wire _5463_;
  wire _5464_;
  wire _5465_;
  wire _5466_;
  wire _5467_;
  wire _5468_;
  wire _5469_;
  wire _5470_;
  wire _5471_;
  wire _5472_;
  wire _5473_;
  wire _5474_;
  wire _5475_;
  wire _5476_;
  wire _5477_;
  wire _5478_;
  wire _5479_;
  wire _5480_;
  wire _5481_;
  wire _5482_;
  wire _5483_;
  wire _5484_;
  wire _5485_;
  wire _5486_;
  wire _5487_;
  wire _5488_;
  wire _5489_;
  wire _5490_;
  wire _5491_;
  wire _5492_;
  wire _5493_;
  wire _5494_;
  wire _5495_;
  wire _5496_;
  wire _5497_;
  wire _5498_;
  wire _5499_;
  wire _5500_;
  wire _5501_;
  wire _5502_;
  wire _5503_;
  wire _5504_;
  wire _5505_;
  wire _5506_;
  wire _5507_;
  wire _5508_;
  wire _5509_;
  wire _5510_;
  wire _5511_;
  wire _5512_;
  wire _5513_;
  wire _5514_;
  wire _5515_;
  wire _5516_;
  wire _5517_;
  wire _5518_;
  wire _5519_;
  wire _5520_;
  wire _5521_;
  wire _5522_;
  wire _5523_;
  wire _5524_;
  wire _5525_;
  wire _5526_;
  wire _5527_;
  wire _5528_;
  wire _5529_;
  wire _5530_;
  wire _5531_;
  wire _5532_;
  wire _5533_;
  wire _5534_;
  wire _5535_;
  wire _5536_;
  wire _5537_;
  wire _5538_;
  wire _5539_;
  wire _5540_;
  wire _5541_;
  wire _5542_;
  wire _5543_;
  wire _5544_;
  wire _5545_;
  wire _5546_;
  wire _5547_;
  wire _5548_;
  wire _5549_;
  wire _5550_;
  wire _5551_;
  wire _5552_;
  wire _5553_;
  wire _5554_;
  wire _5555_;
  wire _5556_;
  wire _5557_;
  wire _5558_;
  wire _5559_;
  wire _5560_;
  wire _5561_;
  wire _5562_;
  wire _5563_;
  wire _5564_;
  wire _5565_;
  wire _5566_;
  wire _5567_;
  wire _5568_;
  wire _5569_;
  wire _5570_;
  wire _5571_;
  wire _5572_;
  wire _5573_;
  wire _5574_;
  wire _5575_;
  wire _5576_;
  wire _5577_;
  wire _5578_;
  wire _5579_;
  wire _5580_;
  wire _5581_;
  wire _5582_;
  wire _5583_;
  wire _5584_;
  wire _5585_;
  wire _5586_;
  wire _5587_;
  wire _5588_;
  wire _5589_;
  wire _5590_;
  wire _5591_;
  wire _5592_;
  wire _5593_;
  wire _5594_;
  wire _5595_;
  wire _5596_;
  wire _5597_;
  wire _5598_;
  wire _5599_;
  wire _5600_;
  wire _5601_;
  wire _5602_;
  wire _5603_;
  wire _5604_;
  wire _5605_;
  wire _5606_;
  wire _5607_;
  wire _5608_;
  wire _5609_;
  wire _5610_;
  wire _5611_;
  wire _5612_;
  wire _5613_;
  wire _5614_;
  wire _5615_;
  wire _5616_;
  wire _5617_;
  wire _5618_;
  wire _5619_;
  wire _5620_;
  wire _5621_;
  wire _5622_;
  wire _5623_;
  wire _5624_;
  wire _5625_;
  wire _5626_;
  wire _5627_;
  wire _5628_;
  wire _5629_;
  wire _5630_;
  wire _5631_;
  wire _5632_;
  wire _5633_;
  wire _5634_;
  wire _5635_;
  wire _5636_;
  wire _5637_;
  wire _5638_;
  wire _5639_;
  wire _5640_;
  wire _5641_;
  wire _5642_;
  wire _5643_;
  wire _5644_;
  wire _5645_;
  wire _5646_;
  wire _5647_;
  wire _5648_;
  wire _5649_;
  wire _5650_;
  wire _5651_;
  wire _5652_;
  wire _5653_;
  wire _5654_;
  wire _5655_;
  wire _5656_;
  wire _5657_;
  wire _5658_;
  wire _5659_;
  wire _5660_;
  wire _5661_;
  wire _5662_;
  wire _5663_;
  wire _5664_;
  wire _5665_;
  wire _5666_;
  wire _5667_;
  wire _5668_;
  wire _5669_;
  wire _5670_;
  wire _5671_;
  wire _5672_;
  wire _5673_;
  wire _5674_;
  wire _5675_;
  wire _5676_;
  wire _5677_;
  wire _5678_;
  wire _5679_;
  wire _5680_;
  wire _5681_;
  wire _5682_;
  wire _5683_;
  wire _5684_;
  wire _5685_;
  wire _5686_;
  wire _5687_;
  wire _5688_;
  wire _5689_;
  wire _5690_;
  wire _5691_;
  wire _5692_;
  wire _5693_;
  wire _5694_;
  wire _5695_;
  wire _5696_;
  wire _5697_;
  wire _5698_;
  wire _5699_;
  wire _5700_;
  wire _5701_;
  wire _5702_;
  wire _5703_;
  wire _5704_;
  wire _5705_;
  wire _5706_;
  wire _5707_;
  wire _5708_;
  wire _5709_;
  wire _5710_;
  wire _5711_;
  wire _5712_;
  wire _5713_;
  wire _5714_;
  wire _5715_;
  wire _5716_;
  wire _5717_;
  wire _5718_;
  wire _5719_;
  wire _5720_;
  wire _5721_;
  wire _5722_;
  wire _5723_;
  wire _5724_;
  wire _5725_;
  wire _5726_;
  wire _5727_;
  wire _5728_;
  wire _5729_;
  wire _5730_;
  wire _5731_;
  wire _5732_;
  wire _5733_;
  wire _5734_;
  wire _5735_;
  wire _5736_;
  wire _5737_;
  wire _5738_;
  wire _5739_;
  wire _5740_;
  wire _5741_;
  wire _5742_;
  wire _5743_;
  wire _5744_;
  wire _5745_;
  wire _5746_;
  wire _5747_;
  wire _5748_;
  wire _5749_;
  wire _5750_;
  wire _5751_;
  wire _5752_;
  wire _5753_;
  wire _5754_;
  wire _5755_;
  wire _5756_;
  wire _5757_;
  wire _5758_;
  wire _5759_;
  wire _5760_;
  wire _5761_;
  wire _5762_;
  wire _5763_;
  wire _5764_;
  wire _5765_;
  wire _5766_;
  wire _5767_;
  wire _5768_;
  wire _5769_;
  wire _5770_;
  wire _5771_;
  wire _5772_;
  wire _5773_;
  wire _5774_;
  wire _5775_;
  wire _5776_;
  wire _5777_;
  wire _5778_;
  wire _5779_;
  wire _5780_;
  wire _5781_;
  wire _5782_;
  wire _5783_;
  wire _5784_;
  wire _5785_;
  wire _5786_;
  wire _5787_;
  wire _5788_;
  wire _5789_;
  wire _5790_;
  wire _5791_;
  wire _5792_;
  wire _5793_;
  wire _5794_;
  wire _5795_;
  wire _5796_;
  wire _5797_;
  wire _5798_;
  wire _5799_;
  wire _5800_;
  wire _5801_;
  wire _5802_;
  wire _5803_;
  wire _5804_;
  wire _5805_;
  wire _5806_;
  wire _5807_;
  wire _5808_;
  wire _5809_;
  wire _5810_;
  wire _5811_;
  wire _5812_;
  wire _5813_;
  wire _5814_;
  wire _5815_;
  wire _5816_;
  wire _5817_;
  wire _5818_;
  wire _5819_;
  wire _5820_;
  wire _5821_;
  wire _5822_;
  wire _5823_;
  wire _5824_;
  wire _5825_;
  wire _5826_;
  wire _5827_;
  wire _5828_;
  wire _5829_;
  wire _5830_;
  wire _5831_;
  wire _5832_;
  wire _5833_;
  wire _5834_;
  wire _5835_;
  wire _5836_;
  wire _5837_;
  wire _5838_;
  wire _5839_;
  wire _5840_;
  wire _5841_;
  wire _5842_;
  wire _5843_;
  wire _5844_;
  wire _5845_;
  wire _5846_;
  wire _5847_;
  wire _5848_;
  wire _5849_;
  wire _5850_;
  wire _5851_;
  wire _5852_;
  wire _5853_;
  wire _5854_;
  wire _5855_;
  wire _5856_;
  wire _5857_;
  wire _5858_;
  wire _5859_;
  wire _5860_;
  wire _5861_;
  wire _5862_;
  wire _5863_;
  wire _5864_;
  wire _5865_;
  wire _5866_;
  wire _5867_;
  wire _5868_;
  wire _5869_;
  wire _5870_;
  wire _5871_;
  wire _5872_;
  wire _5873_;
  wire _5874_;
  wire _5875_;
  wire _5876_;
  wire _5877_;
  wire _5878_;
  wire _5879_;
  wire _5880_;
  wire _5881_;
  wire _5882_;
  wire _5883_;
  wire _5884_;
  wire _5885_;
  wire _5886_;
  wire _5887_;
  wire _5888_;
  wire _5889_;
  wire _5890_;
  wire _5891_;
  wire _5892_;
  wire _5893_;
  wire _5894_;
  wire _5895_;
  wire _5896_;
  wire _5897_;
  wire _5898_;
  wire _5899_;
  wire _5900_;
  wire _5901_;
  wire _5902_;
  wire _5903_;
  wire _5904_;
  wire _5905_;
  wire _5906_;
  wire _5907_;
  wire _5908_;
  wire _5909_;
  wire _5910_;
  wire _5911_;
  wire _5912_;
  wire _5913_;
  wire _5914_;
  wire _5915_;
  wire _5916_;
  wire _5917_;
  wire _5918_;
  wire _5919_;
  wire _5920_;
  wire _5921_;
  wire _5922_;
  wire _5923_;
  wire _5924_;
  wire _5925_;
  wire _5926_;
  wire _5927_;
  wire _5928_;
  wire _5929_;
  wire _5930_;
  wire _5931_;
  wire _5932_;
  wire _5933_;
  wire _5934_;
  wire _5935_;
  wire _5936_;
  wire _5937_;
  wire _5938_;
  wire _5939_;
  wire _5940_;
  wire _5941_;
  wire _5942_;
  wire _5943_;
  wire _5944_;
  wire _5945_;
  wire _5946_;
  wire _5947_;
  wire _5948_;
  wire _5949_;
  wire _5950_;
  wire _5951_;
  wire _5952_;
  wire _5953_;
  wire _5954_;
  wire _5955_;
  wire _5956_;
  wire _5957_;
  wire _5958_;
  wire _5959_;
  wire _5960_;
  wire _5961_;
  wire _5962_;
  wire _5963_;
  wire _5964_;
  wire _5965_;
  wire _5966_;
  wire _5967_;
  wire _5968_;
  wire _5969_;
  wire _5970_;
  wire _5971_;
  wire _5972_;
  wire _5973_;
  wire _5974_;
  wire _5975_;
  wire _5976_;
  wire _5977_;
  wire _5978_;
  wire _5979_;
  wire _5980_;
  wire _5981_;
  wire _5982_;
  wire _5983_;
  wire _5984_;
  wire _5985_;
  wire _5986_;
  wire _5987_;
  wire _5988_;
  wire _5989_;
  wire _5990_;
  wire _5991_;
  wire _5992_;
  wire _5993_;
  wire _5994_;
  wire _5995_;
  wire _5996_;
  wire _5997_;
  wire _5998_;
  wire _5999_;
  wire _6000_;
  wire _6001_;
  wire _6002_;
  wire _6003_;
  wire _6004_;
  wire _6005_;
  wire _6006_;
  wire _6007_;
  wire _6008_;
  wire _6009_;
  wire _6010_;
  wire _6011_;
  wire _6012_;
  wire _6013_;
  wire _6014_;
  wire _6015_;
  wire _6016_;
  wire _6017_;
  wire _6018_;
  wire _6019_;
  wire _6020_;
  wire _6021_;
  wire _6022_;
  wire _6023_;
  wire _6024_;
  wire _6025_;
  wire _6026_;
  wire _6027_;
  wire _6028_;
  wire _6029_;
  wire _6030_;
  wire _6031_;
  wire _6032_;
  wire _6033_;
  wire _6034_;
  wire _6035_;
  wire _6036_;
  wire _6037_;
  wire _6038_;
  wire _6039_;
  wire _6040_;
  wire _6041_;
  wire _6042_;
  wire _6043_;
  wire _6044_;
  wire _6045_;
  wire _6046_;
  wire _6047_;
  wire _6048_;
  wire _6049_;
  wire _6050_;
  wire _6051_;
  wire _6052_;
  wire _6053_;
  wire _6054_;
  wire _6055_;
  wire _6056_;
  wire _6057_;
  wire _6058_;
  wire _6059_;
  wire _6060_;
  wire _6061_;
  wire _6062_;
  wire _6063_;
  wire _6064_;
  wire _6065_;
  wire _6066_;
  wire _6067_;
  wire _6068_;
  wire _6069_;
  wire _6070_;
  wire _6071_;
  wire _6072_;
  wire _6073_;
  wire _6074_;
  wire _6075_;
  wire _6076_;
  wire _6077_;
  wire _6078_;
  wire _6079_;
  wire _6080_;
  wire _6081_;
  wire _6082_;
  wire _6083_;
  wire _6084_;
  wire _6085_;
  wire _6086_;
  wire _6087_;
  wire _6088_;
  wire _6089_;
  wire _6090_;
  wire _6091_;
  wire _6092_;
  wire _6093_;
  wire _6094_;
  wire _6095_;
  wire _6096_;
  wire _6097_;
  wire _6098_;
  wire _6099_;
  wire _6100_;
  wire _6101_;
  wire _6102_;
  wire _6103_;
  wire _6104_;
  wire _6105_;
  wire _6106_;
  wire _6107_;
  wire _6108_;
  wire _6109_;
  wire _6110_;
  wire _6111_;
  wire _6112_;
  wire _6113_;
  wire _6114_;
  wire _6115_;
  wire _6116_;
  wire _6117_;
  wire _6118_;
  wire _6119_;
  wire _6120_;
  wire _6121_;
  wire _6122_;
  wire _6123_;
  wire _6124_;
  wire _6125_;
  wire _6126_;
  wire _6127_;
  wire _6128_;
  wire _6129_;
  wire _6130_;
  wire _6131_;
  wire _6132_;
  wire _6133_;
  wire _6134_;
  wire _6135_;
  wire _6136_;
  wire _6137_;
  wire _6138_;
  wire _6139_;
  wire _6140_;
  wire _6141_;
  wire _6142_;
  wire _6143_;
  wire _6144_;
  wire _6145_;
  wire _6146_;
  wire _6147_;
  wire _6148_;
  wire _6149_;
  wire _6150_;
  wire _6151_;
  wire _6152_;
  wire _6153_;
  wire _6154_;
  wire _6155_;
  wire _6156_;
  wire _6157_;
  wire _6158_;
  wire _6159_;
  wire _6160_;
  wire _6161_;
  wire _6162_;
  wire _6163_;
  wire _6164_;
  wire _6165_;
  wire _6166_;
  wire _6167_;
  wire _6168_;
  wire _6169_;
  wire _6170_;
  wire _6171_;
  wire _6172_;
  wire _6173_;
  wire _6174_;
  wire _6175_;
  wire _6176_;
  wire _6177_;
  wire _6178_;
  wire _6179_;
  wire _6180_;
  wire _6181_;
  wire _6182_;
  wire _6183_;
  wire _6184_;
  wire _6185_;
  wire _6186_;
  wire _6187_;
  wire _6188_;
  wire _6189_;
  wire _6190_;
  wire _6191_;
  wire _6192_;
  wire _6193_;
  wire _6194_;
  wire _6195_;
  wire _6196_;
  wire _6197_;
  wire _6198_;
  wire _6199_;
  wire _6200_;
  wire _6201_;
  wire _6202_;
  wire _6203_;
  wire _6204_;
  wire _6205_;
  wire _6206_;
  wire _6207_;
  wire _6208_;
  wire _6209_;
  wire _6210_;
  wire _6211_;
  wire _6212_;
  wire _6213_;
  wire _6214_;
  wire _6215_;
  wire _6216_;
  wire _6217_;
  wire _6218_;
  wire _6219_;
  wire _6220_;
  wire _6221_;
  wire _6222_;
  wire _6223_;
  wire _6224_;
  wire _6225_;
  wire _6226_;
  wire _6227_;
  wire _6228_;
  wire _6229_;
  wire _6230_;
  wire _6231_;
  wire _6232_;
  wire _6233_;
  wire _6234_;
  wire _6235_;
  wire _6236_;
  wire _6237_;
  wire _6238_;
  wire _6239_;
  wire _6240_;
  wire _6241_;
  wire _6242_;
  wire _6243_;
  wire _6244_;
  wire _6245_;
  wire _6246_;
  wire _6247_;
  wire _6248_;
  wire _6249_;
  wire _6250_;
  wire _6251_;
  wire _6252_;
  wire _6253_;
  wire _6254_;
  wire _6255_;
  wire _6256_;
  wire _6257_;
  wire _6258_;
  wire _6259_;
  wire _6260_;
  wire _6261_;
  wire _6262_;
  wire _6263_;
  wire _6264_;
  wire _6265_;
  wire _6266_;
  wire _6267_;
  wire _6268_;
  wire _6269_;
  wire _6270_;
  wire _6271_;
  wire _6272_;
  wire _6273_;
  wire _6274_;
  wire _6275_;
  wire _6276_;
  wire _6277_;
  wire _6278_;
  wire _6279_;
  wire _6280_;
  wire _6281_;
  wire _6282_;
  wire _6283_;
  wire _6284_;
  wire _6285_;
  wire _6286_;
  wire _6287_;
  wire _6288_;
  wire _6289_;
  wire _6290_;
  wire _6291_;
  wire _6292_;
  wire _6293_;
  wire _6294_;
  wire _6295_;
  wire _6296_;
  wire _6297_;
  wire _6298_;
  wire _6299_;
  wire _6300_;
  wire _6301_;
  wire _6302_;
  wire _6303_;
  wire _6304_;
  wire _6305_;
  wire _6306_;
  wire _6307_;
  wire _6308_;
  wire _6309_;
  wire _6310_;
  wire _6311_;
  wire _6312_;
  wire _6313_;
  wire _6314_;
  wire _6315_;
  wire _6316_;
  wire _6317_;
  wire _6318_;
  wire _6319_;
  wire _6320_;
  wire _6321_;
  wire _6322_;
  wire _6323_;
  wire _6324_;
  wire _6325_;
  wire _6326_;
  wire _6327_;
  wire _6328_;
  wire _6329_;
  wire _6330_;
  wire _6331_;
  wire _6332_;
  wire _6333_;
  wire _6334_;
  wire _6335_;
  wire _6336_;
  wire _6337_;
  wire _6338_;
  wire _6339_;
  wire _6340_;
  wire _6341_;
  wire _6342_;
  wire _6343_;
  wire _6344_;
  wire _6345_;
  wire _6346_;
  wire _6347_;
  wire _6348_;
  wire _6349_;
  wire _6350_;
  wire _6351_;
  wire _6352_;
  wire _6353_;
  wire _6354_;
  wire _6355_;
  wire _6356_;
  wire _6357_;
  wire _6358_;
  wire _6359_;
  wire _6360_;
  wire _6361_;
  wire _6362_;
  wire _6363_;
  wire _6364_;
  wire _6365_;
  wire _6366_;
  wire _6367_;
  wire _6368_;
  wire _6369_;
  wire _6370_;
  wire _6371_;
  wire _6372_;
  wire _6373_;
  wire _6374_;
  wire _6375_;
  wire _6376_;
  wire _6377_;
  wire _6378_;
  wire _6379_;
  wire _6380_;
  wire _6381_;
  wire _6382_;
  wire _6383_;
  wire _6384_;
  wire _6385_;
  wire _6386_;
  wire _6387_;
  wire _6388_;
  wire _6389_;
  wire _6390_;
  wire _6391_;
  wire _6392_;
  wire _6393_;
  wire _6394_;
  wire _6395_;
  wire _6396_;
  wire _6397_;
  wire _6398_;
  wire _6399_;
  wire _6400_;
  wire _6401_;
  wire _6402_;
  wire _6403_;
  wire _6404_;
  wire _6405_;
  wire _6406_;
  wire _6407_;
  wire _6408_;
  wire _6409_;
  wire _6410_;
  wire _6411_;
  wire _6412_;
  wire _6413_;
  wire _6414_;
  wire _6415_;
  wire _6416_;
  wire _6417_;
  wire _6418_;
  wire _6419_;
  wire _6420_;
  wire _6421_;
  wire _6422_;
  wire _6423_;
  wire _6424_;
  wire _6425_;
  wire _6426_;
  wire _6427_;
  wire _6428_;
  wire _6429_;
  wire _6430_;
  wire _6431_;
  wire _6432_;
  wire _6433_;
  wire _6434_;
  wire _6435_;
  wire _6436_;
  wire _6437_;
  wire _6438_;
  wire _6439_;
  wire _6440_;
  wire _6441_;
  wire _6442_;
  wire _6443_;
  wire _6444_;
  wire _6445_;
  wire _6446_;
  wire _6447_;
  wire _6448_;
  wire _6449_;
  wire _6450_;
  wire _6451_;
  wire _6452_;
  wire _6453_;
  wire _6454_;
  wire _6455_;
  wire _6456_;
  wire _6457_;
  wire _6458_;
  wire _6459_;
  wire _6460_;
  wire _6461_;
  wire _6462_;
  wire _6463_;
  wire _6464_;
  wire _6465_;
  wire _6466_;
  wire _6467_;
  wire _6468_;
  wire _6469_;
  wire _6470_;
  wire _6471_;
  wire _6472_;
  wire _6473_;
  wire _6474_;
  wire _6475_;
  wire _6476_;
  wire _6477_;
  wire _6478_;
  wire _6479_;
  wire _6480_;
  wire _6481_;
  wire _6482_;
  wire _6483_;
  wire _6484_;
  wire _6485_;
  wire _6486_;
  wire _6487_;
  wire _6488_;
  wire _6489_;
  wire _6490_;
  wire _6491_;
  wire _6492_;
  wire _6493_;
  wire _6494_;
  wire _6495_;
  wire _6496_;
  wire _6497_;
  wire _6498_;
  wire _6499_;
  wire _6500_;
  wire _6501_;
  wire _6502_;
  wire _6503_;
  wire _6504_;
  wire _6505_;
  wire _6506_;
  wire _6507_;
  wire _6508_;
  wire _6509_;
  wire _6510_;
  wire _6511_;
  wire _6512_;
  wire _6513_;
  wire _6514_;
  wire _6515_;
  wire _6516_;
  wire _6517_;
  wire _6518_;
  wire _6519_;
  wire _6520_;
  wire _6521_;
  wire _6522_;
  wire _6523_;
  wire _6524_;
  wire _6525_;
  wire _6526_;
  wire _6527_;
  wire _6528_;
  wire _6529_;
  wire _6530_;
  wire _6531_;
  wire _6532_;
  wire _6533_;
  wire _6534_;
  wire _6535_;
  wire _6536_;
  wire _6537_;
  wire _6538_;
  wire _6539_;
  wire _6540_;
  wire _6541_;
  wire _6542_;
  wire _6543_;
  wire _6544_;
  wire _6545_;
  wire _6546_;
  wire _6547_;
  wire _6548_;
  wire _6549_;
  wire _6550_;
  wire _6551_;
  wire _6552_;
  wire _6553_;
  wire _6554_;
  wire _6555_;
  wire _6556_;
  wire _6557_;
  wire _6558_;
  wire _6559_;
  wire _6560_;
  wire _6561_;
  wire _6562_;
  wire _6563_;
  wire _6564_;
  wire _6565_;
  wire _6566_;
  wire _6567_;
  wire _6568_;
  wire _6569_;
  wire _6570_;
  wire _6571_;
  wire _6572_;
  wire _6573_;
  wire _6574_;
  wire _6575_;
  wire _6576_;
  wire _6577_;
  wire _6578_;
  wire _6579_;
  wire _6580_;
  wire _6581_;
  wire _6582_;
  wire _6583_;
  wire _6584_;
  wire _6585_;
  wire _6586_;
  wire _6587_;
  wire _6588_;
  wire _6589_;
  wire _6590_;
  wire _6591_;
  wire _6592_;
  wire _6593_;
  wire _6594_;
  wire _6595_;
  wire _6596_;
  wire _6597_;
  wire _6598_;
  wire _6599_;
  wire _6600_;
  wire _6601_;
  wire _6602_;
  wire _6603_;
  wire _6604_;
  wire _6605_;
  wire _6606_;
  wire _6607_;
  wire _6608_;
  wire _6609_;
  wire _6610_;
  wire _6611_;
  wire _6612_;
  wire _6613_;
  wire _6614_;
  wire _6615_;
  wire _6616_;
  wire _6617_;
  wire _6618_;
  wire _6619_;
  wire _6620_;
  wire _6621_;
  wire _6622_;
  wire _6623_;
  wire _6624_;
  wire _6625_;
  wire _6626_;
  wire _6627_;
  wire _6628_;
  wire _6629_;
  wire _6630_;
  wire _6631_;
  wire _6632_;
  wire _6633_;
  wire _6634_;
  wire _6635_;
  wire _6636_;
  wire _6637_;
  wire _6638_;
  wire _6639_;
  wire _6640_;
  wire _6641_;
  wire _6642_;
  wire _6643_;
  wire _6644_;
  wire _6645_;
  wire _6646_;
  wire _6647_;
  wire _6648_;
  wire _6649_;
  wire _6650_;
  wire _6651_;
  wire _6652_;
  wire _6653_;
  wire _6654_;
  wire _6655_;
  wire _6656_;
  wire _6657_;
  wire _6658_;
  wire _6659_;
  wire _6660_;
  wire _6661_;
  wire _6662_;
  wire _6663_;
  wire _6664_;
  wire _6665_;
  wire _6666_;
  wire _6667_;
  wire _6668_;
  wire _6669_;
  wire _6670_;
  wire _6671_;
  wire _6672_;
  wire _6673_;
  wire _6674_;
  wire _6675_;
  wire _6676_;
  wire _6677_;
  wire _6678_;
  wire _6679_;
  wire _6680_;
  wire _6681_;
  wire _6682_;
  wire _6683_;
  wire _6684_;
  wire _6685_;
  wire _6686_;
  wire _6687_;
  wire _6688_;
  wire _6689_;
  wire _6690_;
  wire _6691_;
  wire _6692_;
  wire _6693_;
  wire _6694_;
  wire _6695_;
  wire _6696_;
  wire _6697_;
  wire _6698_;
  wire _6699_;
  wire _6700_;
  wire _6701_;
  wire _6702_;
  wire _6703_;
  wire _6704_;
  wire _6705_;
  wire _6706_;
  wire _6707_;
  wire _6708_;
  wire _6709_;
  wire _6710_;
  wire _6711_;
  wire _6712_;
  wire _6713_;
  wire _6714_;
  wire _6715_;
  wire _6716_;
  wire _6717_;
  wire _6718_;
  wire _6719_;
  wire _6720_;
  wire _6721_;
  wire _6722_;
  wire _6723_;
  wire _6724_;
  wire _6725_;
  wire _6726_;
  wire _6727_;
  wire _6728_;
  wire _6729_;
  wire _6730_;
  wire _6731_;
  wire _6732_;
  wire _6733_;
  wire _6734_;
  wire _6735_;
  wire _6736_;
  wire _6737_;
  wire _6738_;
  wire _6739_;
  wire _6740_;
  wire _6741_;
  wire _6742_;
  wire _6743_;
  wire _6744_;
  wire _6745_;
  wire _6746_;
  wire _6747_;
  wire _6748_;
  wire _6749_;
  wire _6750_;
  wire _6751_;
  wire _6752_;
  wire _6753_;
  wire _6754_;
  wire _6755_;
  wire _6756_;
  wire _6757_;
  wire _6758_;
  wire _6759_;
  wire _6760_;
  wire _6761_;
  wire _6762_;
  wire _6763_;
  wire _6764_;
  wire _6765_;
  wire _6766_;
  wire _6767_;
  wire _6768_;
  wire _6769_;
  wire _6770_;
  wire _6771_;
  wire _6772_;
  wire _6773_;
  wire _6774_;
  wire _6775_;
  wire _6776_;
  wire _6777_;
  wire _6778_;
  wire _6779_;
  wire _6780_;
  wire _6781_;
  wire _6782_;
  wire _6783_;
  wire _6784_;
  wire _6785_;
  wire _6786_;
  wire _6787_;
  wire _6788_;
  wire _6789_;
  wire _6790_;
  wire _6791_;
  wire _6792_;
  wire _6793_;
  wire _6794_;
  wire _6795_;
  wire _6796_;
  wire _6797_;
  wire _6798_;
  wire _6799_;
  wire _6800_;
  wire _6801_;
  wire _6802_;
  wire _6803_;
  wire _6804_;
  wire _6805_;
  wire _6806_;
  wire _6807_;
  wire _6808_;
  wire _6809_;
  wire _6810_;
  wire _6811_;
  wire _6812_;
  wire _6813_;
  wire _6814_;
  wire _6815_;
  wire _6816_;
  wire _6817_;
  wire _6818_;
  wire _6819_;
  wire _6820_;
  wire _6821_;
  wire _6822_;
  wire _6823_;
  wire _6824_;
  wire _6825_;
  wire _6826_;
  wire _6827_;
  wire _6828_;
  wire _6829_;
  wire _6830_;
  wire _6831_;
  wire _6832_;
  wire _6833_;
  wire _6834_;
  wire _6835_;
  wire _6836_;
  wire _6837_;
  wire _6838_;
  wire _6839_;
  wire _6840_;
  wire _6841_;
  wire _6842_;
  wire _6843_;
  wire _6844_;
  wire _6845_;
  wire _6846_;
  wire _6847_;
  wire _6848_;
  wire _6849_;
  wire _6850_;
  wire _6851_;
  wire _6852_;
  wire _6853_;
  wire _6854_;
  wire _6855_;
  wire _6856_;
  wire _6857_;
  wire _6858_;
  wire _6859_;
  wire _6860_;
  wire _6861_;
  wire _6862_;
  wire _6863_;
  wire _6864_;
  wire _6865_;
  wire _6866_;
  wire _6867_;
  wire _6868_;
  wire _6869_;
  wire _6870_;
  wire _6871_;
  wire _6872_;
  wire _6873_;
  wire _6874_;
  wire _6875_;
  wire _6876_;
  wire _6877_;
  wire _6878_;
  wire _6879_;
  wire _6880_;
  wire _6881_;
  wire _6882_;
  wire _6883_;
  wire _6884_;
  wire _6885_;
  wire _6886_;
  wire _6887_;
  wire _6888_;
  wire _6889_;
  wire _6890_;
  wire _6891_;
  wire _6892_;
  wire _6893_;
  wire _6894_;
  wire _6895_;
  wire _6896_;
  wire _6897_;
  wire _6898_;
  wire _6899_;
  wire _6900_;
  wire _6901_;
  wire _6902_;
  wire _6903_;
  wire _6904_;
  wire _6905_;
  wire _6906_;
  wire _6907_;
  wire _6908_;
  wire _6909_;
  wire _6910_;
  wire _6911_;
  wire _6912_;
  wire _6913_;
  wire _6914_;
  wire _6915_;
  wire _6916_;
  wire _6917_;
  wire _6918_;
  wire _6919_;
  wire _6920_;
  wire _6921_;
  wire _6922_;
  wire _6923_;
  wire _6924_;
  wire _6925_;
  wire _6926_;
  wire _6927_;
  wire _6928_;
  wire _6929_;
  wire _6930_;
  wire _6931_;
  wire _6932_;
  wire _6933_;
  wire _6934_;
  wire _6935_;
  wire _6936_;
  wire _6937_;
  wire _6938_;
  wire _6939_;
  wire _6940_;
  wire _6941_;
  wire _6942_;
  wire _6943_;
  wire _6944_;
  wire _6945_;
  wire _6946_;
  wire _6947_;
  wire _6948_;
  wire _6949_;
  wire _6950_;
  wire _6951_;
  wire _6952_;
  wire _6953_;
  wire _6954_;
  wire _6955_;
  wire _6956_;
  wire _6957_;
  wire _6958_;
  wire _6959_;
  wire _6960_;
  wire _6961_;
  wire _6962_;
  wire _6963_;
  wire _6964_;
  wire _6965_;
  wire _6966_;
  wire _6967_;
  wire _6968_;
  wire _6969_;
  wire _6970_;
  wire _6971_;
  wire _6972_;
  wire _6973_;
  wire _6974_;
  wire _6975_;
  wire _6976_;
  wire _6977_;
  wire _6978_;
  wire _6979_;
  wire _6980_;
  wire _6981_;
  wire _6982_;
  wire _6983_;
  wire _6984_;
  wire _6985_;
  wire _6986_;
  wire _6987_;
  wire _6988_;
  wire _6989_;
  wire _6990_;
  wire _6991_;
  wire _6992_;
  wire _6993_;
  wire _6994_;
  wire _6995_;
  wire _6996_;
  wire _6997_;
  wire _6998_;
  wire _6999_;
  wire _7000_;
  wire _7001_;
  wire _7002_;
  wire _7003_;
  wire _7004_;
  wire _7005_;
  wire _7006_;
  wire _7007_;
  wire _7008_;
  wire _7009_;
  wire _7010_;
  wire _7011_;
  wire _7012_;
  wire _7013_;
  wire _7014_;
  wire _7015_;
  wire _7016_;
  wire _7017_;
  wire _7018_;
  wire _7019_;
  wire _7020_;
  wire _7021_;
  wire _7022_;
  wire _7023_;
  wire _7024_;
  wire _7025_;
  wire _7026_;
  wire _7027_;
  wire _7028_;
  wire _7029_;
  wire _7030_;
  wire _7031_;
  wire _7032_;
  wire _7033_;
  wire _7034_;
  wire _7035_;
  wire _7036_;
  wire _7037_;
  wire _7038_;
  wire _7039_;
  wire _7040_;
  wire _7041_;
  wire _7042_;
  wire _7043_;
  wire _7044_;
  wire _7045_;
  wire _7046_;
  wire _7047_;
  wire _7048_;
  wire _7049_;
  wire _7050_;
  wire _7051_;
  wire _7052_;
  wire _7053_;
  wire _7054_;
  wire _7055_;
  wire _7056_;
  wire _7057_;
  wire _7058_;
  wire _7059_;
  wire _7060_;
  wire _7061_;
  wire _7062_;
  wire _7063_;
  wire _7064_;
  wire _7065_;
  wire _7066_;
  wire _7067_;
  wire _7068_;
  wire _7069_;
  wire _7070_;
  wire _7071_;
  wire _7072_;
  wire _7073_;
  wire _7074_;
  wire _7075_;
  wire _7076_;
  wire _7077_;
  wire _7078_;
  wire _7079_;
  wire _7080_;
  wire _7081_;
  wire _7082_;
  wire _7083_;
  wire _7084_;
  wire _7085_;
  wire _7086_;
  wire _7087_;
  wire _7088_;
  wire _7089_;
  wire _7090_;
  wire _7091_;
  wire _7092_;
  wire _7093_;
  wire _7094_;
  wire _7095_;
  wire _7096_;
  wire _7097_;
  wire _7098_;
  wire _7099_;
  wire _7100_;
  wire _7101_;
  wire _7102_;
  wire _7103_;
  wire _7104_;
  wire _7105_;
  wire _7106_;
  wire _7107_;
  wire _7108_;
  wire _7109_;
  wire _7110_;
  wire _7111_;
  wire _7112_;
  wire _7113_;
  wire _7114_;
  wire _7115_;
  wire _7116_;
  wire _7117_;
  wire _7118_;
  wire _7119_;
  wire _7120_;
  wire _7121_;
  wire _7122_;
  wire _7123_;
  wire _7124_;
  wire _7125_;
  wire _7126_;
  wire _7127_;
  wire _7128_;
  wire _7129_;
  wire _7130_;
  wire _7131_;
  wire _7132_;
  wire _7133_;
  wire _7134_;
  wire _7135_;
  wire _7136_;
  wire _7137_;
  wire _7138_;
  wire _7139_;
  wire _7140_;
  wire _7141_;
  wire _7142_;
  wire _7143_;
  wire _7144_;
  wire _7145_;
  wire _7146_;
  wire _7147_;
  wire _7148_;
  wire _7149_;
  wire _7150_;
  wire _7151_;
  wire _7152_;
  wire _7153_;
  wire _7154_;
  wire _7155_;
  wire _7156_;
  wire _7157_;
  wire _7158_;
  wire _7159_;
  wire _7160_;
  wire _7161_;
  wire _7162_;
  wire _7163_;
  wire _7164_;
  wire _7165_;
  wire _7166_;
  wire _7167_;
  wire _7168_;
  wire _7169_;
  wire _7170_;
  wire _7171_;
  wire _7172_;
  wire _7173_;
  wire _7174_;
  wire _7175_;
  wire _7176_;
  wire _7177_;
  wire _7178_;
  wire _7179_;
  wire _7180_;
  wire _7181_;
  wire _7182_;
  wire _7183_;
  wire _7184_;
  wire _7185_;
  wire _7186_;
  wire _7187_;
  wire _7188_;
  wire _7189_;
  wire _7190_;
  wire _7191_;
  wire _7192_;
  wire _7193_;
  wire _7194_;
  wire _7195_;
  wire _7196_;
  wire _7197_;
  wire _7198_;
  wire _7199_;
  wire _7200_;
  wire _7201_;
  wire _7202_;
  wire _7203_;
  wire _7204_;
  wire _7205_;
  wire _7206_;
  wire _7207_;
  wire _7208_;
  wire _7209_;
  wire _7210_;
  wire _7211_;
  wire _7212_;
  wire _7213_;
  wire _7214_;
  wire _7215_;
  wire _7216_;
  wire _7217_;
  wire _7218_;
  wire _7219_;
  wire _7220_;
  wire _7221_;
  wire _7222_;
  wire _7223_;
  wire _7224_;
  wire _7225_;
  wire _7226_;
  wire _7227_;
  wire _7228_;
  wire _7229_;
  wire _7230_;
  wire _7231_;
  wire _7232_;
  wire _7233_;
  wire _7234_;
  wire _7235_;
  wire _7236_;
  wire _7237_;
  wire _7238_;
  wire _7239_;
  wire _7240_;
  wire _7241_;
  wire _7242_;
  wire _7243_;
  wire _7244_;
  wire _7245_;
  wire _7246_;
  wire _7247_;
  wire _7248_;
  wire _7249_;
  wire _7250_;
  wire _7251_;
  wire _7252_;
  wire _7253_;
  wire _7254_;
  wire _7255_;
  wire _7256_;
  wire _7257_;
  wire _7258_;
  wire _7259_;
  wire _7260_;
  wire _7261_;
  wire _7262_;
  wire _7263_;
  wire _7264_;
  wire _7265_;
  wire _7266_;
  wire _7267_;
  wire _7268_;
  wire _7269_;
  wire _7270_;
  wire _7271_;
  wire _7272_;
  wire _7273_;
  wire _7274_;
  wire _7275_;
  wire _7276_;
  wire _7277_;
  wire _7278_;
  wire _7279_;
  wire _7280_;
  wire _7281_;
  wire _7282_;
  wire _7283_;
  wire _7284_;
  wire _7285_;
  wire _7286_;
  wire _7287_;
  wire _7288_;
  wire _7289_;
  wire _7290_;
  wire _7291_;
  wire _7292_;
  wire _7293_;
  wire _7294_;
  wire _7295_;
  wire _7296_;
  wire _7297_;
  wire _7298_;
  wire _7299_;
  wire _7300_;
  wire _7301_;
  wire _7302_;
  wire _7303_;
  wire _7304_;
  wire _7305_;
  wire _7306_;
  wire _7307_;
  wire _7308_;
  wire _7309_;
  wire _7310_;
  wire _7311_;
  wire _7312_;
  wire _7313_;
  wire _7314_;
  wire _7315_;
  wire _7316_;
  wire _7317_;
  wire _7318_;
  wire _7319_;
  wire _7320_;
  wire _7321_;
  wire _7322_;
  wire _7323_;
  wire _7324_;
  wire _7325_;
  wire _7326_;
  wire _7327_;
  wire _7328_;
  wire _7329_;
  wire _7330_;
  wire _7331_;
  wire _7332_;
  wire _7333_;
  wire _7334_;
  wire _7335_;
  wire _7336_;
  wire _7337_;
  wire _7338_;
  wire _7339_;
  wire _7340_;
  wire _7341_;
  wire _7342_;
  wire _7343_;
  wire _7344_;
  wire _7345_;
  wire _7346_;
  wire _7347_;
  wire _7348_;
  wire _7349_;
  wire _7350_;
  wire _7351_;
  wire _7352_;
  wire _7353_;
  wire _7354_;
  wire _7355_;
  wire _7356_;
  wire _7357_;
  wire _7358_;
  wire _7359_;
  wire _7360_;
  wire _7361_;
  wire _7362_;
  wire _7363_;
  wire _7364_;
  wire _7365_;
  wire _7366_;
  wire _7367_;
  wire _7368_;
  wire _7369_;
  wire _7370_;
  wire _7371_;
  wire _7372_;
  wire _7373_;
  wire _7374_;
  wire _7375_;
  wire _7376_;
  wire _7377_;
  wire _7378_;
  wire _7379_;
  wire _7380_;
  wire _7381_;
  wire _7382_;
  wire _7383_;
  wire _7384_;
  wire _7385_;
  wire _7386_;
  wire _7387_;
  wire _7388_;
  wire _7389_;
  wire _7390_;
  wire _7391_;
  wire _7392_;
  wire _7393_;
  wire _7394_;
  wire _7395_;
  wire _7396_;
  wire _7397_;
  wire _7398_;
  wire _7399_;
  wire _7400_;
  wire _7401_;
  wire _7402_;
  wire _7403_;
  wire _7404_;
  wire _7405_;
  wire _7406_;
  wire _7407_;
  wire _7408_;
  wire _7409_;
  wire _7410_;
  wire _7411_;
  wire _7412_;
  wire _7413_;
  wire _7414_;
  wire _7415_;
  wire _7416_;
  wire _7417_;
  wire _7418_;
  wire _7419_;
  wire _7420_;
  wire _7421_;
  wire _7422_;
  wire _7423_;
  wire _7424_;
  wire _7425_;
  wire _7426_;
  wire _7427_;
  wire _7428_;
  wire _7429_;
  wire _7430_;
  wire _7431_;
  wire _7432_;
  wire _7433_;
  wire _7434_;
  wire _7435_;
  wire _7436_;
  wire _7437_;
  wire _7438_;
  wire _7439_;
  wire _7440_;
  wire _7441_;
  wire _7442_;
  wire _7443_;
  wire _7444_;
  wire _7445_;
  wire _7446_;
  wire _7447_;
  wire _7448_;
  wire _7449_;
  wire _7450_;
  wire _7451_;
  wire _7452_;
  wire _7453_;
  wire _7454_;
  wire _7455_;
  wire _7456_;
  wire _7457_;
  wire _7458_;
  wire _7459_;
  wire _7460_;
  wire _7461_;
  wire _7462_;
  wire _7463_;
  wire _7464_;
  wire _7465_;
  wire _7466_;
  wire _7467_;
  wire _7468_;
  wire _7469_;
  wire _7470_;
  wire _7471_;
  wire _7472_;
  wire _7473_;
  wire _7474_;
  wire _7475_;
  wire _7476_;
  wire _7477_;
  wire _7478_;
  wire _7479_;
  wire _7480_;
  wire _7481_;
  wire _7482_;
  wire _7483_;
  wire _7484_;
  wire _7485_;
  wire _7486_;
  wire _7487_;
  wire _7488_;
  wire _7489_;
  wire _7490_;
  wire _7491_;
  wire _7492_;
  wire _7493_;
  wire _7494_;
  wire _7495_;
  wire _7496_;
  wire _7497_;
  wire _7498_;
  wire _7499_;
  wire _7500_;
  wire _7501_;
  wire _7502_;
  wire _7503_;
  wire _7504_;
  wire _7505_;
  wire _7506_;
  wire _7507_;
  wire _7508_;
  wire _7509_;
  wire _7510_;
  wire _7511_;
  wire _7512_;
  wire _7513_;
  wire _7514_;
  wire _7515_;
  wire _7516_;
  wire _7517_;
  wire _7518_;
  wire _7519_;
  wire _7520_;
  wire _7521_;
  wire _7522_;
  wire _7523_;
  wire _7524_;
  wire _7525_;
  wire _7526_;
  wire _7527_;
  wire _7528_;
  wire _7529_;
  wire _7530_;
  wire _7531_;
  wire _7532_;
  wire _7533_;
  wire _7534_;
  wire _7535_;
  wire _7536_;
  wire _7537_;
  wire _7538_;
  wire _7539_;
  wire _7540_;
  wire _7541_;
  wire _7542_;
  wire _7543_;
  wire _7544_;
  wire _7545_;
  wire _7546_;
  wire _7547_;
  wire _7548_;
  wire _7549_;
  wire _7550_;
  wire _7551_;
  wire _7552_;
  wire _7553_;
  wire _7554_;
  wire _7555_;
  wire _7556_;
  wire _7557_;
  wire _7558_;
  wire _7559_;
  wire _7560_;
  wire _7561_;
  wire _7562_;
  wire _7563_;
  wire _7564_;
  wire _7565_;
  wire _7566_;
  wire _7567_;
  wire _7568_;
  wire _7569_;
  wire _7570_;
  wire _7571_;
  wire _7572_;
  wire _7573_;
  wire _7574_;
  wire _7575_;
  wire _7576_;
  wire _7577_;
  wire _7578_;
  wire _7579_;
  wire _7580_;
  wire _7581_;
  wire _7582_;
  wire _7583_;
  wire _7584_;
  wire _7585_;
  wire _7586_;
  wire _7587_;
  wire _7588_;
  wire _7589_;
  wire _7590_;
  wire _7591_;
  wire _7592_;
  wire _7593_;
  wire _7594_;
  wire _7595_;
  wire _7596_;
  wire _7597_;
  wire _7598_;
  wire _7599_;
  wire _7600_;
  wire _7601_;
  wire _7602_;
  wire _7603_;
  wire _7604_;
  wire _7605_;
  wire _7606_;
  wire _7607_;
  wire _7608_;
  wire _7609_;
  wire _7610_;
  wire _7611_;
  wire _7612_;
  wire _7613_;
  wire _7614_;
  wire _7615_;
  wire _7616_;
  wire _7617_;
  wire _7618_;
  wire _7619_;
  wire _7620_;
  wire _7621_;
  wire _7622_;
  wire _7623_;
  wire _7624_;
  wire _7625_;
  wire _7626_;
  wire _7627_;
  wire _7628_;
  wire _7629_;
  wire _7630_;
  wire _7631_;
  wire _7632_;
  wire _7633_;
  wire _7634_;
  wire _7635_;
  wire _7636_;
  wire _7637_;
  wire _7638_;
  wire _7639_;
  wire _7640_;
  wire _7641_;
  wire _7642_;
  wire _7643_;
  wire _7644_;
  wire _7645_;
  wire _7646_;
  wire _7647_;
  wire _7648_;
  wire _7649_;
  wire _7650_;
  wire _7651_;
  wire _7652_;
  wire _7653_;
  wire _7654_;
  wire _7655_;
  wire _7656_;
  wire _7657_;
  wire _7658_;
  wire _7659_;
  wire _7660_;
  wire _7661_;
  wire _7662_;
  wire _7663_;
  wire _7664_;
  wire _7665_;
  wire _7666_;
  wire _7667_;
  wire _7668_;
  wire _7669_;
  wire _7670_;
  wire _7671_;
  wire _7672_;
  wire _7673_;
  wire _7674_;
  wire _7675_;
  wire _7676_;
  wire _7677_;
  wire _7678_;
  wire _7679_;
  wire _7680_;
  wire _7681_;
  wire _7682_;
  wire _7683_;
  wire _7684_;
  wire _7685_;
  wire _7686_;
  wire _7687_;
  wire _7688_;
  wire _7689_;
  wire _7690_;
  wire _7691_;
  wire _7692_;
  wire _7693_;
  wire _7694_;
  wire _7695_;
  wire _7696_;
  wire _7697_;
  wire _7698_;
  wire _7699_;
  wire _7700_;
  wire _7701_;
  wire _7702_;
  wire _7703_;
  wire _7704_;
  wire _7705_;
  wire _7706_;
  wire _7707_;
  wire _7708_;
  wire _7709_;
  wire _7710_;
  wire _7711_;
  wire _7712_;
  wire _7713_;
  wire _7714_;
  wire _7715_;
  wire _7716_;
  wire _7717_;
  wire _7718_;
  wire _7719_;
  wire _7720_;
  wire _7721_;
  wire _7722_;
  wire _7723_;
  wire _7724_;
  wire _7725_;
  wire _7726_;
  wire _7727_;
  wire _7728_;
  wire _7729_;
  wire _7730_;
  wire _7731_;
  wire _7732_;
  wire _7733_;
  wire _7734_;
  wire _7735_;
  wire _7736_;
  wire _7737_;
  wire _7738_;
  wire _7739_;
  wire _7740_;
  wire _7741_;
  wire _7742_;
  wire _7743_;
  wire _7744_;
  wire _7745_;
  wire _7746_;
  wire _7747_;
  wire _7748_;
  wire _7749_;
  wire _7750_;
  wire _7751_;
  wire _7752_;
  wire _7753_;
  wire _7754_;
  wire _7755_;
  wire _7756_;
  wire _7757_;
  wire _7758_;
  wire _7759_;
  wire _7760_;
  wire _7761_;
  wire _7762_;
  wire _7763_;
  wire _7764_;
  wire _7765_;
  wire _7766_;
  wire _7767_;
  wire _7768_;
  wire _7769_;
  wire _7770_;
  wire _7771_;
  wire _7772_;
  wire _7773_;
  wire _7774_;
  wire _7775_;
  wire _7776_;
  wire _7777_;
  wire _7778_;
  wire _7779_;
  wire _7780_;
  wire _7781_;
  wire _7782_;
  wire _7783_;
  wire _7784_;
  wire _7785_;
  wire _7786_;
  wire _7787_;
  wire _7788_;
  wire _7789_;
  wire _7790_;
  wire _7791_;
  wire _7792_;
  wire _7793_;
  wire _7794_;
  wire _7795_;
  wire _7796_;
  wire _7797_;
  wire _7798_;
  wire _7799_;
  wire _7800_;
  wire _7801_;
  wire _7802_;
  wire _7803_;
  wire _7804_;
  wire _7805_;
  wire _7806_;
  wire _7807_;
  wire _7808_;
  wire _7809_;
  wire _7810_;
  wire _7811_;
  wire _7812_;
  wire _7813_;
  wire _7814_;
  wire _7815_;
  wire _7816_;
  wire _7817_;
  wire _7818_;
  wire _7819_;
  wire _7820_;
  wire _7821_;
  wire _7822_;
  wire _7823_;
  wire _7824_;
  wire _7825_;
  wire _7826_;
  wire _7827_;
  wire _7828_;
  wire _7829_;
  wire _7830_;
  wire _7831_;
  wire _7832_;
  wire _7833_;
  wire _7834_;
  wire _7835_;
  wire _7836_;
  wire _7837_;
  wire _7838_;
  wire _7839_;
  wire _7840_;
  wire _7841_;
  wire _7842_;
  wire _7843_;
  wire _7844_;
  wire _7845_;
  wire _7846_;
  wire _7847_;
  wire _7848_;
  wire _7849_;
  wire _7850_;
  wire _7851_;
  wire _7852_;
  wire _7853_;
  wire _7854_;
  wire _7855_;
  wire _7856_;
  wire _7857_;
  wire _7858_;
  wire _7859_;
  wire _7860_;
  wire _7861_;
  wire _7862_;
  wire _7863_;
  wire _7864_;
  wire _7865_;
  wire _7866_;
  wire _7867_;
  wire _7868_;
  wire _7869_;
  wire _7870_;
  wire _7871_;
  wire _7872_;
  wire _7873_;
  wire _7874_;
  wire _7875_;
  wire _7876_;
  wire _7877_;
  wire _7878_;
  wire _7879_;
  wire _7880_;
  wire _7881_;
  wire _7882_;
  wire _7883_;
  wire _7884_;
  wire _7885_;
  wire _7886_;
  wire _7887_;
  wire _7888_;
  wire _7889_;
  wire _7890_;
  wire _7891_;
  wire _7892_;
  wire _7893_;
  wire _7894_;
  wire _7895_;
  wire _7896_;
  wire _7897_;
  wire _7898_;
  wire _7899_;
  wire _7900_;
  wire _7901_;
  wire _7902_;
  wire _7903_;
  wire _7904_;
  wire _7905_;
  wire _7906_;
  wire _7907_;
  wire _7908_;
  wire _7909_;
  wire _7910_;
  wire _7911_;
  wire _7912_;
  wire _7913_;
  wire _7914_;
  wire _7915_;
  wire _7916_;
  wire _7917_;
  wire _7918_;
  wire _7919_;
  wire _7920_;
  wire _7921_;
  wire _7922_;
  wire _7923_;
  wire _7924_;
  wire _7925_;
  wire _7926_;
  wire _7927_;
  wire _7928_;
  wire _7929_;
  wire _7930_;
  wire _7931_;
  wire _7932_;
  wire _7933_;
  wire _7934_;
  wire _7935_;
  wire _7936_;
  wire _7937_;
  wire _7938_;
  wire _7939_;
  wire _7940_;
  wire _7941_;
  wire _7942_;
  wire _7943_;
  wire _7944_;
  wire _7945_;
  wire _7946_;
  wire _7947_;
  wire _7948_;
  wire _7949_;
  wire _7950_;
  wire _7951_;
  wire _7952_;
  wire _7953_;
  wire _7954_;
  wire _7955_;
  wire _7956_;
  wire _7957_;
  wire _7958_;
  wire _7959_;
  wire _7960_;
  wire _7961_;
  wire _7962_;
  wire _7963_;
  wire _7964_;
  wire _7965_;
  wire _7966_;
  wire _7967_;
  wire _7968_;
  wire _7969_;
  wire _7970_;
  wire _7971_;
  wire _7972_;
  wire _7973_;
  wire _7974_;
  wire _7975_;
  wire _7976_;
  wire _7977_;
  wire _7978_;
  wire _7979_;
  wire _7980_;
  wire _7981_;
  wire _7982_;
  wire _7983_;
  wire _7984_;
  wire _7985_;
  wire _7986_;
  wire _7987_;
  wire _7988_;
  wire _7989_;
  wire _7990_;
  wire _7991_;
  wire _7992_;
  wire _7993_;
  wire _7994_;
  wire _7995_;
  wire _7996_;
  wire _7997_;
  wire _7998_;
  wire _7999_;
  wire _8000_;
  wire _8001_;
  wire _8002_;
  wire _8003_;
  wire _8004_;
  wire _8005_;
  wire _8006_;
  wire _8007_;
  wire _8008_;
  wire _8009_;
  wire _8010_;
  wire _8011_;
  wire _8012_;
  wire _8013_;
  wire _8014_;
  wire _8015_;
  wire _8016_;
  wire _8017_;
  wire _8018_;
  wire _8019_;
  wire _8020_;
  wire _8021_;
  wire _8022_;
  wire _8023_;
  wire _8024_;
  wire _8025_;
  wire _8026_;
  wire _8027_;
  wire _8028_;
  wire _8029_;
  wire _8030_;
  wire _8031_;
  wire _8032_;
  wire _8033_;
  wire _8034_;
  wire _8035_;
  wire _8036_;
  wire _8037_;
  wire _8038_;
  wire _8039_;
  wire _8040_;
  wire _8041_;
  wire _8042_;
  wire _8043_;
  wire _8044_;
  wire _8045_;
  wire _8046_;
  wire _8047_;
  wire _8048_;
  wire _8049_;
  wire _8050_;
  wire _8051_;
  wire _8052_;
  wire _8053_;
  wire _8054_;
  wire _8055_;
  wire _8056_;
  wire _8057_;
  wire _8058_;
  wire _8059_;
  wire _8060_;
  wire _8061_;
  wire _8062_;
  wire _8063_;
  wire _8064_;
  wire _8065_;
  wire _8066_;
  wire _8067_;
  wire _8068_;
  wire _8069_;
  wire _8070_;
  wire _8071_;
  wire _8072_;
  wire _8073_;
  wire _8074_;
  wire _8075_;
  wire _8076_;
  wire _8077_;
  wire _8078_;
  wire _8079_;
  wire _8080_;
  wire _8081_;
  wire _8082_;
  wire _8083_;
  wire _8084_;
  wire _8085_;
  wire _8086_;
  wire _8087_;
  wire _8088_;
  wire _8089_;
  wire _8090_;
  wire _8091_;
  wire _8092_;
  wire _8093_;
  wire _8094_;
  wire _8095_;
  wire _8096_;
  wire _8097_;
  wire _8098_;
  wire _8099_;
  wire _8100_;
  wire _8101_;
  wire _8102_;
  wire _8103_;
  wire _8104_;
  wire _8105_;
  wire _8106_;
  wire _8107_;
  wire _8108_;
  wire _8109_;
  wire _8110_;
  wire _8111_;
  wire _8112_;
  wire _8113_;
  wire _8114_;
  wire _8115_;
  wire _8116_;
  wire _8117_;
  wire _8118_;
  wire _8119_;
  wire _8120_;
  wire _8121_;
  wire _8122_;
  wire _8123_;
  wire _8124_;
  wire _8125_;
  wire _8126_;
  wire _8127_;
  wire _8128_;
  wire _8129_;
  wire _8130_;
  wire _8131_;
  wire _8132_;
  wire _8133_;
  wire _8134_;
  wire _8135_;
  wire _8136_;
  wire _8137_;
  wire _8138_;
  wire _8139_;
  wire _8140_;
  wire _8141_;
  wire _8142_;
  wire _8143_;
  wire _8144_;
  wire _8145_;
  wire _8146_;
  wire _8147_;
  wire _8148_;
  wire _8149_;
  wire _8150_;
  wire _8151_;
  wire _8152_;
  wire _8153_;
  wire _8154_;
  wire _8155_;
  wire _8156_;
  wire _8157_;
  wire _8158_;
  wire _8159_;
  wire _8160_;
  wire _8161_;
  wire _8162_;
  wire _8163_;
  wire _8164_;
  wire _8165_;
  wire _8166_;
  wire _8167_;
  wire _8168_;
  wire _8169_;
  wire _8170_;
  wire _8171_;
  wire _8172_;
  wire _8173_;
  wire _8174_;
  wire _8175_;
  wire _8176_;
  wire _8177_;
  wire _8178_;
  wire _8179_;
  wire _8180_;
  wire _8181_;
  wire _8182_;
  wire _8183_;
  wire _8184_;
  wire _8185_;
  wire _8186_;
  wire _8187_;
  wire _8188_;
  wire _8189_;
  wire _8190_;
  wire _8191_;
  wire _8192_;
  wire _8193_;
  wire _8194_;
  wire _8195_;
  wire _8196_;
  wire _8197_;
  wire _8198_;
  wire _8199_;
  wire _8200_;
  wire _8201_;
  wire _8202_;
  wire _8203_;
  wire _8204_;
  wire _8205_;
  wire _8206_;
  wire _8207_;
  wire _8208_;
  wire _8209_;
  wire _8210_;
  wire _8211_;
  wire _8212_;
  wire _8213_;
  wire _8214_;
  wire _8215_;
  wire _8216_;
  wire _8217_;
  wire _8218_;
  wire _8219_;
  wire _8220_;
  wire _8221_;
  wire _8222_;
  wire _8223_;
  wire _8224_;
  wire _8225_;
  wire _8226_;
  wire _8227_;
  wire _8228_;
  wire _8229_;
  wire _8230_;
  wire _8231_;
  wire _8232_;
  wire _8233_;
  wire _8234_;
  wire _8235_;
  wire _8236_;
  wire _8237_;
  wire _8238_;
  wire _8239_;
  wire _8240_;
  wire _8241_;
  wire _8242_;
  wire _8243_;
  wire _8244_;
  wire _8245_;
  wire _8246_;
  wire _8247_;
  wire _8248_;
  wire _8249_;
  wire _8250_;
  wire _8251_;
  wire _8252_;
  wire _8253_;
  wire _8254_;
  wire _8255_;
  wire _8256_;
  wire _8257_;
  wire _8258_;
  wire _8259_;
  wire _8260_;
  wire _8261_;
  wire _8262_;
  wire _8263_;
  wire _8264_;
  wire _8265_;
  wire _8266_;
  wire _8267_;
  wire _8268_;
  wire _8269_;
  wire _8270_;
  wire _8271_;
  wire _8272_;
  wire _8273_;
  wire _8274_;
  wire _8275_;
  wire _8276_;
  wire _8277_;
  wire _8278_;
  wire _8279_;
  wire _8280_;
  wire _8281_;
  wire _8282_;
  wire _8283_;
  wire _8284_;
  wire _8285_;
  wire _8286_;
  wire _8287_;
  wire _8288_;
  wire _8289_;
  wire _8290_;
  wire _8291_;
  wire _8292_;
  wire _8293_;
  wire _8294_;
  wire _8295_;
  wire _8296_;
  wire _8297_;
  wire _8298_;
  wire _8299_;
  wire _8300_;
  wire _8301_;
  wire _8302_;
  wire _8303_;
  wire _8304_;
  wire _8305_;
  wire _8306_;
  wire _8307_;
  wire _8308_;
  wire _8309_;
  wire _8310_;
  wire _8311_;
  wire _8312_;
  wire _8313_;
  wire _8314_;
  wire _8315_;
  wire _8316_;
  wire _8317_;
  wire _8318_;
  wire _8319_;
  wire _8320_;
  wire _8321_;
  wire _8322_;
  wire _8323_;
  wire _8324_;
  wire _8325_;
  wire _8326_;
  wire _8327_;
  wire _8328_;
  wire _8329_;
  wire _8330_;
  wire _8331_;
  wire _8332_;
  wire _8333_;
  wire _8334_;
  wire _8335_;
  wire _8336_;
  wire _8337_;
  wire _8338_;
  wire _8339_;
  wire _8340_;
  wire _8341_;
  wire _8342_;
  wire _8343_;
  wire _8344_;
  wire _8345_;
  wire _8346_;
  wire _8347_;
  wire _8348_;
  wire _8349_;
  wire _8350_;
  wire _8351_;
  wire _8352_;
  wire _8353_;
  wire _8354_;
  wire _8355_;
  wire _8356_;
  wire _8357_;
  wire _8358_;
  wire _8359_;
  wire _8360_;
  wire _8361_;
  wire _8362_;
  wire _8363_;
  wire _8364_;
  wire _8365_;
  wire _8366_;
  wire _8367_;
  wire _8368_;
  wire _8369_;
  wire _8370_;
  wire _8371_;
  wire _8372_;
  wire _8373_;
  wire _8374_;
  wire _8375_;
  wire _8376_;
  wire _8377_;
  wire _8378_;
  wire _8379_;
  wire _8380_;
  wire _8381_;
  wire _8382_;
  wire _8383_;
  wire _8384_;
  wire _8385_;
  wire _8386_;
  wire _8387_;
  wire _8388_;
  wire _8389_;
  wire _8390_;
  wire _8391_;
  wire _8392_;
  wire _8393_;
  wire _8394_;
  wire _8395_;
  wire _8396_;
  wire _8397_;
  wire _8398_;
  wire _8399_;
  wire _8400_;
  wire _8401_;
  wire _8402_;
  wire _8403_;
  wire _8404_;
  wire _8405_;
  wire _8406_;
  wire _8407_;
  wire _8408_;
  wire _8409_;
  wire _8410_;
  wire _8411_;
  wire _8412_;
  wire _8413_;
  wire _8414_;
  wire _8415_;
  wire _8416_;
  wire _8417_;
  wire _8418_;
  wire _8419_;
  wire _8420_;
  wire _8421_;
  wire _8422_;
  wire _8423_;
  wire _8424_;
  wire _8425_;
  wire _8426_;
  wire _8427_;
  wire _8428_;
  wire _8429_;
  wire _8430_;
  wire _8431_;
  wire _8432_;
  wire _8433_;
  wire _8434_;
  wire _8435_;
  wire _8436_;
  wire _8437_;
  wire _8438_;
  wire _8439_;
  wire _8440_;
  wire _8441_;
  wire _8442_;
  wire _8443_;
  wire _8444_;
  wire _8445_;
  wire _8446_;
  wire _8447_;
  wire _8448_;
  wire _8449_;
  wire _8450_;
  wire _8451_;
  wire _8452_;
  wire _8453_;
  wire _8454_;
  wire _8455_;
  wire _8456_;
  wire _8457_;
  wire _8458_;
  wire _8459_;
  wire _8460_;
  wire _8461_;
  wire _8462_;
  wire _8463_;
  wire _8464_;
  wire _8465_;
  wire _8466_;
  wire _8467_;
  wire _8468_;
  wire _8469_;
  wire _8470_;
  wire _8471_;
  wire _8472_;
  wire _8473_;
  wire _8474_;
  wire _8475_;
  wire _8476_;
  wire _8477_;
  wire _8478_;
  wire _8479_;
  wire _8480_;
  wire _8481_;
  wire _8482_;
  wire _8483_;
  wire _8484_;
  wire _8485_;
  wire _8486_;
  wire _8487_;
  wire _8488_;
  wire _8489_;
  wire _8490_;
  wire _8491_;
  wire _8492_;
  wire _8493_;
  wire _8494_;
  wire _8495_;
  wire _8496_;
  wire _8497_;
  wire _8498_;
  wire _8499_;
  wire _8500_;
  wire _8501_;
  wire _8502_;
  wire _8503_;
  wire _8504_;
  wire _8505_;
  wire _8506_;
  wire _8507_;
  wire _8508_;
  wire _8509_;
  wire _8510_;
  wire _8511_;
  wire _8512_;
  wire _8513_;
  wire _8514_;
  wire _8515_;
  wire _8516_;
  wire _8517_;
  wire _8518_;
  wire _8519_;
  wire _8520_;
  wire _8521_;
  wire _8522_;
  wire _8523_;
  wire _8524_;
  wire _8525_;
  wire _8526_;
  wire _8527_;
  wire _8528_;
  wire _8529_;
  wire _8530_;
  wire _8531_;
  wire _8532_;
  wire _8533_;
  wire _8534_;
  wire _8535_;
  wire _8536_;
  wire _8537_;
  wire _8538_;
  wire _8539_;
  wire _8540_;
  wire _8541_;
  wire _8542_;
  wire _8543_;
  wire _8544_;
  wire _8545_;
  wire _8546_;
  wire _8547_;
  wire _8548_;
  wire _8549_;
  wire _8550_;
  wire _8551_;
  wire _8552_;
  wire _8553_;
  wire _8554_;
  wire _8555_;
  wire _8556_;
  wire _8557_;
  wire _8558_;
  wire _8559_;
  wire _8560_;
  wire _8561_;
  wire _8562_;
  wire _8563_;
  wire _8564_;
  wire _8565_;
  wire _8566_;
  wire _8567_;
  wire _8568_;
  wire _8569_;
  wire _8570_;
  wire _8571_;
  wire _8572_;
  wire _8573_;
  wire _8574_;
  wire _8575_;
  wire _8576_;
  wire _8577_;
  wire _8578_;
  wire _8579_;
  wire _8580_;
  wire _8581_;
  wire _8582_;
  wire _8583_;
  wire _8584_;
  wire _8585_;
  wire _8586_;
  wire _8587_;
  wire _8588_;
  wire _8589_;
  wire _8590_;
  wire _8591_;
  wire _8592_;
  wire _8593_;
  wire _8594_;
  wire _8595_;
  wire _8596_;
  wire _8597_;
  wire _8598_;
  wire _8599_;
  wire _8600_;
  wire _8601_;
  wire _8602_;
  wire _8603_;
  wire _8604_;
  wire _8605_;
  wire _8606_;
  wire _8607_;
  wire _8608_;
  wire _8609_;
  wire _8610_;
  wire _8611_;
  wire _8612_;
  wire _8613_;
  wire _8614_;
  wire _8615_;
  wire _8616_;
  wire _8617_;
  wire _8618_;
  wire _8619_;
  wire _8620_;
  wire _8621_;
  wire _8622_;
  wire _8623_;
  wire _8624_;
  wire _8625_;
  wire _8626_;
  wire _8627_;
  wire _8628_;
  wire _8629_;
  wire _8630_;
  wire _8631_;
  wire _8632_;
  wire _8633_;
  wire _8634_;
  wire _8635_;
  wire _8636_;
  wire _8637_;
  wire _8638_;
  wire _8639_;
  wire _8640_;
  wire _8641_;
  wire _8642_;
  wire _8643_;
  wire _8644_;
  wire _8645_;
  wire _8646_;
  wire _8647_;
  wire _8648_;
  wire _8649_;
  wire _8650_;
  wire _8651_;
  wire _8652_;
  wire _8653_;
  wire _8654_;
  wire _8655_;
  wire _8656_;
  wire _8657_;
  wire _8658_;
  wire _8659_;
  wire _8660_;
  wire _8661_;
  wire _8662_;
  wire _8663_;
  wire _8664_;
  wire _8665_;
  wire _8666_;
  wire _8667_;
  wire _8668_;
  wire _8669_;
  wire _8670_;
  wire _8671_;
  wire _8672_;
  wire _8673_;
  wire _8674_;
  wire _8675_;
  wire _8676_;
  wire _8677_;
  wire _8678_;
  wire _8679_;
  wire _8680_;
  wire _8681_;
  wire _8682_;
  wire _8683_;
  wire _8684_;
  wire _8685_;
  wire _8686_;
  wire _8687_;
  wire _8688_;
  wire _8689_;
  wire _8690_;
  wire _8691_;
  wire _8692_;
  wire _8693_;
  wire _8694_;
  wire _8695_;
  wire _8696_;
  wire _8697_;
  wire _8698_;
  wire _8699_;
  wire _8700_;
  wire _8701_;
  wire _8702_;
  wire _8703_;
  wire _8704_;
  wire _8705_;
  wire _8706_;
  wire _8707_;
  wire _8708_;
  wire _8709_;
  wire _8710_;
  wire _8711_;
  wire _8712_;
  wire _8713_;
  wire _8714_;
  wire _8715_;
  wire _8716_;
  wire _8717_;
  wire _8718_;
  wire _8719_;
  wire _8720_;
  wire _8721_;
  wire _8722_;
  wire _8723_;
  wire _8724_;
  wire _8725_;
  wire _8726_;
  wire _8727_;
  wire _8728_;
  wire _8729_;
  wire _8730_;
  wire _8731_;
  wire _8732_;
  wire _8733_;
  wire _8734_;
  wire _8735_;
  wire _8736_;
  wire _8737_;
  wire _8738_;
  wire _8739_;
  wire _8740_;
  wire _8741_;
  wire _8742_;
  wire _8743_;
  wire _8744_;
  wire _8745_;
  wire _8746_;
  wire _8747_;
  wire _8748_;
  wire _8749_;
  wire _8750_;
  wire _8751_;
  wire _8752_;
  wire _8753_;
  wire _8754_;
  wire _8755_;
  wire _8756_;
  wire _8757_;
  wire _8758_;
  wire _8759_;
  wire _8760_;
  wire _8761_;
  wire _8762_;
  wire _8763_;
  wire _8764_;
  wire _8765_;
  wire _8766_;
  wire _8767_;
  wire _8768_;
  wire _8769_;
  wire _8770_;
  wire _8771_;
  wire _8772_;
  wire _8773_;
  wire _8774_;
  wire _8775_;
  wire _8776_;
  wire _8777_;
  wire _8778_;
  wire _8779_;
  wire _8780_;
  wire _8781_;
  wire _8782_;
  wire _8783_;
  wire _8784_;
  wire _8785_;
  wire _8786_;
  wire _8787_;
  wire _8788_;
  wire _8789_;
  wire _8790_;
  wire _8791_;
  wire _8792_;
  wire _8793_;
  wire _8794_;
  wire _8795_;
  wire _8796_;
  wire _8797_;
  wire _8798_;
  wire _8799_;
  wire _8800_;
  wire _8801_;
  wire _8802_;
  wire _8803_;
  wire _8804_;
  wire _8805_;
  wire _8806_;
  wire _8807_;
  wire _8808_;
  wire _8809_;
  wire _8810_;
  wire _8811_;
  wire _8812_;
  wire _8813_;
  wire _8814_;
  wire _8815_;
  wire _8816_;
  wire _8817_;
  wire _8818_;
  wire _8819_;
  wire _8820_;
  wire _8821_;
  wire _8822_;
  wire _8823_;
  wire _8824_;
  wire _8825_;
  wire _8826_;
  wire _8827_;
  wire _8828_;
  wire _8829_;
  wire _8830_;
  wire _8831_;
  wire _8832_;
  wire _8833_;
  wire _8834_;
  wire _8835_;
  wire _8836_;
  wire _8837_;
  wire _8838_;
  wire _8839_;
  wire _8840_;
  wire _8841_;
  wire _8842_;
  wire _8843_;
  wire _8844_;
  wire _8845_;
  wire _8846_;
  wire _8847_;
  wire _8848_;
  wire _8849_;
  wire _8850_;
  wire _8851_;
  wire _8852_;
  wire _8853_;
  wire _8854_;
  wire _8855_;
  wire _8856_;
  wire _8857_;
  wire _8858_;
  wire _8859_;
  wire _8860_;
  wire _8861_;
  wire _8862_;
  wire _8863_;
  wire _8864_;
  wire _8865_;
  wire _8866_;
  wire _8867_;
  wire _8868_;
  wire _8869_;
  wire _8870_;
  wire _8871_;
  wire _8872_;
  wire _8873_;
  wire _8874_;
  wire _8875_;
  wire _8876_;
  wire _8877_;
  wire _8878_;
  wire _8879_;
  wire _8880_;
  wire _8881_;
  wire _8882_;
  wire _8883_;
  wire _8884_;
  wire _8885_;
  wire _8886_;
  wire _8887_;
  wire _8888_;
  wire _8889_;
  wire _8890_;
  wire _8891_;
  wire _8892_;
  wire _8893_;
  wire _8894_;
  wire _8895_;
  wire _8896_;
  wire _8897_;
  wire _8898_;
  wire _8899_;
  wire _8900_;
  wire _8901_;
  wire _8902_;
  wire _8903_;
  wire _8904_;
  wire _8905_;
  wire _8906_;
  wire _8907_;
  wire _8908_;
  wire _8909_;
  wire _8910_;
  wire _8911_;
  wire _8912_;
  wire _8913_;
  wire _8914_;
  wire _8915_;
  wire _8916_;
  wire _8917_;
  wire _8918_;
  wire _8919_;
  wire _8920_;
  wire _8921_;
  wire _8922_;
  wire _8923_;
  wire _8924_;
  wire _8925_;
  wire _8926_;
  wire _8927_;
  wire _8928_;
  wire _8929_;
  wire _8930_;
  wire _8931_;
  wire _8932_;
  wire _8933_;
  wire _8934_;
  wire _8935_;
  wire _8936_;
  wire _8937_;
  wire _8938_;
  wire _8939_;
  wire _8940_;
  wire _8941_;
  wire _8942_;
  wire _8943_;
  wire _8944_;
  wire _8945_;
  wire _8946_;
  wire _8947_;
  wire _8948_;
  wire _8949_;
  wire _8950_;
  wire _8951_;
  wire _8952_;
  wire _8953_;
  wire _8954_;
  wire _8955_;
  wire _8956_;
  wire _8957_;
  wire _8958_;
  wire _8959_;
  wire _8960_;
  wire _8961_;
  wire _8962_;
  wire _8963_;
  wire _8964_;
  wire _8965_;
  wire _8966_;
  wire _8967_;
  wire _8968_;
  wire _8969_;
  wire _8970_;
  wire _8971_;
  wire _8972_;
  wire _8973_;
  wire _8974_;
  wire _8975_;
  wire _8976_;
  wire _8977_;
  wire _8978_;
  wire _8979_;
  wire _8980_;
  wire _8981_;
  wire _8982_;
  wire _8983_;
  wire _8984_;
  wire _8985_;
  wire _8986_;
  wire _8987_;
  wire _8988_;
  wire _8989_;
  wire _8990_;
  wire _8991_;
  wire _8992_;
  wire _8993_;
  wire _8994_;
  wire _8995_;
  wire _8996_;
  wire _8997_;
  wire _8998_;
  wire _8999_;
  wire _9000_;
  wire _9001_;
  wire _9002_;
  wire _9003_;
  wire _9004_;
  wire _9005_;
  wire _9006_;
  wire _9007_;
  wire _9008_;
  wire _9009_;
  wire _9010_;
  wire _9011_;
  wire _9012_;
  wire _9013_;
  wire _9014_;
  wire _9015_;
  wire _9016_;
  wire _9017_;
  wire _9018_;
  wire _9019_;
  wire _9020_;
  wire _9021_;
  wire _9022_;
  wire _9023_;
  wire _9024_;
  wire _9025_;
  wire _9026_;
  wire _9027_;
  wire _9028_;
  wire _9029_;
  wire _9030_;
  wire _9031_;
  wire _9032_;
  wire _9033_;
  wire _9034_;
  wire _9035_;
  wire _9036_;
  wire _9037_;
  wire _9038_;
  wire _9039_;
  wire _9040_;
  wire _9041_;
  wire _9042_;
  wire _9043_;
  wire _9044_;
  wire _9045_;
  wire _9046_;
  wire _9047_;
  wire _9048_;
  wire _9049_;
  wire _9050_;
  wire _9051_;
  wire _9052_;
  wire _9053_;
  wire _9054_;
  wire _9055_;
  wire _9056_;
  wire _9057_;
  wire _9058_;
  wire _9059_;
  wire _9060_;
  wire _9061_;
  wire _9062_;
  wire _9063_;
  wire _9064_;
  wire _9065_;
  wire _9066_;
  wire _9067_;
  wire _9068_;
  wire _9069_;
  wire _9070_;
  wire _9071_;
  wire _9072_;
  wire _9073_;
  wire _9074_;
  wire _9075_;
  wire _9076_;
  wire _9077_;
  wire _9078_;
  wire _9079_;
  wire _9080_;
  wire _9081_;
  wire _9082_;
  wire _9083_;
  wire _9084_;
  wire _9085_;
  wire _9086_;
  wire _9087_;
  wire _9088_;
  wire _9089_;
  wire _9090_;
  wire _9091_;
  wire _9092_;
  wire _9093_;
  wire _9094_;
  wire _9095_;
  wire _9096_;
  wire _9097_;
  wire _9098_;
  wire _9099_;
  wire _9100_;
  wire _9101_;
  wire _9102_;
  wire _9103_;
  wire _9104_;
  wire _9105_;
  wire _9106_;
  wire _9107_;
  wire _9108_;
  wire _9109_;
  wire _9110_;
  wire _9111_;
  wire _9112_;
  wire _9113_;
  wire _9114_;
  wire _9115_;
  wire _9116_;
  wire _9117_;
  wire _9118_;
  wire _9119_;
  wire _9120_;
  wire _9121_;
  wire _9122_;
  wire _9123_;
  wire _9124_;
  wire _9125_;
  wire _9126_;
  wire _9127_;
  wire _9128_;
  wire _9129_;
  wire _9130_;
  wire _9131_;
  wire _9132_;
  wire _9133_;
  wire _9134_;
  wire _9135_;
  wire _9136_;
  wire _9137_;
  wire _9138_;
  wire _9139_;
  wire _9140_;
  wire _9141_;
  wire _9142_;
  wire _9143_;
  wire _9144_;
  wire _9145_;
  wire _9146_;
  wire _9147_;
  wire _9148_;
  wire _9149_;
  wire _9150_;
  wire _9151_;
  wire _9152_;
  wire _9153_;
  wire _9154_;
  wire _9155_;
  wire _9156_;
  wire _9157_;
  wire _9158_;
  wire _9159_;
  wire _9160_;
  wire _9161_;
  wire _9162_;
  wire _9163_;
  wire _9164_;
  wire _9165_;
  wire _9166_;
  wire _9167_;
  wire _9168_;
  wire _9169_;
  wire _9170_;
  wire _9171_;
  wire _9172_;
  wire _9173_;
  wire _9174_;
  wire _9175_;
  wire _9176_;
  wire _9177_;
  wire _9178_;
  wire _9179_;
  wire _9180_;
  wire _9181_;
  wire _9182_;
  wire _9183_;
  wire _9184_;
  wire _9185_;
  wire _9186_;
  wire _9187_;
  wire _9188_;
  wire _9189_;
  wire _9190_;
  wire _9191_;
  wire _9192_;
  wire _9193_;
  wire _9194_;
  wire _9195_;
  wire _9196_;
  wire _9197_;
  wire _9198_;
  wire _9199_;
  wire _9200_;
  wire _9201_;
  wire _9202_;
  wire _9203_;
  wire _9204_;
  wire _9205_;
  wire _9206_;
  wire _9207_;
  wire _9208_;
  wire _9209_;
  wire _9210_;
  wire _9211_;
  wire _9212_;
  wire _9213_;
  wire _9214_;
  wire _9215_;
  wire _9216_;
  wire _9217_;
  wire _9218_;
  wire _9219_;
  wire _9220_;
  wire _9221_;
  wire _9222_;
  wire _9223_;
  wire _9224_;
  wire _9225_;
  wire _9226_;
  wire _9227_;
  wire _9228_;
  wire _9229_;
  wire _9230_;
  wire _9231_;
  wire _9232_;
  wire _9233_;
  wire _9234_;
  wire _9235_;
  wire _9236_;
  wire _9237_;
  wire _9238_;
  wire _9239_;
  wire _9240_;
  wire _9241_;
  wire _9242_;
  wire _9243_;
  wire _9244_;
  wire _9245_;
  wire _9246_;
  wire _9247_;
  wire _9248_;
  wire _9249_;
  wire _9250_;
  wire _9251_;
  wire _9252_;
  wire _9253_;
  wire _9254_;
  wire _9255_;
  wire _9256_;
  wire _9257_;
  wire _9258_;
  wire _9259_;
  wire _9260_;
  wire _9261_;
  wire _9262_;
  wire _9263_;
  wire _9264_;
  wire _9265_;
  wire _9266_;
  wire _9267_;
  wire _9268_;
  wire _9269_;
  wire _9270_;
  wire _9271_;
  wire _9272_;
  wire _9273_;
  wire _9274_;
  wire _9275_;
  wire _9276_;
  wire _9277_;
  wire _9278_;
  wire _9279_;
  wire _9280_;
  wire _9281_;
  wire _9282_;
  wire _9283_;
  wire _9284_;
  wire _9285_;
  wire _9286_;
  wire _9287_;
  wire _9288_;
  wire _9289_;
  wire _9290_;
  wire _9291_;
  wire _9292_;
  wire _9293_;
  wire _9294_;
  wire _9295_;
  wire _9296_;
  wire _9297_;
  wire _9298_;
  wire _9299_;
  wire _9300_;
  wire _9301_;
  wire _9302_;
  wire _9303_;
  wire _9304_;
  wire _9305_;
  wire _9306_;
  wire _9307_;
  wire _9308_;
  wire _9309_;
  wire _9310_;
  wire _9311_;
  wire _9312_;
  wire _9313_;
  wire _9314_;
  wire _9315_;
  wire _9316_;
  wire _9317_;
  wire _9318_;
  wire _9319_;
  wire _9320_;
  wire _9321_;
  wire _9322_;
  wire _9323_;
  wire _9324_;
  wire _9325_;
  wire _9326_;
  wire _9327_;
  wire _9328_;
  wire _9329_;
  wire _9330_;
  wire _9331_;
  wire _9332_;
  wire _9333_;
  wire _9334_;
  wire _9335_;
  wire _9336_;
  wire _9337_;
  wire _9338_;
  wire _9339_;
  wire _9340_;
  wire _9341_;
  wire _9342_;
  wire _9343_;
  wire _9344_;
  wire _9345_;
  wire _9346_;
  wire _9347_;
  wire _9348_;
  wire _9349_;
  wire _9350_;
  wire _9351_;
  wire _9352_;
  wire _9353_;
  wire _9354_;
  wire _9355_;
  wire _9356_;
  wire _9357_;
  wire _9358_;
  wire _9359_;
  wire _9360_;
  wire _9361_;
  wire _9362_;
  wire _9363_;
  wire _9364_;
  wire _9365_;
  wire _9366_;
  wire _9367_;
  wire _9368_;
  wire _9369_;
  wire _9370_;
  wire _9371_;
  wire _9372_;
  wire _9373_;
  wire _9374_;
  wire _9375_;
  wire _9376_;
  wire _9377_;
  wire _9378_;
  wire _9379_;
  wire _9380_;
  wire _9381_;
  wire _9382_;
  wire _9383_;
  wire _9384_;
  wire _9385_;
  wire _9386_;
  wire _9387_;
  wire _9388_;
  wire _9389_;
  wire _9390_;
  wire _9391_;
  wire _9392_;
  wire _9393_;
  wire _9394_;
  wire _9395_;
  wire _9396_;
  wire _9397_;
  wire _9398_;
  wire _9399_;
  wire _9400_;
  wire _9401_;
  wire _9402_;
  wire _9403_;
  wire _9404_;
  wire _9405_;
  wire _9406_;
  wire _9407_;
  wire _9408_;
  wire _9409_;
  wire _9410_;
  wire _9411_;
  wire _9412_;
  wire _9413_;
  wire _9414_;
  wire _9415_;
  wire _9416_;
  wire _9417_;
  wire _9418_;
  wire _9419_;
  wire _9420_;
  wire _9421_;
  wire _9422_;
  wire _9423_;
  wire _9424_;
  wire _9425_;
  wire _9426_;
  wire _9427_;
  wire _9428_;
  wire _9429_;
  wire _9430_;
  wire _9431_;
  wire _9432_;
  wire _9433_;
  wire _9434_;
  wire _9435_;
  wire _9436_;
  wire _9437_;
  wire _9438_;
  wire _9439_;
  wire _9440_;
  wire _9441_;
  wire _9442_;
  wire _9443_;
  wire _9444_;
  wire _9445_;
  wire _9446_;
  wire _9447_;
  wire _9448_;
  wire _9449_;
  wire _9450_;
  wire _9451_;
  wire _9452_;
  wire _9453_;
  wire _9454_;
  wire _9455_;
  wire _9456_;
  wire _9457_;
  wire _9458_;
  wire _9459_;
  wire _9460_;
  wire _9461_;
  wire _9462_;
  wire _9463_;
  wire _9464_;
  wire _9465_;
  wire _9466_;
  wire _9467_;
  wire _9468_;
  wire _9469_;
  wire _9470_;
  wire _9471_;
  wire _9472_;
  wire _9473_;
  wire _9474_;
  wire _9475_;
  wire _9476_;
  wire _9477_;
  wire _9478_;
  wire _9479_;
  wire _9480_;
  wire _9481_;
  wire _9482_;
  wire _9483_;
  wire _9484_;
  wire _9485_;
  wire _9486_;
  wire _9487_;
  wire _9488_;
  wire _9489_;
  wire _9490_;
  wire _9491_;
  wire _9492_;
  wire _9493_;
  wire _9494_;
  wire _9495_;
  wire _9496_;
  wire _9497_;
  wire _9498_;
  wire _9499_;
  wire _9500_;
  wire _9501_;
  wire _9502_;
  wire _9503_;
  wire _9504_;
  wire _9505_;
  wire _9506_;
  wire _9507_;
  wire _9508_;
  wire _9509_;
  wire _9510_;
  wire _9511_;
  wire _9512_;
  wire _9513_;
  wire _9514_;
  wire _9515_;
  wire _9516_;
  wire _9517_;
  wire _9518_;
  wire _9519_;
  wire _9520_;
  wire _9521_;
  wire _9522_;
  wire _9523_;
  wire _9524_;
  wire _9525_;
  wire _9526_;
  wire _9527_;
  wire _9528_;
  wire _9529_;
  wire _9530_;
  wire _9531_;
  wire _9532_;
  wire _9533_;
  wire _9534_;
  wire _9535_;
  wire _9536_;
  wire _9537_;
  wire _9538_;
  wire _9539_;
  wire _9540_;
  wire _9541_;
  wire _9542_;
  wire _9543_;
  wire _9544_;
  wire _9545_;
  wire _9546_;
  wire _9547_;
  wire _9548_;
  wire _9549_;
  wire _9550_;
  wire _9551_;
  wire _9552_;
  wire _9553_;
  wire _9554_;
  wire _9555_;
  wire _9556_;
  wire _9557_;
  wire _9558_;
  wire _9559_;
  wire _9560_;
  wire _9561_;
  wire _9562_;
  wire _9563_;
  wire _9564_;
  wire _9565_;
  wire _9566_;
  wire _9567_;
  wire _9568_;
  wire _9569_;
  wire _9570_;
  wire _9571_;
  wire _9572_;
  wire _9573_;
  wire _9574_;
  wire _9575_;
  wire _9576_;
  wire _9577_;
  wire _9578_;
  wire _9579_;
  wire _9580_;
  wire _9581_;
  wire _9582_;
  wire _9583_;
  wire _9584_;
  wire _9585_;
  wire _9586_;
  wire _9587_;
  wire _9588_;
  wire _9589_;
  wire _9590_;
  wire _9591_;
  wire _9592_;
  wire _9593_;
  wire _9594_;
  wire _9595_;
  wire _9596_;
  wire _9597_;
  wire _9598_;
  wire _9599_;
  wire _9600_;
  wire _9601_;
  wire _9602_;
  wire _9603_;
  wire _9604_;
  wire _9605_;
  wire _9606_;
  wire _9607_;
  wire _9608_;
  wire _9609_;
  wire _9610_;
  wire _9611_;
  wire _9612_;
  wire _9613_;
  wire _9614_;
  wire _9615_;
  wire _9616_;
  wire _9617_;
  wire _9618_;
  wire _9619_;
  wire _9620_;
  wire _9621_;
  wire _9622_;
  wire _9623_;
  wire _9624_;
  wire _9625_;
  wire _9626_;
  wire _9627_;
  wire _9628_;
  wire _9629_;
  wire _9630_;
  wire _9631_;
  wire _9632_;
  wire _9633_;
  wire _9634_;
  wire _9635_;
  wire _9636_;
  wire _9637_;
  wire _9638_;
  wire _9639_;
  wire _9640_;
  wire _9641_;
  wire _9642_;
  wire _9643_;
  wire _9644_;
  wire _9645_;
  wire _9646_;
  wire _9647_;
  wire _9648_;
  wire _9649_;
  wire _9650_;
  wire _9651_;
  wire _9652_;
  wire _9653_;
  wire _9654_;
  wire _9655_;
  wire _9656_;
  wire _9657_;
  wire _9658_;
  wire _9659_;
  wire _9660_;
  wire _9661_;
  wire _9662_;
  wire _9663_;
  wire _9664_;
  wire _9665_;
  wire _9666_;
  wire _9667_;
  wire _9668_;
  wire _9669_;
  wire _9670_;
  wire _9671_;
  wire _9672_;
  wire _9673_;
  wire _9674_;
  wire _9675_;
  wire _9676_;
  wire _9677_;
  wire _9678_;
  wire _9679_;
  wire _9680_;
  wire _9681_;
  wire _9682_;
  wire _9683_;
  wire _9684_;
  wire _9685_;
  wire _9686_;
  wire _9687_;
  wire _9688_;
  wire _9689_;
  wire _9690_;
  wire _9691_;
  wire _9692_;
  wire _9693_;
  wire _9694_;
  wire _9695_;
  wire _9696_;
  wire _9697_;
  wire _9698_;
  wire _9699_;
  wire _9700_;
  wire _9701_;
  wire _9702_;
  wire _9703_;
  wire _9704_;
  wire _9705_;
  wire _9706_;
  wire _9707_;
  wire _9708_;
  wire _9709_;
  wire _9710_;
  wire _9711_;
  wire _9712_;
  wire _9713_;
  wire _9714_;
  wire _9715_;
  wire _9716_;
  wire _9717_;
  wire _9718_;
  wire _9719_;
  wire _9720_;
  wire _9721_;
  wire _9722_;
  wire _9723_;
  wire _9724_;
  wire _9725_;
  wire _9726_;
  wire _9727_;
  wire _9728_;
  wire _9729_;
  wire _9730_;
  wire _9731_;
  wire _9732_;
  wire _9733_;
  wire _9734_;
  wire _9735_;
  wire _9736_;
  wire _9737_;
  wire _9738_;
  wire _9739_;
  wire _9740_;
  wire _9741_;
  wire _9742_;
  wire _9743_;
  wire _9744_;
  wire _9745_;
  wire _9746_;
  wire _9747_;
  wire _9748_;
  wire _9749_;
  wire _9750_;
  wire _9751_;
  wire _9752_;
  wire _9753_;
  wire _9754_;
  wire _9755_;
  wire _9756_;
  wire _9757_;
  wire _9758_;
  wire _9759_;
  wire _9760_;
  wire _9761_;
  wire _9762_;
  wire _9763_;
  wire _9764_;
  wire _9765_;
  wire _9766_;
  wire _9767_;
  wire _9768_;
  wire _9769_;
  wire _9770_;
  wire _9771_;
  wire _9772_;
  wire _9773_;
  wire _9774_;
  wire _9775_;
  wire _9776_;
  wire _9777_;
  wire _9778_;
  wire _9779_;
  wire _9780_;
  wire _9781_;
  wire _9782_;
  wire _9783_;
  wire _9784_;
  wire _9785_;
  wire _9786_;
  wire _9787_;
  wire _9788_;
  wire _9789_;
  wire _9790_;
  wire _9791_;
  wire _9792_;
  wire _9793_;
  wire _9794_;
  wire _9795_;
  wire _9796_;
  wire _9797_;
  wire _9798_;
  wire _9799_;
  wire _9800_;
  wire _9801_;
  wire _9802_;
  wire _9803_;
  wire _9804_;
  wire _9805_;
  wire _9806_;
  wire _9807_;
  wire _9808_;
  wire _9809_;
  wire _9810_;
  wire _9811_;
  wire _9812_;
  wire _9813_;
  wire _9814_;
  wire _9815_;
  wire _9816_;
  wire _9817_;
  wire _9818_;
  wire _9819_;
  wire _9820_;
  wire _9821_;
  wire _9822_;
  wire _9823_;
  wire _9824_;
  wire _9825_;
  wire _9826_;
  wire _9827_;
  wire _9828_;
  wire _9829_;
  wire _9830_;
  wire _9831_;
  wire _9832_;
  wire _9833_;
  wire _9834_;
  wire _9835_;
  wire _9836_;
  wire _9837_;
  wire _9838_;
  wire _9839_;
  wire _9840_;
  wire _9841_;
  wire _9842_;
  wire _9843_;
  wire _9844_;
  wire _9845_;
  wire _9846_;
  wire _9847_;
  wire _9848_;
  wire _9849_;
  wire _9850_;
  wire _9851_;
  wire _9852_;
  wire _9853_;
  wire _9854_;
  wire _9855_;
  wire _9856_;
  wire _9857_;
  wire _9858_;
  wire _9859_;
  wire _9860_;
  wire _9861_;
  wire _9862_;
  wire _9863_;
  wire _9864_;
  wire _9865_;
  wire _9866_;
  wire _9867_;
  wire _9868_;
  wire _9869_;
  wire _9870_;
  wire _9871_;
  wire _9872_;
  wire _9873_;
  wire _9874_;
  wire _9875_;
  wire _9876_;
  wire _9877_;
  wire _9878_;
  wire _9879_;
  wire _9880_;
  wire _9881_;
  wire _9882_;
  wire _9883_;
  wire _9884_;
  wire _9885_;
  wire _9886_;
  wire _9887_;
  wire _9888_;
  wire _9889_;
  wire _9890_;
  wire _9891_;
  wire _9892_;
  wire _9893_;
  wire _9894_;
  wire _9895_;
  wire _9896_;
  wire _9897_;
  wire _9898_;
  wire _9899_;
  wire _9900_;
  wire _9901_;
  wire _9902_;
  wire _9903_;
  wire _9904_;
  wire _9905_;
  wire _9906_;
  wire _9907_;
  wire _9908_;
  wire _9909_;
  wire _9910_;
  wire _9911_;
  wire _9912_;
  wire _9913_;
  wire _9914_;
  wire _9915_;
  wire _9916_;
  wire _9917_;
  wire _9918_;
  wire _9919_;
  wire _9920_;
  wire _9921_;
  wire _9922_;
  wire _9923_;
  wire _9924_;
  wire _9925_;
  wire _9926_;
  wire _9927_;
  wire _9928_;
  wire _9929_;
  wire _9930_;
  wire _9931_;
  wire _9932_;
  wire _9933_;
  wire _9934_;
  wire _9935_;
  wire _9936_;
  wire _9937_;
  wire _9938_;
  wire _9939_;
  wire _9940_;
  wire _9941_;
  wire _9942_;
  wire _9943_;
  wire _9944_;
  wire _9945_;
  wire _9946_;
  wire _9947_;
  wire _9948_;
  wire _9949_;
  wire _9950_;
  wire _9951_;
  wire _9952_;
  wire _9953_;
  wire _9954_;
  wire _9955_;
  wire _9956_;
  wire _9957_;
  wire _9958_;
  wire _9959_;
  wire _9960_;
  wire _9961_;
  wire _9962_;
  wire _9963_;
  wire _9964_;
  wire _9965_;
  wire _9966_;
  wire _9967_;
  wire _9968_;
  wire _9969_;
  wire _9970_;
  wire _9971_;
  wire _9972_;
  wire _9973_;
  wire _9974_;
  wire _9975_;
  wire _9976_;
  wire _9977_;
  wire _9978_;
  wire _9979_;
  wire _9980_;
  wire _9981_;
  wire _9982_;
  wire _9983_;
  wire _9984_;
  wire _9985_;
  wire _9986_;
  wire _9987_;
  wire _9988_;
  wire _9989_;
  wire _9990_;
  wire _9991_;
  wire _9992_;
  wire _9993_;
  wire _9994_;
  wire _9995_;
  wire _9996_;
  wire _9997_;
  wire _9998_;
  wire _9999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire [62:0] r_0;
  wire [63:0] r_1;
  wire [63:0] m_1;
  wire [63:0] sum_1;
  wire [62:0] inv_1;
  wire [64:0] r_2;
  wire [64:0] m_2;
  wire [64:0] sum_2;
  wire [63:0] inv_2;
  wire [65:0] r_3;
  wire [65:0] m_3;
  wire [65:0] sum_3;
  wire [64:0] inv_3;
  wire [66:0] r_4;
  wire [66:0] m_4;
  wire [66:0] sum_4;
  wire [65:0] inv_4;
  wire [67:0] r_5;
  wire [67:0] m_5;
  wire [67:0] sum_5;
  wire [66:0] inv_5;
  wire [68:0] r_6;
  wire [68:0] m_6;
  wire [68:0] sum_6;
  wire [67:0] inv_6;
  wire [69:0] r_7;
  wire [69:0] m_7;
  wire [69:0] sum_7;
  wire [68:0] inv_7;
  wire [70:0] r_8;
  wire [70:0] m_8;
  wire [70:0] sum_8;
  wire [69:0] inv_8;
  wire [71:0] r_9;
  wire [71:0] m_9;
  wire [71:0] sum_9;
  wire [70:0] inv_9;
  wire [72:0] r_10;
  wire [72:0] m_10;
  wire [72:0] sum_10;
  wire [71:0] inv_10;
  wire [73:0] r_11;
  wire [73:0] m_11;
  wire [73:0] sum_11;
  wire [72:0] inv_11;
  wire [74:0] r_12;
  wire [74:0] m_12;
  wire [74:0] sum_12;
  wire [73:0] inv_12;
  wire [75:0] r_13;
  wire [75:0] m_13;
  wire [75:0] sum_13;
  wire [74:0] inv_13;
  wire [76:0] r_14;
  wire [76:0] m_14;
  wire [76:0] sum_14;
  wire [75:0] inv_14;
  wire [77:0] r_15;
  wire [77:0] m_15;
  wire [77:0] sum_15;
  wire [76:0] inv_15;
  wire [78:0] r_16;
  wire [78:0] m_16;
  wire [78:0] sum_16;
  wire [77:0] inv_16;
  wire [79:0] r_17;
  wire [79:0] m_17;
  wire [79:0] sum_17;
  wire [78:0] inv_17;
  wire [80:0] r_18;
  wire [80:0] m_18;
  wire [80:0] sum_18;
  wire [79:0] inv_18;
  wire [81:0] r_19;
  wire [81:0] m_19;
  wire [81:0] sum_19;
  wire [80:0] inv_19;
  wire [82:0] r_20;
  wire [82:0] m_20;
  wire [82:0] sum_20;
  wire [81:0] inv_20;
  wire [83:0] r_21;
  wire [83:0] m_21;
  wire [83:0] sum_21;
  wire [82:0] inv_21;
  wire [84:0] r_22;
  wire [84:0] m_22;
  wire [84:0] sum_22;
  wire [83:0] inv_22;
  wire [85:0] r_23;
  wire [85:0] m_23;
  wire [85:0] sum_23;
  wire [84:0] inv_23;
  wire [86:0] r_24;
  wire [86:0] m_24;
  wire [86:0] sum_24;
  wire [85:0] inv_24;
  wire [87:0] r_25;
  wire [87:0] m_25;
  wire [87:0] sum_25;
  wire [86:0] inv_25;
  wire [88:0] r_26;
  wire [88:0] m_26;
  wire [88:0] sum_26;
  wire [87:0] inv_26;
  wire [89:0] r_27;
  wire [89:0] m_27;
  wire [89:0] sum_27;
  wire [88:0] inv_27;
  wire [90:0] r_28;
  wire [90:0] m_28;
  wire [90:0] sum_28;
  wire [89:0] inv_28;
  wire [91:0] r_29;
  wire [91:0] m_29;
  wire [91:0] sum_29;
  wire [90:0] inv_29;
  wire [92:0] r_30;
  wire [92:0] m_30;
  wire [92:0] sum_30;
  wire [91:0] inv_30;
  wire [93:0] r_31;
  wire [93:0] m_31;
  wire [93:0] sum_31;
  wire [92:0] inv_31;
  wire [94:0] r_32;
  wire [94:0] m_32;
  wire [94:0] sum_32;
  wire [93:0] inv_32;
  wire zeroWire;
  wire oneWire;
  input [61:0] rin;
  input [30:0] div;
  output [31:0] q;
  output [94:0] rout;
  assign zeroWire = 1'b0 /*0*/;
  assign oneWire = 1'b1 /*0*/;
  assign r_0[0] = rin[0] /*35744*/;
  assign r_0[1] = rin[1] /*35743*/;
  assign r_0[2] = rin[2] /*35742*/;
  assign r_0[3] = rin[3] /*35741*/;
  assign r_0[4] = rin[4] /*35740*/;
  assign r_0[5] = rin[5] /*35739*/;
  assign r_0[6] = rin[6] /*35738*/;
  assign r_0[7] = rin[7] /*35737*/;
  assign r_0[8] = rin[8] /*35736*/;
  assign r_0[9] = rin[9] /*35735*/;
  assign r_0[10] = rin[10] /*35734*/;
  assign r_0[11] = rin[11] /*35733*/;
  assign r_0[12] = rin[12] /*35732*/;
  assign r_0[13] = rin[13] /*35731*/;
  assign r_0[14] = rin[14] /*35730*/;
  assign r_0[15] = rin[15] /*35729*/;
  assign r_0[16] = rin[16] /*35728*/;
  assign r_0[17] = rin[17] /*35727*/;
  assign r_0[18] = rin[18] /*35726*/;
  assign r_0[19] = rin[19] /*35725*/;
  assign r_0[20] = rin[20] /*35724*/;
  assign r_0[21] = rin[21] /*35723*/;
  assign r_0[22] = rin[22] /*35722*/;
  assign r_0[23] = rin[23] /*35721*/;
  assign r_0[24] = rin[24] /*35720*/;
  assign r_0[25] = rin[25] /*35719*/;
  assign r_0[26] = rin[26] /*35718*/;
  assign r_0[27] = rin[27] /*35717*/;
  assign r_0[28] = rin[28] /*35716*/;
  assign r_0[29] = rin[29] /*35715*/;
  assign r_0[30] = rin[30] /*35714*/;
  assign r_0[31] = rin[31] /*35713*/;
  assign r_0[32] = rin[32] /*35712*/;
  assign r_0[33] = rin[33] /*35711*/;
  assign r_0[34] = rin[34] /*35710*/;
  assign r_0[35] = rin[35] /*35709*/;
  assign r_0[36] = rin[36] /*35708*/;
  assign r_0[37] = rin[37] /*35707*/;
  assign r_0[38] = rin[38] /*35706*/;
  assign r_0[39] = rin[39] /*35705*/;
  assign r_0[40] = rin[40] /*35704*/;
  assign r_0[41] = rin[41] /*35703*/;
  assign r_0[42] = rin[42] /*35702*/;
  assign r_0[43] = rin[43] /*35701*/;
  assign r_0[44] = rin[44] /*35700*/;
  assign r_0[45] = rin[45] /*35699*/;
  assign r_0[46] = rin[46] /*35698*/;
  assign r_0[47] = rin[47] /*35697*/;
  assign r_0[48] = rin[48] /*35696*/;
  assign r_0[49] = rin[49] /*35695*/;
  assign r_0[50] = rin[50] /*35694*/;
  assign r_0[51] = rin[51] /*35693*/;
  assign r_0[52] = rin[52] /*35692*/;
  assign r_0[53] = rin[53] /*35691*/;
  assign r_0[54] = rin[54] /*35690*/;
  assign r_0[55] = rin[55] /*35689*/;
  assign r_0[56] = rin[56] /*35688*/;
  assign r_0[57] = rin[57] /*35687*/;
  assign r_0[58] = rin[58] /*35686*/;
  assign r_0[59] = rin[59] /*35685*/;
  assign r_0[60] = rin[60] /*35684*/;
  assign r_0[61] = rin[61] /*35683*/;
  assign r_0[62] = zeroWire /*35682*/;
  assign inv_1[0] = oneWire /*34496*/;
  assign inv_1[1] = oneWire /*34490*/;
  assign inv_1[2] = oneWire /*34484*/;
  assign inv_1[3] = oneWire /*34478*/;
  assign inv_1[4] = oneWire /*34472*/;
  assign inv_1[5] = oneWire /*34466*/;
  assign inv_1[6] = oneWire /*34460*/;
  assign inv_1[7] = oneWire /*34454*/;
  assign inv_1[8] = oneWire /*34448*/;
  assign inv_1[9] = oneWire /*34442*/;
  assign inv_1[10] = oneWire /*34436*/;
  assign inv_1[11] = oneWire /*34430*/;
  assign inv_1[12] = oneWire /*34424*/;
  assign inv_1[13] = oneWire /*34418*/;
  assign inv_1[14] = oneWire /*34412*/;
  assign inv_1[15] = oneWire /*34406*/;
  assign inv_1[16] = oneWire /*34400*/;
  assign inv_1[17] = oneWire /*34394*/;
  assign inv_1[18] = oneWire /*34388*/;
  assign inv_1[19] = oneWire /*34382*/;
  assign inv_1[20] = oneWire /*34376*/;
  assign inv_1[21] = oneWire /*34370*/;
  assign inv_1[22] = oneWire /*34364*/;
  assign inv_1[23] = oneWire /*34358*/;
  assign inv_1[24] = oneWire /*34352*/;
  assign inv_1[25] = oneWire /*34346*/;
  assign inv_1[26] = oneWire /*34340*/;
  assign inv_1[27] = oneWire /*34334*/;
  assign inv_1[28] = oneWire /*34328*/;
  assign inv_1[29] = oneWire /*34322*/;
  assign inv_1[30] = oneWire /*34316*/;
  assign inv_1[31] = ~div[0] /*34310*/;
  assign inv_1[32] = ~div[1] /*34304*/;
  assign inv_1[33] = ~div[2] /*34298*/;
  assign inv_1[34] = ~div[3] /*34292*/;
  assign inv_1[35] = ~div[4] /*34286*/;
  assign inv_1[36] = ~div[5] /*34280*/;
  assign inv_1[37] = ~div[6] /*34274*/;
  assign inv_1[38] = ~div[7] /*34268*/;
  assign inv_1[39] = ~div[8] /*34262*/;
  assign inv_1[40] = ~div[9] /*34256*/;
  assign inv_1[41] = ~div[10] /*34250*/;
  assign inv_1[42] = ~div[11] /*34244*/;
  assign inv_1[43] = ~div[12] /*34238*/;
  assign inv_1[44] = ~div[13] /*34232*/;
  assign inv_1[45] = ~div[14] /*34226*/;
  assign inv_1[46] = ~div[15] /*34220*/;
  assign inv_1[47] = ~div[16] /*34214*/;
  assign inv_1[48] = ~div[17] /*34208*/;
  assign inv_1[49] = ~div[18] /*34202*/;
  assign inv_1[50] = ~div[19] /*34196*/;
  assign inv_1[51] = ~div[20] /*34190*/;
  assign inv_1[52] = ~div[21] /*34184*/;
  assign inv_1[53] = ~div[22] /*34178*/;
  assign inv_1[54] = ~div[23] /*34172*/;
  assign inv_1[55] = ~div[24] /*34166*/;
  assign inv_1[56] = ~div[25] /*34160*/;
  assign inv_1[57] = ~div[26] /*34154*/;
  assign inv_1[58] = ~div[27] /*34148*/;
  assign inv_1[59] = ~div[28] /*34142*/;
  assign inv_1[60] = ~div[29] /*34136*/;
  assign inv_1[61] = ~div[30] /*34130*/;
  assign inv_1[62] = oneWire /*34124*/;
  assign _0_ = inv_1[0] ^ r_0[0] /*34495*/;
  assign sum_1[0] = _0_ ^ oneWire /*34494*/;
  assign _1_ = _0_ & oneWire /*34493*/;
  assign _2_ = inv_1[0] & r_0[0] /*34492*/;
  assign _3_ = _1_ | _2_ /*34491*/;
  assign _4_ = inv_1[1] ^ r_0[1] /*34489*/;
  assign sum_1[1] = _4_ ^ _3_ /*34488*/;
  assign _5_ = _4_ & _3_ /*34487*/;
  assign _6_ = inv_1[1] & r_0[1] /*34486*/;
  assign _7_ = _5_ | _6_ /*34485*/;
  assign _8_ = inv_1[2] ^ r_0[2] /*34483*/;
  assign sum_1[2] = _8_ ^ _7_ /*34482*/;
  assign _9_ = _8_ & _7_ /*34481*/;
  assign _10_ = inv_1[2] & r_0[2] /*34480*/;
  assign _11_ = _9_ | _10_ /*34479*/;
  assign _12_ = inv_1[3] ^ r_0[3] /*34477*/;
  assign sum_1[3] = _12_ ^ _11_ /*34476*/;
  assign _13_ = _12_ & _11_ /*34475*/;
  assign _14_ = inv_1[3] & r_0[3] /*34474*/;
  assign _15_ = _13_ | _14_ /*34473*/;
  assign _16_ = inv_1[4] ^ r_0[4] /*34471*/;
  assign sum_1[4] = _16_ ^ _15_ /*34470*/;
  assign _17_ = _16_ & _15_ /*34469*/;
  assign _18_ = inv_1[4] & r_0[4] /*34468*/;
  assign _19_ = _17_ | _18_ /*34467*/;
  assign _20_ = inv_1[5] ^ r_0[5] /*34465*/;
  assign sum_1[5] = _20_ ^ _19_ /*34464*/;
  assign _21_ = _20_ & _19_ /*34463*/;
  assign _22_ = inv_1[5] & r_0[5] /*34462*/;
  assign _23_ = _21_ | _22_ /*34461*/;
  assign _24_ = inv_1[6] ^ r_0[6] /*34459*/;
  assign sum_1[6] = _24_ ^ _23_ /*34458*/;
  assign _25_ = _24_ & _23_ /*34457*/;
  assign _26_ = inv_1[6] & r_0[6] /*34456*/;
  assign _27_ = _25_ | _26_ /*34455*/;
  assign _28_ = inv_1[7] ^ r_0[7] /*34453*/;
  assign sum_1[7] = _28_ ^ _27_ /*34452*/;
  assign _29_ = _28_ & _27_ /*34451*/;
  assign _30_ = inv_1[7] & r_0[7] /*34450*/;
  assign _31_ = _29_ | _30_ /*34449*/;
  assign _32_ = inv_1[8] ^ r_0[8] /*34447*/;
  assign sum_1[8] = _32_ ^ _31_ /*34446*/;
  assign _33_ = _32_ & _31_ /*34445*/;
  assign _34_ = inv_1[8] & r_0[8] /*34444*/;
  assign _35_ = _33_ | _34_ /*34443*/;
  assign _36_ = inv_1[9] ^ r_0[9] /*34441*/;
  assign sum_1[9] = _36_ ^ _35_ /*34440*/;
  assign _37_ = _36_ & _35_ /*34439*/;
  assign _38_ = inv_1[9] & r_0[9] /*34438*/;
  assign _39_ = _37_ | _38_ /*34437*/;
  assign _40_ = inv_1[10] ^ r_0[10] /*34435*/;
  assign sum_1[10] = _40_ ^ _39_ /*34434*/;
  assign _41_ = _40_ & _39_ /*34433*/;
  assign _42_ = inv_1[10] & r_0[10] /*34432*/;
  assign _43_ = _41_ | _42_ /*34431*/;
  assign _44_ = inv_1[11] ^ r_0[11] /*34429*/;
  assign sum_1[11] = _44_ ^ _43_ /*34428*/;
  assign _45_ = _44_ & _43_ /*34427*/;
  assign _46_ = inv_1[11] & r_0[11] /*34426*/;
  assign _47_ = _45_ | _46_ /*34425*/;
  assign _48_ = inv_1[12] ^ r_0[12] /*34423*/;
  assign sum_1[12] = _48_ ^ _47_ /*34422*/;
  assign _49_ = _48_ & _47_ /*34421*/;
  assign _50_ = inv_1[12] & r_0[12] /*34420*/;
  assign _51_ = _49_ | _50_ /*34419*/;
  assign _52_ = inv_1[13] ^ r_0[13] /*34417*/;
  assign sum_1[13] = _52_ ^ _51_ /*34416*/;
  assign _53_ = _52_ & _51_ /*34415*/;
  assign _54_ = inv_1[13] & r_0[13] /*34414*/;
  assign _55_ = _53_ | _54_ /*34413*/;
  assign _56_ = inv_1[14] ^ r_0[14] /*34411*/;
  assign sum_1[14] = _56_ ^ _55_ /*34410*/;
  assign _57_ = _56_ & _55_ /*34409*/;
  assign _58_ = inv_1[14] & r_0[14] /*34408*/;
  assign _59_ = _57_ | _58_ /*34407*/;
  assign _60_ = inv_1[15] ^ r_0[15] /*34405*/;
  assign sum_1[15] = _60_ ^ _59_ /*34404*/;
  assign _61_ = _60_ & _59_ /*34403*/;
  assign _62_ = inv_1[15] & r_0[15] /*34402*/;
  assign _63_ = _61_ | _62_ /*34401*/;
  assign _64_ = inv_1[16] ^ r_0[16] /*34399*/;
  assign sum_1[16] = _64_ ^ _63_ /*34398*/;
  assign _65_ = _64_ & _63_ /*34397*/;
  assign _66_ = inv_1[16] & r_0[16] /*34396*/;
  assign _67_ = _65_ | _66_ /*34395*/;
  assign _68_ = inv_1[17] ^ r_0[17] /*34393*/;
  assign sum_1[17] = _68_ ^ _67_ /*34392*/;
  assign _69_ = _68_ & _67_ /*34391*/;
  assign _70_ = inv_1[17] & r_0[17] /*34390*/;
  assign _71_ = _69_ | _70_ /*34389*/;
  assign _72_ = inv_1[18] ^ r_0[18] /*34387*/;
  assign sum_1[18] = _72_ ^ _71_ /*34386*/;
  assign _73_ = _72_ & _71_ /*34385*/;
  assign _74_ = inv_1[18] & r_0[18] /*34384*/;
  assign _75_ = _73_ | _74_ /*34383*/;
  assign _76_ = inv_1[19] ^ r_0[19] /*34381*/;
  assign sum_1[19] = _76_ ^ _75_ /*34380*/;
  assign _77_ = _76_ & _75_ /*34379*/;
  assign _78_ = inv_1[19] & r_0[19] /*34378*/;
  assign _79_ = _77_ | _78_ /*34377*/;
  assign _80_ = inv_1[20] ^ r_0[20] /*34375*/;
  assign sum_1[20] = _80_ ^ _79_ /*34374*/;
  assign _81_ = _80_ & _79_ /*34373*/;
  assign _82_ = inv_1[20] & r_0[20] /*34372*/;
  assign _83_ = _81_ | _82_ /*34371*/;
  assign _84_ = inv_1[21] ^ r_0[21] /*34369*/;
  assign sum_1[21] = _84_ ^ _83_ /*34368*/;
  assign _85_ = _84_ & _83_ /*34367*/;
  assign _86_ = inv_1[21] & r_0[21] /*34366*/;
  assign _87_ = _85_ | _86_ /*34365*/;
  assign _88_ = inv_1[22] ^ r_0[22] /*34363*/;
  assign sum_1[22] = _88_ ^ _87_ /*34362*/;
  assign _89_ = _88_ & _87_ /*34361*/;
  assign _90_ = inv_1[22] & r_0[22] /*34360*/;
  assign _91_ = _89_ | _90_ /*34359*/;
  assign _92_ = inv_1[23] ^ r_0[23] /*34357*/;
  assign sum_1[23] = _92_ ^ _91_ /*34356*/;
  assign _93_ = _92_ & _91_ /*34355*/;
  assign _94_ = inv_1[23] & r_0[23] /*34354*/;
  assign _95_ = _93_ | _94_ /*34353*/;
  assign _96_ = inv_1[24] ^ r_0[24] /*34351*/;
  assign sum_1[24] = _96_ ^ _95_ /*34350*/;
  assign _97_ = _96_ & _95_ /*34349*/;
  assign _98_ = inv_1[24] & r_0[24] /*34348*/;
  assign _99_ = _97_ | _98_ /*34347*/;
  assign _100_ = inv_1[25] ^ r_0[25] /*34345*/;
  assign sum_1[25] = _100_ ^ _99_ /*34344*/;
  assign _101_ = _100_ & _99_ /*34343*/;
  assign _102_ = inv_1[25] & r_0[25] /*34342*/;
  assign _103_ = _101_ | _102_ /*34341*/;
  assign _104_ = inv_1[26] ^ r_0[26] /*34339*/;
  assign sum_1[26] = _104_ ^ _103_ /*34338*/;
  assign _105_ = _104_ & _103_ /*34337*/;
  assign _106_ = inv_1[26] & r_0[26] /*34336*/;
  assign _107_ = _105_ | _106_ /*34335*/;
  assign _108_ = inv_1[27] ^ r_0[27] /*34333*/;
  assign sum_1[27] = _108_ ^ _107_ /*34332*/;
  assign _109_ = _108_ & _107_ /*34331*/;
  assign _110_ = inv_1[27] & r_0[27] /*34330*/;
  assign _111_ = _109_ | _110_ /*34329*/;
  assign _112_ = inv_1[28] ^ r_0[28] /*34327*/;
  assign sum_1[28] = _112_ ^ _111_ /*34326*/;
  assign _113_ = _112_ & _111_ /*34325*/;
  assign _114_ = inv_1[28] & r_0[28] /*34324*/;
  assign _115_ = _113_ | _114_ /*34323*/;
  assign _116_ = inv_1[29] ^ r_0[29] /*34321*/;
  assign sum_1[29] = _116_ ^ _115_ /*34320*/;
  assign _117_ = _116_ & _115_ /*34319*/;
  assign _118_ = inv_1[29] & r_0[29] /*34318*/;
  assign _119_ = _117_ | _118_ /*34317*/;
  assign _120_ = inv_1[30] ^ r_0[30] /*34315*/;
  assign sum_1[30] = _120_ ^ _119_ /*34314*/;
  assign _121_ = _120_ & _119_ /*34313*/;
  assign _122_ = inv_1[30] & r_0[30] /*34312*/;
  assign _123_ = _121_ | _122_ /*34311*/;
  assign _124_ = inv_1[31] ^ r_0[31] /*34309*/;
  assign sum_1[31] = _124_ ^ _123_ /*34308*/;
  assign _125_ = _124_ & _123_ /*34307*/;
  assign _126_ = inv_1[31] & r_0[31] /*34306*/;
  assign _127_ = _125_ | _126_ /*34305*/;
  assign _128_ = inv_1[32] ^ r_0[32] /*34303*/;
  assign sum_1[32] = _128_ ^ _127_ /*34302*/;
  assign _129_ = _128_ & _127_ /*34301*/;
  assign _130_ = inv_1[32] & r_0[32] /*34300*/;
  assign _131_ = _129_ | _130_ /*34299*/;
  assign _132_ = inv_1[33] ^ r_0[33] /*34297*/;
  assign sum_1[33] = _132_ ^ _131_ /*34296*/;
  assign _133_ = _132_ & _131_ /*34295*/;
  assign _134_ = inv_1[33] & r_0[33] /*34294*/;
  assign _135_ = _133_ | _134_ /*34293*/;
  assign _136_ = inv_1[34] ^ r_0[34] /*34291*/;
  assign sum_1[34] = _136_ ^ _135_ /*34290*/;
  assign _137_ = _136_ & _135_ /*34289*/;
  assign _138_ = inv_1[34] & r_0[34] /*34288*/;
  assign _139_ = _137_ | _138_ /*34287*/;
  assign _140_ = inv_1[35] ^ r_0[35] /*34285*/;
  assign sum_1[35] = _140_ ^ _139_ /*34284*/;
  assign _141_ = _140_ & _139_ /*34283*/;
  assign _142_ = inv_1[35] & r_0[35] /*34282*/;
  assign _143_ = _141_ | _142_ /*34281*/;
  assign _144_ = inv_1[36] ^ r_0[36] /*34279*/;
  assign sum_1[36] = _144_ ^ _143_ /*34278*/;
  assign _145_ = _144_ & _143_ /*34277*/;
  assign _146_ = inv_1[36] & r_0[36] /*34276*/;
  assign _147_ = _145_ | _146_ /*34275*/;
  assign _148_ = inv_1[37] ^ r_0[37] /*34273*/;
  assign sum_1[37] = _148_ ^ _147_ /*34272*/;
  assign _149_ = _148_ & _147_ /*34271*/;
  assign _150_ = inv_1[37] & r_0[37] /*34270*/;
  assign _151_ = _149_ | _150_ /*34269*/;
  assign _152_ = inv_1[38] ^ r_0[38] /*34267*/;
  assign sum_1[38] = _152_ ^ _151_ /*34266*/;
  assign _153_ = _152_ & _151_ /*34265*/;
  assign _154_ = inv_1[38] & r_0[38] /*34264*/;
  assign _155_ = _153_ | _154_ /*34263*/;
  assign _156_ = inv_1[39] ^ r_0[39] /*34261*/;
  assign sum_1[39] = _156_ ^ _155_ /*34260*/;
  assign _157_ = _156_ & _155_ /*34259*/;
  assign _158_ = inv_1[39] & r_0[39] /*34258*/;
  assign _159_ = _157_ | _158_ /*34257*/;
  assign _160_ = inv_1[40] ^ r_0[40] /*34255*/;
  assign sum_1[40] = _160_ ^ _159_ /*34254*/;
  assign _161_ = _160_ & _159_ /*34253*/;
  assign _162_ = inv_1[40] & r_0[40] /*34252*/;
  assign _163_ = _161_ | _162_ /*34251*/;
  assign _164_ = inv_1[41] ^ r_0[41] /*34249*/;
  assign sum_1[41] = _164_ ^ _163_ /*34248*/;
  assign _165_ = _164_ & _163_ /*34247*/;
  assign _166_ = inv_1[41] & r_0[41] /*34246*/;
  assign _167_ = _165_ | _166_ /*34245*/;
  assign _168_ = inv_1[42] ^ r_0[42] /*34243*/;
  assign sum_1[42] = _168_ ^ _167_ /*34242*/;
  assign _169_ = _168_ & _167_ /*34241*/;
  assign _170_ = inv_1[42] & r_0[42] /*34240*/;
  assign _171_ = _169_ | _170_ /*34239*/;
  assign _172_ = inv_1[43] ^ r_0[43] /*34237*/;
  assign sum_1[43] = _172_ ^ _171_ /*34236*/;
  assign _173_ = _172_ & _171_ /*34235*/;
  assign _174_ = inv_1[43] & r_0[43] /*34234*/;
  assign _175_ = _173_ | _174_ /*34233*/;
  assign _176_ = inv_1[44] ^ r_0[44] /*34231*/;
  assign sum_1[44] = _176_ ^ _175_ /*34230*/;
  assign _177_ = _176_ & _175_ /*34229*/;
  assign _178_ = inv_1[44] & r_0[44] /*34228*/;
  assign _179_ = _177_ | _178_ /*34227*/;
  assign _180_ = inv_1[45] ^ r_0[45] /*34225*/;
  assign sum_1[45] = _180_ ^ _179_ /*34224*/;
  assign _181_ = _180_ & _179_ /*34223*/;
  assign _182_ = inv_1[45] & r_0[45] /*34222*/;
  assign _183_ = _181_ | _182_ /*34221*/;
  assign _184_ = inv_1[46] ^ r_0[46] /*34219*/;
  assign sum_1[46] = _184_ ^ _183_ /*34218*/;
  assign _185_ = _184_ & _183_ /*34217*/;
  assign _186_ = inv_1[46] & r_0[46] /*34216*/;
  assign _187_ = _185_ | _186_ /*34215*/;
  assign _188_ = inv_1[47] ^ r_0[47] /*34213*/;
  assign sum_1[47] = _188_ ^ _187_ /*34212*/;
  assign _189_ = _188_ & _187_ /*34211*/;
  assign _190_ = inv_1[47] & r_0[47] /*34210*/;
  assign _191_ = _189_ | _190_ /*34209*/;
  assign _192_ = inv_1[48] ^ r_0[48] /*34207*/;
  assign sum_1[48] = _192_ ^ _191_ /*34206*/;
  assign _193_ = _192_ & _191_ /*34205*/;
  assign _194_ = inv_1[48] & r_0[48] /*34204*/;
  assign _195_ = _193_ | _194_ /*34203*/;
  assign _196_ = inv_1[49] ^ r_0[49] /*34201*/;
  assign sum_1[49] = _196_ ^ _195_ /*34200*/;
  assign _197_ = _196_ & _195_ /*34199*/;
  assign _198_ = inv_1[49] & r_0[49] /*34198*/;
  assign _199_ = _197_ | _198_ /*34197*/;
  assign _200_ = inv_1[50] ^ r_0[50] /*34195*/;
  assign sum_1[50] = _200_ ^ _199_ /*34194*/;
  assign _201_ = _200_ & _199_ /*34193*/;
  assign _202_ = inv_1[50] & r_0[50] /*34192*/;
  assign _203_ = _201_ | _202_ /*34191*/;
  assign _204_ = inv_1[51] ^ r_0[51] /*34189*/;
  assign sum_1[51] = _204_ ^ _203_ /*34188*/;
  assign _205_ = _204_ & _203_ /*34187*/;
  assign _206_ = inv_1[51] & r_0[51] /*34186*/;
  assign _207_ = _205_ | _206_ /*34185*/;
  assign _208_ = inv_1[52] ^ r_0[52] /*34183*/;
  assign sum_1[52] = _208_ ^ _207_ /*34182*/;
  assign _209_ = _208_ & _207_ /*34181*/;
  assign _210_ = inv_1[52] & r_0[52] /*34180*/;
  assign _211_ = _209_ | _210_ /*34179*/;
  assign _212_ = inv_1[53] ^ r_0[53] /*34177*/;
  assign sum_1[53] = _212_ ^ _211_ /*34176*/;
  assign _213_ = _212_ & _211_ /*34175*/;
  assign _214_ = inv_1[53] & r_0[53] /*34174*/;
  assign _215_ = _213_ | _214_ /*34173*/;
  assign _216_ = inv_1[54] ^ r_0[54] /*34171*/;
  assign sum_1[54] = _216_ ^ _215_ /*34170*/;
  assign _217_ = _216_ & _215_ /*34169*/;
  assign _218_ = inv_1[54] & r_0[54] /*34168*/;
  assign _219_ = _217_ | _218_ /*34167*/;
  assign _220_ = inv_1[55] ^ r_0[55] /*34165*/;
  assign sum_1[55] = _220_ ^ _219_ /*34164*/;
  assign _221_ = _220_ & _219_ /*34163*/;
  assign _222_ = inv_1[55] & r_0[55] /*34162*/;
  assign _223_ = _221_ | _222_ /*34161*/;
  assign _224_ = inv_1[56] ^ r_0[56] /*34159*/;
  assign sum_1[56] = _224_ ^ _223_ /*34158*/;
  assign _225_ = _224_ & _223_ /*34157*/;
  assign _226_ = inv_1[56] & r_0[56] /*34156*/;
  assign _227_ = _225_ | _226_ /*34155*/;
  assign _228_ = inv_1[57] ^ r_0[57] /*34153*/;
  assign sum_1[57] = _228_ ^ _227_ /*34152*/;
  assign _229_ = _228_ & _227_ /*34151*/;
  assign _230_ = inv_1[57] & r_0[57] /*34150*/;
  assign _231_ = _229_ | _230_ /*34149*/;
  assign _232_ = inv_1[58] ^ r_0[58] /*34147*/;
  assign sum_1[58] = _232_ ^ _231_ /*34146*/;
  assign _233_ = _232_ & _231_ /*34145*/;
  assign _234_ = inv_1[58] & r_0[58] /*34144*/;
  assign _235_ = _233_ | _234_ /*34143*/;
  assign _236_ = inv_1[59] ^ r_0[59] /*34141*/;
  assign sum_1[59] = _236_ ^ _235_ /*34140*/;
  assign _237_ = _236_ & _235_ /*34139*/;
  assign _238_ = inv_1[59] & r_0[59] /*34138*/;
  assign _239_ = _237_ | _238_ /*34137*/;
  assign _240_ = inv_1[60] ^ r_0[60] /*34135*/;
  assign sum_1[60] = _240_ ^ _239_ /*34134*/;
  assign _241_ = _240_ & _239_ /*34133*/;
  assign _242_ = inv_1[60] & r_0[60] /*34132*/;
  assign _243_ = _241_ | _242_ /*34131*/;
  assign _244_ = inv_1[61] ^ r_0[61] /*34129*/;
  assign sum_1[61] = _244_ ^ _243_ /*34128*/;
  assign _245_ = _244_ & _243_ /*34127*/;
  assign _246_ = inv_1[61] & r_0[61] /*34126*/;
  assign _247_ = _245_ | _246_ /*34125*/;
  assign _248_ = inv_1[62] ^ r_0[62] /*34123*/;
  assign sum_1[62] = _248_ ^ _247_ /*34122*/;
  assign _249_ = _248_ & _247_ /*34121*/;
  assign _250_ = inv_1[62] & r_0[62] /*34120*/;
  assign _251_ = _249_ | _250_ /*34119*/;
  assign _252_ = _251_ ^ _247_ /*34118*/;
  assign _253_ = ~_252_ /*34117*/;
  assign _254_ = sum_1[62] & _253_ /*34116*/;
  assign _255_ = _252_ & _251_ /*34115*/;
  assign sum_1[63] = _255_ | _254_ /*34114*/;
  assign q[31] = ~sum_1[63] /*34113*/;
  assign m_1[0] = r_0[0] /*34112*/;
  assign m_1[1] = r_0[1] /*34111*/;
  assign m_1[2] = r_0[2] /*34110*/;
  assign m_1[3] = r_0[3] /*34109*/;
  assign m_1[4] = r_0[4] /*34108*/;
  assign m_1[5] = r_0[5] /*34107*/;
  assign m_1[6] = r_0[6] /*34106*/;
  assign m_1[7] = r_0[7] /*34105*/;
  assign m_1[8] = r_0[8] /*34104*/;
  assign m_1[9] = r_0[9] /*34103*/;
  assign m_1[10] = r_0[10] /*34102*/;
  assign m_1[11] = r_0[11] /*34101*/;
  assign m_1[12] = r_0[12] /*34100*/;
  assign m_1[13] = r_0[13] /*34099*/;
  assign m_1[14] = r_0[14] /*34098*/;
  assign m_1[15] = r_0[15] /*34097*/;
  assign m_1[16] = r_0[16] /*34096*/;
  assign m_1[17] = r_0[17] /*34095*/;
  assign m_1[18] = r_0[18] /*34094*/;
  assign m_1[19] = r_0[19] /*34093*/;
  assign m_1[20] = r_0[20] /*34092*/;
  assign m_1[21] = r_0[21] /*34091*/;
  assign m_1[22] = r_0[22] /*34090*/;
  assign m_1[23] = r_0[23] /*34089*/;
  assign m_1[24] = r_0[24] /*34088*/;
  assign m_1[25] = r_0[25] /*34087*/;
  assign m_1[26] = r_0[26] /*34086*/;
  assign m_1[27] = r_0[27] /*34085*/;
  assign m_1[28] = r_0[28] /*34084*/;
  assign m_1[29] = r_0[29] /*34083*/;
  assign m_1[30] = r_0[30] /*34082*/;
  assign m_1[31] = r_0[31] /*34081*/;
  assign m_1[32] = r_0[32] /*34080*/;
  assign m_1[33] = r_0[33] /*34079*/;
  assign m_1[34] = r_0[34] /*34078*/;
  assign m_1[35] = r_0[35] /*34077*/;
  assign m_1[36] = r_0[36] /*34076*/;
  assign m_1[37] = r_0[37] /*34075*/;
  assign m_1[38] = r_0[38] /*34074*/;
  assign m_1[39] = r_0[39] /*34073*/;
  assign m_1[40] = r_0[40] /*34072*/;
  assign m_1[41] = r_0[41] /*34071*/;
  assign m_1[42] = r_0[42] /*34070*/;
  assign m_1[43] = r_0[43] /*34069*/;
  assign m_1[44] = r_0[44] /*34068*/;
  assign m_1[45] = r_0[45] /*34067*/;
  assign m_1[46] = r_0[46] /*34066*/;
  assign m_1[47] = r_0[47] /*34065*/;
  assign m_1[48] = r_0[48] /*34064*/;
  assign m_1[49] = r_0[49] /*34063*/;
  assign m_1[50] = r_0[50] /*34062*/;
  assign m_1[51] = r_0[51] /*34061*/;
  assign m_1[52] = r_0[52] /*34060*/;
  assign m_1[53] = r_0[53] /*34059*/;
  assign m_1[54] = r_0[54] /*34058*/;
  assign m_1[55] = r_0[55] /*34057*/;
  assign m_1[56] = r_0[56] /*34056*/;
  assign m_1[57] = r_0[57] /*34055*/;
  assign m_1[58] = r_0[58] /*34054*/;
  assign m_1[59] = r_0[59] /*34053*/;
  assign m_1[60] = r_0[60] /*34052*/;
  assign m_1[61] = r_0[61] /*34051*/;
  assign m_1[62] = r_0[62] /*34050*/;
  assign m_1[63] = r_0[62] /*34049*/;
  assign _257_ = ~q[31] /*34048*/;
  assign _258_ = sum_1[0] & q[31] /*34047*/;
  assign _259_ = m_1[0] & _257_ /*34046*/;
  assign r_1[0] = _259_ | _258_ /*34045*/;
  assign _260_ = ~q[31] /*34044*/;
  assign _261_ = sum_1[1] & q[31] /*34043*/;
  assign _262_ = m_1[1] & _260_ /*34042*/;
  assign r_1[1] = _262_ | _261_ /*34041*/;
  assign _263_ = ~q[31] /*34040*/;
  assign _264_ = sum_1[2] & q[31] /*34039*/;
  assign _265_ = m_1[2] & _263_ /*34038*/;
  assign r_1[2] = _265_ | _264_ /*34037*/;
  assign _266_ = ~q[31] /*34036*/;
  assign _267_ = sum_1[3] & q[31] /*34035*/;
  assign _268_ = m_1[3] & _266_ /*34034*/;
  assign r_1[3] = _268_ | _267_ /*34033*/;
  assign _269_ = ~q[31] /*34032*/;
  assign _270_ = sum_1[4] & q[31] /*34031*/;
  assign _271_ = m_1[4] & _269_ /*34030*/;
  assign r_1[4] = _271_ | _270_ /*34029*/;
  assign _272_ = ~q[31] /*34028*/;
  assign _273_ = sum_1[5] & q[31] /*34027*/;
  assign _274_ = m_1[5] & _272_ /*34026*/;
  assign r_1[5] = _274_ | _273_ /*34025*/;
  assign _275_ = ~q[31] /*34024*/;
  assign _276_ = sum_1[6] & q[31] /*34023*/;
  assign _277_ = m_1[6] & _275_ /*34022*/;
  assign r_1[6] = _277_ | _276_ /*34021*/;
  assign _278_ = ~q[31] /*34020*/;
  assign _279_ = sum_1[7] & q[31] /*34019*/;
  assign _280_ = m_1[7] & _278_ /*34018*/;
  assign r_1[7] = _280_ | _279_ /*34017*/;
  assign _281_ = ~q[31] /*34016*/;
  assign _282_ = sum_1[8] & q[31] /*34015*/;
  assign _283_ = m_1[8] & _281_ /*34014*/;
  assign r_1[8] = _283_ | _282_ /*34013*/;
  assign _284_ = ~q[31] /*34012*/;
  assign _285_ = sum_1[9] & q[31] /*34011*/;
  assign _286_ = m_1[9] & _284_ /*34010*/;
  assign r_1[9] = _286_ | _285_ /*34009*/;
  assign _287_ = ~q[31] /*34008*/;
  assign _288_ = sum_1[10] & q[31] /*34007*/;
  assign _289_ = m_1[10] & _287_ /*34006*/;
  assign r_1[10] = _289_ | _288_ /*34005*/;
  assign _290_ = ~q[31] /*34004*/;
  assign _291_ = sum_1[11] & q[31] /*34003*/;
  assign _292_ = m_1[11] & _290_ /*34002*/;
  assign r_1[11] = _292_ | _291_ /*34001*/;
  assign _293_ = ~q[31] /*34000*/;
  assign _294_ = sum_1[12] & q[31] /*33999*/;
  assign _295_ = m_1[12] & _293_ /*33998*/;
  assign r_1[12] = _295_ | _294_ /*33997*/;
  assign _296_ = ~q[31] /*33996*/;
  assign _297_ = sum_1[13] & q[31] /*33995*/;
  assign _298_ = m_1[13] & _296_ /*33994*/;
  assign r_1[13] = _298_ | _297_ /*33993*/;
  assign _299_ = ~q[31] /*33992*/;
  assign _300_ = sum_1[14] & q[31] /*33991*/;
  assign _301_ = m_1[14] & _299_ /*33990*/;
  assign r_1[14] = _301_ | _300_ /*33989*/;
  assign _302_ = ~q[31] /*33988*/;
  assign _303_ = sum_1[15] & q[31] /*33987*/;
  assign _304_ = m_1[15] & _302_ /*33986*/;
  assign r_1[15] = _304_ | _303_ /*33985*/;
  assign _305_ = ~q[31] /*33984*/;
  assign _306_ = sum_1[16] & q[31] /*33983*/;
  assign _307_ = m_1[16] & _305_ /*33982*/;
  assign r_1[16] = _307_ | _306_ /*33981*/;
  assign _308_ = ~q[31] /*33980*/;
  assign _309_ = sum_1[17] & q[31] /*33979*/;
  assign _310_ = m_1[17] & _308_ /*33978*/;
  assign r_1[17] = _310_ | _309_ /*33977*/;
  assign _311_ = ~q[31] /*33976*/;
  assign _312_ = sum_1[18] & q[31] /*33975*/;
  assign _313_ = m_1[18] & _311_ /*33974*/;
  assign r_1[18] = _313_ | _312_ /*33973*/;
  assign _314_ = ~q[31] /*33972*/;
  assign _315_ = sum_1[19] & q[31] /*33971*/;
  assign _316_ = m_1[19] & _314_ /*33970*/;
  assign r_1[19] = _316_ | _315_ /*33969*/;
  assign _317_ = ~q[31] /*33968*/;
  assign _318_ = sum_1[20] & q[31] /*33967*/;
  assign _319_ = m_1[20] & _317_ /*33966*/;
  assign r_1[20] = _319_ | _318_ /*33965*/;
  assign _320_ = ~q[31] /*33964*/;
  assign _321_ = sum_1[21] & q[31] /*33963*/;
  assign _322_ = m_1[21] & _320_ /*33962*/;
  assign r_1[21] = _322_ | _321_ /*33961*/;
  assign _323_ = ~q[31] /*33960*/;
  assign _324_ = sum_1[22] & q[31] /*33959*/;
  assign _325_ = m_1[22] & _323_ /*33958*/;
  assign r_1[22] = _325_ | _324_ /*33957*/;
  assign _326_ = ~q[31] /*33956*/;
  assign _327_ = sum_1[23] & q[31] /*33955*/;
  assign _328_ = m_1[23] & _326_ /*33954*/;
  assign r_1[23] = _328_ | _327_ /*33953*/;
  assign _329_ = ~q[31] /*33952*/;
  assign _330_ = sum_1[24] & q[31] /*33951*/;
  assign _331_ = m_1[24] & _329_ /*33950*/;
  assign r_1[24] = _331_ | _330_ /*33949*/;
  assign _332_ = ~q[31] /*33948*/;
  assign _333_ = sum_1[25] & q[31] /*33947*/;
  assign _334_ = m_1[25] & _332_ /*33946*/;
  assign r_1[25] = _334_ | _333_ /*33945*/;
  assign _335_ = ~q[31] /*33944*/;
  assign _336_ = sum_1[26] & q[31] /*33943*/;
  assign _337_ = m_1[26] & _335_ /*33942*/;
  assign r_1[26] = _337_ | _336_ /*33941*/;
  assign _338_ = ~q[31] /*33940*/;
  assign _339_ = sum_1[27] & q[31] /*33939*/;
  assign _340_ = m_1[27] & _338_ /*33938*/;
  assign r_1[27] = _340_ | _339_ /*33937*/;
  assign _341_ = ~q[31] /*33936*/;
  assign _342_ = sum_1[28] & q[31] /*33935*/;
  assign _343_ = m_1[28] & _341_ /*33934*/;
  assign r_1[28] = _343_ | _342_ /*33933*/;
  assign _344_ = ~q[31] /*33932*/;
  assign _345_ = sum_1[29] & q[31] /*33931*/;
  assign _346_ = m_1[29] & _344_ /*33930*/;
  assign r_1[29] = _346_ | _345_ /*33929*/;
  assign _347_ = ~q[31] /*33928*/;
  assign _348_ = sum_1[30] & q[31] /*33927*/;
  assign _349_ = m_1[30] & _347_ /*33926*/;
  assign r_1[30] = _349_ | _348_ /*33925*/;
  assign _350_ = ~q[31] /*33924*/;
  assign _351_ = sum_1[31] & q[31] /*33923*/;
  assign _352_ = m_1[31] & _350_ /*33922*/;
  assign r_1[31] = _352_ | _351_ /*33921*/;
  assign _353_ = ~q[31] /*33920*/;
  assign _354_ = sum_1[32] & q[31] /*33919*/;
  assign _355_ = m_1[32] & _353_ /*33918*/;
  assign r_1[32] = _355_ | _354_ /*33917*/;
  assign _356_ = ~q[31] /*33916*/;
  assign _357_ = sum_1[33] & q[31] /*33915*/;
  assign _358_ = m_1[33] & _356_ /*33914*/;
  assign r_1[33] = _358_ | _357_ /*33913*/;
  assign _359_ = ~q[31] /*33912*/;
  assign _360_ = sum_1[34] & q[31] /*33911*/;
  assign _361_ = m_1[34] & _359_ /*33910*/;
  assign r_1[34] = _361_ | _360_ /*33909*/;
  assign _362_ = ~q[31] /*33908*/;
  assign _363_ = sum_1[35] & q[31] /*33907*/;
  assign _364_ = m_1[35] & _362_ /*33906*/;
  assign r_1[35] = _364_ | _363_ /*33905*/;
  assign _365_ = ~q[31] /*33904*/;
  assign _366_ = sum_1[36] & q[31] /*33903*/;
  assign _367_ = m_1[36] & _365_ /*33902*/;
  assign r_1[36] = _367_ | _366_ /*33901*/;
  assign _368_ = ~q[31] /*33900*/;
  assign _369_ = sum_1[37] & q[31] /*33899*/;
  assign _370_ = m_1[37] & _368_ /*33898*/;
  assign r_1[37] = _370_ | _369_ /*33897*/;
  assign _371_ = ~q[31] /*33896*/;
  assign _372_ = sum_1[38] & q[31] /*33895*/;
  assign _373_ = m_1[38] & _371_ /*33894*/;
  assign r_1[38] = _373_ | _372_ /*33893*/;
  assign _374_ = ~q[31] /*33892*/;
  assign _375_ = sum_1[39] & q[31] /*33891*/;
  assign _376_ = m_1[39] & _374_ /*33890*/;
  assign r_1[39] = _376_ | _375_ /*33889*/;
  assign _377_ = ~q[31] /*33888*/;
  assign _378_ = sum_1[40] & q[31] /*33887*/;
  assign _379_ = m_1[40] & _377_ /*33886*/;
  assign r_1[40] = _379_ | _378_ /*33885*/;
  assign _380_ = ~q[31] /*33884*/;
  assign _381_ = sum_1[41] & q[31] /*33883*/;
  assign _382_ = m_1[41] & _380_ /*33882*/;
  assign r_1[41] = _382_ | _381_ /*33881*/;
  assign _383_ = ~q[31] /*33880*/;
  assign _384_ = sum_1[42] & q[31] /*33879*/;
  assign _385_ = m_1[42] & _383_ /*33878*/;
  assign r_1[42] = _385_ | _384_ /*33877*/;
  assign _386_ = ~q[31] /*33876*/;
  assign _387_ = sum_1[43] & q[31] /*33875*/;
  assign _388_ = m_1[43] & _386_ /*33874*/;
  assign r_1[43] = _388_ | _387_ /*33873*/;
  assign _389_ = ~q[31] /*33872*/;
  assign _390_ = sum_1[44] & q[31] /*33871*/;
  assign _391_ = m_1[44] & _389_ /*33870*/;
  assign r_1[44] = _391_ | _390_ /*33869*/;
  assign _392_ = ~q[31] /*33868*/;
  assign _393_ = sum_1[45] & q[31] /*33867*/;
  assign _394_ = m_1[45] & _392_ /*33866*/;
  assign r_1[45] = _394_ | _393_ /*33865*/;
  assign _395_ = ~q[31] /*33864*/;
  assign _396_ = sum_1[46] & q[31] /*33863*/;
  assign _397_ = m_1[46] & _395_ /*33862*/;
  assign r_1[46] = _397_ | _396_ /*33861*/;
  assign _398_ = ~q[31] /*33860*/;
  assign _399_ = sum_1[47] & q[31] /*33859*/;
  assign _400_ = m_1[47] & _398_ /*33858*/;
  assign r_1[47] = _400_ | _399_ /*33857*/;
  assign _401_ = ~q[31] /*33856*/;
  assign _402_ = sum_1[48] & q[31] /*33855*/;
  assign _403_ = m_1[48] & _401_ /*33854*/;
  assign r_1[48] = _403_ | _402_ /*33853*/;
  assign _404_ = ~q[31] /*33852*/;
  assign _405_ = sum_1[49] & q[31] /*33851*/;
  assign _406_ = m_1[49] & _404_ /*33850*/;
  assign r_1[49] = _406_ | _405_ /*33849*/;
  assign _407_ = ~q[31] /*33848*/;
  assign _408_ = sum_1[50] & q[31] /*33847*/;
  assign _409_ = m_1[50] & _407_ /*33846*/;
  assign r_1[50] = _409_ | _408_ /*33845*/;
  assign _410_ = ~q[31] /*33844*/;
  assign _411_ = sum_1[51] & q[31] /*33843*/;
  assign _412_ = m_1[51] & _410_ /*33842*/;
  assign r_1[51] = _412_ | _411_ /*33841*/;
  assign _413_ = ~q[31] /*33840*/;
  assign _414_ = sum_1[52] & q[31] /*33839*/;
  assign _415_ = m_1[52] & _413_ /*33838*/;
  assign r_1[52] = _415_ | _414_ /*33837*/;
  assign _416_ = ~q[31] /*33836*/;
  assign _417_ = sum_1[53] & q[31] /*33835*/;
  assign _418_ = m_1[53] & _416_ /*33834*/;
  assign r_1[53] = _418_ | _417_ /*33833*/;
  assign _419_ = ~q[31] /*33832*/;
  assign _420_ = sum_1[54] & q[31] /*33831*/;
  assign _421_ = m_1[54] & _419_ /*33830*/;
  assign r_1[54] = _421_ | _420_ /*33829*/;
  assign _422_ = ~q[31] /*33828*/;
  assign _423_ = sum_1[55] & q[31] /*33827*/;
  assign _424_ = m_1[55] & _422_ /*33826*/;
  assign r_1[55] = _424_ | _423_ /*33825*/;
  assign _425_ = ~q[31] /*33824*/;
  assign _426_ = sum_1[56] & q[31] /*33823*/;
  assign _427_ = m_1[56] & _425_ /*33822*/;
  assign r_1[56] = _427_ | _426_ /*33821*/;
  assign _428_ = ~q[31] /*33820*/;
  assign _429_ = sum_1[57] & q[31] /*33819*/;
  assign _430_ = m_1[57] & _428_ /*33818*/;
  assign r_1[57] = _430_ | _429_ /*33817*/;
  assign _431_ = ~q[31] /*33816*/;
  assign _432_ = sum_1[58] & q[31] /*33815*/;
  assign _433_ = m_1[58] & _431_ /*33814*/;
  assign r_1[58] = _433_ | _432_ /*33813*/;
  assign _434_ = ~q[31] /*33812*/;
  assign _435_ = sum_1[59] & q[31] /*33811*/;
  assign _436_ = m_1[59] & _434_ /*33810*/;
  assign r_1[59] = _436_ | _435_ /*33809*/;
  assign _437_ = ~q[31] /*33808*/;
  assign _438_ = sum_1[60] & q[31] /*33807*/;
  assign _439_ = m_1[60] & _437_ /*33806*/;
  assign r_1[60] = _439_ | _438_ /*33805*/;
  assign _440_ = ~q[31] /*33804*/;
  assign _441_ = sum_1[61] & q[31] /*33803*/;
  assign _442_ = m_1[61] & _440_ /*33802*/;
  assign r_1[61] = _442_ | _441_ /*33801*/;
  assign _443_ = ~q[31] /*33800*/;
  assign _444_ = sum_1[62] & q[31] /*33799*/;
  assign _445_ = m_1[62] & _443_ /*33798*/;
  assign r_1[62] = _445_ | _444_ /*33797*/;
  assign _446_ = ~q[31] /*33796*/;
  assign _447_ = sum_1[63] & q[31] /*33795*/;
  assign _448_ = m_1[63] & _446_ /*33794*/;
  assign r_1[63] = _448_ | _447_ /*33793*/;
  assign inv_2[0] = oneWire /*33420*/;
  assign inv_2[1] = oneWire /*33414*/;
  assign inv_2[2] = oneWire /*33408*/;
  assign inv_2[3] = oneWire /*33402*/;
  assign inv_2[4] = oneWire /*33396*/;
  assign inv_2[5] = oneWire /*33390*/;
  assign inv_2[6] = oneWire /*33384*/;
  assign inv_2[7] = oneWire /*33378*/;
  assign inv_2[8] = oneWire /*33372*/;
  assign inv_2[9] = oneWire /*33366*/;
  assign inv_2[10] = oneWire /*33360*/;
  assign inv_2[11] = oneWire /*33354*/;
  assign inv_2[12] = oneWire /*33348*/;
  assign inv_2[13] = oneWire /*33342*/;
  assign inv_2[14] = oneWire /*33336*/;
  assign inv_2[15] = oneWire /*33330*/;
  assign inv_2[16] = oneWire /*33324*/;
  assign inv_2[17] = oneWire /*33318*/;
  assign inv_2[18] = oneWire /*33312*/;
  assign inv_2[19] = oneWire /*33306*/;
  assign inv_2[20] = oneWire /*33300*/;
  assign inv_2[21] = oneWire /*33294*/;
  assign inv_2[22] = oneWire /*33288*/;
  assign inv_2[23] = oneWire /*33282*/;
  assign inv_2[24] = oneWire /*33276*/;
  assign inv_2[25] = oneWire /*33270*/;
  assign inv_2[26] = oneWire /*33264*/;
  assign inv_2[27] = oneWire /*33258*/;
  assign inv_2[28] = oneWire /*33252*/;
  assign inv_2[29] = oneWire /*33246*/;
  assign inv_2[30] = ~div[0] /*33240*/;
  assign inv_2[31] = ~div[1] /*33234*/;
  assign inv_2[32] = ~div[2] /*33228*/;
  assign inv_2[33] = ~div[3] /*33222*/;
  assign inv_2[34] = ~div[4] /*33216*/;
  assign inv_2[35] = ~div[5] /*33210*/;
  assign inv_2[36] = ~div[6] /*33204*/;
  assign inv_2[37] = ~div[7] /*33198*/;
  assign inv_2[38] = ~div[8] /*33192*/;
  assign inv_2[39] = ~div[9] /*33186*/;
  assign inv_2[40] = ~div[10] /*33180*/;
  assign inv_2[41] = ~div[11] /*33174*/;
  assign inv_2[42] = ~div[12] /*33168*/;
  assign inv_2[43] = ~div[13] /*33162*/;
  assign inv_2[44] = ~div[14] /*33156*/;
  assign inv_2[45] = ~div[15] /*33150*/;
  assign inv_2[46] = ~div[16] /*33144*/;
  assign inv_2[47] = ~div[17] /*33138*/;
  assign inv_2[48] = ~div[18] /*33132*/;
  assign inv_2[49] = ~div[19] /*33126*/;
  assign inv_2[50] = ~div[20] /*33120*/;
  assign inv_2[51] = ~div[21] /*33114*/;
  assign inv_2[52] = ~div[22] /*33108*/;
  assign inv_2[53] = ~div[23] /*33102*/;
  assign inv_2[54] = ~div[24] /*33096*/;
  assign inv_2[55] = ~div[25] /*33090*/;
  assign inv_2[56] = ~div[26] /*33084*/;
  assign inv_2[57] = ~div[27] /*33078*/;
  assign inv_2[58] = ~div[28] /*33072*/;
  assign inv_2[59] = ~div[29] /*33066*/;
  assign inv_2[60] = ~div[30] /*33060*/;
  assign inv_2[61] = oneWire /*33054*/;
  assign inv_2[62] = oneWire /*33048*/;
  assign inv_2[63] = oneWire /*33042*/;
  assign _449_ = inv_2[0] ^ r_1[0] /*33419*/;
  assign sum_2[0] = _449_ ^ oneWire /*33418*/;
  assign _450_ = _449_ & oneWire /*33417*/;
  assign _451_ = inv_2[0] & r_1[0] /*33416*/;
  assign _452_ = _450_ | _451_ /*33415*/;
  assign _453_ = inv_2[1] ^ r_1[1] /*33413*/;
  assign sum_2[1] = _453_ ^ _452_ /*33412*/;
  assign _454_ = _453_ & _452_ /*33411*/;
  assign _455_ = inv_2[1] & r_1[1] /*33410*/;
  assign _456_ = _454_ | _455_ /*33409*/;
  assign _457_ = inv_2[2] ^ r_1[2] /*33407*/;
  assign sum_2[2] = _457_ ^ _456_ /*33406*/;
  assign _458_ = _457_ & _456_ /*33405*/;
  assign _459_ = inv_2[2] & r_1[2] /*33404*/;
  assign _460_ = _458_ | _459_ /*33403*/;
  assign _461_ = inv_2[3] ^ r_1[3] /*33401*/;
  assign sum_2[3] = _461_ ^ _460_ /*33400*/;
  assign _462_ = _461_ & _460_ /*33399*/;
  assign _463_ = inv_2[3] & r_1[3] /*33398*/;
  assign _464_ = _462_ | _463_ /*33397*/;
  assign _465_ = inv_2[4] ^ r_1[4] /*33395*/;
  assign sum_2[4] = _465_ ^ _464_ /*33394*/;
  assign _466_ = _465_ & _464_ /*33393*/;
  assign _467_ = inv_2[4] & r_1[4] /*33392*/;
  assign _468_ = _466_ | _467_ /*33391*/;
  assign _469_ = inv_2[5] ^ r_1[5] /*33389*/;
  assign sum_2[5] = _469_ ^ _468_ /*33388*/;
  assign _470_ = _469_ & _468_ /*33387*/;
  assign _471_ = inv_2[5] & r_1[5] /*33386*/;
  assign _472_ = _470_ | _471_ /*33385*/;
  assign _473_ = inv_2[6] ^ r_1[6] /*33383*/;
  assign sum_2[6] = _473_ ^ _472_ /*33382*/;
  assign _474_ = _473_ & _472_ /*33381*/;
  assign _475_ = inv_2[6] & r_1[6] /*33380*/;
  assign _476_ = _474_ | _475_ /*33379*/;
  assign _477_ = inv_2[7] ^ r_1[7] /*33377*/;
  assign sum_2[7] = _477_ ^ _476_ /*33376*/;
  assign _478_ = _477_ & _476_ /*33375*/;
  assign _479_ = inv_2[7] & r_1[7] /*33374*/;
  assign _480_ = _478_ | _479_ /*33373*/;
  assign _481_ = inv_2[8] ^ r_1[8] /*33371*/;
  assign sum_2[8] = _481_ ^ _480_ /*33370*/;
  assign _482_ = _481_ & _480_ /*33369*/;
  assign _483_ = inv_2[8] & r_1[8] /*33368*/;
  assign _484_ = _482_ | _483_ /*33367*/;
  assign _485_ = inv_2[9] ^ r_1[9] /*33365*/;
  assign sum_2[9] = _485_ ^ _484_ /*33364*/;
  assign _486_ = _485_ & _484_ /*33363*/;
  assign _487_ = inv_2[9] & r_1[9] /*33362*/;
  assign _488_ = _486_ | _487_ /*33361*/;
  assign _489_ = inv_2[10] ^ r_1[10] /*33359*/;
  assign sum_2[10] = _489_ ^ _488_ /*33358*/;
  assign _490_ = _489_ & _488_ /*33357*/;
  assign _491_ = inv_2[10] & r_1[10] /*33356*/;
  assign _492_ = _490_ | _491_ /*33355*/;
  assign _493_ = inv_2[11] ^ r_1[11] /*33353*/;
  assign sum_2[11] = _493_ ^ _492_ /*33352*/;
  assign _494_ = _493_ & _492_ /*33351*/;
  assign _495_ = inv_2[11] & r_1[11] /*33350*/;
  assign _496_ = _494_ | _495_ /*33349*/;
  assign _497_ = inv_2[12] ^ r_1[12] /*33347*/;
  assign sum_2[12] = _497_ ^ _496_ /*33346*/;
  assign _498_ = _497_ & _496_ /*33345*/;
  assign _499_ = inv_2[12] & r_1[12] /*33344*/;
  assign _500_ = _498_ | _499_ /*33343*/;
  assign _501_ = inv_2[13] ^ r_1[13] /*33341*/;
  assign sum_2[13] = _501_ ^ _500_ /*33340*/;
  assign _502_ = _501_ & _500_ /*33339*/;
  assign _503_ = inv_2[13] & r_1[13] /*33338*/;
  assign _504_ = _502_ | _503_ /*33337*/;
  assign _505_ = inv_2[14] ^ r_1[14] /*33335*/;
  assign sum_2[14] = _505_ ^ _504_ /*33334*/;
  assign _506_ = _505_ & _504_ /*33333*/;
  assign _507_ = inv_2[14] & r_1[14] /*33332*/;
  assign _508_ = _506_ | _507_ /*33331*/;
  assign _509_ = inv_2[15] ^ r_1[15] /*33329*/;
  assign sum_2[15] = _509_ ^ _508_ /*33328*/;
  assign _510_ = _509_ & _508_ /*33327*/;
  assign _511_ = inv_2[15] & r_1[15] /*33326*/;
  assign _512_ = _510_ | _511_ /*33325*/;
  assign _513_ = inv_2[16] ^ r_1[16] /*33323*/;
  assign sum_2[16] = _513_ ^ _512_ /*33322*/;
  assign _514_ = _513_ & _512_ /*33321*/;
  assign _515_ = inv_2[16] & r_1[16] /*33320*/;
  assign _516_ = _514_ | _515_ /*33319*/;
  assign _517_ = inv_2[17] ^ r_1[17] /*33317*/;
  assign sum_2[17] = _517_ ^ _516_ /*33316*/;
  assign _518_ = _517_ & _516_ /*33315*/;
  assign _519_ = inv_2[17] & r_1[17] /*33314*/;
  assign _520_ = _518_ | _519_ /*33313*/;
  assign _521_ = inv_2[18] ^ r_1[18] /*33311*/;
  assign sum_2[18] = _521_ ^ _520_ /*33310*/;
  assign _522_ = _521_ & _520_ /*33309*/;
  assign _523_ = inv_2[18] & r_1[18] /*33308*/;
  assign _524_ = _522_ | _523_ /*33307*/;
  assign _525_ = inv_2[19] ^ r_1[19] /*33305*/;
  assign sum_2[19] = _525_ ^ _524_ /*33304*/;
  assign _526_ = _525_ & _524_ /*33303*/;
  assign _527_ = inv_2[19] & r_1[19] /*33302*/;
  assign _528_ = _526_ | _527_ /*33301*/;
  assign _529_ = inv_2[20] ^ r_1[20] /*33299*/;
  assign sum_2[20] = _529_ ^ _528_ /*33298*/;
  assign _530_ = _529_ & _528_ /*33297*/;
  assign _531_ = inv_2[20] & r_1[20] /*33296*/;
  assign _532_ = _530_ | _531_ /*33295*/;
  assign _533_ = inv_2[21] ^ r_1[21] /*33293*/;
  assign sum_2[21] = _533_ ^ _532_ /*33292*/;
  assign _534_ = _533_ & _532_ /*33291*/;
  assign _535_ = inv_2[21] & r_1[21] /*33290*/;
  assign _536_ = _534_ | _535_ /*33289*/;
  assign _537_ = inv_2[22] ^ r_1[22] /*33287*/;
  assign sum_2[22] = _537_ ^ _536_ /*33286*/;
  assign _538_ = _537_ & _536_ /*33285*/;
  assign _539_ = inv_2[22] & r_1[22] /*33284*/;
  assign _540_ = _538_ | _539_ /*33283*/;
  assign _541_ = inv_2[23] ^ r_1[23] /*33281*/;
  assign sum_2[23] = _541_ ^ _540_ /*33280*/;
  assign _542_ = _541_ & _540_ /*33279*/;
  assign _543_ = inv_2[23] & r_1[23] /*33278*/;
  assign _544_ = _542_ | _543_ /*33277*/;
  assign _545_ = inv_2[24] ^ r_1[24] /*33275*/;
  assign sum_2[24] = _545_ ^ _544_ /*33274*/;
  assign _546_ = _545_ & _544_ /*33273*/;
  assign _547_ = inv_2[24] & r_1[24] /*33272*/;
  assign _548_ = _546_ | _547_ /*33271*/;
  assign _549_ = inv_2[25] ^ r_1[25] /*33269*/;
  assign sum_2[25] = _549_ ^ _548_ /*33268*/;
  assign _550_ = _549_ & _548_ /*33267*/;
  assign _551_ = inv_2[25] & r_1[25] /*33266*/;
  assign _552_ = _550_ | _551_ /*33265*/;
  assign _553_ = inv_2[26] ^ r_1[26] /*33263*/;
  assign sum_2[26] = _553_ ^ _552_ /*33262*/;
  assign _554_ = _553_ & _552_ /*33261*/;
  assign _555_ = inv_2[26] & r_1[26] /*33260*/;
  assign _556_ = _554_ | _555_ /*33259*/;
  assign _557_ = inv_2[27] ^ r_1[27] /*33257*/;
  assign sum_2[27] = _557_ ^ _556_ /*33256*/;
  assign _558_ = _557_ & _556_ /*33255*/;
  assign _559_ = inv_2[27] & r_1[27] /*33254*/;
  assign _560_ = _558_ | _559_ /*33253*/;
  assign _561_ = inv_2[28] ^ r_1[28] /*33251*/;
  assign sum_2[28] = _561_ ^ _560_ /*33250*/;
  assign _562_ = _561_ & _560_ /*33249*/;
  assign _563_ = inv_2[28] & r_1[28] /*33248*/;
  assign _564_ = _562_ | _563_ /*33247*/;
  assign _565_ = inv_2[29] ^ r_1[29] /*33245*/;
  assign sum_2[29] = _565_ ^ _564_ /*33244*/;
  assign _566_ = _565_ & _564_ /*33243*/;
  assign _567_ = inv_2[29] & r_1[29] /*33242*/;
  assign _568_ = _566_ | _567_ /*33241*/;
  assign _569_ = inv_2[30] ^ r_1[30] /*33239*/;
  assign sum_2[30] = _569_ ^ _568_ /*33238*/;
  assign _570_ = _569_ & _568_ /*33237*/;
  assign _571_ = inv_2[30] & r_1[30] /*33236*/;
  assign _572_ = _570_ | _571_ /*33235*/;
  assign _573_ = inv_2[31] ^ r_1[31] /*33233*/;
  assign sum_2[31] = _573_ ^ _572_ /*33232*/;
  assign _574_ = _573_ & _572_ /*33231*/;
  assign _575_ = inv_2[31] & r_1[31] /*33230*/;
  assign _576_ = _574_ | _575_ /*33229*/;
  assign _577_ = inv_2[32] ^ r_1[32] /*33227*/;
  assign sum_2[32] = _577_ ^ _576_ /*33226*/;
  assign _578_ = _577_ & _576_ /*33225*/;
  assign _579_ = inv_2[32] & r_1[32] /*33224*/;
  assign _580_ = _578_ | _579_ /*33223*/;
  assign _581_ = inv_2[33] ^ r_1[33] /*33221*/;
  assign sum_2[33] = _581_ ^ _580_ /*33220*/;
  assign _582_ = _581_ & _580_ /*33219*/;
  assign _583_ = inv_2[33] & r_1[33] /*33218*/;
  assign _584_ = _582_ | _583_ /*33217*/;
  assign _585_ = inv_2[34] ^ r_1[34] /*33215*/;
  assign sum_2[34] = _585_ ^ _584_ /*33214*/;
  assign _586_ = _585_ & _584_ /*33213*/;
  assign _587_ = inv_2[34] & r_1[34] /*33212*/;
  assign _588_ = _586_ | _587_ /*33211*/;
  assign _589_ = inv_2[35] ^ r_1[35] /*33209*/;
  assign sum_2[35] = _589_ ^ _588_ /*33208*/;
  assign _590_ = _589_ & _588_ /*33207*/;
  assign _591_ = inv_2[35] & r_1[35] /*33206*/;
  assign _592_ = _590_ | _591_ /*33205*/;
  assign _593_ = inv_2[36] ^ r_1[36] /*33203*/;
  assign sum_2[36] = _593_ ^ _592_ /*33202*/;
  assign _594_ = _593_ & _592_ /*33201*/;
  assign _595_ = inv_2[36] & r_1[36] /*33200*/;
  assign _596_ = _594_ | _595_ /*33199*/;
  assign _597_ = inv_2[37] ^ r_1[37] /*33197*/;
  assign sum_2[37] = _597_ ^ _596_ /*33196*/;
  assign _598_ = _597_ & _596_ /*33195*/;
  assign _599_ = inv_2[37] & r_1[37] /*33194*/;
  assign _600_ = _598_ | _599_ /*33193*/;
  assign _601_ = inv_2[38] ^ r_1[38] /*33191*/;
  assign sum_2[38] = _601_ ^ _600_ /*33190*/;
  assign _602_ = _601_ & _600_ /*33189*/;
  assign _603_ = inv_2[38] & r_1[38] /*33188*/;
  assign _604_ = _602_ | _603_ /*33187*/;
  assign _605_ = inv_2[39] ^ r_1[39] /*33185*/;
  assign sum_2[39] = _605_ ^ _604_ /*33184*/;
  assign _606_ = _605_ & _604_ /*33183*/;
  assign _607_ = inv_2[39] & r_1[39] /*33182*/;
  assign _608_ = _606_ | _607_ /*33181*/;
  assign _609_ = inv_2[40] ^ r_1[40] /*33179*/;
  assign sum_2[40] = _609_ ^ _608_ /*33178*/;
  assign _610_ = _609_ & _608_ /*33177*/;
  assign _611_ = inv_2[40] & r_1[40] /*33176*/;
  assign _612_ = _610_ | _611_ /*33175*/;
  assign _613_ = inv_2[41] ^ r_1[41] /*33173*/;
  assign sum_2[41] = _613_ ^ _612_ /*33172*/;
  assign _614_ = _613_ & _612_ /*33171*/;
  assign _615_ = inv_2[41] & r_1[41] /*33170*/;
  assign _616_ = _614_ | _615_ /*33169*/;
  assign _617_ = inv_2[42] ^ r_1[42] /*33167*/;
  assign sum_2[42] = _617_ ^ _616_ /*33166*/;
  assign _618_ = _617_ & _616_ /*33165*/;
  assign _619_ = inv_2[42] & r_1[42] /*33164*/;
  assign _620_ = _618_ | _619_ /*33163*/;
  assign _621_ = inv_2[43] ^ r_1[43] /*33161*/;
  assign sum_2[43] = _621_ ^ _620_ /*33160*/;
  assign _622_ = _621_ & _620_ /*33159*/;
  assign _623_ = inv_2[43] & r_1[43] /*33158*/;
  assign _624_ = _622_ | _623_ /*33157*/;
  assign _625_ = inv_2[44] ^ r_1[44] /*33155*/;
  assign sum_2[44] = _625_ ^ _624_ /*33154*/;
  assign _626_ = _625_ & _624_ /*33153*/;
  assign _627_ = inv_2[44] & r_1[44] /*33152*/;
  assign _628_ = _626_ | _627_ /*33151*/;
  assign _629_ = inv_2[45] ^ r_1[45] /*33149*/;
  assign sum_2[45] = _629_ ^ _628_ /*33148*/;
  assign _630_ = _629_ & _628_ /*33147*/;
  assign _631_ = inv_2[45] & r_1[45] /*33146*/;
  assign _632_ = _630_ | _631_ /*33145*/;
  assign _633_ = inv_2[46] ^ r_1[46] /*33143*/;
  assign sum_2[46] = _633_ ^ _632_ /*33142*/;
  assign _634_ = _633_ & _632_ /*33141*/;
  assign _635_ = inv_2[46] & r_1[46] /*33140*/;
  assign _636_ = _634_ | _635_ /*33139*/;
  assign _637_ = inv_2[47] ^ r_1[47] /*33137*/;
  assign sum_2[47] = _637_ ^ _636_ /*33136*/;
  assign _638_ = _637_ & _636_ /*33135*/;
  assign _639_ = inv_2[47] & r_1[47] /*33134*/;
  assign _640_ = _638_ | _639_ /*33133*/;
  assign _641_ = inv_2[48] ^ r_1[48] /*33131*/;
  assign sum_2[48] = _641_ ^ _640_ /*33130*/;
  assign _642_ = _641_ & _640_ /*33129*/;
  assign _643_ = inv_2[48] & r_1[48] /*33128*/;
  assign _644_ = _642_ | _643_ /*33127*/;
  assign _645_ = inv_2[49] ^ r_1[49] /*33125*/;
  assign sum_2[49] = _645_ ^ _644_ /*33124*/;
  assign _646_ = _645_ & _644_ /*33123*/;
  assign _647_ = inv_2[49] & r_1[49] /*33122*/;
  assign _648_ = _646_ | _647_ /*33121*/;
  assign _649_ = inv_2[50] ^ r_1[50] /*33119*/;
  assign sum_2[50] = _649_ ^ _648_ /*33118*/;
  assign _650_ = _649_ & _648_ /*33117*/;
  assign _651_ = inv_2[50] & r_1[50] /*33116*/;
  assign _652_ = _650_ | _651_ /*33115*/;
  assign _653_ = inv_2[51] ^ r_1[51] /*33113*/;
  assign sum_2[51] = _653_ ^ _652_ /*33112*/;
  assign _654_ = _653_ & _652_ /*33111*/;
  assign _655_ = inv_2[51] & r_1[51] /*33110*/;
  assign _656_ = _654_ | _655_ /*33109*/;
  assign _657_ = inv_2[52] ^ r_1[52] /*33107*/;
  assign sum_2[52] = _657_ ^ _656_ /*33106*/;
  assign _658_ = _657_ & _656_ /*33105*/;
  assign _659_ = inv_2[52] & r_1[52] /*33104*/;
  assign _660_ = _658_ | _659_ /*33103*/;
  assign _661_ = inv_2[53] ^ r_1[53] /*33101*/;
  assign sum_2[53] = _661_ ^ _660_ /*33100*/;
  assign _662_ = _661_ & _660_ /*33099*/;
  assign _663_ = inv_2[53] & r_1[53] /*33098*/;
  assign _664_ = _662_ | _663_ /*33097*/;
  assign _665_ = inv_2[54] ^ r_1[54] /*33095*/;
  assign sum_2[54] = _665_ ^ _664_ /*33094*/;
  assign _666_ = _665_ & _664_ /*33093*/;
  assign _667_ = inv_2[54] & r_1[54] /*33092*/;
  assign _668_ = _666_ | _667_ /*33091*/;
  assign _669_ = inv_2[55] ^ r_1[55] /*33089*/;
  assign sum_2[55] = _669_ ^ _668_ /*33088*/;
  assign _670_ = _669_ & _668_ /*33087*/;
  assign _671_ = inv_2[55] & r_1[55] /*33086*/;
  assign _672_ = _670_ | _671_ /*33085*/;
  assign _673_ = inv_2[56] ^ r_1[56] /*33083*/;
  assign sum_2[56] = _673_ ^ _672_ /*33082*/;
  assign _674_ = _673_ & _672_ /*33081*/;
  assign _675_ = inv_2[56] & r_1[56] /*33080*/;
  assign _676_ = _674_ | _675_ /*33079*/;
  assign _677_ = inv_2[57] ^ r_1[57] /*33077*/;
  assign sum_2[57] = _677_ ^ _676_ /*33076*/;
  assign _678_ = _677_ & _676_ /*33075*/;
  assign _679_ = inv_2[57] & r_1[57] /*33074*/;
  assign _680_ = _678_ | _679_ /*33073*/;
  assign _681_ = inv_2[58] ^ r_1[58] /*33071*/;
  assign sum_2[58] = _681_ ^ _680_ /*33070*/;
  assign _682_ = _681_ & _680_ /*33069*/;
  assign _683_ = inv_2[58] & r_1[58] /*33068*/;
  assign _684_ = _682_ | _683_ /*33067*/;
  assign _685_ = inv_2[59] ^ r_1[59] /*33065*/;
  assign sum_2[59] = _685_ ^ _684_ /*33064*/;
  assign _686_ = _685_ & _684_ /*33063*/;
  assign _687_ = inv_2[59] & r_1[59] /*33062*/;
  assign _688_ = _686_ | _687_ /*33061*/;
  assign _689_ = inv_2[60] ^ r_1[60] /*33059*/;
  assign sum_2[60] = _689_ ^ _688_ /*33058*/;
  assign _690_ = _689_ & _688_ /*33057*/;
  assign _691_ = inv_2[60] & r_1[60] /*33056*/;
  assign _692_ = _690_ | _691_ /*33055*/;
  assign _693_ = inv_2[61] ^ r_1[61] /*33053*/;
  assign sum_2[61] = _693_ ^ _692_ /*33052*/;
  assign _694_ = _693_ & _692_ /*33051*/;
  assign _695_ = inv_2[61] & r_1[61] /*33050*/;
  assign _696_ = _694_ | _695_ /*33049*/;
  assign _697_ = inv_2[62] ^ r_1[62] /*33047*/;
  assign sum_2[62] = _697_ ^ _696_ /*33046*/;
  assign _698_ = _697_ & _696_ /*33045*/;
  assign _699_ = inv_2[62] & r_1[62] /*33044*/;
  assign _700_ = _698_ | _699_ /*33043*/;
  assign _701_ = inv_2[63] ^ r_1[63] /*33041*/;
  assign sum_2[63] = _701_ ^ _700_ /*33040*/;
  assign _702_ = _701_ & _700_ /*33039*/;
  assign _703_ = inv_2[63] & r_1[63] /*33038*/;
  assign _704_ = _702_ | _703_ /*33037*/;
  assign _705_ = _704_ ^ _700_ /*33036*/;
  assign _706_ = ~_705_ /*33035*/;
  assign _707_ = sum_2[63] & _706_ /*33034*/;
  assign _708_ = _705_ & _704_ /*33033*/;
  assign sum_2[64] = _708_ | _707_ /*33032*/;
  assign q[30] = ~sum_2[64] /*33031*/;
  assign m_2[0] = r_1[0] /*33030*/;
  assign m_2[1] = r_1[1] /*33029*/;
  assign m_2[2] = r_1[2] /*33028*/;
  assign m_2[3] = r_1[3] /*33027*/;
  assign m_2[4] = r_1[4] /*33026*/;
  assign m_2[5] = r_1[5] /*33025*/;
  assign m_2[6] = r_1[6] /*33024*/;
  assign m_2[7] = r_1[7] /*33023*/;
  assign m_2[8] = r_1[8] /*33022*/;
  assign m_2[9] = r_1[9] /*33021*/;
  assign m_2[10] = r_1[10] /*33020*/;
  assign m_2[11] = r_1[11] /*33019*/;
  assign m_2[12] = r_1[12] /*33018*/;
  assign m_2[13] = r_1[13] /*33017*/;
  assign m_2[14] = r_1[14] /*33016*/;
  assign m_2[15] = r_1[15] /*33015*/;
  assign m_2[16] = r_1[16] /*33014*/;
  assign m_2[17] = r_1[17] /*33013*/;
  assign m_2[18] = r_1[18] /*33012*/;
  assign m_2[19] = r_1[19] /*33011*/;
  assign m_2[20] = r_1[20] /*33010*/;
  assign m_2[21] = r_1[21] /*33009*/;
  assign m_2[22] = r_1[22] /*33008*/;
  assign m_2[23] = r_1[23] /*33007*/;
  assign m_2[24] = r_1[24] /*33006*/;
  assign m_2[25] = r_1[25] /*33005*/;
  assign m_2[26] = r_1[26] /*33004*/;
  assign m_2[27] = r_1[27] /*33003*/;
  assign m_2[28] = r_1[28] /*33002*/;
  assign m_2[29] = r_1[29] /*33001*/;
  assign m_2[30] = r_1[30] /*33000*/;
  assign m_2[31] = r_1[31] /*32999*/;
  assign m_2[32] = r_1[32] /*32998*/;
  assign m_2[33] = r_1[33] /*32997*/;
  assign m_2[34] = r_1[34] /*32996*/;
  assign m_2[35] = r_1[35] /*32995*/;
  assign m_2[36] = r_1[36] /*32994*/;
  assign m_2[37] = r_1[37] /*32993*/;
  assign m_2[38] = r_1[38] /*32992*/;
  assign m_2[39] = r_1[39] /*32991*/;
  assign m_2[40] = r_1[40] /*32990*/;
  assign m_2[41] = r_1[41] /*32989*/;
  assign m_2[42] = r_1[42] /*32988*/;
  assign m_2[43] = r_1[43] /*32987*/;
  assign m_2[44] = r_1[44] /*32986*/;
  assign m_2[45] = r_1[45] /*32985*/;
  assign m_2[46] = r_1[46] /*32984*/;
  assign m_2[47] = r_1[47] /*32983*/;
  assign m_2[48] = r_1[48] /*32982*/;
  assign m_2[49] = r_1[49] /*32981*/;
  assign m_2[50] = r_1[50] /*32980*/;
  assign m_2[51] = r_1[51] /*32979*/;
  assign m_2[52] = r_1[52] /*32978*/;
  assign m_2[53] = r_1[53] /*32977*/;
  assign m_2[54] = r_1[54] /*32976*/;
  assign m_2[55] = r_1[55] /*32975*/;
  assign m_2[56] = r_1[56] /*32974*/;
  assign m_2[57] = r_1[57] /*32973*/;
  assign m_2[58] = r_1[58] /*32972*/;
  assign m_2[59] = r_1[59] /*32971*/;
  assign m_2[60] = r_1[60] /*32970*/;
  assign m_2[61] = r_1[61] /*32969*/;
  assign m_2[62] = r_1[62] /*32968*/;
  assign m_2[63] = r_1[63] /*32967*/;
  assign m_2[64] = r_1[63] /*32966*/;
  assign _710_ = ~q[30] /*32965*/;
  assign _711_ = sum_2[0] & q[30] /*32964*/;
  assign _712_ = m_2[0] & _710_ /*32963*/;
  assign r_2[0] = _712_ | _711_ /*32962*/;
  assign _713_ = ~q[30] /*32961*/;
  assign _714_ = sum_2[1] & q[30] /*32960*/;
  assign _715_ = m_2[1] & _713_ /*32959*/;
  assign r_2[1] = _715_ | _714_ /*32958*/;
  assign _716_ = ~q[30] /*32957*/;
  assign _717_ = sum_2[2] & q[30] /*32956*/;
  assign _718_ = m_2[2] & _716_ /*32955*/;
  assign r_2[2] = _718_ | _717_ /*32954*/;
  assign _719_ = ~q[30] /*32953*/;
  assign _720_ = sum_2[3] & q[30] /*32952*/;
  assign _721_ = m_2[3] & _719_ /*32951*/;
  assign r_2[3] = _721_ | _720_ /*32950*/;
  assign _722_ = ~q[30] /*32949*/;
  assign _723_ = sum_2[4] & q[30] /*32948*/;
  assign _724_ = m_2[4] & _722_ /*32947*/;
  assign r_2[4] = _724_ | _723_ /*32946*/;
  assign _725_ = ~q[30] /*32945*/;
  assign _726_ = sum_2[5] & q[30] /*32944*/;
  assign _727_ = m_2[5] & _725_ /*32943*/;
  assign r_2[5] = _727_ | _726_ /*32942*/;
  assign _728_ = ~q[30] /*32941*/;
  assign _729_ = sum_2[6] & q[30] /*32940*/;
  assign _730_ = m_2[6] & _728_ /*32939*/;
  assign r_2[6] = _730_ | _729_ /*32938*/;
  assign _731_ = ~q[30] /*32937*/;
  assign _732_ = sum_2[7] & q[30] /*32936*/;
  assign _733_ = m_2[7] & _731_ /*32935*/;
  assign r_2[7] = _733_ | _732_ /*32934*/;
  assign _734_ = ~q[30] /*32933*/;
  assign _735_ = sum_2[8] & q[30] /*32932*/;
  assign _736_ = m_2[8] & _734_ /*32931*/;
  assign r_2[8] = _736_ | _735_ /*32930*/;
  assign _737_ = ~q[30] /*32929*/;
  assign _738_ = sum_2[9] & q[30] /*32928*/;
  assign _739_ = m_2[9] & _737_ /*32927*/;
  assign r_2[9] = _739_ | _738_ /*32926*/;
  assign _740_ = ~q[30] /*32925*/;
  assign _741_ = sum_2[10] & q[30] /*32924*/;
  assign _742_ = m_2[10] & _740_ /*32923*/;
  assign r_2[10] = _742_ | _741_ /*32922*/;
  assign _743_ = ~q[30] /*32921*/;
  assign _744_ = sum_2[11] & q[30] /*32920*/;
  assign _745_ = m_2[11] & _743_ /*32919*/;
  assign r_2[11] = _745_ | _744_ /*32918*/;
  assign _746_ = ~q[30] /*32917*/;
  assign _747_ = sum_2[12] & q[30] /*32916*/;
  assign _748_ = m_2[12] & _746_ /*32915*/;
  assign r_2[12] = _748_ | _747_ /*32914*/;
  assign _749_ = ~q[30] /*32913*/;
  assign _750_ = sum_2[13] & q[30] /*32912*/;
  assign _751_ = m_2[13] & _749_ /*32911*/;
  assign r_2[13] = _751_ | _750_ /*32910*/;
  assign _752_ = ~q[30] /*32909*/;
  assign _753_ = sum_2[14] & q[30] /*32908*/;
  assign _754_ = m_2[14] & _752_ /*32907*/;
  assign r_2[14] = _754_ | _753_ /*32906*/;
  assign _755_ = ~q[30] /*32905*/;
  assign _756_ = sum_2[15] & q[30] /*32904*/;
  assign _757_ = m_2[15] & _755_ /*32903*/;
  assign r_2[15] = _757_ | _756_ /*32902*/;
  assign _758_ = ~q[30] /*32901*/;
  assign _759_ = sum_2[16] & q[30] /*32900*/;
  assign _760_ = m_2[16] & _758_ /*32899*/;
  assign r_2[16] = _760_ | _759_ /*32898*/;
  assign _761_ = ~q[30] /*32897*/;
  assign _762_ = sum_2[17] & q[30] /*32896*/;
  assign _763_ = m_2[17] & _761_ /*32895*/;
  assign r_2[17] = _763_ | _762_ /*32894*/;
  assign _764_ = ~q[30] /*32893*/;
  assign _765_ = sum_2[18] & q[30] /*32892*/;
  assign _766_ = m_2[18] & _764_ /*32891*/;
  assign r_2[18] = _766_ | _765_ /*32890*/;
  assign _767_ = ~q[30] /*32889*/;
  assign _768_ = sum_2[19] & q[30] /*32888*/;
  assign _769_ = m_2[19] & _767_ /*32887*/;
  assign r_2[19] = _769_ | _768_ /*32886*/;
  assign _770_ = ~q[30] /*32885*/;
  assign _771_ = sum_2[20] & q[30] /*32884*/;
  assign _772_ = m_2[20] & _770_ /*32883*/;
  assign r_2[20] = _772_ | _771_ /*32882*/;
  assign _773_ = ~q[30] /*32881*/;
  assign _774_ = sum_2[21] & q[30] /*32880*/;
  assign _775_ = m_2[21] & _773_ /*32879*/;
  assign r_2[21] = _775_ | _774_ /*32878*/;
  assign _776_ = ~q[30] /*32877*/;
  assign _777_ = sum_2[22] & q[30] /*32876*/;
  assign _778_ = m_2[22] & _776_ /*32875*/;
  assign r_2[22] = _778_ | _777_ /*32874*/;
  assign _779_ = ~q[30] /*32873*/;
  assign _780_ = sum_2[23] & q[30] /*32872*/;
  assign _781_ = m_2[23] & _779_ /*32871*/;
  assign r_2[23] = _781_ | _780_ /*32870*/;
  assign _782_ = ~q[30] /*32869*/;
  assign _783_ = sum_2[24] & q[30] /*32868*/;
  assign _784_ = m_2[24] & _782_ /*32867*/;
  assign r_2[24] = _784_ | _783_ /*32866*/;
  assign _785_ = ~q[30] /*32865*/;
  assign _786_ = sum_2[25] & q[30] /*32864*/;
  assign _787_ = m_2[25] & _785_ /*32863*/;
  assign r_2[25] = _787_ | _786_ /*32862*/;
  assign _788_ = ~q[30] /*32861*/;
  assign _789_ = sum_2[26] & q[30] /*32860*/;
  assign _790_ = m_2[26] & _788_ /*32859*/;
  assign r_2[26] = _790_ | _789_ /*32858*/;
  assign _791_ = ~q[30] /*32857*/;
  assign _792_ = sum_2[27] & q[30] /*32856*/;
  assign _793_ = m_2[27] & _791_ /*32855*/;
  assign r_2[27] = _793_ | _792_ /*32854*/;
  assign _794_ = ~q[30] /*32853*/;
  assign _795_ = sum_2[28] & q[30] /*32852*/;
  assign _796_ = m_2[28] & _794_ /*32851*/;
  assign r_2[28] = _796_ | _795_ /*32850*/;
  assign _797_ = ~q[30] /*32849*/;
  assign _798_ = sum_2[29] & q[30] /*32848*/;
  assign _799_ = m_2[29] & _797_ /*32847*/;
  assign r_2[29] = _799_ | _798_ /*32846*/;
  assign _800_ = ~q[30] /*32845*/;
  assign _801_ = sum_2[30] & q[30] /*32844*/;
  assign _802_ = m_2[30] & _800_ /*32843*/;
  assign r_2[30] = _802_ | _801_ /*32842*/;
  assign _803_ = ~q[30] /*32841*/;
  assign _804_ = sum_2[31] & q[30] /*32840*/;
  assign _805_ = m_2[31] & _803_ /*32839*/;
  assign r_2[31] = _805_ | _804_ /*32838*/;
  assign _806_ = ~q[30] /*32837*/;
  assign _807_ = sum_2[32] & q[30] /*32836*/;
  assign _808_ = m_2[32] & _806_ /*32835*/;
  assign r_2[32] = _808_ | _807_ /*32834*/;
  assign _809_ = ~q[30] /*32833*/;
  assign _810_ = sum_2[33] & q[30] /*32832*/;
  assign _811_ = m_2[33] & _809_ /*32831*/;
  assign r_2[33] = _811_ | _810_ /*32830*/;
  assign _812_ = ~q[30] /*32829*/;
  assign _813_ = sum_2[34] & q[30] /*32828*/;
  assign _814_ = m_2[34] & _812_ /*32827*/;
  assign r_2[34] = _814_ | _813_ /*32826*/;
  assign _815_ = ~q[30] /*32825*/;
  assign _816_ = sum_2[35] & q[30] /*32824*/;
  assign _817_ = m_2[35] & _815_ /*32823*/;
  assign r_2[35] = _817_ | _816_ /*32822*/;
  assign _818_ = ~q[30] /*32821*/;
  assign _819_ = sum_2[36] & q[30] /*32820*/;
  assign _820_ = m_2[36] & _818_ /*32819*/;
  assign r_2[36] = _820_ | _819_ /*32818*/;
  assign _821_ = ~q[30] /*32817*/;
  assign _822_ = sum_2[37] & q[30] /*32816*/;
  assign _823_ = m_2[37] & _821_ /*32815*/;
  assign r_2[37] = _823_ | _822_ /*32814*/;
  assign _824_ = ~q[30] /*32813*/;
  assign _825_ = sum_2[38] & q[30] /*32812*/;
  assign _826_ = m_2[38] & _824_ /*32811*/;
  assign r_2[38] = _826_ | _825_ /*32810*/;
  assign _827_ = ~q[30] /*32809*/;
  assign _828_ = sum_2[39] & q[30] /*32808*/;
  assign _829_ = m_2[39] & _827_ /*32807*/;
  assign r_2[39] = _829_ | _828_ /*32806*/;
  assign _830_ = ~q[30] /*32805*/;
  assign _831_ = sum_2[40] & q[30] /*32804*/;
  assign _832_ = m_2[40] & _830_ /*32803*/;
  assign r_2[40] = _832_ | _831_ /*32802*/;
  assign _833_ = ~q[30] /*32801*/;
  assign _834_ = sum_2[41] & q[30] /*32800*/;
  assign _835_ = m_2[41] & _833_ /*32799*/;
  assign r_2[41] = _835_ | _834_ /*32798*/;
  assign _836_ = ~q[30] /*32797*/;
  assign _837_ = sum_2[42] & q[30] /*32796*/;
  assign _838_ = m_2[42] & _836_ /*32795*/;
  assign r_2[42] = _838_ | _837_ /*32794*/;
  assign _839_ = ~q[30] /*32793*/;
  assign _840_ = sum_2[43] & q[30] /*32792*/;
  assign _841_ = m_2[43] & _839_ /*32791*/;
  assign r_2[43] = _841_ | _840_ /*32790*/;
  assign _842_ = ~q[30] /*32789*/;
  assign _843_ = sum_2[44] & q[30] /*32788*/;
  assign _844_ = m_2[44] & _842_ /*32787*/;
  assign r_2[44] = _844_ | _843_ /*32786*/;
  assign _845_ = ~q[30] /*32785*/;
  assign _846_ = sum_2[45] & q[30] /*32784*/;
  assign _847_ = m_2[45] & _845_ /*32783*/;
  assign r_2[45] = _847_ | _846_ /*32782*/;
  assign _848_ = ~q[30] /*32781*/;
  assign _849_ = sum_2[46] & q[30] /*32780*/;
  assign _850_ = m_2[46] & _848_ /*32779*/;
  assign r_2[46] = _850_ | _849_ /*32778*/;
  assign _851_ = ~q[30] /*32777*/;
  assign _852_ = sum_2[47] & q[30] /*32776*/;
  assign _853_ = m_2[47] & _851_ /*32775*/;
  assign r_2[47] = _853_ | _852_ /*32774*/;
  assign _854_ = ~q[30] /*32773*/;
  assign _855_ = sum_2[48] & q[30] /*32772*/;
  assign _856_ = m_2[48] & _854_ /*32771*/;
  assign r_2[48] = _856_ | _855_ /*32770*/;
  assign _857_ = ~q[30] /*32769*/;
  assign _858_ = sum_2[49] & q[30] /*32768*/;
  assign _859_ = m_2[49] & _857_ /*32767*/;
  assign r_2[49] = _859_ | _858_ /*32766*/;
  assign _860_ = ~q[30] /*32765*/;
  assign _861_ = sum_2[50] & q[30] /*32764*/;
  assign _862_ = m_2[50] & _860_ /*32763*/;
  assign r_2[50] = _862_ | _861_ /*32762*/;
  assign _863_ = ~q[30] /*32761*/;
  assign _864_ = sum_2[51] & q[30] /*32760*/;
  assign _865_ = m_2[51] & _863_ /*32759*/;
  assign r_2[51] = _865_ | _864_ /*32758*/;
  assign _866_ = ~q[30] /*32757*/;
  assign _867_ = sum_2[52] & q[30] /*32756*/;
  assign _868_ = m_2[52] & _866_ /*32755*/;
  assign r_2[52] = _868_ | _867_ /*32754*/;
  assign _869_ = ~q[30] /*32753*/;
  assign _870_ = sum_2[53] & q[30] /*32752*/;
  assign _871_ = m_2[53] & _869_ /*32751*/;
  assign r_2[53] = _871_ | _870_ /*32750*/;
  assign _872_ = ~q[30] /*32749*/;
  assign _873_ = sum_2[54] & q[30] /*32748*/;
  assign _874_ = m_2[54] & _872_ /*32747*/;
  assign r_2[54] = _874_ | _873_ /*32746*/;
  assign _875_ = ~q[30] /*32745*/;
  assign _876_ = sum_2[55] & q[30] /*32744*/;
  assign _877_ = m_2[55] & _875_ /*32743*/;
  assign r_2[55] = _877_ | _876_ /*32742*/;
  assign _878_ = ~q[30] /*32741*/;
  assign _879_ = sum_2[56] & q[30] /*32740*/;
  assign _880_ = m_2[56] & _878_ /*32739*/;
  assign r_2[56] = _880_ | _879_ /*32738*/;
  assign _881_ = ~q[30] /*32737*/;
  assign _882_ = sum_2[57] & q[30] /*32736*/;
  assign _883_ = m_2[57] & _881_ /*32735*/;
  assign r_2[57] = _883_ | _882_ /*32734*/;
  assign _884_ = ~q[30] /*32733*/;
  assign _885_ = sum_2[58] & q[30] /*32732*/;
  assign _886_ = m_2[58] & _884_ /*32731*/;
  assign r_2[58] = _886_ | _885_ /*32730*/;
  assign _887_ = ~q[30] /*32729*/;
  assign _888_ = sum_2[59] & q[30] /*32728*/;
  assign _889_ = m_2[59] & _887_ /*32727*/;
  assign r_2[59] = _889_ | _888_ /*32726*/;
  assign _890_ = ~q[30] /*32725*/;
  assign _891_ = sum_2[60] & q[30] /*32724*/;
  assign _892_ = m_2[60] & _890_ /*32723*/;
  assign r_2[60] = _892_ | _891_ /*32722*/;
  assign _893_ = ~q[30] /*32721*/;
  assign _894_ = sum_2[61] & q[30] /*32720*/;
  assign _895_ = m_2[61] & _893_ /*32719*/;
  assign r_2[61] = _895_ | _894_ /*32718*/;
  assign _896_ = ~q[30] /*32717*/;
  assign _897_ = sum_2[62] & q[30] /*32716*/;
  assign _898_ = m_2[62] & _896_ /*32715*/;
  assign r_2[62] = _898_ | _897_ /*32714*/;
  assign _899_ = ~q[30] /*32713*/;
  assign _900_ = sum_2[63] & q[30] /*32712*/;
  assign _901_ = m_2[63] & _899_ /*32711*/;
  assign r_2[63] = _901_ | _900_ /*32710*/;
  assign _902_ = ~q[30] /*32709*/;
  assign _903_ = sum_2[64] & q[30] /*32708*/;
  assign _904_ = m_2[64] & _902_ /*32707*/;
  assign r_2[64] = _904_ | _903_ /*32706*/;
  assign inv_3[0] = oneWire /*32344*/;
  assign inv_3[1] = oneWire /*32338*/;
  assign inv_3[2] = oneWire /*32332*/;
  assign inv_3[3] = oneWire /*32326*/;
  assign inv_3[4] = oneWire /*32320*/;
  assign inv_3[5] = oneWire /*32314*/;
  assign inv_3[6] = oneWire /*32308*/;
  assign inv_3[7] = oneWire /*32302*/;
  assign inv_3[8] = oneWire /*32296*/;
  assign inv_3[9] = oneWire /*32290*/;
  assign inv_3[10] = oneWire /*32284*/;
  assign inv_3[11] = oneWire /*32278*/;
  assign inv_3[12] = oneWire /*32272*/;
  assign inv_3[13] = oneWire /*32266*/;
  assign inv_3[14] = oneWire /*32260*/;
  assign inv_3[15] = oneWire /*32254*/;
  assign inv_3[16] = oneWire /*32248*/;
  assign inv_3[17] = oneWire /*32242*/;
  assign inv_3[18] = oneWire /*32236*/;
  assign inv_3[19] = oneWire /*32230*/;
  assign inv_3[20] = oneWire /*32224*/;
  assign inv_3[21] = oneWire /*32218*/;
  assign inv_3[22] = oneWire /*32212*/;
  assign inv_3[23] = oneWire /*32206*/;
  assign inv_3[24] = oneWire /*32200*/;
  assign inv_3[25] = oneWire /*32194*/;
  assign inv_3[26] = oneWire /*32188*/;
  assign inv_3[27] = oneWire /*32182*/;
  assign inv_3[28] = oneWire /*32176*/;
  assign inv_3[29] = ~div[0] /*32170*/;
  assign inv_3[30] = ~div[1] /*32164*/;
  assign inv_3[31] = ~div[2] /*32158*/;
  assign inv_3[32] = ~div[3] /*32152*/;
  assign inv_3[33] = ~div[4] /*32146*/;
  assign inv_3[34] = ~div[5] /*32140*/;
  assign inv_3[35] = ~div[6] /*32134*/;
  assign inv_3[36] = ~div[7] /*32128*/;
  assign inv_3[37] = ~div[8] /*32122*/;
  assign inv_3[38] = ~div[9] /*32116*/;
  assign inv_3[39] = ~div[10] /*32110*/;
  assign inv_3[40] = ~div[11] /*32104*/;
  assign inv_3[41] = ~div[12] /*32098*/;
  assign inv_3[42] = ~div[13] /*32092*/;
  assign inv_3[43] = ~div[14] /*32086*/;
  assign inv_3[44] = ~div[15] /*32080*/;
  assign inv_3[45] = ~div[16] /*32074*/;
  assign inv_3[46] = ~div[17] /*32068*/;
  assign inv_3[47] = ~div[18] /*32062*/;
  assign inv_3[48] = ~div[19] /*32056*/;
  assign inv_3[49] = ~div[20] /*32050*/;
  assign inv_3[50] = ~div[21] /*32044*/;
  assign inv_3[51] = ~div[22] /*32038*/;
  assign inv_3[52] = ~div[23] /*32032*/;
  assign inv_3[53] = ~div[24] /*32026*/;
  assign inv_3[54] = ~div[25] /*32020*/;
  assign inv_3[55] = ~div[26] /*32014*/;
  assign inv_3[56] = ~div[27] /*32008*/;
  assign inv_3[57] = ~div[28] /*32002*/;
  assign inv_3[58] = ~div[29] /*31996*/;
  assign inv_3[59] = ~div[30] /*31990*/;
  assign inv_3[60] = oneWire /*31984*/;
  assign inv_3[61] = oneWire /*31978*/;
  assign inv_3[62] = oneWire /*31972*/;
  assign inv_3[63] = oneWire /*31966*/;
  assign inv_3[64] = oneWire /*31960*/;
  assign _905_ = inv_3[0] ^ r_2[0] /*32343*/;
  assign sum_3[0] = _905_ ^ oneWire /*32342*/;
  assign _906_ = _905_ & oneWire /*32341*/;
  assign _907_ = inv_3[0] & r_2[0] /*32340*/;
  assign _908_ = _906_ | _907_ /*32339*/;
  assign _909_ = inv_3[1] ^ r_2[1] /*32337*/;
  assign sum_3[1] = _909_ ^ _908_ /*32336*/;
  assign _910_ = _909_ & _908_ /*32335*/;
  assign _911_ = inv_3[1] & r_2[1] /*32334*/;
  assign _912_ = _910_ | _911_ /*32333*/;
  assign _913_ = inv_3[2] ^ r_2[2] /*32331*/;
  assign sum_3[2] = _913_ ^ _912_ /*32330*/;
  assign _914_ = _913_ & _912_ /*32329*/;
  assign _915_ = inv_3[2] & r_2[2] /*32328*/;
  assign _916_ = _914_ | _915_ /*32327*/;
  assign _917_ = inv_3[3] ^ r_2[3] /*32325*/;
  assign sum_3[3] = _917_ ^ _916_ /*32324*/;
  assign _918_ = _917_ & _916_ /*32323*/;
  assign _919_ = inv_3[3] & r_2[3] /*32322*/;
  assign _920_ = _918_ | _919_ /*32321*/;
  assign _921_ = inv_3[4] ^ r_2[4] /*32319*/;
  assign sum_3[4] = _921_ ^ _920_ /*32318*/;
  assign _922_ = _921_ & _920_ /*32317*/;
  assign _923_ = inv_3[4] & r_2[4] /*32316*/;
  assign _924_ = _922_ | _923_ /*32315*/;
  assign _925_ = inv_3[5] ^ r_2[5] /*32313*/;
  assign sum_3[5] = _925_ ^ _924_ /*32312*/;
  assign _926_ = _925_ & _924_ /*32311*/;
  assign _927_ = inv_3[5] & r_2[5] /*32310*/;
  assign _928_ = _926_ | _927_ /*32309*/;
  assign _929_ = inv_3[6] ^ r_2[6] /*32307*/;
  assign sum_3[6] = _929_ ^ _928_ /*32306*/;
  assign _930_ = _929_ & _928_ /*32305*/;
  assign _931_ = inv_3[6] & r_2[6] /*32304*/;
  assign _932_ = _930_ | _931_ /*32303*/;
  assign _933_ = inv_3[7] ^ r_2[7] /*32301*/;
  assign sum_3[7] = _933_ ^ _932_ /*32300*/;
  assign _934_ = _933_ & _932_ /*32299*/;
  assign _935_ = inv_3[7] & r_2[7] /*32298*/;
  assign _936_ = _934_ | _935_ /*32297*/;
  assign _937_ = inv_3[8] ^ r_2[8] /*32295*/;
  assign sum_3[8] = _937_ ^ _936_ /*32294*/;
  assign _938_ = _937_ & _936_ /*32293*/;
  assign _939_ = inv_3[8] & r_2[8] /*32292*/;
  assign _940_ = _938_ | _939_ /*32291*/;
  assign _941_ = inv_3[9] ^ r_2[9] /*32289*/;
  assign sum_3[9] = _941_ ^ _940_ /*32288*/;
  assign _942_ = _941_ & _940_ /*32287*/;
  assign _943_ = inv_3[9] & r_2[9] /*32286*/;
  assign _944_ = _942_ | _943_ /*32285*/;
  assign _945_ = inv_3[10] ^ r_2[10] /*32283*/;
  assign sum_3[10] = _945_ ^ _944_ /*32282*/;
  assign _946_ = _945_ & _944_ /*32281*/;
  assign _947_ = inv_3[10] & r_2[10] /*32280*/;
  assign _948_ = _946_ | _947_ /*32279*/;
  assign _949_ = inv_3[11] ^ r_2[11] /*32277*/;
  assign sum_3[11] = _949_ ^ _948_ /*32276*/;
  assign _950_ = _949_ & _948_ /*32275*/;
  assign _951_ = inv_3[11] & r_2[11] /*32274*/;
  assign _952_ = _950_ | _951_ /*32273*/;
  assign _953_ = inv_3[12] ^ r_2[12] /*32271*/;
  assign sum_3[12] = _953_ ^ _952_ /*32270*/;
  assign _954_ = _953_ & _952_ /*32269*/;
  assign _955_ = inv_3[12] & r_2[12] /*32268*/;
  assign _956_ = _954_ | _955_ /*32267*/;
  assign _957_ = inv_3[13] ^ r_2[13] /*32265*/;
  assign sum_3[13] = _957_ ^ _956_ /*32264*/;
  assign _958_ = _957_ & _956_ /*32263*/;
  assign _959_ = inv_3[13] & r_2[13] /*32262*/;
  assign _960_ = _958_ | _959_ /*32261*/;
  assign _961_ = inv_3[14] ^ r_2[14] /*32259*/;
  assign sum_3[14] = _961_ ^ _960_ /*32258*/;
  assign _962_ = _961_ & _960_ /*32257*/;
  assign _963_ = inv_3[14] & r_2[14] /*32256*/;
  assign _964_ = _962_ | _963_ /*32255*/;
  assign _965_ = inv_3[15] ^ r_2[15] /*32253*/;
  assign sum_3[15] = _965_ ^ _964_ /*32252*/;
  assign _966_ = _965_ & _964_ /*32251*/;
  assign _967_ = inv_3[15] & r_2[15] /*32250*/;
  assign _968_ = _966_ | _967_ /*32249*/;
  assign _969_ = inv_3[16] ^ r_2[16] /*32247*/;
  assign sum_3[16] = _969_ ^ _968_ /*32246*/;
  assign _970_ = _969_ & _968_ /*32245*/;
  assign _971_ = inv_3[16] & r_2[16] /*32244*/;
  assign _972_ = _970_ | _971_ /*32243*/;
  assign _973_ = inv_3[17] ^ r_2[17] /*32241*/;
  assign sum_3[17] = _973_ ^ _972_ /*32240*/;
  assign _974_ = _973_ & _972_ /*32239*/;
  assign _975_ = inv_3[17] & r_2[17] /*32238*/;
  assign _976_ = _974_ | _975_ /*32237*/;
  assign _977_ = inv_3[18] ^ r_2[18] /*32235*/;
  assign sum_3[18] = _977_ ^ _976_ /*32234*/;
  assign _978_ = _977_ & _976_ /*32233*/;
  assign _979_ = inv_3[18] & r_2[18] /*32232*/;
  assign _980_ = _978_ | _979_ /*32231*/;
  assign _981_ = inv_3[19] ^ r_2[19] /*32229*/;
  assign sum_3[19] = _981_ ^ _980_ /*32228*/;
  assign _982_ = _981_ & _980_ /*32227*/;
  assign _983_ = inv_3[19] & r_2[19] /*32226*/;
  assign _984_ = _982_ | _983_ /*32225*/;
  assign _985_ = inv_3[20] ^ r_2[20] /*32223*/;
  assign sum_3[20] = _985_ ^ _984_ /*32222*/;
  assign _986_ = _985_ & _984_ /*32221*/;
  assign _987_ = inv_3[20] & r_2[20] /*32220*/;
  assign _988_ = _986_ | _987_ /*32219*/;
  assign _989_ = inv_3[21] ^ r_2[21] /*32217*/;
  assign sum_3[21] = _989_ ^ _988_ /*32216*/;
  assign _990_ = _989_ & _988_ /*32215*/;
  assign _991_ = inv_3[21] & r_2[21] /*32214*/;
  assign _992_ = _990_ | _991_ /*32213*/;
  assign _993_ = inv_3[22] ^ r_2[22] /*32211*/;
  assign sum_3[22] = _993_ ^ _992_ /*32210*/;
  assign _994_ = _993_ & _992_ /*32209*/;
  assign _995_ = inv_3[22] & r_2[22] /*32208*/;
  assign _996_ = _994_ | _995_ /*32207*/;
  assign _997_ = inv_3[23] ^ r_2[23] /*32205*/;
  assign sum_3[23] = _997_ ^ _996_ /*32204*/;
  assign _998_ = _997_ & _996_ /*32203*/;
  assign _999_ = inv_3[23] & r_2[23] /*32202*/;
  assign _1000_ = _998_ | _999_ /*32201*/;
  assign _1001_ = inv_3[24] ^ r_2[24] /*32199*/;
  assign sum_3[24] = _1001_ ^ _1000_ /*32198*/;
  assign _1002_ = _1001_ & _1000_ /*32197*/;
  assign _1003_ = inv_3[24] & r_2[24] /*32196*/;
  assign _1004_ = _1002_ | _1003_ /*32195*/;
  assign _1005_ = inv_3[25] ^ r_2[25] /*32193*/;
  assign sum_3[25] = _1005_ ^ _1004_ /*32192*/;
  assign _1006_ = _1005_ & _1004_ /*32191*/;
  assign _1007_ = inv_3[25] & r_2[25] /*32190*/;
  assign _1008_ = _1006_ | _1007_ /*32189*/;
  assign _1009_ = inv_3[26] ^ r_2[26] /*32187*/;
  assign sum_3[26] = _1009_ ^ _1008_ /*32186*/;
  assign _1010_ = _1009_ & _1008_ /*32185*/;
  assign _1011_ = inv_3[26] & r_2[26] /*32184*/;
  assign _1012_ = _1010_ | _1011_ /*32183*/;
  assign _1013_ = inv_3[27] ^ r_2[27] /*32181*/;
  assign sum_3[27] = _1013_ ^ _1012_ /*32180*/;
  assign _1014_ = _1013_ & _1012_ /*32179*/;
  assign _1015_ = inv_3[27] & r_2[27] /*32178*/;
  assign _1016_ = _1014_ | _1015_ /*32177*/;
  assign _1017_ = inv_3[28] ^ r_2[28] /*32175*/;
  assign sum_3[28] = _1017_ ^ _1016_ /*32174*/;
  assign _1018_ = _1017_ & _1016_ /*32173*/;
  assign _1019_ = inv_3[28] & r_2[28] /*32172*/;
  assign _1020_ = _1018_ | _1019_ /*32171*/;
  assign _1021_ = inv_3[29] ^ r_2[29] /*32169*/;
  assign sum_3[29] = _1021_ ^ _1020_ /*32168*/;
  assign _1022_ = _1021_ & _1020_ /*32167*/;
  assign _1023_ = inv_3[29] & r_2[29] /*32166*/;
  assign _1024_ = _1022_ | _1023_ /*32165*/;
  assign _1025_ = inv_3[30] ^ r_2[30] /*32163*/;
  assign sum_3[30] = _1025_ ^ _1024_ /*32162*/;
  assign _1026_ = _1025_ & _1024_ /*32161*/;
  assign _1027_ = inv_3[30] & r_2[30] /*32160*/;
  assign _1028_ = _1026_ | _1027_ /*32159*/;
  assign _1029_ = inv_3[31] ^ r_2[31] /*32157*/;
  assign sum_3[31] = _1029_ ^ _1028_ /*32156*/;
  assign _1030_ = _1029_ & _1028_ /*32155*/;
  assign _1031_ = inv_3[31] & r_2[31] /*32154*/;
  assign _1032_ = _1030_ | _1031_ /*32153*/;
  assign _1033_ = inv_3[32] ^ r_2[32] /*32151*/;
  assign sum_3[32] = _1033_ ^ _1032_ /*32150*/;
  assign _1034_ = _1033_ & _1032_ /*32149*/;
  assign _1035_ = inv_3[32] & r_2[32] /*32148*/;
  assign _1036_ = _1034_ | _1035_ /*32147*/;
  assign _1037_ = inv_3[33] ^ r_2[33] /*32145*/;
  assign sum_3[33] = _1037_ ^ _1036_ /*32144*/;
  assign _1038_ = _1037_ & _1036_ /*32143*/;
  assign _1039_ = inv_3[33] & r_2[33] /*32142*/;
  assign _1040_ = _1038_ | _1039_ /*32141*/;
  assign _1041_ = inv_3[34] ^ r_2[34] /*32139*/;
  assign sum_3[34] = _1041_ ^ _1040_ /*32138*/;
  assign _1042_ = _1041_ & _1040_ /*32137*/;
  assign _1043_ = inv_3[34] & r_2[34] /*32136*/;
  assign _1044_ = _1042_ | _1043_ /*32135*/;
  assign _1045_ = inv_3[35] ^ r_2[35] /*32133*/;
  assign sum_3[35] = _1045_ ^ _1044_ /*32132*/;
  assign _1046_ = _1045_ & _1044_ /*32131*/;
  assign _1047_ = inv_3[35] & r_2[35] /*32130*/;
  assign _1048_ = _1046_ | _1047_ /*32129*/;
  assign _1049_ = inv_3[36] ^ r_2[36] /*32127*/;
  assign sum_3[36] = _1049_ ^ _1048_ /*32126*/;
  assign _1050_ = _1049_ & _1048_ /*32125*/;
  assign _1051_ = inv_3[36] & r_2[36] /*32124*/;
  assign _1052_ = _1050_ | _1051_ /*32123*/;
  assign _1053_ = inv_3[37] ^ r_2[37] /*32121*/;
  assign sum_3[37] = _1053_ ^ _1052_ /*32120*/;
  assign _1054_ = _1053_ & _1052_ /*32119*/;
  assign _1055_ = inv_3[37] & r_2[37] /*32118*/;
  assign _1056_ = _1054_ | _1055_ /*32117*/;
  assign _1057_ = inv_3[38] ^ r_2[38] /*32115*/;
  assign sum_3[38] = _1057_ ^ _1056_ /*32114*/;
  assign _1058_ = _1057_ & _1056_ /*32113*/;
  assign _1059_ = inv_3[38] & r_2[38] /*32112*/;
  assign _1060_ = _1058_ | _1059_ /*32111*/;
  assign _1061_ = inv_3[39] ^ r_2[39] /*32109*/;
  assign sum_3[39] = _1061_ ^ _1060_ /*32108*/;
  assign _1062_ = _1061_ & _1060_ /*32107*/;
  assign _1063_ = inv_3[39] & r_2[39] /*32106*/;
  assign _1064_ = _1062_ | _1063_ /*32105*/;
  assign _1065_ = inv_3[40] ^ r_2[40] /*32103*/;
  assign sum_3[40] = _1065_ ^ _1064_ /*32102*/;
  assign _1066_ = _1065_ & _1064_ /*32101*/;
  assign _1067_ = inv_3[40] & r_2[40] /*32100*/;
  assign _1068_ = _1066_ | _1067_ /*32099*/;
  assign _1069_ = inv_3[41] ^ r_2[41] /*32097*/;
  assign sum_3[41] = _1069_ ^ _1068_ /*32096*/;
  assign _1070_ = _1069_ & _1068_ /*32095*/;
  assign _1071_ = inv_3[41] & r_2[41] /*32094*/;
  assign _1072_ = _1070_ | _1071_ /*32093*/;
  assign _1073_ = inv_3[42] ^ r_2[42] /*32091*/;
  assign sum_3[42] = _1073_ ^ _1072_ /*32090*/;
  assign _1074_ = _1073_ & _1072_ /*32089*/;
  assign _1075_ = inv_3[42] & r_2[42] /*32088*/;
  assign _1076_ = _1074_ | _1075_ /*32087*/;
  assign _1077_ = inv_3[43] ^ r_2[43] /*32085*/;
  assign sum_3[43] = _1077_ ^ _1076_ /*32084*/;
  assign _1078_ = _1077_ & _1076_ /*32083*/;
  assign _1079_ = inv_3[43] & r_2[43] /*32082*/;
  assign _1080_ = _1078_ | _1079_ /*32081*/;
  assign _1081_ = inv_3[44] ^ r_2[44] /*32079*/;
  assign sum_3[44] = _1081_ ^ _1080_ /*32078*/;
  assign _1082_ = _1081_ & _1080_ /*32077*/;
  assign _1083_ = inv_3[44] & r_2[44] /*32076*/;
  assign _1084_ = _1082_ | _1083_ /*32075*/;
  assign _1085_ = inv_3[45] ^ r_2[45] /*32073*/;
  assign sum_3[45] = _1085_ ^ _1084_ /*32072*/;
  assign _1086_ = _1085_ & _1084_ /*32071*/;
  assign _1087_ = inv_3[45] & r_2[45] /*32070*/;
  assign _1088_ = _1086_ | _1087_ /*32069*/;
  assign _1089_ = inv_3[46] ^ r_2[46] /*32067*/;
  assign sum_3[46] = _1089_ ^ _1088_ /*32066*/;
  assign _1090_ = _1089_ & _1088_ /*32065*/;
  assign _1091_ = inv_3[46] & r_2[46] /*32064*/;
  assign _1092_ = _1090_ | _1091_ /*32063*/;
  assign _1093_ = inv_3[47] ^ r_2[47] /*32061*/;
  assign sum_3[47] = _1093_ ^ _1092_ /*32060*/;
  assign _1094_ = _1093_ & _1092_ /*32059*/;
  assign _1095_ = inv_3[47] & r_2[47] /*32058*/;
  assign _1096_ = _1094_ | _1095_ /*32057*/;
  assign _1097_ = inv_3[48] ^ r_2[48] /*32055*/;
  assign sum_3[48] = _1097_ ^ _1096_ /*32054*/;
  assign _1098_ = _1097_ & _1096_ /*32053*/;
  assign _1099_ = inv_3[48] & r_2[48] /*32052*/;
  assign _1100_ = _1098_ | _1099_ /*32051*/;
  assign _1101_ = inv_3[49] ^ r_2[49] /*32049*/;
  assign sum_3[49] = _1101_ ^ _1100_ /*32048*/;
  assign _1102_ = _1101_ & _1100_ /*32047*/;
  assign _1103_ = inv_3[49] & r_2[49] /*32046*/;
  assign _1104_ = _1102_ | _1103_ /*32045*/;
  assign _1105_ = inv_3[50] ^ r_2[50] /*32043*/;
  assign sum_3[50] = _1105_ ^ _1104_ /*32042*/;
  assign _1106_ = _1105_ & _1104_ /*32041*/;
  assign _1107_ = inv_3[50] & r_2[50] /*32040*/;
  assign _1108_ = _1106_ | _1107_ /*32039*/;
  assign _1109_ = inv_3[51] ^ r_2[51] /*32037*/;
  assign sum_3[51] = _1109_ ^ _1108_ /*32036*/;
  assign _1110_ = _1109_ & _1108_ /*32035*/;
  assign _1111_ = inv_3[51] & r_2[51] /*32034*/;
  assign _1112_ = _1110_ | _1111_ /*32033*/;
  assign _1113_ = inv_3[52] ^ r_2[52] /*32031*/;
  assign sum_3[52] = _1113_ ^ _1112_ /*32030*/;
  assign _1114_ = _1113_ & _1112_ /*32029*/;
  assign _1115_ = inv_3[52] & r_2[52] /*32028*/;
  assign _1116_ = _1114_ | _1115_ /*32027*/;
  assign _1117_ = inv_3[53] ^ r_2[53] /*32025*/;
  assign sum_3[53] = _1117_ ^ _1116_ /*32024*/;
  assign _1118_ = _1117_ & _1116_ /*32023*/;
  assign _1119_ = inv_3[53] & r_2[53] /*32022*/;
  assign _1120_ = _1118_ | _1119_ /*32021*/;
  assign _1121_ = inv_3[54] ^ r_2[54] /*32019*/;
  assign sum_3[54] = _1121_ ^ _1120_ /*32018*/;
  assign _1122_ = _1121_ & _1120_ /*32017*/;
  assign _1123_ = inv_3[54] & r_2[54] /*32016*/;
  assign _1124_ = _1122_ | _1123_ /*32015*/;
  assign _1125_ = inv_3[55] ^ r_2[55] /*32013*/;
  assign sum_3[55] = _1125_ ^ _1124_ /*32012*/;
  assign _1126_ = _1125_ & _1124_ /*32011*/;
  assign _1127_ = inv_3[55] & r_2[55] /*32010*/;
  assign _1128_ = _1126_ | _1127_ /*32009*/;
  assign _1129_ = inv_3[56] ^ r_2[56] /*32007*/;
  assign sum_3[56] = _1129_ ^ _1128_ /*32006*/;
  assign _1130_ = _1129_ & _1128_ /*32005*/;
  assign _1131_ = inv_3[56] & r_2[56] /*32004*/;
  assign _1132_ = _1130_ | _1131_ /*32003*/;
  assign _1133_ = inv_3[57] ^ r_2[57] /*32001*/;
  assign sum_3[57] = _1133_ ^ _1132_ /*32000*/;
  assign _1134_ = _1133_ & _1132_ /*31999*/;
  assign _1135_ = inv_3[57] & r_2[57] /*31998*/;
  assign _1136_ = _1134_ | _1135_ /*31997*/;
  assign _1137_ = inv_3[58] ^ r_2[58] /*31995*/;
  assign sum_3[58] = _1137_ ^ _1136_ /*31994*/;
  assign _1138_ = _1137_ & _1136_ /*31993*/;
  assign _1139_ = inv_3[58] & r_2[58] /*31992*/;
  assign _1140_ = _1138_ | _1139_ /*31991*/;
  assign _1141_ = inv_3[59] ^ r_2[59] /*31989*/;
  assign sum_3[59] = _1141_ ^ _1140_ /*31988*/;
  assign _1142_ = _1141_ & _1140_ /*31987*/;
  assign _1143_ = inv_3[59] & r_2[59] /*31986*/;
  assign _1144_ = _1142_ | _1143_ /*31985*/;
  assign _1145_ = inv_3[60] ^ r_2[60] /*31983*/;
  assign sum_3[60] = _1145_ ^ _1144_ /*31982*/;
  assign _1146_ = _1145_ & _1144_ /*31981*/;
  assign _1147_ = inv_3[60] & r_2[60] /*31980*/;
  assign _1148_ = _1146_ | _1147_ /*31979*/;
  assign _1149_ = inv_3[61] ^ r_2[61] /*31977*/;
  assign sum_3[61] = _1149_ ^ _1148_ /*31976*/;
  assign _1150_ = _1149_ & _1148_ /*31975*/;
  assign _1151_ = inv_3[61] & r_2[61] /*31974*/;
  assign _1152_ = _1150_ | _1151_ /*31973*/;
  assign _1153_ = inv_3[62] ^ r_2[62] /*31971*/;
  assign sum_3[62] = _1153_ ^ _1152_ /*31970*/;
  assign _1154_ = _1153_ & _1152_ /*31969*/;
  assign _1155_ = inv_3[62] & r_2[62] /*31968*/;
  assign _1156_ = _1154_ | _1155_ /*31967*/;
  assign _1157_ = inv_3[63] ^ r_2[63] /*31965*/;
  assign sum_3[63] = _1157_ ^ _1156_ /*31964*/;
  assign _1158_ = _1157_ & _1156_ /*31963*/;
  assign _1159_ = inv_3[63] & r_2[63] /*31962*/;
  assign _1160_ = _1158_ | _1159_ /*31961*/;
  assign _1161_ = inv_3[64] ^ r_2[64] /*31959*/;
  assign sum_3[64] = _1161_ ^ _1160_ /*31958*/;
  assign _1162_ = _1161_ & _1160_ /*31957*/;
  assign _1163_ = inv_3[64] & r_2[64] /*31956*/;
  assign _1164_ = _1162_ | _1163_ /*31955*/;
  assign _1165_ = _1164_ ^ _1160_ /*31954*/;
  assign _1166_ = ~_1165_ /*31953*/;
  assign _1167_ = sum_3[64] & _1166_ /*31952*/;
  assign _1168_ = _1165_ & _1164_ /*31951*/;
  assign sum_3[65] = _1168_ | _1167_ /*31950*/;
  assign q[29] = ~sum_3[65] /*31949*/;
  assign m_3[0] = r_2[0] /*31948*/;
  assign m_3[1] = r_2[1] /*31947*/;
  assign m_3[2] = r_2[2] /*31946*/;
  assign m_3[3] = r_2[3] /*31945*/;
  assign m_3[4] = r_2[4] /*31944*/;
  assign m_3[5] = r_2[5] /*31943*/;
  assign m_3[6] = r_2[6] /*31942*/;
  assign m_3[7] = r_2[7] /*31941*/;
  assign m_3[8] = r_2[8] /*31940*/;
  assign m_3[9] = r_2[9] /*31939*/;
  assign m_3[10] = r_2[10] /*31938*/;
  assign m_3[11] = r_2[11] /*31937*/;
  assign m_3[12] = r_2[12] /*31936*/;
  assign m_3[13] = r_2[13] /*31935*/;
  assign m_3[14] = r_2[14] /*31934*/;
  assign m_3[15] = r_2[15] /*31933*/;
  assign m_3[16] = r_2[16] /*31932*/;
  assign m_3[17] = r_2[17] /*31931*/;
  assign m_3[18] = r_2[18] /*31930*/;
  assign m_3[19] = r_2[19] /*31929*/;
  assign m_3[20] = r_2[20] /*31928*/;
  assign m_3[21] = r_2[21] /*31927*/;
  assign m_3[22] = r_2[22] /*31926*/;
  assign m_3[23] = r_2[23] /*31925*/;
  assign m_3[24] = r_2[24] /*31924*/;
  assign m_3[25] = r_2[25] /*31923*/;
  assign m_3[26] = r_2[26] /*31922*/;
  assign m_3[27] = r_2[27] /*31921*/;
  assign m_3[28] = r_2[28] /*31920*/;
  assign m_3[29] = r_2[29] /*31919*/;
  assign m_3[30] = r_2[30] /*31918*/;
  assign m_3[31] = r_2[31] /*31917*/;
  assign m_3[32] = r_2[32] /*31916*/;
  assign m_3[33] = r_2[33] /*31915*/;
  assign m_3[34] = r_2[34] /*31914*/;
  assign m_3[35] = r_2[35] /*31913*/;
  assign m_3[36] = r_2[36] /*31912*/;
  assign m_3[37] = r_2[37] /*31911*/;
  assign m_3[38] = r_2[38] /*31910*/;
  assign m_3[39] = r_2[39] /*31909*/;
  assign m_3[40] = r_2[40] /*31908*/;
  assign m_3[41] = r_2[41] /*31907*/;
  assign m_3[42] = r_2[42] /*31906*/;
  assign m_3[43] = r_2[43] /*31905*/;
  assign m_3[44] = r_2[44] /*31904*/;
  assign m_3[45] = r_2[45] /*31903*/;
  assign m_3[46] = r_2[46] /*31902*/;
  assign m_3[47] = r_2[47] /*31901*/;
  assign m_3[48] = r_2[48] /*31900*/;
  assign m_3[49] = r_2[49] /*31899*/;
  assign m_3[50] = r_2[50] /*31898*/;
  assign m_3[51] = r_2[51] /*31897*/;
  assign m_3[52] = r_2[52] /*31896*/;
  assign m_3[53] = r_2[53] /*31895*/;
  assign m_3[54] = r_2[54] /*31894*/;
  assign m_3[55] = r_2[55] /*31893*/;
  assign m_3[56] = r_2[56] /*31892*/;
  assign m_3[57] = r_2[57] /*31891*/;
  assign m_3[58] = r_2[58] /*31890*/;
  assign m_3[59] = r_2[59] /*31889*/;
  assign m_3[60] = r_2[60] /*31888*/;
  assign m_3[61] = r_2[61] /*31887*/;
  assign m_3[62] = r_2[62] /*31886*/;
  assign m_3[63] = r_2[63] /*31885*/;
  assign m_3[64] = r_2[64] /*31884*/;
  assign m_3[65] = r_2[64] /*31883*/;
  assign _1170_ = ~q[29] /*31882*/;
  assign _1171_ = sum_3[0] & q[29] /*31881*/;
  assign _1172_ = m_3[0] & _1170_ /*31880*/;
  assign r_3[0] = _1172_ | _1171_ /*31879*/;
  assign _1173_ = ~q[29] /*31878*/;
  assign _1174_ = sum_3[1] & q[29] /*31877*/;
  assign _1175_ = m_3[1] & _1173_ /*31876*/;
  assign r_3[1] = _1175_ | _1174_ /*31875*/;
  assign _1176_ = ~q[29] /*31874*/;
  assign _1177_ = sum_3[2] & q[29] /*31873*/;
  assign _1178_ = m_3[2] & _1176_ /*31872*/;
  assign r_3[2] = _1178_ | _1177_ /*31871*/;
  assign _1179_ = ~q[29] /*31870*/;
  assign _1180_ = sum_3[3] & q[29] /*31869*/;
  assign _1181_ = m_3[3] & _1179_ /*31868*/;
  assign r_3[3] = _1181_ | _1180_ /*31867*/;
  assign _1182_ = ~q[29] /*31866*/;
  assign _1183_ = sum_3[4] & q[29] /*31865*/;
  assign _1184_ = m_3[4] & _1182_ /*31864*/;
  assign r_3[4] = _1184_ | _1183_ /*31863*/;
  assign _1185_ = ~q[29] /*31862*/;
  assign _1186_ = sum_3[5] & q[29] /*31861*/;
  assign _1187_ = m_3[5] & _1185_ /*31860*/;
  assign r_3[5] = _1187_ | _1186_ /*31859*/;
  assign _1188_ = ~q[29] /*31858*/;
  assign _1189_ = sum_3[6] & q[29] /*31857*/;
  assign _1190_ = m_3[6] & _1188_ /*31856*/;
  assign r_3[6] = _1190_ | _1189_ /*31855*/;
  assign _1191_ = ~q[29] /*31854*/;
  assign _1192_ = sum_3[7] & q[29] /*31853*/;
  assign _1193_ = m_3[7] & _1191_ /*31852*/;
  assign r_3[7] = _1193_ | _1192_ /*31851*/;
  assign _1194_ = ~q[29] /*31850*/;
  assign _1195_ = sum_3[8] & q[29] /*31849*/;
  assign _1196_ = m_3[8] & _1194_ /*31848*/;
  assign r_3[8] = _1196_ | _1195_ /*31847*/;
  assign _1197_ = ~q[29] /*31846*/;
  assign _1198_ = sum_3[9] & q[29] /*31845*/;
  assign _1199_ = m_3[9] & _1197_ /*31844*/;
  assign r_3[9] = _1199_ | _1198_ /*31843*/;
  assign _1200_ = ~q[29] /*31842*/;
  assign _1201_ = sum_3[10] & q[29] /*31841*/;
  assign _1202_ = m_3[10] & _1200_ /*31840*/;
  assign r_3[10] = _1202_ | _1201_ /*31839*/;
  assign _1203_ = ~q[29] /*31838*/;
  assign _1204_ = sum_3[11] & q[29] /*31837*/;
  assign _1205_ = m_3[11] & _1203_ /*31836*/;
  assign r_3[11] = _1205_ | _1204_ /*31835*/;
  assign _1206_ = ~q[29] /*31834*/;
  assign _1207_ = sum_3[12] & q[29] /*31833*/;
  assign _1208_ = m_3[12] & _1206_ /*31832*/;
  assign r_3[12] = _1208_ | _1207_ /*31831*/;
  assign _1209_ = ~q[29] /*31830*/;
  assign _1210_ = sum_3[13] & q[29] /*31829*/;
  assign _1211_ = m_3[13] & _1209_ /*31828*/;
  assign r_3[13] = _1211_ | _1210_ /*31827*/;
  assign _1212_ = ~q[29] /*31826*/;
  assign _1213_ = sum_3[14] & q[29] /*31825*/;
  assign _1214_ = m_3[14] & _1212_ /*31824*/;
  assign r_3[14] = _1214_ | _1213_ /*31823*/;
  assign _1215_ = ~q[29] /*31822*/;
  assign _1216_ = sum_3[15] & q[29] /*31821*/;
  assign _1217_ = m_3[15] & _1215_ /*31820*/;
  assign r_3[15] = _1217_ | _1216_ /*31819*/;
  assign _1218_ = ~q[29] /*31818*/;
  assign _1219_ = sum_3[16] & q[29] /*31817*/;
  assign _1220_ = m_3[16] & _1218_ /*31816*/;
  assign r_3[16] = _1220_ | _1219_ /*31815*/;
  assign _1221_ = ~q[29] /*31814*/;
  assign _1222_ = sum_3[17] & q[29] /*31813*/;
  assign _1223_ = m_3[17] & _1221_ /*31812*/;
  assign r_3[17] = _1223_ | _1222_ /*31811*/;
  assign _1224_ = ~q[29] /*31810*/;
  assign _1225_ = sum_3[18] & q[29] /*31809*/;
  assign _1226_ = m_3[18] & _1224_ /*31808*/;
  assign r_3[18] = _1226_ | _1225_ /*31807*/;
  assign _1227_ = ~q[29] /*31806*/;
  assign _1228_ = sum_3[19] & q[29] /*31805*/;
  assign _1229_ = m_3[19] & _1227_ /*31804*/;
  assign r_3[19] = _1229_ | _1228_ /*31803*/;
  assign _1230_ = ~q[29] /*31802*/;
  assign _1231_ = sum_3[20] & q[29] /*31801*/;
  assign _1232_ = m_3[20] & _1230_ /*31800*/;
  assign r_3[20] = _1232_ | _1231_ /*31799*/;
  assign _1233_ = ~q[29] /*31798*/;
  assign _1234_ = sum_3[21] & q[29] /*31797*/;
  assign _1235_ = m_3[21] & _1233_ /*31796*/;
  assign r_3[21] = _1235_ | _1234_ /*31795*/;
  assign _1236_ = ~q[29] /*31794*/;
  assign _1237_ = sum_3[22] & q[29] /*31793*/;
  assign _1238_ = m_3[22] & _1236_ /*31792*/;
  assign r_3[22] = _1238_ | _1237_ /*31791*/;
  assign _1239_ = ~q[29] /*31790*/;
  assign _1240_ = sum_3[23] & q[29] /*31789*/;
  assign _1241_ = m_3[23] & _1239_ /*31788*/;
  assign r_3[23] = _1241_ | _1240_ /*31787*/;
  assign _1242_ = ~q[29] /*31786*/;
  assign _1243_ = sum_3[24] & q[29] /*31785*/;
  assign _1244_ = m_3[24] & _1242_ /*31784*/;
  assign r_3[24] = _1244_ | _1243_ /*31783*/;
  assign _1245_ = ~q[29] /*31782*/;
  assign _1246_ = sum_3[25] & q[29] /*31781*/;
  assign _1247_ = m_3[25] & _1245_ /*31780*/;
  assign r_3[25] = _1247_ | _1246_ /*31779*/;
  assign _1248_ = ~q[29] /*31778*/;
  assign _1249_ = sum_3[26] & q[29] /*31777*/;
  assign _1250_ = m_3[26] & _1248_ /*31776*/;
  assign r_3[26] = _1250_ | _1249_ /*31775*/;
  assign _1251_ = ~q[29] /*31774*/;
  assign _1252_ = sum_3[27] & q[29] /*31773*/;
  assign _1253_ = m_3[27] & _1251_ /*31772*/;
  assign r_3[27] = _1253_ | _1252_ /*31771*/;
  assign _1254_ = ~q[29] /*31770*/;
  assign _1255_ = sum_3[28] & q[29] /*31769*/;
  assign _1256_ = m_3[28] & _1254_ /*31768*/;
  assign r_3[28] = _1256_ | _1255_ /*31767*/;
  assign _1257_ = ~q[29] /*31766*/;
  assign _1258_ = sum_3[29] & q[29] /*31765*/;
  assign _1259_ = m_3[29] & _1257_ /*31764*/;
  assign r_3[29] = _1259_ | _1258_ /*31763*/;
  assign _1260_ = ~q[29] /*31762*/;
  assign _1261_ = sum_3[30] & q[29] /*31761*/;
  assign _1262_ = m_3[30] & _1260_ /*31760*/;
  assign r_3[30] = _1262_ | _1261_ /*31759*/;
  assign _1263_ = ~q[29] /*31758*/;
  assign _1264_ = sum_3[31] & q[29] /*31757*/;
  assign _1265_ = m_3[31] & _1263_ /*31756*/;
  assign r_3[31] = _1265_ | _1264_ /*31755*/;
  assign _1266_ = ~q[29] /*31754*/;
  assign _1267_ = sum_3[32] & q[29] /*31753*/;
  assign _1268_ = m_3[32] & _1266_ /*31752*/;
  assign r_3[32] = _1268_ | _1267_ /*31751*/;
  assign _1269_ = ~q[29] /*31750*/;
  assign _1270_ = sum_3[33] & q[29] /*31749*/;
  assign _1271_ = m_3[33] & _1269_ /*31748*/;
  assign r_3[33] = _1271_ | _1270_ /*31747*/;
  assign _1272_ = ~q[29] /*31746*/;
  assign _1273_ = sum_3[34] & q[29] /*31745*/;
  assign _1274_ = m_3[34] & _1272_ /*31744*/;
  assign r_3[34] = _1274_ | _1273_ /*31743*/;
  assign _1275_ = ~q[29] /*31742*/;
  assign _1276_ = sum_3[35] & q[29] /*31741*/;
  assign _1277_ = m_3[35] & _1275_ /*31740*/;
  assign r_3[35] = _1277_ | _1276_ /*31739*/;
  assign _1278_ = ~q[29] /*31738*/;
  assign _1279_ = sum_3[36] & q[29] /*31737*/;
  assign _1280_ = m_3[36] & _1278_ /*31736*/;
  assign r_3[36] = _1280_ | _1279_ /*31735*/;
  assign _1281_ = ~q[29] /*31734*/;
  assign _1282_ = sum_3[37] & q[29] /*31733*/;
  assign _1283_ = m_3[37] & _1281_ /*31732*/;
  assign r_3[37] = _1283_ | _1282_ /*31731*/;
  assign _1284_ = ~q[29] /*31730*/;
  assign _1285_ = sum_3[38] & q[29] /*31729*/;
  assign _1286_ = m_3[38] & _1284_ /*31728*/;
  assign r_3[38] = _1286_ | _1285_ /*31727*/;
  assign _1287_ = ~q[29] /*31726*/;
  assign _1288_ = sum_3[39] & q[29] /*31725*/;
  assign _1289_ = m_3[39] & _1287_ /*31724*/;
  assign r_3[39] = _1289_ | _1288_ /*31723*/;
  assign _1290_ = ~q[29] /*31722*/;
  assign _1291_ = sum_3[40] & q[29] /*31721*/;
  assign _1292_ = m_3[40] & _1290_ /*31720*/;
  assign r_3[40] = _1292_ | _1291_ /*31719*/;
  assign _1293_ = ~q[29] /*31718*/;
  assign _1294_ = sum_3[41] & q[29] /*31717*/;
  assign _1295_ = m_3[41] & _1293_ /*31716*/;
  assign r_3[41] = _1295_ | _1294_ /*31715*/;
  assign _1296_ = ~q[29] /*31714*/;
  assign _1297_ = sum_3[42] & q[29] /*31713*/;
  assign _1298_ = m_3[42] & _1296_ /*31712*/;
  assign r_3[42] = _1298_ | _1297_ /*31711*/;
  assign _1299_ = ~q[29] /*31710*/;
  assign _1300_ = sum_3[43] & q[29] /*31709*/;
  assign _1301_ = m_3[43] & _1299_ /*31708*/;
  assign r_3[43] = _1301_ | _1300_ /*31707*/;
  assign _1302_ = ~q[29] /*31706*/;
  assign _1303_ = sum_3[44] & q[29] /*31705*/;
  assign _1304_ = m_3[44] & _1302_ /*31704*/;
  assign r_3[44] = _1304_ | _1303_ /*31703*/;
  assign _1305_ = ~q[29] /*31702*/;
  assign _1306_ = sum_3[45] & q[29] /*31701*/;
  assign _1307_ = m_3[45] & _1305_ /*31700*/;
  assign r_3[45] = _1307_ | _1306_ /*31699*/;
  assign _1308_ = ~q[29] /*31698*/;
  assign _1309_ = sum_3[46] & q[29] /*31697*/;
  assign _1310_ = m_3[46] & _1308_ /*31696*/;
  assign r_3[46] = _1310_ | _1309_ /*31695*/;
  assign _1311_ = ~q[29] /*31694*/;
  assign _1312_ = sum_3[47] & q[29] /*31693*/;
  assign _1313_ = m_3[47] & _1311_ /*31692*/;
  assign r_3[47] = _1313_ | _1312_ /*31691*/;
  assign _1314_ = ~q[29] /*31690*/;
  assign _1315_ = sum_3[48] & q[29] /*31689*/;
  assign _1316_ = m_3[48] & _1314_ /*31688*/;
  assign r_3[48] = _1316_ | _1315_ /*31687*/;
  assign _1317_ = ~q[29] /*31686*/;
  assign _1318_ = sum_3[49] & q[29] /*31685*/;
  assign _1319_ = m_3[49] & _1317_ /*31684*/;
  assign r_3[49] = _1319_ | _1318_ /*31683*/;
  assign _1320_ = ~q[29] /*31682*/;
  assign _1321_ = sum_3[50] & q[29] /*31681*/;
  assign _1322_ = m_3[50] & _1320_ /*31680*/;
  assign r_3[50] = _1322_ | _1321_ /*31679*/;
  assign _1323_ = ~q[29] /*31678*/;
  assign _1324_ = sum_3[51] & q[29] /*31677*/;
  assign _1325_ = m_3[51] & _1323_ /*31676*/;
  assign r_3[51] = _1325_ | _1324_ /*31675*/;
  assign _1326_ = ~q[29] /*31674*/;
  assign _1327_ = sum_3[52] & q[29] /*31673*/;
  assign _1328_ = m_3[52] & _1326_ /*31672*/;
  assign r_3[52] = _1328_ | _1327_ /*31671*/;
  assign _1329_ = ~q[29] /*31670*/;
  assign _1330_ = sum_3[53] & q[29] /*31669*/;
  assign _1331_ = m_3[53] & _1329_ /*31668*/;
  assign r_3[53] = _1331_ | _1330_ /*31667*/;
  assign _1332_ = ~q[29] /*31666*/;
  assign _1333_ = sum_3[54] & q[29] /*31665*/;
  assign _1334_ = m_3[54] & _1332_ /*31664*/;
  assign r_3[54] = _1334_ | _1333_ /*31663*/;
  assign _1335_ = ~q[29] /*31662*/;
  assign _1336_ = sum_3[55] & q[29] /*31661*/;
  assign _1337_ = m_3[55] & _1335_ /*31660*/;
  assign r_3[55] = _1337_ | _1336_ /*31659*/;
  assign _1338_ = ~q[29] /*31658*/;
  assign _1339_ = sum_3[56] & q[29] /*31657*/;
  assign _1340_ = m_3[56] & _1338_ /*31656*/;
  assign r_3[56] = _1340_ | _1339_ /*31655*/;
  assign _1341_ = ~q[29] /*31654*/;
  assign _1342_ = sum_3[57] & q[29] /*31653*/;
  assign _1343_ = m_3[57] & _1341_ /*31652*/;
  assign r_3[57] = _1343_ | _1342_ /*31651*/;
  assign _1344_ = ~q[29] /*31650*/;
  assign _1345_ = sum_3[58] & q[29] /*31649*/;
  assign _1346_ = m_3[58] & _1344_ /*31648*/;
  assign r_3[58] = _1346_ | _1345_ /*31647*/;
  assign _1347_ = ~q[29] /*31646*/;
  assign _1348_ = sum_3[59] & q[29] /*31645*/;
  assign _1349_ = m_3[59] & _1347_ /*31644*/;
  assign r_3[59] = _1349_ | _1348_ /*31643*/;
  assign _1350_ = ~q[29] /*31642*/;
  assign _1351_ = sum_3[60] & q[29] /*31641*/;
  assign _1352_ = m_3[60] & _1350_ /*31640*/;
  assign r_3[60] = _1352_ | _1351_ /*31639*/;
  assign _1353_ = ~q[29] /*31638*/;
  assign _1354_ = sum_3[61] & q[29] /*31637*/;
  assign _1355_ = m_3[61] & _1353_ /*31636*/;
  assign r_3[61] = _1355_ | _1354_ /*31635*/;
  assign _1356_ = ~q[29] /*31634*/;
  assign _1357_ = sum_3[62] & q[29] /*31633*/;
  assign _1358_ = m_3[62] & _1356_ /*31632*/;
  assign r_3[62] = _1358_ | _1357_ /*31631*/;
  assign _1359_ = ~q[29] /*31630*/;
  assign _1360_ = sum_3[63] & q[29] /*31629*/;
  assign _1361_ = m_3[63] & _1359_ /*31628*/;
  assign r_3[63] = _1361_ | _1360_ /*31627*/;
  assign _1362_ = ~q[29] /*31626*/;
  assign _1363_ = sum_3[64] & q[29] /*31625*/;
  assign _1364_ = m_3[64] & _1362_ /*31624*/;
  assign r_3[64] = _1364_ | _1363_ /*31623*/;
  assign _1365_ = ~q[29] /*31622*/;
  assign _1366_ = sum_3[65] & q[29] /*31621*/;
  assign _1367_ = m_3[65] & _1365_ /*31620*/;
  assign r_3[65] = _1367_ | _1366_ /*31619*/;
  assign inv_4[0] = oneWire /*31268*/;
  assign inv_4[1] = oneWire /*31262*/;
  assign inv_4[2] = oneWire /*31256*/;
  assign inv_4[3] = oneWire /*31250*/;
  assign inv_4[4] = oneWire /*31244*/;
  assign inv_4[5] = oneWire /*31238*/;
  assign inv_4[6] = oneWire /*31232*/;
  assign inv_4[7] = oneWire /*31226*/;
  assign inv_4[8] = oneWire /*31220*/;
  assign inv_4[9] = oneWire /*31214*/;
  assign inv_4[10] = oneWire /*31208*/;
  assign inv_4[11] = oneWire /*31202*/;
  assign inv_4[12] = oneWire /*31196*/;
  assign inv_4[13] = oneWire /*31190*/;
  assign inv_4[14] = oneWire /*31184*/;
  assign inv_4[15] = oneWire /*31178*/;
  assign inv_4[16] = oneWire /*31172*/;
  assign inv_4[17] = oneWire /*31166*/;
  assign inv_4[18] = oneWire /*31160*/;
  assign inv_4[19] = oneWire /*31154*/;
  assign inv_4[20] = oneWire /*31148*/;
  assign inv_4[21] = oneWire /*31142*/;
  assign inv_4[22] = oneWire /*31136*/;
  assign inv_4[23] = oneWire /*31130*/;
  assign inv_4[24] = oneWire /*31124*/;
  assign inv_4[25] = oneWire /*31118*/;
  assign inv_4[26] = oneWire /*31112*/;
  assign inv_4[27] = oneWire /*31106*/;
  assign inv_4[28] = ~div[0] /*31100*/;
  assign inv_4[29] = ~div[1] /*31094*/;
  assign inv_4[30] = ~div[2] /*31088*/;
  assign inv_4[31] = ~div[3] /*31082*/;
  assign inv_4[32] = ~div[4] /*31076*/;
  assign inv_4[33] = ~div[5] /*31070*/;
  assign inv_4[34] = ~div[6] /*31064*/;
  assign inv_4[35] = ~div[7] /*31058*/;
  assign inv_4[36] = ~div[8] /*31052*/;
  assign inv_4[37] = ~div[9] /*31046*/;
  assign inv_4[38] = ~div[10] /*31040*/;
  assign inv_4[39] = ~div[11] /*31034*/;
  assign inv_4[40] = ~div[12] /*31028*/;
  assign inv_4[41] = ~div[13] /*31022*/;
  assign inv_4[42] = ~div[14] /*31016*/;
  assign inv_4[43] = ~div[15] /*31010*/;
  assign inv_4[44] = ~div[16] /*31004*/;
  assign inv_4[45] = ~div[17] /*30998*/;
  assign inv_4[46] = ~div[18] /*30992*/;
  assign inv_4[47] = ~div[19] /*30986*/;
  assign inv_4[48] = ~div[20] /*30980*/;
  assign inv_4[49] = ~div[21] /*30974*/;
  assign inv_4[50] = ~div[22] /*30968*/;
  assign inv_4[51] = ~div[23] /*30962*/;
  assign inv_4[52] = ~div[24] /*30956*/;
  assign inv_4[53] = ~div[25] /*30950*/;
  assign inv_4[54] = ~div[26] /*30944*/;
  assign inv_4[55] = ~div[27] /*30938*/;
  assign inv_4[56] = ~div[28] /*30932*/;
  assign inv_4[57] = ~div[29] /*30926*/;
  assign inv_4[58] = ~div[30] /*30920*/;
  assign inv_4[59] = oneWire /*30914*/;
  assign inv_4[60] = oneWire /*30908*/;
  assign inv_4[61] = oneWire /*30902*/;
  assign inv_4[62] = oneWire /*30896*/;
  assign inv_4[63] = oneWire /*30890*/;
  assign inv_4[64] = oneWire /*30884*/;
  assign inv_4[65] = oneWire /*30878*/;
  assign _1368_ = inv_4[0] ^ r_3[0] /*31267*/;
  assign sum_4[0] = _1368_ ^ oneWire /*31266*/;
  assign _1369_ = _1368_ & oneWire /*31265*/;
  assign _1370_ = inv_4[0] & r_3[0] /*31264*/;
  assign _1371_ = _1369_ | _1370_ /*31263*/;
  assign _1372_ = inv_4[1] ^ r_3[1] /*31261*/;
  assign sum_4[1] = _1372_ ^ _1371_ /*31260*/;
  assign _1373_ = _1372_ & _1371_ /*31259*/;
  assign _1374_ = inv_4[1] & r_3[1] /*31258*/;
  assign _1375_ = _1373_ | _1374_ /*31257*/;
  assign _1376_ = inv_4[2] ^ r_3[2] /*31255*/;
  assign sum_4[2] = _1376_ ^ _1375_ /*31254*/;
  assign _1377_ = _1376_ & _1375_ /*31253*/;
  assign _1378_ = inv_4[2] & r_3[2] /*31252*/;
  assign _1379_ = _1377_ | _1378_ /*31251*/;
  assign _1380_ = inv_4[3] ^ r_3[3] /*31249*/;
  assign sum_4[3] = _1380_ ^ _1379_ /*31248*/;
  assign _1381_ = _1380_ & _1379_ /*31247*/;
  assign _1382_ = inv_4[3] & r_3[3] /*31246*/;
  assign _1383_ = _1381_ | _1382_ /*31245*/;
  assign _1384_ = inv_4[4] ^ r_3[4] /*31243*/;
  assign sum_4[4] = _1384_ ^ _1383_ /*31242*/;
  assign _1385_ = _1384_ & _1383_ /*31241*/;
  assign _1386_ = inv_4[4] & r_3[4] /*31240*/;
  assign _1387_ = _1385_ | _1386_ /*31239*/;
  assign _1388_ = inv_4[5] ^ r_3[5] /*31237*/;
  assign sum_4[5] = _1388_ ^ _1387_ /*31236*/;
  assign _1389_ = _1388_ & _1387_ /*31235*/;
  assign _1390_ = inv_4[5] & r_3[5] /*31234*/;
  assign _1391_ = _1389_ | _1390_ /*31233*/;
  assign _1392_ = inv_4[6] ^ r_3[6] /*31231*/;
  assign sum_4[6] = _1392_ ^ _1391_ /*31230*/;
  assign _1393_ = _1392_ & _1391_ /*31229*/;
  assign _1394_ = inv_4[6] & r_3[6] /*31228*/;
  assign _1395_ = _1393_ | _1394_ /*31227*/;
  assign _1396_ = inv_4[7] ^ r_3[7] /*31225*/;
  assign sum_4[7] = _1396_ ^ _1395_ /*31224*/;
  assign _1397_ = _1396_ & _1395_ /*31223*/;
  assign _1398_ = inv_4[7] & r_3[7] /*31222*/;
  assign _1399_ = _1397_ | _1398_ /*31221*/;
  assign _1400_ = inv_4[8] ^ r_3[8] /*31219*/;
  assign sum_4[8] = _1400_ ^ _1399_ /*31218*/;
  assign _1401_ = _1400_ & _1399_ /*31217*/;
  assign _1402_ = inv_4[8] & r_3[8] /*31216*/;
  assign _1403_ = _1401_ | _1402_ /*31215*/;
  assign _1404_ = inv_4[9] ^ r_3[9] /*31213*/;
  assign sum_4[9] = _1404_ ^ _1403_ /*31212*/;
  assign _1405_ = _1404_ & _1403_ /*31211*/;
  assign _1406_ = inv_4[9] & r_3[9] /*31210*/;
  assign _1407_ = _1405_ | _1406_ /*31209*/;
  assign _1408_ = inv_4[10] ^ r_3[10] /*31207*/;
  assign sum_4[10] = _1408_ ^ _1407_ /*31206*/;
  assign _1409_ = _1408_ & _1407_ /*31205*/;
  assign _1410_ = inv_4[10] & r_3[10] /*31204*/;
  assign _1411_ = _1409_ | _1410_ /*31203*/;
  assign _1412_ = inv_4[11] ^ r_3[11] /*31201*/;
  assign sum_4[11] = _1412_ ^ _1411_ /*31200*/;
  assign _1413_ = _1412_ & _1411_ /*31199*/;
  assign _1414_ = inv_4[11] & r_3[11] /*31198*/;
  assign _1415_ = _1413_ | _1414_ /*31197*/;
  assign _1416_ = inv_4[12] ^ r_3[12] /*31195*/;
  assign sum_4[12] = _1416_ ^ _1415_ /*31194*/;
  assign _1417_ = _1416_ & _1415_ /*31193*/;
  assign _1418_ = inv_4[12] & r_3[12] /*31192*/;
  assign _1419_ = _1417_ | _1418_ /*31191*/;
  assign _1420_ = inv_4[13] ^ r_3[13] /*31189*/;
  assign sum_4[13] = _1420_ ^ _1419_ /*31188*/;
  assign _1421_ = _1420_ & _1419_ /*31187*/;
  assign _1422_ = inv_4[13] & r_3[13] /*31186*/;
  assign _1423_ = _1421_ | _1422_ /*31185*/;
  assign _1424_ = inv_4[14] ^ r_3[14] /*31183*/;
  assign sum_4[14] = _1424_ ^ _1423_ /*31182*/;
  assign _1425_ = _1424_ & _1423_ /*31181*/;
  assign _1426_ = inv_4[14] & r_3[14] /*31180*/;
  assign _1427_ = _1425_ | _1426_ /*31179*/;
  assign _1428_ = inv_4[15] ^ r_3[15] /*31177*/;
  assign sum_4[15] = _1428_ ^ _1427_ /*31176*/;
  assign _1429_ = _1428_ & _1427_ /*31175*/;
  assign _1430_ = inv_4[15] & r_3[15] /*31174*/;
  assign _1431_ = _1429_ | _1430_ /*31173*/;
  assign _1432_ = inv_4[16] ^ r_3[16] /*31171*/;
  assign sum_4[16] = _1432_ ^ _1431_ /*31170*/;
  assign _1433_ = _1432_ & _1431_ /*31169*/;
  assign _1434_ = inv_4[16] & r_3[16] /*31168*/;
  assign _1435_ = _1433_ | _1434_ /*31167*/;
  assign _1436_ = inv_4[17] ^ r_3[17] /*31165*/;
  assign sum_4[17] = _1436_ ^ _1435_ /*31164*/;
  assign _1437_ = _1436_ & _1435_ /*31163*/;
  assign _1438_ = inv_4[17] & r_3[17] /*31162*/;
  assign _1439_ = _1437_ | _1438_ /*31161*/;
  assign _1440_ = inv_4[18] ^ r_3[18] /*31159*/;
  assign sum_4[18] = _1440_ ^ _1439_ /*31158*/;
  assign _1441_ = _1440_ & _1439_ /*31157*/;
  assign _1442_ = inv_4[18] & r_3[18] /*31156*/;
  assign _1443_ = _1441_ | _1442_ /*31155*/;
  assign _1444_ = inv_4[19] ^ r_3[19] /*31153*/;
  assign sum_4[19] = _1444_ ^ _1443_ /*31152*/;
  assign _1445_ = _1444_ & _1443_ /*31151*/;
  assign _1446_ = inv_4[19] & r_3[19] /*31150*/;
  assign _1447_ = _1445_ | _1446_ /*31149*/;
  assign _1448_ = inv_4[20] ^ r_3[20] /*31147*/;
  assign sum_4[20] = _1448_ ^ _1447_ /*31146*/;
  assign _1449_ = _1448_ & _1447_ /*31145*/;
  assign _1450_ = inv_4[20] & r_3[20] /*31144*/;
  assign _1451_ = _1449_ | _1450_ /*31143*/;
  assign _1452_ = inv_4[21] ^ r_3[21] /*31141*/;
  assign sum_4[21] = _1452_ ^ _1451_ /*31140*/;
  assign _1453_ = _1452_ & _1451_ /*31139*/;
  assign _1454_ = inv_4[21] & r_3[21] /*31138*/;
  assign _1455_ = _1453_ | _1454_ /*31137*/;
  assign _1456_ = inv_4[22] ^ r_3[22] /*31135*/;
  assign sum_4[22] = _1456_ ^ _1455_ /*31134*/;
  assign _1457_ = _1456_ & _1455_ /*31133*/;
  assign _1458_ = inv_4[22] & r_3[22] /*31132*/;
  assign _1459_ = _1457_ | _1458_ /*31131*/;
  assign _1460_ = inv_4[23] ^ r_3[23] /*31129*/;
  assign sum_4[23] = _1460_ ^ _1459_ /*31128*/;
  assign _1461_ = _1460_ & _1459_ /*31127*/;
  assign _1462_ = inv_4[23] & r_3[23] /*31126*/;
  assign _1463_ = _1461_ | _1462_ /*31125*/;
  assign _1464_ = inv_4[24] ^ r_3[24] /*31123*/;
  assign sum_4[24] = _1464_ ^ _1463_ /*31122*/;
  assign _1465_ = _1464_ & _1463_ /*31121*/;
  assign _1466_ = inv_4[24] & r_3[24] /*31120*/;
  assign _1467_ = _1465_ | _1466_ /*31119*/;
  assign _1468_ = inv_4[25] ^ r_3[25] /*31117*/;
  assign sum_4[25] = _1468_ ^ _1467_ /*31116*/;
  assign _1469_ = _1468_ & _1467_ /*31115*/;
  assign _1470_ = inv_4[25] & r_3[25] /*31114*/;
  assign _1471_ = _1469_ | _1470_ /*31113*/;
  assign _1472_ = inv_4[26] ^ r_3[26] /*31111*/;
  assign sum_4[26] = _1472_ ^ _1471_ /*31110*/;
  assign _1473_ = _1472_ & _1471_ /*31109*/;
  assign _1474_ = inv_4[26] & r_3[26] /*31108*/;
  assign _1475_ = _1473_ | _1474_ /*31107*/;
  assign _1476_ = inv_4[27] ^ r_3[27] /*31105*/;
  assign sum_4[27] = _1476_ ^ _1475_ /*31104*/;
  assign _1477_ = _1476_ & _1475_ /*31103*/;
  assign _1478_ = inv_4[27] & r_3[27] /*31102*/;
  assign _1479_ = _1477_ | _1478_ /*31101*/;
  assign _1480_ = inv_4[28] ^ r_3[28] /*31099*/;
  assign sum_4[28] = _1480_ ^ _1479_ /*31098*/;
  assign _1481_ = _1480_ & _1479_ /*31097*/;
  assign _1482_ = inv_4[28] & r_3[28] /*31096*/;
  assign _1483_ = _1481_ | _1482_ /*31095*/;
  assign _1484_ = inv_4[29] ^ r_3[29] /*31093*/;
  assign sum_4[29] = _1484_ ^ _1483_ /*31092*/;
  assign _1485_ = _1484_ & _1483_ /*31091*/;
  assign _1486_ = inv_4[29] & r_3[29] /*31090*/;
  assign _1487_ = _1485_ | _1486_ /*31089*/;
  assign _1488_ = inv_4[30] ^ r_3[30] /*31087*/;
  assign sum_4[30] = _1488_ ^ _1487_ /*31086*/;
  assign _1489_ = _1488_ & _1487_ /*31085*/;
  assign _1490_ = inv_4[30] & r_3[30] /*31084*/;
  assign _1491_ = _1489_ | _1490_ /*31083*/;
  assign _1492_ = inv_4[31] ^ r_3[31] /*31081*/;
  assign sum_4[31] = _1492_ ^ _1491_ /*31080*/;
  assign _1493_ = _1492_ & _1491_ /*31079*/;
  assign _1494_ = inv_4[31] & r_3[31] /*31078*/;
  assign _1495_ = _1493_ | _1494_ /*31077*/;
  assign _1496_ = inv_4[32] ^ r_3[32] /*31075*/;
  assign sum_4[32] = _1496_ ^ _1495_ /*31074*/;
  assign _1497_ = _1496_ & _1495_ /*31073*/;
  assign _1498_ = inv_4[32] & r_3[32] /*31072*/;
  assign _1499_ = _1497_ | _1498_ /*31071*/;
  assign _1500_ = inv_4[33] ^ r_3[33] /*31069*/;
  assign sum_4[33] = _1500_ ^ _1499_ /*31068*/;
  assign _1501_ = _1500_ & _1499_ /*31067*/;
  assign _1502_ = inv_4[33] & r_3[33] /*31066*/;
  assign _1503_ = _1501_ | _1502_ /*31065*/;
  assign _1504_ = inv_4[34] ^ r_3[34] /*31063*/;
  assign sum_4[34] = _1504_ ^ _1503_ /*31062*/;
  assign _1505_ = _1504_ & _1503_ /*31061*/;
  assign _1506_ = inv_4[34] & r_3[34] /*31060*/;
  assign _1507_ = _1505_ | _1506_ /*31059*/;
  assign _1508_ = inv_4[35] ^ r_3[35] /*31057*/;
  assign sum_4[35] = _1508_ ^ _1507_ /*31056*/;
  assign _1509_ = _1508_ & _1507_ /*31055*/;
  assign _1510_ = inv_4[35] & r_3[35] /*31054*/;
  assign _1511_ = _1509_ | _1510_ /*31053*/;
  assign _1512_ = inv_4[36] ^ r_3[36] /*31051*/;
  assign sum_4[36] = _1512_ ^ _1511_ /*31050*/;
  assign _1513_ = _1512_ & _1511_ /*31049*/;
  assign _1514_ = inv_4[36] & r_3[36] /*31048*/;
  assign _1515_ = _1513_ | _1514_ /*31047*/;
  assign _1516_ = inv_4[37] ^ r_3[37] /*31045*/;
  assign sum_4[37] = _1516_ ^ _1515_ /*31044*/;
  assign _1517_ = _1516_ & _1515_ /*31043*/;
  assign _1518_ = inv_4[37] & r_3[37] /*31042*/;
  assign _1519_ = _1517_ | _1518_ /*31041*/;
  assign _1520_ = inv_4[38] ^ r_3[38] /*31039*/;
  assign sum_4[38] = _1520_ ^ _1519_ /*31038*/;
  assign _1521_ = _1520_ & _1519_ /*31037*/;
  assign _1522_ = inv_4[38] & r_3[38] /*31036*/;
  assign _1523_ = _1521_ | _1522_ /*31035*/;
  assign _1524_ = inv_4[39] ^ r_3[39] /*31033*/;
  assign sum_4[39] = _1524_ ^ _1523_ /*31032*/;
  assign _1525_ = _1524_ & _1523_ /*31031*/;
  assign _1526_ = inv_4[39] & r_3[39] /*31030*/;
  assign _1527_ = _1525_ | _1526_ /*31029*/;
  assign _1528_ = inv_4[40] ^ r_3[40] /*31027*/;
  assign sum_4[40] = _1528_ ^ _1527_ /*31026*/;
  assign _1529_ = _1528_ & _1527_ /*31025*/;
  assign _1530_ = inv_4[40] & r_3[40] /*31024*/;
  assign _1531_ = _1529_ | _1530_ /*31023*/;
  assign _1532_ = inv_4[41] ^ r_3[41] /*31021*/;
  assign sum_4[41] = _1532_ ^ _1531_ /*31020*/;
  assign _1533_ = _1532_ & _1531_ /*31019*/;
  assign _1534_ = inv_4[41] & r_3[41] /*31018*/;
  assign _1535_ = _1533_ | _1534_ /*31017*/;
  assign _1536_ = inv_4[42] ^ r_3[42] /*31015*/;
  assign sum_4[42] = _1536_ ^ _1535_ /*31014*/;
  assign _1537_ = _1536_ & _1535_ /*31013*/;
  assign _1538_ = inv_4[42] & r_3[42] /*31012*/;
  assign _1539_ = _1537_ | _1538_ /*31011*/;
  assign _1540_ = inv_4[43] ^ r_3[43] /*31009*/;
  assign sum_4[43] = _1540_ ^ _1539_ /*31008*/;
  assign _1541_ = _1540_ & _1539_ /*31007*/;
  assign _1542_ = inv_4[43] & r_3[43] /*31006*/;
  assign _1543_ = _1541_ | _1542_ /*31005*/;
  assign _1544_ = inv_4[44] ^ r_3[44] /*31003*/;
  assign sum_4[44] = _1544_ ^ _1543_ /*31002*/;
  assign _1545_ = _1544_ & _1543_ /*31001*/;
  assign _1546_ = inv_4[44] & r_3[44] /*31000*/;
  assign _1547_ = _1545_ | _1546_ /*30999*/;
  assign _1548_ = inv_4[45] ^ r_3[45] /*30997*/;
  assign sum_4[45] = _1548_ ^ _1547_ /*30996*/;
  assign _1549_ = _1548_ & _1547_ /*30995*/;
  assign _1550_ = inv_4[45] & r_3[45] /*30994*/;
  assign _1551_ = _1549_ | _1550_ /*30993*/;
  assign _1552_ = inv_4[46] ^ r_3[46] /*30991*/;
  assign sum_4[46] = _1552_ ^ _1551_ /*30990*/;
  assign _1553_ = _1552_ & _1551_ /*30989*/;
  assign _1554_ = inv_4[46] & r_3[46] /*30988*/;
  assign _1555_ = _1553_ | _1554_ /*30987*/;
  assign _1556_ = inv_4[47] ^ r_3[47] /*30985*/;
  assign sum_4[47] = _1556_ ^ _1555_ /*30984*/;
  assign _1557_ = _1556_ & _1555_ /*30983*/;
  assign _1558_ = inv_4[47] & r_3[47] /*30982*/;
  assign _1559_ = _1557_ | _1558_ /*30981*/;
  assign _1560_ = inv_4[48] ^ r_3[48] /*30979*/;
  assign sum_4[48] = _1560_ ^ _1559_ /*30978*/;
  assign _1561_ = _1560_ & _1559_ /*30977*/;
  assign _1562_ = inv_4[48] & r_3[48] /*30976*/;
  assign _1563_ = _1561_ | _1562_ /*30975*/;
  assign _1564_ = inv_4[49] ^ r_3[49] /*30973*/;
  assign sum_4[49] = _1564_ ^ _1563_ /*30972*/;
  assign _1565_ = _1564_ & _1563_ /*30971*/;
  assign _1566_ = inv_4[49] & r_3[49] /*30970*/;
  assign _1567_ = _1565_ | _1566_ /*30969*/;
  assign _1568_ = inv_4[50] ^ r_3[50] /*30967*/;
  assign sum_4[50] = _1568_ ^ _1567_ /*30966*/;
  assign _1569_ = _1568_ & _1567_ /*30965*/;
  assign _1570_ = inv_4[50] & r_3[50] /*30964*/;
  assign _1571_ = _1569_ | _1570_ /*30963*/;
  assign _1572_ = inv_4[51] ^ r_3[51] /*30961*/;
  assign sum_4[51] = _1572_ ^ _1571_ /*30960*/;
  assign _1573_ = _1572_ & _1571_ /*30959*/;
  assign _1574_ = inv_4[51] & r_3[51] /*30958*/;
  assign _1575_ = _1573_ | _1574_ /*30957*/;
  assign _1576_ = inv_4[52] ^ r_3[52] /*30955*/;
  assign sum_4[52] = _1576_ ^ _1575_ /*30954*/;
  assign _1577_ = _1576_ & _1575_ /*30953*/;
  assign _1578_ = inv_4[52] & r_3[52] /*30952*/;
  assign _1579_ = _1577_ | _1578_ /*30951*/;
  assign _1580_ = inv_4[53] ^ r_3[53] /*30949*/;
  assign sum_4[53] = _1580_ ^ _1579_ /*30948*/;
  assign _1581_ = _1580_ & _1579_ /*30947*/;
  assign _1582_ = inv_4[53] & r_3[53] /*30946*/;
  assign _1583_ = _1581_ | _1582_ /*30945*/;
  assign _1584_ = inv_4[54] ^ r_3[54] /*30943*/;
  assign sum_4[54] = _1584_ ^ _1583_ /*30942*/;
  assign _1585_ = _1584_ & _1583_ /*30941*/;
  assign _1586_ = inv_4[54] & r_3[54] /*30940*/;
  assign _1587_ = _1585_ | _1586_ /*30939*/;
  assign _1588_ = inv_4[55] ^ r_3[55] /*30937*/;
  assign sum_4[55] = _1588_ ^ _1587_ /*30936*/;
  assign _1589_ = _1588_ & _1587_ /*30935*/;
  assign _1590_ = inv_4[55] & r_3[55] /*30934*/;
  assign _1591_ = _1589_ | _1590_ /*30933*/;
  assign _1592_ = inv_4[56] ^ r_3[56] /*30931*/;
  assign sum_4[56] = _1592_ ^ _1591_ /*30930*/;
  assign _1593_ = _1592_ & _1591_ /*30929*/;
  assign _1594_ = inv_4[56] & r_3[56] /*30928*/;
  assign _1595_ = _1593_ | _1594_ /*30927*/;
  assign _1596_ = inv_4[57] ^ r_3[57] /*30925*/;
  assign sum_4[57] = _1596_ ^ _1595_ /*30924*/;
  assign _1597_ = _1596_ & _1595_ /*30923*/;
  assign _1598_ = inv_4[57] & r_3[57] /*30922*/;
  assign _1599_ = _1597_ | _1598_ /*30921*/;
  assign _1600_ = inv_4[58] ^ r_3[58] /*30919*/;
  assign sum_4[58] = _1600_ ^ _1599_ /*30918*/;
  assign _1601_ = _1600_ & _1599_ /*30917*/;
  assign _1602_ = inv_4[58] & r_3[58] /*30916*/;
  assign _1603_ = _1601_ | _1602_ /*30915*/;
  assign _1604_ = inv_4[59] ^ r_3[59] /*30913*/;
  assign sum_4[59] = _1604_ ^ _1603_ /*30912*/;
  assign _1605_ = _1604_ & _1603_ /*30911*/;
  assign _1606_ = inv_4[59] & r_3[59] /*30910*/;
  assign _1607_ = _1605_ | _1606_ /*30909*/;
  assign _1608_ = inv_4[60] ^ r_3[60] /*30907*/;
  assign sum_4[60] = _1608_ ^ _1607_ /*30906*/;
  assign _1609_ = _1608_ & _1607_ /*30905*/;
  assign _1610_ = inv_4[60] & r_3[60] /*30904*/;
  assign _1611_ = _1609_ | _1610_ /*30903*/;
  assign _1612_ = inv_4[61] ^ r_3[61] /*30901*/;
  assign sum_4[61] = _1612_ ^ _1611_ /*30900*/;
  assign _1613_ = _1612_ & _1611_ /*30899*/;
  assign _1614_ = inv_4[61] & r_3[61] /*30898*/;
  assign _1615_ = _1613_ | _1614_ /*30897*/;
  assign _1616_ = inv_4[62] ^ r_3[62] /*30895*/;
  assign sum_4[62] = _1616_ ^ _1615_ /*30894*/;
  assign _1617_ = _1616_ & _1615_ /*30893*/;
  assign _1618_ = inv_4[62] & r_3[62] /*30892*/;
  assign _1619_ = _1617_ | _1618_ /*30891*/;
  assign _1620_ = inv_4[63] ^ r_3[63] /*30889*/;
  assign sum_4[63] = _1620_ ^ _1619_ /*30888*/;
  assign _1621_ = _1620_ & _1619_ /*30887*/;
  assign _1622_ = inv_4[63] & r_3[63] /*30886*/;
  assign _1623_ = _1621_ | _1622_ /*30885*/;
  assign _1624_ = inv_4[64] ^ r_3[64] /*30883*/;
  assign sum_4[64] = _1624_ ^ _1623_ /*30882*/;
  assign _1625_ = _1624_ & _1623_ /*30881*/;
  assign _1626_ = inv_4[64] & r_3[64] /*30880*/;
  assign _1627_ = _1625_ | _1626_ /*30879*/;
  assign _1628_ = inv_4[65] ^ r_3[65] /*30877*/;
  assign sum_4[65] = _1628_ ^ _1627_ /*30876*/;
  assign _1629_ = _1628_ & _1627_ /*30875*/;
  assign _1630_ = inv_4[65] & r_3[65] /*30874*/;
  assign _1631_ = _1629_ | _1630_ /*30873*/;
  assign _1632_ = _1631_ ^ _1627_ /*30872*/;
  assign _1633_ = ~_1632_ /*30871*/;
  assign _1634_ = sum_4[65] & _1633_ /*30870*/;
  assign _1635_ = _1632_ & _1631_ /*30869*/;
  assign sum_4[66] = _1635_ | _1634_ /*30868*/;
  assign q[28] = ~sum_4[66] /*30867*/;
  assign m_4[0] = r_3[0] /*30866*/;
  assign m_4[1] = r_3[1] /*30865*/;
  assign m_4[2] = r_3[2] /*30864*/;
  assign m_4[3] = r_3[3] /*30863*/;
  assign m_4[4] = r_3[4] /*30862*/;
  assign m_4[5] = r_3[5] /*30861*/;
  assign m_4[6] = r_3[6] /*30860*/;
  assign m_4[7] = r_3[7] /*30859*/;
  assign m_4[8] = r_3[8] /*30858*/;
  assign m_4[9] = r_3[9] /*30857*/;
  assign m_4[10] = r_3[10] /*30856*/;
  assign m_4[11] = r_3[11] /*30855*/;
  assign m_4[12] = r_3[12] /*30854*/;
  assign m_4[13] = r_3[13] /*30853*/;
  assign m_4[14] = r_3[14] /*30852*/;
  assign m_4[15] = r_3[15] /*30851*/;
  assign m_4[16] = r_3[16] /*30850*/;
  assign m_4[17] = r_3[17] /*30849*/;
  assign m_4[18] = r_3[18] /*30848*/;
  assign m_4[19] = r_3[19] /*30847*/;
  assign m_4[20] = r_3[20] /*30846*/;
  assign m_4[21] = r_3[21] /*30845*/;
  assign m_4[22] = r_3[22] /*30844*/;
  assign m_4[23] = r_3[23] /*30843*/;
  assign m_4[24] = r_3[24] /*30842*/;
  assign m_4[25] = r_3[25] /*30841*/;
  assign m_4[26] = r_3[26] /*30840*/;
  assign m_4[27] = r_3[27] /*30839*/;
  assign m_4[28] = r_3[28] /*30838*/;
  assign m_4[29] = r_3[29] /*30837*/;
  assign m_4[30] = r_3[30] /*30836*/;
  assign m_4[31] = r_3[31] /*30835*/;
  assign m_4[32] = r_3[32] /*30834*/;
  assign m_4[33] = r_3[33] /*30833*/;
  assign m_4[34] = r_3[34] /*30832*/;
  assign m_4[35] = r_3[35] /*30831*/;
  assign m_4[36] = r_3[36] /*30830*/;
  assign m_4[37] = r_3[37] /*30829*/;
  assign m_4[38] = r_3[38] /*30828*/;
  assign m_4[39] = r_3[39] /*30827*/;
  assign m_4[40] = r_3[40] /*30826*/;
  assign m_4[41] = r_3[41] /*30825*/;
  assign m_4[42] = r_3[42] /*30824*/;
  assign m_4[43] = r_3[43] /*30823*/;
  assign m_4[44] = r_3[44] /*30822*/;
  assign m_4[45] = r_3[45] /*30821*/;
  assign m_4[46] = r_3[46] /*30820*/;
  assign m_4[47] = r_3[47] /*30819*/;
  assign m_4[48] = r_3[48] /*30818*/;
  assign m_4[49] = r_3[49] /*30817*/;
  assign m_4[50] = r_3[50] /*30816*/;
  assign m_4[51] = r_3[51] /*30815*/;
  assign m_4[52] = r_3[52] /*30814*/;
  assign m_4[53] = r_3[53] /*30813*/;
  assign m_4[54] = r_3[54] /*30812*/;
  assign m_4[55] = r_3[55] /*30811*/;
  assign m_4[56] = r_3[56] /*30810*/;
  assign m_4[57] = r_3[57] /*30809*/;
  assign m_4[58] = r_3[58] /*30808*/;
  assign m_4[59] = r_3[59] /*30807*/;
  assign m_4[60] = r_3[60] /*30806*/;
  assign m_4[61] = r_3[61] /*30805*/;
  assign m_4[62] = r_3[62] /*30804*/;
  assign m_4[63] = r_3[63] /*30803*/;
  assign m_4[64] = r_3[64] /*30802*/;
  assign m_4[65] = r_3[65] /*30801*/;
  assign m_4[66] = r_3[65] /*30800*/;
  assign _1637_ = ~q[28] /*30799*/;
  assign _1638_ = sum_4[0] & q[28] /*30798*/;
  assign _1639_ = m_4[0] & _1637_ /*30797*/;
  assign r_4[0] = _1639_ | _1638_ /*30796*/;
  assign _1640_ = ~q[28] /*30795*/;
  assign _1641_ = sum_4[1] & q[28] /*30794*/;
  assign _1642_ = m_4[1] & _1640_ /*30793*/;
  assign r_4[1] = _1642_ | _1641_ /*30792*/;
  assign _1643_ = ~q[28] /*30791*/;
  assign _1644_ = sum_4[2] & q[28] /*30790*/;
  assign _1645_ = m_4[2] & _1643_ /*30789*/;
  assign r_4[2] = _1645_ | _1644_ /*30788*/;
  assign _1646_ = ~q[28] /*30787*/;
  assign _1647_ = sum_4[3] & q[28] /*30786*/;
  assign _1648_ = m_4[3] & _1646_ /*30785*/;
  assign r_4[3] = _1648_ | _1647_ /*30784*/;
  assign _1649_ = ~q[28] /*30783*/;
  assign _1650_ = sum_4[4] & q[28] /*30782*/;
  assign _1651_ = m_4[4] & _1649_ /*30781*/;
  assign r_4[4] = _1651_ | _1650_ /*30780*/;
  assign _1652_ = ~q[28] /*30779*/;
  assign _1653_ = sum_4[5] & q[28] /*30778*/;
  assign _1654_ = m_4[5] & _1652_ /*30777*/;
  assign r_4[5] = _1654_ | _1653_ /*30776*/;
  assign _1655_ = ~q[28] /*30775*/;
  assign _1656_ = sum_4[6] & q[28] /*30774*/;
  assign _1657_ = m_4[6] & _1655_ /*30773*/;
  assign r_4[6] = _1657_ | _1656_ /*30772*/;
  assign _1658_ = ~q[28] /*30771*/;
  assign _1659_ = sum_4[7] & q[28] /*30770*/;
  assign _1660_ = m_4[7] & _1658_ /*30769*/;
  assign r_4[7] = _1660_ | _1659_ /*30768*/;
  assign _1661_ = ~q[28] /*30767*/;
  assign _1662_ = sum_4[8] & q[28] /*30766*/;
  assign _1663_ = m_4[8] & _1661_ /*30765*/;
  assign r_4[8] = _1663_ | _1662_ /*30764*/;
  assign _1664_ = ~q[28] /*30763*/;
  assign _1665_ = sum_4[9] & q[28] /*30762*/;
  assign _1666_ = m_4[9] & _1664_ /*30761*/;
  assign r_4[9] = _1666_ | _1665_ /*30760*/;
  assign _1667_ = ~q[28] /*30759*/;
  assign _1668_ = sum_4[10] & q[28] /*30758*/;
  assign _1669_ = m_4[10] & _1667_ /*30757*/;
  assign r_4[10] = _1669_ | _1668_ /*30756*/;
  assign _1670_ = ~q[28] /*30755*/;
  assign _1671_ = sum_4[11] & q[28] /*30754*/;
  assign _1672_ = m_4[11] & _1670_ /*30753*/;
  assign r_4[11] = _1672_ | _1671_ /*30752*/;
  assign _1673_ = ~q[28] /*30751*/;
  assign _1674_ = sum_4[12] & q[28] /*30750*/;
  assign _1675_ = m_4[12] & _1673_ /*30749*/;
  assign r_4[12] = _1675_ | _1674_ /*30748*/;
  assign _1676_ = ~q[28] /*30747*/;
  assign _1677_ = sum_4[13] & q[28] /*30746*/;
  assign _1678_ = m_4[13] & _1676_ /*30745*/;
  assign r_4[13] = _1678_ | _1677_ /*30744*/;
  assign _1679_ = ~q[28] /*30743*/;
  assign _1680_ = sum_4[14] & q[28] /*30742*/;
  assign _1681_ = m_4[14] & _1679_ /*30741*/;
  assign r_4[14] = _1681_ | _1680_ /*30740*/;
  assign _1682_ = ~q[28] /*30739*/;
  assign _1683_ = sum_4[15] & q[28] /*30738*/;
  assign _1684_ = m_4[15] & _1682_ /*30737*/;
  assign r_4[15] = _1684_ | _1683_ /*30736*/;
  assign _1685_ = ~q[28] /*30735*/;
  assign _1686_ = sum_4[16] & q[28] /*30734*/;
  assign _1687_ = m_4[16] & _1685_ /*30733*/;
  assign r_4[16] = _1687_ | _1686_ /*30732*/;
  assign _1688_ = ~q[28] /*30731*/;
  assign _1689_ = sum_4[17] & q[28] /*30730*/;
  assign _1690_ = m_4[17] & _1688_ /*30729*/;
  assign r_4[17] = _1690_ | _1689_ /*30728*/;
  assign _1691_ = ~q[28] /*30727*/;
  assign _1692_ = sum_4[18] & q[28] /*30726*/;
  assign _1693_ = m_4[18] & _1691_ /*30725*/;
  assign r_4[18] = _1693_ | _1692_ /*30724*/;
  assign _1694_ = ~q[28] /*30723*/;
  assign _1695_ = sum_4[19] & q[28] /*30722*/;
  assign _1696_ = m_4[19] & _1694_ /*30721*/;
  assign r_4[19] = _1696_ | _1695_ /*30720*/;
  assign _1697_ = ~q[28] /*30719*/;
  assign _1698_ = sum_4[20] & q[28] /*30718*/;
  assign _1699_ = m_4[20] & _1697_ /*30717*/;
  assign r_4[20] = _1699_ | _1698_ /*30716*/;
  assign _1700_ = ~q[28] /*30715*/;
  assign _1701_ = sum_4[21] & q[28] /*30714*/;
  assign _1702_ = m_4[21] & _1700_ /*30713*/;
  assign r_4[21] = _1702_ | _1701_ /*30712*/;
  assign _1703_ = ~q[28] /*30711*/;
  assign _1704_ = sum_4[22] & q[28] /*30710*/;
  assign _1705_ = m_4[22] & _1703_ /*30709*/;
  assign r_4[22] = _1705_ | _1704_ /*30708*/;
  assign _1706_ = ~q[28] /*30707*/;
  assign _1707_ = sum_4[23] & q[28] /*30706*/;
  assign _1708_ = m_4[23] & _1706_ /*30705*/;
  assign r_4[23] = _1708_ | _1707_ /*30704*/;
  assign _1709_ = ~q[28] /*30703*/;
  assign _1710_ = sum_4[24] & q[28] /*30702*/;
  assign _1711_ = m_4[24] & _1709_ /*30701*/;
  assign r_4[24] = _1711_ | _1710_ /*30700*/;
  assign _1712_ = ~q[28] /*30699*/;
  assign _1713_ = sum_4[25] & q[28] /*30698*/;
  assign _1714_ = m_4[25] & _1712_ /*30697*/;
  assign r_4[25] = _1714_ | _1713_ /*30696*/;
  assign _1715_ = ~q[28] /*30695*/;
  assign _1716_ = sum_4[26] & q[28] /*30694*/;
  assign _1717_ = m_4[26] & _1715_ /*30693*/;
  assign r_4[26] = _1717_ | _1716_ /*30692*/;
  assign _1718_ = ~q[28] /*30691*/;
  assign _1719_ = sum_4[27] & q[28] /*30690*/;
  assign _1720_ = m_4[27] & _1718_ /*30689*/;
  assign r_4[27] = _1720_ | _1719_ /*30688*/;
  assign _1721_ = ~q[28] /*30687*/;
  assign _1722_ = sum_4[28] & q[28] /*30686*/;
  assign _1723_ = m_4[28] & _1721_ /*30685*/;
  assign r_4[28] = _1723_ | _1722_ /*30684*/;
  assign _1724_ = ~q[28] /*30683*/;
  assign _1725_ = sum_4[29] & q[28] /*30682*/;
  assign _1726_ = m_4[29] & _1724_ /*30681*/;
  assign r_4[29] = _1726_ | _1725_ /*30680*/;
  assign _1727_ = ~q[28] /*30679*/;
  assign _1728_ = sum_4[30] & q[28] /*30678*/;
  assign _1729_ = m_4[30] & _1727_ /*30677*/;
  assign r_4[30] = _1729_ | _1728_ /*30676*/;
  assign _1730_ = ~q[28] /*30675*/;
  assign _1731_ = sum_4[31] & q[28] /*30674*/;
  assign _1732_ = m_4[31] & _1730_ /*30673*/;
  assign r_4[31] = _1732_ | _1731_ /*30672*/;
  assign _1733_ = ~q[28] /*30671*/;
  assign _1734_ = sum_4[32] & q[28] /*30670*/;
  assign _1735_ = m_4[32] & _1733_ /*30669*/;
  assign r_4[32] = _1735_ | _1734_ /*30668*/;
  assign _1736_ = ~q[28] /*30667*/;
  assign _1737_ = sum_4[33] & q[28] /*30666*/;
  assign _1738_ = m_4[33] & _1736_ /*30665*/;
  assign r_4[33] = _1738_ | _1737_ /*30664*/;
  assign _1739_ = ~q[28] /*30663*/;
  assign _1740_ = sum_4[34] & q[28] /*30662*/;
  assign _1741_ = m_4[34] & _1739_ /*30661*/;
  assign r_4[34] = _1741_ | _1740_ /*30660*/;
  assign _1742_ = ~q[28] /*30659*/;
  assign _1743_ = sum_4[35] & q[28] /*30658*/;
  assign _1744_ = m_4[35] & _1742_ /*30657*/;
  assign r_4[35] = _1744_ | _1743_ /*30656*/;
  assign _1745_ = ~q[28] /*30655*/;
  assign _1746_ = sum_4[36] & q[28] /*30654*/;
  assign _1747_ = m_4[36] & _1745_ /*30653*/;
  assign r_4[36] = _1747_ | _1746_ /*30652*/;
  assign _1748_ = ~q[28] /*30651*/;
  assign _1749_ = sum_4[37] & q[28] /*30650*/;
  assign _1750_ = m_4[37] & _1748_ /*30649*/;
  assign r_4[37] = _1750_ | _1749_ /*30648*/;
  assign _1751_ = ~q[28] /*30647*/;
  assign _1752_ = sum_4[38] & q[28] /*30646*/;
  assign _1753_ = m_4[38] & _1751_ /*30645*/;
  assign r_4[38] = _1753_ | _1752_ /*30644*/;
  assign _1754_ = ~q[28] /*30643*/;
  assign _1755_ = sum_4[39] & q[28] /*30642*/;
  assign _1756_ = m_4[39] & _1754_ /*30641*/;
  assign r_4[39] = _1756_ | _1755_ /*30640*/;
  assign _1757_ = ~q[28] /*30639*/;
  assign _1758_ = sum_4[40] & q[28] /*30638*/;
  assign _1759_ = m_4[40] & _1757_ /*30637*/;
  assign r_4[40] = _1759_ | _1758_ /*30636*/;
  assign _1760_ = ~q[28] /*30635*/;
  assign _1761_ = sum_4[41] & q[28] /*30634*/;
  assign _1762_ = m_4[41] & _1760_ /*30633*/;
  assign r_4[41] = _1762_ | _1761_ /*30632*/;
  assign _1763_ = ~q[28] /*30631*/;
  assign _1764_ = sum_4[42] & q[28] /*30630*/;
  assign _1765_ = m_4[42] & _1763_ /*30629*/;
  assign r_4[42] = _1765_ | _1764_ /*30628*/;
  assign _1766_ = ~q[28] /*30627*/;
  assign _1767_ = sum_4[43] & q[28] /*30626*/;
  assign _1768_ = m_4[43] & _1766_ /*30625*/;
  assign r_4[43] = _1768_ | _1767_ /*30624*/;
  assign _1769_ = ~q[28] /*30623*/;
  assign _1770_ = sum_4[44] & q[28] /*30622*/;
  assign _1771_ = m_4[44] & _1769_ /*30621*/;
  assign r_4[44] = _1771_ | _1770_ /*30620*/;
  assign _1772_ = ~q[28] /*30619*/;
  assign _1773_ = sum_4[45] & q[28] /*30618*/;
  assign _1774_ = m_4[45] & _1772_ /*30617*/;
  assign r_4[45] = _1774_ | _1773_ /*30616*/;
  assign _1775_ = ~q[28] /*30615*/;
  assign _1776_ = sum_4[46] & q[28] /*30614*/;
  assign _1777_ = m_4[46] & _1775_ /*30613*/;
  assign r_4[46] = _1777_ | _1776_ /*30612*/;
  assign _1778_ = ~q[28] /*30611*/;
  assign _1779_ = sum_4[47] & q[28] /*30610*/;
  assign _1780_ = m_4[47] & _1778_ /*30609*/;
  assign r_4[47] = _1780_ | _1779_ /*30608*/;
  assign _1781_ = ~q[28] /*30607*/;
  assign _1782_ = sum_4[48] & q[28] /*30606*/;
  assign _1783_ = m_4[48] & _1781_ /*30605*/;
  assign r_4[48] = _1783_ | _1782_ /*30604*/;
  assign _1784_ = ~q[28] /*30603*/;
  assign _1785_ = sum_4[49] & q[28] /*30602*/;
  assign _1786_ = m_4[49] & _1784_ /*30601*/;
  assign r_4[49] = _1786_ | _1785_ /*30600*/;
  assign _1787_ = ~q[28] /*30599*/;
  assign _1788_ = sum_4[50] & q[28] /*30598*/;
  assign _1789_ = m_4[50] & _1787_ /*30597*/;
  assign r_4[50] = _1789_ | _1788_ /*30596*/;
  assign _1790_ = ~q[28] /*30595*/;
  assign _1791_ = sum_4[51] & q[28] /*30594*/;
  assign _1792_ = m_4[51] & _1790_ /*30593*/;
  assign r_4[51] = _1792_ | _1791_ /*30592*/;
  assign _1793_ = ~q[28] /*30591*/;
  assign _1794_ = sum_4[52] & q[28] /*30590*/;
  assign _1795_ = m_4[52] & _1793_ /*30589*/;
  assign r_4[52] = _1795_ | _1794_ /*30588*/;
  assign _1796_ = ~q[28] /*30587*/;
  assign _1797_ = sum_4[53] & q[28] /*30586*/;
  assign _1798_ = m_4[53] & _1796_ /*30585*/;
  assign r_4[53] = _1798_ | _1797_ /*30584*/;
  assign _1799_ = ~q[28] /*30583*/;
  assign _1800_ = sum_4[54] & q[28] /*30582*/;
  assign _1801_ = m_4[54] & _1799_ /*30581*/;
  assign r_4[54] = _1801_ | _1800_ /*30580*/;
  assign _1802_ = ~q[28] /*30579*/;
  assign _1803_ = sum_4[55] & q[28] /*30578*/;
  assign _1804_ = m_4[55] & _1802_ /*30577*/;
  assign r_4[55] = _1804_ | _1803_ /*30576*/;
  assign _1805_ = ~q[28] /*30575*/;
  assign _1806_ = sum_4[56] & q[28] /*30574*/;
  assign _1807_ = m_4[56] & _1805_ /*30573*/;
  assign r_4[56] = _1807_ | _1806_ /*30572*/;
  assign _1808_ = ~q[28] /*30571*/;
  assign _1809_ = sum_4[57] & q[28] /*30570*/;
  assign _1810_ = m_4[57] & _1808_ /*30569*/;
  assign r_4[57] = _1810_ | _1809_ /*30568*/;
  assign _1811_ = ~q[28] /*30567*/;
  assign _1812_ = sum_4[58] & q[28] /*30566*/;
  assign _1813_ = m_4[58] & _1811_ /*30565*/;
  assign r_4[58] = _1813_ | _1812_ /*30564*/;
  assign _1814_ = ~q[28] /*30563*/;
  assign _1815_ = sum_4[59] & q[28] /*30562*/;
  assign _1816_ = m_4[59] & _1814_ /*30561*/;
  assign r_4[59] = _1816_ | _1815_ /*30560*/;
  assign _1817_ = ~q[28] /*30559*/;
  assign _1818_ = sum_4[60] & q[28] /*30558*/;
  assign _1819_ = m_4[60] & _1817_ /*30557*/;
  assign r_4[60] = _1819_ | _1818_ /*30556*/;
  assign _1820_ = ~q[28] /*30555*/;
  assign _1821_ = sum_4[61] & q[28] /*30554*/;
  assign _1822_ = m_4[61] & _1820_ /*30553*/;
  assign r_4[61] = _1822_ | _1821_ /*30552*/;
  assign _1823_ = ~q[28] /*30551*/;
  assign _1824_ = sum_4[62] & q[28] /*30550*/;
  assign _1825_ = m_4[62] & _1823_ /*30549*/;
  assign r_4[62] = _1825_ | _1824_ /*30548*/;
  assign _1826_ = ~q[28] /*30547*/;
  assign _1827_ = sum_4[63] & q[28] /*30546*/;
  assign _1828_ = m_4[63] & _1826_ /*30545*/;
  assign r_4[63] = _1828_ | _1827_ /*30544*/;
  assign _1829_ = ~q[28] /*30543*/;
  assign _1830_ = sum_4[64] & q[28] /*30542*/;
  assign _1831_ = m_4[64] & _1829_ /*30541*/;
  assign r_4[64] = _1831_ | _1830_ /*30540*/;
  assign _1832_ = ~q[28] /*30539*/;
  assign _1833_ = sum_4[65] & q[28] /*30538*/;
  assign _1834_ = m_4[65] & _1832_ /*30537*/;
  assign r_4[65] = _1834_ | _1833_ /*30536*/;
  assign _1835_ = ~q[28] /*30535*/;
  assign _1836_ = sum_4[66] & q[28] /*30534*/;
  assign _1837_ = m_4[66] & _1835_ /*30533*/;
  assign r_4[66] = _1837_ | _1836_ /*30532*/;
  assign inv_5[0] = oneWire /*30192*/;
  assign inv_5[1] = oneWire /*30186*/;
  assign inv_5[2] = oneWire /*30180*/;
  assign inv_5[3] = oneWire /*30174*/;
  assign inv_5[4] = oneWire /*30168*/;
  assign inv_5[5] = oneWire /*30162*/;
  assign inv_5[6] = oneWire /*30156*/;
  assign inv_5[7] = oneWire /*30150*/;
  assign inv_5[8] = oneWire /*30144*/;
  assign inv_5[9] = oneWire /*30138*/;
  assign inv_5[10] = oneWire /*30132*/;
  assign inv_5[11] = oneWire /*30126*/;
  assign inv_5[12] = oneWire /*30120*/;
  assign inv_5[13] = oneWire /*30114*/;
  assign inv_5[14] = oneWire /*30108*/;
  assign inv_5[15] = oneWire /*30102*/;
  assign inv_5[16] = oneWire /*30096*/;
  assign inv_5[17] = oneWire /*30090*/;
  assign inv_5[18] = oneWire /*30084*/;
  assign inv_5[19] = oneWire /*30078*/;
  assign inv_5[20] = oneWire /*30072*/;
  assign inv_5[21] = oneWire /*30066*/;
  assign inv_5[22] = oneWire /*30060*/;
  assign inv_5[23] = oneWire /*30054*/;
  assign inv_5[24] = oneWire /*30048*/;
  assign inv_5[25] = oneWire /*30042*/;
  assign inv_5[26] = oneWire /*30036*/;
  assign inv_5[27] = ~div[0] /*30030*/;
  assign inv_5[28] = ~div[1] /*30024*/;
  assign inv_5[29] = ~div[2] /*30018*/;
  assign inv_5[30] = ~div[3] /*30012*/;
  assign inv_5[31] = ~div[4] /*30006*/;
  assign inv_5[32] = ~div[5] /*30000*/;
  assign inv_5[33] = ~div[6] /*29994*/;
  assign inv_5[34] = ~div[7] /*29988*/;
  assign inv_5[35] = ~div[8] /*29982*/;
  assign inv_5[36] = ~div[9] /*29976*/;
  assign inv_5[37] = ~div[10] /*29970*/;
  assign inv_5[38] = ~div[11] /*29964*/;
  assign inv_5[39] = ~div[12] /*29958*/;
  assign inv_5[40] = ~div[13] /*29952*/;
  assign inv_5[41] = ~div[14] /*29946*/;
  assign inv_5[42] = ~div[15] /*29940*/;
  assign inv_5[43] = ~div[16] /*29934*/;
  assign inv_5[44] = ~div[17] /*29928*/;
  assign inv_5[45] = ~div[18] /*29922*/;
  assign inv_5[46] = ~div[19] /*29916*/;
  assign inv_5[47] = ~div[20] /*29910*/;
  assign inv_5[48] = ~div[21] /*29904*/;
  assign inv_5[49] = ~div[22] /*29898*/;
  assign inv_5[50] = ~div[23] /*29892*/;
  assign inv_5[51] = ~div[24] /*29886*/;
  assign inv_5[52] = ~div[25] /*29880*/;
  assign inv_5[53] = ~div[26] /*29874*/;
  assign inv_5[54] = ~div[27] /*29868*/;
  assign inv_5[55] = ~div[28] /*29862*/;
  assign inv_5[56] = ~div[29] /*29856*/;
  assign inv_5[57] = ~div[30] /*29850*/;
  assign inv_5[58] = oneWire /*29844*/;
  assign inv_5[59] = oneWire /*29838*/;
  assign inv_5[60] = oneWire /*29832*/;
  assign inv_5[61] = oneWire /*29826*/;
  assign inv_5[62] = oneWire /*29820*/;
  assign inv_5[63] = oneWire /*29814*/;
  assign inv_5[64] = oneWire /*29808*/;
  assign inv_5[65] = oneWire /*29802*/;
  assign inv_5[66] = oneWire /*29796*/;
  assign _1838_ = inv_5[0] ^ r_4[0] /*30191*/;
  assign sum_5[0] = _1838_ ^ oneWire /*30190*/;
  assign _1839_ = _1838_ & oneWire /*30189*/;
  assign _1840_ = inv_5[0] & r_4[0] /*30188*/;
  assign _1841_ = _1839_ | _1840_ /*30187*/;
  assign _1842_ = inv_5[1] ^ r_4[1] /*30185*/;
  assign sum_5[1] = _1842_ ^ _1841_ /*30184*/;
  assign _1843_ = _1842_ & _1841_ /*30183*/;
  assign _1844_ = inv_5[1] & r_4[1] /*30182*/;
  assign _1845_ = _1843_ | _1844_ /*30181*/;
  assign _1846_ = inv_5[2] ^ r_4[2] /*30179*/;
  assign sum_5[2] = _1846_ ^ _1845_ /*30178*/;
  assign _1847_ = _1846_ & _1845_ /*30177*/;
  assign _1848_ = inv_5[2] & r_4[2] /*30176*/;
  assign _1849_ = _1847_ | _1848_ /*30175*/;
  assign _1850_ = inv_5[3] ^ r_4[3] /*30173*/;
  assign sum_5[3] = _1850_ ^ _1849_ /*30172*/;
  assign _1851_ = _1850_ & _1849_ /*30171*/;
  assign _1852_ = inv_5[3] & r_4[3] /*30170*/;
  assign _1853_ = _1851_ | _1852_ /*30169*/;
  assign _1854_ = inv_5[4] ^ r_4[4] /*30167*/;
  assign sum_5[4] = _1854_ ^ _1853_ /*30166*/;
  assign _1855_ = _1854_ & _1853_ /*30165*/;
  assign _1856_ = inv_5[4] & r_4[4] /*30164*/;
  assign _1857_ = _1855_ | _1856_ /*30163*/;
  assign _1858_ = inv_5[5] ^ r_4[5] /*30161*/;
  assign sum_5[5] = _1858_ ^ _1857_ /*30160*/;
  assign _1859_ = _1858_ & _1857_ /*30159*/;
  assign _1860_ = inv_5[5] & r_4[5] /*30158*/;
  assign _1861_ = _1859_ | _1860_ /*30157*/;
  assign _1862_ = inv_5[6] ^ r_4[6] /*30155*/;
  assign sum_5[6] = _1862_ ^ _1861_ /*30154*/;
  assign _1863_ = _1862_ & _1861_ /*30153*/;
  assign _1864_ = inv_5[6] & r_4[6] /*30152*/;
  assign _1865_ = _1863_ | _1864_ /*30151*/;
  assign _1866_ = inv_5[7] ^ r_4[7] /*30149*/;
  assign sum_5[7] = _1866_ ^ _1865_ /*30148*/;
  assign _1867_ = _1866_ & _1865_ /*30147*/;
  assign _1868_ = inv_5[7] & r_4[7] /*30146*/;
  assign _1869_ = _1867_ | _1868_ /*30145*/;
  assign _1870_ = inv_5[8] ^ r_4[8] /*30143*/;
  assign sum_5[8] = _1870_ ^ _1869_ /*30142*/;
  assign _1871_ = _1870_ & _1869_ /*30141*/;
  assign _1872_ = inv_5[8] & r_4[8] /*30140*/;
  assign _1873_ = _1871_ | _1872_ /*30139*/;
  assign _1874_ = inv_5[9] ^ r_4[9] /*30137*/;
  assign sum_5[9] = _1874_ ^ _1873_ /*30136*/;
  assign _1875_ = _1874_ & _1873_ /*30135*/;
  assign _1876_ = inv_5[9] & r_4[9] /*30134*/;
  assign _1877_ = _1875_ | _1876_ /*30133*/;
  assign _1878_ = inv_5[10] ^ r_4[10] /*30131*/;
  assign sum_5[10] = _1878_ ^ _1877_ /*30130*/;
  assign _1879_ = _1878_ & _1877_ /*30129*/;
  assign _1880_ = inv_5[10] & r_4[10] /*30128*/;
  assign _1881_ = _1879_ | _1880_ /*30127*/;
  assign _1882_ = inv_5[11] ^ r_4[11] /*30125*/;
  assign sum_5[11] = _1882_ ^ _1881_ /*30124*/;
  assign _1883_ = _1882_ & _1881_ /*30123*/;
  assign _1884_ = inv_5[11] & r_4[11] /*30122*/;
  assign _1885_ = _1883_ | _1884_ /*30121*/;
  assign _1886_ = inv_5[12] ^ r_4[12] /*30119*/;
  assign sum_5[12] = _1886_ ^ _1885_ /*30118*/;
  assign _1887_ = _1886_ & _1885_ /*30117*/;
  assign _1888_ = inv_5[12] & r_4[12] /*30116*/;
  assign _1889_ = _1887_ | _1888_ /*30115*/;
  assign _1890_ = inv_5[13] ^ r_4[13] /*30113*/;
  assign sum_5[13] = _1890_ ^ _1889_ /*30112*/;
  assign _1891_ = _1890_ & _1889_ /*30111*/;
  assign _1892_ = inv_5[13] & r_4[13] /*30110*/;
  assign _1893_ = _1891_ | _1892_ /*30109*/;
  assign _1894_ = inv_5[14] ^ r_4[14] /*30107*/;
  assign sum_5[14] = _1894_ ^ _1893_ /*30106*/;
  assign _1895_ = _1894_ & _1893_ /*30105*/;
  assign _1896_ = inv_5[14] & r_4[14] /*30104*/;
  assign _1897_ = _1895_ | _1896_ /*30103*/;
  assign _1898_ = inv_5[15] ^ r_4[15] /*30101*/;
  assign sum_5[15] = _1898_ ^ _1897_ /*30100*/;
  assign _1899_ = _1898_ & _1897_ /*30099*/;
  assign _1900_ = inv_5[15] & r_4[15] /*30098*/;
  assign _1901_ = _1899_ | _1900_ /*30097*/;
  assign _1902_ = inv_5[16] ^ r_4[16] /*30095*/;
  assign sum_5[16] = _1902_ ^ _1901_ /*30094*/;
  assign _1903_ = _1902_ & _1901_ /*30093*/;
  assign _1904_ = inv_5[16] & r_4[16] /*30092*/;
  assign _1905_ = _1903_ | _1904_ /*30091*/;
  assign _1906_ = inv_5[17] ^ r_4[17] /*30089*/;
  assign sum_5[17] = _1906_ ^ _1905_ /*30088*/;
  assign _1907_ = _1906_ & _1905_ /*30087*/;
  assign _1908_ = inv_5[17] & r_4[17] /*30086*/;
  assign _1909_ = _1907_ | _1908_ /*30085*/;
  assign _1910_ = inv_5[18] ^ r_4[18] /*30083*/;
  assign sum_5[18] = _1910_ ^ _1909_ /*30082*/;
  assign _1911_ = _1910_ & _1909_ /*30081*/;
  assign _1912_ = inv_5[18] & r_4[18] /*30080*/;
  assign _1913_ = _1911_ | _1912_ /*30079*/;
  assign _1914_ = inv_5[19] ^ r_4[19] /*30077*/;
  assign sum_5[19] = _1914_ ^ _1913_ /*30076*/;
  assign _1915_ = _1914_ & _1913_ /*30075*/;
  assign _1916_ = inv_5[19] & r_4[19] /*30074*/;
  assign _1917_ = _1915_ | _1916_ /*30073*/;
  assign _1918_ = inv_5[20] ^ r_4[20] /*30071*/;
  assign sum_5[20] = _1918_ ^ _1917_ /*30070*/;
  assign _1919_ = _1918_ & _1917_ /*30069*/;
  assign _1920_ = inv_5[20] & r_4[20] /*30068*/;
  assign _1921_ = _1919_ | _1920_ /*30067*/;
  assign _1922_ = inv_5[21] ^ r_4[21] /*30065*/;
  assign sum_5[21] = _1922_ ^ _1921_ /*30064*/;
  assign _1923_ = _1922_ & _1921_ /*30063*/;
  assign _1924_ = inv_5[21] & r_4[21] /*30062*/;
  assign _1925_ = _1923_ | _1924_ /*30061*/;
  assign _1926_ = inv_5[22] ^ r_4[22] /*30059*/;
  assign sum_5[22] = _1926_ ^ _1925_ /*30058*/;
  assign _1927_ = _1926_ & _1925_ /*30057*/;
  assign _1928_ = inv_5[22] & r_4[22] /*30056*/;
  assign _1929_ = _1927_ | _1928_ /*30055*/;
  assign _1930_ = inv_5[23] ^ r_4[23] /*30053*/;
  assign sum_5[23] = _1930_ ^ _1929_ /*30052*/;
  assign _1931_ = _1930_ & _1929_ /*30051*/;
  assign _1932_ = inv_5[23] & r_4[23] /*30050*/;
  assign _1933_ = _1931_ | _1932_ /*30049*/;
  assign _1934_ = inv_5[24] ^ r_4[24] /*30047*/;
  assign sum_5[24] = _1934_ ^ _1933_ /*30046*/;
  assign _1935_ = _1934_ & _1933_ /*30045*/;
  assign _1936_ = inv_5[24] & r_4[24] /*30044*/;
  assign _1937_ = _1935_ | _1936_ /*30043*/;
  assign _1938_ = inv_5[25] ^ r_4[25] /*30041*/;
  assign sum_5[25] = _1938_ ^ _1937_ /*30040*/;
  assign _1939_ = _1938_ & _1937_ /*30039*/;
  assign _1940_ = inv_5[25] & r_4[25] /*30038*/;
  assign _1941_ = _1939_ | _1940_ /*30037*/;
  assign _1942_ = inv_5[26] ^ r_4[26] /*30035*/;
  assign sum_5[26] = _1942_ ^ _1941_ /*30034*/;
  assign _1943_ = _1942_ & _1941_ /*30033*/;
  assign _1944_ = inv_5[26] & r_4[26] /*30032*/;
  assign _1945_ = _1943_ | _1944_ /*30031*/;
  assign _1946_ = inv_5[27] ^ r_4[27] /*30029*/;
  assign sum_5[27] = _1946_ ^ _1945_ /*30028*/;
  assign _1947_ = _1946_ & _1945_ /*30027*/;
  assign _1948_ = inv_5[27] & r_4[27] /*30026*/;
  assign _1949_ = _1947_ | _1948_ /*30025*/;
  assign _1950_ = inv_5[28] ^ r_4[28] /*30023*/;
  assign sum_5[28] = _1950_ ^ _1949_ /*30022*/;
  assign _1951_ = _1950_ & _1949_ /*30021*/;
  assign _1952_ = inv_5[28] & r_4[28] /*30020*/;
  assign _1953_ = _1951_ | _1952_ /*30019*/;
  assign _1954_ = inv_5[29] ^ r_4[29] /*30017*/;
  assign sum_5[29] = _1954_ ^ _1953_ /*30016*/;
  assign _1955_ = _1954_ & _1953_ /*30015*/;
  assign _1956_ = inv_5[29] & r_4[29] /*30014*/;
  assign _1957_ = _1955_ | _1956_ /*30013*/;
  assign _1958_ = inv_5[30] ^ r_4[30] /*30011*/;
  assign sum_5[30] = _1958_ ^ _1957_ /*30010*/;
  assign _1959_ = _1958_ & _1957_ /*30009*/;
  assign _1960_ = inv_5[30] & r_4[30] /*30008*/;
  assign _1961_ = _1959_ | _1960_ /*30007*/;
  assign _1962_ = inv_5[31] ^ r_4[31] /*30005*/;
  assign sum_5[31] = _1962_ ^ _1961_ /*30004*/;
  assign _1963_ = _1962_ & _1961_ /*30003*/;
  assign _1964_ = inv_5[31] & r_4[31] /*30002*/;
  assign _1965_ = _1963_ | _1964_ /*30001*/;
  assign _1966_ = inv_5[32] ^ r_4[32] /*29999*/;
  assign sum_5[32] = _1966_ ^ _1965_ /*29998*/;
  assign _1967_ = _1966_ & _1965_ /*29997*/;
  assign _1968_ = inv_5[32] & r_4[32] /*29996*/;
  assign _1969_ = _1967_ | _1968_ /*29995*/;
  assign _1970_ = inv_5[33] ^ r_4[33] /*29993*/;
  assign sum_5[33] = _1970_ ^ _1969_ /*29992*/;
  assign _1971_ = _1970_ & _1969_ /*29991*/;
  assign _1972_ = inv_5[33] & r_4[33] /*29990*/;
  assign _1973_ = _1971_ | _1972_ /*29989*/;
  assign _1974_ = inv_5[34] ^ r_4[34] /*29987*/;
  assign sum_5[34] = _1974_ ^ _1973_ /*29986*/;
  assign _1975_ = _1974_ & _1973_ /*29985*/;
  assign _1976_ = inv_5[34] & r_4[34] /*29984*/;
  assign _1977_ = _1975_ | _1976_ /*29983*/;
  assign _1978_ = inv_5[35] ^ r_4[35] /*29981*/;
  assign sum_5[35] = _1978_ ^ _1977_ /*29980*/;
  assign _1979_ = _1978_ & _1977_ /*29979*/;
  assign _1980_ = inv_5[35] & r_4[35] /*29978*/;
  assign _1981_ = _1979_ | _1980_ /*29977*/;
  assign _1982_ = inv_5[36] ^ r_4[36] /*29975*/;
  assign sum_5[36] = _1982_ ^ _1981_ /*29974*/;
  assign _1983_ = _1982_ & _1981_ /*29973*/;
  assign _1984_ = inv_5[36] & r_4[36] /*29972*/;
  assign _1985_ = _1983_ | _1984_ /*29971*/;
  assign _1986_ = inv_5[37] ^ r_4[37] /*29969*/;
  assign sum_5[37] = _1986_ ^ _1985_ /*29968*/;
  assign _1987_ = _1986_ & _1985_ /*29967*/;
  assign _1988_ = inv_5[37] & r_4[37] /*29966*/;
  assign _1989_ = _1987_ | _1988_ /*29965*/;
  assign _1990_ = inv_5[38] ^ r_4[38] /*29963*/;
  assign sum_5[38] = _1990_ ^ _1989_ /*29962*/;
  assign _1991_ = _1990_ & _1989_ /*29961*/;
  assign _1992_ = inv_5[38] & r_4[38] /*29960*/;
  assign _1993_ = _1991_ | _1992_ /*29959*/;
  assign _1994_ = inv_5[39] ^ r_4[39] /*29957*/;
  assign sum_5[39] = _1994_ ^ _1993_ /*29956*/;
  assign _1995_ = _1994_ & _1993_ /*29955*/;
  assign _1996_ = inv_5[39] & r_4[39] /*29954*/;
  assign _1997_ = _1995_ | _1996_ /*29953*/;
  assign _1998_ = inv_5[40] ^ r_4[40] /*29951*/;
  assign sum_5[40] = _1998_ ^ _1997_ /*29950*/;
  assign _1999_ = _1998_ & _1997_ /*29949*/;
  assign _2000_ = inv_5[40] & r_4[40] /*29948*/;
  assign _2001_ = _1999_ | _2000_ /*29947*/;
  assign _2002_ = inv_5[41] ^ r_4[41] /*29945*/;
  assign sum_5[41] = _2002_ ^ _2001_ /*29944*/;
  assign _2003_ = _2002_ & _2001_ /*29943*/;
  assign _2004_ = inv_5[41] & r_4[41] /*29942*/;
  assign _2005_ = _2003_ | _2004_ /*29941*/;
  assign _2006_ = inv_5[42] ^ r_4[42] /*29939*/;
  assign sum_5[42] = _2006_ ^ _2005_ /*29938*/;
  assign _2007_ = _2006_ & _2005_ /*29937*/;
  assign _2008_ = inv_5[42] & r_4[42] /*29936*/;
  assign _2009_ = _2007_ | _2008_ /*29935*/;
  assign _2010_ = inv_5[43] ^ r_4[43] /*29933*/;
  assign sum_5[43] = _2010_ ^ _2009_ /*29932*/;
  assign _2011_ = _2010_ & _2009_ /*29931*/;
  assign _2012_ = inv_5[43] & r_4[43] /*29930*/;
  assign _2013_ = _2011_ | _2012_ /*29929*/;
  assign _2014_ = inv_5[44] ^ r_4[44] /*29927*/;
  assign sum_5[44] = _2014_ ^ _2013_ /*29926*/;
  assign _2015_ = _2014_ & _2013_ /*29925*/;
  assign _2016_ = inv_5[44] & r_4[44] /*29924*/;
  assign _2017_ = _2015_ | _2016_ /*29923*/;
  assign _2018_ = inv_5[45] ^ r_4[45] /*29921*/;
  assign sum_5[45] = _2018_ ^ _2017_ /*29920*/;
  assign _2019_ = _2018_ & _2017_ /*29919*/;
  assign _2020_ = inv_5[45] & r_4[45] /*29918*/;
  assign _2021_ = _2019_ | _2020_ /*29917*/;
  assign _2022_ = inv_5[46] ^ r_4[46] /*29915*/;
  assign sum_5[46] = _2022_ ^ _2021_ /*29914*/;
  assign _2023_ = _2022_ & _2021_ /*29913*/;
  assign _2024_ = inv_5[46] & r_4[46] /*29912*/;
  assign _2025_ = _2023_ | _2024_ /*29911*/;
  assign _2026_ = inv_5[47] ^ r_4[47] /*29909*/;
  assign sum_5[47] = _2026_ ^ _2025_ /*29908*/;
  assign _2027_ = _2026_ & _2025_ /*29907*/;
  assign _2028_ = inv_5[47] & r_4[47] /*29906*/;
  assign _2029_ = _2027_ | _2028_ /*29905*/;
  assign _2030_ = inv_5[48] ^ r_4[48] /*29903*/;
  assign sum_5[48] = _2030_ ^ _2029_ /*29902*/;
  assign _2031_ = _2030_ & _2029_ /*29901*/;
  assign _2032_ = inv_5[48] & r_4[48] /*29900*/;
  assign _2033_ = _2031_ | _2032_ /*29899*/;
  assign _2034_ = inv_5[49] ^ r_4[49] /*29897*/;
  assign sum_5[49] = _2034_ ^ _2033_ /*29896*/;
  assign _2035_ = _2034_ & _2033_ /*29895*/;
  assign _2036_ = inv_5[49] & r_4[49] /*29894*/;
  assign _2037_ = _2035_ | _2036_ /*29893*/;
  assign _2038_ = inv_5[50] ^ r_4[50] /*29891*/;
  assign sum_5[50] = _2038_ ^ _2037_ /*29890*/;
  assign _2039_ = _2038_ & _2037_ /*29889*/;
  assign _2040_ = inv_5[50] & r_4[50] /*29888*/;
  assign _2041_ = _2039_ | _2040_ /*29887*/;
  assign _2042_ = inv_5[51] ^ r_4[51] /*29885*/;
  assign sum_5[51] = _2042_ ^ _2041_ /*29884*/;
  assign _2043_ = _2042_ & _2041_ /*29883*/;
  assign _2044_ = inv_5[51] & r_4[51] /*29882*/;
  assign _2045_ = _2043_ | _2044_ /*29881*/;
  assign _2046_ = inv_5[52] ^ r_4[52] /*29879*/;
  assign sum_5[52] = _2046_ ^ _2045_ /*29878*/;
  assign _2047_ = _2046_ & _2045_ /*29877*/;
  assign _2048_ = inv_5[52] & r_4[52] /*29876*/;
  assign _2049_ = _2047_ | _2048_ /*29875*/;
  assign _2050_ = inv_5[53] ^ r_4[53] /*29873*/;
  assign sum_5[53] = _2050_ ^ _2049_ /*29872*/;
  assign _2051_ = _2050_ & _2049_ /*29871*/;
  assign _2052_ = inv_5[53] & r_4[53] /*29870*/;
  assign _2053_ = _2051_ | _2052_ /*29869*/;
  assign _2054_ = inv_5[54] ^ r_4[54] /*29867*/;
  assign sum_5[54] = _2054_ ^ _2053_ /*29866*/;
  assign _2055_ = _2054_ & _2053_ /*29865*/;
  assign _2056_ = inv_5[54] & r_4[54] /*29864*/;
  assign _2057_ = _2055_ | _2056_ /*29863*/;
  assign _2058_ = inv_5[55] ^ r_4[55] /*29861*/;
  assign sum_5[55] = _2058_ ^ _2057_ /*29860*/;
  assign _2059_ = _2058_ & _2057_ /*29859*/;
  assign _2060_ = inv_5[55] & r_4[55] /*29858*/;
  assign _2061_ = _2059_ | _2060_ /*29857*/;
  assign _2062_ = inv_5[56] ^ r_4[56] /*29855*/;
  assign sum_5[56] = _2062_ ^ _2061_ /*29854*/;
  assign _2063_ = _2062_ & _2061_ /*29853*/;
  assign _2064_ = inv_5[56] & r_4[56] /*29852*/;
  assign _2065_ = _2063_ | _2064_ /*29851*/;
  assign _2066_ = inv_5[57] ^ r_4[57] /*29849*/;
  assign sum_5[57] = _2066_ ^ _2065_ /*29848*/;
  assign _2067_ = _2066_ & _2065_ /*29847*/;
  assign _2068_ = inv_5[57] & r_4[57] /*29846*/;
  assign _2069_ = _2067_ | _2068_ /*29845*/;
  assign _2070_ = inv_5[58] ^ r_4[58] /*29843*/;
  assign sum_5[58] = _2070_ ^ _2069_ /*29842*/;
  assign _2071_ = _2070_ & _2069_ /*29841*/;
  assign _2072_ = inv_5[58] & r_4[58] /*29840*/;
  assign _2073_ = _2071_ | _2072_ /*29839*/;
  assign _2074_ = inv_5[59] ^ r_4[59] /*29837*/;
  assign sum_5[59] = _2074_ ^ _2073_ /*29836*/;
  assign _2075_ = _2074_ & _2073_ /*29835*/;
  assign _2076_ = inv_5[59] & r_4[59] /*29834*/;
  assign _2077_ = _2075_ | _2076_ /*29833*/;
  assign _2078_ = inv_5[60] ^ r_4[60] /*29831*/;
  assign sum_5[60] = _2078_ ^ _2077_ /*29830*/;
  assign _2079_ = _2078_ & _2077_ /*29829*/;
  assign _2080_ = inv_5[60] & r_4[60] /*29828*/;
  assign _2081_ = _2079_ | _2080_ /*29827*/;
  assign _2082_ = inv_5[61] ^ r_4[61] /*29825*/;
  assign sum_5[61] = _2082_ ^ _2081_ /*29824*/;
  assign _2083_ = _2082_ & _2081_ /*29823*/;
  assign _2084_ = inv_5[61] & r_4[61] /*29822*/;
  assign _2085_ = _2083_ | _2084_ /*29821*/;
  assign _2086_ = inv_5[62] ^ r_4[62] /*29819*/;
  assign sum_5[62] = _2086_ ^ _2085_ /*29818*/;
  assign _2087_ = _2086_ & _2085_ /*29817*/;
  assign _2088_ = inv_5[62] & r_4[62] /*29816*/;
  assign _2089_ = _2087_ | _2088_ /*29815*/;
  assign _2090_ = inv_5[63] ^ r_4[63] /*29813*/;
  assign sum_5[63] = _2090_ ^ _2089_ /*29812*/;
  assign _2091_ = _2090_ & _2089_ /*29811*/;
  assign _2092_ = inv_5[63] & r_4[63] /*29810*/;
  assign _2093_ = _2091_ | _2092_ /*29809*/;
  assign _2094_ = inv_5[64] ^ r_4[64] /*29807*/;
  assign sum_5[64] = _2094_ ^ _2093_ /*29806*/;
  assign _2095_ = _2094_ & _2093_ /*29805*/;
  assign _2096_ = inv_5[64] & r_4[64] /*29804*/;
  assign _2097_ = _2095_ | _2096_ /*29803*/;
  assign _2098_ = inv_5[65] ^ r_4[65] /*29801*/;
  assign sum_5[65] = _2098_ ^ _2097_ /*29800*/;
  assign _2099_ = _2098_ & _2097_ /*29799*/;
  assign _2100_ = inv_5[65] & r_4[65] /*29798*/;
  assign _2101_ = _2099_ | _2100_ /*29797*/;
  assign _2102_ = inv_5[66] ^ r_4[66] /*29795*/;
  assign sum_5[66] = _2102_ ^ _2101_ /*29794*/;
  assign _2103_ = _2102_ & _2101_ /*29793*/;
  assign _2104_ = inv_5[66] & r_4[66] /*29792*/;
  assign _2105_ = _2103_ | _2104_ /*29791*/;
  assign _2106_ = _2105_ ^ _2101_ /*29790*/;
  assign _2107_ = ~_2106_ /*29789*/;
  assign _2108_ = sum_5[66] & _2107_ /*29788*/;
  assign _2109_ = _2106_ & _2105_ /*29787*/;
  assign sum_5[67] = _2109_ | _2108_ /*29786*/;
  assign q[27] = ~sum_5[67] /*29785*/;
  assign m_5[0] = r_4[0] /*29784*/;
  assign m_5[1] = r_4[1] /*29783*/;
  assign m_5[2] = r_4[2] /*29782*/;
  assign m_5[3] = r_4[3] /*29781*/;
  assign m_5[4] = r_4[4] /*29780*/;
  assign m_5[5] = r_4[5] /*29779*/;
  assign m_5[6] = r_4[6] /*29778*/;
  assign m_5[7] = r_4[7] /*29777*/;
  assign m_5[8] = r_4[8] /*29776*/;
  assign m_5[9] = r_4[9] /*29775*/;
  assign m_5[10] = r_4[10] /*29774*/;
  assign m_5[11] = r_4[11] /*29773*/;
  assign m_5[12] = r_4[12] /*29772*/;
  assign m_5[13] = r_4[13] /*29771*/;
  assign m_5[14] = r_4[14] /*29770*/;
  assign m_5[15] = r_4[15] /*29769*/;
  assign m_5[16] = r_4[16] /*29768*/;
  assign m_5[17] = r_4[17] /*29767*/;
  assign m_5[18] = r_4[18] /*29766*/;
  assign m_5[19] = r_4[19] /*29765*/;
  assign m_5[20] = r_4[20] /*29764*/;
  assign m_5[21] = r_4[21] /*29763*/;
  assign m_5[22] = r_4[22] /*29762*/;
  assign m_5[23] = r_4[23] /*29761*/;
  assign m_5[24] = r_4[24] /*29760*/;
  assign m_5[25] = r_4[25] /*29759*/;
  assign m_5[26] = r_4[26] /*29758*/;
  assign m_5[27] = r_4[27] /*29757*/;
  assign m_5[28] = r_4[28] /*29756*/;
  assign m_5[29] = r_4[29] /*29755*/;
  assign m_5[30] = r_4[30] /*29754*/;
  assign m_5[31] = r_4[31] /*29753*/;
  assign m_5[32] = r_4[32] /*29752*/;
  assign m_5[33] = r_4[33] /*29751*/;
  assign m_5[34] = r_4[34] /*29750*/;
  assign m_5[35] = r_4[35] /*29749*/;
  assign m_5[36] = r_4[36] /*29748*/;
  assign m_5[37] = r_4[37] /*29747*/;
  assign m_5[38] = r_4[38] /*29746*/;
  assign m_5[39] = r_4[39] /*29745*/;
  assign m_5[40] = r_4[40] /*29744*/;
  assign m_5[41] = r_4[41] /*29743*/;
  assign m_5[42] = r_4[42] /*29742*/;
  assign m_5[43] = r_4[43] /*29741*/;
  assign m_5[44] = r_4[44] /*29740*/;
  assign m_5[45] = r_4[45] /*29739*/;
  assign m_5[46] = r_4[46] /*29738*/;
  assign m_5[47] = r_4[47] /*29737*/;
  assign m_5[48] = r_4[48] /*29736*/;
  assign m_5[49] = r_4[49] /*29735*/;
  assign m_5[50] = r_4[50] /*29734*/;
  assign m_5[51] = r_4[51] /*29733*/;
  assign m_5[52] = r_4[52] /*29732*/;
  assign m_5[53] = r_4[53] /*29731*/;
  assign m_5[54] = r_4[54] /*29730*/;
  assign m_5[55] = r_4[55] /*29729*/;
  assign m_5[56] = r_4[56] /*29728*/;
  assign m_5[57] = r_4[57] /*29727*/;
  assign m_5[58] = r_4[58] /*29726*/;
  assign m_5[59] = r_4[59] /*29725*/;
  assign m_5[60] = r_4[60] /*29724*/;
  assign m_5[61] = r_4[61] /*29723*/;
  assign m_5[62] = r_4[62] /*29722*/;
  assign m_5[63] = r_4[63] /*29721*/;
  assign m_5[64] = r_4[64] /*29720*/;
  assign m_5[65] = r_4[65] /*29719*/;
  assign m_5[66] = r_4[66] /*29718*/;
  assign m_5[67] = r_4[66] /*29717*/;
  assign _2111_ = ~q[27] /*29716*/;
  assign _2112_ = sum_5[0] & q[27] /*29715*/;
  assign _2113_ = m_5[0] & _2111_ /*29714*/;
  assign r_5[0] = _2113_ | _2112_ /*29713*/;
  assign _2114_ = ~q[27] /*29712*/;
  assign _2115_ = sum_5[1] & q[27] /*29711*/;
  assign _2116_ = m_5[1] & _2114_ /*29710*/;
  assign r_5[1] = _2116_ | _2115_ /*29709*/;
  assign _2117_ = ~q[27] /*29708*/;
  assign _2118_ = sum_5[2] & q[27] /*29707*/;
  assign _2119_ = m_5[2] & _2117_ /*29706*/;
  assign r_5[2] = _2119_ | _2118_ /*29705*/;
  assign _2120_ = ~q[27] /*29704*/;
  assign _2121_ = sum_5[3] & q[27] /*29703*/;
  assign _2122_ = m_5[3] & _2120_ /*29702*/;
  assign r_5[3] = _2122_ | _2121_ /*29701*/;
  assign _2123_ = ~q[27] /*29700*/;
  assign _2124_ = sum_5[4] & q[27] /*29699*/;
  assign _2125_ = m_5[4] & _2123_ /*29698*/;
  assign r_5[4] = _2125_ | _2124_ /*29697*/;
  assign _2126_ = ~q[27] /*29696*/;
  assign _2127_ = sum_5[5] & q[27] /*29695*/;
  assign _2128_ = m_5[5] & _2126_ /*29694*/;
  assign r_5[5] = _2128_ | _2127_ /*29693*/;
  assign _2129_ = ~q[27] /*29692*/;
  assign _2130_ = sum_5[6] & q[27] /*29691*/;
  assign _2131_ = m_5[6] & _2129_ /*29690*/;
  assign r_5[6] = _2131_ | _2130_ /*29689*/;
  assign _2132_ = ~q[27] /*29688*/;
  assign _2133_ = sum_5[7] & q[27] /*29687*/;
  assign _2134_ = m_5[7] & _2132_ /*29686*/;
  assign r_5[7] = _2134_ | _2133_ /*29685*/;
  assign _2135_ = ~q[27] /*29684*/;
  assign _2136_ = sum_5[8] & q[27] /*29683*/;
  assign _2137_ = m_5[8] & _2135_ /*29682*/;
  assign r_5[8] = _2137_ | _2136_ /*29681*/;
  assign _2138_ = ~q[27] /*29680*/;
  assign _2139_ = sum_5[9] & q[27] /*29679*/;
  assign _2140_ = m_5[9] & _2138_ /*29678*/;
  assign r_5[9] = _2140_ | _2139_ /*29677*/;
  assign _2141_ = ~q[27] /*29676*/;
  assign _2142_ = sum_5[10] & q[27] /*29675*/;
  assign _2143_ = m_5[10] & _2141_ /*29674*/;
  assign r_5[10] = _2143_ | _2142_ /*29673*/;
  assign _2144_ = ~q[27] /*29672*/;
  assign _2145_ = sum_5[11] & q[27] /*29671*/;
  assign _2146_ = m_5[11] & _2144_ /*29670*/;
  assign r_5[11] = _2146_ | _2145_ /*29669*/;
  assign _2147_ = ~q[27] /*29668*/;
  assign _2148_ = sum_5[12] & q[27] /*29667*/;
  assign _2149_ = m_5[12] & _2147_ /*29666*/;
  assign r_5[12] = _2149_ | _2148_ /*29665*/;
  assign _2150_ = ~q[27] /*29664*/;
  assign _2151_ = sum_5[13] & q[27] /*29663*/;
  assign _2152_ = m_5[13] & _2150_ /*29662*/;
  assign r_5[13] = _2152_ | _2151_ /*29661*/;
  assign _2153_ = ~q[27] /*29660*/;
  assign _2154_ = sum_5[14] & q[27] /*29659*/;
  assign _2155_ = m_5[14] & _2153_ /*29658*/;
  assign r_5[14] = _2155_ | _2154_ /*29657*/;
  assign _2156_ = ~q[27] /*29656*/;
  assign _2157_ = sum_5[15] & q[27] /*29655*/;
  assign _2158_ = m_5[15] & _2156_ /*29654*/;
  assign r_5[15] = _2158_ | _2157_ /*29653*/;
  assign _2159_ = ~q[27] /*29652*/;
  assign _2160_ = sum_5[16] & q[27] /*29651*/;
  assign _2161_ = m_5[16] & _2159_ /*29650*/;
  assign r_5[16] = _2161_ | _2160_ /*29649*/;
  assign _2162_ = ~q[27] /*29648*/;
  assign _2163_ = sum_5[17] & q[27] /*29647*/;
  assign _2164_ = m_5[17] & _2162_ /*29646*/;
  assign r_5[17] = _2164_ | _2163_ /*29645*/;
  assign _2165_ = ~q[27] /*29644*/;
  assign _2166_ = sum_5[18] & q[27] /*29643*/;
  assign _2167_ = m_5[18] & _2165_ /*29642*/;
  assign r_5[18] = _2167_ | _2166_ /*29641*/;
  assign _2168_ = ~q[27] /*29640*/;
  assign _2169_ = sum_5[19] & q[27] /*29639*/;
  assign _2170_ = m_5[19] & _2168_ /*29638*/;
  assign r_5[19] = _2170_ | _2169_ /*29637*/;
  assign _2171_ = ~q[27] /*29636*/;
  assign _2172_ = sum_5[20] & q[27] /*29635*/;
  assign _2173_ = m_5[20] & _2171_ /*29634*/;
  assign r_5[20] = _2173_ | _2172_ /*29633*/;
  assign _2174_ = ~q[27] /*29632*/;
  assign _2175_ = sum_5[21] & q[27] /*29631*/;
  assign _2176_ = m_5[21] & _2174_ /*29630*/;
  assign r_5[21] = _2176_ | _2175_ /*29629*/;
  assign _2177_ = ~q[27] /*29628*/;
  assign _2178_ = sum_5[22] & q[27] /*29627*/;
  assign _2179_ = m_5[22] & _2177_ /*29626*/;
  assign r_5[22] = _2179_ | _2178_ /*29625*/;
  assign _2180_ = ~q[27] /*29624*/;
  assign _2181_ = sum_5[23] & q[27] /*29623*/;
  assign _2182_ = m_5[23] & _2180_ /*29622*/;
  assign r_5[23] = _2182_ | _2181_ /*29621*/;
  assign _2183_ = ~q[27] /*29620*/;
  assign _2184_ = sum_5[24] & q[27] /*29619*/;
  assign _2185_ = m_5[24] & _2183_ /*29618*/;
  assign r_5[24] = _2185_ | _2184_ /*29617*/;
  assign _2186_ = ~q[27] /*29616*/;
  assign _2187_ = sum_5[25] & q[27] /*29615*/;
  assign _2188_ = m_5[25] & _2186_ /*29614*/;
  assign r_5[25] = _2188_ | _2187_ /*29613*/;
  assign _2189_ = ~q[27] /*29612*/;
  assign _2190_ = sum_5[26] & q[27] /*29611*/;
  assign _2191_ = m_5[26] & _2189_ /*29610*/;
  assign r_5[26] = _2191_ | _2190_ /*29609*/;
  assign _2192_ = ~q[27] /*29608*/;
  assign _2193_ = sum_5[27] & q[27] /*29607*/;
  assign _2194_ = m_5[27] & _2192_ /*29606*/;
  assign r_5[27] = _2194_ | _2193_ /*29605*/;
  assign _2195_ = ~q[27] /*29604*/;
  assign _2196_ = sum_5[28] & q[27] /*29603*/;
  assign _2197_ = m_5[28] & _2195_ /*29602*/;
  assign r_5[28] = _2197_ | _2196_ /*29601*/;
  assign _2198_ = ~q[27] /*29600*/;
  assign _2199_ = sum_5[29] & q[27] /*29599*/;
  assign _2200_ = m_5[29] & _2198_ /*29598*/;
  assign r_5[29] = _2200_ | _2199_ /*29597*/;
  assign _2201_ = ~q[27] /*29596*/;
  assign _2202_ = sum_5[30] & q[27] /*29595*/;
  assign _2203_ = m_5[30] & _2201_ /*29594*/;
  assign r_5[30] = _2203_ | _2202_ /*29593*/;
  assign _2204_ = ~q[27] /*29592*/;
  assign _2205_ = sum_5[31] & q[27] /*29591*/;
  assign _2206_ = m_5[31] & _2204_ /*29590*/;
  assign r_5[31] = _2206_ | _2205_ /*29589*/;
  assign _2207_ = ~q[27] /*29588*/;
  assign _2208_ = sum_5[32] & q[27] /*29587*/;
  assign _2209_ = m_5[32] & _2207_ /*29586*/;
  assign r_5[32] = _2209_ | _2208_ /*29585*/;
  assign _2210_ = ~q[27] /*29584*/;
  assign _2211_ = sum_5[33] & q[27] /*29583*/;
  assign _2212_ = m_5[33] & _2210_ /*29582*/;
  assign r_5[33] = _2212_ | _2211_ /*29581*/;
  assign _2213_ = ~q[27] /*29580*/;
  assign _2214_ = sum_5[34] & q[27] /*29579*/;
  assign _2215_ = m_5[34] & _2213_ /*29578*/;
  assign r_5[34] = _2215_ | _2214_ /*29577*/;
  assign _2216_ = ~q[27] /*29576*/;
  assign _2217_ = sum_5[35] & q[27] /*29575*/;
  assign _2218_ = m_5[35] & _2216_ /*29574*/;
  assign r_5[35] = _2218_ | _2217_ /*29573*/;
  assign _2219_ = ~q[27] /*29572*/;
  assign _2220_ = sum_5[36] & q[27] /*29571*/;
  assign _2221_ = m_5[36] & _2219_ /*29570*/;
  assign r_5[36] = _2221_ | _2220_ /*29569*/;
  assign _2222_ = ~q[27] /*29568*/;
  assign _2223_ = sum_5[37] & q[27] /*29567*/;
  assign _2224_ = m_5[37] & _2222_ /*29566*/;
  assign r_5[37] = _2224_ | _2223_ /*29565*/;
  assign _2225_ = ~q[27] /*29564*/;
  assign _2226_ = sum_5[38] & q[27] /*29563*/;
  assign _2227_ = m_5[38] & _2225_ /*29562*/;
  assign r_5[38] = _2227_ | _2226_ /*29561*/;
  assign _2228_ = ~q[27] /*29560*/;
  assign _2229_ = sum_5[39] & q[27] /*29559*/;
  assign _2230_ = m_5[39] & _2228_ /*29558*/;
  assign r_5[39] = _2230_ | _2229_ /*29557*/;
  assign _2231_ = ~q[27] /*29556*/;
  assign _2232_ = sum_5[40] & q[27] /*29555*/;
  assign _2233_ = m_5[40] & _2231_ /*29554*/;
  assign r_5[40] = _2233_ | _2232_ /*29553*/;
  assign _2234_ = ~q[27] /*29552*/;
  assign _2235_ = sum_5[41] & q[27] /*29551*/;
  assign _2236_ = m_5[41] & _2234_ /*29550*/;
  assign r_5[41] = _2236_ | _2235_ /*29549*/;
  assign _2237_ = ~q[27] /*29548*/;
  assign _2238_ = sum_5[42] & q[27] /*29547*/;
  assign _2239_ = m_5[42] & _2237_ /*29546*/;
  assign r_5[42] = _2239_ | _2238_ /*29545*/;
  assign _2240_ = ~q[27] /*29544*/;
  assign _2241_ = sum_5[43] & q[27] /*29543*/;
  assign _2242_ = m_5[43] & _2240_ /*29542*/;
  assign r_5[43] = _2242_ | _2241_ /*29541*/;
  assign _2243_ = ~q[27] /*29540*/;
  assign _2244_ = sum_5[44] & q[27] /*29539*/;
  assign _2245_ = m_5[44] & _2243_ /*29538*/;
  assign r_5[44] = _2245_ | _2244_ /*29537*/;
  assign _2246_ = ~q[27] /*29536*/;
  assign _2247_ = sum_5[45] & q[27] /*29535*/;
  assign _2248_ = m_5[45] & _2246_ /*29534*/;
  assign r_5[45] = _2248_ | _2247_ /*29533*/;
  assign _2249_ = ~q[27] /*29532*/;
  assign _2250_ = sum_5[46] & q[27] /*29531*/;
  assign _2251_ = m_5[46] & _2249_ /*29530*/;
  assign r_5[46] = _2251_ | _2250_ /*29529*/;
  assign _2252_ = ~q[27] /*29528*/;
  assign _2253_ = sum_5[47] & q[27] /*29527*/;
  assign _2254_ = m_5[47] & _2252_ /*29526*/;
  assign r_5[47] = _2254_ | _2253_ /*29525*/;
  assign _2255_ = ~q[27] /*29524*/;
  assign _2256_ = sum_5[48] & q[27] /*29523*/;
  assign _2257_ = m_5[48] & _2255_ /*29522*/;
  assign r_5[48] = _2257_ | _2256_ /*29521*/;
  assign _2258_ = ~q[27] /*29520*/;
  assign _2259_ = sum_5[49] & q[27] /*29519*/;
  assign _2260_ = m_5[49] & _2258_ /*29518*/;
  assign r_5[49] = _2260_ | _2259_ /*29517*/;
  assign _2261_ = ~q[27] /*29516*/;
  assign _2262_ = sum_5[50] & q[27] /*29515*/;
  assign _2263_ = m_5[50] & _2261_ /*29514*/;
  assign r_5[50] = _2263_ | _2262_ /*29513*/;
  assign _2264_ = ~q[27] /*29512*/;
  assign _2265_ = sum_5[51] & q[27] /*29511*/;
  assign _2266_ = m_5[51] & _2264_ /*29510*/;
  assign r_5[51] = _2266_ | _2265_ /*29509*/;
  assign _2267_ = ~q[27] /*29508*/;
  assign _2268_ = sum_5[52] & q[27] /*29507*/;
  assign _2269_ = m_5[52] & _2267_ /*29506*/;
  assign r_5[52] = _2269_ | _2268_ /*29505*/;
  assign _2270_ = ~q[27] /*29504*/;
  assign _2271_ = sum_5[53] & q[27] /*29503*/;
  assign _2272_ = m_5[53] & _2270_ /*29502*/;
  assign r_5[53] = _2272_ | _2271_ /*29501*/;
  assign _2273_ = ~q[27] /*29500*/;
  assign _2274_ = sum_5[54] & q[27] /*29499*/;
  assign _2275_ = m_5[54] & _2273_ /*29498*/;
  assign r_5[54] = _2275_ | _2274_ /*29497*/;
  assign _2276_ = ~q[27] /*29496*/;
  assign _2277_ = sum_5[55] & q[27] /*29495*/;
  assign _2278_ = m_5[55] & _2276_ /*29494*/;
  assign r_5[55] = _2278_ | _2277_ /*29493*/;
  assign _2279_ = ~q[27] /*29492*/;
  assign _2280_ = sum_5[56] & q[27] /*29491*/;
  assign _2281_ = m_5[56] & _2279_ /*29490*/;
  assign r_5[56] = _2281_ | _2280_ /*29489*/;
  assign _2282_ = ~q[27] /*29488*/;
  assign _2283_ = sum_5[57] & q[27] /*29487*/;
  assign _2284_ = m_5[57] & _2282_ /*29486*/;
  assign r_5[57] = _2284_ | _2283_ /*29485*/;
  assign _2285_ = ~q[27] /*29484*/;
  assign _2286_ = sum_5[58] & q[27] /*29483*/;
  assign _2287_ = m_5[58] & _2285_ /*29482*/;
  assign r_5[58] = _2287_ | _2286_ /*29481*/;
  assign _2288_ = ~q[27] /*29480*/;
  assign _2289_ = sum_5[59] & q[27] /*29479*/;
  assign _2290_ = m_5[59] & _2288_ /*29478*/;
  assign r_5[59] = _2290_ | _2289_ /*29477*/;
  assign _2291_ = ~q[27] /*29476*/;
  assign _2292_ = sum_5[60] & q[27] /*29475*/;
  assign _2293_ = m_5[60] & _2291_ /*29474*/;
  assign r_5[60] = _2293_ | _2292_ /*29473*/;
  assign _2294_ = ~q[27] /*29472*/;
  assign _2295_ = sum_5[61] & q[27] /*29471*/;
  assign _2296_ = m_5[61] & _2294_ /*29470*/;
  assign r_5[61] = _2296_ | _2295_ /*29469*/;
  assign _2297_ = ~q[27] /*29468*/;
  assign _2298_ = sum_5[62] & q[27] /*29467*/;
  assign _2299_ = m_5[62] & _2297_ /*29466*/;
  assign r_5[62] = _2299_ | _2298_ /*29465*/;
  assign _2300_ = ~q[27] /*29464*/;
  assign _2301_ = sum_5[63] & q[27] /*29463*/;
  assign _2302_ = m_5[63] & _2300_ /*29462*/;
  assign r_5[63] = _2302_ | _2301_ /*29461*/;
  assign _2303_ = ~q[27] /*29460*/;
  assign _2304_ = sum_5[64] & q[27] /*29459*/;
  assign _2305_ = m_5[64] & _2303_ /*29458*/;
  assign r_5[64] = _2305_ | _2304_ /*29457*/;
  assign _2306_ = ~q[27] /*29456*/;
  assign _2307_ = sum_5[65] & q[27] /*29455*/;
  assign _2308_ = m_5[65] & _2306_ /*29454*/;
  assign r_5[65] = _2308_ | _2307_ /*29453*/;
  assign _2309_ = ~q[27] /*29452*/;
  assign _2310_ = sum_5[66] & q[27] /*29451*/;
  assign _2311_ = m_5[66] & _2309_ /*29450*/;
  assign r_5[66] = _2311_ | _2310_ /*29449*/;
  assign _2312_ = ~q[27] /*29448*/;
  assign _2313_ = sum_5[67] & q[27] /*29447*/;
  assign _2314_ = m_5[67] & _2312_ /*29446*/;
  assign r_5[67] = _2314_ | _2313_ /*29445*/;
  assign inv_6[0] = oneWire /*29116*/;
  assign inv_6[1] = oneWire /*29110*/;
  assign inv_6[2] = oneWire /*29104*/;
  assign inv_6[3] = oneWire /*29098*/;
  assign inv_6[4] = oneWire /*29092*/;
  assign inv_6[5] = oneWire /*29086*/;
  assign inv_6[6] = oneWire /*29080*/;
  assign inv_6[7] = oneWire /*29074*/;
  assign inv_6[8] = oneWire /*29068*/;
  assign inv_6[9] = oneWire /*29062*/;
  assign inv_6[10] = oneWire /*29056*/;
  assign inv_6[11] = oneWire /*29050*/;
  assign inv_6[12] = oneWire /*29044*/;
  assign inv_6[13] = oneWire /*29038*/;
  assign inv_6[14] = oneWire /*29032*/;
  assign inv_6[15] = oneWire /*29026*/;
  assign inv_6[16] = oneWire /*29020*/;
  assign inv_6[17] = oneWire /*29014*/;
  assign inv_6[18] = oneWire /*29008*/;
  assign inv_6[19] = oneWire /*29002*/;
  assign inv_6[20] = oneWire /*28996*/;
  assign inv_6[21] = oneWire /*28990*/;
  assign inv_6[22] = oneWire /*28984*/;
  assign inv_6[23] = oneWire /*28978*/;
  assign inv_6[24] = oneWire /*28972*/;
  assign inv_6[25] = oneWire /*28966*/;
  assign inv_6[26] = ~div[0] /*28960*/;
  assign inv_6[27] = ~div[1] /*28954*/;
  assign inv_6[28] = ~div[2] /*28948*/;
  assign inv_6[29] = ~div[3] /*28942*/;
  assign inv_6[30] = ~div[4] /*28936*/;
  assign inv_6[31] = ~div[5] /*28930*/;
  assign inv_6[32] = ~div[6] /*28924*/;
  assign inv_6[33] = ~div[7] /*28918*/;
  assign inv_6[34] = ~div[8] /*28912*/;
  assign inv_6[35] = ~div[9] /*28906*/;
  assign inv_6[36] = ~div[10] /*28900*/;
  assign inv_6[37] = ~div[11] /*28894*/;
  assign inv_6[38] = ~div[12] /*28888*/;
  assign inv_6[39] = ~div[13] /*28882*/;
  assign inv_6[40] = ~div[14] /*28876*/;
  assign inv_6[41] = ~div[15] /*28870*/;
  assign inv_6[42] = ~div[16] /*28864*/;
  assign inv_6[43] = ~div[17] /*28858*/;
  assign inv_6[44] = ~div[18] /*28852*/;
  assign inv_6[45] = ~div[19] /*28846*/;
  assign inv_6[46] = ~div[20] /*28840*/;
  assign inv_6[47] = ~div[21] /*28834*/;
  assign inv_6[48] = ~div[22] /*28828*/;
  assign inv_6[49] = ~div[23] /*28822*/;
  assign inv_6[50] = ~div[24] /*28816*/;
  assign inv_6[51] = ~div[25] /*28810*/;
  assign inv_6[52] = ~div[26] /*28804*/;
  assign inv_6[53] = ~div[27] /*28798*/;
  assign inv_6[54] = ~div[28] /*28792*/;
  assign inv_6[55] = ~div[29] /*28786*/;
  assign inv_6[56] = ~div[30] /*28780*/;
  assign inv_6[57] = oneWire /*28774*/;
  assign inv_6[58] = oneWire /*28768*/;
  assign inv_6[59] = oneWire /*28762*/;
  assign inv_6[60] = oneWire /*28756*/;
  assign inv_6[61] = oneWire /*28750*/;
  assign inv_6[62] = oneWire /*28744*/;
  assign inv_6[63] = oneWire /*28738*/;
  assign inv_6[64] = oneWire /*28732*/;
  assign inv_6[65] = oneWire /*28726*/;
  assign inv_6[66] = oneWire /*28720*/;
  assign inv_6[67] = oneWire /*28714*/;
  assign _2315_ = inv_6[0] ^ r_5[0] /*29115*/;
  assign sum_6[0] = _2315_ ^ oneWire /*29114*/;
  assign _2316_ = _2315_ & oneWire /*29113*/;
  assign _2317_ = inv_6[0] & r_5[0] /*29112*/;
  assign _2318_ = _2316_ | _2317_ /*29111*/;
  assign _2319_ = inv_6[1] ^ r_5[1] /*29109*/;
  assign sum_6[1] = _2319_ ^ _2318_ /*29108*/;
  assign _2320_ = _2319_ & _2318_ /*29107*/;
  assign _2321_ = inv_6[1] & r_5[1] /*29106*/;
  assign _2322_ = _2320_ | _2321_ /*29105*/;
  assign _2323_ = inv_6[2] ^ r_5[2] /*29103*/;
  assign sum_6[2] = _2323_ ^ _2322_ /*29102*/;
  assign _2324_ = _2323_ & _2322_ /*29101*/;
  assign _2325_ = inv_6[2] & r_5[2] /*29100*/;
  assign _2326_ = _2324_ | _2325_ /*29099*/;
  assign _2327_ = inv_6[3] ^ r_5[3] /*29097*/;
  assign sum_6[3] = _2327_ ^ _2326_ /*29096*/;
  assign _2328_ = _2327_ & _2326_ /*29095*/;
  assign _2329_ = inv_6[3] & r_5[3] /*29094*/;
  assign _2330_ = _2328_ | _2329_ /*29093*/;
  assign _2331_ = inv_6[4] ^ r_5[4] /*29091*/;
  assign sum_6[4] = _2331_ ^ _2330_ /*29090*/;
  assign _2332_ = _2331_ & _2330_ /*29089*/;
  assign _2333_ = inv_6[4] & r_5[4] /*29088*/;
  assign _2334_ = _2332_ | _2333_ /*29087*/;
  assign _2335_ = inv_6[5] ^ r_5[5] /*29085*/;
  assign sum_6[5] = _2335_ ^ _2334_ /*29084*/;
  assign _2336_ = _2335_ & _2334_ /*29083*/;
  assign _2337_ = inv_6[5] & r_5[5] /*29082*/;
  assign _2338_ = _2336_ | _2337_ /*29081*/;
  assign _2339_ = inv_6[6] ^ r_5[6] /*29079*/;
  assign sum_6[6] = _2339_ ^ _2338_ /*29078*/;
  assign _2340_ = _2339_ & _2338_ /*29077*/;
  assign _2341_ = inv_6[6] & r_5[6] /*29076*/;
  assign _2342_ = _2340_ | _2341_ /*29075*/;
  assign _2343_ = inv_6[7] ^ r_5[7] /*29073*/;
  assign sum_6[7] = _2343_ ^ _2342_ /*29072*/;
  assign _2344_ = _2343_ & _2342_ /*29071*/;
  assign _2345_ = inv_6[7] & r_5[7] /*29070*/;
  assign _2346_ = _2344_ | _2345_ /*29069*/;
  assign _2347_ = inv_6[8] ^ r_5[8] /*29067*/;
  assign sum_6[8] = _2347_ ^ _2346_ /*29066*/;
  assign _2348_ = _2347_ & _2346_ /*29065*/;
  assign _2349_ = inv_6[8] & r_5[8] /*29064*/;
  assign _2350_ = _2348_ | _2349_ /*29063*/;
  assign _2351_ = inv_6[9] ^ r_5[9] /*29061*/;
  assign sum_6[9] = _2351_ ^ _2350_ /*29060*/;
  assign _2352_ = _2351_ & _2350_ /*29059*/;
  assign _2353_ = inv_6[9] & r_5[9] /*29058*/;
  assign _2354_ = _2352_ | _2353_ /*29057*/;
  assign _2355_ = inv_6[10] ^ r_5[10] /*29055*/;
  assign sum_6[10] = _2355_ ^ _2354_ /*29054*/;
  assign _2356_ = _2355_ & _2354_ /*29053*/;
  assign _2357_ = inv_6[10] & r_5[10] /*29052*/;
  assign _2358_ = _2356_ | _2357_ /*29051*/;
  assign _2359_ = inv_6[11] ^ r_5[11] /*29049*/;
  assign sum_6[11] = _2359_ ^ _2358_ /*29048*/;
  assign _2360_ = _2359_ & _2358_ /*29047*/;
  assign _2361_ = inv_6[11] & r_5[11] /*29046*/;
  assign _2362_ = _2360_ | _2361_ /*29045*/;
  assign _2363_ = inv_6[12] ^ r_5[12] /*29043*/;
  assign sum_6[12] = _2363_ ^ _2362_ /*29042*/;
  assign _2364_ = _2363_ & _2362_ /*29041*/;
  assign _2365_ = inv_6[12] & r_5[12] /*29040*/;
  assign _2366_ = _2364_ | _2365_ /*29039*/;
  assign _2367_ = inv_6[13] ^ r_5[13] /*29037*/;
  assign sum_6[13] = _2367_ ^ _2366_ /*29036*/;
  assign _2368_ = _2367_ & _2366_ /*29035*/;
  assign _2369_ = inv_6[13] & r_5[13] /*29034*/;
  assign _2370_ = _2368_ | _2369_ /*29033*/;
  assign _2371_ = inv_6[14] ^ r_5[14] /*29031*/;
  assign sum_6[14] = _2371_ ^ _2370_ /*29030*/;
  assign _2372_ = _2371_ & _2370_ /*29029*/;
  assign _2373_ = inv_6[14] & r_5[14] /*29028*/;
  assign _2374_ = _2372_ | _2373_ /*29027*/;
  assign _2375_ = inv_6[15] ^ r_5[15] /*29025*/;
  assign sum_6[15] = _2375_ ^ _2374_ /*29024*/;
  assign _2376_ = _2375_ & _2374_ /*29023*/;
  assign _2377_ = inv_6[15] & r_5[15] /*29022*/;
  assign _2378_ = _2376_ | _2377_ /*29021*/;
  assign _2379_ = inv_6[16] ^ r_5[16] /*29019*/;
  assign sum_6[16] = _2379_ ^ _2378_ /*29018*/;
  assign _2380_ = _2379_ & _2378_ /*29017*/;
  assign _2381_ = inv_6[16] & r_5[16] /*29016*/;
  assign _2382_ = _2380_ | _2381_ /*29015*/;
  assign _2383_ = inv_6[17] ^ r_5[17] /*29013*/;
  assign sum_6[17] = _2383_ ^ _2382_ /*29012*/;
  assign _2384_ = _2383_ & _2382_ /*29011*/;
  assign _2385_ = inv_6[17] & r_5[17] /*29010*/;
  assign _2386_ = _2384_ | _2385_ /*29009*/;
  assign _2387_ = inv_6[18] ^ r_5[18] /*29007*/;
  assign sum_6[18] = _2387_ ^ _2386_ /*29006*/;
  assign _2388_ = _2387_ & _2386_ /*29005*/;
  assign _2389_ = inv_6[18] & r_5[18] /*29004*/;
  assign _2390_ = _2388_ | _2389_ /*29003*/;
  assign _2391_ = inv_6[19] ^ r_5[19] /*29001*/;
  assign sum_6[19] = _2391_ ^ _2390_ /*29000*/;
  assign _2392_ = _2391_ & _2390_ /*28999*/;
  assign _2393_ = inv_6[19] & r_5[19] /*28998*/;
  assign _2394_ = _2392_ | _2393_ /*28997*/;
  assign _2395_ = inv_6[20] ^ r_5[20] /*28995*/;
  assign sum_6[20] = _2395_ ^ _2394_ /*28994*/;
  assign _2396_ = _2395_ & _2394_ /*28993*/;
  assign _2397_ = inv_6[20] & r_5[20] /*28992*/;
  assign _2398_ = _2396_ | _2397_ /*28991*/;
  assign _2399_ = inv_6[21] ^ r_5[21] /*28989*/;
  assign sum_6[21] = _2399_ ^ _2398_ /*28988*/;
  assign _2400_ = _2399_ & _2398_ /*28987*/;
  assign _2401_ = inv_6[21] & r_5[21] /*28986*/;
  assign _2402_ = _2400_ | _2401_ /*28985*/;
  assign _2403_ = inv_6[22] ^ r_5[22] /*28983*/;
  assign sum_6[22] = _2403_ ^ _2402_ /*28982*/;
  assign _2404_ = _2403_ & _2402_ /*28981*/;
  assign _2405_ = inv_6[22] & r_5[22] /*28980*/;
  assign _2406_ = _2404_ | _2405_ /*28979*/;
  assign _2407_ = inv_6[23] ^ r_5[23] /*28977*/;
  assign sum_6[23] = _2407_ ^ _2406_ /*28976*/;
  assign _2408_ = _2407_ & _2406_ /*28975*/;
  assign _2409_ = inv_6[23] & r_5[23] /*28974*/;
  assign _2410_ = _2408_ | _2409_ /*28973*/;
  assign _2411_ = inv_6[24] ^ r_5[24] /*28971*/;
  assign sum_6[24] = _2411_ ^ _2410_ /*28970*/;
  assign _2412_ = _2411_ & _2410_ /*28969*/;
  assign _2413_ = inv_6[24] & r_5[24] /*28968*/;
  assign _2414_ = _2412_ | _2413_ /*28967*/;
  assign _2415_ = inv_6[25] ^ r_5[25] /*28965*/;
  assign sum_6[25] = _2415_ ^ _2414_ /*28964*/;
  assign _2416_ = _2415_ & _2414_ /*28963*/;
  assign _2417_ = inv_6[25] & r_5[25] /*28962*/;
  assign _2418_ = _2416_ | _2417_ /*28961*/;
  assign _2419_ = inv_6[26] ^ r_5[26] /*28959*/;
  assign sum_6[26] = _2419_ ^ _2418_ /*28958*/;
  assign _2420_ = _2419_ & _2418_ /*28957*/;
  assign _2421_ = inv_6[26] & r_5[26] /*28956*/;
  assign _2422_ = _2420_ | _2421_ /*28955*/;
  assign _2423_ = inv_6[27] ^ r_5[27] /*28953*/;
  assign sum_6[27] = _2423_ ^ _2422_ /*28952*/;
  assign _2424_ = _2423_ & _2422_ /*28951*/;
  assign _2425_ = inv_6[27] & r_5[27] /*28950*/;
  assign _2426_ = _2424_ | _2425_ /*28949*/;
  assign _2427_ = inv_6[28] ^ r_5[28] /*28947*/;
  assign sum_6[28] = _2427_ ^ _2426_ /*28946*/;
  assign _2428_ = _2427_ & _2426_ /*28945*/;
  assign _2429_ = inv_6[28] & r_5[28] /*28944*/;
  assign _2430_ = _2428_ | _2429_ /*28943*/;
  assign _2431_ = inv_6[29] ^ r_5[29] /*28941*/;
  assign sum_6[29] = _2431_ ^ _2430_ /*28940*/;
  assign _2432_ = _2431_ & _2430_ /*28939*/;
  assign _2433_ = inv_6[29] & r_5[29] /*28938*/;
  assign _2434_ = _2432_ | _2433_ /*28937*/;
  assign _2435_ = inv_6[30] ^ r_5[30] /*28935*/;
  assign sum_6[30] = _2435_ ^ _2434_ /*28934*/;
  assign _2436_ = _2435_ & _2434_ /*28933*/;
  assign _2437_ = inv_6[30] & r_5[30] /*28932*/;
  assign _2438_ = _2436_ | _2437_ /*28931*/;
  assign _2439_ = inv_6[31] ^ r_5[31] /*28929*/;
  assign sum_6[31] = _2439_ ^ _2438_ /*28928*/;
  assign _2440_ = _2439_ & _2438_ /*28927*/;
  assign _2441_ = inv_6[31] & r_5[31] /*28926*/;
  assign _2442_ = _2440_ | _2441_ /*28925*/;
  assign _2443_ = inv_6[32] ^ r_5[32] /*28923*/;
  assign sum_6[32] = _2443_ ^ _2442_ /*28922*/;
  assign _2444_ = _2443_ & _2442_ /*28921*/;
  assign _2445_ = inv_6[32] & r_5[32] /*28920*/;
  assign _2446_ = _2444_ | _2445_ /*28919*/;
  assign _2447_ = inv_6[33] ^ r_5[33] /*28917*/;
  assign sum_6[33] = _2447_ ^ _2446_ /*28916*/;
  assign _2448_ = _2447_ & _2446_ /*28915*/;
  assign _2449_ = inv_6[33] & r_5[33] /*28914*/;
  assign _2450_ = _2448_ | _2449_ /*28913*/;
  assign _2451_ = inv_6[34] ^ r_5[34] /*28911*/;
  assign sum_6[34] = _2451_ ^ _2450_ /*28910*/;
  assign _2452_ = _2451_ & _2450_ /*28909*/;
  assign _2453_ = inv_6[34] & r_5[34] /*28908*/;
  assign _2454_ = _2452_ | _2453_ /*28907*/;
  assign _2455_ = inv_6[35] ^ r_5[35] /*28905*/;
  assign sum_6[35] = _2455_ ^ _2454_ /*28904*/;
  assign _2456_ = _2455_ & _2454_ /*28903*/;
  assign _2457_ = inv_6[35] & r_5[35] /*28902*/;
  assign _2458_ = _2456_ | _2457_ /*28901*/;
  assign _2459_ = inv_6[36] ^ r_5[36] /*28899*/;
  assign sum_6[36] = _2459_ ^ _2458_ /*28898*/;
  assign _2460_ = _2459_ & _2458_ /*28897*/;
  assign _2461_ = inv_6[36] & r_5[36] /*28896*/;
  assign _2462_ = _2460_ | _2461_ /*28895*/;
  assign _2463_ = inv_6[37] ^ r_5[37] /*28893*/;
  assign sum_6[37] = _2463_ ^ _2462_ /*28892*/;
  assign _2464_ = _2463_ & _2462_ /*28891*/;
  assign _2465_ = inv_6[37] & r_5[37] /*28890*/;
  assign _2466_ = _2464_ | _2465_ /*28889*/;
  assign _2467_ = inv_6[38] ^ r_5[38] /*28887*/;
  assign sum_6[38] = _2467_ ^ _2466_ /*28886*/;
  assign _2468_ = _2467_ & _2466_ /*28885*/;
  assign _2469_ = inv_6[38] & r_5[38] /*28884*/;
  assign _2470_ = _2468_ | _2469_ /*28883*/;
  assign _2471_ = inv_6[39] ^ r_5[39] /*28881*/;
  assign sum_6[39] = _2471_ ^ _2470_ /*28880*/;
  assign _2472_ = _2471_ & _2470_ /*28879*/;
  assign _2473_ = inv_6[39] & r_5[39] /*28878*/;
  assign _2474_ = _2472_ | _2473_ /*28877*/;
  assign _2475_ = inv_6[40] ^ r_5[40] /*28875*/;
  assign sum_6[40] = _2475_ ^ _2474_ /*28874*/;
  assign _2476_ = _2475_ & _2474_ /*28873*/;
  assign _2477_ = inv_6[40] & r_5[40] /*28872*/;
  assign _2478_ = _2476_ | _2477_ /*28871*/;
  assign _2479_ = inv_6[41] ^ r_5[41] /*28869*/;
  assign sum_6[41] = _2479_ ^ _2478_ /*28868*/;
  assign _2480_ = _2479_ & _2478_ /*28867*/;
  assign _2481_ = inv_6[41] & r_5[41] /*28866*/;
  assign _2482_ = _2480_ | _2481_ /*28865*/;
  assign _2483_ = inv_6[42] ^ r_5[42] /*28863*/;
  assign sum_6[42] = _2483_ ^ _2482_ /*28862*/;
  assign _2484_ = _2483_ & _2482_ /*28861*/;
  assign _2485_ = inv_6[42] & r_5[42] /*28860*/;
  assign _2486_ = _2484_ | _2485_ /*28859*/;
  assign _2487_ = inv_6[43] ^ r_5[43] /*28857*/;
  assign sum_6[43] = _2487_ ^ _2486_ /*28856*/;
  assign _2488_ = _2487_ & _2486_ /*28855*/;
  assign _2489_ = inv_6[43] & r_5[43] /*28854*/;
  assign _2490_ = _2488_ | _2489_ /*28853*/;
  assign _2491_ = inv_6[44] ^ r_5[44] /*28851*/;
  assign sum_6[44] = _2491_ ^ _2490_ /*28850*/;
  assign _2492_ = _2491_ & _2490_ /*28849*/;
  assign _2493_ = inv_6[44] & r_5[44] /*28848*/;
  assign _2494_ = _2492_ | _2493_ /*28847*/;
  assign _2495_ = inv_6[45] ^ r_5[45] /*28845*/;
  assign sum_6[45] = _2495_ ^ _2494_ /*28844*/;
  assign _2496_ = _2495_ & _2494_ /*28843*/;
  assign _2497_ = inv_6[45] & r_5[45] /*28842*/;
  assign _2498_ = _2496_ | _2497_ /*28841*/;
  assign _2499_ = inv_6[46] ^ r_5[46] /*28839*/;
  assign sum_6[46] = _2499_ ^ _2498_ /*28838*/;
  assign _2500_ = _2499_ & _2498_ /*28837*/;
  assign _2501_ = inv_6[46] & r_5[46] /*28836*/;
  assign _2502_ = _2500_ | _2501_ /*28835*/;
  assign _2503_ = inv_6[47] ^ r_5[47] /*28833*/;
  assign sum_6[47] = _2503_ ^ _2502_ /*28832*/;
  assign _2504_ = _2503_ & _2502_ /*28831*/;
  assign _2505_ = inv_6[47] & r_5[47] /*28830*/;
  assign _2506_ = _2504_ | _2505_ /*28829*/;
  assign _2507_ = inv_6[48] ^ r_5[48] /*28827*/;
  assign sum_6[48] = _2507_ ^ _2506_ /*28826*/;
  assign _2508_ = _2507_ & _2506_ /*28825*/;
  assign _2509_ = inv_6[48] & r_5[48] /*28824*/;
  assign _2510_ = _2508_ | _2509_ /*28823*/;
  assign _2511_ = inv_6[49] ^ r_5[49] /*28821*/;
  assign sum_6[49] = _2511_ ^ _2510_ /*28820*/;
  assign _2512_ = _2511_ & _2510_ /*28819*/;
  assign _2513_ = inv_6[49] & r_5[49] /*28818*/;
  assign _2514_ = _2512_ | _2513_ /*28817*/;
  assign _2515_ = inv_6[50] ^ r_5[50] /*28815*/;
  assign sum_6[50] = _2515_ ^ _2514_ /*28814*/;
  assign _2516_ = _2515_ & _2514_ /*28813*/;
  assign _2517_ = inv_6[50] & r_5[50] /*28812*/;
  assign _2518_ = _2516_ | _2517_ /*28811*/;
  assign _2519_ = inv_6[51] ^ r_5[51] /*28809*/;
  assign sum_6[51] = _2519_ ^ _2518_ /*28808*/;
  assign _2520_ = _2519_ & _2518_ /*28807*/;
  assign _2521_ = inv_6[51] & r_5[51] /*28806*/;
  assign _2522_ = _2520_ | _2521_ /*28805*/;
  assign _2523_ = inv_6[52] ^ r_5[52] /*28803*/;
  assign sum_6[52] = _2523_ ^ _2522_ /*28802*/;
  assign _2524_ = _2523_ & _2522_ /*28801*/;
  assign _2525_ = inv_6[52] & r_5[52] /*28800*/;
  assign _2526_ = _2524_ | _2525_ /*28799*/;
  assign _2527_ = inv_6[53] ^ r_5[53] /*28797*/;
  assign sum_6[53] = _2527_ ^ _2526_ /*28796*/;
  assign _2528_ = _2527_ & _2526_ /*28795*/;
  assign _2529_ = inv_6[53] & r_5[53] /*28794*/;
  assign _2530_ = _2528_ | _2529_ /*28793*/;
  assign _2531_ = inv_6[54] ^ r_5[54] /*28791*/;
  assign sum_6[54] = _2531_ ^ _2530_ /*28790*/;
  assign _2532_ = _2531_ & _2530_ /*28789*/;
  assign _2533_ = inv_6[54] & r_5[54] /*28788*/;
  assign _2534_ = _2532_ | _2533_ /*28787*/;
  assign _2535_ = inv_6[55] ^ r_5[55] /*28785*/;
  assign sum_6[55] = _2535_ ^ _2534_ /*28784*/;
  assign _2536_ = _2535_ & _2534_ /*28783*/;
  assign _2537_ = inv_6[55] & r_5[55] /*28782*/;
  assign _2538_ = _2536_ | _2537_ /*28781*/;
  assign _2539_ = inv_6[56] ^ r_5[56] /*28779*/;
  assign sum_6[56] = _2539_ ^ _2538_ /*28778*/;
  assign _2540_ = _2539_ & _2538_ /*28777*/;
  assign _2541_ = inv_6[56] & r_5[56] /*28776*/;
  assign _2542_ = _2540_ | _2541_ /*28775*/;
  assign _2543_ = inv_6[57] ^ r_5[57] /*28773*/;
  assign sum_6[57] = _2543_ ^ _2542_ /*28772*/;
  assign _2544_ = _2543_ & _2542_ /*28771*/;
  assign _2545_ = inv_6[57] & r_5[57] /*28770*/;
  assign _2546_ = _2544_ | _2545_ /*28769*/;
  assign _2547_ = inv_6[58] ^ r_5[58] /*28767*/;
  assign sum_6[58] = _2547_ ^ _2546_ /*28766*/;
  assign _2548_ = _2547_ & _2546_ /*28765*/;
  assign _2549_ = inv_6[58] & r_5[58] /*28764*/;
  assign _2550_ = _2548_ | _2549_ /*28763*/;
  assign _2551_ = inv_6[59] ^ r_5[59] /*28761*/;
  assign sum_6[59] = _2551_ ^ _2550_ /*28760*/;
  assign _2552_ = _2551_ & _2550_ /*28759*/;
  assign _2553_ = inv_6[59] & r_5[59] /*28758*/;
  assign _2554_ = _2552_ | _2553_ /*28757*/;
  assign _2555_ = inv_6[60] ^ r_5[60] /*28755*/;
  assign sum_6[60] = _2555_ ^ _2554_ /*28754*/;
  assign _2556_ = _2555_ & _2554_ /*28753*/;
  assign _2557_ = inv_6[60] & r_5[60] /*28752*/;
  assign _2558_ = _2556_ | _2557_ /*28751*/;
  assign _2559_ = inv_6[61] ^ r_5[61] /*28749*/;
  assign sum_6[61] = _2559_ ^ _2558_ /*28748*/;
  assign _2560_ = _2559_ & _2558_ /*28747*/;
  assign _2561_ = inv_6[61] & r_5[61] /*28746*/;
  assign _2562_ = _2560_ | _2561_ /*28745*/;
  assign _2563_ = inv_6[62] ^ r_5[62] /*28743*/;
  assign sum_6[62] = _2563_ ^ _2562_ /*28742*/;
  assign _2564_ = _2563_ & _2562_ /*28741*/;
  assign _2565_ = inv_6[62] & r_5[62] /*28740*/;
  assign _2566_ = _2564_ | _2565_ /*28739*/;
  assign _2567_ = inv_6[63] ^ r_5[63] /*28737*/;
  assign sum_6[63] = _2567_ ^ _2566_ /*28736*/;
  assign _2568_ = _2567_ & _2566_ /*28735*/;
  assign _2569_ = inv_6[63] & r_5[63] /*28734*/;
  assign _2570_ = _2568_ | _2569_ /*28733*/;
  assign _2571_ = inv_6[64] ^ r_5[64] /*28731*/;
  assign sum_6[64] = _2571_ ^ _2570_ /*28730*/;
  assign _2572_ = _2571_ & _2570_ /*28729*/;
  assign _2573_ = inv_6[64] & r_5[64] /*28728*/;
  assign _2574_ = _2572_ | _2573_ /*28727*/;
  assign _2575_ = inv_6[65] ^ r_5[65] /*28725*/;
  assign sum_6[65] = _2575_ ^ _2574_ /*28724*/;
  assign _2576_ = _2575_ & _2574_ /*28723*/;
  assign _2577_ = inv_6[65] & r_5[65] /*28722*/;
  assign _2578_ = _2576_ | _2577_ /*28721*/;
  assign _2579_ = inv_6[66] ^ r_5[66] /*28719*/;
  assign sum_6[66] = _2579_ ^ _2578_ /*28718*/;
  assign _2580_ = _2579_ & _2578_ /*28717*/;
  assign _2581_ = inv_6[66] & r_5[66] /*28716*/;
  assign _2582_ = _2580_ | _2581_ /*28715*/;
  assign _2583_ = inv_6[67] ^ r_5[67] /*28713*/;
  assign sum_6[67] = _2583_ ^ _2582_ /*28712*/;
  assign _2584_ = _2583_ & _2582_ /*28711*/;
  assign _2585_ = inv_6[67] & r_5[67] /*28710*/;
  assign _2586_ = _2584_ | _2585_ /*28709*/;
  assign _2587_ = _2586_ ^ _2582_ /*28708*/;
  assign _2588_ = ~_2587_ /*28707*/;
  assign _2589_ = sum_6[67] & _2588_ /*28706*/;
  assign _2590_ = _2587_ & _2586_ /*28705*/;
  assign sum_6[68] = _2590_ | _2589_ /*28704*/;
  assign q[26] = ~sum_6[68] /*28703*/;
  assign m_6[0] = r_5[0] /*28702*/;
  assign m_6[1] = r_5[1] /*28701*/;
  assign m_6[2] = r_5[2] /*28700*/;
  assign m_6[3] = r_5[3] /*28699*/;
  assign m_6[4] = r_5[4] /*28698*/;
  assign m_6[5] = r_5[5] /*28697*/;
  assign m_6[6] = r_5[6] /*28696*/;
  assign m_6[7] = r_5[7] /*28695*/;
  assign m_6[8] = r_5[8] /*28694*/;
  assign m_6[9] = r_5[9] /*28693*/;
  assign m_6[10] = r_5[10] /*28692*/;
  assign m_6[11] = r_5[11] /*28691*/;
  assign m_6[12] = r_5[12] /*28690*/;
  assign m_6[13] = r_5[13] /*28689*/;
  assign m_6[14] = r_5[14] /*28688*/;
  assign m_6[15] = r_5[15] /*28687*/;
  assign m_6[16] = r_5[16] /*28686*/;
  assign m_6[17] = r_5[17] /*28685*/;
  assign m_6[18] = r_5[18] /*28684*/;
  assign m_6[19] = r_5[19] /*28683*/;
  assign m_6[20] = r_5[20] /*28682*/;
  assign m_6[21] = r_5[21] /*28681*/;
  assign m_6[22] = r_5[22] /*28680*/;
  assign m_6[23] = r_5[23] /*28679*/;
  assign m_6[24] = r_5[24] /*28678*/;
  assign m_6[25] = r_5[25] /*28677*/;
  assign m_6[26] = r_5[26] /*28676*/;
  assign m_6[27] = r_5[27] /*28675*/;
  assign m_6[28] = r_5[28] /*28674*/;
  assign m_6[29] = r_5[29] /*28673*/;
  assign m_6[30] = r_5[30] /*28672*/;
  assign m_6[31] = r_5[31] /*28671*/;
  assign m_6[32] = r_5[32] /*28670*/;
  assign m_6[33] = r_5[33] /*28669*/;
  assign m_6[34] = r_5[34] /*28668*/;
  assign m_6[35] = r_5[35] /*28667*/;
  assign m_6[36] = r_5[36] /*28666*/;
  assign m_6[37] = r_5[37] /*28665*/;
  assign m_6[38] = r_5[38] /*28664*/;
  assign m_6[39] = r_5[39] /*28663*/;
  assign m_6[40] = r_5[40] /*28662*/;
  assign m_6[41] = r_5[41] /*28661*/;
  assign m_6[42] = r_5[42] /*28660*/;
  assign m_6[43] = r_5[43] /*28659*/;
  assign m_6[44] = r_5[44] /*28658*/;
  assign m_6[45] = r_5[45] /*28657*/;
  assign m_6[46] = r_5[46] /*28656*/;
  assign m_6[47] = r_5[47] /*28655*/;
  assign m_6[48] = r_5[48] /*28654*/;
  assign m_6[49] = r_5[49] /*28653*/;
  assign m_6[50] = r_5[50] /*28652*/;
  assign m_6[51] = r_5[51] /*28651*/;
  assign m_6[52] = r_5[52] /*28650*/;
  assign m_6[53] = r_5[53] /*28649*/;
  assign m_6[54] = r_5[54] /*28648*/;
  assign m_6[55] = r_5[55] /*28647*/;
  assign m_6[56] = r_5[56] /*28646*/;
  assign m_6[57] = r_5[57] /*28645*/;
  assign m_6[58] = r_5[58] /*28644*/;
  assign m_6[59] = r_5[59] /*28643*/;
  assign m_6[60] = r_5[60] /*28642*/;
  assign m_6[61] = r_5[61] /*28641*/;
  assign m_6[62] = r_5[62] /*28640*/;
  assign m_6[63] = r_5[63] /*28639*/;
  assign m_6[64] = r_5[64] /*28638*/;
  assign m_6[65] = r_5[65] /*28637*/;
  assign m_6[66] = r_5[66] /*28636*/;
  assign m_6[67] = r_5[67] /*28635*/;
  assign m_6[68] = r_5[67] /*28634*/;
  assign _2592_ = ~q[26] /*28633*/;
  assign _2593_ = sum_6[0] & q[26] /*28632*/;
  assign _2594_ = m_6[0] & _2592_ /*28631*/;
  assign r_6[0] = _2594_ | _2593_ /*28630*/;
  assign _2595_ = ~q[26] /*28629*/;
  assign _2596_ = sum_6[1] & q[26] /*28628*/;
  assign _2597_ = m_6[1] & _2595_ /*28627*/;
  assign r_6[1] = _2597_ | _2596_ /*28626*/;
  assign _2598_ = ~q[26] /*28625*/;
  assign _2599_ = sum_6[2] & q[26] /*28624*/;
  assign _2600_ = m_6[2] & _2598_ /*28623*/;
  assign r_6[2] = _2600_ | _2599_ /*28622*/;
  assign _2601_ = ~q[26] /*28621*/;
  assign _2602_ = sum_6[3] & q[26] /*28620*/;
  assign _2603_ = m_6[3] & _2601_ /*28619*/;
  assign r_6[3] = _2603_ | _2602_ /*28618*/;
  assign _2604_ = ~q[26] /*28617*/;
  assign _2605_ = sum_6[4] & q[26] /*28616*/;
  assign _2606_ = m_6[4] & _2604_ /*28615*/;
  assign r_6[4] = _2606_ | _2605_ /*28614*/;
  assign _2607_ = ~q[26] /*28613*/;
  assign _2608_ = sum_6[5] & q[26] /*28612*/;
  assign _2609_ = m_6[5] & _2607_ /*28611*/;
  assign r_6[5] = _2609_ | _2608_ /*28610*/;
  assign _2610_ = ~q[26] /*28609*/;
  assign _2611_ = sum_6[6] & q[26] /*28608*/;
  assign _2612_ = m_6[6] & _2610_ /*28607*/;
  assign r_6[6] = _2612_ | _2611_ /*28606*/;
  assign _2613_ = ~q[26] /*28605*/;
  assign _2614_ = sum_6[7] & q[26] /*28604*/;
  assign _2615_ = m_6[7] & _2613_ /*28603*/;
  assign r_6[7] = _2615_ | _2614_ /*28602*/;
  assign _2616_ = ~q[26] /*28601*/;
  assign _2617_ = sum_6[8] & q[26] /*28600*/;
  assign _2618_ = m_6[8] & _2616_ /*28599*/;
  assign r_6[8] = _2618_ | _2617_ /*28598*/;
  assign _2619_ = ~q[26] /*28597*/;
  assign _2620_ = sum_6[9] & q[26] /*28596*/;
  assign _2621_ = m_6[9] & _2619_ /*28595*/;
  assign r_6[9] = _2621_ | _2620_ /*28594*/;
  assign _2622_ = ~q[26] /*28593*/;
  assign _2623_ = sum_6[10] & q[26] /*28592*/;
  assign _2624_ = m_6[10] & _2622_ /*28591*/;
  assign r_6[10] = _2624_ | _2623_ /*28590*/;
  assign _2625_ = ~q[26] /*28589*/;
  assign _2626_ = sum_6[11] & q[26] /*28588*/;
  assign _2627_ = m_6[11] & _2625_ /*28587*/;
  assign r_6[11] = _2627_ | _2626_ /*28586*/;
  assign _2628_ = ~q[26] /*28585*/;
  assign _2629_ = sum_6[12] & q[26] /*28584*/;
  assign _2630_ = m_6[12] & _2628_ /*28583*/;
  assign r_6[12] = _2630_ | _2629_ /*28582*/;
  assign _2631_ = ~q[26] /*28581*/;
  assign _2632_ = sum_6[13] & q[26] /*28580*/;
  assign _2633_ = m_6[13] & _2631_ /*28579*/;
  assign r_6[13] = _2633_ | _2632_ /*28578*/;
  assign _2634_ = ~q[26] /*28577*/;
  assign _2635_ = sum_6[14] & q[26] /*28576*/;
  assign _2636_ = m_6[14] & _2634_ /*28575*/;
  assign r_6[14] = _2636_ | _2635_ /*28574*/;
  assign _2637_ = ~q[26] /*28573*/;
  assign _2638_ = sum_6[15] & q[26] /*28572*/;
  assign _2639_ = m_6[15] & _2637_ /*28571*/;
  assign r_6[15] = _2639_ | _2638_ /*28570*/;
  assign _2640_ = ~q[26] /*28569*/;
  assign _2641_ = sum_6[16] & q[26] /*28568*/;
  assign _2642_ = m_6[16] & _2640_ /*28567*/;
  assign r_6[16] = _2642_ | _2641_ /*28566*/;
  assign _2643_ = ~q[26] /*28565*/;
  assign _2644_ = sum_6[17] & q[26] /*28564*/;
  assign _2645_ = m_6[17] & _2643_ /*28563*/;
  assign r_6[17] = _2645_ | _2644_ /*28562*/;
  assign _2646_ = ~q[26] /*28561*/;
  assign _2647_ = sum_6[18] & q[26] /*28560*/;
  assign _2648_ = m_6[18] & _2646_ /*28559*/;
  assign r_6[18] = _2648_ | _2647_ /*28558*/;
  assign _2649_ = ~q[26] /*28557*/;
  assign _2650_ = sum_6[19] & q[26] /*28556*/;
  assign _2651_ = m_6[19] & _2649_ /*28555*/;
  assign r_6[19] = _2651_ | _2650_ /*28554*/;
  assign _2652_ = ~q[26] /*28553*/;
  assign _2653_ = sum_6[20] & q[26] /*28552*/;
  assign _2654_ = m_6[20] & _2652_ /*28551*/;
  assign r_6[20] = _2654_ | _2653_ /*28550*/;
  assign _2655_ = ~q[26] /*28549*/;
  assign _2656_ = sum_6[21] & q[26] /*28548*/;
  assign _2657_ = m_6[21] & _2655_ /*28547*/;
  assign r_6[21] = _2657_ | _2656_ /*28546*/;
  assign _2658_ = ~q[26] /*28545*/;
  assign _2659_ = sum_6[22] & q[26] /*28544*/;
  assign _2660_ = m_6[22] & _2658_ /*28543*/;
  assign r_6[22] = _2660_ | _2659_ /*28542*/;
  assign _2661_ = ~q[26] /*28541*/;
  assign _2662_ = sum_6[23] & q[26] /*28540*/;
  assign _2663_ = m_6[23] & _2661_ /*28539*/;
  assign r_6[23] = _2663_ | _2662_ /*28538*/;
  assign _2664_ = ~q[26] /*28537*/;
  assign _2665_ = sum_6[24] & q[26] /*28536*/;
  assign _2666_ = m_6[24] & _2664_ /*28535*/;
  assign r_6[24] = _2666_ | _2665_ /*28534*/;
  assign _2667_ = ~q[26] /*28533*/;
  assign _2668_ = sum_6[25] & q[26] /*28532*/;
  assign _2669_ = m_6[25] & _2667_ /*28531*/;
  assign r_6[25] = _2669_ | _2668_ /*28530*/;
  assign _2670_ = ~q[26] /*28529*/;
  assign _2671_ = sum_6[26] & q[26] /*28528*/;
  assign _2672_ = m_6[26] & _2670_ /*28527*/;
  assign r_6[26] = _2672_ | _2671_ /*28526*/;
  assign _2673_ = ~q[26] /*28525*/;
  assign _2674_ = sum_6[27] & q[26] /*28524*/;
  assign _2675_ = m_6[27] & _2673_ /*28523*/;
  assign r_6[27] = _2675_ | _2674_ /*28522*/;
  assign _2676_ = ~q[26] /*28521*/;
  assign _2677_ = sum_6[28] & q[26] /*28520*/;
  assign _2678_ = m_6[28] & _2676_ /*28519*/;
  assign r_6[28] = _2678_ | _2677_ /*28518*/;
  assign _2679_ = ~q[26] /*28517*/;
  assign _2680_ = sum_6[29] & q[26] /*28516*/;
  assign _2681_ = m_6[29] & _2679_ /*28515*/;
  assign r_6[29] = _2681_ | _2680_ /*28514*/;
  assign _2682_ = ~q[26] /*28513*/;
  assign _2683_ = sum_6[30] & q[26] /*28512*/;
  assign _2684_ = m_6[30] & _2682_ /*28511*/;
  assign r_6[30] = _2684_ | _2683_ /*28510*/;
  assign _2685_ = ~q[26] /*28509*/;
  assign _2686_ = sum_6[31] & q[26] /*28508*/;
  assign _2687_ = m_6[31] & _2685_ /*28507*/;
  assign r_6[31] = _2687_ | _2686_ /*28506*/;
  assign _2688_ = ~q[26] /*28505*/;
  assign _2689_ = sum_6[32] & q[26] /*28504*/;
  assign _2690_ = m_6[32] & _2688_ /*28503*/;
  assign r_6[32] = _2690_ | _2689_ /*28502*/;
  assign _2691_ = ~q[26] /*28501*/;
  assign _2692_ = sum_6[33] & q[26] /*28500*/;
  assign _2693_ = m_6[33] & _2691_ /*28499*/;
  assign r_6[33] = _2693_ | _2692_ /*28498*/;
  assign _2694_ = ~q[26] /*28497*/;
  assign _2695_ = sum_6[34] & q[26] /*28496*/;
  assign _2696_ = m_6[34] & _2694_ /*28495*/;
  assign r_6[34] = _2696_ | _2695_ /*28494*/;
  assign _2697_ = ~q[26] /*28493*/;
  assign _2698_ = sum_6[35] & q[26] /*28492*/;
  assign _2699_ = m_6[35] & _2697_ /*28491*/;
  assign r_6[35] = _2699_ | _2698_ /*28490*/;
  assign _2700_ = ~q[26] /*28489*/;
  assign _2701_ = sum_6[36] & q[26] /*28488*/;
  assign _2702_ = m_6[36] & _2700_ /*28487*/;
  assign r_6[36] = _2702_ | _2701_ /*28486*/;
  assign _2703_ = ~q[26] /*28485*/;
  assign _2704_ = sum_6[37] & q[26] /*28484*/;
  assign _2705_ = m_6[37] & _2703_ /*28483*/;
  assign r_6[37] = _2705_ | _2704_ /*28482*/;
  assign _2706_ = ~q[26] /*28481*/;
  assign _2707_ = sum_6[38] & q[26] /*28480*/;
  assign _2708_ = m_6[38] & _2706_ /*28479*/;
  assign r_6[38] = _2708_ | _2707_ /*28478*/;
  assign _2709_ = ~q[26] /*28477*/;
  assign _2710_ = sum_6[39] & q[26] /*28476*/;
  assign _2711_ = m_6[39] & _2709_ /*28475*/;
  assign r_6[39] = _2711_ | _2710_ /*28474*/;
  assign _2712_ = ~q[26] /*28473*/;
  assign _2713_ = sum_6[40] & q[26] /*28472*/;
  assign _2714_ = m_6[40] & _2712_ /*28471*/;
  assign r_6[40] = _2714_ | _2713_ /*28470*/;
  assign _2715_ = ~q[26] /*28469*/;
  assign _2716_ = sum_6[41] & q[26] /*28468*/;
  assign _2717_ = m_6[41] & _2715_ /*28467*/;
  assign r_6[41] = _2717_ | _2716_ /*28466*/;
  assign _2718_ = ~q[26] /*28465*/;
  assign _2719_ = sum_6[42] & q[26] /*28464*/;
  assign _2720_ = m_6[42] & _2718_ /*28463*/;
  assign r_6[42] = _2720_ | _2719_ /*28462*/;
  assign _2721_ = ~q[26] /*28461*/;
  assign _2722_ = sum_6[43] & q[26] /*28460*/;
  assign _2723_ = m_6[43] & _2721_ /*28459*/;
  assign r_6[43] = _2723_ | _2722_ /*28458*/;
  assign _2724_ = ~q[26] /*28457*/;
  assign _2725_ = sum_6[44] & q[26] /*28456*/;
  assign _2726_ = m_6[44] & _2724_ /*28455*/;
  assign r_6[44] = _2726_ | _2725_ /*28454*/;
  assign _2727_ = ~q[26] /*28453*/;
  assign _2728_ = sum_6[45] & q[26] /*28452*/;
  assign _2729_ = m_6[45] & _2727_ /*28451*/;
  assign r_6[45] = _2729_ | _2728_ /*28450*/;
  assign _2730_ = ~q[26] /*28449*/;
  assign _2731_ = sum_6[46] & q[26] /*28448*/;
  assign _2732_ = m_6[46] & _2730_ /*28447*/;
  assign r_6[46] = _2732_ | _2731_ /*28446*/;
  assign _2733_ = ~q[26] /*28445*/;
  assign _2734_ = sum_6[47] & q[26] /*28444*/;
  assign _2735_ = m_6[47] & _2733_ /*28443*/;
  assign r_6[47] = _2735_ | _2734_ /*28442*/;
  assign _2736_ = ~q[26] /*28441*/;
  assign _2737_ = sum_6[48] & q[26] /*28440*/;
  assign _2738_ = m_6[48] & _2736_ /*28439*/;
  assign r_6[48] = _2738_ | _2737_ /*28438*/;
  assign _2739_ = ~q[26] /*28437*/;
  assign _2740_ = sum_6[49] & q[26] /*28436*/;
  assign _2741_ = m_6[49] & _2739_ /*28435*/;
  assign r_6[49] = _2741_ | _2740_ /*28434*/;
  assign _2742_ = ~q[26] /*28433*/;
  assign _2743_ = sum_6[50] & q[26] /*28432*/;
  assign _2744_ = m_6[50] & _2742_ /*28431*/;
  assign r_6[50] = _2744_ | _2743_ /*28430*/;
  assign _2745_ = ~q[26] /*28429*/;
  assign _2746_ = sum_6[51] & q[26] /*28428*/;
  assign _2747_ = m_6[51] & _2745_ /*28427*/;
  assign r_6[51] = _2747_ | _2746_ /*28426*/;
  assign _2748_ = ~q[26] /*28425*/;
  assign _2749_ = sum_6[52] & q[26] /*28424*/;
  assign _2750_ = m_6[52] & _2748_ /*28423*/;
  assign r_6[52] = _2750_ | _2749_ /*28422*/;
  assign _2751_ = ~q[26] /*28421*/;
  assign _2752_ = sum_6[53] & q[26] /*28420*/;
  assign _2753_ = m_6[53] & _2751_ /*28419*/;
  assign r_6[53] = _2753_ | _2752_ /*28418*/;
  assign _2754_ = ~q[26] /*28417*/;
  assign _2755_ = sum_6[54] & q[26] /*28416*/;
  assign _2756_ = m_6[54] & _2754_ /*28415*/;
  assign r_6[54] = _2756_ | _2755_ /*28414*/;
  assign _2757_ = ~q[26] /*28413*/;
  assign _2758_ = sum_6[55] & q[26] /*28412*/;
  assign _2759_ = m_6[55] & _2757_ /*28411*/;
  assign r_6[55] = _2759_ | _2758_ /*28410*/;
  assign _2760_ = ~q[26] /*28409*/;
  assign _2761_ = sum_6[56] & q[26] /*28408*/;
  assign _2762_ = m_6[56] & _2760_ /*28407*/;
  assign r_6[56] = _2762_ | _2761_ /*28406*/;
  assign _2763_ = ~q[26] /*28405*/;
  assign _2764_ = sum_6[57] & q[26] /*28404*/;
  assign _2765_ = m_6[57] & _2763_ /*28403*/;
  assign r_6[57] = _2765_ | _2764_ /*28402*/;
  assign _2766_ = ~q[26] /*28401*/;
  assign _2767_ = sum_6[58] & q[26] /*28400*/;
  assign _2768_ = m_6[58] & _2766_ /*28399*/;
  assign r_6[58] = _2768_ | _2767_ /*28398*/;
  assign _2769_ = ~q[26] /*28397*/;
  assign _2770_ = sum_6[59] & q[26] /*28396*/;
  assign _2771_ = m_6[59] & _2769_ /*28395*/;
  assign r_6[59] = _2771_ | _2770_ /*28394*/;
  assign _2772_ = ~q[26] /*28393*/;
  assign _2773_ = sum_6[60] & q[26] /*28392*/;
  assign _2774_ = m_6[60] & _2772_ /*28391*/;
  assign r_6[60] = _2774_ | _2773_ /*28390*/;
  assign _2775_ = ~q[26] /*28389*/;
  assign _2776_ = sum_6[61] & q[26] /*28388*/;
  assign _2777_ = m_6[61] & _2775_ /*28387*/;
  assign r_6[61] = _2777_ | _2776_ /*28386*/;
  assign _2778_ = ~q[26] /*28385*/;
  assign _2779_ = sum_6[62] & q[26] /*28384*/;
  assign _2780_ = m_6[62] & _2778_ /*28383*/;
  assign r_6[62] = _2780_ | _2779_ /*28382*/;
  assign _2781_ = ~q[26] /*28381*/;
  assign _2782_ = sum_6[63] & q[26] /*28380*/;
  assign _2783_ = m_6[63] & _2781_ /*28379*/;
  assign r_6[63] = _2783_ | _2782_ /*28378*/;
  assign _2784_ = ~q[26] /*28377*/;
  assign _2785_ = sum_6[64] & q[26] /*28376*/;
  assign _2786_ = m_6[64] & _2784_ /*28375*/;
  assign r_6[64] = _2786_ | _2785_ /*28374*/;
  assign _2787_ = ~q[26] /*28373*/;
  assign _2788_ = sum_6[65] & q[26] /*28372*/;
  assign _2789_ = m_6[65] & _2787_ /*28371*/;
  assign r_6[65] = _2789_ | _2788_ /*28370*/;
  assign _2790_ = ~q[26] /*28369*/;
  assign _2791_ = sum_6[66] & q[26] /*28368*/;
  assign _2792_ = m_6[66] & _2790_ /*28367*/;
  assign r_6[66] = _2792_ | _2791_ /*28366*/;
  assign _2793_ = ~q[26] /*28365*/;
  assign _2794_ = sum_6[67] & q[26] /*28364*/;
  assign _2795_ = m_6[67] & _2793_ /*28363*/;
  assign r_6[67] = _2795_ | _2794_ /*28362*/;
  assign _2796_ = ~q[26] /*28361*/;
  assign _2797_ = sum_6[68] & q[26] /*28360*/;
  assign _2798_ = m_6[68] & _2796_ /*28359*/;
  assign r_6[68] = _2798_ | _2797_ /*28358*/;
  assign inv_7[0] = oneWire /*28040*/;
  assign inv_7[1] = oneWire /*28034*/;
  assign inv_7[2] = oneWire /*28028*/;
  assign inv_7[3] = oneWire /*28022*/;
  assign inv_7[4] = oneWire /*28016*/;
  assign inv_7[5] = oneWire /*28010*/;
  assign inv_7[6] = oneWire /*28004*/;
  assign inv_7[7] = oneWire /*27998*/;
  assign inv_7[8] = oneWire /*27992*/;
  assign inv_7[9] = oneWire /*27986*/;
  assign inv_7[10] = oneWire /*27980*/;
  assign inv_7[11] = oneWire /*27974*/;
  assign inv_7[12] = oneWire /*27968*/;
  assign inv_7[13] = oneWire /*27962*/;
  assign inv_7[14] = oneWire /*27956*/;
  assign inv_7[15] = oneWire /*27950*/;
  assign inv_7[16] = oneWire /*27944*/;
  assign inv_7[17] = oneWire /*27938*/;
  assign inv_7[18] = oneWire /*27932*/;
  assign inv_7[19] = oneWire /*27926*/;
  assign inv_7[20] = oneWire /*27920*/;
  assign inv_7[21] = oneWire /*27914*/;
  assign inv_7[22] = oneWire /*27908*/;
  assign inv_7[23] = oneWire /*27902*/;
  assign inv_7[24] = oneWire /*27896*/;
  assign inv_7[25] = ~div[0] /*27890*/;
  assign inv_7[26] = ~div[1] /*27884*/;
  assign inv_7[27] = ~div[2] /*27878*/;
  assign inv_7[28] = ~div[3] /*27872*/;
  assign inv_7[29] = ~div[4] /*27866*/;
  assign inv_7[30] = ~div[5] /*27860*/;
  assign inv_7[31] = ~div[6] /*27854*/;
  assign inv_7[32] = ~div[7] /*27848*/;
  assign inv_7[33] = ~div[8] /*27842*/;
  assign inv_7[34] = ~div[9] /*27836*/;
  assign inv_7[35] = ~div[10] /*27830*/;
  assign inv_7[36] = ~div[11] /*27824*/;
  assign inv_7[37] = ~div[12] /*27818*/;
  assign inv_7[38] = ~div[13] /*27812*/;
  assign inv_7[39] = ~div[14] /*27806*/;
  assign inv_7[40] = ~div[15] /*27800*/;
  assign inv_7[41] = ~div[16] /*27794*/;
  assign inv_7[42] = ~div[17] /*27788*/;
  assign inv_7[43] = ~div[18] /*27782*/;
  assign inv_7[44] = ~div[19] /*27776*/;
  assign inv_7[45] = ~div[20] /*27770*/;
  assign inv_7[46] = ~div[21] /*27764*/;
  assign inv_7[47] = ~div[22] /*27758*/;
  assign inv_7[48] = ~div[23] /*27752*/;
  assign inv_7[49] = ~div[24] /*27746*/;
  assign inv_7[50] = ~div[25] /*27740*/;
  assign inv_7[51] = ~div[26] /*27734*/;
  assign inv_7[52] = ~div[27] /*27728*/;
  assign inv_7[53] = ~div[28] /*27722*/;
  assign inv_7[54] = ~div[29] /*27716*/;
  assign inv_7[55] = ~div[30] /*27710*/;
  assign inv_7[56] = oneWire /*27704*/;
  assign inv_7[57] = oneWire /*27698*/;
  assign inv_7[58] = oneWire /*27692*/;
  assign inv_7[59] = oneWire /*27686*/;
  assign inv_7[60] = oneWire /*27680*/;
  assign inv_7[61] = oneWire /*27674*/;
  assign inv_7[62] = oneWire /*27668*/;
  assign inv_7[63] = oneWire /*27662*/;
  assign inv_7[64] = oneWire /*27656*/;
  assign inv_7[65] = oneWire /*27650*/;
  assign inv_7[66] = oneWire /*27644*/;
  assign inv_7[67] = oneWire /*27638*/;
  assign inv_7[68] = oneWire /*27632*/;
  assign _2799_ = inv_7[0] ^ r_6[0] /*28039*/;
  assign sum_7[0] = _2799_ ^ oneWire /*28038*/;
  assign _2800_ = _2799_ & oneWire /*28037*/;
  assign _2801_ = inv_7[0] & r_6[0] /*28036*/;
  assign _2802_ = _2800_ | _2801_ /*28035*/;
  assign _2803_ = inv_7[1] ^ r_6[1] /*28033*/;
  assign sum_7[1] = _2803_ ^ _2802_ /*28032*/;
  assign _2804_ = _2803_ & _2802_ /*28031*/;
  assign _2805_ = inv_7[1] & r_6[1] /*28030*/;
  assign _2806_ = _2804_ | _2805_ /*28029*/;
  assign _2807_ = inv_7[2] ^ r_6[2] /*28027*/;
  assign sum_7[2] = _2807_ ^ _2806_ /*28026*/;
  assign _2808_ = _2807_ & _2806_ /*28025*/;
  assign _2809_ = inv_7[2] & r_6[2] /*28024*/;
  assign _2810_ = _2808_ | _2809_ /*28023*/;
  assign _2811_ = inv_7[3] ^ r_6[3] /*28021*/;
  assign sum_7[3] = _2811_ ^ _2810_ /*28020*/;
  assign _2812_ = _2811_ & _2810_ /*28019*/;
  assign _2813_ = inv_7[3] & r_6[3] /*28018*/;
  assign _2814_ = _2812_ | _2813_ /*28017*/;
  assign _2815_ = inv_7[4] ^ r_6[4] /*28015*/;
  assign sum_7[4] = _2815_ ^ _2814_ /*28014*/;
  assign _2816_ = _2815_ & _2814_ /*28013*/;
  assign _2817_ = inv_7[4] & r_6[4] /*28012*/;
  assign _2818_ = _2816_ | _2817_ /*28011*/;
  assign _2819_ = inv_7[5] ^ r_6[5] /*28009*/;
  assign sum_7[5] = _2819_ ^ _2818_ /*28008*/;
  assign _2820_ = _2819_ & _2818_ /*28007*/;
  assign _2821_ = inv_7[5] & r_6[5] /*28006*/;
  assign _2822_ = _2820_ | _2821_ /*28005*/;
  assign _2823_ = inv_7[6] ^ r_6[6] /*28003*/;
  assign sum_7[6] = _2823_ ^ _2822_ /*28002*/;
  assign _2824_ = _2823_ & _2822_ /*28001*/;
  assign _2825_ = inv_7[6] & r_6[6] /*28000*/;
  assign _2826_ = _2824_ | _2825_ /*27999*/;
  assign _2827_ = inv_7[7] ^ r_6[7] /*27997*/;
  assign sum_7[7] = _2827_ ^ _2826_ /*27996*/;
  assign _2828_ = _2827_ & _2826_ /*27995*/;
  assign _2829_ = inv_7[7] & r_6[7] /*27994*/;
  assign _2830_ = _2828_ | _2829_ /*27993*/;
  assign _2831_ = inv_7[8] ^ r_6[8] /*27991*/;
  assign sum_7[8] = _2831_ ^ _2830_ /*27990*/;
  assign _2832_ = _2831_ & _2830_ /*27989*/;
  assign _2833_ = inv_7[8] & r_6[8] /*27988*/;
  assign _2834_ = _2832_ | _2833_ /*27987*/;
  assign _2835_ = inv_7[9] ^ r_6[9] /*27985*/;
  assign sum_7[9] = _2835_ ^ _2834_ /*27984*/;
  assign _2836_ = _2835_ & _2834_ /*27983*/;
  assign _2837_ = inv_7[9] & r_6[9] /*27982*/;
  assign _2838_ = _2836_ | _2837_ /*27981*/;
  assign _2839_ = inv_7[10] ^ r_6[10] /*27979*/;
  assign sum_7[10] = _2839_ ^ _2838_ /*27978*/;
  assign _2840_ = _2839_ & _2838_ /*27977*/;
  assign _2841_ = inv_7[10] & r_6[10] /*27976*/;
  assign _2842_ = _2840_ | _2841_ /*27975*/;
  assign _2843_ = inv_7[11] ^ r_6[11] /*27973*/;
  assign sum_7[11] = _2843_ ^ _2842_ /*27972*/;
  assign _2844_ = _2843_ & _2842_ /*27971*/;
  assign _2845_ = inv_7[11] & r_6[11] /*27970*/;
  assign _2846_ = _2844_ | _2845_ /*27969*/;
  assign _2847_ = inv_7[12] ^ r_6[12] /*27967*/;
  assign sum_7[12] = _2847_ ^ _2846_ /*27966*/;
  assign _2848_ = _2847_ & _2846_ /*27965*/;
  assign _2849_ = inv_7[12] & r_6[12] /*27964*/;
  assign _2850_ = _2848_ | _2849_ /*27963*/;
  assign _2851_ = inv_7[13] ^ r_6[13] /*27961*/;
  assign sum_7[13] = _2851_ ^ _2850_ /*27960*/;
  assign _2852_ = _2851_ & _2850_ /*27959*/;
  assign _2853_ = inv_7[13] & r_6[13] /*27958*/;
  assign _2854_ = _2852_ | _2853_ /*27957*/;
  assign _2855_ = inv_7[14] ^ r_6[14] /*27955*/;
  assign sum_7[14] = _2855_ ^ _2854_ /*27954*/;
  assign _2856_ = _2855_ & _2854_ /*27953*/;
  assign _2857_ = inv_7[14] & r_6[14] /*27952*/;
  assign _2858_ = _2856_ | _2857_ /*27951*/;
  assign _2859_ = inv_7[15] ^ r_6[15] /*27949*/;
  assign sum_7[15] = _2859_ ^ _2858_ /*27948*/;
  assign _2860_ = _2859_ & _2858_ /*27947*/;
  assign _2861_ = inv_7[15] & r_6[15] /*27946*/;
  assign _2862_ = _2860_ | _2861_ /*27945*/;
  assign _2863_ = inv_7[16] ^ r_6[16] /*27943*/;
  assign sum_7[16] = _2863_ ^ _2862_ /*27942*/;
  assign _2864_ = _2863_ & _2862_ /*27941*/;
  assign _2865_ = inv_7[16] & r_6[16] /*27940*/;
  assign _2866_ = _2864_ | _2865_ /*27939*/;
  assign _2867_ = inv_7[17] ^ r_6[17] /*27937*/;
  assign sum_7[17] = _2867_ ^ _2866_ /*27936*/;
  assign _2868_ = _2867_ & _2866_ /*27935*/;
  assign _2869_ = inv_7[17] & r_6[17] /*27934*/;
  assign _2870_ = _2868_ | _2869_ /*27933*/;
  assign _2871_ = inv_7[18] ^ r_6[18] /*27931*/;
  assign sum_7[18] = _2871_ ^ _2870_ /*27930*/;
  assign _2872_ = _2871_ & _2870_ /*27929*/;
  assign _2873_ = inv_7[18] & r_6[18] /*27928*/;
  assign _2874_ = _2872_ | _2873_ /*27927*/;
  assign _2875_ = inv_7[19] ^ r_6[19] /*27925*/;
  assign sum_7[19] = _2875_ ^ _2874_ /*27924*/;
  assign _2876_ = _2875_ & _2874_ /*27923*/;
  assign _2877_ = inv_7[19] & r_6[19] /*27922*/;
  assign _2878_ = _2876_ | _2877_ /*27921*/;
  assign _2879_ = inv_7[20] ^ r_6[20] /*27919*/;
  assign sum_7[20] = _2879_ ^ _2878_ /*27918*/;
  assign _2880_ = _2879_ & _2878_ /*27917*/;
  assign _2881_ = inv_7[20] & r_6[20] /*27916*/;
  assign _2882_ = _2880_ | _2881_ /*27915*/;
  assign _2883_ = inv_7[21] ^ r_6[21] /*27913*/;
  assign sum_7[21] = _2883_ ^ _2882_ /*27912*/;
  assign _2884_ = _2883_ & _2882_ /*27911*/;
  assign _2885_ = inv_7[21] & r_6[21] /*27910*/;
  assign _2886_ = _2884_ | _2885_ /*27909*/;
  assign _2887_ = inv_7[22] ^ r_6[22] /*27907*/;
  assign sum_7[22] = _2887_ ^ _2886_ /*27906*/;
  assign _2888_ = _2887_ & _2886_ /*27905*/;
  assign _2889_ = inv_7[22] & r_6[22] /*27904*/;
  assign _2890_ = _2888_ | _2889_ /*27903*/;
  assign _2891_ = inv_7[23] ^ r_6[23] /*27901*/;
  assign sum_7[23] = _2891_ ^ _2890_ /*27900*/;
  assign _2892_ = _2891_ & _2890_ /*27899*/;
  assign _2893_ = inv_7[23] & r_6[23] /*27898*/;
  assign _2894_ = _2892_ | _2893_ /*27897*/;
  assign _2895_ = inv_7[24] ^ r_6[24] /*27895*/;
  assign sum_7[24] = _2895_ ^ _2894_ /*27894*/;
  assign _2896_ = _2895_ & _2894_ /*27893*/;
  assign _2897_ = inv_7[24] & r_6[24] /*27892*/;
  assign _2898_ = _2896_ | _2897_ /*27891*/;
  assign _2899_ = inv_7[25] ^ r_6[25] /*27889*/;
  assign sum_7[25] = _2899_ ^ _2898_ /*27888*/;
  assign _2900_ = _2899_ & _2898_ /*27887*/;
  assign _2901_ = inv_7[25] & r_6[25] /*27886*/;
  assign _2902_ = _2900_ | _2901_ /*27885*/;
  assign _2903_ = inv_7[26] ^ r_6[26] /*27883*/;
  assign sum_7[26] = _2903_ ^ _2902_ /*27882*/;
  assign _2904_ = _2903_ & _2902_ /*27881*/;
  assign _2905_ = inv_7[26] & r_6[26] /*27880*/;
  assign _2906_ = _2904_ | _2905_ /*27879*/;
  assign _2907_ = inv_7[27] ^ r_6[27] /*27877*/;
  assign sum_7[27] = _2907_ ^ _2906_ /*27876*/;
  assign _2908_ = _2907_ & _2906_ /*27875*/;
  assign _2909_ = inv_7[27] & r_6[27] /*27874*/;
  assign _2910_ = _2908_ | _2909_ /*27873*/;
  assign _2911_ = inv_7[28] ^ r_6[28] /*27871*/;
  assign sum_7[28] = _2911_ ^ _2910_ /*27870*/;
  assign _2912_ = _2911_ & _2910_ /*27869*/;
  assign _2913_ = inv_7[28] & r_6[28] /*27868*/;
  assign _2914_ = _2912_ | _2913_ /*27867*/;
  assign _2915_ = inv_7[29] ^ r_6[29] /*27865*/;
  assign sum_7[29] = _2915_ ^ _2914_ /*27864*/;
  assign _2916_ = _2915_ & _2914_ /*27863*/;
  assign _2917_ = inv_7[29] & r_6[29] /*27862*/;
  assign _2918_ = _2916_ | _2917_ /*27861*/;
  assign _2919_ = inv_7[30] ^ r_6[30] /*27859*/;
  assign sum_7[30] = _2919_ ^ _2918_ /*27858*/;
  assign _2920_ = _2919_ & _2918_ /*27857*/;
  assign _2921_ = inv_7[30] & r_6[30] /*27856*/;
  assign _2922_ = _2920_ | _2921_ /*27855*/;
  assign _2923_ = inv_7[31] ^ r_6[31] /*27853*/;
  assign sum_7[31] = _2923_ ^ _2922_ /*27852*/;
  assign _2924_ = _2923_ & _2922_ /*27851*/;
  assign _2925_ = inv_7[31] & r_6[31] /*27850*/;
  assign _2926_ = _2924_ | _2925_ /*27849*/;
  assign _2927_ = inv_7[32] ^ r_6[32] /*27847*/;
  assign sum_7[32] = _2927_ ^ _2926_ /*27846*/;
  assign _2928_ = _2927_ & _2926_ /*27845*/;
  assign _2929_ = inv_7[32] & r_6[32] /*27844*/;
  assign _2930_ = _2928_ | _2929_ /*27843*/;
  assign _2931_ = inv_7[33] ^ r_6[33] /*27841*/;
  assign sum_7[33] = _2931_ ^ _2930_ /*27840*/;
  assign _2932_ = _2931_ & _2930_ /*27839*/;
  assign _2933_ = inv_7[33] & r_6[33] /*27838*/;
  assign _2934_ = _2932_ | _2933_ /*27837*/;
  assign _2935_ = inv_7[34] ^ r_6[34] /*27835*/;
  assign sum_7[34] = _2935_ ^ _2934_ /*27834*/;
  assign _2936_ = _2935_ & _2934_ /*27833*/;
  assign _2937_ = inv_7[34] & r_6[34] /*27832*/;
  assign _2938_ = _2936_ | _2937_ /*27831*/;
  assign _2939_ = inv_7[35] ^ r_6[35] /*27829*/;
  assign sum_7[35] = _2939_ ^ _2938_ /*27828*/;
  assign _2940_ = _2939_ & _2938_ /*27827*/;
  assign _2941_ = inv_7[35] & r_6[35] /*27826*/;
  assign _2942_ = _2940_ | _2941_ /*27825*/;
  assign _2943_ = inv_7[36] ^ r_6[36] /*27823*/;
  assign sum_7[36] = _2943_ ^ _2942_ /*27822*/;
  assign _2944_ = _2943_ & _2942_ /*27821*/;
  assign _2945_ = inv_7[36] & r_6[36] /*27820*/;
  assign _2946_ = _2944_ | _2945_ /*27819*/;
  assign _2947_ = inv_7[37] ^ r_6[37] /*27817*/;
  assign sum_7[37] = _2947_ ^ _2946_ /*27816*/;
  assign _2948_ = _2947_ & _2946_ /*27815*/;
  assign _2949_ = inv_7[37] & r_6[37] /*27814*/;
  assign _2950_ = _2948_ | _2949_ /*27813*/;
  assign _2951_ = inv_7[38] ^ r_6[38] /*27811*/;
  assign sum_7[38] = _2951_ ^ _2950_ /*27810*/;
  assign _2952_ = _2951_ & _2950_ /*27809*/;
  assign _2953_ = inv_7[38] & r_6[38] /*27808*/;
  assign _2954_ = _2952_ | _2953_ /*27807*/;
  assign _2955_ = inv_7[39] ^ r_6[39] /*27805*/;
  assign sum_7[39] = _2955_ ^ _2954_ /*27804*/;
  assign _2956_ = _2955_ & _2954_ /*27803*/;
  assign _2957_ = inv_7[39] & r_6[39] /*27802*/;
  assign _2958_ = _2956_ | _2957_ /*27801*/;
  assign _2959_ = inv_7[40] ^ r_6[40] /*27799*/;
  assign sum_7[40] = _2959_ ^ _2958_ /*27798*/;
  assign _2960_ = _2959_ & _2958_ /*27797*/;
  assign _2961_ = inv_7[40] & r_6[40] /*27796*/;
  assign _2962_ = _2960_ | _2961_ /*27795*/;
  assign _2963_ = inv_7[41] ^ r_6[41] /*27793*/;
  assign sum_7[41] = _2963_ ^ _2962_ /*27792*/;
  assign _2964_ = _2963_ & _2962_ /*27791*/;
  assign _2965_ = inv_7[41] & r_6[41] /*27790*/;
  assign _2966_ = _2964_ | _2965_ /*27789*/;
  assign _2967_ = inv_7[42] ^ r_6[42] /*27787*/;
  assign sum_7[42] = _2967_ ^ _2966_ /*27786*/;
  assign _2968_ = _2967_ & _2966_ /*27785*/;
  assign _2969_ = inv_7[42] & r_6[42] /*27784*/;
  assign _2970_ = _2968_ | _2969_ /*27783*/;
  assign _2971_ = inv_7[43] ^ r_6[43] /*27781*/;
  assign sum_7[43] = _2971_ ^ _2970_ /*27780*/;
  assign _2972_ = _2971_ & _2970_ /*27779*/;
  assign _2973_ = inv_7[43] & r_6[43] /*27778*/;
  assign _2974_ = _2972_ | _2973_ /*27777*/;
  assign _2975_ = inv_7[44] ^ r_6[44] /*27775*/;
  assign sum_7[44] = _2975_ ^ _2974_ /*27774*/;
  assign _2976_ = _2975_ & _2974_ /*27773*/;
  assign _2977_ = inv_7[44] & r_6[44] /*27772*/;
  assign _2978_ = _2976_ | _2977_ /*27771*/;
  assign _2979_ = inv_7[45] ^ r_6[45] /*27769*/;
  assign sum_7[45] = _2979_ ^ _2978_ /*27768*/;
  assign _2980_ = _2979_ & _2978_ /*27767*/;
  assign _2981_ = inv_7[45] & r_6[45] /*27766*/;
  assign _2982_ = _2980_ | _2981_ /*27765*/;
  assign _2983_ = inv_7[46] ^ r_6[46] /*27763*/;
  assign sum_7[46] = _2983_ ^ _2982_ /*27762*/;
  assign _2984_ = _2983_ & _2982_ /*27761*/;
  assign _2985_ = inv_7[46] & r_6[46] /*27760*/;
  assign _2986_ = _2984_ | _2985_ /*27759*/;
  assign _2987_ = inv_7[47] ^ r_6[47] /*27757*/;
  assign sum_7[47] = _2987_ ^ _2986_ /*27756*/;
  assign _2988_ = _2987_ & _2986_ /*27755*/;
  assign _2989_ = inv_7[47] & r_6[47] /*27754*/;
  assign _2990_ = _2988_ | _2989_ /*27753*/;
  assign _2991_ = inv_7[48] ^ r_6[48] /*27751*/;
  assign sum_7[48] = _2991_ ^ _2990_ /*27750*/;
  assign _2992_ = _2991_ & _2990_ /*27749*/;
  assign _2993_ = inv_7[48] & r_6[48] /*27748*/;
  assign _2994_ = _2992_ | _2993_ /*27747*/;
  assign _2995_ = inv_7[49] ^ r_6[49] /*27745*/;
  assign sum_7[49] = _2995_ ^ _2994_ /*27744*/;
  assign _2996_ = _2995_ & _2994_ /*27743*/;
  assign _2997_ = inv_7[49] & r_6[49] /*27742*/;
  assign _2998_ = _2996_ | _2997_ /*27741*/;
  assign _2999_ = inv_7[50] ^ r_6[50] /*27739*/;
  assign sum_7[50] = _2999_ ^ _2998_ /*27738*/;
  assign _3000_ = _2999_ & _2998_ /*27737*/;
  assign _3001_ = inv_7[50] & r_6[50] /*27736*/;
  assign _3002_ = _3000_ | _3001_ /*27735*/;
  assign _3003_ = inv_7[51] ^ r_6[51] /*27733*/;
  assign sum_7[51] = _3003_ ^ _3002_ /*27732*/;
  assign _3004_ = _3003_ & _3002_ /*27731*/;
  assign _3005_ = inv_7[51] & r_6[51] /*27730*/;
  assign _3006_ = _3004_ | _3005_ /*27729*/;
  assign _3007_ = inv_7[52] ^ r_6[52] /*27727*/;
  assign sum_7[52] = _3007_ ^ _3006_ /*27726*/;
  assign _3008_ = _3007_ & _3006_ /*27725*/;
  assign _3009_ = inv_7[52] & r_6[52] /*27724*/;
  assign _3010_ = _3008_ | _3009_ /*27723*/;
  assign _3011_ = inv_7[53] ^ r_6[53] /*27721*/;
  assign sum_7[53] = _3011_ ^ _3010_ /*27720*/;
  assign _3012_ = _3011_ & _3010_ /*27719*/;
  assign _3013_ = inv_7[53] & r_6[53] /*27718*/;
  assign _3014_ = _3012_ | _3013_ /*27717*/;
  assign _3015_ = inv_7[54] ^ r_6[54] /*27715*/;
  assign sum_7[54] = _3015_ ^ _3014_ /*27714*/;
  assign _3016_ = _3015_ & _3014_ /*27713*/;
  assign _3017_ = inv_7[54] & r_6[54] /*27712*/;
  assign _3018_ = _3016_ | _3017_ /*27711*/;
  assign _3019_ = inv_7[55] ^ r_6[55] /*27709*/;
  assign sum_7[55] = _3019_ ^ _3018_ /*27708*/;
  assign _3020_ = _3019_ & _3018_ /*27707*/;
  assign _3021_ = inv_7[55] & r_6[55] /*27706*/;
  assign _3022_ = _3020_ | _3021_ /*27705*/;
  assign _3023_ = inv_7[56] ^ r_6[56] /*27703*/;
  assign sum_7[56] = _3023_ ^ _3022_ /*27702*/;
  assign _3024_ = _3023_ & _3022_ /*27701*/;
  assign _3025_ = inv_7[56] & r_6[56] /*27700*/;
  assign _3026_ = _3024_ | _3025_ /*27699*/;
  assign _3027_ = inv_7[57] ^ r_6[57] /*27697*/;
  assign sum_7[57] = _3027_ ^ _3026_ /*27696*/;
  assign _3028_ = _3027_ & _3026_ /*27695*/;
  assign _3029_ = inv_7[57] & r_6[57] /*27694*/;
  assign _3030_ = _3028_ | _3029_ /*27693*/;
  assign _3031_ = inv_7[58] ^ r_6[58] /*27691*/;
  assign sum_7[58] = _3031_ ^ _3030_ /*27690*/;
  assign _3032_ = _3031_ & _3030_ /*27689*/;
  assign _3033_ = inv_7[58] & r_6[58] /*27688*/;
  assign _3034_ = _3032_ | _3033_ /*27687*/;
  assign _3035_ = inv_7[59] ^ r_6[59] /*27685*/;
  assign sum_7[59] = _3035_ ^ _3034_ /*27684*/;
  assign _3036_ = _3035_ & _3034_ /*27683*/;
  assign _3037_ = inv_7[59] & r_6[59] /*27682*/;
  assign _3038_ = _3036_ | _3037_ /*27681*/;
  assign _3039_ = inv_7[60] ^ r_6[60] /*27679*/;
  assign sum_7[60] = _3039_ ^ _3038_ /*27678*/;
  assign _3040_ = _3039_ & _3038_ /*27677*/;
  assign _3041_ = inv_7[60] & r_6[60] /*27676*/;
  assign _3042_ = _3040_ | _3041_ /*27675*/;
  assign _3043_ = inv_7[61] ^ r_6[61] /*27673*/;
  assign sum_7[61] = _3043_ ^ _3042_ /*27672*/;
  assign _3044_ = _3043_ & _3042_ /*27671*/;
  assign _3045_ = inv_7[61] & r_6[61] /*27670*/;
  assign _3046_ = _3044_ | _3045_ /*27669*/;
  assign _3047_ = inv_7[62] ^ r_6[62] /*27667*/;
  assign sum_7[62] = _3047_ ^ _3046_ /*27666*/;
  assign _3048_ = _3047_ & _3046_ /*27665*/;
  assign _3049_ = inv_7[62] & r_6[62] /*27664*/;
  assign _3050_ = _3048_ | _3049_ /*27663*/;
  assign _3051_ = inv_7[63] ^ r_6[63] /*27661*/;
  assign sum_7[63] = _3051_ ^ _3050_ /*27660*/;
  assign _3052_ = _3051_ & _3050_ /*27659*/;
  assign _3053_ = inv_7[63] & r_6[63] /*27658*/;
  assign _3054_ = _3052_ | _3053_ /*27657*/;
  assign _3055_ = inv_7[64] ^ r_6[64] /*27655*/;
  assign sum_7[64] = _3055_ ^ _3054_ /*27654*/;
  assign _3056_ = _3055_ & _3054_ /*27653*/;
  assign _3057_ = inv_7[64] & r_6[64] /*27652*/;
  assign _3058_ = _3056_ | _3057_ /*27651*/;
  assign _3059_ = inv_7[65] ^ r_6[65] /*27649*/;
  assign sum_7[65] = _3059_ ^ _3058_ /*27648*/;
  assign _3060_ = _3059_ & _3058_ /*27647*/;
  assign _3061_ = inv_7[65] & r_6[65] /*27646*/;
  assign _3062_ = _3060_ | _3061_ /*27645*/;
  assign _3063_ = inv_7[66] ^ r_6[66] /*27643*/;
  assign sum_7[66] = _3063_ ^ _3062_ /*27642*/;
  assign _3064_ = _3063_ & _3062_ /*27641*/;
  assign _3065_ = inv_7[66] & r_6[66] /*27640*/;
  assign _3066_ = _3064_ | _3065_ /*27639*/;
  assign _3067_ = inv_7[67] ^ r_6[67] /*27637*/;
  assign sum_7[67] = _3067_ ^ _3066_ /*27636*/;
  assign _3068_ = _3067_ & _3066_ /*27635*/;
  assign _3069_ = inv_7[67] & r_6[67] /*27634*/;
  assign _3070_ = _3068_ | _3069_ /*27633*/;
  assign _3071_ = inv_7[68] ^ r_6[68] /*27631*/;
  assign sum_7[68] = _3071_ ^ _3070_ /*27630*/;
  assign _3072_ = _3071_ & _3070_ /*27629*/;
  assign _3073_ = inv_7[68] & r_6[68] /*27628*/;
  assign _3074_ = _3072_ | _3073_ /*27627*/;
  assign _3075_ = _3074_ ^ _3070_ /*27626*/;
  assign _3076_ = ~_3075_ /*27625*/;
  assign _3077_ = sum_7[68] & _3076_ /*27624*/;
  assign _3078_ = _3075_ & _3074_ /*27623*/;
  assign sum_7[69] = _3078_ | _3077_ /*27622*/;
  assign q[25] = ~sum_7[69] /*27621*/;
  assign m_7[0] = r_6[0] /*27620*/;
  assign m_7[1] = r_6[1] /*27619*/;
  assign m_7[2] = r_6[2] /*27618*/;
  assign m_7[3] = r_6[3] /*27617*/;
  assign m_7[4] = r_6[4] /*27616*/;
  assign m_7[5] = r_6[5] /*27615*/;
  assign m_7[6] = r_6[6] /*27614*/;
  assign m_7[7] = r_6[7] /*27613*/;
  assign m_7[8] = r_6[8] /*27612*/;
  assign m_7[9] = r_6[9] /*27611*/;
  assign m_7[10] = r_6[10] /*27610*/;
  assign m_7[11] = r_6[11] /*27609*/;
  assign m_7[12] = r_6[12] /*27608*/;
  assign m_7[13] = r_6[13] /*27607*/;
  assign m_7[14] = r_6[14] /*27606*/;
  assign m_7[15] = r_6[15] /*27605*/;
  assign m_7[16] = r_6[16] /*27604*/;
  assign m_7[17] = r_6[17] /*27603*/;
  assign m_7[18] = r_6[18] /*27602*/;
  assign m_7[19] = r_6[19] /*27601*/;
  assign m_7[20] = r_6[20] /*27600*/;
  assign m_7[21] = r_6[21] /*27599*/;
  assign m_7[22] = r_6[22] /*27598*/;
  assign m_7[23] = r_6[23] /*27597*/;
  assign m_7[24] = r_6[24] /*27596*/;
  assign m_7[25] = r_6[25] /*27595*/;
  assign m_7[26] = r_6[26] /*27594*/;
  assign m_7[27] = r_6[27] /*27593*/;
  assign m_7[28] = r_6[28] /*27592*/;
  assign m_7[29] = r_6[29] /*27591*/;
  assign m_7[30] = r_6[30] /*27590*/;
  assign m_7[31] = r_6[31] /*27589*/;
  assign m_7[32] = r_6[32] /*27588*/;
  assign m_7[33] = r_6[33] /*27587*/;
  assign m_7[34] = r_6[34] /*27586*/;
  assign m_7[35] = r_6[35] /*27585*/;
  assign m_7[36] = r_6[36] /*27584*/;
  assign m_7[37] = r_6[37] /*27583*/;
  assign m_7[38] = r_6[38] /*27582*/;
  assign m_7[39] = r_6[39] /*27581*/;
  assign m_7[40] = r_6[40] /*27580*/;
  assign m_7[41] = r_6[41] /*27579*/;
  assign m_7[42] = r_6[42] /*27578*/;
  assign m_7[43] = r_6[43] /*27577*/;
  assign m_7[44] = r_6[44] /*27576*/;
  assign m_7[45] = r_6[45] /*27575*/;
  assign m_7[46] = r_6[46] /*27574*/;
  assign m_7[47] = r_6[47] /*27573*/;
  assign m_7[48] = r_6[48] /*27572*/;
  assign m_7[49] = r_6[49] /*27571*/;
  assign m_7[50] = r_6[50] /*27570*/;
  assign m_7[51] = r_6[51] /*27569*/;
  assign m_7[52] = r_6[52] /*27568*/;
  assign m_7[53] = r_6[53] /*27567*/;
  assign m_7[54] = r_6[54] /*27566*/;
  assign m_7[55] = r_6[55] /*27565*/;
  assign m_7[56] = r_6[56] /*27564*/;
  assign m_7[57] = r_6[57] /*27563*/;
  assign m_7[58] = r_6[58] /*27562*/;
  assign m_7[59] = r_6[59] /*27561*/;
  assign m_7[60] = r_6[60] /*27560*/;
  assign m_7[61] = r_6[61] /*27559*/;
  assign m_7[62] = r_6[62] /*27558*/;
  assign m_7[63] = r_6[63] /*27557*/;
  assign m_7[64] = r_6[64] /*27556*/;
  assign m_7[65] = r_6[65] /*27555*/;
  assign m_7[66] = r_6[66] /*27554*/;
  assign m_7[67] = r_6[67] /*27553*/;
  assign m_7[68] = r_6[68] /*27552*/;
  assign m_7[69] = r_6[68] /*27551*/;
  assign _3080_ = ~q[25] /*27550*/;
  assign _3081_ = sum_7[0] & q[25] /*27549*/;
  assign _3082_ = m_7[0] & _3080_ /*27548*/;
  assign r_7[0] = _3082_ | _3081_ /*27547*/;
  assign _3083_ = ~q[25] /*27546*/;
  assign _3084_ = sum_7[1] & q[25] /*27545*/;
  assign _3085_ = m_7[1] & _3083_ /*27544*/;
  assign r_7[1] = _3085_ | _3084_ /*27543*/;
  assign _3086_ = ~q[25] /*27542*/;
  assign _3087_ = sum_7[2] & q[25] /*27541*/;
  assign _3088_ = m_7[2] & _3086_ /*27540*/;
  assign r_7[2] = _3088_ | _3087_ /*27539*/;
  assign _3089_ = ~q[25] /*27538*/;
  assign _3090_ = sum_7[3] & q[25] /*27537*/;
  assign _3091_ = m_7[3] & _3089_ /*27536*/;
  assign r_7[3] = _3091_ | _3090_ /*27535*/;
  assign _3092_ = ~q[25] /*27534*/;
  assign _3093_ = sum_7[4] & q[25] /*27533*/;
  assign _3094_ = m_7[4] & _3092_ /*27532*/;
  assign r_7[4] = _3094_ | _3093_ /*27531*/;
  assign _3095_ = ~q[25] /*27530*/;
  assign _3096_ = sum_7[5] & q[25] /*27529*/;
  assign _3097_ = m_7[5] & _3095_ /*27528*/;
  assign r_7[5] = _3097_ | _3096_ /*27527*/;
  assign _3098_ = ~q[25] /*27526*/;
  assign _3099_ = sum_7[6] & q[25] /*27525*/;
  assign _3100_ = m_7[6] & _3098_ /*27524*/;
  assign r_7[6] = _3100_ | _3099_ /*27523*/;
  assign _3101_ = ~q[25] /*27522*/;
  assign _3102_ = sum_7[7] & q[25] /*27521*/;
  assign _3103_ = m_7[7] & _3101_ /*27520*/;
  assign r_7[7] = _3103_ | _3102_ /*27519*/;
  assign _3104_ = ~q[25] /*27518*/;
  assign _3105_ = sum_7[8] & q[25] /*27517*/;
  assign _3106_ = m_7[8] & _3104_ /*27516*/;
  assign r_7[8] = _3106_ | _3105_ /*27515*/;
  assign _3107_ = ~q[25] /*27514*/;
  assign _3108_ = sum_7[9] & q[25] /*27513*/;
  assign _3109_ = m_7[9] & _3107_ /*27512*/;
  assign r_7[9] = _3109_ | _3108_ /*27511*/;
  assign _3110_ = ~q[25] /*27510*/;
  assign _3111_ = sum_7[10] & q[25] /*27509*/;
  assign _3112_ = m_7[10] & _3110_ /*27508*/;
  assign r_7[10] = _3112_ | _3111_ /*27507*/;
  assign _3113_ = ~q[25] /*27506*/;
  assign _3114_ = sum_7[11] & q[25] /*27505*/;
  assign _3115_ = m_7[11] & _3113_ /*27504*/;
  assign r_7[11] = _3115_ | _3114_ /*27503*/;
  assign _3116_ = ~q[25] /*27502*/;
  assign _3117_ = sum_7[12] & q[25] /*27501*/;
  assign _3118_ = m_7[12] & _3116_ /*27500*/;
  assign r_7[12] = _3118_ | _3117_ /*27499*/;
  assign _3119_ = ~q[25] /*27498*/;
  assign _3120_ = sum_7[13] & q[25] /*27497*/;
  assign _3121_ = m_7[13] & _3119_ /*27496*/;
  assign r_7[13] = _3121_ | _3120_ /*27495*/;
  assign _3122_ = ~q[25] /*27494*/;
  assign _3123_ = sum_7[14] & q[25] /*27493*/;
  assign _3124_ = m_7[14] & _3122_ /*27492*/;
  assign r_7[14] = _3124_ | _3123_ /*27491*/;
  assign _3125_ = ~q[25] /*27490*/;
  assign _3126_ = sum_7[15] & q[25] /*27489*/;
  assign _3127_ = m_7[15] & _3125_ /*27488*/;
  assign r_7[15] = _3127_ | _3126_ /*27487*/;
  assign _3128_ = ~q[25] /*27486*/;
  assign _3129_ = sum_7[16] & q[25] /*27485*/;
  assign _3130_ = m_7[16] & _3128_ /*27484*/;
  assign r_7[16] = _3130_ | _3129_ /*27483*/;
  assign _3131_ = ~q[25] /*27482*/;
  assign _3132_ = sum_7[17] & q[25] /*27481*/;
  assign _3133_ = m_7[17] & _3131_ /*27480*/;
  assign r_7[17] = _3133_ | _3132_ /*27479*/;
  assign _3134_ = ~q[25] /*27478*/;
  assign _3135_ = sum_7[18] & q[25] /*27477*/;
  assign _3136_ = m_7[18] & _3134_ /*27476*/;
  assign r_7[18] = _3136_ | _3135_ /*27475*/;
  assign _3137_ = ~q[25] /*27474*/;
  assign _3138_ = sum_7[19] & q[25] /*27473*/;
  assign _3139_ = m_7[19] & _3137_ /*27472*/;
  assign r_7[19] = _3139_ | _3138_ /*27471*/;
  assign _3140_ = ~q[25] /*27470*/;
  assign _3141_ = sum_7[20] & q[25] /*27469*/;
  assign _3142_ = m_7[20] & _3140_ /*27468*/;
  assign r_7[20] = _3142_ | _3141_ /*27467*/;
  assign _3143_ = ~q[25] /*27466*/;
  assign _3144_ = sum_7[21] & q[25] /*27465*/;
  assign _3145_ = m_7[21] & _3143_ /*27464*/;
  assign r_7[21] = _3145_ | _3144_ /*27463*/;
  assign _3146_ = ~q[25] /*27462*/;
  assign _3147_ = sum_7[22] & q[25] /*27461*/;
  assign _3148_ = m_7[22] & _3146_ /*27460*/;
  assign r_7[22] = _3148_ | _3147_ /*27459*/;
  assign _3149_ = ~q[25] /*27458*/;
  assign _3150_ = sum_7[23] & q[25] /*27457*/;
  assign _3151_ = m_7[23] & _3149_ /*27456*/;
  assign r_7[23] = _3151_ | _3150_ /*27455*/;
  assign _3152_ = ~q[25] /*27454*/;
  assign _3153_ = sum_7[24] & q[25] /*27453*/;
  assign _3154_ = m_7[24] & _3152_ /*27452*/;
  assign r_7[24] = _3154_ | _3153_ /*27451*/;
  assign _3155_ = ~q[25] /*27450*/;
  assign _3156_ = sum_7[25] & q[25] /*27449*/;
  assign _3157_ = m_7[25] & _3155_ /*27448*/;
  assign r_7[25] = _3157_ | _3156_ /*27447*/;
  assign _3158_ = ~q[25] /*27446*/;
  assign _3159_ = sum_7[26] & q[25] /*27445*/;
  assign _3160_ = m_7[26] & _3158_ /*27444*/;
  assign r_7[26] = _3160_ | _3159_ /*27443*/;
  assign _3161_ = ~q[25] /*27442*/;
  assign _3162_ = sum_7[27] & q[25] /*27441*/;
  assign _3163_ = m_7[27] & _3161_ /*27440*/;
  assign r_7[27] = _3163_ | _3162_ /*27439*/;
  assign _3164_ = ~q[25] /*27438*/;
  assign _3165_ = sum_7[28] & q[25] /*27437*/;
  assign _3166_ = m_7[28] & _3164_ /*27436*/;
  assign r_7[28] = _3166_ | _3165_ /*27435*/;
  assign _3167_ = ~q[25] /*27434*/;
  assign _3168_ = sum_7[29] & q[25] /*27433*/;
  assign _3169_ = m_7[29] & _3167_ /*27432*/;
  assign r_7[29] = _3169_ | _3168_ /*27431*/;
  assign _3170_ = ~q[25] /*27430*/;
  assign _3171_ = sum_7[30] & q[25] /*27429*/;
  assign _3172_ = m_7[30] & _3170_ /*27428*/;
  assign r_7[30] = _3172_ | _3171_ /*27427*/;
  assign _3173_ = ~q[25] /*27426*/;
  assign _3174_ = sum_7[31] & q[25] /*27425*/;
  assign _3175_ = m_7[31] & _3173_ /*27424*/;
  assign r_7[31] = _3175_ | _3174_ /*27423*/;
  assign _3176_ = ~q[25] /*27422*/;
  assign _3177_ = sum_7[32] & q[25] /*27421*/;
  assign _3178_ = m_7[32] & _3176_ /*27420*/;
  assign r_7[32] = _3178_ | _3177_ /*27419*/;
  assign _3179_ = ~q[25] /*27418*/;
  assign _3180_ = sum_7[33] & q[25] /*27417*/;
  assign _3181_ = m_7[33] & _3179_ /*27416*/;
  assign r_7[33] = _3181_ | _3180_ /*27415*/;
  assign _3182_ = ~q[25] /*27414*/;
  assign _3183_ = sum_7[34] & q[25] /*27413*/;
  assign _3184_ = m_7[34] & _3182_ /*27412*/;
  assign r_7[34] = _3184_ | _3183_ /*27411*/;
  assign _3185_ = ~q[25] /*27410*/;
  assign _3186_ = sum_7[35] & q[25] /*27409*/;
  assign _3187_ = m_7[35] & _3185_ /*27408*/;
  assign r_7[35] = _3187_ | _3186_ /*27407*/;
  assign _3188_ = ~q[25] /*27406*/;
  assign _3189_ = sum_7[36] & q[25] /*27405*/;
  assign _3190_ = m_7[36] & _3188_ /*27404*/;
  assign r_7[36] = _3190_ | _3189_ /*27403*/;
  assign _3191_ = ~q[25] /*27402*/;
  assign _3192_ = sum_7[37] & q[25] /*27401*/;
  assign _3193_ = m_7[37] & _3191_ /*27400*/;
  assign r_7[37] = _3193_ | _3192_ /*27399*/;
  assign _3194_ = ~q[25] /*27398*/;
  assign _3195_ = sum_7[38] & q[25] /*27397*/;
  assign _3196_ = m_7[38] & _3194_ /*27396*/;
  assign r_7[38] = _3196_ | _3195_ /*27395*/;
  assign _3197_ = ~q[25] /*27394*/;
  assign _3198_ = sum_7[39] & q[25] /*27393*/;
  assign _3199_ = m_7[39] & _3197_ /*27392*/;
  assign r_7[39] = _3199_ | _3198_ /*27391*/;
  assign _3200_ = ~q[25] /*27390*/;
  assign _3201_ = sum_7[40] & q[25] /*27389*/;
  assign _3202_ = m_7[40] & _3200_ /*27388*/;
  assign r_7[40] = _3202_ | _3201_ /*27387*/;
  assign _3203_ = ~q[25] /*27386*/;
  assign _3204_ = sum_7[41] & q[25] /*27385*/;
  assign _3205_ = m_7[41] & _3203_ /*27384*/;
  assign r_7[41] = _3205_ | _3204_ /*27383*/;
  assign _3206_ = ~q[25] /*27382*/;
  assign _3207_ = sum_7[42] & q[25] /*27381*/;
  assign _3208_ = m_7[42] & _3206_ /*27380*/;
  assign r_7[42] = _3208_ | _3207_ /*27379*/;
  assign _3209_ = ~q[25] /*27378*/;
  assign _3210_ = sum_7[43] & q[25] /*27377*/;
  assign _3211_ = m_7[43] & _3209_ /*27376*/;
  assign r_7[43] = _3211_ | _3210_ /*27375*/;
  assign _3212_ = ~q[25] /*27374*/;
  assign _3213_ = sum_7[44] & q[25] /*27373*/;
  assign _3214_ = m_7[44] & _3212_ /*27372*/;
  assign r_7[44] = _3214_ | _3213_ /*27371*/;
  assign _3215_ = ~q[25] /*27370*/;
  assign _3216_ = sum_7[45] & q[25] /*27369*/;
  assign _3217_ = m_7[45] & _3215_ /*27368*/;
  assign r_7[45] = _3217_ | _3216_ /*27367*/;
  assign _3218_ = ~q[25] /*27366*/;
  assign _3219_ = sum_7[46] & q[25] /*27365*/;
  assign _3220_ = m_7[46] & _3218_ /*27364*/;
  assign r_7[46] = _3220_ | _3219_ /*27363*/;
  assign _3221_ = ~q[25] /*27362*/;
  assign _3222_ = sum_7[47] & q[25] /*27361*/;
  assign _3223_ = m_7[47] & _3221_ /*27360*/;
  assign r_7[47] = _3223_ | _3222_ /*27359*/;
  assign _3224_ = ~q[25] /*27358*/;
  assign _3225_ = sum_7[48] & q[25] /*27357*/;
  assign _3226_ = m_7[48] & _3224_ /*27356*/;
  assign r_7[48] = _3226_ | _3225_ /*27355*/;
  assign _3227_ = ~q[25] /*27354*/;
  assign _3228_ = sum_7[49] & q[25] /*27353*/;
  assign _3229_ = m_7[49] & _3227_ /*27352*/;
  assign r_7[49] = _3229_ | _3228_ /*27351*/;
  assign _3230_ = ~q[25] /*27350*/;
  assign _3231_ = sum_7[50] & q[25] /*27349*/;
  assign _3232_ = m_7[50] & _3230_ /*27348*/;
  assign r_7[50] = _3232_ | _3231_ /*27347*/;
  assign _3233_ = ~q[25] /*27346*/;
  assign _3234_ = sum_7[51] & q[25] /*27345*/;
  assign _3235_ = m_7[51] & _3233_ /*27344*/;
  assign r_7[51] = _3235_ | _3234_ /*27343*/;
  assign _3236_ = ~q[25] /*27342*/;
  assign _3237_ = sum_7[52] & q[25] /*27341*/;
  assign _3238_ = m_7[52] & _3236_ /*27340*/;
  assign r_7[52] = _3238_ | _3237_ /*27339*/;
  assign _3239_ = ~q[25] /*27338*/;
  assign _3240_ = sum_7[53] & q[25] /*27337*/;
  assign _3241_ = m_7[53] & _3239_ /*27336*/;
  assign r_7[53] = _3241_ | _3240_ /*27335*/;
  assign _3242_ = ~q[25] /*27334*/;
  assign _3243_ = sum_7[54] & q[25] /*27333*/;
  assign _3244_ = m_7[54] & _3242_ /*27332*/;
  assign r_7[54] = _3244_ | _3243_ /*27331*/;
  assign _3245_ = ~q[25] /*27330*/;
  assign _3246_ = sum_7[55] & q[25] /*27329*/;
  assign _3247_ = m_7[55] & _3245_ /*27328*/;
  assign r_7[55] = _3247_ | _3246_ /*27327*/;
  assign _3248_ = ~q[25] /*27326*/;
  assign _3249_ = sum_7[56] & q[25] /*27325*/;
  assign _3250_ = m_7[56] & _3248_ /*27324*/;
  assign r_7[56] = _3250_ | _3249_ /*27323*/;
  assign _3251_ = ~q[25] /*27322*/;
  assign _3252_ = sum_7[57] & q[25] /*27321*/;
  assign _3253_ = m_7[57] & _3251_ /*27320*/;
  assign r_7[57] = _3253_ | _3252_ /*27319*/;
  assign _3254_ = ~q[25] /*27318*/;
  assign _3255_ = sum_7[58] & q[25] /*27317*/;
  assign _3256_ = m_7[58] & _3254_ /*27316*/;
  assign r_7[58] = _3256_ | _3255_ /*27315*/;
  assign _3257_ = ~q[25] /*27314*/;
  assign _3258_ = sum_7[59] & q[25] /*27313*/;
  assign _3259_ = m_7[59] & _3257_ /*27312*/;
  assign r_7[59] = _3259_ | _3258_ /*27311*/;
  assign _3260_ = ~q[25] /*27310*/;
  assign _3261_ = sum_7[60] & q[25] /*27309*/;
  assign _3262_ = m_7[60] & _3260_ /*27308*/;
  assign r_7[60] = _3262_ | _3261_ /*27307*/;
  assign _3263_ = ~q[25] /*27306*/;
  assign _3264_ = sum_7[61] & q[25] /*27305*/;
  assign _3265_ = m_7[61] & _3263_ /*27304*/;
  assign r_7[61] = _3265_ | _3264_ /*27303*/;
  assign _3266_ = ~q[25] /*27302*/;
  assign _3267_ = sum_7[62] & q[25] /*27301*/;
  assign _3268_ = m_7[62] & _3266_ /*27300*/;
  assign r_7[62] = _3268_ | _3267_ /*27299*/;
  assign _3269_ = ~q[25] /*27298*/;
  assign _3270_ = sum_7[63] & q[25] /*27297*/;
  assign _3271_ = m_7[63] & _3269_ /*27296*/;
  assign r_7[63] = _3271_ | _3270_ /*27295*/;
  assign _3272_ = ~q[25] /*27294*/;
  assign _3273_ = sum_7[64] & q[25] /*27293*/;
  assign _3274_ = m_7[64] & _3272_ /*27292*/;
  assign r_7[64] = _3274_ | _3273_ /*27291*/;
  assign _3275_ = ~q[25] /*27290*/;
  assign _3276_ = sum_7[65] & q[25] /*27289*/;
  assign _3277_ = m_7[65] & _3275_ /*27288*/;
  assign r_7[65] = _3277_ | _3276_ /*27287*/;
  assign _3278_ = ~q[25] /*27286*/;
  assign _3279_ = sum_7[66] & q[25] /*27285*/;
  assign _3280_ = m_7[66] & _3278_ /*27284*/;
  assign r_7[66] = _3280_ | _3279_ /*27283*/;
  assign _3281_ = ~q[25] /*27282*/;
  assign _3282_ = sum_7[67] & q[25] /*27281*/;
  assign _3283_ = m_7[67] & _3281_ /*27280*/;
  assign r_7[67] = _3283_ | _3282_ /*27279*/;
  assign _3284_ = ~q[25] /*27278*/;
  assign _3285_ = sum_7[68] & q[25] /*27277*/;
  assign _3286_ = m_7[68] & _3284_ /*27276*/;
  assign r_7[68] = _3286_ | _3285_ /*27275*/;
  assign _3287_ = ~q[25] /*27274*/;
  assign _3288_ = sum_7[69] & q[25] /*27273*/;
  assign _3289_ = m_7[69] & _3287_ /*27272*/;
  assign r_7[69] = _3289_ | _3288_ /*27271*/;
  assign inv_8[0] = oneWire /*26964*/;
  assign inv_8[1] = oneWire /*26958*/;
  assign inv_8[2] = oneWire /*26952*/;
  assign inv_8[3] = oneWire /*26946*/;
  assign inv_8[4] = oneWire /*26940*/;
  assign inv_8[5] = oneWire /*26934*/;
  assign inv_8[6] = oneWire /*26928*/;
  assign inv_8[7] = oneWire /*26922*/;
  assign inv_8[8] = oneWire /*26916*/;
  assign inv_8[9] = oneWire /*26910*/;
  assign inv_8[10] = oneWire /*26904*/;
  assign inv_8[11] = oneWire /*26898*/;
  assign inv_8[12] = oneWire /*26892*/;
  assign inv_8[13] = oneWire /*26886*/;
  assign inv_8[14] = oneWire /*26880*/;
  assign inv_8[15] = oneWire /*26874*/;
  assign inv_8[16] = oneWire /*26868*/;
  assign inv_8[17] = oneWire /*26862*/;
  assign inv_8[18] = oneWire /*26856*/;
  assign inv_8[19] = oneWire /*26850*/;
  assign inv_8[20] = oneWire /*26844*/;
  assign inv_8[21] = oneWire /*26838*/;
  assign inv_8[22] = oneWire /*26832*/;
  assign inv_8[23] = oneWire /*26826*/;
  assign inv_8[24] = ~div[0] /*26820*/;
  assign inv_8[25] = ~div[1] /*26814*/;
  assign inv_8[26] = ~div[2] /*26808*/;
  assign inv_8[27] = ~div[3] /*26802*/;
  assign inv_8[28] = ~div[4] /*26796*/;
  assign inv_8[29] = ~div[5] /*26790*/;
  assign inv_8[30] = ~div[6] /*26784*/;
  assign inv_8[31] = ~div[7] /*26778*/;
  assign inv_8[32] = ~div[8] /*26772*/;
  assign inv_8[33] = ~div[9] /*26766*/;
  assign inv_8[34] = ~div[10] /*26760*/;
  assign inv_8[35] = ~div[11] /*26754*/;
  assign inv_8[36] = ~div[12] /*26748*/;
  assign inv_8[37] = ~div[13] /*26742*/;
  assign inv_8[38] = ~div[14] /*26736*/;
  assign inv_8[39] = ~div[15] /*26730*/;
  assign inv_8[40] = ~div[16] /*26724*/;
  assign inv_8[41] = ~div[17] /*26718*/;
  assign inv_8[42] = ~div[18] /*26712*/;
  assign inv_8[43] = ~div[19] /*26706*/;
  assign inv_8[44] = ~div[20] /*26700*/;
  assign inv_8[45] = ~div[21] /*26694*/;
  assign inv_8[46] = ~div[22] /*26688*/;
  assign inv_8[47] = ~div[23] /*26682*/;
  assign inv_8[48] = ~div[24] /*26676*/;
  assign inv_8[49] = ~div[25] /*26670*/;
  assign inv_8[50] = ~div[26] /*26664*/;
  assign inv_8[51] = ~div[27] /*26658*/;
  assign inv_8[52] = ~div[28] /*26652*/;
  assign inv_8[53] = ~div[29] /*26646*/;
  assign inv_8[54] = ~div[30] /*26640*/;
  assign inv_8[55] = oneWire /*26634*/;
  assign inv_8[56] = oneWire /*26628*/;
  assign inv_8[57] = oneWire /*26622*/;
  assign inv_8[58] = oneWire /*26616*/;
  assign inv_8[59] = oneWire /*26610*/;
  assign inv_8[60] = oneWire /*26604*/;
  assign inv_8[61] = oneWire /*26598*/;
  assign inv_8[62] = oneWire /*26592*/;
  assign inv_8[63] = oneWire /*26586*/;
  assign inv_8[64] = oneWire /*26580*/;
  assign inv_8[65] = oneWire /*26574*/;
  assign inv_8[66] = oneWire /*26568*/;
  assign inv_8[67] = oneWire /*26562*/;
  assign inv_8[68] = oneWire /*26556*/;
  assign inv_8[69] = oneWire /*26550*/;
  assign _3290_ = inv_8[0] ^ r_7[0] /*26963*/;
  assign sum_8[0] = _3290_ ^ oneWire /*26962*/;
  assign _3291_ = _3290_ & oneWire /*26961*/;
  assign _3292_ = inv_8[0] & r_7[0] /*26960*/;
  assign _3293_ = _3291_ | _3292_ /*26959*/;
  assign _3294_ = inv_8[1] ^ r_7[1] /*26957*/;
  assign sum_8[1] = _3294_ ^ _3293_ /*26956*/;
  assign _3295_ = _3294_ & _3293_ /*26955*/;
  assign _3296_ = inv_8[1] & r_7[1] /*26954*/;
  assign _3297_ = _3295_ | _3296_ /*26953*/;
  assign _3298_ = inv_8[2] ^ r_7[2] /*26951*/;
  assign sum_8[2] = _3298_ ^ _3297_ /*26950*/;
  assign _3299_ = _3298_ & _3297_ /*26949*/;
  assign _3300_ = inv_8[2] & r_7[2] /*26948*/;
  assign _3301_ = _3299_ | _3300_ /*26947*/;
  assign _3302_ = inv_8[3] ^ r_7[3] /*26945*/;
  assign sum_8[3] = _3302_ ^ _3301_ /*26944*/;
  assign _3303_ = _3302_ & _3301_ /*26943*/;
  assign _3304_ = inv_8[3] & r_7[3] /*26942*/;
  assign _3305_ = _3303_ | _3304_ /*26941*/;
  assign _3306_ = inv_8[4] ^ r_7[4] /*26939*/;
  assign sum_8[4] = _3306_ ^ _3305_ /*26938*/;
  assign _3307_ = _3306_ & _3305_ /*26937*/;
  assign _3308_ = inv_8[4] & r_7[4] /*26936*/;
  assign _3309_ = _3307_ | _3308_ /*26935*/;
  assign _3310_ = inv_8[5] ^ r_7[5] /*26933*/;
  assign sum_8[5] = _3310_ ^ _3309_ /*26932*/;
  assign _3311_ = _3310_ & _3309_ /*26931*/;
  assign _3312_ = inv_8[5] & r_7[5] /*26930*/;
  assign _3313_ = _3311_ | _3312_ /*26929*/;
  assign _3314_ = inv_8[6] ^ r_7[6] /*26927*/;
  assign sum_8[6] = _3314_ ^ _3313_ /*26926*/;
  assign _3315_ = _3314_ & _3313_ /*26925*/;
  assign _3316_ = inv_8[6] & r_7[6] /*26924*/;
  assign _3317_ = _3315_ | _3316_ /*26923*/;
  assign _3318_ = inv_8[7] ^ r_7[7] /*26921*/;
  assign sum_8[7] = _3318_ ^ _3317_ /*26920*/;
  assign _3319_ = _3318_ & _3317_ /*26919*/;
  assign _3320_ = inv_8[7] & r_7[7] /*26918*/;
  assign _3321_ = _3319_ | _3320_ /*26917*/;
  assign _3322_ = inv_8[8] ^ r_7[8] /*26915*/;
  assign sum_8[8] = _3322_ ^ _3321_ /*26914*/;
  assign _3323_ = _3322_ & _3321_ /*26913*/;
  assign _3324_ = inv_8[8] & r_7[8] /*26912*/;
  assign _3325_ = _3323_ | _3324_ /*26911*/;
  assign _3326_ = inv_8[9] ^ r_7[9] /*26909*/;
  assign sum_8[9] = _3326_ ^ _3325_ /*26908*/;
  assign _3327_ = _3326_ & _3325_ /*26907*/;
  assign _3328_ = inv_8[9] & r_7[9] /*26906*/;
  assign _3329_ = _3327_ | _3328_ /*26905*/;
  assign _3330_ = inv_8[10] ^ r_7[10] /*26903*/;
  assign sum_8[10] = _3330_ ^ _3329_ /*26902*/;
  assign _3331_ = _3330_ & _3329_ /*26901*/;
  assign _3332_ = inv_8[10] & r_7[10] /*26900*/;
  assign _3333_ = _3331_ | _3332_ /*26899*/;
  assign _3334_ = inv_8[11] ^ r_7[11] /*26897*/;
  assign sum_8[11] = _3334_ ^ _3333_ /*26896*/;
  assign _3335_ = _3334_ & _3333_ /*26895*/;
  assign _3336_ = inv_8[11] & r_7[11] /*26894*/;
  assign _3337_ = _3335_ | _3336_ /*26893*/;
  assign _3338_ = inv_8[12] ^ r_7[12] /*26891*/;
  assign sum_8[12] = _3338_ ^ _3337_ /*26890*/;
  assign _3339_ = _3338_ & _3337_ /*26889*/;
  assign _3340_ = inv_8[12] & r_7[12] /*26888*/;
  assign _3341_ = _3339_ | _3340_ /*26887*/;
  assign _3342_ = inv_8[13] ^ r_7[13] /*26885*/;
  assign sum_8[13] = _3342_ ^ _3341_ /*26884*/;
  assign _3343_ = _3342_ & _3341_ /*26883*/;
  assign _3344_ = inv_8[13] & r_7[13] /*26882*/;
  assign _3345_ = _3343_ | _3344_ /*26881*/;
  assign _3346_ = inv_8[14] ^ r_7[14] /*26879*/;
  assign sum_8[14] = _3346_ ^ _3345_ /*26878*/;
  assign _3347_ = _3346_ & _3345_ /*26877*/;
  assign _3348_ = inv_8[14] & r_7[14] /*26876*/;
  assign _3349_ = _3347_ | _3348_ /*26875*/;
  assign _3350_ = inv_8[15] ^ r_7[15] /*26873*/;
  assign sum_8[15] = _3350_ ^ _3349_ /*26872*/;
  assign _3351_ = _3350_ & _3349_ /*26871*/;
  assign _3352_ = inv_8[15] & r_7[15] /*26870*/;
  assign _3353_ = _3351_ | _3352_ /*26869*/;
  assign _3354_ = inv_8[16] ^ r_7[16] /*26867*/;
  assign sum_8[16] = _3354_ ^ _3353_ /*26866*/;
  assign _3355_ = _3354_ & _3353_ /*26865*/;
  assign _3356_ = inv_8[16] & r_7[16] /*26864*/;
  assign _3357_ = _3355_ | _3356_ /*26863*/;
  assign _3358_ = inv_8[17] ^ r_7[17] /*26861*/;
  assign sum_8[17] = _3358_ ^ _3357_ /*26860*/;
  assign _3359_ = _3358_ & _3357_ /*26859*/;
  assign _3360_ = inv_8[17] & r_7[17] /*26858*/;
  assign _3361_ = _3359_ | _3360_ /*26857*/;
  assign _3362_ = inv_8[18] ^ r_7[18] /*26855*/;
  assign sum_8[18] = _3362_ ^ _3361_ /*26854*/;
  assign _3363_ = _3362_ & _3361_ /*26853*/;
  assign _3364_ = inv_8[18] & r_7[18] /*26852*/;
  assign _3365_ = _3363_ | _3364_ /*26851*/;
  assign _3366_ = inv_8[19] ^ r_7[19] /*26849*/;
  assign sum_8[19] = _3366_ ^ _3365_ /*26848*/;
  assign _3367_ = _3366_ & _3365_ /*26847*/;
  assign _3368_ = inv_8[19] & r_7[19] /*26846*/;
  assign _3369_ = _3367_ | _3368_ /*26845*/;
  assign _3370_ = inv_8[20] ^ r_7[20] /*26843*/;
  assign sum_8[20] = _3370_ ^ _3369_ /*26842*/;
  assign _3371_ = _3370_ & _3369_ /*26841*/;
  assign _3372_ = inv_8[20] & r_7[20] /*26840*/;
  assign _3373_ = _3371_ | _3372_ /*26839*/;
  assign _3374_ = inv_8[21] ^ r_7[21] /*26837*/;
  assign sum_8[21] = _3374_ ^ _3373_ /*26836*/;
  assign _3375_ = _3374_ & _3373_ /*26835*/;
  assign _3376_ = inv_8[21] & r_7[21] /*26834*/;
  assign _3377_ = _3375_ | _3376_ /*26833*/;
  assign _3378_ = inv_8[22] ^ r_7[22] /*26831*/;
  assign sum_8[22] = _3378_ ^ _3377_ /*26830*/;
  assign _3379_ = _3378_ & _3377_ /*26829*/;
  assign _3380_ = inv_8[22] & r_7[22] /*26828*/;
  assign _3381_ = _3379_ | _3380_ /*26827*/;
  assign _3382_ = inv_8[23] ^ r_7[23] /*26825*/;
  assign sum_8[23] = _3382_ ^ _3381_ /*26824*/;
  assign _3383_ = _3382_ & _3381_ /*26823*/;
  assign _3384_ = inv_8[23] & r_7[23] /*26822*/;
  assign _3385_ = _3383_ | _3384_ /*26821*/;
  assign _3386_ = inv_8[24] ^ r_7[24] /*26819*/;
  assign sum_8[24] = _3386_ ^ _3385_ /*26818*/;
  assign _3387_ = _3386_ & _3385_ /*26817*/;
  assign _3388_ = inv_8[24] & r_7[24] /*26816*/;
  assign _3389_ = _3387_ | _3388_ /*26815*/;
  assign _3390_ = inv_8[25] ^ r_7[25] /*26813*/;
  assign sum_8[25] = _3390_ ^ _3389_ /*26812*/;
  assign _3391_ = _3390_ & _3389_ /*26811*/;
  assign _3392_ = inv_8[25] & r_7[25] /*26810*/;
  assign _3393_ = _3391_ | _3392_ /*26809*/;
  assign _3394_ = inv_8[26] ^ r_7[26] /*26807*/;
  assign sum_8[26] = _3394_ ^ _3393_ /*26806*/;
  assign _3395_ = _3394_ & _3393_ /*26805*/;
  assign _3396_ = inv_8[26] & r_7[26] /*26804*/;
  assign _3397_ = _3395_ | _3396_ /*26803*/;
  assign _3398_ = inv_8[27] ^ r_7[27] /*26801*/;
  assign sum_8[27] = _3398_ ^ _3397_ /*26800*/;
  assign _3399_ = _3398_ & _3397_ /*26799*/;
  assign _3400_ = inv_8[27] & r_7[27] /*26798*/;
  assign _3401_ = _3399_ | _3400_ /*26797*/;
  assign _3402_ = inv_8[28] ^ r_7[28] /*26795*/;
  assign sum_8[28] = _3402_ ^ _3401_ /*26794*/;
  assign _3403_ = _3402_ & _3401_ /*26793*/;
  assign _3404_ = inv_8[28] & r_7[28] /*26792*/;
  assign _3405_ = _3403_ | _3404_ /*26791*/;
  assign _3406_ = inv_8[29] ^ r_7[29] /*26789*/;
  assign sum_8[29] = _3406_ ^ _3405_ /*26788*/;
  assign _3407_ = _3406_ & _3405_ /*26787*/;
  assign _3408_ = inv_8[29] & r_7[29] /*26786*/;
  assign _3409_ = _3407_ | _3408_ /*26785*/;
  assign _3410_ = inv_8[30] ^ r_7[30] /*26783*/;
  assign sum_8[30] = _3410_ ^ _3409_ /*26782*/;
  assign _3411_ = _3410_ & _3409_ /*26781*/;
  assign _3412_ = inv_8[30] & r_7[30] /*26780*/;
  assign _3413_ = _3411_ | _3412_ /*26779*/;
  assign _3414_ = inv_8[31] ^ r_7[31] /*26777*/;
  assign sum_8[31] = _3414_ ^ _3413_ /*26776*/;
  assign _3415_ = _3414_ & _3413_ /*26775*/;
  assign _3416_ = inv_8[31] & r_7[31] /*26774*/;
  assign _3417_ = _3415_ | _3416_ /*26773*/;
  assign _3418_ = inv_8[32] ^ r_7[32] /*26771*/;
  assign sum_8[32] = _3418_ ^ _3417_ /*26770*/;
  assign _3419_ = _3418_ & _3417_ /*26769*/;
  assign _3420_ = inv_8[32] & r_7[32] /*26768*/;
  assign _3421_ = _3419_ | _3420_ /*26767*/;
  assign _3422_ = inv_8[33] ^ r_7[33] /*26765*/;
  assign sum_8[33] = _3422_ ^ _3421_ /*26764*/;
  assign _3423_ = _3422_ & _3421_ /*26763*/;
  assign _3424_ = inv_8[33] & r_7[33] /*26762*/;
  assign _3425_ = _3423_ | _3424_ /*26761*/;
  assign _3426_ = inv_8[34] ^ r_7[34] /*26759*/;
  assign sum_8[34] = _3426_ ^ _3425_ /*26758*/;
  assign _3427_ = _3426_ & _3425_ /*26757*/;
  assign _3428_ = inv_8[34] & r_7[34] /*26756*/;
  assign _3429_ = _3427_ | _3428_ /*26755*/;
  assign _3430_ = inv_8[35] ^ r_7[35] /*26753*/;
  assign sum_8[35] = _3430_ ^ _3429_ /*26752*/;
  assign _3431_ = _3430_ & _3429_ /*26751*/;
  assign _3432_ = inv_8[35] & r_7[35] /*26750*/;
  assign _3433_ = _3431_ | _3432_ /*26749*/;
  assign _3434_ = inv_8[36] ^ r_7[36] /*26747*/;
  assign sum_8[36] = _3434_ ^ _3433_ /*26746*/;
  assign _3435_ = _3434_ & _3433_ /*26745*/;
  assign _3436_ = inv_8[36] & r_7[36] /*26744*/;
  assign _3437_ = _3435_ | _3436_ /*26743*/;
  assign _3438_ = inv_8[37] ^ r_7[37] /*26741*/;
  assign sum_8[37] = _3438_ ^ _3437_ /*26740*/;
  assign _3439_ = _3438_ & _3437_ /*26739*/;
  assign _3440_ = inv_8[37] & r_7[37] /*26738*/;
  assign _3441_ = _3439_ | _3440_ /*26737*/;
  assign _3442_ = inv_8[38] ^ r_7[38] /*26735*/;
  assign sum_8[38] = _3442_ ^ _3441_ /*26734*/;
  assign _3443_ = _3442_ & _3441_ /*26733*/;
  assign _3444_ = inv_8[38] & r_7[38] /*26732*/;
  assign _3445_ = _3443_ | _3444_ /*26731*/;
  assign _3446_ = inv_8[39] ^ r_7[39] /*26729*/;
  assign sum_8[39] = _3446_ ^ _3445_ /*26728*/;
  assign _3447_ = _3446_ & _3445_ /*26727*/;
  assign _3448_ = inv_8[39] & r_7[39] /*26726*/;
  assign _3449_ = _3447_ | _3448_ /*26725*/;
  assign _3450_ = inv_8[40] ^ r_7[40] /*26723*/;
  assign sum_8[40] = _3450_ ^ _3449_ /*26722*/;
  assign _3451_ = _3450_ & _3449_ /*26721*/;
  assign _3452_ = inv_8[40] & r_7[40] /*26720*/;
  assign _3453_ = _3451_ | _3452_ /*26719*/;
  assign _3454_ = inv_8[41] ^ r_7[41] /*26717*/;
  assign sum_8[41] = _3454_ ^ _3453_ /*26716*/;
  assign _3455_ = _3454_ & _3453_ /*26715*/;
  assign _3456_ = inv_8[41] & r_7[41] /*26714*/;
  assign _3457_ = _3455_ | _3456_ /*26713*/;
  assign _3458_ = inv_8[42] ^ r_7[42] /*26711*/;
  assign sum_8[42] = _3458_ ^ _3457_ /*26710*/;
  assign _3459_ = _3458_ & _3457_ /*26709*/;
  assign _3460_ = inv_8[42] & r_7[42] /*26708*/;
  assign _3461_ = _3459_ | _3460_ /*26707*/;
  assign _3462_ = inv_8[43] ^ r_7[43] /*26705*/;
  assign sum_8[43] = _3462_ ^ _3461_ /*26704*/;
  assign _3463_ = _3462_ & _3461_ /*26703*/;
  assign _3464_ = inv_8[43] & r_7[43] /*26702*/;
  assign _3465_ = _3463_ | _3464_ /*26701*/;
  assign _3466_ = inv_8[44] ^ r_7[44] /*26699*/;
  assign sum_8[44] = _3466_ ^ _3465_ /*26698*/;
  assign _3467_ = _3466_ & _3465_ /*26697*/;
  assign _3468_ = inv_8[44] & r_7[44] /*26696*/;
  assign _3469_ = _3467_ | _3468_ /*26695*/;
  assign _3470_ = inv_8[45] ^ r_7[45] /*26693*/;
  assign sum_8[45] = _3470_ ^ _3469_ /*26692*/;
  assign _3471_ = _3470_ & _3469_ /*26691*/;
  assign _3472_ = inv_8[45] & r_7[45] /*26690*/;
  assign _3473_ = _3471_ | _3472_ /*26689*/;
  assign _3474_ = inv_8[46] ^ r_7[46] /*26687*/;
  assign sum_8[46] = _3474_ ^ _3473_ /*26686*/;
  assign _3475_ = _3474_ & _3473_ /*26685*/;
  assign _3476_ = inv_8[46] & r_7[46] /*26684*/;
  assign _3477_ = _3475_ | _3476_ /*26683*/;
  assign _3478_ = inv_8[47] ^ r_7[47] /*26681*/;
  assign sum_8[47] = _3478_ ^ _3477_ /*26680*/;
  assign _3479_ = _3478_ & _3477_ /*26679*/;
  assign _3480_ = inv_8[47] & r_7[47] /*26678*/;
  assign _3481_ = _3479_ | _3480_ /*26677*/;
  assign _3482_ = inv_8[48] ^ r_7[48] /*26675*/;
  assign sum_8[48] = _3482_ ^ _3481_ /*26674*/;
  assign _3483_ = _3482_ & _3481_ /*26673*/;
  assign _3484_ = inv_8[48] & r_7[48] /*26672*/;
  assign _3485_ = _3483_ | _3484_ /*26671*/;
  assign _3486_ = inv_8[49] ^ r_7[49] /*26669*/;
  assign sum_8[49] = _3486_ ^ _3485_ /*26668*/;
  assign _3487_ = _3486_ & _3485_ /*26667*/;
  assign _3488_ = inv_8[49] & r_7[49] /*26666*/;
  assign _3489_ = _3487_ | _3488_ /*26665*/;
  assign _3490_ = inv_8[50] ^ r_7[50] /*26663*/;
  assign sum_8[50] = _3490_ ^ _3489_ /*26662*/;
  assign _3491_ = _3490_ & _3489_ /*26661*/;
  assign _3492_ = inv_8[50] & r_7[50] /*26660*/;
  assign _3493_ = _3491_ | _3492_ /*26659*/;
  assign _3494_ = inv_8[51] ^ r_7[51] /*26657*/;
  assign sum_8[51] = _3494_ ^ _3493_ /*26656*/;
  assign _3495_ = _3494_ & _3493_ /*26655*/;
  assign _3496_ = inv_8[51] & r_7[51] /*26654*/;
  assign _3497_ = _3495_ | _3496_ /*26653*/;
  assign _3498_ = inv_8[52] ^ r_7[52] /*26651*/;
  assign sum_8[52] = _3498_ ^ _3497_ /*26650*/;
  assign _3499_ = _3498_ & _3497_ /*26649*/;
  assign _3500_ = inv_8[52] & r_7[52] /*26648*/;
  assign _3501_ = _3499_ | _3500_ /*26647*/;
  assign _3502_ = inv_8[53] ^ r_7[53] /*26645*/;
  assign sum_8[53] = _3502_ ^ _3501_ /*26644*/;
  assign _3503_ = _3502_ & _3501_ /*26643*/;
  assign _3504_ = inv_8[53] & r_7[53] /*26642*/;
  assign _3505_ = _3503_ | _3504_ /*26641*/;
  assign _3506_ = inv_8[54] ^ r_7[54] /*26639*/;
  assign sum_8[54] = _3506_ ^ _3505_ /*26638*/;
  assign _3507_ = _3506_ & _3505_ /*26637*/;
  assign _3508_ = inv_8[54] & r_7[54] /*26636*/;
  assign _3509_ = _3507_ | _3508_ /*26635*/;
  assign _3510_ = inv_8[55] ^ r_7[55] /*26633*/;
  assign sum_8[55] = _3510_ ^ _3509_ /*26632*/;
  assign _3511_ = _3510_ & _3509_ /*26631*/;
  assign _3512_ = inv_8[55] & r_7[55] /*26630*/;
  assign _3513_ = _3511_ | _3512_ /*26629*/;
  assign _3514_ = inv_8[56] ^ r_7[56] /*26627*/;
  assign sum_8[56] = _3514_ ^ _3513_ /*26626*/;
  assign _3515_ = _3514_ & _3513_ /*26625*/;
  assign _3516_ = inv_8[56] & r_7[56] /*26624*/;
  assign _3517_ = _3515_ | _3516_ /*26623*/;
  assign _3518_ = inv_8[57] ^ r_7[57] /*26621*/;
  assign sum_8[57] = _3518_ ^ _3517_ /*26620*/;
  assign _3519_ = _3518_ & _3517_ /*26619*/;
  assign _3520_ = inv_8[57] & r_7[57] /*26618*/;
  assign _3521_ = _3519_ | _3520_ /*26617*/;
  assign _3522_ = inv_8[58] ^ r_7[58] /*26615*/;
  assign sum_8[58] = _3522_ ^ _3521_ /*26614*/;
  assign _3523_ = _3522_ & _3521_ /*26613*/;
  assign _3524_ = inv_8[58] & r_7[58] /*26612*/;
  assign _3525_ = _3523_ | _3524_ /*26611*/;
  assign _3526_ = inv_8[59] ^ r_7[59] /*26609*/;
  assign sum_8[59] = _3526_ ^ _3525_ /*26608*/;
  assign _3527_ = _3526_ & _3525_ /*26607*/;
  assign _3528_ = inv_8[59] & r_7[59] /*26606*/;
  assign _3529_ = _3527_ | _3528_ /*26605*/;
  assign _3530_ = inv_8[60] ^ r_7[60] /*26603*/;
  assign sum_8[60] = _3530_ ^ _3529_ /*26602*/;
  assign _3531_ = _3530_ & _3529_ /*26601*/;
  assign _3532_ = inv_8[60] & r_7[60] /*26600*/;
  assign _3533_ = _3531_ | _3532_ /*26599*/;
  assign _3534_ = inv_8[61] ^ r_7[61] /*26597*/;
  assign sum_8[61] = _3534_ ^ _3533_ /*26596*/;
  assign _3535_ = _3534_ & _3533_ /*26595*/;
  assign _3536_ = inv_8[61] & r_7[61] /*26594*/;
  assign _3537_ = _3535_ | _3536_ /*26593*/;
  assign _3538_ = inv_8[62] ^ r_7[62] /*26591*/;
  assign sum_8[62] = _3538_ ^ _3537_ /*26590*/;
  assign _3539_ = _3538_ & _3537_ /*26589*/;
  assign _3540_ = inv_8[62] & r_7[62] /*26588*/;
  assign _3541_ = _3539_ | _3540_ /*26587*/;
  assign _3542_ = inv_8[63] ^ r_7[63] /*26585*/;
  assign sum_8[63] = _3542_ ^ _3541_ /*26584*/;
  assign _3543_ = _3542_ & _3541_ /*26583*/;
  assign _3544_ = inv_8[63] & r_7[63] /*26582*/;
  assign _3545_ = _3543_ | _3544_ /*26581*/;
  assign _3546_ = inv_8[64] ^ r_7[64] /*26579*/;
  assign sum_8[64] = _3546_ ^ _3545_ /*26578*/;
  assign _3547_ = _3546_ & _3545_ /*26577*/;
  assign _3548_ = inv_8[64] & r_7[64] /*26576*/;
  assign _3549_ = _3547_ | _3548_ /*26575*/;
  assign _3550_ = inv_8[65] ^ r_7[65] /*26573*/;
  assign sum_8[65] = _3550_ ^ _3549_ /*26572*/;
  assign _3551_ = _3550_ & _3549_ /*26571*/;
  assign _3552_ = inv_8[65] & r_7[65] /*26570*/;
  assign _3553_ = _3551_ | _3552_ /*26569*/;
  assign _3554_ = inv_8[66] ^ r_7[66] /*26567*/;
  assign sum_8[66] = _3554_ ^ _3553_ /*26566*/;
  assign _3555_ = _3554_ & _3553_ /*26565*/;
  assign _3556_ = inv_8[66] & r_7[66] /*26564*/;
  assign _3557_ = _3555_ | _3556_ /*26563*/;
  assign _3558_ = inv_8[67] ^ r_7[67] /*26561*/;
  assign sum_8[67] = _3558_ ^ _3557_ /*26560*/;
  assign _3559_ = _3558_ & _3557_ /*26559*/;
  assign _3560_ = inv_8[67] & r_7[67] /*26558*/;
  assign _3561_ = _3559_ | _3560_ /*26557*/;
  assign _3562_ = inv_8[68] ^ r_7[68] /*26555*/;
  assign sum_8[68] = _3562_ ^ _3561_ /*26554*/;
  assign _3563_ = _3562_ & _3561_ /*26553*/;
  assign _3564_ = inv_8[68] & r_7[68] /*26552*/;
  assign _3565_ = _3563_ | _3564_ /*26551*/;
  assign _3566_ = inv_8[69] ^ r_7[69] /*26549*/;
  assign sum_8[69] = _3566_ ^ _3565_ /*26548*/;
  assign _3567_ = _3566_ & _3565_ /*26547*/;
  assign _3568_ = inv_8[69] & r_7[69] /*26546*/;
  assign _3569_ = _3567_ | _3568_ /*26545*/;
  assign _3570_ = _3569_ ^ _3565_ /*26544*/;
  assign _3571_ = ~_3570_ /*26543*/;
  assign _3572_ = sum_8[69] & _3571_ /*26542*/;
  assign _3573_ = _3570_ & _3569_ /*26541*/;
  assign sum_8[70] = _3573_ | _3572_ /*26540*/;
  assign q[24] = ~sum_8[70] /*26539*/;
  assign m_8[0] = r_7[0] /*26538*/;
  assign m_8[1] = r_7[1] /*26537*/;
  assign m_8[2] = r_7[2] /*26536*/;
  assign m_8[3] = r_7[3] /*26535*/;
  assign m_8[4] = r_7[4] /*26534*/;
  assign m_8[5] = r_7[5] /*26533*/;
  assign m_8[6] = r_7[6] /*26532*/;
  assign m_8[7] = r_7[7] /*26531*/;
  assign m_8[8] = r_7[8] /*26530*/;
  assign m_8[9] = r_7[9] /*26529*/;
  assign m_8[10] = r_7[10] /*26528*/;
  assign m_8[11] = r_7[11] /*26527*/;
  assign m_8[12] = r_7[12] /*26526*/;
  assign m_8[13] = r_7[13] /*26525*/;
  assign m_8[14] = r_7[14] /*26524*/;
  assign m_8[15] = r_7[15] /*26523*/;
  assign m_8[16] = r_7[16] /*26522*/;
  assign m_8[17] = r_7[17] /*26521*/;
  assign m_8[18] = r_7[18] /*26520*/;
  assign m_8[19] = r_7[19] /*26519*/;
  assign m_8[20] = r_7[20] /*26518*/;
  assign m_8[21] = r_7[21] /*26517*/;
  assign m_8[22] = r_7[22] /*26516*/;
  assign m_8[23] = r_7[23] /*26515*/;
  assign m_8[24] = r_7[24] /*26514*/;
  assign m_8[25] = r_7[25] /*26513*/;
  assign m_8[26] = r_7[26] /*26512*/;
  assign m_8[27] = r_7[27] /*26511*/;
  assign m_8[28] = r_7[28] /*26510*/;
  assign m_8[29] = r_7[29] /*26509*/;
  assign m_8[30] = r_7[30] /*26508*/;
  assign m_8[31] = r_7[31] /*26507*/;
  assign m_8[32] = r_7[32] /*26506*/;
  assign m_8[33] = r_7[33] /*26505*/;
  assign m_8[34] = r_7[34] /*26504*/;
  assign m_8[35] = r_7[35] /*26503*/;
  assign m_8[36] = r_7[36] /*26502*/;
  assign m_8[37] = r_7[37] /*26501*/;
  assign m_8[38] = r_7[38] /*26500*/;
  assign m_8[39] = r_7[39] /*26499*/;
  assign m_8[40] = r_7[40] /*26498*/;
  assign m_8[41] = r_7[41] /*26497*/;
  assign m_8[42] = r_7[42] /*26496*/;
  assign m_8[43] = r_7[43] /*26495*/;
  assign m_8[44] = r_7[44] /*26494*/;
  assign m_8[45] = r_7[45] /*26493*/;
  assign m_8[46] = r_7[46] /*26492*/;
  assign m_8[47] = r_7[47] /*26491*/;
  assign m_8[48] = r_7[48] /*26490*/;
  assign m_8[49] = r_7[49] /*26489*/;
  assign m_8[50] = r_7[50] /*26488*/;
  assign m_8[51] = r_7[51] /*26487*/;
  assign m_8[52] = r_7[52] /*26486*/;
  assign m_8[53] = r_7[53] /*26485*/;
  assign m_8[54] = r_7[54] /*26484*/;
  assign m_8[55] = r_7[55] /*26483*/;
  assign m_8[56] = r_7[56] /*26482*/;
  assign m_8[57] = r_7[57] /*26481*/;
  assign m_8[58] = r_7[58] /*26480*/;
  assign m_8[59] = r_7[59] /*26479*/;
  assign m_8[60] = r_7[60] /*26478*/;
  assign m_8[61] = r_7[61] /*26477*/;
  assign m_8[62] = r_7[62] /*26476*/;
  assign m_8[63] = r_7[63] /*26475*/;
  assign m_8[64] = r_7[64] /*26474*/;
  assign m_8[65] = r_7[65] /*26473*/;
  assign m_8[66] = r_7[66] /*26472*/;
  assign m_8[67] = r_7[67] /*26471*/;
  assign m_8[68] = r_7[68] /*26470*/;
  assign m_8[69] = r_7[69] /*26469*/;
  assign m_8[70] = r_7[69] /*26468*/;
  assign _3575_ = ~q[24] /*26467*/;
  assign _3576_ = sum_8[0] & q[24] /*26466*/;
  assign _3577_ = m_8[0] & _3575_ /*26465*/;
  assign r_8[0] = _3577_ | _3576_ /*26464*/;
  assign _3578_ = ~q[24] /*26463*/;
  assign _3579_ = sum_8[1] & q[24] /*26462*/;
  assign _3580_ = m_8[1] & _3578_ /*26461*/;
  assign r_8[1] = _3580_ | _3579_ /*26460*/;
  assign _3581_ = ~q[24] /*26459*/;
  assign _3582_ = sum_8[2] & q[24] /*26458*/;
  assign _3583_ = m_8[2] & _3581_ /*26457*/;
  assign r_8[2] = _3583_ | _3582_ /*26456*/;
  assign _3584_ = ~q[24] /*26455*/;
  assign _3585_ = sum_8[3] & q[24] /*26454*/;
  assign _3586_ = m_8[3] & _3584_ /*26453*/;
  assign r_8[3] = _3586_ | _3585_ /*26452*/;
  assign _3587_ = ~q[24] /*26451*/;
  assign _3588_ = sum_8[4] & q[24] /*26450*/;
  assign _3589_ = m_8[4] & _3587_ /*26449*/;
  assign r_8[4] = _3589_ | _3588_ /*26448*/;
  assign _3590_ = ~q[24] /*26447*/;
  assign _3591_ = sum_8[5] & q[24] /*26446*/;
  assign _3592_ = m_8[5] & _3590_ /*26445*/;
  assign r_8[5] = _3592_ | _3591_ /*26444*/;
  assign _3593_ = ~q[24] /*26443*/;
  assign _3594_ = sum_8[6] & q[24] /*26442*/;
  assign _3595_ = m_8[6] & _3593_ /*26441*/;
  assign r_8[6] = _3595_ | _3594_ /*26440*/;
  assign _3596_ = ~q[24] /*26439*/;
  assign _3597_ = sum_8[7] & q[24] /*26438*/;
  assign _3598_ = m_8[7] & _3596_ /*26437*/;
  assign r_8[7] = _3598_ | _3597_ /*26436*/;
  assign _3599_ = ~q[24] /*26435*/;
  assign _3600_ = sum_8[8] & q[24] /*26434*/;
  assign _3601_ = m_8[8] & _3599_ /*26433*/;
  assign r_8[8] = _3601_ | _3600_ /*26432*/;
  assign _3602_ = ~q[24] /*26431*/;
  assign _3603_ = sum_8[9] & q[24] /*26430*/;
  assign _3604_ = m_8[9] & _3602_ /*26429*/;
  assign r_8[9] = _3604_ | _3603_ /*26428*/;
  assign _3605_ = ~q[24] /*26427*/;
  assign _3606_ = sum_8[10] & q[24] /*26426*/;
  assign _3607_ = m_8[10] & _3605_ /*26425*/;
  assign r_8[10] = _3607_ | _3606_ /*26424*/;
  assign _3608_ = ~q[24] /*26423*/;
  assign _3609_ = sum_8[11] & q[24] /*26422*/;
  assign _3610_ = m_8[11] & _3608_ /*26421*/;
  assign r_8[11] = _3610_ | _3609_ /*26420*/;
  assign _3611_ = ~q[24] /*26419*/;
  assign _3612_ = sum_8[12] & q[24] /*26418*/;
  assign _3613_ = m_8[12] & _3611_ /*26417*/;
  assign r_8[12] = _3613_ | _3612_ /*26416*/;
  assign _3614_ = ~q[24] /*26415*/;
  assign _3615_ = sum_8[13] & q[24] /*26414*/;
  assign _3616_ = m_8[13] & _3614_ /*26413*/;
  assign r_8[13] = _3616_ | _3615_ /*26412*/;
  assign _3617_ = ~q[24] /*26411*/;
  assign _3618_ = sum_8[14] & q[24] /*26410*/;
  assign _3619_ = m_8[14] & _3617_ /*26409*/;
  assign r_8[14] = _3619_ | _3618_ /*26408*/;
  assign _3620_ = ~q[24] /*26407*/;
  assign _3621_ = sum_8[15] & q[24] /*26406*/;
  assign _3622_ = m_8[15] & _3620_ /*26405*/;
  assign r_8[15] = _3622_ | _3621_ /*26404*/;
  assign _3623_ = ~q[24] /*26403*/;
  assign _3624_ = sum_8[16] & q[24] /*26402*/;
  assign _3625_ = m_8[16] & _3623_ /*26401*/;
  assign r_8[16] = _3625_ | _3624_ /*26400*/;
  assign _3626_ = ~q[24] /*26399*/;
  assign _3627_ = sum_8[17] & q[24] /*26398*/;
  assign _3628_ = m_8[17] & _3626_ /*26397*/;
  assign r_8[17] = _3628_ | _3627_ /*26396*/;
  assign _3629_ = ~q[24] /*26395*/;
  assign _3630_ = sum_8[18] & q[24] /*26394*/;
  assign _3631_ = m_8[18] & _3629_ /*26393*/;
  assign r_8[18] = _3631_ | _3630_ /*26392*/;
  assign _3632_ = ~q[24] /*26391*/;
  assign _3633_ = sum_8[19] & q[24] /*26390*/;
  assign _3634_ = m_8[19] & _3632_ /*26389*/;
  assign r_8[19] = _3634_ | _3633_ /*26388*/;
  assign _3635_ = ~q[24] /*26387*/;
  assign _3636_ = sum_8[20] & q[24] /*26386*/;
  assign _3637_ = m_8[20] & _3635_ /*26385*/;
  assign r_8[20] = _3637_ | _3636_ /*26384*/;
  assign _3638_ = ~q[24] /*26383*/;
  assign _3639_ = sum_8[21] & q[24] /*26382*/;
  assign _3640_ = m_8[21] & _3638_ /*26381*/;
  assign r_8[21] = _3640_ | _3639_ /*26380*/;
  assign _3641_ = ~q[24] /*26379*/;
  assign _3642_ = sum_8[22] & q[24] /*26378*/;
  assign _3643_ = m_8[22] & _3641_ /*26377*/;
  assign r_8[22] = _3643_ | _3642_ /*26376*/;
  assign _3644_ = ~q[24] /*26375*/;
  assign _3645_ = sum_8[23] & q[24] /*26374*/;
  assign _3646_ = m_8[23] & _3644_ /*26373*/;
  assign r_8[23] = _3646_ | _3645_ /*26372*/;
  assign _3647_ = ~q[24] /*26371*/;
  assign _3648_ = sum_8[24] & q[24] /*26370*/;
  assign _3649_ = m_8[24] & _3647_ /*26369*/;
  assign r_8[24] = _3649_ | _3648_ /*26368*/;
  assign _3650_ = ~q[24] /*26367*/;
  assign _3651_ = sum_8[25] & q[24] /*26366*/;
  assign _3652_ = m_8[25] & _3650_ /*26365*/;
  assign r_8[25] = _3652_ | _3651_ /*26364*/;
  assign _3653_ = ~q[24] /*26363*/;
  assign _3654_ = sum_8[26] & q[24] /*26362*/;
  assign _3655_ = m_8[26] & _3653_ /*26361*/;
  assign r_8[26] = _3655_ | _3654_ /*26360*/;
  assign _3656_ = ~q[24] /*26359*/;
  assign _3657_ = sum_8[27] & q[24] /*26358*/;
  assign _3658_ = m_8[27] & _3656_ /*26357*/;
  assign r_8[27] = _3658_ | _3657_ /*26356*/;
  assign _3659_ = ~q[24] /*26355*/;
  assign _3660_ = sum_8[28] & q[24] /*26354*/;
  assign _3661_ = m_8[28] & _3659_ /*26353*/;
  assign r_8[28] = _3661_ | _3660_ /*26352*/;
  assign _3662_ = ~q[24] /*26351*/;
  assign _3663_ = sum_8[29] & q[24] /*26350*/;
  assign _3664_ = m_8[29] & _3662_ /*26349*/;
  assign r_8[29] = _3664_ | _3663_ /*26348*/;
  assign _3665_ = ~q[24] /*26347*/;
  assign _3666_ = sum_8[30] & q[24] /*26346*/;
  assign _3667_ = m_8[30] & _3665_ /*26345*/;
  assign r_8[30] = _3667_ | _3666_ /*26344*/;
  assign _3668_ = ~q[24] /*26343*/;
  assign _3669_ = sum_8[31] & q[24] /*26342*/;
  assign _3670_ = m_8[31] & _3668_ /*26341*/;
  assign r_8[31] = _3670_ | _3669_ /*26340*/;
  assign _3671_ = ~q[24] /*26339*/;
  assign _3672_ = sum_8[32] & q[24] /*26338*/;
  assign _3673_ = m_8[32] & _3671_ /*26337*/;
  assign r_8[32] = _3673_ | _3672_ /*26336*/;
  assign _3674_ = ~q[24] /*26335*/;
  assign _3675_ = sum_8[33] & q[24] /*26334*/;
  assign _3676_ = m_8[33] & _3674_ /*26333*/;
  assign r_8[33] = _3676_ | _3675_ /*26332*/;
  assign _3677_ = ~q[24] /*26331*/;
  assign _3678_ = sum_8[34] & q[24] /*26330*/;
  assign _3679_ = m_8[34] & _3677_ /*26329*/;
  assign r_8[34] = _3679_ | _3678_ /*26328*/;
  assign _3680_ = ~q[24] /*26327*/;
  assign _3681_ = sum_8[35] & q[24] /*26326*/;
  assign _3682_ = m_8[35] & _3680_ /*26325*/;
  assign r_8[35] = _3682_ | _3681_ /*26324*/;
  assign _3683_ = ~q[24] /*26323*/;
  assign _3684_ = sum_8[36] & q[24] /*26322*/;
  assign _3685_ = m_8[36] & _3683_ /*26321*/;
  assign r_8[36] = _3685_ | _3684_ /*26320*/;
  assign _3686_ = ~q[24] /*26319*/;
  assign _3687_ = sum_8[37] & q[24] /*26318*/;
  assign _3688_ = m_8[37] & _3686_ /*26317*/;
  assign r_8[37] = _3688_ | _3687_ /*26316*/;
  assign _3689_ = ~q[24] /*26315*/;
  assign _3690_ = sum_8[38] & q[24] /*26314*/;
  assign _3691_ = m_8[38] & _3689_ /*26313*/;
  assign r_8[38] = _3691_ | _3690_ /*26312*/;
  assign _3692_ = ~q[24] /*26311*/;
  assign _3693_ = sum_8[39] & q[24] /*26310*/;
  assign _3694_ = m_8[39] & _3692_ /*26309*/;
  assign r_8[39] = _3694_ | _3693_ /*26308*/;
  assign _3695_ = ~q[24] /*26307*/;
  assign _3696_ = sum_8[40] & q[24] /*26306*/;
  assign _3697_ = m_8[40] & _3695_ /*26305*/;
  assign r_8[40] = _3697_ | _3696_ /*26304*/;
  assign _3698_ = ~q[24] /*26303*/;
  assign _3699_ = sum_8[41] & q[24] /*26302*/;
  assign _3700_ = m_8[41] & _3698_ /*26301*/;
  assign r_8[41] = _3700_ | _3699_ /*26300*/;
  assign _3701_ = ~q[24] /*26299*/;
  assign _3702_ = sum_8[42] & q[24] /*26298*/;
  assign _3703_ = m_8[42] & _3701_ /*26297*/;
  assign r_8[42] = _3703_ | _3702_ /*26296*/;
  assign _3704_ = ~q[24] /*26295*/;
  assign _3705_ = sum_8[43] & q[24] /*26294*/;
  assign _3706_ = m_8[43] & _3704_ /*26293*/;
  assign r_8[43] = _3706_ | _3705_ /*26292*/;
  assign _3707_ = ~q[24] /*26291*/;
  assign _3708_ = sum_8[44] & q[24] /*26290*/;
  assign _3709_ = m_8[44] & _3707_ /*26289*/;
  assign r_8[44] = _3709_ | _3708_ /*26288*/;
  assign _3710_ = ~q[24] /*26287*/;
  assign _3711_ = sum_8[45] & q[24] /*26286*/;
  assign _3712_ = m_8[45] & _3710_ /*26285*/;
  assign r_8[45] = _3712_ | _3711_ /*26284*/;
  assign _3713_ = ~q[24] /*26283*/;
  assign _3714_ = sum_8[46] & q[24] /*26282*/;
  assign _3715_ = m_8[46] & _3713_ /*26281*/;
  assign r_8[46] = _3715_ | _3714_ /*26280*/;
  assign _3716_ = ~q[24] /*26279*/;
  assign _3717_ = sum_8[47] & q[24] /*26278*/;
  assign _3718_ = m_8[47] & _3716_ /*26277*/;
  assign r_8[47] = _3718_ | _3717_ /*26276*/;
  assign _3719_ = ~q[24] /*26275*/;
  assign _3720_ = sum_8[48] & q[24] /*26274*/;
  assign _3721_ = m_8[48] & _3719_ /*26273*/;
  assign r_8[48] = _3721_ | _3720_ /*26272*/;
  assign _3722_ = ~q[24] /*26271*/;
  assign _3723_ = sum_8[49] & q[24] /*26270*/;
  assign _3724_ = m_8[49] & _3722_ /*26269*/;
  assign r_8[49] = _3724_ | _3723_ /*26268*/;
  assign _3725_ = ~q[24] /*26267*/;
  assign _3726_ = sum_8[50] & q[24] /*26266*/;
  assign _3727_ = m_8[50] & _3725_ /*26265*/;
  assign r_8[50] = _3727_ | _3726_ /*26264*/;
  assign _3728_ = ~q[24] /*26263*/;
  assign _3729_ = sum_8[51] & q[24] /*26262*/;
  assign _3730_ = m_8[51] & _3728_ /*26261*/;
  assign r_8[51] = _3730_ | _3729_ /*26260*/;
  assign _3731_ = ~q[24] /*26259*/;
  assign _3732_ = sum_8[52] & q[24] /*26258*/;
  assign _3733_ = m_8[52] & _3731_ /*26257*/;
  assign r_8[52] = _3733_ | _3732_ /*26256*/;
  assign _3734_ = ~q[24] /*26255*/;
  assign _3735_ = sum_8[53] & q[24] /*26254*/;
  assign _3736_ = m_8[53] & _3734_ /*26253*/;
  assign r_8[53] = _3736_ | _3735_ /*26252*/;
  assign _3737_ = ~q[24] /*26251*/;
  assign _3738_ = sum_8[54] & q[24] /*26250*/;
  assign _3739_ = m_8[54] & _3737_ /*26249*/;
  assign r_8[54] = _3739_ | _3738_ /*26248*/;
  assign _3740_ = ~q[24] /*26247*/;
  assign _3741_ = sum_8[55] & q[24] /*26246*/;
  assign _3742_ = m_8[55] & _3740_ /*26245*/;
  assign r_8[55] = _3742_ | _3741_ /*26244*/;
  assign _3743_ = ~q[24] /*26243*/;
  assign _3744_ = sum_8[56] & q[24] /*26242*/;
  assign _3745_ = m_8[56] & _3743_ /*26241*/;
  assign r_8[56] = _3745_ | _3744_ /*26240*/;
  assign _3746_ = ~q[24] /*26239*/;
  assign _3747_ = sum_8[57] & q[24] /*26238*/;
  assign _3748_ = m_8[57] & _3746_ /*26237*/;
  assign r_8[57] = _3748_ | _3747_ /*26236*/;
  assign _3749_ = ~q[24] /*26235*/;
  assign _3750_ = sum_8[58] & q[24] /*26234*/;
  assign _3751_ = m_8[58] & _3749_ /*26233*/;
  assign r_8[58] = _3751_ | _3750_ /*26232*/;
  assign _3752_ = ~q[24] /*26231*/;
  assign _3753_ = sum_8[59] & q[24] /*26230*/;
  assign _3754_ = m_8[59] & _3752_ /*26229*/;
  assign r_8[59] = _3754_ | _3753_ /*26228*/;
  assign _3755_ = ~q[24] /*26227*/;
  assign _3756_ = sum_8[60] & q[24] /*26226*/;
  assign _3757_ = m_8[60] & _3755_ /*26225*/;
  assign r_8[60] = _3757_ | _3756_ /*26224*/;
  assign _3758_ = ~q[24] /*26223*/;
  assign _3759_ = sum_8[61] & q[24] /*26222*/;
  assign _3760_ = m_8[61] & _3758_ /*26221*/;
  assign r_8[61] = _3760_ | _3759_ /*26220*/;
  assign _3761_ = ~q[24] /*26219*/;
  assign _3762_ = sum_8[62] & q[24] /*26218*/;
  assign _3763_ = m_8[62] & _3761_ /*26217*/;
  assign r_8[62] = _3763_ | _3762_ /*26216*/;
  assign _3764_ = ~q[24] /*26215*/;
  assign _3765_ = sum_8[63] & q[24] /*26214*/;
  assign _3766_ = m_8[63] & _3764_ /*26213*/;
  assign r_8[63] = _3766_ | _3765_ /*26212*/;
  assign _3767_ = ~q[24] /*26211*/;
  assign _3768_ = sum_8[64] & q[24] /*26210*/;
  assign _3769_ = m_8[64] & _3767_ /*26209*/;
  assign r_8[64] = _3769_ | _3768_ /*26208*/;
  assign _3770_ = ~q[24] /*26207*/;
  assign _3771_ = sum_8[65] & q[24] /*26206*/;
  assign _3772_ = m_8[65] & _3770_ /*26205*/;
  assign r_8[65] = _3772_ | _3771_ /*26204*/;
  assign _3773_ = ~q[24] /*26203*/;
  assign _3774_ = sum_8[66] & q[24] /*26202*/;
  assign _3775_ = m_8[66] & _3773_ /*26201*/;
  assign r_8[66] = _3775_ | _3774_ /*26200*/;
  assign _3776_ = ~q[24] /*26199*/;
  assign _3777_ = sum_8[67] & q[24] /*26198*/;
  assign _3778_ = m_8[67] & _3776_ /*26197*/;
  assign r_8[67] = _3778_ | _3777_ /*26196*/;
  assign _3779_ = ~q[24] /*26195*/;
  assign _3780_ = sum_8[68] & q[24] /*26194*/;
  assign _3781_ = m_8[68] & _3779_ /*26193*/;
  assign r_8[68] = _3781_ | _3780_ /*26192*/;
  assign _3782_ = ~q[24] /*26191*/;
  assign _3783_ = sum_8[69] & q[24] /*26190*/;
  assign _3784_ = m_8[69] & _3782_ /*26189*/;
  assign r_8[69] = _3784_ | _3783_ /*26188*/;
  assign _3785_ = ~q[24] /*26187*/;
  assign _3786_ = sum_8[70] & q[24] /*26186*/;
  assign _3787_ = m_8[70] & _3785_ /*26185*/;
  assign r_8[70] = _3787_ | _3786_ /*26184*/;
  assign inv_9[0] = oneWire /*25888*/;
  assign inv_9[1] = oneWire /*25882*/;
  assign inv_9[2] = oneWire /*25876*/;
  assign inv_9[3] = oneWire /*25870*/;
  assign inv_9[4] = oneWire /*25864*/;
  assign inv_9[5] = oneWire /*25858*/;
  assign inv_9[6] = oneWire /*25852*/;
  assign inv_9[7] = oneWire /*25846*/;
  assign inv_9[8] = oneWire /*25840*/;
  assign inv_9[9] = oneWire /*25834*/;
  assign inv_9[10] = oneWire /*25828*/;
  assign inv_9[11] = oneWire /*25822*/;
  assign inv_9[12] = oneWire /*25816*/;
  assign inv_9[13] = oneWire /*25810*/;
  assign inv_9[14] = oneWire /*25804*/;
  assign inv_9[15] = oneWire /*25798*/;
  assign inv_9[16] = oneWire /*25792*/;
  assign inv_9[17] = oneWire /*25786*/;
  assign inv_9[18] = oneWire /*25780*/;
  assign inv_9[19] = oneWire /*25774*/;
  assign inv_9[20] = oneWire /*25768*/;
  assign inv_9[21] = oneWire /*25762*/;
  assign inv_9[22] = oneWire /*25756*/;
  assign inv_9[23] = ~div[0] /*25750*/;
  assign inv_9[24] = ~div[1] /*25744*/;
  assign inv_9[25] = ~div[2] /*25738*/;
  assign inv_9[26] = ~div[3] /*25732*/;
  assign inv_9[27] = ~div[4] /*25726*/;
  assign inv_9[28] = ~div[5] /*25720*/;
  assign inv_9[29] = ~div[6] /*25714*/;
  assign inv_9[30] = ~div[7] /*25708*/;
  assign inv_9[31] = ~div[8] /*25702*/;
  assign inv_9[32] = ~div[9] /*25696*/;
  assign inv_9[33] = ~div[10] /*25690*/;
  assign inv_9[34] = ~div[11] /*25684*/;
  assign inv_9[35] = ~div[12] /*25678*/;
  assign inv_9[36] = ~div[13] /*25672*/;
  assign inv_9[37] = ~div[14] /*25666*/;
  assign inv_9[38] = ~div[15] /*25660*/;
  assign inv_9[39] = ~div[16] /*25654*/;
  assign inv_9[40] = ~div[17] /*25648*/;
  assign inv_9[41] = ~div[18] /*25642*/;
  assign inv_9[42] = ~div[19] /*25636*/;
  assign inv_9[43] = ~div[20] /*25630*/;
  assign inv_9[44] = ~div[21] /*25624*/;
  assign inv_9[45] = ~div[22] /*25618*/;
  assign inv_9[46] = ~div[23] /*25612*/;
  assign inv_9[47] = ~div[24] /*25606*/;
  assign inv_9[48] = ~div[25] /*25600*/;
  assign inv_9[49] = ~div[26] /*25594*/;
  assign inv_9[50] = ~div[27] /*25588*/;
  assign inv_9[51] = ~div[28] /*25582*/;
  assign inv_9[52] = ~div[29] /*25576*/;
  assign inv_9[53] = ~div[30] /*25570*/;
  assign inv_9[54] = oneWire /*25564*/;
  assign inv_9[55] = oneWire /*25558*/;
  assign inv_9[56] = oneWire /*25552*/;
  assign inv_9[57] = oneWire /*25546*/;
  assign inv_9[58] = oneWire /*25540*/;
  assign inv_9[59] = oneWire /*25534*/;
  assign inv_9[60] = oneWire /*25528*/;
  assign inv_9[61] = oneWire /*25522*/;
  assign inv_9[62] = oneWire /*25516*/;
  assign inv_9[63] = oneWire /*25510*/;
  assign inv_9[64] = oneWire /*25504*/;
  assign inv_9[65] = oneWire /*25498*/;
  assign inv_9[66] = oneWire /*25492*/;
  assign inv_9[67] = oneWire /*25486*/;
  assign inv_9[68] = oneWire /*25480*/;
  assign inv_9[69] = oneWire /*25474*/;
  assign inv_9[70] = oneWire /*25468*/;
  assign _3788_ = inv_9[0] ^ r_8[0] /*25887*/;
  assign sum_9[0] = _3788_ ^ oneWire /*25886*/;
  assign _3789_ = _3788_ & oneWire /*25885*/;
  assign _3790_ = inv_9[0] & r_8[0] /*25884*/;
  assign _3791_ = _3789_ | _3790_ /*25883*/;
  assign _3792_ = inv_9[1] ^ r_8[1] /*25881*/;
  assign sum_9[1] = _3792_ ^ _3791_ /*25880*/;
  assign _3793_ = _3792_ & _3791_ /*25879*/;
  assign _3794_ = inv_9[1] & r_8[1] /*25878*/;
  assign _3795_ = _3793_ | _3794_ /*25877*/;
  assign _3796_ = inv_9[2] ^ r_8[2] /*25875*/;
  assign sum_9[2] = _3796_ ^ _3795_ /*25874*/;
  assign _3797_ = _3796_ & _3795_ /*25873*/;
  assign _3798_ = inv_9[2] & r_8[2] /*25872*/;
  assign _3799_ = _3797_ | _3798_ /*25871*/;
  assign _3800_ = inv_9[3] ^ r_8[3] /*25869*/;
  assign sum_9[3] = _3800_ ^ _3799_ /*25868*/;
  assign _3801_ = _3800_ & _3799_ /*25867*/;
  assign _3802_ = inv_9[3] & r_8[3] /*25866*/;
  assign _3803_ = _3801_ | _3802_ /*25865*/;
  assign _3804_ = inv_9[4] ^ r_8[4] /*25863*/;
  assign sum_9[4] = _3804_ ^ _3803_ /*25862*/;
  assign _3805_ = _3804_ & _3803_ /*25861*/;
  assign _3806_ = inv_9[4] & r_8[4] /*25860*/;
  assign _3807_ = _3805_ | _3806_ /*25859*/;
  assign _3808_ = inv_9[5] ^ r_8[5] /*25857*/;
  assign sum_9[5] = _3808_ ^ _3807_ /*25856*/;
  assign _3809_ = _3808_ & _3807_ /*25855*/;
  assign _3810_ = inv_9[5] & r_8[5] /*25854*/;
  assign _3811_ = _3809_ | _3810_ /*25853*/;
  assign _3812_ = inv_9[6] ^ r_8[6] /*25851*/;
  assign sum_9[6] = _3812_ ^ _3811_ /*25850*/;
  assign _3813_ = _3812_ & _3811_ /*25849*/;
  assign _3814_ = inv_9[6] & r_8[6] /*25848*/;
  assign _3815_ = _3813_ | _3814_ /*25847*/;
  assign _3816_ = inv_9[7] ^ r_8[7] /*25845*/;
  assign sum_9[7] = _3816_ ^ _3815_ /*25844*/;
  assign _3817_ = _3816_ & _3815_ /*25843*/;
  assign _3818_ = inv_9[7] & r_8[7] /*25842*/;
  assign _3819_ = _3817_ | _3818_ /*25841*/;
  assign _3820_ = inv_9[8] ^ r_8[8] /*25839*/;
  assign sum_9[8] = _3820_ ^ _3819_ /*25838*/;
  assign _3821_ = _3820_ & _3819_ /*25837*/;
  assign _3822_ = inv_9[8] & r_8[8] /*25836*/;
  assign _3823_ = _3821_ | _3822_ /*25835*/;
  assign _3824_ = inv_9[9] ^ r_8[9] /*25833*/;
  assign sum_9[9] = _3824_ ^ _3823_ /*25832*/;
  assign _3825_ = _3824_ & _3823_ /*25831*/;
  assign _3826_ = inv_9[9] & r_8[9] /*25830*/;
  assign _3827_ = _3825_ | _3826_ /*25829*/;
  assign _3828_ = inv_9[10] ^ r_8[10] /*25827*/;
  assign sum_9[10] = _3828_ ^ _3827_ /*25826*/;
  assign _3829_ = _3828_ & _3827_ /*25825*/;
  assign _3830_ = inv_9[10] & r_8[10] /*25824*/;
  assign _3831_ = _3829_ | _3830_ /*25823*/;
  assign _3832_ = inv_9[11] ^ r_8[11] /*25821*/;
  assign sum_9[11] = _3832_ ^ _3831_ /*25820*/;
  assign _3833_ = _3832_ & _3831_ /*25819*/;
  assign _3834_ = inv_9[11] & r_8[11] /*25818*/;
  assign _3835_ = _3833_ | _3834_ /*25817*/;
  assign _3836_ = inv_9[12] ^ r_8[12] /*25815*/;
  assign sum_9[12] = _3836_ ^ _3835_ /*25814*/;
  assign _3837_ = _3836_ & _3835_ /*25813*/;
  assign _3838_ = inv_9[12] & r_8[12] /*25812*/;
  assign _3839_ = _3837_ | _3838_ /*25811*/;
  assign _3840_ = inv_9[13] ^ r_8[13] /*25809*/;
  assign sum_9[13] = _3840_ ^ _3839_ /*25808*/;
  assign _3841_ = _3840_ & _3839_ /*25807*/;
  assign _3842_ = inv_9[13] & r_8[13] /*25806*/;
  assign _3843_ = _3841_ | _3842_ /*25805*/;
  assign _3844_ = inv_9[14] ^ r_8[14] /*25803*/;
  assign sum_9[14] = _3844_ ^ _3843_ /*25802*/;
  assign _3845_ = _3844_ & _3843_ /*25801*/;
  assign _3846_ = inv_9[14] & r_8[14] /*25800*/;
  assign _3847_ = _3845_ | _3846_ /*25799*/;
  assign _3848_ = inv_9[15] ^ r_8[15] /*25797*/;
  assign sum_9[15] = _3848_ ^ _3847_ /*25796*/;
  assign _3849_ = _3848_ & _3847_ /*25795*/;
  assign _3850_ = inv_9[15] & r_8[15] /*25794*/;
  assign _3851_ = _3849_ | _3850_ /*25793*/;
  assign _3852_ = inv_9[16] ^ r_8[16] /*25791*/;
  assign sum_9[16] = _3852_ ^ _3851_ /*25790*/;
  assign _3853_ = _3852_ & _3851_ /*25789*/;
  assign _3854_ = inv_9[16] & r_8[16] /*25788*/;
  assign _3855_ = _3853_ | _3854_ /*25787*/;
  assign _3856_ = inv_9[17] ^ r_8[17] /*25785*/;
  assign sum_9[17] = _3856_ ^ _3855_ /*25784*/;
  assign _3857_ = _3856_ & _3855_ /*25783*/;
  assign _3858_ = inv_9[17] & r_8[17] /*25782*/;
  assign _3859_ = _3857_ | _3858_ /*25781*/;
  assign _3860_ = inv_9[18] ^ r_8[18] /*25779*/;
  assign sum_9[18] = _3860_ ^ _3859_ /*25778*/;
  assign _3861_ = _3860_ & _3859_ /*25777*/;
  assign _3862_ = inv_9[18] & r_8[18] /*25776*/;
  assign _3863_ = _3861_ | _3862_ /*25775*/;
  assign _3864_ = inv_9[19] ^ r_8[19] /*25773*/;
  assign sum_9[19] = _3864_ ^ _3863_ /*25772*/;
  assign _3865_ = _3864_ & _3863_ /*25771*/;
  assign _3866_ = inv_9[19] & r_8[19] /*25770*/;
  assign _3867_ = _3865_ | _3866_ /*25769*/;
  assign _3868_ = inv_9[20] ^ r_8[20] /*25767*/;
  assign sum_9[20] = _3868_ ^ _3867_ /*25766*/;
  assign _3869_ = _3868_ & _3867_ /*25765*/;
  assign _3870_ = inv_9[20] & r_8[20] /*25764*/;
  assign _3871_ = _3869_ | _3870_ /*25763*/;
  assign _3872_ = inv_9[21] ^ r_8[21] /*25761*/;
  assign sum_9[21] = _3872_ ^ _3871_ /*25760*/;
  assign _3873_ = _3872_ & _3871_ /*25759*/;
  assign _3874_ = inv_9[21] & r_8[21] /*25758*/;
  assign _3875_ = _3873_ | _3874_ /*25757*/;
  assign _3876_ = inv_9[22] ^ r_8[22] /*25755*/;
  assign sum_9[22] = _3876_ ^ _3875_ /*25754*/;
  assign _3877_ = _3876_ & _3875_ /*25753*/;
  assign _3878_ = inv_9[22] & r_8[22] /*25752*/;
  assign _3879_ = _3877_ | _3878_ /*25751*/;
  assign _3880_ = inv_9[23] ^ r_8[23] /*25749*/;
  assign sum_9[23] = _3880_ ^ _3879_ /*25748*/;
  assign _3881_ = _3880_ & _3879_ /*25747*/;
  assign _3882_ = inv_9[23] & r_8[23] /*25746*/;
  assign _3883_ = _3881_ | _3882_ /*25745*/;
  assign _3884_ = inv_9[24] ^ r_8[24] /*25743*/;
  assign sum_9[24] = _3884_ ^ _3883_ /*25742*/;
  assign _3885_ = _3884_ & _3883_ /*25741*/;
  assign _3886_ = inv_9[24] & r_8[24] /*25740*/;
  assign _3887_ = _3885_ | _3886_ /*25739*/;
  assign _3888_ = inv_9[25] ^ r_8[25] /*25737*/;
  assign sum_9[25] = _3888_ ^ _3887_ /*25736*/;
  assign _3889_ = _3888_ & _3887_ /*25735*/;
  assign _3890_ = inv_9[25] & r_8[25] /*25734*/;
  assign _3891_ = _3889_ | _3890_ /*25733*/;
  assign _3892_ = inv_9[26] ^ r_8[26] /*25731*/;
  assign sum_9[26] = _3892_ ^ _3891_ /*25730*/;
  assign _3893_ = _3892_ & _3891_ /*25729*/;
  assign _3894_ = inv_9[26] & r_8[26] /*25728*/;
  assign _3895_ = _3893_ | _3894_ /*25727*/;
  assign _3896_ = inv_9[27] ^ r_8[27] /*25725*/;
  assign sum_9[27] = _3896_ ^ _3895_ /*25724*/;
  assign _3897_ = _3896_ & _3895_ /*25723*/;
  assign _3898_ = inv_9[27] & r_8[27] /*25722*/;
  assign _3899_ = _3897_ | _3898_ /*25721*/;
  assign _3900_ = inv_9[28] ^ r_8[28] /*25719*/;
  assign sum_9[28] = _3900_ ^ _3899_ /*25718*/;
  assign _3901_ = _3900_ & _3899_ /*25717*/;
  assign _3902_ = inv_9[28] & r_8[28] /*25716*/;
  assign _3903_ = _3901_ | _3902_ /*25715*/;
  assign _3904_ = inv_9[29] ^ r_8[29] /*25713*/;
  assign sum_9[29] = _3904_ ^ _3903_ /*25712*/;
  assign _3905_ = _3904_ & _3903_ /*25711*/;
  assign _3906_ = inv_9[29] & r_8[29] /*25710*/;
  assign _3907_ = _3905_ | _3906_ /*25709*/;
  assign _3908_ = inv_9[30] ^ r_8[30] /*25707*/;
  assign sum_9[30] = _3908_ ^ _3907_ /*25706*/;
  assign _3909_ = _3908_ & _3907_ /*25705*/;
  assign _3910_ = inv_9[30] & r_8[30] /*25704*/;
  assign _3911_ = _3909_ | _3910_ /*25703*/;
  assign _3912_ = inv_9[31] ^ r_8[31] /*25701*/;
  assign sum_9[31] = _3912_ ^ _3911_ /*25700*/;
  assign _3913_ = _3912_ & _3911_ /*25699*/;
  assign _3914_ = inv_9[31] & r_8[31] /*25698*/;
  assign _3915_ = _3913_ | _3914_ /*25697*/;
  assign _3916_ = inv_9[32] ^ r_8[32] /*25695*/;
  assign sum_9[32] = _3916_ ^ _3915_ /*25694*/;
  assign _3917_ = _3916_ & _3915_ /*25693*/;
  assign _3918_ = inv_9[32] & r_8[32] /*25692*/;
  assign _3919_ = _3917_ | _3918_ /*25691*/;
  assign _3920_ = inv_9[33] ^ r_8[33] /*25689*/;
  assign sum_9[33] = _3920_ ^ _3919_ /*25688*/;
  assign _3921_ = _3920_ & _3919_ /*25687*/;
  assign _3922_ = inv_9[33] & r_8[33] /*25686*/;
  assign _3923_ = _3921_ | _3922_ /*25685*/;
  assign _3924_ = inv_9[34] ^ r_8[34] /*25683*/;
  assign sum_9[34] = _3924_ ^ _3923_ /*25682*/;
  assign _3925_ = _3924_ & _3923_ /*25681*/;
  assign _3926_ = inv_9[34] & r_8[34] /*25680*/;
  assign _3927_ = _3925_ | _3926_ /*25679*/;
  assign _3928_ = inv_9[35] ^ r_8[35] /*25677*/;
  assign sum_9[35] = _3928_ ^ _3927_ /*25676*/;
  assign _3929_ = _3928_ & _3927_ /*25675*/;
  assign _3930_ = inv_9[35] & r_8[35] /*25674*/;
  assign _3931_ = _3929_ | _3930_ /*25673*/;
  assign _3932_ = inv_9[36] ^ r_8[36] /*25671*/;
  assign sum_9[36] = _3932_ ^ _3931_ /*25670*/;
  assign _3933_ = _3932_ & _3931_ /*25669*/;
  assign _3934_ = inv_9[36] & r_8[36] /*25668*/;
  assign _3935_ = _3933_ | _3934_ /*25667*/;
  assign _3936_ = inv_9[37] ^ r_8[37] /*25665*/;
  assign sum_9[37] = _3936_ ^ _3935_ /*25664*/;
  assign _3937_ = _3936_ & _3935_ /*25663*/;
  assign _3938_ = inv_9[37] & r_8[37] /*25662*/;
  assign _3939_ = _3937_ | _3938_ /*25661*/;
  assign _3940_ = inv_9[38] ^ r_8[38] /*25659*/;
  assign sum_9[38] = _3940_ ^ _3939_ /*25658*/;
  assign _3941_ = _3940_ & _3939_ /*25657*/;
  assign _3942_ = inv_9[38] & r_8[38] /*25656*/;
  assign _3943_ = _3941_ | _3942_ /*25655*/;
  assign _3944_ = inv_9[39] ^ r_8[39] /*25653*/;
  assign sum_9[39] = _3944_ ^ _3943_ /*25652*/;
  assign _3945_ = _3944_ & _3943_ /*25651*/;
  assign _3946_ = inv_9[39] & r_8[39] /*25650*/;
  assign _3947_ = _3945_ | _3946_ /*25649*/;
  assign _3948_ = inv_9[40] ^ r_8[40] /*25647*/;
  assign sum_9[40] = _3948_ ^ _3947_ /*25646*/;
  assign _3949_ = _3948_ & _3947_ /*25645*/;
  assign _3950_ = inv_9[40] & r_8[40] /*25644*/;
  assign _3951_ = _3949_ | _3950_ /*25643*/;
  assign _3952_ = inv_9[41] ^ r_8[41] /*25641*/;
  assign sum_9[41] = _3952_ ^ _3951_ /*25640*/;
  assign _3953_ = _3952_ & _3951_ /*25639*/;
  assign _3954_ = inv_9[41] & r_8[41] /*25638*/;
  assign _3955_ = _3953_ | _3954_ /*25637*/;
  assign _3956_ = inv_9[42] ^ r_8[42] /*25635*/;
  assign sum_9[42] = _3956_ ^ _3955_ /*25634*/;
  assign _3957_ = _3956_ & _3955_ /*25633*/;
  assign _3958_ = inv_9[42] & r_8[42] /*25632*/;
  assign _3959_ = _3957_ | _3958_ /*25631*/;
  assign _3960_ = inv_9[43] ^ r_8[43] /*25629*/;
  assign sum_9[43] = _3960_ ^ _3959_ /*25628*/;
  assign _3961_ = _3960_ & _3959_ /*25627*/;
  assign _3962_ = inv_9[43] & r_8[43] /*25626*/;
  assign _3963_ = _3961_ | _3962_ /*25625*/;
  assign _3964_ = inv_9[44] ^ r_8[44] /*25623*/;
  assign sum_9[44] = _3964_ ^ _3963_ /*25622*/;
  assign _3965_ = _3964_ & _3963_ /*25621*/;
  assign _3966_ = inv_9[44] & r_8[44] /*25620*/;
  assign _3967_ = _3965_ | _3966_ /*25619*/;
  assign _3968_ = inv_9[45] ^ r_8[45] /*25617*/;
  assign sum_9[45] = _3968_ ^ _3967_ /*25616*/;
  assign _3969_ = _3968_ & _3967_ /*25615*/;
  assign _3970_ = inv_9[45] & r_8[45] /*25614*/;
  assign _3971_ = _3969_ | _3970_ /*25613*/;
  assign _3972_ = inv_9[46] ^ r_8[46] /*25611*/;
  assign sum_9[46] = _3972_ ^ _3971_ /*25610*/;
  assign _3973_ = _3972_ & _3971_ /*25609*/;
  assign _3974_ = inv_9[46] & r_8[46] /*25608*/;
  assign _3975_ = _3973_ | _3974_ /*25607*/;
  assign _3976_ = inv_9[47] ^ r_8[47] /*25605*/;
  assign sum_9[47] = _3976_ ^ _3975_ /*25604*/;
  assign _3977_ = _3976_ & _3975_ /*25603*/;
  assign _3978_ = inv_9[47] & r_8[47] /*25602*/;
  assign _3979_ = _3977_ | _3978_ /*25601*/;
  assign _3980_ = inv_9[48] ^ r_8[48] /*25599*/;
  assign sum_9[48] = _3980_ ^ _3979_ /*25598*/;
  assign _3981_ = _3980_ & _3979_ /*25597*/;
  assign _3982_ = inv_9[48] & r_8[48] /*25596*/;
  assign _3983_ = _3981_ | _3982_ /*25595*/;
  assign _3984_ = inv_9[49] ^ r_8[49] /*25593*/;
  assign sum_9[49] = _3984_ ^ _3983_ /*25592*/;
  assign _3985_ = _3984_ & _3983_ /*25591*/;
  assign _3986_ = inv_9[49] & r_8[49] /*25590*/;
  assign _3987_ = _3985_ | _3986_ /*25589*/;
  assign _3988_ = inv_9[50] ^ r_8[50] /*25587*/;
  assign sum_9[50] = _3988_ ^ _3987_ /*25586*/;
  assign _3989_ = _3988_ & _3987_ /*25585*/;
  assign _3990_ = inv_9[50] & r_8[50] /*25584*/;
  assign _3991_ = _3989_ | _3990_ /*25583*/;
  assign _3992_ = inv_9[51] ^ r_8[51] /*25581*/;
  assign sum_9[51] = _3992_ ^ _3991_ /*25580*/;
  assign _3993_ = _3992_ & _3991_ /*25579*/;
  assign _3994_ = inv_9[51] & r_8[51] /*25578*/;
  assign _3995_ = _3993_ | _3994_ /*25577*/;
  assign _3996_ = inv_9[52] ^ r_8[52] /*25575*/;
  assign sum_9[52] = _3996_ ^ _3995_ /*25574*/;
  assign _3997_ = _3996_ & _3995_ /*25573*/;
  assign _3998_ = inv_9[52] & r_8[52] /*25572*/;
  assign _3999_ = _3997_ | _3998_ /*25571*/;
  assign _4000_ = inv_9[53] ^ r_8[53] /*25569*/;
  assign sum_9[53] = _4000_ ^ _3999_ /*25568*/;
  assign _4001_ = _4000_ & _3999_ /*25567*/;
  assign _4002_ = inv_9[53] & r_8[53] /*25566*/;
  assign _4003_ = _4001_ | _4002_ /*25565*/;
  assign _4004_ = inv_9[54] ^ r_8[54] /*25563*/;
  assign sum_9[54] = _4004_ ^ _4003_ /*25562*/;
  assign _4005_ = _4004_ & _4003_ /*25561*/;
  assign _4006_ = inv_9[54] & r_8[54] /*25560*/;
  assign _4007_ = _4005_ | _4006_ /*25559*/;
  assign _4008_ = inv_9[55] ^ r_8[55] /*25557*/;
  assign sum_9[55] = _4008_ ^ _4007_ /*25556*/;
  assign _4009_ = _4008_ & _4007_ /*25555*/;
  assign _4010_ = inv_9[55] & r_8[55] /*25554*/;
  assign _4011_ = _4009_ | _4010_ /*25553*/;
  assign _4012_ = inv_9[56] ^ r_8[56] /*25551*/;
  assign sum_9[56] = _4012_ ^ _4011_ /*25550*/;
  assign _4013_ = _4012_ & _4011_ /*25549*/;
  assign _4014_ = inv_9[56] & r_8[56] /*25548*/;
  assign _4015_ = _4013_ | _4014_ /*25547*/;
  assign _4016_ = inv_9[57] ^ r_8[57] /*25545*/;
  assign sum_9[57] = _4016_ ^ _4015_ /*25544*/;
  assign _4017_ = _4016_ & _4015_ /*25543*/;
  assign _4018_ = inv_9[57] & r_8[57] /*25542*/;
  assign _4019_ = _4017_ | _4018_ /*25541*/;
  assign _4020_ = inv_9[58] ^ r_8[58] /*25539*/;
  assign sum_9[58] = _4020_ ^ _4019_ /*25538*/;
  assign _4021_ = _4020_ & _4019_ /*25537*/;
  assign _4022_ = inv_9[58] & r_8[58] /*25536*/;
  assign _4023_ = _4021_ | _4022_ /*25535*/;
  assign _4024_ = inv_9[59] ^ r_8[59] /*25533*/;
  assign sum_9[59] = _4024_ ^ _4023_ /*25532*/;
  assign _4025_ = _4024_ & _4023_ /*25531*/;
  assign _4026_ = inv_9[59] & r_8[59] /*25530*/;
  assign _4027_ = _4025_ | _4026_ /*25529*/;
  assign _4028_ = inv_9[60] ^ r_8[60] /*25527*/;
  assign sum_9[60] = _4028_ ^ _4027_ /*25526*/;
  assign _4029_ = _4028_ & _4027_ /*25525*/;
  assign _4030_ = inv_9[60] & r_8[60] /*25524*/;
  assign _4031_ = _4029_ | _4030_ /*25523*/;
  assign _4032_ = inv_9[61] ^ r_8[61] /*25521*/;
  assign sum_9[61] = _4032_ ^ _4031_ /*25520*/;
  assign _4033_ = _4032_ & _4031_ /*25519*/;
  assign _4034_ = inv_9[61] & r_8[61] /*25518*/;
  assign _4035_ = _4033_ | _4034_ /*25517*/;
  assign _4036_ = inv_9[62] ^ r_8[62] /*25515*/;
  assign sum_9[62] = _4036_ ^ _4035_ /*25514*/;
  assign _4037_ = _4036_ & _4035_ /*25513*/;
  assign _4038_ = inv_9[62] & r_8[62] /*25512*/;
  assign _4039_ = _4037_ | _4038_ /*25511*/;
  assign _4040_ = inv_9[63] ^ r_8[63] /*25509*/;
  assign sum_9[63] = _4040_ ^ _4039_ /*25508*/;
  assign _4041_ = _4040_ & _4039_ /*25507*/;
  assign _4042_ = inv_9[63] & r_8[63] /*25506*/;
  assign _4043_ = _4041_ | _4042_ /*25505*/;
  assign _4044_ = inv_9[64] ^ r_8[64] /*25503*/;
  assign sum_9[64] = _4044_ ^ _4043_ /*25502*/;
  assign _4045_ = _4044_ & _4043_ /*25501*/;
  assign _4046_ = inv_9[64] & r_8[64] /*25500*/;
  assign _4047_ = _4045_ | _4046_ /*25499*/;
  assign _4048_ = inv_9[65] ^ r_8[65] /*25497*/;
  assign sum_9[65] = _4048_ ^ _4047_ /*25496*/;
  assign _4049_ = _4048_ & _4047_ /*25495*/;
  assign _4050_ = inv_9[65] & r_8[65] /*25494*/;
  assign _4051_ = _4049_ | _4050_ /*25493*/;
  assign _4052_ = inv_9[66] ^ r_8[66] /*25491*/;
  assign sum_9[66] = _4052_ ^ _4051_ /*25490*/;
  assign _4053_ = _4052_ & _4051_ /*25489*/;
  assign _4054_ = inv_9[66] & r_8[66] /*25488*/;
  assign _4055_ = _4053_ | _4054_ /*25487*/;
  assign _4056_ = inv_9[67] ^ r_8[67] /*25485*/;
  assign sum_9[67] = _4056_ ^ _4055_ /*25484*/;
  assign _4057_ = _4056_ & _4055_ /*25483*/;
  assign _4058_ = inv_9[67] & r_8[67] /*25482*/;
  assign _4059_ = _4057_ | _4058_ /*25481*/;
  assign _4060_ = inv_9[68] ^ r_8[68] /*25479*/;
  assign sum_9[68] = _4060_ ^ _4059_ /*25478*/;
  assign _4061_ = _4060_ & _4059_ /*25477*/;
  assign _4062_ = inv_9[68] & r_8[68] /*25476*/;
  assign _4063_ = _4061_ | _4062_ /*25475*/;
  assign _4064_ = inv_9[69] ^ r_8[69] /*25473*/;
  assign sum_9[69] = _4064_ ^ _4063_ /*25472*/;
  assign _4065_ = _4064_ & _4063_ /*25471*/;
  assign _4066_ = inv_9[69] & r_8[69] /*25470*/;
  assign _4067_ = _4065_ | _4066_ /*25469*/;
  assign _4068_ = inv_9[70] ^ r_8[70] /*25467*/;
  assign sum_9[70] = _4068_ ^ _4067_ /*25466*/;
  assign _4069_ = _4068_ & _4067_ /*25465*/;
  assign _4070_ = inv_9[70] & r_8[70] /*25464*/;
  assign _4071_ = _4069_ | _4070_ /*25463*/;
  assign _4072_ = _4071_ ^ _4067_ /*25462*/;
  assign _4073_ = ~_4072_ /*25461*/;
  assign _4074_ = sum_9[70] & _4073_ /*25460*/;
  assign _4075_ = _4072_ & _4071_ /*25459*/;
  assign sum_9[71] = _4075_ | _4074_ /*25458*/;
  assign q[23] = ~sum_9[71] /*25457*/;
  assign m_9[0] = r_8[0] /*25456*/;
  assign m_9[1] = r_8[1] /*25455*/;
  assign m_9[2] = r_8[2] /*25454*/;
  assign m_9[3] = r_8[3] /*25453*/;
  assign m_9[4] = r_8[4] /*25452*/;
  assign m_9[5] = r_8[5] /*25451*/;
  assign m_9[6] = r_8[6] /*25450*/;
  assign m_9[7] = r_8[7] /*25449*/;
  assign m_9[8] = r_8[8] /*25448*/;
  assign m_9[9] = r_8[9] /*25447*/;
  assign m_9[10] = r_8[10] /*25446*/;
  assign m_9[11] = r_8[11] /*25445*/;
  assign m_9[12] = r_8[12] /*25444*/;
  assign m_9[13] = r_8[13] /*25443*/;
  assign m_9[14] = r_8[14] /*25442*/;
  assign m_9[15] = r_8[15] /*25441*/;
  assign m_9[16] = r_8[16] /*25440*/;
  assign m_9[17] = r_8[17] /*25439*/;
  assign m_9[18] = r_8[18] /*25438*/;
  assign m_9[19] = r_8[19] /*25437*/;
  assign m_9[20] = r_8[20] /*25436*/;
  assign m_9[21] = r_8[21] /*25435*/;
  assign m_9[22] = r_8[22] /*25434*/;
  assign m_9[23] = r_8[23] /*25433*/;
  assign m_9[24] = r_8[24] /*25432*/;
  assign m_9[25] = r_8[25] /*25431*/;
  assign m_9[26] = r_8[26] /*25430*/;
  assign m_9[27] = r_8[27] /*25429*/;
  assign m_9[28] = r_8[28] /*25428*/;
  assign m_9[29] = r_8[29] /*25427*/;
  assign m_9[30] = r_8[30] /*25426*/;
  assign m_9[31] = r_8[31] /*25425*/;
  assign m_9[32] = r_8[32] /*25424*/;
  assign m_9[33] = r_8[33] /*25423*/;
  assign m_9[34] = r_8[34] /*25422*/;
  assign m_9[35] = r_8[35] /*25421*/;
  assign m_9[36] = r_8[36] /*25420*/;
  assign m_9[37] = r_8[37] /*25419*/;
  assign m_9[38] = r_8[38] /*25418*/;
  assign m_9[39] = r_8[39] /*25417*/;
  assign m_9[40] = r_8[40] /*25416*/;
  assign m_9[41] = r_8[41] /*25415*/;
  assign m_9[42] = r_8[42] /*25414*/;
  assign m_9[43] = r_8[43] /*25413*/;
  assign m_9[44] = r_8[44] /*25412*/;
  assign m_9[45] = r_8[45] /*25411*/;
  assign m_9[46] = r_8[46] /*25410*/;
  assign m_9[47] = r_8[47] /*25409*/;
  assign m_9[48] = r_8[48] /*25408*/;
  assign m_9[49] = r_8[49] /*25407*/;
  assign m_9[50] = r_8[50] /*25406*/;
  assign m_9[51] = r_8[51] /*25405*/;
  assign m_9[52] = r_8[52] /*25404*/;
  assign m_9[53] = r_8[53] /*25403*/;
  assign m_9[54] = r_8[54] /*25402*/;
  assign m_9[55] = r_8[55] /*25401*/;
  assign m_9[56] = r_8[56] /*25400*/;
  assign m_9[57] = r_8[57] /*25399*/;
  assign m_9[58] = r_8[58] /*25398*/;
  assign m_9[59] = r_8[59] /*25397*/;
  assign m_9[60] = r_8[60] /*25396*/;
  assign m_9[61] = r_8[61] /*25395*/;
  assign m_9[62] = r_8[62] /*25394*/;
  assign m_9[63] = r_8[63] /*25393*/;
  assign m_9[64] = r_8[64] /*25392*/;
  assign m_9[65] = r_8[65] /*25391*/;
  assign m_9[66] = r_8[66] /*25390*/;
  assign m_9[67] = r_8[67] /*25389*/;
  assign m_9[68] = r_8[68] /*25388*/;
  assign m_9[69] = r_8[69] /*25387*/;
  assign m_9[70] = r_8[70] /*25386*/;
  assign m_9[71] = r_8[70] /*25385*/;
  assign _4077_ = ~q[23] /*25384*/;
  assign _4078_ = sum_9[0] & q[23] /*25383*/;
  assign _4079_ = m_9[0] & _4077_ /*25382*/;
  assign r_9[0] = _4079_ | _4078_ /*25381*/;
  assign _4080_ = ~q[23] /*25380*/;
  assign _4081_ = sum_9[1] & q[23] /*25379*/;
  assign _4082_ = m_9[1] & _4080_ /*25378*/;
  assign r_9[1] = _4082_ | _4081_ /*25377*/;
  assign _4083_ = ~q[23] /*25376*/;
  assign _4084_ = sum_9[2] & q[23] /*25375*/;
  assign _4085_ = m_9[2] & _4083_ /*25374*/;
  assign r_9[2] = _4085_ | _4084_ /*25373*/;
  assign _4086_ = ~q[23] /*25372*/;
  assign _4087_ = sum_9[3] & q[23] /*25371*/;
  assign _4088_ = m_9[3] & _4086_ /*25370*/;
  assign r_9[3] = _4088_ | _4087_ /*25369*/;
  assign _4089_ = ~q[23] /*25368*/;
  assign _4090_ = sum_9[4] & q[23] /*25367*/;
  assign _4091_ = m_9[4] & _4089_ /*25366*/;
  assign r_9[4] = _4091_ | _4090_ /*25365*/;
  assign _4092_ = ~q[23] /*25364*/;
  assign _4093_ = sum_9[5] & q[23] /*25363*/;
  assign _4094_ = m_9[5] & _4092_ /*25362*/;
  assign r_9[5] = _4094_ | _4093_ /*25361*/;
  assign _4095_ = ~q[23] /*25360*/;
  assign _4096_ = sum_9[6] & q[23] /*25359*/;
  assign _4097_ = m_9[6] & _4095_ /*25358*/;
  assign r_9[6] = _4097_ | _4096_ /*25357*/;
  assign _4098_ = ~q[23] /*25356*/;
  assign _4099_ = sum_9[7] & q[23] /*25355*/;
  assign _4100_ = m_9[7] & _4098_ /*25354*/;
  assign r_9[7] = _4100_ | _4099_ /*25353*/;
  assign _4101_ = ~q[23] /*25352*/;
  assign _4102_ = sum_9[8] & q[23] /*25351*/;
  assign _4103_ = m_9[8] & _4101_ /*25350*/;
  assign r_9[8] = _4103_ | _4102_ /*25349*/;
  assign _4104_ = ~q[23] /*25348*/;
  assign _4105_ = sum_9[9] & q[23] /*25347*/;
  assign _4106_ = m_9[9] & _4104_ /*25346*/;
  assign r_9[9] = _4106_ | _4105_ /*25345*/;
  assign _4107_ = ~q[23] /*25344*/;
  assign _4108_ = sum_9[10] & q[23] /*25343*/;
  assign _4109_ = m_9[10] & _4107_ /*25342*/;
  assign r_9[10] = _4109_ | _4108_ /*25341*/;
  assign _4110_ = ~q[23] /*25340*/;
  assign _4111_ = sum_9[11] & q[23] /*25339*/;
  assign _4112_ = m_9[11] & _4110_ /*25338*/;
  assign r_9[11] = _4112_ | _4111_ /*25337*/;
  assign _4113_ = ~q[23] /*25336*/;
  assign _4114_ = sum_9[12] & q[23] /*25335*/;
  assign _4115_ = m_9[12] & _4113_ /*25334*/;
  assign r_9[12] = _4115_ | _4114_ /*25333*/;
  assign _4116_ = ~q[23] /*25332*/;
  assign _4117_ = sum_9[13] & q[23] /*25331*/;
  assign _4118_ = m_9[13] & _4116_ /*25330*/;
  assign r_9[13] = _4118_ | _4117_ /*25329*/;
  assign _4119_ = ~q[23] /*25328*/;
  assign _4120_ = sum_9[14] & q[23] /*25327*/;
  assign _4121_ = m_9[14] & _4119_ /*25326*/;
  assign r_9[14] = _4121_ | _4120_ /*25325*/;
  assign _4122_ = ~q[23] /*25324*/;
  assign _4123_ = sum_9[15] & q[23] /*25323*/;
  assign _4124_ = m_9[15] & _4122_ /*25322*/;
  assign r_9[15] = _4124_ | _4123_ /*25321*/;
  assign _4125_ = ~q[23] /*25320*/;
  assign _4126_ = sum_9[16] & q[23] /*25319*/;
  assign _4127_ = m_9[16] & _4125_ /*25318*/;
  assign r_9[16] = _4127_ | _4126_ /*25317*/;
  assign _4128_ = ~q[23] /*25316*/;
  assign _4129_ = sum_9[17] & q[23] /*25315*/;
  assign _4130_ = m_9[17] & _4128_ /*25314*/;
  assign r_9[17] = _4130_ | _4129_ /*25313*/;
  assign _4131_ = ~q[23] /*25312*/;
  assign _4132_ = sum_9[18] & q[23] /*25311*/;
  assign _4133_ = m_9[18] & _4131_ /*25310*/;
  assign r_9[18] = _4133_ | _4132_ /*25309*/;
  assign _4134_ = ~q[23] /*25308*/;
  assign _4135_ = sum_9[19] & q[23] /*25307*/;
  assign _4136_ = m_9[19] & _4134_ /*25306*/;
  assign r_9[19] = _4136_ | _4135_ /*25305*/;
  assign _4137_ = ~q[23] /*25304*/;
  assign _4138_ = sum_9[20] & q[23] /*25303*/;
  assign _4139_ = m_9[20] & _4137_ /*25302*/;
  assign r_9[20] = _4139_ | _4138_ /*25301*/;
  assign _4140_ = ~q[23] /*25300*/;
  assign _4141_ = sum_9[21] & q[23] /*25299*/;
  assign _4142_ = m_9[21] & _4140_ /*25298*/;
  assign r_9[21] = _4142_ | _4141_ /*25297*/;
  assign _4143_ = ~q[23] /*25296*/;
  assign _4144_ = sum_9[22] & q[23] /*25295*/;
  assign _4145_ = m_9[22] & _4143_ /*25294*/;
  assign r_9[22] = _4145_ | _4144_ /*25293*/;
  assign _4146_ = ~q[23] /*25292*/;
  assign _4147_ = sum_9[23] & q[23] /*25291*/;
  assign _4148_ = m_9[23] & _4146_ /*25290*/;
  assign r_9[23] = _4148_ | _4147_ /*25289*/;
  assign _4149_ = ~q[23] /*25288*/;
  assign _4150_ = sum_9[24] & q[23] /*25287*/;
  assign _4151_ = m_9[24] & _4149_ /*25286*/;
  assign r_9[24] = _4151_ | _4150_ /*25285*/;
  assign _4152_ = ~q[23] /*25284*/;
  assign _4153_ = sum_9[25] & q[23] /*25283*/;
  assign _4154_ = m_9[25] & _4152_ /*25282*/;
  assign r_9[25] = _4154_ | _4153_ /*25281*/;
  assign _4155_ = ~q[23] /*25280*/;
  assign _4156_ = sum_9[26] & q[23] /*25279*/;
  assign _4157_ = m_9[26] & _4155_ /*25278*/;
  assign r_9[26] = _4157_ | _4156_ /*25277*/;
  assign _4158_ = ~q[23] /*25276*/;
  assign _4159_ = sum_9[27] & q[23] /*25275*/;
  assign _4160_ = m_9[27] & _4158_ /*25274*/;
  assign r_9[27] = _4160_ | _4159_ /*25273*/;
  assign _4161_ = ~q[23] /*25272*/;
  assign _4162_ = sum_9[28] & q[23] /*25271*/;
  assign _4163_ = m_9[28] & _4161_ /*25270*/;
  assign r_9[28] = _4163_ | _4162_ /*25269*/;
  assign _4164_ = ~q[23] /*25268*/;
  assign _4165_ = sum_9[29] & q[23] /*25267*/;
  assign _4166_ = m_9[29] & _4164_ /*25266*/;
  assign r_9[29] = _4166_ | _4165_ /*25265*/;
  assign _4167_ = ~q[23] /*25264*/;
  assign _4168_ = sum_9[30] & q[23] /*25263*/;
  assign _4169_ = m_9[30] & _4167_ /*25262*/;
  assign r_9[30] = _4169_ | _4168_ /*25261*/;
  assign _4170_ = ~q[23] /*25260*/;
  assign _4171_ = sum_9[31] & q[23] /*25259*/;
  assign _4172_ = m_9[31] & _4170_ /*25258*/;
  assign r_9[31] = _4172_ | _4171_ /*25257*/;
  assign _4173_ = ~q[23] /*25256*/;
  assign _4174_ = sum_9[32] & q[23] /*25255*/;
  assign _4175_ = m_9[32] & _4173_ /*25254*/;
  assign r_9[32] = _4175_ | _4174_ /*25253*/;
  assign _4176_ = ~q[23] /*25252*/;
  assign _4177_ = sum_9[33] & q[23] /*25251*/;
  assign _4178_ = m_9[33] & _4176_ /*25250*/;
  assign r_9[33] = _4178_ | _4177_ /*25249*/;
  assign _4179_ = ~q[23] /*25248*/;
  assign _4180_ = sum_9[34] & q[23] /*25247*/;
  assign _4181_ = m_9[34] & _4179_ /*25246*/;
  assign r_9[34] = _4181_ | _4180_ /*25245*/;
  assign _4182_ = ~q[23] /*25244*/;
  assign _4183_ = sum_9[35] & q[23] /*25243*/;
  assign _4184_ = m_9[35] & _4182_ /*25242*/;
  assign r_9[35] = _4184_ | _4183_ /*25241*/;
  assign _4185_ = ~q[23] /*25240*/;
  assign _4186_ = sum_9[36] & q[23] /*25239*/;
  assign _4187_ = m_9[36] & _4185_ /*25238*/;
  assign r_9[36] = _4187_ | _4186_ /*25237*/;
  assign _4188_ = ~q[23] /*25236*/;
  assign _4189_ = sum_9[37] & q[23] /*25235*/;
  assign _4190_ = m_9[37] & _4188_ /*25234*/;
  assign r_9[37] = _4190_ | _4189_ /*25233*/;
  assign _4191_ = ~q[23] /*25232*/;
  assign _4192_ = sum_9[38] & q[23] /*25231*/;
  assign _4193_ = m_9[38] & _4191_ /*25230*/;
  assign r_9[38] = _4193_ | _4192_ /*25229*/;
  assign _4194_ = ~q[23] /*25228*/;
  assign _4195_ = sum_9[39] & q[23] /*25227*/;
  assign _4196_ = m_9[39] & _4194_ /*25226*/;
  assign r_9[39] = _4196_ | _4195_ /*25225*/;
  assign _4197_ = ~q[23] /*25224*/;
  assign _4198_ = sum_9[40] & q[23] /*25223*/;
  assign _4199_ = m_9[40] & _4197_ /*25222*/;
  assign r_9[40] = _4199_ | _4198_ /*25221*/;
  assign _4200_ = ~q[23] /*25220*/;
  assign _4201_ = sum_9[41] & q[23] /*25219*/;
  assign _4202_ = m_9[41] & _4200_ /*25218*/;
  assign r_9[41] = _4202_ | _4201_ /*25217*/;
  assign _4203_ = ~q[23] /*25216*/;
  assign _4204_ = sum_9[42] & q[23] /*25215*/;
  assign _4205_ = m_9[42] & _4203_ /*25214*/;
  assign r_9[42] = _4205_ | _4204_ /*25213*/;
  assign _4206_ = ~q[23] /*25212*/;
  assign _4207_ = sum_9[43] & q[23] /*25211*/;
  assign _4208_ = m_9[43] & _4206_ /*25210*/;
  assign r_9[43] = _4208_ | _4207_ /*25209*/;
  assign _4209_ = ~q[23] /*25208*/;
  assign _4210_ = sum_9[44] & q[23] /*25207*/;
  assign _4211_ = m_9[44] & _4209_ /*25206*/;
  assign r_9[44] = _4211_ | _4210_ /*25205*/;
  assign _4212_ = ~q[23] /*25204*/;
  assign _4213_ = sum_9[45] & q[23] /*25203*/;
  assign _4214_ = m_9[45] & _4212_ /*25202*/;
  assign r_9[45] = _4214_ | _4213_ /*25201*/;
  assign _4215_ = ~q[23] /*25200*/;
  assign _4216_ = sum_9[46] & q[23] /*25199*/;
  assign _4217_ = m_9[46] & _4215_ /*25198*/;
  assign r_9[46] = _4217_ | _4216_ /*25197*/;
  assign _4218_ = ~q[23] /*25196*/;
  assign _4219_ = sum_9[47] & q[23] /*25195*/;
  assign _4220_ = m_9[47] & _4218_ /*25194*/;
  assign r_9[47] = _4220_ | _4219_ /*25193*/;
  assign _4221_ = ~q[23] /*25192*/;
  assign _4222_ = sum_9[48] & q[23] /*25191*/;
  assign _4223_ = m_9[48] & _4221_ /*25190*/;
  assign r_9[48] = _4223_ | _4222_ /*25189*/;
  assign _4224_ = ~q[23] /*25188*/;
  assign _4225_ = sum_9[49] & q[23] /*25187*/;
  assign _4226_ = m_9[49] & _4224_ /*25186*/;
  assign r_9[49] = _4226_ | _4225_ /*25185*/;
  assign _4227_ = ~q[23] /*25184*/;
  assign _4228_ = sum_9[50] & q[23] /*25183*/;
  assign _4229_ = m_9[50] & _4227_ /*25182*/;
  assign r_9[50] = _4229_ | _4228_ /*25181*/;
  assign _4230_ = ~q[23] /*25180*/;
  assign _4231_ = sum_9[51] & q[23] /*25179*/;
  assign _4232_ = m_9[51] & _4230_ /*25178*/;
  assign r_9[51] = _4232_ | _4231_ /*25177*/;
  assign _4233_ = ~q[23] /*25176*/;
  assign _4234_ = sum_9[52] & q[23] /*25175*/;
  assign _4235_ = m_9[52] & _4233_ /*25174*/;
  assign r_9[52] = _4235_ | _4234_ /*25173*/;
  assign _4236_ = ~q[23] /*25172*/;
  assign _4237_ = sum_9[53] & q[23] /*25171*/;
  assign _4238_ = m_9[53] & _4236_ /*25170*/;
  assign r_9[53] = _4238_ | _4237_ /*25169*/;
  assign _4239_ = ~q[23] /*25168*/;
  assign _4240_ = sum_9[54] & q[23] /*25167*/;
  assign _4241_ = m_9[54] & _4239_ /*25166*/;
  assign r_9[54] = _4241_ | _4240_ /*25165*/;
  assign _4242_ = ~q[23] /*25164*/;
  assign _4243_ = sum_9[55] & q[23] /*25163*/;
  assign _4244_ = m_9[55] & _4242_ /*25162*/;
  assign r_9[55] = _4244_ | _4243_ /*25161*/;
  assign _4245_ = ~q[23] /*25160*/;
  assign _4246_ = sum_9[56] & q[23] /*25159*/;
  assign _4247_ = m_9[56] & _4245_ /*25158*/;
  assign r_9[56] = _4247_ | _4246_ /*25157*/;
  assign _4248_ = ~q[23] /*25156*/;
  assign _4249_ = sum_9[57] & q[23] /*25155*/;
  assign _4250_ = m_9[57] & _4248_ /*25154*/;
  assign r_9[57] = _4250_ | _4249_ /*25153*/;
  assign _4251_ = ~q[23] /*25152*/;
  assign _4252_ = sum_9[58] & q[23] /*25151*/;
  assign _4253_ = m_9[58] & _4251_ /*25150*/;
  assign r_9[58] = _4253_ | _4252_ /*25149*/;
  assign _4254_ = ~q[23] /*25148*/;
  assign _4255_ = sum_9[59] & q[23] /*25147*/;
  assign _4256_ = m_9[59] & _4254_ /*25146*/;
  assign r_9[59] = _4256_ | _4255_ /*25145*/;
  assign _4257_ = ~q[23] /*25144*/;
  assign _4258_ = sum_9[60] & q[23] /*25143*/;
  assign _4259_ = m_9[60] & _4257_ /*25142*/;
  assign r_9[60] = _4259_ | _4258_ /*25141*/;
  assign _4260_ = ~q[23] /*25140*/;
  assign _4261_ = sum_9[61] & q[23] /*25139*/;
  assign _4262_ = m_9[61] & _4260_ /*25138*/;
  assign r_9[61] = _4262_ | _4261_ /*25137*/;
  assign _4263_ = ~q[23] /*25136*/;
  assign _4264_ = sum_9[62] & q[23] /*25135*/;
  assign _4265_ = m_9[62] & _4263_ /*25134*/;
  assign r_9[62] = _4265_ | _4264_ /*25133*/;
  assign _4266_ = ~q[23] /*25132*/;
  assign _4267_ = sum_9[63] & q[23] /*25131*/;
  assign _4268_ = m_9[63] & _4266_ /*25130*/;
  assign r_9[63] = _4268_ | _4267_ /*25129*/;
  assign _4269_ = ~q[23] /*25128*/;
  assign _4270_ = sum_9[64] & q[23] /*25127*/;
  assign _4271_ = m_9[64] & _4269_ /*25126*/;
  assign r_9[64] = _4271_ | _4270_ /*25125*/;
  assign _4272_ = ~q[23] /*25124*/;
  assign _4273_ = sum_9[65] & q[23] /*25123*/;
  assign _4274_ = m_9[65] & _4272_ /*25122*/;
  assign r_9[65] = _4274_ | _4273_ /*25121*/;
  assign _4275_ = ~q[23] /*25120*/;
  assign _4276_ = sum_9[66] & q[23] /*25119*/;
  assign _4277_ = m_9[66] & _4275_ /*25118*/;
  assign r_9[66] = _4277_ | _4276_ /*25117*/;
  assign _4278_ = ~q[23] /*25116*/;
  assign _4279_ = sum_9[67] & q[23] /*25115*/;
  assign _4280_ = m_9[67] & _4278_ /*25114*/;
  assign r_9[67] = _4280_ | _4279_ /*25113*/;
  assign _4281_ = ~q[23] /*25112*/;
  assign _4282_ = sum_9[68] & q[23] /*25111*/;
  assign _4283_ = m_9[68] & _4281_ /*25110*/;
  assign r_9[68] = _4283_ | _4282_ /*25109*/;
  assign _4284_ = ~q[23] /*25108*/;
  assign _4285_ = sum_9[69] & q[23] /*25107*/;
  assign _4286_ = m_9[69] & _4284_ /*25106*/;
  assign r_9[69] = _4286_ | _4285_ /*25105*/;
  assign _4287_ = ~q[23] /*25104*/;
  assign _4288_ = sum_9[70] & q[23] /*25103*/;
  assign _4289_ = m_9[70] & _4287_ /*25102*/;
  assign r_9[70] = _4289_ | _4288_ /*25101*/;
  assign _4290_ = ~q[23] /*25100*/;
  assign _4291_ = sum_9[71] & q[23] /*25099*/;
  assign _4292_ = m_9[71] & _4290_ /*25098*/;
  assign r_9[71] = _4292_ | _4291_ /*25097*/;
  assign inv_10[0] = oneWire /*24812*/;
  assign inv_10[1] = oneWire /*24806*/;
  assign inv_10[2] = oneWire /*24800*/;
  assign inv_10[3] = oneWire /*24794*/;
  assign inv_10[4] = oneWire /*24788*/;
  assign inv_10[5] = oneWire /*24782*/;
  assign inv_10[6] = oneWire /*24776*/;
  assign inv_10[7] = oneWire /*24770*/;
  assign inv_10[8] = oneWire /*24764*/;
  assign inv_10[9] = oneWire /*24758*/;
  assign inv_10[10] = oneWire /*24752*/;
  assign inv_10[11] = oneWire /*24746*/;
  assign inv_10[12] = oneWire /*24740*/;
  assign inv_10[13] = oneWire /*24734*/;
  assign inv_10[14] = oneWire /*24728*/;
  assign inv_10[15] = oneWire /*24722*/;
  assign inv_10[16] = oneWire /*24716*/;
  assign inv_10[17] = oneWire /*24710*/;
  assign inv_10[18] = oneWire /*24704*/;
  assign inv_10[19] = oneWire /*24698*/;
  assign inv_10[20] = oneWire /*24692*/;
  assign inv_10[21] = oneWire /*24686*/;
  assign inv_10[22] = ~div[0] /*24680*/;
  assign inv_10[23] = ~div[1] /*24674*/;
  assign inv_10[24] = ~div[2] /*24668*/;
  assign inv_10[25] = ~div[3] /*24662*/;
  assign inv_10[26] = ~div[4] /*24656*/;
  assign inv_10[27] = ~div[5] /*24650*/;
  assign inv_10[28] = ~div[6] /*24644*/;
  assign inv_10[29] = ~div[7] /*24638*/;
  assign inv_10[30] = ~div[8] /*24632*/;
  assign inv_10[31] = ~div[9] /*24626*/;
  assign inv_10[32] = ~div[10] /*24620*/;
  assign inv_10[33] = ~div[11] /*24614*/;
  assign inv_10[34] = ~div[12] /*24608*/;
  assign inv_10[35] = ~div[13] /*24602*/;
  assign inv_10[36] = ~div[14] /*24596*/;
  assign inv_10[37] = ~div[15] /*24590*/;
  assign inv_10[38] = ~div[16] /*24584*/;
  assign inv_10[39] = ~div[17] /*24578*/;
  assign inv_10[40] = ~div[18] /*24572*/;
  assign inv_10[41] = ~div[19] /*24566*/;
  assign inv_10[42] = ~div[20] /*24560*/;
  assign inv_10[43] = ~div[21] /*24554*/;
  assign inv_10[44] = ~div[22] /*24548*/;
  assign inv_10[45] = ~div[23] /*24542*/;
  assign inv_10[46] = ~div[24] /*24536*/;
  assign inv_10[47] = ~div[25] /*24530*/;
  assign inv_10[48] = ~div[26] /*24524*/;
  assign inv_10[49] = ~div[27] /*24518*/;
  assign inv_10[50] = ~div[28] /*24512*/;
  assign inv_10[51] = ~div[29] /*24506*/;
  assign inv_10[52] = ~div[30] /*24500*/;
  assign inv_10[53] = oneWire /*24494*/;
  assign inv_10[54] = oneWire /*24488*/;
  assign inv_10[55] = oneWire /*24482*/;
  assign inv_10[56] = oneWire /*24476*/;
  assign inv_10[57] = oneWire /*24470*/;
  assign inv_10[58] = oneWire /*24464*/;
  assign inv_10[59] = oneWire /*24458*/;
  assign inv_10[60] = oneWire /*24452*/;
  assign inv_10[61] = oneWire /*24446*/;
  assign inv_10[62] = oneWire /*24440*/;
  assign inv_10[63] = oneWire /*24434*/;
  assign inv_10[64] = oneWire /*24428*/;
  assign inv_10[65] = oneWire /*24422*/;
  assign inv_10[66] = oneWire /*24416*/;
  assign inv_10[67] = oneWire /*24410*/;
  assign inv_10[68] = oneWire /*24404*/;
  assign inv_10[69] = oneWire /*24398*/;
  assign inv_10[70] = oneWire /*24392*/;
  assign inv_10[71] = oneWire /*24386*/;
  assign _4293_ = inv_10[0] ^ r_9[0] /*24811*/;
  assign sum_10[0] = _4293_ ^ oneWire /*24810*/;
  assign _4294_ = _4293_ & oneWire /*24809*/;
  assign _4295_ = inv_10[0] & r_9[0] /*24808*/;
  assign _4296_ = _4294_ | _4295_ /*24807*/;
  assign _4297_ = inv_10[1] ^ r_9[1] /*24805*/;
  assign sum_10[1] = _4297_ ^ _4296_ /*24804*/;
  assign _4298_ = _4297_ & _4296_ /*24803*/;
  assign _4299_ = inv_10[1] & r_9[1] /*24802*/;
  assign _4300_ = _4298_ | _4299_ /*24801*/;
  assign _4301_ = inv_10[2] ^ r_9[2] /*24799*/;
  assign sum_10[2] = _4301_ ^ _4300_ /*24798*/;
  assign _4302_ = _4301_ & _4300_ /*24797*/;
  assign _4303_ = inv_10[2] & r_9[2] /*24796*/;
  assign _4304_ = _4302_ | _4303_ /*24795*/;
  assign _4305_ = inv_10[3] ^ r_9[3] /*24793*/;
  assign sum_10[3] = _4305_ ^ _4304_ /*24792*/;
  assign _4306_ = _4305_ & _4304_ /*24791*/;
  assign _4307_ = inv_10[3] & r_9[3] /*24790*/;
  assign _4308_ = _4306_ | _4307_ /*24789*/;
  assign _4309_ = inv_10[4] ^ r_9[4] /*24787*/;
  assign sum_10[4] = _4309_ ^ _4308_ /*24786*/;
  assign _4310_ = _4309_ & _4308_ /*24785*/;
  assign _4311_ = inv_10[4] & r_9[4] /*24784*/;
  assign _4312_ = _4310_ | _4311_ /*24783*/;
  assign _4313_ = inv_10[5] ^ r_9[5] /*24781*/;
  assign sum_10[5] = _4313_ ^ _4312_ /*24780*/;
  assign _4314_ = _4313_ & _4312_ /*24779*/;
  assign _4315_ = inv_10[5] & r_9[5] /*24778*/;
  assign _4316_ = _4314_ | _4315_ /*24777*/;
  assign _4317_ = inv_10[6] ^ r_9[6] /*24775*/;
  assign sum_10[6] = _4317_ ^ _4316_ /*24774*/;
  assign _4318_ = _4317_ & _4316_ /*24773*/;
  assign _4319_ = inv_10[6] & r_9[6] /*24772*/;
  assign _4320_ = _4318_ | _4319_ /*24771*/;
  assign _4321_ = inv_10[7] ^ r_9[7] /*24769*/;
  assign sum_10[7] = _4321_ ^ _4320_ /*24768*/;
  assign _4322_ = _4321_ & _4320_ /*24767*/;
  assign _4323_ = inv_10[7] & r_9[7] /*24766*/;
  assign _4324_ = _4322_ | _4323_ /*24765*/;
  assign _4325_ = inv_10[8] ^ r_9[8] /*24763*/;
  assign sum_10[8] = _4325_ ^ _4324_ /*24762*/;
  assign _4326_ = _4325_ & _4324_ /*24761*/;
  assign _4327_ = inv_10[8] & r_9[8] /*24760*/;
  assign _4328_ = _4326_ | _4327_ /*24759*/;
  assign _4329_ = inv_10[9] ^ r_9[9] /*24757*/;
  assign sum_10[9] = _4329_ ^ _4328_ /*24756*/;
  assign _4330_ = _4329_ & _4328_ /*24755*/;
  assign _4331_ = inv_10[9] & r_9[9] /*24754*/;
  assign _4332_ = _4330_ | _4331_ /*24753*/;
  assign _4333_ = inv_10[10] ^ r_9[10] /*24751*/;
  assign sum_10[10] = _4333_ ^ _4332_ /*24750*/;
  assign _4334_ = _4333_ & _4332_ /*24749*/;
  assign _4335_ = inv_10[10] & r_9[10] /*24748*/;
  assign _4336_ = _4334_ | _4335_ /*24747*/;
  assign _4337_ = inv_10[11] ^ r_9[11] /*24745*/;
  assign sum_10[11] = _4337_ ^ _4336_ /*24744*/;
  assign _4338_ = _4337_ & _4336_ /*24743*/;
  assign _4339_ = inv_10[11] & r_9[11] /*24742*/;
  assign _4340_ = _4338_ | _4339_ /*24741*/;
  assign _4341_ = inv_10[12] ^ r_9[12] /*24739*/;
  assign sum_10[12] = _4341_ ^ _4340_ /*24738*/;
  assign _4342_ = _4341_ & _4340_ /*24737*/;
  assign _4343_ = inv_10[12] & r_9[12] /*24736*/;
  assign _4344_ = _4342_ | _4343_ /*24735*/;
  assign _4345_ = inv_10[13] ^ r_9[13] /*24733*/;
  assign sum_10[13] = _4345_ ^ _4344_ /*24732*/;
  assign _4346_ = _4345_ & _4344_ /*24731*/;
  assign _4347_ = inv_10[13] & r_9[13] /*24730*/;
  assign _4348_ = _4346_ | _4347_ /*24729*/;
  assign _4349_ = inv_10[14] ^ r_9[14] /*24727*/;
  assign sum_10[14] = _4349_ ^ _4348_ /*24726*/;
  assign _4350_ = _4349_ & _4348_ /*24725*/;
  assign _4351_ = inv_10[14] & r_9[14] /*24724*/;
  assign _4352_ = _4350_ | _4351_ /*24723*/;
  assign _4353_ = inv_10[15] ^ r_9[15] /*24721*/;
  assign sum_10[15] = _4353_ ^ _4352_ /*24720*/;
  assign _4354_ = _4353_ & _4352_ /*24719*/;
  assign _4355_ = inv_10[15] & r_9[15] /*24718*/;
  assign _4356_ = _4354_ | _4355_ /*24717*/;
  assign _4357_ = inv_10[16] ^ r_9[16] /*24715*/;
  assign sum_10[16] = _4357_ ^ _4356_ /*24714*/;
  assign _4358_ = _4357_ & _4356_ /*24713*/;
  assign _4359_ = inv_10[16] & r_9[16] /*24712*/;
  assign _4360_ = _4358_ | _4359_ /*24711*/;
  assign _4361_ = inv_10[17] ^ r_9[17] /*24709*/;
  assign sum_10[17] = _4361_ ^ _4360_ /*24708*/;
  assign _4362_ = _4361_ & _4360_ /*24707*/;
  assign _4363_ = inv_10[17] & r_9[17] /*24706*/;
  assign _4364_ = _4362_ | _4363_ /*24705*/;
  assign _4365_ = inv_10[18] ^ r_9[18] /*24703*/;
  assign sum_10[18] = _4365_ ^ _4364_ /*24702*/;
  assign _4366_ = _4365_ & _4364_ /*24701*/;
  assign _4367_ = inv_10[18] & r_9[18] /*24700*/;
  assign _4368_ = _4366_ | _4367_ /*24699*/;
  assign _4369_ = inv_10[19] ^ r_9[19] /*24697*/;
  assign sum_10[19] = _4369_ ^ _4368_ /*24696*/;
  assign _4370_ = _4369_ & _4368_ /*24695*/;
  assign _4371_ = inv_10[19] & r_9[19] /*24694*/;
  assign _4372_ = _4370_ | _4371_ /*24693*/;
  assign _4373_ = inv_10[20] ^ r_9[20] /*24691*/;
  assign sum_10[20] = _4373_ ^ _4372_ /*24690*/;
  assign _4374_ = _4373_ & _4372_ /*24689*/;
  assign _4375_ = inv_10[20] & r_9[20] /*24688*/;
  assign _4376_ = _4374_ | _4375_ /*24687*/;
  assign _4377_ = inv_10[21] ^ r_9[21] /*24685*/;
  assign sum_10[21] = _4377_ ^ _4376_ /*24684*/;
  assign _4378_ = _4377_ & _4376_ /*24683*/;
  assign _4379_ = inv_10[21] & r_9[21] /*24682*/;
  assign _4380_ = _4378_ | _4379_ /*24681*/;
  assign _4381_ = inv_10[22] ^ r_9[22] /*24679*/;
  assign sum_10[22] = _4381_ ^ _4380_ /*24678*/;
  assign _4382_ = _4381_ & _4380_ /*24677*/;
  assign _4383_ = inv_10[22] & r_9[22] /*24676*/;
  assign _4384_ = _4382_ | _4383_ /*24675*/;
  assign _4385_ = inv_10[23] ^ r_9[23] /*24673*/;
  assign sum_10[23] = _4385_ ^ _4384_ /*24672*/;
  assign _4386_ = _4385_ & _4384_ /*24671*/;
  assign _4387_ = inv_10[23] & r_9[23] /*24670*/;
  assign _4388_ = _4386_ | _4387_ /*24669*/;
  assign _4389_ = inv_10[24] ^ r_9[24] /*24667*/;
  assign sum_10[24] = _4389_ ^ _4388_ /*24666*/;
  assign _4390_ = _4389_ & _4388_ /*24665*/;
  assign _4391_ = inv_10[24] & r_9[24] /*24664*/;
  assign _4392_ = _4390_ | _4391_ /*24663*/;
  assign _4393_ = inv_10[25] ^ r_9[25] /*24661*/;
  assign sum_10[25] = _4393_ ^ _4392_ /*24660*/;
  assign _4394_ = _4393_ & _4392_ /*24659*/;
  assign _4395_ = inv_10[25] & r_9[25] /*24658*/;
  assign _4396_ = _4394_ | _4395_ /*24657*/;
  assign _4397_ = inv_10[26] ^ r_9[26] /*24655*/;
  assign sum_10[26] = _4397_ ^ _4396_ /*24654*/;
  assign _4398_ = _4397_ & _4396_ /*24653*/;
  assign _4399_ = inv_10[26] & r_9[26] /*24652*/;
  assign _4400_ = _4398_ | _4399_ /*24651*/;
  assign _4401_ = inv_10[27] ^ r_9[27] /*24649*/;
  assign sum_10[27] = _4401_ ^ _4400_ /*24648*/;
  assign _4402_ = _4401_ & _4400_ /*24647*/;
  assign _4403_ = inv_10[27] & r_9[27] /*24646*/;
  assign _4404_ = _4402_ | _4403_ /*24645*/;
  assign _4405_ = inv_10[28] ^ r_9[28] /*24643*/;
  assign sum_10[28] = _4405_ ^ _4404_ /*24642*/;
  assign _4406_ = _4405_ & _4404_ /*24641*/;
  assign _4407_ = inv_10[28] & r_9[28] /*24640*/;
  assign _4408_ = _4406_ | _4407_ /*24639*/;
  assign _4409_ = inv_10[29] ^ r_9[29] /*24637*/;
  assign sum_10[29] = _4409_ ^ _4408_ /*24636*/;
  assign _4410_ = _4409_ & _4408_ /*24635*/;
  assign _4411_ = inv_10[29] & r_9[29] /*24634*/;
  assign _4412_ = _4410_ | _4411_ /*24633*/;
  assign _4413_ = inv_10[30] ^ r_9[30] /*24631*/;
  assign sum_10[30] = _4413_ ^ _4412_ /*24630*/;
  assign _4414_ = _4413_ & _4412_ /*24629*/;
  assign _4415_ = inv_10[30] & r_9[30] /*24628*/;
  assign _4416_ = _4414_ | _4415_ /*24627*/;
  assign _4417_ = inv_10[31] ^ r_9[31] /*24625*/;
  assign sum_10[31] = _4417_ ^ _4416_ /*24624*/;
  assign _4418_ = _4417_ & _4416_ /*24623*/;
  assign _4419_ = inv_10[31] & r_9[31] /*24622*/;
  assign _4420_ = _4418_ | _4419_ /*24621*/;
  assign _4421_ = inv_10[32] ^ r_9[32] /*24619*/;
  assign sum_10[32] = _4421_ ^ _4420_ /*24618*/;
  assign _4422_ = _4421_ & _4420_ /*24617*/;
  assign _4423_ = inv_10[32] & r_9[32] /*24616*/;
  assign _4424_ = _4422_ | _4423_ /*24615*/;
  assign _4425_ = inv_10[33] ^ r_9[33] /*24613*/;
  assign sum_10[33] = _4425_ ^ _4424_ /*24612*/;
  assign _4426_ = _4425_ & _4424_ /*24611*/;
  assign _4427_ = inv_10[33] & r_9[33] /*24610*/;
  assign _4428_ = _4426_ | _4427_ /*24609*/;
  assign _4429_ = inv_10[34] ^ r_9[34] /*24607*/;
  assign sum_10[34] = _4429_ ^ _4428_ /*24606*/;
  assign _4430_ = _4429_ & _4428_ /*24605*/;
  assign _4431_ = inv_10[34] & r_9[34] /*24604*/;
  assign _4432_ = _4430_ | _4431_ /*24603*/;
  assign _4433_ = inv_10[35] ^ r_9[35] /*24601*/;
  assign sum_10[35] = _4433_ ^ _4432_ /*24600*/;
  assign _4434_ = _4433_ & _4432_ /*24599*/;
  assign _4435_ = inv_10[35] & r_9[35] /*24598*/;
  assign _4436_ = _4434_ | _4435_ /*24597*/;
  assign _4437_ = inv_10[36] ^ r_9[36] /*24595*/;
  assign sum_10[36] = _4437_ ^ _4436_ /*24594*/;
  assign _4438_ = _4437_ & _4436_ /*24593*/;
  assign _4439_ = inv_10[36] & r_9[36] /*24592*/;
  assign _4440_ = _4438_ | _4439_ /*24591*/;
  assign _4441_ = inv_10[37] ^ r_9[37] /*24589*/;
  assign sum_10[37] = _4441_ ^ _4440_ /*24588*/;
  assign _4442_ = _4441_ & _4440_ /*24587*/;
  assign _4443_ = inv_10[37] & r_9[37] /*24586*/;
  assign _4444_ = _4442_ | _4443_ /*24585*/;
  assign _4445_ = inv_10[38] ^ r_9[38] /*24583*/;
  assign sum_10[38] = _4445_ ^ _4444_ /*24582*/;
  assign _4446_ = _4445_ & _4444_ /*24581*/;
  assign _4447_ = inv_10[38] & r_9[38] /*24580*/;
  assign _4448_ = _4446_ | _4447_ /*24579*/;
  assign _4449_ = inv_10[39] ^ r_9[39] /*24577*/;
  assign sum_10[39] = _4449_ ^ _4448_ /*24576*/;
  assign _4450_ = _4449_ & _4448_ /*24575*/;
  assign _4451_ = inv_10[39] & r_9[39] /*24574*/;
  assign _4452_ = _4450_ | _4451_ /*24573*/;
  assign _4453_ = inv_10[40] ^ r_9[40] /*24571*/;
  assign sum_10[40] = _4453_ ^ _4452_ /*24570*/;
  assign _4454_ = _4453_ & _4452_ /*24569*/;
  assign _4455_ = inv_10[40] & r_9[40] /*24568*/;
  assign _4456_ = _4454_ | _4455_ /*24567*/;
  assign _4457_ = inv_10[41] ^ r_9[41] /*24565*/;
  assign sum_10[41] = _4457_ ^ _4456_ /*24564*/;
  assign _4458_ = _4457_ & _4456_ /*24563*/;
  assign _4459_ = inv_10[41] & r_9[41] /*24562*/;
  assign _4460_ = _4458_ | _4459_ /*24561*/;
  assign _4461_ = inv_10[42] ^ r_9[42] /*24559*/;
  assign sum_10[42] = _4461_ ^ _4460_ /*24558*/;
  assign _4462_ = _4461_ & _4460_ /*24557*/;
  assign _4463_ = inv_10[42] & r_9[42] /*24556*/;
  assign _4464_ = _4462_ | _4463_ /*24555*/;
  assign _4465_ = inv_10[43] ^ r_9[43] /*24553*/;
  assign sum_10[43] = _4465_ ^ _4464_ /*24552*/;
  assign _4466_ = _4465_ & _4464_ /*24551*/;
  assign _4467_ = inv_10[43] & r_9[43] /*24550*/;
  assign _4468_ = _4466_ | _4467_ /*24549*/;
  assign _4469_ = inv_10[44] ^ r_9[44] /*24547*/;
  assign sum_10[44] = _4469_ ^ _4468_ /*24546*/;
  assign _4470_ = _4469_ & _4468_ /*24545*/;
  assign _4471_ = inv_10[44] & r_9[44] /*24544*/;
  assign _4472_ = _4470_ | _4471_ /*24543*/;
  assign _4473_ = inv_10[45] ^ r_9[45] /*24541*/;
  assign sum_10[45] = _4473_ ^ _4472_ /*24540*/;
  assign _4474_ = _4473_ & _4472_ /*24539*/;
  assign _4475_ = inv_10[45] & r_9[45] /*24538*/;
  assign _4476_ = _4474_ | _4475_ /*24537*/;
  assign _4477_ = inv_10[46] ^ r_9[46] /*24535*/;
  assign sum_10[46] = _4477_ ^ _4476_ /*24534*/;
  assign _4478_ = _4477_ & _4476_ /*24533*/;
  assign _4479_ = inv_10[46] & r_9[46] /*24532*/;
  assign _4480_ = _4478_ | _4479_ /*24531*/;
  assign _4481_ = inv_10[47] ^ r_9[47] /*24529*/;
  assign sum_10[47] = _4481_ ^ _4480_ /*24528*/;
  assign _4482_ = _4481_ & _4480_ /*24527*/;
  assign _4483_ = inv_10[47] & r_9[47] /*24526*/;
  assign _4484_ = _4482_ | _4483_ /*24525*/;
  assign _4485_ = inv_10[48] ^ r_9[48] /*24523*/;
  assign sum_10[48] = _4485_ ^ _4484_ /*24522*/;
  assign _4486_ = _4485_ & _4484_ /*24521*/;
  assign _4487_ = inv_10[48] & r_9[48] /*24520*/;
  assign _4488_ = _4486_ | _4487_ /*24519*/;
  assign _4489_ = inv_10[49] ^ r_9[49] /*24517*/;
  assign sum_10[49] = _4489_ ^ _4488_ /*24516*/;
  assign _4490_ = _4489_ & _4488_ /*24515*/;
  assign _4491_ = inv_10[49] & r_9[49] /*24514*/;
  assign _4492_ = _4490_ | _4491_ /*24513*/;
  assign _4493_ = inv_10[50] ^ r_9[50] /*24511*/;
  assign sum_10[50] = _4493_ ^ _4492_ /*24510*/;
  assign _4494_ = _4493_ & _4492_ /*24509*/;
  assign _4495_ = inv_10[50] & r_9[50] /*24508*/;
  assign _4496_ = _4494_ | _4495_ /*24507*/;
  assign _4497_ = inv_10[51] ^ r_9[51] /*24505*/;
  assign sum_10[51] = _4497_ ^ _4496_ /*24504*/;
  assign _4498_ = _4497_ & _4496_ /*24503*/;
  assign _4499_ = inv_10[51] & r_9[51] /*24502*/;
  assign _4500_ = _4498_ | _4499_ /*24501*/;
  assign _4501_ = inv_10[52] ^ r_9[52] /*24499*/;
  assign sum_10[52] = _4501_ ^ _4500_ /*24498*/;
  assign _4502_ = _4501_ & _4500_ /*24497*/;
  assign _4503_ = inv_10[52] & r_9[52] /*24496*/;
  assign _4504_ = _4502_ | _4503_ /*24495*/;
  assign _4505_ = inv_10[53] ^ r_9[53] /*24493*/;
  assign sum_10[53] = _4505_ ^ _4504_ /*24492*/;
  assign _4506_ = _4505_ & _4504_ /*24491*/;
  assign _4507_ = inv_10[53] & r_9[53] /*24490*/;
  assign _4508_ = _4506_ | _4507_ /*24489*/;
  assign _4509_ = inv_10[54] ^ r_9[54] /*24487*/;
  assign sum_10[54] = _4509_ ^ _4508_ /*24486*/;
  assign _4510_ = _4509_ & _4508_ /*24485*/;
  assign _4511_ = inv_10[54] & r_9[54] /*24484*/;
  assign _4512_ = _4510_ | _4511_ /*24483*/;
  assign _4513_ = inv_10[55] ^ r_9[55] /*24481*/;
  assign sum_10[55] = _4513_ ^ _4512_ /*24480*/;
  assign _4514_ = _4513_ & _4512_ /*24479*/;
  assign _4515_ = inv_10[55] & r_9[55] /*24478*/;
  assign _4516_ = _4514_ | _4515_ /*24477*/;
  assign _4517_ = inv_10[56] ^ r_9[56] /*24475*/;
  assign sum_10[56] = _4517_ ^ _4516_ /*24474*/;
  assign _4518_ = _4517_ & _4516_ /*24473*/;
  assign _4519_ = inv_10[56] & r_9[56] /*24472*/;
  assign _4520_ = _4518_ | _4519_ /*24471*/;
  assign _4521_ = inv_10[57] ^ r_9[57] /*24469*/;
  assign sum_10[57] = _4521_ ^ _4520_ /*24468*/;
  assign _4522_ = _4521_ & _4520_ /*24467*/;
  assign _4523_ = inv_10[57] & r_9[57] /*24466*/;
  assign _4524_ = _4522_ | _4523_ /*24465*/;
  assign _4525_ = inv_10[58] ^ r_9[58] /*24463*/;
  assign sum_10[58] = _4525_ ^ _4524_ /*24462*/;
  assign _4526_ = _4525_ & _4524_ /*24461*/;
  assign _4527_ = inv_10[58] & r_9[58] /*24460*/;
  assign _4528_ = _4526_ | _4527_ /*24459*/;
  assign _4529_ = inv_10[59] ^ r_9[59] /*24457*/;
  assign sum_10[59] = _4529_ ^ _4528_ /*24456*/;
  assign _4530_ = _4529_ & _4528_ /*24455*/;
  assign _4531_ = inv_10[59] & r_9[59] /*24454*/;
  assign _4532_ = _4530_ | _4531_ /*24453*/;
  assign _4533_ = inv_10[60] ^ r_9[60] /*24451*/;
  assign sum_10[60] = _4533_ ^ _4532_ /*24450*/;
  assign _4534_ = _4533_ & _4532_ /*24449*/;
  assign _4535_ = inv_10[60] & r_9[60] /*24448*/;
  assign _4536_ = _4534_ | _4535_ /*24447*/;
  assign _4537_ = inv_10[61] ^ r_9[61] /*24445*/;
  assign sum_10[61] = _4537_ ^ _4536_ /*24444*/;
  assign _4538_ = _4537_ & _4536_ /*24443*/;
  assign _4539_ = inv_10[61] & r_9[61] /*24442*/;
  assign _4540_ = _4538_ | _4539_ /*24441*/;
  assign _4541_ = inv_10[62] ^ r_9[62] /*24439*/;
  assign sum_10[62] = _4541_ ^ _4540_ /*24438*/;
  assign _4542_ = _4541_ & _4540_ /*24437*/;
  assign _4543_ = inv_10[62] & r_9[62] /*24436*/;
  assign _4544_ = _4542_ | _4543_ /*24435*/;
  assign _4545_ = inv_10[63] ^ r_9[63] /*24433*/;
  assign sum_10[63] = _4545_ ^ _4544_ /*24432*/;
  assign _4546_ = _4545_ & _4544_ /*24431*/;
  assign _4547_ = inv_10[63] & r_9[63] /*24430*/;
  assign _4548_ = _4546_ | _4547_ /*24429*/;
  assign _4549_ = inv_10[64] ^ r_9[64] /*24427*/;
  assign sum_10[64] = _4549_ ^ _4548_ /*24426*/;
  assign _4550_ = _4549_ & _4548_ /*24425*/;
  assign _4551_ = inv_10[64] & r_9[64] /*24424*/;
  assign _4552_ = _4550_ | _4551_ /*24423*/;
  assign _4553_ = inv_10[65] ^ r_9[65] /*24421*/;
  assign sum_10[65] = _4553_ ^ _4552_ /*24420*/;
  assign _4554_ = _4553_ & _4552_ /*24419*/;
  assign _4555_ = inv_10[65] & r_9[65] /*24418*/;
  assign _4556_ = _4554_ | _4555_ /*24417*/;
  assign _4557_ = inv_10[66] ^ r_9[66] /*24415*/;
  assign sum_10[66] = _4557_ ^ _4556_ /*24414*/;
  assign _4558_ = _4557_ & _4556_ /*24413*/;
  assign _4559_ = inv_10[66] & r_9[66] /*24412*/;
  assign _4560_ = _4558_ | _4559_ /*24411*/;
  assign _4561_ = inv_10[67] ^ r_9[67] /*24409*/;
  assign sum_10[67] = _4561_ ^ _4560_ /*24408*/;
  assign _4562_ = _4561_ & _4560_ /*24407*/;
  assign _4563_ = inv_10[67] & r_9[67] /*24406*/;
  assign _4564_ = _4562_ | _4563_ /*24405*/;
  assign _4565_ = inv_10[68] ^ r_9[68] /*24403*/;
  assign sum_10[68] = _4565_ ^ _4564_ /*24402*/;
  assign _4566_ = _4565_ & _4564_ /*24401*/;
  assign _4567_ = inv_10[68] & r_9[68] /*24400*/;
  assign _4568_ = _4566_ | _4567_ /*24399*/;
  assign _4569_ = inv_10[69] ^ r_9[69] /*24397*/;
  assign sum_10[69] = _4569_ ^ _4568_ /*24396*/;
  assign _4570_ = _4569_ & _4568_ /*24395*/;
  assign _4571_ = inv_10[69] & r_9[69] /*24394*/;
  assign _4572_ = _4570_ | _4571_ /*24393*/;
  assign _4573_ = inv_10[70] ^ r_9[70] /*24391*/;
  assign sum_10[70] = _4573_ ^ _4572_ /*24390*/;
  assign _4574_ = _4573_ & _4572_ /*24389*/;
  assign _4575_ = inv_10[70] & r_9[70] /*24388*/;
  assign _4576_ = _4574_ | _4575_ /*24387*/;
  assign _4577_ = inv_10[71] ^ r_9[71] /*24385*/;
  assign sum_10[71] = _4577_ ^ _4576_ /*24384*/;
  assign _4578_ = _4577_ & _4576_ /*24383*/;
  assign _4579_ = inv_10[71] & r_9[71] /*24382*/;
  assign _4580_ = _4578_ | _4579_ /*24381*/;
  assign _4581_ = _4580_ ^ _4576_ /*24380*/;
  assign _4582_ = ~_4581_ /*24379*/;
  assign _4583_ = sum_10[71] & _4582_ /*24378*/;
  assign _4584_ = _4581_ & _4580_ /*24377*/;
  assign sum_10[72] = _4584_ | _4583_ /*24376*/;
  assign q[22] = ~sum_10[72] /*24375*/;
  assign m_10[0] = r_9[0] /*24374*/;
  assign m_10[1] = r_9[1] /*24373*/;
  assign m_10[2] = r_9[2] /*24372*/;
  assign m_10[3] = r_9[3] /*24371*/;
  assign m_10[4] = r_9[4] /*24370*/;
  assign m_10[5] = r_9[5] /*24369*/;
  assign m_10[6] = r_9[6] /*24368*/;
  assign m_10[7] = r_9[7] /*24367*/;
  assign m_10[8] = r_9[8] /*24366*/;
  assign m_10[9] = r_9[9] /*24365*/;
  assign m_10[10] = r_9[10] /*24364*/;
  assign m_10[11] = r_9[11] /*24363*/;
  assign m_10[12] = r_9[12] /*24362*/;
  assign m_10[13] = r_9[13] /*24361*/;
  assign m_10[14] = r_9[14] /*24360*/;
  assign m_10[15] = r_9[15] /*24359*/;
  assign m_10[16] = r_9[16] /*24358*/;
  assign m_10[17] = r_9[17] /*24357*/;
  assign m_10[18] = r_9[18] /*24356*/;
  assign m_10[19] = r_9[19] /*24355*/;
  assign m_10[20] = r_9[20] /*24354*/;
  assign m_10[21] = r_9[21] /*24353*/;
  assign m_10[22] = r_9[22] /*24352*/;
  assign m_10[23] = r_9[23] /*24351*/;
  assign m_10[24] = r_9[24] /*24350*/;
  assign m_10[25] = r_9[25] /*24349*/;
  assign m_10[26] = r_9[26] /*24348*/;
  assign m_10[27] = r_9[27] /*24347*/;
  assign m_10[28] = r_9[28] /*24346*/;
  assign m_10[29] = r_9[29] /*24345*/;
  assign m_10[30] = r_9[30] /*24344*/;
  assign m_10[31] = r_9[31] /*24343*/;
  assign m_10[32] = r_9[32] /*24342*/;
  assign m_10[33] = r_9[33] /*24341*/;
  assign m_10[34] = r_9[34] /*24340*/;
  assign m_10[35] = r_9[35] /*24339*/;
  assign m_10[36] = r_9[36] /*24338*/;
  assign m_10[37] = r_9[37] /*24337*/;
  assign m_10[38] = r_9[38] /*24336*/;
  assign m_10[39] = r_9[39] /*24335*/;
  assign m_10[40] = r_9[40] /*24334*/;
  assign m_10[41] = r_9[41] /*24333*/;
  assign m_10[42] = r_9[42] /*24332*/;
  assign m_10[43] = r_9[43] /*24331*/;
  assign m_10[44] = r_9[44] /*24330*/;
  assign m_10[45] = r_9[45] /*24329*/;
  assign m_10[46] = r_9[46] /*24328*/;
  assign m_10[47] = r_9[47] /*24327*/;
  assign m_10[48] = r_9[48] /*24326*/;
  assign m_10[49] = r_9[49] /*24325*/;
  assign m_10[50] = r_9[50] /*24324*/;
  assign m_10[51] = r_9[51] /*24323*/;
  assign m_10[52] = r_9[52] /*24322*/;
  assign m_10[53] = r_9[53] /*24321*/;
  assign m_10[54] = r_9[54] /*24320*/;
  assign m_10[55] = r_9[55] /*24319*/;
  assign m_10[56] = r_9[56] /*24318*/;
  assign m_10[57] = r_9[57] /*24317*/;
  assign m_10[58] = r_9[58] /*24316*/;
  assign m_10[59] = r_9[59] /*24315*/;
  assign m_10[60] = r_9[60] /*24314*/;
  assign m_10[61] = r_9[61] /*24313*/;
  assign m_10[62] = r_9[62] /*24312*/;
  assign m_10[63] = r_9[63] /*24311*/;
  assign m_10[64] = r_9[64] /*24310*/;
  assign m_10[65] = r_9[65] /*24309*/;
  assign m_10[66] = r_9[66] /*24308*/;
  assign m_10[67] = r_9[67] /*24307*/;
  assign m_10[68] = r_9[68] /*24306*/;
  assign m_10[69] = r_9[69] /*24305*/;
  assign m_10[70] = r_9[70] /*24304*/;
  assign m_10[71] = r_9[71] /*24303*/;
  assign m_10[72] = r_9[71] /*24302*/;
  assign _4586_ = ~q[22] /*24301*/;
  assign _4587_ = sum_10[0] & q[22] /*24300*/;
  assign _4588_ = m_10[0] & _4586_ /*24299*/;
  assign r_10[0] = _4588_ | _4587_ /*24298*/;
  assign _4589_ = ~q[22] /*24297*/;
  assign _4590_ = sum_10[1] & q[22] /*24296*/;
  assign _4591_ = m_10[1] & _4589_ /*24295*/;
  assign r_10[1] = _4591_ | _4590_ /*24294*/;
  assign _4592_ = ~q[22] /*24293*/;
  assign _4593_ = sum_10[2] & q[22] /*24292*/;
  assign _4594_ = m_10[2] & _4592_ /*24291*/;
  assign r_10[2] = _4594_ | _4593_ /*24290*/;
  assign _4595_ = ~q[22] /*24289*/;
  assign _4596_ = sum_10[3] & q[22] /*24288*/;
  assign _4597_ = m_10[3] & _4595_ /*24287*/;
  assign r_10[3] = _4597_ | _4596_ /*24286*/;
  assign _4598_ = ~q[22] /*24285*/;
  assign _4599_ = sum_10[4] & q[22] /*24284*/;
  assign _4600_ = m_10[4] & _4598_ /*24283*/;
  assign r_10[4] = _4600_ | _4599_ /*24282*/;
  assign _4601_ = ~q[22] /*24281*/;
  assign _4602_ = sum_10[5] & q[22] /*24280*/;
  assign _4603_ = m_10[5] & _4601_ /*24279*/;
  assign r_10[5] = _4603_ | _4602_ /*24278*/;
  assign _4604_ = ~q[22] /*24277*/;
  assign _4605_ = sum_10[6] & q[22] /*24276*/;
  assign _4606_ = m_10[6] & _4604_ /*24275*/;
  assign r_10[6] = _4606_ | _4605_ /*24274*/;
  assign _4607_ = ~q[22] /*24273*/;
  assign _4608_ = sum_10[7] & q[22] /*24272*/;
  assign _4609_ = m_10[7] & _4607_ /*24271*/;
  assign r_10[7] = _4609_ | _4608_ /*24270*/;
  assign _4610_ = ~q[22] /*24269*/;
  assign _4611_ = sum_10[8] & q[22] /*24268*/;
  assign _4612_ = m_10[8] & _4610_ /*24267*/;
  assign r_10[8] = _4612_ | _4611_ /*24266*/;
  assign _4613_ = ~q[22] /*24265*/;
  assign _4614_ = sum_10[9] & q[22] /*24264*/;
  assign _4615_ = m_10[9] & _4613_ /*24263*/;
  assign r_10[9] = _4615_ | _4614_ /*24262*/;
  assign _4616_ = ~q[22] /*24261*/;
  assign _4617_ = sum_10[10] & q[22] /*24260*/;
  assign _4618_ = m_10[10] & _4616_ /*24259*/;
  assign r_10[10] = _4618_ | _4617_ /*24258*/;
  assign _4619_ = ~q[22] /*24257*/;
  assign _4620_ = sum_10[11] & q[22] /*24256*/;
  assign _4621_ = m_10[11] & _4619_ /*24255*/;
  assign r_10[11] = _4621_ | _4620_ /*24254*/;
  assign _4622_ = ~q[22] /*24253*/;
  assign _4623_ = sum_10[12] & q[22] /*24252*/;
  assign _4624_ = m_10[12] & _4622_ /*24251*/;
  assign r_10[12] = _4624_ | _4623_ /*24250*/;
  assign _4625_ = ~q[22] /*24249*/;
  assign _4626_ = sum_10[13] & q[22] /*24248*/;
  assign _4627_ = m_10[13] & _4625_ /*24247*/;
  assign r_10[13] = _4627_ | _4626_ /*24246*/;
  assign _4628_ = ~q[22] /*24245*/;
  assign _4629_ = sum_10[14] & q[22] /*24244*/;
  assign _4630_ = m_10[14] & _4628_ /*24243*/;
  assign r_10[14] = _4630_ | _4629_ /*24242*/;
  assign _4631_ = ~q[22] /*24241*/;
  assign _4632_ = sum_10[15] & q[22] /*24240*/;
  assign _4633_ = m_10[15] & _4631_ /*24239*/;
  assign r_10[15] = _4633_ | _4632_ /*24238*/;
  assign _4634_ = ~q[22] /*24237*/;
  assign _4635_ = sum_10[16] & q[22] /*24236*/;
  assign _4636_ = m_10[16] & _4634_ /*24235*/;
  assign r_10[16] = _4636_ | _4635_ /*24234*/;
  assign _4637_ = ~q[22] /*24233*/;
  assign _4638_ = sum_10[17] & q[22] /*24232*/;
  assign _4639_ = m_10[17] & _4637_ /*24231*/;
  assign r_10[17] = _4639_ | _4638_ /*24230*/;
  assign _4640_ = ~q[22] /*24229*/;
  assign _4641_ = sum_10[18] & q[22] /*24228*/;
  assign _4642_ = m_10[18] & _4640_ /*24227*/;
  assign r_10[18] = _4642_ | _4641_ /*24226*/;
  assign _4643_ = ~q[22] /*24225*/;
  assign _4644_ = sum_10[19] & q[22] /*24224*/;
  assign _4645_ = m_10[19] & _4643_ /*24223*/;
  assign r_10[19] = _4645_ | _4644_ /*24222*/;
  assign _4646_ = ~q[22] /*24221*/;
  assign _4647_ = sum_10[20] & q[22] /*24220*/;
  assign _4648_ = m_10[20] & _4646_ /*24219*/;
  assign r_10[20] = _4648_ | _4647_ /*24218*/;
  assign _4649_ = ~q[22] /*24217*/;
  assign _4650_ = sum_10[21] & q[22] /*24216*/;
  assign _4651_ = m_10[21] & _4649_ /*24215*/;
  assign r_10[21] = _4651_ | _4650_ /*24214*/;
  assign _4652_ = ~q[22] /*24213*/;
  assign _4653_ = sum_10[22] & q[22] /*24212*/;
  assign _4654_ = m_10[22] & _4652_ /*24211*/;
  assign r_10[22] = _4654_ | _4653_ /*24210*/;
  assign _4655_ = ~q[22] /*24209*/;
  assign _4656_ = sum_10[23] & q[22] /*24208*/;
  assign _4657_ = m_10[23] & _4655_ /*24207*/;
  assign r_10[23] = _4657_ | _4656_ /*24206*/;
  assign _4658_ = ~q[22] /*24205*/;
  assign _4659_ = sum_10[24] & q[22] /*24204*/;
  assign _4660_ = m_10[24] & _4658_ /*24203*/;
  assign r_10[24] = _4660_ | _4659_ /*24202*/;
  assign _4661_ = ~q[22] /*24201*/;
  assign _4662_ = sum_10[25] & q[22] /*24200*/;
  assign _4663_ = m_10[25] & _4661_ /*24199*/;
  assign r_10[25] = _4663_ | _4662_ /*24198*/;
  assign _4664_ = ~q[22] /*24197*/;
  assign _4665_ = sum_10[26] & q[22] /*24196*/;
  assign _4666_ = m_10[26] & _4664_ /*24195*/;
  assign r_10[26] = _4666_ | _4665_ /*24194*/;
  assign _4667_ = ~q[22] /*24193*/;
  assign _4668_ = sum_10[27] & q[22] /*24192*/;
  assign _4669_ = m_10[27] & _4667_ /*24191*/;
  assign r_10[27] = _4669_ | _4668_ /*24190*/;
  assign _4670_ = ~q[22] /*24189*/;
  assign _4671_ = sum_10[28] & q[22] /*24188*/;
  assign _4672_ = m_10[28] & _4670_ /*24187*/;
  assign r_10[28] = _4672_ | _4671_ /*24186*/;
  assign _4673_ = ~q[22] /*24185*/;
  assign _4674_ = sum_10[29] & q[22] /*24184*/;
  assign _4675_ = m_10[29] & _4673_ /*24183*/;
  assign r_10[29] = _4675_ | _4674_ /*24182*/;
  assign _4676_ = ~q[22] /*24181*/;
  assign _4677_ = sum_10[30] & q[22] /*24180*/;
  assign _4678_ = m_10[30] & _4676_ /*24179*/;
  assign r_10[30] = _4678_ | _4677_ /*24178*/;
  assign _4679_ = ~q[22] /*24177*/;
  assign _4680_ = sum_10[31] & q[22] /*24176*/;
  assign _4681_ = m_10[31] & _4679_ /*24175*/;
  assign r_10[31] = _4681_ | _4680_ /*24174*/;
  assign _4682_ = ~q[22] /*24173*/;
  assign _4683_ = sum_10[32] & q[22] /*24172*/;
  assign _4684_ = m_10[32] & _4682_ /*24171*/;
  assign r_10[32] = _4684_ | _4683_ /*24170*/;
  assign _4685_ = ~q[22] /*24169*/;
  assign _4686_ = sum_10[33] & q[22] /*24168*/;
  assign _4687_ = m_10[33] & _4685_ /*24167*/;
  assign r_10[33] = _4687_ | _4686_ /*24166*/;
  assign _4688_ = ~q[22] /*24165*/;
  assign _4689_ = sum_10[34] & q[22] /*24164*/;
  assign _4690_ = m_10[34] & _4688_ /*24163*/;
  assign r_10[34] = _4690_ | _4689_ /*24162*/;
  assign _4691_ = ~q[22] /*24161*/;
  assign _4692_ = sum_10[35] & q[22] /*24160*/;
  assign _4693_ = m_10[35] & _4691_ /*24159*/;
  assign r_10[35] = _4693_ | _4692_ /*24158*/;
  assign _4694_ = ~q[22] /*24157*/;
  assign _4695_ = sum_10[36] & q[22] /*24156*/;
  assign _4696_ = m_10[36] & _4694_ /*24155*/;
  assign r_10[36] = _4696_ | _4695_ /*24154*/;
  assign _4697_ = ~q[22] /*24153*/;
  assign _4698_ = sum_10[37] & q[22] /*24152*/;
  assign _4699_ = m_10[37] & _4697_ /*24151*/;
  assign r_10[37] = _4699_ | _4698_ /*24150*/;
  assign _4700_ = ~q[22] /*24149*/;
  assign _4701_ = sum_10[38] & q[22] /*24148*/;
  assign _4702_ = m_10[38] & _4700_ /*24147*/;
  assign r_10[38] = _4702_ | _4701_ /*24146*/;
  assign _4703_ = ~q[22] /*24145*/;
  assign _4704_ = sum_10[39] & q[22] /*24144*/;
  assign _4705_ = m_10[39] & _4703_ /*24143*/;
  assign r_10[39] = _4705_ | _4704_ /*24142*/;
  assign _4706_ = ~q[22] /*24141*/;
  assign _4707_ = sum_10[40] & q[22] /*24140*/;
  assign _4708_ = m_10[40] & _4706_ /*24139*/;
  assign r_10[40] = _4708_ | _4707_ /*24138*/;
  assign _4709_ = ~q[22] /*24137*/;
  assign _4710_ = sum_10[41] & q[22] /*24136*/;
  assign _4711_ = m_10[41] & _4709_ /*24135*/;
  assign r_10[41] = _4711_ | _4710_ /*24134*/;
  assign _4712_ = ~q[22] /*24133*/;
  assign _4713_ = sum_10[42] & q[22] /*24132*/;
  assign _4714_ = m_10[42] & _4712_ /*24131*/;
  assign r_10[42] = _4714_ | _4713_ /*24130*/;
  assign _4715_ = ~q[22] /*24129*/;
  assign _4716_ = sum_10[43] & q[22] /*24128*/;
  assign _4717_ = m_10[43] & _4715_ /*24127*/;
  assign r_10[43] = _4717_ | _4716_ /*24126*/;
  assign _4718_ = ~q[22] /*24125*/;
  assign _4719_ = sum_10[44] & q[22] /*24124*/;
  assign _4720_ = m_10[44] & _4718_ /*24123*/;
  assign r_10[44] = _4720_ | _4719_ /*24122*/;
  assign _4721_ = ~q[22] /*24121*/;
  assign _4722_ = sum_10[45] & q[22] /*24120*/;
  assign _4723_ = m_10[45] & _4721_ /*24119*/;
  assign r_10[45] = _4723_ | _4722_ /*24118*/;
  assign _4724_ = ~q[22] /*24117*/;
  assign _4725_ = sum_10[46] & q[22] /*24116*/;
  assign _4726_ = m_10[46] & _4724_ /*24115*/;
  assign r_10[46] = _4726_ | _4725_ /*24114*/;
  assign _4727_ = ~q[22] /*24113*/;
  assign _4728_ = sum_10[47] & q[22] /*24112*/;
  assign _4729_ = m_10[47] & _4727_ /*24111*/;
  assign r_10[47] = _4729_ | _4728_ /*24110*/;
  assign _4730_ = ~q[22] /*24109*/;
  assign _4731_ = sum_10[48] & q[22] /*24108*/;
  assign _4732_ = m_10[48] & _4730_ /*24107*/;
  assign r_10[48] = _4732_ | _4731_ /*24106*/;
  assign _4733_ = ~q[22] /*24105*/;
  assign _4734_ = sum_10[49] & q[22] /*24104*/;
  assign _4735_ = m_10[49] & _4733_ /*24103*/;
  assign r_10[49] = _4735_ | _4734_ /*24102*/;
  assign _4736_ = ~q[22] /*24101*/;
  assign _4737_ = sum_10[50] & q[22] /*24100*/;
  assign _4738_ = m_10[50] & _4736_ /*24099*/;
  assign r_10[50] = _4738_ | _4737_ /*24098*/;
  assign _4739_ = ~q[22] /*24097*/;
  assign _4740_ = sum_10[51] & q[22] /*24096*/;
  assign _4741_ = m_10[51] & _4739_ /*24095*/;
  assign r_10[51] = _4741_ | _4740_ /*24094*/;
  assign _4742_ = ~q[22] /*24093*/;
  assign _4743_ = sum_10[52] & q[22] /*24092*/;
  assign _4744_ = m_10[52] & _4742_ /*24091*/;
  assign r_10[52] = _4744_ | _4743_ /*24090*/;
  assign _4745_ = ~q[22] /*24089*/;
  assign _4746_ = sum_10[53] & q[22] /*24088*/;
  assign _4747_ = m_10[53] & _4745_ /*24087*/;
  assign r_10[53] = _4747_ | _4746_ /*24086*/;
  assign _4748_ = ~q[22] /*24085*/;
  assign _4749_ = sum_10[54] & q[22] /*24084*/;
  assign _4750_ = m_10[54] & _4748_ /*24083*/;
  assign r_10[54] = _4750_ | _4749_ /*24082*/;
  assign _4751_ = ~q[22] /*24081*/;
  assign _4752_ = sum_10[55] & q[22] /*24080*/;
  assign _4753_ = m_10[55] & _4751_ /*24079*/;
  assign r_10[55] = _4753_ | _4752_ /*24078*/;
  assign _4754_ = ~q[22] /*24077*/;
  assign _4755_ = sum_10[56] & q[22] /*24076*/;
  assign _4756_ = m_10[56] & _4754_ /*24075*/;
  assign r_10[56] = _4756_ | _4755_ /*24074*/;
  assign _4757_ = ~q[22] /*24073*/;
  assign _4758_ = sum_10[57] & q[22] /*24072*/;
  assign _4759_ = m_10[57] & _4757_ /*24071*/;
  assign r_10[57] = _4759_ | _4758_ /*24070*/;
  assign _4760_ = ~q[22] /*24069*/;
  assign _4761_ = sum_10[58] & q[22] /*24068*/;
  assign _4762_ = m_10[58] & _4760_ /*24067*/;
  assign r_10[58] = _4762_ | _4761_ /*24066*/;
  assign _4763_ = ~q[22] /*24065*/;
  assign _4764_ = sum_10[59] & q[22] /*24064*/;
  assign _4765_ = m_10[59] & _4763_ /*24063*/;
  assign r_10[59] = _4765_ | _4764_ /*24062*/;
  assign _4766_ = ~q[22] /*24061*/;
  assign _4767_ = sum_10[60] & q[22] /*24060*/;
  assign _4768_ = m_10[60] & _4766_ /*24059*/;
  assign r_10[60] = _4768_ | _4767_ /*24058*/;
  assign _4769_ = ~q[22] /*24057*/;
  assign _4770_ = sum_10[61] & q[22] /*24056*/;
  assign _4771_ = m_10[61] & _4769_ /*24055*/;
  assign r_10[61] = _4771_ | _4770_ /*24054*/;
  assign _4772_ = ~q[22] /*24053*/;
  assign _4773_ = sum_10[62] & q[22] /*24052*/;
  assign _4774_ = m_10[62] & _4772_ /*24051*/;
  assign r_10[62] = _4774_ | _4773_ /*24050*/;
  assign _4775_ = ~q[22] /*24049*/;
  assign _4776_ = sum_10[63] & q[22] /*24048*/;
  assign _4777_ = m_10[63] & _4775_ /*24047*/;
  assign r_10[63] = _4777_ | _4776_ /*24046*/;
  assign _4778_ = ~q[22] /*24045*/;
  assign _4779_ = sum_10[64] & q[22] /*24044*/;
  assign _4780_ = m_10[64] & _4778_ /*24043*/;
  assign r_10[64] = _4780_ | _4779_ /*24042*/;
  assign _4781_ = ~q[22] /*24041*/;
  assign _4782_ = sum_10[65] & q[22] /*24040*/;
  assign _4783_ = m_10[65] & _4781_ /*24039*/;
  assign r_10[65] = _4783_ | _4782_ /*24038*/;
  assign _4784_ = ~q[22] /*24037*/;
  assign _4785_ = sum_10[66] & q[22] /*24036*/;
  assign _4786_ = m_10[66] & _4784_ /*24035*/;
  assign r_10[66] = _4786_ | _4785_ /*24034*/;
  assign _4787_ = ~q[22] /*24033*/;
  assign _4788_ = sum_10[67] & q[22] /*24032*/;
  assign _4789_ = m_10[67] & _4787_ /*24031*/;
  assign r_10[67] = _4789_ | _4788_ /*24030*/;
  assign _4790_ = ~q[22] /*24029*/;
  assign _4791_ = sum_10[68] & q[22] /*24028*/;
  assign _4792_ = m_10[68] & _4790_ /*24027*/;
  assign r_10[68] = _4792_ | _4791_ /*24026*/;
  assign _4793_ = ~q[22] /*24025*/;
  assign _4794_ = sum_10[69] & q[22] /*24024*/;
  assign _4795_ = m_10[69] & _4793_ /*24023*/;
  assign r_10[69] = _4795_ | _4794_ /*24022*/;
  assign _4796_ = ~q[22] /*24021*/;
  assign _4797_ = sum_10[70] & q[22] /*24020*/;
  assign _4798_ = m_10[70] & _4796_ /*24019*/;
  assign r_10[70] = _4798_ | _4797_ /*24018*/;
  assign _4799_ = ~q[22] /*24017*/;
  assign _4800_ = sum_10[71] & q[22] /*24016*/;
  assign _4801_ = m_10[71] & _4799_ /*24015*/;
  assign r_10[71] = _4801_ | _4800_ /*24014*/;
  assign _4802_ = ~q[22] /*24013*/;
  assign _4803_ = sum_10[72] & q[22] /*24012*/;
  assign _4804_ = m_10[72] & _4802_ /*24011*/;
  assign r_10[72] = _4804_ | _4803_ /*24010*/;
  assign inv_11[0] = oneWire /*23736*/;
  assign inv_11[1] = oneWire /*23730*/;
  assign inv_11[2] = oneWire /*23724*/;
  assign inv_11[3] = oneWire /*23718*/;
  assign inv_11[4] = oneWire /*23712*/;
  assign inv_11[5] = oneWire /*23706*/;
  assign inv_11[6] = oneWire /*23700*/;
  assign inv_11[7] = oneWire /*23694*/;
  assign inv_11[8] = oneWire /*23688*/;
  assign inv_11[9] = oneWire /*23682*/;
  assign inv_11[10] = oneWire /*23676*/;
  assign inv_11[11] = oneWire /*23670*/;
  assign inv_11[12] = oneWire /*23664*/;
  assign inv_11[13] = oneWire /*23658*/;
  assign inv_11[14] = oneWire /*23652*/;
  assign inv_11[15] = oneWire /*23646*/;
  assign inv_11[16] = oneWire /*23640*/;
  assign inv_11[17] = oneWire /*23634*/;
  assign inv_11[18] = oneWire /*23628*/;
  assign inv_11[19] = oneWire /*23622*/;
  assign inv_11[20] = oneWire /*23616*/;
  assign inv_11[21] = ~div[0] /*23610*/;
  assign inv_11[22] = ~div[1] /*23604*/;
  assign inv_11[23] = ~div[2] /*23598*/;
  assign inv_11[24] = ~div[3] /*23592*/;
  assign inv_11[25] = ~div[4] /*23586*/;
  assign inv_11[26] = ~div[5] /*23580*/;
  assign inv_11[27] = ~div[6] /*23574*/;
  assign inv_11[28] = ~div[7] /*23568*/;
  assign inv_11[29] = ~div[8] /*23562*/;
  assign inv_11[30] = ~div[9] /*23556*/;
  assign inv_11[31] = ~div[10] /*23550*/;
  assign inv_11[32] = ~div[11] /*23544*/;
  assign inv_11[33] = ~div[12] /*23538*/;
  assign inv_11[34] = ~div[13] /*23532*/;
  assign inv_11[35] = ~div[14] /*23526*/;
  assign inv_11[36] = ~div[15] /*23520*/;
  assign inv_11[37] = ~div[16] /*23514*/;
  assign inv_11[38] = ~div[17] /*23508*/;
  assign inv_11[39] = ~div[18] /*23502*/;
  assign inv_11[40] = ~div[19] /*23496*/;
  assign inv_11[41] = ~div[20] /*23490*/;
  assign inv_11[42] = ~div[21] /*23484*/;
  assign inv_11[43] = ~div[22] /*23478*/;
  assign inv_11[44] = ~div[23] /*23472*/;
  assign inv_11[45] = ~div[24] /*23466*/;
  assign inv_11[46] = ~div[25] /*23460*/;
  assign inv_11[47] = ~div[26] /*23454*/;
  assign inv_11[48] = ~div[27] /*23448*/;
  assign inv_11[49] = ~div[28] /*23442*/;
  assign inv_11[50] = ~div[29] /*23436*/;
  assign inv_11[51] = ~div[30] /*23430*/;
  assign inv_11[52] = oneWire /*23424*/;
  assign inv_11[53] = oneWire /*23418*/;
  assign inv_11[54] = oneWire /*23412*/;
  assign inv_11[55] = oneWire /*23406*/;
  assign inv_11[56] = oneWire /*23400*/;
  assign inv_11[57] = oneWire /*23394*/;
  assign inv_11[58] = oneWire /*23388*/;
  assign inv_11[59] = oneWire /*23382*/;
  assign inv_11[60] = oneWire /*23376*/;
  assign inv_11[61] = oneWire /*23370*/;
  assign inv_11[62] = oneWire /*23364*/;
  assign inv_11[63] = oneWire /*23358*/;
  assign inv_11[64] = oneWire /*23352*/;
  assign inv_11[65] = oneWire /*23346*/;
  assign inv_11[66] = oneWire /*23340*/;
  assign inv_11[67] = oneWire /*23334*/;
  assign inv_11[68] = oneWire /*23328*/;
  assign inv_11[69] = oneWire /*23322*/;
  assign inv_11[70] = oneWire /*23316*/;
  assign inv_11[71] = oneWire /*23310*/;
  assign inv_11[72] = oneWire /*23304*/;
  assign _4805_ = inv_11[0] ^ r_10[0] /*23735*/;
  assign sum_11[0] = _4805_ ^ oneWire /*23734*/;
  assign _4806_ = _4805_ & oneWire /*23733*/;
  assign _4807_ = inv_11[0] & r_10[0] /*23732*/;
  assign _4808_ = _4806_ | _4807_ /*23731*/;
  assign _4809_ = inv_11[1] ^ r_10[1] /*23729*/;
  assign sum_11[1] = _4809_ ^ _4808_ /*23728*/;
  assign _4810_ = _4809_ & _4808_ /*23727*/;
  assign _4811_ = inv_11[1] & r_10[1] /*23726*/;
  assign _4812_ = _4810_ | _4811_ /*23725*/;
  assign _4813_ = inv_11[2] ^ r_10[2] /*23723*/;
  assign sum_11[2] = _4813_ ^ _4812_ /*23722*/;
  assign _4814_ = _4813_ & _4812_ /*23721*/;
  assign _4815_ = inv_11[2] & r_10[2] /*23720*/;
  assign _4816_ = _4814_ | _4815_ /*23719*/;
  assign _4817_ = inv_11[3] ^ r_10[3] /*23717*/;
  assign sum_11[3] = _4817_ ^ _4816_ /*23716*/;
  assign _4818_ = _4817_ & _4816_ /*23715*/;
  assign _4819_ = inv_11[3] & r_10[3] /*23714*/;
  assign _4820_ = _4818_ | _4819_ /*23713*/;
  assign _4821_ = inv_11[4] ^ r_10[4] /*23711*/;
  assign sum_11[4] = _4821_ ^ _4820_ /*23710*/;
  assign _4822_ = _4821_ & _4820_ /*23709*/;
  assign _4823_ = inv_11[4] & r_10[4] /*23708*/;
  assign _4824_ = _4822_ | _4823_ /*23707*/;
  assign _4825_ = inv_11[5] ^ r_10[5] /*23705*/;
  assign sum_11[5] = _4825_ ^ _4824_ /*23704*/;
  assign _4826_ = _4825_ & _4824_ /*23703*/;
  assign _4827_ = inv_11[5] & r_10[5] /*23702*/;
  assign _4828_ = _4826_ | _4827_ /*23701*/;
  assign _4829_ = inv_11[6] ^ r_10[6] /*23699*/;
  assign sum_11[6] = _4829_ ^ _4828_ /*23698*/;
  assign _4830_ = _4829_ & _4828_ /*23697*/;
  assign _4831_ = inv_11[6] & r_10[6] /*23696*/;
  assign _4832_ = _4830_ | _4831_ /*23695*/;
  assign _4833_ = inv_11[7] ^ r_10[7] /*23693*/;
  assign sum_11[7] = _4833_ ^ _4832_ /*23692*/;
  assign _4834_ = _4833_ & _4832_ /*23691*/;
  assign _4835_ = inv_11[7] & r_10[7] /*23690*/;
  assign _4836_ = _4834_ | _4835_ /*23689*/;
  assign _4837_ = inv_11[8] ^ r_10[8] /*23687*/;
  assign sum_11[8] = _4837_ ^ _4836_ /*23686*/;
  assign _4838_ = _4837_ & _4836_ /*23685*/;
  assign _4839_ = inv_11[8] & r_10[8] /*23684*/;
  assign _4840_ = _4838_ | _4839_ /*23683*/;
  assign _4841_ = inv_11[9] ^ r_10[9] /*23681*/;
  assign sum_11[9] = _4841_ ^ _4840_ /*23680*/;
  assign _4842_ = _4841_ & _4840_ /*23679*/;
  assign _4843_ = inv_11[9] & r_10[9] /*23678*/;
  assign _4844_ = _4842_ | _4843_ /*23677*/;
  assign _4845_ = inv_11[10] ^ r_10[10] /*23675*/;
  assign sum_11[10] = _4845_ ^ _4844_ /*23674*/;
  assign _4846_ = _4845_ & _4844_ /*23673*/;
  assign _4847_ = inv_11[10] & r_10[10] /*23672*/;
  assign _4848_ = _4846_ | _4847_ /*23671*/;
  assign _4849_ = inv_11[11] ^ r_10[11] /*23669*/;
  assign sum_11[11] = _4849_ ^ _4848_ /*23668*/;
  assign _4850_ = _4849_ & _4848_ /*23667*/;
  assign _4851_ = inv_11[11] & r_10[11] /*23666*/;
  assign _4852_ = _4850_ | _4851_ /*23665*/;
  assign _4853_ = inv_11[12] ^ r_10[12] /*23663*/;
  assign sum_11[12] = _4853_ ^ _4852_ /*23662*/;
  assign _4854_ = _4853_ & _4852_ /*23661*/;
  assign _4855_ = inv_11[12] & r_10[12] /*23660*/;
  assign _4856_ = _4854_ | _4855_ /*23659*/;
  assign _4857_ = inv_11[13] ^ r_10[13] /*23657*/;
  assign sum_11[13] = _4857_ ^ _4856_ /*23656*/;
  assign _4858_ = _4857_ & _4856_ /*23655*/;
  assign _4859_ = inv_11[13] & r_10[13] /*23654*/;
  assign _4860_ = _4858_ | _4859_ /*23653*/;
  assign _4861_ = inv_11[14] ^ r_10[14] /*23651*/;
  assign sum_11[14] = _4861_ ^ _4860_ /*23650*/;
  assign _4862_ = _4861_ & _4860_ /*23649*/;
  assign _4863_ = inv_11[14] & r_10[14] /*23648*/;
  assign _4864_ = _4862_ | _4863_ /*23647*/;
  assign _4865_ = inv_11[15] ^ r_10[15] /*23645*/;
  assign sum_11[15] = _4865_ ^ _4864_ /*23644*/;
  assign _4866_ = _4865_ & _4864_ /*23643*/;
  assign _4867_ = inv_11[15] & r_10[15] /*23642*/;
  assign _4868_ = _4866_ | _4867_ /*23641*/;
  assign _4869_ = inv_11[16] ^ r_10[16] /*23639*/;
  assign sum_11[16] = _4869_ ^ _4868_ /*23638*/;
  assign _4870_ = _4869_ & _4868_ /*23637*/;
  assign _4871_ = inv_11[16] & r_10[16] /*23636*/;
  assign _4872_ = _4870_ | _4871_ /*23635*/;
  assign _4873_ = inv_11[17] ^ r_10[17] /*23633*/;
  assign sum_11[17] = _4873_ ^ _4872_ /*23632*/;
  assign _4874_ = _4873_ & _4872_ /*23631*/;
  assign _4875_ = inv_11[17] & r_10[17] /*23630*/;
  assign _4876_ = _4874_ | _4875_ /*23629*/;
  assign _4877_ = inv_11[18] ^ r_10[18] /*23627*/;
  assign sum_11[18] = _4877_ ^ _4876_ /*23626*/;
  assign _4878_ = _4877_ & _4876_ /*23625*/;
  assign _4879_ = inv_11[18] & r_10[18] /*23624*/;
  assign _4880_ = _4878_ | _4879_ /*23623*/;
  assign _4881_ = inv_11[19] ^ r_10[19] /*23621*/;
  assign sum_11[19] = _4881_ ^ _4880_ /*23620*/;
  assign _4882_ = _4881_ & _4880_ /*23619*/;
  assign _4883_ = inv_11[19] & r_10[19] /*23618*/;
  assign _4884_ = _4882_ | _4883_ /*23617*/;
  assign _4885_ = inv_11[20] ^ r_10[20] /*23615*/;
  assign sum_11[20] = _4885_ ^ _4884_ /*23614*/;
  assign _4886_ = _4885_ & _4884_ /*23613*/;
  assign _4887_ = inv_11[20] & r_10[20] /*23612*/;
  assign _4888_ = _4886_ | _4887_ /*23611*/;
  assign _4889_ = inv_11[21] ^ r_10[21] /*23609*/;
  assign sum_11[21] = _4889_ ^ _4888_ /*23608*/;
  assign _4890_ = _4889_ & _4888_ /*23607*/;
  assign _4891_ = inv_11[21] & r_10[21] /*23606*/;
  assign _4892_ = _4890_ | _4891_ /*23605*/;
  assign _4893_ = inv_11[22] ^ r_10[22] /*23603*/;
  assign sum_11[22] = _4893_ ^ _4892_ /*23602*/;
  assign _4894_ = _4893_ & _4892_ /*23601*/;
  assign _4895_ = inv_11[22] & r_10[22] /*23600*/;
  assign _4896_ = _4894_ | _4895_ /*23599*/;
  assign _4897_ = inv_11[23] ^ r_10[23] /*23597*/;
  assign sum_11[23] = _4897_ ^ _4896_ /*23596*/;
  assign _4898_ = _4897_ & _4896_ /*23595*/;
  assign _4899_ = inv_11[23] & r_10[23] /*23594*/;
  assign _4900_ = _4898_ | _4899_ /*23593*/;
  assign _4901_ = inv_11[24] ^ r_10[24] /*23591*/;
  assign sum_11[24] = _4901_ ^ _4900_ /*23590*/;
  assign _4902_ = _4901_ & _4900_ /*23589*/;
  assign _4903_ = inv_11[24] & r_10[24] /*23588*/;
  assign _4904_ = _4902_ | _4903_ /*23587*/;
  assign _4905_ = inv_11[25] ^ r_10[25] /*23585*/;
  assign sum_11[25] = _4905_ ^ _4904_ /*23584*/;
  assign _4906_ = _4905_ & _4904_ /*23583*/;
  assign _4907_ = inv_11[25] & r_10[25] /*23582*/;
  assign _4908_ = _4906_ | _4907_ /*23581*/;
  assign _4909_ = inv_11[26] ^ r_10[26] /*23579*/;
  assign sum_11[26] = _4909_ ^ _4908_ /*23578*/;
  assign _4910_ = _4909_ & _4908_ /*23577*/;
  assign _4911_ = inv_11[26] & r_10[26] /*23576*/;
  assign _4912_ = _4910_ | _4911_ /*23575*/;
  assign _4913_ = inv_11[27] ^ r_10[27] /*23573*/;
  assign sum_11[27] = _4913_ ^ _4912_ /*23572*/;
  assign _4914_ = _4913_ & _4912_ /*23571*/;
  assign _4915_ = inv_11[27] & r_10[27] /*23570*/;
  assign _4916_ = _4914_ | _4915_ /*23569*/;
  assign _4917_ = inv_11[28] ^ r_10[28] /*23567*/;
  assign sum_11[28] = _4917_ ^ _4916_ /*23566*/;
  assign _4918_ = _4917_ & _4916_ /*23565*/;
  assign _4919_ = inv_11[28] & r_10[28] /*23564*/;
  assign _4920_ = _4918_ | _4919_ /*23563*/;
  assign _4921_ = inv_11[29] ^ r_10[29] /*23561*/;
  assign sum_11[29] = _4921_ ^ _4920_ /*23560*/;
  assign _4922_ = _4921_ & _4920_ /*23559*/;
  assign _4923_ = inv_11[29] & r_10[29] /*23558*/;
  assign _4924_ = _4922_ | _4923_ /*23557*/;
  assign _4925_ = inv_11[30] ^ r_10[30] /*23555*/;
  assign sum_11[30] = _4925_ ^ _4924_ /*23554*/;
  assign _4926_ = _4925_ & _4924_ /*23553*/;
  assign _4927_ = inv_11[30] & r_10[30] /*23552*/;
  assign _4928_ = _4926_ | _4927_ /*23551*/;
  assign _4929_ = inv_11[31] ^ r_10[31] /*23549*/;
  assign sum_11[31] = _4929_ ^ _4928_ /*23548*/;
  assign _4930_ = _4929_ & _4928_ /*23547*/;
  assign _4931_ = inv_11[31] & r_10[31] /*23546*/;
  assign _4932_ = _4930_ | _4931_ /*23545*/;
  assign _4933_ = inv_11[32] ^ r_10[32] /*23543*/;
  assign sum_11[32] = _4933_ ^ _4932_ /*23542*/;
  assign _4934_ = _4933_ & _4932_ /*23541*/;
  assign _4935_ = inv_11[32] & r_10[32] /*23540*/;
  assign _4936_ = _4934_ | _4935_ /*23539*/;
  assign _4937_ = inv_11[33] ^ r_10[33] /*23537*/;
  assign sum_11[33] = _4937_ ^ _4936_ /*23536*/;
  assign _4938_ = _4937_ & _4936_ /*23535*/;
  assign _4939_ = inv_11[33] & r_10[33] /*23534*/;
  assign _4940_ = _4938_ | _4939_ /*23533*/;
  assign _4941_ = inv_11[34] ^ r_10[34] /*23531*/;
  assign sum_11[34] = _4941_ ^ _4940_ /*23530*/;
  assign _4942_ = _4941_ & _4940_ /*23529*/;
  assign _4943_ = inv_11[34] & r_10[34] /*23528*/;
  assign _4944_ = _4942_ | _4943_ /*23527*/;
  assign _4945_ = inv_11[35] ^ r_10[35] /*23525*/;
  assign sum_11[35] = _4945_ ^ _4944_ /*23524*/;
  assign _4946_ = _4945_ & _4944_ /*23523*/;
  assign _4947_ = inv_11[35] & r_10[35] /*23522*/;
  assign _4948_ = _4946_ | _4947_ /*23521*/;
  assign _4949_ = inv_11[36] ^ r_10[36] /*23519*/;
  assign sum_11[36] = _4949_ ^ _4948_ /*23518*/;
  assign _4950_ = _4949_ & _4948_ /*23517*/;
  assign _4951_ = inv_11[36] & r_10[36] /*23516*/;
  assign _4952_ = _4950_ | _4951_ /*23515*/;
  assign _4953_ = inv_11[37] ^ r_10[37] /*23513*/;
  assign sum_11[37] = _4953_ ^ _4952_ /*23512*/;
  assign _4954_ = _4953_ & _4952_ /*23511*/;
  assign _4955_ = inv_11[37] & r_10[37] /*23510*/;
  assign _4956_ = _4954_ | _4955_ /*23509*/;
  assign _4957_ = inv_11[38] ^ r_10[38] /*23507*/;
  assign sum_11[38] = _4957_ ^ _4956_ /*23506*/;
  assign _4958_ = _4957_ & _4956_ /*23505*/;
  assign _4959_ = inv_11[38] & r_10[38] /*23504*/;
  assign _4960_ = _4958_ | _4959_ /*23503*/;
  assign _4961_ = inv_11[39] ^ r_10[39] /*23501*/;
  assign sum_11[39] = _4961_ ^ _4960_ /*23500*/;
  assign _4962_ = _4961_ & _4960_ /*23499*/;
  assign _4963_ = inv_11[39] & r_10[39] /*23498*/;
  assign _4964_ = _4962_ | _4963_ /*23497*/;
  assign _4965_ = inv_11[40] ^ r_10[40] /*23495*/;
  assign sum_11[40] = _4965_ ^ _4964_ /*23494*/;
  assign _4966_ = _4965_ & _4964_ /*23493*/;
  assign _4967_ = inv_11[40] & r_10[40] /*23492*/;
  assign _4968_ = _4966_ | _4967_ /*23491*/;
  assign _4969_ = inv_11[41] ^ r_10[41] /*23489*/;
  assign sum_11[41] = _4969_ ^ _4968_ /*23488*/;
  assign _4970_ = _4969_ & _4968_ /*23487*/;
  assign _4971_ = inv_11[41] & r_10[41] /*23486*/;
  assign _4972_ = _4970_ | _4971_ /*23485*/;
  assign _4973_ = inv_11[42] ^ r_10[42] /*23483*/;
  assign sum_11[42] = _4973_ ^ _4972_ /*23482*/;
  assign _4974_ = _4973_ & _4972_ /*23481*/;
  assign _4975_ = inv_11[42] & r_10[42] /*23480*/;
  assign _4976_ = _4974_ | _4975_ /*23479*/;
  assign _4977_ = inv_11[43] ^ r_10[43] /*23477*/;
  assign sum_11[43] = _4977_ ^ _4976_ /*23476*/;
  assign _4978_ = _4977_ & _4976_ /*23475*/;
  assign _4979_ = inv_11[43] & r_10[43] /*23474*/;
  assign _4980_ = _4978_ | _4979_ /*23473*/;
  assign _4981_ = inv_11[44] ^ r_10[44] /*23471*/;
  assign sum_11[44] = _4981_ ^ _4980_ /*23470*/;
  assign _4982_ = _4981_ & _4980_ /*23469*/;
  assign _4983_ = inv_11[44] & r_10[44] /*23468*/;
  assign _4984_ = _4982_ | _4983_ /*23467*/;
  assign _4985_ = inv_11[45] ^ r_10[45] /*23465*/;
  assign sum_11[45] = _4985_ ^ _4984_ /*23464*/;
  assign _4986_ = _4985_ & _4984_ /*23463*/;
  assign _4987_ = inv_11[45] & r_10[45] /*23462*/;
  assign _4988_ = _4986_ | _4987_ /*23461*/;
  assign _4989_ = inv_11[46] ^ r_10[46] /*23459*/;
  assign sum_11[46] = _4989_ ^ _4988_ /*23458*/;
  assign _4990_ = _4989_ & _4988_ /*23457*/;
  assign _4991_ = inv_11[46] & r_10[46] /*23456*/;
  assign _4992_ = _4990_ | _4991_ /*23455*/;
  assign _4993_ = inv_11[47] ^ r_10[47] /*23453*/;
  assign sum_11[47] = _4993_ ^ _4992_ /*23452*/;
  assign _4994_ = _4993_ & _4992_ /*23451*/;
  assign _4995_ = inv_11[47] & r_10[47] /*23450*/;
  assign _4996_ = _4994_ | _4995_ /*23449*/;
  assign _4997_ = inv_11[48] ^ r_10[48] /*23447*/;
  assign sum_11[48] = _4997_ ^ _4996_ /*23446*/;
  assign _4998_ = _4997_ & _4996_ /*23445*/;
  assign _4999_ = inv_11[48] & r_10[48] /*23444*/;
  assign _5000_ = _4998_ | _4999_ /*23443*/;
  assign _5001_ = inv_11[49] ^ r_10[49] /*23441*/;
  assign sum_11[49] = _5001_ ^ _5000_ /*23440*/;
  assign _5002_ = _5001_ & _5000_ /*23439*/;
  assign _5003_ = inv_11[49] & r_10[49] /*23438*/;
  assign _5004_ = _5002_ | _5003_ /*23437*/;
  assign _5005_ = inv_11[50] ^ r_10[50] /*23435*/;
  assign sum_11[50] = _5005_ ^ _5004_ /*23434*/;
  assign _5006_ = _5005_ & _5004_ /*23433*/;
  assign _5007_ = inv_11[50] & r_10[50] /*23432*/;
  assign _5008_ = _5006_ | _5007_ /*23431*/;
  assign _5009_ = inv_11[51] ^ r_10[51] /*23429*/;
  assign sum_11[51] = _5009_ ^ _5008_ /*23428*/;
  assign _5010_ = _5009_ & _5008_ /*23427*/;
  assign _5011_ = inv_11[51] & r_10[51] /*23426*/;
  assign _5012_ = _5010_ | _5011_ /*23425*/;
  assign _5013_ = inv_11[52] ^ r_10[52] /*23423*/;
  assign sum_11[52] = _5013_ ^ _5012_ /*23422*/;
  assign _5014_ = _5013_ & _5012_ /*23421*/;
  assign _5015_ = inv_11[52] & r_10[52] /*23420*/;
  assign _5016_ = _5014_ | _5015_ /*23419*/;
  assign _5017_ = inv_11[53] ^ r_10[53] /*23417*/;
  assign sum_11[53] = _5017_ ^ _5016_ /*23416*/;
  assign _5018_ = _5017_ & _5016_ /*23415*/;
  assign _5019_ = inv_11[53] & r_10[53] /*23414*/;
  assign _5020_ = _5018_ | _5019_ /*23413*/;
  assign _5021_ = inv_11[54] ^ r_10[54] /*23411*/;
  assign sum_11[54] = _5021_ ^ _5020_ /*23410*/;
  assign _5022_ = _5021_ & _5020_ /*23409*/;
  assign _5023_ = inv_11[54] & r_10[54] /*23408*/;
  assign _5024_ = _5022_ | _5023_ /*23407*/;
  assign _5025_ = inv_11[55] ^ r_10[55] /*23405*/;
  assign sum_11[55] = _5025_ ^ _5024_ /*23404*/;
  assign _5026_ = _5025_ & _5024_ /*23403*/;
  assign _5027_ = inv_11[55] & r_10[55] /*23402*/;
  assign _5028_ = _5026_ | _5027_ /*23401*/;
  assign _5029_ = inv_11[56] ^ r_10[56] /*23399*/;
  assign sum_11[56] = _5029_ ^ _5028_ /*23398*/;
  assign _5030_ = _5029_ & _5028_ /*23397*/;
  assign _5031_ = inv_11[56] & r_10[56] /*23396*/;
  assign _5032_ = _5030_ | _5031_ /*23395*/;
  assign _5033_ = inv_11[57] ^ r_10[57] /*23393*/;
  assign sum_11[57] = _5033_ ^ _5032_ /*23392*/;
  assign _5034_ = _5033_ & _5032_ /*23391*/;
  assign _5035_ = inv_11[57] & r_10[57] /*23390*/;
  assign _5036_ = _5034_ | _5035_ /*23389*/;
  assign _5037_ = inv_11[58] ^ r_10[58] /*23387*/;
  assign sum_11[58] = _5037_ ^ _5036_ /*23386*/;
  assign _5038_ = _5037_ & _5036_ /*23385*/;
  assign _5039_ = inv_11[58] & r_10[58] /*23384*/;
  assign _5040_ = _5038_ | _5039_ /*23383*/;
  assign _5041_ = inv_11[59] ^ r_10[59] /*23381*/;
  assign sum_11[59] = _5041_ ^ _5040_ /*23380*/;
  assign _5042_ = _5041_ & _5040_ /*23379*/;
  assign _5043_ = inv_11[59] & r_10[59] /*23378*/;
  assign _5044_ = _5042_ | _5043_ /*23377*/;
  assign _5045_ = inv_11[60] ^ r_10[60] /*23375*/;
  assign sum_11[60] = _5045_ ^ _5044_ /*23374*/;
  assign _5046_ = _5045_ & _5044_ /*23373*/;
  assign _5047_ = inv_11[60] & r_10[60] /*23372*/;
  assign _5048_ = _5046_ | _5047_ /*23371*/;
  assign _5049_ = inv_11[61] ^ r_10[61] /*23369*/;
  assign sum_11[61] = _5049_ ^ _5048_ /*23368*/;
  assign _5050_ = _5049_ & _5048_ /*23367*/;
  assign _5051_ = inv_11[61] & r_10[61] /*23366*/;
  assign _5052_ = _5050_ | _5051_ /*23365*/;
  assign _5053_ = inv_11[62] ^ r_10[62] /*23363*/;
  assign sum_11[62] = _5053_ ^ _5052_ /*23362*/;
  assign _5054_ = _5053_ & _5052_ /*23361*/;
  assign _5055_ = inv_11[62] & r_10[62] /*23360*/;
  assign _5056_ = _5054_ | _5055_ /*23359*/;
  assign _5057_ = inv_11[63] ^ r_10[63] /*23357*/;
  assign sum_11[63] = _5057_ ^ _5056_ /*23356*/;
  assign _5058_ = _5057_ & _5056_ /*23355*/;
  assign _5059_ = inv_11[63] & r_10[63] /*23354*/;
  assign _5060_ = _5058_ | _5059_ /*23353*/;
  assign _5061_ = inv_11[64] ^ r_10[64] /*23351*/;
  assign sum_11[64] = _5061_ ^ _5060_ /*23350*/;
  assign _5062_ = _5061_ & _5060_ /*23349*/;
  assign _5063_ = inv_11[64] & r_10[64] /*23348*/;
  assign _5064_ = _5062_ | _5063_ /*23347*/;
  assign _5065_ = inv_11[65] ^ r_10[65] /*23345*/;
  assign sum_11[65] = _5065_ ^ _5064_ /*23344*/;
  assign _5066_ = _5065_ & _5064_ /*23343*/;
  assign _5067_ = inv_11[65] & r_10[65] /*23342*/;
  assign _5068_ = _5066_ | _5067_ /*23341*/;
  assign _5069_ = inv_11[66] ^ r_10[66] /*23339*/;
  assign sum_11[66] = _5069_ ^ _5068_ /*23338*/;
  assign _5070_ = _5069_ & _5068_ /*23337*/;
  assign _5071_ = inv_11[66] & r_10[66] /*23336*/;
  assign _5072_ = _5070_ | _5071_ /*23335*/;
  assign _5073_ = inv_11[67] ^ r_10[67] /*23333*/;
  assign sum_11[67] = _5073_ ^ _5072_ /*23332*/;
  assign _5074_ = _5073_ & _5072_ /*23331*/;
  assign _5075_ = inv_11[67] & r_10[67] /*23330*/;
  assign _5076_ = _5074_ | _5075_ /*23329*/;
  assign _5077_ = inv_11[68] ^ r_10[68] /*23327*/;
  assign sum_11[68] = _5077_ ^ _5076_ /*23326*/;
  assign _5078_ = _5077_ & _5076_ /*23325*/;
  assign _5079_ = inv_11[68] & r_10[68] /*23324*/;
  assign _5080_ = _5078_ | _5079_ /*23323*/;
  assign _5081_ = inv_11[69] ^ r_10[69] /*23321*/;
  assign sum_11[69] = _5081_ ^ _5080_ /*23320*/;
  assign _5082_ = _5081_ & _5080_ /*23319*/;
  assign _5083_ = inv_11[69] & r_10[69] /*23318*/;
  assign _5084_ = _5082_ | _5083_ /*23317*/;
  assign _5085_ = inv_11[70] ^ r_10[70] /*23315*/;
  assign sum_11[70] = _5085_ ^ _5084_ /*23314*/;
  assign _5086_ = _5085_ & _5084_ /*23313*/;
  assign _5087_ = inv_11[70] & r_10[70] /*23312*/;
  assign _5088_ = _5086_ | _5087_ /*23311*/;
  assign _5089_ = inv_11[71] ^ r_10[71] /*23309*/;
  assign sum_11[71] = _5089_ ^ _5088_ /*23308*/;
  assign _5090_ = _5089_ & _5088_ /*23307*/;
  assign _5091_ = inv_11[71] & r_10[71] /*23306*/;
  assign _5092_ = _5090_ | _5091_ /*23305*/;
  assign _5093_ = inv_11[72] ^ r_10[72] /*23303*/;
  assign sum_11[72] = _5093_ ^ _5092_ /*23302*/;
  assign _5094_ = _5093_ & _5092_ /*23301*/;
  assign _5095_ = inv_11[72] & r_10[72] /*23300*/;
  assign _5096_ = _5094_ | _5095_ /*23299*/;
  assign _5097_ = _5096_ ^ _5092_ /*23298*/;
  assign _5098_ = ~_5097_ /*23297*/;
  assign _5099_ = sum_11[72] & _5098_ /*23296*/;
  assign _5100_ = _5097_ & _5096_ /*23295*/;
  assign sum_11[73] = _5100_ | _5099_ /*23294*/;
  assign q[21] = ~sum_11[73] /*23293*/;
  assign m_11[0] = r_10[0] /*23292*/;
  assign m_11[1] = r_10[1] /*23291*/;
  assign m_11[2] = r_10[2] /*23290*/;
  assign m_11[3] = r_10[3] /*23289*/;
  assign m_11[4] = r_10[4] /*23288*/;
  assign m_11[5] = r_10[5] /*23287*/;
  assign m_11[6] = r_10[6] /*23286*/;
  assign m_11[7] = r_10[7] /*23285*/;
  assign m_11[8] = r_10[8] /*23284*/;
  assign m_11[9] = r_10[9] /*23283*/;
  assign m_11[10] = r_10[10] /*23282*/;
  assign m_11[11] = r_10[11] /*23281*/;
  assign m_11[12] = r_10[12] /*23280*/;
  assign m_11[13] = r_10[13] /*23279*/;
  assign m_11[14] = r_10[14] /*23278*/;
  assign m_11[15] = r_10[15] /*23277*/;
  assign m_11[16] = r_10[16] /*23276*/;
  assign m_11[17] = r_10[17] /*23275*/;
  assign m_11[18] = r_10[18] /*23274*/;
  assign m_11[19] = r_10[19] /*23273*/;
  assign m_11[20] = r_10[20] /*23272*/;
  assign m_11[21] = r_10[21] /*23271*/;
  assign m_11[22] = r_10[22] /*23270*/;
  assign m_11[23] = r_10[23] /*23269*/;
  assign m_11[24] = r_10[24] /*23268*/;
  assign m_11[25] = r_10[25] /*23267*/;
  assign m_11[26] = r_10[26] /*23266*/;
  assign m_11[27] = r_10[27] /*23265*/;
  assign m_11[28] = r_10[28] /*23264*/;
  assign m_11[29] = r_10[29] /*23263*/;
  assign m_11[30] = r_10[30] /*23262*/;
  assign m_11[31] = r_10[31] /*23261*/;
  assign m_11[32] = r_10[32] /*23260*/;
  assign m_11[33] = r_10[33] /*23259*/;
  assign m_11[34] = r_10[34] /*23258*/;
  assign m_11[35] = r_10[35] /*23257*/;
  assign m_11[36] = r_10[36] /*23256*/;
  assign m_11[37] = r_10[37] /*23255*/;
  assign m_11[38] = r_10[38] /*23254*/;
  assign m_11[39] = r_10[39] /*23253*/;
  assign m_11[40] = r_10[40] /*23252*/;
  assign m_11[41] = r_10[41] /*23251*/;
  assign m_11[42] = r_10[42] /*23250*/;
  assign m_11[43] = r_10[43] /*23249*/;
  assign m_11[44] = r_10[44] /*23248*/;
  assign m_11[45] = r_10[45] /*23247*/;
  assign m_11[46] = r_10[46] /*23246*/;
  assign m_11[47] = r_10[47] /*23245*/;
  assign m_11[48] = r_10[48] /*23244*/;
  assign m_11[49] = r_10[49] /*23243*/;
  assign m_11[50] = r_10[50] /*23242*/;
  assign m_11[51] = r_10[51] /*23241*/;
  assign m_11[52] = r_10[52] /*23240*/;
  assign m_11[53] = r_10[53] /*23239*/;
  assign m_11[54] = r_10[54] /*23238*/;
  assign m_11[55] = r_10[55] /*23237*/;
  assign m_11[56] = r_10[56] /*23236*/;
  assign m_11[57] = r_10[57] /*23235*/;
  assign m_11[58] = r_10[58] /*23234*/;
  assign m_11[59] = r_10[59] /*23233*/;
  assign m_11[60] = r_10[60] /*23232*/;
  assign m_11[61] = r_10[61] /*23231*/;
  assign m_11[62] = r_10[62] /*23230*/;
  assign m_11[63] = r_10[63] /*23229*/;
  assign m_11[64] = r_10[64] /*23228*/;
  assign m_11[65] = r_10[65] /*23227*/;
  assign m_11[66] = r_10[66] /*23226*/;
  assign m_11[67] = r_10[67] /*23225*/;
  assign m_11[68] = r_10[68] /*23224*/;
  assign m_11[69] = r_10[69] /*23223*/;
  assign m_11[70] = r_10[70] /*23222*/;
  assign m_11[71] = r_10[71] /*23221*/;
  assign m_11[72] = r_10[72] /*23220*/;
  assign m_11[73] = r_10[72] /*23219*/;
  assign _5102_ = ~q[21] /*23218*/;
  assign _5103_ = sum_11[0] & q[21] /*23217*/;
  assign _5104_ = m_11[0] & _5102_ /*23216*/;
  assign r_11[0] = _5104_ | _5103_ /*23215*/;
  assign _5105_ = ~q[21] /*23214*/;
  assign _5106_ = sum_11[1] & q[21] /*23213*/;
  assign _5107_ = m_11[1] & _5105_ /*23212*/;
  assign r_11[1] = _5107_ | _5106_ /*23211*/;
  assign _5108_ = ~q[21] /*23210*/;
  assign _5109_ = sum_11[2] & q[21] /*23209*/;
  assign _5110_ = m_11[2] & _5108_ /*23208*/;
  assign r_11[2] = _5110_ | _5109_ /*23207*/;
  assign _5111_ = ~q[21] /*23206*/;
  assign _5112_ = sum_11[3] & q[21] /*23205*/;
  assign _5113_ = m_11[3] & _5111_ /*23204*/;
  assign r_11[3] = _5113_ | _5112_ /*23203*/;
  assign _5114_ = ~q[21] /*23202*/;
  assign _5115_ = sum_11[4] & q[21] /*23201*/;
  assign _5116_ = m_11[4] & _5114_ /*23200*/;
  assign r_11[4] = _5116_ | _5115_ /*23199*/;
  assign _5117_ = ~q[21] /*23198*/;
  assign _5118_ = sum_11[5] & q[21] /*23197*/;
  assign _5119_ = m_11[5] & _5117_ /*23196*/;
  assign r_11[5] = _5119_ | _5118_ /*23195*/;
  assign _5120_ = ~q[21] /*23194*/;
  assign _5121_ = sum_11[6] & q[21] /*23193*/;
  assign _5122_ = m_11[6] & _5120_ /*23192*/;
  assign r_11[6] = _5122_ | _5121_ /*23191*/;
  assign _5123_ = ~q[21] /*23190*/;
  assign _5124_ = sum_11[7] & q[21] /*23189*/;
  assign _5125_ = m_11[7] & _5123_ /*23188*/;
  assign r_11[7] = _5125_ | _5124_ /*23187*/;
  assign _5126_ = ~q[21] /*23186*/;
  assign _5127_ = sum_11[8] & q[21] /*23185*/;
  assign _5128_ = m_11[8] & _5126_ /*23184*/;
  assign r_11[8] = _5128_ | _5127_ /*23183*/;
  assign _5129_ = ~q[21] /*23182*/;
  assign _5130_ = sum_11[9] & q[21] /*23181*/;
  assign _5131_ = m_11[9] & _5129_ /*23180*/;
  assign r_11[9] = _5131_ | _5130_ /*23179*/;
  assign _5132_ = ~q[21] /*23178*/;
  assign _5133_ = sum_11[10] & q[21] /*23177*/;
  assign _5134_ = m_11[10] & _5132_ /*23176*/;
  assign r_11[10] = _5134_ | _5133_ /*23175*/;
  assign _5135_ = ~q[21] /*23174*/;
  assign _5136_ = sum_11[11] & q[21] /*23173*/;
  assign _5137_ = m_11[11] & _5135_ /*23172*/;
  assign r_11[11] = _5137_ | _5136_ /*23171*/;
  assign _5138_ = ~q[21] /*23170*/;
  assign _5139_ = sum_11[12] & q[21] /*23169*/;
  assign _5140_ = m_11[12] & _5138_ /*23168*/;
  assign r_11[12] = _5140_ | _5139_ /*23167*/;
  assign _5141_ = ~q[21] /*23166*/;
  assign _5142_ = sum_11[13] & q[21] /*23165*/;
  assign _5143_ = m_11[13] & _5141_ /*23164*/;
  assign r_11[13] = _5143_ | _5142_ /*23163*/;
  assign _5144_ = ~q[21] /*23162*/;
  assign _5145_ = sum_11[14] & q[21] /*23161*/;
  assign _5146_ = m_11[14] & _5144_ /*23160*/;
  assign r_11[14] = _5146_ | _5145_ /*23159*/;
  assign _5147_ = ~q[21] /*23158*/;
  assign _5148_ = sum_11[15] & q[21] /*23157*/;
  assign _5149_ = m_11[15] & _5147_ /*23156*/;
  assign r_11[15] = _5149_ | _5148_ /*23155*/;
  assign _5150_ = ~q[21] /*23154*/;
  assign _5151_ = sum_11[16] & q[21] /*23153*/;
  assign _5152_ = m_11[16] & _5150_ /*23152*/;
  assign r_11[16] = _5152_ | _5151_ /*23151*/;
  assign _5153_ = ~q[21] /*23150*/;
  assign _5154_ = sum_11[17] & q[21] /*23149*/;
  assign _5155_ = m_11[17] & _5153_ /*23148*/;
  assign r_11[17] = _5155_ | _5154_ /*23147*/;
  assign _5156_ = ~q[21] /*23146*/;
  assign _5157_ = sum_11[18] & q[21] /*23145*/;
  assign _5158_ = m_11[18] & _5156_ /*23144*/;
  assign r_11[18] = _5158_ | _5157_ /*23143*/;
  assign _5159_ = ~q[21] /*23142*/;
  assign _5160_ = sum_11[19] & q[21] /*23141*/;
  assign _5161_ = m_11[19] & _5159_ /*23140*/;
  assign r_11[19] = _5161_ | _5160_ /*23139*/;
  assign _5162_ = ~q[21] /*23138*/;
  assign _5163_ = sum_11[20] & q[21] /*23137*/;
  assign _5164_ = m_11[20] & _5162_ /*23136*/;
  assign r_11[20] = _5164_ | _5163_ /*23135*/;
  assign _5165_ = ~q[21] /*23134*/;
  assign _5166_ = sum_11[21] & q[21] /*23133*/;
  assign _5167_ = m_11[21] & _5165_ /*23132*/;
  assign r_11[21] = _5167_ | _5166_ /*23131*/;
  assign _5168_ = ~q[21] /*23130*/;
  assign _5169_ = sum_11[22] & q[21] /*23129*/;
  assign _5170_ = m_11[22] & _5168_ /*23128*/;
  assign r_11[22] = _5170_ | _5169_ /*23127*/;
  assign _5171_ = ~q[21] /*23126*/;
  assign _5172_ = sum_11[23] & q[21] /*23125*/;
  assign _5173_ = m_11[23] & _5171_ /*23124*/;
  assign r_11[23] = _5173_ | _5172_ /*23123*/;
  assign _5174_ = ~q[21] /*23122*/;
  assign _5175_ = sum_11[24] & q[21] /*23121*/;
  assign _5176_ = m_11[24] & _5174_ /*23120*/;
  assign r_11[24] = _5176_ | _5175_ /*23119*/;
  assign _5177_ = ~q[21] /*23118*/;
  assign _5178_ = sum_11[25] & q[21] /*23117*/;
  assign _5179_ = m_11[25] & _5177_ /*23116*/;
  assign r_11[25] = _5179_ | _5178_ /*23115*/;
  assign _5180_ = ~q[21] /*23114*/;
  assign _5181_ = sum_11[26] & q[21] /*23113*/;
  assign _5182_ = m_11[26] & _5180_ /*23112*/;
  assign r_11[26] = _5182_ | _5181_ /*23111*/;
  assign _5183_ = ~q[21] /*23110*/;
  assign _5184_ = sum_11[27] & q[21] /*23109*/;
  assign _5185_ = m_11[27] & _5183_ /*23108*/;
  assign r_11[27] = _5185_ | _5184_ /*23107*/;
  assign _5186_ = ~q[21] /*23106*/;
  assign _5187_ = sum_11[28] & q[21] /*23105*/;
  assign _5188_ = m_11[28] & _5186_ /*23104*/;
  assign r_11[28] = _5188_ | _5187_ /*23103*/;
  assign _5189_ = ~q[21] /*23102*/;
  assign _5190_ = sum_11[29] & q[21] /*23101*/;
  assign _5191_ = m_11[29] & _5189_ /*23100*/;
  assign r_11[29] = _5191_ | _5190_ /*23099*/;
  assign _5192_ = ~q[21] /*23098*/;
  assign _5193_ = sum_11[30] & q[21] /*23097*/;
  assign _5194_ = m_11[30] & _5192_ /*23096*/;
  assign r_11[30] = _5194_ | _5193_ /*23095*/;
  assign _5195_ = ~q[21] /*23094*/;
  assign _5196_ = sum_11[31] & q[21] /*23093*/;
  assign _5197_ = m_11[31] & _5195_ /*23092*/;
  assign r_11[31] = _5197_ | _5196_ /*23091*/;
  assign _5198_ = ~q[21] /*23090*/;
  assign _5199_ = sum_11[32] & q[21] /*23089*/;
  assign _5200_ = m_11[32] & _5198_ /*23088*/;
  assign r_11[32] = _5200_ | _5199_ /*23087*/;
  assign _5201_ = ~q[21] /*23086*/;
  assign _5202_ = sum_11[33] & q[21] /*23085*/;
  assign _5203_ = m_11[33] & _5201_ /*23084*/;
  assign r_11[33] = _5203_ | _5202_ /*23083*/;
  assign _5204_ = ~q[21] /*23082*/;
  assign _5205_ = sum_11[34] & q[21] /*23081*/;
  assign _5206_ = m_11[34] & _5204_ /*23080*/;
  assign r_11[34] = _5206_ | _5205_ /*23079*/;
  assign _5207_ = ~q[21] /*23078*/;
  assign _5208_ = sum_11[35] & q[21] /*23077*/;
  assign _5209_ = m_11[35] & _5207_ /*23076*/;
  assign r_11[35] = _5209_ | _5208_ /*23075*/;
  assign _5210_ = ~q[21] /*23074*/;
  assign _5211_ = sum_11[36] & q[21] /*23073*/;
  assign _5212_ = m_11[36] & _5210_ /*23072*/;
  assign r_11[36] = _5212_ | _5211_ /*23071*/;
  assign _5213_ = ~q[21] /*23070*/;
  assign _5214_ = sum_11[37] & q[21] /*23069*/;
  assign _5215_ = m_11[37] & _5213_ /*23068*/;
  assign r_11[37] = _5215_ | _5214_ /*23067*/;
  assign _5216_ = ~q[21] /*23066*/;
  assign _5217_ = sum_11[38] & q[21] /*23065*/;
  assign _5218_ = m_11[38] & _5216_ /*23064*/;
  assign r_11[38] = _5218_ | _5217_ /*23063*/;
  assign _5219_ = ~q[21] /*23062*/;
  assign _5220_ = sum_11[39] & q[21] /*23061*/;
  assign _5221_ = m_11[39] & _5219_ /*23060*/;
  assign r_11[39] = _5221_ | _5220_ /*23059*/;
  assign _5222_ = ~q[21] /*23058*/;
  assign _5223_ = sum_11[40] & q[21] /*23057*/;
  assign _5224_ = m_11[40] & _5222_ /*23056*/;
  assign r_11[40] = _5224_ | _5223_ /*23055*/;
  assign _5225_ = ~q[21] /*23054*/;
  assign _5226_ = sum_11[41] & q[21] /*23053*/;
  assign _5227_ = m_11[41] & _5225_ /*23052*/;
  assign r_11[41] = _5227_ | _5226_ /*23051*/;
  assign _5228_ = ~q[21] /*23050*/;
  assign _5229_ = sum_11[42] & q[21] /*23049*/;
  assign _5230_ = m_11[42] & _5228_ /*23048*/;
  assign r_11[42] = _5230_ | _5229_ /*23047*/;
  assign _5231_ = ~q[21] /*23046*/;
  assign _5232_ = sum_11[43] & q[21] /*23045*/;
  assign _5233_ = m_11[43] & _5231_ /*23044*/;
  assign r_11[43] = _5233_ | _5232_ /*23043*/;
  assign _5234_ = ~q[21] /*23042*/;
  assign _5235_ = sum_11[44] & q[21] /*23041*/;
  assign _5236_ = m_11[44] & _5234_ /*23040*/;
  assign r_11[44] = _5236_ | _5235_ /*23039*/;
  assign _5237_ = ~q[21] /*23038*/;
  assign _5238_ = sum_11[45] & q[21] /*23037*/;
  assign _5239_ = m_11[45] & _5237_ /*23036*/;
  assign r_11[45] = _5239_ | _5238_ /*23035*/;
  assign _5240_ = ~q[21] /*23034*/;
  assign _5241_ = sum_11[46] & q[21] /*23033*/;
  assign _5242_ = m_11[46] & _5240_ /*23032*/;
  assign r_11[46] = _5242_ | _5241_ /*23031*/;
  assign _5243_ = ~q[21] /*23030*/;
  assign _5244_ = sum_11[47] & q[21] /*23029*/;
  assign _5245_ = m_11[47] & _5243_ /*23028*/;
  assign r_11[47] = _5245_ | _5244_ /*23027*/;
  assign _5246_ = ~q[21] /*23026*/;
  assign _5247_ = sum_11[48] & q[21] /*23025*/;
  assign _5248_ = m_11[48] & _5246_ /*23024*/;
  assign r_11[48] = _5248_ | _5247_ /*23023*/;
  assign _5249_ = ~q[21] /*23022*/;
  assign _5250_ = sum_11[49] & q[21] /*23021*/;
  assign _5251_ = m_11[49] & _5249_ /*23020*/;
  assign r_11[49] = _5251_ | _5250_ /*23019*/;
  assign _5252_ = ~q[21] /*23018*/;
  assign _5253_ = sum_11[50] & q[21] /*23017*/;
  assign _5254_ = m_11[50] & _5252_ /*23016*/;
  assign r_11[50] = _5254_ | _5253_ /*23015*/;
  assign _5255_ = ~q[21] /*23014*/;
  assign _5256_ = sum_11[51] & q[21] /*23013*/;
  assign _5257_ = m_11[51] & _5255_ /*23012*/;
  assign r_11[51] = _5257_ | _5256_ /*23011*/;
  assign _5258_ = ~q[21] /*23010*/;
  assign _5259_ = sum_11[52] & q[21] /*23009*/;
  assign _5260_ = m_11[52] & _5258_ /*23008*/;
  assign r_11[52] = _5260_ | _5259_ /*23007*/;
  assign _5261_ = ~q[21] /*23006*/;
  assign _5262_ = sum_11[53] & q[21] /*23005*/;
  assign _5263_ = m_11[53] & _5261_ /*23004*/;
  assign r_11[53] = _5263_ | _5262_ /*23003*/;
  assign _5264_ = ~q[21] /*23002*/;
  assign _5265_ = sum_11[54] & q[21] /*23001*/;
  assign _5266_ = m_11[54] & _5264_ /*23000*/;
  assign r_11[54] = _5266_ | _5265_ /*22999*/;
  assign _5267_ = ~q[21] /*22998*/;
  assign _5268_ = sum_11[55] & q[21] /*22997*/;
  assign _5269_ = m_11[55] & _5267_ /*22996*/;
  assign r_11[55] = _5269_ | _5268_ /*22995*/;
  assign _5270_ = ~q[21] /*22994*/;
  assign _5271_ = sum_11[56] & q[21] /*22993*/;
  assign _5272_ = m_11[56] & _5270_ /*22992*/;
  assign r_11[56] = _5272_ | _5271_ /*22991*/;
  assign _5273_ = ~q[21] /*22990*/;
  assign _5274_ = sum_11[57] & q[21] /*22989*/;
  assign _5275_ = m_11[57] & _5273_ /*22988*/;
  assign r_11[57] = _5275_ | _5274_ /*22987*/;
  assign _5276_ = ~q[21] /*22986*/;
  assign _5277_ = sum_11[58] & q[21] /*22985*/;
  assign _5278_ = m_11[58] & _5276_ /*22984*/;
  assign r_11[58] = _5278_ | _5277_ /*22983*/;
  assign _5279_ = ~q[21] /*22982*/;
  assign _5280_ = sum_11[59] & q[21] /*22981*/;
  assign _5281_ = m_11[59] & _5279_ /*22980*/;
  assign r_11[59] = _5281_ | _5280_ /*22979*/;
  assign _5282_ = ~q[21] /*22978*/;
  assign _5283_ = sum_11[60] & q[21] /*22977*/;
  assign _5284_ = m_11[60] & _5282_ /*22976*/;
  assign r_11[60] = _5284_ | _5283_ /*22975*/;
  assign _5285_ = ~q[21] /*22974*/;
  assign _5286_ = sum_11[61] & q[21] /*22973*/;
  assign _5287_ = m_11[61] & _5285_ /*22972*/;
  assign r_11[61] = _5287_ | _5286_ /*22971*/;
  assign _5288_ = ~q[21] /*22970*/;
  assign _5289_ = sum_11[62] & q[21] /*22969*/;
  assign _5290_ = m_11[62] & _5288_ /*22968*/;
  assign r_11[62] = _5290_ | _5289_ /*22967*/;
  assign _5291_ = ~q[21] /*22966*/;
  assign _5292_ = sum_11[63] & q[21] /*22965*/;
  assign _5293_ = m_11[63] & _5291_ /*22964*/;
  assign r_11[63] = _5293_ | _5292_ /*22963*/;
  assign _5294_ = ~q[21] /*22962*/;
  assign _5295_ = sum_11[64] & q[21] /*22961*/;
  assign _5296_ = m_11[64] & _5294_ /*22960*/;
  assign r_11[64] = _5296_ | _5295_ /*22959*/;
  assign _5297_ = ~q[21] /*22958*/;
  assign _5298_ = sum_11[65] & q[21] /*22957*/;
  assign _5299_ = m_11[65] & _5297_ /*22956*/;
  assign r_11[65] = _5299_ | _5298_ /*22955*/;
  assign _5300_ = ~q[21] /*22954*/;
  assign _5301_ = sum_11[66] & q[21] /*22953*/;
  assign _5302_ = m_11[66] & _5300_ /*22952*/;
  assign r_11[66] = _5302_ | _5301_ /*22951*/;
  assign _5303_ = ~q[21] /*22950*/;
  assign _5304_ = sum_11[67] & q[21] /*22949*/;
  assign _5305_ = m_11[67] & _5303_ /*22948*/;
  assign r_11[67] = _5305_ | _5304_ /*22947*/;
  assign _5306_ = ~q[21] /*22946*/;
  assign _5307_ = sum_11[68] & q[21] /*22945*/;
  assign _5308_ = m_11[68] & _5306_ /*22944*/;
  assign r_11[68] = _5308_ | _5307_ /*22943*/;
  assign _5309_ = ~q[21] /*22942*/;
  assign _5310_ = sum_11[69] & q[21] /*22941*/;
  assign _5311_ = m_11[69] & _5309_ /*22940*/;
  assign r_11[69] = _5311_ | _5310_ /*22939*/;
  assign _5312_ = ~q[21] /*22938*/;
  assign _5313_ = sum_11[70] & q[21] /*22937*/;
  assign _5314_ = m_11[70] & _5312_ /*22936*/;
  assign r_11[70] = _5314_ | _5313_ /*22935*/;
  assign _5315_ = ~q[21] /*22934*/;
  assign _5316_ = sum_11[71] & q[21] /*22933*/;
  assign _5317_ = m_11[71] & _5315_ /*22932*/;
  assign r_11[71] = _5317_ | _5316_ /*22931*/;
  assign _5318_ = ~q[21] /*22930*/;
  assign _5319_ = sum_11[72] & q[21] /*22929*/;
  assign _5320_ = m_11[72] & _5318_ /*22928*/;
  assign r_11[72] = _5320_ | _5319_ /*22927*/;
  assign _5321_ = ~q[21] /*22926*/;
  assign _5322_ = sum_11[73] & q[21] /*22925*/;
  assign _5323_ = m_11[73] & _5321_ /*22924*/;
  assign r_11[73] = _5323_ | _5322_ /*22923*/;
  assign inv_12[0] = oneWire /*22660*/;
  assign inv_12[1] = oneWire /*22654*/;
  assign inv_12[2] = oneWire /*22648*/;
  assign inv_12[3] = oneWire /*22642*/;
  assign inv_12[4] = oneWire /*22636*/;
  assign inv_12[5] = oneWire /*22630*/;
  assign inv_12[6] = oneWire /*22624*/;
  assign inv_12[7] = oneWire /*22618*/;
  assign inv_12[8] = oneWire /*22612*/;
  assign inv_12[9] = oneWire /*22606*/;
  assign inv_12[10] = oneWire /*22600*/;
  assign inv_12[11] = oneWire /*22594*/;
  assign inv_12[12] = oneWire /*22588*/;
  assign inv_12[13] = oneWire /*22582*/;
  assign inv_12[14] = oneWire /*22576*/;
  assign inv_12[15] = oneWire /*22570*/;
  assign inv_12[16] = oneWire /*22564*/;
  assign inv_12[17] = oneWire /*22558*/;
  assign inv_12[18] = oneWire /*22552*/;
  assign inv_12[19] = oneWire /*22546*/;
  assign inv_12[20] = ~div[0] /*22540*/;
  assign inv_12[21] = ~div[1] /*22534*/;
  assign inv_12[22] = ~div[2] /*22528*/;
  assign inv_12[23] = ~div[3] /*22522*/;
  assign inv_12[24] = ~div[4] /*22516*/;
  assign inv_12[25] = ~div[5] /*22510*/;
  assign inv_12[26] = ~div[6] /*22504*/;
  assign inv_12[27] = ~div[7] /*22498*/;
  assign inv_12[28] = ~div[8] /*22492*/;
  assign inv_12[29] = ~div[9] /*22486*/;
  assign inv_12[30] = ~div[10] /*22480*/;
  assign inv_12[31] = ~div[11] /*22474*/;
  assign inv_12[32] = ~div[12] /*22468*/;
  assign inv_12[33] = ~div[13] /*22462*/;
  assign inv_12[34] = ~div[14] /*22456*/;
  assign inv_12[35] = ~div[15] /*22450*/;
  assign inv_12[36] = ~div[16] /*22444*/;
  assign inv_12[37] = ~div[17] /*22438*/;
  assign inv_12[38] = ~div[18] /*22432*/;
  assign inv_12[39] = ~div[19] /*22426*/;
  assign inv_12[40] = ~div[20] /*22420*/;
  assign inv_12[41] = ~div[21] /*22414*/;
  assign inv_12[42] = ~div[22] /*22408*/;
  assign inv_12[43] = ~div[23] /*22402*/;
  assign inv_12[44] = ~div[24] /*22396*/;
  assign inv_12[45] = ~div[25] /*22390*/;
  assign inv_12[46] = ~div[26] /*22384*/;
  assign inv_12[47] = ~div[27] /*22378*/;
  assign inv_12[48] = ~div[28] /*22372*/;
  assign inv_12[49] = ~div[29] /*22366*/;
  assign inv_12[50] = ~div[30] /*22360*/;
  assign inv_12[51] = oneWire /*22354*/;
  assign inv_12[52] = oneWire /*22348*/;
  assign inv_12[53] = oneWire /*22342*/;
  assign inv_12[54] = oneWire /*22336*/;
  assign inv_12[55] = oneWire /*22330*/;
  assign inv_12[56] = oneWire /*22324*/;
  assign inv_12[57] = oneWire /*22318*/;
  assign inv_12[58] = oneWire /*22312*/;
  assign inv_12[59] = oneWire /*22306*/;
  assign inv_12[60] = oneWire /*22300*/;
  assign inv_12[61] = oneWire /*22294*/;
  assign inv_12[62] = oneWire /*22288*/;
  assign inv_12[63] = oneWire /*22282*/;
  assign inv_12[64] = oneWire /*22276*/;
  assign inv_12[65] = oneWire /*22270*/;
  assign inv_12[66] = oneWire /*22264*/;
  assign inv_12[67] = oneWire /*22258*/;
  assign inv_12[68] = oneWire /*22252*/;
  assign inv_12[69] = oneWire /*22246*/;
  assign inv_12[70] = oneWire /*22240*/;
  assign inv_12[71] = oneWire /*22234*/;
  assign inv_12[72] = oneWire /*22228*/;
  assign inv_12[73] = oneWire /*22222*/;
  assign _5324_ = inv_12[0] ^ r_11[0] /*22659*/;
  assign sum_12[0] = _5324_ ^ oneWire /*22658*/;
  assign _5325_ = _5324_ & oneWire /*22657*/;
  assign _5326_ = inv_12[0] & r_11[0] /*22656*/;
  assign _5327_ = _5325_ | _5326_ /*22655*/;
  assign _5328_ = inv_12[1] ^ r_11[1] /*22653*/;
  assign sum_12[1] = _5328_ ^ _5327_ /*22652*/;
  assign _5329_ = _5328_ & _5327_ /*22651*/;
  assign _5330_ = inv_12[1] & r_11[1] /*22650*/;
  assign _5331_ = _5329_ | _5330_ /*22649*/;
  assign _5332_ = inv_12[2] ^ r_11[2] /*22647*/;
  assign sum_12[2] = _5332_ ^ _5331_ /*22646*/;
  assign _5333_ = _5332_ & _5331_ /*22645*/;
  assign _5334_ = inv_12[2] & r_11[2] /*22644*/;
  assign _5335_ = _5333_ | _5334_ /*22643*/;
  assign _5336_ = inv_12[3] ^ r_11[3] /*22641*/;
  assign sum_12[3] = _5336_ ^ _5335_ /*22640*/;
  assign _5337_ = _5336_ & _5335_ /*22639*/;
  assign _5338_ = inv_12[3] & r_11[3] /*22638*/;
  assign _5339_ = _5337_ | _5338_ /*22637*/;
  assign _5340_ = inv_12[4] ^ r_11[4] /*22635*/;
  assign sum_12[4] = _5340_ ^ _5339_ /*22634*/;
  assign _5341_ = _5340_ & _5339_ /*22633*/;
  assign _5342_ = inv_12[4] & r_11[4] /*22632*/;
  assign _5343_ = _5341_ | _5342_ /*22631*/;
  assign _5344_ = inv_12[5] ^ r_11[5] /*22629*/;
  assign sum_12[5] = _5344_ ^ _5343_ /*22628*/;
  assign _5345_ = _5344_ & _5343_ /*22627*/;
  assign _5346_ = inv_12[5] & r_11[5] /*22626*/;
  assign _5347_ = _5345_ | _5346_ /*22625*/;
  assign _5348_ = inv_12[6] ^ r_11[6] /*22623*/;
  assign sum_12[6] = _5348_ ^ _5347_ /*22622*/;
  assign _5349_ = _5348_ & _5347_ /*22621*/;
  assign _5350_ = inv_12[6] & r_11[6] /*22620*/;
  assign _5351_ = _5349_ | _5350_ /*22619*/;
  assign _5352_ = inv_12[7] ^ r_11[7] /*22617*/;
  assign sum_12[7] = _5352_ ^ _5351_ /*22616*/;
  assign _5353_ = _5352_ & _5351_ /*22615*/;
  assign _5354_ = inv_12[7] & r_11[7] /*22614*/;
  assign _5355_ = _5353_ | _5354_ /*22613*/;
  assign _5356_ = inv_12[8] ^ r_11[8] /*22611*/;
  assign sum_12[8] = _5356_ ^ _5355_ /*22610*/;
  assign _5357_ = _5356_ & _5355_ /*22609*/;
  assign _5358_ = inv_12[8] & r_11[8] /*22608*/;
  assign _5359_ = _5357_ | _5358_ /*22607*/;
  assign _5360_ = inv_12[9] ^ r_11[9] /*22605*/;
  assign sum_12[9] = _5360_ ^ _5359_ /*22604*/;
  assign _5361_ = _5360_ & _5359_ /*22603*/;
  assign _5362_ = inv_12[9] & r_11[9] /*22602*/;
  assign _5363_ = _5361_ | _5362_ /*22601*/;
  assign _5364_ = inv_12[10] ^ r_11[10] /*22599*/;
  assign sum_12[10] = _5364_ ^ _5363_ /*22598*/;
  assign _5365_ = _5364_ & _5363_ /*22597*/;
  assign _5366_ = inv_12[10] & r_11[10] /*22596*/;
  assign _5367_ = _5365_ | _5366_ /*22595*/;
  assign _5368_ = inv_12[11] ^ r_11[11] /*22593*/;
  assign sum_12[11] = _5368_ ^ _5367_ /*22592*/;
  assign _5369_ = _5368_ & _5367_ /*22591*/;
  assign _5370_ = inv_12[11] & r_11[11] /*22590*/;
  assign _5371_ = _5369_ | _5370_ /*22589*/;
  assign _5372_ = inv_12[12] ^ r_11[12] /*22587*/;
  assign sum_12[12] = _5372_ ^ _5371_ /*22586*/;
  assign _5373_ = _5372_ & _5371_ /*22585*/;
  assign _5374_ = inv_12[12] & r_11[12] /*22584*/;
  assign _5375_ = _5373_ | _5374_ /*22583*/;
  assign _5376_ = inv_12[13] ^ r_11[13] /*22581*/;
  assign sum_12[13] = _5376_ ^ _5375_ /*22580*/;
  assign _5377_ = _5376_ & _5375_ /*22579*/;
  assign _5378_ = inv_12[13] & r_11[13] /*22578*/;
  assign _5379_ = _5377_ | _5378_ /*22577*/;
  assign _5380_ = inv_12[14] ^ r_11[14] /*22575*/;
  assign sum_12[14] = _5380_ ^ _5379_ /*22574*/;
  assign _5381_ = _5380_ & _5379_ /*22573*/;
  assign _5382_ = inv_12[14] & r_11[14] /*22572*/;
  assign _5383_ = _5381_ | _5382_ /*22571*/;
  assign _5384_ = inv_12[15] ^ r_11[15] /*22569*/;
  assign sum_12[15] = _5384_ ^ _5383_ /*22568*/;
  assign _5385_ = _5384_ & _5383_ /*22567*/;
  assign _5386_ = inv_12[15] & r_11[15] /*22566*/;
  assign _5387_ = _5385_ | _5386_ /*22565*/;
  assign _5388_ = inv_12[16] ^ r_11[16] /*22563*/;
  assign sum_12[16] = _5388_ ^ _5387_ /*22562*/;
  assign _5389_ = _5388_ & _5387_ /*22561*/;
  assign _5390_ = inv_12[16] & r_11[16] /*22560*/;
  assign _5391_ = _5389_ | _5390_ /*22559*/;
  assign _5392_ = inv_12[17] ^ r_11[17] /*22557*/;
  assign sum_12[17] = _5392_ ^ _5391_ /*22556*/;
  assign _5393_ = _5392_ & _5391_ /*22555*/;
  assign _5394_ = inv_12[17] & r_11[17] /*22554*/;
  assign _5395_ = _5393_ | _5394_ /*22553*/;
  assign _5396_ = inv_12[18] ^ r_11[18] /*22551*/;
  assign sum_12[18] = _5396_ ^ _5395_ /*22550*/;
  assign _5397_ = _5396_ & _5395_ /*22549*/;
  assign _5398_ = inv_12[18] & r_11[18] /*22548*/;
  assign _5399_ = _5397_ | _5398_ /*22547*/;
  assign _5400_ = inv_12[19] ^ r_11[19] /*22545*/;
  assign sum_12[19] = _5400_ ^ _5399_ /*22544*/;
  assign _5401_ = _5400_ & _5399_ /*22543*/;
  assign _5402_ = inv_12[19] & r_11[19] /*22542*/;
  assign _5403_ = _5401_ | _5402_ /*22541*/;
  assign _5404_ = inv_12[20] ^ r_11[20] /*22539*/;
  assign sum_12[20] = _5404_ ^ _5403_ /*22538*/;
  assign _5405_ = _5404_ & _5403_ /*22537*/;
  assign _5406_ = inv_12[20] & r_11[20] /*22536*/;
  assign _5407_ = _5405_ | _5406_ /*22535*/;
  assign _5408_ = inv_12[21] ^ r_11[21] /*22533*/;
  assign sum_12[21] = _5408_ ^ _5407_ /*22532*/;
  assign _5409_ = _5408_ & _5407_ /*22531*/;
  assign _5410_ = inv_12[21] & r_11[21] /*22530*/;
  assign _5411_ = _5409_ | _5410_ /*22529*/;
  assign _5412_ = inv_12[22] ^ r_11[22] /*22527*/;
  assign sum_12[22] = _5412_ ^ _5411_ /*22526*/;
  assign _5413_ = _5412_ & _5411_ /*22525*/;
  assign _5414_ = inv_12[22] & r_11[22] /*22524*/;
  assign _5415_ = _5413_ | _5414_ /*22523*/;
  assign _5416_ = inv_12[23] ^ r_11[23] /*22521*/;
  assign sum_12[23] = _5416_ ^ _5415_ /*22520*/;
  assign _5417_ = _5416_ & _5415_ /*22519*/;
  assign _5418_ = inv_12[23] & r_11[23] /*22518*/;
  assign _5419_ = _5417_ | _5418_ /*22517*/;
  assign _5420_ = inv_12[24] ^ r_11[24] /*22515*/;
  assign sum_12[24] = _5420_ ^ _5419_ /*22514*/;
  assign _5421_ = _5420_ & _5419_ /*22513*/;
  assign _5422_ = inv_12[24] & r_11[24] /*22512*/;
  assign _5423_ = _5421_ | _5422_ /*22511*/;
  assign _5424_ = inv_12[25] ^ r_11[25] /*22509*/;
  assign sum_12[25] = _5424_ ^ _5423_ /*22508*/;
  assign _5425_ = _5424_ & _5423_ /*22507*/;
  assign _5426_ = inv_12[25] & r_11[25] /*22506*/;
  assign _5427_ = _5425_ | _5426_ /*22505*/;
  assign _5428_ = inv_12[26] ^ r_11[26] /*22503*/;
  assign sum_12[26] = _5428_ ^ _5427_ /*22502*/;
  assign _5429_ = _5428_ & _5427_ /*22501*/;
  assign _5430_ = inv_12[26] & r_11[26] /*22500*/;
  assign _5431_ = _5429_ | _5430_ /*22499*/;
  assign _5432_ = inv_12[27] ^ r_11[27] /*22497*/;
  assign sum_12[27] = _5432_ ^ _5431_ /*22496*/;
  assign _5433_ = _5432_ & _5431_ /*22495*/;
  assign _5434_ = inv_12[27] & r_11[27] /*22494*/;
  assign _5435_ = _5433_ | _5434_ /*22493*/;
  assign _5436_ = inv_12[28] ^ r_11[28] /*22491*/;
  assign sum_12[28] = _5436_ ^ _5435_ /*22490*/;
  assign _5437_ = _5436_ & _5435_ /*22489*/;
  assign _5438_ = inv_12[28] & r_11[28] /*22488*/;
  assign _5439_ = _5437_ | _5438_ /*22487*/;
  assign _5440_ = inv_12[29] ^ r_11[29] /*22485*/;
  assign sum_12[29] = _5440_ ^ _5439_ /*22484*/;
  assign _5441_ = _5440_ & _5439_ /*22483*/;
  assign _5442_ = inv_12[29] & r_11[29] /*22482*/;
  assign _5443_ = _5441_ | _5442_ /*22481*/;
  assign _5444_ = inv_12[30] ^ r_11[30] /*22479*/;
  assign sum_12[30] = _5444_ ^ _5443_ /*22478*/;
  assign _5445_ = _5444_ & _5443_ /*22477*/;
  assign _5446_ = inv_12[30] & r_11[30] /*22476*/;
  assign _5447_ = _5445_ | _5446_ /*22475*/;
  assign _5448_ = inv_12[31] ^ r_11[31] /*22473*/;
  assign sum_12[31] = _5448_ ^ _5447_ /*22472*/;
  assign _5449_ = _5448_ & _5447_ /*22471*/;
  assign _5450_ = inv_12[31] & r_11[31] /*22470*/;
  assign _5451_ = _5449_ | _5450_ /*22469*/;
  assign _5452_ = inv_12[32] ^ r_11[32] /*22467*/;
  assign sum_12[32] = _5452_ ^ _5451_ /*22466*/;
  assign _5453_ = _5452_ & _5451_ /*22465*/;
  assign _5454_ = inv_12[32] & r_11[32] /*22464*/;
  assign _5455_ = _5453_ | _5454_ /*22463*/;
  assign _5456_ = inv_12[33] ^ r_11[33] /*22461*/;
  assign sum_12[33] = _5456_ ^ _5455_ /*22460*/;
  assign _5457_ = _5456_ & _5455_ /*22459*/;
  assign _5458_ = inv_12[33] & r_11[33] /*22458*/;
  assign _5459_ = _5457_ | _5458_ /*22457*/;
  assign _5460_ = inv_12[34] ^ r_11[34] /*22455*/;
  assign sum_12[34] = _5460_ ^ _5459_ /*22454*/;
  assign _5461_ = _5460_ & _5459_ /*22453*/;
  assign _5462_ = inv_12[34] & r_11[34] /*22452*/;
  assign _5463_ = _5461_ | _5462_ /*22451*/;
  assign _5464_ = inv_12[35] ^ r_11[35] /*22449*/;
  assign sum_12[35] = _5464_ ^ _5463_ /*22448*/;
  assign _5465_ = _5464_ & _5463_ /*22447*/;
  assign _5466_ = inv_12[35] & r_11[35] /*22446*/;
  assign _5467_ = _5465_ | _5466_ /*22445*/;
  assign _5468_ = inv_12[36] ^ r_11[36] /*22443*/;
  assign sum_12[36] = _5468_ ^ _5467_ /*22442*/;
  assign _5469_ = _5468_ & _5467_ /*22441*/;
  assign _5470_ = inv_12[36] & r_11[36] /*22440*/;
  assign _5471_ = _5469_ | _5470_ /*22439*/;
  assign _5472_ = inv_12[37] ^ r_11[37] /*22437*/;
  assign sum_12[37] = _5472_ ^ _5471_ /*22436*/;
  assign _5473_ = _5472_ & _5471_ /*22435*/;
  assign _5474_ = inv_12[37] & r_11[37] /*22434*/;
  assign _5475_ = _5473_ | _5474_ /*22433*/;
  assign _5476_ = inv_12[38] ^ r_11[38] /*22431*/;
  assign sum_12[38] = _5476_ ^ _5475_ /*22430*/;
  assign _5477_ = _5476_ & _5475_ /*22429*/;
  assign _5478_ = inv_12[38] & r_11[38] /*22428*/;
  assign _5479_ = _5477_ | _5478_ /*22427*/;
  assign _5480_ = inv_12[39] ^ r_11[39] /*22425*/;
  assign sum_12[39] = _5480_ ^ _5479_ /*22424*/;
  assign _5481_ = _5480_ & _5479_ /*22423*/;
  assign _5482_ = inv_12[39] & r_11[39] /*22422*/;
  assign _5483_ = _5481_ | _5482_ /*22421*/;
  assign _5484_ = inv_12[40] ^ r_11[40] /*22419*/;
  assign sum_12[40] = _5484_ ^ _5483_ /*22418*/;
  assign _5485_ = _5484_ & _5483_ /*22417*/;
  assign _5486_ = inv_12[40] & r_11[40] /*22416*/;
  assign _5487_ = _5485_ | _5486_ /*22415*/;
  assign _5488_ = inv_12[41] ^ r_11[41] /*22413*/;
  assign sum_12[41] = _5488_ ^ _5487_ /*22412*/;
  assign _5489_ = _5488_ & _5487_ /*22411*/;
  assign _5490_ = inv_12[41] & r_11[41] /*22410*/;
  assign _5491_ = _5489_ | _5490_ /*22409*/;
  assign _5492_ = inv_12[42] ^ r_11[42] /*22407*/;
  assign sum_12[42] = _5492_ ^ _5491_ /*22406*/;
  assign _5493_ = _5492_ & _5491_ /*22405*/;
  assign _5494_ = inv_12[42] & r_11[42] /*22404*/;
  assign _5495_ = _5493_ | _5494_ /*22403*/;
  assign _5496_ = inv_12[43] ^ r_11[43] /*22401*/;
  assign sum_12[43] = _5496_ ^ _5495_ /*22400*/;
  assign _5497_ = _5496_ & _5495_ /*22399*/;
  assign _5498_ = inv_12[43] & r_11[43] /*22398*/;
  assign _5499_ = _5497_ | _5498_ /*22397*/;
  assign _5500_ = inv_12[44] ^ r_11[44] /*22395*/;
  assign sum_12[44] = _5500_ ^ _5499_ /*22394*/;
  assign _5501_ = _5500_ & _5499_ /*22393*/;
  assign _5502_ = inv_12[44] & r_11[44] /*22392*/;
  assign _5503_ = _5501_ | _5502_ /*22391*/;
  assign _5504_ = inv_12[45] ^ r_11[45] /*22389*/;
  assign sum_12[45] = _5504_ ^ _5503_ /*22388*/;
  assign _5505_ = _5504_ & _5503_ /*22387*/;
  assign _5506_ = inv_12[45] & r_11[45] /*22386*/;
  assign _5507_ = _5505_ | _5506_ /*22385*/;
  assign _5508_ = inv_12[46] ^ r_11[46] /*22383*/;
  assign sum_12[46] = _5508_ ^ _5507_ /*22382*/;
  assign _5509_ = _5508_ & _5507_ /*22381*/;
  assign _5510_ = inv_12[46] & r_11[46] /*22380*/;
  assign _5511_ = _5509_ | _5510_ /*22379*/;
  assign _5512_ = inv_12[47] ^ r_11[47] /*22377*/;
  assign sum_12[47] = _5512_ ^ _5511_ /*22376*/;
  assign _5513_ = _5512_ & _5511_ /*22375*/;
  assign _5514_ = inv_12[47] & r_11[47] /*22374*/;
  assign _5515_ = _5513_ | _5514_ /*22373*/;
  assign _5516_ = inv_12[48] ^ r_11[48] /*22371*/;
  assign sum_12[48] = _5516_ ^ _5515_ /*22370*/;
  assign _5517_ = _5516_ & _5515_ /*22369*/;
  assign _5518_ = inv_12[48] & r_11[48] /*22368*/;
  assign _5519_ = _5517_ | _5518_ /*22367*/;
  assign _5520_ = inv_12[49] ^ r_11[49] /*22365*/;
  assign sum_12[49] = _5520_ ^ _5519_ /*22364*/;
  assign _5521_ = _5520_ & _5519_ /*22363*/;
  assign _5522_ = inv_12[49] & r_11[49] /*22362*/;
  assign _5523_ = _5521_ | _5522_ /*22361*/;
  assign _5524_ = inv_12[50] ^ r_11[50] /*22359*/;
  assign sum_12[50] = _5524_ ^ _5523_ /*22358*/;
  assign _5525_ = _5524_ & _5523_ /*22357*/;
  assign _5526_ = inv_12[50] & r_11[50] /*22356*/;
  assign _5527_ = _5525_ | _5526_ /*22355*/;
  assign _5528_ = inv_12[51] ^ r_11[51] /*22353*/;
  assign sum_12[51] = _5528_ ^ _5527_ /*22352*/;
  assign _5529_ = _5528_ & _5527_ /*22351*/;
  assign _5530_ = inv_12[51] & r_11[51] /*22350*/;
  assign _5531_ = _5529_ | _5530_ /*22349*/;
  assign _5532_ = inv_12[52] ^ r_11[52] /*22347*/;
  assign sum_12[52] = _5532_ ^ _5531_ /*22346*/;
  assign _5533_ = _5532_ & _5531_ /*22345*/;
  assign _5534_ = inv_12[52] & r_11[52] /*22344*/;
  assign _5535_ = _5533_ | _5534_ /*22343*/;
  assign _5536_ = inv_12[53] ^ r_11[53] /*22341*/;
  assign sum_12[53] = _5536_ ^ _5535_ /*22340*/;
  assign _5537_ = _5536_ & _5535_ /*22339*/;
  assign _5538_ = inv_12[53] & r_11[53] /*22338*/;
  assign _5539_ = _5537_ | _5538_ /*22337*/;
  assign _5540_ = inv_12[54] ^ r_11[54] /*22335*/;
  assign sum_12[54] = _5540_ ^ _5539_ /*22334*/;
  assign _5541_ = _5540_ & _5539_ /*22333*/;
  assign _5542_ = inv_12[54] & r_11[54] /*22332*/;
  assign _5543_ = _5541_ | _5542_ /*22331*/;
  assign _5544_ = inv_12[55] ^ r_11[55] /*22329*/;
  assign sum_12[55] = _5544_ ^ _5543_ /*22328*/;
  assign _5545_ = _5544_ & _5543_ /*22327*/;
  assign _5546_ = inv_12[55] & r_11[55] /*22326*/;
  assign _5547_ = _5545_ | _5546_ /*22325*/;
  assign _5548_ = inv_12[56] ^ r_11[56] /*22323*/;
  assign sum_12[56] = _5548_ ^ _5547_ /*22322*/;
  assign _5549_ = _5548_ & _5547_ /*22321*/;
  assign _5550_ = inv_12[56] & r_11[56] /*22320*/;
  assign _5551_ = _5549_ | _5550_ /*22319*/;
  assign _5552_ = inv_12[57] ^ r_11[57] /*22317*/;
  assign sum_12[57] = _5552_ ^ _5551_ /*22316*/;
  assign _5553_ = _5552_ & _5551_ /*22315*/;
  assign _5554_ = inv_12[57] & r_11[57] /*22314*/;
  assign _5555_ = _5553_ | _5554_ /*22313*/;
  assign _5556_ = inv_12[58] ^ r_11[58] /*22311*/;
  assign sum_12[58] = _5556_ ^ _5555_ /*22310*/;
  assign _5557_ = _5556_ & _5555_ /*22309*/;
  assign _5558_ = inv_12[58] & r_11[58] /*22308*/;
  assign _5559_ = _5557_ | _5558_ /*22307*/;
  assign _5560_ = inv_12[59] ^ r_11[59] /*22305*/;
  assign sum_12[59] = _5560_ ^ _5559_ /*22304*/;
  assign _5561_ = _5560_ & _5559_ /*22303*/;
  assign _5562_ = inv_12[59] & r_11[59] /*22302*/;
  assign _5563_ = _5561_ | _5562_ /*22301*/;
  assign _5564_ = inv_12[60] ^ r_11[60] /*22299*/;
  assign sum_12[60] = _5564_ ^ _5563_ /*22298*/;
  assign _5565_ = _5564_ & _5563_ /*22297*/;
  assign _5566_ = inv_12[60] & r_11[60] /*22296*/;
  assign _5567_ = _5565_ | _5566_ /*22295*/;
  assign _5568_ = inv_12[61] ^ r_11[61] /*22293*/;
  assign sum_12[61] = _5568_ ^ _5567_ /*22292*/;
  assign _5569_ = _5568_ & _5567_ /*22291*/;
  assign _5570_ = inv_12[61] & r_11[61] /*22290*/;
  assign _5571_ = _5569_ | _5570_ /*22289*/;
  assign _5572_ = inv_12[62] ^ r_11[62] /*22287*/;
  assign sum_12[62] = _5572_ ^ _5571_ /*22286*/;
  assign _5573_ = _5572_ & _5571_ /*22285*/;
  assign _5574_ = inv_12[62] & r_11[62] /*22284*/;
  assign _5575_ = _5573_ | _5574_ /*22283*/;
  assign _5576_ = inv_12[63] ^ r_11[63] /*22281*/;
  assign sum_12[63] = _5576_ ^ _5575_ /*22280*/;
  assign _5577_ = _5576_ & _5575_ /*22279*/;
  assign _5578_ = inv_12[63] & r_11[63] /*22278*/;
  assign _5579_ = _5577_ | _5578_ /*22277*/;
  assign _5580_ = inv_12[64] ^ r_11[64] /*22275*/;
  assign sum_12[64] = _5580_ ^ _5579_ /*22274*/;
  assign _5581_ = _5580_ & _5579_ /*22273*/;
  assign _5582_ = inv_12[64] & r_11[64] /*22272*/;
  assign _5583_ = _5581_ | _5582_ /*22271*/;
  assign _5584_ = inv_12[65] ^ r_11[65] /*22269*/;
  assign sum_12[65] = _5584_ ^ _5583_ /*22268*/;
  assign _5585_ = _5584_ & _5583_ /*22267*/;
  assign _5586_ = inv_12[65] & r_11[65] /*22266*/;
  assign _5587_ = _5585_ | _5586_ /*22265*/;
  assign _5588_ = inv_12[66] ^ r_11[66] /*22263*/;
  assign sum_12[66] = _5588_ ^ _5587_ /*22262*/;
  assign _5589_ = _5588_ & _5587_ /*22261*/;
  assign _5590_ = inv_12[66] & r_11[66] /*22260*/;
  assign _5591_ = _5589_ | _5590_ /*22259*/;
  assign _5592_ = inv_12[67] ^ r_11[67] /*22257*/;
  assign sum_12[67] = _5592_ ^ _5591_ /*22256*/;
  assign _5593_ = _5592_ & _5591_ /*22255*/;
  assign _5594_ = inv_12[67] & r_11[67] /*22254*/;
  assign _5595_ = _5593_ | _5594_ /*22253*/;
  assign _5596_ = inv_12[68] ^ r_11[68] /*22251*/;
  assign sum_12[68] = _5596_ ^ _5595_ /*22250*/;
  assign _5597_ = _5596_ & _5595_ /*22249*/;
  assign _5598_ = inv_12[68] & r_11[68] /*22248*/;
  assign _5599_ = _5597_ | _5598_ /*22247*/;
  assign _5600_ = inv_12[69] ^ r_11[69] /*22245*/;
  assign sum_12[69] = _5600_ ^ _5599_ /*22244*/;
  assign _5601_ = _5600_ & _5599_ /*22243*/;
  assign _5602_ = inv_12[69] & r_11[69] /*22242*/;
  assign _5603_ = _5601_ | _5602_ /*22241*/;
  assign _5604_ = inv_12[70] ^ r_11[70] /*22239*/;
  assign sum_12[70] = _5604_ ^ _5603_ /*22238*/;
  assign _5605_ = _5604_ & _5603_ /*22237*/;
  assign _5606_ = inv_12[70] & r_11[70] /*22236*/;
  assign _5607_ = _5605_ | _5606_ /*22235*/;
  assign _5608_ = inv_12[71] ^ r_11[71] /*22233*/;
  assign sum_12[71] = _5608_ ^ _5607_ /*22232*/;
  assign _5609_ = _5608_ & _5607_ /*22231*/;
  assign _5610_ = inv_12[71] & r_11[71] /*22230*/;
  assign _5611_ = _5609_ | _5610_ /*22229*/;
  assign _5612_ = inv_12[72] ^ r_11[72] /*22227*/;
  assign sum_12[72] = _5612_ ^ _5611_ /*22226*/;
  assign _5613_ = _5612_ & _5611_ /*22225*/;
  assign _5614_ = inv_12[72] & r_11[72] /*22224*/;
  assign _5615_ = _5613_ | _5614_ /*22223*/;
  assign _5616_ = inv_12[73] ^ r_11[73] /*22221*/;
  assign sum_12[73] = _5616_ ^ _5615_ /*22220*/;
  assign _5617_ = _5616_ & _5615_ /*22219*/;
  assign _5618_ = inv_12[73] & r_11[73] /*22218*/;
  assign _5619_ = _5617_ | _5618_ /*22217*/;
  assign _5620_ = _5619_ ^ _5615_ /*22216*/;
  assign _5621_ = ~_5620_ /*22215*/;
  assign _5622_ = sum_12[73] & _5621_ /*22214*/;
  assign _5623_ = _5620_ & _5619_ /*22213*/;
  assign sum_12[74] = _5623_ | _5622_ /*22212*/;
  assign q[20] = ~sum_12[74] /*22211*/;
  assign m_12[0] = r_11[0] /*22210*/;
  assign m_12[1] = r_11[1] /*22209*/;
  assign m_12[2] = r_11[2] /*22208*/;
  assign m_12[3] = r_11[3] /*22207*/;
  assign m_12[4] = r_11[4] /*22206*/;
  assign m_12[5] = r_11[5] /*22205*/;
  assign m_12[6] = r_11[6] /*22204*/;
  assign m_12[7] = r_11[7] /*22203*/;
  assign m_12[8] = r_11[8] /*22202*/;
  assign m_12[9] = r_11[9] /*22201*/;
  assign m_12[10] = r_11[10] /*22200*/;
  assign m_12[11] = r_11[11] /*22199*/;
  assign m_12[12] = r_11[12] /*22198*/;
  assign m_12[13] = r_11[13] /*22197*/;
  assign m_12[14] = r_11[14] /*22196*/;
  assign m_12[15] = r_11[15] /*22195*/;
  assign m_12[16] = r_11[16] /*22194*/;
  assign m_12[17] = r_11[17] /*22193*/;
  assign m_12[18] = r_11[18] /*22192*/;
  assign m_12[19] = r_11[19] /*22191*/;
  assign m_12[20] = r_11[20] /*22190*/;
  assign m_12[21] = r_11[21] /*22189*/;
  assign m_12[22] = r_11[22] /*22188*/;
  assign m_12[23] = r_11[23] /*22187*/;
  assign m_12[24] = r_11[24] /*22186*/;
  assign m_12[25] = r_11[25] /*22185*/;
  assign m_12[26] = r_11[26] /*22184*/;
  assign m_12[27] = r_11[27] /*22183*/;
  assign m_12[28] = r_11[28] /*22182*/;
  assign m_12[29] = r_11[29] /*22181*/;
  assign m_12[30] = r_11[30] /*22180*/;
  assign m_12[31] = r_11[31] /*22179*/;
  assign m_12[32] = r_11[32] /*22178*/;
  assign m_12[33] = r_11[33] /*22177*/;
  assign m_12[34] = r_11[34] /*22176*/;
  assign m_12[35] = r_11[35] /*22175*/;
  assign m_12[36] = r_11[36] /*22174*/;
  assign m_12[37] = r_11[37] /*22173*/;
  assign m_12[38] = r_11[38] /*22172*/;
  assign m_12[39] = r_11[39] /*22171*/;
  assign m_12[40] = r_11[40] /*22170*/;
  assign m_12[41] = r_11[41] /*22169*/;
  assign m_12[42] = r_11[42] /*22168*/;
  assign m_12[43] = r_11[43] /*22167*/;
  assign m_12[44] = r_11[44] /*22166*/;
  assign m_12[45] = r_11[45] /*22165*/;
  assign m_12[46] = r_11[46] /*22164*/;
  assign m_12[47] = r_11[47] /*22163*/;
  assign m_12[48] = r_11[48] /*22162*/;
  assign m_12[49] = r_11[49] /*22161*/;
  assign m_12[50] = r_11[50] /*22160*/;
  assign m_12[51] = r_11[51] /*22159*/;
  assign m_12[52] = r_11[52] /*22158*/;
  assign m_12[53] = r_11[53] /*22157*/;
  assign m_12[54] = r_11[54] /*22156*/;
  assign m_12[55] = r_11[55] /*22155*/;
  assign m_12[56] = r_11[56] /*22154*/;
  assign m_12[57] = r_11[57] /*22153*/;
  assign m_12[58] = r_11[58] /*22152*/;
  assign m_12[59] = r_11[59] /*22151*/;
  assign m_12[60] = r_11[60] /*22150*/;
  assign m_12[61] = r_11[61] /*22149*/;
  assign m_12[62] = r_11[62] /*22148*/;
  assign m_12[63] = r_11[63] /*22147*/;
  assign m_12[64] = r_11[64] /*22146*/;
  assign m_12[65] = r_11[65] /*22145*/;
  assign m_12[66] = r_11[66] /*22144*/;
  assign m_12[67] = r_11[67] /*22143*/;
  assign m_12[68] = r_11[68] /*22142*/;
  assign m_12[69] = r_11[69] /*22141*/;
  assign m_12[70] = r_11[70] /*22140*/;
  assign m_12[71] = r_11[71] /*22139*/;
  assign m_12[72] = r_11[72] /*22138*/;
  assign m_12[73] = r_11[73] /*22137*/;
  assign m_12[74] = r_11[73] /*22136*/;
  assign _5625_ = ~q[20] /*22135*/;
  assign _5626_ = sum_12[0] & q[20] /*22134*/;
  assign _5627_ = m_12[0] & _5625_ /*22133*/;
  assign r_12[0] = _5627_ | _5626_ /*22132*/;
  assign _5628_ = ~q[20] /*22131*/;
  assign _5629_ = sum_12[1] & q[20] /*22130*/;
  assign _5630_ = m_12[1] & _5628_ /*22129*/;
  assign r_12[1] = _5630_ | _5629_ /*22128*/;
  assign _5631_ = ~q[20] /*22127*/;
  assign _5632_ = sum_12[2] & q[20] /*22126*/;
  assign _5633_ = m_12[2] & _5631_ /*22125*/;
  assign r_12[2] = _5633_ | _5632_ /*22124*/;
  assign _5634_ = ~q[20] /*22123*/;
  assign _5635_ = sum_12[3] & q[20] /*22122*/;
  assign _5636_ = m_12[3] & _5634_ /*22121*/;
  assign r_12[3] = _5636_ | _5635_ /*22120*/;
  assign _5637_ = ~q[20] /*22119*/;
  assign _5638_ = sum_12[4] & q[20] /*22118*/;
  assign _5639_ = m_12[4] & _5637_ /*22117*/;
  assign r_12[4] = _5639_ | _5638_ /*22116*/;
  assign _5640_ = ~q[20] /*22115*/;
  assign _5641_ = sum_12[5] & q[20] /*22114*/;
  assign _5642_ = m_12[5] & _5640_ /*22113*/;
  assign r_12[5] = _5642_ | _5641_ /*22112*/;
  assign _5643_ = ~q[20] /*22111*/;
  assign _5644_ = sum_12[6] & q[20] /*22110*/;
  assign _5645_ = m_12[6] & _5643_ /*22109*/;
  assign r_12[6] = _5645_ | _5644_ /*22108*/;
  assign _5646_ = ~q[20] /*22107*/;
  assign _5647_ = sum_12[7] & q[20] /*22106*/;
  assign _5648_ = m_12[7] & _5646_ /*22105*/;
  assign r_12[7] = _5648_ | _5647_ /*22104*/;
  assign _5649_ = ~q[20] /*22103*/;
  assign _5650_ = sum_12[8] & q[20] /*22102*/;
  assign _5651_ = m_12[8] & _5649_ /*22101*/;
  assign r_12[8] = _5651_ | _5650_ /*22100*/;
  assign _5652_ = ~q[20] /*22099*/;
  assign _5653_ = sum_12[9] & q[20] /*22098*/;
  assign _5654_ = m_12[9] & _5652_ /*22097*/;
  assign r_12[9] = _5654_ | _5653_ /*22096*/;
  assign _5655_ = ~q[20] /*22095*/;
  assign _5656_ = sum_12[10] & q[20] /*22094*/;
  assign _5657_ = m_12[10] & _5655_ /*22093*/;
  assign r_12[10] = _5657_ | _5656_ /*22092*/;
  assign _5658_ = ~q[20] /*22091*/;
  assign _5659_ = sum_12[11] & q[20] /*22090*/;
  assign _5660_ = m_12[11] & _5658_ /*22089*/;
  assign r_12[11] = _5660_ | _5659_ /*22088*/;
  assign _5661_ = ~q[20] /*22087*/;
  assign _5662_ = sum_12[12] & q[20] /*22086*/;
  assign _5663_ = m_12[12] & _5661_ /*22085*/;
  assign r_12[12] = _5663_ | _5662_ /*22084*/;
  assign _5664_ = ~q[20] /*22083*/;
  assign _5665_ = sum_12[13] & q[20] /*22082*/;
  assign _5666_ = m_12[13] & _5664_ /*22081*/;
  assign r_12[13] = _5666_ | _5665_ /*22080*/;
  assign _5667_ = ~q[20] /*22079*/;
  assign _5668_ = sum_12[14] & q[20] /*22078*/;
  assign _5669_ = m_12[14] & _5667_ /*22077*/;
  assign r_12[14] = _5669_ | _5668_ /*22076*/;
  assign _5670_ = ~q[20] /*22075*/;
  assign _5671_ = sum_12[15] & q[20] /*22074*/;
  assign _5672_ = m_12[15] & _5670_ /*22073*/;
  assign r_12[15] = _5672_ | _5671_ /*22072*/;
  assign _5673_ = ~q[20] /*22071*/;
  assign _5674_ = sum_12[16] & q[20] /*22070*/;
  assign _5675_ = m_12[16] & _5673_ /*22069*/;
  assign r_12[16] = _5675_ | _5674_ /*22068*/;
  assign _5676_ = ~q[20] /*22067*/;
  assign _5677_ = sum_12[17] & q[20] /*22066*/;
  assign _5678_ = m_12[17] & _5676_ /*22065*/;
  assign r_12[17] = _5678_ | _5677_ /*22064*/;
  assign _5679_ = ~q[20] /*22063*/;
  assign _5680_ = sum_12[18] & q[20] /*22062*/;
  assign _5681_ = m_12[18] & _5679_ /*22061*/;
  assign r_12[18] = _5681_ | _5680_ /*22060*/;
  assign _5682_ = ~q[20] /*22059*/;
  assign _5683_ = sum_12[19] & q[20] /*22058*/;
  assign _5684_ = m_12[19] & _5682_ /*22057*/;
  assign r_12[19] = _5684_ | _5683_ /*22056*/;
  assign _5685_ = ~q[20] /*22055*/;
  assign _5686_ = sum_12[20] & q[20] /*22054*/;
  assign _5687_ = m_12[20] & _5685_ /*22053*/;
  assign r_12[20] = _5687_ | _5686_ /*22052*/;
  assign _5688_ = ~q[20] /*22051*/;
  assign _5689_ = sum_12[21] & q[20] /*22050*/;
  assign _5690_ = m_12[21] & _5688_ /*22049*/;
  assign r_12[21] = _5690_ | _5689_ /*22048*/;
  assign _5691_ = ~q[20] /*22047*/;
  assign _5692_ = sum_12[22] & q[20] /*22046*/;
  assign _5693_ = m_12[22] & _5691_ /*22045*/;
  assign r_12[22] = _5693_ | _5692_ /*22044*/;
  assign _5694_ = ~q[20] /*22043*/;
  assign _5695_ = sum_12[23] & q[20] /*22042*/;
  assign _5696_ = m_12[23] & _5694_ /*22041*/;
  assign r_12[23] = _5696_ | _5695_ /*22040*/;
  assign _5697_ = ~q[20] /*22039*/;
  assign _5698_ = sum_12[24] & q[20] /*22038*/;
  assign _5699_ = m_12[24] & _5697_ /*22037*/;
  assign r_12[24] = _5699_ | _5698_ /*22036*/;
  assign _5700_ = ~q[20] /*22035*/;
  assign _5701_ = sum_12[25] & q[20] /*22034*/;
  assign _5702_ = m_12[25] & _5700_ /*22033*/;
  assign r_12[25] = _5702_ | _5701_ /*22032*/;
  assign _5703_ = ~q[20] /*22031*/;
  assign _5704_ = sum_12[26] & q[20] /*22030*/;
  assign _5705_ = m_12[26] & _5703_ /*22029*/;
  assign r_12[26] = _5705_ | _5704_ /*22028*/;
  assign _5706_ = ~q[20] /*22027*/;
  assign _5707_ = sum_12[27] & q[20] /*22026*/;
  assign _5708_ = m_12[27] & _5706_ /*22025*/;
  assign r_12[27] = _5708_ | _5707_ /*22024*/;
  assign _5709_ = ~q[20] /*22023*/;
  assign _5710_ = sum_12[28] & q[20] /*22022*/;
  assign _5711_ = m_12[28] & _5709_ /*22021*/;
  assign r_12[28] = _5711_ | _5710_ /*22020*/;
  assign _5712_ = ~q[20] /*22019*/;
  assign _5713_ = sum_12[29] & q[20] /*22018*/;
  assign _5714_ = m_12[29] & _5712_ /*22017*/;
  assign r_12[29] = _5714_ | _5713_ /*22016*/;
  assign _5715_ = ~q[20] /*22015*/;
  assign _5716_ = sum_12[30] & q[20] /*22014*/;
  assign _5717_ = m_12[30] & _5715_ /*22013*/;
  assign r_12[30] = _5717_ | _5716_ /*22012*/;
  assign _5718_ = ~q[20] /*22011*/;
  assign _5719_ = sum_12[31] & q[20] /*22010*/;
  assign _5720_ = m_12[31] & _5718_ /*22009*/;
  assign r_12[31] = _5720_ | _5719_ /*22008*/;
  assign _5721_ = ~q[20] /*22007*/;
  assign _5722_ = sum_12[32] & q[20] /*22006*/;
  assign _5723_ = m_12[32] & _5721_ /*22005*/;
  assign r_12[32] = _5723_ | _5722_ /*22004*/;
  assign _5724_ = ~q[20] /*22003*/;
  assign _5725_ = sum_12[33] & q[20] /*22002*/;
  assign _5726_ = m_12[33] & _5724_ /*22001*/;
  assign r_12[33] = _5726_ | _5725_ /*22000*/;
  assign _5727_ = ~q[20] /*21999*/;
  assign _5728_ = sum_12[34] & q[20] /*21998*/;
  assign _5729_ = m_12[34] & _5727_ /*21997*/;
  assign r_12[34] = _5729_ | _5728_ /*21996*/;
  assign _5730_ = ~q[20] /*21995*/;
  assign _5731_ = sum_12[35] & q[20] /*21994*/;
  assign _5732_ = m_12[35] & _5730_ /*21993*/;
  assign r_12[35] = _5732_ | _5731_ /*21992*/;
  assign _5733_ = ~q[20] /*21991*/;
  assign _5734_ = sum_12[36] & q[20] /*21990*/;
  assign _5735_ = m_12[36] & _5733_ /*21989*/;
  assign r_12[36] = _5735_ | _5734_ /*21988*/;
  assign _5736_ = ~q[20] /*21987*/;
  assign _5737_ = sum_12[37] & q[20] /*21986*/;
  assign _5738_ = m_12[37] & _5736_ /*21985*/;
  assign r_12[37] = _5738_ | _5737_ /*21984*/;
  assign _5739_ = ~q[20] /*21983*/;
  assign _5740_ = sum_12[38] & q[20] /*21982*/;
  assign _5741_ = m_12[38] & _5739_ /*21981*/;
  assign r_12[38] = _5741_ | _5740_ /*21980*/;
  assign _5742_ = ~q[20] /*21979*/;
  assign _5743_ = sum_12[39] & q[20] /*21978*/;
  assign _5744_ = m_12[39] & _5742_ /*21977*/;
  assign r_12[39] = _5744_ | _5743_ /*21976*/;
  assign _5745_ = ~q[20] /*21975*/;
  assign _5746_ = sum_12[40] & q[20] /*21974*/;
  assign _5747_ = m_12[40] & _5745_ /*21973*/;
  assign r_12[40] = _5747_ | _5746_ /*21972*/;
  assign _5748_ = ~q[20] /*21971*/;
  assign _5749_ = sum_12[41] & q[20] /*21970*/;
  assign _5750_ = m_12[41] & _5748_ /*21969*/;
  assign r_12[41] = _5750_ | _5749_ /*21968*/;
  assign _5751_ = ~q[20] /*21967*/;
  assign _5752_ = sum_12[42] & q[20] /*21966*/;
  assign _5753_ = m_12[42] & _5751_ /*21965*/;
  assign r_12[42] = _5753_ | _5752_ /*21964*/;
  assign _5754_ = ~q[20] /*21963*/;
  assign _5755_ = sum_12[43] & q[20] /*21962*/;
  assign _5756_ = m_12[43] & _5754_ /*21961*/;
  assign r_12[43] = _5756_ | _5755_ /*21960*/;
  assign _5757_ = ~q[20] /*21959*/;
  assign _5758_ = sum_12[44] & q[20] /*21958*/;
  assign _5759_ = m_12[44] & _5757_ /*21957*/;
  assign r_12[44] = _5759_ | _5758_ /*21956*/;
  assign _5760_ = ~q[20] /*21955*/;
  assign _5761_ = sum_12[45] & q[20] /*21954*/;
  assign _5762_ = m_12[45] & _5760_ /*21953*/;
  assign r_12[45] = _5762_ | _5761_ /*21952*/;
  assign _5763_ = ~q[20] /*21951*/;
  assign _5764_ = sum_12[46] & q[20] /*21950*/;
  assign _5765_ = m_12[46] & _5763_ /*21949*/;
  assign r_12[46] = _5765_ | _5764_ /*21948*/;
  assign _5766_ = ~q[20] /*21947*/;
  assign _5767_ = sum_12[47] & q[20] /*21946*/;
  assign _5768_ = m_12[47] & _5766_ /*21945*/;
  assign r_12[47] = _5768_ | _5767_ /*21944*/;
  assign _5769_ = ~q[20] /*21943*/;
  assign _5770_ = sum_12[48] & q[20] /*21942*/;
  assign _5771_ = m_12[48] & _5769_ /*21941*/;
  assign r_12[48] = _5771_ | _5770_ /*21940*/;
  assign _5772_ = ~q[20] /*21939*/;
  assign _5773_ = sum_12[49] & q[20] /*21938*/;
  assign _5774_ = m_12[49] & _5772_ /*21937*/;
  assign r_12[49] = _5774_ | _5773_ /*21936*/;
  assign _5775_ = ~q[20] /*21935*/;
  assign _5776_ = sum_12[50] & q[20] /*21934*/;
  assign _5777_ = m_12[50] & _5775_ /*21933*/;
  assign r_12[50] = _5777_ | _5776_ /*21932*/;
  assign _5778_ = ~q[20] /*21931*/;
  assign _5779_ = sum_12[51] & q[20] /*21930*/;
  assign _5780_ = m_12[51] & _5778_ /*21929*/;
  assign r_12[51] = _5780_ | _5779_ /*21928*/;
  assign _5781_ = ~q[20] /*21927*/;
  assign _5782_ = sum_12[52] & q[20] /*21926*/;
  assign _5783_ = m_12[52] & _5781_ /*21925*/;
  assign r_12[52] = _5783_ | _5782_ /*21924*/;
  assign _5784_ = ~q[20] /*21923*/;
  assign _5785_ = sum_12[53] & q[20] /*21922*/;
  assign _5786_ = m_12[53] & _5784_ /*21921*/;
  assign r_12[53] = _5786_ | _5785_ /*21920*/;
  assign _5787_ = ~q[20] /*21919*/;
  assign _5788_ = sum_12[54] & q[20] /*21918*/;
  assign _5789_ = m_12[54] & _5787_ /*21917*/;
  assign r_12[54] = _5789_ | _5788_ /*21916*/;
  assign _5790_ = ~q[20] /*21915*/;
  assign _5791_ = sum_12[55] & q[20] /*21914*/;
  assign _5792_ = m_12[55] & _5790_ /*21913*/;
  assign r_12[55] = _5792_ | _5791_ /*21912*/;
  assign _5793_ = ~q[20] /*21911*/;
  assign _5794_ = sum_12[56] & q[20] /*21910*/;
  assign _5795_ = m_12[56] & _5793_ /*21909*/;
  assign r_12[56] = _5795_ | _5794_ /*21908*/;
  assign _5796_ = ~q[20] /*21907*/;
  assign _5797_ = sum_12[57] & q[20] /*21906*/;
  assign _5798_ = m_12[57] & _5796_ /*21905*/;
  assign r_12[57] = _5798_ | _5797_ /*21904*/;
  assign _5799_ = ~q[20] /*21903*/;
  assign _5800_ = sum_12[58] & q[20] /*21902*/;
  assign _5801_ = m_12[58] & _5799_ /*21901*/;
  assign r_12[58] = _5801_ | _5800_ /*21900*/;
  assign _5802_ = ~q[20] /*21899*/;
  assign _5803_ = sum_12[59] & q[20] /*21898*/;
  assign _5804_ = m_12[59] & _5802_ /*21897*/;
  assign r_12[59] = _5804_ | _5803_ /*21896*/;
  assign _5805_ = ~q[20] /*21895*/;
  assign _5806_ = sum_12[60] & q[20] /*21894*/;
  assign _5807_ = m_12[60] & _5805_ /*21893*/;
  assign r_12[60] = _5807_ | _5806_ /*21892*/;
  assign _5808_ = ~q[20] /*21891*/;
  assign _5809_ = sum_12[61] & q[20] /*21890*/;
  assign _5810_ = m_12[61] & _5808_ /*21889*/;
  assign r_12[61] = _5810_ | _5809_ /*21888*/;
  assign _5811_ = ~q[20] /*21887*/;
  assign _5812_ = sum_12[62] & q[20] /*21886*/;
  assign _5813_ = m_12[62] & _5811_ /*21885*/;
  assign r_12[62] = _5813_ | _5812_ /*21884*/;
  assign _5814_ = ~q[20] /*21883*/;
  assign _5815_ = sum_12[63] & q[20] /*21882*/;
  assign _5816_ = m_12[63] & _5814_ /*21881*/;
  assign r_12[63] = _5816_ | _5815_ /*21880*/;
  assign _5817_ = ~q[20] /*21879*/;
  assign _5818_ = sum_12[64] & q[20] /*21878*/;
  assign _5819_ = m_12[64] & _5817_ /*21877*/;
  assign r_12[64] = _5819_ | _5818_ /*21876*/;
  assign _5820_ = ~q[20] /*21875*/;
  assign _5821_ = sum_12[65] & q[20] /*21874*/;
  assign _5822_ = m_12[65] & _5820_ /*21873*/;
  assign r_12[65] = _5822_ | _5821_ /*21872*/;
  assign _5823_ = ~q[20] /*21871*/;
  assign _5824_ = sum_12[66] & q[20] /*21870*/;
  assign _5825_ = m_12[66] & _5823_ /*21869*/;
  assign r_12[66] = _5825_ | _5824_ /*21868*/;
  assign _5826_ = ~q[20] /*21867*/;
  assign _5827_ = sum_12[67] & q[20] /*21866*/;
  assign _5828_ = m_12[67] & _5826_ /*21865*/;
  assign r_12[67] = _5828_ | _5827_ /*21864*/;
  assign _5829_ = ~q[20] /*21863*/;
  assign _5830_ = sum_12[68] & q[20] /*21862*/;
  assign _5831_ = m_12[68] & _5829_ /*21861*/;
  assign r_12[68] = _5831_ | _5830_ /*21860*/;
  assign _5832_ = ~q[20] /*21859*/;
  assign _5833_ = sum_12[69] & q[20] /*21858*/;
  assign _5834_ = m_12[69] & _5832_ /*21857*/;
  assign r_12[69] = _5834_ | _5833_ /*21856*/;
  assign _5835_ = ~q[20] /*21855*/;
  assign _5836_ = sum_12[70] & q[20] /*21854*/;
  assign _5837_ = m_12[70] & _5835_ /*21853*/;
  assign r_12[70] = _5837_ | _5836_ /*21852*/;
  assign _5838_ = ~q[20] /*21851*/;
  assign _5839_ = sum_12[71] & q[20] /*21850*/;
  assign _5840_ = m_12[71] & _5838_ /*21849*/;
  assign r_12[71] = _5840_ | _5839_ /*21848*/;
  assign _5841_ = ~q[20] /*21847*/;
  assign _5842_ = sum_12[72] & q[20] /*21846*/;
  assign _5843_ = m_12[72] & _5841_ /*21845*/;
  assign r_12[72] = _5843_ | _5842_ /*21844*/;
  assign _5844_ = ~q[20] /*21843*/;
  assign _5845_ = sum_12[73] & q[20] /*21842*/;
  assign _5846_ = m_12[73] & _5844_ /*21841*/;
  assign r_12[73] = _5846_ | _5845_ /*21840*/;
  assign _5847_ = ~q[20] /*21839*/;
  assign _5848_ = sum_12[74] & q[20] /*21838*/;
  assign _5849_ = m_12[74] & _5847_ /*21837*/;
  assign r_12[74] = _5849_ | _5848_ /*21836*/;
  assign inv_13[0] = oneWire /*21584*/;
  assign inv_13[1] = oneWire /*21578*/;
  assign inv_13[2] = oneWire /*21572*/;
  assign inv_13[3] = oneWire /*21566*/;
  assign inv_13[4] = oneWire /*21560*/;
  assign inv_13[5] = oneWire /*21554*/;
  assign inv_13[6] = oneWire /*21548*/;
  assign inv_13[7] = oneWire /*21542*/;
  assign inv_13[8] = oneWire /*21536*/;
  assign inv_13[9] = oneWire /*21530*/;
  assign inv_13[10] = oneWire /*21524*/;
  assign inv_13[11] = oneWire /*21518*/;
  assign inv_13[12] = oneWire /*21512*/;
  assign inv_13[13] = oneWire /*21506*/;
  assign inv_13[14] = oneWire /*21500*/;
  assign inv_13[15] = oneWire /*21494*/;
  assign inv_13[16] = oneWire /*21488*/;
  assign inv_13[17] = oneWire /*21482*/;
  assign inv_13[18] = oneWire /*21476*/;
  assign inv_13[19] = ~div[0] /*21470*/;
  assign inv_13[20] = ~div[1] /*21464*/;
  assign inv_13[21] = ~div[2] /*21458*/;
  assign inv_13[22] = ~div[3] /*21452*/;
  assign inv_13[23] = ~div[4] /*21446*/;
  assign inv_13[24] = ~div[5] /*21440*/;
  assign inv_13[25] = ~div[6] /*21434*/;
  assign inv_13[26] = ~div[7] /*21428*/;
  assign inv_13[27] = ~div[8] /*21422*/;
  assign inv_13[28] = ~div[9] /*21416*/;
  assign inv_13[29] = ~div[10] /*21410*/;
  assign inv_13[30] = ~div[11] /*21404*/;
  assign inv_13[31] = ~div[12] /*21398*/;
  assign inv_13[32] = ~div[13] /*21392*/;
  assign inv_13[33] = ~div[14] /*21386*/;
  assign inv_13[34] = ~div[15] /*21380*/;
  assign inv_13[35] = ~div[16] /*21374*/;
  assign inv_13[36] = ~div[17] /*21368*/;
  assign inv_13[37] = ~div[18] /*21362*/;
  assign inv_13[38] = ~div[19] /*21356*/;
  assign inv_13[39] = ~div[20] /*21350*/;
  assign inv_13[40] = ~div[21] /*21344*/;
  assign inv_13[41] = ~div[22] /*21338*/;
  assign inv_13[42] = ~div[23] /*21332*/;
  assign inv_13[43] = ~div[24] /*21326*/;
  assign inv_13[44] = ~div[25] /*21320*/;
  assign inv_13[45] = ~div[26] /*21314*/;
  assign inv_13[46] = ~div[27] /*21308*/;
  assign inv_13[47] = ~div[28] /*21302*/;
  assign inv_13[48] = ~div[29] /*21296*/;
  assign inv_13[49] = ~div[30] /*21290*/;
  assign inv_13[50] = oneWire /*21284*/;
  assign inv_13[51] = oneWire /*21278*/;
  assign inv_13[52] = oneWire /*21272*/;
  assign inv_13[53] = oneWire /*21266*/;
  assign inv_13[54] = oneWire /*21260*/;
  assign inv_13[55] = oneWire /*21254*/;
  assign inv_13[56] = oneWire /*21248*/;
  assign inv_13[57] = oneWire /*21242*/;
  assign inv_13[58] = oneWire /*21236*/;
  assign inv_13[59] = oneWire /*21230*/;
  assign inv_13[60] = oneWire /*21224*/;
  assign inv_13[61] = oneWire /*21218*/;
  assign inv_13[62] = oneWire /*21212*/;
  assign inv_13[63] = oneWire /*21206*/;
  assign inv_13[64] = oneWire /*21200*/;
  assign inv_13[65] = oneWire /*21194*/;
  assign inv_13[66] = oneWire /*21188*/;
  assign inv_13[67] = oneWire /*21182*/;
  assign inv_13[68] = oneWire /*21176*/;
  assign inv_13[69] = oneWire /*21170*/;
  assign inv_13[70] = oneWire /*21164*/;
  assign inv_13[71] = oneWire /*21158*/;
  assign inv_13[72] = oneWire /*21152*/;
  assign inv_13[73] = oneWire /*21146*/;
  assign inv_13[74] = oneWire /*21140*/;
  assign _5850_ = inv_13[0] ^ r_12[0] /*21583*/;
  assign sum_13[0] = _5850_ ^ oneWire /*21582*/;
  assign _5851_ = _5850_ & oneWire /*21581*/;
  assign _5852_ = inv_13[0] & r_12[0] /*21580*/;
  assign _5853_ = _5851_ | _5852_ /*21579*/;
  assign _5854_ = inv_13[1] ^ r_12[1] /*21577*/;
  assign sum_13[1] = _5854_ ^ _5853_ /*21576*/;
  assign _5855_ = _5854_ & _5853_ /*21575*/;
  assign _5856_ = inv_13[1] & r_12[1] /*21574*/;
  assign _5857_ = _5855_ | _5856_ /*21573*/;
  assign _5858_ = inv_13[2] ^ r_12[2] /*21571*/;
  assign sum_13[2] = _5858_ ^ _5857_ /*21570*/;
  assign _5859_ = _5858_ & _5857_ /*21569*/;
  assign _5860_ = inv_13[2] & r_12[2] /*21568*/;
  assign _5861_ = _5859_ | _5860_ /*21567*/;
  assign _5862_ = inv_13[3] ^ r_12[3] /*21565*/;
  assign sum_13[3] = _5862_ ^ _5861_ /*21564*/;
  assign _5863_ = _5862_ & _5861_ /*21563*/;
  assign _5864_ = inv_13[3] & r_12[3] /*21562*/;
  assign _5865_ = _5863_ | _5864_ /*21561*/;
  assign _5866_ = inv_13[4] ^ r_12[4] /*21559*/;
  assign sum_13[4] = _5866_ ^ _5865_ /*21558*/;
  assign _5867_ = _5866_ & _5865_ /*21557*/;
  assign _5868_ = inv_13[4] & r_12[4] /*21556*/;
  assign _5869_ = _5867_ | _5868_ /*21555*/;
  assign _5870_ = inv_13[5] ^ r_12[5] /*21553*/;
  assign sum_13[5] = _5870_ ^ _5869_ /*21552*/;
  assign _5871_ = _5870_ & _5869_ /*21551*/;
  assign _5872_ = inv_13[5] & r_12[5] /*21550*/;
  assign _5873_ = _5871_ | _5872_ /*21549*/;
  assign _5874_ = inv_13[6] ^ r_12[6] /*21547*/;
  assign sum_13[6] = _5874_ ^ _5873_ /*21546*/;
  assign _5875_ = _5874_ & _5873_ /*21545*/;
  assign _5876_ = inv_13[6] & r_12[6] /*21544*/;
  assign _5877_ = _5875_ | _5876_ /*21543*/;
  assign _5878_ = inv_13[7] ^ r_12[7] /*21541*/;
  assign sum_13[7] = _5878_ ^ _5877_ /*21540*/;
  assign _5879_ = _5878_ & _5877_ /*21539*/;
  assign _5880_ = inv_13[7] & r_12[7] /*21538*/;
  assign _5881_ = _5879_ | _5880_ /*21537*/;
  assign _5882_ = inv_13[8] ^ r_12[8] /*21535*/;
  assign sum_13[8] = _5882_ ^ _5881_ /*21534*/;
  assign _5883_ = _5882_ & _5881_ /*21533*/;
  assign _5884_ = inv_13[8] & r_12[8] /*21532*/;
  assign _5885_ = _5883_ | _5884_ /*21531*/;
  assign _5886_ = inv_13[9] ^ r_12[9] /*21529*/;
  assign sum_13[9] = _5886_ ^ _5885_ /*21528*/;
  assign _5887_ = _5886_ & _5885_ /*21527*/;
  assign _5888_ = inv_13[9] & r_12[9] /*21526*/;
  assign _5889_ = _5887_ | _5888_ /*21525*/;
  assign _5890_ = inv_13[10] ^ r_12[10] /*21523*/;
  assign sum_13[10] = _5890_ ^ _5889_ /*21522*/;
  assign _5891_ = _5890_ & _5889_ /*21521*/;
  assign _5892_ = inv_13[10] & r_12[10] /*21520*/;
  assign _5893_ = _5891_ | _5892_ /*21519*/;
  assign _5894_ = inv_13[11] ^ r_12[11] /*21517*/;
  assign sum_13[11] = _5894_ ^ _5893_ /*21516*/;
  assign _5895_ = _5894_ & _5893_ /*21515*/;
  assign _5896_ = inv_13[11] & r_12[11] /*21514*/;
  assign _5897_ = _5895_ | _5896_ /*21513*/;
  assign _5898_ = inv_13[12] ^ r_12[12] /*21511*/;
  assign sum_13[12] = _5898_ ^ _5897_ /*21510*/;
  assign _5899_ = _5898_ & _5897_ /*21509*/;
  assign _5900_ = inv_13[12] & r_12[12] /*21508*/;
  assign _5901_ = _5899_ | _5900_ /*21507*/;
  assign _5902_ = inv_13[13] ^ r_12[13] /*21505*/;
  assign sum_13[13] = _5902_ ^ _5901_ /*21504*/;
  assign _5903_ = _5902_ & _5901_ /*21503*/;
  assign _5904_ = inv_13[13] & r_12[13] /*21502*/;
  assign _5905_ = _5903_ | _5904_ /*21501*/;
  assign _5906_ = inv_13[14] ^ r_12[14] /*21499*/;
  assign sum_13[14] = _5906_ ^ _5905_ /*21498*/;
  assign _5907_ = _5906_ & _5905_ /*21497*/;
  assign _5908_ = inv_13[14] & r_12[14] /*21496*/;
  assign _5909_ = _5907_ | _5908_ /*21495*/;
  assign _5910_ = inv_13[15] ^ r_12[15] /*21493*/;
  assign sum_13[15] = _5910_ ^ _5909_ /*21492*/;
  assign _5911_ = _5910_ & _5909_ /*21491*/;
  assign _5912_ = inv_13[15] & r_12[15] /*21490*/;
  assign _5913_ = _5911_ | _5912_ /*21489*/;
  assign _5914_ = inv_13[16] ^ r_12[16] /*21487*/;
  assign sum_13[16] = _5914_ ^ _5913_ /*21486*/;
  assign _5915_ = _5914_ & _5913_ /*21485*/;
  assign _5916_ = inv_13[16] & r_12[16] /*21484*/;
  assign _5917_ = _5915_ | _5916_ /*21483*/;
  assign _5918_ = inv_13[17] ^ r_12[17] /*21481*/;
  assign sum_13[17] = _5918_ ^ _5917_ /*21480*/;
  assign _5919_ = _5918_ & _5917_ /*21479*/;
  assign _5920_ = inv_13[17] & r_12[17] /*21478*/;
  assign _5921_ = _5919_ | _5920_ /*21477*/;
  assign _5922_ = inv_13[18] ^ r_12[18] /*21475*/;
  assign sum_13[18] = _5922_ ^ _5921_ /*21474*/;
  assign _5923_ = _5922_ & _5921_ /*21473*/;
  assign _5924_ = inv_13[18] & r_12[18] /*21472*/;
  assign _5925_ = _5923_ | _5924_ /*21471*/;
  assign _5926_ = inv_13[19] ^ r_12[19] /*21469*/;
  assign sum_13[19] = _5926_ ^ _5925_ /*21468*/;
  assign _5927_ = _5926_ & _5925_ /*21467*/;
  assign _5928_ = inv_13[19] & r_12[19] /*21466*/;
  assign _5929_ = _5927_ | _5928_ /*21465*/;
  assign _5930_ = inv_13[20] ^ r_12[20] /*21463*/;
  assign sum_13[20] = _5930_ ^ _5929_ /*21462*/;
  assign _5931_ = _5930_ & _5929_ /*21461*/;
  assign _5932_ = inv_13[20] & r_12[20] /*21460*/;
  assign _5933_ = _5931_ | _5932_ /*21459*/;
  assign _5934_ = inv_13[21] ^ r_12[21] /*21457*/;
  assign sum_13[21] = _5934_ ^ _5933_ /*21456*/;
  assign _5935_ = _5934_ & _5933_ /*21455*/;
  assign _5936_ = inv_13[21] & r_12[21] /*21454*/;
  assign _5937_ = _5935_ | _5936_ /*21453*/;
  assign _5938_ = inv_13[22] ^ r_12[22] /*21451*/;
  assign sum_13[22] = _5938_ ^ _5937_ /*21450*/;
  assign _5939_ = _5938_ & _5937_ /*21449*/;
  assign _5940_ = inv_13[22] & r_12[22] /*21448*/;
  assign _5941_ = _5939_ | _5940_ /*21447*/;
  assign _5942_ = inv_13[23] ^ r_12[23] /*21445*/;
  assign sum_13[23] = _5942_ ^ _5941_ /*21444*/;
  assign _5943_ = _5942_ & _5941_ /*21443*/;
  assign _5944_ = inv_13[23] & r_12[23] /*21442*/;
  assign _5945_ = _5943_ | _5944_ /*21441*/;
  assign _5946_ = inv_13[24] ^ r_12[24] /*21439*/;
  assign sum_13[24] = _5946_ ^ _5945_ /*21438*/;
  assign _5947_ = _5946_ & _5945_ /*21437*/;
  assign _5948_ = inv_13[24] & r_12[24] /*21436*/;
  assign _5949_ = _5947_ | _5948_ /*21435*/;
  assign _5950_ = inv_13[25] ^ r_12[25] /*21433*/;
  assign sum_13[25] = _5950_ ^ _5949_ /*21432*/;
  assign _5951_ = _5950_ & _5949_ /*21431*/;
  assign _5952_ = inv_13[25] & r_12[25] /*21430*/;
  assign _5953_ = _5951_ | _5952_ /*21429*/;
  assign _5954_ = inv_13[26] ^ r_12[26] /*21427*/;
  assign sum_13[26] = _5954_ ^ _5953_ /*21426*/;
  assign _5955_ = _5954_ & _5953_ /*21425*/;
  assign _5956_ = inv_13[26] & r_12[26] /*21424*/;
  assign _5957_ = _5955_ | _5956_ /*21423*/;
  assign _5958_ = inv_13[27] ^ r_12[27] /*21421*/;
  assign sum_13[27] = _5958_ ^ _5957_ /*21420*/;
  assign _5959_ = _5958_ & _5957_ /*21419*/;
  assign _5960_ = inv_13[27] & r_12[27] /*21418*/;
  assign _5961_ = _5959_ | _5960_ /*21417*/;
  assign _5962_ = inv_13[28] ^ r_12[28] /*21415*/;
  assign sum_13[28] = _5962_ ^ _5961_ /*21414*/;
  assign _5963_ = _5962_ & _5961_ /*21413*/;
  assign _5964_ = inv_13[28] & r_12[28] /*21412*/;
  assign _5965_ = _5963_ | _5964_ /*21411*/;
  assign _5966_ = inv_13[29] ^ r_12[29] /*21409*/;
  assign sum_13[29] = _5966_ ^ _5965_ /*21408*/;
  assign _5967_ = _5966_ & _5965_ /*21407*/;
  assign _5968_ = inv_13[29] & r_12[29] /*21406*/;
  assign _5969_ = _5967_ | _5968_ /*21405*/;
  assign _5970_ = inv_13[30] ^ r_12[30] /*21403*/;
  assign sum_13[30] = _5970_ ^ _5969_ /*21402*/;
  assign _5971_ = _5970_ & _5969_ /*21401*/;
  assign _5972_ = inv_13[30] & r_12[30] /*21400*/;
  assign _5973_ = _5971_ | _5972_ /*21399*/;
  assign _5974_ = inv_13[31] ^ r_12[31] /*21397*/;
  assign sum_13[31] = _5974_ ^ _5973_ /*21396*/;
  assign _5975_ = _5974_ & _5973_ /*21395*/;
  assign _5976_ = inv_13[31] & r_12[31] /*21394*/;
  assign _5977_ = _5975_ | _5976_ /*21393*/;
  assign _5978_ = inv_13[32] ^ r_12[32] /*21391*/;
  assign sum_13[32] = _5978_ ^ _5977_ /*21390*/;
  assign _5979_ = _5978_ & _5977_ /*21389*/;
  assign _5980_ = inv_13[32] & r_12[32] /*21388*/;
  assign _5981_ = _5979_ | _5980_ /*21387*/;
  assign _5982_ = inv_13[33] ^ r_12[33] /*21385*/;
  assign sum_13[33] = _5982_ ^ _5981_ /*21384*/;
  assign _5983_ = _5982_ & _5981_ /*21383*/;
  assign _5984_ = inv_13[33] & r_12[33] /*21382*/;
  assign _5985_ = _5983_ | _5984_ /*21381*/;
  assign _5986_ = inv_13[34] ^ r_12[34] /*21379*/;
  assign sum_13[34] = _5986_ ^ _5985_ /*21378*/;
  assign _5987_ = _5986_ & _5985_ /*21377*/;
  assign _5988_ = inv_13[34] & r_12[34] /*21376*/;
  assign _5989_ = _5987_ | _5988_ /*21375*/;
  assign _5990_ = inv_13[35] ^ r_12[35] /*21373*/;
  assign sum_13[35] = _5990_ ^ _5989_ /*21372*/;
  assign _5991_ = _5990_ & _5989_ /*21371*/;
  assign _5992_ = inv_13[35] & r_12[35] /*21370*/;
  assign _5993_ = _5991_ | _5992_ /*21369*/;
  assign _5994_ = inv_13[36] ^ r_12[36] /*21367*/;
  assign sum_13[36] = _5994_ ^ _5993_ /*21366*/;
  assign _5995_ = _5994_ & _5993_ /*21365*/;
  assign _5996_ = inv_13[36] & r_12[36] /*21364*/;
  assign _5997_ = _5995_ | _5996_ /*21363*/;
  assign _5998_ = inv_13[37] ^ r_12[37] /*21361*/;
  assign sum_13[37] = _5998_ ^ _5997_ /*21360*/;
  assign _5999_ = _5998_ & _5997_ /*21359*/;
  assign _6000_ = inv_13[37] & r_12[37] /*21358*/;
  assign _6001_ = _5999_ | _6000_ /*21357*/;
  assign _6002_ = inv_13[38] ^ r_12[38] /*21355*/;
  assign sum_13[38] = _6002_ ^ _6001_ /*21354*/;
  assign _6003_ = _6002_ & _6001_ /*21353*/;
  assign _6004_ = inv_13[38] & r_12[38] /*21352*/;
  assign _6005_ = _6003_ | _6004_ /*21351*/;
  assign _6006_ = inv_13[39] ^ r_12[39] /*21349*/;
  assign sum_13[39] = _6006_ ^ _6005_ /*21348*/;
  assign _6007_ = _6006_ & _6005_ /*21347*/;
  assign _6008_ = inv_13[39] & r_12[39] /*21346*/;
  assign _6009_ = _6007_ | _6008_ /*21345*/;
  assign _6010_ = inv_13[40] ^ r_12[40] /*21343*/;
  assign sum_13[40] = _6010_ ^ _6009_ /*21342*/;
  assign _6011_ = _6010_ & _6009_ /*21341*/;
  assign _6012_ = inv_13[40] & r_12[40] /*21340*/;
  assign _6013_ = _6011_ | _6012_ /*21339*/;
  assign _6014_ = inv_13[41] ^ r_12[41] /*21337*/;
  assign sum_13[41] = _6014_ ^ _6013_ /*21336*/;
  assign _6015_ = _6014_ & _6013_ /*21335*/;
  assign _6016_ = inv_13[41] & r_12[41] /*21334*/;
  assign _6017_ = _6015_ | _6016_ /*21333*/;
  assign _6018_ = inv_13[42] ^ r_12[42] /*21331*/;
  assign sum_13[42] = _6018_ ^ _6017_ /*21330*/;
  assign _6019_ = _6018_ & _6017_ /*21329*/;
  assign _6020_ = inv_13[42] & r_12[42] /*21328*/;
  assign _6021_ = _6019_ | _6020_ /*21327*/;
  assign _6022_ = inv_13[43] ^ r_12[43] /*21325*/;
  assign sum_13[43] = _6022_ ^ _6021_ /*21324*/;
  assign _6023_ = _6022_ & _6021_ /*21323*/;
  assign _6024_ = inv_13[43] & r_12[43] /*21322*/;
  assign _6025_ = _6023_ | _6024_ /*21321*/;
  assign _6026_ = inv_13[44] ^ r_12[44] /*21319*/;
  assign sum_13[44] = _6026_ ^ _6025_ /*21318*/;
  assign _6027_ = _6026_ & _6025_ /*21317*/;
  assign _6028_ = inv_13[44] & r_12[44] /*21316*/;
  assign _6029_ = _6027_ | _6028_ /*21315*/;
  assign _6030_ = inv_13[45] ^ r_12[45] /*21313*/;
  assign sum_13[45] = _6030_ ^ _6029_ /*21312*/;
  assign _6031_ = _6030_ & _6029_ /*21311*/;
  assign _6032_ = inv_13[45] & r_12[45] /*21310*/;
  assign _6033_ = _6031_ | _6032_ /*21309*/;
  assign _6034_ = inv_13[46] ^ r_12[46] /*21307*/;
  assign sum_13[46] = _6034_ ^ _6033_ /*21306*/;
  assign _6035_ = _6034_ & _6033_ /*21305*/;
  assign _6036_ = inv_13[46] & r_12[46] /*21304*/;
  assign _6037_ = _6035_ | _6036_ /*21303*/;
  assign _6038_ = inv_13[47] ^ r_12[47] /*21301*/;
  assign sum_13[47] = _6038_ ^ _6037_ /*21300*/;
  assign _6039_ = _6038_ & _6037_ /*21299*/;
  assign _6040_ = inv_13[47] & r_12[47] /*21298*/;
  assign _6041_ = _6039_ | _6040_ /*21297*/;
  assign _6042_ = inv_13[48] ^ r_12[48] /*21295*/;
  assign sum_13[48] = _6042_ ^ _6041_ /*21294*/;
  assign _6043_ = _6042_ & _6041_ /*21293*/;
  assign _6044_ = inv_13[48] & r_12[48] /*21292*/;
  assign _6045_ = _6043_ | _6044_ /*21291*/;
  assign _6046_ = inv_13[49] ^ r_12[49] /*21289*/;
  assign sum_13[49] = _6046_ ^ _6045_ /*21288*/;
  assign _6047_ = _6046_ & _6045_ /*21287*/;
  assign _6048_ = inv_13[49] & r_12[49] /*21286*/;
  assign _6049_ = _6047_ | _6048_ /*21285*/;
  assign _6050_ = inv_13[50] ^ r_12[50] /*21283*/;
  assign sum_13[50] = _6050_ ^ _6049_ /*21282*/;
  assign _6051_ = _6050_ & _6049_ /*21281*/;
  assign _6052_ = inv_13[50] & r_12[50] /*21280*/;
  assign _6053_ = _6051_ | _6052_ /*21279*/;
  assign _6054_ = inv_13[51] ^ r_12[51] /*21277*/;
  assign sum_13[51] = _6054_ ^ _6053_ /*21276*/;
  assign _6055_ = _6054_ & _6053_ /*21275*/;
  assign _6056_ = inv_13[51] & r_12[51] /*21274*/;
  assign _6057_ = _6055_ | _6056_ /*21273*/;
  assign _6058_ = inv_13[52] ^ r_12[52] /*21271*/;
  assign sum_13[52] = _6058_ ^ _6057_ /*21270*/;
  assign _6059_ = _6058_ & _6057_ /*21269*/;
  assign _6060_ = inv_13[52] & r_12[52] /*21268*/;
  assign _6061_ = _6059_ | _6060_ /*21267*/;
  assign _6062_ = inv_13[53] ^ r_12[53] /*21265*/;
  assign sum_13[53] = _6062_ ^ _6061_ /*21264*/;
  assign _6063_ = _6062_ & _6061_ /*21263*/;
  assign _6064_ = inv_13[53] & r_12[53] /*21262*/;
  assign _6065_ = _6063_ | _6064_ /*21261*/;
  assign _6066_ = inv_13[54] ^ r_12[54] /*21259*/;
  assign sum_13[54] = _6066_ ^ _6065_ /*21258*/;
  assign _6067_ = _6066_ & _6065_ /*21257*/;
  assign _6068_ = inv_13[54] & r_12[54] /*21256*/;
  assign _6069_ = _6067_ | _6068_ /*21255*/;
  assign _6070_ = inv_13[55] ^ r_12[55] /*21253*/;
  assign sum_13[55] = _6070_ ^ _6069_ /*21252*/;
  assign _6071_ = _6070_ & _6069_ /*21251*/;
  assign _6072_ = inv_13[55] & r_12[55] /*21250*/;
  assign _6073_ = _6071_ | _6072_ /*21249*/;
  assign _6074_ = inv_13[56] ^ r_12[56] /*21247*/;
  assign sum_13[56] = _6074_ ^ _6073_ /*21246*/;
  assign _6075_ = _6074_ & _6073_ /*21245*/;
  assign _6076_ = inv_13[56] & r_12[56] /*21244*/;
  assign _6077_ = _6075_ | _6076_ /*21243*/;
  assign _6078_ = inv_13[57] ^ r_12[57] /*21241*/;
  assign sum_13[57] = _6078_ ^ _6077_ /*21240*/;
  assign _6079_ = _6078_ & _6077_ /*21239*/;
  assign _6080_ = inv_13[57] & r_12[57] /*21238*/;
  assign _6081_ = _6079_ | _6080_ /*21237*/;
  assign _6082_ = inv_13[58] ^ r_12[58] /*21235*/;
  assign sum_13[58] = _6082_ ^ _6081_ /*21234*/;
  assign _6083_ = _6082_ & _6081_ /*21233*/;
  assign _6084_ = inv_13[58] & r_12[58] /*21232*/;
  assign _6085_ = _6083_ | _6084_ /*21231*/;
  assign _6086_ = inv_13[59] ^ r_12[59] /*21229*/;
  assign sum_13[59] = _6086_ ^ _6085_ /*21228*/;
  assign _6087_ = _6086_ & _6085_ /*21227*/;
  assign _6088_ = inv_13[59] & r_12[59] /*21226*/;
  assign _6089_ = _6087_ | _6088_ /*21225*/;
  assign _6090_ = inv_13[60] ^ r_12[60] /*21223*/;
  assign sum_13[60] = _6090_ ^ _6089_ /*21222*/;
  assign _6091_ = _6090_ & _6089_ /*21221*/;
  assign _6092_ = inv_13[60] & r_12[60] /*21220*/;
  assign _6093_ = _6091_ | _6092_ /*21219*/;
  assign _6094_ = inv_13[61] ^ r_12[61] /*21217*/;
  assign sum_13[61] = _6094_ ^ _6093_ /*21216*/;
  assign _6095_ = _6094_ & _6093_ /*21215*/;
  assign _6096_ = inv_13[61] & r_12[61] /*21214*/;
  assign _6097_ = _6095_ | _6096_ /*21213*/;
  assign _6098_ = inv_13[62] ^ r_12[62] /*21211*/;
  assign sum_13[62] = _6098_ ^ _6097_ /*21210*/;
  assign _6099_ = _6098_ & _6097_ /*21209*/;
  assign _6100_ = inv_13[62] & r_12[62] /*21208*/;
  assign _6101_ = _6099_ | _6100_ /*21207*/;
  assign _6102_ = inv_13[63] ^ r_12[63] /*21205*/;
  assign sum_13[63] = _6102_ ^ _6101_ /*21204*/;
  assign _6103_ = _6102_ & _6101_ /*21203*/;
  assign _6104_ = inv_13[63] & r_12[63] /*21202*/;
  assign _6105_ = _6103_ | _6104_ /*21201*/;
  assign _6106_ = inv_13[64] ^ r_12[64] /*21199*/;
  assign sum_13[64] = _6106_ ^ _6105_ /*21198*/;
  assign _6107_ = _6106_ & _6105_ /*21197*/;
  assign _6108_ = inv_13[64] & r_12[64] /*21196*/;
  assign _6109_ = _6107_ | _6108_ /*21195*/;
  assign _6110_ = inv_13[65] ^ r_12[65] /*21193*/;
  assign sum_13[65] = _6110_ ^ _6109_ /*21192*/;
  assign _6111_ = _6110_ & _6109_ /*21191*/;
  assign _6112_ = inv_13[65] & r_12[65] /*21190*/;
  assign _6113_ = _6111_ | _6112_ /*21189*/;
  assign _6114_ = inv_13[66] ^ r_12[66] /*21187*/;
  assign sum_13[66] = _6114_ ^ _6113_ /*21186*/;
  assign _6115_ = _6114_ & _6113_ /*21185*/;
  assign _6116_ = inv_13[66] & r_12[66] /*21184*/;
  assign _6117_ = _6115_ | _6116_ /*21183*/;
  assign _6118_ = inv_13[67] ^ r_12[67] /*21181*/;
  assign sum_13[67] = _6118_ ^ _6117_ /*21180*/;
  assign _6119_ = _6118_ & _6117_ /*21179*/;
  assign _6120_ = inv_13[67] & r_12[67] /*21178*/;
  assign _6121_ = _6119_ | _6120_ /*21177*/;
  assign _6122_ = inv_13[68] ^ r_12[68] /*21175*/;
  assign sum_13[68] = _6122_ ^ _6121_ /*21174*/;
  assign _6123_ = _6122_ & _6121_ /*21173*/;
  assign _6124_ = inv_13[68] & r_12[68] /*21172*/;
  assign _6125_ = _6123_ | _6124_ /*21171*/;
  assign _6126_ = inv_13[69] ^ r_12[69] /*21169*/;
  assign sum_13[69] = _6126_ ^ _6125_ /*21168*/;
  assign _6127_ = _6126_ & _6125_ /*21167*/;
  assign _6128_ = inv_13[69] & r_12[69] /*21166*/;
  assign _6129_ = _6127_ | _6128_ /*21165*/;
  assign _6130_ = inv_13[70] ^ r_12[70] /*21163*/;
  assign sum_13[70] = _6130_ ^ _6129_ /*21162*/;
  assign _6131_ = _6130_ & _6129_ /*21161*/;
  assign _6132_ = inv_13[70] & r_12[70] /*21160*/;
  assign _6133_ = _6131_ | _6132_ /*21159*/;
  assign _6134_ = inv_13[71] ^ r_12[71] /*21157*/;
  assign sum_13[71] = _6134_ ^ _6133_ /*21156*/;
  assign _6135_ = _6134_ & _6133_ /*21155*/;
  assign _6136_ = inv_13[71] & r_12[71] /*21154*/;
  assign _6137_ = _6135_ | _6136_ /*21153*/;
  assign _6138_ = inv_13[72] ^ r_12[72] /*21151*/;
  assign sum_13[72] = _6138_ ^ _6137_ /*21150*/;
  assign _6139_ = _6138_ & _6137_ /*21149*/;
  assign _6140_ = inv_13[72] & r_12[72] /*21148*/;
  assign _6141_ = _6139_ | _6140_ /*21147*/;
  assign _6142_ = inv_13[73] ^ r_12[73] /*21145*/;
  assign sum_13[73] = _6142_ ^ _6141_ /*21144*/;
  assign _6143_ = _6142_ & _6141_ /*21143*/;
  assign _6144_ = inv_13[73] & r_12[73] /*21142*/;
  assign _6145_ = _6143_ | _6144_ /*21141*/;
  assign _6146_ = inv_13[74] ^ r_12[74] /*21139*/;
  assign sum_13[74] = _6146_ ^ _6145_ /*21138*/;
  assign _6147_ = _6146_ & _6145_ /*21137*/;
  assign _6148_ = inv_13[74] & r_12[74] /*21136*/;
  assign _6149_ = _6147_ | _6148_ /*21135*/;
  assign _6150_ = _6149_ ^ _6145_ /*21134*/;
  assign _6151_ = ~_6150_ /*21133*/;
  assign _6152_ = sum_13[74] & _6151_ /*21132*/;
  assign _6153_ = _6150_ & _6149_ /*21131*/;
  assign sum_13[75] = _6153_ | _6152_ /*21130*/;
  assign q[19] = ~sum_13[75] /*21129*/;
  assign m_13[0] = r_12[0] /*21128*/;
  assign m_13[1] = r_12[1] /*21127*/;
  assign m_13[2] = r_12[2] /*21126*/;
  assign m_13[3] = r_12[3] /*21125*/;
  assign m_13[4] = r_12[4] /*21124*/;
  assign m_13[5] = r_12[5] /*21123*/;
  assign m_13[6] = r_12[6] /*21122*/;
  assign m_13[7] = r_12[7] /*21121*/;
  assign m_13[8] = r_12[8] /*21120*/;
  assign m_13[9] = r_12[9] /*21119*/;
  assign m_13[10] = r_12[10] /*21118*/;
  assign m_13[11] = r_12[11] /*21117*/;
  assign m_13[12] = r_12[12] /*21116*/;
  assign m_13[13] = r_12[13] /*21115*/;
  assign m_13[14] = r_12[14] /*21114*/;
  assign m_13[15] = r_12[15] /*21113*/;
  assign m_13[16] = r_12[16] /*21112*/;
  assign m_13[17] = r_12[17] /*21111*/;
  assign m_13[18] = r_12[18] /*21110*/;
  assign m_13[19] = r_12[19] /*21109*/;
  assign m_13[20] = r_12[20] /*21108*/;
  assign m_13[21] = r_12[21] /*21107*/;
  assign m_13[22] = r_12[22] /*21106*/;
  assign m_13[23] = r_12[23] /*21105*/;
  assign m_13[24] = r_12[24] /*21104*/;
  assign m_13[25] = r_12[25] /*21103*/;
  assign m_13[26] = r_12[26] /*21102*/;
  assign m_13[27] = r_12[27] /*21101*/;
  assign m_13[28] = r_12[28] /*21100*/;
  assign m_13[29] = r_12[29] /*21099*/;
  assign m_13[30] = r_12[30] /*21098*/;
  assign m_13[31] = r_12[31] /*21097*/;
  assign m_13[32] = r_12[32] /*21096*/;
  assign m_13[33] = r_12[33] /*21095*/;
  assign m_13[34] = r_12[34] /*21094*/;
  assign m_13[35] = r_12[35] /*21093*/;
  assign m_13[36] = r_12[36] /*21092*/;
  assign m_13[37] = r_12[37] /*21091*/;
  assign m_13[38] = r_12[38] /*21090*/;
  assign m_13[39] = r_12[39] /*21089*/;
  assign m_13[40] = r_12[40] /*21088*/;
  assign m_13[41] = r_12[41] /*21087*/;
  assign m_13[42] = r_12[42] /*21086*/;
  assign m_13[43] = r_12[43] /*21085*/;
  assign m_13[44] = r_12[44] /*21084*/;
  assign m_13[45] = r_12[45] /*21083*/;
  assign m_13[46] = r_12[46] /*21082*/;
  assign m_13[47] = r_12[47] /*21081*/;
  assign m_13[48] = r_12[48] /*21080*/;
  assign m_13[49] = r_12[49] /*21079*/;
  assign m_13[50] = r_12[50] /*21078*/;
  assign m_13[51] = r_12[51] /*21077*/;
  assign m_13[52] = r_12[52] /*21076*/;
  assign m_13[53] = r_12[53] /*21075*/;
  assign m_13[54] = r_12[54] /*21074*/;
  assign m_13[55] = r_12[55] /*21073*/;
  assign m_13[56] = r_12[56] /*21072*/;
  assign m_13[57] = r_12[57] /*21071*/;
  assign m_13[58] = r_12[58] /*21070*/;
  assign m_13[59] = r_12[59] /*21069*/;
  assign m_13[60] = r_12[60] /*21068*/;
  assign m_13[61] = r_12[61] /*21067*/;
  assign m_13[62] = r_12[62] /*21066*/;
  assign m_13[63] = r_12[63] /*21065*/;
  assign m_13[64] = r_12[64] /*21064*/;
  assign m_13[65] = r_12[65] /*21063*/;
  assign m_13[66] = r_12[66] /*21062*/;
  assign m_13[67] = r_12[67] /*21061*/;
  assign m_13[68] = r_12[68] /*21060*/;
  assign m_13[69] = r_12[69] /*21059*/;
  assign m_13[70] = r_12[70] /*21058*/;
  assign m_13[71] = r_12[71] /*21057*/;
  assign m_13[72] = r_12[72] /*21056*/;
  assign m_13[73] = r_12[73] /*21055*/;
  assign m_13[74] = r_12[74] /*21054*/;
  assign m_13[75] = r_12[74] /*21053*/;
  assign _6155_ = ~q[19] /*21052*/;
  assign _6156_ = sum_13[0] & q[19] /*21051*/;
  assign _6157_ = m_13[0] & _6155_ /*21050*/;
  assign r_13[0] = _6157_ | _6156_ /*21049*/;
  assign _6158_ = ~q[19] /*21048*/;
  assign _6159_ = sum_13[1] & q[19] /*21047*/;
  assign _6160_ = m_13[1] & _6158_ /*21046*/;
  assign r_13[1] = _6160_ | _6159_ /*21045*/;
  assign _6161_ = ~q[19] /*21044*/;
  assign _6162_ = sum_13[2] & q[19] /*21043*/;
  assign _6163_ = m_13[2] & _6161_ /*21042*/;
  assign r_13[2] = _6163_ | _6162_ /*21041*/;
  assign _6164_ = ~q[19] /*21040*/;
  assign _6165_ = sum_13[3] & q[19] /*21039*/;
  assign _6166_ = m_13[3] & _6164_ /*21038*/;
  assign r_13[3] = _6166_ | _6165_ /*21037*/;
  assign _6167_ = ~q[19] /*21036*/;
  assign _6168_ = sum_13[4] & q[19] /*21035*/;
  assign _6169_ = m_13[4] & _6167_ /*21034*/;
  assign r_13[4] = _6169_ | _6168_ /*21033*/;
  assign _6170_ = ~q[19] /*21032*/;
  assign _6171_ = sum_13[5] & q[19] /*21031*/;
  assign _6172_ = m_13[5] & _6170_ /*21030*/;
  assign r_13[5] = _6172_ | _6171_ /*21029*/;
  assign _6173_ = ~q[19] /*21028*/;
  assign _6174_ = sum_13[6] & q[19] /*21027*/;
  assign _6175_ = m_13[6] & _6173_ /*21026*/;
  assign r_13[6] = _6175_ | _6174_ /*21025*/;
  assign _6176_ = ~q[19] /*21024*/;
  assign _6177_ = sum_13[7] & q[19] /*21023*/;
  assign _6178_ = m_13[7] & _6176_ /*21022*/;
  assign r_13[7] = _6178_ | _6177_ /*21021*/;
  assign _6179_ = ~q[19] /*21020*/;
  assign _6180_ = sum_13[8] & q[19] /*21019*/;
  assign _6181_ = m_13[8] & _6179_ /*21018*/;
  assign r_13[8] = _6181_ | _6180_ /*21017*/;
  assign _6182_ = ~q[19] /*21016*/;
  assign _6183_ = sum_13[9] & q[19] /*21015*/;
  assign _6184_ = m_13[9] & _6182_ /*21014*/;
  assign r_13[9] = _6184_ | _6183_ /*21013*/;
  assign _6185_ = ~q[19] /*21012*/;
  assign _6186_ = sum_13[10] & q[19] /*21011*/;
  assign _6187_ = m_13[10] & _6185_ /*21010*/;
  assign r_13[10] = _6187_ | _6186_ /*21009*/;
  assign _6188_ = ~q[19] /*21008*/;
  assign _6189_ = sum_13[11] & q[19] /*21007*/;
  assign _6190_ = m_13[11] & _6188_ /*21006*/;
  assign r_13[11] = _6190_ | _6189_ /*21005*/;
  assign _6191_ = ~q[19] /*21004*/;
  assign _6192_ = sum_13[12] & q[19] /*21003*/;
  assign _6193_ = m_13[12] & _6191_ /*21002*/;
  assign r_13[12] = _6193_ | _6192_ /*21001*/;
  assign _6194_ = ~q[19] /*21000*/;
  assign _6195_ = sum_13[13] & q[19] /*20999*/;
  assign _6196_ = m_13[13] & _6194_ /*20998*/;
  assign r_13[13] = _6196_ | _6195_ /*20997*/;
  assign _6197_ = ~q[19] /*20996*/;
  assign _6198_ = sum_13[14] & q[19] /*20995*/;
  assign _6199_ = m_13[14] & _6197_ /*20994*/;
  assign r_13[14] = _6199_ | _6198_ /*20993*/;
  assign _6200_ = ~q[19] /*20992*/;
  assign _6201_ = sum_13[15] & q[19] /*20991*/;
  assign _6202_ = m_13[15] & _6200_ /*20990*/;
  assign r_13[15] = _6202_ | _6201_ /*20989*/;
  assign _6203_ = ~q[19] /*20988*/;
  assign _6204_ = sum_13[16] & q[19] /*20987*/;
  assign _6205_ = m_13[16] & _6203_ /*20986*/;
  assign r_13[16] = _6205_ | _6204_ /*20985*/;
  assign _6206_ = ~q[19] /*20984*/;
  assign _6207_ = sum_13[17] & q[19] /*20983*/;
  assign _6208_ = m_13[17] & _6206_ /*20982*/;
  assign r_13[17] = _6208_ | _6207_ /*20981*/;
  assign _6209_ = ~q[19] /*20980*/;
  assign _6210_ = sum_13[18] & q[19] /*20979*/;
  assign _6211_ = m_13[18] & _6209_ /*20978*/;
  assign r_13[18] = _6211_ | _6210_ /*20977*/;
  assign _6212_ = ~q[19] /*20976*/;
  assign _6213_ = sum_13[19] & q[19] /*20975*/;
  assign _6214_ = m_13[19] & _6212_ /*20974*/;
  assign r_13[19] = _6214_ | _6213_ /*20973*/;
  assign _6215_ = ~q[19] /*20972*/;
  assign _6216_ = sum_13[20] & q[19] /*20971*/;
  assign _6217_ = m_13[20] & _6215_ /*20970*/;
  assign r_13[20] = _6217_ | _6216_ /*20969*/;
  assign _6218_ = ~q[19] /*20968*/;
  assign _6219_ = sum_13[21] & q[19] /*20967*/;
  assign _6220_ = m_13[21] & _6218_ /*20966*/;
  assign r_13[21] = _6220_ | _6219_ /*20965*/;
  assign _6221_ = ~q[19] /*20964*/;
  assign _6222_ = sum_13[22] & q[19] /*20963*/;
  assign _6223_ = m_13[22] & _6221_ /*20962*/;
  assign r_13[22] = _6223_ | _6222_ /*20961*/;
  assign _6224_ = ~q[19] /*20960*/;
  assign _6225_ = sum_13[23] & q[19] /*20959*/;
  assign _6226_ = m_13[23] & _6224_ /*20958*/;
  assign r_13[23] = _6226_ | _6225_ /*20957*/;
  assign _6227_ = ~q[19] /*20956*/;
  assign _6228_ = sum_13[24] & q[19] /*20955*/;
  assign _6229_ = m_13[24] & _6227_ /*20954*/;
  assign r_13[24] = _6229_ | _6228_ /*20953*/;
  assign _6230_ = ~q[19] /*20952*/;
  assign _6231_ = sum_13[25] & q[19] /*20951*/;
  assign _6232_ = m_13[25] & _6230_ /*20950*/;
  assign r_13[25] = _6232_ | _6231_ /*20949*/;
  assign _6233_ = ~q[19] /*20948*/;
  assign _6234_ = sum_13[26] & q[19] /*20947*/;
  assign _6235_ = m_13[26] & _6233_ /*20946*/;
  assign r_13[26] = _6235_ | _6234_ /*20945*/;
  assign _6236_ = ~q[19] /*20944*/;
  assign _6237_ = sum_13[27] & q[19] /*20943*/;
  assign _6238_ = m_13[27] & _6236_ /*20942*/;
  assign r_13[27] = _6238_ | _6237_ /*20941*/;
  assign _6239_ = ~q[19] /*20940*/;
  assign _6240_ = sum_13[28] & q[19] /*20939*/;
  assign _6241_ = m_13[28] & _6239_ /*20938*/;
  assign r_13[28] = _6241_ | _6240_ /*20937*/;
  assign _6242_ = ~q[19] /*20936*/;
  assign _6243_ = sum_13[29] & q[19] /*20935*/;
  assign _6244_ = m_13[29] & _6242_ /*20934*/;
  assign r_13[29] = _6244_ | _6243_ /*20933*/;
  assign _6245_ = ~q[19] /*20932*/;
  assign _6246_ = sum_13[30] & q[19] /*20931*/;
  assign _6247_ = m_13[30] & _6245_ /*20930*/;
  assign r_13[30] = _6247_ | _6246_ /*20929*/;
  assign _6248_ = ~q[19] /*20928*/;
  assign _6249_ = sum_13[31] & q[19] /*20927*/;
  assign _6250_ = m_13[31] & _6248_ /*20926*/;
  assign r_13[31] = _6250_ | _6249_ /*20925*/;
  assign _6251_ = ~q[19] /*20924*/;
  assign _6252_ = sum_13[32] & q[19] /*20923*/;
  assign _6253_ = m_13[32] & _6251_ /*20922*/;
  assign r_13[32] = _6253_ | _6252_ /*20921*/;
  assign _6254_ = ~q[19] /*20920*/;
  assign _6255_ = sum_13[33] & q[19] /*20919*/;
  assign _6256_ = m_13[33] & _6254_ /*20918*/;
  assign r_13[33] = _6256_ | _6255_ /*20917*/;
  assign _6257_ = ~q[19] /*20916*/;
  assign _6258_ = sum_13[34] & q[19] /*20915*/;
  assign _6259_ = m_13[34] & _6257_ /*20914*/;
  assign r_13[34] = _6259_ | _6258_ /*20913*/;
  assign _6260_ = ~q[19] /*20912*/;
  assign _6261_ = sum_13[35] & q[19] /*20911*/;
  assign _6262_ = m_13[35] & _6260_ /*20910*/;
  assign r_13[35] = _6262_ | _6261_ /*20909*/;
  assign _6263_ = ~q[19] /*20908*/;
  assign _6264_ = sum_13[36] & q[19] /*20907*/;
  assign _6265_ = m_13[36] & _6263_ /*20906*/;
  assign r_13[36] = _6265_ | _6264_ /*20905*/;
  assign _6266_ = ~q[19] /*20904*/;
  assign _6267_ = sum_13[37] & q[19] /*20903*/;
  assign _6268_ = m_13[37] & _6266_ /*20902*/;
  assign r_13[37] = _6268_ | _6267_ /*20901*/;
  assign _6269_ = ~q[19] /*20900*/;
  assign _6270_ = sum_13[38] & q[19] /*20899*/;
  assign _6271_ = m_13[38] & _6269_ /*20898*/;
  assign r_13[38] = _6271_ | _6270_ /*20897*/;
  assign _6272_ = ~q[19] /*20896*/;
  assign _6273_ = sum_13[39] & q[19] /*20895*/;
  assign _6274_ = m_13[39] & _6272_ /*20894*/;
  assign r_13[39] = _6274_ | _6273_ /*20893*/;
  assign _6275_ = ~q[19] /*20892*/;
  assign _6276_ = sum_13[40] & q[19] /*20891*/;
  assign _6277_ = m_13[40] & _6275_ /*20890*/;
  assign r_13[40] = _6277_ | _6276_ /*20889*/;
  assign _6278_ = ~q[19] /*20888*/;
  assign _6279_ = sum_13[41] & q[19] /*20887*/;
  assign _6280_ = m_13[41] & _6278_ /*20886*/;
  assign r_13[41] = _6280_ | _6279_ /*20885*/;
  assign _6281_ = ~q[19] /*20884*/;
  assign _6282_ = sum_13[42] & q[19] /*20883*/;
  assign _6283_ = m_13[42] & _6281_ /*20882*/;
  assign r_13[42] = _6283_ | _6282_ /*20881*/;
  assign _6284_ = ~q[19] /*20880*/;
  assign _6285_ = sum_13[43] & q[19] /*20879*/;
  assign _6286_ = m_13[43] & _6284_ /*20878*/;
  assign r_13[43] = _6286_ | _6285_ /*20877*/;
  assign _6287_ = ~q[19] /*20876*/;
  assign _6288_ = sum_13[44] & q[19] /*20875*/;
  assign _6289_ = m_13[44] & _6287_ /*20874*/;
  assign r_13[44] = _6289_ | _6288_ /*20873*/;
  assign _6290_ = ~q[19] /*20872*/;
  assign _6291_ = sum_13[45] & q[19] /*20871*/;
  assign _6292_ = m_13[45] & _6290_ /*20870*/;
  assign r_13[45] = _6292_ | _6291_ /*20869*/;
  assign _6293_ = ~q[19] /*20868*/;
  assign _6294_ = sum_13[46] & q[19] /*20867*/;
  assign _6295_ = m_13[46] & _6293_ /*20866*/;
  assign r_13[46] = _6295_ | _6294_ /*20865*/;
  assign _6296_ = ~q[19] /*20864*/;
  assign _6297_ = sum_13[47] & q[19] /*20863*/;
  assign _6298_ = m_13[47] & _6296_ /*20862*/;
  assign r_13[47] = _6298_ | _6297_ /*20861*/;
  assign _6299_ = ~q[19] /*20860*/;
  assign _6300_ = sum_13[48] & q[19] /*20859*/;
  assign _6301_ = m_13[48] & _6299_ /*20858*/;
  assign r_13[48] = _6301_ | _6300_ /*20857*/;
  assign _6302_ = ~q[19] /*20856*/;
  assign _6303_ = sum_13[49] & q[19] /*20855*/;
  assign _6304_ = m_13[49] & _6302_ /*20854*/;
  assign r_13[49] = _6304_ | _6303_ /*20853*/;
  assign _6305_ = ~q[19] /*20852*/;
  assign _6306_ = sum_13[50] & q[19] /*20851*/;
  assign _6307_ = m_13[50] & _6305_ /*20850*/;
  assign r_13[50] = _6307_ | _6306_ /*20849*/;
  assign _6308_ = ~q[19] /*20848*/;
  assign _6309_ = sum_13[51] & q[19] /*20847*/;
  assign _6310_ = m_13[51] & _6308_ /*20846*/;
  assign r_13[51] = _6310_ | _6309_ /*20845*/;
  assign _6311_ = ~q[19] /*20844*/;
  assign _6312_ = sum_13[52] & q[19] /*20843*/;
  assign _6313_ = m_13[52] & _6311_ /*20842*/;
  assign r_13[52] = _6313_ | _6312_ /*20841*/;
  assign _6314_ = ~q[19] /*20840*/;
  assign _6315_ = sum_13[53] & q[19] /*20839*/;
  assign _6316_ = m_13[53] & _6314_ /*20838*/;
  assign r_13[53] = _6316_ | _6315_ /*20837*/;
  assign _6317_ = ~q[19] /*20836*/;
  assign _6318_ = sum_13[54] & q[19] /*20835*/;
  assign _6319_ = m_13[54] & _6317_ /*20834*/;
  assign r_13[54] = _6319_ | _6318_ /*20833*/;
  assign _6320_ = ~q[19] /*20832*/;
  assign _6321_ = sum_13[55] & q[19] /*20831*/;
  assign _6322_ = m_13[55] & _6320_ /*20830*/;
  assign r_13[55] = _6322_ | _6321_ /*20829*/;
  assign _6323_ = ~q[19] /*20828*/;
  assign _6324_ = sum_13[56] & q[19] /*20827*/;
  assign _6325_ = m_13[56] & _6323_ /*20826*/;
  assign r_13[56] = _6325_ | _6324_ /*20825*/;
  assign _6326_ = ~q[19] /*20824*/;
  assign _6327_ = sum_13[57] & q[19] /*20823*/;
  assign _6328_ = m_13[57] & _6326_ /*20822*/;
  assign r_13[57] = _6328_ | _6327_ /*20821*/;
  assign _6329_ = ~q[19] /*20820*/;
  assign _6330_ = sum_13[58] & q[19] /*20819*/;
  assign _6331_ = m_13[58] & _6329_ /*20818*/;
  assign r_13[58] = _6331_ | _6330_ /*20817*/;
  assign _6332_ = ~q[19] /*20816*/;
  assign _6333_ = sum_13[59] & q[19] /*20815*/;
  assign _6334_ = m_13[59] & _6332_ /*20814*/;
  assign r_13[59] = _6334_ | _6333_ /*20813*/;
  assign _6335_ = ~q[19] /*20812*/;
  assign _6336_ = sum_13[60] & q[19] /*20811*/;
  assign _6337_ = m_13[60] & _6335_ /*20810*/;
  assign r_13[60] = _6337_ | _6336_ /*20809*/;
  assign _6338_ = ~q[19] /*20808*/;
  assign _6339_ = sum_13[61] & q[19] /*20807*/;
  assign _6340_ = m_13[61] & _6338_ /*20806*/;
  assign r_13[61] = _6340_ | _6339_ /*20805*/;
  assign _6341_ = ~q[19] /*20804*/;
  assign _6342_ = sum_13[62] & q[19] /*20803*/;
  assign _6343_ = m_13[62] & _6341_ /*20802*/;
  assign r_13[62] = _6343_ | _6342_ /*20801*/;
  assign _6344_ = ~q[19] /*20800*/;
  assign _6345_ = sum_13[63] & q[19] /*20799*/;
  assign _6346_ = m_13[63] & _6344_ /*20798*/;
  assign r_13[63] = _6346_ | _6345_ /*20797*/;
  assign _6347_ = ~q[19] /*20796*/;
  assign _6348_ = sum_13[64] & q[19] /*20795*/;
  assign _6349_ = m_13[64] & _6347_ /*20794*/;
  assign r_13[64] = _6349_ | _6348_ /*20793*/;
  assign _6350_ = ~q[19] /*20792*/;
  assign _6351_ = sum_13[65] & q[19] /*20791*/;
  assign _6352_ = m_13[65] & _6350_ /*20790*/;
  assign r_13[65] = _6352_ | _6351_ /*20789*/;
  assign _6353_ = ~q[19] /*20788*/;
  assign _6354_ = sum_13[66] & q[19] /*20787*/;
  assign _6355_ = m_13[66] & _6353_ /*20786*/;
  assign r_13[66] = _6355_ | _6354_ /*20785*/;
  assign _6356_ = ~q[19] /*20784*/;
  assign _6357_ = sum_13[67] & q[19] /*20783*/;
  assign _6358_ = m_13[67] & _6356_ /*20782*/;
  assign r_13[67] = _6358_ | _6357_ /*20781*/;
  assign _6359_ = ~q[19] /*20780*/;
  assign _6360_ = sum_13[68] & q[19] /*20779*/;
  assign _6361_ = m_13[68] & _6359_ /*20778*/;
  assign r_13[68] = _6361_ | _6360_ /*20777*/;
  assign _6362_ = ~q[19] /*20776*/;
  assign _6363_ = sum_13[69] & q[19] /*20775*/;
  assign _6364_ = m_13[69] & _6362_ /*20774*/;
  assign r_13[69] = _6364_ | _6363_ /*20773*/;
  assign _6365_ = ~q[19] /*20772*/;
  assign _6366_ = sum_13[70] & q[19] /*20771*/;
  assign _6367_ = m_13[70] & _6365_ /*20770*/;
  assign r_13[70] = _6367_ | _6366_ /*20769*/;
  assign _6368_ = ~q[19] /*20768*/;
  assign _6369_ = sum_13[71] & q[19] /*20767*/;
  assign _6370_ = m_13[71] & _6368_ /*20766*/;
  assign r_13[71] = _6370_ | _6369_ /*20765*/;
  assign _6371_ = ~q[19] /*20764*/;
  assign _6372_ = sum_13[72] & q[19] /*20763*/;
  assign _6373_ = m_13[72] & _6371_ /*20762*/;
  assign r_13[72] = _6373_ | _6372_ /*20761*/;
  assign _6374_ = ~q[19] /*20760*/;
  assign _6375_ = sum_13[73] & q[19] /*20759*/;
  assign _6376_ = m_13[73] & _6374_ /*20758*/;
  assign r_13[73] = _6376_ | _6375_ /*20757*/;
  assign _6377_ = ~q[19] /*20756*/;
  assign _6378_ = sum_13[74] & q[19] /*20755*/;
  assign _6379_ = m_13[74] & _6377_ /*20754*/;
  assign r_13[74] = _6379_ | _6378_ /*20753*/;
  assign _6380_ = ~q[19] /*20752*/;
  assign _6381_ = sum_13[75] & q[19] /*20751*/;
  assign _6382_ = m_13[75] & _6380_ /*20750*/;
  assign r_13[75] = _6382_ | _6381_ /*20749*/;
  assign inv_14[0] = oneWire /*20508*/;
  assign inv_14[1] = oneWire /*20502*/;
  assign inv_14[2] = oneWire /*20496*/;
  assign inv_14[3] = oneWire /*20490*/;
  assign inv_14[4] = oneWire /*20484*/;
  assign inv_14[5] = oneWire /*20478*/;
  assign inv_14[6] = oneWire /*20472*/;
  assign inv_14[7] = oneWire /*20466*/;
  assign inv_14[8] = oneWire /*20460*/;
  assign inv_14[9] = oneWire /*20454*/;
  assign inv_14[10] = oneWire /*20448*/;
  assign inv_14[11] = oneWire /*20442*/;
  assign inv_14[12] = oneWire /*20436*/;
  assign inv_14[13] = oneWire /*20430*/;
  assign inv_14[14] = oneWire /*20424*/;
  assign inv_14[15] = oneWire /*20418*/;
  assign inv_14[16] = oneWire /*20412*/;
  assign inv_14[17] = oneWire /*20406*/;
  assign inv_14[18] = ~div[0] /*20400*/;
  assign inv_14[19] = ~div[1] /*20394*/;
  assign inv_14[20] = ~div[2] /*20388*/;
  assign inv_14[21] = ~div[3] /*20382*/;
  assign inv_14[22] = ~div[4] /*20376*/;
  assign inv_14[23] = ~div[5] /*20370*/;
  assign inv_14[24] = ~div[6] /*20364*/;
  assign inv_14[25] = ~div[7] /*20358*/;
  assign inv_14[26] = ~div[8] /*20352*/;
  assign inv_14[27] = ~div[9] /*20346*/;
  assign inv_14[28] = ~div[10] /*20340*/;
  assign inv_14[29] = ~div[11] /*20334*/;
  assign inv_14[30] = ~div[12] /*20328*/;
  assign inv_14[31] = ~div[13] /*20322*/;
  assign inv_14[32] = ~div[14] /*20316*/;
  assign inv_14[33] = ~div[15] /*20310*/;
  assign inv_14[34] = ~div[16] /*20304*/;
  assign inv_14[35] = ~div[17] /*20298*/;
  assign inv_14[36] = ~div[18] /*20292*/;
  assign inv_14[37] = ~div[19] /*20286*/;
  assign inv_14[38] = ~div[20] /*20280*/;
  assign inv_14[39] = ~div[21] /*20274*/;
  assign inv_14[40] = ~div[22] /*20268*/;
  assign inv_14[41] = ~div[23] /*20262*/;
  assign inv_14[42] = ~div[24] /*20256*/;
  assign inv_14[43] = ~div[25] /*20250*/;
  assign inv_14[44] = ~div[26] /*20244*/;
  assign inv_14[45] = ~div[27] /*20238*/;
  assign inv_14[46] = ~div[28] /*20232*/;
  assign inv_14[47] = ~div[29] /*20226*/;
  assign inv_14[48] = ~div[30] /*20220*/;
  assign inv_14[49] = oneWire /*20214*/;
  assign inv_14[50] = oneWire /*20208*/;
  assign inv_14[51] = oneWire /*20202*/;
  assign inv_14[52] = oneWire /*20196*/;
  assign inv_14[53] = oneWire /*20190*/;
  assign inv_14[54] = oneWire /*20184*/;
  assign inv_14[55] = oneWire /*20178*/;
  assign inv_14[56] = oneWire /*20172*/;
  assign inv_14[57] = oneWire /*20166*/;
  assign inv_14[58] = oneWire /*20160*/;
  assign inv_14[59] = oneWire /*20154*/;
  assign inv_14[60] = oneWire /*20148*/;
  assign inv_14[61] = oneWire /*20142*/;
  assign inv_14[62] = oneWire /*20136*/;
  assign inv_14[63] = oneWire /*20130*/;
  assign inv_14[64] = oneWire /*20124*/;
  assign inv_14[65] = oneWire /*20118*/;
  assign inv_14[66] = oneWire /*20112*/;
  assign inv_14[67] = oneWire /*20106*/;
  assign inv_14[68] = oneWire /*20100*/;
  assign inv_14[69] = oneWire /*20094*/;
  assign inv_14[70] = oneWire /*20088*/;
  assign inv_14[71] = oneWire /*20082*/;
  assign inv_14[72] = oneWire /*20076*/;
  assign inv_14[73] = oneWire /*20070*/;
  assign inv_14[74] = oneWire /*20064*/;
  assign inv_14[75] = oneWire /*20058*/;
  assign _6383_ = inv_14[0] ^ r_13[0] /*20507*/;
  assign sum_14[0] = _6383_ ^ oneWire /*20506*/;
  assign _6384_ = _6383_ & oneWire /*20505*/;
  assign _6385_ = inv_14[0] & r_13[0] /*20504*/;
  assign _6386_ = _6384_ | _6385_ /*20503*/;
  assign _6387_ = inv_14[1] ^ r_13[1] /*20501*/;
  assign sum_14[1] = _6387_ ^ _6386_ /*20500*/;
  assign _6388_ = _6387_ & _6386_ /*20499*/;
  assign _6389_ = inv_14[1] & r_13[1] /*20498*/;
  assign _6390_ = _6388_ | _6389_ /*20497*/;
  assign _6391_ = inv_14[2] ^ r_13[2] /*20495*/;
  assign sum_14[2] = _6391_ ^ _6390_ /*20494*/;
  assign _6392_ = _6391_ & _6390_ /*20493*/;
  assign _6393_ = inv_14[2] & r_13[2] /*20492*/;
  assign _6394_ = _6392_ | _6393_ /*20491*/;
  assign _6395_ = inv_14[3] ^ r_13[3] /*20489*/;
  assign sum_14[3] = _6395_ ^ _6394_ /*20488*/;
  assign _6396_ = _6395_ & _6394_ /*20487*/;
  assign _6397_ = inv_14[3] & r_13[3] /*20486*/;
  assign _6398_ = _6396_ | _6397_ /*20485*/;
  assign _6399_ = inv_14[4] ^ r_13[4] /*20483*/;
  assign sum_14[4] = _6399_ ^ _6398_ /*20482*/;
  assign _6400_ = _6399_ & _6398_ /*20481*/;
  assign _6401_ = inv_14[4] & r_13[4] /*20480*/;
  assign _6402_ = _6400_ | _6401_ /*20479*/;
  assign _6403_ = inv_14[5] ^ r_13[5] /*20477*/;
  assign sum_14[5] = _6403_ ^ _6402_ /*20476*/;
  assign _6404_ = _6403_ & _6402_ /*20475*/;
  assign _6405_ = inv_14[5] & r_13[5] /*20474*/;
  assign _6406_ = _6404_ | _6405_ /*20473*/;
  assign _6407_ = inv_14[6] ^ r_13[6] /*20471*/;
  assign sum_14[6] = _6407_ ^ _6406_ /*20470*/;
  assign _6408_ = _6407_ & _6406_ /*20469*/;
  assign _6409_ = inv_14[6] & r_13[6] /*20468*/;
  assign _6410_ = _6408_ | _6409_ /*20467*/;
  assign _6411_ = inv_14[7] ^ r_13[7] /*20465*/;
  assign sum_14[7] = _6411_ ^ _6410_ /*20464*/;
  assign _6412_ = _6411_ & _6410_ /*20463*/;
  assign _6413_ = inv_14[7] & r_13[7] /*20462*/;
  assign _6414_ = _6412_ | _6413_ /*20461*/;
  assign _6415_ = inv_14[8] ^ r_13[8] /*20459*/;
  assign sum_14[8] = _6415_ ^ _6414_ /*20458*/;
  assign _6416_ = _6415_ & _6414_ /*20457*/;
  assign _6417_ = inv_14[8] & r_13[8] /*20456*/;
  assign _6418_ = _6416_ | _6417_ /*20455*/;
  assign _6419_ = inv_14[9] ^ r_13[9] /*20453*/;
  assign sum_14[9] = _6419_ ^ _6418_ /*20452*/;
  assign _6420_ = _6419_ & _6418_ /*20451*/;
  assign _6421_ = inv_14[9] & r_13[9] /*20450*/;
  assign _6422_ = _6420_ | _6421_ /*20449*/;
  assign _6423_ = inv_14[10] ^ r_13[10] /*20447*/;
  assign sum_14[10] = _6423_ ^ _6422_ /*20446*/;
  assign _6424_ = _6423_ & _6422_ /*20445*/;
  assign _6425_ = inv_14[10] & r_13[10] /*20444*/;
  assign _6426_ = _6424_ | _6425_ /*20443*/;
  assign _6427_ = inv_14[11] ^ r_13[11] /*20441*/;
  assign sum_14[11] = _6427_ ^ _6426_ /*20440*/;
  assign _6428_ = _6427_ & _6426_ /*20439*/;
  assign _6429_ = inv_14[11] & r_13[11] /*20438*/;
  assign _6430_ = _6428_ | _6429_ /*20437*/;
  assign _6431_ = inv_14[12] ^ r_13[12] /*20435*/;
  assign sum_14[12] = _6431_ ^ _6430_ /*20434*/;
  assign _6432_ = _6431_ & _6430_ /*20433*/;
  assign _6433_ = inv_14[12] & r_13[12] /*20432*/;
  assign _6434_ = _6432_ | _6433_ /*20431*/;
  assign _6435_ = inv_14[13] ^ r_13[13] /*20429*/;
  assign sum_14[13] = _6435_ ^ _6434_ /*20428*/;
  assign _6436_ = _6435_ & _6434_ /*20427*/;
  assign _6437_ = inv_14[13] & r_13[13] /*20426*/;
  assign _6438_ = _6436_ | _6437_ /*20425*/;
  assign _6439_ = inv_14[14] ^ r_13[14] /*20423*/;
  assign sum_14[14] = _6439_ ^ _6438_ /*20422*/;
  assign _6440_ = _6439_ & _6438_ /*20421*/;
  assign _6441_ = inv_14[14] & r_13[14] /*20420*/;
  assign _6442_ = _6440_ | _6441_ /*20419*/;
  assign _6443_ = inv_14[15] ^ r_13[15] /*20417*/;
  assign sum_14[15] = _6443_ ^ _6442_ /*20416*/;
  assign _6444_ = _6443_ & _6442_ /*20415*/;
  assign _6445_ = inv_14[15] & r_13[15] /*20414*/;
  assign _6446_ = _6444_ | _6445_ /*20413*/;
  assign _6447_ = inv_14[16] ^ r_13[16] /*20411*/;
  assign sum_14[16] = _6447_ ^ _6446_ /*20410*/;
  assign _6448_ = _6447_ & _6446_ /*20409*/;
  assign _6449_ = inv_14[16] & r_13[16] /*20408*/;
  assign _6450_ = _6448_ | _6449_ /*20407*/;
  assign _6451_ = inv_14[17] ^ r_13[17] /*20405*/;
  assign sum_14[17] = _6451_ ^ _6450_ /*20404*/;
  assign _6452_ = _6451_ & _6450_ /*20403*/;
  assign _6453_ = inv_14[17] & r_13[17] /*20402*/;
  assign _6454_ = _6452_ | _6453_ /*20401*/;
  assign _6455_ = inv_14[18] ^ r_13[18] /*20399*/;
  assign sum_14[18] = _6455_ ^ _6454_ /*20398*/;
  assign _6456_ = _6455_ & _6454_ /*20397*/;
  assign _6457_ = inv_14[18] & r_13[18] /*20396*/;
  assign _6458_ = _6456_ | _6457_ /*20395*/;
  assign _6459_ = inv_14[19] ^ r_13[19] /*20393*/;
  assign sum_14[19] = _6459_ ^ _6458_ /*20392*/;
  assign _6460_ = _6459_ & _6458_ /*20391*/;
  assign _6461_ = inv_14[19] & r_13[19] /*20390*/;
  assign _6462_ = _6460_ | _6461_ /*20389*/;
  assign _6463_ = inv_14[20] ^ r_13[20] /*20387*/;
  assign sum_14[20] = _6463_ ^ _6462_ /*20386*/;
  assign _6464_ = _6463_ & _6462_ /*20385*/;
  assign _6465_ = inv_14[20] & r_13[20] /*20384*/;
  assign _6466_ = _6464_ | _6465_ /*20383*/;
  assign _6467_ = inv_14[21] ^ r_13[21] /*20381*/;
  assign sum_14[21] = _6467_ ^ _6466_ /*20380*/;
  assign _6468_ = _6467_ & _6466_ /*20379*/;
  assign _6469_ = inv_14[21] & r_13[21] /*20378*/;
  assign _6470_ = _6468_ | _6469_ /*20377*/;
  assign _6471_ = inv_14[22] ^ r_13[22] /*20375*/;
  assign sum_14[22] = _6471_ ^ _6470_ /*20374*/;
  assign _6472_ = _6471_ & _6470_ /*20373*/;
  assign _6473_ = inv_14[22] & r_13[22] /*20372*/;
  assign _6474_ = _6472_ | _6473_ /*20371*/;
  assign _6475_ = inv_14[23] ^ r_13[23] /*20369*/;
  assign sum_14[23] = _6475_ ^ _6474_ /*20368*/;
  assign _6476_ = _6475_ & _6474_ /*20367*/;
  assign _6477_ = inv_14[23] & r_13[23] /*20366*/;
  assign _6478_ = _6476_ | _6477_ /*20365*/;
  assign _6479_ = inv_14[24] ^ r_13[24] /*20363*/;
  assign sum_14[24] = _6479_ ^ _6478_ /*20362*/;
  assign _6480_ = _6479_ & _6478_ /*20361*/;
  assign _6481_ = inv_14[24] & r_13[24] /*20360*/;
  assign _6482_ = _6480_ | _6481_ /*20359*/;
  assign _6483_ = inv_14[25] ^ r_13[25] /*20357*/;
  assign sum_14[25] = _6483_ ^ _6482_ /*20356*/;
  assign _6484_ = _6483_ & _6482_ /*20355*/;
  assign _6485_ = inv_14[25] & r_13[25] /*20354*/;
  assign _6486_ = _6484_ | _6485_ /*20353*/;
  assign _6487_ = inv_14[26] ^ r_13[26] /*20351*/;
  assign sum_14[26] = _6487_ ^ _6486_ /*20350*/;
  assign _6488_ = _6487_ & _6486_ /*20349*/;
  assign _6489_ = inv_14[26] & r_13[26] /*20348*/;
  assign _6490_ = _6488_ | _6489_ /*20347*/;
  assign _6491_ = inv_14[27] ^ r_13[27] /*20345*/;
  assign sum_14[27] = _6491_ ^ _6490_ /*20344*/;
  assign _6492_ = _6491_ & _6490_ /*20343*/;
  assign _6493_ = inv_14[27] & r_13[27] /*20342*/;
  assign _6494_ = _6492_ | _6493_ /*20341*/;
  assign _6495_ = inv_14[28] ^ r_13[28] /*20339*/;
  assign sum_14[28] = _6495_ ^ _6494_ /*20338*/;
  assign _6496_ = _6495_ & _6494_ /*20337*/;
  assign _6497_ = inv_14[28] & r_13[28] /*20336*/;
  assign _6498_ = _6496_ | _6497_ /*20335*/;
  assign _6499_ = inv_14[29] ^ r_13[29] /*20333*/;
  assign sum_14[29] = _6499_ ^ _6498_ /*20332*/;
  assign _6500_ = _6499_ & _6498_ /*20331*/;
  assign _6501_ = inv_14[29] & r_13[29] /*20330*/;
  assign _6502_ = _6500_ | _6501_ /*20329*/;
  assign _6503_ = inv_14[30] ^ r_13[30] /*20327*/;
  assign sum_14[30] = _6503_ ^ _6502_ /*20326*/;
  assign _6504_ = _6503_ & _6502_ /*20325*/;
  assign _6505_ = inv_14[30] & r_13[30] /*20324*/;
  assign _6506_ = _6504_ | _6505_ /*20323*/;
  assign _6507_ = inv_14[31] ^ r_13[31] /*20321*/;
  assign sum_14[31] = _6507_ ^ _6506_ /*20320*/;
  assign _6508_ = _6507_ & _6506_ /*20319*/;
  assign _6509_ = inv_14[31] & r_13[31] /*20318*/;
  assign _6510_ = _6508_ | _6509_ /*20317*/;
  assign _6511_ = inv_14[32] ^ r_13[32] /*20315*/;
  assign sum_14[32] = _6511_ ^ _6510_ /*20314*/;
  assign _6512_ = _6511_ & _6510_ /*20313*/;
  assign _6513_ = inv_14[32] & r_13[32] /*20312*/;
  assign _6514_ = _6512_ | _6513_ /*20311*/;
  assign _6515_ = inv_14[33] ^ r_13[33] /*20309*/;
  assign sum_14[33] = _6515_ ^ _6514_ /*20308*/;
  assign _6516_ = _6515_ & _6514_ /*20307*/;
  assign _6517_ = inv_14[33] & r_13[33] /*20306*/;
  assign _6518_ = _6516_ | _6517_ /*20305*/;
  assign _6519_ = inv_14[34] ^ r_13[34] /*20303*/;
  assign sum_14[34] = _6519_ ^ _6518_ /*20302*/;
  assign _6520_ = _6519_ & _6518_ /*20301*/;
  assign _6521_ = inv_14[34] & r_13[34] /*20300*/;
  assign _6522_ = _6520_ | _6521_ /*20299*/;
  assign _6523_ = inv_14[35] ^ r_13[35] /*20297*/;
  assign sum_14[35] = _6523_ ^ _6522_ /*20296*/;
  assign _6524_ = _6523_ & _6522_ /*20295*/;
  assign _6525_ = inv_14[35] & r_13[35] /*20294*/;
  assign _6526_ = _6524_ | _6525_ /*20293*/;
  assign _6527_ = inv_14[36] ^ r_13[36] /*20291*/;
  assign sum_14[36] = _6527_ ^ _6526_ /*20290*/;
  assign _6528_ = _6527_ & _6526_ /*20289*/;
  assign _6529_ = inv_14[36] & r_13[36] /*20288*/;
  assign _6530_ = _6528_ | _6529_ /*20287*/;
  assign _6531_ = inv_14[37] ^ r_13[37] /*20285*/;
  assign sum_14[37] = _6531_ ^ _6530_ /*20284*/;
  assign _6532_ = _6531_ & _6530_ /*20283*/;
  assign _6533_ = inv_14[37] & r_13[37] /*20282*/;
  assign _6534_ = _6532_ | _6533_ /*20281*/;
  assign _6535_ = inv_14[38] ^ r_13[38] /*20279*/;
  assign sum_14[38] = _6535_ ^ _6534_ /*20278*/;
  assign _6536_ = _6535_ & _6534_ /*20277*/;
  assign _6537_ = inv_14[38] & r_13[38] /*20276*/;
  assign _6538_ = _6536_ | _6537_ /*20275*/;
  assign _6539_ = inv_14[39] ^ r_13[39] /*20273*/;
  assign sum_14[39] = _6539_ ^ _6538_ /*20272*/;
  assign _6540_ = _6539_ & _6538_ /*20271*/;
  assign _6541_ = inv_14[39] & r_13[39] /*20270*/;
  assign _6542_ = _6540_ | _6541_ /*20269*/;
  assign _6543_ = inv_14[40] ^ r_13[40] /*20267*/;
  assign sum_14[40] = _6543_ ^ _6542_ /*20266*/;
  assign _6544_ = _6543_ & _6542_ /*20265*/;
  assign _6545_ = inv_14[40] & r_13[40] /*20264*/;
  assign _6546_ = _6544_ | _6545_ /*20263*/;
  assign _6547_ = inv_14[41] ^ r_13[41] /*20261*/;
  assign sum_14[41] = _6547_ ^ _6546_ /*20260*/;
  assign _6548_ = _6547_ & _6546_ /*20259*/;
  assign _6549_ = inv_14[41] & r_13[41] /*20258*/;
  assign _6550_ = _6548_ | _6549_ /*20257*/;
  assign _6551_ = inv_14[42] ^ r_13[42] /*20255*/;
  assign sum_14[42] = _6551_ ^ _6550_ /*20254*/;
  assign _6552_ = _6551_ & _6550_ /*20253*/;
  assign _6553_ = inv_14[42] & r_13[42] /*20252*/;
  assign _6554_ = _6552_ | _6553_ /*20251*/;
  assign _6555_ = inv_14[43] ^ r_13[43] /*20249*/;
  assign sum_14[43] = _6555_ ^ _6554_ /*20248*/;
  assign _6556_ = _6555_ & _6554_ /*20247*/;
  assign _6557_ = inv_14[43] & r_13[43] /*20246*/;
  assign _6558_ = _6556_ | _6557_ /*20245*/;
  assign _6559_ = inv_14[44] ^ r_13[44] /*20243*/;
  assign sum_14[44] = _6559_ ^ _6558_ /*20242*/;
  assign _6560_ = _6559_ & _6558_ /*20241*/;
  assign _6561_ = inv_14[44] & r_13[44] /*20240*/;
  assign _6562_ = _6560_ | _6561_ /*20239*/;
  assign _6563_ = inv_14[45] ^ r_13[45] /*20237*/;
  assign sum_14[45] = _6563_ ^ _6562_ /*20236*/;
  assign _6564_ = _6563_ & _6562_ /*20235*/;
  assign _6565_ = inv_14[45] & r_13[45] /*20234*/;
  assign _6566_ = _6564_ | _6565_ /*20233*/;
  assign _6567_ = inv_14[46] ^ r_13[46] /*20231*/;
  assign sum_14[46] = _6567_ ^ _6566_ /*20230*/;
  assign _6568_ = _6567_ & _6566_ /*20229*/;
  assign _6569_ = inv_14[46] & r_13[46] /*20228*/;
  assign _6570_ = _6568_ | _6569_ /*20227*/;
  assign _6571_ = inv_14[47] ^ r_13[47] /*20225*/;
  assign sum_14[47] = _6571_ ^ _6570_ /*20224*/;
  assign _6572_ = _6571_ & _6570_ /*20223*/;
  assign _6573_ = inv_14[47] & r_13[47] /*20222*/;
  assign _6574_ = _6572_ | _6573_ /*20221*/;
  assign _6575_ = inv_14[48] ^ r_13[48] /*20219*/;
  assign sum_14[48] = _6575_ ^ _6574_ /*20218*/;
  assign _6576_ = _6575_ & _6574_ /*20217*/;
  assign _6577_ = inv_14[48] & r_13[48] /*20216*/;
  assign _6578_ = _6576_ | _6577_ /*20215*/;
  assign _6579_ = inv_14[49] ^ r_13[49] /*20213*/;
  assign sum_14[49] = _6579_ ^ _6578_ /*20212*/;
  assign _6580_ = _6579_ & _6578_ /*20211*/;
  assign _6581_ = inv_14[49] & r_13[49] /*20210*/;
  assign _6582_ = _6580_ | _6581_ /*20209*/;
  assign _6583_ = inv_14[50] ^ r_13[50] /*20207*/;
  assign sum_14[50] = _6583_ ^ _6582_ /*20206*/;
  assign _6584_ = _6583_ & _6582_ /*20205*/;
  assign _6585_ = inv_14[50] & r_13[50] /*20204*/;
  assign _6586_ = _6584_ | _6585_ /*20203*/;
  assign _6587_ = inv_14[51] ^ r_13[51] /*20201*/;
  assign sum_14[51] = _6587_ ^ _6586_ /*20200*/;
  assign _6588_ = _6587_ & _6586_ /*20199*/;
  assign _6589_ = inv_14[51] & r_13[51] /*20198*/;
  assign _6590_ = _6588_ | _6589_ /*20197*/;
  assign _6591_ = inv_14[52] ^ r_13[52] /*20195*/;
  assign sum_14[52] = _6591_ ^ _6590_ /*20194*/;
  assign _6592_ = _6591_ & _6590_ /*20193*/;
  assign _6593_ = inv_14[52] & r_13[52] /*20192*/;
  assign _6594_ = _6592_ | _6593_ /*20191*/;
  assign _6595_ = inv_14[53] ^ r_13[53] /*20189*/;
  assign sum_14[53] = _6595_ ^ _6594_ /*20188*/;
  assign _6596_ = _6595_ & _6594_ /*20187*/;
  assign _6597_ = inv_14[53] & r_13[53] /*20186*/;
  assign _6598_ = _6596_ | _6597_ /*20185*/;
  assign _6599_ = inv_14[54] ^ r_13[54] /*20183*/;
  assign sum_14[54] = _6599_ ^ _6598_ /*20182*/;
  assign _6600_ = _6599_ & _6598_ /*20181*/;
  assign _6601_ = inv_14[54] & r_13[54] /*20180*/;
  assign _6602_ = _6600_ | _6601_ /*20179*/;
  assign _6603_ = inv_14[55] ^ r_13[55] /*20177*/;
  assign sum_14[55] = _6603_ ^ _6602_ /*20176*/;
  assign _6604_ = _6603_ & _6602_ /*20175*/;
  assign _6605_ = inv_14[55] & r_13[55] /*20174*/;
  assign _6606_ = _6604_ | _6605_ /*20173*/;
  assign _6607_ = inv_14[56] ^ r_13[56] /*20171*/;
  assign sum_14[56] = _6607_ ^ _6606_ /*20170*/;
  assign _6608_ = _6607_ & _6606_ /*20169*/;
  assign _6609_ = inv_14[56] & r_13[56] /*20168*/;
  assign _6610_ = _6608_ | _6609_ /*20167*/;
  assign _6611_ = inv_14[57] ^ r_13[57] /*20165*/;
  assign sum_14[57] = _6611_ ^ _6610_ /*20164*/;
  assign _6612_ = _6611_ & _6610_ /*20163*/;
  assign _6613_ = inv_14[57] & r_13[57] /*20162*/;
  assign _6614_ = _6612_ | _6613_ /*20161*/;
  assign _6615_ = inv_14[58] ^ r_13[58] /*20159*/;
  assign sum_14[58] = _6615_ ^ _6614_ /*20158*/;
  assign _6616_ = _6615_ & _6614_ /*20157*/;
  assign _6617_ = inv_14[58] & r_13[58] /*20156*/;
  assign _6618_ = _6616_ | _6617_ /*20155*/;
  assign _6619_ = inv_14[59] ^ r_13[59] /*20153*/;
  assign sum_14[59] = _6619_ ^ _6618_ /*20152*/;
  assign _6620_ = _6619_ & _6618_ /*20151*/;
  assign _6621_ = inv_14[59] & r_13[59] /*20150*/;
  assign _6622_ = _6620_ | _6621_ /*20149*/;
  assign _6623_ = inv_14[60] ^ r_13[60] /*20147*/;
  assign sum_14[60] = _6623_ ^ _6622_ /*20146*/;
  assign _6624_ = _6623_ & _6622_ /*20145*/;
  assign _6625_ = inv_14[60] & r_13[60] /*20144*/;
  assign _6626_ = _6624_ | _6625_ /*20143*/;
  assign _6627_ = inv_14[61] ^ r_13[61] /*20141*/;
  assign sum_14[61] = _6627_ ^ _6626_ /*20140*/;
  assign _6628_ = _6627_ & _6626_ /*20139*/;
  assign _6629_ = inv_14[61] & r_13[61] /*20138*/;
  assign _6630_ = _6628_ | _6629_ /*20137*/;
  assign _6631_ = inv_14[62] ^ r_13[62] /*20135*/;
  assign sum_14[62] = _6631_ ^ _6630_ /*20134*/;
  assign _6632_ = _6631_ & _6630_ /*20133*/;
  assign _6633_ = inv_14[62] & r_13[62] /*20132*/;
  assign _6634_ = _6632_ | _6633_ /*20131*/;
  assign _6635_ = inv_14[63] ^ r_13[63] /*20129*/;
  assign sum_14[63] = _6635_ ^ _6634_ /*20128*/;
  assign _6636_ = _6635_ & _6634_ /*20127*/;
  assign _6637_ = inv_14[63] & r_13[63] /*20126*/;
  assign _6638_ = _6636_ | _6637_ /*20125*/;
  assign _6639_ = inv_14[64] ^ r_13[64] /*20123*/;
  assign sum_14[64] = _6639_ ^ _6638_ /*20122*/;
  assign _6640_ = _6639_ & _6638_ /*20121*/;
  assign _6641_ = inv_14[64] & r_13[64] /*20120*/;
  assign _6642_ = _6640_ | _6641_ /*20119*/;
  assign _6643_ = inv_14[65] ^ r_13[65] /*20117*/;
  assign sum_14[65] = _6643_ ^ _6642_ /*20116*/;
  assign _6644_ = _6643_ & _6642_ /*20115*/;
  assign _6645_ = inv_14[65] & r_13[65] /*20114*/;
  assign _6646_ = _6644_ | _6645_ /*20113*/;
  assign _6647_ = inv_14[66] ^ r_13[66] /*20111*/;
  assign sum_14[66] = _6647_ ^ _6646_ /*20110*/;
  assign _6648_ = _6647_ & _6646_ /*20109*/;
  assign _6649_ = inv_14[66] & r_13[66] /*20108*/;
  assign _6650_ = _6648_ | _6649_ /*20107*/;
  assign _6651_ = inv_14[67] ^ r_13[67] /*20105*/;
  assign sum_14[67] = _6651_ ^ _6650_ /*20104*/;
  assign _6652_ = _6651_ & _6650_ /*20103*/;
  assign _6653_ = inv_14[67] & r_13[67] /*20102*/;
  assign _6654_ = _6652_ | _6653_ /*20101*/;
  assign _6655_ = inv_14[68] ^ r_13[68] /*20099*/;
  assign sum_14[68] = _6655_ ^ _6654_ /*20098*/;
  assign _6656_ = _6655_ & _6654_ /*20097*/;
  assign _6657_ = inv_14[68] & r_13[68] /*20096*/;
  assign _6658_ = _6656_ | _6657_ /*20095*/;
  assign _6659_ = inv_14[69] ^ r_13[69] /*20093*/;
  assign sum_14[69] = _6659_ ^ _6658_ /*20092*/;
  assign _6660_ = _6659_ & _6658_ /*20091*/;
  assign _6661_ = inv_14[69] & r_13[69] /*20090*/;
  assign _6662_ = _6660_ | _6661_ /*20089*/;
  assign _6663_ = inv_14[70] ^ r_13[70] /*20087*/;
  assign sum_14[70] = _6663_ ^ _6662_ /*20086*/;
  assign _6664_ = _6663_ & _6662_ /*20085*/;
  assign _6665_ = inv_14[70] & r_13[70] /*20084*/;
  assign _6666_ = _6664_ | _6665_ /*20083*/;
  assign _6667_ = inv_14[71] ^ r_13[71] /*20081*/;
  assign sum_14[71] = _6667_ ^ _6666_ /*20080*/;
  assign _6668_ = _6667_ & _6666_ /*20079*/;
  assign _6669_ = inv_14[71] & r_13[71] /*20078*/;
  assign _6670_ = _6668_ | _6669_ /*20077*/;
  assign _6671_ = inv_14[72] ^ r_13[72] /*20075*/;
  assign sum_14[72] = _6671_ ^ _6670_ /*20074*/;
  assign _6672_ = _6671_ & _6670_ /*20073*/;
  assign _6673_ = inv_14[72] & r_13[72] /*20072*/;
  assign _6674_ = _6672_ | _6673_ /*20071*/;
  assign _6675_ = inv_14[73] ^ r_13[73] /*20069*/;
  assign sum_14[73] = _6675_ ^ _6674_ /*20068*/;
  assign _6676_ = _6675_ & _6674_ /*20067*/;
  assign _6677_ = inv_14[73] & r_13[73] /*20066*/;
  assign _6678_ = _6676_ | _6677_ /*20065*/;
  assign _6679_ = inv_14[74] ^ r_13[74] /*20063*/;
  assign sum_14[74] = _6679_ ^ _6678_ /*20062*/;
  assign _6680_ = _6679_ & _6678_ /*20061*/;
  assign _6681_ = inv_14[74] & r_13[74] /*20060*/;
  assign _6682_ = _6680_ | _6681_ /*20059*/;
  assign _6683_ = inv_14[75] ^ r_13[75] /*20057*/;
  assign sum_14[75] = _6683_ ^ _6682_ /*20056*/;
  assign _6684_ = _6683_ & _6682_ /*20055*/;
  assign _6685_ = inv_14[75] & r_13[75] /*20054*/;
  assign _6686_ = _6684_ | _6685_ /*20053*/;
  assign _6687_ = _6686_ ^ _6682_ /*20052*/;
  assign _6688_ = ~_6687_ /*20051*/;
  assign _6689_ = sum_14[75] & _6688_ /*20050*/;
  assign _6690_ = _6687_ & _6686_ /*20049*/;
  assign sum_14[76] = _6690_ | _6689_ /*20048*/;
  assign q[18] = ~sum_14[76] /*20047*/;
  assign m_14[0] = r_13[0] /*20046*/;
  assign m_14[1] = r_13[1] /*20045*/;
  assign m_14[2] = r_13[2] /*20044*/;
  assign m_14[3] = r_13[3] /*20043*/;
  assign m_14[4] = r_13[4] /*20042*/;
  assign m_14[5] = r_13[5] /*20041*/;
  assign m_14[6] = r_13[6] /*20040*/;
  assign m_14[7] = r_13[7] /*20039*/;
  assign m_14[8] = r_13[8] /*20038*/;
  assign m_14[9] = r_13[9] /*20037*/;
  assign m_14[10] = r_13[10] /*20036*/;
  assign m_14[11] = r_13[11] /*20035*/;
  assign m_14[12] = r_13[12] /*20034*/;
  assign m_14[13] = r_13[13] /*20033*/;
  assign m_14[14] = r_13[14] /*20032*/;
  assign m_14[15] = r_13[15] /*20031*/;
  assign m_14[16] = r_13[16] /*20030*/;
  assign m_14[17] = r_13[17] /*20029*/;
  assign m_14[18] = r_13[18] /*20028*/;
  assign m_14[19] = r_13[19] /*20027*/;
  assign m_14[20] = r_13[20] /*20026*/;
  assign m_14[21] = r_13[21] /*20025*/;
  assign m_14[22] = r_13[22] /*20024*/;
  assign m_14[23] = r_13[23] /*20023*/;
  assign m_14[24] = r_13[24] /*20022*/;
  assign m_14[25] = r_13[25] /*20021*/;
  assign m_14[26] = r_13[26] /*20020*/;
  assign m_14[27] = r_13[27] /*20019*/;
  assign m_14[28] = r_13[28] /*20018*/;
  assign m_14[29] = r_13[29] /*20017*/;
  assign m_14[30] = r_13[30] /*20016*/;
  assign m_14[31] = r_13[31] /*20015*/;
  assign m_14[32] = r_13[32] /*20014*/;
  assign m_14[33] = r_13[33] /*20013*/;
  assign m_14[34] = r_13[34] /*20012*/;
  assign m_14[35] = r_13[35] /*20011*/;
  assign m_14[36] = r_13[36] /*20010*/;
  assign m_14[37] = r_13[37] /*20009*/;
  assign m_14[38] = r_13[38] /*20008*/;
  assign m_14[39] = r_13[39] /*20007*/;
  assign m_14[40] = r_13[40] /*20006*/;
  assign m_14[41] = r_13[41] /*20005*/;
  assign m_14[42] = r_13[42] /*20004*/;
  assign m_14[43] = r_13[43] /*20003*/;
  assign m_14[44] = r_13[44] /*20002*/;
  assign m_14[45] = r_13[45] /*20001*/;
  assign m_14[46] = r_13[46] /*20000*/;
  assign m_14[47] = r_13[47] /*19999*/;
  assign m_14[48] = r_13[48] /*19998*/;
  assign m_14[49] = r_13[49] /*19997*/;
  assign m_14[50] = r_13[50] /*19996*/;
  assign m_14[51] = r_13[51] /*19995*/;
  assign m_14[52] = r_13[52] /*19994*/;
  assign m_14[53] = r_13[53] /*19993*/;
  assign m_14[54] = r_13[54] /*19992*/;
  assign m_14[55] = r_13[55] /*19991*/;
  assign m_14[56] = r_13[56] /*19990*/;
  assign m_14[57] = r_13[57] /*19989*/;
  assign m_14[58] = r_13[58] /*19988*/;
  assign m_14[59] = r_13[59] /*19987*/;
  assign m_14[60] = r_13[60] /*19986*/;
  assign m_14[61] = r_13[61] /*19985*/;
  assign m_14[62] = r_13[62] /*19984*/;
  assign m_14[63] = r_13[63] /*19983*/;
  assign m_14[64] = r_13[64] /*19982*/;
  assign m_14[65] = r_13[65] /*19981*/;
  assign m_14[66] = r_13[66] /*19980*/;
  assign m_14[67] = r_13[67] /*19979*/;
  assign m_14[68] = r_13[68] /*19978*/;
  assign m_14[69] = r_13[69] /*19977*/;
  assign m_14[70] = r_13[70] /*19976*/;
  assign m_14[71] = r_13[71] /*19975*/;
  assign m_14[72] = r_13[72] /*19974*/;
  assign m_14[73] = r_13[73] /*19973*/;
  assign m_14[74] = r_13[74] /*19972*/;
  assign m_14[75] = r_13[75] /*19971*/;
  assign m_14[76] = r_13[75] /*19970*/;
  assign _6692_ = ~q[18] /*19969*/;
  assign _6693_ = sum_14[0] & q[18] /*19968*/;
  assign _6694_ = m_14[0] & _6692_ /*19967*/;
  assign r_14[0] = _6694_ | _6693_ /*19966*/;
  assign _6695_ = ~q[18] /*19965*/;
  assign _6696_ = sum_14[1] & q[18] /*19964*/;
  assign _6697_ = m_14[1] & _6695_ /*19963*/;
  assign r_14[1] = _6697_ | _6696_ /*19962*/;
  assign _6698_ = ~q[18] /*19961*/;
  assign _6699_ = sum_14[2] & q[18] /*19960*/;
  assign _6700_ = m_14[2] & _6698_ /*19959*/;
  assign r_14[2] = _6700_ | _6699_ /*19958*/;
  assign _6701_ = ~q[18] /*19957*/;
  assign _6702_ = sum_14[3] & q[18] /*19956*/;
  assign _6703_ = m_14[3] & _6701_ /*19955*/;
  assign r_14[3] = _6703_ | _6702_ /*19954*/;
  assign _6704_ = ~q[18] /*19953*/;
  assign _6705_ = sum_14[4] & q[18] /*19952*/;
  assign _6706_ = m_14[4] & _6704_ /*19951*/;
  assign r_14[4] = _6706_ | _6705_ /*19950*/;
  assign _6707_ = ~q[18] /*19949*/;
  assign _6708_ = sum_14[5] & q[18] /*19948*/;
  assign _6709_ = m_14[5] & _6707_ /*19947*/;
  assign r_14[5] = _6709_ | _6708_ /*19946*/;
  assign _6710_ = ~q[18] /*19945*/;
  assign _6711_ = sum_14[6] & q[18] /*19944*/;
  assign _6712_ = m_14[6] & _6710_ /*19943*/;
  assign r_14[6] = _6712_ | _6711_ /*19942*/;
  assign _6713_ = ~q[18] /*19941*/;
  assign _6714_ = sum_14[7] & q[18] /*19940*/;
  assign _6715_ = m_14[7] & _6713_ /*19939*/;
  assign r_14[7] = _6715_ | _6714_ /*19938*/;
  assign _6716_ = ~q[18] /*19937*/;
  assign _6717_ = sum_14[8] & q[18] /*19936*/;
  assign _6718_ = m_14[8] & _6716_ /*19935*/;
  assign r_14[8] = _6718_ | _6717_ /*19934*/;
  assign _6719_ = ~q[18] /*19933*/;
  assign _6720_ = sum_14[9] & q[18] /*19932*/;
  assign _6721_ = m_14[9] & _6719_ /*19931*/;
  assign r_14[9] = _6721_ | _6720_ /*19930*/;
  assign _6722_ = ~q[18] /*19929*/;
  assign _6723_ = sum_14[10] & q[18] /*19928*/;
  assign _6724_ = m_14[10] & _6722_ /*19927*/;
  assign r_14[10] = _6724_ | _6723_ /*19926*/;
  assign _6725_ = ~q[18] /*19925*/;
  assign _6726_ = sum_14[11] & q[18] /*19924*/;
  assign _6727_ = m_14[11] & _6725_ /*19923*/;
  assign r_14[11] = _6727_ | _6726_ /*19922*/;
  assign _6728_ = ~q[18] /*19921*/;
  assign _6729_ = sum_14[12] & q[18] /*19920*/;
  assign _6730_ = m_14[12] & _6728_ /*19919*/;
  assign r_14[12] = _6730_ | _6729_ /*19918*/;
  assign _6731_ = ~q[18] /*19917*/;
  assign _6732_ = sum_14[13] & q[18] /*19916*/;
  assign _6733_ = m_14[13] & _6731_ /*19915*/;
  assign r_14[13] = _6733_ | _6732_ /*19914*/;
  assign _6734_ = ~q[18] /*19913*/;
  assign _6735_ = sum_14[14] & q[18] /*19912*/;
  assign _6736_ = m_14[14] & _6734_ /*19911*/;
  assign r_14[14] = _6736_ | _6735_ /*19910*/;
  assign _6737_ = ~q[18] /*19909*/;
  assign _6738_ = sum_14[15] & q[18] /*19908*/;
  assign _6739_ = m_14[15] & _6737_ /*19907*/;
  assign r_14[15] = _6739_ | _6738_ /*19906*/;
  assign _6740_ = ~q[18] /*19905*/;
  assign _6741_ = sum_14[16] & q[18] /*19904*/;
  assign _6742_ = m_14[16] & _6740_ /*19903*/;
  assign r_14[16] = _6742_ | _6741_ /*19902*/;
  assign _6743_ = ~q[18] /*19901*/;
  assign _6744_ = sum_14[17] & q[18] /*19900*/;
  assign _6745_ = m_14[17] & _6743_ /*19899*/;
  assign r_14[17] = _6745_ | _6744_ /*19898*/;
  assign _6746_ = ~q[18] /*19897*/;
  assign _6747_ = sum_14[18] & q[18] /*19896*/;
  assign _6748_ = m_14[18] & _6746_ /*19895*/;
  assign r_14[18] = _6748_ | _6747_ /*19894*/;
  assign _6749_ = ~q[18] /*19893*/;
  assign _6750_ = sum_14[19] & q[18] /*19892*/;
  assign _6751_ = m_14[19] & _6749_ /*19891*/;
  assign r_14[19] = _6751_ | _6750_ /*19890*/;
  assign _6752_ = ~q[18] /*19889*/;
  assign _6753_ = sum_14[20] & q[18] /*19888*/;
  assign _6754_ = m_14[20] & _6752_ /*19887*/;
  assign r_14[20] = _6754_ | _6753_ /*19886*/;
  assign _6755_ = ~q[18] /*19885*/;
  assign _6756_ = sum_14[21] & q[18] /*19884*/;
  assign _6757_ = m_14[21] & _6755_ /*19883*/;
  assign r_14[21] = _6757_ | _6756_ /*19882*/;
  assign _6758_ = ~q[18] /*19881*/;
  assign _6759_ = sum_14[22] & q[18] /*19880*/;
  assign _6760_ = m_14[22] & _6758_ /*19879*/;
  assign r_14[22] = _6760_ | _6759_ /*19878*/;
  assign _6761_ = ~q[18] /*19877*/;
  assign _6762_ = sum_14[23] & q[18] /*19876*/;
  assign _6763_ = m_14[23] & _6761_ /*19875*/;
  assign r_14[23] = _6763_ | _6762_ /*19874*/;
  assign _6764_ = ~q[18] /*19873*/;
  assign _6765_ = sum_14[24] & q[18] /*19872*/;
  assign _6766_ = m_14[24] & _6764_ /*19871*/;
  assign r_14[24] = _6766_ | _6765_ /*19870*/;
  assign _6767_ = ~q[18] /*19869*/;
  assign _6768_ = sum_14[25] & q[18] /*19868*/;
  assign _6769_ = m_14[25] & _6767_ /*19867*/;
  assign r_14[25] = _6769_ | _6768_ /*19866*/;
  assign _6770_ = ~q[18] /*19865*/;
  assign _6771_ = sum_14[26] & q[18] /*19864*/;
  assign _6772_ = m_14[26] & _6770_ /*19863*/;
  assign r_14[26] = _6772_ | _6771_ /*19862*/;
  assign _6773_ = ~q[18] /*19861*/;
  assign _6774_ = sum_14[27] & q[18] /*19860*/;
  assign _6775_ = m_14[27] & _6773_ /*19859*/;
  assign r_14[27] = _6775_ | _6774_ /*19858*/;
  assign _6776_ = ~q[18] /*19857*/;
  assign _6777_ = sum_14[28] & q[18] /*19856*/;
  assign _6778_ = m_14[28] & _6776_ /*19855*/;
  assign r_14[28] = _6778_ | _6777_ /*19854*/;
  assign _6779_ = ~q[18] /*19853*/;
  assign _6780_ = sum_14[29] & q[18] /*19852*/;
  assign _6781_ = m_14[29] & _6779_ /*19851*/;
  assign r_14[29] = _6781_ | _6780_ /*19850*/;
  assign _6782_ = ~q[18] /*19849*/;
  assign _6783_ = sum_14[30] & q[18] /*19848*/;
  assign _6784_ = m_14[30] & _6782_ /*19847*/;
  assign r_14[30] = _6784_ | _6783_ /*19846*/;
  assign _6785_ = ~q[18] /*19845*/;
  assign _6786_ = sum_14[31] & q[18] /*19844*/;
  assign _6787_ = m_14[31] & _6785_ /*19843*/;
  assign r_14[31] = _6787_ | _6786_ /*19842*/;
  assign _6788_ = ~q[18] /*19841*/;
  assign _6789_ = sum_14[32] & q[18] /*19840*/;
  assign _6790_ = m_14[32] & _6788_ /*19839*/;
  assign r_14[32] = _6790_ | _6789_ /*19838*/;
  assign _6791_ = ~q[18] /*19837*/;
  assign _6792_ = sum_14[33] & q[18] /*19836*/;
  assign _6793_ = m_14[33] & _6791_ /*19835*/;
  assign r_14[33] = _6793_ | _6792_ /*19834*/;
  assign _6794_ = ~q[18] /*19833*/;
  assign _6795_ = sum_14[34] & q[18] /*19832*/;
  assign _6796_ = m_14[34] & _6794_ /*19831*/;
  assign r_14[34] = _6796_ | _6795_ /*19830*/;
  assign _6797_ = ~q[18] /*19829*/;
  assign _6798_ = sum_14[35] & q[18] /*19828*/;
  assign _6799_ = m_14[35] & _6797_ /*19827*/;
  assign r_14[35] = _6799_ | _6798_ /*19826*/;
  assign _6800_ = ~q[18] /*19825*/;
  assign _6801_ = sum_14[36] & q[18] /*19824*/;
  assign _6802_ = m_14[36] & _6800_ /*19823*/;
  assign r_14[36] = _6802_ | _6801_ /*19822*/;
  assign _6803_ = ~q[18] /*19821*/;
  assign _6804_ = sum_14[37] & q[18] /*19820*/;
  assign _6805_ = m_14[37] & _6803_ /*19819*/;
  assign r_14[37] = _6805_ | _6804_ /*19818*/;
  assign _6806_ = ~q[18] /*19817*/;
  assign _6807_ = sum_14[38] & q[18] /*19816*/;
  assign _6808_ = m_14[38] & _6806_ /*19815*/;
  assign r_14[38] = _6808_ | _6807_ /*19814*/;
  assign _6809_ = ~q[18] /*19813*/;
  assign _6810_ = sum_14[39] & q[18] /*19812*/;
  assign _6811_ = m_14[39] & _6809_ /*19811*/;
  assign r_14[39] = _6811_ | _6810_ /*19810*/;
  assign _6812_ = ~q[18] /*19809*/;
  assign _6813_ = sum_14[40] & q[18] /*19808*/;
  assign _6814_ = m_14[40] & _6812_ /*19807*/;
  assign r_14[40] = _6814_ | _6813_ /*19806*/;
  assign _6815_ = ~q[18] /*19805*/;
  assign _6816_ = sum_14[41] & q[18] /*19804*/;
  assign _6817_ = m_14[41] & _6815_ /*19803*/;
  assign r_14[41] = _6817_ | _6816_ /*19802*/;
  assign _6818_ = ~q[18] /*19801*/;
  assign _6819_ = sum_14[42] & q[18] /*19800*/;
  assign _6820_ = m_14[42] & _6818_ /*19799*/;
  assign r_14[42] = _6820_ | _6819_ /*19798*/;
  assign _6821_ = ~q[18] /*19797*/;
  assign _6822_ = sum_14[43] & q[18] /*19796*/;
  assign _6823_ = m_14[43] & _6821_ /*19795*/;
  assign r_14[43] = _6823_ | _6822_ /*19794*/;
  assign _6824_ = ~q[18] /*19793*/;
  assign _6825_ = sum_14[44] & q[18] /*19792*/;
  assign _6826_ = m_14[44] & _6824_ /*19791*/;
  assign r_14[44] = _6826_ | _6825_ /*19790*/;
  assign _6827_ = ~q[18] /*19789*/;
  assign _6828_ = sum_14[45] & q[18] /*19788*/;
  assign _6829_ = m_14[45] & _6827_ /*19787*/;
  assign r_14[45] = _6829_ | _6828_ /*19786*/;
  assign _6830_ = ~q[18] /*19785*/;
  assign _6831_ = sum_14[46] & q[18] /*19784*/;
  assign _6832_ = m_14[46] & _6830_ /*19783*/;
  assign r_14[46] = _6832_ | _6831_ /*19782*/;
  assign _6833_ = ~q[18] /*19781*/;
  assign _6834_ = sum_14[47] & q[18] /*19780*/;
  assign _6835_ = m_14[47] & _6833_ /*19779*/;
  assign r_14[47] = _6835_ | _6834_ /*19778*/;
  assign _6836_ = ~q[18] /*19777*/;
  assign _6837_ = sum_14[48] & q[18] /*19776*/;
  assign _6838_ = m_14[48] & _6836_ /*19775*/;
  assign r_14[48] = _6838_ | _6837_ /*19774*/;
  assign _6839_ = ~q[18] /*19773*/;
  assign _6840_ = sum_14[49] & q[18] /*19772*/;
  assign _6841_ = m_14[49] & _6839_ /*19771*/;
  assign r_14[49] = _6841_ | _6840_ /*19770*/;
  assign _6842_ = ~q[18] /*19769*/;
  assign _6843_ = sum_14[50] & q[18] /*19768*/;
  assign _6844_ = m_14[50] & _6842_ /*19767*/;
  assign r_14[50] = _6844_ | _6843_ /*19766*/;
  assign _6845_ = ~q[18] /*19765*/;
  assign _6846_ = sum_14[51] & q[18] /*19764*/;
  assign _6847_ = m_14[51] & _6845_ /*19763*/;
  assign r_14[51] = _6847_ | _6846_ /*19762*/;
  assign _6848_ = ~q[18] /*19761*/;
  assign _6849_ = sum_14[52] & q[18] /*19760*/;
  assign _6850_ = m_14[52] & _6848_ /*19759*/;
  assign r_14[52] = _6850_ | _6849_ /*19758*/;
  assign _6851_ = ~q[18] /*19757*/;
  assign _6852_ = sum_14[53] & q[18] /*19756*/;
  assign _6853_ = m_14[53] & _6851_ /*19755*/;
  assign r_14[53] = _6853_ | _6852_ /*19754*/;
  assign _6854_ = ~q[18] /*19753*/;
  assign _6855_ = sum_14[54] & q[18] /*19752*/;
  assign _6856_ = m_14[54] & _6854_ /*19751*/;
  assign r_14[54] = _6856_ | _6855_ /*19750*/;
  assign _6857_ = ~q[18] /*19749*/;
  assign _6858_ = sum_14[55] & q[18] /*19748*/;
  assign _6859_ = m_14[55] & _6857_ /*19747*/;
  assign r_14[55] = _6859_ | _6858_ /*19746*/;
  assign _6860_ = ~q[18] /*19745*/;
  assign _6861_ = sum_14[56] & q[18] /*19744*/;
  assign _6862_ = m_14[56] & _6860_ /*19743*/;
  assign r_14[56] = _6862_ | _6861_ /*19742*/;
  assign _6863_ = ~q[18] /*19741*/;
  assign _6864_ = sum_14[57] & q[18] /*19740*/;
  assign _6865_ = m_14[57] & _6863_ /*19739*/;
  assign r_14[57] = _6865_ | _6864_ /*19738*/;
  assign _6866_ = ~q[18] /*19737*/;
  assign _6867_ = sum_14[58] & q[18] /*19736*/;
  assign _6868_ = m_14[58] & _6866_ /*19735*/;
  assign r_14[58] = _6868_ | _6867_ /*19734*/;
  assign _6869_ = ~q[18] /*19733*/;
  assign _6870_ = sum_14[59] & q[18] /*19732*/;
  assign _6871_ = m_14[59] & _6869_ /*19731*/;
  assign r_14[59] = _6871_ | _6870_ /*19730*/;
  assign _6872_ = ~q[18] /*19729*/;
  assign _6873_ = sum_14[60] & q[18] /*19728*/;
  assign _6874_ = m_14[60] & _6872_ /*19727*/;
  assign r_14[60] = _6874_ | _6873_ /*19726*/;
  assign _6875_ = ~q[18] /*19725*/;
  assign _6876_ = sum_14[61] & q[18] /*19724*/;
  assign _6877_ = m_14[61] & _6875_ /*19723*/;
  assign r_14[61] = _6877_ | _6876_ /*19722*/;
  assign _6878_ = ~q[18] /*19721*/;
  assign _6879_ = sum_14[62] & q[18] /*19720*/;
  assign _6880_ = m_14[62] & _6878_ /*19719*/;
  assign r_14[62] = _6880_ | _6879_ /*19718*/;
  assign _6881_ = ~q[18] /*19717*/;
  assign _6882_ = sum_14[63] & q[18] /*19716*/;
  assign _6883_ = m_14[63] & _6881_ /*19715*/;
  assign r_14[63] = _6883_ | _6882_ /*19714*/;
  assign _6884_ = ~q[18] /*19713*/;
  assign _6885_ = sum_14[64] & q[18] /*19712*/;
  assign _6886_ = m_14[64] & _6884_ /*19711*/;
  assign r_14[64] = _6886_ | _6885_ /*19710*/;
  assign _6887_ = ~q[18] /*19709*/;
  assign _6888_ = sum_14[65] & q[18] /*19708*/;
  assign _6889_ = m_14[65] & _6887_ /*19707*/;
  assign r_14[65] = _6889_ | _6888_ /*19706*/;
  assign _6890_ = ~q[18] /*19705*/;
  assign _6891_ = sum_14[66] & q[18] /*19704*/;
  assign _6892_ = m_14[66] & _6890_ /*19703*/;
  assign r_14[66] = _6892_ | _6891_ /*19702*/;
  assign _6893_ = ~q[18] /*19701*/;
  assign _6894_ = sum_14[67] & q[18] /*19700*/;
  assign _6895_ = m_14[67] & _6893_ /*19699*/;
  assign r_14[67] = _6895_ | _6894_ /*19698*/;
  assign _6896_ = ~q[18] /*19697*/;
  assign _6897_ = sum_14[68] & q[18] /*19696*/;
  assign _6898_ = m_14[68] & _6896_ /*19695*/;
  assign r_14[68] = _6898_ | _6897_ /*19694*/;
  assign _6899_ = ~q[18] /*19693*/;
  assign _6900_ = sum_14[69] & q[18] /*19692*/;
  assign _6901_ = m_14[69] & _6899_ /*19691*/;
  assign r_14[69] = _6901_ | _6900_ /*19690*/;
  assign _6902_ = ~q[18] /*19689*/;
  assign _6903_ = sum_14[70] & q[18] /*19688*/;
  assign _6904_ = m_14[70] & _6902_ /*19687*/;
  assign r_14[70] = _6904_ | _6903_ /*19686*/;
  assign _6905_ = ~q[18] /*19685*/;
  assign _6906_ = sum_14[71] & q[18] /*19684*/;
  assign _6907_ = m_14[71] & _6905_ /*19683*/;
  assign r_14[71] = _6907_ | _6906_ /*19682*/;
  assign _6908_ = ~q[18] /*19681*/;
  assign _6909_ = sum_14[72] & q[18] /*19680*/;
  assign _6910_ = m_14[72] & _6908_ /*19679*/;
  assign r_14[72] = _6910_ | _6909_ /*19678*/;
  assign _6911_ = ~q[18] /*19677*/;
  assign _6912_ = sum_14[73] & q[18] /*19676*/;
  assign _6913_ = m_14[73] & _6911_ /*19675*/;
  assign r_14[73] = _6913_ | _6912_ /*19674*/;
  assign _6914_ = ~q[18] /*19673*/;
  assign _6915_ = sum_14[74] & q[18] /*19672*/;
  assign _6916_ = m_14[74] & _6914_ /*19671*/;
  assign r_14[74] = _6916_ | _6915_ /*19670*/;
  assign _6917_ = ~q[18] /*19669*/;
  assign _6918_ = sum_14[75] & q[18] /*19668*/;
  assign _6919_ = m_14[75] & _6917_ /*19667*/;
  assign r_14[75] = _6919_ | _6918_ /*19666*/;
  assign _6920_ = ~q[18] /*19665*/;
  assign _6921_ = sum_14[76] & q[18] /*19664*/;
  assign _6922_ = m_14[76] & _6920_ /*19663*/;
  assign r_14[76] = _6922_ | _6921_ /*19662*/;
  assign inv_15[0] = oneWire /*19432*/;
  assign inv_15[1] = oneWire /*19426*/;
  assign inv_15[2] = oneWire /*19420*/;
  assign inv_15[3] = oneWire /*19414*/;
  assign inv_15[4] = oneWire /*19408*/;
  assign inv_15[5] = oneWire /*19402*/;
  assign inv_15[6] = oneWire /*19396*/;
  assign inv_15[7] = oneWire /*19390*/;
  assign inv_15[8] = oneWire /*19384*/;
  assign inv_15[9] = oneWire /*19378*/;
  assign inv_15[10] = oneWire /*19372*/;
  assign inv_15[11] = oneWire /*19366*/;
  assign inv_15[12] = oneWire /*19360*/;
  assign inv_15[13] = oneWire /*19354*/;
  assign inv_15[14] = oneWire /*19348*/;
  assign inv_15[15] = oneWire /*19342*/;
  assign inv_15[16] = oneWire /*19336*/;
  assign inv_15[17] = ~div[0] /*19330*/;
  assign inv_15[18] = ~div[1] /*19324*/;
  assign inv_15[19] = ~div[2] /*19318*/;
  assign inv_15[20] = ~div[3] /*19312*/;
  assign inv_15[21] = ~div[4] /*19306*/;
  assign inv_15[22] = ~div[5] /*19300*/;
  assign inv_15[23] = ~div[6] /*19294*/;
  assign inv_15[24] = ~div[7] /*19288*/;
  assign inv_15[25] = ~div[8] /*19282*/;
  assign inv_15[26] = ~div[9] /*19276*/;
  assign inv_15[27] = ~div[10] /*19270*/;
  assign inv_15[28] = ~div[11] /*19264*/;
  assign inv_15[29] = ~div[12] /*19258*/;
  assign inv_15[30] = ~div[13] /*19252*/;
  assign inv_15[31] = ~div[14] /*19246*/;
  assign inv_15[32] = ~div[15] /*19240*/;
  assign inv_15[33] = ~div[16] /*19234*/;
  assign inv_15[34] = ~div[17] /*19228*/;
  assign inv_15[35] = ~div[18] /*19222*/;
  assign inv_15[36] = ~div[19] /*19216*/;
  assign inv_15[37] = ~div[20] /*19210*/;
  assign inv_15[38] = ~div[21] /*19204*/;
  assign inv_15[39] = ~div[22] /*19198*/;
  assign inv_15[40] = ~div[23] /*19192*/;
  assign inv_15[41] = ~div[24] /*19186*/;
  assign inv_15[42] = ~div[25] /*19180*/;
  assign inv_15[43] = ~div[26] /*19174*/;
  assign inv_15[44] = ~div[27] /*19168*/;
  assign inv_15[45] = ~div[28] /*19162*/;
  assign inv_15[46] = ~div[29] /*19156*/;
  assign inv_15[47] = ~div[30] /*19150*/;
  assign inv_15[48] = oneWire /*19144*/;
  assign inv_15[49] = oneWire /*19138*/;
  assign inv_15[50] = oneWire /*19132*/;
  assign inv_15[51] = oneWire /*19126*/;
  assign inv_15[52] = oneWire /*19120*/;
  assign inv_15[53] = oneWire /*19114*/;
  assign inv_15[54] = oneWire /*19108*/;
  assign inv_15[55] = oneWire /*19102*/;
  assign inv_15[56] = oneWire /*19096*/;
  assign inv_15[57] = oneWire /*19090*/;
  assign inv_15[58] = oneWire /*19084*/;
  assign inv_15[59] = oneWire /*19078*/;
  assign inv_15[60] = oneWire /*19072*/;
  assign inv_15[61] = oneWire /*19066*/;
  assign inv_15[62] = oneWire /*19060*/;
  assign inv_15[63] = oneWire /*19054*/;
  assign inv_15[64] = oneWire /*19048*/;
  assign inv_15[65] = oneWire /*19042*/;
  assign inv_15[66] = oneWire /*19036*/;
  assign inv_15[67] = oneWire /*19030*/;
  assign inv_15[68] = oneWire /*19024*/;
  assign inv_15[69] = oneWire /*19018*/;
  assign inv_15[70] = oneWire /*19012*/;
  assign inv_15[71] = oneWire /*19006*/;
  assign inv_15[72] = oneWire /*19000*/;
  assign inv_15[73] = oneWire /*18994*/;
  assign inv_15[74] = oneWire /*18988*/;
  assign inv_15[75] = oneWire /*18982*/;
  assign inv_15[76] = oneWire /*18976*/;
  assign _6923_ = inv_15[0] ^ r_14[0] /*19431*/;
  assign sum_15[0] = _6923_ ^ oneWire /*19430*/;
  assign _6924_ = _6923_ & oneWire /*19429*/;
  assign _6925_ = inv_15[0] & r_14[0] /*19428*/;
  assign _6926_ = _6924_ | _6925_ /*19427*/;
  assign _6927_ = inv_15[1] ^ r_14[1] /*19425*/;
  assign sum_15[1] = _6927_ ^ _6926_ /*19424*/;
  assign _6928_ = _6927_ & _6926_ /*19423*/;
  assign _6929_ = inv_15[1] & r_14[1] /*19422*/;
  assign _6930_ = _6928_ | _6929_ /*19421*/;
  assign _6931_ = inv_15[2] ^ r_14[2] /*19419*/;
  assign sum_15[2] = _6931_ ^ _6930_ /*19418*/;
  assign _6932_ = _6931_ & _6930_ /*19417*/;
  assign _6933_ = inv_15[2] & r_14[2] /*19416*/;
  assign _6934_ = _6932_ | _6933_ /*19415*/;
  assign _6935_ = inv_15[3] ^ r_14[3] /*19413*/;
  assign sum_15[3] = _6935_ ^ _6934_ /*19412*/;
  assign _6936_ = _6935_ & _6934_ /*19411*/;
  assign _6937_ = inv_15[3] & r_14[3] /*19410*/;
  assign _6938_ = _6936_ | _6937_ /*19409*/;
  assign _6939_ = inv_15[4] ^ r_14[4] /*19407*/;
  assign sum_15[4] = _6939_ ^ _6938_ /*19406*/;
  assign _6940_ = _6939_ & _6938_ /*19405*/;
  assign _6941_ = inv_15[4] & r_14[4] /*19404*/;
  assign _6942_ = _6940_ | _6941_ /*19403*/;
  assign _6943_ = inv_15[5] ^ r_14[5] /*19401*/;
  assign sum_15[5] = _6943_ ^ _6942_ /*19400*/;
  assign _6944_ = _6943_ & _6942_ /*19399*/;
  assign _6945_ = inv_15[5] & r_14[5] /*19398*/;
  assign _6946_ = _6944_ | _6945_ /*19397*/;
  assign _6947_ = inv_15[6] ^ r_14[6] /*19395*/;
  assign sum_15[6] = _6947_ ^ _6946_ /*19394*/;
  assign _6948_ = _6947_ & _6946_ /*19393*/;
  assign _6949_ = inv_15[6] & r_14[6] /*19392*/;
  assign _6950_ = _6948_ | _6949_ /*19391*/;
  assign _6951_ = inv_15[7] ^ r_14[7] /*19389*/;
  assign sum_15[7] = _6951_ ^ _6950_ /*19388*/;
  assign _6952_ = _6951_ & _6950_ /*19387*/;
  assign _6953_ = inv_15[7] & r_14[7] /*19386*/;
  assign _6954_ = _6952_ | _6953_ /*19385*/;
  assign _6955_ = inv_15[8] ^ r_14[8] /*19383*/;
  assign sum_15[8] = _6955_ ^ _6954_ /*19382*/;
  assign _6956_ = _6955_ & _6954_ /*19381*/;
  assign _6957_ = inv_15[8] & r_14[8] /*19380*/;
  assign _6958_ = _6956_ | _6957_ /*19379*/;
  assign _6959_ = inv_15[9] ^ r_14[9] /*19377*/;
  assign sum_15[9] = _6959_ ^ _6958_ /*19376*/;
  assign _6960_ = _6959_ & _6958_ /*19375*/;
  assign _6961_ = inv_15[9] & r_14[9] /*19374*/;
  assign _6962_ = _6960_ | _6961_ /*19373*/;
  assign _6963_ = inv_15[10] ^ r_14[10] /*19371*/;
  assign sum_15[10] = _6963_ ^ _6962_ /*19370*/;
  assign _6964_ = _6963_ & _6962_ /*19369*/;
  assign _6965_ = inv_15[10] & r_14[10] /*19368*/;
  assign _6966_ = _6964_ | _6965_ /*19367*/;
  assign _6967_ = inv_15[11] ^ r_14[11] /*19365*/;
  assign sum_15[11] = _6967_ ^ _6966_ /*19364*/;
  assign _6968_ = _6967_ & _6966_ /*19363*/;
  assign _6969_ = inv_15[11] & r_14[11] /*19362*/;
  assign _6970_ = _6968_ | _6969_ /*19361*/;
  assign _6971_ = inv_15[12] ^ r_14[12] /*19359*/;
  assign sum_15[12] = _6971_ ^ _6970_ /*19358*/;
  assign _6972_ = _6971_ & _6970_ /*19357*/;
  assign _6973_ = inv_15[12] & r_14[12] /*19356*/;
  assign _6974_ = _6972_ | _6973_ /*19355*/;
  assign _6975_ = inv_15[13] ^ r_14[13] /*19353*/;
  assign sum_15[13] = _6975_ ^ _6974_ /*19352*/;
  assign _6976_ = _6975_ & _6974_ /*19351*/;
  assign _6977_ = inv_15[13] & r_14[13] /*19350*/;
  assign _6978_ = _6976_ | _6977_ /*19349*/;
  assign _6979_ = inv_15[14] ^ r_14[14] /*19347*/;
  assign sum_15[14] = _6979_ ^ _6978_ /*19346*/;
  assign _6980_ = _6979_ & _6978_ /*19345*/;
  assign _6981_ = inv_15[14] & r_14[14] /*19344*/;
  assign _6982_ = _6980_ | _6981_ /*19343*/;
  assign _6983_ = inv_15[15] ^ r_14[15] /*19341*/;
  assign sum_15[15] = _6983_ ^ _6982_ /*19340*/;
  assign _6984_ = _6983_ & _6982_ /*19339*/;
  assign _6985_ = inv_15[15] & r_14[15] /*19338*/;
  assign _6986_ = _6984_ | _6985_ /*19337*/;
  assign _6987_ = inv_15[16] ^ r_14[16] /*19335*/;
  assign sum_15[16] = _6987_ ^ _6986_ /*19334*/;
  assign _6988_ = _6987_ & _6986_ /*19333*/;
  assign _6989_ = inv_15[16] & r_14[16] /*19332*/;
  assign _6990_ = _6988_ | _6989_ /*19331*/;
  assign _6991_ = inv_15[17] ^ r_14[17] /*19329*/;
  assign sum_15[17] = _6991_ ^ _6990_ /*19328*/;
  assign _6992_ = _6991_ & _6990_ /*19327*/;
  assign _6993_ = inv_15[17] & r_14[17] /*19326*/;
  assign _6994_ = _6992_ | _6993_ /*19325*/;
  assign _6995_ = inv_15[18] ^ r_14[18] /*19323*/;
  assign sum_15[18] = _6995_ ^ _6994_ /*19322*/;
  assign _6996_ = _6995_ & _6994_ /*19321*/;
  assign _6997_ = inv_15[18] & r_14[18] /*19320*/;
  assign _6998_ = _6996_ | _6997_ /*19319*/;
  assign _6999_ = inv_15[19] ^ r_14[19] /*19317*/;
  assign sum_15[19] = _6999_ ^ _6998_ /*19316*/;
  assign _7000_ = _6999_ & _6998_ /*19315*/;
  assign _7001_ = inv_15[19] & r_14[19] /*19314*/;
  assign _7002_ = _7000_ | _7001_ /*19313*/;
  assign _7003_ = inv_15[20] ^ r_14[20] /*19311*/;
  assign sum_15[20] = _7003_ ^ _7002_ /*19310*/;
  assign _7004_ = _7003_ & _7002_ /*19309*/;
  assign _7005_ = inv_15[20] & r_14[20] /*19308*/;
  assign _7006_ = _7004_ | _7005_ /*19307*/;
  assign _7007_ = inv_15[21] ^ r_14[21] /*19305*/;
  assign sum_15[21] = _7007_ ^ _7006_ /*19304*/;
  assign _7008_ = _7007_ & _7006_ /*19303*/;
  assign _7009_ = inv_15[21] & r_14[21] /*19302*/;
  assign _7010_ = _7008_ | _7009_ /*19301*/;
  assign _7011_ = inv_15[22] ^ r_14[22] /*19299*/;
  assign sum_15[22] = _7011_ ^ _7010_ /*19298*/;
  assign _7012_ = _7011_ & _7010_ /*19297*/;
  assign _7013_ = inv_15[22] & r_14[22] /*19296*/;
  assign _7014_ = _7012_ | _7013_ /*19295*/;
  assign _7015_ = inv_15[23] ^ r_14[23] /*19293*/;
  assign sum_15[23] = _7015_ ^ _7014_ /*19292*/;
  assign _7016_ = _7015_ & _7014_ /*19291*/;
  assign _7017_ = inv_15[23] & r_14[23] /*19290*/;
  assign _7018_ = _7016_ | _7017_ /*19289*/;
  assign _7019_ = inv_15[24] ^ r_14[24] /*19287*/;
  assign sum_15[24] = _7019_ ^ _7018_ /*19286*/;
  assign _7020_ = _7019_ & _7018_ /*19285*/;
  assign _7021_ = inv_15[24] & r_14[24] /*19284*/;
  assign _7022_ = _7020_ | _7021_ /*19283*/;
  assign _7023_ = inv_15[25] ^ r_14[25] /*19281*/;
  assign sum_15[25] = _7023_ ^ _7022_ /*19280*/;
  assign _7024_ = _7023_ & _7022_ /*19279*/;
  assign _7025_ = inv_15[25] & r_14[25] /*19278*/;
  assign _7026_ = _7024_ | _7025_ /*19277*/;
  assign _7027_ = inv_15[26] ^ r_14[26] /*19275*/;
  assign sum_15[26] = _7027_ ^ _7026_ /*19274*/;
  assign _7028_ = _7027_ & _7026_ /*19273*/;
  assign _7029_ = inv_15[26] & r_14[26] /*19272*/;
  assign _7030_ = _7028_ | _7029_ /*19271*/;
  assign _7031_ = inv_15[27] ^ r_14[27] /*19269*/;
  assign sum_15[27] = _7031_ ^ _7030_ /*19268*/;
  assign _7032_ = _7031_ & _7030_ /*19267*/;
  assign _7033_ = inv_15[27] & r_14[27] /*19266*/;
  assign _7034_ = _7032_ | _7033_ /*19265*/;
  assign _7035_ = inv_15[28] ^ r_14[28] /*19263*/;
  assign sum_15[28] = _7035_ ^ _7034_ /*19262*/;
  assign _7036_ = _7035_ & _7034_ /*19261*/;
  assign _7037_ = inv_15[28] & r_14[28] /*19260*/;
  assign _7038_ = _7036_ | _7037_ /*19259*/;
  assign _7039_ = inv_15[29] ^ r_14[29] /*19257*/;
  assign sum_15[29] = _7039_ ^ _7038_ /*19256*/;
  assign _7040_ = _7039_ & _7038_ /*19255*/;
  assign _7041_ = inv_15[29] & r_14[29] /*19254*/;
  assign _7042_ = _7040_ | _7041_ /*19253*/;
  assign _7043_ = inv_15[30] ^ r_14[30] /*19251*/;
  assign sum_15[30] = _7043_ ^ _7042_ /*19250*/;
  assign _7044_ = _7043_ & _7042_ /*19249*/;
  assign _7045_ = inv_15[30] & r_14[30] /*19248*/;
  assign _7046_ = _7044_ | _7045_ /*19247*/;
  assign _7047_ = inv_15[31] ^ r_14[31] /*19245*/;
  assign sum_15[31] = _7047_ ^ _7046_ /*19244*/;
  assign _7048_ = _7047_ & _7046_ /*19243*/;
  assign _7049_ = inv_15[31] & r_14[31] /*19242*/;
  assign _7050_ = _7048_ | _7049_ /*19241*/;
  assign _7051_ = inv_15[32] ^ r_14[32] /*19239*/;
  assign sum_15[32] = _7051_ ^ _7050_ /*19238*/;
  assign _7052_ = _7051_ & _7050_ /*19237*/;
  assign _7053_ = inv_15[32] & r_14[32] /*19236*/;
  assign _7054_ = _7052_ | _7053_ /*19235*/;
  assign _7055_ = inv_15[33] ^ r_14[33] /*19233*/;
  assign sum_15[33] = _7055_ ^ _7054_ /*19232*/;
  assign _7056_ = _7055_ & _7054_ /*19231*/;
  assign _7057_ = inv_15[33] & r_14[33] /*19230*/;
  assign _7058_ = _7056_ | _7057_ /*19229*/;
  assign _7059_ = inv_15[34] ^ r_14[34] /*19227*/;
  assign sum_15[34] = _7059_ ^ _7058_ /*19226*/;
  assign _7060_ = _7059_ & _7058_ /*19225*/;
  assign _7061_ = inv_15[34] & r_14[34] /*19224*/;
  assign _7062_ = _7060_ | _7061_ /*19223*/;
  assign _7063_ = inv_15[35] ^ r_14[35] /*19221*/;
  assign sum_15[35] = _7063_ ^ _7062_ /*19220*/;
  assign _7064_ = _7063_ & _7062_ /*19219*/;
  assign _7065_ = inv_15[35] & r_14[35] /*19218*/;
  assign _7066_ = _7064_ | _7065_ /*19217*/;
  assign _7067_ = inv_15[36] ^ r_14[36] /*19215*/;
  assign sum_15[36] = _7067_ ^ _7066_ /*19214*/;
  assign _7068_ = _7067_ & _7066_ /*19213*/;
  assign _7069_ = inv_15[36] & r_14[36] /*19212*/;
  assign _7070_ = _7068_ | _7069_ /*19211*/;
  assign _7071_ = inv_15[37] ^ r_14[37] /*19209*/;
  assign sum_15[37] = _7071_ ^ _7070_ /*19208*/;
  assign _7072_ = _7071_ & _7070_ /*19207*/;
  assign _7073_ = inv_15[37] & r_14[37] /*19206*/;
  assign _7074_ = _7072_ | _7073_ /*19205*/;
  assign _7075_ = inv_15[38] ^ r_14[38] /*19203*/;
  assign sum_15[38] = _7075_ ^ _7074_ /*19202*/;
  assign _7076_ = _7075_ & _7074_ /*19201*/;
  assign _7077_ = inv_15[38] & r_14[38] /*19200*/;
  assign _7078_ = _7076_ | _7077_ /*19199*/;
  assign _7079_ = inv_15[39] ^ r_14[39] /*19197*/;
  assign sum_15[39] = _7079_ ^ _7078_ /*19196*/;
  assign _7080_ = _7079_ & _7078_ /*19195*/;
  assign _7081_ = inv_15[39] & r_14[39] /*19194*/;
  assign _7082_ = _7080_ | _7081_ /*19193*/;
  assign _7083_ = inv_15[40] ^ r_14[40] /*19191*/;
  assign sum_15[40] = _7083_ ^ _7082_ /*19190*/;
  assign _7084_ = _7083_ & _7082_ /*19189*/;
  assign _7085_ = inv_15[40] & r_14[40] /*19188*/;
  assign _7086_ = _7084_ | _7085_ /*19187*/;
  assign _7087_ = inv_15[41] ^ r_14[41] /*19185*/;
  assign sum_15[41] = _7087_ ^ _7086_ /*19184*/;
  assign _7088_ = _7087_ & _7086_ /*19183*/;
  assign _7089_ = inv_15[41] & r_14[41] /*19182*/;
  assign _7090_ = _7088_ | _7089_ /*19181*/;
  assign _7091_ = inv_15[42] ^ r_14[42] /*19179*/;
  assign sum_15[42] = _7091_ ^ _7090_ /*19178*/;
  assign _7092_ = _7091_ & _7090_ /*19177*/;
  assign _7093_ = inv_15[42] & r_14[42] /*19176*/;
  assign _7094_ = _7092_ | _7093_ /*19175*/;
  assign _7095_ = inv_15[43] ^ r_14[43] /*19173*/;
  assign sum_15[43] = _7095_ ^ _7094_ /*19172*/;
  assign _7096_ = _7095_ & _7094_ /*19171*/;
  assign _7097_ = inv_15[43] & r_14[43] /*19170*/;
  assign _7098_ = _7096_ | _7097_ /*19169*/;
  assign _7099_ = inv_15[44] ^ r_14[44] /*19167*/;
  assign sum_15[44] = _7099_ ^ _7098_ /*19166*/;
  assign _7100_ = _7099_ & _7098_ /*19165*/;
  assign _7101_ = inv_15[44] & r_14[44] /*19164*/;
  assign _7102_ = _7100_ | _7101_ /*19163*/;
  assign _7103_ = inv_15[45] ^ r_14[45] /*19161*/;
  assign sum_15[45] = _7103_ ^ _7102_ /*19160*/;
  assign _7104_ = _7103_ & _7102_ /*19159*/;
  assign _7105_ = inv_15[45] & r_14[45] /*19158*/;
  assign _7106_ = _7104_ | _7105_ /*19157*/;
  assign _7107_ = inv_15[46] ^ r_14[46] /*19155*/;
  assign sum_15[46] = _7107_ ^ _7106_ /*19154*/;
  assign _7108_ = _7107_ & _7106_ /*19153*/;
  assign _7109_ = inv_15[46] & r_14[46] /*19152*/;
  assign _7110_ = _7108_ | _7109_ /*19151*/;
  assign _7111_ = inv_15[47] ^ r_14[47] /*19149*/;
  assign sum_15[47] = _7111_ ^ _7110_ /*19148*/;
  assign _7112_ = _7111_ & _7110_ /*19147*/;
  assign _7113_ = inv_15[47] & r_14[47] /*19146*/;
  assign _7114_ = _7112_ | _7113_ /*19145*/;
  assign _7115_ = inv_15[48] ^ r_14[48] /*19143*/;
  assign sum_15[48] = _7115_ ^ _7114_ /*19142*/;
  assign _7116_ = _7115_ & _7114_ /*19141*/;
  assign _7117_ = inv_15[48] & r_14[48] /*19140*/;
  assign _7118_ = _7116_ | _7117_ /*19139*/;
  assign _7119_ = inv_15[49] ^ r_14[49] /*19137*/;
  assign sum_15[49] = _7119_ ^ _7118_ /*19136*/;
  assign _7120_ = _7119_ & _7118_ /*19135*/;
  assign _7121_ = inv_15[49] & r_14[49] /*19134*/;
  assign _7122_ = _7120_ | _7121_ /*19133*/;
  assign _7123_ = inv_15[50] ^ r_14[50] /*19131*/;
  assign sum_15[50] = _7123_ ^ _7122_ /*19130*/;
  assign _7124_ = _7123_ & _7122_ /*19129*/;
  assign _7125_ = inv_15[50] & r_14[50] /*19128*/;
  assign _7126_ = _7124_ | _7125_ /*19127*/;
  assign _7127_ = inv_15[51] ^ r_14[51] /*19125*/;
  assign sum_15[51] = _7127_ ^ _7126_ /*19124*/;
  assign _7128_ = _7127_ & _7126_ /*19123*/;
  assign _7129_ = inv_15[51] & r_14[51] /*19122*/;
  assign _7130_ = _7128_ | _7129_ /*19121*/;
  assign _7131_ = inv_15[52] ^ r_14[52] /*19119*/;
  assign sum_15[52] = _7131_ ^ _7130_ /*19118*/;
  assign _7132_ = _7131_ & _7130_ /*19117*/;
  assign _7133_ = inv_15[52] & r_14[52] /*19116*/;
  assign _7134_ = _7132_ | _7133_ /*19115*/;
  assign _7135_ = inv_15[53] ^ r_14[53] /*19113*/;
  assign sum_15[53] = _7135_ ^ _7134_ /*19112*/;
  assign _7136_ = _7135_ & _7134_ /*19111*/;
  assign _7137_ = inv_15[53] & r_14[53] /*19110*/;
  assign _7138_ = _7136_ | _7137_ /*19109*/;
  assign _7139_ = inv_15[54] ^ r_14[54] /*19107*/;
  assign sum_15[54] = _7139_ ^ _7138_ /*19106*/;
  assign _7140_ = _7139_ & _7138_ /*19105*/;
  assign _7141_ = inv_15[54] & r_14[54] /*19104*/;
  assign _7142_ = _7140_ | _7141_ /*19103*/;
  assign _7143_ = inv_15[55] ^ r_14[55] /*19101*/;
  assign sum_15[55] = _7143_ ^ _7142_ /*19100*/;
  assign _7144_ = _7143_ & _7142_ /*19099*/;
  assign _7145_ = inv_15[55] & r_14[55] /*19098*/;
  assign _7146_ = _7144_ | _7145_ /*19097*/;
  assign _7147_ = inv_15[56] ^ r_14[56] /*19095*/;
  assign sum_15[56] = _7147_ ^ _7146_ /*19094*/;
  assign _7148_ = _7147_ & _7146_ /*19093*/;
  assign _7149_ = inv_15[56] & r_14[56] /*19092*/;
  assign _7150_ = _7148_ | _7149_ /*19091*/;
  assign _7151_ = inv_15[57] ^ r_14[57] /*19089*/;
  assign sum_15[57] = _7151_ ^ _7150_ /*19088*/;
  assign _7152_ = _7151_ & _7150_ /*19087*/;
  assign _7153_ = inv_15[57] & r_14[57] /*19086*/;
  assign _7154_ = _7152_ | _7153_ /*19085*/;
  assign _7155_ = inv_15[58] ^ r_14[58] /*19083*/;
  assign sum_15[58] = _7155_ ^ _7154_ /*19082*/;
  assign _7156_ = _7155_ & _7154_ /*19081*/;
  assign _7157_ = inv_15[58] & r_14[58] /*19080*/;
  assign _7158_ = _7156_ | _7157_ /*19079*/;
  assign _7159_ = inv_15[59] ^ r_14[59] /*19077*/;
  assign sum_15[59] = _7159_ ^ _7158_ /*19076*/;
  assign _7160_ = _7159_ & _7158_ /*19075*/;
  assign _7161_ = inv_15[59] & r_14[59] /*19074*/;
  assign _7162_ = _7160_ | _7161_ /*19073*/;
  assign _7163_ = inv_15[60] ^ r_14[60] /*19071*/;
  assign sum_15[60] = _7163_ ^ _7162_ /*19070*/;
  assign _7164_ = _7163_ & _7162_ /*19069*/;
  assign _7165_ = inv_15[60] & r_14[60] /*19068*/;
  assign _7166_ = _7164_ | _7165_ /*19067*/;
  assign _7167_ = inv_15[61] ^ r_14[61] /*19065*/;
  assign sum_15[61] = _7167_ ^ _7166_ /*19064*/;
  assign _7168_ = _7167_ & _7166_ /*19063*/;
  assign _7169_ = inv_15[61] & r_14[61] /*19062*/;
  assign _7170_ = _7168_ | _7169_ /*19061*/;
  assign _7171_ = inv_15[62] ^ r_14[62] /*19059*/;
  assign sum_15[62] = _7171_ ^ _7170_ /*19058*/;
  assign _7172_ = _7171_ & _7170_ /*19057*/;
  assign _7173_ = inv_15[62] & r_14[62] /*19056*/;
  assign _7174_ = _7172_ | _7173_ /*19055*/;
  assign _7175_ = inv_15[63] ^ r_14[63] /*19053*/;
  assign sum_15[63] = _7175_ ^ _7174_ /*19052*/;
  assign _7176_ = _7175_ & _7174_ /*19051*/;
  assign _7177_ = inv_15[63] & r_14[63] /*19050*/;
  assign _7178_ = _7176_ | _7177_ /*19049*/;
  assign _7179_ = inv_15[64] ^ r_14[64] /*19047*/;
  assign sum_15[64] = _7179_ ^ _7178_ /*19046*/;
  assign _7180_ = _7179_ & _7178_ /*19045*/;
  assign _7181_ = inv_15[64] & r_14[64] /*19044*/;
  assign _7182_ = _7180_ | _7181_ /*19043*/;
  assign _7183_ = inv_15[65] ^ r_14[65] /*19041*/;
  assign sum_15[65] = _7183_ ^ _7182_ /*19040*/;
  assign _7184_ = _7183_ & _7182_ /*19039*/;
  assign _7185_ = inv_15[65] & r_14[65] /*19038*/;
  assign _7186_ = _7184_ | _7185_ /*19037*/;
  assign _7187_ = inv_15[66] ^ r_14[66] /*19035*/;
  assign sum_15[66] = _7187_ ^ _7186_ /*19034*/;
  assign _7188_ = _7187_ & _7186_ /*19033*/;
  assign _7189_ = inv_15[66] & r_14[66] /*19032*/;
  assign _7190_ = _7188_ | _7189_ /*19031*/;
  assign _7191_ = inv_15[67] ^ r_14[67] /*19029*/;
  assign sum_15[67] = _7191_ ^ _7190_ /*19028*/;
  assign _7192_ = _7191_ & _7190_ /*19027*/;
  assign _7193_ = inv_15[67] & r_14[67] /*19026*/;
  assign _7194_ = _7192_ | _7193_ /*19025*/;
  assign _7195_ = inv_15[68] ^ r_14[68] /*19023*/;
  assign sum_15[68] = _7195_ ^ _7194_ /*19022*/;
  assign _7196_ = _7195_ & _7194_ /*19021*/;
  assign _7197_ = inv_15[68] & r_14[68] /*19020*/;
  assign _7198_ = _7196_ | _7197_ /*19019*/;
  assign _7199_ = inv_15[69] ^ r_14[69] /*19017*/;
  assign sum_15[69] = _7199_ ^ _7198_ /*19016*/;
  assign _7200_ = _7199_ & _7198_ /*19015*/;
  assign _7201_ = inv_15[69] & r_14[69] /*19014*/;
  assign _7202_ = _7200_ | _7201_ /*19013*/;
  assign _7203_ = inv_15[70] ^ r_14[70] /*19011*/;
  assign sum_15[70] = _7203_ ^ _7202_ /*19010*/;
  assign _7204_ = _7203_ & _7202_ /*19009*/;
  assign _7205_ = inv_15[70] & r_14[70] /*19008*/;
  assign _7206_ = _7204_ | _7205_ /*19007*/;
  assign _7207_ = inv_15[71] ^ r_14[71] /*19005*/;
  assign sum_15[71] = _7207_ ^ _7206_ /*19004*/;
  assign _7208_ = _7207_ & _7206_ /*19003*/;
  assign _7209_ = inv_15[71] & r_14[71] /*19002*/;
  assign _7210_ = _7208_ | _7209_ /*19001*/;
  assign _7211_ = inv_15[72] ^ r_14[72] /*18999*/;
  assign sum_15[72] = _7211_ ^ _7210_ /*18998*/;
  assign _7212_ = _7211_ & _7210_ /*18997*/;
  assign _7213_ = inv_15[72] & r_14[72] /*18996*/;
  assign _7214_ = _7212_ | _7213_ /*18995*/;
  assign _7215_ = inv_15[73] ^ r_14[73] /*18993*/;
  assign sum_15[73] = _7215_ ^ _7214_ /*18992*/;
  assign _7216_ = _7215_ & _7214_ /*18991*/;
  assign _7217_ = inv_15[73] & r_14[73] /*18990*/;
  assign _7218_ = _7216_ | _7217_ /*18989*/;
  assign _7219_ = inv_15[74] ^ r_14[74] /*18987*/;
  assign sum_15[74] = _7219_ ^ _7218_ /*18986*/;
  assign _7220_ = _7219_ & _7218_ /*18985*/;
  assign _7221_ = inv_15[74] & r_14[74] /*18984*/;
  assign _7222_ = _7220_ | _7221_ /*18983*/;
  assign _7223_ = inv_15[75] ^ r_14[75] /*18981*/;
  assign sum_15[75] = _7223_ ^ _7222_ /*18980*/;
  assign _7224_ = _7223_ & _7222_ /*18979*/;
  assign _7225_ = inv_15[75] & r_14[75] /*18978*/;
  assign _7226_ = _7224_ | _7225_ /*18977*/;
  assign _7227_ = inv_15[76] ^ r_14[76] /*18975*/;
  assign sum_15[76] = _7227_ ^ _7226_ /*18974*/;
  assign _7228_ = _7227_ & _7226_ /*18973*/;
  assign _7229_ = inv_15[76] & r_14[76] /*18972*/;
  assign _7230_ = _7228_ | _7229_ /*18971*/;
  assign _7231_ = _7230_ ^ _7226_ /*18970*/;
  assign _7232_ = ~_7231_ /*18969*/;
  assign _7233_ = sum_15[76] & _7232_ /*18968*/;
  assign _7234_ = _7231_ & _7230_ /*18967*/;
  assign sum_15[77] = _7234_ | _7233_ /*18966*/;
  assign q[17] = ~sum_15[77] /*18965*/;
  assign m_15[0] = r_14[0] /*18964*/;
  assign m_15[1] = r_14[1] /*18963*/;
  assign m_15[2] = r_14[2] /*18962*/;
  assign m_15[3] = r_14[3] /*18961*/;
  assign m_15[4] = r_14[4] /*18960*/;
  assign m_15[5] = r_14[5] /*18959*/;
  assign m_15[6] = r_14[6] /*18958*/;
  assign m_15[7] = r_14[7] /*18957*/;
  assign m_15[8] = r_14[8] /*18956*/;
  assign m_15[9] = r_14[9] /*18955*/;
  assign m_15[10] = r_14[10] /*18954*/;
  assign m_15[11] = r_14[11] /*18953*/;
  assign m_15[12] = r_14[12] /*18952*/;
  assign m_15[13] = r_14[13] /*18951*/;
  assign m_15[14] = r_14[14] /*18950*/;
  assign m_15[15] = r_14[15] /*18949*/;
  assign m_15[16] = r_14[16] /*18948*/;
  assign m_15[17] = r_14[17] /*18947*/;
  assign m_15[18] = r_14[18] /*18946*/;
  assign m_15[19] = r_14[19] /*18945*/;
  assign m_15[20] = r_14[20] /*18944*/;
  assign m_15[21] = r_14[21] /*18943*/;
  assign m_15[22] = r_14[22] /*18942*/;
  assign m_15[23] = r_14[23] /*18941*/;
  assign m_15[24] = r_14[24] /*18940*/;
  assign m_15[25] = r_14[25] /*18939*/;
  assign m_15[26] = r_14[26] /*18938*/;
  assign m_15[27] = r_14[27] /*18937*/;
  assign m_15[28] = r_14[28] /*18936*/;
  assign m_15[29] = r_14[29] /*18935*/;
  assign m_15[30] = r_14[30] /*18934*/;
  assign m_15[31] = r_14[31] /*18933*/;
  assign m_15[32] = r_14[32] /*18932*/;
  assign m_15[33] = r_14[33] /*18931*/;
  assign m_15[34] = r_14[34] /*18930*/;
  assign m_15[35] = r_14[35] /*18929*/;
  assign m_15[36] = r_14[36] /*18928*/;
  assign m_15[37] = r_14[37] /*18927*/;
  assign m_15[38] = r_14[38] /*18926*/;
  assign m_15[39] = r_14[39] /*18925*/;
  assign m_15[40] = r_14[40] /*18924*/;
  assign m_15[41] = r_14[41] /*18923*/;
  assign m_15[42] = r_14[42] /*18922*/;
  assign m_15[43] = r_14[43] /*18921*/;
  assign m_15[44] = r_14[44] /*18920*/;
  assign m_15[45] = r_14[45] /*18919*/;
  assign m_15[46] = r_14[46] /*18918*/;
  assign m_15[47] = r_14[47] /*18917*/;
  assign m_15[48] = r_14[48] /*18916*/;
  assign m_15[49] = r_14[49] /*18915*/;
  assign m_15[50] = r_14[50] /*18914*/;
  assign m_15[51] = r_14[51] /*18913*/;
  assign m_15[52] = r_14[52] /*18912*/;
  assign m_15[53] = r_14[53] /*18911*/;
  assign m_15[54] = r_14[54] /*18910*/;
  assign m_15[55] = r_14[55] /*18909*/;
  assign m_15[56] = r_14[56] /*18908*/;
  assign m_15[57] = r_14[57] /*18907*/;
  assign m_15[58] = r_14[58] /*18906*/;
  assign m_15[59] = r_14[59] /*18905*/;
  assign m_15[60] = r_14[60] /*18904*/;
  assign m_15[61] = r_14[61] /*18903*/;
  assign m_15[62] = r_14[62] /*18902*/;
  assign m_15[63] = r_14[63] /*18901*/;
  assign m_15[64] = r_14[64] /*18900*/;
  assign m_15[65] = r_14[65] /*18899*/;
  assign m_15[66] = r_14[66] /*18898*/;
  assign m_15[67] = r_14[67] /*18897*/;
  assign m_15[68] = r_14[68] /*18896*/;
  assign m_15[69] = r_14[69] /*18895*/;
  assign m_15[70] = r_14[70] /*18894*/;
  assign m_15[71] = r_14[71] /*18893*/;
  assign m_15[72] = r_14[72] /*18892*/;
  assign m_15[73] = r_14[73] /*18891*/;
  assign m_15[74] = r_14[74] /*18890*/;
  assign m_15[75] = r_14[75] /*18889*/;
  assign m_15[76] = r_14[76] /*18888*/;
  assign m_15[77] = r_14[76] /*18887*/;
  assign _7236_ = ~q[17] /*18886*/;
  assign _7237_ = sum_15[0] & q[17] /*18885*/;
  assign _7238_ = m_15[0] & _7236_ /*18884*/;
  assign r_15[0] = _7238_ | _7237_ /*18883*/;
  assign _7239_ = ~q[17] /*18882*/;
  assign _7240_ = sum_15[1] & q[17] /*18881*/;
  assign _7241_ = m_15[1] & _7239_ /*18880*/;
  assign r_15[1] = _7241_ | _7240_ /*18879*/;
  assign _7242_ = ~q[17] /*18878*/;
  assign _7243_ = sum_15[2] & q[17] /*18877*/;
  assign _7244_ = m_15[2] & _7242_ /*18876*/;
  assign r_15[2] = _7244_ | _7243_ /*18875*/;
  assign _7245_ = ~q[17] /*18874*/;
  assign _7246_ = sum_15[3] & q[17] /*18873*/;
  assign _7247_ = m_15[3] & _7245_ /*18872*/;
  assign r_15[3] = _7247_ | _7246_ /*18871*/;
  assign _7248_ = ~q[17] /*18870*/;
  assign _7249_ = sum_15[4] & q[17] /*18869*/;
  assign _7250_ = m_15[4] & _7248_ /*18868*/;
  assign r_15[4] = _7250_ | _7249_ /*18867*/;
  assign _7251_ = ~q[17] /*18866*/;
  assign _7252_ = sum_15[5] & q[17] /*18865*/;
  assign _7253_ = m_15[5] & _7251_ /*18864*/;
  assign r_15[5] = _7253_ | _7252_ /*18863*/;
  assign _7254_ = ~q[17] /*18862*/;
  assign _7255_ = sum_15[6] & q[17] /*18861*/;
  assign _7256_ = m_15[6] & _7254_ /*18860*/;
  assign r_15[6] = _7256_ | _7255_ /*18859*/;
  assign _7257_ = ~q[17] /*18858*/;
  assign _7258_ = sum_15[7] & q[17] /*18857*/;
  assign _7259_ = m_15[7] & _7257_ /*18856*/;
  assign r_15[7] = _7259_ | _7258_ /*18855*/;
  assign _7260_ = ~q[17] /*18854*/;
  assign _7261_ = sum_15[8] & q[17] /*18853*/;
  assign _7262_ = m_15[8] & _7260_ /*18852*/;
  assign r_15[8] = _7262_ | _7261_ /*18851*/;
  assign _7263_ = ~q[17] /*18850*/;
  assign _7264_ = sum_15[9] & q[17] /*18849*/;
  assign _7265_ = m_15[9] & _7263_ /*18848*/;
  assign r_15[9] = _7265_ | _7264_ /*18847*/;
  assign _7266_ = ~q[17] /*18846*/;
  assign _7267_ = sum_15[10] & q[17] /*18845*/;
  assign _7268_ = m_15[10] & _7266_ /*18844*/;
  assign r_15[10] = _7268_ | _7267_ /*18843*/;
  assign _7269_ = ~q[17] /*18842*/;
  assign _7270_ = sum_15[11] & q[17] /*18841*/;
  assign _7271_ = m_15[11] & _7269_ /*18840*/;
  assign r_15[11] = _7271_ | _7270_ /*18839*/;
  assign _7272_ = ~q[17] /*18838*/;
  assign _7273_ = sum_15[12] & q[17] /*18837*/;
  assign _7274_ = m_15[12] & _7272_ /*18836*/;
  assign r_15[12] = _7274_ | _7273_ /*18835*/;
  assign _7275_ = ~q[17] /*18834*/;
  assign _7276_ = sum_15[13] & q[17] /*18833*/;
  assign _7277_ = m_15[13] & _7275_ /*18832*/;
  assign r_15[13] = _7277_ | _7276_ /*18831*/;
  assign _7278_ = ~q[17] /*18830*/;
  assign _7279_ = sum_15[14] & q[17] /*18829*/;
  assign _7280_ = m_15[14] & _7278_ /*18828*/;
  assign r_15[14] = _7280_ | _7279_ /*18827*/;
  assign _7281_ = ~q[17] /*18826*/;
  assign _7282_ = sum_15[15] & q[17] /*18825*/;
  assign _7283_ = m_15[15] & _7281_ /*18824*/;
  assign r_15[15] = _7283_ | _7282_ /*18823*/;
  assign _7284_ = ~q[17] /*18822*/;
  assign _7285_ = sum_15[16] & q[17] /*18821*/;
  assign _7286_ = m_15[16] & _7284_ /*18820*/;
  assign r_15[16] = _7286_ | _7285_ /*18819*/;
  assign _7287_ = ~q[17] /*18818*/;
  assign _7288_ = sum_15[17] & q[17] /*18817*/;
  assign _7289_ = m_15[17] & _7287_ /*18816*/;
  assign r_15[17] = _7289_ | _7288_ /*18815*/;
  assign _7290_ = ~q[17] /*18814*/;
  assign _7291_ = sum_15[18] & q[17] /*18813*/;
  assign _7292_ = m_15[18] & _7290_ /*18812*/;
  assign r_15[18] = _7292_ | _7291_ /*18811*/;
  assign _7293_ = ~q[17] /*18810*/;
  assign _7294_ = sum_15[19] & q[17] /*18809*/;
  assign _7295_ = m_15[19] & _7293_ /*18808*/;
  assign r_15[19] = _7295_ | _7294_ /*18807*/;
  assign _7296_ = ~q[17] /*18806*/;
  assign _7297_ = sum_15[20] & q[17] /*18805*/;
  assign _7298_ = m_15[20] & _7296_ /*18804*/;
  assign r_15[20] = _7298_ | _7297_ /*18803*/;
  assign _7299_ = ~q[17] /*18802*/;
  assign _7300_ = sum_15[21] & q[17] /*18801*/;
  assign _7301_ = m_15[21] & _7299_ /*18800*/;
  assign r_15[21] = _7301_ | _7300_ /*18799*/;
  assign _7302_ = ~q[17] /*18798*/;
  assign _7303_ = sum_15[22] & q[17] /*18797*/;
  assign _7304_ = m_15[22] & _7302_ /*18796*/;
  assign r_15[22] = _7304_ | _7303_ /*18795*/;
  assign _7305_ = ~q[17] /*18794*/;
  assign _7306_ = sum_15[23] & q[17] /*18793*/;
  assign _7307_ = m_15[23] & _7305_ /*18792*/;
  assign r_15[23] = _7307_ | _7306_ /*18791*/;
  assign _7308_ = ~q[17] /*18790*/;
  assign _7309_ = sum_15[24] & q[17] /*18789*/;
  assign _7310_ = m_15[24] & _7308_ /*18788*/;
  assign r_15[24] = _7310_ | _7309_ /*18787*/;
  assign _7311_ = ~q[17] /*18786*/;
  assign _7312_ = sum_15[25] & q[17] /*18785*/;
  assign _7313_ = m_15[25] & _7311_ /*18784*/;
  assign r_15[25] = _7313_ | _7312_ /*18783*/;
  assign _7314_ = ~q[17] /*18782*/;
  assign _7315_ = sum_15[26] & q[17] /*18781*/;
  assign _7316_ = m_15[26] & _7314_ /*18780*/;
  assign r_15[26] = _7316_ | _7315_ /*18779*/;
  assign _7317_ = ~q[17] /*18778*/;
  assign _7318_ = sum_15[27] & q[17] /*18777*/;
  assign _7319_ = m_15[27] & _7317_ /*18776*/;
  assign r_15[27] = _7319_ | _7318_ /*18775*/;
  assign _7320_ = ~q[17] /*18774*/;
  assign _7321_ = sum_15[28] & q[17] /*18773*/;
  assign _7322_ = m_15[28] & _7320_ /*18772*/;
  assign r_15[28] = _7322_ | _7321_ /*18771*/;
  assign _7323_ = ~q[17] /*18770*/;
  assign _7324_ = sum_15[29] & q[17] /*18769*/;
  assign _7325_ = m_15[29] & _7323_ /*18768*/;
  assign r_15[29] = _7325_ | _7324_ /*18767*/;
  assign _7326_ = ~q[17] /*18766*/;
  assign _7327_ = sum_15[30] & q[17] /*18765*/;
  assign _7328_ = m_15[30] & _7326_ /*18764*/;
  assign r_15[30] = _7328_ | _7327_ /*18763*/;
  assign _7329_ = ~q[17] /*18762*/;
  assign _7330_ = sum_15[31] & q[17] /*18761*/;
  assign _7331_ = m_15[31] & _7329_ /*18760*/;
  assign r_15[31] = _7331_ | _7330_ /*18759*/;
  assign _7332_ = ~q[17] /*18758*/;
  assign _7333_ = sum_15[32] & q[17] /*18757*/;
  assign _7334_ = m_15[32] & _7332_ /*18756*/;
  assign r_15[32] = _7334_ | _7333_ /*18755*/;
  assign _7335_ = ~q[17] /*18754*/;
  assign _7336_ = sum_15[33] & q[17] /*18753*/;
  assign _7337_ = m_15[33] & _7335_ /*18752*/;
  assign r_15[33] = _7337_ | _7336_ /*18751*/;
  assign _7338_ = ~q[17] /*18750*/;
  assign _7339_ = sum_15[34] & q[17] /*18749*/;
  assign _7340_ = m_15[34] & _7338_ /*18748*/;
  assign r_15[34] = _7340_ | _7339_ /*18747*/;
  assign _7341_ = ~q[17] /*18746*/;
  assign _7342_ = sum_15[35] & q[17] /*18745*/;
  assign _7343_ = m_15[35] & _7341_ /*18744*/;
  assign r_15[35] = _7343_ | _7342_ /*18743*/;
  assign _7344_ = ~q[17] /*18742*/;
  assign _7345_ = sum_15[36] & q[17] /*18741*/;
  assign _7346_ = m_15[36] & _7344_ /*18740*/;
  assign r_15[36] = _7346_ | _7345_ /*18739*/;
  assign _7347_ = ~q[17] /*18738*/;
  assign _7348_ = sum_15[37] & q[17] /*18737*/;
  assign _7349_ = m_15[37] & _7347_ /*18736*/;
  assign r_15[37] = _7349_ | _7348_ /*18735*/;
  assign _7350_ = ~q[17] /*18734*/;
  assign _7351_ = sum_15[38] & q[17] /*18733*/;
  assign _7352_ = m_15[38] & _7350_ /*18732*/;
  assign r_15[38] = _7352_ | _7351_ /*18731*/;
  assign _7353_ = ~q[17] /*18730*/;
  assign _7354_ = sum_15[39] & q[17] /*18729*/;
  assign _7355_ = m_15[39] & _7353_ /*18728*/;
  assign r_15[39] = _7355_ | _7354_ /*18727*/;
  assign _7356_ = ~q[17] /*18726*/;
  assign _7357_ = sum_15[40] & q[17] /*18725*/;
  assign _7358_ = m_15[40] & _7356_ /*18724*/;
  assign r_15[40] = _7358_ | _7357_ /*18723*/;
  assign _7359_ = ~q[17] /*18722*/;
  assign _7360_ = sum_15[41] & q[17] /*18721*/;
  assign _7361_ = m_15[41] & _7359_ /*18720*/;
  assign r_15[41] = _7361_ | _7360_ /*18719*/;
  assign _7362_ = ~q[17] /*18718*/;
  assign _7363_ = sum_15[42] & q[17] /*18717*/;
  assign _7364_ = m_15[42] & _7362_ /*18716*/;
  assign r_15[42] = _7364_ | _7363_ /*18715*/;
  assign _7365_ = ~q[17] /*18714*/;
  assign _7366_ = sum_15[43] & q[17] /*18713*/;
  assign _7367_ = m_15[43] & _7365_ /*18712*/;
  assign r_15[43] = _7367_ | _7366_ /*18711*/;
  assign _7368_ = ~q[17] /*18710*/;
  assign _7369_ = sum_15[44] & q[17] /*18709*/;
  assign _7370_ = m_15[44] & _7368_ /*18708*/;
  assign r_15[44] = _7370_ | _7369_ /*18707*/;
  assign _7371_ = ~q[17] /*18706*/;
  assign _7372_ = sum_15[45] & q[17] /*18705*/;
  assign _7373_ = m_15[45] & _7371_ /*18704*/;
  assign r_15[45] = _7373_ | _7372_ /*18703*/;
  assign _7374_ = ~q[17] /*18702*/;
  assign _7375_ = sum_15[46] & q[17] /*18701*/;
  assign _7376_ = m_15[46] & _7374_ /*18700*/;
  assign r_15[46] = _7376_ | _7375_ /*18699*/;
  assign _7377_ = ~q[17] /*18698*/;
  assign _7378_ = sum_15[47] & q[17] /*18697*/;
  assign _7379_ = m_15[47] & _7377_ /*18696*/;
  assign r_15[47] = _7379_ | _7378_ /*18695*/;
  assign _7380_ = ~q[17] /*18694*/;
  assign _7381_ = sum_15[48] & q[17] /*18693*/;
  assign _7382_ = m_15[48] & _7380_ /*18692*/;
  assign r_15[48] = _7382_ | _7381_ /*18691*/;
  assign _7383_ = ~q[17] /*18690*/;
  assign _7384_ = sum_15[49] & q[17] /*18689*/;
  assign _7385_ = m_15[49] & _7383_ /*18688*/;
  assign r_15[49] = _7385_ | _7384_ /*18687*/;
  assign _7386_ = ~q[17] /*18686*/;
  assign _7387_ = sum_15[50] & q[17] /*18685*/;
  assign _7388_ = m_15[50] & _7386_ /*18684*/;
  assign r_15[50] = _7388_ | _7387_ /*18683*/;
  assign _7389_ = ~q[17] /*18682*/;
  assign _7390_ = sum_15[51] & q[17] /*18681*/;
  assign _7391_ = m_15[51] & _7389_ /*18680*/;
  assign r_15[51] = _7391_ | _7390_ /*18679*/;
  assign _7392_ = ~q[17] /*18678*/;
  assign _7393_ = sum_15[52] & q[17] /*18677*/;
  assign _7394_ = m_15[52] & _7392_ /*18676*/;
  assign r_15[52] = _7394_ | _7393_ /*18675*/;
  assign _7395_ = ~q[17] /*18674*/;
  assign _7396_ = sum_15[53] & q[17] /*18673*/;
  assign _7397_ = m_15[53] & _7395_ /*18672*/;
  assign r_15[53] = _7397_ | _7396_ /*18671*/;
  assign _7398_ = ~q[17] /*18670*/;
  assign _7399_ = sum_15[54] & q[17] /*18669*/;
  assign _7400_ = m_15[54] & _7398_ /*18668*/;
  assign r_15[54] = _7400_ | _7399_ /*18667*/;
  assign _7401_ = ~q[17] /*18666*/;
  assign _7402_ = sum_15[55] & q[17] /*18665*/;
  assign _7403_ = m_15[55] & _7401_ /*18664*/;
  assign r_15[55] = _7403_ | _7402_ /*18663*/;
  assign _7404_ = ~q[17] /*18662*/;
  assign _7405_ = sum_15[56] & q[17] /*18661*/;
  assign _7406_ = m_15[56] & _7404_ /*18660*/;
  assign r_15[56] = _7406_ | _7405_ /*18659*/;
  assign _7407_ = ~q[17] /*18658*/;
  assign _7408_ = sum_15[57] & q[17] /*18657*/;
  assign _7409_ = m_15[57] & _7407_ /*18656*/;
  assign r_15[57] = _7409_ | _7408_ /*18655*/;
  assign _7410_ = ~q[17] /*18654*/;
  assign _7411_ = sum_15[58] & q[17] /*18653*/;
  assign _7412_ = m_15[58] & _7410_ /*18652*/;
  assign r_15[58] = _7412_ | _7411_ /*18651*/;
  assign _7413_ = ~q[17] /*18650*/;
  assign _7414_ = sum_15[59] & q[17] /*18649*/;
  assign _7415_ = m_15[59] & _7413_ /*18648*/;
  assign r_15[59] = _7415_ | _7414_ /*18647*/;
  assign _7416_ = ~q[17] /*18646*/;
  assign _7417_ = sum_15[60] & q[17] /*18645*/;
  assign _7418_ = m_15[60] & _7416_ /*18644*/;
  assign r_15[60] = _7418_ | _7417_ /*18643*/;
  assign _7419_ = ~q[17] /*18642*/;
  assign _7420_ = sum_15[61] & q[17] /*18641*/;
  assign _7421_ = m_15[61] & _7419_ /*18640*/;
  assign r_15[61] = _7421_ | _7420_ /*18639*/;
  assign _7422_ = ~q[17] /*18638*/;
  assign _7423_ = sum_15[62] & q[17] /*18637*/;
  assign _7424_ = m_15[62] & _7422_ /*18636*/;
  assign r_15[62] = _7424_ | _7423_ /*18635*/;
  assign _7425_ = ~q[17] /*18634*/;
  assign _7426_ = sum_15[63] & q[17] /*18633*/;
  assign _7427_ = m_15[63] & _7425_ /*18632*/;
  assign r_15[63] = _7427_ | _7426_ /*18631*/;
  assign _7428_ = ~q[17] /*18630*/;
  assign _7429_ = sum_15[64] & q[17] /*18629*/;
  assign _7430_ = m_15[64] & _7428_ /*18628*/;
  assign r_15[64] = _7430_ | _7429_ /*18627*/;
  assign _7431_ = ~q[17] /*18626*/;
  assign _7432_ = sum_15[65] & q[17] /*18625*/;
  assign _7433_ = m_15[65] & _7431_ /*18624*/;
  assign r_15[65] = _7433_ | _7432_ /*18623*/;
  assign _7434_ = ~q[17] /*18622*/;
  assign _7435_ = sum_15[66] & q[17] /*18621*/;
  assign _7436_ = m_15[66] & _7434_ /*18620*/;
  assign r_15[66] = _7436_ | _7435_ /*18619*/;
  assign _7437_ = ~q[17] /*18618*/;
  assign _7438_ = sum_15[67] & q[17] /*18617*/;
  assign _7439_ = m_15[67] & _7437_ /*18616*/;
  assign r_15[67] = _7439_ | _7438_ /*18615*/;
  assign _7440_ = ~q[17] /*18614*/;
  assign _7441_ = sum_15[68] & q[17] /*18613*/;
  assign _7442_ = m_15[68] & _7440_ /*18612*/;
  assign r_15[68] = _7442_ | _7441_ /*18611*/;
  assign _7443_ = ~q[17] /*18610*/;
  assign _7444_ = sum_15[69] & q[17] /*18609*/;
  assign _7445_ = m_15[69] & _7443_ /*18608*/;
  assign r_15[69] = _7445_ | _7444_ /*18607*/;
  assign _7446_ = ~q[17] /*18606*/;
  assign _7447_ = sum_15[70] & q[17] /*18605*/;
  assign _7448_ = m_15[70] & _7446_ /*18604*/;
  assign r_15[70] = _7448_ | _7447_ /*18603*/;
  assign _7449_ = ~q[17] /*18602*/;
  assign _7450_ = sum_15[71] & q[17] /*18601*/;
  assign _7451_ = m_15[71] & _7449_ /*18600*/;
  assign r_15[71] = _7451_ | _7450_ /*18599*/;
  assign _7452_ = ~q[17] /*18598*/;
  assign _7453_ = sum_15[72] & q[17] /*18597*/;
  assign _7454_ = m_15[72] & _7452_ /*18596*/;
  assign r_15[72] = _7454_ | _7453_ /*18595*/;
  assign _7455_ = ~q[17] /*18594*/;
  assign _7456_ = sum_15[73] & q[17] /*18593*/;
  assign _7457_ = m_15[73] & _7455_ /*18592*/;
  assign r_15[73] = _7457_ | _7456_ /*18591*/;
  assign _7458_ = ~q[17] /*18590*/;
  assign _7459_ = sum_15[74] & q[17] /*18589*/;
  assign _7460_ = m_15[74] & _7458_ /*18588*/;
  assign r_15[74] = _7460_ | _7459_ /*18587*/;
  assign _7461_ = ~q[17] /*18586*/;
  assign _7462_ = sum_15[75] & q[17] /*18585*/;
  assign _7463_ = m_15[75] & _7461_ /*18584*/;
  assign r_15[75] = _7463_ | _7462_ /*18583*/;
  assign _7464_ = ~q[17] /*18582*/;
  assign _7465_ = sum_15[76] & q[17] /*18581*/;
  assign _7466_ = m_15[76] & _7464_ /*18580*/;
  assign r_15[76] = _7466_ | _7465_ /*18579*/;
  assign _7467_ = ~q[17] /*18578*/;
  assign _7468_ = sum_15[77] & q[17] /*18577*/;
  assign _7469_ = m_15[77] & _7467_ /*18576*/;
  assign r_15[77] = _7469_ | _7468_ /*18575*/;
  assign inv_16[0] = oneWire /*18356*/;
  assign inv_16[1] = oneWire /*18350*/;
  assign inv_16[2] = oneWire /*18344*/;
  assign inv_16[3] = oneWire /*18338*/;
  assign inv_16[4] = oneWire /*18332*/;
  assign inv_16[5] = oneWire /*18326*/;
  assign inv_16[6] = oneWire /*18320*/;
  assign inv_16[7] = oneWire /*18314*/;
  assign inv_16[8] = oneWire /*18308*/;
  assign inv_16[9] = oneWire /*18302*/;
  assign inv_16[10] = oneWire /*18296*/;
  assign inv_16[11] = oneWire /*18290*/;
  assign inv_16[12] = oneWire /*18284*/;
  assign inv_16[13] = oneWire /*18278*/;
  assign inv_16[14] = oneWire /*18272*/;
  assign inv_16[15] = oneWire /*18266*/;
  assign inv_16[16] = ~div[0] /*18260*/;
  assign inv_16[17] = ~div[1] /*18254*/;
  assign inv_16[18] = ~div[2] /*18248*/;
  assign inv_16[19] = ~div[3] /*18242*/;
  assign inv_16[20] = ~div[4] /*18236*/;
  assign inv_16[21] = ~div[5] /*18230*/;
  assign inv_16[22] = ~div[6] /*18224*/;
  assign inv_16[23] = ~div[7] /*18218*/;
  assign inv_16[24] = ~div[8] /*18212*/;
  assign inv_16[25] = ~div[9] /*18206*/;
  assign inv_16[26] = ~div[10] /*18200*/;
  assign inv_16[27] = ~div[11] /*18194*/;
  assign inv_16[28] = ~div[12] /*18188*/;
  assign inv_16[29] = ~div[13] /*18182*/;
  assign inv_16[30] = ~div[14] /*18176*/;
  assign inv_16[31] = ~div[15] /*18170*/;
  assign inv_16[32] = ~div[16] /*18164*/;
  assign inv_16[33] = ~div[17] /*18158*/;
  assign inv_16[34] = ~div[18] /*18152*/;
  assign inv_16[35] = ~div[19] /*18146*/;
  assign inv_16[36] = ~div[20] /*18140*/;
  assign inv_16[37] = ~div[21] /*18134*/;
  assign inv_16[38] = ~div[22] /*18128*/;
  assign inv_16[39] = ~div[23] /*18122*/;
  assign inv_16[40] = ~div[24] /*18116*/;
  assign inv_16[41] = ~div[25] /*18110*/;
  assign inv_16[42] = ~div[26] /*18104*/;
  assign inv_16[43] = ~div[27] /*18098*/;
  assign inv_16[44] = ~div[28] /*18092*/;
  assign inv_16[45] = ~div[29] /*18086*/;
  assign inv_16[46] = ~div[30] /*18080*/;
  assign inv_16[47] = oneWire /*18074*/;
  assign inv_16[48] = oneWire /*18068*/;
  assign inv_16[49] = oneWire /*18062*/;
  assign inv_16[50] = oneWire /*18056*/;
  assign inv_16[51] = oneWire /*18050*/;
  assign inv_16[52] = oneWire /*18044*/;
  assign inv_16[53] = oneWire /*18038*/;
  assign inv_16[54] = oneWire /*18032*/;
  assign inv_16[55] = oneWire /*18026*/;
  assign inv_16[56] = oneWire /*18020*/;
  assign inv_16[57] = oneWire /*18014*/;
  assign inv_16[58] = oneWire /*18008*/;
  assign inv_16[59] = oneWire /*18002*/;
  assign inv_16[60] = oneWire /*17996*/;
  assign inv_16[61] = oneWire /*17990*/;
  assign inv_16[62] = oneWire /*17984*/;
  assign inv_16[63] = oneWire /*17978*/;
  assign inv_16[64] = oneWire /*17972*/;
  assign inv_16[65] = oneWire /*17966*/;
  assign inv_16[66] = oneWire /*17960*/;
  assign inv_16[67] = oneWire /*17954*/;
  assign inv_16[68] = oneWire /*17948*/;
  assign inv_16[69] = oneWire /*17942*/;
  assign inv_16[70] = oneWire /*17936*/;
  assign inv_16[71] = oneWire /*17930*/;
  assign inv_16[72] = oneWire /*17924*/;
  assign inv_16[73] = oneWire /*17918*/;
  assign inv_16[74] = oneWire /*17912*/;
  assign inv_16[75] = oneWire /*17906*/;
  assign inv_16[76] = oneWire /*17900*/;
  assign inv_16[77] = oneWire /*17894*/;
  assign _7470_ = inv_16[0] ^ r_15[0] /*18355*/;
  assign sum_16[0] = _7470_ ^ oneWire /*18354*/;
  assign _7471_ = _7470_ & oneWire /*18353*/;
  assign _7472_ = inv_16[0] & r_15[0] /*18352*/;
  assign _7473_ = _7471_ | _7472_ /*18351*/;
  assign _7474_ = inv_16[1] ^ r_15[1] /*18349*/;
  assign sum_16[1] = _7474_ ^ _7473_ /*18348*/;
  assign _7475_ = _7474_ & _7473_ /*18347*/;
  assign _7476_ = inv_16[1] & r_15[1] /*18346*/;
  assign _7477_ = _7475_ | _7476_ /*18345*/;
  assign _7478_ = inv_16[2] ^ r_15[2] /*18343*/;
  assign sum_16[2] = _7478_ ^ _7477_ /*18342*/;
  assign _7479_ = _7478_ & _7477_ /*18341*/;
  assign _7480_ = inv_16[2] & r_15[2] /*18340*/;
  assign _7481_ = _7479_ | _7480_ /*18339*/;
  assign _7482_ = inv_16[3] ^ r_15[3] /*18337*/;
  assign sum_16[3] = _7482_ ^ _7481_ /*18336*/;
  assign _7483_ = _7482_ & _7481_ /*18335*/;
  assign _7484_ = inv_16[3] & r_15[3] /*18334*/;
  assign _7485_ = _7483_ | _7484_ /*18333*/;
  assign _7486_ = inv_16[4] ^ r_15[4] /*18331*/;
  assign sum_16[4] = _7486_ ^ _7485_ /*18330*/;
  assign _7487_ = _7486_ & _7485_ /*18329*/;
  assign _7488_ = inv_16[4] & r_15[4] /*18328*/;
  assign _7489_ = _7487_ | _7488_ /*18327*/;
  assign _7490_ = inv_16[5] ^ r_15[5] /*18325*/;
  assign sum_16[5] = _7490_ ^ _7489_ /*18324*/;
  assign _7491_ = _7490_ & _7489_ /*18323*/;
  assign _7492_ = inv_16[5] & r_15[5] /*18322*/;
  assign _7493_ = _7491_ | _7492_ /*18321*/;
  assign _7494_ = inv_16[6] ^ r_15[6] /*18319*/;
  assign sum_16[6] = _7494_ ^ _7493_ /*18318*/;
  assign _7495_ = _7494_ & _7493_ /*18317*/;
  assign _7496_ = inv_16[6] & r_15[6] /*18316*/;
  assign _7497_ = _7495_ | _7496_ /*18315*/;
  assign _7498_ = inv_16[7] ^ r_15[7] /*18313*/;
  assign sum_16[7] = _7498_ ^ _7497_ /*18312*/;
  assign _7499_ = _7498_ & _7497_ /*18311*/;
  assign _7500_ = inv_16[7] & r_15[7] /*18310*/;
  assign _7501_ = _7499_ | _7500_ /*18309*/;
  assign _7502_ = inv_16[8] ^ r_15[8] /*18307*/;
  assign sum_16[8] = _7502_ ^ _7501_ /*18306*/;
  assign _7503_ = _7502_ & _7501_ /*18305*/;
  assign _7504_ = inv_16[8] & r_15[8] /*18304*/;
  assign _7505_ = _7503_ | _7504_ /*18303*/;
  assign _7506_ = inv_16[9] ^ r_15[9] /*18301*/;
  assign sum_16[9] = _7506_ ^ _7505_ /*18300*/;
  assign _7507_ = _7506_ & _7505_ /*18299*/;
  assign _7508_ = inv_16[9] & r_15[9] /*18298*/;
  assign _7509_ = _7507_ | _7508_ /*18297*/;
  assign _7510_ = inv_16[10] ^ r_15[10] /*18295*/;
  assign sum_16[10] = _7510_ ^ _7509_ /*18294*/;
  assign _7511_ = _7510_ & _7509_ /*18293*/;
  assign _7512_ = inv_16[10] & r_15[10] /*18292*/;
  assign _7513_ = _7511_ | _7512_ /*18291*/;
  assign _7514_ = inv_16[11] ^ r_15[11] /*18289*/;
  assign sum_16[11] = _7514_ ^ _7513_ /*18288*/;
  assign _7515_ = _7514_ & _7513_ /*18287*/;
  assign _7516_ = inv_16[11] & r_15[11] /*18286*/;
  assign _7517_ = _7515_ | _7516_ /*18285*/;
  assign _7518_ = inv_16[12] ^ r_15[12] /*18283*/;
  assign sum_16[12] = _7518_ ^ _7517_ /*18282*/;
  assign _7519_ = _7518_ & _7517_ /*18281*/;
  assign _7520_ = inv_16[12] & r_15[12] /*18280*/;
  assign _7521_ = _7519_ | _7520_ /*18279*/;
  assign _7522_ = inv_16[13] ^ r_15[13] /*18277*/;
  assign sum_16[13] = _7522_ ^ _7521_ /*18276*/;
  assign _7523_ = _7522_ & _7521_ /*18275*/;
  assign _7524_ = inv_16[13] & r_15[13] /*18274*/;
  assign _7525_ = _7523_ | _7524_ /*18273*/;
  assign _7526_ = inv_16[14] ^ r_15[14] /*18271*/;
  assign sum_16[14] = _7526_ ^ _7525_ /*18270*/;
  assign _7527_ = _7526_ & _7525_ /*18269*/;
  assign _7528_ = inv_16[14] & r_15[14] /*18268*/;
  assign _7529_ = _7527_ | _7528_ /*18267*/;
  assign _7530_ = inv_16[15] ^ r_15[15] /*18265*/;
  assign sum_16[15] = _7530_ ^ _7529_ /*18264*/;
  assign _7531_ = _7530_ & _7529_ /*18263*/;
  assign _7532_ = inv_16[15] & r_15[15] /*18262*/;
  assign _7533_ = _7531_ | _7532_ /*18261*/;
  assign _7534_ = inv_16[16] ^ r_15[16] /*18259*/;
  assign sum_16[16] = _7534_ ^ _7533_ /*18258*/;
  assign _7535_ = _7534_ & _7533_ /*18257*/;
  assign _7536_ = inv_16[16] & r_15[16] /*18256*/;
  assign _7537_ = _7535_ | _7536_ /*18255*/;
  assign _7538_ = inv_16[17] ^ r_15[17] /*18253*/;
  assign sum_16[17] = _7538_ ^ _7537_ /*18252*/;
  assign _7539_ = _7538_ & _7537_ /*18251*/;
  assign _7540_ = inv_16[17] & r_15[17] /*18250*/;
  assign _7541_ = _7539_ | _7540_ /*18249*/;
  assign _7542_ = inv_16[18] ^ r_15[18] /*18247*/;
  assign sum_16[18] = _7542_ ^ _7541_ /*18246*/;
  assign _7543_ = _7542_ & _7541_ /*18245*/;
  assign _7544_ = inv_16[18] & r_15[18] /*18244*/;
  assign _7545_ = _7543_ | _7544_ /*18243*/;
  assign _7546_ = inv_16[19] ^ r_15[19] /*18241*/;
  assign sum_16[19] = _7546_ ^ _7545_ /*18240*/;
  assign _7547_ = _7546_ & _7545_ /*18239*/;
  assign _7548_ = inv_16[19] & r_15[19] /*18238*/;
  assign _7549_ = _7547_ | _7548_ /*18237*/;
  assign _7550_ = inv_16[20] ^ r_15[20] /*18235*/;
  assign sum_16[20] = _7550_ ^ _7549_ /*18234*/;
  assign _7551_ = _7550_ & _7549_ /*18233*/;
  assign _7552_ = inv_16[20] & r_15[20] /*18232*/;
  assign _7553_ = _7551_ | _7552_ /*18231*/;
  assign _7554_ = inv_16[21] ^ r_15[21] /*18229*/;
  assign sum_16[21] = _7554_ ^ _7553_ /*18228*/;
  assign _7555_ = _7554_ & _7553_ /*18227*/;
  assign _7556_ = inv_16[21] & r_15[21] /*18226*/;
  assign _7557_ = _7555_ | _7556_ /*18225*/;
  assign _7558_ = inv_16[22] ^ r_15[22] /*18223*/;
  assign sum_16[22] = _7558_ ^ _7557_ /*18222*/;
  assign _7559_ = _7558_ & _7557_ /*18221*/;
  assign _7560_ = inv_16[22] & r_15[22] /*18220*/;
  assign _7561_ = _7559_ | _7560_ /*18219*/;
  assign _7562_ = inv_16[23] ^ r_15[23] /*18217*/;
  assign sum_16[23] = _7562_ ^ _7561_ /*18216*/;
  assign _7563_ = _7562_ & _7561_ /*18215*/;
  assign _7564_ = inv_16[23] & r_15[23] /*18214*/;
  assign _7565_ = _7563_ | _7564_ /*18213*/;
  assign _7566_ = inv_16[24] ^ r_15[24] /*18211*/;
  assign sum_16[24] = _7566_ ^ _7565_ /*18210*/;
  assign _7567_ = _7566_ & _7565_ /*18209*/;
  assign _7568_ = inv_16[24] & r_15[24] /*18208*/;
  assign _7569_ = _7567_ | _7568_ /*18207*/;
  assign _7570_ = inv_16[25] ^ r_15[25] /*18205*/;
  assign sum_16[25] = _7570_ ^ _7569_ /*18204*/;
  assign _7571_ = _7570_ & _7569_ /*18203*/;
  assign _7572_ = inv_16[25] & r_15[25] /*18202*/;
  assign _7573_ = _7571_ | _7572_ /*18201*/;
  assign _7574_ = inv_16[26] ^ r_15[26] /*18199*/;
  assign sum_16[26] = _7574_ ^ _7573_ /*18198*/;
  assign _7575_ = _7574_ & _7573_ /*18197*/;
  assign _7576_ = inv_16[26] & r_15[26] /*18196*/;
  assign _7577_ = _7575_ | _7576_ /*18195*/;
  assign _7578_ = inv_16[27] ^ r_15[27] /*18193*/;
  assign sum_16[27] = _7578_ ^ _7577_ /*18192*/;
  assign _7579_ = _7578_ & _7577_ /*18191*/;
  assign _7580_ = inv_16[27] & r_15[27] /*18190*/;
  assign _7581_ = _7579_ | _7580_ /*18189*/;
  assign _7582_ = inv_16[28] ^ r_15[28] /*18187*/;
  assign sum_16[28] = _7582_ ^ _7581_ /*18186*/;
  assign _7583_ = _7582_ & _7581_ /*18185*/;
  assign _7584_ = inv_16[28] & r_15[28] /*18184*/;
  assign _7585_ = _7583_ | _7584_ /*18183*/;
  assign _7586_ = inv_16[29] ^ r_15[29] /*18181*/;
  assign sum_16[29] = _7586_ ^ _7585_ /*18180*/;
  assign _7587_ = _7586_ & _7585_ /*18179*/;
  assign _7588_ = inv_16[29] & r_15[29] /*18178*/;
  assign _7589_ = _7587_ | _7588_ /*18177*/;
  assign _7590_ = inv_16[30] ^ r_15[30] /*18175*/;
  assign sum_16[30] = _7590_ ^ _7589_ /*18174*/;
  assign _7591_ = _7590_ & _7589_ /*18173*/;
  assign _7592_ = inv_16[30] & r_15[30] /*18172*/;
  assign _7593_ = _7591_ | _7592_ /*18171*/;
  assign _7594_ = inv_16[31] ^ r_15[31] /*18169*/;
  assign sum_16[31] = _7594_ ^ _7593_ /*18168*/;
  assign _7595_ = _7594_ & _7593_ /*18167*/;
  assign _7596_ = inv_16[31] & r_15[31] /*18166*/;
  assign _7597_ = _7595_ | _7596_ /*18165*/;
  assign _7598_ = inv_16[32] ^ r_15[32] /*18163*/;
  assign sum_16[32] = _7598_ ^ _7597_ /*18162*/;
  assign _7599_ = _7598_ & _7597_ /*18161*/;
  assign _7600_ = inv_16[32] & r_15[32] /*18160*/;
  assign _7601_ = _7599_ | _7600_ /*18159*/;
  assign _7602_ = inv_16[33] ^ r_15[33] /*18157*/;
  assign sum_16[33] = _7602_ ^ _7601_ /*18156*/;
  assign _7603_ = _7602_ & _7601_ /*18155*/;
  assign _7604_ = inv_16[33] & r_15[33] /*18154*/;
  assign _7605_ = _7603_ | _7604_ /*18153*/;
  assign _7606_ = inv_16[34] ^ r_15[34] /*18151*/;
  assign sum_16[34] = _7606_ ^ _7605_ /*18150*/;
  assign _7607_ = _7606_ & _7605_ /*18149*/;
  assign _7608_ = inv_16[34] & r_15[34] /*18148*/;
  assign _7609_ = _7607_ | _7608_ /*18147*/;
  assign _7610_ = inv_16[35] ^ r_15[35] /*18145*/;
  assign sum_16[35] = _7610_ ^ _7609_ /*18144*/;
  assign _7611_ = _7610_ & _7609_ /*18143*/;
  assign _7612_ = inv_16[35] & r_15[35] /*18142*/;
  assign _7613_ = _7611_ | _7612_ /*18141*/;
  assign _7614_ = inv_16[36] ^ r_15[36] /*18139*/;
  assign sum_16[36] = _7614_ ^ _7613_ /*18138*/;
  assign _7615_ = _7614_ & _7613_ /*18137*/;
  assign _7616_ = inv_16[36] & r_15[36] /*18136*/;
  assign _7617_ = _7615_ | _7616_ /*18135*/;
  assign _7618_ = inv_16[37] ^ r_15[37] /*18133*/;
  assign sum_16[37] = _7618_ ^ _7617_ /*18132*/;
  assign _7619_ = _7618_ & _7617_ /*18131*/;
  assign _7620_ = inv_16[37] & r_15[37] /*18130*/;
  assign _7621_ = _7619_ | _7620_ /*18129*/;
  assign _7622_ = inv_16[38] ^ r_15[38] /*18127*/;
  assign sum_16[38] = _7622_ ^ _7621_ /*18126*/;
  assign _7623_ = _7622_ & _7621_ /*18125*/;
  assign _7624_ = inv_16[38] & r_15[38] /*18124*/;
  assign _7625_ = _7623_ | _7624_ /*18123*/;
  assign _7626_ = inv_16[39] ^ r_15[39] /*18121*/;
  assign sum_16[39] = _7626_ ^ _7625_ /*18120*/;
  assign _7627_ = _7626_ & _7625_ /*18119*/;
  assign _7628_ = inv_16[39] & r_15[39] /*18118*/;
  assign _7629_ = _7627_ | _7628_ /*18117*/;
  assign _7630_ = inv_16[40] ^ r_15[40] /*18115*/;
  assign sum_16[40] = _7630_ ^ _7629_ /*18114*/;
  assign _7631_ = _7630_ & _7629_ /*18113*/;
  assign _7632_ = inv_16[40] & r_15[40] /*18112*/;
  assign _7633_ = _7631_ | _7632_ /*18111*/;
  assign _7634_ = inv_16[41] ^ r_15[41] /*18109*/;
  assign sum_16[41] = _7634_ ^ _7633_ /*18108*/;
  assign _7635_ = _7634_ & _7633_ /*18107*/;
  assign _7636_ = inv_16[41] & r_15[41] /*18106*/;
  assign _7637_ = _7635_ | _7636_ /*18105*/;
  assign _7638_ = inv_16[42] ^ r_15[42] /*18103*/;
  assign sum_16[42] = _7638_ ^ _7637_ /*18102*/;
  assign _7639_ = _7638_ & _7637_ /*18101*/;
  assign _7640_ = inv_16[42] & r_15[42] /*18100*/;
  assign _7641_ = _7639_ | _7640_ /*18099*/;
  assign _7642_ = inv_16[43] ^ r_15[43] /*18097*/;
  assign sum_16[43] = _7642_ ^ _7641_ /*18096*/;
  assign _7643_ = _7642_ & _7641_ /*18095*/;
  assign _7644_ = inv_16[43] & r_15[43] /*18094*/;
  assign _7645_ = _7643_ | _7644_ /*18093*/;
  assign _7646_ = inv_16[44] ^ r_15[44] /*18091*/;
  assign sum_16[44] = _7646_ ^ _7645_ /*18090*/;
  assign _7647_ = _7646_ & _7645_ /*18089*/;
  assign _7648_ = inv_16[44] & r_15[44] /*18088*/;
  assign _7649_ = _7647_ | _7648_ /*18087*/;
  assign _7650_ = inv_16[45] ^ r_15[45] /*18085*/;
  assign sum_16[45] = _7650_ ^ _7649_ /*18084*/;
  assign _7651_ = _7650_ & _7649_ /*18083*/;
  assign _7652_ = inv_16[45] & r_15[45] /*18082*/;
  assign _7653_ = _7651_ | _7652_ /*18081*/;
  assign _7654_ = inv_16[46] ^ r_15[46] /*18079*/;
  assign sum_16[46] = _7654_ ^ _7653_ /*18078*/;
  assign _7655_ = _7654_ & _7653_ /*18077*/;
  assign _7656_ = inv_16[46] & r_15[46] /*18076*/;
  assign _7657_ = _7655_ | _7656_ /*18075*/;
  assign _7658_ = inv_16[47] ^ r_15[47] /*18073*/;
  assign sum_16[47] = _7658_ ^ _7657_ /*18072*/;
  assign _7659_ = _7658_ & _7657_ /*18071*/;
  assign _7660_ = inv_16[47] & r_15[47] /*18070*/;
  assign _7661_ = _7659_ | _7660_ /*18069*/;
  assign _7662_ = inv_16[48] ^ r_15[48] /*18067*/;
  assign sum_16[48] = _7662_ ^ _7661_ /*18066*/;
  assign _7663_ = _7662_ & _7661_ /*18065*/;
  assign _7664_ = inv_16[48] & r_15[48] /*18064*/;
  assign _7665_ = _7663_ | _7664_ /*18063*/;
  assign _7666_ = inv_16[49] ^ r_15[49] /*18061*/;
  assign sum_16[49] = _7666_ ^ _7665_ /*18060*/;
  assign _7667_ = _7666_ & _7665_ /*18059*/;
  assign _7668_ = inv_16[49] & r_15[49] /*18058*/;
  assign _7669_ = _7667_ | _7668_ /*18057*/;
  assign _7670_ = inv_16[50] ^ r_15[50] /*18055*/;
  assign sum_16[50] = _7670_ ^ _7669_ /*18054*/;
  assign _7671_ = _7670_ & _7669_ /*18053*/;
  assign _7672_ = inv_16[50] & r_15[50] /*18052*/;
  assign _7673_ = _7671_ | _7672_ /*18051*/;
  assign _7674_ = inv_16[51] ^ r_15[51] /*18049*/;
  assign sum_16[51] = _7674_ ^ _7673_ /*18048*/;
  assign _7675_ = _7674_ & _7673_ /*18047*/;
  assign _7676_ = inv_16[51] & r_15[51] /*18046*/;
  assign _7677_ = _7675_ | _7676_ /*18045*/;
  assign _7678_ = inv_16[52] ^ r_15[52] /*18043*/;
  assign sum_16[52] = _7678_ ^ _7677_ /*18042*/;
  assign _7679_ = _7678_ & _7677_ /*18041*/;
  assign _7680_ = inv_16[52] & r_15[52] /*18040*/;
  assign _7681_ = _7679_ | _7680_ /*18039*/;
  assign _7682_ = inv_16[53] ^ r_15[53] /*18037*/;
  assign sum_16[53] = _7682_ ^ _7681_ /*18036*/;
  assign _7683_ = _7682_ & _7681_ /*18035*/;
  assign _7684_ = inv_16[53] & r_15[53] /*18034*/;
  assign _7685_ = _7683_ | _7684_ /*18033*/;
  assign _7686_ = inv_16[54] ^ r_15[54] /*18031*/;
  assign sum_16[54] = _7686_ ^ _7685_ /*18030*/;
  assign _7687_ = _7686_ & _7685_ /*18029*/;
  assign _7688_ = inv_16[54] & r_15[54] /*18028*/;
  assign _7689_ = _7687_ | _7688_ /*18027*/;
  assign _7690_ = inv_16[55] ^ r_15[55] /*18025*/;
  assign sum_16[55] = _7690_ ^ _7689_ /*18024*/;
  assign _7691_ = _7690_ & _7689_ /*18023*/;
  assign _7692_ = inv_16[55] & r_15[55] /*18022*/;
  assign _7693_ = _7691_ | _7692_ /*18021*/;
  assign _7694_ = inv_16[56] ^ r_15[56] /*18019*/;
  assign sum_16[56] = _7694_ ^ _7693_ /*18018*/;
  assign _7695_ = _7694_ & _7693_ /*18017*/;
  assign _7696_ = inv_16[56] & r_15[56] /*18016*/;
  assign _7697_ = _7695_ | _7696_ /*18015*/;
  assign _7698_ = inv_16[57] ^ r_15[57] /*18013*/;
  assign sum_16[57] = _7698_ ^ _7697_ /*18012*/;
  assign _7699_ = _7698_ & _7697_ /*18011*/;
  assign _7700_ = inv_16[57] & r_15[57] /*18010*/;
  assign _7701_ = _7699_ | _7700_ /*18009*/;
  assign _7702_ = inv_16[58] ^ r_15[58] /*18007*/;
  assign sum_16[58] = _7702_ ^ _7701_ /*18006*/;
  assign _7703_ = _7702_ & _7701_ /*18005*/;
  assign _7704_ = inv_16[58] & r_15[58] /*18004*/;
  assign _7705_ = _7703_ | _7704_ /*18003*/;
  assign _7706_ = inv_16[59] ^ r_15[59] /*18001*/;
  assign sum_16[59] = _7706_ ^ _7705_ /*18000*/;
  assign _7707_ = _7706_ & _7705_ /*17999*/;
  assign _7708_ = inv_16[59] & r_15[59] /*17998*/;
  assign _7709_ = _7707_ | _7708_ /*17997*/;
  assign _7710_ = inv_16[60] ^ r_15[60] /*17995*/;
  assign sum_16[60] = _7710_ ^ _7709_ /*17994*/;
  assign _7711_ = _7710_ & _7709_ /*17993*/;
  assign _7712_ = inv_16[60] & r_15[60] /*17992*/;
  assign _7713_ = _7711_ | _7712_ /*17991*/;
  assign _7714_ = inv_16[61] ^ r_15[61] /*17989*/;
  assign sum_16[61] = _7714_ ^ _7713_ /*17988*/;
  assign _7715_ = _7714_ & _7713_ /*17987*/;
  assign _7716_ = inv_16[61] & r_15[61] /*17986*/;
  assign _7717_ = _7715_ | _7716_ /*17985*/;
  assign _7718_ = inv_16[62] ^ r_15[62] /*17983*/;
  assign sum_16[62] = _7718_ ^ _7717_ /*17982*/;
  assign _7719_ = _7718_ & _7717_ /*17981*/;
  assign _7720_ = inv_16[62] & r_15[62] /*17980*/;
  assign _7721_ = _7719_ | _7720_ /*17979*/;
  assign _7722_ = inv_16[63] ^ r_15[63] /*17977*/;
  assign sum_16[63] = _7722_ ^ _7721_ /*17976*/;
  assign _7723_ = _7722_ & _7721_ /*17975*/;
  assign _7724_ = inv_16[63] & r_15[63] /*17974*/;
  assign _7725_ = _7723_ | _7724_ /*17973*/;
  assign _7726_ = inv_16[64] ^ r_15[64] /*17971*/;
  assign sum_16[64] = _7726_ ^ _7725_ /*17970*/;
  assign _7727_ = _7726_ & _7725_ /*17969*/;
  assign _7728_ = inv_16[64] & r_15[64] /*17968*/;
  assign _7729_ = _7727_ | _7728_ /*17967*/;
  assign _7730_ = inv_16[65] ^ r_15[65] /*17965*/;
  assign sum_16[65] = _7730_ ^ _7729_ /*17964*/;
  assign _7731_ = _7730_ & _7729_ /*17963*/;
  assign _7732_ = inv_16[65] & r_15[65] /*17962*/;
  assign _7733_ = _7731_ | _7732_ /*17961*/;
  assign _7734_ = inv_16[66] ^ r_15[66] /*17959*/;
  assign sum_16[66] = _7734_ ^ _7733_ /*17958*/;
  assign _7735_ = _7734_ & _7733_ /*17957*/;
  assign _7736_ = inv_16[66] & r_15[66] /*17956*/;
  assign _7737_ = _7735_ | _7736_ /*17955*/;
  assign _7738_ = inv_16[67] ^ r_15[67] /*17953*/;
  assign sum_16[67] = _7738_ ^ _7737_ /*17952*/;
  assign _7739_ = _7738_ & _7737_ /*17951*/;
  assign _7740_ = inv_16[67] & r_15[67] /*17950*/;
  assign _7741_ = _7739_ | _7740_ /*17949*/;
  assign _7742_ = inv_16[68] ^ r_15[68] /*17947*/;
  assign sum_16[68] = _7742_ ^ _7741_ /*17946*/;
  assign _7743_ = _7742_ & _7741_ /*17945*/;
  assign _7744_ = inv_16[68] & r_15[68] /*17944*/;
  assign _7745_ = _7743_ | _7744_ /*17943*/;
  assign _7746_ = inv_16[69] ^ r_15[69] /*17941*/;
  assign sum_16[69] = _7746_ ^ _7745_ /*17940*/;
  assign _7747_ = _7746_ & _7745_ /*17939*/;
  assign _7748_ = inv_16[69] & r_15[69] /*17938*/;
  assign _7749_ = _7747_ | _7748_ /*17937*/;
  assign _7750_ = inv_16[70] ^ r_15[70] /*17935*/;
  assign sum_16[70] = _7750_ ^ _7749_ /*17934*/;
  assign _7751_ = _7750_ & _7749_ /*17933*/;
  assign _7752_ = inv_16[70] & r_15[70] /*17932*/;
  assign _7753_ = _7751_ | _7752_ /*17931*/;
  assign _7754_ = inv_16[71] ^ r_15[71] /*17929*/;
  assign sum_16[71] = _7754_ ^ _7753_ /*17928*/;
  assign _7755_ = _7754_ & _7753_ /*17927*/;
  assign _7756_ = inv_16[71] & r_15[71] /*17926*/;
  assign _7757_ = _7755_ | _7756_ /*17925*/;
  assign _7758_ = inv_16[72] ^ r_15[72] /*17923*/;
  assign sum_16[72] = _7758_ ^ _7757_ /*17922*/;
  assign _7759_ = _7758_ & _7757_ /*17921*/;
  assign _7760_ = inv_16[72] & r_15[72] /*17920*/;
  assign _7761_ = _7759_ | _7760_ /*17919*/;
  assign _7762_ = inv_16[73] ^ r_15[73] /*17917*/;
  assign sum_16[73] = _7762_ ^ _7761_ /*17916*/;
  assign _7763_ = _7762_ & _7761_ /*17915*/;
  assign _7764_ = inv_16[73] & r_15[73] /*17914*/;
  assign _7765_ = _7763_ | _7764_ /*17913*/;
  assign _7766_ = inv_16[74] ^ r_15[74] /*17911*/;
  assign sum_16[74] = _7766_ ^ _7765_ /*17910*/;
  assign _7767_ = _7766_ & _7765_ /*17909*/;
  assign _7768_ = inv_16[74] & r_15[74] /*17908*/;
  assign _7769_ = _7767_ | _7768_ /*17907*/;
  assign _7770_ = inv_16[75] ^ r_15[75] /*17905*/;
  assign sum_16[75] = _7770_ ^ _7769_ /*17904*/;
  assign _7771_ = _7770_ & _7769_ /*17903*/;
  assign _7772_ = inv_16[75] & r_15[75] /*17902*/;
  assign _7773_ = _7771_ | _7772_ /*17901*/;
  assign _7774_ = inv_16[76] ^ r_15[76] /*17899*/;
  assign sum_16[76] = _7774_ ^ _7773_ /*17898*/;
  assign _7775_ = _7774_ & _7773_ /*17897*/;
  assign _7776_ = inv_16[76] & r_15[76] /*17896*/;
  assign _7777_ = _7775_ | _7776_ /*17895*/;
  assign _7778_ = inv_16[77] ^ r_15[77] /*17893*/;
  assign sum_16[77] = _7778_ ^ _7777_ /*17892*/;
  assign _7779_ = _7778_ & _7777_ /*17891*/;
  assign _7780_ = inv_16[77] & r_15[77] /*17890*/;
  assign _7781_ = _7779_ | _7780_ /*17889*/;
  assign _7782_ = _7781_ ^ _7777_ /*17888*/;
  assign _7783_ = ~_7782_ /*17887*/;
  assign _7784_ = sum_16[77] & _7783_ /*17886*/;
  assign _7785_ = _7782_ & _7781_ /*17885*/;
  assign sum_16[78] = _7785_ | _7784_ /*17884*/;
  assign q[16] = ~sum_16[78] /*17883*/;
  assign m_16[0] = r_15[0] /*17882*/;
  assign m_16[1] = r_15[1] /*17881*/;
  assign m_16[2] = r_15[2] /*17880*/;
  assign m_16[3] = r_15[3] /*17879*/;
  assign m_16[4] = r_15[4] /*17878*/;
  assign m_16[5] = r_15[5] /*17877*/;
  assign m_16[6] = r_15[6] /*17876*/;
  assign m_16[7] = r_15[7] /*17875*/;
  assign m_16[8] = r_15[8] /*17874*/;
  assign m_16[9] = r_15[9] /*17873*/;
  assign m_16[10] = r_15[10] /*17872*/;
  assign m_16[11] = r_15[11] /*17871*/;
  assign m_16[12] = r_15[12] /*17870*/;
  assign m_16[13] = r_15[13] /*17869*/;
  assign m_16[14] = r_15[14] /*17868*/;
  assign m_16[15] = r_15[15] /*17867*/;
  assign m_16[16] = r_15[16] /*17866*/;
  assign m_16[17] = r_15[17] /*17865*/;
  assign m_16[18] = r_15[18] /*17864*/;
  assign m_16[19] = r_15[19] /*17863*/;
  assign m_16[20] = r_15[20] /*17862*/;
  assign m_16[21] = r_15[21] /*17861*/;
  assign m_16[22] = r_15[22] /*17860*/;
  assign m_16[23] = r_15[23] /*17859*/;
  assign m_16[24] = r_15[24] /*17858*/;
  assign m_16[25] = r_15[25] /*17857*/;
  assign m_16[26] = r_15[26] /*17856*/;
  assign m_16[27] = r_15[27] /*17855*/;
  assign m_16[28] = r_15[28] /*17854*/;
  assign m_16[29] = r_15[29] /*17853*/;
  assign m_16[30] = r_15[30] /*17852*/;
  assign m_16[31] = r_15[31] /*17851*/;
  assign m_16[32] = r_15[32] /*17850*/;
  assign m_16[33] = r_15[33] /*17849*/;
  assign m_16[34] = r_15[34] /*17848*/;
  assign m_16[35] = r_15[35] /*17847*/;
  assign m_16[36] = r_15[36] /*17846*/;
  assign m_16[37] = r_15[37] /*17845*/;
  assign m_16[38] = r_15[38] /*17844*/;
  assign m_16[39] = r_15[39] /*17843*/;
  assign m_16[40] = r_15[40] /*17842*/;
  assign m_16[41] = r_15[41] /*17841*/;
  assign m_16[42] = r_15[42] /*17840*/;
  assign m_16[43] = r_15[43] /*17839*/;
  assign m_16[44] = r_15[44] /*17838*/;
  assign m_16[45] = r_15[45] /*17837*/;
  assign m_16[46] = r_15[46] /*17836*/;
  assign m_16[47] = r_15[47] /*17835*/;
  assign m_16[48] = r_15[48] /*17834*/;
  assign m_16[49] = r_15[49] /*17833*/;
  assign m_16[50] = r_15[50] /*17832*/;
  assign m_16[51] = r_15[51] /*17831*/;
  assign m_16[52] = r_15[52] /*17830*/;
  assign m_16[53] = r_15[53] /*17829*/;
  assign m_16[54] = r_15[54] /*17828*/;
  assign m_16[55] = r_15[55] /*17827*/;
  assign m_16[56] = r_15[56] /*17826*/;
  assign m_16[57] = r_15[57] /*17825*/;
  assign m_16[58] = r_15[58] /*17824*/;
  assign m_16[59] = r_15[59] /*17823*/;
  assign m_16[60] = r_15[60] /*17822*/;
  assign m_16[61] = r_15[61] /*17821*/;
  assign m_16[62] = r_15[62] /*17820*/;
  assign m_16[63] = r_15[63] /*17819*/;
  assign m_16[64] = r_15[64] /*17818*/;
  assign m_16[65] = r_15[65] /*17817*/;
  assign m_16[66] = r_15[66] /*17816*/;
  assign m_16[67] = r_15[67] /*17815*/;
  assign m_16[68] = r_15[68] /*17814*/;
  assign m_16[69] = r_15[69] /*17813*/;
  assign m_16[70] = r_15[70] /*17812*/;
  assign m_16[71] = r_15[71] /*17811*/;
  assign m_16[72] = r_15[72] /*17810*/;
  assign m_16[73] = r_15[73] /*17809*/;
  assign m_16[74] = r_15[74] /*17808*/;
  assign m_16[75] = r_15[75] /*17807*/;
  assign m_16[76] = r_15[76] /*17806*/;
  assign m_16[77] = r_15[77] /*17805*/;
  assign m_16[78] = r_15[77] /*17804*/;
  assign _7787_ = ~q[16] /*17803*/;
  assign _7788_ = sum_16[0] & q[16] /*17802*/;
  assign _7789_ = m_16[0] & _7787_ /*17801*/;
  assign r_16[0] = _7789_ | _7788_ /*17800*/;
  assign _7790_ = ~q[16] /*17799*/;
  assign _7791_ = sum_16[1] & q[16] /*17798*/;
  assign _7792_ = m_16[1] & _7790_ /*17797*/;
  assign r_16[1] = _7792_ | _7791_ /*17796*/;
  assign _7793_ = ~q[16] /*17795*/;
  assign _7794_ = sum_16[2] & q[16] /*17794*/;
  assign _7795_ = m_16[2] & _7793_ /*17793*/;
  assign r_16[2] = _7795_ | _7794_ /*17792*/;
  assign _7796_ = ~q[16] /*17791*/;
  assign _7797_ = sum_16[3] & q[16] /*17790*/;
  assign _7798_ = m_16[3] & _7796_ /*17789*/;
  assign r_16[3] = _7798_ | _7797_ /*17788*/;
  assign _7799_ = ~q[16] /*17787*/;
  assign _7800_ = sum_16[4] & q[16] /*17786*/;
  assign _7801_ = m_16[4] & _7799_ /*17785*/;
  assign r_16[4] = _7801_ | _7800_ /*17784*/;
  assign _7802_ = ~q[16] /*17783*/;
  assign _7803_ = sum_16[5] & q[16] /*17782*/;
  assign _7804_ = m_16[5] & _7802_ /*17781*/;
  assign r_16[5] = _7804_ | _7803_ /*17780*/;
  assign _7805_ = ~q[16] /*17779*/;
  assign _7806_ = sum_16[6] & q[16] /*17778*/;
  assign _7807_ = m_16[6] & _7805_ /*17777*/;
  assign r_16[6] = _7807_ | _7806_ /*17776*/;
  assign _7808_ = ~q[16] /*17775*/;
  assign _7809_ = sum_16[7] & q[16] /*17774*/;
  assign _7810_ = m_16[7] & _7808_ /*17773*/;
  assign r_16[7] = _7810_ | _7809_ /*17772*/;
  assign _7811_ = ~q[16] /*17771*/;
  assign _7812_ = sum_16[8] & q[16] /*17770*/;
  assign _7813_ = m_16[8] & _7811_ /*17769*/;
  assign r_16[8] = _7813_ | _7812_ /*17768*/;
  assign _7814_ = ~q[16] /*17767*/;
  assign _7815_ = sum_16[9] & q[16] /*17766*/;
  assign _7816_ = m_16[9] & _7814_ /*17765*/;
  assign r_16[9] = _7816_ | _7815_ /*17764*/;
  assign _7817_ = ~q[16] /*17763*/;
  assign _7818_ = sum_16[10] & q[16] /*17762*/;
  assign _7819_ = m_16[10] & _7817_ /*17761*/;
  assign r_16[10] = _7819_ | _7818_ /*17760*/;
  assign _7820_ = ~q[16] /*17759*/;
  assign _7821_ = sum_16[11] & q[16] /*17758*/;
  assign _7822_ = m_16[11] & _7820_ /*17757*/;
  assign r_16[11] = _7822_ | _7821_ /*17756*/;
  assign _7823_ = ~q[16] /*17755*/;
  assign _7824_ = sum_16[12] & q[16] /*17754*/;
  assign _7825_ = m_16[12] & _7823_ /*17753*/;
  assign r_16[12] = _7825_ | _7824_ /*17752*/;
  assign _7826_ = ~q[16] /*17751*/;
  assign _7827_ = sum_16[13] & q[16] /*17750*/;
  assign _7828_ = m_16[13] & _7826_ /*17749*/;
  assign r_16[13] = _7828_ | _7827_ /*17748*/;
  assign _7829_ = ~q[16] /*17747*/;
  assign _7830_ = sum_16[14] & q[16] /*17746*/;
  assign _7831_ = m_16[14] & _7829_ /*17745*/;
  assign r_16[14] = _7831_ | _7830_ /*17744*/;
  assign _7832_ = ~q[16] /*17743*/;
  assign _7833_ = sum_16[15] & q[16] /*17742*/;
  assign _7834_ = m_16[15] & _7832_ /*17741*/;
  assign r_16[15] = _7834_ | _7833_ /*17740*/;
  assign _7835_ = ~q[16] /*17739*/;
  assign _7836_ = sum_16[16] & q[16] /*17738*/;
  assign _7837_ = m_16[16] & _7835_ /*17737*/;
  assign r_16[16] = _7837_ | _7836_ /*17736*/;
  assign _7838_ = ~q[16] /*17735*/;
  assign _7839_ = sum_16[17] & q[16] /*17734*/;
  assign _7840_ = m_16[17] & _7838_ /*17733*/;
  assign r_16[17] = _7840_ | _7839_ /*17732*/;
  assign _7841_ = ~q[16] /*17731*/;
  assign _7842_ = sum_16[18] & q[16] /*17730*/;
  assign _7843_ = m_16[18] & _7841_ /*17729*/;
  assign r_16[18] = _7843_ | _7842_ /*17728*/;
  assign _7844_ = ~q[16] /*17727*/;
  assign _7845_ = sum_16[19] & q[16] /*17726*/;
  assign _7846_ = m_16[19] & _7844_ /*17725*/;
  assign r_16[19] = _7846_ | _7845_ /*17724*/;
  assign _7847_ = ~q[16] /*17723*/;
  assign _7848_ = sum_16[20] & q[16] /*17722*/;
  assign _7849_ = m_16[20] & _7847_ /*17721*/;
  assign r_16[20] = _7849_ | _7848_ /*17720*/;
  assign _7850_ = ~q[16] /*17719*/;
  assign _7851_ = sum_16[21] & q[16] /*17718*/;
  assign _7852_ = m_16[21] & _7850_ /*17717*/;
  assign r_16[21] = _7852_ | _7851_ /*17716*/;
  assign _7853_ = ~q[16] /*17715*/;
  assign _7854_ = sum_16[22] & q[16] /*17714*/;
  assign _7855_ = m_16[22] & _7853_ /*17713*/;
  assign r_16[22] = _7855_ | _7854_ /*17712*/;
  assign _7856_ = ~q[16] /*17711*/;
  assign _7857_ = sum_16[23] & q[16] /*17710*/;
  assign _7858_ = m_16[23] & _7856_ /*17709*/;
  assign r_16[23] = _7858_ | _7857_ /*17708*/;
  assign _7859_ = ~q[16] /*17707*/;
  assign _7860_ = sum_16[24] & q[16] /*17706*/;
  assign _7861_ = m_16[24] & _7859_ /*17705*/;
  assign r_16[24] = _7861_ | _7860_ /*17704*/;
  assign _7862_ = ~q[16] /*17703*/;
  assign _7863_ = sum_16[25] & q[16] /*17702*/;
  assign _7864_ = m_16[25] & _7862_ /*17701*/;
  assign r_16[25] = _7864_ | _7863_ /*17700*/;
  assign _7865_ = ~q[16] /*17699*/;
  assign _7866_ = sum_16[26] & q[16] /*17698*/;
  assign _7867_ = m_16[26] & _7865_ /*17697*/;
  assign r_16[26] = _7867_ | _7866_ /*17696*/;
  assign _7868_ = ~q[16] /*17695*/;
  assign _7869_ = sum_16[27] & q[16] /*17694*/;
  assign _7870_ = m_16[27] & _7868_ /*17693*/;
  assign r_16[27] = _7870_ | _7869_ /*17692*/;
  assign _7871_ = ~q[16] /*17691*/;
  assign _7872_ = sum_16[28] & q[16] /*17690*/;
  assign _7873_ = m_16[28] & _7871_ /*17689*/;
  assign r_16[28] = _7873_ | _7872_ /*17688*/;
  assign _7874_ = ~q[16] /*17687*/;
  assign _7875_ = sum_16[29] & q[16] /*17686*/;
  assign _7876_ = m_16[29] & _7874_ /*17685*/;
  assign r_16[29] = _7876_ | _7875_ /*17684*/;
  assign _7877_ = ~q[16] /*17683*/;
  assign _7878_ = sum_16[30] & q[16] /*17682*/;
  assign _7879_ = m_16[30] & _7877_ /*17681*/;
  assign r_16[30] = _7879_ | _7878_ /*17680*/;
  assign _7880_ = ~q[16] /*17679*/;
  assign _7881_ = sum_16[31] & q[16] /*17678*/;
  assign _7882_ = m_16[31] & _7880_ /*17677*/;
  assign r_16[31] = _7882_ | _7881_ /*17676*/;
  assign _7883_ = ~q[16] /*17675*/;
  assign _7884_ = sum_16[32] & q[16] /*17674*/;
  assign _7885_ = m_16[32] & _7883_ /*17673*/;
  assign r_16[32] = _7885_ | _7884_ /*17672*/;
  assign _7886_ = ~q[16] /*17671*/;
  assign _7887_ = sum_16[33] & q[16] /*17670*/;
  assign _7888_ = m_16[33] & _7886_ /*17669*/;
  assign r_16[33] = _7888_ | _7887_ /*17668*/;
  assign _7889_ = ~q[16] /*17667*/;
  assign _7890_ = sum_16[34] & q[16] /*17666*/;
  assign _7891_ = m_16[34] & _7889_ /*17665*/;
  assign r_16[34] = _7891_ | _7890_ /*17664*/;
  assign _7892_ = ~q[16] /*17663*/;
  assign _7893_ = sum_16[35] & q[16] /*17662*/;
  assign _7894_ = m_16[35] & _7892_ /*17661*/;
  assign r_16[35] = _7894_ | _7893_ /*17660*/;
  assign _7895_ = ~q[16] /*17659*/;
  assign _7896_ = sum_16[36] & q[16] /*17658*/;
  assign _7897_ = m_16[36] & _7895_ /*17657*/;
  assign r_16[36] = _7897_ | _7896_ /*17656*/;
  assign _7898_ = ~q[16] /*17655*/;
  assign _7899_ = sum_16[37] & q[16] /*17654*/;
  assign _7900_ = m_16[37] & _7898_ /*17653*/;
  assign r_16[37] = _7900_ | _7899_ /*17652*/;
  assign _7901_ = ~q[16] /*17651*/;
  assign _7902_ = sum_16[38] & q[16] /*17650*/;
  assign _7903_ = m_16[38] & _7901_ /*17649*/;
  assign r_16[38] = _7903_ | _7902_ /*17648*/;
  assign _7904_ = ~q[16] /*17647*/;
  assign _7905_ = sum_16[39] & q[16] /*17646*/;
  assign _7906_ = m_16[39] & _7904_ /*17645*/;
  assign r_16[39] = _7906_ | _7905_ /*17644*/;
  assign _7907_ = ~q[16] /*17643*/;
  assign _7908_ = sum_16[40] & q[16] /*17642*/;
  assign _7909_ = m_16[40] & _7907_ /*17641*/;
  assign r_16[40] = _7909_ | _7908_ /*17640*/;
  assign _7910_ = ~q[16] /*17639*/;
  assign _7911_ = sum_16[41] & q[16] /*17638*/;
  assign _7912_ = m_16[41] & _7910_ /*17637*/;
  assign r_16[41] = _7912_ | _7911_ /*17636*/;
  assign _7913_ = ~q[16] /*17635*/;
  assign _7914_ = sum_16[42] & q[16] /*17634*/;
  assign _7915_ = m_16[42] & _7913_ /*17633*/;
  assign r_16[42] = _7915_ | _7914_ /*17632*/;
  assign _7916_ = ~q[16] /*17631*/;
  assign _7917_ = sum_16[43] & q[16] /*17630*/;
  assign _7918_ = m_16[43] & _7916_ /*17629*/;
  assign r_16[43] = _7918_ | _7917_ /*17628*/;
  assign _7919_ = ~q[16] /*17627*/;
  assign _7920_ = sum_16[44] & q[16] /*17626*/;
  assign _7921_ = m_16[44] & _7919_ /*17625*/;
  assign r_16[44] = _7921_ | _7920_ /*17624*/;
  assign _7922_ = ~q[16] /*17623*/;
  assign _7923_ = sum_16[45] & q[16] /*17622*/;
  assign _7924_ = m_16[45] & _7922_ /*17621*/;
  assign r_16[45] = _7924_ | _7923_ /*17620*/;
  assign _7925_ = ~q[16] /*17619*/;
  assign _7926_ = sum_16[46] & q[16] /*17618*/;
  assign _7927_ = m_16[46] & _7925_ /*17617*/;
  assign r_16[46] = _7927_ | _7926_ /*17616*/;
  assign _7928_ = ~q[16] /*17615*/;
  assign _7929_ = sum_16[47] & q[16] /*17614*/;
  assign _7930_ = m_16[47] & _7928_ /*17613*/;
  assign r_16[47] = _7930_ | _7929_ /*17612*/;
  assign _7931_ = ~q[16] /*17611*/;
  assign _7932_ = sum_16[48] & q[16] /*17610*/;
  assign _7933_ = m_16[48] & _7931_ /*17609*/;
  assign r_16[48] = _7933_ | _7932_ /*17608*/;
  assign _7934_ = ~q[16] /*17607*/;
  assign _7935_ = sum_16[49] & q[16] /*17606*/;
  assign _7936_ = m_16[49] & _7934_ /*17605*/;
  assign r_16[49] = _7936_ | _7935_ /*17604*/;
  assign _7937_ = ~q[16] /*17603*/;
  assign _7938_ = sum_16[50] & q[16] /*17602*/;
  assign _7939_ = m_16[50] & _7937_ /*17601*/;
  assign r_16[50] = _7939_ | _7938_ /*17600*/;
  assign _7940_ = ~q[16] /*17599*/;
  assign _7941_ = sum_16[51] & q[16] /*17598*/;
  assign _7942_ = m_16[51] & _7940_ /*17597*/;
  assign r_16[51] = _7942_ | _7941_ /*17596*/;
  assign _7943_ = ~q[16] /*17595*/;
  assign _7944_ = sum_16[52] & q[16] /*17594*/;
  assign _7945_ = m_16[52] & _7943_ /*17593*/;
  assign r_16[52] = _7945_ | _7944_ /*17592*/;
  assign _7946_ = ~q[16] /*17591*/;
  assign _7947_ = sum_16[53] & q[16] /*17590*/;
  assign _7948_ = m_16[53] & _7946_ /*17589*/;
  assign r_16[53] = _7948_ | _7947_ /*17588*/;
  assign _7949_ = ~q[16] /*17587*/;
  assign _7950_ = sum_16[54] & q[16] /*17586*/;
  assign _7951_ = m_16[54] & _7949_ /*17585*/;
  assign r_16[54] = _7951_ | _7950_ /*17584*/;
  assign _7952_ = ~q[16] /*17583*/;
  assign _7953_ = sum_16[55] & q[16] /*17582*/;
  assign _7954_ = m_16[55] & _7952_ /*17581*/;
  assign r_16[55] = _7954_ | _7953_ /*17580*/;
  assign _7955_ = ~q[16] /*17579*/;
  assign _7956_ = sum_16[56] & q[16] /*17578*/;
  assign _7957_ = m_16[56] & _7955_ /*17577*/;
  assign r_16[56] = _7957_ | _7956_ /*17576*/;
  assign _7958_ = ~q[16] /*17575*/;
  assign _7959_ = sum_16[57] & q[16] /*17574*/;
  assign _7960_ = m_16[57] & _7958_ /*17573*/;
  assign r_16[57] = _7960_ | _7959_ /*17572*/;
  assign _7961_ = ~q[16] /*17571*/;
  assign _7962_ = sum_16[58] & q[16] /*17570*/;
  assign _7963_ = m_16[58] & _7961_ /*17569*/;
  assign r_16[58] = _7963_ | _7962_ /*17568*/;
  assign _7964_ = ~q[16] /*17567*/;
  assign _7965_ = sum_16[59] & q[16] /*17566*/;
  assign _7966_ = m_16[59] & _7964_ /*17565*/;
  assign r_16[59] = _7966_ | _7965_ /*17564*/;
  assign _7967_ = ~q[16] /*17563*/;
  assign _7968_ = sum_16[60] & q[16] /*17562*/;
  assign _7969_ = m_16[60] & _7967_ /*17561*/;
  assign r_16[60] = _7969_ | _7968_ /*17560*/;
  assign _7970_ = ~q[16] /*17559*/;
  assign _7971_ = sum_16[61] & q[16] /*17558*/;
  assign _7972_ = m_16[61] & _7970_ /*17557*/;
  assign r_16[61] = _7972_ | _7971_ /*17556*/;
  assign _7973_ = ~q[16] /*17555*/;
  assign _7974_ = sum_16[62] & q[16] /*17554*/;
  assign _7975_ = m_16[62] & _7973_ /*17553*/;
  assign r_16[62] = _7975_ | _7974_ /*17552*/;
  assign _7976_ = ~q[16] /*17551*/;
  assign _7977_ = sum_16[63] & q[16] /*17550*/;
  assign _7978_ = m_16[63] & _7976_ /*17549*/;
  assign r_16[63] = _7978_ | _7977_ /*17548*/;
  assign _7979_ = ~q[16] /*17547*/;
  assign _7980_ = sum_16[64] & q[16] /*17546*/;
  assign _7981_ = m_16[64] & _7979_ /*17545*/;
  assign r_16[64] = _7981_ | _7980_ /*17544*/;
  assign _7982_ = ~q[16] /*17543*/;
  assign _7983_ = sum_16[65] & q[16] /*17542*/;
  assign _7984_ = m_16[65] & _7982_ /*17541*/;
  assign r_16[65] = _7984_ | _7983_ /*17540*/;
  assign _7985_ = ~q[16] /*17539*/;
  assign _7986_ = sum_16[66] & q[16] /*17538*/;
  assign _7987_ = m_16[66] & _7985_ /*17537*/;
  assign r_16[66] = _7987_ | _7986_ /*17536*/;
  assign _7988_ = ~q[16] /*17535*/;
  assign _7989_ = sum_16[67] & q[16] /*17534*/;
  assign _7990_ = m_16[67] & _7988_ /*17533*/;
  assign r_16[67] = _7990_ | _7989_ /*17532*/;
  assign _7991_ = ~q[16] /*17531*/;
  assign _7992_ = sum_16[68] & q[16] /*17530*/;
  assign _7993_ = m_16[68] & _7991_ /*17529*/;
  assign r_16[68] = _7993_ | _7992_ /*17528*/;
  assign _7994_ = ~q[16] /*17527*/;
  assign _7995_ = sum_16[69] & q[16] /*17526*/;
  assign _7996_ = m_16[69] & _7994_ /*17525*/;
  assign r_16[69] = _7996_ | _7995_ /*17524*/;
  assign _7997_ = ~q[16] /*17523*/;
  assign _7998_ = sum_16[70] & q[16] /*17522*/;
  assign _7999_ = m_16[70] & _7997_ /*17521*/;
  assign r_16[70] = _7999_ | _7998_ /*17520*/;
  assign _8000_ = ~q[16] /*17519*/;
  assign _8001_ = sum_16[71] & q[16] /*17518*/;
  assign _8002_ = m_16[71] & _8000_ /*17517*/;
  assign r_16[71] = _8002_ | _8001_ /*17516*/;
  assign _8003_ = ~q[16] /*17515*/;
  assign _8004_ = sum_16[72] & q[16] /*17514*/;
  assign _8005_ = m_16[72] & _8003_ /*17513*/;
  assign r_16[72] = _8005_ | _8004_ /*17512*/;
  assign _8006_ = ~q[16] /*17511*/;
  assign _8007_ = sum_16[73] & q[16] /*17510*/;
  assign _8008_ = m_16[73] & _8006_ /*17509*/;
  assign r_16[73] = _8008_ | _8007_ /*17508*/;
  assign _8009_ = ~q[16] /*17507*/;
  assign _8010_ = sum_16[74] & q[16] /*17506*/;
  assign _8011_ = m_16[74] & _8009_ /*17505*/;
  assign r_16[74] = _8011_ | _8010_ /*17504*/;
  assign _8012_ = ~q[16] /*17503*/;
  assign _8013_ = sum_16[75] & q[16] /*17502*/;
  assign _8014_ = m_16[75] & _8012_ /*17501*/;
  assign r_16[75] = _8014_ | _8013_ /*17500*/;
  assign _8015_ = ~q[16] /*17499*/;
  assign _8016_ = sum_16[76] & q[16] /*17498*/;
  assign _8017_ = m_16[76] & _8015_ /*17497*/;
  assign r_16[76] = _8017_ | _8016_ /*17496*/;
  assign _8018_ = ~q[16] /*17495*/;
  assign _8019_ = sum_16[77] & q[16] /*17494*/;
  assign _8020_ = m_16[77] & _8018_ /*17493*/;
  assign r_16[77] = _8020_ | _8019_ /*17492*/;
  assign _8021_ = ~q[16] /*17491*/;
  assign _8022_ = sum_16[78] & q[16] /*17490*/;
  assign _8023_ = m_16[78] & _8021_ /*17489*/;
  assign r_16[78] = _8023_ | _8022_ /*17488*/;
  assign inv_17[0] = oneWire /*17280*/;
  assign inv_17[1] = oneWire /*17274*/;
  assign inv_17[2] = oneWire /*17268*/;
  assign inv_17[3] = oneWire /*17262*/;
  assign inv_17[4] = oneWire /*17256*/;
  assign inv_17[5] = oneWire /*17250*/;
  assign inv_17[6] = oneWire /*17244*/;
  assign inv_17[7] = oneWire /*17238*/;
  assign inv_17[8] = oneWire /*17232*/;
  assign inv_17[9] = oneWire /*17226*/;
  assign inv_17[10] = oneWire /*17220*/;
  assign inv_17[11] = oneWire /*17214*/;
  assign inv_17[12] = oneWire /*17208*/;
  assign inv_17[13] = oneWire /*17202*/;
  assign inv_17[14] = oneWire /*17196*/;
  assign inv_17[15] = ~div[0] /*17190*/;
  assign inv_17[16] = ~div[1] /*17184*/;
  assign inv_17[17] = ~div[2] /*17178*/;
  assign inv_17[18] = ~div[3] /*17172*/;
  assign inv_17[19] = ~div[4] /*17166*/;
  assign inv_17[20] = ~div[5] /*17160*/;
  assign inv_17[21] = ~div[6] /*17154*/;
  assign inv_17[22] = ~div[7] /*17148*/;
  assign inv_17[23] = ~div[8] /*17142*/;
  assign inv_17[24] = ~div[9] /*17136*/;
  assign inv_17[25] = ~div[10] /*17130*/;
  assign inv_17[26] = ~div[11] /*17124*/;
  assign inv_17[27] = ~div[12] /*17118*/;
  assign inv_17[28] = ~div[13] /*17112*/;
  assign inv_17[29] = ~div[14] /*17106*/;
  assign inv_17[30] = ~div[15] /*17100*/;
  assign inv_17[31] = ~div[16] /*17094*/;
  assign inv_17[32] = ~div[17] /*17088*/;
  assign inv_17[33] = ~div[18] /*17082*/;
  assign inv_17[34] = ~div[19] /*17076*/;
  assign inv_17[35] = ~div[20] /*17070*/;
  assign inv_17[36] = ~div[21] /*17064*/;
  assign inv_17[37] = ~div[22] /*17058*/;
  assign inv_17[38] = ~div[23] /*17052*/;
  assign inv_17[39] = ~div[24] /*17046*/;
  assign inv_17[40] = ~div[25] /*17040*/;
  assign inv_17[41] = ~div[26] /*17034*/;
  assign inv_17[42] = ~div[27] /*17028*/;
  assign inv_17[43] = ~div[28] /*17022*/;
  assign inv_17[44] = ~div[29] /*17016*/;
  assign inv_17[45] = ~div[30] /*17010*/;
  assign inv_17[46] = oneWire /*17004*/;
  assign inv_17[47] = oneWire /*16998*/;
  assign inv_17[48] = oneWire /*16992*/;
  assign inv_17[49] = oneWire /*16986*/;
  assign inv_17[50] = oneWire /*16980*/;
  assign inv_17[51] = oneWire /*16974*/;
  assign inv_17[52] = oneWire /*16968*/;
  assign inv_17[53] = oneWire /*16962*/;
  assign inv_17[54] = oneWire /*16956*/;
  assign inv_17[55] = oneWire /*16950*/;
  assign inv_17[56] = oneWire /*16944*/;
  assign inv_17[57] = oneWire /*16938*/;
  assign inv_17[58] = oneWire /*16932*/;
  assign inv_17[59] = oneWire /*16926*/;
  assign inv_17[60] = oneWire /*16920*/;
  assign inv_17[61] = oneWire /*16914*/;
  assign inv_17[62] = oneWire /*16908*/;
  assign inv_17[63] = oneWire /*16902*/;
  assign inv_17[64] = oneWire /*16896*/;
  assign inv_17[65] = oneWire /*16890*/;
  assign inv_17[66] = oneWire /*16884*/;
  assign inv_17[67] = oneWire /*16878*/;
  assign inv_17[68] = oneWire /*16872*/;
  assign inv_17[69] = oneWire /*16866*/;
  assign inv_17[70] = oneWire /*16860*/;
  assign inv_17[71] = oneWire /*16854*/;
  assign inv_17[72] = oneWire /*16848*/;
  assign inv_17[73] = oneWire /*16842*/;
  assign inv_17[74] = oneWire /*16836*/;
  assign inv_17[75] = oneWire /*16830*/;
  assign inv_17[76] = oneWire /*16824*/;
  assign inv_17[77] = oneWire /*16818*/;
  assign inv_17[78] = oneWire /*16812*/;
  assign _8024_ = inv_17[0] ^ r_16[0] /*17279*/;
  assign sum_17[0] = _8024_ ^ oneWire /*17278*/;
  assign _8025_ = _8024_ & oneWire /*17277*/;
  assign _8026_ = inv_17[0] & r_16[0] /*17276*/;
  assign _8027_ = _8025_ | _8026_ /*17275*/;
  assign _8028_ = inv_17[1] ^ r_16[1] /*17273*/;
  assign sum_17[1] = _8028_ ^ _8027_ /*17272*/;
  assign _8029_ = _8028_ & _8027_ /*17271*/;
  assign _8030_ = inv_17[1] & r_16[1] /*17270*/;
  assign _8031_ = _8029_ | _8030_ /*17269*/;
  assign _8032_ = inv_17[2] ^ r_16[2] /*17267*/;
  assign sum_17[2] = _8032_ ^ _8031_ /*17266*/;
  assign _8033_ = _8032_ & _8031_ /*17265*/;
  assign _8034_ = inv_17[2] & r_16[2] /*17264*/;
  assign _8035_ = _8033_ | _8034_ /*17263*/;
  assign _8036_ = inv_17[3] ^ r_16[3] /*17261*/;
  assign sum_17[3] = _8036_ ^ _8035_ /*17260*/;
  assign _8037_ = _8036_ & _8035_ /*17259*/;
  assign _8038_ = inv_17[3] & r_16[3] /*17258*/;
  assign _8039_ = _8037_ | _8038_ /*17257*/;
  assign _8040_ = inv_17[4] ^ r_16[4] /*17255*/;
  assign sum_17[4] = _8040_ ^ _8039_ /*17254*/;
  assign _8041_ = _8040_ & _8039_ /*17253*/;
  assign _8042_ = inv_17[4] & r_16[4] /*17252*/;
  assign _8043_ = _8041_ | _8042_ /*17251*/;
  assign _8044_ = inv_17[5] ^ r_16[5] /*17249*/;
  assign sum_17[5] = _8044_ ^ _8043_ /*17248*/;
  assign _8045_ = _8044_ & _8043_ /*17247*/;
  assign _8046_ = inv_17[5] & r_16[5] /*17246*/;
  assign _8047_ = _8045_ | _8046_ /*17245*/;
  assign _8048_ = inv_17[6] ^ r_16[6] /*17243*/;
  assign sum_17[6] = _8048_ ^ _8047_ /*17242*/;
  assign _8049_ = _8048_ & _8047_ /*17241*/;
  assign _8050_ = inv_17[6] & r_16[6] /*17240*/;
  assign _8051_ = _8049_ | _8050_ /*17239*/;
  assign _8052_ = inv_17[7] ^ r_16[7] /*17237*/;
  assign sum_17[7] = _8052_ ^ _8051_ /*17236*/;
  assign _8053_ = _8052_ & _8051_ /*17235*/;
  assign _8054_ = inv_17[7] & r_16[7] /*17234*/;
  assign _8055_ = _8053_ | _8054_ /*17233*/;
  assign _8056_ = inv_17[8] ^ r_16[8] /*17231*/;
  assign sum_17[8] = _8056_ ^ _8055_ /*17230*/;
  assign _8057_ = _8056_ & _8055_ /*17229*/;
  assign _8058_ = inv_17[8] & r_16[8] /*17228*/;
  assign _8059_ = _8057_ | _8058_ /*17227*/;
  assign _8060_ = inv_17[9] ^ r_16[9] /*17225*/;
  assign sum_17[9] = _8060_ ^ _8059_ /*17224*/;
  assign _8061_ = _8060_ & _8059_ /*17223*/;
  assign _8062_ = inv_17[9] & r_16[9] /*17222*/;
  assign _8063_ = _8061_ | _8062_ /*17221*/;
  assign _8064_ = inv_17[10] ^ r_16[10] /*17219*/;
  assign sum_17[10] = _8064_ ^ _8063_ /*17218*/;
  assign _8065_ = _8064_ & _8063_ /*17217*/;
  assign _8066_ = inv_17[10] & r_16[10] /*17216*/;
  assign _8067_ = _8065_ | _8066_ /*17215*/;
  assign _8068_ = inv_17[11] ^ r_16[11] /*17213*/;
  assign sum_17[11] = _8068_ ^ _8067_ /*17212*/;
  assign _8069_ = _8068_ & _8067_ /*17211*/;
  assign _8070_ = inv_17[11] & r_16[11] /*17210*/;
  assign _8071_ = _8069_ | _8070_ /*17209*/;
  assign _8072_ = inv_17[12] ^ r_16[12] /*17207*/;
  assign sum_17[12] = _8072_ ^ _8071_ /*17206*/;
  assign _8073_ = _8072_ & _8071_ /*17205*/;
  assign _8074_ = inv_17[12] & r_16[12] /*17204*/;
  assign _8075_ = _8073_ | _8074_ /*17203*/;
  assign _8076_ = inv_17[13] ^ r_16[13] /*17201*/;
  assign sum_17[13] = _8076_ ^ _8075_ /*17200*/;
  assign _8077_ = _8076_ & _8075_ /*17199*/;
  assign _8078_ = inv_17[13] & r_16[13] /*17198*/;
  assign _8079_ = _8077_ | _8078_ /*17197*/;
  assign _8080_ = inv_17[14] ^ r_16[14] /*17195*/;
  assign sum_17[14] = _8080_ ^ _8079_ /*17194*/;
  assign _8081_ = _8080_ & _8079_ /*17193*/;
  assign _8082_ = inv_17[14] & r_16[14] /*17192*/;
  assign _8083_ = _8081_ | _8082_ /*17191*/;
  assign _8084_ = inv_17[15] ^ r_16[15] /*17189*/;
  assign sum_17[15] = _8084_ ^ _8083_ /*17188*/;
  assign _8085_ = _8084_ & _8083_ /*17187*/;
  assign _8086_ = inv_17[15] & r_16[15] /*17186*/;
  assign _8087_ = _8085_ | _8086_ /*17185*/;
  assign _8088_ = inv_17[16] ^ r_16[16] /*17183*/;
  assign sum_17[16] = _8088_ ^ _8087_ /*17182*/;
  assign _8089_ = _8088_ & _8087_ /*17181*/;
  assign _8090_ = inv_17[16] & r_16[16] /*17180*/;
  assign _8091_ = _8089_ | _8090_ /*17179*/;
  assign _8092_ = inv_17[17] ^ r_16[17] /*17177*/;
  assign sum_17[17] = _8092_ ^ _8091_ /*17176*/;
  assign _8093_ = _8092_ & _8091_ /*17175*/;
  assign _8094_ = inv_17[17] & r_16[17] /*17174*/;
  assign _8095_ = _8093_ | _8094_ /*17173*/;
  assign _8096_ = inv_17[18] ^ r_16[18] /*17171*/;
  assign sum_17[18] = _8096_ ^ _8095_ /*17170*/;
  assign _8097_ = _8096_ & _8095_ /*17169*/;
  assign _8098_ = inv_17[18] & r_16[18] /*17168*/;
  assign _8099_ = _8097_ | _8098_ /*17167*/;
  assign _8100_ = inv_17[19] ^ r_16[19] /*17165*/;
  assign sum_17[19] = _8100_ ^ _8099_ /*17164*/;
  assign _8101_ = _8100_ & _8099_ /*17163*/;
  assign _8102_ = inv_17[19] & r_16[19] /*17162*/;
  assign _8103_ = _8101_ | _8102_ /*17161*/;
  assign _8104_ = inv_17[20] ^ r_16[20] /*17159*/;
  assign sum_17[20] = _8104_ ^ _8103_ /*17158*/;
  assign _8105_ = _8104_ & _8103_ /*17157*/;
  assign _8106_ = inv_17[20] & r_16[20] /*17156*/;
  assign _8107_ = _8105_ | _8106_ /*17155*/;
  assign _8108_ = inv_17[21] ^ r_16[21] /*17153*/;
  assign sum_17[21] = _8108_ ^ _8107_ /*17152*/;
  assign _8109_ = _8108_ & _8107_ /*17151*/;
  assign _8110_ = inv_17[21] & r_16[21] /*17150*/;
  assign _8111_ = _8109_ | _8110_ /*17149*/;
  assign _8112_ = inv_17[22] ^ r_16[22] /*17147*/;
  assign sum_17[22] = _8112_ ^ _8111_ /*17146*/;
  assign _8113_ = _8112_ & _8111_ /*17145*/;
  assign _8114_ = inv_17[22] & r_16[22] /*17144*/;
  assign _8115_ = _8113_ | _8114_ /*17143*/;
  assign _8116_ = inv_17[23] ^ r_16[23] /*17141*/;
  assign sum_17[23] = _8116_ ^ _8115_ /*17140*/;
  assign _8117_ = _8116_ & _8115_ /*17139*/;
  assign _8118_ = inv_17[23] & r_16[23] /*17138*/;
  assign _8119_ = _8117_ | _8118_ /*17137*/;
  assign _8120_ = inv_17[24] ^ r_16[24] /*17135*/;
  assign sum_17[24] = _8120_ ^ _8119_ /*17134*/;
  assign _8121_ = _8120_ & _8119_ /*17133*/;
  assign _8122_ = inv_17[24] & r_16[24] /*17132*/;
  assign _8123_ = _8121_ | _8122_ /*17131*/;
  assign _8124_ = inv_17[25] ^ r_16[25] /*17129*/;
  assign sum_17[25] = _8124_ ^ _8123_ /*17128*/;
  assign _8125_ = _8124_ & _8123_ /*17127*/;
  assign _8126_ = inv_17[25] & r_16[25] /*17126*/;
  assign _8127_ = _8125_ | _8126_ /*17125*/;
  assign _8128_ = inv_17[26] ^ r_16[26] /*17123*/;
  assign sum_17[26] = _8128_ ^ _8127_ /*17122*/;
  assign _8129_ = _8128_ & _8127_ /*17121*/;
  assign _8130_ = inv_17[26] & r_16[26] /*17120*/;
  assign _8131_ = _8129_ | _8130_ /*17119*/;
  assign _8132_ = inv_17[27] ^ r_16[27] /*17117*/;
  assign sum_17[27] = _8132_ ^ _8131_ /*17116*/;
  assign _8133_ = _8132_ & _8131_ /*17115*/;
  assign _8134_ = inv_17[27] & r_16[27] /*17114*/;
  assign _8135_ = _8133_ | _8134_ /*17113*/;
  assign _8136_ = inv_17[28] ^ r_16[28] /*17111*/;
  assign sum_17[28] = _8136_ ^ _8135_ /*17110*/;
  assign _8137_ = _8136_ & _8135_ /*17109*/;
  assign _8138_ = inv_17[28] & r_16[28] /*17108*/;
  assign _8139_ = _8137_ | _8138_ /*17107*/;
  assign _8140_ = inv_17[29] ^ r_16[29] /*17105*/;
  assign sum_17[29] = _8140_ ^ _8139_ /*17104*/;
  assign _8141_ = _8140_ & _8139_ /*17103*/;
  assign _8142_ = inv_17[29] & r_16[29] /*17102*/;
  assign _8143_ = _8141_ | _8142_ /*17101*/;
  assign _8144_ = inv_17[30] ^ r_16[30] /*17099*/;
  assign sum_17[30] = _8144_ ^ _8143_ /*17098*/;
  assign _8145_ = _8144_ & _8143_ /*17097*/;
  assign _8146_ = inv_17[30] & r_16[30] /*17096*/;
  assign _8147_ = _8145_ | _8146_ /*17095*/;
  assign _8148_ = inv_17[31] ^ r_16[31] /*17093*/;
  assign sum_17[31] = _8148_ ^ _8147_ /*17092*/;
  assign _8149_ = _8148_ & _8147_ /*17091*/;
  assign _8150_ = inv_17[31] & r_16[31] /*17090*/;
  assign _8151_ = _8149_ | _8150_ /*17089*/;
  assign _8152_ = inv_17[32] ^ r_16[32] /*17087*/;
  assign sum_17[32] = _8152_ ^ _8151_ /*17086*/;
  assign _8153_ = _8152_ & _8151_ /*17085*/;
  assign _8154_ = inv_17[32] & r_16[32] /*17084*/;
  assign _8155_ = _8153_ | _8154_ /*17083*/;
  assign _8156_ = inv_17[33] ^ r_16[33] /*17081*/;
  assign sum_17[33] = _8156_ ^ _8155_ /*17080*/;
  assign _8157_ = _8156_ & _8155_ /*17079*/;
  assign _8158_ = inv_17[33] & r_16[33] /*17078*/;
  assign _8159_ = _8157_ | _8158_ /*17077*/;
  assign _8160_ = inv_17[34] ^ r_16[34] /*17075*/;
  assign sum_17[34] = _8160_ ^ _8159_ /*17074*/;
  assign _8161_ = _8160_ & _8159_ /*17073*/;
  assign _8162_ = inv_17[34] & r_16[34] /*17072*/;
  assign _8163_ = _8161_ | _8162_ /*17071*/;
  assign _8164_ = inv_17[35] ^ r_16[35] /*17069*/;
  assign sum_17[35] = _8164_ ^ _8163_ /*17068*/;
  assign _8165_ = _8164_ & _8163_ /*17067*/;
  assign _8166_ = inv_17[35] & r_16[35] /*17066*/;
  assign _8167_ = _8165_ | _8166_ /*17065*/;
  assign _8168_ = inv_17[36] ^ r_16[36] /*17063*/;
  assign sum_17[36] = _8168_ ^ _8167_ /*17062*/;
  assign _8169_ = _8168_ & _8167_ /*17061*/;
  assign _8170_ = inv_17[36] & r_16[36] /*17060*/;
  assign _8171_ = _8169_ | _8170_ /*17059*/;
  assign _8172_ = inv_17[37] ^ r_16[37] /*17057*/;
  assign sum_17[37] = _8172_ ^ _8171_ /*17056*/;
  assign _8173_ = _8172_ & _8171_ /*17055*/;
  assign _8174_ = inv_17[37] & r_16[37] /*17054*/;
  assign _8175_ = _8173_ | _8174_ /*17053*/;
  assign _8176_ = inv_17[38] ^ r_16[38] /*17051*/;
  assign sum_17[38] = _8176_ ^ _8175_ /*17050*/;
  assign _8177_ = _8176_ & _8175_ /*17049*/;
  assign _8178_ = inv_17[38] & r_16[38] /*17048*/;
  assign _8179_ = _8177_ | _8178_ /*17047*/;
  assign _8180_ = inv_17[39] ^ r_16[39] /*17045*/;
  assign sum_17[39] = _8180_ ^ _8179_ /*17044*/;
  assign _8181_ = _8180_ & _8179_ /*17043*/;
  assign _8182_ = inv_17[39] & r_16[39] /*17042*/;
  assign _8183_ = _8181_ | _8182_ /*17041*/;
  assign _8184_ = inv_17[40] ^ r_16[40] /*17039*/;
  assign sum_17[40] = _8184_ ^ _8183_ /*17038*/;
  assign _8185_ = _8184_ & _8183_ /*17037*/;
  assign _8186_ = inv_17[40] & r_16[40] /*17036*/;
  assign _8187_ = _8185_ | _8186_ /*17035*/;
  assign _8188_ = inv_17[41] ^ r_16[41] /*17033*/;
  assign sum_17[41] = _8188_ ^ _8187_ /*17032*/;
  assign _8189_ = _8188_ & _8187_ /*17031*/;
  assign _8190_ = inv_17[41] & r_16[41] /*17030*/;
  assign _8191_ = _8189_ | _8190_ /*17029*/;
  assign _8192_ = inv_17[42] ^ r_16[42] /*17027*/;
  assign sum_17[42] = _8192_ ^ _8191_ /*17026*/;
  assign _8193_ = _8192_ & _8191_ /*17025*/;
  assign _8194_ = inv_17[42] & r_16[42] /*17024*/;
  assign _8195_ = _8193_ | _8194_ /*17023*/;
  assign _8196_ = inv_17[43] ^ r_16[43] /*17021*/;
  assign sum_17[43] = _8196_ ^ _8195_ /*17020*/;
  assign _8197_ = _8196_ & _8195_ /*17019*/;
  assign _8198_ = inv_17[43] & r_16[43] /*17018*/;
  assign _8199_ = _8197_ | _8198_ /*17017*/;
  assign _8200_ = inv_17[44] ^ r_16[44] /*17015*/;
  assign sum_17[44] = _8200_ ^ _8199_ /*17014*/;
  assign _8201_ = _8200_ & _8199_ /*17013*/;
  assign _8202_ = inv_17[44] & r_16[44] /*17012*/;
  assign _8203_ = _8201_ | _8202_ /*17011*/;
  assign _8204_ = inv_17[45] ^ r_16[45] /*17009*/;
  assign sum_17[45] = _8204_ ^ _8203_ /*17008*/;
  assign _8205_ = _8204_ & _8203_ /*17007*/;
  assign _8206_ = inv_17[45] & r_16[45] /*17006*/;
  assign _8207_ = _8205_ | _8206_ /*17005*/;
  assign _8208_ = inv_17[46] ^ r_16[46] /*17003*/;
  assign sum_17[46] = _8208_ ^ _8207_ /*17002*/;
  assign _8209_ = _8208_ & _8207_ /*17001*/;
  assign _8210_ = inv_17[46] & r_16[46] /*17000*/;
  assign _8211_ = _8209_ | _8210_ /*16999*/;
  assign _8212_ = inv_17[47] ^ r_16[47] /*16997*/;
  assign sum_17[47] = _8212_ ^ _8211_ /*16996*/;
  assign _8213_ = _8212_ & _8211_ /*16995*/;
  assign _8214_ = inv_17[47] & r_16[47] /*16994*/;
  assign _8215_ = _8213_ | _8214_ /*16993*/;
  assign _8216_ = inv_17[48] ^ r_16[48] /*16991*/;
  assign sum_17[48] = _8216_ ^ _8215_ /*16990*/;
  assign _8217_ = _8216_ & _8215_ /*16989*/;
  assign _8218_ = inv_17[48] & r_16[48] /*16988*/;
  assign _8219_ = _8217_ | _8218_ /*16987*/;
  assign _8220_ = inv_17[49] ^ r_16[49] /*16985*/;
  assign sum_17[49] = _8220_ ^ _8219_ /*16984*/;
  assign _8221_ = _8220_ & _8219_ /*16983*/;
  assign _8222_ = inv_17[49] & r_16[49] /*16982*/;
  assign _8223_ = _8221_ | _8222_ /*16981*/;
  assign _8224_ = inv_17[50] ^ r_16[50] /*16979*/;
  assign sum_17[50] = _8224_ ^ _8223_ /*16978*/;
  assign _8225_ = _8224_ & _8223_ /*16977*/;
  assign _8226_ = inv_17[50] & r_16[50] /*16976*/;
  assign _8227_ = _8225_ | _8226_ /*16975*/;
  assign _8228_ = inv_17[51] ^ r_16[51] /*16973*/;
  assign sum_17[51] = _8228_ ^ _8227_ /*16972*/;
  assign _8229_ = _8228_ & _8227_ /*16971*/;
  assign _8230_ = inv_17[51] & r_16[51] /*16970*/;
  assign _8231_ = _8229_ | _8230_ /*16969*/;
  assign _8232_ = inv_17[52] ^ r_16[52] /*16967*/;
  assign sum_17[52] = _8232_ ^ _8231_ /*16966*/;
  assign _8233_ = _8232_ & _8231_ /*16965*/;
  assign _8234_ = inv_17[52] & r_16[52] /*16964*/;
  assign _8235_ = _8233_ | _8234_ /*16963*/;
  assign _8236_ = inv_17[53] ^ r_16[53] /*16961*/;
  assign sum_17[53] = _8236_ ^ _8235_ /*16960*/;
  assign _8237_ = _8236_ & _8235_ /*16959*/;
  assign _8238_ = inv_17[53] & r_16[53] /*16958*/;
  assign _8239_ = _8237_ | _8238_ /*16957*/;
  assign _8240_ = inv_17[54] ^ r_16[54] /*16955*/;
  assign sum_17[54] = _8240_ ^ _8239_ /*16954*/;
  assign _8241_ = _8240_ & _8239_ /*16953*/;
  assign _8242_ = inv_17[54] & r_16[54] /*16952*/;
  assign _8243_ = _8241_ | _8242_ /*16951*/;
  assign _8244_ = inv_17[55] ^ r_16[55] /*16949*/;
  assign sum_17[55] = _8244_ ^ _8243_ /*16948*/;
  assign _8245_ = _8244_ & _8243_ /*16947*/;
  assign _8246_ = inv_17[55] & r_16[55] /*16946*/;
  assign _8247_ = _8245_ | _8246_ /*16945*/;
  assign _8248_ = inv_17[56] ^ r_16[56] /*16943*/;
  assign sum_17[56] = _8248_ ^ _8247_ /*16942*/;
  assign _8249_ = _8248_ & _8247_ /*16941*/;
  assign _8250_ = inv_17[56] & r_16[56] /*16940*/;
  assign _8251_ = _8249_ | _8250_ /*16939*/;
  assign _8252_ = inv_17[57] ^ r_16[57] /*16937*/;
  assign sum_17[57] = _8252_ ^ _8251_ /*16936*/;
  assign _8253_ = _8252_ & _8251_ /*16935*/;
  assign _8254_ = inv_17[57] & r_16[57] /*16934*/;
  assign _8255_ = _8253_ | _8254_ /*16933*/;
  assign _8256_ = inv_17[58] ^ r_16[58] /*16931*/;
  assign sum_17[58] = _8256_ ^ _8255_ /*16930*/;
  assign _8257_ = _8256_ & _8255_ /*16929*/;
  assign _8258_ = inv_17[58] & r_16[58] /*16928*/;
  assign _8259_ = _8257_ | _8258_ /*16927*/;
  assign _8260_ = inv_17[59] ^ r_16[59] /*16925*/;
  assign sum_17[59] = _8260_ ^ _8259_ /*16924*/;
  assign _8261_ = _8260_ & _8259_ /*16923*/;
  assign _8262_ = inv_17[59] & r_16[59] /*16922*/;
  assign _8263_ = _8261_ | _8262_ /*16921*/;
  assign _8264_ = inv_17[60] ^ r_16[60] /*16919*/;
  assign sum_17[60] = _8264_ ^ _8263_ /*16918*/;
  assign _8265_ = _8264_ & _8263_ /*16917*/;
  assign _8266_ = inv_17[60] & r_16[60] /*16916*/;
  assign _8267_ = _8265_ | _8266_ /*16915*/;
  assign _8268_ = inv_17[61] ^ r_16[61] /*16913*/;
  assign sum_17[61] = _8268_ ^ _8267_ /*16912*/;
  assign _8269_ = _8268_ & _8267_ /*16911*/;
  assign _8270_ = inv_17[61] & r_16[61] /*16910*/;
  assign _8271_ = _8269_ | _8270_ /*16909*/;
  assign _8272_ = inv_17[62] ^ r_16[62] /*16907*/;
  assign sum_17[62] = _8272_ ^ _8271_ /*16906*/;
  assign _8273_ = _8272_ & _8271_ /*16905*/;
  assign _8274_ = inv_17[62] & r_16[62] /*16904*/;
  assign _8275_ = _8273_ | _8274_ /*16903*/;
  assign _8276_ = inv_17[63] ^ r_16[63] /*16901*/;
  assign sum_17[63] = _8276_ ^ _8275_ /*16900*/;
  assign _8277_ = _8276_ & _8275_ /*16899*/;
  assign _8278_ = inv_17[63] & r_16[63] /*16898*/;
  assign _8279_ = _8277_ | _8278_ /*16897*/;
  assign _8280_ = inv_17[64] ^ r_16[64] /*16895*/;
  assign sum_17[64] = _8280_ ^ _8279_ /*16894*/;
  assign _8281_ = _8280_ & _8279_ /*16893*/;
  assign _8282_ = inv_17[64] & r_16[64] /*16892*/;
  assign _8283_ = _8281_ | _8282_ /*16891*/;
  assign _8284_ = inv_17[65] ^ r_16[65] /*16889*/;
  assign sum_17[65] = _8284_ ^ _8283_ /*16888*/;
  assign _8285_ = _8284_ & _8283_ /*16887*/;
  assign _8286_ = inv_17[65] & r_16[65] /*16886*/;
  assign _8287_ = _8285_ | _8286_ /*16885*/;
  assign _8288_ = inv_17[66] ^ r_16[66] /*16883*/;
  assign sum_17[66] = _8288_ ^ _8287_ /*16882*/;
  assign _8289_ = _8288_ & _8287_ /*16881*/;
  assign _8290_ = inv_17[66] & r_16[66] /*16880*/;
  assign _8291_ = _8289_ | _8290_ /*16879*/;
  assign _8292_ = inv_17[67] ^ r_16[67] /*16877*/;
  assign sum_17[67] = _8292_ ^ _8291_ /*16876*/;
  assign _8293_ = _8292_ & _8291_ /*16875*/;
  assign _8294_ = inv_17[67] & r_16[67] /*16874*/;
  assign _8295_ = _8293_ | _8294_ /*16873*/;
  assign _8296_ = inv_17[68] ^ r_16[68] /*16871*/;
  assign sum_17[68] = _8296_ ^ _8295_ /*16870*/;
  assign _8297_ = _8296_ & _8295_ /*16869*/;
  assign _8298_ = inv_17[68] & r_16[68] /*16868*/;
  assign _8299_ = _8297_ | _8298_ /*16867*/;
  assign _8300_ = inv_17[69] ^ r_16[69] /*16865*/;
  assign sum_17[69] = _8300_ ^ _8299_ /*16864*/;
  assign _8301_ = _8300_ & _8299_ /*16863*/;
  assign _8302_ = inv_17[69] & r_16[69] /*16862*/;
  assign _8303_ = _8301_ | _8302_ /*16861*/;
  assign _8304_ = inv_17[70] ^ r_16[70] /*16859*/;
  assign sum_17[70] = _8304_ ^ _8303_ /*16858*/;
  assign _8305_ = _8304_ & _8303_ /*16857*/;
  assign _8306_ = inv_17[70] & r_16[70] /*16856*/;
  assign _8307_ = _8305_ | _8306_ /*16855*/;
  assign _8308_ = inv_17[71] ^ r_16[71] /*16853*/;
  assign sum_17[71] = _8308_ ^ _8307_ /*16852*/;
  assign _8309_ = _8308_ & _8307_ /*16851*/;
  assign _8310_ = inv_17[71] & r_16[71] /*16850*/;
  assign _8311_ = _8309_ | _8310_ /*16849*/;
  assign _8312_ = inv_17[72] ^ r_16[72] /*16847*/;
  assign sum_17[72] = _8312_ ^ _8311_ /*16846*/;
  assign _8313_ = _8312_ & _8311_ /*16845*/;
  assign _8314_ = inv_17[72] & r_16[72] /*16844*/;
  assign _8315_ = _8313_ | _8314_ /*16843*/;
  assign _8316_ = inv_17[73] ^ r_16[73] /*16841*/;
  assign sum_17[73] = _8316_ ^ _8315_ /*16840*/;
  assign _8317_ = _8316_ & _8315_ /*16839*/;
  assign _8318_ = inv_17[73] & r_16[73] /*16838*/;
  assign _8319_ = _8317_ | _8318_ /*16837*/;
  assign _8320_ = inv_17[74] ^ r_16[74] /*16835*/;
  assign sum_17[74] = _8320_ ^ _8319_ /*16834*/;
  assign _8321_ = _8320_ & _8319_ /*16833*/;
  assign _8322_ = inv_17[74] & r_16[74] /*16832*/;
  assign _8323_ = _8321_ | _8322_ /*16831*/;
  assign _8324_ = inv_17[75] ^ r_16[75] /*16829*/;
  assign sum_17[75] = _8324_ ^ _8323_ /*16828*/;
  assign _8325_ = _8324_ & _8323_ /*16827*/;
  assign _8326_ = inv_17[75] & r_16[75] /*16826*/;
  assign _8327_ = _8325_ | _8326_ /*16825*/;
  assign _8328_ = inv_17[76] ^ r_16[76] /*16823*/;
  assign sum_17[76] = _8328_ ^ _8327_ /*16822*/;
  assign _8329_ = _8328_ & _8327_ /*16821*/;
  assign _8330_ = inv_17[76] & r_16[76] /*16820*/;
  assign _8331_ = _8329_ | _8330_ /*16819*/;
  assign _8332_ = inv_17[77] ^ r_16[77] /*16817*/;
  assign sum_17[77] = _8332_ ^ _8331_ /*16816*/;
  assign _8333_ = _8332_ & _8331_ /*16815*/;
  assign _8334_ = inv_17[77] & r_16[77] /*16814*/;
  assign _8335_ = _8333_ | _8334_ /*16813*/;
  assign _8336_ = inv_17[78] ^ r_16[78] /*16811*/;
  assign sum_17[78] = _8336_ ^ _8335_ /*16810*/;
  assign _8337_ = _8336_ & _8335_ /*16809*/;
  assign _8338_ = inv_17[78] & r_16[78] /*16808*/;
  assign _8339_ = _8337_ | _8338_ /*16807*/;
  assign _8340_ = _8339_ ^ _8335_ /*16806*/;
  assign _8341_ = ~_8340_ /*16805*/;
  assign _8342_ = sum_17[78] & _8341_ /*16804*/;
  assign _8343_ = _8340_ & _8339_ /*16803*/;
  assign sum_17[79] = _8343_ | _8342_ /*16802*/;
  assign q[15] = ~sum_17[79] /*16801*/;
  assign m_17[0] = r_16[0] /*16800*/;
  assign m_17[1] = r_16[1] /*16799*/;
  assign m_17[2] = r_16[2] /*16798*/;
  assign m_17[3] = r_16[3] /*16797*/;
  assign m_17[4] = r_16[4] /*16796*/;
  assign m_17[5] = r_16[5] /*16795*/;
  assign m_17[6] = r_16[6] /*16794*/;
  assign m_17[7] = r_16[7] /*16793*/;
  assign m_17[8] = r_16[8] /*16792*/;
  assign m_17[9] = r_16[9] /*16791*/;
  assign m_17[10] = r_16[10] /*16790*/;
  assign m_17[11] = r_16[11] /*16789*/;
  assign m_17[12] = r_16[12] /*16788*/;
  assign m_17[13] = r_16[13] /*16787*/;
  assign m_17[14] = r_16[14] /*16786*/;
  assign m_17[15] = r_16[15] /*16785*/;
  assign m_17[16] = r_16[16] /*16784*/;
  assign m_17[17] = r_16[17] /*16783*/;
  assign m_17[18] = r_16[18] /*16782*/;
  assign m_17[19] = r_16[19] /*16781*/;
  assign m_17[20] = r_16[20] /*16780*/;
  assign m_17[21] = r_16[21] /*16779*/;
  assign m_17[22] = r_16[22] /*16778*/;
  assign m_17[23] = r_16[23] /*16777*/;
  assign m_17[24] = r_16[24] /*16776*/;
  assign m_17[25] = r_16[25] /*16775*/;
  assign m_17[26] = r_16[26] /*16774*/;
  assign m_17[27] = r_16[27] /*16773*/;
  assign m_17[28] = r_16[28] /*16772*/;
  assign m_17[29] = r_16[29] /*16771*/;
  assign m_17[30] = r_16[30] /*16770*/;
  assign m_17[31] = r_16[31] /*16769*/;
  assign m_17[32] = r_16[32] /*16768*/;
  assign m_17[33] = r_16[33] /*16767*/;
  assign m_17[34] = r_16[34] /*16766*/;
  assign m_17[35] = r_16[35] /*16765*/;
  assign m_17[36] = r_16[36] /*16764*/;
  assign m_17[37] = r_16[37] /*16763*/;
  assign m_17[38] = r_16[38] /*16762*/;
  assign m_17[39] = r_16[39] /*16761*/;
  assign m_17[40] = r_16[40] /*16760*/;
  assign m_17[41] = r_16[41] /*16759*/;
  assign m_17[42] = r_16[42] /*16758*/;
  assign m_17[43] = r_16[43] /*16757*/;
  assign m_17[44] = r_16[44] /*16756*/;
  assign m_17[45] = r_16[45] /*16755*/;
  assign m_17[46] = r_16[46] /*16754*/;
  assign m_17[47] = r_16[47] /*16753*/;
  assign m_17[48] = r_16[48] /*16752*/;
  assign m_17[49] = r_16[49] /*16751*/;
  assign m_17[50] = r_16[50] /*16750*/;
  assign m_17[51] = r_16[51] /*16749*/;
  assign m_17[52] = r_16[52] /*16748*/;
  assign m_17[53] = r_16[53] /*16747*/;
  assign m_17[54] = r_16[54] /*16746*/;
  assign m_17[55] = r_16[55] /*16745*/;
  assign m_17[56] = r_16[56] /*16744*/;
  assign m_17[57] = r_16[57] /*16743*/;
  assign m_17[58] = r_16[58] /*16742*/;
  assign m_17[59] = r_16[59] /*16741*/;
  assign m_17[60] = r_16[60] /*16740*/;
  assign m_17[61] = r_16[61] /*16739*/;
  assign m_17[62] = r_16[62] /*16738*/;
  assign m_17[63] = r_16[63] /*16737*/;
  assign m_17[64] = r_16[64] /*16736*/;
  assign m_17[65] = r_16[65] /*16735*/;
  assign m_17[66] = r_16[66] /*16734*/;
  assign m_17[67] = r_16[67] /*16733*/;
  assign m_17[68] = r_16[68] /*16732*/;
  assign m_17[69] = r_16[69] /*16731*/;
  assign m_17[70] = r_16[70] /*16730*/;
  assign m_17[71] = r_16[71] /*16729*/;
  assign m_17[72] = r_16[72] /*16728*/;
  assign m_17[73] = r_16[73] /*16727*/;
  assign m_17[74] = r_16[74] /*16726*/;
  assign m_17[75] = r_16[75] /*16725*/;
  assign m_17[76] = r_16[76] /*16724*/;
  assign m_17[77] = r_16[77] /*16723*/;
  assign m_17[78] = r_16[78] /*16722*/;
  assign m_17[79] = r_16[78] /*16721*/;
  assign _8345_ = ~q[15] /*16720*/;
  assign _8346_ = sum_17[0] & q[15] /*16719*/;
  assign _8347_ = m_17[0] & _8345_ /*16718*/;
  assign r_17[0] = _8347_ | _8346_ /*16717*/;
  assign _8348_ = ~q[15] /*16716*/;
  assign _8349_ = sum_17[1] & q[15] /*16715*/;
  assign _8350_ = m_17[1] & _8348_ /*16714*/;
  assign r_17[1] = _8350_ | _8349_ /*16713*/;
  assign _8351_ = ~q[15] /*16712*/;
  assign _8352_ = sum_17[2] & q[15] /*16711*/;
  assign _8353_ = m_17[2] & _8351_ /*16710*/;
  assign r_17[2] = _8353_ | _8352_ /*16709*/;
  assign _8354_ = ~q[15] /*16708*/;
  assign _8355_ = sum_17[3] & q[15] /*16707*/;
  assign _8356_ = m_17[3] & _8354_ /*16706*/;
  assign r_17[3] = _8356_ | _8355_ /*16705*/;
  assign _8357_ = ~q[15] /*16704*/;
  assign _8358_ = sum_17[4] & q[15] /*16703*/;
  assign _8359_ = m_17[4] & _8357_ /*16702*/;
  assign r_17[4] = _8359_ | _8358_ /*16701*/;
  assign _8360_ = ~q[15] /*16700*/;
  assign _8361_ = sum_17[5] & q[15] /*16699*/;
  assign _8362_ = m_17[5] & _8360_ /*16698*/;
  assign r_17[5] = _8362_ | _8361_ /*16697*/;
  assign _8363_ = ~q[15] /*16696*/;
  assign _8364_ = sum_17[6] & q[15] /*16695*/;
  assign _8365_ = m_17[6] & _8363_ /*16694*/;
  assign r_17[6] = _8365_ | _8364_ /*16693*/;
  assign _8366_ = ~q[15] /*16692*/;
  assign _8367_ = sum_17[7] & q[15] /*16691*/;
  assign _8368_ = m_17[7] & _8366_ /*16690*/;
  assign r_17[7] = _8368_ | _8367_ /*16689*/;
  assign _8369_ = ~q[15] /*16688*/;
  assign _8370_ = sum_17[8] & q[15] /*16687*/;
  assign _8371_ = m_17[8] & _8369_ /*16686*/;
  assign r_17[8] = _8371_ | _8370_ /*16685*/;
  assign _8372_ = ~q[15] /*16684*/;
  assign _8373_ = sum_17[9] & q[15] /*16683*/;
  assign _8374_ = m_17[9] & _8372_ /*16682*/;
  assign r_17[9] = _8374_ | _8373_ /*16681*/;
  assign _8375_ = ~q[15] /*16680*/;
  assign _8376_ = sum_17[10] & q[15] /*16679*/;
  assign _8377_ = m_17[10] & _8375_ /*16678*/;
  assign r_17[10] = _8377_ | _8376_ /*16677*/;
  assign _8378_ = ~q[15] /*16676*/;
  assign _8379_ = sum_17[11] & q[15] /*16675*/;
  assign _8380_ = m_17[11] & _8378_ /*16674*/;
  assign r_17[11] = _8380_ | _8379_ /*16673*/;
  assign _8381_ = ~q[15] /*16672*/;
  assign _8382_ = sum_17[12] & q[15] /*16671*/;
  assign _8383_ = m_17[12] & _8381_ /*16670*/;
  assign r_17[12] = _8383_ | _8382_ /*16669*/;
  assign _8384_ = ~q[15] /*16668*/;
  assign _8385_ = sum_17[13] & q[15] /*16667*/;
  assign _8386_ = m_17[13] & _8384_ /*16666*/;
  assign r_17[13] = _8386_ | _8385_ /*16665*/;
  assign _8387_ = ~q[15] /*16664*/;
  assign _8388_ = sum_17[14] & q[15] /*16663*/;
  assign _8389_ = m_17[14] & _8387_ /*16662*/;
  assign r_17[14] = _8389_ | _8388_ /*16661*/;
  assign _8390_ = ~q[15] /*16660*/;
  assign _8391_ = sum_17[15] & q[15] /*16659*/;
  assign _8392_ = m_17[15] & _8390_ /*16658*/;
  assign r_17[15] = _8392_ | _8391_ /*16657*/;
  assign _8393_ = ~q[15] /*16656*/;
  assign _8394_ = sum_17[16] & q[15] /*16655*/;
  assign _8395_ = m_17[16] & _8393_ /*16654*/;
  assign r_17[16] = _8395_ | _8394_ /*16653*/;
  assign _8396_ = ~q[15] /*16652*/;
  assign _8397_ = sum_17[17] & q[15] /*16651*/;
  assign _8398_ = m_17[17] & _8396_ /*16650*/;
  assign r_17[17] = _8398_ | _8397_ /*16649*/;
  assign _8399_ = ~q[15] /*16648*/;
  assign _8400_ = sum_17[18] & q[15] /*16647*/;
  assign _8401_ = m_17[18] & _8399_ /*16646*/;
  assign r_17[18] = _8401_ | _8400_ /*16645*/;
  assign _8402_ = ~q[15] /*16644*/;
  assign _8403_ = sum_17[19] & q[15] /*16643*/;
  assign _8404_ = m_17[19] & _8402_ /*16642*/;
  assign r_17[19] = _8404_ | _8403_ /*16641*/;
  assign _8405_ = ~q[15] /*16640*/;
  assign _8406_ = sum_17[20] & q[15] /*16639*/;
  assign _8407_ = m_17[20] & _8405_ /*16638*/;
  assign r_17[20] = _8407_ | _8406_ /*16637*/;
  assign _8408_ = ~q[15] /*16636*/;
  assign _8409_ = sum_17[21] & q[15] /*16635*/;
  assign _8410_ = m_17[21] & _8408_ /*16634*/;
  assign r_17[21] = _8410_ | _8409_ /*16633*/;
  assign _8411_ = ~q[15] /*16632*/;
  assign _8412_ = sum_17[22] & q[15] /*16631*/;
  assign _8413_ = m_17[22] & _8411_ /*16630*/;
  assign r_17[22] = _8413_ | _8412_ /*16629*/;
  assign _8414_ = ~q[15] /*16628*/;
  assign _8415_ = sum_17[23] & q[15] /*16627*/;
  assign _8416_ = m_17[23] & _8414_ /*16626*/;
  assign r_17[23] = _8416_ | _8415_ /*16625*/;
  assign _8417_ = ~q[15] /*16624*/;
  assign _8418_ = sum_17[24] & q[15] /*16623*/;
  assign _8419_ = m_17[24] & _8417_ /*16622*/;
  assign r_17[24] = _8419_ | _8418_ /*16621*/;
  assign _8420_ = ~q[15] /*16620*/;
  assign _8421_ = sum_17[25] & q[15] /*16619*/;
  assign _8422_ = m_17[25] & _8420_ /*16618*/;
  assign r_17[25] = _8422_ | _8421_ /*16617*/;
  assign _8423_ = ~q[15] /*16616*/;
  assign _8424_ = sum_17[26] & q[15] /*16615*/;
  assign _8425_ = m_17[26] & _8423_ /*16614*/;
  assign r_17[26] = _8425_ | _8424_ /*16613*/;
  assign _8426_ = ~q[15] /*16612*/;
  assign _8427_ = sum_17[27] & q[15] /*16611*/;
  assign _8428_ = m_17[27] & _8426_ /*16610*/;
  assign r_17[27] = _8428_ | _8427_ /*16609*/;
  assign _8429_ = ~q[15] /*16608*/;
  assign _8430_ = sum_17[28] & q[15] /*16607*/;
  assign _8431_ = m_17[28] & _8429_ /*16606*/;
  assign r_17[28] = _8431_ | _8430_ /*16605*/;
  assign _8432_ = ~q[15] /*16604*/;
  assign _8433_ = sum_17[29] & q[15] /*16603*/;
  assign _8434_ = m_17[29] & _8432_ /*16602*/;
  assign r_17[29] = _8434_ | _8433_ /*16601*/;
  assign _8435_ = ~q[15] /*16600*/;
  assign _8436_ = sum_17[30] & q[15] /*16599*/;
  assign _8437_ = m_17[30] & _8435_ /*16598*/;
  assign r_17[30] = _8437_ | _8436_ /*16597*/;
  assign _8438_ = ~q[15] /*16596*/;
  assign _8439_ = sum_17[31] & q[15] /*16595*/;
  assign _8440_ = m_17[31] & _8438_ /*16594*/;
  assign r_17[31] = _8440_ | _8439_ /*16593*/;
  assign _8441_ = ~q[15] /*16592*/;
  assign _8442_ = sum_17[32] & q[15] /*16591*/;
  assign _8443_ = m_17[32] & _8441_ /*16590*/;
  assign r_17[32] = _8443_ | _8442_ /*16589*/;
  assign _8444_ = ~q[15] /*16588*/;
  assign _8445_ = sum_17[33] & q[15] /*16587*/;
  assign _8446_ = m_17[33] & _8444_ /*16586*/;
  assign r_17[33] = _8446_ | _8445_ /*16585*/;
  assign _8447_ = ~q[15] /*16584*/;
  assign _8448_ = sum_17[34] & q[15] /*16583*/;
  assign _8449_ = m_17[34] & _8447_ /*16582*/;
  assign r_17[34] = _8449_ | _8448_ /*16581*/;
  assign _8450_ = ~q[15] /*16580*/;
  assign _8451_ = sum_17[35] & q[15] /*16579*/;
  assign _8452_ = m_17[35] & _8450_ /*16578*/;
  assign r_17[35] = _8452_ | _8451_ /*16577*/;
  assign _8453_ = ~q[15] /*16576*/;
  assign _8454_ = sum_17[36] & q[15] /*16575*/;
  assign _8455_ = m_17[36] & _8453_ /*16574*/;
  assign r_17[36] = _8455_ | _8454_ /*16573*/;
  assign _8456_ = ~q[15] /*16572*/;
  assign _8457_ = sum_17[37] & q[15] /*16571*/;
  assign _8458_ = m_17[37] & _8456_ /*16570*/;
  assign r_17[37] = _8458_ | _8457_ /*16569*/;
  assign _8459_ = ~q[15] /*16568*/;
  assign _8460_ = sum_17[38] & q[15] /*16567*/;
  assign _8461_ = m_17[38] & _8459_ /*16566*/;
  assign r_17[38] = _8461_ | _8460_ /*16565*/;
  assign _8462_ = ~q[15] /*16564*/;
  assign _8463_ = sum_17[39] & q[15] /*16563*/;
  assign _8464_ = m_17[39] & _8462_ /*16562*/;
  assign r_17[39] = _8464_ | _8463_ /*16561*/;
  assign _8465_ = ~q[15] /*16560*/;
  assign _8466_ = sum_17[40] & q[15] /*16559*/;
  assign _8467_ = m_17[40] & _8465_ /*16558*/;
  assign r_17[40] = _8467_ | _8466_ /*16557*/;
  assign _8468_ = ~q[15] /*16556*/;
  assign _8469_ = sum_17[41] & q[15] /*16555*/;
  assign _8470_ = m_17[41] & _8468_ /*16554*/;
  assign r_17[41] = _8470_ | _8469_ /*16553*/;
  assign _8471_ = ~q[15] /*16552*/;
  assign _8472_ = sum_17[42] & q[15] /*16551*/;
  assign _8473_ = m_17[42] & _8471_ /*16550*/;
  assign r_17[42] = _8473_ | _8472_ /*16549*/;
  assign _8474_ = ~q[15] /*16548*/;
  assign _8475_ = sum_17[43] & q[15] /*16547*/;
  assign _8476_ = m_17[43] & _8474_ /*16546*/;
  assign r_17[43] = _8476_ | _8475_ /*16545*/;
  assign _8477_ = ~q[15] /*16544*/;
  assign _8478_ = sum_17[44] & q[15] /*16543*/;
  assign _8479_ = m_17[44] & _8477_ /*16542*/;
  assign r_17[44] = _8479_ | _8478_ /*16541*/;
  assign _8480_ = ~q[15] /*16540*/;
  assign _8481_ = sum_17[45] & q[15] /*16539*/;
  assign _8482_ = m_17[45] & _8480_ /*16538*/;
  assign r_17[45] = _8482_ | _8481_ /*16537*/;
  assign _8483_ = ~q[15] /*16536*/;
  assign _8484_ = sum_17[46] & q[15] /*16535*/;
  assign _8485_ = m_17[46] & _8483_ /*16534*/;
  assign r_17[46] = _8485_ | _8484_ /*16533*/;
  assign _8486_ = ~q[15] /*16532*/;
  assign _8487_ = sum_17[47] & q[15] /*16531*/;
  assign _8488_ = m_17[47] & _8486_ /*16530*/;
  assign r_17[47] = _8488_ | _8487_ /*16529*/;
  assign _8489_ = ~q[15] /*16528*/;
  assign _8490_ = sum_17[48] & q[15] /*16527*/;
  assign _8491_ = m_17[48] & _8489_ /*16526*/;
  assign r_17[48] = _8491_ | _8490_ /*16525*/;
  assign _8492_ = ~q[15] /*16524*/;
  assign _8493_ = sum_17[49] & q[15] /*16523*/;
  assign _8494_ = m_17[49] & _8492_ /*16522*/;
  assign r_17[49] = _8494_ | _8493_ /*16521*/;
  assign _8495_ = ~q[15] /*16520*/;
  assign _8496_ = sum_17[50] & q[15] /*16519*/;
  assign _8497_ = m_17[50] & _8495_ /*16518*/;
  assign r_17[50] = _8497_ | _8496_ /*16517*/;
  assign _8498_ = ~q[15] /*16516*/;
  assign _8499_ = sum_17[51] & q[15] /*16515*/;
  assign _8500_ = m_17[51] & _8498_ /*16514*/;
  assign r_17[51] = _8500_ | _8499_ /*16513*/;
  assign _8501_ = ~q[15] /*16512*/;
  assign _8502_ = sum_17[52] & q[15] /*16511*/;
  assign _8503_ = m_17[52] & _8501_ /*16510*/;
  assign r_17[52] = _8503_ | _8502_ /*16509*/;
  assign _8504_ = ~q[15] /*16508*/;
  assign _8505_ = sum_17[53] & q[15] /*16507*/;
  assign _8506_ = m_17[53] & _8504_ /*16506*/;
  assign r_17[53] = _8506_ | _8505_ /*16505*/;
  assign _8507_ = ~q[15] /*16504*/;
  assign _8508_ = sum_17[54] & q[15] /*16503*/;
  assign _8509_ = m_17[54] & _8507_ /*16502*/;
  assign r_17[54] = _8509_ | _8508_ /*16501*/;
  assign _8510_ = ~q[15] /*16500*/;
  assign _8511_ = sum_17[55] & q[15] /*16499*/;
  assign _8512_ = m_17[55] & _8510_ /*16498*/;
  assign r_17[55] = _8512_ | _8511_ /*16497*/;
  assign _8513_ = ~q[15] /*16496*/;
  assign _8514_ = sum_17[56] & q[15] /*16495*/;
  assign _8515_ = m_17[56] & _8513_ /*16494*/;
  assign r_17[56] = _8515_ | _8514_ /*16493*/;
  assign _8516_ = ~q[15] /*16492*/;
  assign _8517_ = sum_17[57] & q[15] /*16491*/;
  assign _8518_ = m_17[57] & _8516_ /*16490*/;
  assign r_17[57] = _8518_ | _8517_ /*16489*/;
  assign _8519_ = ~q[15] /*16488*/;
  assign _8520_ = sum_17[58] & q[15] /*16487*/;
  assign _8521_ = m_17[58] & _8519_ /*16486*/;
  assign r_17[58] = _8521_ | _8520_ /*16485*/;
  assign _8522_ = ~q[15] /*16484*/;
  assign _8523_ = sum_17[59] & q[15] /*16483*/;
  assign _8524_ = m_17[59] & _8522_ /*16482*/;
  assign r_17[59] = _8524_ | _8523_ /*16481*/;
  assign _8525_ = ~q[15] /*16480*/;
  assign _8526_ = sum_17[60] & q[15] /*16479*/;
  assign _8527_ = m_17[60] & _8525_ /*16478*/;
  assign r_17[60] = _8527_ | _8526_ /*16477*/;
  assign _8528_ = ~q[15] /*16476*/;
  assign _8529_ = sum_17[61] & q[15] /*16475*/;
  assign _8530_ = m_17[61] & _8528_ /*16474*/;
  assign r_17[61] = _8530_ | _8529_ /*16473*/;
  assign _8531_ = ~q[15] /*16472*/;
  assign _8532_ = sum_17[62] & q[15] /*16471*/;
  assign _8533_ = m_17[62] & _8531_ /*16470*/;
  assign r_17[62] = _8533_ | _8532_ /*16469*/;
  assign _8534_ = ~q[15] /*16468*/;
  assign _8535_ = sum_17[63] & q[15] /*16467*/;
  assign _8536_ = m_17[63] & _8534_ /*16466*/;
  assign r_17[63] = _8536_ | _8535_ /*16465*/;
  assign _8537_ = ~q[15] /*16464*/;
  assign _8538_ = sum_17[64] & q[15] /*16463*/;
  assign _8539_ = m_17[64] & _8537_ /*16462*/;
  assign r_17[64] = _8539_ | _8538_ /*16461*/;
  assign _8540_ = ~q[15] /*16460*/;
  assign _8541_ = sum_17[65] & q[15] /*16459*/;
  assign _8542_ = m_17[65] & _8540_ /*16458*/;
  assign r_17[65] = _8542_ | _8541_ /*16457*/;
  assign _8543_ = ~q[15] /*16456*/;
  assign _8544_ = sum_17[66] & q[15] /*16455*/;
  assign _8545_ = m_17[66] & _8543_ /*16454*/;
  assign r_17[66] = _8545_ | _8544_ /*16453*/;
  assign _8546_ = ~q[15] /*16452*/;
  assign _8547_ = sum_17[67] & q[15] /*16451*/;
  assign _8548_ = m_17[67] & _8546_ /*16450*/;
  assign r_17[67] = _8548_ | _8547_ /*16449*/;
  assign _8549_ = ~q[15] /*16448*/;
  assign _8550_ = sum_17[68] & q[15] /*16447*/;
  assign _8551_ = m_17[68] & _8549_ /*16446*/;
  assign r_17[68] = _8551_ | _8550_ /*16445*/;
  assign _8552_ = ~q[15] /*16444*/;
  assign _8553_ = sum_17[69] & q[15] /*16443*/;
  assign _8554_ = m_17[69] & _8552_ /*16442*/;
  assign r_17[69] = _8554_ | _8553_ /*16441*/;
  assign _8555_ = ~q[15] /*16440*/;
  assign _8556_ = sum_17[70] & q[15] /*16439*/;
  assign _8557_ = m_17[70] & _8555_ /*16438*/;
  assign r_17[70] = _8557_ | _8556_ /*16437*/;
  assign _8558_ = ~q[15] /*16436*/;
  assign _8559_ = sum_17[71] & q[15] /*16435*/;
  assign _8560_ = m_17[71] & _8558_ /*16434*/;
  assign r_17[71] = _8560_ | _8559_ /*16433*/;
  assign _8561_ = ~q[15] /*16432*/;
  assign _8562_ = sum_17[72] & q[15] /*16431*/;
  assign _8563_ = m_17[72] & _8561_ /*16430*/;
  assign r_17[72] = _8563_ | _8562_ /*16429*/;
  assign _8564_ = ~q[15] /*16428*/;
  assign _8565_ = sum_17[73] & q[15] /*16427*/;
  assign _8566_ = m_17[73] & _8564_ /*16426*/;
  assign r_17[73] = _8566_ | _8565_ /*16425*/;
  assign _8567_ = ~q[15] /*16424*/;
  assign _8568_ = sum_17[74] & q[15] /*16423*/;
  assign _8569_ = m_17[74] & _8567_ /*16422*/;
  assign r_17[74] = _8569_ | _8568_ /*16421*/;
  assign _8570_ = ~q[15] /*16420*/;
  assign _8571_ = sum_17[75] & q[15] /*16419*/;
  assign _8572_ = m_17[75] & _8570_ /*16418*/;
  assign r_17[75] = _8572_ | _8571_ /*16417*/;
  assign _8573_ = ~q[15] /*16416*/;
  assign _8574_ = sum_17[76] & q[15] /*16415*/;
  assign _8575_ = m_17[76] & _8573_ /*16414*/;
  assign r_17[76] = _8575_ | _8574_ /*16413*/;
  assign _8576_ = ~q[15] /*16412*/;
  assign _8577_ = sum_17[77] & q[15] /*16411*/;
  assign _8578_ = m_17[77] & _8576_ /*16410*/;
  assign r_17[77] = _8578_ | _8577_ /*16409*/;
  assign _8579_ = ~q[15] /*16408*/;
  assign _8580_ = sum_17[78] & q[15] /*16407*/;
  assign _8581_ = m_17[78] & _8579_ /*16406*/;
  assign r_17[78] = _8581_ | _8580_ /*16405*/;
  assign _8582_ = ~q[15] /*16404*/;
  assign _8583_ = sum_17[79] & q[15] /*16403*/;
  assign _8584_ = m_17[79] & _8582_ /*16402*/;
  assign r_17[79] = _8584_ | _8583_ /*16401*/;
  assign inv_18[0] = oneWire /*16204*/;
  assign inv_18[1] = oneWire /*16198*/;
  assign inv_18[2] = oneWire /*16192*/;
  assign inv_18[3] = oneWire /*16186*/;
  assign inv_18[4] = oneWire /*16180*/;
  assign inv_18[5] = oneWire /*16174*/;
  assign inv_18[6] = oneWire /*16168*/;
  assign inv_18[7] = oneWire /*16162*/;
  assign inv_18[8] = oneWire /*16156*/;
  assign inv_18[9] = oneWire /*16150*/;
  assign inv_18[10] = oneWire /*16144*/;
  assign inv_18[11] = oneWire /*16138*/;
  assign inv_18[12] = oneWire /*16132*/;
  assign inv_18[13] = oneWire /*16126*/;
  assign inv_18[14] = ~div[0] /*16120*/;
  assign inv_18[15] = ~div[1] /*16114*/;
  assign inv_18[16] = ~div[2] /*16108*/;
  assign inv_18[17] = ~div[3] /*16102*/;
  assign inv_18[18] = ~div[4] /*16096*/;
  assign inv_18[19] = ~div[5] /*16090*/;
  assign inv_18[20] = ~div[6] /*16084*/;
  assign inv_18[21] = ~div[7] /*16078*/;
  assign inv_18[22] = ~div[8] /*16072*/;
  assign inv_18[23] = ~div[9] /*16066*/;
  assign inv_18[24] = ~div[10] /*16060*/;
  assign inv_18[25] = ~div[11] /*16054*/;
  assign inv_18[26] = ~div[12] /*16048*/;
  assign inv_18[27] = ~div[13] /*16042*/;
  assign inv_18[28] = ~div[14] /*16036*/;
  assign inv_18[29] = ~div[15] /*16030*/;
  assign inv_18[30] = ~div[16] /*16024*/;
  assign inv_18[31] = ~div[17] /*16018*/;
  assign inv_18[32] = ~div[18] /*16012*/;
  assign inv_18[33] = ~div[19] /*16006*/;
  assign inv_18[34] = ~div[20] /*16000*/;
  assign inv_18[35] = ~div[21] /*15994*/;
  assign inv_18[36] = ~div[22] /*15988*/;
  assign inv_18[37] = ~div[23] /*15982*/;
  assign inv_18[38] = ~div[24] /*15976*/;
  assign inv_18[39] = ~div[25] /*15970*/;
  assign inv_18[40] = ~div[26] /*15964*/;
  assign inv_18[41] = ~div[27] /*15958*/;
  assign inv_18[42] = ~div[28] /*15952*/;
  assign inv_18[43] = ~div[29] /*15946*/;
  assign inv_18[44] = ~div[30] /*15940*/;
  assign inv_18[45] = oneWire /*15934*/;
  assign inv_18[46] = oneWire /*15928*/;
  assign inv_18[47] = oneWire /*15922*/;
  assign inv_18[48] = oneWire /*15916*/;
  assign inv_18[49] = oneWire /*15910*/;
  assign inv_18[50] = oneWire /*15904*/;
  assign inv_18[51] = oneWire /*15898*/;
  assign inv_18[52] = oneWire /*15892*/;
  assign inv_18[53] = oneWire /*15886*/;
  assign inv_18[54] = oneWire /*15880*/;
  assign inv_18[55] = oneWire /*15874*/;
  assign inv_18[56] = oneWire /*15868*/;
  assign inv_18[57] = oneWire /*15862*/;
  assign inv_18[58] = oneWire /*15856*/;
  assign inv_18[59] = oneWire /*15850*/;
  assign inv_18[60] = oneWire /*15844*/;
  assign inv_18[61] = oneWire /*15838*/;
  assign inv_18[62] = oneWire /*15832*/;
  assign inv_18[63] = oneWire /*15826*/;
  assign inv_18[64] = oneWire /*15820*/;
  assign inv_18[65] = oneWire /*15814*/;
  assign inv_18[66] = oneWire /*15808*/;
  assign inv_18[67] = oneWire /*15802*/;
  assign inv_18[68] = oneWire /*15796*/;
  assign inv_18[69] = oneWire /*15790*/;
  assign inv_18[70] = oneWire /*15784*/;
  assign inv_18[71] = oneWire /*15778*/;
  assign inv_18[72] = oneWire /*15772*/;
  assign inv_18[73] = oneWire /*15766*/;
  assign inv_18[74] = oneWire /*15760*/;
  assign inv_18[75] = oneWire /*15754*/;
  assign inv_18[76] = oneWire /*15748*/;
  assign inv_18[77] = oneWire /*15742*/;
  assign inv_18[78] = oneWire /*15736*/;
  assign inv_18[79] = oneWire /*15730*/;
  assign _8585_ = inv_18[0] ^ r_17[0] /*16203*/;
  assign sum_18[0] = _8585_ ^ oneWire /*16202*/;
  assign _8586_ = _8585_ & oneWire /*16201*/;
  assign _8587_ = inv_18[0] & r_17[0] /*16200*/;
  assign _8588_ = _8586_ | _8587_ /*16199*/;
  assign _8589_ = inv_18[1] ^ r_17[1] /*16197*/;
  assign sum_18[1] = _8589_ ^ _8588_ /*16196*/;
  assign _8590_ = _8589_ & _8588_ /*16195*/;
  assign _8591_ = inv_18[1] & r_17[1] /*16194*/;
  assign _8592_ = _8590_ | _8591_ /*16193*/;
  assign _8593_ = inv_18[2] ^ r_17[2] /*16191*/;
  assign sum_18[2] = _8593_ ^ _8592_ /*16190*/;
  assign _8594_ = _8593_ & _8592_ /*16189*/;
  assign _8595_ = inv_18[2] & r_17[2] /*16188*/;
  assign _8596_ = _8594_ | _8595_ /*16187*/;
  assign _8597_ = inv_18[3] ^ r_17[3] /*16185*/;
  assign sum_18[3] = _8597_ ^ _8596_ /*16184*/;
  assign _8598_ = _8597_ & _8596_ /*16183*/;
  assign _8599_ = inv_18[3] & r_17[3] /*16182*/;
  assign _8600_ = _8598_ | _8599_ /*16181*/;
  assign _8601_ = inv_18[4] ^ r_17[4] /*16179*/;
  assign sum_18[4] = _8601_ ^ _8600_ /*16178*/;
  assign _8602_ = _8601_ & _8600_ /*16177*/;
  assign _8603_ = inv_18[4] & r_17[4] /*16176*/;
  assign _8604_ = _8602_ | _8603_ /*16175*/;
  assign _8605_ = inv_18[5] ^ r_17[5] /*16173*/;
  assign sum_18[5] = _8605_ ^ _8604_ /*16172*/;
  assign _8606_ = _8605_ & _8604_ /*16171*/;
  assign _8607_ = inv_18[5] & r_17[5] /*16170*/;
  assign _8608_ = _8606_ | _8607_ /*16169*/;
  assign _8609_ = inv_18[6] ^ r_17[6] /*16167*/;
  assign sum_18[6] = _8609_ ^ _8608_ /*16166*/;
  assign _8610_ = _8609_ & _8608_ /*16165*/;
  assign _8611_ = inv_18[6] & r_17[6] /*16164*/;
  assign _8612_ = _8610_ | _8611_ /*16163*/;
  assign _8613_ = inv_18[7] ^ r_17[7] /*16161*/;
  assign sum_18[7] = _8613_ ^ _8612_ /*16160*/;
  assign _8614_ = _8613_ & _8612_ /*16159*/;
  assign _8615_ = inv_18[7] & r_17[7] /*16158*/;
  assign _8616_ = _8614_ | _8615_ /*16157*/;
  assign _8617_ = inv_18[8] ^ r_17[8] /*16155*/;
  assign sum_18[8] = _8617_ ^ _8616_ /*16154*/;
  assign _8618_ = _8617_ & _8616_ /*16153*/;
  assign _8619_ = inv_18[8] & r_17[8] /*16152*/;
  assign _8620_ = _8618_ | _8619_ /*16151*/;
  assign _8621_ = inv_18[9] ^ r_17[9] /*16149*/;
  assign sum_18[9] = _8621_ ^ _8620_ /*16148*/;
  assign _8622_ = _8621_ & _8620_ /*16147*/;
  assign _8623_ = inv_18[9] & r_17[9] /*16146*/;
  assign _8624_ = _8622_ | _8623_ /*16145*/;
  assign _8625_ = inv_18[10] ^ r_17[10] /*16143*/;
  assign sum_18[10] = _8625_ ^ _8624_ /*16142*/;
  assign _8626_ = _8625_ & _8624_ /*16141*/;
  assign _8627_ = inv_18[10] & r_17[10] /*16140*/;
  assign _8628_ = _8626_ | _8627_ /*16139*/;
  assign _8629_ = inv_18[11] ^ r_17[11] /*16137*/;
  assign sum_18[11] = _8629_ ^ _8628_ /*16136*/;
  assign _8630_ = _8629_ & _8628_ /*16135*/;
  assign _8631_ = inv_18[11] & r_17[11] /*16134*/;
  assign _8632_ = _8630_ | _8631_ /*16133*/;
  assign _8633_ = inv_18[12] ^ r_17[12] /*16131*/;
  assign sum_18[12] = _8633_ ^ _8632_ /*16130*/;
  assign _8634_ = _8633_ & _8632_ /*16129*/;
  assign _8635_ = inv_18[12] & r_17[12] /*16128*/;
  assign _8636_ = _8634_ | _8635_ /*16127*/;
  assign _8637_ = inv_18[13] ^ r_17[13] /*16125*/;
  assign sum_18[13] = _8637_ ^ _8636_ /*16124*/;
  assign _8638_ = _8637_ & _8636_ /*16123*/;
  assign _8639_ = inv_18[13] & r_17[13] /*16122*/;
  assign _8640_ = _8638_ | _8639_ /*16121*/;
  assign _8641_ = inv_18[14] ^ r_17[14] /*16119*/;
  assign sum_18[14] = _8641_ ^ _8640_ /*16118*/;
  assign _8642_ = _8641_ & _8640_ /*16117*/;
  assign _8643_ = inv_18[14] & r_17[14] /*16116*/;
  assign _8644_ = _8642_ | _8643_ /*16115*/;
  assign _8645_ = inv_18[15] ^ r_17[15] /*16113*/;
  assign sum_18[15] = _8645_ ^ _8644_ /*16112*/;
  assign _8646_ = _8645_ & _8644_ /*16111*/;
  assign _8647_ = inv_18[15] & r_17[15] /*16110*/;
  assign _8648_ = _8646_ | _8647_ /*16109*/;
  assign _8649_ = inv_18[16] ^ r_17[16] /*16107*/;
  assign sum_18[16] = _8649_ ^ _8648_ /*16106*/;
  assign _8650_ = _8649_ & _8648_ /*16105*/;
  assign _8651_ = inv_18[16] & r_17[16] /*16104*/;
  assign _8652_ = _8650_ | _8651_ /*16103*/;
  assign _8653_ = inv_18[17] ^ r_17[17] /*16101*/;
  assign sum_18[17] = _8653_ ^ _8652_ /*16100*/;
  assign _8654_ = _8653_ & _8652_ /*16099*/;
  assign _8655_ = inv_18[17] & r_17[17] /*16098*/;
  assign _8656_ = _8654_ | _8655_ /*16097*/;
  assign _8657_ = inv_18[18] ^ r_17[18] /*16095*/;
  assign sum_18[18] = _8657_ ^ _8656_ /*16094*/;
  assign _8658_ = _8657_ & _8656_ /*16093*/;
  assign _8659_ = inv_18[18] & r_17[18] /*16092*/;
  assign _8660_ = _8658_ | _8659_ /*16091*/;
  assign _8661_ = inv_18[19] ^ r_17[19] /*16089*/;
  assign sum_18[19] = _8661_ ^ _8660_ /*16088*/;
  assign _8662_ = _8661_ & _8660_ /*16087*/;
  assign _8663_ = inv_18[19] & r_17[19] /*16086*/;
  assign _8664_ = _8662_ | _8663_ /*16085*/;
  assign _8665_ = inv_18[20] ^ r_17[20] /*16083*/;
  assign sum_18[20] = _8665_ ^ _8664_ /*16082*/;
  assign _8666_ = _8665_ & _8664_ /*16081*/;
  assign _8667_ = inv_18[20] & r_17[20] /*16080*/;
  assign _8668_ = _8666_ | _8667_ /*16079*/;
  assign _8669_ = inv_18[21] ^ r_17[21] /*16077*/;
  assign sum_18[21] = _8669_ ^ _8668_ /*16076*/;
  assign _8670_ = _8669_ & _8668_ /*16075*/;
  assign _8671_ = inv_18[21] & r_17[21] /*16074*/;
  assign _8672_ = _8670_ | _8671_ /*16073*/;
  assign _8673_ = inv_18[22] ^ r_17[22] /*16071*/;
  assign sum_18[22] = _8673_ ^ _8672_ /*16070*/;
  assign _8674_ = _8673_ & _8672_ /*16069*/;
  assign _8675_ = inv_18[22] & r_17[22] /*16068*/;
  assign _8676_ = _8674_ | _8675_ /*16067*/;
  assign _8677_ = inv_18[23] ^ r_17[23] /*16065*/;
  assign sum_18[23] = _8677_ ^ _8676_ /*16064*/;
  assign _8678_ = _8677_ & _8676_ /*16063*/;
  assign _8679_ = inv_18[23] & r_17[23] /*16062*/;
  assign _8680_ = _8678_ | _8679_ /*16061*/;
  assign _8681_ = inv_18[24] ^ r_17[24] /*16059*/;
  assign sum_18[24] = _8681_ ^ _8680_ /*16058*/;
  assign _8682_ = _8681_ & _8680_ /*16057*/;
  assign _8683_ = inv_18[24] & r_17[24] /*16056*/;
  assign _8684_ = _8682_ | _8683_ /*16055*/;
  assign _8685_ = inv_18[25] ^ r_17[25] /*16053*/;
  assign sum_18[25] = _8685_ ^ _8684_ /*16052*/;
  assign _8686_ = _8685_ & _8684_ /*16051*/;
  assign _8687_ = inv_18[25] & r_17[25] /*16050*/;
  assign _8688_ = _8686_ | _8687_ /*16049*/;
  assign _8689_ = inv_18[26] ^ r_17[26] /*16047*/;
  assign sum_18[26] = _8689_ ^ _8688_ /*16046*/;
  assign _8690_ = _8689_ & _8688_ /*16045*/;
  assign _8691_ = inv_18[26] & r_17[26] /*16044*/;
  assign _8692_ = _8690_ | _8691_ /*16043*/;
  assign _8693_ = inv_18[27] ^ r_17[27] /*16041*/;
  assign sum_18[27] = _8693_ ^ _8692_ /*16040*/;
  assign _8694_ = _8693_ & _8692_ /*16039*/;
  assign _8695_ = inv_18[27] & r_17[27] /*16038*/;
  assign _8696_ = _8694_ | _8695_ /*16037*/;
  assign _8697_ = inv_18[28] ^ r_17[28] /*16035*/;
  assign sum_18[28] = _8697_ ^ _8696_ /*16034*/;
  assign _8698_ = _8697_ & _8696_ /*16033*/;
  assign _8699_ = inv_18[28] & r_17[28] /*16032*/;
  assign _8700_ = _8698_ | _8699_ /*16031*/;
  assign _8701_ = inv_18[29] ^ r_17[29] /*16029*/;
  assign sum_18[29] = _8701_ ^ _8700_ /*16028*/;
  assign _8702_ = _8701_ & _8700_ /*16027*/;
  assign _8703_ = inv_18[29] & r_17[29] /*16026*/;
  assign _8704_ = _8702_ | _8703_ /*16025*/;
  assign _8705_ = inv_18[30] ^ r_17[30] /*16023*/;
  assign sum_18[30] = _8705_ ^ _8704_ /*16022*/;
  assign _8706_ = _8705_ & _8704_ /*16021*/;
  assign _8707_ = inv_18[30] & r_17[30] /*16020*/;
  assign _8708_ = _8706_ | _8707_ /*16019*/;
  assign _8709_ = inv_18[31] ^ r_17[31] /*16017*/;
  assign sum_18[31] = _8709_ ^ _8708_ /*16016*/;
  assign _8710_ = _8709_ & _8708_ /*16015*/;
  assign _8711_ = inv_18[31] & r_17[31] /*16014*/;
  assign _8712_ = _8710_ | _8711_ /*16013*/;
  assign _8713_ = inv_18[32] ^ r_17[32] /*16011*/;
  assign sum_18[32] = _8713_ ^ _8712_ /*16010*/;
  assign _8714_ = _8713_ & _8712_ /*16009*/;
  assign _8715_ = inv_18[32] & r_17[32] /*16008*/;
  assign _8716_ = _8714_ | _8715_ /*16007*/;
  assign _8717_ = inv_18[33] ^ r_17[33] /*16005*/;
  assign sum_18[33] = _8717_ ^ _8716_ /*16004*/;
  assign _8718_ = _8717_ & _8716_ /*16003*/;
  assign _8719_ = inv_18[33] & r_17[33] /*16002*/;
  assign _8720_ = _8718_ | _8719_ /*16001*/;
  assign _8721_ = inv_18[34] ^ r_17[34] /*15999*/;
  assign sum_18[34] = _8721_ ^ _8720_ /*15998*/;
  assign _8722_ = _8721_ & _8720_ /*15997*/;
  assign _8723_ = inv_18[34] & r_17[34] /*15996*/;
  assign _8724_ = _8722_ | _8723_ /*15995*/;
  assign _8725_ = inv_18[35] ^ r_17[35] /*15993*/;
  assign sum_18[35] = _8725_ ^ _8724_ /*15992*/;
  assign _8726_ = _8725_ & _8724_ /*15991*/;
  assign _8727_ = inv_18[35] & r_17[35] /*15990*/;
  assign _8728_ = _8726_ | _8727_ /*15989*/;
  assign _8729_ = inv_18[36] ^ r_17[36] /*15987*/;
  assign sum_18[36] = _8729_ ^ _8728_ /*15986*/;
  assign _8730_ = _8729_ & _8728_ /*15985*/;
  assign _8731_ = inv_18[36] & r_17[36] /*15984*/;
  assign _8732_ = _8730_ | _8731_ /*15983*/;
  assign _8733_ = inv_18[37] ^ r_17[37] /*15981*/;
  assign sum_18[37] = _8733_ ^ _8732_ /*15980*/;
  assign _8734_ = _8733_ & _8732_ /*15979*/;
  assign _8735_ = inv_18[37] & r_17[37] /*15978*/;
  assign _8736_ = _8734_ | _8735_ /*15977*/;
  assign _8737_ = inv_18[38] ^ r_17[38] /*15975*/;
  assign sum_18[38] = _8737_ ^ _8736_ /*15974*/;
  assign _8738_ = _8737_ & _8736_ /*15973*/;
  assign _8739_ = inv_18[38] & r_17[38] /*15972*/;
  assign _8740_ = _8738_ | _8739_ /*15971*/;
  assign _8741_ = inv_18[39] ^ r_17[39] /*15969*/;
  assign sum_18[39] = _8741_ ^ _8740_ /*15968*/;
  assign _8742_ = _8741_ & _8740_ /*15967*/;
  assign _8743_ = inv_18[39] & r_17[39] /*15966*/;
  assign _8744_ = _8742_ | _8743_ /*15965*/;
  assign _8745_ = inv_18[40] ^ r_17[40] /*15963*/;
  assign sum_18[40] = _8745_ ^ _8744_ /*15962*/;
  assign _8746_ = _8745_ & _8744_ /*15961*/;
  assign _8747_ = inv_18[40] & r_17[40] /*15960*/;
  assign _8748_ = _8746_ | _8747_ /*15959*/;
  assign _8749_ = inv_18[41] ^ r_17[41] /*15957*/;
  assign sum_18[41] = _8749_ ^ _8748_ /*15956*/;
  assign _8750_ = _8749_ & _8748_ /*15955*/;
  assign _8751_ = inv_18[41] & r_17[41] /*15954*/;
  assign _8752_ = _8750_ | _8751_ /*15953*/;
  assign _8753_ = inv_18[42] ^ r_17[42] /*15951*/;
  assign sum_18[42] = _8753_ ^ _8752_ /*15950*/;
  assign _8754_ = _8753_ & _8752_ /*15949*/;
  assign _8755_ = inv_18[42] & r_17[42] /*15948*/;
  assign _8756_ = _8754_ | _8755_ /*15947*/;
  assign _8757_ = inv_18[43] ^ r_17[43] /*15945*/;
  assign sum_18[43] = _8757_ ^ _8756_ /*15944*/;
  assign _8758_ = _8757_ & _8756_ /*15943*/;
  assign _8759_ = inv_18[43] & r_17[43] /*15942*/;
  assign _8760_ = _8758_ | _8759_ /*15941*/;
  assign _8761_ = inv_18[44] ^ r_17[44] /*15939*/;
  assign sum_18[44] = _8761_ ^ _8760_ /*15938*/;
  assign _8762_ = _8761_ & _8760_ /*15937*/;
  assign _8763_ = inv_18[44] & r_17[44] /*15936*/;
  assign _8764_ = _8762_ | _8763_ /*15935*/;
  assign _8765_ = inv_18[45] ^ r_17[45] /*15933*/;
  assign sum_18[45] = _8765_ ^ _8764_ /*15932*/;
  assign _8766_ = _8765_ & _8764_ /*15931*/;
  assign _8767_ = inv_18[45] & r_17[45] /*15930*/;
  assign _8768_ = _8766_ | _8767_ /*15929*/;
  assign _8769_ = inv_18[46] ^ r_17[46] /*15927*/;
  assign sum_18[46] = _8769_ ^ _8768_ /*15926*/;
  assign _8770_ = _8769_ & _8768_ /*15925*/;
  assign _8771_ = inv_18[46] & r_17[46] /*15924*/;
  assign _8772_ = _8770_ | _8771_ /*15923*/;
  assign _8773_ = inv_18[47] ^ r_17[47] /*15921*/;
  assign sum_18[47] = _8773_ ^ _8772_ /*15920*/;
  assign _8774_ = _8773_ & _8772_ /*15919*/;
  assign _8775_ = inv_18[47] & r_17[47] /*15918*/;
  assign _8776_ = _8774_ | _8775_ /*15917*/;
  assign _8777_ = inv_18[48] ^ r_17[48] /*15915*/;
  assign sum_18[48] = _8777_ ^ _8776_ /*15914*/;
  assign _8778_ = _8777_ & _8776_ /*15913*/;
  assign _8779_ = inv_18[48] & r_17[48] /*15912*/;
  assign _8780_ = _8778_ | _8779_ /*15911*/;
  assign _8781_ = inv_18[49] ^ r_17[49] /*15909*/;
  assign sum_18[49] = _8781_ ^ _8780_ /*15908*/;
  assign _8782_ = _8781_ & _8780_ /*15907*/;
  assign _8783_ = inv_18[49] & r_17[49] /*15906*/;
  assign _8784_ = _8782_ | _8783_ /*15905*/;
  assign _8785_ = inv_18[50] ^ r_17[50] /*15903*/;
  assign sum_18[50] = _8785_ ^ _8784_ /*15902*/;
  assign _8786_ = _8785_ & _8784_ /*15901*/;
  assign _8787_ = inv_18[50] & r_17[50] /*15900*/;
  assign _8788_ = _8786_ | _8787_ /*15899*/;
  assign _8789_ = inv_18[51] ^ r_17[51] /*15897*/;
  assign sum_18[51] = _8789_ ^ _8788_ /*15896*/;
  assign _8790_ = _8789_ & _8788_ /*15895*/;
  assign _8791_ = inv_18[51] & r_17[51] /*15894*/;
  assign _8792_ = _8790_ | _8791_ /*15893*/;
  assign _8793_ = inv_18[52] ^ r_17[52] /*15891*/;
  assign sum_18[52] = _8793_ ^ _8792_ /*15890*/;
  assign _8794_ = _8793_ & _8792_ /*15889*/;
  assign _8795_ = inv_18[52] & r_17[52] /*15888*/;
  assign _8796_ = _8794_ | _8795_ /*15887*/;
  assign _8797_ = inv_18[53] ^ r_17[53] /*15885*/;
  assign sum_18[53] = _8797_ ^ _8796_ /*15884*/;
  assign _8798_ = _8797_ & _8796_ /*15883*/;
  assign _8799_ = inv_18[53] & r_17[53] /*15882*/;
  assign _8800_ = _8798_ | _8799_ /*15881*/;
  assign _8801_ = inv_18[54] ^ r_17[54] /*15879*/;
  assign sum_18[54] = _8801_ ^ _8800_ /*15878*/;
  assign _8802_ = _8801_ & _8800_ /*15877*/;
  assign _8803_ = inv_18[54] & r_17[54] /*15876*/;
  assign _8804_ = _8802_ | _8803_ /*15875*/;
  assign _8805_ = inv_18[55] ^ r_17[55] /*15873*/;
  assign sum_18[55] = _8805_ ^ _8804_ /*15872*/;
  assign _8806_ = _8805_ & _8804_ /*15871*/;
  assign _8807_ = inv_18[55] & r_17[55] /*15870*/;
  assign _8808_ = _8806_ | _8807_ /*15869*/;
  assign _8809_ = inv_18[56] ^ r_17[56] /*15867*/;
  assign sum_18[56] = _8809_ ^ _8808_ /*15866*/;
  assign _8810_ = _8809_ & _8808_ /*15865*/;
  assign _8811_ = inv_18[56] & r_17[56] /*15864*/;
  assign _8812_ = _8810_ | _8811_ /*15863*/;
  assign _8813_ = inv_18[57] ^ r_17[57] /*15861*/;
  assign sum_18[57] = _8813_ ^ _8812_ /*15860*/;
  assign _8814_ = _8813_ & _8812_ /*15859*/;
  assign _8815_ = inv_18[57] & r_17[57] /*15858*/;
  assign _8816_ = _8814_ | _8815_ /*15857*/;
  assign _8817_ = inv_18[58] ^ r_17[58] /*15855*/;
  assign sum_18[58] = _8817_ ^ _8816_ /*15854*/;
  assign _8818_ = _8817_ & _8816_ /*15853*/;
  assign _8819_ = inv_18[58] & r_17[58] /*15852*/;
  assign _8820_ = _8818_ | _8819_ /*15851*/;
  assign _8821_ = inv_18[59] ^ r_17[59] /*15849*/;
  assign sum_18[59] = _8821_ ^ _8820_ /*15848*/;
  assign _8822_ = _8821_ & _8820_ /*15847*/;
  assign _8823_ = inv_18[59] & r_17[59] /*15846*/;
  assign _8824_ = _8822_ | _8823_ /*15845*/;
  assign _8825_ = inv_18[60] ^ r_17[60] /*15843*/;
  assign sum_18[60] = _8825_ ^ _8824_ /*15842*/;
  assign _8826_ = _8825_ & _8824_ /*15841*/;
  assign _8827_ = inv_18[60] & r_17[60] /*15840*/;
  assign _8828_ = _8826_ | _8827_ /*15839*/;
  assign _8829_ = inv_18[61] ^ r_17[61] /*15837*/;
  assign sum_18[61] = _8829_ ^ _8828_ /*15836*/;
  assign _8830_ = _8829_ & _8828_ /*15835*/;
  assign _8831_ = inv_18[61] & r_17[61] /*15834*/;
  assign _8832_ = _8830_ | _8831_ /*15833*/;
  assign _8833_ = inv_18[62] ^ r_17[62] /*15831*/;
  assign sum_18[62] = _8833_ ^ _8832_ /*15830*/;
  assign _8834_ = _8833_ & _8832_ /*15829*/;
  assign _8835_ = inv_18[62] & r_17[62] /*15828*/;
  assign _8836_ = _8834_ | _8835_ /*15827*/;
  assign _8837_ = inv_18[63] ^ r_17[63] /*15825*/;
  assign sum_18[63] = _8837_ ^ _8836_ /*15824*/;
  assign _8838_ = _8837_ & _8836_ /*15823*/;
  assign _8839_ = inv_18[63] & r_17[63] /*15822*/;
  assign _8840_ = _8838_ | _8839_ /*15821*/;
  assign _8841_ = inv_18[64] ^ r_17[64] /*15819*/;
  assign sum_18[64] = _8841_ ^ _8840_ /*15818*/;
  assign _8842_ = _8841_ & _8840_ /*15817*/;
  assign _8843_ = inv_18[64] & r_17[64] /*15816*/;
  assign _8844_ = _8842_ | _8843_ /*15815*/;
  assign _8845_ = inv_18[65] ^ r_17[65] /*15813*/;
  assign sum_18[65] = _8845_ ^ _8844_ /*15812*/;
  assign _8846_ = _8845_ & _8844_ /*15811*/;
  assign _8847_ = inv_18[65] & r_17[65] /*15810*/;
  assign _8848_ = _8846_ | _8847_ /*15809*/;
  assign _8849_ = inv_18[66] ^ r_17[66] /*15807*/;
  assign sum_18[66] = _8849_ ^ _8848_ /*15806*/;
  assign _8850_ = _8849_ & _8848_ /*15805*/;
  assign _8851_ = inv_18[66] & r_17[66] /*15804*/;
  assign _8852_ = _8850_ | _8851_ /*15803*/;
  assign _8853_ = inv_18[67] ^ r_17[67] /*15801*/;
  assign sum_18[67] = _8853_ ^ _8852_ /*15800*/;
  assign _8854_ = _8853_ & _8852_ /*15799*/;
  assign _8855_ = inv_18[67] & r_17[67] /*15798*/;
  assign _8856_ = _8854_ | _8855_ /*15797*/;
  assign _8857_ = inv_18[68] ^ r_17[68] /*15795*/;
  assign sum_18[68] = _8857_ ^ _8856_ /*15794*/;
  assign _8858_ = _8857_ & _8856_ /*15793*/;
  assign _8859_ = inv_18[68] & r_17[68] /*15792*/;
  assign _8860_ = _8858_ | _8859_ /*15791*/;
  assign _8861_ = inv_18[69] ^ r_17[69] /*15789*/;
  assign sum_18[69] = _8861_ ^ _8860_ /*15788*/;
  assign _8862_ = _8861_ & _8860_ /*15787*/;
  assign _8863_ = inv_18[69] & r_17[69] /*15786*/;
  assign _8864_ = _8862_ | _8863_ /*15785*/;
  assign _8865_ = inv_18[70] ^ r_17[70] /*15783*/;
  assign sum_18[70] = _8865_ ^ _8864_ /*15782*/;
  assign _8866_ = _8865_ & _8864_ /*15781*/;
  assign _8867_ = inv_18[70] & r_17[70] /*15780*/;
  assign _8868_ = _8866_ | _8867_ /*15779*/;
  assign _8869_ = inv_18[71] ^ r_17[71] /*15777*/;
  assign sum_18[71] = _8869_ ^ _8868_ /*15776*/;
  assign _8870_ = _8869_ & _8868_ /*15775*/;
  assign _8871_ = inv_18[71] & r_17[71] /*15774*/;
  assign _8872_ = _8870_ | _8871_ /*15773*/;
  assign _8873_ = inv_18[72] ^ r_17[72] /*15771*/;
  assign sum_18[72] = _8873_ ^ _8872_ /*15770*/;
  assign _8874_ = _8873_ & _8872_ /*15769*/;
  assign _8875_ = inv_18[72] & r_17[72] /*15768*/;
  assign _8876_ = _8874_ | _8875_ /*15767*/;
  assign _8877_ = inv_18[73] ^ r_17[73] /*15765*/;
  assign sum_18[73] = _8877_ ^ _8876_ /*15764*/;
  assign _8878_ = _8877_ & _8876_ /*15763*/;
  assign _8879_ = inv_18[73] & r_17[73] /*15762*/;
  assign _8880_ = _8878_ | _8879_ /*15761*/;
  assign _8881_ = inv_18[74] ^ r_17[74] /*15759*/;
  assign sum_18[74] = _8881_ ^ _8880_ /*15758*/;
  assign _8882_ = _8881_ & _8880_ /*15757*/;
  assign _8883_ = inv_18[74] & r_17[74] /*15756*/;
  assign _8884_ = _8882_ | _8883_ /*15755*/;
  assign _8885_ = inv_18[75] ^ r_17[75] /*15753*/;
  assign sum_18[75] = _8885_ ^ _8884_ /*15752*/;
  assign _8886_ = _8885_ & _8884_ /*15751*/;
  assign _8887_ = inv_18[75] & r_17[75] /*15750*/;
  assign _8888_ = _8886_ | _8887_ /*15749*/;
  assign _8889_ = inv_18[76] ^ r_17[76] /*15747*/;
  assign sum_18[76] = _8889_ ^ _8888_ /*15746*/;
  assign _8890_ = _8889_ & _8888_ /*15745*/;
  assign _8891_ = inv_18[76] & r_17[76] /*15744*/;
  assign _8892_ = _8890_ | _8891_ /*15743*/;
  assign _8893_ = inv_18[77] ^ r_17[77] /*15741*/;
  assign sum_18[77] = _8893_ ^ _8892_ /*15740*/;
  assign _8894_ = _8893_ & _8892_ /*15739*/;
  assign _8895_ = inv_18[77] & r_17[77] /*15738*/;
  assign _8896_ = _8894_ | _8895_ /*15737*/;
  assign _8897_ = inv_18[78] ^ r_17[78] /*15735*/;
  assign sum_18[78] = _8897_ ^ _8896_ /*15734*/;
  assign _8898_ = _8897_ & _8896_ /*15733*/;
  assign _8899_ = inv_18[78] & r_17[78] /*15732*/;
  assign _8900_ = _8898_ | _8899_ /*15731*/;
  assign _8901_ = inv_18[79] ^ r_17[79] /*15729*/;
  assign sum_18[79] = _8901_ ^ _8900_ /*15728*/;
  assign _8902_ = _8901_ & _8900_ /*15727*/;
  assign _8903_ = inv_18[79] & r_17[79] /*15726*/;
  assign _8904_ = _8902_ | _8903_ /*15725*/;
  assign _8905_ = _8904_ ^ _8900_ /*15724*/;
  assign _8906_ = ~_8905_ /*15723*/;
  assign _8907_ = sum_18[79] & _8906_ /*15722*/;
  assign _8908_ = _8905_ & _8904_ /*15721*/;
  assign sum_18[80] = _8908_ | _8907_ /*15720*/;
  assign q[14] = ~sum_18[80] /*15719*/;
  assign m_18[0] = r_17[0] /*15718*/;
  assign m_18[1] = r_17[1] /*15717*/;
  assign m_18[2] = r_17[2] /*15716*/;
  assign m_18[3] = r_17[3] /*15715*/;
  assign m_18[4] = r_17[4] /*15714*/;
  assign m_18[5] = r_17[5] /*15713*/;
  assign m_18[6] = r_17[6] /*15712*/;
  assign m_18[7] = r_17[7] /*15711*/;
  assign m_18[8] = r_17[8] /*15710*/;
  assign m_18[9] = r_17[9] /*15709*/;
  assign m_18[10] = r_17[10] /*15708*/;
  assign m_18[11] = r_17[11] /*15707*/;
  assign m_18[12] = r_17[12] /*15706*/;
  assign m_18[13] = r_17[13] /*15705*/;
  assign m_18[14] = r_17[14] /*15704*/;
  assign m_18[15] = r_17[15] /*15703*/;
  assign m_18[16] = r_17[16] /*15702*/;
  assign m_18[17] = r_17[17] /*15701*/;
  assign m_18[18] = r_17[18] /*15700*/;
  assign m_18[19] = r_17[19] /*15699*/;
  assign m_18[20] = r_17[20] /*15698*/;
  assign m_18[21] = r_17[21] /*15697*/;
  assign m_18[22] = r_17[22] /*15696*/;
  assign m_18[23] = r_17[23] /*15695*/;
  assign m_18[24] = r_17[24] /*15694*/;
  assign m_18[25] = r_17[25] /*15693*/;
  assign m_18[26] = r_17[26] /*15692*/;
  assign m_18[27] = r_17[27] /*15691*/;
  assign m_18[28] = r_17[28] /*15690*/;
  assign m_18[29] = r_17[29] /*15689*/;
  assign m_18[30] = r_17[30] /*15688*/;
  assign m_18[31] = r_17[31] /*15687*/;
  assign m_18[32] = r_17[32] /*15686*/;
  assign m_18[33] = r_17[33] /*15685*/;
  assign m_18[34] = r_17[34] /*15684*/;
  assign m_18[35] = r_17[35] /*15683*/;
  assign m_18[36] = r_17[36] /*15682*/;
  assign m_18[37] = r_17[37] /*15681*/;
  assign m_18[38] = r_17[38] /*15680*/;
  assign m_18[39] = r_17[39] /*15679*/;
  assign m_18[40] = r_17[40] /*15678*/;
  assign m_18[41] = r_17[41] /*15677*/;
  assign m_18[42] = r_17[42] /*15676*/;
  assign m_18[43] = r_17[43] /*15675*/;
  assign m_18[44] = r_17[44] /*15674*/;
  assign m_18[45] = r_17[45] /*15673*/;
  assign m_18[46] = r_17[46] /*15672*/;
  assign m_18[47] = r_17[47] /*15671*/;
  assign m_18[48] = r_17[48] /*15670*/;
  assign m_18[49] = r_17[49] /*15669*/;
  assign m_18[50] = r_17[50] /*15668*/;
  assign m_18[51] = r_17[51] /*15667*/;
  assign m_18[52] = r_17[52] /*15666*/;
  assign m_18[53] = r_17[53] /*15665*/;
  assign m_18[54] = r_17[54] /*15664*/;
  assign m_18[55] = r_17[55] /*15663*/;
  assign m_18[56] = r_17[56] /*15662*/;
  assign m_18[57] = r_17[57] /*15661*/;
  assign m_18[58] = r_17[58] /*15660*/;
  assign m_18[59] = r_17[59] /*15659*/;
  assign m_18[60] = r_17[60] /*15658*/;
  assign m_18[61] = r_17[61] /*15657*/;
  assign m_18[62] = r_17[62] /*15656*/;
  assign m_18[63] = r_17[63] /*15655*/;
  assign m_18[64] = r_17[64] /*15654*/;
  assign m_18[65] = r_17[65] /*15653*/;
  assign m_18[66] = r_17[66] /*15652*/;
  assign m_18[67] = r_17[67] /*15651*/;
  assign m_18[68] = r_17[68] /*15650*/;
  assign m_18[69] = r_17[69] /*15649*/;
  assign m_18[70] = r_17[70] /*15648*/;
  assign m_18[71] = r_17[71] /*15647*/;
  assign m_18[72] = r_17[72] /*15646*/;
  assign m_18[73] = r_17[73] /*15645*/;
  assign m_18[74] = r_17[74] /*15644*/;
  assign m_18[75] = r_17[75] /*15643*/;
  assign m_18[76] = r_17[76] /*15642*/;
  assign m_18[77] = r_17[77] /*15641*/;
  assign m_18[78] = r_17[78] /*15640*/;
  assign m_18[79] = r_17[79] /*15639*/;
  assign m_18[80] = r_17[79] /*15638*/;
  assign _8910_ = ~q[14] /*15637*/;
  assign _8911_ = sum_18[0] & q[14] /*15636*/;
  assign _8912_ = m_18[0] & _8910_ /*15635*/;
  assign r_18[0] = _8912_ | _8911_ /*15634*/;
  assign _8913_ = ~q[14] /*15633*/;
  assign _8914_ = sum_18[1] & q[14] /*15632*/;
  assign _8915_ = m_18[1] & _8913_ /*15631*/;
  assign r_18[1] = _8915_ | _8914_ /*15630*/;
  assign _8916_ = ~q[14] /*15629*/;
  assign _8917_ = sum_18[2] & q[14] /*15628*/;
  assign _8918_ = m_18[2] & _8916_ /*15627*/;
  assign r_18[2] = _8918_ | _8917_ /*15626*/;
  assign _8919_ = ~q[14] /*15625*/;
  assign _8920_ = sum_18[3] & q[14] /*15624*/;
  assign _8921_ = m_18[3] & _8919_ /*15623*/;
  assign r_18[3] = _8921_ | _8920_ /*15622*/;
  assign _8922_ = ~q[14] /*15621*/;
  assign _8923_ = sum_18[4] & q[14] /*15620*/;
  assign _8924_ = m_18[4] & _8922_ /*15619*/;
  assign r_18[4] = _8924_ | _8923_ /*15618*/;
  assign _8925_ = ~q[14] /*15617*/;
  assign _8926_ = sum_18[5] & q[14] /*15616*/;
  assign _8927_ = m_18[5] & _8925_ /*15615*/;
  assign r_18[5] = _8927_ | _8926_ /*15614*/;
  assign _8928_ = ~q[14] /*15613*/;
  assign _8929_ = sum_18[6] & q[14] /*15612*/;
  assign _8930_ = m_18[6] & _8928_ /*15611*/;
  assign r_18[6] = _8930_ | _8929_ /*15610*/;
  assign _8931_ = ~q[14] /*15609*/;
  assign _8932_ = sum_18[7] & q[14] /*15608*/;
  assign _8933_ = m_18[7] & _8931_ /*15607*/;
  assign r_18[7] = _8933_ | _8932_ /*15606*/;
  assign _8934_ = ~q[14] /*15605*/;
  assign _8935_ = sum_18[8] & q[14] /*15604*/;
  assign _8936_ = m_18[8] & _8934_ /*15603*/;
  assign r_18[8] = _8936_ | _8935_ /*15602*/;
  assign _8937_ = ~q[14] /*15601*/;
  assign _8938_ = sum_18[9] & q[14] /*15600*/;
  assign _8939_ = m_18[9] & _8937_ /*15599*/;
  assign r_18[9] = _8939_ | _8938_ /*15598*/;
  assign _8940_ = ~q[14] /*15597*/;
  assign _8941_ = sum_18[10] & q[14] /*15596*/;
  assign _8942_ = m_18[10] & _8940_ /*15595*/;
  assign r_18[10] = _8942_ | _8941_ /*15594*/;
  assign _8943_ = ~q[14] /*15593*/;
  assign _8944_ = sum_18[11] & q[14] /*15592*/;
  assign _8945_ = m_18[11] & _8943_ /*15591*/;
  assign r_18[11] = _8945_ | _8944_ /*15590*/;
  assign _8946_ = ~q[14] /*15589*/;
  assign _8947_ = sum_18[12] & q[14] /*15588*/;
  assign _8948_ = m_18[12] & _8946_ /*15587*/;
  assign r_18[12] = _8948_ | _8947_ /*15586*/;
  assign _8949_ = ~q[14] /*15585*/;
  assign _8950_ = sum_18[13] & q[14] /*15584*/;
  assign _8951_ = m_18[13] & _8949_ /*15583*/;
  assign r_18[13] = _8951_ | _8950_ /*15582*/;
  assign _8952_ = ~q[14] /*15581*/;
  assign _8953_ = sum_18[14] & q[14] /*15580*/;
  assign _8954_ = m_18[14] & _8952_ /*15579*/;
  assign r_18[14] = _8954_ | _8953_ /*15578*/;
  assign _8955_ = ~q[14] /*15577*/;
  assign _8956_ = sum_18[15] & q[14] /*15576*/;
  assign _8957_ = m_18[15] & _8955_ /*15575*/;
  assign r_18[15] = _8957_ | _8956_ /*15574*/;
  assign _8958_ = ~q[14] /*15573*/;
  assign _8959_ = sum_18[16] & q[14] /*15572*/;
  assign _8960_ = m_18[16] & _8958_ /*15571*/;
  assign r_18[16] = _8960_ | _8959_ /*15570*/;
  assign _8961_ = ~q[14] /*15569*/;
  assign _8962_ = sum_18[17] & q[14] /*15568*/;
  assign _8963_ = m_18[17] & _8961_ /*15567*/;
  assign r_18[17] = _8963_ | _8962_ /*15566*/;
  assign _8964_ = ~q[14] /*15565*/;
  assign _8965_ = sum_18[18] & q[14] /*15564*/;
  assign _8966_ = m_18[18] & _8964_ /*15563*/;
  assign r_18[18] = _8966_ | _8965_ /*15562*/;
  assign _8967_ = ~q[14] /*15561*/;
  assign _8968_ = sum_18[19] & q[14] /*15560*/;
  assign _8969_ = m_18[19] & _8967_ /*15559*/;
  assign r_18[19] = _8969_ | _8968_ /*15558*/;
  assign _8970_ = ~q[14] /*15557*/;
  assign _8971_ = sum_18[20] & q[14] /*15556*/;
  assign _8972_ = m_18[20] & _8970_ /*15555*/;
  assign r_18[20] = _8972_ | _8971_ /*15554*/;
  assign _8973_ = ~q[14] /*15553*/;
  assign _8974_ = sum_18[21] & q[14] /*15552*/;
  assign _8975_ = m_18[21] & _8973_ /*15551*/;
  assign r_18[21] = _8975_ | _8974_ /*15550*/;
  assign _8976_ = ~q[14] /*15549*/;
  assign _8977_ = sum_18[22] & q[14] /*15548*/;
  assign _8978_ = m_18[22] & _8976_ /*15547*/;
  assign r_18[22] = _8978_ | _8977_ /*15546*/;
  assign _8979_ = ~q[14] /*15545*/;
  assign _8980_ = sum_18[23] & q[14] /*15544*/;
  assign _8981_ = m_18[23] & _8979_ /*15543*/;
  assign r_18[23] = _8981_ | _8980_ /*15542*/;
  assign _8982_ = ~q[14] /*15541*/;
  assign _8983_ = sum_18[24] & q[14] /*15540*/;
  assign _8984_ = m_18[24] & _8982_ /*15539*/;
  assign r_18[24] = _8984_ | _8983_ /*15538*/;
  assign _8985_ = ~q[14] /*15537*/;
  assign _8986_ = sum_18[25] & q[14] /*15536*/;
  assign _8987_ = m_18[25] & _8985_ /*15535*/;
  assign r_18[25] = _8987_ | _8986_ /*15534*/;
  assign _8988_ = ~q[14] /*15533*/;
  assign _8989_ = sum_18[26] & q[14] /*15532*/;
  assign _8990_ = m_18[26] & _8988_ /*15531*/;
  assign r_18[26] = _8990_ | _8989_ /*15530*/;
  assign _8991_ = ~q[14] /*15529*/;
  assign _8992_ = sum_18[27] & q[14] /*15528*/;
  assign _8993_ = m_18[27] & _8991_ /*15527*/;
  assign r_18[27] = _8993_ | _8992_ /*15526*/;
  assign _8994_ = ~q[14] /*15525*/;
  assign _8995_ = sum_18[28] & q[14] /*15524*/;
  assign _8996_ = m_18[28] & _8994_ /*15523*/;
  assign r_18[28] = _8996_ | _8995_ /*15522*/;
  assign _8997_ = ~q[14] /*15521*/;
  assign _8998_ = sum_18[29] & q[14] /*15520*/;
  assign _8999_ = m_18[29] & _8997_ /*15519*/;
  assign r_18[29] = _8999_ | _8998_ /*15518*/;
  assign _9000_ = ~q[14] /*15517*/;
  assign _9001_ = sum_18[30] & q[14] /*15516*/;
  assign _9002_ = m_18[30] & _9000_ /*15515*/;
  assign r_18[30] = _9002_ | _9001_ /*15514*/;
  assign _9003_ = ~q[14] /*15513*/;
  assign _9004_ = sum_18[31] & q[14] /*15512*/;
  assign _9005_ = m_18[31] & _9003_ /*15511*/;
  assign r_18[31] = _9005_ | _9004_ /*15510*/;
  assign _9006_ = ~q[14] /*15509*/;
  assign _9007_ = sum_18[32] & q[14] /*15508*/;
  assign _9008_ = m_18[32] & _9006_ /*15507*/;
  assign r_18[32] = _9008_ | _9007_ /*15506*/;
  assign _9009_ = ~q[14] /*15505*/;
  assign _9010_ = sum_18[33] & q[14] /*15504*/;
  assign _9011_ = m_18[33] & _9009_ /*15503*/;
  assign r_18[33] = _9011_ | _9010_ /*15502*/;
  assign _9012_ = ~q[14] /*15501*/;
  assign _9013_ = sum_18[34] & q[14] /*15500*/;
  assign _9014_ = m_18[34] & _9012_ /*15499*/;
  assign r_18[34] = _9014_ | _9013_ /*15498*/;
  assign _9015_ = ~q[14] /*15497*/;
  assign _9016_ = sum_18[35] & q[14] /*15496*/;
  assign _9017_ = m_18[35] & _9015_ /*15495*/;
  assign r_18[35] = _9017_ | _9016_ /*15494*/;
  assign _9018_ = ~q[14] /*15493*/;
  assign _9019_ = sum_18[36] & q[14] /*15492*/;
  assign _9020_ = m_18[36] & _9018_ /*15491*/;
  assign r_18[36] = _9020_ | _9019_ /*15490*/;
  assign _9021_ = ~q[14] /*15489*/;
  assign _9022_ = sum_18[37] & q[14] /*15488*/;
  assign _9023_ = m_18[37] & _9021_ /*15487*/;
  assign r_18[37] = _9023_ | _9022_ /*15486*/;
  assign _9024_ = ~q[14] /*15485*/;
  assign _9025_ = sum_18[38] & q[14] /*15484*/;
  assign _9026_ = m_18[38] & _9024_ /*15483*/;
  assign r_18[38] = _9026_ | _9025_ /*15482*/;
  assign _9027_ = ~q[14] /*15481*/;
  assign _9028_ = sum_18[39] & q[14] /*15480*/;
  assign _9029_ = m_18[39] & _9027_ /*15479*/;
  assign r_18[39] = _9029_ | _9028_ /*15478*/;
  assign _9030_ = ~q[14] /*15477*/;
  assign _9031_ = sum_18[40] & q[14] /*15476*/;
  assign _9032_ = m_18[40] & _9030_ /*15475*/;
  assign r_18[40] = _9032_ | _9031_ /*15474*/;
  assign _9033_ = ~q[14] /*15473*/;
  assign _9034_ = sum_18[41] & q[14] /*15472*/;
  assign _9035_ = m_18[41] & _9033_ /*15471*/;
  assign r_18[41] = _9035_ | _9034_ /*15470*/;
  assign _9036_ = ~q[14] /*15469*/;
  assign _9037_ = sum_18[42] & q[14] /*15468*/;
  assign _9038_ = m_18[42] & _9036_ /*15467*/;
  assign r_18[42] = _9038_ | _9037_ /*15466*/;
  assign _9039_ = ~q[14] /*15465*/;
  assign _9040_ = sum_18[43] & q[14] /*15464*/;
  assign _9041_ = m_18[43] & _9039_ /*15463*/;
  assign r_18[43] = _9041_ | _9040_ /*15462*/;
  assign _9042_ = ~q[14] /*15461*/;
  assign _9043_ = sum_18[44] & q[14] /*15460*/;
  assign _9044_ = m_18[44] & _9042_ /*15459*/;
  assign r_18[44] = _9044_ | _9043_ /*15458*/;
  assign _9045_ = ~q[14] /*15457*/;
  assign _9046_ = sum_18[45] & q[14] /*15456*/;
  assign _9047_ = m_18[45] & _9045_ /*15455*/;
  assign r_18[45] = _9047_ | _9046_ /*15454*/;
  assign _9048_ = ~q[14] /*15453*/;
  assign _9049_ = sum_18[46] & q[14] /*15452*/;
  assign _9050_ = m_18[46] & _9048_ /*15451*/;
  assign r_18[46] = _9050_ | _9049_ /*15450*/;
  assign _9051_ = ~q[14] /*15449*/;
  assign _9052_ = sum_18[47] & q[14] /*15448*/;
  assign _9053_ = m_18[47] & _9051_ /*15447*/;
  assign r_18[47] = _9053_ | _9052_ /*15446*/;
  assign _9054_ = ~q[14] /*15445*/;
  assign _9055_ = sum_18[48] & q[14] /*15444*/;
  assign _9056_ = m_18[48] & _9054_ /*15443*/;
  assign r_18[48] = _9056_ | _9055_ /*15442*/;
  assign _9057_ = ~q[14] /*15441*/;
  assign _9058_ = sum_18[49] & q[14] /*15440*/;
  assign _9059_ = m_18[49] & _9057_ /*15439*/;
  assign r_18[49] = _9059_ | _9058_ /*15438*/;
  assign _9060_ = ~q[14] /*15437*/;
  assign _9061_ = sum_18[50] & q[14] /*15436*/;
  assign _9062_ = m_18[50] & _9060_ /*15435*/;
  assign r_18[50] = _9062_ | _9061_ /*15434*/;
  assign _9063_ = ~q[14] /*15433*/;
  assign _9064_ = sum_18[51] & q[14] /*15432*/;
  assign _9065_ = m_18[51] & _9063_ /*15431*/;
  assign r_18[51] = _9065_ | _9064_ /*15430*/;
  assign _9066_ = ~q[14] /*15429*/;
  assign _9067_ = sum_18[52] & q[14] /*15428*/;
  assign _9068_ = m_18[52] & _9066_ /*15427*/;
  assign r_18[52] = _9068_ | _9067_ /*15426*/;
  assign _9069_ = ~q[14] /*15425*/;
  assign _9070_ = sum_18[53] & q[14] /*15424*/;
  assign _9071_ = m_18[53] & _9069_ /*15423*/;
  assign r_18[53] = _9071_ | _9070_ /*15422*/;
  assign _9072_ = ~q[14] /*15421*/;
  assign _9073_ = sum_18[54] & q[14] /*15420*/;
  assign _9074_ = m_18[54] & _9072_ /*15419*/;
  assign r_18[54] = _9074_ | _9073_ /*15418*/;
  assign _9075_ = ~q[14] /*15417*/;
  assign _9076_ = sum_18[55] & q[14] /*15416*/;
  assign _9077_ = m_18[55] & _9075_ /*15415*/;
  assign r_18[55] = _9077_ | _9076_ /*15414*/;
  assign _9078_ = ~q[14] /*15413*/;
  assign _9079_ = sum_18[56] & q[14] /*15412*/;
  assign _9080_ = m_18[56] & _9078_ /*15411*/;
  assign r_18[56] = _9080_ | _9079_ /*15410*/;
  assign _9081_ = ~q[14] /*15409*/;
  assign _9082_ = sum_18[57] & q[14] /*15408*/;
  assign _9083_ = m_18[57] & _9081_ /*15407*/;
  assign r_18[57] = _9083_ | _9082_ /*15406*/;
  assign _9084_ = ~q[14] /*15405*/;
  assign _9085_ = sum_18[58] & q[14] /*15404*/;
  assign _9086_ = m_18[58] & _9084_ /*15403*/;
  assign r_18[58] = _9086_ | _9085_ /*15402*/;
  assign _9087_ = ~q[14] /*15401*/;
  assign _9088_ = sum_18[59] & q[14] /*15400*/;
  assign _9089_ = m_18[59] & _9087_ /*15399*/;
  assign r_18[59] = _9089_ | _9088_ /*15398*/;
  assign _9090_ = ~q[14] /*15397*/;
  assign _9091_ = sum_18[60] & q[14] /*15396*/;
  assign _9092_ = m_18[60] & _9090_ /*15395*/;
  assign r_18[60] = _9092_ | _9091_ /*15394*/;
  assign _9093_ = ~q[14] /*15393*/;
  assign _9094_ = sum_18[61] & q[14] /*15392*/;
  assign _9095_ = m_18[61] & _9093_ /*15391*/;
  assign r_18[61] = _9095_ | _9094_ /*15390*/;
  assign _9096_ = ~q[14] /*15389*/;
  assign _9097_ = sum_18[62] & q[14] /*15388*/;
  assign _9098_ = m_18[62] & _9096_ /*15387*/;
  assign r_18[62] = _9098_ | _9097_ /*15386*/;
  assign _9099_ = ~q[14] /*15385*/;
  assign _9100_ = sum_18[63] & q[14] /*15384*/;
  assign _9101_ = m_18[63] & _9099_ /*15383*/;
  assign r_18[63] = _9101_ | _9100_ /*15382*/;
  assign _9102_ = ~q[14] /*15381*/;
  assign _9103_ = sum_18[64] & q[14] /*15380*/;
  assign _9104_ = m_18[64] & _9102_ /*15379*/;
  assign r_18[64] = _9104_ | _9103_ /*15378*/;
  assign _9105_ = ~q[14] /*15377*/;
  assign _9106_ = sum_18[65] & q[14] /*15376*/;
  assign _9107_ = m_18[65] & _9105_ /*15375*/;
  assign r_18[65] = _9107_ | _9106_ /*15374*/;
  assign _9108_ = ~q[14] /*15373*/;
  assign _9109_ = sum_18[66] & q[14] /*15372*/;
  assign _9110_ = m_18[66] & _9108_ /*15371*/;
  assign r_18[66] = _9110_ | _9109_ /*15370*/;
  assign _9111_ = ~q[14] /*15369*/;
  assign _9112_ = sum_18[67] & q[14] /*15368*/;
  assign _9113_ = m_18[67] & _9111_ /*15367*/;
  assign r_18[67] = _9113_ | _9112_ /*15366*/;
  assign _9114_ = ~q[14] /*15365*/;
  assign _9115_ = sum_18[68] & q[14] /*15364*/;
  assign _9116_ = m_18[68] & _9114_ /*15363*/;
  assign r_18[68] = _9116_ | _9115_ /*15362*/;
  assign _9117_ = ~q[14] /*15361*/;
  assign _9118_ = sum_18[69] & q[14] /*15360*/;
  assign _9119_ = m_18[69] & _9117_ /*15359*/;
  assign r_18[69] = _9119_ | _9118_ /*15358*/;
  assign _9120_ = ~q[14] /*15357*/;
  assign _9121_ = sum_18[70] & q[14] /*15356*/;
  assign _9122_ = m_18[70] & _9120_ /*15355*/;
  assign r_18[70] = _9122_ | _9121_ /*15354*/;
  assign _9123_ = ~q[14] /*15353*/;
  assign _9124_ = sum_18[71] & q[14] /*15352*/;
  assign _9125_ = m_18[71] & _9123_ /*15351*/;
  assign r_18[71] = _9125_ | _9124_ /*15350*/;
  assign _9126_ = ~q[14] /*15349*/;
  assign _9127_ = sum_18[72] & q[14] /*15348*/;
  assign _9128_ = m_18[72] & _9126_ /*15347*/;
  assign r_18[72] = _9128_ | _9127_ /*15346*/;
  assign _9129_ = ~q[14] /*15345*/;
  assign _9130_ = sum_18[73] & q[14] /*15344*/;
  assign _9131_ = m_18[73] & _9129_ /*15343*/;
  assign r_18[73] = _9131_ | _9130_ /*15342*/;
  assign _9132_ = ~q[14] /*15341*/;
  assign _9133_ = sum_18[74] & q[14] /*15340*/;
  assign _9134_ = m_18[74] & _9132_ /*15339*/;
  assign r_18[74] = _9134_ | _9133_ /*15338*/;
  assign _9135_ = ~q[14] /*15337*/;
  assign _9136_ = sum_18[75] & q[14] /*15336*/;
  assign _9137_ = m_18[75] & _9135_ /*15335*/;
  assign r_18[75] = _9137_ | _9136_ /*15334*/;
  assign _9138_ = ~q[14] /*15333*/;
  assign _9139_ = sum_18[76] & q[14] /*15332*/;
  assign _9140_ = m_18[76] & _9138_ /*15331*/;
  assign r_18[76] = _9140_ | _9139_ /*15330*/;
  assign _9141_ = ~q[14] /*15329*/;
  assign _9142_ = sum_18[77] & q[14] /*15328*/;
  assign _9143_ = m_18[77] & _9141_ /*15327*/;
  assign r_18[77] = _9143_ | _9142_ /*15326*/;
  assign _9144_ = ~q[14] /*15325*/;
  assign _9145_ = sum_18[78] & q[14] /*15324*/;
  assign _9146_ = m_18[78] & _9144_ /*15323*/;
  assign r_18[78] = _9146_ | _9145_ /*15322*/;
  assign _9147_ = ~q[14] /*15321*/;
  assign _9148_ = sum_18[79] & q[14] /*15320*/;
  assign _9149_ = m_18[79] & _9147_ /*15319*/;
  assign r_18[79] = _9149_ | _9148_ /*15318*/;
  assign _9150_ = ~q[14] /*15317*/;
  assign _9151_ = sum_18[80] & q[14] /*15316*/;
  assign _9152_ = m_18[80] & _9150_ /*15315*/;
  assign r_18[80] = _9152_ | _9151_ /*15314*/;
  assign inv_19[0] = oneWire /*15128*/;
  assign inv_19[1] = oneWire /*15122*/;
  assign inv_19[2] = oneWire /*15116*/;
  assign inv_19[3] = oneWire /*15110*/;
  assign inv_19[4] = oneWire /*15104*/;
  assign inv_19[5] = oneWire /*15098*/;
  assign inv_19[6] = oneWire /*15092*/;
  assign inv_19[7] = oneWire /*15086*/;
  assign inv_19[8] = oneWire /*15080*/;
  assign inv_19[9] = oneWire /*15074*/;
  assign inv_19[10] = oneWire /*15068*/;
  assign inv_19[11] = oneWire /*15062*/;
  assign inv_19[12] = oneWire /*15056*/;
  assign inv_19[13] = ~div[0] /*15050*/;
  assign inv_19[14] = ~div[1] /*15044*/;
  assign inv_19[15] = ~div[2] /*15038*/;
  assign inv_19[16] = ~div[3] /*15032*/;
  assign inv_19[17] = ~div[4] /*15026*/;
  assign inv_19[18] = ~div[5] /*15020*/;
  assign inv_19[19] = ~div[6] /*15014*/;
  assign inv_19[20] = ~div[7] /*15008*/;
  assign inv_19[21] = ~div[8] /*15002*/;
  assign inv_19[22] = ~div[9] /*14996*/;
  assign inv_19[23] = ~div[10] /*14990*/;
  assign inv_19[24] = ~div[11] /*14984*/;
  assign inv_19[25] = ~div[12] /*14978*/;
  assign inv_19[26] = ~div[13] /*14972*/;
  assign inv_19[27] = ~div[14] /*14966*/;
  assign inv_19[28] = ~div[15] /*14960*/;
  assign inv_19[29] = ~div[16] /*14954*/;
  assign inv_19[30] = ~div[17] /*14948*/;
  assign inv_19[31] = ~div[18] /*14942*/;
  assign inv_19[32] = ~div[19] /*14936*/;
  assign inv_19[33] = ~div[20] /*14930*/;
  assign inv_19[34] = ~div[21] /*14924*/;
  assign inv_19[35] = ~div[22] /*14918*/;
  assign inv_19[36] = ~div[23] /*14912*/;
  assign inv_19[37] = ~div[24] /*14906*/;
  assign inv_19[38] = ~div[25] /*14900*/;
  assign inv_19[39] = ~div[26] /*14894*/;
  assign inv_19[40] = ~div[27] /*14888*/;
  assign inv_19[41] = ~div[28] /*14882*/;
  assign inv_19[42] = ~div[29] /*14876*/;
  assign inv_19[43] = ~div[30] /*14870*/;
  assign inv_19[44] = oneWire /*14864*/;
  assign inv_19[45] = oneWire /*14858*/;
  assign inv_19[46] = oneWire /*14852*/;
  assign inv_19[47] = oneWire /*14846*/;
  assign inv_19[48] = oneWire /*14840*/;
  assign inv_19[49] = oneWire /*14834*/;
  assign inv_19[50] = oneWire /*14828*/;
  assign inv_19[51] = oneWire /*14822*/;
  assign inv_19[52] = oneWire /*14816*/;
  assign inv_19[53] = oneWire /*14810*/;
  assign inv_19[54] = oneWire /*14804*/;
  assign inv_19[55] = oneWire /*14798*/;
  assign inv_19[56] = oneWire /*14792*/;
  assign inv_19[57] = oneWire /*14786*/;
  assign inv_19[58] = oneWire /*14780*/;
  assign inv_19[59] = oneWire /*14774*/;
  assign inv_19[60] = oneWire /*14768*/;
  assign inv_19[61] = oneWire /*14762*/;
  assign inv_19[62] = oneWire /*14756*/;
  assign inv_19[63] = oneWire /*14750*/;
  assign inv_19[64] = oneWire /*14744*/;
  assign inv_19[65] = oneWire /*14738*/;
  assign inv_19[66] = oneWire /*14732*/;
  assign inv_19[67] = oneWire /*14726*/;
  assign inv_19[68] = oneWire /*14720*/;
  assign inv_19[69] = oneWire /*14714*/;
  assign inv_19[70] = oneWire /*14708*/;
  assign inv_19[71] = oneWire /*14702*/;
  assign inv_19[72] = oneWire /*14696*/;
  assign inv_19[73] = oneWire /*14690*/;
  assign inv_19[74] = oneWire /*14684*/;
  assign inv_19[75] = oneWire /*14678*/;
  assign inv_19[76] = oneWire /*14672*/;
  assign inv_19[77] = oneWire /*14666*/;
  assign inv_19[78] = oneWire /*14660*/;
  assign inv_19[79] = oneWire /*14654*/;
  assign inv_19[80] = oneWire /*14648*/;
  assign _9153_ = inv_19[0] ^ r_18[0] /*15127*/;
  assign sum_19[0] = _9153_ ^ oneWire /*15126*/;
  assign _9154_ = _9153_ & oneWire /*15125*/;
  assign _9155_ = inv_19[0] & r_18[0] /*15124*/;
  assign _9156_ = _9154_ | _9155_ /*15123*/;
  assign _9157_ = inv_19[1] ^ r_18[1] /*15121*/;
  assign sum_19[1] = _9157_ ^ _9156_ /*15120*/;
  assign _9158_ = _9157_ & _9156_ /*15119*/;
  assign _9159_ = inv_19[1] & r_18[1] /*15118*/;
  assign _9160_ = _9158_ | _9159_ /*15117*/;
  assign _9161_ = inv_19[2] ^ r_18[2] /*15115*/;
  assign sum_19[2] = _9161_ ^ _9160_ /*15114*/;
  assign _9162_ = _9161_ & _9160_ /*15113*/;
  assign _9163_ = inv_19[2] & r_18[2] /*15112*/;
  assign _9164_ = _9162_ | _9163_ /*15111*/;
  assign _9165_ = inv_19[3] ^ r_18[3] /*15109*/;
  assign sum_19[3] = _9165_ ^ _9164_ /*15108*/;
  assign _9166_ = _9165_ & _9164_ /*15107*/;
  assign _9167_ = inv_19[3] & r_18[3] /*15106*/;
  assign _9168_ = _9166_ | _9167_ /*15105*/;
  assign _9169_ = inv_19[4] ^ r_18[4] /*15103*/;
  assign sum_19[4] = _9169_ ^ _9168_ /*15102*/;
  assign _9170_ = _9169_ & _9168_ /*15101*/;
  assign _9171_ = inv_19[4] & r_18[4] /*15100*/;
  assign _9172_ = _9170_ | _9171_ /*15099*/;
  assign _9173_ = inv_19[5] ^ r_18[5] /*15097*/;
  assign sum_19[5] = _9173_ ^ _9172_ /*15096*/;
  assign _9174_ = _9173_ & _9172_ /*15095*/;
  assign _9175_ = inv_19[5] & r_18[5] /*15094*/;
  assign _9176_ = _9174_ | _9175_ /*15093*/;
  assign _9177_ = inv_19[6] ^ r_18[6] /*15091*/;
  assign sum_19[6] = _9177_ ^ _9176_ /*15090*/;
  assign _9178_ = _9177_ & _9176_ /*15089*/;
  assign _9179_ = inv_19[6] & r_18[6] /*15088*/;
  assign _9180_ = _9178_ | _9179_ /*15087*/;
  assign _9181_ = inv_19[7] ^ r_18[7] /*15085*/;
  assign sum_19[7] = _9181_ ^ _9180_ /*15084*/;
  assign _9182_ = _9181_ & _9180_ /*15083*/;
  assign _9183_ = inv_19[7] & r_18[7] /*15082*/;
  assign _9184_ = _9182_ | _9183_ /*15081*/;
  assign _9185_ = inv_19[8] ^ r_18[8] /*15079*/;
  assign sum_19[8] = _9185_ ^ _9184_ /*15078*/;
  assign _9186_ = _9185_ & _9184_ /*15077*/;
  assign _9187_ = inv_19[8] & r_18[8] /*15076*/;
  assign _9188_ = _9186_ | _9187_ /*15075*/;
  assign _9189_ = inv_19[9] ^ r_18[9] /*15073*/;
  assign sum_19[9] = _9189_ ^ _9188_ /*15072*/;
  assign _9190_ = _9189_ & _9188_ /*15071*/;
  assign _9191_ = inv_19[9] & r_18[9] /*15070*/;
  assign _9192_ = _9190_ | _9191_ /*15069*/;
  assign _9193_ = inv_19[10] ^ r_18[10] /*15067*/;
  assign sum_19[10] = _9193_ ^ _9192_ /*15066*/;
  assign _9194_ = _9193_ & _9192_ /*15065*/;
  assign _9195_ = inv_19[10] & r_18[10] /*15064*/;
  assign _9196_ = _9194_ | _9195_ /*15063*/;
  assign _9197_ = inv_19[11] ^ r_18[11] /*15061*/;
  assign sum_19[11] = _9197_ ^ _9196_ /*15060*/;
  assign _9198_ = _9197_ & _9196_ /*15059*/;
  assign _9199_ = inv_19[11] & r_18[11] /*15058*/;
  assign _9200_ = _9198_ | _9199_ /*15057*/;
  assign _9201_ = inv_19[12] ^ r_18[12] /*15055*/;
  assign sum_19[12] = _9201_ ^ _9200_ /*15054*/;
  assign _9202_ = _9201_ & _9200_ /*15053*/;
  assign _9203_ = inv_19[12] & r_18[12] /*15052*/;
  assign _9204_ = _9202_ | _9203_ /*15051*/;
  assign _9205_ = inv_19[13] ^ r_18[13] /*15049*/;
  assign sum_19[13] = _9205_ ^ _9204_ /*15048*/;
  assign _9206_ = _9205_ & _9204_ /*15047*/;
  assign _9207_ = inv_19[13] & r_18[13] /*15046*/;
  assign _9208_ = _9206_ | _9207_ /*15045*/;
  assign _9209_ = inv_19[14] ^ r_18[14] /*15043*/;
  assign sum_19[14] = _9209_ ^ _9208_ /*15042*/;
  assign _9210_ = _9209_ & _9208_ /*15041*/;
  assign _9211_ = inv_19[14] & r_18[14] /*15040*/;
  assign _9212_ = _9210_ | _9211_ /*15039*/;
  assign _9213_ = inv_19[15] ^ r_18[15] /*15037*/;
  assign sum_19[15] = _9213_ ^ _9212_ /*15036*/;
  assign _9214_ = _9213_ & _9212_ /*15035*/;
  assign _9215_ = inv_19[15] & r_18[15] /*15034*/;
  assign _9216_ = _9214_ | _9215_ /*15033*/;
  assign _9217_ = inv_19[16] ^ r_18[16] /*15031*/;
  assign sum_19[16] = _9217_ ^ _9216_ /*15030*/;
  assign _9218_ = _9217_ & _9216_ /*15029*/;
  assign _9219_ = inv_19[16] & r_18[16] /*15028*/;
  assign _9220_ = _9218_ | _9219_ /*15027*/;
  assign _9221_ = inv_19[17] ^ r_18[17] /*15025*/;
  assign sum_19[17] = _9221_ ^ _9220_ /*15024*/;
  assign _9222_ = _9221_ & _9220_ /*15023*/;
  assign _9223_ = inv_19[17] & r_18[17] /*15022*/;
  assign _9224_ = _9222_ | _9223_ /*15021*/;
  assign _9225_ = inv_19[18] ^ r_18[18] /*15019*/;
  assign sum_19[18] = _9225_ ^ _9224_ /*15018*/;
  assign _9226_ = _9225_ & _9224_ /*15017*/;
  assign _9227_ = inv_19[18] & r_18[18] /*15016*/;
  assign _9228_ = _9226_ | _9227_ /*15015*/;
  assign _9229_ = inv_19[19] ^ r_18[19] /*15013*/;
  assign sum_19[19] = _9229_ ^ _9228_ /*15012*/;
  assign _9230_ = _9229_ & _9228_ /*15011*/;
  assign _9231_ = inv_19[19] & r_18[19] /*15010*/;
  assign _9232_ = _9230_ | _9231_ /*15009*/;
  assign _9233_ = inv_19[20] ^ r_18[20] /*15007*/;
  assign sum_19[20] = _9233_ ^ _9232_ /*15006*/;
  assign _9234_ = _9233_ & _9232_ /*15005*/;
  assign _9235_ = inv_19[20] & r_18[20] /*15004*/;
  assign _9236_ = _9234_ | _9235_ /*15003*/;
  assign _9237_ = inv_19[21] ^ r_18[21] /*15001*/;
  assign sum_19[21] = _9237_ ^ _9236_ /*15000*/;
  assign _9238_ = _9237_ & _9236_ /*14999*/;
  assign _9239_ = inv_19[21] & r_18[21] /*14998*/;
  assign _9240_ = _9238_ | _9239_ /*14997*/;
  assign _9241_ = inv_19[22] ^ r_18[22] /*14995*/;
  assign sum_19[22] = _9241_ ^ _9240_ /*14994*/;
  assign _9242_ = _9241_ & _9240_ /*14993*/;
  assign _9243_ = inv_19[22] & r_18[22] /*14992*/;
  assign _9244_ = _9242_ | _9243_ /*14991*/;
  assign _9245_ = inv_19[23] ^ r_18[23] /*14989*/;
  assign sum_19[23] = _9245_ ^ _9244_ /*14988*/;
  assign _9246_ = _9245_ & _9244_ /*14987*/;
  assign _9247_ = inv_19[23] & r_18[23] /*14986*/;
  assign _9248_ = _9246_ | _9247_ /*14985*/;
  assign _9249_ = inv_19[24] ^ r_18[24] /*14983*/;
  assign sum_19[24] = _9249_ ^ _9248_ /*14982*/;
  assign _9250_ = _9249_ & _9248_ /*14981*/;
  assign _9251_ = inv_19[24] & r_18[24] /*14980*/;
  assign _9252_ = _9250_ | _9251_ /*14979*/;
  assign _9253_ = inv_19[25] ^ r_18[25] /*14977*/;
  assign sum_19[25] = _9253_ ^ _9252_ /*14976*/;
  assign _9254_ = _9253_ & _9252_ /*14975*/;
  assign _9255_ = inv_19[25] & r_18[25] /*14974*/;
  assign _9256_ = _9254_ | _9255_ /*14973*/;
  assign _9257_ = inv_19[26] ^ r_18[26] /*14971*/;
  assign sum_19[26] = _9257_ ^ _9256_ /*14970*/;
  assign _9258_ = _9257_ & _9256_ /*14969*/;
  assign _9259_ = inv_19[26] & r_18[26] /*14968*/;
  assign _9260_ = _9258_ | _9259_ /*14967*/;
  assign _9261_ = inv_19[27] ^ r_18[27] /*14965*/;
  assign sum_19[27] = _9261_ ^ _9260_ /*14964*/;
  assign _9262_ = _9261_ & _9260_ /*14963*/;
  assign _9263_ = inv_19[27] & r_18[27] /*14962*/;
  assign _9264_ = _9262_ | _9263_ /*14961*/;
  assign _9265_ = inv_19[28] ^ r_18[28] /*14959*/;
  assign sum_19[28] = _9265_ ^ _9264_ /*14958*/;
  assign _9266_ = _9265_ & _9264_ /*14957*/;
  assign _9267_ = inv_19[28] & r_18[28] /*14956*/;
  assign _9268_ = _9266_ | _9267_ /*14955*/;
  assign _9269_ = inv_19[29] ^ r_18[29] /*14953*/;
  assign sum_19[29] = _9269_ ^ _9268_ /*14952*/;
  assign _9270_ = _9269_ & _9268_ /*14951*/;
  assign _9271_ = inv_19[29] & r_18[29] /*14950*/;
  assign _9272_ = _9270_ | _9271_ /*14949*/;
  assign _9273_ = inv_19[30] ^ r_18[30] /*14947*/;
  assign sum_19[30] = _9273_ ^ _9272_ /*14946*/;
  assign _9274_ = _9273_ & _9272_ /*14945*/;
  assign _9275_ = inv_19[30] & r_18[30] /*14944*/;
  assign _9276_ = _9274_ | _9275_ /*14943*/;
  assign _9277_ = inv_19[31] ^ r_18[31] /*14941*/;
  assign sum_19[31] = _9277_ ^ _9276_ /*14940*/;
  assign _9278_ = _9277_ & _9276_ /*14939*/;
  assign _9279_ = inv_19[31] & r_18[31] /*14938*/;
  assign _9280_ = _9278_ | _9279_ /*14937*/;
  assign _9281_ = inv_19[32] ^ r_18[32] /*14935*/;
  assign sum_19[32] = _9281_ ^ _9280_ /*14934*/;
  assign _9282_ = _9281_ & _9280_ /*14933*/;
  assign _9283_ = inv_19[32] & r_18[32] /*14932*/;
  assign _9284_ = _9282_ | _9283_ /*14931*/;
  assign _9285_ = inv_19[33] ^ r_18[33] /*14929*/;
  assign sum_19[33] = _9285_ ^ _9284_ /*14928*/;
  assign _9286_ = _9285_ & _9284_ /*14927*/;
  assign _9287_ = inv_19[33] & r_18[33] /*14926*/;
  assign _9288_ = _9286_ | _9287_ /*14925*/;
  assign _9289_ = inv_19[34] ^ r_18[34] /*14923*/;
  assign sum_19[34] = _9289_ ^ _9288_ /*14922*/;
  assign _9290_ = _9289_ & _9288_ /*14921*/;
  assign _9291_ = inv_19[34] & r_18[34] /*14920*/;
  assign _9292_ = _9290_ | _9291_ /*14919*/;
  assign _9293_ = inv_19[35] ^ r_18[35] /*14917*/;
  assign sum_19[35] = _9293_ ^ _9292_ /*14916*/;
  assign _9294_ = _9293_ & _9292_ /*14915*/;
  assign _9295_ = inv_19[35] & r_18[35] /*14914*/;
  assign _9296_ = _9294_ | _9295_ /*14913*/;
  assign _9297_ = inv_19[36] ^ r_18[36] /*14911*/;
  assign sum_19[36] = _9297_ ^ _9296_ /*14910*/;
  assign _9298_ = _9297_ & _9296_ /*14909*/;
  assign _9299_ = inv_19[36] & r_18[36] /*14908*/;
  assign _9300_ = _9298_ | _9299_ /*14907*/;
  assign _9301_ = inv_19[37] ^ r_18[37] /*14905*/;
  assign sum_19[37] = _9301_ ^ _9300_ /*14904*/;
  assign _9302_ = _9301_ & _9300_ /*14903*/;
  assign _9303_ = inv_19[37] & r_18[37] /*14902*/;
  assign _9304_ = _9302_ | _9303_ /*14901*/;
  assign _9305_ = inv_19[38] ^ r_18[38] /*14899*/;
  assign sum_19[38] = _9305_ ^ _9304_ /*14898*/;
  assign _9306_ = _9305_ & _9304_ /*14897*/;
  assign _9307_ = inv_19[38] & r_18[38] /*14896*/;
  assign _9308_ = _9306_ | _9307_ /*14895*/;
  assign _9309_ = inv_19[39] ^ r_18[39] /*14893*/;
  assign sum_19[39] = _9309_ ^ _9308_ /*14892*/;
  assign _9310_ = _9309_ & _9308_ /*14891*/;
  assign _9311_ = inv_19[39] & r_18[39] /*14890*/;
  assign _9312_ = _9310_ | _9311_ /*14889*/;
  assign _9313_ = inv_19[40] ^ r_18[40] /*14887*/;
  assign sum_19[40] = _9313_ ^ _9312_ /*14886*/;
  assign _9314_ = _9313_ & _9312_ /*14885*/;
  assign _9315_ = inv_19[40] & r_18[40] /*14884*/;
  assign _9316_ = _9314_ | _9315_ /*14883*/;
  assign _9317_ = inv_19[41] ^ r_18[41] /*14881*/;
  assign sum_19[41] = _9317_ ^ _9316_ /*14880*/;
  assign _9318_ = _9317_ & _9316_ /*14879*/;
  assign _9319_ = inv_19[41] & r_18[41] /*14878*/;
  assign _9320_ = _9318_ | _9319_ /*14877*/;
  assign _9321_ = inv_19[42] ^ r_18[42] /*14875*/;
  assign sum_19[42] = _9321_ ^ _9320_ /*14874*/;
  assign _9322_ = _9321_ & _9320_ /*14873*/;
  assign _9323_ = inv_19[42] & r_18[42] /*14872*/;
  assign _9324_ = _9322_ | _9323_ /*14871*/;
  assign _9325_ = inv_19[43] ^ r_18[43] /*14869*/;
  assign sum_19[43] = _9325_ ^ _9324_ /*14868*/;
  assign _9326_ = _9325_ & _9324_ /*14867*/;
  assign _9327_ = inv_19[43] & r_18[43] /*14866*/;
  assign _9328_ = _9326_ | _9327_ /*14865*/;
  assign _9329_ = inv_19[44] ^ r_18[44] /*14863*/;
  assign sum_19[44] = _9329_ ^ _9328_ /*14862*/;
  assign _9330_ = _9329_ & _9328_ /*14861*/;
  assign _9331_ = inv_19[44] & r_18[44] /*14860*/;
  assign _9332_ = _9330_ | _9331_ /*14859*/;
  assign _9333_ = inv_19[45] ^ r_18[45] /*14857*/;
  assign sum_19[45] = _9333_ ^ _9332_ /*14856*/;
  assign _9334_ = _9333_ & _9332_ /*14855*/;
  assign _9335_ = inv_19[45] & r_18[45] /*14854*/;
  assign _9336_ = _9334_ | _9335_ /*14853*/;
  assign _9337_ = inv_19[46] ^ r_18[46] /*14851*/;
  assign sum_19[46] = _9337_ ^ _9336_ /*14850*/;
  assign _9338_ = _9337_ & _9336_ /*14849*/;
  assign _9339_ = inv_19[46] & r_18[46] /*14848*/;
  assign _9340_ = _9338_ | _9339_ /*14847*/;
  assign _9341_ = inv_19[47] ^ r_18[47] /*14845*/;
  assign sum_19[47] = _9341_ ^ _9340_ /*14844*/;
  assign _9342_ = _9341_ & _9340_ /*14843*/;
  assign _9343_ = inv_19[47] & r_18[47] /*14842*/;
  assign _9344_ = _9342_ | _9343_ /*14841*/;
  assign _9345_ = inv_19[48] ^ r_18[48] /*14839*/;
  assign sum_19[48] = _9345_ ^ _9344_ /*14838*/;
  assign _9346_ = _9345_ & _9344_ /*14837*/;
  assign _9347_ = inv_19[48] & r_18[48] /*14836*/;
  assign _9348_ = _9346_ | _9347_ /*14835*/;
  assign _9349_ = inv_19[49] ^ r_18[49] /*14833*/;
  assign sum_19[49] = _9349_ ^ _9348_ /*14832*/;
  assign _9350_ = _9349_ & _9348_ /*14831*/;
  assign _9351_ = inv_19[49] & r_18[49] /*14830*/;
  assign _9352_ = _9350_ | _9351_ /*14829*/;
  assign _9353_ = inv_19[50] ^ r_18[50] /*14827*/;
  assign sum_19[50] = _9353_ ^ _9352_ /*14826*/;
  assign _9354_ = _9353_ & _9352_ /*14825*/;
  assign _9355_ = inv_19[50] & r_18[50] /*14824*/;
  assign _9356_ = _9354_ | _9355_ /*14823*/;
  assign _9357_ = inv_19[51] ^ r_18[51] /*14821*/;
  assign sum_19[51] = _9357_ ^ _9356_ /*14820*/;
  assign _9358_ = _9357_ & _9356_ /*14819*/;
  assign _9359_ = inv_19[51] & r_18[51] /*14818*/;
  assign _9360_ = _9358_ | _9359_ /*14817*/;
  assign _9361_ = inv_19[52] ^ r_18[52] /*14815*/;
  assign sum_19[52] = _9361_ ^ _9360_ /*14814*/;
  assign _9362_ = _9361_ & _9360_ /*14813*/;
  assign _9363_ = inv_19[52] & r_18[52] /*14812*/;
  assign _9364_ = _9362_ | _9363_ /*14811*/;
  assign _9365_ = inv_19[53] ^ r_18[53] /*14809*/;
  assign sum_19[53] = _9365_ ^ _9364_ /*14808*/;
  assign _9366_ = _9365_ & _9364_ /*14807*/;
  assign _9367_ = inv_19[53] & r_18[53] /*14806*/;
  assign _9368_ = _9366_ | _9367_ /*14805*/;
  assign _9369_ = inv_19[54] ^ r_18[54] /*14803*/;
  assign sum_19[54] = _9369_ ^ _9368_ /*14802*/;
  assign _9370_ = _9369_ & _9368_ /*14801*/;
  assign _9371_ = inv_19[54] & r_18[54] /*14800*/;
  assign _9372_ = _9370_ | _9371_ /*14799*/;
  assign _9373_ = inv_19[55] ^ r_18[55] /*14797*/;
  assign sum_19[55] = _9373_ ^ _9372_ /*14796*/;
  assign _9374_ = _9373_ & _9372_ /*14795*/;
  assign _9375_ = inv_19[55] & r_18[55] /*14794*/;
  assign _9376_ = _9374_ | _9375_ /*14793*/;
  assign _9377_ = inv_19[56] ^ r_18[56] /*14791*/;
  assign sum_19[56] = _9377_ ^ _9376_ /*14790*/;
  assign _9378_ = _9377_ & _9376_ /*14789*/;
  assign _9379_ = inv_19[56] & r_18[56] /*14788*/;
  assign _9380_ = _9378_ | _9379_ /*14787*/;
  assign _9381_ = inv_19[57] ^ r_18[57] /*14785*/;
  assign sum_19[57] = _9381_ ^ _9380_ /*14784*/;
  assign _9382_ = _9381_ & _9380_ /*14783*/;
  assign _9383_ = inv_19[57] & r_18[57] /*14782*/;
  assign _9384_ = _9382_ | _9383_ /*14781*/;
  assign _9385_ = inv_19[58] ^ r_18[58] /*14779*/;
  assign sum_19[58] = _9385_ ^ _9384_ /*14778*/;
  assign _9386_ = _9385_ & _9384_ /*14777*/;
  assign _9387_ = inv_19[58] & r_18[58] /*14776*/;
  assign _9388_ = _9386_ | _9387_ /*14775*/;
  assign _9389_ = inv_19[59] ^ r_18[59] /*14773*/;
  assign sum_19[59] = _9389_ ^ _9388_ /*14772*/;
  assign _9390_ = _9389_ & _9388_ /*14771*/;
  assign _9391_ = inv_19[59] & r_18[59] /*14770*/;
  assign _9392_ = _9390_ | _9391_ /*14769*/;
  assign _9393_ = inv_19[60] ^ r_18[60] /*14767*/;
  assign sum_19[60] = _9393_ ^ _9392_ /*14766*/;
  assign _9394_ = _9393_ & _9392_ /*14765*/;
  assign _9395_ = inv_19[60] & r_18[60] /*14764*/;
  assign _9396_ = _9394_ | _9395_ /*14763*/;
  assign _9397_ = inv_19[61] ^ r_18[61] /*14761*/;
  assign sum_19[61] = _9397_ ^ _9396_ /*14760*/;
  assign _9398_ = _9397_ & _9396_ /*14759*/;
  assign _9399_ = inv_19[61] & r_18[61] /*14758*/;
  assign _9400_ = _9398_ | _9399_ /*14757*/;
  assign _9401_ = inv_19[62] ^ r_18[62] /*14755*/;
  assign sum_19[62] = _9401_ ^ _9400_ /*14754*/;
  assign _9402_ = _9401_ & _9400_ /*14753*/;
  assign _9403_ = inv_19[62] & r_18[62] /*14752*/;
  assign _9404_ = _9402_ | _9403_ /*14751*/;
  assign _9405_ = inv_19[63] ^ r_18[63] /*14749*/;
  assign sum_19[63] = _9405_ ^ _9404_ /*14748*/;
  assign _9406_ = _9405_ & _9404_ /*14747*/;
  assign _9407_ = inv_19[63] & r_18[63] /*14746*/;
  assign _9408_ = _9406_ | _9407_ /*14745*/;
  assign _9409_ = inv_19[64] ^ r_18[64] /*14743*/;
  assign sum_19[64] = _9409_ ^ _9408_ /*14742*/;
  assign _9410_ = _9409_ & _9408_ /*14741*/;
  assign _9411_ = inv_19[64] & r_18[64] /*14740*/;
  assign _9412_ = _9410_ | _9411_ /*14739*/;
  assign _9413_ = inv_19[65] ^ r_18[65] /*14737*/;
  assign sum_19[65] = _9413_ ^ _9412_ /*14736*/;
  assign _9414_ = _9413_ & _9412_ /*14735*/;
  assign _9415_ = inv_19[65] & r_18[65] /*14734*/;
  assign _9416_ = _9414_ | _9415_ /*14733*/;
  assign _9417_ = inv_19[66] ^ r_18[66] /*14731*/;
  assign sum_19[66] = _9417_ ^ _9416_ /*14730*/;
  assign _9418_ = _9417_ & _9416_ /*14729*/;
  assign _9419_ = inv_19[66] & r_18[66] /*14728*/;
  assign _9420_ = _9418_ | _9419_ /*14727*/;
  assign _9421_ = inv_19[67] ^ r_18[67] /*14725*/;
  assign sum_19[67] = _9421_ ^ _9420_ /*14724*/;
  assign _9422_ = _9421_ & _9420_ /*14723*/;
  assign _9423_ = inv_19[67] & r_18[67] /*14722*/;
  assign _9424_ = _9422_ | _9423_ /*14721*/;
  assign _9425_ = inv_19[68] ^ r_18[68] /*14719*/;
  assign sum_19[68] = _9425_ ^ _9424_ /*14718*/;
  assign _9426_ = _9425_ & _9424_ /*14717*/;
  assign _9427_ = inv_19[68] & r_18[68] /*14716*/;
  assign _9428_ = _9426_ | _9427_ /*14715*/;
  assign _9429_ = inv_19[69] ^ r_18[69] /*14713*/;
  assign sum_19[69] = _9429_ ^ _9428_ /*14712*/;
  assign _9430_ = _9429_ & _9428_ /*14711*/;
  assign _9431_ = inv_19[69] & r_18[69] /*14710*/;
  assign _9432_ = _9430_ | _9431_ /*14709*/;
  assign _9433_ = inv_19[70] ^ r_18[70] /*14707*/;
  assign sum_19[70] = _9433_ ^ _9432_ /*14706*/;
  assign _9434_ = _9433_ & _9432_ /*14705*/;
  assign _9435_ = inv_19[70] & r_18[70] /*14704*/;
  assign _9436_ = _9434_ | _9435_ /*14703*/;
  assign _9437_ = inv_19[71] ^ r_18[71] /*14701*/;
  assign sum_19[71] = _9437_ ^ _9436_ /*14700*/;
  assign _9438_ = _9437_ & _9436_ /*14699*/;
  assign _9439_ = inv_19[71] & r_18[71] /*14698*/;
  assign _9440_ = _9438_ | _9439_ /*14697*/;
  assign _9441_ = inv_19[72] ^ r_18[72] /*14695*/;
  assign sum_19[72] = _9441_ ^ _9440_ /*14694*/;
  assign _9442_ = _9441_ & _9440_ /*14693*/;
  assign _9443_ = inv_19[72] & r_18[72] /*14692*/;
  assign _9444_ = _9442_ | _9443_ /*14691*/;
  assign _9445_ = inv_19[73] ^ r_18[73] /*14689*/;
  assign sum_19[73] = _9445_ ^ _9444_ /*14688*/;
  assign _9446_ = _9445_ & _9444_ /*14687*/;
  assign _9447_ = inv_19[73] & r_18[73] /*14686*/;
  assign _9448_ = _9446_ | _9447_ /*14685*/;
  assign _9449_ = inv_19[74] ^ r_18[74] /*14683*/;
  assign sum_19[74] = _9449_ ^ _9448_ /*14682*/;
  assign _9450_ = _9449_ & _9448_ /*14681*/;
  assign _9451_ = inv_19[74] & r_18[74] /*14680*/;
  assign _9452_ = _9450_ | _9451_ /*14679*/;
  assign _9453_ = inv_19[75] ^ r_18[75] /*14677*/;
  assign sum_19[75] = _9453_ ^ _9452_ /*14676*/;
  assign _9454_ = _9453_ & _9452_ /*14675*/;
  assign _9455_ = inv_19[75] & r_18[75] /*14674*/;
  assign _9456_ = _9454_ | _9455_ /*14673*/;
  assign _9457_ = inv_19[76] ^ r_18[76] /*14671*/;
  assign sum_19[76] = _9457_ ^ _9456_ /*14670*/;
  assign _9458_ = _9457_ & _9456_ /*14669*/;
  assign _9459_ = inv_19[76] & r_18[76] /*14668*/;
  assign _9460_ = _9458_ | _9459_ /*14667*/;
  assign _9461_ = inv_19[77] ^ r_18[77] /*14665*/;
  assign sum_19[77] = _9461_ ^ _9460_ /*14664*/;
  assign _9462_ = _9461_ & _9460_ /*14663*/;
  assign _9463_ = inv_19[77] & r_18[77] /*14662*/;
  assign _9464_ = _9462_ | _9463_ /*14661*/;
  assign _9465_ = inv_19[78] ^ r_18[78] /*14659*/;
  assign sum_19[78] = _9465_ ^ _9464_ /*14658*/;
  assign _9466_ = _9465_ & _9464_ /*14657*/;
  assign _9467_ = inv_19[78] & r_18[78] /*14656*/;
  assign _9468_ = _9466_ | _9467_ /*14655*/;
  assign _9469_ = inv_19[79] ^ r_18[79] /*14653*/;
  assign sum_19[79] = _9469_ ^ _9468_ /*14652*/;
  assign _9470_ = _9469_ & _9468_ /*14651*/;
  assign _9471_ = inv_19[79] & r_18[79] /*14650*/;
  assign _9472_ = _9470_ | _9471_ /*14649*/;
  assign _9473_ = inv_19[80] ^ r_18[80] /*14647*/;
  assign sum_19[80] = _9473_ ^ _9472_ /*14646*/;
  assign _9474_ = _9473_ & _9472_ /*14645*/;
  assign _9475_ = inv_19[80] & r_18[80] /*14644*/;
  assign _9476_ = _9474_ | _9475_ /*14643*/;
  assign _9477_ = _9476_ ^ _9472_ /*14642*/;
  assign _9478_ = ~_9477_ /*14641*/;
  assign _9479_ = sum_19[80] & _9478_ /*14640*/;
  assign _9480_ = _9477_ & _9476_ /*14639*/;
  assign sum_19[81] = _9480_ | _9479_ /*14638*/;
  assign q[13] = ~sum_19[81] /*14637*/;
  assign m_19[0] = r_18[0] /*14636*/;
  assign m_19[1] = r_18[1] /*14635*/;
  assign m_19[2] = r_18[2] /*14634*/;
  assign m_19[3] = r_18[3] /*14633*/;
  assign m_19[4] = r_18[4] /*14632*/;
  assign m_19[5] = r_18[5] /*14631*/;
  assign m_19[6] = r_18[6] /*14630*/;
  assign m_19[7] = r_18[7] /*14629*/;
  assign m_19[8] = r_18[8] /*14628*/;
  assign m_19[9] = r_18[9] /*14627*/;
  assign m_19[10] = r_18[10] /*14626*/;
  assign m_19[11] = r_18[11] /*14625*/;
  assign m_19[12] = r_18[12] /*14624*/;
  assign m_19[13] = r_18[13] /*14623*/;
  assign m_19[14] = r_18[14] /*14622*/;
  assign m_19[15] = r_18[15] /*14621*/;
  assign m_19[16] = r_18[16] /*14620*/;
  assign m_19[17] = r_18[17] /*14619*/;
  assign m_19[18] = r_18[18] /*14618*/;
  assign m_19[19] = r_18[19] /*14617*/;
  assign m_19[20] = r_18[20] /*14616*/;
  assign m_19[21] = r_18[21] /*14615*/;
  assign m_19[22] = r_18[22] /*14614*/;
  assign m_19[23] = r_18[23] /*14613*/;
  assign m_19[24] = r_18[24] /*14612*/;
  assign m_19[25] = r_18[25] /*14611*/;
  assign m_19[26] = r_18[26] /*14610*/;
  assign m_19[27] = r_18[27] /*14609*/;
  assign m_19[28] = r_18[28] /*14608*/;
  assign m_19[29] = r_18[29] /*14607*/;
  assign m_19[30] = r_18[30] /*14606*/;
  assign m_19[31] = r_18[31] /*14605*/;
  assign m_19[32] = r_18[32] /*14604*/;
  assign m_19[33] = r_18[33] /*14603*/;
  assign m_19[34] = r_18[34] /*14602*/;
  assign m_19[35] = r_18[35] /*14601*/;
  assign m_19[36] = r_18[36] /*14600*/;
  assign m_19[37] = r_18[37] /*14599*/;
  assign m_19[38] = r_18[38] /*14598*/;
  assign m_19[39] = r_18[39] /*14597*/;
  assign m_19[40] = r_18[40] /*14596*/;
  assign m_19[41] = r_18[41] /*14595*/;
  assign m_19[42] = r_18[42] /*14594*/;
  assign m_19[43] = r_18[43] /*14593*/;
  assign m_19[44] = r_18[44] /*14592*/;
  assign m_19[45] = r_18[45] /*14591*/;
  assign m_19[46] = r_18[46] /*14590*/;
  assign m_19[47] = r_18[47] /*14589*/;
  assign m_19[48] = r_18[48] /*14588*/;
  assign m_19[49] = r_18[49] /*14587*/;
  assign m_19[50] = r_18[50] /*14586*/;
  assign m_19[51] = r_18[51] /*14585*/;
  assign m_19[52] = r_18[52] /*14584*/;
  assign m_19[53] = r_18[53] /*14583*/;
  assign m_19[54] = r_18[54] /*14582*/;
  assign m_19[55] = r_18[55] /*14581*/;
  assign m_19[56] = r_18[56] /*14580*/;
  assign m_19[57] = r_18[57] /*14579*/;
  assign m_19[58] = r_18[58] /*14578*/;
  assign m_19[59] = r_18[59] /*14577*/;
  assign m_19[60] = r_18[60] /*14576*/;
  assign m_19[61] = r_18[61] /*14575*/;
  assign m_19[62] = r_18[62] /*14574*/;
  assign m_19[63] = r_18[63] /*14573*/;
  assign m_19[64] = r_18[64] /*14572*/;
  assign m_19[65] = r_18[65] /*14571*/;
  assign m_19[66] = r_18[66] /*14570*/;
  assign m_19[67] = r_18[67] /*14569*/;
  assign m_19[68] = r_18[68] /*14568*/;
  assign m_19[69] = r_18[69] /*14567*/;
  assign m_19[70] = r_18[70] /*14566*/;
  assign m_19[71] = r_18[71] /*14565*/;
  assign m_19[72] = r_18[72] /*14564*/;
  assign m_19[73] = r_18[73] /*14563*/;
  assign m_19[74] = r_18[74] /*14562*/;
  assign m_19[75] = r_18[75] /*14561*/;
  assign m_19[76] = r_18[76] /*14560*/;
  assign m_19[77] = r_18[77] /*14559*/;
  assign m_19[78] = r_18[78] /*14558*/;
  assign m_19[79] = r_18[79] /*14557*/;
  assign m_19[80] = r_18[80] /*14556*/;
  assign m_19[81] = r_18[80] /*14555*/;
  assign _9482_ = ~q[13] /*14554*/;
  assign _9483_ = sum_19[0] & q[13] /*14553*/;
  assign _9484_ = m_19[0] & _9482_ /*14552*/;
  assign r_19[0] = _9484_ | _9483_ /*14551*/;
  assign _9485_ = ~q[13] /*14550*/;
  assign _9486_ = sum_19[1] & q[13] /*14549*/;
  assign _9487_ = m_19[1] & _9485_ /*14548*/;
  assign r_19[1] = _9487_ | _9486_ /*14547*/;
  assign _9488_ = ~q[13] /*14546*/;
  assign _9489_ = sum_19[2] & q[13] /*14545*/;
  assign _9490_ = m_19[2] & _9488_ /*14544*/;
  assign r_19[2] = _9490_ | _9489_ /*14543*/;
  assign _9491_ = ~q[13] /*14542*/;
  assign _9492_ = sum_19[3] & q[13] /*14541*/;
  assign _9493_ = m_19[3] & _9491_ /*14540*/;
  assign r_19[3] = _9493_ | _9492_ /*14539*/;
  assign _9494_ = ~q[13] /*14538*/;
  assign _9495_ = sum_19[4] & q[13] /*14537*/;
  assign _9496_ = m_19[4] & _9494_ /*14536*/;
  assign r_19[4] = _9496_ | _9495_ /*14535*/;
  assign _9497_ = ~q[13] /*14534*/;
  assign _9498_ = sum_19[5] & q[13] /*14533*/;
  assign _9499_ = m_19[5] & _9497_ /*14532*/;
  assign r_19[5] = _9499_ | _9498_ /*14531*/;
  assign _9500_ = ~q[13] /*14530*/;
  assign _9501_ = sum_19[6] & q[13] /*14529*/;
  assign _9502_ = m_19[6] & _9500_ /*14528*/;
  assign r_19[6] = _9502_ | _9501_ /*14527*/;
  assign _9503_ = ~q[13] /*14526*/;
  assign _9504_ = sum_19[7] & q[13] /*14525*/;
  assign _9505_ = m_19[7] & _9503_ /*14524*/;
  assign r_19[7] = _9505_ | _9504_ /*14523*/;
  assign _9506_ = ~q[13] /*14522*/;
  assign _9507_ = sum_19[8] & q[13] /*14521*/;
  assign _9508_ = m_19[8] & _9506_ /*14520*/;
  assign r_19[8] = _9508_ | _9507_ /*14519*/;
  assign _9509_ = ~q[13] /*14518*/;
  assign _9510_ = sum_19[9] & q[13] /*14517*/;
  assign _9511_ = m_19[9] & _9509_ /*14516*/;
  assign r_19[9] = _9511_ | _9510_ /*14515*/;
  assign _9512_ = ~q[13] /*14514*/;
  assign _9513_ = sum_19[10] & q[13] /*14513*/;
  assign _9514_ = m_19[10] & _9512_ /*14512*/;
  assign r_19[10] = _9514_ | _9513_ /*14511*/;
  assign _9515_ = ~q[13] /*14510*/;
  assign _9516_ = sum_19[11] & q[13] /*14509*/;
  assign _9517_ = m_19[11] & _9515_ /*14508*/;
  assign r_19[11] = _9517_ | _9516_ /*14507*/;
  assign _9518_ = ~q[13] /*14506*/;
  assign _9519_ = sum_19[12] & q[13] /*14505*/;
  assign _9520_ = m_19[12] & _9518_ /*14504*/;
  assign r_19[12] = _9520_ | _9519_ /*14503*/;
  assign _9521_ = ~q[13] /*14502*/;
  assign _9522_ = sum_19[13] & q[13] /*14501*/;
  assign _9523_ = m_19[13] & _9521_ /*14500*/;
  assign r_19[13] = _9523_ | _9522_ /*14499*/;
  assign _9524_ = ~q[13] /*14498*/;
  assign _9525_ = sum_19[14] & q[13] /*14497*/;
  assign _9526_ = m_19[14] & _9524_ /*14496*/;
  assign r_19[14] = _9526_ | _9525_ /*14495*/;
  assign _9527_ = ~q[13] /*14494*/;
  assign _9528_ = sum_19[15] & q[13] /*14493*/;
  assign _9529_ = m_19[15] & _9527_ /*14492*/;
  assign r_19[15] = _9529_ | _9528_ /*14491*/;
  assign _9530_ = ~q[13] /*14490*/;
  assign _9531_ = sum_19[16] & q[13] /*14489*/;
  assign _9532_ = m_19[16] & _9530_ /*14488*/;
  assign r_19[16] = _9532_ | _9531_ /*14487*/;
  assign _9533_ = ~q[13] /*14486*/;
  assign _9534_ = sum_19[17] & q[13] /*14485*/;
  assign _9535_ = m_19[17] & _9533_ /*14484*/;
  assign r_19[17] = _9535_ | _9534_ /*14483*/;
  assign _9536_ = ~q[13] /*14482*/;
  assign _9537_ = sum_19[18] & q[13] /*14481*/;
  assign _9538_ = m_19[18] & _9536_ /*14480*/;
  assign r_19[18] = _9538_ | _9537_ /*14479*/;
  assign _9539_ = ~q[13] /*14478*/;
  assign _9540_ = sum_19[19] & q[13] /*14477*/;
  assign _9541_ = m_19[19] & _9539_ /*14476*/;
  assign r_19[19] = _9541_ | _9540_ /*14475*/;
  assign _9542_ = ~q[13] /*14474*/;
  assign _9543_ = sum_19[20] & q[13] /*14473*/;
  assign _9544_ = m_19[20] & _9542_ /*14472*/;
  assign r_19[20] = _9544_ | _9543_ /*14471*/;
  assign _9545_ = ~q[13] /*14470*/;
  assign _9546_ = sum_19[21] & q[13] /*14469*/;
  assign _9547_ = m_19[21] & _9545_ /*14468*/;
  assign r_19[21] = _9547_ | _9546_ /*14467*/;
  assign _9548_ = ~q[13] /*14466*/;
  assign _9549_ = sum_19[22] & q[13] /*14465*/;
  assign _9550_ = m_19[22] & _9548_ /*14464*/;
  assign r_19[22] = _9550_ | _9549_ /*14463*/;
  assign _9551_ = ~q[13] /*14462*/;
  assign _9552_ = sum_19[23] & q[13] /*14461*/;
  assign _9553_ = m_19[23] & _9551_ /*14460*/;
  assign r_19[23] = _9553_ | _9552_ /*14459*/;
  assign _9554_ = ~q[13] /*14458*/;
  assign _9555_ = sum_19[24] & q[13] /*14457*/;
  assign _9556_ = m_19[24] & _9554_ /*14456*/;
  assign r_19[24] = _9556_ | _9555_ /*14455*/;
  assign _9557_ = ~q[13] /*14454*/;
  assign _9558_ = sum_19[25] & q[13] /*14453*/;
  assign _9559_ = m_19[25] & _9557_ /*14452*/;
  assign r_19[25] = _9559_ | _9558_ /*14451*/;
  assign _9560_ = ~q[13] /*14450*/;
  assign _9561_ = sum_19[26] & q[13] /*14449*/;
  assign _9562_ = m_19[26] & _9560_ /*14448*/;
  assign r_19[26] = _9562_ | _9561_ /*14447*/;
  assign _9563_ = ~q[13] /*14446*/;
  assign _9564_ = sum_19[27] & q[13] /*14445*/;
  assign _9565_ = m_19[27] & _9563_ /*14444*/;
  assign r_19[27] = _9565_ | _9564_ /*14443*/;
  assign _9566_ = ~q[13] /*14442*/;
  assign _9567_ = sum_19[28] & q[13] /*14441*/;
  assign _9568_ = m_19[28] & _9566_ /*14440*/;
  assign r_19[28] = _9568_ | _9567_ /*14439*/;
  assign _9569_ = ~q[13] /*14438*/;
  assign _9570_ = sum_19[29] & q[13] /*14437*/;
  assign _9571_ = m_19[29] & _9569_ /*14436*/;
  assign r_19[29] = _9571_ | _9570_ /*14435*/;
  assign _9572_ = ~q[13] /*14434*/;
  assign _9573_ = sum_19[30] & q[13] /*14433*/;
  assign _9574_ = m_19[30] & _9572_ /*14432*/;
  assign r_19[30] = _9574_ | _9573_ /*14431*/;
  assign _9575_ = ~q[13] /*14430*/;
  assign _9576_ = sum_19[31] & q[13] /*14429*/;
  assign _9577_ = m_19[31] & _9575_ /*14428*/;
  assign r_19[31] = _9577_ | _9576_ /*14427*/;
  assign _9578_ = ~q[13] /*14426*/;
  assign _9579_ = sum_19[32] & q[13] /*14425*/;
  assign _9580_ = m_19[32] & _9578_ /*14424*/;
  assign r_19[32] = _9580_ | _9579_ /*14423*/;
  assign _9581_ = ~q[13] /*14422*/;
  assign _9582_ = sum_19[33] & q[13] /*14421*/;
  assign _9583_ = m_19[33] & _9581_ /*14420*/;
  assign r_19[33] = _9583_ | _9582_ /*14419*/;
  assign _9584_ = ~q[13] /*14418*/;
  assign _9585_ = sum_19[34] & q[13] /*14417*/;
  assign _9586_ = m_19[34] & _9584_ /*14416*/;
  assign r_19[34] = _9586_ | _9585_ /*14415*/;
  assign _9587_ = ~q[13] /*14414*/;
  assign _9588_ = sum_19[35] & q[13] /*14413*/;
  assign _9589_ = m_19[35] & _9587_ /*14412*/;
  assign r_19[35] = _9589_ | _9588_ /*14411*/;
  assign _9590_ = ~q[13] /*14410*/;
  assign _9591_ = sum_19[36] & q[13] /*14409*/;
  assign _9592_ = m_19[36] & _9590_ /*14408*/;
  assign r_19[36] = _9592_ | _9591_ /*14407*/;
  assign _9593_ = ~q[13] /*14406*/;
  assign _9594_ = sum_19[37] & q[13] /*14405*/;
  assign _9595_ = m_19[37] & _9593_ /*14404*/;
  assign r_19[37] = _9595_ | _9594_ /*14403*/;
  assign _9596_ = ~q[13] /*14402*/;
  assign _9597_ = sum_19[38] & q[13] /*14401*/;
  assign _9598_ = m_19[38] & _9596_ /*14400*/;
  assign r_19[38] = _9598_ | _9597_ /*14399*/;
  assign _9599_ = ~q[13] /*14398*/;
  assign _9600_ = sum_19[39] & q[13] /*14397*/;
  assign _9601_ = m_19[39] & _9599_ /*14396*/;
  assign r_19[39] = _9601_ | _9600_ /*14395*/;
  assign _9602_ = ~q[13] /*14394*/;
  assign _9603_ = sum_19[40] & q[13] /*14393*/;
  assign _9604_ = m_19[40] & _9602_ /*14392*/;
  assign r_19[40] = _9604_ | _9603_ /*14391*/;
  assign _9605_ = ~q[13] /*14390*/;
  assign _9606_ = sum_19[41] & q[13] /*14389*/;
  assign _9607_ = m_19[41] & _9605_ /*14388*/;
  assign r_19[41] = _9607_ | _9606_ /*14387*/;
  assign _9608_ = ~q[13] /*14386*/;
  assign _9609_ = sum_19[42] & q[13] /*14385*/;
  assign _9610_ = m_19[42] & _9608_ /*14384*/;
  assign r_19[42] = _9610_ | _9609_ /*14383*/;
  assign _9611_ = ~q[13] /*14382*/;
  assign _9612_ = sum_19[43] & q[13] /*14381*/;
  assign _9613_ = m_19[43] & _9611_ /*14380*/;
  assign r_19[43] = _9613_ | _9612_ /*14379*/;
  assign _9614_ = ~q[13] /*14378*/;
  assign _9615_ = sum_19[44] & q[13] /*14377*/;
  assign _9616_ = m_19[44] & _9614_ /*14376*/;
  assign r_19[44] = _9616_ | _9615_ /*14375*/;
  assign _9617_ = ~q[13] /*14374*/;
  assign _9618_ = sum_19[45] & q[13] /*14373*/;
  assign _9619_ = m_19[45] & _9617_ /*14372*/;
  assign r_19[45] = _9619_ | _9618_ /*14371*/;
  assign _9620_ = ~q[13] /*14370*/;
  assign _9621_ = sum_19[46] & q[13] /*14369*/;
  assign _9622_ = m_19[46] & _9620_ /*14368*/;
  assign r_19[46] = _9622_ | _9621_ /*14367*/;
  assign _9623_ = ~q[13] /*14366*/;
  assign _9624_ = sum_19[47] & q[13] /*14365*/;
  assign _9625_ = m_19[47] & _9623_ /*14364*/;
  assign r_19[47] = _9625_ | _9624_ /*14363*/;
  assign _9626_ = ~q[13] /*14362*/;
  assign _9627_ = sum_19[48] & q[13] /*14361*/;
  assign _9628_ = m_19[48] & _9626_ /*14360*/;
  assign r_19[48] = _9628_ | _9627_ /*14359*/;
  assign _9629_ = ~q[13] /*14358*/;
  assign _9630_ = sum_19[49] & q[13] /*14357*/;
  assign _9631_ = m_19[49] & _9629_ /*14356*/;
  assign r_19[49] = _9631_ | _9630_ /*14355*/;
  assign _9632_ = ~q[13] /*14354*/;
  assign _9633_ = sum_19[50] & q[13] /*14353*/;
  assign _9634_ = m_19[50] & _9632_ /*14352*/;
  assign r_19[50] = _9634_ | _9633_ /*14351*/;
  assign _9635_ = ~q[13] /*14350*/;
  assign _9636_ = sum_19[51] & q[13] /*14349*/;
  assign _9637_ = m_19[51] & _9635_ /*14348*/;
  assign r_19[51] = _9637_ | _9636_ /*14347*/;
  assign _9638_ = ~q[13] /*14346*/;
  assign _9639_ = sum_19[52] & q[13] /*14345*/;
  assign _9640_ = m_19[52] & _9638_ /*14344*/;
  assign r_19[52] = _9640_ | _9639_ /*14343*/;
  assign _9641_ = ~q[13] /*14342*/;
  assign _9642_ = sum_19[53] & q[13] /*14341*/;
  assign _9643_ = m_19[53] & _9641_ /*14340*/;
  assign r_19[53] = _9643_ | _9642_ /*14339*/;
  assign _9644_ = ~q[13] /*14338*/;
  assign _9645_ = sum_19[54] & q[13] /*14337*/;
  assign _9646_ = m_19[54] & _9644_ /*14336*/;
  assign r_19[54] = _9646_ | _9645_ /*14335*/;
  assign _9647_ = ~q[13] /*14334*/;
  assign _9648_ = sum_19[55] & q[13] /*14333*/;
  assign _9649_ = m_19[55] & _9647_ /*14332*/;
  assign r_19[55] = _9649_ | _9648_ /*14331*/;
  assign _9650_ = ~q[13] /*14330*/;
  assign _9651_ = sum_19[56] & q[13] /*14329*/;
  assign _9652_ = m_19[56] & _9650_ /*14328*/;
  assign r_19[56] = _9652_ | _9651_ /*14327*/;
  assign _9653_ = ~q[13] /*14326*/;
  assign _9654_ = sum_19[57] & q[13] /*14325*/;
  assign _9655_ = m_19[57] & _9653_ /*14324*/;
  assign r_19[57] = _9655_ | _9654_ /*14323*/;
  assign _9656_ = ~q[13] /*14322*/;
  assign _9657_ = sum_19[58] & q[13] /*14321*/;
  assign _9658_ = m_19[58] & _9656_ /*14320*/;
  assign r_19[58] = _9658_ | _9657_ /*14319*/;
  assign _9659_ = ~q[13] /*14318*/;
  assign _9660_ = sum_19[59] & q[13] /*14317*/;
  assign _9661_ = m_19[59] & _9659_ /*14316*/;
  assign r_19[59] = _9661_ | _9660_ /*14315*/;
  assign _9662_ = ~q[13] /*14314*/;
  assign _9663_ = sum_19[60] & q[13] /*14313*/;
  assign _9664_ = m_19[60] & _9662_ /*14312*/;
  assign r_19[60] = _9664_ | _9663_ /*14311*/;
  assign _9665_ = ~q[13] /*14310*/;
  assign _9666_ = sum_19[61] & q[13] /*14309*/;
  assign _9667_ = m_19[61] & _9665_ /*14308*/;
  assign r_19[61] = _9667_ | _9666_ /*14307*/;
  assign _9668_ = ~q[13] /*14306*/;
  assign _9669_ = sum_19[62] & q[13] /*14305*/;
  assign _9670_ = m_19[62] & _9668_ /*14304*/;
  assign r_19[62] = _9670_ | _9669_ /*14303*/;
  assign _9671_ = ~q[13] /*14302*/;
  assign _9672_ = sum_19[63] & q[13] /*14301*/;
  assign _9673_ = m_19[63] & _9671_ /*14300*/;
  assign r_19[63] = _9673_ | _9672_ /*14299*/;
  assign _9674_ = ~q[13] /*14298*/;
  assign _9675_ = sum_19[64] & q[13] /*14297*/;
  assign _9676_ = m_19[64] & _9674_ /*14296*/;
  assign r_19[64] = _9676_ | _9675_ /*14295*/;
  assign _9677_ = ~q[13] /*14294*/;
  assign _9678_ = sum_19[65] & q[13] /*14293*/;
  assign _9679_ = m_19[65] & _9677_ /*14292*/;
  assign r_19[65] = _9679_ | _9678_ /*14291*/;
  assign _9680_ = ~q[13] /*14290*/;
  assign _9681_ = sum_19[66] & q[13] /*14289*/;
  assign _9682_ = m_19[66] & _9680_ /*14288*/;
  assign r_19[66] = _9682_ | _9681_ /*14287*/;
  assign _9683_ = ~q[13] /*14286*/;
  assign _9684_ = sum_19[67] & q[13] /*14285*/;
  assign _9685_ = m_19[67] & _9683_ /*14284*/;
  assign r_19[67] = _9685_ | _9684_ /*14283*/;
  assign _9686_ = ~q[13] /*14282*/;
  assign _9687_ = sum_19[68] & q[13] /*14281*/;
  assign _9688_ = m_19[68] & _9686_ /*14280*/;
  assign r_19[68] = _9688_ | _9687_ /*14279*/;
  assign _9689_ = ~q[13] /*14278*/;
  assign _9690_ = sum_19[69] & q[13] /*14277*/;
  assign _9691_ = m_19[69] & _9689_ /*14276*/;
  assign r_19[69] = _9691_ | _9690_ /*14275*/;
  assign _9692_ = ~q[13] /*14274*/;
  assign _9693_ = sum_19[70] & q[13] /*14273*/;
  assign _9694_ = m_19[70] & _9692_ /*14272*/;
  assign r_19[70] = _9694_ | _9693_ /*14271*/;
  assign _9695_ = ~q[13] /*14270*/;
  assign _9696_ = sum_19[71] & q[13] /*14269*/;
  assign _9697_ = m_19[71] & _9695_ /*14268*/;
  assign r_19[71] = _9697_ | _9696_ /*14267*/;
  assign _9698_ = ~q[13] /*14266*/;
  assign _9699_ = sum_19[72] & q[13] /*14265*/;
  assign _9700_ = m_19[72] & _9698_ /*14264*/;
  assign r_19[72] = _9700_ | _9699_ /*14263*/;
  assign _9701_ = ~q[13] /*14262*/;
  assign _9702_ = sum_19[73] & q[13] /*14261*/;
  assign _9703_ = m_19[73] & _9701_ /*14260*/;
  assign r_19[73] = _9703_ | _9702_ /*14259*/;
  assign _9704_ = ~q[13] /*14258*/;
  assign _9705_ = sum_19[74] & q[13] /*14257*/;
  assign _9706_ = m_19[74] & _9704_ /*14256*/;
  assign r_19[74] = _9706_ | _9705_ /*14255*/;
  assign _9707_ = ~q[13] /*14254*/;
  assign _9708_ = sum_19[75] & q[13] /*14253*/;
  assign _9709_ = m_19[75] & _9707_ /*14252*/;
  assign r_19[75] = _9709_ | _9708_ /*14251*/;
  assign _9710_ = ~q[13] /*14250*/;
  assign _9711_ = sum_19[76] & q[13] /*14249*/;
  assign _9712_ = m_19[76] & _9710_ /*14248*/;
  assign r_19[76] = _9712_ | _9711_ /*14247*/;
  assign _9713_ = ~q[13] /*14246*/;
  assign _9714_ = sum_19[77] & q[13] /*14245*/;
  assign _9715_ = m_19[77] & _9713_ /*14244*/;
  assign r_19[77] = _9715_ | _9714_ /*14243*/;
  assign _9716_ = ~q[13] /*14242*/;
  assign _9717_ = sum_19[78] & q[13] /*14241*/;
  assign _9718_ = m_19[78] & _9716_ /*14240*/;
  assign r_19[78] = _9718_ | _9717_ /*14239*/;
  assign _9719_ = ~q[13] /*14238*/;
  assign _9720_ = sum_19[79] & q[13] /*14237*/;
  assign _9721_ = m_19[79] & _9719_ /*14236*/;
  assign r_19[79] = _9721_ | _9720_ /*14235*/;
  assign _9722_ = ~q[13] /*14234*/;
  assign _9723_ = sum_19[80] & q[13] /*14233*/;
  assign _9724_ = m_19[80] & _9722_ /*14232*/;
  assign r_19[80] = _9724_ | _9723_ /*14231*/;
  assign _9725_ = ~q[13] /*14230*/;
  assign _9726_ = sum_19[81] & q[13] /*14229*/;
  assign _9727_ = m_19[81] & _9725_ /*14228*/;
  assign r_19[81] = _9727_ | _9726_ /*14227*/;
  assign inv_20[0] = oneWire /*14052*/;
  assign inv_20[1] = oneWire /*14046*/;
  assign inv_20[2] = oneWire /*14040*/;
  assign inv_20[3] = oneWire /*14034*/;
  assign inv_20[4] = oneWire /*14028*/;
  assign inv_20[5] = oneWire /*14022*/;
  assign inv_20[6] = oneWire /*14016*/;
  assign inv_20[7] = oneWire /*14010*/;
  assign inv_20[8] = oneWire /*14004*/;
  assign inv_20[9] = oneWire /*13998*/;
  assign inv_20[10] = oneWire /*13992*/;
  assign inv_20[11] = oneWire /*13986*/;
  assign inv_20[12] = ~div[0] /*13980*/;
  assign inv_20[13] = ~div[1] /*13974*/;
  assign inv_20[14] = ~div[2] /*13968*/;
  assign inv_20[15] = ~div[3] /*13962*/;
  assign inv_20[16] = ~div[4] /*13956*/;
  assign inv_20[17] = ~div[5] /*13950*/;
  assign inv_20[18] = ~div[6] /*13944*/;
  assign inv_20[19] = ~div[7] /*13938*/;
  assign inv_20[20] = ~div[8] /*13932*/;
  assign inv_20[21] = ~div[9] /*13926*/;
  assign inv_20[22] = ~div[10] /*13920*/;
  assign inv_20[23] = ~div[11] /*13914*/;
  assign inv_20[24] = ~div[12] /*13908*/;
  assign inv_20[25] = ~div[13] /*13902*/;
  assign inv_20[26] = ~div[14] /*13896*/;
  assign inv_20[27] = ~div[15] /*13890*/;
  assign inv_20[28] = ~div[16] /*13884*/;
  assign inv_20[29] = ~div[17] /*13878*/;
  assign inv_20[30] = ~div[18] /*13872*/;
  assign inv_20[31] = ~div[19] /*13866*/;
  assign inv_20[32] = ~div[20] /*13860*/;
  assign inv_20[33] = ~div[21] /*13854*/;
  assign inv_20[34] = ~div[22] /*13848*/;
  assign inv_20[35] = ~div[23] /*13842*/;
  assign inv_20[36] = ~div[24] /*13836*/;
  assign inv_20[37] = ~div[25] /*13830*/;
  assign inv_20[38] = ~div[26] /*13824*/;
  assign inv_20[39] = ~div[27] /*13818*/;
  assign inv_20[40] = ~div[28] /*13812*/;
  assign inv_20[41] = ~div[29] /*13806*/;
  assign inv_20[42] = ~div[30] /*13800*/;
  assign inv_20[43] = oneWire /*13794*/;
  assign inv_20[44] = oneWire /*13788*/;
  assign inv_20[45] = oneWire /*13782*/;
  assign inv_20[46] = oneWire /*13776*/;
  assign inv_20[47] = oneWire /*13770*/;
  assign inv_20[48] = oneWire /*13764*/;
  assign inv_20[49] = oneWire /*13758*/;
  assign inv_20[50] = oneWire /*13752*/;
  assign inv_20[51] = oneWire /*13746*/;
  assign inv_20[52] = oneWire /*13740*/;
  assign inv_20[53] = oneWire /*13734*/;
  assign inv_20[54] = oneWire /*13728*/;
  assign inv_20[55] = oneWire /*13722*/;
  assign inv_20[56] = oneWire /*13716*/;
  assign inv_20[57] = oneWire /*13710*/;
  assign inv_20[58] = oneWire /*13704*/;
  assign inv_20[59] = oneWire /*13698*/;
  assign inv_20[60] = oneWire /*13692*/;
  assign inv_20[61] = oneWire /*13686*/;
  assign inv_20[62] = oneWire /*13680*/;
  assign inv_20[63] = oneWire /*13674*/;
  assign inv_20[64] = oneWire /*13668*/;
  assign inv_20[65] = oneWire /*13662*/;
  assign inv_20[66] = oneWire /*13656*/;
  assign inv_20[67] = oneWire /*13650*/;
  assign inv_20[68] = oneWire /*13644*/;
  assign inv_20[69] = oneWire /*13638*/;
  assign inv_20[70] = oneWire /*13632*/;
  assign inv_20[71] = oneWire /*13626*/;
  assign inv_20[72] = oneWire /*13620*/;
  assign inv_20[73] = oneWire /*13614*/;
  assign inv_20[74] = oneWire /*13608*/;
  assign inv_20[75] = oneWire /*13602*/;
  assign inv_20[76] = oneWire /*13596*/;
  assign inv_20[77] = oneWire /*13590*/;
  assign inv_20[78] = oneWire /*13584*/;
  assign inv_20[79] = oneWire /*13578*/;
  assign inv_20[80] = oneWire /*13572*/;
  assign inv_20[81] = oneWire /*13566*/;
  assign _9728_ = inv_20[0] ^ r_19[0] /*14051*/;
  assign sum_20[0] = _9728_ ^ oneWire /*14050*/;
  assign _9729_ = _9728_ & oneWire /*14049*/;
  assign _9730_ = inv_20[0] & r_19[0] /*14048*/;
  assign _9731_ = _9729_ | _9730_ /*14047*/;
  assign _9732_ = inv_20[1] ^ r_19[1] /*14045*/;
  assign sum_20[1] = _9732_ ^ _9731_ /*14044*/;
  assign _9733_ = _9732_ & _9731_ /*14043*/;
  assign _9734_ = inv_20[1] & r_19[1] /*14042*/;
  assign _9735_ = _9733_ | _9734_ /*14041*/;
  assign _9736_ = inv_20[2] ^ r_19[2] /*14039*/;
  assign sum_20[2] = _9736_ ^ _9735_ /*14038*/;
  assign _9737_ = _9736_ & _9735_ /*14037*/;
  assign _9738_ = inv_20[2] & r_19[2] /*14036*/;
  assign _9739_ = _9737_ | _9738_ /*14035*/;
  assign _9740_ = inv_20[3] ^ r_19[3] /*14033*/;
  assign sum_20[3] = _9740_ ^ _9739_ /*14032*/;
  assign _9741_ = _9740_ & _9739_ /*14031*/;
  assign _9742_ = inv_20[3] & r_19[3] /*14030*/;
  assign _9743_ = _9741_ | _9742_ /*14029*/;
  assign _9744_ = inv_20[4] ^ r_19[4] /*14027*/;
  assign sum_20[4] = _9744_ ^ _9743_ /*14026*/;
  assign _9745_ = _9744_ & _9743_ /*14025*/;
  assign _9746_ = inv_20[4] & r_19[4] /*14024*/;
  assign _9747_ = _9745_ | _9746_ /*14023*/;
  assign _9748_ = inv_20[5] ^ r_19[5] /*14021*/;
  assign sum_20[5] = _9748_ ^ _9747_ /*14020*/;
  assign _9749_ = _9748_ & _9747_ /*14019*/;
  assign _9750_ = inv_20[5] & r_19[5] /*14018*/;
  assign _9751_ = _9749_ | _9750_ /*14017*/;
  assign _9752_ = inv_20[6] ^ r_19[6] /*14015*/;
  assign sum_20[6] = _9752_ ^ _9751_ /*14014*/;
  assign _9753_ = _9752_ & _9751_ /*14013*/;
  assign _9754_ = inv_20[6] & r_19[6] /*14012*/;
  assign _9755_ = _9753_ | _9754_ /*14011*/;
  assign _9756_ = inv_20[7] ^ r_19[7] /*14009*/;
  assign sum_20[7] = _9756_ ^ _9755_ /*14008*/;
  assign _9757_ = _9756_ & _9755_ /*14007*/;
  assign _9758_ = inv_20[7] & r_19[7] /*14006*/;
  assign _9759_ = _9757_ | _9758_ /*14005*/;
  assign _9760_ = inv_20[8] ^ r_19[8] /*14003*/;
  assign sum_20[8] = _9760_ ^ _9759_ /*14002*/;
  assign _9761_ = _9760_ & _9759_ /*14001*/;
  assign _9762_ = inv_20[8] & r_19[8] /*14000*/;
  assign _9763_ = _9761_ | _9762_ /*13999*/;
  assign _9764_ = inv_20[9] ^ r_19[9] /*13997*/;
  assign sum_20[9] = _9764_ ^ _9763_ /*13996*/;
  assign _9765_ = _9764_ & _9763_ /*13995*/;
  assign _9766_ = inv_20[9] & r_19[9] /*13994*/;
  assign _9767_ = _9765_ | _9766_ /*13993*/;
  assign _9768_ = inv_20[10] ^ r_19[10] /*13991*/;
  assign sum_20[10] = _9768_ ^ _9767_ /*13990*/;
  assign _9769_ = _9768_ & _9767_ /*13989*/;
  assign _9770_ = inv_20[10] & r_19[10] /*13988*/;
  assign _9771_ = _9769_ | _9770_ /*13987*/;
  assign _9772_ = inv_20[11] ^ r_19[11] /*13985*/;
  assign sum_20[11] = _9772_ ^ _9771_ /*13984*/;
  assign _9773_ = _9772_ & _9771_ /*13983*/;
  assign _9774_ = inv_20[11] & r_19[11] /*13982*/;
  assign _9775_ = _9773_ | _9774_ /*13981*/;
  assign _9776_ = inv_20[12] ^ r_19[12] /*13979*/;
  assign sum_20[12] = _9776_ ^ _9775_ /*13978*/;
  assign _9777_ = _9776_ & _9775_ /*13977*/;
  assign _9778_ = inv_20[12] & r_19[12] /*13976*/;
  assign _9779_ = _9777_ | _9778_ /*13975*/;
  assign _9780_ = inv_20[13] ^ r_19[13] /*13973*/;
  assign sum_20[13] = _9780_ ^ _9779_ /*13972*/;
  assign _9781_ = _9780_ & _9779_ /*13971*/;
  assign _9782_ = inv_20[13] & r_19[13] /*13970*/;
  assign _9783_ = _9781_ | _9782_ /*13969*/;
  assign _9784_ = inv_20[14] ^ r_19[14] /*13967*/;
  assign sum_20[14] = _9784_ ^ _9783_ /*13966*/;
  assign _9785_ = _9784_ & _9783_ /*13965*/;
  assign _9786_ = inv_20[14] & r_19[14] /*13964*/;
  assign _9787_ = _9785_ | _9786_ /*13963*/;
  assign _9788_ = inv_20[15] ^ r_19[15] /*13961*/;
  assign sum_20[15] = _9788_ ^ _9787_ /*13960*/;
  assign _9789_ = _9788_ & _9787_ /*13959*/;
  assign _9790_ = inv_20[15] & r_19[15] /*13958*/;
  assign _9791_ = _9789_ | _9790_ /*13957*/;
  assign _9792_ = inv_20[16] ^ r_19[16] /*13955*/;
  assign sum_20[16] = _9792_ ^ _9791_ /*13954*/;
  assign _9793_ = _9792_ & _9791_ /*13953*/;
  assign _9794_ = inv_20[16] & r_19[16] /*13952*/;
  assign _9795_ = _9793_ | _9794_ /*13951*/;
  assign _9796_ = inv_20[17] ^ r_19[17] /*13949*/;
  assign sum_20[17] = _9796_ ^ _9795_ /*13948*/;
  assign _9797_ = _9796_ & _9795_ /*13947*/;
  assign _9798_ = inv_20[17] & r_19[17] /*13946*/;
  assign _9799_ = _9797_ | _9798_ /*13945*/;
  assign _9800_ = inv_20[18] ^ r_19[18] /*13943*/;
  assign sum_20[18] = _9800_ ^ _9799_ /*13942*/;
  assign _9801_ = _9800_ & _9799_ /*13941*/;
  assign _9802_ = inv_20[18] & r_19[18] /*13940*/;
  assign _9803_ = _9801_ | _9802_ /*13939*/;
  assign _9804_ = inv_20[19] ^ r_19[19] /*13937*/;
  assign sum_20[19] = _9804_ ^ _9803_ /*13936*/;
  assign _9805_ = _9804_ & _9803_ /*13935*/;
  assign _9806_ = inv_20[19] & r_19[19] /*13934*/;
  assign _9807_ = _9805_ | _9806_ /*13933*/;
  assign _9808_ = inv_20[20] ^ r_19[20] /*13931*/;
  assign sum_20[20] = _9808_ ^ _9807_ /*13930*/;
  assign _9809_ = _9808_ & _9807_ /*13929*/;
  assign _9810_ = inv_20[20] & r_19[20] /*13928*/;
  assign _9811_ = _9809_ | _9810_ /*13927*/;
  assign _9812_ = inv_20[21] ^ r_19[21] /*13925*/;
  assign sum_20[21] = _9812_ ^ _9811_ /*13924*/;
  assign _9813_ = _9812_ & _9811_ /*13923*/;
  assign _9814_ = inv_20[21] & r_19[21] /*13922*/;
  assign _9815_ = _9813_ | _9814_ /*13921*/;
  assign _9816_ = inv_20[22] ^ r_19[22] /*13919*/;
  assign sum_20[22] = _9816_ ^ _9815_ /*13918*/;
  assign _9817_ = _9816_ & _9815_ /*13917*/;
  assign _9818_ = inv_20[22] & r_19[22] /*13916*/;
  assign _9819_ = _9817_ | _9818_ /*13915*/;
  assign _9820_ = inv_20[23] ^ r_19[23] /*13913*/;
  assign sum_20[23] = _9820_ ^ _9819_ /*13912*/;
  assign _9821_ = _9820_ & _9819_ /*13911*/;
  assign _9822_ = inv_20[23] & r_19[23] /*13910*/;
  assign _9823_ = _9821_ | _9822_ /*13909*/;
  assign _9824_ = inv_20[24] ^ r_19[24] /*13907*/;
  assign sum_20[24] = _9824_ ^ _9823_ /*13906*/;
  assign _9825_ = _9824_ & _9823_ /*13905*/;
  assign _9826_ = inv_20[24] & r_19[24] /*13904*/;
  assign _9827_ = _9825_ | _9826_ /*13903*/;
  assign _9828_ = inv_20[25] ^ r_19[25] /*13901*/;
  assign sum_20[25] = _9828_ ^ _9827_ /*13900*/;
  assign _9829_ = _9828_ & _9827_ /*13899*/;
  assign _9830_ = inv_20[25] & r_19[25] /*13898*/;
  assign _9831_ = _9829_ | _9830_ /*13897*/;
  assign _9832_ = inv_20[26] ^ r_19[26] /*13895*/;
  assign sum_20[26] = _9832_ ^ _9831_ /*13894*/;
  assign _9833_ = _9832_ & _9831_ /*13893*/;
  assign _9834_ = inv_20[26] & r_19[26] /*13892*/;
  assign _9835_ = _9833_ | _9834_ /*13891*/;
  assign _9836_ = inv_20[27] ^ r_19[27] /*13889*/;
  assign sum_20[27] = _9836_ ^ _9835_ /*13888*/;
  assign _9837_ = _9836_ & _9835_ /*13887*/;
  assign _9838_ = inv_20[27] & r_19[27] /*13886*/;
  assign _9839_ = _9837_ | _9838_ /*13885*/;
  assign _9840_ = inv_20[28] ^ r_19[28] /*13883*/;
  assign sum_20[28] = _9840_ ^ _9839_ /*13882*/;
  assign _9841_ = _9840_ & _9839_ /*13881*/;
  assign _9842_ = inv_20[28] & r_19[28] /*13880*/;
  assign _9843_ = _9841_ | _9842_ /*13879*/;
  assign _9844_ = inv_20[29] ^ r_19[29] /*13877*/;
  assign sum_20[29] = _9844_ ^ _9843_ /*13876*/;
  assign _9845_ = _9844_ & _9843_ /*13875*/;
  assign _9846_ = inv_20[29] & r_19[29] /*13874*/;
  assign _9847_ = _9845_ | _9846_ /*13873*/;
  assign _9848_ = inv_20[30] ^ r_19[30] /*13871*/;
  assign sum_20[30] = _9848_ ^ _9847_ /*13870*/;
  assign _9849_ = _9848_ & _9847_ /*13869*/;
  assign _9850_ = inv_20[30] & r_19[30] /*13868*/;
  assign _9851_ = _9849_ | _9850_ /*13867*/;
  assign _9852_ = inv_20[31] ^ r_19[31] /*13865*/;
  assign sum_20[31] = _9852_ ^ _9851_ /*13864*/;
  assign _9853_ = _9852_ & _9851_ /*13863*/;
  assign _9854_ = inv_20[31] & r_19[31] /*13862*/;
  assign _9855_ = _9853_ | _9854_ /*13861*/;
  assign _9856_ = inv_20[32] ^ r_19[32] /*13859*/;
  assign sum_20[32] = _9856_ ^ _9855_ /*13858*/;
  assign _9857_ = _9856_ & _9855_ /*13857*/;
  assign _9858_ = inv_20[32] & r_19[32] /*13856*/;
  assign _9859_ = _9857_ | _9858_ /*13855*/;
  assign _9860_ = inv_20[33] ^ r_19[33] /*13853*/;
  assign sum_20[33] = _9860_ ^ _9859_ /*13852*/;
  assign _9861_ = _9860_ & _9859_ /*13851*/;
  assign _9862_ = inv_20[33] & r_19[33] /*13850*/;
  assign _9863_ = _9861_ | _9862_ /*13849*/;
  assign _9864_ = inv_20[34] ^ r_19[34] /*13847*/;
  assign sum_20[34] = _9864_ ^ _9863_ /*13846*/;
  assign _9865_ = _9864_ & _9863_ /*13845*/;
  assign _9866_ = inv_20[34] & r_19[34] /*13844*/;
  assign _9867_ = _9865_ | _9866_ /*13843*/;
  assign _9868_ = inv_20[35] ^ r_19[35] /*13841*/;
  assign sum_20[35] = _9868_ ^ _9867_ /*13840*/;
  assign _9869_ = _9868_ & _9867_ /*13839*/;
  assign _9870_ = inv_20[35] & r_19[35] /*13838*/;
  assign _9871_ = _9869_ | _9870_ /*13837*/;
  assign _9872_ = inv_20[36] ^ r_19[36] /*13835*/;
  assign sum_20[36] = _9872_ ^ _9871_ /*13834*/;
  assign _9873_ = _9872_ & _9871_ /*13833*/;
  assign _9874_ = inv_20[36] & r_19[36] /*13832*/;
  assign _9875_ = _9873_ | _9874_ /*13831*/;
  assign _9876_ = inv_20[37] ^ r_19[37] /*13829*/;
  assign sum_20[37] = _9876_ ^ _9875_ /*13828*/;
  assign _9877_ = _9876_ & _9875_ /*13827*/;
  assign _9878_ = inv_20[37] & r_19[37] /*13826*/;
  assign _9879_ = _9877_ | _9878_ /*13825*/;
  assign _9880_ = inv_20[38] ^ r_19[38] /*13823*/;
  assign sum_20[38] = _9880_ ^ _9879_ /*13822*/;
  assign _9881_ = _9880_ & _9879_ /*13821*/;
  assign _9882_ = inv_20[38] & r_19[38] /*13820*/;
  assign _9883_ = _9881_ | _9882_ /*13819*/;
  assign _9884_ = inv_20[39] ^ r_19[39] /*13817*/;
  assign sum_20[39] = _9884_ ^ _9883_ /*13816*/;
  assign _9885_ = _9884_ & _9883_ /*13815*/;
  assign _9886_ = inv_20[39] & r_19[39] /*13814*/;
  assign _9887_ = _9885_ | _9886_ /*13813*/;
  assign _9888_ = inv_20[40] ^ r_19[40] /*13811*/;
  assign sum_20[40] = _9888_ ^ _9887_ /*13810*/;
  assign _9889_ = _9888_ & _9887_ /*13809*/;
  assign _9890_ = inv_20[40] & r_19[40] /*13808*/;
  assign _9891_ = _9889_ | _9890_ /*13807*/;
  assign _9892_ = inv_20[41] ^ r_19[41] /*13805*/;
  assign sum_20[41] = _9892_ ^ _9891_ /*13804*/;
  assign _9893_ = _9892_ & _9891_ /*13803*/;
  assign _9894_ = inv_20[41] & r_19[41] /*13802*/;
  assign _9895_ = _9893_ | _9894_ /*13801*/;
  assign _9896_ = inv_20[42] ^ r_19[42] /*13799*/;
  assign sum_20[42] = _9896_ ^ _9895_ /*13798*/;
  assign _9897_ = _9896_ & _9895_ /*13797*/;
  assign _9898_ = inv_20[42] & r_19[42] /*13796*/;
  assign _9899_ = _9897_ | _9898_ /*13795*/;
  assign _9900_ = inv_20[43] ^ r_19[43] /*13793*/;
  assign sum_20[43] = _9900_ ^ _9899_ /*13792*/;
  assign _9901_ = _9900_ & _9899_ /*13791*/;
  assign _9902_ = inv_20[43] & r_19[43] /*13790*/;
  assign _9903_ = _9901_ | _9902_ /*13789*/;
  assign _9904_ = inv_20[44] ^ r_19[44] /*13787*/;
  assign sum_20[44] = _9904_ ^ _9903_ /*13786*/;
  assign _9905_ = _9904_ & _9903_ /*13785*/;
  assign _9906_ = inv_20[44] & r_19[44] /*13784*/;
  assign _9907_ = _9905_ | _9906_ /*13783*/;
  assign _9908_ = inv_20[45] ^ r_19[45] /*13781*/;
  assign sum_20[45] = _9908_ ^ _9907_ /*13780*/;
  assign _9909_ = _9908_ & _9907_ /*13779*/;
  assign _9910_ = inv_20[45] & r_19[45] /*13778*/;
  assign _9911_ = _9909_ | _9910_ /*13777*/;
  assign _9912_ = inv_20[46] ^ r_19[46] /*13775*/;
  assign sum_20[46] = _9912_ ^ _9911_ /*13774*/;
  assign _9913_ = _9912_ & _9911_ /*13773*/;
  assign _9914_ = inv_20[46] & r_19[46] /*13772*/;
  assign _9915_ = _9913_ | _9914_ /*13771*/;
  assign _9916_ = inv_20[47] ^ r_19[47] /*13769*/;
  assign sum_20[47] = _9916_ ^ _9915_ /*13768*/;
  assign _9917_ = _9916_ & _9915_ /*13767*/;
  assign _9918_ = inv_20[47] & r_19[47] /*13766*/;
  assign _9919_ = _9917_ | _9918_ /*13765*/;
  assign _9920_ = inv_20[48] ^ r_19[48] /*13763*/;
  assign sum_20[48] = _9920_ ^ _9919_ /*13762*/;
  assign _9921_ = _9920_ & _9919_ /*13761*/;
  assign _9922_ = inv_20[48] & r_19[48] /*13760*/;
  assign _9923_ = _9921_ | _9922_ /*13759*/;
  assign _9924_ = inv_20[49] ^ r_19[49] /*13757*/;
  assign sum_20[49] = _9924_ ^ _9923_ /*13756*/;
  assign _9925_ = _9924_ & _9923_ /*13755*/;
  assign _9926_ = inv_20[49] & r_19[49] /*13754*/;
  assign _9927_ = _9925_ | _9926_ /*13753*/;
  assign _9928_ = inv_20[50] ^ r_19[50] /*13751*/;
  assign sum_20[50] = _9928_ ^ _9927_ /*13750*/;
  assign _9929_ = _9928_ & _9927_ /*13749*/;
  assign _9930_ = inv_20[50] & r_19[50] /*13748*/;
  assign _9931_ = _9929_ | _9930_ /*13747*/;
  assign _9932_ = inv_20[51] ^ r_19[51] /*13745*/;
  assign sum_20[51] = _9932_ ^ _9931_ /*13744*/;
  assign _9933_ = _9932_ & _9931_ /*13743*/;
  assign _9934_ = inv_20[51] & r_19[51] /*13742*/;
  assign _9935_ = _9933_ | _9934_ /*13741*/;
  assign _9936_ = inv_20[52] ^ r_19[52] /*13739*/;
  assign sum_20[52] = _9936_ ^ _9935_ /*13738*/;
  assign _9937_ = _9936_ & _9935_ /*13737*/;
  assign _9938_ = inv_20[52] & r_19[52] /*13736*/;
  assign _9939_ = _9937_ | _9938_ /*13735*/;
  assign _9940_ = inv_20[53] ^ r_19[53] /*13733*/;
  assign sum_20[53] = _9940_ ^ _9939_ /*13732*/;
  assign _9941_ = _9940_ & _9939_ /*13731*/;
  assign _9942_ = inv_20[53] & r_19[53] /*13730*/;
  assign _9943_ = _9941_ | _9942_ /*13729*/;
  assign _9944_ = inv_20[54] ^ r_19[54] /*13727*/;
  assign sum_20[54] = _9944_ ^ _9943_ /*13726*/;
  assign _9945_ = _9944_ & _9943_ /*13725*/;
  assign _9946_ = inv_20[54] & r_19[54] /*13724*/;
  assign _9947_ = _9945_ | _9946_ /*13723*/;
  assign _9948_ = inv_20[55] ^ r_19[55] /*13721*/;
  assign sum_20[55] = _9948_ ^ _9947_ /*13720*/;
  assign _9949_ = _9948_ & _9947_ /*13719*/;
  assign _9950_ = inv_20[55] & r_19[55] /*13718*/;
  assign _9951_ = _9949_ | _9950_ /*13717*/;
  assign _9952_ = inv_20[56] ^ r_19[56] /*13715*/;
  assign sum_20[56] = _9952_ ^ _9951_ /*13714*/;
  assign _9953_ = _9952_ & _9951_ /*13713*/;
  assign _9954_ = inv_20[56] & r_19[56] /*13712*/;
  assign _9955_ = _9953_ | _9954_ /*13711*/;
  assign _9956_ = inv_20[57] ^ r_19[57] /*13709*/;
  assign sum_20[57] = _9956_ ^ _9955_ /*13708*/;
  assign _9957_ = _9956_ & _9955_ /*13707*/;
  assign _9958_ = inv_20[57] & r_19[57] /*13706*/;
  assign _9959_ = _9957_ | _9958_ /*13705*/;
  assign _9960_ = inv_20[58] ^ r_19[58] /*13703*/;
  assign sum_20[58] = _9960_ ^ _9959_ /*13702*/;
  assign _9961_ = _9960_ & _9959_ /*13701*/;
  assign _9962_ = inv_20[58] & r_19[58] /*13700*/;
  assign _9963_ = _9961_ | _9962_ /*13699*/;
  assign _9964_ = inv_20[59] ^ r_19[59] /*13697*/;
  assign sum_20[59] = _9964_ ^ _9963_ /*13696*/;
  assign _9965_ = _9964_ & _9963_ /*13695*/;
  assign _9966_ = inv_20[59] & r_19[59] /*13694*/;
  assign _9967_ = _9965_ | _9966_ /*13693*/;
  assign _9968_ = inv_20[60] ^ r_19[60] /*13691*/;
  assign sum_20[60] = _9968_ ^ _9967_ /*13690*/;
  assign _9969_ = _9968_ & _9967_ /*13689*/;
  assign _9970_ = inv_20[60] & r_19[60] /*13688*/;
  assign _9971_ = _9969_ | _9970_ /*13687*/;
  assign _9972_ = inv_20[61] ^ r_19[61] /*13685*/;
  assign sum_20[61] = _9972_ ^ _9971_ /*13684*/;
  assign _9973_ = _9972_ & _9971_ /*13683*/;
  assign _9974_ = inv_20[61] & r_19[61] /*13682*/;
  assign _9975_ = _9973_ | _9974_ /*13681*/;
  assign _9976_ = inv_20[62] ^ r_19[62] /*13679*/;
  assign sum_20[62] = _9976_ ^ _9975_ /*13678*/;
  assign _9977_ = _9976_ & _9975_ /*13677*/;
  assign _9978_ = inv_20[62] & r_19[62] /*13676*/;
  assign _9979_ = _9977_ | _9978_ /*13675*/;
  assign _9980_ = inv_20[63] ^ r_19[63] /*13673*/;
  assign sum_20[63] = _9980_ ^ _9979_ /*13672*/;
  assign _9981_ = _9980_ & _9979_ /*13671*/;
  assign _9982_ = inv_20[63] & r_19[63] /*13670*/;
  assign _9983_ = _9981_ | _9982_ /*13669*/;
  assign _9984_ = inv_20[64] ^ r_19[64] /*13667*/;
  assign sum_20[64] = _9984_ ^ _9983_ /*13666*/;
  assign _9985_ = _9984_ & _9983_ /*13665*/;
  assign _9986_ = inv_20[64] & r_19[64] /*13664*/;
  assign _9987_ = _9985_ | _9986_ /*13663*/;
  assign _9988_ = inv_20[65] ^ r_19[65] /*13661*/;
  assign sum_20[65] = _9988_ ^ _9987_ /*13660*/;
  assign _9989_ = _9988_ & _9987_ /*13659*/;
  assign _9990_ = inv_20[65] & r_19[65] /*13658*/;
  assign _9991_ = _9989_ | _9990_ /*13657*/;
  assign _9992_ = inv_20[66] ^ r_19[66] /*13655*/;
  assign sum_20[66] = _9992_ ^ _9991_ /*13654*/;
  assign _9993_ = _9992_ & _9991_ /*13653*/;
  assign _9994_ = inv_20[66] & r_19[66] /*13652*/;
  assign _9995_ = _9993_ | _9994_ /*13651*/;
  assign _9996_ = inv_20[67] ^ r_19[67] /*13649*/;
  assign sum_20[67] = _9996_ ^ _9995_ /*13648*/;
  assign _9997_ = _9996_ & _9995_ /*13647*/;
  assign _9998_ = inv_20[67] & r_19[67] /*13646*/;
  assign _9999_ = _9997_ | _9998_ /*13645*/;
  assign _10000_ = inv_20[68] ^ r_19[68] /*13643*/;
  assign sum_20[68] = _10000_ ^ _9999_ /*13642*/;
  assign _10001_ = _10000_ & _9999_ /*13641*/;
  assign _10002_ = inv_20[68] & r_19[68] /*13640*/;
  assign _10003_ = _10001_ | _10002_ /*13639*/;
  assign _10004_ = inv_20[69] ^ r_19[69] /*13637*/;
  assign sum_20[69] = _10004_ ^ _10003_ /*13636*/;
  assign _10005_ = _10004_ & _10003_ /*13635*/;
  assign _10006_ = inv_20[69] & r_19[69] /*13634*/;
  assign _10007_ = _10005_ | _10006_ /*13633*/;
  assign _10008_ = inv_20[70] ^ r_19[70] /*13631*/;
  assign sum_20[70] = _10008_ ^ _10007_ /*13630*/;
  assign _10009_ = _10008_ & _10007_ /*13629*/;
  assign _10010_ = inv_20[70] & r_19[70] /*13628*/;
  assign _10011_ = _10009_ | _10010_ /*13627*/;
  assign _10012_ = inv_20[71] ^ r_19[71] /*13625*/;
  assign sum_20[71] = _10012_ ^ _10011_ /*13624*/;
  assign _10013_ = _10012_ & _10011_ /*13623*/;
  assign _10014_ = inv_20[71] & r_19[71] /*13622*/;
  assign _10015_ = _10013_ | _10014_ /*13621*/;
  assign _10016_ = inv_20[72] ^ r_19[72] /*13619*/;
  assign sum_20[72] = _10016_ ^ _10015_ /*13618*/;
  assign _10017_ = _10016_ & _10015_ /*13617*/;
  assign _10018_ = inv_20[72] & r_19[72] /*13616*/;
  assign _10019_ = _10017_ | _10018_ /*13615*/;
  assign _10020_ = inv_20[73] ^ r_19[73] /*13613*/;
  assign sum_20[73] = _10020_ ^ _10019_ /*13612*/;
  assign _10021_ = _10020_ & _10019_ /*13611*/;
  assign _10022_ = inv_20[73] & r_19[73] /*13610*/;
  assign _10023_ = _10021_ | _10022_ /*13609*/;
  assign _10024_ = inv_20[74] ^ r_19[74] /*13607*/;
  assign sum_20[74] = _10024_ ^ _10023_ /*13606*/;
  assign _10025_ = _10024_ & _10023_ /*13605*/;
  assign _10026_ = inv_20[74] & r_19[74] /*13604*/;
  assign _10027_ = _10025_ | _10026_ /*13603*/;
  assign _10028_ = inv_20[75] ^ r_19[75] /*13601*/;
  assign sum_20[75] = _10028_ ^ _10027_ /*13600*/;
  assign _10029_ = _10028_ & _10027_ /*13599*/;
  assign _10030_ = inv_20[75] & r_19[75] /*13598*/;
  assign _10031_ = _10029_ | _10030_ /*13597*/;
  assign _10032_ = inv_20[76] ^ r_19[76] /*13595*/;
  assign sum_20[76] = _10032_ ^ _10031_ /*13594*/;
  assign _10033_ = _10032_ & _10031_ /*13593*/;
  assign _10034_ = inv_20[76] & r_19[76] /*13592*/;
  assign _10035_ = _10033_ | _10034_ /*13591*/;
  assign _10036_ = inv_20[77] ^ r_19[77] /*13589*/;
  assign sum_20[77] = _10036_ ^ _10035_ /*13588*/;
  assign _10037_ = _10036_ & _10035_ /*13587*/;
  assign _10038_ = inv_20[77] & r_19[77] /*13586*/;
  assign _10039_ = _10037_ | _10038_ /*13585*/;
  assign _10040_ = inv_20[78] ^ r_19[78] /*13583*/;
  assign sum_20[78] = _10040_ ^ _10039_ /*13582*/;
  assign _10041_ = _10040_ & _10039_ /*13581*/;
  assign _10042_ = inv_20[78] & r_19[78] /*13580*/;
  assign _10043_ = _10041_ | _10042_ /*13579*/;
  assign _10044_ = inv_20[79] ^ r_19[79] /*13577*/;
  assign sum_20[79] = _10044_ ^ _10043_ /*13576*/;
  assign _10045_ = _10044_ & _10043_ /*13575*/;
  assign _10046_ = inv_20[79] & r_19[79] /*13574*/;
  assign _10047_ = _10045_ | _10046_ /*13573*/;
  assign _10048_ = inv_20[80] ^ r_19[80] /*13571*/;
  assign sum_20[80] = _10048_ ^ _10047_ /*13570*/;
  assign _10049_ = _10048_ & _10047_ /*13569*/;
  assign _10050_ = inv_20[80] & r_19[80] /*13568*/;
  assign _10051_ = _10049_ | _10050_ /*13567*/;
  assign _10052_ = inv_20[81] ^ r_19[81] /*13565*/;
  assign sum_20[81] = _10052_ ^ _10051_ /*13564*/;
  assign _10053_ = _10052_ & _10051_ /*13563*/;
  assign _10054_ = inv_20[81] & r_19[81] /*13562*/;
  assign _10055_ = _10053_ | _10054_ /*13561*/;
  assign _10056_ = _10055_ ^ _10051_ /*13560*/;
  assign _10057_ = ~_10056_ /*13559*/;
  assign _10058_ = sum_20[81] & _10057_ /*13558*/;
  assign _10059_ = _10056_ & _10055_ /*13557*/;
  assign sum_20[82] = _10059_ | _10058_ /*13556*/;
  assign q[12] = ~sum_20[82] /*13555*/;
  assign m_20[0] = r_19[0] /*13554*/;
  assign m_20[1] = r_19[1] /*13553*/;
  assign m_20[2] = r_19[2] /*13552*/;
  assign m_20[3] = r_19[3] /*13551*/;
  assign m_20[4] = r_19[4] /*13550*/;
  assign m_20[5] = r_19[5] /*13549*/;
  assign m_20[6] = r_19[6] /*13548*/;
  assign m_20[7] = r_19[7] /*13547*/;
  assign m_20[8] = r_19[8] /*13546*/;
  assign m_20[9] = r_19[9] /*13545*/;
  assign m_20[10] = r_19[10] /*13544*/;
  assign m_20[11] = r_19[11] /*13543*/;
  assign m_20[12] = r_19[12] /*13542*/;
  assign m_20[13] = r_19[13] /*13541*/;
  assign m_20[14] = r_19[14] /*13540*/;
  assign m_20[15] = r_19[15] /*13539*/;
  assign m_20[16] = r_19[16] /*13538*/;
  assign m_20[17] = r_19[17] /*13537*/;
  assign m_20[18] = r_19[18] /*13536*/;
  assign m_20[19] = r_19[19] /*13535*/;
  assign m_20[20] = r_19[20] /*13534*/;
  assign m_20[21] = r_19[21] /*13533*/;
  assign m_20[22] = r_19[22] /*13532*/;
  assign m_20[23] = r_19[23] /*13531*/;
  assign m_20[24] = r_19[24] /*13530*/;
  assign m_20[25] = r_19[25] /*13529*/;
  assign m_20[26] = r_19[26] /*13528*/;
  assign m_20[27] = r_19[27] /*13527*/;
  assign m_20[28] = r_19[28] /*13526*/;
  assign m_20[29] = r_19[29] /*13525*/;
  assign m_20[30] = r_19[30] /*13524*/;
  assign m_20[31] = r_19[31] /*13523*/;
  assign m_20[32] = r_19[32] /*13522*/;
  assign m_20[33] = r_19[33] /*13521*/;
  assign m_20[34] = r_19[34] /*13520*/;
  assign m_20[35] = r_19[35] /*13519*/;
  assign m_20[36] = r_19[36] /*13518*/;
  assign m_20[37] = r_19[37] /*13517*/;
  assign m_20[38] = r_19[38] /*13516*/;
  assign m_20[39] = r_19[39] /*13515*/;
  assign m_20[40] = r_19[40] /*13514*/;
  assign m_20[41] = r_19[41] /*13513*/;
  assign m_20[42] = r_19[42] /*13512*/;
  assign m_20[43] = r_19[43] /*13511*/;
  assign m_20[44] = r_19[44] /*13510*/;
  assign m_20[45] = r_19[45] /*13509*/;
  assign m_20[46] = r_19[46] /*13508*/;
  assign m_20[47] = r_19[47] /*13507*/;
  assign m_20[48] = r_19[48] /*13506*/;
  assign m_20[49] = r_19[49] /*13505*/;
  assign m_20[50] = r_19[50] /*13504*/;
  assign m_20[51] = r_19[51] /*13503*/;
  assign m_20[52] = r_19[52] /*13502*/;
  assign m_20[53] = r_19[53] /*13501*/;
  assign m_20[54] = r_19[54] /*13500*/;
  assign m_20[55] = r_19[55] /*13499*/;
  assign m_20[56] = r_19[56] /*13498*/;
  assign m_20[57] = r_19[57] /*13497*/;
  assign m_20[58] = r_19[58] /*13496*/;
  assign m_20[59] = r_19[59] /*13495*/;
  assign m_20[60] = r_19[60] /*13494*/;
  assign m_20[61] = r_19[61] /*13493*/;
  assign m_20[62] = r_19[62] /*13492*/;
  assign m_20[63] = r_19[63] /*13491*/;
  assign m_20[64] = r_19[64] /*13490*/;
  assign m_20[65] = r_19[65] /*13489*/;
  assign m_20[66] = r_19[66] /*13488*/;
  assign m_20[67] = r_19[67] /*13487*/;
  assign m_20[68] = r_19[68] /*13486*/;
  assign m_20[69] = r_19[69] /*13485*/;
  assign m_20[70] = r_19[70] /*13484*/;
  assign m_20[71] = r_19[71] /*13483*/;
  assign m_20[72] = r_19[72] /*13482*/;
  assign m_20[73] = r_19[73] /*13481*/;
  assign m_20[74] = r_19[74] /*13480*/;
  assign m_20[75] = r_19[75] /*13479*/;
  assign m_20[76] = r_19[76] /*13478*/;
  assign m_20[77] = r_19[77] /*13477*/;
  assign m_20[78] = r_19[78] /*13476*/;
  assign m_20[79] = r_19[79] /*13475*/;
  assign m_20[80] = r_19[80] /*13474*/;
  assign m_20[81] = r_19[81] /*13473*/;
  assign m_20[82] = r_19[81] /*13472*/;
  assign _10061_ = ~q[12] /*13471*/;
  assign _10062_ = sum_20[0] & q[12] /*13470*/;
  assign _10063_ = m_20[0] & _10061_ /*13469*/;
  assign r_20[0] = _10063_ | _10062_ /*13468*/;
  assign _10064_ = ~q[12] /*13467*/;
  assign _10065_ = sum_20[1] & q[12] /*13466*/;
  assign _10066_ = m_20[1] & _10064_ /*13465*/;
  assign r_20[1] = _10066_ | _10065_ /*13464*/;
  assign _10067_ = ~q[12] /*13463*/;
  assign _10068_ = sum_20[2] & q[12] /*13462*/;
  assign _10069_ = m_20[2] & _10067_ /*13461*/;
  assign r_20[2] = _10069_ | _10068_ /*13460*/;
  assign _10070_ = ~q[12] /*13459*/;
  assign _10071_ = sum_20[3] & q[12] /*13458*/;
  assign _10072_ = m_20[3] & _10070_ /*13457*/;
  assign r_20[3] = _10072_ | _10071_ /*13456*/;
  assign _10073_ = ~q[12] /*13455*/;
  assign _10074_ = sum_20[4] & q[12] /*13454*/;
  assign _10075_ = m_20[4] & _10073_ /*13453*/;
  assign r_20[4] = _10075_ | _10074_ /*13452*/;
  assign _10076_ = ~q[12] /*13451*/;
  assign _10077_ = sum_20[5] & q[12] /*13450*/;
  assign _10078_ = m_20[5] & _10076_ /*13449*/;
  assign r_20[5] = _10078_ | _10077_ /*13448*/;
  assign _10079_ = ~q[12] /*13447*/;
  assign _10080_ = sum_20[6] & q[12] /*13446*/;
  assign _10081_ = m_20[6] & _10079_ /*13445*/;
  assign r_20[6] = _10081_ | _10080_ /*13444*/;
  assign _10082_ = ~q[12] /*13443*/;
  assign _10083_ = sum_20[7] & q[12] /*13442*/;
  assign _10084_ = m_20[7] & _10082_ /*13441*/;
  assign r_20[7] = _10084_ | _10083_ /*13440*/;
  assign _10085_ = ~q[12] /*13439*/;
  assign _10086_ = sum_20[8] & q[12] /*13438*/;
  assign _10087_ = m_20[8] & _10085_ /*13437*/;
  assign r_20[8] = _10087_ | _10086_ /*13436*/;
  assign _10088_ = ~q[12] /*13435*/;
  assign _10089_ = sum_20[9] & q[12] /*13434*/;
  assign _10090_ = m_20[9] & _10088_ /*13433*/;
  assign r_20[9] = _10090_ | _10089_ /*13432*/;
  assign _10091_ = ~q[12] /*13431*/;
  assign _10092_ = sum_20[10] & q[12] /*13430*/;
  assign _10093_ = m_20[10] & _10091_ /*13429*/;
  assign r_20[10] = _10093_ | _10092_ /*13428*/;
  assign _10094_ = ~q[12] /*13427*/;
  assign _10095_ = sum_20[11] & q[12] /*13426*/;
  assign _10096_ = m_20[11] & _10094_ /*13425*/;
  assign r_20[11] = _10096_ | _10095_ /*13424*/;
  assign _10097_ = ~q[12] /*13423*/;
  assign _10098_ = sum_20[12] & q[12] /*13422*/;
  assign _10099_ = m_20[12] & _10097_ /*13421*/;
  assign r_20[12] = _10099_ | _10098_ /*13420*/;
  assign _10100_ = ~q[12] /*13419*/;
  assign _10101_ = sum_20[13] & q[12] /*13418*/;
  assign _10102_ = m_20[13] & _10100_ /*13417*/;
  assign r_20[13] = _10102_ | _10101_ /*13416*/;
  assign _10103_ = ~q[12] /*13415*/;
  assign _10104_ = sum_20[14] & q[12] /*13414*/;
  assign _10105_ = m_20[14] & _10103_ /*13413*/;
  assign r_20[14] = _10105_ | _10104_ /*13412*/;
  assign _10106_ = ~q[12] /*13411*/;
  assign _10107_ = sum_20[15] & q[12] /*13410*/;
  assign _10108_ = m_20[15] & _10106_ /*13409*/;
  assign r_20[15] = _10108_ | _10107_ /*13408*/;
  assign _10109_ = ~q[12] /*13407*/;
  assign _10110_ = sum_20[16] & q[12] /*13406*/;
  assign _10111_ = m_20[16] & _10109_ /*13405*/;
  assign r_20[16] = _10111_ | _10110_ /*13404*/;
  assign _10112_ = ~q[12] /*13403*/;
  assign _10113_ = sum_20[17] & q[12] /*13402*/;
  assign _10114_ = m_20[17] & _10112_ /*13401*/;
  assign r_20[17] = _10114_ | _10113_ /*13400*/;
  assign _10115_ = ~q[12] /*13399*/;
  assign _10116_ = sum_20[18] & q[12] /*13398*/;
  assign _10117_ = m_20[18] & _10115_ /*13397*/;
  assign r_20[18] = _10117_ | _10116_ /*13396*/;
  assign _10118_ = ~q[12] /*13395*/;
  assign _10119_ = sum_20[19] & q[12] /*13394*/;
  assign _10120_ = m_20[19] & _10118_ /*13393*/;
  assign r_20[19] = _10120_ | _10119_ /*13392*/;
  assign _10121_ = ~q[12] /*13391*/;
  assign _10122_ = sum_20[20] & q[12] /*13390*/;
  assign _10123_ = m_20[20] & _10121_ /*13389*/;
  assign r_20[20] = _10123_ | _10122_ /*13388*/;
  assign _10124_ = ~q[12] /*13387*/;
  assign _10125_ = sum_20[21] & q[12] /*13386*/;
  assign _10126_ = m_20[21] & _10124_ /*13385*/;
  assign r_20[21] = _10126_ | _10125_ /*13384*/;
  assign _10127_ = ~q[12] /*13383*/;
  assign _10128_ = sum_20[22] & q[12] /*13382*/;
  assign _10129_ = m_20[22] & _10127_ /*13381*/;
  assign r_20[22] = _10129_ | _10128_ /*13380*/;
  assign _10130_ = ~q[12] /*13379*/;
  assign _10131_ = sum_20[23] & q[12] /*13378*/;
  assign _10132_ = m_20[23] & _10130_ /*13377*/;
  assign r_20[23] = _10132_ | _10131_ /*13376*/;
  assign _10133_ = ~q[12] /*13375*/;
  assign _10134_ = sum_20[24] & q[12] /*13374*/;
  assign _10135_ = m_20[24] & _10133_ /*13373*/;
  assign r_20[24] = _10135_ | _10134_ /*13372*/;
  assign _10136_ = ~q[12] /*13371*/;
  assign _10137_ = sum_20[25] & q[12] /*13370*/;
  assign _10138_ = m_20[25] & _10136_ /*13369*/;
  assign r_20[25] = _10138_ | _10137_ /*13368*/;
  assign _10139_ = ~q[12] /*13367*/;
  assign _10140_ = sum_20[26] & q[12] /*13366*/;
  assign _10141_ = m_20[26] & _10139_ /*13365*/;
  assign r_20[26] = _10141_ | _10140_ /*13364*/;
  assign _10142_ = ~q[12] /*13363*/;
  assign _10143_ = sum_20[27] & q[12] /*13362*/;
  assign _10144_ = m_20[27] & _10142_ /*13361*/;
  assign r_20[27] = _10144_ | _10143_ /*13360*/;
  assign _10145_ = ~q[12] /*13359*/;
  assign _10146_ = sum_20[28] & q[12] /*13358*/;
  assign _10147_ = m_20[28] & _10145_ /*13357*/;
  assign r_20[28] = _10147_ | _10146_ /*13356*/;
  assign _10148_ = ~q[12] /*13355*/;
  assign _10149_ = sum_20[29] & q[12] /*13354*/;
  assign _10150_ = m_20[29] & _10148_ /*13353*/;
  assign r_20[29] = _10150_ | _10149_ /*13352*/;
  assign _10151_ = ~q[12] /*13351*/;
  assign _10152_ = sum_20[30] & q[12] /*13350*/;
  assign _10153_ = m_20[30] & _10151_ /*13349*/;
  assign r_20[30] = _10153_ | _10152_ /*13348*/;
  assign _10154_ = ~q[12] /*13347*/;
  assign _10155_ = sum_20[31] & q[12] /*13346*/;
  assign _10156_ = m_20[31] & _10154_ /*13345*/;
  assign r_20[31] = _10156_ | _10155_ /*13344*/;
  assign _10157_ = ~q[12] /*13343*/;
  assign _10158_ = sum_20[32] & q[12] /*13342*/;
  assign _10159_ = m_20[32] & _10157_ /*13341*/;
  assign r_20[32] = _10159_ | _10158_ /*13340*/;
  assign _10160_ = ~q[12] /*13339*/;
  assign _10161_ = sum_20[33] & q[12] /*13338*/;
  assign _10162_ = m_20[33] & _10160_ /*13337*/;
  assign r_20[33] = _10162_ | _10161_ /*13336*/;
  assign _10163_ = ~q[12] /*13335*/;
  assign _10164_ = sum_20[34] & q[12] /*13334*/;
  assign _10165_ = m_20[34] & _10163_ /*13333*/;
  assign r_20[34] = _10165_ | _10164_ /*13332*/;
  assign _10166_ = ~q[12] /*13331*/;
  assign _10167_ = sum_20[35] & q[12] /*13330*/;
  assign _10168_ = m_20[35] & _10166_ /*13329*/;
  assign r_20[35] = _10168_ | _10167_ /*13328*/;
  assign _10169_ = ~q[12] /*13327*/;
  assign _10170_ = sum_20[36] & q[12] /*13326*/;
  assign _10171_ = m_20[36] & _10169_ /*13325*/;
  assign r_20[36] = _10171_ | _10170_ /*13324*/;
  assign _10172_ = ~q[12] /*13323*/;
  assign _10173_ = sum_20[37] & q[12] /*13322*/;
  assign _10174_ = m_20[37] & _10172_ /*13321*/;
  assign r_20[37] = _10174_ | _10173_ /*13320*/;
  assign _10175_ = ~q[12] /*13319*/;
  assign _10176_ = sum_20[38] & q[12] /*13318*/;
  assign _10177_ = m_20[38] & _10175_ /*13317*/;
  assign r_20[38] = _10177_ | _10176_ /*13316*/;
  assign _10178_ = ~q[12] /*13315*/;
  assign _10179_ = sum_20[39] & q[12] /*13314*/;
  assign _10180_ = m_20[39] & _10178_ /*13313*/;
  assign r_20[39] = _10180_ | _10179_ /*13312*/;
  assign _10181_ = ~q[12] /*13311*/;
  assign _10182_ = sum_20[40] & q[12] /*13310*/;
  assign _10183_ = m_20[40] & _10181_ /*13309*/;
  assign r_20[40] = _10183_ | _10182_ /*13308*/;
  assign _10184_ = ~q[12] /*13307*/;
  assign _10185_ = sum_20[41] & q[12] /*13306*/;
  assign _10186_ = m_20[41] & _10184_ /*13305*/;
  assign r_20[41] = _10186_ | _10185_ /*13304*/;
  assign _10187_ = ~q[12] /*13303*/;
  assign _10188_ = sum_20[42] & q[12] /*13302*/;
  assign _10189_ = m_20[42] & _10187_ /*13301*/;
  assign r_20[42] = _10189_ | _10188_ /*13300*/;
  assign _10190_ = ~q[12] /*13299*/;
  assign _10191_ = sum_20[43] & q[12] /*13298*/;
  assign _10192_ = m_20[43] & _10190_ /*13297*/;
  assign r_20[43] = _10192_ | _10191_ /*13296*/;
  assign _10193_ = ~q[12] /*13295*/;
  assign _10194_ = sum_20[44] & q[12] /*13294*/;
  assign _10195_ = m_20[44] & _10193_ /*13293*/;
  assign r_20[44] = _10195_ | _10194_ /*13292*/;
  assign _10196_ = ~q[12] /*13291*/;
  assign _10197_ = sum_20[45] & q[12] /*13290*/;
  assign _10198_ = m_20[45] & _10196_ /*13289*/;
  assign r_20[45] = _10198_ | _10197_ /*13288*/;
  assign _10199_ = ~q[12] /*13287*/;
  assign _10200_ = sum_20[46] & q[12] /*13286*/;
  assign _10201_ = m_20[46] & _10199_ /*13285*/;
  assign r_20[46] = _10201_ | _10200_ /*13284*/;
  assign _10202_ = ~q[12] /*13283*/;
  assign _10203_ = sum_20[47] & q[12] /*13282*/;
  assign _10204_ = m_20[47] & _10202_ /*13281*/;
  assign r_20[47] = _10204_ | _10203_ /*13280*/;
  assign _10205_ = ~q[12] /*13279*/;
  assign _10206_ = sum_20[48] & q[12] /*13278*/;
  assign _10207_ = m_20[48] & _10205_ /*13277*/;
  assign r_20[48] = _10207_ | _10206_ /*13276*/;
  assign _10208_ = ~q[12] /*13275*/;
  assign _10209_ = sum_20[49] & q[12] /*13274*/;
  assign _10210_ = m_20[49] & _10208_ /*13273*/;
  assign r_20[49] = _10210_ | _10209_ /*13272*/;
  assign _10211_ = ~q[12] /*13271*/;
  assign _10212_ = sum_20[50] & q[12] /*13270*/;
  assign _10213_ = m_20[50] & _10211_ /*13269*/;
  assign r_20[50] = _10213_ | _10212_ /*13268*/;
  assign _10214_ = ~q[12] /*13267*/;
  assign _10215_ = sum_20[51] & q[12] /*13266*/;
  assign _10216_ = m_20[51] & _10214_ /*13265*/;
  assign r_20[51] = _10216_ | _10215_ /*13264*/;
  assign _10217_ = ~q[12] /*13263*/;
  assign _10218_ = sum_20[52] & q[12] /*13262*/;
  assign _10219_ = m_20[52] & _10217_ /*13261*/;
  assign r_20[52] = _10219_ | _10218_ /*13260*/;
  assign _10220_ = ~q[12] /*13259*/;
  assign _10221_ = sum_20[53] & q[12] /*13258*/;
  assign _10222_ = m_20[53] & _10220_ /*13257*/;
  assign r_20[53] = _10222_ | _10221_ /*13256*/;
  assign _10223_ = ~q[12] /*13255*/;
  assign _10224_ = sum_20[54] & q[12] /*13254*/;
  assign _10225_ = m_20[54] & _10223_ /*13253*/;
  assign r_20[54] = _10225_ | _10224_ /*13252*/;
  assign _10226_ = ~q[12] /*13251*/;
  assign _10227_ = sum_20[55] & q[12] /*13250*/;
  assign _10228_ = m_20[55] & _10226_ /*13249*/;
  assign r_20[55] = _10228_ | _10227_ /*13248*/;
  assign _10229_ = ~q[12] /*13247*/;
  assign _10230_ = sum_20[56] & q[12] /*13246*/;
  assign _10231_ = m_20[56] & _10229_ /*13245*/;
  assign r_20[56] = _10231_ | _10230_ /*13244*/;
  assign _10232_ = ~q[12] /*13243*/;
  assign _10233_ = sum_20[57] & q[12] /*13242*/;
  assign _10234_ = m_20[57] & _10232_ /*13241*/;
  assign r_20[57] = _10234_ | _10233_ /*13240*/;
  assign _10235_ = ~q[12] /*13239*/;
  assign _10236_ = sum_20[58] & q[12] /*13238*/;
  assign _10237_ = m_20[58] & _10235_ /*13237*/;
  assign r_20[58] = _10237_ | _10236_ /*13236*/;
  assign _10238_ = ~q[12] /*13235*/;
  assign _10239_ = sum_20[59] & q[12] /*13234*/;
  assign _10240_ = m_20[59] & _10238_ /*13233*/;
  assign r_20[59] = _10240_ | _10239_ /*13232*/;
  assign _10241_ = ~q[12] /*13231*/;
  assign _10242_ = sum_20[60] & q[12] /*13230*/;
  assign _10243_ = m_20[60] & _10241_ /*13229*/;
  assign r_20[60] = _10243_ | _10242_ /*13228*/;
  assign _10244_ = ~q[12] /*13227*/;
  assign _10245_ = sum_20[61] & q[12] /*13226*/;
  assign _10246_ = m_20[61] & _10244_ /*13225*/;
  assign r_20[61] = _10246_ | _10245_ /*13224*/;
  assign _10247_ = ~q[12] /*13223*/;
  assign _10248_ = sum_20[62] & q[12] /*13222*/;
  assign _10249_ = m_20[62] & _10247_ /*13221*/;
  assign r_20[62] = _10249_ | _10248_ /*13220*/;
  assign _10250_ = ~q[12] /*13219*/;
  assign _10251_ = sum_20[63] & q[12] /*13218*/;
  assign _10252_ = m_20[63] & _10250_ /*13217*/;
  assign r_20[63] = _10252_ | _10251_ /*13216*/;
  assign _10253_ = ~q[12] /*13215*/;
  assign _10254_ = sum_20[64] & q[12] /*13214*/;
  assign _10255_ = m_20[64] & _10253_ /*13213*/;
  assign r_20[64] = _10255_ | _10254_ /*13212*/;
  assign _10256_ = ~q[12] /*13211*/;
  assign _10257_ = sum_20[65] & q[12] /*13210*/;
  assign _10258_ = m_20[65] & _10256_ /*13209*/;
  assign r_20[65] = _10258_ | _10257_ /*13208*/;
  assign _10259_ = ~q[12] /*13207*/;
  assign _10260_ = sum_20[66] & q[12] /*13206*/;
  assign _10261_ = m_20[66] & _10259_ /*13205*/;
  assign r_20[66] = _10261_ | _10260_ /*13204*/;
  assign _10262_ = ~q[12] /*13203*/;
  assign _10263_ = sum_20[67] & q[12] /*13202*/;
  assign _10264_ = m_20[67] & _10262_ /*13201*/;
  assign r_20[67] = _10264_ | _10263_ /*13200*/;
  assign _10265_ = ~q[12] /*13199*/;
  assign _10266_ = sum_20[68] & q[12] /*13198*/;
  assign _10267_ = m_20[68] & _10265_ /*13197*/;
  assign r_20[68] = _10267_ | _10266_ /*13196*/;
  assign _10268_ = ~q[12] /*13195*/;
  assign _10269_ = sum_20[69] & q[12] /*13194*/;
  assign _10270_ = m_20[69] & _10268_ /*13193*/;
  assign r_20[69] = _10270_ | _10269_ /*13192*/;
  assign _10271_ = ~q[12] /*13191*/;
  assign _10272_ = sum_20[70] & q[12] /*13190*/;
  assign _10273_ = m_20[70] & _10271_ /*13189*/;
  assign r_20[70] = _10273_ | _10272_ /*13188*/;
  assign _10274_ = ~q[12] /*13187*/;
  assign _10275_ = sum_20[71] & q[12] /*13186*/;
  assign _10276_ = m_20[71] & _10274_ /*13185*/;
  assign r_20[71] = _10276_ | _10275_ /*13184*/;
  assign _10277_ = ~q[12] /*13183*/;
  assign _10278_ = sum_20[72] & q[12] /*13182*/;
  assign _10279_ = m_20[72] & _10277_ /*13181*/;
  assign r_20[72] = _10279_ | _10278_ /*13180*/;
  assign _10280_ = ~q[12] /*13179*/;
  assign _10281_ = sum_20[73] & q[12] /*13178*/;
  assign _10282_ = m_20[73] & _10280_ /*13177*/;
  assign r_20[73] = _10282_ | _10281_ /*13176*/;
  assign _10283_ = ~q[12] /*13175*/;
  assign _10284_ = sum_20[74] & q[12] /*13174*/;
  assign _10285_ = m_20[74] & _10283_ /*13173*/;
  assign r_20[74] = _10285_ | _10284_ /*13172*/;
  assign _10286_ = ~q[12] /*13171*/;
  assign _10287_ = sum_20[75] & q[12] /*13170*/;
  assign _10288_ = m_20[75] & _10286_ /*13169*/;
  assign r_20[75] = _10288_ | _10287_ /*13168*/;
  assign _10289_ = ~q[12] /*13167*/;
  assign _10290_ = sum_20[76] & q[12] /*13166*/;
  assign _10291_ = m_20[76] & _10289_ /*13165*/;
  assign r_20[76] = _10291_ | _10290_ /*13164*/;
  assign _10292_ = ~q[12] /*13163*/;
  assign _10293_ = sum_20[77] & q[12] /*13162*/;
  assign _10294_ = m_20[77] & _10292_ /*13161*/;
  assign r_20[77] = _10294_ | _10293_ /*13160*/;
  assign _10295_ = ~q[12] /*13159*/;
  assign _10296_ = sum_20[78] & q[12] /*13158*/;
  assign _10297_ = m_20[78] & _10295_ /*13157*/;
  assign r_20[78] = _10297_ | _10296_ /*13156*/;
  assign _10298_ = ~q[12] /*13155*/;
  assign _10299_ = sum_20[79] & q[12] /*13154*/;
  assign _10300_ = m_20[79] & _10298_ /*13153*/;
  assign r_20[79] = _10300_ | _10299_ /*13152*/;
  assign _10301_ = ~q[12] /*13151*/;
  assign _10302_ = sum_20[80] & q[12] /*13150*/;
  assign _10303_ = m_20[80] & _10301_ /*13149*/;
  assign r_20[80] = _10303_ | _10302_ /*13148*/;
  assign _10304_ = ~q[12] /*13147*/;
  assign _10305_ = sum_20[81] & q[12] /*13146*/;
  assign _10306_ = m_20[81] & _10304_ /*13145*/;
  assign r_20[81] = _10306_ | _10305_ /*13144*/;
  assign _10307_ = ~q[12] /*13143*/;
  assign _10308_ = sum_20[82] & q[12] /*13142*/;
  assign _10309_ = m_20[82] & _10307_ /*13141*/;
  assign r_20[82] = _10309_ | _10308_ /*13140*/;
  assign inv_21[0] = oneWire /*12976*/;
  assign inv_21[1] = oneWire /*12970*/;
  assign inv_21[2] = oneWire /*12964*/;
  assign inv_21[3] = oneWire /*12958*/;
  assign inv_21[4] = oneWire /*12952*/;
  assign inv_21[5] = oneWire /*12946*/;
  assign inv_21[6] = oneWire /*12940*/;
  assign inv_21[7] = oneWire /*12934*/;
  assign inv_21[8] = oneWire /*12928*/;
  assign inv_21[9] = oneWire /*12922*/;
  assign inv_21[10] = oneWire /*12916*/;
  assign inv_21[11] = ~div[0] /*12910*/;
  assign inv_21[12] = ~div[1] /*12904*/;
  assign inv_21[13] = ~div[2] /*12898*/;
  assign inv_21[14] = ~div[3] /*12892*/;
  assign inv_21[15] = ~div[4] /*12886*/;
  assign inv_21[16] = ~div[5] /*12880*/;
  assign inv_21[17] = ~div[6] /*12874*/;
  assign inv_21[18] = ~div[7] /*12868*/;
  assign inv_21[19] = ~div[8] /*12862*/;
  assign inv_21[20] = ~div[9] /*12856*/;
  assign inv_21[21] = ~div[10] /*12850*/;
  assign inv_21[22] = ~div[11] /*12844*/;
  assign inv_21[23] = ~div[12] /*12838*/;
  assign inv_21[24] = ~div[13] /*12832*/;
  assign inv_21[25] = ~div[14] /*12826*/;
  assign inv_21[26] = ~div[15] /*12820*/;
  assign inv_21[27] = ~div[16] /*12814*/;
  assign inv_21[28] = ~div[17] /*12808*/;
  assign inv_21[29] = ~div[18] /*12802*/;
  assign inv_21[30] = ~div[19] /*12796*/;
  assign inv_21[31] = ~div[20] /*12790*/;
  assign inv_21[32] = ~div[21] /*12784*/;
  assign inv_21[33] = ~div[22] /*12778*/;
  assign inv_21[34] = ~div[23] /*12772*/;
  assign inv_21[35] = ~div[24] /*12766*/;
  assign inv_21[36] = ~div[25] /*12760*/;
  assign inv_21[37] = ~div[26] /*12754*/;
  assign inv_21[38] = ~div[27] /*12748*/;
  assign inv_21[39] = ~div[28] /*12742*/;
  assign inv_21[40] = ~div[29] /*12736*/;
  assign inv_21[41] = ~div[30] /*12730*/;
  assign inv_21[42] = oneWire /*12724*/;
  assign inv_21[43] = oneWire /*12718*/;
  assign inv_21[44] = oneWire /*12712*/;
  assign inv_21[45] = oneWire /*12706*/;
  assign inv_21[46] = oneWire /*12700*/;
  assign inv_21[47] = oneWire /*12694*/;
  assign inv_21[48] = oneWire /*12688*/;
  assign inv_21[49] = oneWire /*12682*/;
  assign inv_21[50] = oneWire /*12676*/;
  assign inv_21[51] = oneWire /*12670*/;
  assign inv_21[52] = oneWire /*12664*/;
  assign inv_21[53] = oneWire /*12658*/;
  assign inv_21[54] = oneWire /*12652*/;
  assign inv_21[55] = oneWire /*12646*/;
  assign inv_21[56] = oneWire /*12640*/;
  assign inv_21[57] = oneWire /*12634*/;
  assign inv_21[58] = oneWire /*12628*/;
  assign inv_21[59] = oneWire /*12622*/;
  assign inv_21[60] = oneWire /*12616*/;
  assign inv_21[61] = oneWire /*12610*/;
  assign inv_21[62] = oneWire /*12604*/;
  assign inv_21[63] = oneWire /*12598*/;
  assign inv_21[64] = oneWire /*12592*/;
  assign inv_21[65] = oneWire /*12586*/;
  assign inv_21[66] = oneWire /*12580*/;
  assign inv_21[67] = oneWire /*12574*/;
  assign inv_21[68] = oneWire /*12568*/;
  assign inv_21[69] = oneWire /*12562*/;
  assign inv_21[70] = oneWire /*12556*/;
  assign inv_21[71] = oneWire /*12550*/;
  assign inv_21[72] = oneWire /*12544*/;
  assign inv_21[73] = oneWire /*12538*/;
  assign inv_21[74] = oneWire /*12532*/;
  assign inv_21[75] = oneWire /*12526*/;
  assign inv_21[76] = oneWire /*12520*/;
  assign inv_21[77] = oneWire /*12514*/;
  assign inv_21[78] = oneWire /*12508*/;
  assign inv_21[79] = oneWire /*12502*/;
  assign inv_21[80] = oneWire /*12496*/;
  assign inv_21[81] = oneWire /*12490*/;
  assign inv_21[82] = oneWire /*12484*/;
  assign _10310_ = inv_21[0] ^ r_20[0] /*12975*/;
  assign sum_21[0] = _10310_ ^ oneWire /*12974*/;
  assign _10311_ = _10310_ & oneWire /*12973*/;
  assign _10312_ = inv_21[0] & r_20[0] /*12972*/;
  assign _10313_ = _10311_ | _10312_ /*12971*/;
  assign _10314_ = inv_21[1] ^ r_20[1] /*12969*/;
  assign sum_21[1] = _10314_ ^ _10313_ /*12968*/;
  assign _10315_ = _10314_ & _10313_ /*12967*/;
  assign _10316_ = inv_21[1] & r_20[1] /*12966*/;
  assign _10317_ = _10315_ | _10316_ /*12965*/;
  assign _10318_ = inv_21[2] ^ r_20[2] /*12963*/;
  assign sum_21[2] = _10318_ ^ _10317_ /*12962*/;
  assign _10319_ = _10318_ & _10317_ /*12961*/;
  assign _10320_ = inv_21[2] & r_20[2] /*12960*/;
  assign _10321_ = _10319_ | _10320_ /*12959*/;
  assign _10322_ = inv_21[3] ^ r_20[3] /*12957*/;
  assign sum_21[3] = _10322_ ^ _10321_ /*12956*/;
  assign _10323_ = _10322_ & _10321_ /*12955*/;
  assign _10324_ = inv_21[3] & r_20[3] /*12954*/;
  assign _10325_ = _10323_ | _10324_ /*12953*/;
  assign _10326_ = inv_21[4] ^ r_20[4] /*12951*/;
  assign sum_21[4] = _10326_ ^ _10325_ /*12950*/;
  assign _10327_ = _10326_ & _10325_ /*12949*/;
  assign _10328_ = inv_21[4] & r_20[4] /*12948*/;
  assign _10329_ = _10327_ | _10328_ /*12947*/;
  assign _10330_ = inv_21[5] ^ r_20[5] /*12945*/;
  assign sum_21[5] = _10330_ ^ _10329_ /*12944*/;
  assign _10331_ = _10330_ & _10329_ /*12943*/;
  assign _10332_ = inv_21[5] & r_20[5] /*12942*/;
  assign _10333_ = _10331_ | _10332_ /*12941*/;
  assign _10334_ = inv_21[6] ^ r_20[6] /*12939*/;
  assign sum_21[6] = _10334_ ^ _10333_ /*12938*/;
  assign _10335_ = _10334_ & _10333_ /*12937*/;
  assign _10336_ = inv_21[6] & r_20[6] /*12936*/;
  assign _10337_ = _10335_ | _10336_ /*12935*/;
  assign _10338_ = inv_21[7] ^ r_20[7] /*12933*/;
  assign sum_21[7] = _10338_ ^ _10337_ /*12932*/;
  assign _10339_ = _10338_ & _10337_ /*12931*/;
  assign _10340_ = inv_21[7] & r_20[7] /*12930*/;
  assign _10341_ = _10339_ | _10340_ /*12929*/;
  assign _10342_ = inv_21[8] ^ r_20[8] /*12927*/;
  assign sum_21[8] = _10342_ ^ _10341_ /*12926*/;
  assign _10343_ = _10342_ & _10341_ /*12925*/;
  assign _10344_ = inv_21[8] & r_20[8] /*12924*/;
  assign _10345_ = _10343_ | _10344_ /*12923*/;
  assign _10346_ = inv_21[9] ^ r_20[9] /*12921*/;
  assign sum_21[9] = _10346_ ^ _10345_ /*12920*/;
  assign _10347_ = _10346_ & _10345_ /*12919*/;
  assign _10348_ = inv_21[9] & r_20[9] /*12918*/;
  assign _10349_ = _10347_ | _10348_ /*12917*/;
  assign _10350_ = inv_21[10] ^ r_20[10] /*12915*/;
  assign sum_21[10] = _10350_ ^ _10349_ /*12914*/;
  assign _10351_ = _10350_ & _10349_ /*12913*/;
  assign _10352_ = inv_21[10] & r_20[10] /*12912*/;
  assign _10353_ = _10351_ | _10352_ /*12911*/;
  assign _10354_ = inv_21[11] ^ r_20[11] /*12909*/;
  assign sum_21[11] = _10354_ ^ _10353_ /*12908*/;
  assign _10355_ = _10354_ & _10353_ /*12907*/;
  assign _10356_ = inv_21[11] & r_20[11] /*12906*/;
  assign _10357_ = _10355_ | _10356_ /*12905*/;
  assign _10358_ = inv_21[12] ^ r_20[12] /*12903*/;
  assign sum_21[12] = _10358_ ^ _10357_ /*12902*/;
  assign _10359_ = _10358_ & _10357_ /*12901*/;
  assign _10360_ = inv_21[12] & r_20[12] /*12900*/;
  assign _10361_ = _10359_ | _10360_ /*12899*/;
  assign _10362_ = inv_21[13] ^ r_20[13] /*12897*/;
  assign sum_21[13] = _10362_ ^ _10361_ /*12896*/;
  assign _10363_ = _10362_ & _10361_ /*12895*/;
  assign _10364_ = inv_21[13] & r_20[13] /*12894*/;
  assign _10365_ = _10363_ | _10364_ /*12893*/;
  assign _10366_ = inv_21[14] ^ r_20[14] /*12891*/;
  assign sum_21[14] = _10366_ ^ _10365_ /*12890*/;
  assign _10367_ = _10366_ & _10365_ /*12889*/;
  assign _10368_ = inv_21[14] & r_20[14] /*12888*/;
  assign _10369_ = _10367_ | _10368_ /*12887*/;
  assign _10370_ = inv_21[15] ^ r_20[15] /*12885*/;
  assign sum_21[15] = _10370_ ^ _10369_ /*12884*/;
  assign _10371_ = _10370_ & _10369_ /*12883*/;
  assign _10372_ = inv_21[15] & r_20[15] /*12882*/;
  assign _10373_ = _10371_ | _10372_ /*12881*/;
  assign _10374_ = inv_21[16] ^ r_20[16] /*12879*/;
  assign sum_21[16] = _10374_ ^ _10373_ /*12878*/;
  assign _10375_ = _10374_ & _10373_ /*12877*/;
  assign _10376_ = inv_21[16] & r_20[16] /*12876*/;
  assign _10377_ = _10375_ | _10376_ /*12875*/;
  assign _10378_ = inv_21[17] ^ r_20[17] /*12873*/;
  assign sum_21[17] = _10378_ ^ _10377_ /*12872*/;
  assign _10379_ = _10378_ & _10377_ /*12871*/;
  assign _10380_ = inv_21[17] & r_20[17] /*12870*/;
  assign _10381_ = _10379_ | _10380_ /*12869*/;
  assign _10382_ = inv_21[18] ^ r_20[18] /*12867*/;
  assign sum_21[18] = _10382_ ^ _10381_ /*12866*/;
  assign _10383_ = _10382_ & _10381_ /*12865*/;
  assign _10384_ = inv_21[18] & r_20[18] /*12864*/;
  assign _10385_ = _10383_ | _10384_ /*12863*/;
  assign _10386_ = inv_21[19] ^ r_20[19] /*12861*/;
  assign sum_21[19] = _10386_ ^ _10385_ /*12860*/;
  assign _10387_ = _10386_ & _10385_ /*12859*/;
  assign _10388_ = inv_21[19] & r_20[19] /*12858*/;
  assign _10389_ = _10387_ | _10388_ /*12857*/;
  assign _10390_ = inv_21[20] ^ r_20[20] /*12855*/;
  assign sum_21[20] = _10390_ ^ _10389_ /*12854*/;
  assign _10391_ = _10390_ & _10389_ /*12853*/;
  assign _10392_ = inv_21[20] & r_20[20] /*12852*/;
  assign _10393_ = _10391_ | _10392_ /*12851*/;
  assign _10394_ = inv_21[21] ^ r_20[21] /*12849*/;
  assign sum_21[21] = _10394_ ^ _10393_ /*12848*/;
  assign _10395_ = _10394_ & _10393_ /*12847*/;
  assign _10396_ = inv_21[21] & r_20[21] /*12846*/;
  assign _10397_ = _10395_ | _10396_ /*12845*/;
  assign _10398_ = inv_21[22] ^ r_20[22] /*12843*/;
  assign sum_21[22] = _10398_ ^ _10397_ /*12842*/;
  assign _10399_ = _10398_ & _10397_ /*12841*/;
  assign _10400_ = inv_21[22] & r_20[22] /*12840*/;
  assign _10401_ = _10399_ | _10400_ /*12839*/;
  assign _10402_ = inv_21[23] ^ r_20[23] /*12837*/;
  assign sum_21[23] = _10402_ ^ _10401_ /*12836*/;
  assign _10403_ = _10402_ & _10401_ /*12835*/;
  assign _10404_ = inv_21[23] & r_20[23] /*12834*/;
  assign _10405_ = _10403_ | _10404_ /*12833*/;
  assign _10406_ = inv_21[24] ^ r_20[24] /*12831*/;
  assign sum_21[24] = _10406_ ^ _10405_ /*12830*/;
  assign _10407_ = _10406_ & _10405_ /*12829*/;
  assign _10408_ = inv_21[24] & r_20[24] /*12828*/;
  assign _10409_ = _10407_ | _10408_ /*12827*/;
  assign _10410_ = inv_21[25] ^ r_20[25] /*12825*/;
  assign sum_21[25] = _10410_ ^ _10409_ /*12824*/;
  assign _10411_ = _10410_ & _10409_ /*12823*/;
  assign _10412_ = inv_21[25] & r_20[25] /*12822*/;
  assign _10413_ = _10411_ | _10412_ /*12821*/;
  assign _10414_ = inv_21[26] ^ r_20[26] /*12819*/;
  assign sum_21[26] = _10414_ ^ _10413_ /*12818*/;
  assign _10415_ = _10414_ & _10413_ /*12817*/;
  assign _10416_ = inv_21[26] & r_20[26] /*12816*/;
  assign _10417_ = _10415_ | _10416_ /*12815*/;
  assign _10418_ = inv_21[27] ^ r_20[27] /*12813*/;
  assign sum_21[27] = _10418_ ^ _10417_ /*12812*/;
  assign _10419_ = _10418_ & _10417_ /*12811*/;
  assign _10420_ = inv_21[27] & r_20[27] /*12810*/;
  assign _10421_ = _10419_ | _10420_ /*12809*/;
  assign _10422_ = inv_21[28] ^ r_20[28] /*12807*/;
  assign sum_21[28] = _10422_ ^ _10421_ /*12806*/;
  assign _10423_ = _10422_ & _10421_ /*12805*/;
  assign _10424_ = inv_21[28] & r_20[28] /*12804*/;
  assign _10425_ = _10423_ | _10424_ /*12803*/;
  assign _10426_ = inv_21[29] ^ r_20[29] /*12801*/;
  assign sum_21[29] = _10426_ ^ _10425_ /*12800*/;
  assign _10427_ = _10426_ & _10425_ /*12799*/;
  assign _10428_ = inv_21[29] & r_20[29] /*12798*/;
  assign _10429_ = _10427_ | _10428_ /*12797*/;
  assign _10430_ = inv_21[30] ^ r_20[30] /*12795*/;
  assign sum_21[30] = _10430_ ^ _10429_ /*12794*/;
  assign _10431_ = _10430_ & _10429_ /*12793*/;
  assign _10432_ = inv_21[30] & r_20[30] /*12792*/;
  assign _10433_ = _10431_ | _10432_ /*12791*/;
  assign _10434_ = inv_21[31] ^ r_20[31] /*12789*/;
  assign sum_21[31] = _10434_ ^ _10433_ /*12788*/;
  assign _10435_ = _10434_ & _10433_ /*12787*/;
  assign _10436_ = inv_21[31] & r_20[31] /*12786*/;
  assign _10437_ = _10435_ | _10436_ /*12785*/;
  assign _10438_ = inv_21[32] ^ r_20[32] /*12783*/;
  assign sum_21[32] = _10438_ ^ _10437_ /*12782*/;
  assign _10439_ = _10438_ & _10437_ /*12781*/;
  assign _10440_ = inv_21[32] & r_20[32] /*12780*/;
  assign _10441_ = _10439_ | _10440_ /*12779*/;
  assign _10442_ = inv_21[33] ^ r_20[33] /*12777*/;
  assign sum_21[33] = _10442_ ^ _10441_ /*12776*/;
  assign _10443_ = _10442_ & _10441_ /*12775*/;
  assign _10444_ = inv_21[33] & r_20[33] /*12774*/;
  assign _10445_ = _10443_ | _10444_ /*12773*/;
  assign _10446_ = inv_21[34] ^ r_20[34] /*12771*/;
  assign sum_21[34] = _10446_ ^ _10445_ /*12770*/;
  assign _10447_ = _10446_ & _10445_ /*12769*/;
  assign _10448_ = inv_21[34] & r_20[34] /*12768*/;
  assign _10449_ = _10447_ | _10448_ /*12767*/;
  assign _10450_ = inv_21[35] ^ r_20[35] /*12765*/;
  assign sum_21[35] = _10450_ ^ _10449_ /*12764*/;
  assign _10451_ = _10450_ & _10449_ /*12763*/;
  assign _10452_ = inv_21[35] & r_20[35] /*12762*/;
  assign _10453_ = _10451_ | _10452_ /*12761*/;
  assign _10454_ = inv_21[36] ^ r_20[36] /*12759*/;
  assign sum_21[36] = _10454_ ^ _10453_ /*12758*/;
  assign _10455_ = _10454_ & _10453_ /*12757*/;
  assign _10456_ = inv_21[36] & r_20[36] /*12756*/;
  assign _10457_ = _10455_ | _10456_ /*12755*/;
  assign _10458_ = inv_21[37] ^ r_20[37] /*12753*/;
  assign sum_21[37] = _10458_ ^ _10457_ /*12752*/;
  assign _10459_ = _10458_ & _10457_ /*12751*/;
  assign _10460_ = inv_21[37] & r_20[37] /*12750*/;
  assign _10461_ = _10459_ | _10460_ /*12749*/;
  assign _10462_ = inv_21[38] ^ r_20[38] /*12747*/;
  assign sum_21[38] = _10462_ ^ _10461_ /*12746*/;
  assign _10463_ = _10462_ & _10461_ /*12745*/;
  assign _10464_ = inv_21[38] & r_20[38] /*12744*/;
  assign _10465_ = _10463_ | _10464_ /*12743*/;
  assign _10466_ = inv_21[39] ^ r_20[39] /*12741*/;
  assign sum_21[39] = _10466_ ^ _10465_ /*12740*/;
  assign _10467_ = _10466_ & _10465_ /*12739*/;
  assign _10468_ = inv_21[39] & r_20[39] /*12738*/;
  assign _10469_ = _10467_ | _10468_ /*12737*/;
  assign _10470_ = inv_21[40] ^ r_20[40] /*12735*/;
  assign sum_21[40] = _10470_ ^ _10469_ /*12734*/;
  assign _10471_ = _10470_ & _10469_ /*12733*/;
  assign _10472_ = inv_21[40] & r_20[40] /*12732*/;
  assign _10473_ = _10471_ | _10472_ /*12731*/;
  assign _10474_ = inv_21[41] ^ r_20[41] /*12729*/;
  assign sum_21[41] = _10474_ ^ _10473_ /*12728*/;
  assign _10475_ = _10474_ & _10473_ /*12727*/;
  assign _10476_ = inv_21[41] & r_20[41] /*12726*/;
  assign _10477_ = _10475_ | _10476_ /*12725*/;
  assign _10478_ = inv_21[42] ^ r_20[42] /*12723*/;
  assign sum_21[42] = _10478_ ^ _10477_ /*12722*/;
  assign _10479_ = _10478_ & _10477_ /*12721*/;
  assign _10480_ = inv_21[42] & r_20[42] /*12720*/;
  assign _10481_ = _10479_ | _10480_ /*12719*/;
  assign _10482_ = inv_21[43] ^ r_20[43] /*12717*/;
  assign sum_21[43] = _10482_ ^ _10481_ /*12716*/;
  assign _10483_ = _10482_ & _10481_ /*12715*/;
  assign _10484_ = inv_21[43] & r_20[43] /*12714*/;
  assign _10485_ = _10483_ | _10484_ /*12713*/;
  assign _10486_ = inv_21[44] ^ r_20[44] /*12711*/;
  assign sum_21[44] = _10486_ ^ _10485_ /*12710*/;
  assign _10487_ = _10486_ & _10485_ /*12709*/;
  assign _10488_ = inv_21[44] & r_20[44] /*12708*/;
  assign _10489_ = _10487_ | _10488_ /*12707*/;
  assign _10490_ = inv_21[45] ^ r_20[45] /*12705*/;
  assign sum_21[45] = _10490_ ^ _10489_ /*12704*/;
  assign _10491_ = _10490_ & _10489_ /*12703*/;
  assign _10492_ = inv_21[45] & r_20[45] /*12702*/;
  assign _10493_ = _10491_ | _10492_ /*12701*/;
  assign _10494_ = inv_21[46] ^ r_20[46] /*12699*/;
  assign sum_21[46] = _10494_ ^ _10493_ /*12698*/;
  assign _10495_ = _10494_ & _10493_ /*12697*/;
  assign _10496_ = inv_21[46] & r_20[46] /*12696*/;
  assign _10497_ = _10495_ | _10496_ /*12695*/;
  assign _10498_ = inv_21[47] ^ r_20[47] /*12693*/;
  assign sum_21[47] = _10498_ ^ _10497_ /*12692*/;
  assign _10499_ = _10498_ & _10497_ /*12691*/;
  assign _10500_ = inv_21[47] & r_20[47] /*12690*/;
  assign _10501_ = _10499_ | _10500_ /*12689*/;
  assign _10502_ = inv_21[48] ^ r_20[48] /*12687*/;
  assign sum_21[48] = _10502_ ^ _10501_ /*12686*/;
  assign _10503_ = _10502_ & _10501_ /*12685*/;
  assign _10504_ = inv_21[48] & r_20[48] /*12684*/;
  assign _10505_ = _10503_ | _10504_ /*12683*/;
  assign _10506_ = inv_21[49] ^ r_20[49] /*12681*/;
  assign sum_21[49] = _10506_ ^ _10505_ /*12680*/;
  assign _10507_ = _10506_ & _10505_ /*12679*/;
  assign _10508_ = inv_21[49] & r_20[49] /*12678*/;
  assign _10509_ = _10507_ | _10508_ /*12677*/;
  assign _10510_ = inv_21[50] ^ r_20[50] /*12675*/;
  assign sum_21[50] = _10510_ ^ _10509_ /*12674*/;
  assign _10511_ = _10510_ & _10509_ /*12673*/;
  assign _10512_ = inv_21[50] & r_20[50] /*12672*/;
  assign _10513_ = _10511_ | _10512_ /*12671*/;
  assign _10514_ = inv_21[51] ^ r_20[51] /*12669*/;
  assign sum_21[51] = _10514_ ^ _10513_ /*12668*/;
  assign _10515_ = _10514_ & _10513_ /*12667*/;
  assign _10516_ = inv_21[51] & r_20[51] /*12666*/;
  assign _10517_ = _10515_ | _10516_ /*12665*/;
  assign _10518_ = inv_21[52] ^ r_20[52] /*12663*/;
  assign sum_21[52] = _10518_ ^ _10517_ /*12662*/;
  assign _10519_ = _10518_ & _10517_ /*12661*/;
  assign _10520_ = inv_21[52] & r_20[52] /*12660*/;
  assign _10521_ = _10519_ | _10520_ /*12659*/;
  assign _10522_ = inv_21[53] ^ r_20[53] /*12657*/;
  assign sum_21[53] = _10522_ ^ _10521_ /*12656*/;
  assign _10523_ = _10522_ & _10521_ /*12655*/;
  assign _10524_ = inv_21[53] & r_20[53] /*12654*/;
  assign _10525_ = _10523_ | _10524_ /*12653*/;
  assign _10526_ = inv_21[54] ^ r_20[54] /*12651*/;
  assign sum_21[54] = _10526_ ^ _10525_ /*12650*/;
  assign _10527_ = _10526_ & _10525_ /*12649*/;
  assign _10528_ = inv_21[54] & r_20[54] /*12648*/;
  assign _10529_ = _10527_ | _10528_ /*12647*/;
  assign _10530_ = inv_21[55] ^ r_20[55] /*12645*/;
  assign sum_21[55] = _10530_ ^ _10529_ /*12644*/;
  assign _10531_ = _10530_ & _10529_ /*12643*/;
  assign _10532_ = inv_21[55] & r_20[55] /*12642*/;
  assign _10533_ = _10531_ | _10532_ /*12641*/;
  assign _10534_ = inv_21[56] ^ r_20[56] /*12639*/;
  assign sum_21[56] = _10534_ ^ _10533_ /*12638*/;
  assign _10535_ = _10534_ & _10533_ /*12637*/;
  assign _10536_ = inv_21[56] & r_20[56] /*12636*/;
  assign _10537_ = _10535_ | _10536_ /*12635*/;
  assign _10538_ = inv_21[57] ^ r_20[57] /*12633*/;
  assign sum_21[57] = _10538_ ^ _10537_ /*12632*/;
  assign _10539_ = _10538_ & _10537_ /*12631*/;
  assign _10540_ = inv_21[57] & r_20[57] /*12630*/;
  assign _10541_ = _10539_ | _10540_ /*12629*/;
  assign _10542_ = inv_21[58] ^ r_20[58] /*12627*/;
  assign sum_21[58] = _10542_ ^ _10541_ /*12626*/;
  assign _10543_ = _10542_ & _10541_ /*12625*/;
  assign _10544_ = inv_21[58] & r_20[58] /*12624*/;
  assign _10545_ = _10543_ | _10544_ /*12623*/;
  assign _10546_ = inv_21[59] ^ r_20[59] /*12621*/;
  assign sum_21[59] = _10546_ ^ _10545_ /*12620*/;
  assign _10547_ = _10546_ & _10545_ /*12619*/;
  assign _10548_ = inv_21[59] & r_20[59] /*12618*/;
  assign _10549_ = _10547_ | _10548_ /*12617*/;
  assign _10550_ = inv_21[60] ^ r_20[60] /*12615*/;
  assign sum_21[60] = _10550_ ^ _10549_ /*12614*/;
  assign _10551_ = _10550_ & _10549_ /*12613*/;
  assign _10552_ = inv_21[60] & r_20[60] /*12612*/;
  assign _10553_ = _10551_ | _10552_ /*12611*/;
  assign _10554_ = inv_21[61] ^ r_20[61] /*12609*/;
  assign sum_21[61] = _10554_ ^ _10553_ /*12608*/;
  assign _10555_ = _10554_ & _10553_ /*12607*/;
  assign _10556_ = inv_21[61] & r_20[61] /*12606*/;
  assign _10557_ = _10555_ | _10556_ /*12605*/;
  assign _10558_ = inv_21[62] ^ r_20[62] /*12603*/;
  assign sum_21[62] = _10558_ ^ _10557_ /*12602*/;
  assign _10559_ = _10558_ & _10557_ /*12601*/;
  assign _10560_ = inv_21[62] & r_20[62] /*12600*/;
  assign _10561_ = _10559_ | _10560_ /*12599*/;
  assign _10562_ = inv_21[63] ^ r_20[63] /*12597*/;
  assign sum_21[63] = _10562_ ^ _10561_ /*12596*/;
  assign _10563_ = _10562_ & _10561_ /*12595*/;
  assign _10564_ = inv_21[63] & r_20[63] /*12594*/;
  assign _10565_ = _10563_ | _10564_ /*12593*/;
  assign _10566_ = inv_21[64] ^ r_20[64] /*12591*/;
  assign sum_21[64] = _10566_ ^ _10565_ /*12590*/;
  assign _10567_ = _10566_ & _10565_ /*12589*/;
  assign _10568_ = inv_21[64] & r_20[64] /*12588*/;
  assign _10569_ = _10567_ | _10568_ /*12587*/;
  assign _10570_ = inv_21[65] ^ r_20[65] /*12585*/;
  assign sum_21[65] = _10570_ ^ _10569_ /*12584*/;
  assign _10571_ = _10570_ & _10569_ /*12583*/;
  assign _10572_ = inv_21[65] & r_20[65] /*12582*/;
  assign _10573_ = _10571_ | _10572_ /*12581*/;
  assign _10574_ = inv_21[66] ^ r_20[66] /*12579*/;
  assign sum_21[66] = _10574_ ^ _10573_ /*12578*/;
  assign _10575_ = _10574_ & _10573_ /*12577*/;
  assign _10576_ = inv_21[66] & r_20[66] /*12576*/;
  assign _10577_ = _10575_ | _10576_ /*12575*/;
  assign _10578_ = inv_21[67] ^ r_20[67] /*12573*/;
  assign sum_21[67] = _10578_ ^ _10577_ /*12572*/;
  assign _10579_ = _10578_ & _10577_ /*12571*/;
  assign _10580_ = inv_21[67] & r_20[67] /*12570*/;
  assign _10581_ = _10579_ | _10580_ /*12569*/;
  assign _10582_ = inv_21[68] ^ r_20[68] /*12567*/;
  assign sum_21[68] = _10582_ ^ _10581_ /*12566*/;
  assign _10583_ = _10582_ & _10581_ /*12565*/;
  assign _10584_ = inv_21[68] & r_20[68] /*12564*/;
  assign _10585_ = _10583_ | _10584_ /*12563*/;
  assign _10586_ = inv_21[69] ^ r_20[69] /*12561*/;
  assign sum_21[69] = _10586_ ^ _10585_ /*12560*/;
  assign _10587_ = _10586_ & _10585_ /*12559*/;
  assign _10588_ = inv_21[69] & r_20[69] /*12558*/;
  assign _10589_ = _10587_ | _10588_ /*12557*/;
  assign _10590_ = inv_21[70] ^ r_20[70] /*12555*/;
  assign sum_21[70] = _10590_ ^ _10589_ /*12554*/;
  assign _10591_ = _10590_ & _10589_ /*12553*/;
  assign _10592_ = inv_21[70] & r_20[70] /*12552*/;
  assign _10593_ = _10591_ | _10592_ /*12551*/;
  assign _10594_ = inv_21[71] ^ r_20[71] /*12549*/;
  assign sum_21[71] = _10594_ ^ _10593_ /*12548*/;
  assign _10595_ = _10594_ & _10593_ /*12547*/;
  assign _10596_ = inv_21[71] & r_20[71] /*12546*/;
  assign _10597_ = _10595_ | _10596_ /*12545*/;
  assign _10598_ = inv_21[72] ^ r_20[72] /*12543*/;
  assign sum_21[72] = _10598_ ^ _10597_ /*12542*/;
  assign _10599_ = _10598_ & _10597_ /*12541*/;
  assign _10600_ = inv_21[72] & r_20[72] /*12540*/;
  assign _10601_ = _10599_ | _10600_ /*12539*/;
  assign _10602_ = inv_21[73] ^ r_20[73] /*12537*/;
  assign sum_21[73] = _10602_ ^ _10601_ /*12536*/;
  assign _10603_ = _10602_ & _10601_ /*12535*/;
  assign _10604_ = inv_21[73] & r_20[73] /*12534*/;
  assign _10605_ = _10603_ | _10604_ /*12533*/;
  assign _10606_ = inv_21[74] ^ r_20[74] /*12531*/;
  assign sum_21[74] = _10606_ ^ _10605_ /*12530*/;
  assign _10607_ = _10606_ & _10605_ /*12529*/;
  assign _10608_ = inv_21[74] & r_20[74] /*12528*/;
  assign _10609_ = _10607_ | _10608_ /*12527*/;
  assign _10610_ = inv_21[75] ^ r_20[75] /*12525*/;
  assign sum_21[75] = _10610_ ^ _10609_ /*12524*/;
  assign _10611_ = _10610_ & _10609_ /*12523*/;
  assign _10612_ = inv_21[75] & r_20[75] /*12522*/;
  assign _10613_ = _10611_ | _10612_ /*12521*/;
  assign _10614_ = inv_21[76] ^ r_20[76] /*12519*/;
  assign sum_21[76] = _10614_ ^ _10613_ /*12518*/;
  assign _10615_ = _10614_ & _10613_ /*12517*/;
  assign _10616_ = inv_21[76] & r_20[76] /*12516*/;
  assign _10617_ = _10615_ | _10616_ /*12515*/;
  assign _10618_ = inv_21[77] ^ r_20[77] /*12513*/;
  assign sum_21[77] = _10618_ ^ _10617_ /*12512*/;
  assign _10619_ = _10618_ & _10617_ /*12511*/;
  assign _10620_ = inv_21[77] & r_20[77] /*12510*/;
  assign _10621_ = _10619_ | _10620_ /*12509*/;
  assign _10622_ = inv_21[78] ^ r_20[78] /*12507*/;
  assign sum_21[78] = _10622_ ^ _10621_ /*12506*/;
  assign _10623_ = _10622_ & _10621_ /*12505*/;
  assign _10624_ = inv_21[78] & r_20[78] /*12504*/;
  assign _10625_ = _10623_ | _10624_ /*12503*/;
  assign _10626_ = inv_21[79] ^ r_20[79] /*12501*/;
  assign sum_21[79] = _10626_ ^ _10625_ /*12500*/;
  assign _10627_ = _10626_ & _10625_ /*12499*/;
  assign _10628_ = inv_21[79] & r_20[79] /*12498*/;
  assign _10629_ = _10627_ | _10628_ /*12497*/;
  assign _10630_ = inv_21[80] ^ r_20[80] /*12495*/;
  assign sum_21[80] = _10630_ ^ _10629_ /*12494*/;
  assign _10631_ = _10630_ & _10629_ /*12493*/;
  assign _10632_ = inv_21[80] & r_20[80] /*12492*/;
  assign _10633_ = _10631_ | _10632_ /*12491*/;
  assign _10634_ = inv_21[81] ^ r_20[81] /*12489*/;
  assign sum_21[81] = _10634_ ^ _10633_ /*12488*/;
  assign _10635_ = _10634_ & _10633_ /*12487*/;
  assign _10636_ = inv_21[81] & r_20[81] /*12486*/;
  assign _10637_ = _10635_ | _10636_ /*12485*/;
  assign _10638_ = inv_21[82] ^ r_20[82] /*12483*/;
  assign sum_21[82] = _10638_ ^ _10637_ /*12482*/;
  assign _10639_ = _10638_ & _10637_ /*12481*/;
  assign _10640_ = inv_21[82] & r_20[82] /*12480*/;
  assign _10641_ = _10639_ | _10640_ /*12479*/;
  assign _10642_ = _10641_ ^ _10637_ /*12478*/;
  assign _10643_ = ~_10642_ /*12477*/;
  assign _10644_ = sum_21[82] & _10643_ /*12476*/;
  assign _10645_ = _10642_ & _10641_ /*12475*/;
  assign sum_21[83] = _10645_ | _10644_ /*12474*/;
  assign q[11] = ~sum_21[83] /*12473*/;
  assign m_21[0] = r_20[0] /*12472*/;
  assign m_21[1] = r_20[1] /*12471*/;
  assign m_21[2] = r_20[2] /*12470*/;
  assign m_21[3] = r_20[3] /*12469*/;
  assign m_21[4] = r_20[4] /*12468*/;
  assign m_21[5] = r_20[5] /*12467*/;
  assign m_21[6] = r_20[6] /*12466*/;
  assign m_21[7] = r_20[7] /*12465*/;
  assign m_21[8] = r_20[8] /*12464*/;
  assign m_21[9] = r_20[9] /*12463*/;
  assign m_21[10] = r_20[10] /*12462*/;
  assign m_21[11] = r_20[11] /*12461*/;
  assign m_21[12] = r_20[12] /*12460*/;
  assign m_21[13] = r_20[13] /*12459*/;
  assign m_21[14] = r_20[14] /*12458*/;
  assign m_21[15] = r_20[15] /*12457*/;
  assign m_21[16] = r_20[16] /*12456*/;
  assign m_21[17] = r_20[17] /*12455*/;
  assign m_21[18] = r_20[18] /*12454*/;
  assign m_21[19] = r_20[19] /*12453*/;
  assign m_21[20] = r_20[20] /*12452*/;
  assign m_21[21] = r_20[21] /*12451*/;
  assign m_21[22] = r_20[22] /*12450*/;
  assign m_21[23] = r_20[23] /*12449*/;
  assign m_21[24] = r_20[24] /*12448*/;
  assign m_21[25] = r_20[25] /*12447*/;
  assign m_21[26] = r_20[26] /*12446*/;
  assign m_21[27] = r_20[27] /*12445*/;
  assign m_21[28] = r_20[28] /*12444*/;
  assign m_21[29] = r_20[29] /*12443*/;
  assign m_21[30] = r_20[30] /*12442*/;
  assign m_21[31] = r_20[31] /*12441*/;
  assign m_21[32] = r_20[32] /*12440*/;
  assign m_21[33] = r_20[33] /*12439*/;
  assign m_21[34] = r_20[34] /*12438*/;
  assign m_21[35] = r_20[35] /*12437*/;
  assign m_21[36] = r_20[36] /*12436*/;
  assign m_21[37] = r_20[37] /*12435*/;
  assign m_21[38] = r_20[38] /*12434*/;
  assign m_21[39] = r_20[39] /*12433*/;
  assign m_21[40] = r_20[40] /*12432*/;
  assign m_21[41] = r_20[41] /*12431*/;
  assign m_21[42] = r_20[42] /*12430*/;
  assign m_21[43] = r_20[43] /*12429*/;
  assign m_21[44] = r_20[44] /*12428*/;
  assign m_21[45] = r_20[45] /*12427*/;
  assign m_21[46] = r_20[46] /*12426*/;
  assign m_21[47] = r_20[47] /*12425*/;
  assign m_21[48] = r_20[48] /*12424*/;
  assign m_21[49] = r_20[49] /*12423*/;
  assign m_21[50] = r_20[50] /*12422*/;
  assign m_21[51] = r_20[51] /*12421*/;
  assign m_21[52] = r_20[52] /*12420*/;
  assign m_21[53] = r_20[53] /*12419*/;
  assign m_21[54] = r_20[54] /*12418*/;
  assign m_21[55] = r_20[55] /*12417*/;
  assign m_21[56] = r_20[56] /*12416*/;
  assign m_21[57] = r_20[57] /*12415*/;
  assign m_21[58] = r_20[58] /*12414*/;
  assign m_21[59] = r_20[59] /*12413*/;
  assign m_21[60] = r_20[60] /*12412*/;
  assign m_21[61] = r_20[61] /*12411*/;
  assign m_21[62] = r_20[62] /*12410*/;
  assign m_21[63] = r_20[63] /*12409*/;
  assign m_21[64] = r_20[64] /*12408*/;
  assign m_21[65] = r_20[65] /*12407*/;
  assign m_21[66] = r_20[66] /*12406*/;
  assign m_21[67] = r_20[67] /*12405*/;
  assign m_21[68] = r_20[68] /*12404*/;
  assign m_21[69] = r_20[69] /*12403*/;
  assign m_21[70] = r_20[70] /*12402*/;
  assign m_21[71] = r_20[71] /*12401*/;
  assign m_21[72] = r_20[72] /*12400*/;
  assign m_21[73] = r_20[73] /*12399*/;
  assign m_21[74] = r_20[74] /*12398*/;
  assign m_21[75] = r_20[75] /*12397*/;
  assign m_21[76] = r_20[76] /*12396*/;
  assign m_21[77] = r_20[77] /*12395*/;
  assign m_21[78] = r_20[78] /*12394*/;
  assign m_21[79] = r_20[79] /*12393*/;
  assign m_21[80] = r_20[80] /*12392*/;
  assign m_21[81] = r_20[81] /*12391*/;
  assign m_21[82] = r_20[82] /*12390*/;
  assign m_21[83] = r_20[82] /*12389*/;
  assign _10647_ = ~q[11] /*12388*/;
  assign _10648_ = sum_21[0] & q[11] /*12387*/;
  assign _10649_ = m_21[0] & _10647_ /*12386*/;
  assign r_21[0] = _10649_ | _10648_ /*12385*/;
  assign _10650_ = ~q[11] /*12384*/;
  assign _10651_ = sum_21[1] & q[11] /*12383*/;
  assign _10652_ = m_21[1] & _10650_ /*12382*/;
  assign r_21[1] = _10652_ | _10651_ /*12381*/;
  assign _10653_ = ~q[11] /*12380*/;
  assign _10654_ = sum_21[2] & q[11] /*12379*/;
  assign _10655_ = m_21[2] & _10653_ /*12378*/;
  assign r_21[2] = _10655_ | _10654_ /*12377*/;
  assign _10656_ = ~q[11] /*12376*/;
  assign _10657_ = sum_21[3] & q[11] /*12375*/;
  assign _10658_ = m_21[3] & _10656_ /*12374*/;
  assign r_21[3] = _10658_ | _10657_ /*12373*/;
  assign _10659_ = ~q[11] /*12372*/;
  assign _10660_ = sum_21[4] & q[11] /*12371*/;
  assign _10661_ = m_21[4] & _10659_ /*12370*/;
  assign r_21[4] = _10661_ | _10660_ /*12369*/;
  assign _10662_ = ~q[11] /*12368*/;
  assign _10663_ = sum_21[5] & q[11] /*12367*/;
  assign _10664_ = m_21[5] & _10662_ /*12366*/;
  assign r_21[5] = _10664_ | _10663_ /*12365*/;
  assign _10665_ = ~q[11] /*12364*/;
  assign _10666_ = sum_21[6] & q[11] /*12363*/;
  assign _10667_ = m_21[6] & _10665_ /*12362*/;
  assign r_21[6] = _10667_ | _10666_ /*12361*/;
  assign _10668_ = ~q[11] /*12360*/;
  assign _10669_ = sum_21[7] & q[11] /*12359*/;
  assign _10670_ = m_21[7] & _10668_ /*12358*/;
  assign r_21[7] = _10670_ | _10669_ /*12357*/;
  assign _10671_ = ~q[11] /*12356*/;
  assign _10672_ = sum_21[8] & q[11] /*12355*/;
  assign _10673_ = m_21[8] & _10671_ /*12354*/;
  assign r_21[8] = _10673_ | _10672_ /*12353*/;
  assign _10674_ = ~q[11] /*12352*/;
  assign _10675_ = sum_21[9] & q[11] /*12351*/;
  assign _10676_ = m_21[9] & _10674_ /*12350*/;
  assign r_21[9] = _10676_ | _10675_ /*12349*/;
  assign _10677_ = ~q[11] /*12348*/;
  assign _10678_ = sum_21[10] & q[11] /*12347*/;
  assign _10679_ = m_21[10] & _10677_ /*12346*/;
  assign r_21[10] = _10679_ | _10678_ /*12345*/;
  assign _10680_ = ~q[11] /*12344*/;
  assign _10681_ = sum_21[11] & q[11] /*12343*/;
  assign _10682_ = m_21[11] & _10680_ /*12342*/;
  assign r_21[11] = _10682_ | _10681_ /*12341*/;
  assign _10683_ = ~q[11] /*12340*/;
  assign _10684_ = sum_21[12] & q[11] /*12339*/;
  assign _10685_ = m_21[12] & _10683_ /*12338*/;
  assign r_21[12] = _10685_ | _10684_ /*12337*/;
  assign _10686_ = ~q[11] /*12336*/;
  assign _10687_ = sum_21[13] & q[11] /*12335*/;
  assign _10688_ = m_21[13] & _10686_ /*12334*/;
  assign r_21[13] = _10688_ | _10687_ /*12333*/;
  assign _10689_ = ~q[11] /*12332*/;
  assign _10690_ = sum_21[14] & q[11] /*12331*/;
  assign _10691_ = m_21[14] & _10689_ /*12330*/;
  assign r_21[14] = _10691_ | _10690_ /*12329*/;
  assign _10692_ = ~q[11] /*12328*/;
  assign _10693_ = sum_21[15] & q[11] /*12327*/;
  assign _10694_ = m_21[15] & _10692_ /*12326*/;
  assign r_21[15] = _10694_ | _10693_ /*12325*/;
  assign _10695_ = ~q[11] /*12324*/;
  assign _10696_ = sum_21[16] & q[11] /*12323*/;
  assign _10697_ = m_21[16] & _10695_ /*12322*/;
  assign r_21[16] = _10697_ | _10696_ /*12321*/;
  assign _10698_ = ~q[11] /*12320*/;
  assign _10699_ = sum_21[17] & q[11] /*12319*/;
  assign _10700_ = m_21[17] & _10698_ /*12318*/;
  assign r_21[17] = _10700_ | _10699_ /*12317*/;
  assign _10701_ = ~q[11] /*12316*/;
  assign _10702_ = sum_21[18] & q[11] /*12315*/;
  assign _10703_ = m_21[18] & _10701_ /*12314*/;
  assign r_21[18] = _10703_ | _10702_ /*12313*/;
  assign _10704_ = ~q[11] /*12312*/;
  assign _10705_ = sum_21[19] & q[11] /*12311*/;
  assign _10706_ = m_21[19] & _10704_ /*12310*/;
  assign r_21[19] = _10706_ | _10705_ /*12309*/;
  assign _10707_ = ~q[11] /*12308*/;
  assign _10708_ = sum_21[20] & q[11] /*12307*/;
  assign _10709_ = m_21[20] & _10707_ /*12306*/;
  assign r_21[20] = _10709_ | _10708_ /*12305*/;
  assign _10710_ = ~q[11] /*12304*/;
  assign _10711_ = sum_21[21] & q[11] /*12303*/;
  assign _10712_ = m_21[21] & _10710_ /*12302*/;
  assign r_21[21] = _10712_ | _10711_ /*12301*/;
  assign _10713_ = ~q[11] /*12300*/;
  assign _10714_ = sum_21[22] & q[11] /*12299*/;
  assign _10715_ = m_21[22] & _10713_ /*12298*/;
  assign r_21[22] = _10715_ | _10714_ /*12297*/;
  assign _10716_ = ~q[11] /*12296*/;
  assign _10717_ = sum_21[23] & q[11] /*12295*/;
  assign _10718_ = m_21[23] & _10716_ /*12294*/;
  assign r_21[23] = _10718_ | _10717_ /*12293*/;
  assign _10719_ = ~q[11] /*12292*/;
  assign _10720_ = sum_21[24] & q[11] /*12291*/;
  assign _10721_ = m_21[24] & _10719_ /*12290*/;
  assign r_21[24] = _10721_ | _10720_ /*12289*/;
  assign _10722_ = ~q[11] /*12288*/;
  assign _10723_ = sum_21[25] & q[11] /*12287*/;
  assign _10724_ = m_21[25] & _10722_ /*12286*/;
  assign r_21[25] = _10724_ | _10723_ /*12285*/;
  assign _10725_ = ~q[11] /*12284*/;
  assign _10726_ = sum_21[26] & q[11] /*12283*/;
  assign _10727_ = m_21[26] & _10725_ /*12282*/;
  assign r_21[26] = _10727_ | _10726_ /*12281*/;
  assign _10728_ = ~q[11] /*12280*/;
  assign _10729_ = sum_21[27] & q[11] /*12279*/;
  assign _10730_ = m_21[27] & _10728_ /*12278*/;
  assign r_21[27] = _10730_ | _10729_ /*12277*/;
  assign _10731_ = ~q[11] /*12276*/;
  assign _10732_ = sum_21[28] & q[11] /*12275*/;
  assign _10733_ = m_21[28] & _10731_ /*12274*/;
  assign r_21[28] = _10733_ | _10732_ /*12273*/;
  assign _10734_ = ~q[11] /*12272*/;
  assign _10735_ = sum_21[29] & q[11] /*12271*/;
  assign _10736_ = m_21[29] & _10734_ /*12270*/;
  assign r_21[29] = _10736_ | _10735_ /*12269*/;
  assign _10737_ = ~q[11] /*12268*/;
  assign _10738_ = sum_21[30] & q[11] /*12267*/;
  assign _10739_ = m_21[30] & _10737_ /*12266*/;
  assign r_21[30] = _10739_ | _10738_ /*12265*/;
  assign _10740_ = ~q[11] /*12264*/;
  assign _10741_ = sum_21[31] & q[11] /*12263*/;
  assign _10742_ = m_21[31] & _10740_ /*12262*/;
  assign r_21[31] = _10742_ | _10741_ /*12261*/;
  assign _10743_ = ~q[11] /*12260*/;
  assign _10744_ = sum_21[32] & q[11] /*12259*/;
  assign _10745_ = m_21[32] & _10743_ /*12258*/;
  assign r_21[32] = _10745_ | _10744_ /*12257*/;
  assign _10746_ = ~q[11] /*12256*/;
  assign _10747_ = sum_21[33] & q[11] /*12255*/;
  assign _10748_ = m_21[33] & _10746_ /*12254*/;
  assign r_21[33] = _10748_ | _10747_ /*12253*/;
  assign _10749_ = ~q[11] /*12252*/;
  assign _10750_ = sum_21[34] & q[11] /*12251*/;
  assign _10751_ = m_21[34] & _10749_ /*12250*/;
  assign r_21[34] = _10751_ | _10750_ /*12249*/;
  assign _10752_ = ~q[11] /*12248*/;
  assign _10753_ = sum_21[35] & q[11] /*12247*/;
  assign _10754_ = m_21[35] & _10752_ /*12246*/;
  assign r_21[35] = _10754_ | _10753_ /*12245*/;
  assign _10755_ = ~q[11] /*12244*/;
  assign _10756_ = sum_21[36] & q[11] /*12243*/;
  assign _10757_ = m_21[36] & _10755_ /*12242*/;
  assign r_21[36] = _10757_ | _10756_ /*12241*/;
  assign _10758_ = ~q[11] /*12240*/;
  assign _10759_ = sum_21[37] & q[11] /*12239*/;
  assign _10760_ = m_21[37] & _10758_ /*12238*/;
  assign r_21[37] = _10760_ | _10759_ /*12237*/;
  assign _10761_ = ~q[11] /*12236*/;
  assign _10762_ = sum_21[38] & q[11] /*12235*/;
  assign _10763_ = m_21[38] & _10761_ /*12234*/;
  assign r_21[38] = _10763_ | _10762_ /*12233*/;
  assign _10764_ = ~q[11] /*12232*/;
  assign _10765_ = sum_21[39] & q[11] /*12231*/;
  assign _10766_ = m_21[39] & _10764_ /*12230*/;
  assign r_21[39] = _10766_ | _10765_ /*12229*/;
  assign _10767_ = ~q[11] /*12228*/;
  assign _10768_ = sum_21[40] & q[11] /*12227*/;
  assign _10769_ = m_21[40] & _10767_ /*12226*/;
  assign r_21[40] = _10769_ | _10768_ /*12225*/;
  assign _10770_ = ~q[11] /*12224*/;
  assign _10771_ = sum_21[41] & q[11] /*12223*/;
  assign _10772_ = m_21[41] & _10770_ /*12222*/;
  assign r_21[41] = _10772_ | _10771_ /*12221*/;
  assign _10773_ = ~q[11] /*12220*/;
  assign _10774_ = sum_21[42] & q[11] /*12219*/;
  assign _10775_ = m_21[42] & _10773_ /*12218*/;
  assign r_21[42] = _10775_ | _10774_ /*12217*/;
  assign _10776_ = ~q[11] /*12216*/;
  assign _10777_ = sum_21[43] & q[11] /*12215*/;
  assign _10778_ = m_21[43] & _10776_ /*12214*/;
  assign r_21[43] = _10778_ | _10777_ /*12213*/;
  assign _10779_ = ~q[11] /*12212*/;
  assign _10780_ = sum_21[44] & q[11] /*12211*/;
  assign _10781_ = m_21[44] & _10779_ /*12210*/;
  assign r_21[44] = _10781_ | _10780_ /*12209*/;
  assign _10782_ = ~q[11] /*12208*/;
  assign _10783_ = sum_21[45] & q[11] /*12207*/;
  assign _10784_ = m_21[45] & _10782_ /*12206*/;
  assign r_21[45] = _10784_ | _10783_ /*12205*/;
  assign _10785_ = ~q[11] /*12204*/;
  assign _10786_ = sum_21[46] & q[11] /*12203*/;
  assign _10787_ = m_21[46] & _10785_ /*12202*/;
  assign r_21[46] = _10787_ | _10786_ /*12201*/;
  assign _10788_ = ~q[11] /*12200*/;
  assign _10789_ = sum_21[47] & q[11] /*12199*/;
  assign _10790_ = m_21[47] & _10788_ /*12198*/;
  assign r_21[47] = _10790_ | _10789_ /*12197*/;
  assign _10791_ = ~q[11] /*12196*/;
  assign _10792_ = sum_21[48] & q[11] /*12195*/;
  assign _10793_ = m_21[48] & _10791_ /*12194*/;
  assign r_21[48] = _10793_ | _10792_ /*12193*/;
  assign _10794_ = ~q[11] /*12192*/;
  assign _10795_ = sum_21[49] & q[11] /*12191*/;
  assign _10796_ = m_21[49] & _10794_ /*12190*/;
  assign r_21[49] = _10796_ | _10795_ /*12189*/;
  assign _10797_ = ~q[11] /*12188*/;
  assign _10798_ = sum_21[50] & q[11] /*12187*/;
  assign _10799_ = m_21[50] & _10797_ /*12186*/;
  assign r_21[50] = _10799_ | _10798_ /*12185*/;
  assign _10800_ = ~q[11] /*12184*/;
  assign _10801_ = sum_21[51] & q[11] /*12183*/;
  assign _10802_ = m_21[51] & _10800_ /*12182*/;
  assign r_21[51] = _10802_ | _10801_ /*12181*/;
  assign _10803_ = ~q[11] /*12180*/;
  assign _10804_ = sum_21[52] & q[11] /*12179*/;
  assign _10805_ = m_21[52] & _10803_ /*12178*/;
  assign r_21[52] = _10805_ | _10804_ /*12177*/;
  assign _10806_ = ~q[11] /*12176*/;
  assign _10807_ = sum_21[53] & q[11] /*12175*/;
  assign _10808_ = m_21[53] & _10806_ /*12174*/;
  assign r_21[53] = _10808_ | _10807_ /*12173*/;
  assign _10809_ = ~q[11] /*12172*/;
  assign _10810_ = sum_21[54] & q[11] /*12171*/;
  assign _10811_ = m_21[54] & _10809_ /*12170*/;
  assign r_21[54] = _10811_ | _10810_ /*12169*/;
  assign _10812_ = ~q[11] /*12168*/;
  assign _10813_ = sum_21[55] & q[11] /*12167*/;
  assign _10814_ = m_21[55] & _10812_ /*12166*/;
  assign r_21[55] = _10814_ | _10813_ /*12165*/;
  assign _10815_ = ~q[11] /*12164*/;
  assign _10816_ = sum_21[56] & q[11] /*12163*/;
  assign _10817_ = m_21[56] & _10815_ /*12162*/;
  assign r_21[56] = _10817_ | _10816_ /*12161*/;
  assign _10818_ = ~q[11] /*12160*/;
  assign _10819_ = sum_21[57] & q[11] /*12159*/;
  assign _10820_ = m_21[57] & _10818_ /*12158*/;
  assign r_21[57] = _10820_ | _10819_ /*12157*/;
  assign _10821_ = ~q[11] /*12156*/;
  assign _10822_ = sum_21[58] & q[11] /*12155*/;
  assign _10823_ = m_21[58] & _10821_ /*12154*/;
  assign r_21[58] = _10823_ | _10822_ /*12153*/;
  assign _10824_ = ~q[11] /*12152*/;
  assign _10825_ = sum_21[59] & q[11] /*12151*/;
  assign _10826_ = m_21[59] & _10824_ /*12150*/;
  assign r_21[59] = _10826_ | _10825_ /*12149*/;
  assign _10827_ = ~q[11] /*12148*/;
  assign _10828_ = sum_21[60] & q[11] /*12147*/;
  assign _10829_ = m_21[60] & _10827_ /*12146*/;
  assign r_21[60] = _10829_ | _10828_ /*12145*/;
  assign _10830_ = ~q[11] /*12144*/;
  assign _10831_ = sum_21[61] & q[11] /*12143*/;
  assign _10832_ = m_21[61] & _10830_ /*12142*/;
  assign r_21[61] = _10832_ | _10831_ /*12141*/;
  assign _10833_ = ~q[11] /*12140*/;
  assign _10834_ = sum_21[62] & q[11] /*12139*/;
  assign _10835_ = m_21[62] & _10833_ /*12138*/;
  assign r_21[62] = _10835_ | _10834_ /*12137*/;
  assign _10836_ = ~q[11] /*12136*/;
  assign _10837_ = sum_21[63] & q[11] /*12135*/;
  assign _10838_ = m_21[63] & _10836_ /*12134*/;
  assign r_21[63] = _10838_ | _10837_ /*12133*/;
  assign _10839_ = ~q[11] /*12132*/;
  assign _10840_ = sum_21[64] & q[11] /*12131*/;
  assign _10841_ = m_21[64] & _10839_ /*12130*/;
  assign r_21[64] = _10841_ | _10840_ /*12129*/;
  assign _10842_ = ~q[11] /*12128*/;
  assign _10843_ = sum_21[65] & q[11] /*12127*/;
  assign _10844_ = m_21[65] & _10842_ /*12126*/;
  assign r_21[65] = _10844_ | _10843_ /*12125*/;
  assign _10845_ = ~q[11] /*12124*/;
  assign _10846_ = sum_21[66] & q[11] /*12123*/;
  assign _10847_ = m_21[66] & _10845_ /*12122*/;
  assign r_21[66] = _10847_ | _10846_ /*12121*/;
  assign _10848_ = ~q[11] /*12120*/;
  assign _10849_ = sum_21[67] & q[11] /*12119*/;
  assign _10850_ = m_21[67] & _10848_ /*12118*/;
  assign r_21[67] = _10850_ | _10849_ /*12117*/;
  assign _10851_ = ~q[11] /*12116*/;
  assign _10852_ = sum_21[68] & q[11] /*12115*/;
  assign _10853_ = m_21[68] & _10851_ /*12114*/;
  assign r_21[68] = _10853_ | _10852_ /*12113*/;
  assign _10854_ = ~q[11] /*12112*/;
  assign _10855_ = sum_21[69] & q[11] /*12111*/;
  assign _10856_ = m_21[69] & _10854_ /*12110*/;
  assign r_21[69] = _10856_ | _10855_ /*12109*/;
  assign _10857_ = ~q[11] /*12108*/;
  assign _10858_ = sum_21[70] & q[11] /*12107*/;
  assign _10859_ = m_21[70] & _10857_ /*12106*/;
  assign r_21[70] = _10859_ | _10858_ /*12105*/;
  assign _10860_ = ~q[11] /*12104*/;
  assign _10861_ = sum_21[71] & q[11] /*12103*/;
  assign _10862_ = m_21[71] & _10860_ /*12102*/;
  assign r_21[71] = _10862_ | _10861_ /*12101*/;
  assign _10863_ = ~q[11] /*12100*/;
  assign _10864_ = sum_21[72] & q[11] /*12099*/;
  assign _10865_ = m_21[72] & _10863_ /*12098*/;
  assign r_21[72] = _10865_ | _10864_ /*12097*/;
  assign _10866_ = ~q[11] /*12096*/;
  assign _10867_ = sum_21[73] & q[11] /*12095*/;
  assign _10868_ = m_21[73] & _10866_ /*12094*/;
  assign r_21[73] = _10868_ | _10867_ /*12093*/;
  assign _10869_ = ~q[11] /*12092*/;
  assign _10870_ = sum_21[74] & q[11] /*12091*/;
  assign _10871_ = m_21[74] & _10869_ /*12090*/;
  assign r_21[74] = _10871_ | _10870_ /*12089*/;
  assign _10872_ = ~q[11] /*12088*/;
  assign _10873_ = sum_21[75] & q[11] /*12087*/;
  assign _10874_ = m_21[75] & _10872_ /*12086*/;
  assign r_21[75] = _10874_ | _10873_ /*12085*/;
  assign _10875_ = ~q[11] /*12084*/;
  assign _10876_ = sum_21[76] & q[11] /*12083*/;
  assign _10877_ = m_21[76] & _10875_ /*12082*/;
  assign r_21[76] = _10877_ | _10876_ /*12081*/;
  assign _10878_ = ~q[11] /*12080*/;
  assign _10879_ = sum_21[77] & q[11] /*12079*/;
  assign _10880_ = m_21[77] & _10878_ /*12078*/;
  assign r_21[77] = _10880_ | _10879_ /*12077*/;
  assign _10881_ = ~q[11] /*12076*/;
  assign _10882_ = sum_21[78] & q[11] /*12075*/;
  assign _10883_ = m_21[78] & _10881_ /*12074*/;
  assign r_21[78] = _10883_ | _10882_ /*12073*/;
  assign _10884_ = ~q[11] /*12072*/;
  assign _10885_ = sum_21[79] & q[11] /*12071*/;
  assign _10886_ = m_21[79] & _10884_ /*12070*/;
  assign r_21[79] = _10886_ | _10885_ /*12069*/;
  assign _10887_ = ~q[11] /*12068*/;
  assign _10888_ = sum_21[80] & q[11] /*12067*/;
  assign _10889_ = m_21[80] & _10887_ /*12066*/;
  assign r_21[80] = _10889_ | _10888_ /*12065*/;
  assign _10890_ = ~q[11] /*12064*/;
  assign _10891_ = sum_21[81] & q[11] /*12063*/;
  assign _10892_ = m_21[81] & _10890_ /*12062*/;
  assign r_21[81] = _10892_ | _10891_ /*12061*/;
  assign _10893_ = ~q[11] /*12060*/;
  assign _10894_ = sum_21[82] & q[11] /*12059*/;
  assign _10895_ = m_21[82] & _10893_ /*12058*/;
  assign r_21[82] = _10895_ | _10894_ /*12057*/;
  assign _10896_ = ~q[11] /*12056*/;
  assign _10897_ = sum_21[83] & q[11] /*12055*/;
  assign _10898_ = m_21[83] & _10896_ /*12054*/;
  assign r_21[83] = _10898_ | _10897_ /*12053*/;
  assign inv_22[0] = oneWire /*11900*/;
  assign inv_22[1] = oneWire /*11894*/;
  assign inv_22[2] = oneWire /*11888*/;
  assign inv_22[3] = oneWire /*11882*/;
  assign inv_22[4] = oneWire /*11876*/;
  assign inv_22[5] = oneWire /*11870*/;
  assign inv_22[6] = oneWire /*11864*/;
  assign inv_22[7] = oneWire /*11858*/;
  assign inv_22[8] = oneWire /*11852*/;
  assign inv_22[9] = oneWire /*11846*/;
  assign inv_22[10] = ~div[0] /*11840*/;
  assign inv_22[11] = ~div[1] /*11834*/;
  assign inv_22[12] = ~div[2] /*11828*/;
  assign inv_22[13] = ~div[3] /*11822*/;
  assign inv_22[14] = ~div[4] /*11816*/;
  assign inv_22[15] = ~div[5] /*11810*/;
  assign inv_22[16] = ~div[6] /*11804*/;
  assign inv_22[17] = ~div[7] /*11798*/;
  assign inv_22[18] = ~div[8] /*11792*/;
  assign inv_22[19] = ~div[9] /*11786*/;
  assign inv_22[20] = ~div[10] /*11780*/;
  assign inv_22[21] = ~div[11] /*11774*/;
  assign inv_22[22] = ~div[12] /*11768*/;
  assign inv_22[23] = ~div[13] /*11762*/;
  assign inv_22[24] = ~div[14] /*11756*/;
  assign inv_22[25] = ~div[15] /*11750*/;
  assign inv_22[26] = ~div[16] /*11744*/;
  assign inv_22[27] = ~div[17] /*11738*/;
  assign inv_22[28] = ~div[18] /*11732*/;
  assign inv_22[29] = ~div[19] /*11726*/;
  assign inv_22[30] = ~div[20] /*11720*/;
  assign inv_22[31] = ~div[21] /*11714*/;
  assign inv_22[32] = ~div[22] /*11708*/;
  assign inv_22[33] = ~div[23] /*11702*/;
  assign inv_22[34] = ~div[24] /*11696*/;
  assign inv_22[35] = ~div[25] /*11690*/;
  assign inv_22[36] = ~div[26] /*11684*/;
  assign inv_22[37] = ~div[27] /*11678*/;
  assign inv_22[38] = ~div[28] /*11672*/;
  assign inv_22[39] = ~div[29] /*11666*/;
  assign inv_22[40] = ~div[30] /*11660*/;
  assign inv_22[41] = oneWire /*11654*/;
  assign inv_22[42] = oneWire /*11648*/;
  assign inv_22[43] = oneWire /*11642*/;
  assign inv_22[44] = oneWire /*11636*/;
  assign inv_22[45] = oneWire /*11630*/;
  assign inv_22[46] = oneWire /*11624*/;
  assign inv_22[47] = oneWire /*11618*/;
  assign inv_22[48] = oneWire /*11612*/;
  assign inv_22[49] = oneWire /*11606*/;
  assign inv_22[50] = oneWire /*11600*/;
  assign inv_22[51] = oneWire /*11594*/;
  assign inv_22[52] = oneWire /*11588*/;
  assign inv_22[53] = oneWire /*11582*/;
  assign inv_22[54] = oneWire /*11576*/;
  assign inv_22[55] = oneWire /*11570*/;
  assign inv_22[56] = oneWire /*11564*/;
  assign inv_22[57] = oneWire /*11558*/;
  assign inv_22[58] = oneWire /*11552*/;
  assign inv_22[59] = oneWire /*11546*/;
  assign inv_22[60] = oneWire /*11540*/;
  assign inv_22[61] = oneWire /*11534*/;
  assign inv_22[62] = oneWire /*11528*/;
  assign inv_22[63] = oneWire /*11522*/;
  assign inv_22[64] = oneWire /*11516*/;
  assign inv_22[65] = oneWire /*11510*/;
  assign inv_22[66] = oneWire /*11504*/;
  assign inv_22[67] = oneWire /*11498*/;
  assign inv_22[68] = oneWire /*11492*/;
  assign inv_22[69] = oneWire /*11486*/;
  assign inv_22[70] = oneWire /*11480*/;
  assign inv_22[71] = oneWire /*11474*/;
  assign inv_22[72] = oneWire /*11468*/;
  assign inv_22[73] = oneWire /*11462*/;
  assign inv_22[74] = oneWire /*11456*/;
  assign inv_22[75] = oneWire /*11450*/;
  assign inv_22[76] = oneWire /*11444*/;
  assign inv_22[77] = oneWire /*11438*/;
  assign inv_22[78] = oneWire /*11432*/;
  assign inv_22[79] = oneWire /*11426*/;
  assign inv_22[80] = oneWire /*11420*/;
  assign inv_22[81] = oneWire /*11414*/;
  assign inv_22[82] = oneWire /*11408*/;
  assign inv_22[83] = oneWire /*11402*/;
  assign _10899_ = inv_22[0] ^ r_21[0] /*11899*/;
  assign sum_22[0] = _10899_ ^ oneWire /*11898*/;
  assign _10900_ = _10899_ & oneWire /*11897*/;
  assign _10901_ = inv_22[0] & r_21[0] /*11896*/;
  assign _10902_ = _10900_ | _10901_ /*11895*/;
  assign _10903_ = inv_22[1] ^ r_21[1] /*11893*/;
  assign sum_22[1] = _10903_ ^ _10902_ /*11892*/;
  assign _10904_ = _10903_ & _10902_ /*11891*/;
  assign _10905_ = inv_22[1] & r_21[1] /*11890*/;
  assign _10906_ = _10904_ | _10905_ /*11889*/;
  assign _10907_ = inv_22[2] ^ r_21[2] /*11887*/;
  assign sum_22[2] = _10907_ ^ _10906_ /*11886*/;
  assign _10908_ = _10907_ & _10906_ /*11885*/;
  assign _10909_ = inv_22[2] & r_21[2] /*11884*/;
  assign _10910_ = _10908_ | _10909_ /*11883*/;
  assign _10911_ = inv_22[3] ^ r_21[3] /*11881*/;
  assign sum_22[3] = _10911_ ^ _10910_ /*11880*/;
  assign _10912_ = _10911_ & _10910_ /*11879*/;
  assign _10913_ = inv_22[3] & r_21[3] /*11878*/;
  assign _10914_ = _10912_ | _10913_ /*11877*/;
  assign _10915_ = inv_22[4] ^ r_21[4] /*11875*/;
  assign sum_22[4] = _10915_ ^ _10914_ /*11874*/;
  assign _10916_ = _10915_ & _10914_ /*11873*/;
  assign _10917_ = inv_22[4] & r_21[4] /*11872*/;
  assign _10918_ = _10916_ | _10917_ /*11871*/;
  assign _10919_ = inv_22[5] ^ r_21[5] /*11869*/;
  assign sum_22[5] = _10919_ ^ _10918_ /*11868*/;
  assign _10920_ = _10919_ & _10918_ /*11867*/;
  assign _10921_ = inv_22[5] & r_21[5] /*11866*/;
  assign _10922_ = _10920_ | _10921_ /*11865*/;
  assign _10923_ = inv_22[6] ^ r_21[6] /*11863*/;
  assign sum_22[6] = _10923_ ^ _10922_ /*11862*/;
  assign _10924_ = _10923_ & _10922_ /*11861*/;
  assign _10925_ = inv_22[6] & r_21[6] /*11860*/;
  assign _10926_ = _10924_ | _10925_ /*11859*/;
  assign _10927_ = inv_22[7] ^ r_21[7] /*11857*/;
  assign sum_22[7] = _10927_ ^ _10926_ /*11856*/;
  assign _10928_ = _10927_ & _10926_ /*11855*/;
  assign _10929_ = inv_22[7] & r_21[7] /*11854*/;
  assign _10930_ = _10928_ | _10929_ /*11853*/;
  assign _10931_ = inv_22[8] ^ r_21[8] /*11851*/;
  assign sum_22[8] = _10931_ ^ _10930_ /*11850*/;
  assign _10932_ = _10931_ & _10930_ /*11849*/;
  assign _10933_ = inv_22[8] & r_21[8] /*11848*/;
  assign _10934_ = _10932_ | _10933_ /*11847*/;
  assign _10935_ = inv_22[9] ^ r_21[9] /*11845*/;
  assign sum_22[9] = _10935_ ^ _10934_ /*11844*/;
  assign _10936_ = _10935_ & _10934_ /*11843*/;
  assign _10937_ = inv_22[9] & r_21[9] /*11842*/;
  assign _10938_ = _10936_ | _10937_ /*11841*/;
  assign _10939_ = inv_22[10] ^ r_21[10] /*11839*/;
  assign sum_22[10] = _10939_ ^ _10938_ /*11838*/;
  assign _10940_ = _10939_ & _10938_ /*11837*/;
  assign _10941_ = inv_22[10] & r_21[10] /*11836*/;
  assign _10942_ = _10940_ | _10941_ /*11835*/;
  assign _10943_ = inv_22[11] ^ r_21[11] /*11833*/;
  assign sum_22[11] = _10943_ ^ _10942_ /*11832*/;
  assign _10944_ = _10943_ & _10942_ /*11831*/;
  assign _10945_ = inv_22[11] & r_21[11] /*11830*/;
  assign _10946_ = _10944_ | _10945_ /*11829*/;
  assign _10947_ = inv_22[12] ^ r_21[12] /*11827*/;
  assign sum_22[12] = _10947_ ^ _10946_ /*11826*/;
  assign _10948_ = _10947_ & _10946_ /*11825*/;
  assign _10949_ = inv_22[12] & r_21[12] /*11824*/;
  assign _10950_ = _10948_ | _10949_ /*11823*/;
  assign _10951_ = inv_22[13] ^ r_21[13] /*11821*/;
  assign sum_22[13] = _10951_ ^ _10950_ /*11820*/;
  assign _10952_ = _10951_ & _10950_ /*11819*/;
  assign _10953_ = inv_22[13] & r_21[13] /*11818*/;
  assign _10954_ = _10952_ | _10953_ /*11817*/;
  assign _10955_ = inv_22[14] ^ r_21[14] /*11815*/;
  assign sum_22[14] = _10955_ ^ _10954_ /*11814*/;
  assign _10956_ = _10955_ & _10954_ /*11813*/;
  assign _10957_ = inv_22[14] & r_21[14] /*11812*/;
  assign _10958_ = _10956_ | _10957_ /*11811*/;
  assign _10959_ = inv_22[15] ^ r_21[15] /*11809*/;
  assign sum_22[15] = _10959_ ^ _10958_ /*11808*/;
  assign _10960_ = _10959_ & _10958_ /*11807*/;
  assign _10961_ = inv_22[15] & r_21[15] /*11806*/;
  assign _10962_ = _10960_ | _10961_ /*11805*/;
  assign _10963_ = inv_22[16] ^ r_21[16] /*11803*/;
  assign sum_22[16] = _10963_ ^ _10962_ /*11802*/;
  assign _10964_ = _10963_ & _10962_ /*11801*/;
  assign _10965_ = inv_22[16] & r_21[16] /*11800*/;
  assign _10966_ = _10964_ | _10965_ /*11799*/;
  assign _10967_ = inv_22[17] ^ r_21[17] /*11797*/;
  assign sum_22[17] = _10967_ ^ _10966_ /*11796*/;
  assign _10968_ = _10967_ & _10966_ /*11795*/;
  assign _10969_ = inv_22[17] & r_21[17] /*11794*/;
  assign _10970_ = _10968_ | _10969_ /*11793*/;
  assign _10971_ = inv_22[18] ^ r_21[18] /*11791*/;
  assign sum_22[18] = _10971_ ^ _10970_ /*11790*/;
  assign _10972_ = _10971_ & _10970_ /*11789*/;
  assign _10973_ = inv_22[18] & r_21[18] /*11788*/;
  assign _10974_ = _10972_ | _10973_ /*11787*/;
  assign _10975_ = inv_22[19] ^ r_21[19] /*11785*/;
  assign sum_22[19] = _10975_ ^ _10974_ /*11784*/;
  assign _10976_ = _10975_ & _10974_ /*11783*/;
  assign _10977_ = inv_22[19] & r_21[19] /*11782*/;
  assign _10978_ = _10976_ | _10977_ /*11781*/;
  assign _10979_ = inv_22[20] ^ r_21[20] /*11779*/;
  assign sum_22[20] = _10979_ ^ _10978_ /*11778*/;
  assign _10980_ = _10979_ & _10978_ /*11777*/;
  assign _10981_ = inv_22[20] & r_21[20] /*11776*/;
  assign _10982_ = _10980_ | _10981_ /*11775*/;
  assign _10983_ = inv_22[21] ^ r_21[21] /*11773*/;
  assign sum_22[21] = _10983_ ^ _10982_ /*11772*/;
  assign _10984_ = _10983_ & _10982_ /*11771*/;
  assign _10985_ = inv_22[21] & r_21[21] /*11770*/;
  assign _10986_ = _10984_ | _10985_ /*11769*/;
  assign _10987_ = inv_22[22] ^ r_21[22] /*11767*/;
  assign sum_22[22] = _10987_ ^ _10986_ /*11766*/;
  assign _10988_ = _10987_ & _10986_ /*11765*/;
  assign _10989_ = inv_22[22] & r_21[22] /*11764*/;
  assign _10990_ = _10988_ | _10989_ /*11763*/;
  assign _10991_ = inv_22[23] ^ r_21[23] /*11761*/;
  assign sum_22[23] = _10991_ ^ _10990_ /*11760*/;
  assign _10992_ = _10991_ & _10990_ /*11759*/;
  assign _10993_ = inv_22[23] & r_21[23] /*11758*/;
  assign _10994_ = _10992_ | _10993_ /*11757*/;
  assign _10995_ = inv_22[24] ^ r_21[24] /*11755*/;
  assign sum_22[24] = _10995_ ^ _10994_ /*11754*/;
  assign _10996_ = _10995_ & _10994_ /*11753*/;
  assign _10997_ = inv_22[24] & r_21[24] /*11752*/;
  assign _10998_ = _10996_ | _10997_ /*11751*/;
  assign _10999_ = inv_22[25] ^ r_21[25] /*11749*/;
  assign sum_22[25] = _10999_ ^ _10998_ /*11748*/;
  assign _11000_ = _10999_ & _10998_ /*11747*/;
  assign _11001_ = inv_22[25] & r_21[25] /*11746*/;
  assign _11002_ = _11000_ | _11001_ /*11745*/;
  assign _11003_ = inv_22[26] ^ r_21[26] /*11743*/;
  assign sum_22[26] = _11003_ ^ _11002_ /*11742*/;
  assign _11004_ = _11003_ & _11002_ /*11741*/;
  assign _11005_ = inv_22[26] & r_21[26] /*11740*/;
  assign _11006_ = _11004_ | _11005_ /*11739*/;
  assign _11007_ = inv_22[27] ^ r_21[27] /*11737*/;
  assign sum_22[27] = _11007_ ^ _11006_ /*11736*/;
  assign _11008_ = _11007_ & _11006_ /*11735*/;
  assign _11009_ = inv_22[27] & r_21[27] /*11734*/;
  assign _11010_ = _11008_ | _11009_ /*11733*/;
  assign _11011_ = inv_22[28] ^ r_21[28] /*11731*/;
  assign sum_22[28] = _11011_ ^ _11010_ /*11730*/;
  assign _11012_ = _11011_ & _11010_ /*11729*/;
  assign _11013_ = inv_22[28] & r_21[28] /*11728*/;
  assign _11014_ = _11012_ | _11013_ /*11727*/;
  assign _11015_ = inv_22[29] ^ r_21[29] /*11725*/;
  assign sum_22[29] = _11015_ ^ _11014_ /*11724*/;
  assign _11016_ = _11015_ & _11014_ /*11723*/;
  assign _11017_ = inv_22[29] & r_21[29] /*11722*/;
  assign _11018_ = _11016_ | _11017_ /*11721*/;
  assign _11019_ = inv_22[30] ^ r_21[30] /*11719*/;
  assign sum_22[30] = _11019_ ^ _11018_ /*11718*/;
  assign _11020_ = _11019_ & _11018_ /*11717*/;
  assign _11021_ = inv_22[30] & r_21[30] /*11716*/;
  assign _11022_ = _11020_ | _11021_ /*11715*/;
  assign _11023_ = inv_22[31] ^ r_21[31] /*11713*/;
  assign sum_22[31] = _11023_ ^ _11022_ /*11712*/;
  assign _11024_ = _11023_ & _11022_ /*11711*/;
  assign _11025_ = inv_22[31] & r_21[31] /*11710*/;
  assign _11026_ = _11024_ | _11025_ /*11709*/;
  assign _11027_ = inv_22[32] ^ r_21[32] /*11707*/;
  assign sum_22[32] = _11027_ ^ _11026_ /*11706*/;
  assign _11028_ = _11027_ & _11026_ /*11705*/;
  assign _11029_ = inv_22[32] & r_21[32] /*11704*/;
  assign _11030_ = _11028_ | _11029_ /*11703*/;
  assign _11031_ = inv_22[33] ^ r_21[33] /*11701*/;
  assign sum_22[33] = _11031_ ^ _11030_ /*11700*/;
  assign _11032_ = _11031_ & _11030_ /*11699*/;
  assign _11033_ = inv_22[33] & r_21[33] /*11698*/;
  assign _11034_ = _11032_ | _11033_ /*11697*/;
  assign _11035_ = inv_22[34] ^ r_21[34] /*11695*/;
  assign sum_22[34] = _11035_ ^ _11034_ /*11694*/;
  assign _11036_ = _11035_ & _11034_ /*11693*/;
  assign _11037_ = inv_22[34] & r_21[34] /*11692*/;
  assign _11038_ = _11036_ | _11037_ /*11691*/;
  assign _11039_ = inv_22[35] ^ r_21[35] /*11689*/;
  assign sum_22[35] = _11039_ ^ _11038_ /*11688*/;
  assign _11040_ = _11039_ & _11038_ /*11687*/;
  assign _11041_ = inv_22[35] & r_21[35] /*11686*/;
  assign _11042_ = _11040_ | _11041_ /*11685*/;
  assign _11043_ = inv_22[36] ^ r_21[36] /*11683*/;
  assign sum_22[36] = _11043_ ^ _11042_ /*11682*/;
  assign _11044_ = _11043_ & _11042_ /*11681*/;
  assign _11045_ = inv_22[36] & r_21[36] /*11680*/;
  assign _11046_ = _11044_ | _11045_ /*11679*/;
  assign _11047_ = inv_22[37] ^ r_21[37] /*11677*/;
  assign sum_22[37] = _11047_ ^ _11046_ /*11676*/;
  assign _11048_ = _11047_ & _11046_ /*11675*/;
  assign _11049_ = inv_22[37] & r_21[37] /*11674*/;
  assign _11050_ = _11048_ | _11049_ /*11673*/;
  assign _11051_ = inv_22[38] ^ r_21[38] /*11671*/;
  assign sum_22[38] = _11051_ ^ _11050_ /*11670*/;
  assign _11052_ = _11051_ & _11050_ /*11669*/;
  assign _11053_ = inv_22[38] & r_21[38] /*11668*/;
  assign _11054_ = _11052_ | _11053_ /*11667*/;
  assign _11055_ = inv_22[39] ^ r_21[39] /*11665*/;
  assign sum_22[39] = _11055_ ^ _11054_ /*11664*/;
  assign _11056_ = _11055_ & _11054_ /*11663*/;
  assign _11057_ = inv_22[39] & r_21[39] /*11662*/;
  assign _11058_ = _11056_ | _11057_ /*11661*/;
  assign _11059_ = inv_22[40] ^ r_21[40] /*11659*/;
  assign sum_22[40] = _11059_ ^ _11058_ /*11658*/;
  assign _11060_ = _11059_ & _11058_ /*11657*/;
  assign _11061_ = inv_22[40] & r_21[40] /*11656*/;
  assign _11062_ = _11060_ | _11061_ /*11655*/;
  assign _11063_ = inv_22[41] ^ r_21[41] /*11653*/;
  assign sum_22[41] = _11063_ ^ _11062_ /*11652*/;
  assign _11064_ = _11063_ & _11062_ /*11651*/;
  assign _11065_ = inv_22[41] & r_21[41] /*11650*/;
  assign _11066_ = _11064_ | _11065_ /*11649*/;
  assign _11067_ = inv_22[42] ^ r_21[42] /*11647*/;
  assign sum_22[42] = _11067_ ^ _11066_ /*11646*/;
  assign _11068_ = _11067_ & _11066_ /*11645*/;
  assign _11069_ = inv_22[42] & r_21[42] /*11644*/;
  assign _11070_ = _11068_ | _11069_ /*11643*/;
  assign _11071_ = inv_22[43] ^ r_21[43] /*11641*/;
  assign sum_22[43] = _11071_ ^ _11070_ /*11640*/;
  assign _11072_ = _11071_ & _11070_ /*11639*/;
  assign _11073_ = inv_22[43] & r_21[43] /*11638*/;
  assign _11074_ = _11072_ | _11073_ /*11637*/;
  assign _11075_ = inv_22[44] ^ r_21[44] /*11635*/;
  assign sum_22[44] = _11075_ ^ _11074_ /*11634*/;
  assign _11076_ = _11075_ & _11074_ /*11633*/;
  assign _11077_ = inv_22[44] & r_21[44] /*11632*/;
  assign _11078_ = _11076_ | _11077_ /*11631*/;
  assign _11079_ = inv_22[45] ^ r_21[45] /*11629*/;
  assign sum_22[45] = _11079_ ^ _11078_ /*11628*/;
  assign _11080_ = _11079_ & _11078_ /*11627*/;
  assign _11081_ = inv_22[45] & r_21[45] /*11626*/;
  assign _11082_ = _11080_ | _11081_ /*11625*/;
  assign _11083_ = inv_22[46] ^ r_21[46] /*11623*/;
  assign sum_22[46] = _11083_ ^ _11082_ /*11622*/;
  assign _11084_ = _11083_ & _11082_ /*11621*/;
  assign _11085_ = inv_22[46] & r_21[46] /*11620*/;
  assign _11086_ = _11084_ | _11085_ /*11619*/;
  assign _11087_ = inv_22[47] ^ r_21[47] /*11617*/;
  assign sum_22[47] = _11087_ ^ _11086_ /*11616*/;
  assign _11088_ = _11087_ & _11086_ /*11615*/;
  assign _11089_ = inv_22[47] & r_21[47] /*11614*/;
  assign _11090_ = _11088_ | _11089_ /*11613*/;
  assign _11091_ = inv_22[48] ^ r_21[48] /*11611*/;
  assign sum_22[48] = _11091_ ^ _11090_ /*11610*/;
  assign _11092_ = _11091_ & _11090_ /*11609*/;
  assign _11093_ = inv_22[48] & r_21[48] /*11608*/;
  assign _11094_ = _11092_ | _11093_ /*11607*/;
  assign _11095_ = inv_22[49] ^ r_21[49] /*11605*/;
  assign sum_22[49] = _11095_ ^ _11094_ /*11604*/;
  assign _11096_ = _11095_ & _11094_ /*11603*/;
  assign _11097_ = inv_22[49] & r_21[49] /*11602*/;
  assign _11098_ = _11096_ | _11097_ /*11601*/;
  assign _11099_ = inv_22[50] ^ r_21[50] /*11599*/;
  assign sum_22[50] = _11099_ ^ _11098_ /*11598*/;
  assign _11100_ = _11099_ & _11098_ /*11597*/;
  assign _11101_ = inv_22[50] & r_21[50] /*11596*/;
  assign _11102_ = _11100_ | _11101_ /*11595*/;
  assign _11103_ = inv_22[51] ^ r_21[51] /*11593*/;
  assign sum_22[51] = _11103_ ^ _11102_ /*11592*/;
  assign _11104_ = _11103_ & _11102_ /*11591*/;
  assign _11105_ = inv_22[51] & r_21[51] /*11590*/;
  assign _11106_ = _11104_ | _11105_ /*11589*/;
  assign _11107_ = inv_22[52] ^ r_21[52] /*11587*/;
  assign sum_22[52] = _11107_ ^ _11106_ /*11586*/;
  assign _11108_ = _11107_ & _11106_ /*11585*/;
  assign _11109_ = inv_22[52] & r_21[52] /*11584*/;
  assign _11110_ = _11108_ | _11109_ /*11583*/;
  assign _11111_ = inv_22[53] ^ r_21[53] /*11581*/;
  assign sum_22[53] = _11111_ ^ _11110_ /*11580*/;
  assign _11112_ = _11111_ & _11110_ /*11579*/;
  assign _11113_ = inv_22[53] & r_21[53] /*11578*/;
  assign _11114_ = _11112_ | _11113_ /*11577*/;
  assign _11115_ = inv_22[54] ^ r_21[54] /*11575*/;
  assign sum_22[54] = _11115_ ^ _11114_ /*11574*/;
  assign _11116_ = _11115_ & _11114_ /*11573*/;
  assign _11117_ = inv_22[54] & r_21[54] /*11572*/;
  assign _11118_ = _11116_ | _11117_ /*11571*/;
  assign _11119_ = inv_22[55] ^ r_21[55] /*11569*/;
  assign sum_22[55] = _11119_ ^ _11118_ /*11568*/;
  assign _11120_ = _11119_ & _11118_ /*11567*/;
  assign _11121_ = inv_22[55] & r_21[55] /*11566*/;
  assign _11122_ = _11120_ | _11121_ /*11565*/;
  assign _11123_ = inv_22[56] ^ r_21[56] /*11563*/;
  assign sum_22[56] = _11123_ ^ _11122_ /*11562*/;
  assign _11124_ = _11123_ & _11122_ /*11561*/;
  assign _11125_ = inv_22[56] & r_21[56] /*11560*/;
  assign _11126_ = _11124_ | _11125_ /*11559*/;
  assign _11127_ = inv_22[57] ^ r_21[57] /*11557*/;
  assign sum_22[57] = _11127_ ^ _11126_ /*11556*/;
  assign _11128_ = _11127_ & _11126_ /*11555*/;
  assign _11129_ = inv_22[57] & r_21[57] /*11554*/;
  assign _11130_ = _11128_ | _11129_ /*11553*/;
  assign _11131_ = inv_22[58] ^ r_21[58] /*11551*/;
  assign sum_22[58] = _11131_ ^ _11130_ /*11550*/;
  assign _11132_ = _11131_ & _11130_ /*11549*/;
  assign _11133_ = inv_22[58] & r_21[58] /*11548*/;
  assign _11134_ = _11132_ | _11133_ /*11547*/;
  assign _11135_ = inv_22[59] ^ r_21[59] /*11545*/;
  assign sum_22[59] = _11135_ ^ _11134_ /*11544*/;
  assign _11136_ = _11135_ & _11134_ /*11543*/;
  assign _11137_ = inv_22[59] & r_21[59] /*11542*/;
  assign _11138_ = _11136_ | _11137_ /*11541*/;
  assign _11139_ = inv_22[60] ^ r_21[60] /*11539*/;
  assign sum_22[60] = _11139_ ^ _11138_ /*11538*/;
  assign _11140_ = _11139_ & _11138_ /*11537*/;
  assign _11141_ = inv_22[60] & r_21[60] /*11536*/;
  assign _11142_ = _11140_ | _11141_ /*11535*/;
  assign _11143_ = inv_22[61] ^ r_21[61] /*11533*/;
  assign sum_22[61] = _11143_ ^ _11142_ /*11532*/;
  assign _11144_ = _11143_ & _11142_ /*11531*/;
  assign _11145_ = inv_22[61] & r_21[61] /*11530*/;
  assign _11146_ = _11144_ | _11145_ /*11529*/;
  assign _11147_ = inv_22[62] ^ r_21[62] /*11527*/;
  assign sum_22[62] = _11147_ ^ _11146_ /*11526*/;
  assign _11148_ = _11147_ & _11146_ /*11525*/;
  assign _11149_ = inv_22[62] & r_21[62] /*11524*/;
  assign _11150_ = _11148_ | _11149_ /*11523*/;
  assign _11151_ = inv_22[63] ^ r_21[63] /*11521*/;
  assign sum_22[63] = _11151_ ^ _11150_ /*11520*/;
  assign _11152_ = _11151_ & _11150_ /*11519*/;
  assign _11153_ = inv_22[63] & r_21[63] /*11518*/;
  assign _11154_ = _11152_ | _11153_ /*11517*/;
  assign _11155_ = inv_22[64] ^ r_21[64] /*11515*/;
  assign sum_22[64] = _11155_ ^ _11154_ /*11514*/;
  assign _11156_ = _11155_ & _11154_ /*11513*/;
  assign _11157_ = inv_22[64] & r_21[64] /*11512*/;
  assign _11158_ = _11156_ | _11157_ /*11511*/;
  assign _11159_ = inv_22[65] ^ r_21[65] /*11509*/;
  assign sum_22[65] = _11159_ ^ _11158_ /*11508*/;
  assign _11160_ = _11159_ & _11158_ /*11507*/;
  assign _11161_ = inv_22[65] & r_21[65] /*11506*/;
  assign _11162_ = _11160_ | _11161_ /*11505*/;
  assign _11163_ = inv_22[66] ^ r_21[66] /*11503*/;
  assign sum_22[66] = _11163_ ^ _11162_ /*11502*/;
  assign _11164_ = _11163_ & _11162_ /*11501*/;
  assign _11165_ = inv_22[66] & r_21[66] /*11500*/;
  assign _11166_ = _11164_ | _11165_ /*11499*/;
  assign _11167_ = inv_22[67] ^ r_21[67] /*11497*/;
  assign sum_22[67] = _11167_ ^ _11166_ /*11496*/;
  assign _11168_ = _11167_ & _11166_ /*11495*/;
  assign _11169_ = inv_22[67] & r_21[67] /*11494*/;
  assign _11170_ = _11168_ | _11169_ /*11493*/;
  assign _11171_ = inv_22[68] ^ r_21[68] /*11491*/;
  assign sum_22[68] = _11171_ ^ _11170_ /*11490*/;
  assign _11172_ = _11171_ & _11170_ /*11489*/;
  assign _11173_ = inv_22[68] & r_21[68] /*11488*/;
  assign _11174_ = _11172_ | _11173_ /*11487*/;
  assign _11175_ = inv_22[69] ^ r_21[69] /*11485*/;
  assign sum_22[69] = _11175_ ^ _11174_ /*11484*/;
  assign _11176_ = _11175_ & _11174_ /*11483*/;
  assign _11177_ = inv_22[69] & r_21[69] /*11482*/;
  assign _11178_ = _11176_ | _11177_ /*11481*/;
  assign _11179_ = inv_22[70] ^ r_21[70] /*11479*/;
  assign sum_22[70] = _11179_ ^ _11178_ /*11478*/;
  assign _11180_ = _11179_ & _11178_ /*11477*/;
  assign _11181_ = inv_22[70] & r_21[70] /*11476*/;
  assign _11182_ = _11180_ | _11181_ /*11475*/;
  assign _11183_ = inv_22[71] ^ r_21[71] /*11473*/;
  assign sum_22[71] = _11183_ ^ _11182_ /*11472*/;
  assign _11184_ = _11183_ & _11182_ /*11471*/;
  assign _11185_ = inv_22[71] & r_21[71] /*11470*/;
  assign _11186_ = _11184_ | _11185_ /*11469*/;
  assign _11187_ = inv_22[72] ^ r_21[72] /*11467*/;
  assign sum_22[72] = _11187_ ^ _11186_ /*11466*/;
  assign _11188_ = _11187_ & _11186_ /*11465*/;
  assign _11189_ = inv_22[72] & r_21[72] /*11464*/;
  assign _11190_ = _11188_ | _11189_ /*11463*/;
  assign _11191_ = inv_22[73] ^ r_21[73] /*11461*/;
  assign sum_22[73] = _11191_ ^ _11190_ /*11460*/;
  assign _11192_ = _11191_ & _11190_ /*11459*/;
  assign _11193_ = inv_22[73] & r_21[73] /*11458*/;
  assign _11194_ = _11192_ | _11193_ /*11457*/;
  assign _11195_ = inv_22[74] ^ r_21[74] /*11455*/;
  assign sum_22[74] = _11195_ ^ _11194_ /*11454*/;
  assign _11196_ = _11195_ & _11194_ /*11453*/;
  assign _11197_ = inv_22[74] & r_21[74] /*11452*/;
  assign _11198_ = _11196_ | _11197_ /*11451*/;
  assign _11199_ = inv_22[75] ^ r_21[75] /*11449*/;
  assign sum_22[75] = _11199_ ^ _11198_ /*11448*/;
  assign _11200_ = _11199_ & _11198_ /*11447*/;
  assign _11201_ = inv_22[75] & r_21[75] /*11446*/;
  assign _11202_ = _11200_ | _11201_ /*11445*/;
  assign _11203_ = inv_22[76] ^ r_21[76] /*11443*/;
  assign sum_22[76] = _11203_ ^ _11202_ /*11442*/;
  assign _11204_ = _11203_ & _11202_ /*11441*/;
  assign _11205_ = inv_22[76] & r_21[76] /*11440*/;
  assign _11206_ = _11204_ | _11205_ /*11439*/;
  assign _11207_ = inv_22[77] ^ r_21[77] /*11437*/;
  assign sum_22[77] = _11207_ ^ _11206_ /*11436*/;
  assign _11208_ = _11207_ & _11206_ /*11435*/;
  assign _11209_ = inv_22[77] & r_21[77] /*11434*/;
  assign _11210_ = _11208_ | _11209_ /*11433*/;
  assign _11211_ = inv_22[78] ^ r_21[78] /*11431*/;
  assign sum_22[78] = _11211_ ^ _11210_ /*11430*/;
  assign _11212_ = _11211_ & _11210_ /*11429*/;
  assign _11213_ = inv_22[78] & r_21[78] /*11428*/;
  assign _11214_ = _11212_ | _11213_ /*11427*/;
  assign _11215_ = inv_22[79] ^ r_21[79] /*11425*/;
  assign sum_22[79] = _11215_ ^ _11214_ /*11424*/;
  assign _11216_ = _11215_ & _11214_ /*11423*/;
  assign _11217_ = inv_22[79] & r_21[79] /*11422*/;
  assign _11218_ = _11216_ | _11217_ /*11421*/;
  assign _11219_ = inv_22[80] ^ r_21[80] /*11419*/;
  assign sum_22[80] = _11219_ ^ _11218_ /*11418*/;
  assign _11220_ = _11219_ & _11218_ /*11417*/;
  assign _11221_ = inv_22[80] & r_21[80] /*11416*/;
  assign _11222_ = _11220_ | _11221_ /*11415*/;
  assign _11223_ = inv_22[81] ^ r_21[81] /*11413*/;
  assign sum_22[81] = _11223_ ^ _11222_ /*11412*/;
  assign _11224_ = _11223_ & _11222_ /*11411*/;
  assign _11225_ = inv_22[81] & r_21[81] /*11410*/;
  assign _11226_ = _11224_ | _11225_ /*11409*/;
  assign _11227_ = inv_22[82] ^ r_21[82] /*11407*/;
  assign sum_22[82] = _11227_ ^ _11226_ /*11406*/;
  assign _11228_ = _11227_ & _11226_ /*11405*/;
  assign _11229_ = inv_22[82] & r_21[82] /*11404*/;
  assign _11230_ = _11228_ | _11229_ /*11403*/;
  assign _11231_ = inv_22[83] ^ r_21[83] /*11401*/;
  assign sum_22[83] = _11231_ ^ _11230_ /*11400*/;
  assign _11232_ = _11231_ & _11230_ /*11399*/;
  assign _11233_ = inv_22[83] & r_21[83] /*11398*/;
  assign _11234_ = _11232_ | _11233_ /*11397*/;
  assign _11235_ = _11234_ ^ _11230_ /*11396*/;
  assign _11236_ = ~_11235_ /*11395*/;
  assign _11237_ = sum_22[83] & _11236_ /*11394*/;
  assign _11238_ = _11235_ & _11234_ /*11393*/;
  assign sum_22[84] = _11238_ | _11237_ /*11392*/;
  assign q[10] = ~sum_22[84] /*11391*/;
  assign m_22[0] = r_21[0] /*11390*/;
  assign m_22[1] = r_21[1] /*11389*/;
  assign m_22[2] = r_21[2] /*11388*/;
  assign m_22[3] = r_21[3] /*11387*/;
  assign m_22[4] = r_21[4] /*11386*/;
  assign m_22[5] = r_21[5] /*11385*/;
  assign m_22[6] = r_21[6] /*11384*/;
  assign m_22[7] = r_21[7] /*11383*/;
  assign m_22[8] = r_21[8] /*11382*/;
  assign m_22[9] = r_21[9] /*11381*/;
  assign m_22[10] = r_21[10] /*11380*/;
  assign m_22[11] = r_21[11] /*11379*/;
  assign m_22[12] = r_21[12] /*11378*/;
  assign m_22[13] = r_21[13] /*11377*/;
  assign m_22[14] = r_21[14] /*11376*/;
  assign m_22[15] = r_21[15] /*11375*/;
  assign m_22[16] = r_21[16] /*11374*/;
  assign m_22[17] = r_21[17] /*11373*/;
  assign m_22[18] = r_21[18] /*11372*/;
  assign m_22[19] = r_21[19] /*11371*/;
  assign m_22[20] = r_21[20] /*11370*/;
  assign m_22[21] = r_21[21] /*11369*/;
  assign m_22[22] = r_21[22] /*11368*/;
  assign m_22[23] = r_21[23] /*11367*/;
  assign m_22[24] = r_21[24] /*11366*/;
  assign m_22[25] = r_21[25] /*11365*/;
  assign m_22[26] = r_21[26] /*11364*/;
  assign m_22[27] = r_21[27] /*11363*/;
  assign m_22[28] = r_21[28] /*11362*/;
  assign m_22[29] = r_21[29] /*11361*/;
  assign m_22[30] = r_21[30] /*11360*/;
  assign m_22[31] = r_21[31] /*11359*/;
  assign m_22[32] = r_21[32] /*11358*/;
  assign m_22[33] = r_21[33] /*11357*/;
  assign m_22[34] = r_21[34] /*11356*/;
  assign m_22[35] = r_21[35] /*11355*/;
  assign m_22[36] = r_21[36] /*11354*/;
  assign m_22[37] = r_21[37] /*11353*/;
  assign m_22[38] = r_21[38] /*11352*/;
  assign m_22[39] = r_21[39] /*11351*/;
  assign m_22[40] = r_21[40] /*11350*/;
  assign m_22[41] = r_21[41] /*11349*/;
  assign m_22[42] = r_21[42] /*11348*/;
  assign m_22[43] = r_21[43] /*11347*/;
  assign m_22[44] = r_21[44] /*11346*/;
  assign m_22[45] = r_21[45] /*11345*/;
  assign m_22[46] = r_21[46] /*11344*/;
  assign m_22[47] = r_21[47] /*11343*/;
  assign m_22[48] = r_21[48] /*11342*/;
  assign m_22[49] = r_21[49] /*11341*/;
  assign m_22[50] = r_21[50] /*11340*/;
  assign m_22[51] = r_21[51] /*11339*/;
  assign m_22[52] = r_21[52] /*11338*/;
  assign m_22[53] = r_21[53] /*11337*/;
  assign m_22[54] = r_21[54] /*11336*/;
  assign m_22[55] = r_21[55] /*11335*/;
  assign m_22[56] = r_21[56] /*11334*/;
  assign m_22[57] = r_21[57] /*11333*/;
  assign m_22[58] = r_21[58] /*11332*/;
  assign m_22[59] = r_21[59] /*11331*/;
  assign m_22[60] = r_21[60] /*11330*/;
  assign m_22[61] = r_21[61] /*11329*/;
  assign m_22[62] = r_21[62] /*11328*/;
  assign m_22[63] = r_21[63] /*11327*/;
  assign m_22[64] = r_21[64] /*11326*/;
  assign m_22[65] = r_21[65] /*11325*/;
  assign m_22[66] = r_21[66] /*11324*/;
  assign m_22[67] = r_21[67] /*11323*/;
  assign m_22[68] = r_21[68] /*11322*/;
  assign m_22[69] = r_21[69] /*11321*/;
  assign m_22[70] = r_21[70] /*11320*/;
  assign m_22[71] = r_21[71] /*11319*/;
  assign m_22[72] = r_21[72] /*11318*/;
  assign m_22[73] = r_21[73] /*11317*/;
  assign m_22[74] = r_21[74] /*11316*/;
  assign m_22[75] = r_21[75] /*11315*/;
  assign m_22[76] = r_21[76] /*11314*/;
  assign m_22[77] = r_21[77] /*11313*/;
  assign m_22[78] = r_21[78] /*11312*/;
  assign m_22[79] = r_21[79] /*11311*/;
  assign m_22[80] = r_21[80] /*11310*/;
  assign m_22[81] = r_21[81] /*11309*/;
  assign m_22[82] = r_21[82] /*11308*/;
  assign m_22[83] = r_21[83] /*11307*/;
  assign m_22[84] = r_21[83] /*11306*/;
  assign _11240_ = ~q[10] /*11305*/;
  assign _11241_ = sum_22[0] & q[10] /*11304*/;
  assign _11242_ = m_22[0] & _11240_ /*11303*/;
  assign r_22[0] = _11242_ | _11241_ /*11302*/;
  assign _11243_ = ~q[10] /*11301*/;
  assign _11244_ = sum_22[1] & q[10] /*11300*/;
  assign _11245_ = m_22[1] & _11243_ /*11299*/;
  assign r_22[1] = _11245_ | _11244_ /*11298*/;
  assign _11246_ = ~q[10] /*11297*/;
  assign _11247_ = sum_22[2] & q[10] /*11296*/;
  assign _11248_ = m_22[2] & _11246_ /*11295*/;
  assign r_22[2] = _11248_ | _11247_ /*11294*/;
  assign _11249_ = ~q[10] /*11293*/;
  assign _11250_ = sum_22[3] & q[10] /*11292*/;
  assign _11251_ = m_22[3] & _11249_ /*11291*/;
  assign r_22[3] = _11251_ | _11250_ /*11290*/;
  assign _11252_ = ~q[10] /*11289*/;
  assign _11253_ = sum_22[4] & q[10] /*11288*/;
  assign _11254_ = m_22[4] & _11252_ /*11287*/;
  assign r_22[4] = _11254_ | _11253_ /*11286*/;
  assign _11255_ = ~q[10] /*11285*/;
  assign _11256_ = sum_22[5] & q[10] /*11284*/;
  assign _11257_ = m_22[5] & _11255_ /*11283*/;
  assign r_22[5] = _11257_ | _11256_ /*11282*/;
  assign _11258_ = ~q[10] /*11281*/;
  assign _11259_ = sum_22[6] & q[10] /*11280*/;
  assign _11260_ = m_22[6] & _11258_ /*11279*/;
  assign r_22[6] = _11260_ | _11259_ /*11278*/;
  assign _11261_ = ~q[10] /*11277*/;
  assign _11262_ = sum_22[7] & q[10] /*11276*/;
  assign _11263_ = m_22[7] & _11261_ /*11275*/;
  assign r_22[7] = _11263_ | _11262_ /*11274*/;
  assign _11264_ = ~q[10] /*11273*/;
  assign _11265_ = sum_22[8] & q[10] /*11272*/;
  assign _11266_ = m_22[8] & _11264_ /*11271*/;
  assign r_22[8] = _11266_ | _11265_ /*11270*/;
  assign _11267_ = ~q[10] /*11269*/;
  assign _11268_ = sum_22[9] & q[10] /*11268*/;
  assign _11269_ = m_22[9] & _11267_ /*11267*/;
  assign r_22[9] = _11269_ | _11268_ /*11266*/;
  assign _11270_ = ~q[10] /*11265*/;
  assign _11271_ = sum_22[10] & q[10] /*11264*/;
  assign _11272_ = m_22[10] & _11270_ /*11263*/;
  assign r_22[10] = _11272_ | _11271_ /*11262*/;
  assign _11273_ = ~q[10] /*11261*/;
  assign _11274_ = sum_22[11] & q[10] /*11260*/;
  assign _11275_ = m_22[11] & _11273_ /*11259*/;
  assign r_22[11] = _11275_ | _11274_ /*11258*/;
  assign _11276_ = ~q[10] /*11257*/;
  assign _11277_ = sum_22[12] & q[10] /*11256*/;
  assign _11278_ = m_22[12] & _11276_ /*11255*/;
  assign r_22[12] = _11278_ | _11277_ /*11254*/;
  assign _11279_ = ~q[10] /*11253*/;
  assign _11280_ = sum_22[13] & q[10] /*11252*/;
  assign _11281_ = m_22[13] & _11279_ /*11251*/;
  assign r_22[13] = _11281_ | _11280_ /*11250*/;
  assign _11282_ = ~q[10] /*11249*/;
  assign _11283_ = sum_22[14] & q[10] /*11248*/;
  assign _11284_ = m_22[14] & _11282_ /*11247*/;
  assign r_22[14] = _11284_ | _11283_ /*11246*/;
  assign _11285_ = ~q[10] /*11245*/;
  assign _11286_ = sum_22[15] & q[10] /*11244*/;
  assign _11287_ = m_22[15] & _11285_ /*11243*/;
  assign r_22[15] = _11287_ | _11286_ /*11242*/;
  assign _11288_ = ~q[10] /*11241*/;
  assign _11289_ = sum_22[16] & q[10] /*11240*/;
  assign _11290_ = m_22[16] & _11288_ /*11239*/;
  assign r_22[16] = _11290_ | _11289_ /*11238*/;
  assign _11291_ = ~q[10] /*11237*/;
  assign _11292_ = sum_22[17] & q[10] /*11236*/;
  assign _11293_ = m_22[17] & _11291_ /*11235*/;
  assign r_22[17] = _11293_ | _11292_ /*11234*/;
  assign _11294_ = ~q[10] /*11233*/;
  assign _11295_ = sum_22[18] & q[10] /*11232*/;
  assign _11296_ = m_22[18] & _11294_ /*11231*/;
  assign r_22[18] = _11296_ | _11295_ /*11230*/;
  assign _11297_ = ~q[10] /*11229*/;
  assign _11298_ = sum_22[19] & q[10] /*11228*/;
  assign _11299_ = m_22[19] & _11297_ /*11227*/;
  assign r_22[19] = _11299_ | _11298_ /*11226*/;
  assign _11300_ = ~q[10] /*11225*/;
  assign _11301_ = sum_22[20] & q[10] /*11224*/;
  assign _11302_ = m_22[20] & _11300_ /*11223*/;
  assign r_22[20] = _11302_ | _11301_ /*11222*/;
  assign _11303_ = ~q[10] /*11221*/;
  assign _11304_ = sum_22[21] & q[10] /*11220*/;
  assign _11305_ = m_22[21] & _11303_ /*11219*/;
  assign r_22[21] = _11305_ | _11304_ /*11218*/;
  assign _11306_ = ~q[10] /*11217*/;
  assign _11307_ = sum_22[22] & q[10] /*11216*/;
  assign _11308_ = m_22[22] & _11306_ /*11215*/;
  assign r_22[22] = _11308_ | _11307_ /*11214*/;
  assign _11309_ = ~q[10] /*11213*/;
  assign _11310_ = sum_22[23] & q[10] /*11212*/;
  assign _11311_ = m_22[23] & _11309_ /*11211*/;
  assign r_22[23] = _11311_ | _11310_ /*11210*/;
  assign _11312_ = ~q[10] /*11209*/;
  assign _11313_ = sum_22[24] & q[10] /*11208*/;
  assign _11314_ = m_22[24] & _11312_ /*11207*/;
  assign r_22[24] = _11314_ | _11313_ /*11206*/;
  assign _11315_ = ~q[10] /*11205*/;
  assign _11316_ = sum_22[25] & q[10] /*11204*/;
  assign _11317_ = m_22[25] & _11315_ /*11203*/;
  assign r_22[25] = _11317_ | _11316_ /*11202*/;
  assign _11318_ = ~q[10] /*11201*/;
  assign _11319_ = sum_22[26] & q[10] /*11200*/;
  assign _11320_ = m_22[26] & _11318_ /*11199*/;
  assign r_22[26] = _11320_ | _11319_ /*11198*/;
  assign _11321_ = ~q[10] /*11197*/;
  assign _11322_ = sum_22[27] & q[10] /*11196*/;
  assign _11323_ = m_22[27] & _11321_ /*11195*/;
  assign r_22[27] = _11323_ | _11322_ /*11194*/;
  assign _11324_ = ~q[10] /*11193*/;
  assign _11325_ = sum_22[28] & q[10] /*11192*/;
  assign _11326_ = m_22[28] & _11324_ /*11191*/;
  assign r_22[28] = _11326_ | _11325_ /*11190*/;
  assign _11327_ = ~q[10] /*11189*/;
  assign _11328_ = sum_22[29] & q[10] /*11188*/;
  assign _11329_ = m_22[29] & _11327_ /*11187*/;
  assign r_22[29] = _11329_ | _11328_ /*11186*/;
  assign _11330_ = ~q[10] /*11185*/;
  assign _11331_ = sum_22[30] & q[10] /*11184*/;
  assign _11332_ = m_22[30] & _11330_ /*11183*/;
  assign r_22[30] = _11332_ | _11331_ /*11182*/;
  assign _11333_ = ~q[10] /*11181*/;
  assign _11334_ = sum_22[31] & q[10] /*11180*/;
  assign _11335_ = m_22[31] & _11333_ /*11179*/;
  assign r_22[31] = _11335_ | _11334_ /*11178*/;
  assign _11336_ = ~q[10] /*11177*/;
  assign _11337_ = sum_22[32] & q[10] /*11176*/;
  assign _11338_ = m_22[32] & _11336_ /*11175*/;
  assign r_22[32] = _11338_ | _11337_ /*11174*/;
  assign _11339_ = ~q[10] /*11173*/;
  assign _11340_ = sum_22[33] & q[10] /*11172*/;
  assign _11341_ = m_22[33] & _11339_ /*11171*/;
  assign r_22[33] = _11341_ | _11340_ /*11170*/;
  assign _11342_ = ~q[10] /*11169*/;
  assign _11343_ = sum_22[34] & q[10] /*11168*/;
  assign _11344_ = m_22[34] & _11342_ /*11167*/;
  assign r_22[34] = _11344_ | _11343_ /*11166*/;
  assign _11345_ = ~q[10] /*11165*/;
  assign _11346_ = sum_22[35] & q[10] /*11164*/;
  assign _11347_ = m_22[35] & _11345_ /*11163*/;
  assign r_22[35] = _11347_ | _11346_ /*11162*/;
  assign _11348_ = ~q[10] /*11161*/;
  assign _11349_ = sum_22[36] & q[10] /*11160*/;
  assign _11350_ = m_22[36] & _11348_ /*11159*/;
  assign r_22[36] = _11350_ | _11349_ /*11158*/;
  assign _11351_ = ~q[10] /*11157*/;
  assign _11352_ = sum_22[37] & q[10] /*11156*/;
  assign _11353_ = m_22[37] & _11351_ /*11155*/;
  assign r_22[37] = _11353_ | _11352_ /*11154*/;
  assign _11354_ = ~q[10] /*11153*/;
  assign _11355_ = sum_22[38] & q[10] /*11152*/;
  assign _11356_ = m_22[38] & _11354_ /*11151*/;
  assign r_22[38] = _11356_ | _11355_ /*11150*/;
  assign _11357_ = ~q[10] /*11149*/;
  assign _11358_ = sum_22[39] & q[10] /*11148*/;
  assign _11359_ = m_22[39] & _11357_ /*11147*/;
  assign r_22[39] = _11359_ | _11358_ /*11146*/;
  assign _11360_ = ~q[10] /*11145*/;
  assign _11361_ = sum_22[40] & q[10] /*11144*/;
  assign _11362_ = m_22[40] & _11360_ /*11143*/;
  assign r_22[40] = _11362_ | _11361_ /*11142*/;
  assign _11363_ = ~q[10] /*11141*/;
  assign _11364_ = sum_22[41] & q[10] /*11140*/;
  assign _11365_ = m_22[41] & _11363_ /*11139*/;
  assign r_22[41] = _11365_ | _11364_ /*11138*/;
  assign _11366_ = ~q[10] /*11137*/;
  assign _11367_ = sum_22[42] & q[10] /*11136*/;
  assign _11368_ = m_22[42] & _11366_ /*11135*/;
  assign r_22[42] = _11368_ | _11367_ /*11134*/;
  assign _11369_ = ~q[10] /*11133*/;
  assign _11370_ = sum_22[43] & q[10] /*11132*/;
  assign _11371_ = m_22[43] & _11369_ /*11131*/;
  assign r_22[43] = _11371_ | _11370_ /*11130*/;
  assign _11372_ = ~q[10] /*11129*/;
  assign _11373_ = sum_22[44] & q[10] /*11128*/;
  assign _11374_ = m_22[44] & _11372_ /*11127*/;
  assign r_22[44] = _11374_ | _11373_ /*11126*/;
  assign _11375_ = ~q[10] /*11125*/;
  assign _11376_ = sum_22[45] & q[10] /*11124*/;
  assign _11377_ = m_22[45] & _11375_ /*11123*/;
  assign r_22[45] = _11377_ | _11376_ /*11122*/;
  assign _11378_ = ~q[10] /*11121*/;
  assign _11379_ = sum_22[46] & q[10] /*11120*/;
  assign _11380_ = m_22[46] & _11378_ /*11119*/;
  assign r_22[46] = _11380_ | _11379_ /*11118*/;
  assign _11381_ = ~q[10] /*11117*/;
  assign _11382_ = sum_22[47] & q[10] /*11116*/;
  assign _11383_ = m_22[47] & _11381_ /*11115*/;
  assign r_22[47] = _11383_ | _11382_ /*11114*/;
  assign _11384_ = ~q[10] /*11113*/;
  assign _11385_ = sum_22[48] & q[10] /*11112*/;
  assign _11386_ = m_22[48] & _11384_ /*11111*/;
  assign r_22[48] = _11386_ | _11385_ /*11110*/;
  assign _11387_ = ~q[10] /*11109*/;
  assign _11388_ = sum_22[49] & q[10] /*11108*/;
  assign _11389_ = m_22[49] & _11387_ /*11107*/;
  assign r_22[49] = _11389_ | _11388_ /*11106*/;
  assign _11390_ = ~q[10] /*11105*/;
  assign _11391_ = sum_22[50] & q[10] /*11104*/;
  assign _11392_ = m_22[50] & _11390_ /*11103*/;
  assign r_22[50] = _11392_ | _11391_ /*11102*/;
  assign _11393_ = ~q[10] /*11101*/;
  assign _11394_ = sum_22[51] & q[10] /*11100*/;
  assign _11395_ = m_22[51] & _11393_ /*11099*/;
  assign r_22[51] = _11395_ | _11394_ /*11098*/;
  assign _11396_ = ~q[10] /*11097*/;
  assign _11397_ = sum_22[52] & q[10] /*11096*/;
  assign _11398_ = m_22[52] & _11396_ /*11095*/;
  assign r_22[52] = _11398_ | _11397_ /*11094*/;
  assign _11399_ = ~q[10] /*11093*/;
  assign _11400_ = sum_22[53] & q[10] /*11092*/;
  assign _11401_ = m_22[53] & _11399_ /*11091*/;
  assign r_22[53] = _11401_ | _11400_ /*11090*/;
  assign _11402_ = ~q[10] /*11089*/;
  assign _11403_ = sum_22[54] & q[10] /*11088*/;
  assign _11404_ = m_22[54] & _11402_ /*11087*/;
  assign r_22[54] = _11404_ | _11403_ /*11086*/;
  assign _11405_ = ~q[10] /*11085*/;
  assign _11406_ = sum_22[55] & q[10] /*11084*/;
  assign _11407_ = m_22[55] & _11405_ /*11083*/;
  assign r_22[55] = _11407_ | _11406_ /*11082*/;
  assign _11408_ = ~q[10] /*11081*/;
  assign _11409_ = sum_22[56] & q[10] /*11080*/;
  assign _11410_ = m_22[56] & _11408_ /*11079*/;
  assign r_22[56] = _11410_ | _11409_ /*11078*/;
  assign _11411_ = ~q[10] /*11077*/;
  assign _11412_ = sum_22[57] & q[10] /*11076*/;
  assign _11413_ = m_22[57] & _11411_ /*11075*/;
  assign r_22[57] = _11413_ | _11412_ /*11074*/;
  assign _11414_ = ~q[10] /*11073*/;
  assign _11415_ = sum_22[58] & q[10] /*11072*/;
  assign _11416_ = m_22[58] & _11414_ /*11071*/;
  assign r_22[58] = _11416_ | _11415_ /*11070*/;
  assign _11417_ = ~q[10] /*11069*/;
  assign _11418_ = sum_22[59] & q[10] /*11068*/;
  assign _11419_ = m_22[59] & _11417_ /*11067*/;
  assign r_22[59] = _11419_ | _11418_ /*11066*/;
  assign _11420_ = ~q[10] /*11065*/;
  assign _11421_ = sum_22[60] & q[10] /*11064*/;
  assign _11422_ = m_22[60] & _11420_ /*11063*/;
  assign r_22[60] = _11422_ | _11421_ /*11062*/;
  assign _11423_ = ~q[10] /*11061*/;
  assign _11424_ = sum_22[61] & q[10] /*11060*/;
  assign _11425_ = m_22[61] & _11423_ /*11059*/;
  assign r_22[61] = _11425_ | _11424_ /*11058*/;
  assign _11426_ = ~q[10] /*11057*/;
  assign _11427_ = sum_22[62] & q[10] /*11056*/;
  assign _11428_ = m_22[62] & _11426_ /*11055*/;
  assign r_22[62] = _11428_ | _11427_ /*11054*/;
  assign _11429_ = ~q[10] /*11053*/;
  assign _11430_ = sum_22[63] & q[10] /*11052*/;
  assign _11431_ = m_22[63] & _11429_ /*11051*/;
  assign r_22[63] = _11431_ | _11430_ /*11050*/;
  assign _11432_ = ~q[10] /*11049*/;
  assign _11433_ = sum_22[64] & q[10] /*11048*/;
  assign _11434_ = m_22[64] & _11432_ /*11047*/;
  assign r_22[64] = _11434_ | _11433_ /*11046*/;
  assign _11435_ = ~q[10] /*11045*/;
  assign _11436_ = sum_22[65] & q[10] /*11044*/;
  assign _11437_ = m_22[65] & _11435_ /*11043*/;
  assign r_22[65] = _11437_ | _11436_ /*11042*/;
  assign _11438_ = ~q[10] /*11041*/;
  assign _11439_ = sum_22[66] & q[10] /*11040*/;
  assign _11440_ = m_22[66] & _11438_ /*11039*/;
  assign r_22[66] = _11440_ | _11439_ /*11038*/;
  assign _11441_ = ~q[10] /*11037*/;
  assign _11442_ = sum_22[67] & q[10] /*11036*/;
  assign _11443_ = m_22[67] & _11441_ /*11035*/;
  assign r_22[67] = _11443_ | _11442_ /*11034*/;
  assign _11444_ = ~q[10] /*11033*/;
  assign _11445_ = sum_22[68] & q[10] /*11032*/;
  assign _11446_ = m_22[68] & _11444_ /*11031*/;
  assign r_22[68] = _11446_ | _11445_ /*11030*/;
  assign _11447_ = ~q[10] /*11029*/;
  assign _11448_ = sum_22[69] & q[10] /*11028*/;
  assign _11449_ = m_22[69] & _11447_ /*11027*/;
  assign r_22[69] = _11449_ | _11448_ /*11026*/;
  assign _11450_ = ~q[10] /*11025*/;
  assign _11451_ = sum_22[70] & q[10] /*11024*/;
  assign _11452_ = m_22[70] & _11450_ /*11023*/;
  assign r_22[70] = _11452_ | _11451_ /*11022*/;
  assign _11453_ = ~q[10] /*11021*/;
  assign _11454_ = sum_22[71] & q[10] /*11020*/;
  assign _11455_ = m_22[71] & _11453_ /*11019*/;
  assign r_22[71] = _11455_ | _11454_ /*11018*/;
  assign _11456_ = ~q[10] /*11017*/;
  assign _11457_ = sum_22[72] & q[10] /*11016*/;
  assign _11458_ = m_22[72] & _11456_ /*11015*/;
  assign r_22[72] = _11458_ | _11457_ /*11014*/;
  assign _11459_ = ~q[10] /*11013*/;
  assign _11460_ = sum_22[73] & q[10] /*11012*/;
  assign _11461_ = m_22[73] & _11459_ /*11011*/;
  assign r_22[73] = _11461_ | _11460_ /*11010*/;
  assign _11462_ = ~q[10] /*11009*/;
  assign _11463_ = sum_22[74] & q[10] /*11008*/;
  assign _11464_ = m_22[74] & _11462_ /*11007*/;
  assign r_22[74] = _11464_ | _11463_ /*11006*/;
  assign _11465_ = ~q[10] /*11005*/;
  assign _11466_ = sum_22[75] & q[10] /*11004*/;
  assign _11467_ = m_22[75] & _11465_ /*11003*/;
  assign r_22[75] = _11467_ | _11466_ /*11002*/;
  assign _11468_ = ~q[10] /*11001*/;
  assign _11469_ = sum_22[76] & q[10] /*11000*/;
  assign _11470_ = m_22[76] & _11468_ /*10999*/;
  assign r_22[76] = _11470_ | _11469_ /*10998*/;
  assign _11471_ = ~q[10] /*10997*/;
  assign _11472_ = sum_22[77] & q[10] /*10996*/;
  assign _11473_ = m_22[77] & _11471_ /*10995*/;
  assign r_22[77] = _11473_ | _11472_ /*10994*/;
  assign _11474_ = ~q[10] /*10993*/;
  assign _11475_ = sum_22[78] & q[10] /*10992*/;
  assign _11476_ = m_22[78] & _11474_ /*10991*/;
  assign r_22[78] = _11476_ | _11475_ /*10990*/;
  assign _11477_ = ~q[10] /*10989*/;
  assign _11478_ = sum_22[79] & q[10] /*10988*/;
  assign _11479_ = m_22[79] & _11477_ /*10987*/;
  assign r_22[79] = _11479_ | _11478_ /*10986*/;
  assign _11480_ = ~q[10] /*10985*/;
  assign _11481_ = sum_22[80] & q[10] /*10984*/;
  assign _11482_ = m_22[80] & _11480_ /*10983*/;
  assign r_22[80] = _11482_ | _11481_ /*10982*/;
  assign _11483_ = ~q[10] /*10981*/;
  assign _11484_ = sum_22[81] & q[10] /*10980*/;
  assign _11485_ = m_22[81] & _11483_ /*10979*/;
  assign r_22[81] = _11485_ | _11484_ /*10978*/;
  assign _11486_ = ~q[10] /*10977*/;
  assign _11487_ = sum_22[82] & q[10] /*10976*/;
  assign _11488_ = m_22[82] & _11486_ /*10975*/;
  assign r_22[82] = _11488_ | _11487_ /*10974*/;
  assign _11489_ = ~q[10] /*10973*/;
  assign _11490_ = sum_22[83] & q[10] /*10972*/;
  assign _11491_ = m_22[83] & _11489_ /*10971*/;
  assign r_22[83] = _11491_ | _11490_ /*10970*/;
  assign _11492_ = ~q[10] /*10969*/;
  assign _11493_ = sum_22[84] & q[10] /*10968*/;
  assign _11494_ = m_22[84] & _11492_ /*10967*/;
  assign r_22[84] = _11494_ | _11493_ /*10966*/;
  assign inv_23[0] = oneWire /*10824*/;
  assign inv_23[1] = oneWire /*10818*/;
  assign inv_23[2] = oneWire /*10812*/;
  assign inv_23[3] = oneWire /*10806*/;
  assign inv_23[4] = oneWire /*10800*/;
  assign inv_23[5] = oneWire /*10794*/;
  assign inv_23[6] = oneWire /*10788*/;
  assign inv_23[7] = oneWire /*10782*/;
  assign inv_23[8] = oneWire /*10776*/;
  assign inv_23[9] = ~div[0] /*10770*/;
  assign inv_23[10] = ~div[1] /*10764*/;
  assign inv_23[11] = ~div[2] /*10758*/;
  assign inv_23[12] = ~div[3] /*10752*/;
  assign inv_23[13] = ~div[4] /*10746*/;
  assign inv_23[14] = ~div[5] /*10740*/;
  assign inv_23[15] = ~div[6] /*10734*/;
  assign inv_23[16] = ~div[7] /*10728*/;
  assign inv_23[17] = ~div[8] /*10722*/;
  assign inv_23[18] = ~div[9] /*10716*/;
  assign inv_23[19] = ~div[10] /*10710*/;
  assign inv_23[20] = ~div[11] /*10704*/;
  assign inv_23[21] = ~div[12] /*10698*/;
  assign inv_23[22] = ~div[13] /*10692*/;
  assign inv_23[23] = ~div[14] /*10686*/;
  assign inv_23[24] = ~div[15] /*10680*/;
  assign inv_23[25] = ~div[16] /*10674*/;
  assign inv_23[26] = ~div[17] /*10668*/;
  assign inv_23[27] = ~div[18] /*10662*/;
  assign inv_23[28] = ~div[19] /*10656*/;
  assign inv_23[29] = ~div[20] /*10650*/;
  assign inv_23[30] = ~div[21] /*10644*/;
  assign inv_23[31] = ~div[22] /*10638*/;
  assign inv_23[32] = ~div[23] /*10632*/;
  assign inv_23[33] = ~div[24] /*10626*/;
  assign inv_23[34] = ~div[25] /*10620*/;
  assign inv_23[35] = ~div[26] /*10614*/;
  assign inv_23[36] = ~div[27] /*10608*/;
  assign inv_23[37] = ~div[28] /*10602*/;
  assign inv_23[38] = ~div[29] /*10596*/;
  assign inv_23[39] = ~div[30] /*10590*/;
  assign inv_23[40] = oneWire /*10584*/;
  assign inv_23[41] = oneWire /*10578*/;
  assign inv_23[42] = oneWire /*10572*/;
  assign inv_23[43] = oneWire /*10566*/;
  assign inv_23[44] = oneWire /*10560*/;
  assign inv_23[45] = oneWire /*10554*/;
  assign inv_23[46] = oneWire /*10548*/;
  assign inv_23[47] = oneWire /*10542*/;
  assign inv_23[48] = oneWire /*10536*/;
  assign inv_23[49] = oneWire /*10530*/;
  assign inv_23[50] = oneWire /*10524*/;
  assign inv_23[51] = oneWire /*10518*/;
  assign inv_23[52] = oneWire /*10512*/;
  assign inv_23[53] = oneWire /*10506*/;
  assign inv_23[54] = oneWire /*10500*/;
  assign inv_23[55] = oneWire /*10494*/;
  assign inv_23[56] = oneWire /*10488*/;
  assign inv_23[57] = oneWire /*10482*/;
  assign inv_23[58] = oneWire /*10476*/;
  assign inv_23[59] = oneWire /*10470*/;
  assign inv_23[60] = oneWire /*10464*/;
  assign inv_23[61] = oneWire /*10458*/;
  assign inv_23[62] = oneWire /*10452*/;
  assign inv_23[63] = oneWire /*10446*/;
  assign inv_23[64] = oneWire /*10440*/;
  assign inv_23[65] = oneWire /*10434*/;
  assign inv_23[66] = oneWire /*10428*/;
  assign inv_23[67] = oneWire /*10422*/;
  assign inv_23[68] = oneWire /*10416*/;
  assign inv_23[69] = oneWire /*10410*/;
  assign inv_23[70] = oneWire /*10404*/;
  assign inv_23[71] = oneWire /*10398*/;
  assign inv_23[72] = oneWire /*10392*/;
  assign inv_23[73] = oneWire /*10386*/;
  assign inv_23[74] = oneWire /*10380*/;
  assign inv_23[75] = oneWire /*10374*/;
  assign inv_23[76] = oneWire /*10368*/;
  assign inv_23[77] = oneWire /*10362*/;
  assign inv_23[78] = oneWire /*10356*/;
  assign inv_23[79] = oneWire /*10350*/;
  assign inv_23[80] = oneWire /*10344*/;
  assign inv_23[81] = oneWire /*10338*/;
  assign inv_23[82] = oneWire /*10332*/;
  assign inv_23[83] = oneWire /*10326*/;
  assign inv_23[84] = oneWire /*10320*/;
  assign _11495_ = inv_23[0] ^ r_22[0] /*10823*/;
  assign sum_23[0] = _11495_ ^ oneWire /*10822*/;
  assign _11496_ = _11495_ & oneWire /*10821*/;
  assign _11497_ = inv_23[0] & r_22[0] /*10820*/;
  assign _11498_ = _11496_ | _11497_ /*10819*/;
  assign _11499_ = inv_23[1] ^ r_22[1] /*10817*/;
  assign sum_23[1] = _11499_ ^ _11498_ /*10816*/;
  assign _11500_ = _11499_ & _11498_ /*10815*/;
  assign _11501_ = inv_23[1] & r_22[1] /*10814*/;
  assign _11502_ = _11500_ | _11501_ /*10813*/;
  assign _11503_ = inv_23[2] ^ r_22[2] /*10811*/;
  assign sum_23[2] = _11503_ ^ _11502_ /*10810*/;
  assign _11504_ = _11503_ & _11502_ /*10809*/;
  assign _11505_ = inv_23[2] & r_22[2] /*10808*/;
  assign _11506_ = _11504_ | _11505_ /*10807*/;
  assign _11507_ = inv_23[3] ^ r_22[3] /*10805*/;
  assign sum_23[3] = _11507_ ^ _11506_ /*10804*/;
  assign _11508_ = _11507_ & _11506_ /*10803*/;
  assign _11509_ = inv_23[3] & r_22[3] /*10802*/;
  assign _11510_ = _11508_ | _11509_ /*10801*/;
  assign _11511_ = inv_23[4] ^ r_22[4] /*10799*/;
  assign sum_23[4] = _11511_ ^ _11510_ /*10798*/;
  assign _11512_ = _11511_ & _11510_ /*10797*/;
  assign _11513_ = inv_23[4] & r_22[4] /*10796*/;
  assign _11514_ = _11512_ | _11513_ /*10795*/;
  assign _11515_ = inv_23[5] ^ r_22[5] /*10793*/;
  assign sum_23[5] = _11515_ ^ _11514_ /*10792*/;
  assign _11516_ = _11515_ & _11514_ /*10791*/;
  assign _11517_ = inv_23[5] & r_22[5] /*10790*/;
  assign _11518_ = _11516_ | _11517_ /*10789*/;
  assign _11519_ = inv_23[6] ^ r_22[6] /*10787*/;
  assign sum_23[6] = _11519_ ^ _11518_ /*10786*/;
  assign _11520_ = _11519_ & _11518_ /*10785*/;
  assign _11521_ = inv_23[6] & r_22[6] /*10784*/;
  assign _11522_ = _11520_ | _11521_ /*10783*/;
  assign _11523_ = inv_23[7] ^ r_22[7] /*10781*/;
  assign sum_23[7] = _11523_ ^ _11522_ /*10780*/;
  assign _11524_ = _11523_ & _11522_ /*10779*/;
  assign _11525_ = inv_23[7] & r_22[7] /*10778*/;
  assign _11526_ = _11524_ | _11525_ /*10777*/;
  assign _11527_ = inv_23[8] ^ r_22[8] /*10775*/;
  assign sum_23[8] = _11527_ ^ _11526_ /*10774*/;
  assign _11528_ = _11527_ & _11526_ /*10773*/;
  assign _11529_ = inv_23[8] & r_22[8] /*10772*/;
  assign _11530_ = _11528_ | _11529_ /*10771*/;
  assign _11531_ = inv_23[9] ^ r_22[9] /*10769*/;
  assign sum_23[9] = _11531_ ^ _11530_ /*10768*/;
  assign _11532_ = _11531_ & _11530_ /*10767*/;
  assign _11533_ = inv_23[9] & r_22[9] /*10766*/;
  assign _11534_ = _11532_ | _11533_ /*10765*/;
  assign _11535_ = inv_23[10] ^ r_22[10] /*10763*/;
  assign sum_23[10] = _11535_ ^ _11534_ /*10762*/;
  assign _11536_ = _11535_ & _11534_ /*10761*/;
  assign _11537_ = inv_23[10] & r_22[10] /*10760*/;
  assign _11538_ = _11536_ | _11537_ /*10759*/;
  assign _11539_ = inv_23[11] ^ r_22[11] /*10757*/;
  assign sum_23[11] = _11539_ ^ _11538_ /*10756*/;
  assign _11540_ = _11539_ & _11538_ /*10755*/;
  assign _11541_ = inv_23[11] & r_22[11] /*10754*/;
  assign _11542_ = _11540_ | _11541_ /*10753*/;
  assign _11543_ = inv_23[12] ^ r_22[12] /*10751*/;
  assign sum_23[12] = _11543_ ^ _11542_ /*10750*/;
  assign _11544_ = _11543_ & _11542_ /*10749*/;
  assign _11545_ = inv_23[12] & r_22[12] /*10748*/;
  assign _11546_ = _11544_ | _11545_ /*10747*/;
  assign _11547_ = inv_23[13] ^ r_22[13] /*10745*/;
  assign sum_23[13] = _11547_ ^ _11546_ /*10744*/;
  assign _11548_ = _11547_ & _11546_ /*10743*/;
  assign _11549_ = inv_23[13] & r_22[13] /*10742*/;
  assign _11550_ = _11548_ | _11549_ /*10741*/;
  assign _11551_ = inv_23[14] ^ r_22[14] /*10739*/;
  assign sum_23[14] = _11551_ ^ _11550_ /*10738*/;
  assign _11552_ = _11551_ & _11550_ /*10737*/;
  assign _11553_ = inv_23[14] & r_22[14] /*10736*/;
  assign _11554_ = _11552_ | _11553_ /*10735*/;
  assign _11555_ = inv_23[15] ^ r_22[15] /*10733*/;
  assign sum_23[15] = _11555_ ^ _11554_ /*10732*/;
  assign _11556_ = _11555_ & _11554_ /*10731*/;
  assign _11557_ = inv_23[15] & r_22[15] /*10730*/;
  assign _11558_ = _11556_ | _11557_ /*10729*/;
  assign _11559_ = inv_23[16] ^ r_22[16] /*10727*/;
  assign sum_23[16] = _11559_ ^ _11558_ /*10726*/;
  assign _11560_ = _11559_ & _11558_ /*10725*/;
  assign _11561_ = inv_23[16] & r_22[16] /*10724*/;
  assign _11562_ = _11560_ | _11561_ /*10723*/;
  assign _11563_ = inv_23[17] ^ r_22[17] /*10721*/;
  assign sum_23[17] = _11563_ ^ _11562_ /*10720*/;
  assign _11564_ = _11563_ & _11562_ /*10719*/;
  assign _11565_ = inv_23[17] & r_22[17] /*10718*/;
  assign _11566_ = _11564_ | _11565_ /*10717*/;
  assign _11567_ = inv_23[18] ^ r_22[18] /*10715*/;
  assign sum_23[18] = _11567_ ^ _11566_ /*10714*/;
  assign _11568_ = _11567_ & _11566_ /*10713*/;
  assign _11569_ = inv_23[18] & r_22[18] /*10712*/;
  assign _11570_ = _11568_ | _11569_ /*10711*/;
  assign _11571_ = inv_23[19] ^ r_22[19] /*10709*/;
  assign sum_23[19] = _11571_ ^ _11570_ /*10708*/;
  assign _11572_ = _11571_ & _11570_ /*10707*/;
  assign _11573_ = inv_23[19] & r_22[19] /*10706*/;
  assign _11574_ = _11572_ | _11573_ /*10705*/;
  assign _11575_ = inv_23[20] ^ r_22[20] /*10703*/;
  assign sum_23[20] = _11575_ ^ _11574_ /*10702*/;
  assign _11576_ = _11575_ & _11574_ /*10701*/;
  assign _11577_ = inv_23[20] & r_22[20] /*10700*/;
  assign _11578_ = _11576_ | _11577_ /*10699*/;
  assign _11579_ = inv_23[21] ^ r_22[21] /*10697*/;
  assign sum_23[21] = _11579_ ^ _11578_ /*10696*/;
  assign _11580_ = _11579_ & _11578_ /*10695*/;
  assign _11581_ = inv_23[21] & r_22[21] /*10694*/;
  assign _11582_ = _11580_ | _11581_ /*10693*/;
  assign _11583_ = inv_23[22] ^ r_22[22] /*10691*/;
  assign sum_23[22] = _11583_ ^ _11582_ /*10690*/;
  assign _11584_ = _11583_ & _11582_ /*10689*/;
  assign _11585_ = inv_23[22] & r_22[22] /*10688*/;
  assign _11586_ = _11584_ | _11585_ /*10687*/;
  assign _11587_ = inv_23[23] ^ r_22[23] /*10685*/;
  assign sum_23[23] = _11587_ ^ _11586_ /*10684*/;
  assign _11588_ = _11587_ & _11586_ /*10683*/;
  assign _11589_ = inv_23[23] & r_22[23] /*10682*/;
  assign _11590_ = _11588_ | _11589_ /*10681*/;
  assign _11591_ = inv_23[24] ^ r_22[24] /*10679*/;
  assign sum_23[24] = _11591_ ^ _11590_ /*10678*/;
  assign _11592_ = _11591_ & _11590_ /*10677*/;
  assign _11593_ = inv_23[24] & r_22[24] /*10676*/;
  assign _11594_ = _11592_ | _11593_ /*10675*/;
  assign _11595_ = inv_23[25] ^ r_22[25] /*10673*/;
  assign sum_23[25] = _11595_ ^ _11594_ /*10672*/;
  assign _11596_ = _11595_ & _11594_ /*10671*/;
  assign _11597_ = inv_23[25] & r_22[25] /*10670*/;
  assign _11598_ = _11596_ | _11597_ /*10669*/;
  assign _11599_ = inv_23[26] ^ r_22[26] /*10667*/;
  assign sum_23[26] = _11599_ ^ _11598_ /*10666*/;
  assign _11600_ = _11599_ & _11598_ /*10665*/;
  assign _11601_ = inv_23[26] & r_22[26] /*10664*/;
  assign _11602_ = _11600_ | _11601_ /*10663*/;
  assign _11603_ = inv_23[27] ^ r_22[27] /*10661*/;
  assign sum_23[27] = _11603_ ^ _11602_ /*10660*/;
  assign _11604_ = _11603_ & _11602_ /*10659*/;
  assign _11605_ = inv_23[27] & r_22[27] /*10658*/;
  assign _11606_ = _11604_ | _11605_ /*10657*/;
  assign _11607_ = inv_23[28] ^ r_22[28] /*10655*/;
  assign sum_23[28] = _11607_ ^ _11606_ /*10654*/;
  assign _11608_ = _11607_ & _11606_ /*10653*/;
  assign _11609_ = inv_23[28] & r_22[28] /*10652*/;
  assign _11610_ = _11608_ | _11609_ /*10651*/;
  assign _11611_ = inv_23[29] ^ r_22[29] /*10649*/;
  assign sum_23[29] = _11611_ ^ _11610_ /*10648*/;
  assign _11612_ = _11611_ & _11610_ /*10647*/;
  assign _11613_ = inv_23[29] & r_22[29] /*10646*/;
  assign _11614_ = _11612_ | _11613_ /*10645*/;
  assign _11615_ = inv_23[30] ^ r_22[30] /*10643*/;
  assign sum_23[30] = _11615_ ^ _11614_ /*10642*/;
  assign _11616_ = _11615_ & _11614_ /*10641*/;
  assign _11617_ = inv_23[30] & r_22[30] /*10640*/;
  assign _11618_ = _11616_ | _11617_ /*10639*/;
  assign _11619_ = inv_23[31] ^ r_22[31] /*10637*/;
  assign sum_23[31] = _11619_ ^ _11618_ /*10636*/;
  assign _11620_ = _11619_ & _11618_ /*10635*/;
  assign _11621_ = inv_23[31] & r_22[31] /*10634*/;
  assign _11622_ = _11620_ | _11621_ /*10633*/;
  assign _11623_ = inv_23[32] ^ r_22[32] /*10631*/;
  assign sum_23[32] = _11623_ ^ _11622_ /*10630*/;
  assign _11624_ = _11623_ & _11622_ /*10629*/;
  assign _11625_ = inv_23[32] & r_22[32] /*10628*/;
  assign _11626_ = _11624_ | _11625_ /*10627*/;
  assign _11627_ = inv_23[33] ^ r_22[33] /*10625*/;
  assign sum_23[33] = _11627_ ^ _11626_ /*10624*/;
  assign _11628_ = _11627_ & _11626_ /*10623*/;
  assign _11629_ = inv_23[33] & r_22[33] /*10622*/;
  assign _11630_ = _11628_ | _11629_ /*10621*/;
  assign _11631_ = inv_23[34] ^ r_22[34] /*10619*/;
  assign sum_23[34] = _11631_ ^ _11630_ /*10618*/;
  assign _11632_ = _11631_ & _11630_ /*10617*/;
  assign _11633_ = inv_23[34] & r_22[34] /*10616*/;
  assign _11634_ = _11632_ | _11633_ /*10615*/;
  assign _11635_ = inv_23[35] ^ r_22[35] /*10613*/;
  assign sum_23[35] = _11635_ ^ _11634_ /*10612*/;
  assign _11636_ = _11635_ & _11634_ /*10611*/;
  assign _11637_ = inv_23[35] & r_22[35] /*10610*/;
  assign _11638_ = _11636_ | _11637_ /*10609*/;
  assign _11639_ = inv_23[36] ^ r_22[36] /*10607*/;
  assign sum_23[36] = _11639_ ^ _11638_ /*10606*/;
  assign _11640_ = _11639_ & _11638_ /*10605*/;
  assign _11641_ = inv_23[36] & r_22[36] /*10604*/;
  assign _11642_ = _11640_ | _11641_ /*10603*/;
  assign _11643_ = inv_23[37] ^ r_22[37] /*10601*/;
  assign sum_23[37] = _11643_ ^ _11642_ /*10600*/;
  assign _11644_ = _11643_ & _11642_ /*10599*/;
  assign _11645_ = inv_23[37] & r_22[37] /*10598*/;
  assign _11646_ = _11644_ | _11645_ /*10597*/;
  assign _11647_ = inv_23[38] ^ r_22[38] /*10595*/;
  assign sum_23[38] = _11647_ ^ _11646_ /*10594*/;
  assign _11648_ = _11647_ & _11646_ /*10593*/;
  assign _11649_ = inv_23[38] & r_22[38] /*10592*/;
  assign _11650_ = _11648_ | _11649_ /*10591*/;
  assign _11651_ = inv_23[39] ^ r_22[39] /*10589*/;
  assign sum_23[39] = _11651_ ^ _11650_ /*10588*/;
  assign _11652_ = _11651_ & _11650_ /*10587*/;
  assign _11653_ = inv_23[39] & r_22[39] /*10586*/;
  assign _11654_ = _11652_ | _11653_ /*10585*/;
  assign _11655_ = inv_23[40] ^ r_22[40] /*10583*/;
  assign sum_23[40] = _11655_ ^ _11654_ /*10582*/;
  assign _11656_ = _11655_ & _11654_ /*10581*/;
  assign _11657_ = inv_23[40] & r_22[40] /*10580*/;
  assign _11658_ = _11656_ | _11657_ /*10579*/;
  assign _11659_ = inv_23[41] ^ r_22[41] /*10577*/;
  assign sum_23[41] = _11659_ ^ _11658_ /*10576*/;
  assign _11660_ = _11659_ & _11658_ /*10575*/;
  assign _11661_ = inv_23[41] & r_22[41] /*10574*/;
  assign _11662_ = _11660_ | _11661_ /*10573*/;
  assign _11663_ = inv_23[42] ^ r_22[42] /*10571*/;
  assign sum_23[42] = _11663_ ^ _11662_ /*10570*/;
  assign _11664_ = _11663_ & _11662_ /*10569*/;
  assign _11665_ = inv_23[42] & r_22[42] /*10568*/;
  assign _11666_ = _11664_ | _11665_ /*10567*/;
  assign _11667_ = inv_23[43] ^ r_22[43] /*10565*/;
  assign sum_23[43] = _11667_ ^ _11666_ /*10564*/;
  assign _11668_ = _11667_ & _11666_ /*10563*/;
  assign _11669_ = inv_23[43] & r_22[43] /*10562*/;
  assign _11670_ = _11668_ | _11669_ /*10561*/;
  assign _11671_ = inv_23[44] ^ r_22[44] /*10559*/;
  assign sum_23[44] = _11671_ ^ _11670_ /*10558*/;
  assign _11672_ = _11671_ & _11670_ /*10557*/;
  assign _11673_ = inv_23[44] & r_22[44] /*10556*/;
  assign _11674_ = _11672_ | _11673_ /*10555*/;
  assign _11675_ = inv_23[45] ^ r_22[45] /*10553*/;
  assign sum_23[45] = _11675_ ^ _11674_ /*10552*/;
  assign _11676_ = _11675_ & _11674_ /*10551*/;
  assign _11677_ = inv_23[45] & r_22[45] /*10550*/;
  assign _11678_ = _11676_ | _11677_ /*10549*/;
  assign _11679_ = inv_23[46] ^ r_22[46] /*10547*/;
  assign sum_23[46] = _11679_ ^ _11678_ /*10546*/;
  assign _11680_ = _11679_ & _11678_ /*10545*/;
  assign _11681_ = inv_23[46] & r_22[46] /*10544*/;
  assign _11682_ = _11680_ | _11681_ /*10543*/;
  assign _11683_ = inv_23[47] ^ r_22[47] /*10541*/;
  assign sum_23[47] = _11683_ ^ _11682_ /*10540*/;
  assign _11684_ = _11683_ & _11682_ /*10539*/;
  assign _11685_ = inv_23[47] & r_22[47] /*10538*/;
  assign _11686_ = _11684_ | _11685_ /*10537*/;
  assign _11687_ = inv_23[48] ^ r_22[48] /*10535*/;
  assign sum_23[48] = _11687_ ^ _11686_ /*10534*/;
  assign _11688_ = _11687_ & _11686_ /*10533*/;
  assign _11689_ = inv_23[48] & r_22[48] /*10532*/;
  assign _11690_ = _11688_ | _11689_ /*10531*/;
  assign _11691_ = inv_23[49] ^ r_22[49] /*10529*/;
  assign sum_23[49] = _11691_ ^ _11690_ /*10528*/;
  assign _11692_ = _11691_ & _11690_ /*10527*/;
  assign _11693_ = inv_23[49] & r_22[49] /*10526*/;
  assign _11694_ = _11692_ | _11693_ /*10525*/;
  assign _11695_ = inv_23[50] ^ r_22[50] /*10523*/;
  assign sum_23[50] = _11695_ ^ _11694_ /*10522*/;
  assign _11696_ = _11695_ & _11694_ /*10521*/;
  assign _11697_ = inv_23[50] & r_22[50] /*10520*/;
  assign _11698_ = _11696_ | _11697_ /*10519*/;
  assign _11699_ = inv_23[51] ^ r_22[51] /*10517*/;
  assign sum_23[51] = _11699_ ^ _11698_ /*10516*/;
  assign _11700_ = _11699_ & _11698_ /*10515*/;
  assign _11701_ = inv_23[51] & r_22[51] /*10514*/;
  assign _11702_ = _11700_ | _11701_ /*10513*/;
  assign _11703_ = inv_23[52] ^ r_22[52] /*10511*/;
  assign sum_23[52] = _11703_ ^ _11702_ /*10510*/;
  assign _11704_ = _11703_ & _11702_ /*10509*/;
  assign _11705_ = inv_23[52] & r_22[52] /*10508*/;
  assign _11706_ = _11704_ | _11705_ /*10507*/;
  assign _11707_ = inv_23[53] ^ r_22[53] /*10505*/;
  assign sum_23[53] = _11707_ ^ _11706_ /*10504*/;
  assign _11708_ = _11707_ & _11706_ /*10503*/;
  assign _11709_ = inv_23[53] & r_22[53] /*10502*/;
  assign _11710_ = _11708_ | _11709_ /*10501*/;
  assign _11711_ = inv_23[54] ^ r_22[54] /*10499*/;
  assign sum_23[54] = _11711_ ^ _11710_ /*10498*/;
  assign _11712_ = _11711_ & _11710_ /*10497*/;
  assign _11713_ = inv_23[54] & r_22[54] /*10496*/;
  assign _11714_ = _11712_ | _11713_ /*10495*/;
  assign _11715_ = inv_23[55] ^ r_22[55] /*10493*/;
  assign sum_23[55] = _11715_ ^ _11714_ /*10492*/;
  assign _11716_ = _11715_ & _11714_ /*10491*/;
  assign _11717_ = inv_23[55] & r_22[55] /*10490*/;
  assign _11718_ = _11716_ | _11717_ /*10489*/;
  assign _11719_ = inv_23[56] ^ r_22[56] /*10487*/;
  assign sum_23[56] = _11719_ ^ _11718_ /*10486*/;
  assign _11720_ = _11719_ & _11718_ /*10485*/;
  assign _11721_ = inv_23[56] & r_22[56] /*10484*/;
  assign _11722_ = _11720_ | _11721_ /*10483*/;
  assign _11723_ = inv_23[57] ^ r_22[57] /*10481*/;
  assign sum_23[57] = _11723_ ^ _11722_ /*10480*/;
  assign _11724_ = _11723_ & _11722_ /*10479*/;
  assign _11725_ = inv_23[57] & r_22[57] /*10478*/;
  assign _11726_ = _11724_ | _11725_ /*10477*/;
  assign _11727_ = inv_23[58] ^ r_22[58] /*10475*/;
  assign sum_23[58] = _11727_ ^ _11726_ /*10474*/;
  assign _11728_ = _11727_ & _11726_ /*10473*/;
  assign _11729_ = inv_23[58] & r_22[58] /*10472*/;
  assign _11730_ = _11728_ | _11729_ /*10471*/;
  assign _11731_ = inv_23[59] ^ r_22[59] /*10469*/;
  assign sum_23[59] = _11731_ ^ _11730_ /*10468*/;
  assign _11732_ = _11731_ & _11730_ /*10467*/;
  assign _11733_ = inv_23[59] & r_22[59] /*10466*/;
  assign _11734_ = _11732_ | _11733_ /*10465*/;
  assign _11735_ = inv_23[60] ^ r_22[60] /*10463*/;
  assign sum_23[60] = _11735_ ^ _11734_ /*10462*/;
  assign _11736_ = _11735_ & _11734_ /*10461*/;
  assign _11737_ = inv_23[60] & r_22[60] /*10460*/;
  assign _11738_ = _11736_ | _11737_ /*10459*/;
  assign _11739_ = inv_23[61] ^ r_22[61] /*10457*/;
  assign sum_23[61] = _11739_ ^ _11738_ /*10456*/;
  assign _11740_ = _11739_ & _11738_ /*10455*/;
  assign _11741_ = inv_23[61] & r_22[61] /*10454*/;
  assign _11742_ = _11740_ | _11741_ /*10453*/;
  assign _11743_ = inv_23[62] ^ r_22[62] /*10451*/;
  assign sum_23[62] = _11743_ ^ _11742_ /*10450*/;
  assign _11744_ = _11743_ & _11742_ /*10449*/;
  assign _11745_ = inv_23[62] & r_22[62] /*10448*/;
  assign _11746_ = _11744_ | _11745_ /*10447*/;
  assign _11747_ = inv_23[63] ^ r_22[63] /*10445*/;
  assign sum_23[63] = _11747_ ^ _11746_ /*10444*/;
  assign _11748_ = _11747_ & _11746_ /*10443*/;
  assign _11749_ = inv_23[63] & r_22[63] /*10442*/;
  assign _11750_ = _11748_ | _11749_ /*10441*/;
  assign _11751_ = inv_23[64] ^ r_22[64] /*10439*/;
  assign sum_23[64] = _11751_ ^ _11750_ /*10438*/;
  assign _11752_ = _11751_ & _11750_ /*10437*/;
  assign _11753_ = inv_23[64] & r_22[64] /*10436*/;
  assign _11754_ = _11752_ | _11753_ /*10435*/;
  assign _11755_ = inv_23[65] ^ r_22[65] /*10433*/;
  assign sum_23[65] = _11755_ ^ _11754_ /*10432*/;
  assign _11756_ = _11755_ & _11754_ /*10431*/;
  assign _11757_ = inv_23[65] & r_22[65] /*10430*/;
  assign _11758_ = _11756_ | _11757_ /*10429*/;
  assign _11759_ = inv_23[66] ^ r_22[66] /*10427*/;
  assign sum_23[66] = _11759_ ^ _11758_ /*10426*/;
  assign _11760_ = _11759_ & _11758_ /*10425*/;
  assign _11761_ = inv_23[66] & r_22[66] /*10424*/;
  assign _11762_ = _11760_ | _11761_ /*10423*/;
  assign _11763_ = inv_23[67] ^ r_22[67] /*10421*/;
  assign sum_23[67] = _11763_ ^ _11762_ /*10420*/;
  assign _11764_ = _11763_ & _11762_ /*10419*/;
  assign _11765_ = inv_23[67] & r_22[67] /*10418*/;
  assign _11766_ = _11764_ | _11765_ /*10417*/;
  assign _11767_ = inv_23[68] ^ r_22[68] /*10415*/;
  assign sum_23[68] = _11767_ ^ _11766_ /*10414*/;
  assign _11768_ = _11767_ & _11766_ /*10413*/;
  assign _11769_ = inv_23[68] & r_22[68] /*10412*/;
  assign _11770_ = _11768_ | _11769_ /*10411*/;
  assign _11771_ = inv_23[69] ^ r_22[69] /*10409*/;
  assign sum_23[69] = _11771_ ^ _11770_ /*10408*/;
  assign _11772_ = _11771_ & _11770_ /*10407*/;
  assign _11773_ = inv_23[69] & r_22[69] /*10406*/;
  assign _11774_ = _11772_ | _11773_ /*10405*/;
  assign _11775_ = inv_23[70] ^ r_22[70] /*10403*/;
  assign sum_23[70] = _11775_ ^ _11774_ /*10402*/;
  assign _11776_ = _11775_ & _11774_ /*10401*/;
  assign _11777_ = inv_23[70] & r_22[70] /*10400*/;
  assign _11778_ = _11776_ | _11777_ /*10399*/;
  assign _11779_ = inv_23[71] ^ r_22[71] /*10397*/;
  assign sum_23[71] = _11779_ ^ _11778_ /*10396*/;
  assign _11780_ = _11779_ & _11778_ /*10395*/;
  assign _11781_ = inv_23[71] & r_22[71] /*10394*/;
  assign _11782_ = _11780_ | _11781_ /*10393*/;
  assign _11783_ = inv_23[72] ^ r_22[72] /*10391*/;
  assign sum_23[72] = _11783_ ^ _11782_ /*10390*/;
  assign _11784_ = _11783_ & _11782_ /*10389*/;
  assign _11785_ = inv_23[72] & r_22[72] /*10388*/;
  assign _11786_ = _11784_ | _11785_ /*10387*/;
  assign _11787_ = inv_23[73] ^ r_22[73] /*10385*/;
  assign sum_23[73] = _11787_ ^ _11786_ /*10384*/;
  assign _11788_ = _11787_ & _11786_ /*10383*/;
  assign _11789_ = inv_23[73] & r_22[73] /*10382*/;
  assign _11790_ = _11788_ | _11789_ /*10381*/;
  assign _11791_ = inv_23[74] ^ r_22[74] /*10379*/;
  assign sum_23[74] = _11791_ ^ _11790_ /*10378*/;
  assign _11792_ = _11791_ & _11790_ /*10377*/;
  assign _11793_ = inv_23[74] & r_22[74] /*10376*/;
  assign _11794_ = _11792_ | _11793_ /*10375*/;
  assign _11795_ = inv_23[75] ^ r_22[75] /*10373*/;
  assign sum_23[75] = _11795_ ^ _11794_ /*10372*/;
  assign _11796_ = _11795_ & _11794_ /*10371*/;
  assign _11797_ = inv_23[75] & r_22[75] /*10370*/;
  assign _11798_ = _11796_ | _11797_ /*10369*/;
  assign _11799_ = inv_23[76] ^ r_22[76] /*10367*/;
  assign sum_23[76] = _11799_ ^ _11798_ /*10366*/;
  assign _11800_ = _11799_ & _11798_ /*10365*/;
  assign _11801_ = inv_23[76] & r_22[76] /*10364*/;
  assign _11802_ = _11800_ | _11801_ /*10363*/;
  assign _11803_ = inv_23[77] ^ r_22[77] /*10361*/;
  assign sum_23[77] = _11803_ ^ _11802_ /*10360*/;
  assign _11804_ = _11803_ & _11802_ /*10359*/;
  assign _11805_ = inv_23[77] & r_22[77] /*10358*/;
  assign _11806_ = _11804_ | _11805_ /*10357*/;
  assign _11807_ = inv_23[78] ^ r_22[78] /*10355*/;
  assign sum_23[78] = _11807_ ^ _11806_ /*10354*/;
  assign _11808_ = _11807_ & _11806_ /*10353*/;
  assign _11809_ = inv_23[78] & r_22[78] /*10352*/;
  assign _11810_ = _11808_ | _11809_ /*10351*/;
  assign _11811_ = inv_23[79] ^ r_22[79] /*10349*/;
  assign sum_23[79] = _11811_ ^ _11810_ /*10348*/;
  assign _11812_ = _11811_ & _11810_ /*10347*/;
  assign _11813_ = inv_23[79] & r_22[79] /*10346*/;
  assign _11814_ = _11812_ | _11813_ /*10345*/;
  assign _11815_ = inv_23[80] ^ r_22[80] /*10343*/;
  assign sum_23[80] = _11815_ ^ _11814_ /*10342*/;
  assign _11816_ = _11815_ & _11814_ /*10341*/;
  assign _11817_ = inv_23[80] & r_22[80] /*10340*/;
  assign _11818_ = _11816_ | _11817_ /*10339*/;
  assign _11819_ = inv_23[81] ^ r_22[81] /*10337*/;
  assign sum_23[81] = _11819_ ^ _11818_ /*10336*/;
  assign _11820_ = _11819_ & _11818_ /*10335*/;
  assign _11821_ = inv_23[81] & r_22[81] /*10334*/;
  assign _11822_ = _11820_ | _11821_ /*10333*/;
  assign _11823_ = inv_23[82] ^ r_22[82] /*10331*/;
  assign sum_23[82] = _11823_ ^ _11822_ /*10330*/;
  assign _11824_ = _11823_ & _11822_ /*10329*/;
  assign _11825_ = inv_23[82] & r_22[82] /*10328*/;
  assign _11826_ = _11824_ | _11825_ /*10327*/;
  assign _11827_ = inv_23[83] ^ r_22[83] /*10325*/;
  assign sum_23[83] = _11827_ ^ _11826_ /*10324*/;
  assign _11828_ = _11827_ & _11826_ /*10323*/;
  assign _11829_ = inv_23[83] & r_22[83] /*10322*/;
  assign _11830_ = _11828_ | _11829_ /*10321*/;
  assign _11831_ = inv_23[84] ^ r_22[84] /*10319*/;
  assign sum_23[84] = _11831_ ^ _11830_ /*10318*/;
  assign _11832_ = _11831_ & _11830_ /*10317*/;
  assign _11833_ = inv_23[84] & r_22[84] /*10316*/;
  assign _11834_ = _11832_ | _11833_ /*10315*/;
  assign _11835_ = _11834_ ^ _11830_ /*10314*/;
  assign _11836_ = ~_11835_ /*10313*/;
  assign _11837_ = sum_23[84] & _11836_ /*10312*/;
  assign _11838_ = _11835_ & _11834_ /*10311*/;
  assign sum_23[85] = _11838_ | _11837_ /*10310*/;
  assign q[9] = ~sum_23[85] /*10309*/;
  assign m_23[0] = r_22[0] /*10308*/;
  assign m_23[1] = r_22[1] /*10307*/;
  assign m_23[2] = r_22[2] /*10306*/;
  assign m_23[3] = r_22[3] /*10305*/;
  assign m_23[4] = r_22[4] /*10304*/;
  assign m_23[5] = r_22[5] /*10303*/;
  assign m_23[6] = r_22[6] /*10302*/;
  assign m_23[7] = r_22[7] /*10301*/;
  assign m_23[8] = r_22[8] /*10300*/;
  assign m_23[9] = r_22[9] /*10299*/;
  assign m_23[10] = r_22[10] /*10298*/;
  assign m_23[11] = r_22[11] /*10297*/;
  assign m_23[12] = r_22[12] /*10296*/;
  assign m_23[13] = r_22[13] /*10295*/;
  assign m_23[14] = r_22[14] /*10294*/;
  assign m_23[15] = r_22[15] /*10293*/;
  assign m_23[16] = r_22[16] /*10292*/;
  assign m_23[17] = r_22[17] /*10291*/;
  assign m_23[18] = r_22[18] /*10290*/;
  assign m_23[19] = r_22[19] /*10289*/;
  assign m_23[20] = r_22[20] /*10288*/;
  assign m_23[21] = r_22[21] /*10287*/;
  assign m_23[22] = r_22[22] /*10286*/;
  assign m_23[23] = r_22[23] /*10285*/;
  assign m_23[24] = r_22[24] /*10284*/;
  assign m_23[25] = r_22[25] /*10283*/;
  assign m_23[26] = r_22[26] /*10282*/;
  assign m_23[27] = r_22[27] /*10281*/;
  assign m_23[28] = r_22[28] /*10280*/;
  assign m_23[29] = r_22[29] /*10279*/;
  assign m_23[30] = r_22[30] /*10278*/;
  assign m_23[31] = r_22[31] /*10277*/;
  assign m_23[32] = r_22[32] /*10276*/;
  assign m_23[33] = r_22[33] /*10275*/;
  assign m_23[34] = r_22[34] /*10274*/;
  assign m_23[35] = r_22[35] /*10273*/;
  assign m_23[36] = r_22[36] /*10272*/;
  assign m_23[37] = r_22[37] /*10271*/;
  assign m_23[38] = r_22[38] /*10270*/;
  assign m_23[39] = r_22[39] /*10269*/;
  assign m_23[40] = r_22[40] /*10268*/;
  assign m_23[41] = r_22[41] /*10267*/;
  assign m_23[42] = r_22[42] /*10266*/;
  assign m_23[43] = r_22[43] /*10265*/;
  assign m_23[44] = r_22[44] /*10264*/;
  assign m_23[45] = r_22[45] /*10263*/;
  assign m_23[46] = r_22[46] /*10262*/;
  assign m_23[47] = r_22[47] /*10261*/;
  assign m_23[48] = r_22[48] /*10260*/;
  assign m_23[49] = r_22[49] /*10259*/;
  assign m_23[50] = r_22[50] /*10258*/;
  assign m_23[51] = r_22[51] /*10257*/;
  assign m_23[52] = r_22[52] /*10256*/;
  assign m_23[53] = r_22[53] /*10255*/;
  assign m_23[54] = r_22[54] /*10254*/;
  assign m_23[55] = r_22[55] /*10253*/;
  assign m_23[56] = r_22[56] /*10252*/;
  assign m_23[57] = r_22[57] /*10251*/;
  assign m_23[58] = r_22[58] /*10250*/;
  assign m_23[59] = r_22[59] /*10249*/;
  assign m_23[60] = r_22[60] /*10248*/;
  assign m_23[61] = r_22[61] /*10247*/;
  assign m_23[62] = r_22[62] /*10246*/;
  assign m_23[63] = r_22[63] /*10245*/;
  assign m_23[64] = r_22[64] /*10244*/;
  assign m_23[65] = r_22[65] /*10243*/;
  assign m_23[66] = r_22[66] /*10242*/;
  assign m_23[67] = r_22[67] /*10241*/;
  assign m_23[68] = r_22[68] /*10240*/;
  assign m_23[69] = r_22[69] /*10239*/;
  assign m_23[70] = r_22[70] /*10238*/;
  assign m_23[71] = r_22[71] /*10237*/;
  assign m_23[72] = r_22[72] /*10236*/;
  assign m_23[73] = r_22[73] /*10235*/;
  assign m_23[74] = r_22[74] /*10234*/;
  assign m_23[75] = r_22[75] /*10233*/;
  assign m_23[76] = r_22[76] /*10232*/;
  assign m_23[77] = r_22[77] /*10231*/;
  assign m_23[78] = r_22[78] /*10230*/;
  assign m_23[79] = r_22[79] /*10229*/;
  assign m_23[80] = r_22[80] /*10228*/;
  assign m_23[81] = r_22[81] /*10227*/;
  assign m_23[82] = r_22[82] /*10226*/;
  assign m_23[83] = r_22[83] /*10225*/;
  assign m_23[84] = r_22[84] /*10224*/;
  assign m_23[85] = r_22[84] /*10223*/;
  assign _11840_ = ~q[9] /*10222*/;
  assign _11841_ = sum_23[0] & q[9] /*10221*/;
  assign _11842_ = m_23[0] & _11840_ /*10220*/;
  assign r_23[0] = _11842_ | _11841_ /*10219*/;
  assign _11843_ = ~q[9] /*10218*/;
  assign _11844_ = sum_23[1] & q[9] /*10217*/;
  assign _11845_ = m_23[1] & _11843_ /*10216*/;
  assign r_23[1] = _11845_ | _11844_ /*10215*/;
  assign _11846_ = ~q[9] /*10214*/;
  assign _11847_ = sum_23[2] & q[9] /*10213*/;
  assign _11848_ = m_23[2] & _11846_ /*10212*/;
  assign r_23[2] = _11848_ | _11847_ /*10211*/;
  assign _11849_ = ~q[9] /*10210*/;
  assign _11850_ = sum_23[3] & q[9] /*10209*/;
  assign _11851_ = m_23[3] & _11849_ /*10208*/;
  assign r_23[3] = _11851_ | _11850_ /*10207*/;
  assign _11852_ = ~q[9] /*10206*/;
  assign _11853_ = sum_23[4] & q[9] /*10205*/;
  assign _11854_ = m_23[4] & _11852_ /*10204*/;
  assign r_23[4] = _11854_ | _11853_ /*10203*/;
  assign _11855_ = ~q[9] /*10202*/;
  assign _11856_ = sum_23[5] & q[9] /*10201*/;
  assign _11857_ = m_23[5] & _11855_ /*10200*/;
  assign r_23[5] = _11857_ | _11856_ /*10199*/;
  assign _11858_ = ~q[9] /*10198*/;
  assign _11859_ = sum_23[6] & q[9] /*10197*/;
  assign _11860_ = m_23[6] & _11858_ /*10196*/;
  assign r_23[6] = _11860_ | _11859_ /*10195*/;
  assign _11861_ = ~q[9] /*10194*/;
  assign _11862_ = sum_23[7] & q[9] /*10193*/;
  assign _11863_ = m_23[7] & _11861_ /*10192*/;
  assign r_23[7] = _11863_ | _11862_ /*10191*/;
  assign _11864_ = ~q[9] /*10190*/;
  assign _11865_ = sum_23[8] & q[9] /*10189*/;
  assign _11866_ = m_23[8] & _11864_ /*10188*/;
  assign r_23[8] = _11866_ | _11865_ /*10187*/;
  assign _11867_ = ~q[9] /*10186*/;
  assign _11868_ = sum_23[9] & q[9] /*10185*/;
  assign _11869_ = m_23[9] & _11867_ /*10184*/;
  assign r_23[9] = _11869_ | _11868_ /*10183*/;
  assign _11870_ = ~q[9] /*10182*/;
  assign _11871_ = sum_23[10] & q[9] /*10181*/;
  assign _11872_ = m_23[10] & _11870_ /*10180*/;
  assign r_23[10] = _11872_ | _11871_ /*10179*/;
  assign _11873_ = ~q[9] /*10178*/;
  assign _11874_ = sum_23[11] & q[9] /*10177*/;
  assign _11875_ = m_23[11] & _11873_ /*10176*/;
  assign r_23[11] = _11875_ | _11874_ /*10175*/;
  assign _11876_ = ~q[9] /*10174*/;
  assign _11877_ = sum_23[12] & q[9] /*10173*/;
  assign _11878_ = m_23[12] & _11876_ /*10172*/;
  assign r_23[12] = _11878_ | _11877_ /*10171*/;
  assign _11879_ = ~q[9] /*10170*/;
  assign _11880_ = sum_23[13] & q[9] /*10169*/;
  assign _11881_ = m_23[13] & _11879_ /*10168*/;
  assign r_23[13] = _11881_ | _11880_ /*10167*/;
  assign _11882_ = ~q[9] /*10166*/;
  assign _11883_ = sum_23[14] & q[9] /*10165*/;
  assign _11884_ = m_23[14] & _11882_ /*10164*/;
  assign r_23[14] = _11884_ | _11883_ /*10163*/;
  assign _11885_ = ~q[9] /*10162*/;
  assign _11886_ = sum_23[15] & q[9] /*10161*/;
  assign _11887_ = m_23[15] & _11885_ /*10160*/;
  assign r_23[15] = _11887_ | _11886_ /*10159*/;
  assign _11888_ = ~q[9] /*10158*/;
  assign _11889_ = sum_23[16] & q[9] /*10157*/;
  assign _11890_ = m_23[16] & _11888_ /*10156*/;
  assign r_23[16] = _11890_ | _11889_ /*10155*/;
  assign _11891_ = ~q[9] /*10154*/;
  assign _11892_ = sum_23[17] & q[9] /*10153*/;
  assign _11893_ = m_23[17] & _11891_ /*10152*/;
  assign r_23[17] = _11893_ | _11892_ /*10151*/;
  assign _11894_ = ~q[9] /*10150*/;
  assign _11895_ = sum_23[18] & q[9] /*10149*/;
  assign _11896_ = m_23[18] & _11894_ /*10148*/;
  assign r_23[18] = _11896_ | _11895_ /*10147*/;
  assign _11897_ = ~q[9] /*10146*/;
  assign _11898_ = sum_23[19] & q[9] /*10145*/;
  assign _11899_ = m_23[19] & _11897_ /*10144*/;
  assign r_23[19] = _11899_ | _11898_ /*10143*/;
  assign _11900_ = ~q[9] /*10142*/;
  assign _11901_ = sum_23[20] & q[9] /*10141*/;
  assign _11902_ = m_23[20] & _11900_ /*10140*/;
  assign r_23[20] = _11902_ | _11901_ /*10139*/;
  assign _11903_ = ~q[9] /*10138*/;
  assign _11904_ = sum_23[21] & q[9] /*10137*/;
  assign _11905_ = m_23[21] & _11903_ /*10136*/;
  assign r_23[21] = _11905_ | _11904_ /*10135*/;
  assign _11906_ = ~q[9] /*10134*/;
  assign _11907_ = sum_23[22] & q[9] /*10133*/;
  assign _11908_ = m_23[22] & _11906_ /*10132*/;
  assign r_23[22] = _11908_ | _11907_ /*10131*/;
  assign _11909_ = ~q[9] /*10130*/;
  assign _11910_ = sum_23[23] & q[9] /*10129*/;
  assign _11911_ = m_23[23] & _11909_ /*10128*/;
  assign r_23[23] = _11911_ | _11910_ /*10127*/;
  assign _11912_ = ~q[9] /*10126*/;
  assign _11913_ = sum_23[24] & q[9] /*10125*/;
  assign _11914_ = m_23[24] & _11912_ /*10124*/;
  assign r_23[24] = _11914_ | _11913_ /*10123*/;
  assign _11915_ = ~q[9] /*10122*/;
  assign _11916_ = sum_23[25] & q[9] /*10121*/;
  assign _11917_ = m_23[25] & _11915_ /*10120*/;
  assign r_23[25] = _11917_ | _11916_ /*10119*/;
  assign _11918_ = ~q[9] /*10118*/;
  assign _11919_ = sum_23[26] & q[9] /*10117*/;
  assign _11920_ = m_23[26] & _11918_ /*10116*/;
  assign r_23[26] = _11920_ | _11919_ /*10115*/;
  assign _11921_ = ~q[9] /*10114*/;
  assign _11922_ = sum_23[27] & q[9] /*10113*/;
  assign _11923_ = m_23[27] & _11921_ /*10112*/;
  assign r_23[27] = _11923_ | _11922_ /*10111*/;
  assign _11924_ = ~q[9] /*10110*/;
  assign _11925_ = sum_23[28] & q[9] /*10109*/;
  assign _11926_ = m_23[28] & _11924_ /*10108*/;
  assign r_23[28] = _11926_ | _11925_ /*10107*/;
  assign _11927_ = ~q[9] /*10106*/;
  assign _11928_ = sum_23[29] & q[9] /*10105*/;
  assign _11929_ = m_23[29] & _11927_ /*10104*/;
  assign r_23[29] = _11929_ | _11928_ /*10103*/;
  assign _11930_ = ~q[9] /*10102*/;
  assign _11931_ = sum_23[30] & q[9] /*10101*/;
  assign _11932_ = m_23[30] & _11930_ /*10100*/;
  assign r_23[30] = _11932_ | _11931_ /*10099*/;
  assign _11933_ = ~q[9] /*10098*/;
  assign _11934_ = sum_23[31] & q[9] /*10097*/;
  assign _11935_ = m_23[31] & _11933_ /*10096*/;
  assign r_23[31] = _11935_ | _11934_ /*10095*/;
  assign _11936_ = ~q[9] /*10094*/;
  assign _11937_ = sum_23[32] & q[9] /*10093*/;
  assign _11938_ = m_23[32] & _11936_ /*10092*/;
  assign r_23[32] = _11938_ | _11937_ /*10091*/;
  assign _11939_ = ~q[9] /*10090*/;
  assign _11940_ = sum_23[33] & q[9] /*10089*/;
  assign _11941_ = m_23[33] & _11939_ /*10088*/;
  assign r_23[33] = _11941_ | _11940_ /*10087*/;
  assign _11942_ = ~q[9] /*10086*/;
  assign _11943_ = sum_23[34] & q[9] /*10085*/;
  assign _11944_ = m_23[34] & _11942_ /*10084*/;
  assign r_23[34] = _11944_ | _11943_ /*10083*/;
  assign _11945_ = ~q[9] /*10082*/;
  assign _11946_ = sum_23[35] & q[9] /*10081*/;
  assign _11947_ = m_23[35] & _11945_ /*10080*/;
  assign r_23[35] = _11947_ | _11946_ /*10079*/;
  assign _11948_ = ~q[9] /*10078*/;
  assign _11949_ = sum_23[36] & q[9] /*10077*/;
  assign _11950_ = m_23[36] & _11948_ /*10076*/;
  assign r_23[36] = _11950_ | _11949_ /*10075*/;
  assign _11951_ = ~q[9] /*10074*/;
  assign _11952_ = sum_23[37] & q[9] /*10073*/;
  assign _11953_ = m_23[37] & _11951_ /*10072*/;
  assign r_23[37] = _11953_ | _11952_ /*10071*/;
  assign _11954_ = ~q[9] /*10070*/;
  assign _11955_ = sum_23[38] & q[9] /*10069*/;
  assign _11956_ = m_23[38] & _11954_ /*10068*/;
  assign r_23[38] = _11956_ | _11955_ /*10067*/;
  assign _11957_ = ~q[9] /*10066*/;
  assign _11958_ = sum_23[39] & q[9] /*10065*/;
  assign _11959_ = m_23[39] & _11957_ /*10064*/;
  assign r_23[39] = _11959_ | _11958_ /*10063*/;
  assign _11960_ = ~q[9] /*10062*/;
  assign _11961_ = sum_23[40] & q[9] /*10061*/;
  assign _11962_ = m_23[40] & _11960_ /*10060*/;
  assign r_23[40] = _11962_ | _11961_ /*10059*/;
  assign _11963_ = ~q[9] /*10058*/;
  assign _11964_ = sum_23[41] & q[9] /*10057*/;
  assign _11965_ = m_23[41] & _11963_ /*10056*/;
  assign r_23[41] = _11965_ | _11964_ /*10055*/;
  assign _11966_ = ~q[9] /*10054*/;
  assign _11967_ = sum_23[42] & q[9] /*10053*/;
  assign _11968_ = m_23[42] & _11966_ /*10052*/;
  assign r_23[42] = _11968_ | _11967_ /*10051*/;
  assign _11969_ = ~q[9] /*10050*/;
  assign _11970_ = sum_23[43] & q[9] /*10049*/;
  assign _11971_ = m_23[43] & _11969_ /*10048*/;
  assign r_23[43] = _11971_ | _11970_ /*10047*/;
  assign _11972_ = ~q[9] /*10046*/;
  assign _11973_ = sum_23[44] & q[9] /*10045*/;
  assign _11974_ = m_23[44] & _11972_ /*10044*/;
  assign r_23[44] = _11974_ | _11973_ /*10043*/;
  assign _11975_ = ~q[9] /*10042*/;
  assign _11976_ = sum_23[45] & q[9] /*10041*/;
  assign _11977_ = m_23[45] & _11975_ /*10040*/;
  assign r_23[45] = _11977_ | _11976_ /*10039*/;
  assign _11978_ = ~q[9] /*10038*/;
  assign _11979_ = sum_23[46] & q[9] /*10037*/;
  assign _11980_ = m_23[46] & _11978_ /*10036*/;
  assign r_23[46] = _11980_ | _11979_ /*10035*/;
  assign _11981_ = ~q[9] /*10034*/;
  assign _11982_ = sum_23[47] & q[9] /*10033*/;
  assign _11983_ = m_23[47] & _11981_ /*10032*/;
  assign r_23[47] = _11983_ | _11982_ /*10031*/;
  assign _11984_ = ~q[9] /*10030*/;
  assign _11985_ = sum_23[48] & q[9] /*10029*/;
  assign _11986_ = m_23[48] & _11984_ /*10028*/;
  assign r_23[48] = _11986_ | _11985_ /*10027*/;
  assign _11987_ = ~q[9] /*10026*/;
  assign _11988_ = sum_23[49] & q[9] /*10025*/;
  assign _11989_ = m_23[49] & _11987_ /*10024*/;
  assign r_23[49] = _11989_ | _11988_ /*10023*/;
  assign _11990_ = ~q[9] /*10022*/;
  assign _11991_ = sum_23[50] & q[9] /*10021*/;
  assign _11992_ = m_23[50] & _11990_ /*10020*/;
  assign r_23[50] = _11992_ | _11991_ /*10019*/;
  assign _11993_ = ~q[9] /*10018*/;
  assign _11994_ = sum_23[51] & q[9] /*10017*/;
  assign _11995_ = m_23[51] & _11993_ /*10016*/;
  assign r_23[51] = _11995_ | _11994_ /*10015*/;
  assign _11996_ = ~q[9] /*10014*/;
  assign _11997_ = sum_23[52] & q[9] /*10013*/;
  assign _11998_ = m_23[52] & _11996_ /*10012*/;
  assign r_23[52] = _11998_ | _11997_ /*10011*/;
  assign _11999_ = ~q[9] /*10010*/;
  assign _12000_ = sum_23[53] & q[9] /*10009*/;
  assign _12001_ = m_23[53] & _11999_ /*10008*/;
  assign r_23[53] = _12001_ | _12000_ /*10007*/;
  assign _12002_ = ~q[9] /*10006*/;
  assign _12003_ = sum_23[54] & q[9] /*10005*/;
  assign _12004_ = m_23[54] & _12002_ /*10004*/;
  assign r_23[54] = _12004_ | _12003_ /*10003*/;
  assign _12005_ = ~q[9] /*10002*/;
  assign _12006_ = sum_23[55] & q[9] /*10001*/;
  assign _12007_ = m_23[55] & _12005_ /*10000*/;
  assign r_23[55] = _12007_ | _12006_ /*9999*/;
  assign _12008_ = ~q[9] /*9998*/;
  assign _12009_ = sum_23[56] & q[9] /*9997*/;
  assign _12010_ = m_23[56] & _12008_ /*9996*/;
  assign r_23[56] = _12010_ | _12009_ /*9995*/;
  assign _12011_ = ~q[9] /*9994*/;
  assign _12012_ = sum_23[57] & q[9] /*9993*/;
  assign _12013_ = m_23[57] & _12011_ /*9992*/;
  assign r_23[57] = _12013_ | _12012_ /*9991*/;
  assign _12014_ = ~q[9] /*9990*/;
  assign _12015_ = sum_23[58] & q[9] /*9989*/;
  assign _12016_ = m_23[58] & _12014_ /*9988*/;
  assign r_23[58] = _12016_ | _12015_ /*9987*/;
  assign _12017_ = ~q[9] /*9986*/;
  assign _12018_ = sum_23[59] & q[9] /*9985*/;
  assign _12019_ = m_23[59] & _12017_ /*9984*/;
  assign r_23[59] = _12019_ | _12018_ /*9983*/;
  assign _12020_ = ~q[9] /*9982*/;
  assign _12021_ = sum_23[60] & q[9] /*9981*/;
  assign _12022_ = m_23[60] & _12020_ /*9980*/;
  assign r_23[60] = _12022_ | _12021_ /*9979*/;
  assign _12023_ = ~q[9] /*9978*/;
  assign _12024_ = sum_23[61] & q[9] /*9977*/;
  assign _12025_ = m_23[61] & _12023_ /*9976*/;
  assign r_23[61] = _12025_ | _12024_ /*9975*/;
  assign _12026_ = ~q[9] /*9974*/;
  assign _12027_ = sum_23[62] & q[9] /*9973*/;
  assign _12028_ = m_23[62] & _12026_ /*9972*/;
  assign r_23[62] = _12028_ | _12027_ /*9971*/;
  assign _12029_ = ~q[9] /*9970*/;
  assign _12030_ = sum_23[63] & q[9] /*9969*/;
  assign _12031_ = m_23[63] & _12029_ /*9968*/;
  assign r_23[63] = _12031_ | _12030_ /*9967*/;
  assign _12032_ = ~q[9] /*9966*/;
  assign _12033_ = sum_23[64] & q[9] /*9965*/;
  assign _12034_ = m_23[64] & _12032_ /*9964*/;
  assign r_23[64] = _12034_ | _12033_ /*9963*/;
  assign _12035_ = ~q[9] /*9962*/;
  assign _12036_ = sum_23[65] & q[9] /*9961*/;
  assign _12037_ = m_23[65] & _12035_ /*9960*/;
  assign r_23[65] = _12037_ | _12036_ /*9959*/;
  assign _12038_ = ~q[9] /*9958*/;
  assign _12039_ = sum_23[66] & q[9] /*9957*/;
  assign _12040_ = m_23[66] & _12038_ /*9956*/;
  assign r_23[66] = _12040_ | _12039_ /*9955*/;
  assign _12041_ = ~q[9] /*9954*/;
  assign _12042_ = sum_23[67] & q[9] /*9953*/;
  assign _12043_ = m_23[67] & _12041_ /*9952*/;
  assign r_23[67] = _12043_ | _12042_ /*9951*/;
  assign _12044_ = ~q[9] /*9950*/;
  assign _12045_ = sum_23[68] & q[9] /*9949*/;
  assign _12046_ = m_23[68] & _12044_ /*9948*/;
  assign r_23[68] = _12046_ | _12045_ /*9947*/;
  assign _12047_ = ~q[9] /*9946*/;
  assign _12048_ = sum_23[69] & q[9] /*9945*/;
  assign _12049_ = m_23[69] & _12047_ /*9944*/;
  assign r_23[69] = _12049_ | _12048_ /*9943*/;
  assign _12050_ = ~q[9] /*9942*/;
  assign _12051_ = sum_23[70] & q[9] /*9941*/;
  assign _12052_ = m_23[70] & _12050_ /*9940*/;
  assign r_23[70] = _12052_ | _12051_ /*9939*/;
  assign _12053_ = ~q[9] /*9938*/;
  assign _12054_ = sum_23[71] & q[9] /*9937*/;
  assign _12055_ = m_23[71] & _12053_ /*9936*/;
  assign r_23[71] = _12055_ | _12054_ /*9935*/;
  assign _12056_ = ~q[9] /*9934*/;
  assign _12057_ = sum_23[72] & q[9] /*9933*/;
  assign _12058_ = m_23[72] & _12056_ /*9932*/;
  assign r_23[72] = _12058_ | _12057_ /*9931*/;
  assign _12059_ = ~q[9] /*9930*/;
  assign _12060_ = sum_23[73] & q[9] /*9929*/;
  assign _12061_ = m_23[73] & _12059_ /*9928*/;
  assign r_23[73] = _12061_ | _12060_ /*9927*/;
  assign _12062_ = ~q[9] /*9926*/;
  assign _12063_ = sum_23[74] & q[9] /*9925*/;
  assign _12064_ = m_23[74] & _12062_ /*9924*/;
  assign r_23[74] = _12064_ | _12063_ /*9923*/;
  assign _12065_ = ~q[9] /*9922*/;
  assign _12066_ = sum_23[75] & q[9] /*9921*/;
  assign _12067_ = m_23[75] & _12065_ /*9920*/;
  assign r_23[75] = _12067_ | _12066_ /*9919*/;
  assign _12068_ = ~q[9] /*9918*/;
  assign _12069_ = sum_23[76] & q[9] /*9917*/;
  assign _12070_ = m_23[76] & _12068_ /*9916*/;
  assign r_23[76] = _12070_ | _12069_ /*9915*/;
  assign _12071_ = ~q[9] /*9914*/;
  assign _12072_ = sum_23[77] & q[9] /*9913*/;
  assign _12073_ = m_23[77] & _12071_ /*9912*/;
  assign r_23[77] = _12073_ | _12072_ /*9911*/;
  assign _12074_ = ~q[9] /*9910*/;
  assign _12075_ = sum_23[78] & q[9] /*9909*/;
  assign _12076_ = m_23[78] & _12074_ /*9908*/;
  assign r_23[78] = _12076_ | _12075_ /*9907*/;
  assign _12077_ = ~q[9] /*9906*/;
  assign _12078_ = sum_23[79] & q[9] /*9905*/;
  assign _12079_ = m_23[79] & _12077_ /*9904*/;
  assign r_23[79] = _12079_ | _12078_ /*9903*/;
  assign _12080_ = ~q[9] /*9902*/;
  assign _12081_ = sum_23[80] & q[9] /*9901*/;
  assign _12082_ = m_23[80] & _12080_ /*9900*/;
  assign r_23[80] = _12082_ | _12081_ /*9899*/;
  assign _12083_ = ~q[9] /*9898*/;
  assign _12084_ = sum_23[81] & q[9] /*9897*/;
  assign _12085_ = m_23[81] & _12083_ /*9896*/;
  assign r_23[81] = _12085_ | _12084_ /*9895*/;
  assign _12086_ = ~q[9] /*9894*/;
  assign _12087_ = sum_23[82] & q[9] /*9893*/;
  assign _12088_ = m_23[82] & _12086_ /*9892*/;
  assign r_23[82] = _12088_ | _12087_ /*9891*/;
  assign _12089_ = ~q[9] /*9890*/;
  assign _12090_ = sum_23[83] & q[9] /*9889*/;
  assign _12091_ = m_23[83] & _12089_ /*9888*/;
  assign r_23[83] = _12091_ | _12090_ /*9887*/;
  assign _12092_ = ~q[9] /*9886*/;
  assign _12093_ = sum_23[84] & q[9] /*9885*/;
  assign _12094_ = m_23[84] & _12092_ /*9884*/;
  assign r_23[84] = _12094_ | _12093_ /*9883*/;
  assign _12095_ = ~q[9] /*9882*/;
  assign _12096_ = sum_23[85] & q[9] /*9881*/;
  assign _12097_ = m_23[85] & _12095_ /*9880*/;
  assign r_23[85] = _12097_ | _12096_ /*9879*/;
  assign inv_24[0] = oneWire /*9748*/;
  assign inv_24[1] = oneWire /*9742*/;
  assign inv_24[2] = oneWire /*9736*/;
  assign inv_24[3] = oneWire /*9730*/;
  assign inv_24[4] = oneWire /*9724*/;
  assign inv_24[5] = oneWire /*9718*/;
  assign inv_24[6] = oneWire /*9712*/;
  assign inv_24[7] = oneWire /*9706*/;
  assign inv_24[8] = ~div[0] /*9700*/;
  assign inv_24[9] = ~div[1] /*9694*/;
  assign inv_24[10] = ~div[2] /*9688*/;
  assign inv_24[11] = ~div[3] /*9682*/;
  assign inv_24[12] = ~div[4] /*9676*/;
  assign inv_24[13] = ~div[5] /*9670*/;
  assign inv_24[14] = ~div[6] /*9664*/;
  assign inv_24[15] = ~div[7] /*9658*/;
  assign inv_24[16] = ~div[8] /*9652*/;
  assign inv_24[17] = ~div[9] /*9646*/;
  assign inv_24[18] = ~div[10] /*9640*/;
  assign inv_24[19] = ~div[11] /*9634*/;
  assign inv_24[20] = ~div[12] /*9628*/;
  assign inv_24[21] = ~div[13] /*9622*/;
  assign inv_24[22] = ~div[14] /*9616*/;
  assign inv_24[23] = ~div[15] /*9610*/;
  assign inv_24[24] = ~div[16] /*9604*/;
  assign inv_24[25] = ~div[17] /*9598*/;
  assign inv_24[26] = ~div[18] /*9592*/;
  assign inv_24[27] = ~div[19] /*9586*/;
  assign inv_24[28] = ~div[20] /*9580*/;
  assign inv_24[29] = ~div[21] /*9574*/;
  assign inv_24[30] = ~div[22] /*9568*/;
  assign inv_24[31] = ~div[23] /*9562*/;
  assign inv_24[32] = ~div[24] /*9556*/;
  assign inv_24[33] = ~div[25] /*9550*/;
  assign inv_24[34] = ~div[26] /*9544*/;
  assign inv_24[35] = ~div[27] /*9538*/;
  assign inv_24[36] = ~div[28] /*9532*/;
  assign inv_24[37] = ~div[29] /*9526*/;
  assign inv_24[38] = ~div[30] /*9520*/;
  assign inv_24[39] = oneWire /*9514*/;
  assign inv_24[40] = oneWire /*9508*/;
  assign inv_24[41] = oneWire /*9502*/;
  assign inv_24[42] = oneWire /*9496*/;
  assign inv_24[43] = oneWire /*9490*/;
  assign inv_24[44] = oneWire /*9484*/;
  assign inv_24[45] = oneWire /*9478*/;
  assign inv_24[46] = oneWire /*9472*/;
  assign inv_24[47] = oneWire /*9466*/;
  assign inv_24[48] = oneWire /*9460*/;
  assign inv_24[49] = oneWire /*9454*/;
  assign inv_24[50] = oneWire /*9448*/;
  assign inv_24[51] = oneWire /*9442*/;
  assign inv_24[52] = oneWire /*9436*/;
  assign inv_24[53] = oneWire /*9430*/;
  assign inv_24[54] = oneWire /*9424*/;
  assign inv_24[55] = oneWire /*9418*/;
  assign inv_24[56] = oneWire /*9412*/;
  assign inv_24[57] = oneWire /*9406*/;
  assign inv_24[58] = oneWire /*9400*/;
  assign inv_24[59] = oneWire /*9394*/;
  assign inv_24[60] = oneWire /*9388*/;
  assign inv_24[61] = oneWire /*9382*/;
  assign inv_24[62] = oneWire /*9376*/;
  assign inv_24[63] = oneWire /*9370*/;
  assign inv_24[64] = oneWire /*9364*/;
  assign inv_24[65] = oneWire /*9358*/;
  assign inv_24[66] = oneWire /*9352*/;
  assign inv_24[67] = oneWire /*9346*/;
  assign inv_24[68] = oneWire /*9340*/;
  assign inv_24[69] = oneWire /*9334*/;
  assign inv_24[70] = oneWire /*9328*/;
  assign inv_24[71] = oneWire /*9322*/;
  assign inv_24[72] = oneWire /*9316*/;
  assign inv_24[73] = oneWire /*9310*/;
  assign inv_24[74] = oneWire /*9304*/;
  assign inv_24[75] = oneWire /*9298*/;
  assign inv_24[76] = oneWire /*9292*/;
  assign inv_24[77] = oneWire /*9286*/;
  assign inv_24[78] = oneWire /*9280*/;
  assign inv_24[79] = oneWire /*9274*/;
  assign inv_24[80] = oneWire /*9268*/;
  assign inv_24[81] = oneWire /*9262*/;
  assign inv_24[82] = oneWire /*9256*/;
  assign inv_24[83] = oneWire /*9250*/;
  assign inv_24[84] = oneWire /*9244*/;
  assign inv_24[85] = oneWire /*9238*/;
  assign _12098_ = inv_24[0] ^ r_23[0] /*9747*/;
  assign sum_24[0] = _12098_ ^ oneWire /*9746*/;
  assign _12099_ = _12098_ & oneWire /*9745*/;
  assign _12100_ = inv_24[0] & r_23[0] /*9744*/;
  assign _12101_ = _12099_ | _12100_ /*9743*/;
  assign _12102_ = inv_24[1] ^ r_23[1] /*9741*/;
  assign sum_24[1] = _12102_ ^ _12101_ /*9740*/;
  assign _12103_ = _12102_ & _12101_ /*9739*/;
  assign _12104_ = inv_24[1] & r_23[1] /*9738*/;
  assign _12105_ = _12103_ | _12104_ /*9737*/;
  assign _12106_ = inv_24[2] ^ r_23[2] /*9735*/;
  assign sum_24[2] = _12106_ ^ _12105_ /*9734*/;
  assign _12107_ = _12106_ & _12105_ /*9733*/;
  assign _12108_ = inv_24[2] & r_23[2] /*9732*/;
  assign _12109_ = _12107_ | _12108_ /*9731*/;
  assign _12110_ = inv_24[3] ^ r_23[3] /*9729*/;
  assign sum_24[3] = _12110_ ^ _12109_ /*9728*/;
  assign _12111_ = _12110_ & _12109_ /*9727*/;
  assign _12112_ = inv_24[3] & r_23[3] /*9726*/;
  assign _12113_ = _12111_ | _12112_ /*9725*/;
  assign _12114_ = inv_24[4] ^ r_23[4] /*9723*/;
  assign sum_24[4] = _12114_ ^ _12113_ /*9722*/;
  assign _12115_ = _12114_ & _12113_ /*9721*/;
  assign _12116_ = inv_24[4] & r_23[4] /*9720*/;
  assign _12117_ = _12115_ | _12116_ /*9719*/;
  assign _12118_ = inv_24[5] ^ r_23[5] /*9717*/;
  assign sum_24[5] = _12118_ ^ _12117_ /*9716*/;
  assign _12119_ = _12118_ & _12117_ /*9715*/;
  assign _12120_ = inv_24[5] & r_23[5] /*9714*/;
  assign _12121_ = _12119_ | _12120_ /*9713*/;
  assign _12122_ = inv_24[6] ^ r_23[6] /*9711*/;
  assign sum_24[6] = _12122_ ^ _12121_ /*9710*/;
  assign _12123_ = _12122_ & _12121_ /*9709*/;
  assign _12124_ = inv_24[6] & r_23[6] /*9708*/;
  assign _12125_ = _12123_ | _12124_ /*9707*/;
  assign _12126_ = inv_24[7] ^ r_23[7] /*9705*/;
  assign sum_24[7] = _12126_ ^ _12125_ /*9704*/;
  assign _12127_ = _12126_ & _12125_ /*9703*/;
  assign _12128_ = inv_24[7] & r_23[7] /*9702*/;
  assign _12129_ = _12127_ | _12128_ /*9701*/;
  assign _12130_ = inv_24[8] ^ r_23[8] /*9699*/;
  assign sum_24[8] = _12130_ ^ _12129_ /*9698*/;
  assign _12131_ = _12130_ & _12129_ /*9697*/;
  assign _12132_ = inv_24[8] & r_23[8] /*9696*/;
  assign _12133_ = _12131_ | _12132_ /*9695*/;
  assign _12134_ = inv_24[9] ^ r_23[9] /*9693*/;
  assign sum_24[9] = _12134_ ^ _12133_ /*9692*/;
  assign _12135_ = _12134_ & _12133_ /*9691*/;
  assign _12136_ = inv_24[9] & r_23[9] /*9690*/;
  assign _12137_ = _12135_ | _12136_ /*9689*/;
  assign _12138_ = inv_24[10] ^ r_23[10] /*9687*/;
  assign sum_24[10] = _12138_ ^ _12137_ /*9686*/;
  assign _12139_ = _12138_ & _12137_ /*9685*/;
  assign _12140_ = inv_24[10] & r_23[10] /*9684*/;
  assign _12141_ = _12139_ | _12140_ /*9683*/;
  assign _12142_ = inv_24[11] ^ r_23[11] /*9681*/;
  assign sum_24[11] = _12142_ ^ _12141_ /*9680*/;
  assign _12143_ = _12142_ & _12141_ /*9679*/;
  assign _12144_ = inv_24[11] & r_23[11] /*9678*/;
  assign _12145_ = _12143_ | _12144_ /*9677*/;
  assign _12146_ = inv_24[12] ^ r_23[12] /*9675*/;
  assign sum_24[12] = _12146_ ^ _12145_ /*9674*/;
  assign _12147_ = _12146_ & _12145_ /*9673*/;
  assign _12148_ = inv_24[12] & r_23[12] /*9672*/;
  assign _12149_ = _12147_ | _12148_ /*9671*/;
  assign _12150_ = inv_24[13] ^ r_23[13] /*9669*/;
  assign sum_24[13] = _12150_ ^ _12149_ /*9668*/;
  assign _12151_ = _12150_ & _12149_ /*9667*/;
  assign _12152_ = inv_24[13] & r_23[13] /*9666*/;
  assign _12153_ = _12151_ | _12152_ /*9665*/;
  assign _12154_ = inv_24[14] ^ r_23[14] /*9663*/;
  assign sum_24[14] = _12154_ ^ _12153_ /*9662*/;
  assign _12155_ = _12154_ & _12153_ /*9661*/;
  assign _12156_ = inv_24[14] & r_23[14] /*9660*/;
  assign _12157_ = _12155_ | _12156_ /*9659*/;
  assign _12158_ = inv_24[15] ^ r_23[15] /*9657*/;
  assign sum_24[15] = _12158_ ^ _12157_ /*9656*/;
  assign _12159_ = _12158_ & _12157_ /*9655*/;
  assign _12160_ = inv_24[15] & r_23[15] /*9654*/;
  assign _12161_ = _12159_ | _12160_ /*9653*/;
  assign _12162_ = inv_24[16] ^ r_23[16] /*9651*/;
  assign sum_24[16] = _12162_ ^ _12161_ /*9650*/;
  assign _12163_ = _12162_ & _12161_ /*9649*/;
  assign _12164_ = inv_24[16] & r_23[16] /*9648*/;
  assign _12165_ = _12163_ | _12164_ /*9647*/;
  assign _12166_ = inv_24[17] ^ r_23[17] /*9645*/;
  assign sum_24[17] = _12166_ ^ _12165_ /*9644*/;
  assign _12167_ = _12166_ & _12165_ /*9643*/;
  assign _12168_ = inv_24[17] & r_23[17] /*9642*/;
  assign _12169_ = _12167_ | _12168_ /*9641*/;
  assign _12170_ = inv_24[18] ^ r_23[18] /*9639*/;
  assign sum_24[18] = _12170_ ^ _12169_ /*9638*/;
  assign _12171_ = _12170_ & _12169_ /*9637*/;
  assign _12172_ = inv_24[18] & r_23[18] /*9636*/;
  assign _12173_ = _12171_ | _12172_ /*9635*/;
  assign _12174_ = inv_24[19] ^ r_23[19] /*9633*/;
  assign sum_24[19] = _12174_ ^ _12173_ /*9632*/;
  assign _12175_ = _12174_ & _12173_ /*9631*/;
  assign _12176_ = inv_24[19] & r_23[19] /*9630*/;
  assign _12177_ = _12175_ | _12176_ /*9629*/;
  assign _12178_ = inv_24[20] ^ r_23[20] /*9627*/;
  assign sum_24[20] = _12178_ ^ _12177_ /*9626*/;
  assign _12179_ = _12178_ & _12177_ /*9625*/;
  assign _12180_ = inv_24[20] & r_23[20] /*9624*/;
  assign _12181_ = _12179_ | _12180_ /*9623*/;
  assign _12182_ = inv_24[21] ^ r_23[21] /*9621*/;
  assign sum_24[21] = _12182_ ^ _12181_ /*9620*/;
  assign _12183_ = _12182_ & _12181_ /*9619*/;
  assign _12184_ = inv_24[21] & r_23[21] /*9618*/;
  assign _12185_ = _12183_ | _12184_ /*9617*/;
  assign _12186_ = inv_24[22] ^ r_23[22] /*9615*/;
  assign sum_24[22] = _12186_ ^ _12185_ /*9614*/;
  assign _12187_ = _12186_ & _12185_ /*9613*/;
  assign _12188_ = inv_24[22] & r_23[22] /*9612*/;
  assign _12189_ = _12187_ | _12188_ /*9611*/;
  assign _12190_ = inv_24[23] ^ r_23[23] /*9609*/;
  assign sum_24[23] = _12190_ ^ _12189_ /*9608*/;
  assign _12191_ = _12190_ & _12189_ /*9607*/;
  assign _12192_ = inv_24[23] & r_23[23] /*9606*/;
  assign _12193_ = _12191_ | _12192_ /*9605*/;
  assign _12194_ = inv_24[24] ^ r_23[24] /*9603*/;
  assign sum_24[24] = _12194_ ^ _12193_ /*9602*/;
  assign _12195_ = _12194_ & _12193_ /*9601*/;
  assign _12196_ = inv_24[24] & r_23[24] /*9600*/;
  assign _12197_ = _12195_ | _12196_ /*9599*/;
  assign _12198_ = inv_24[25] ^ r_23[25] /*9597*/;
  assign sum_24[25] = _12198_ ^ _12197_ /*9596*/;
  assign _12199_ = _12198_ & _12197_ /*9595*/;
  assign _12200_ = inv_24[25] & r_23[25] /*9594*/;
  assign _12201_ = _12199_ | _12200_ /*9593*/;
  assign _12202_ = inv_24[26] ^ r_23[26] /*9591*/;
  assign sum_24[26] = _12202_ ^ _12201_ /*9590*/;
  assign _12203_ = _12202_ & _12201_ /*9589*/;
  assign _12204_ = inv_24[26] & r_23[26] /*9588*/;
  assign _12205_ = _12203_ | _12204_ /*9587*/;
  assign _12206_ = inv_24[27] ^ r_23[27] /*9585*/;
  assign sum_24[27] = _12206_ ^ _12205_ /*9584*/;
  assign _12207_ = _12206_ & _12205_ /*9583*/;
  assign _12208_ = inv_24[27] & r_23[27] /*9582*/;
  assign _12209_ = _12207_ | _12208_ /*9581*/;
  assign _12210_ = inv_24[28] ^ r_23[28] /*9579*/;
  assign sum_24[28] = _12210_ ^ _12209_ /*9578*/;
  assign _12211_ = _12210_ & _12209_ /*9577*/;
  assign _12212_ = inv_24[28] & r_23[28] /*9576*/;
  assign _12213_ = _12211_ | _12212_ /*9575*/;
  assign _12214_ = inv_24[29] ^ r_23[29] /*9573*/;
  assign sum_24[29] = _12214_ ^ _12213_ /*9572*/;
  assign _12215_ = _12214_ & _12213_ /*9571*/;
  assign _12216_ = inv_24[29] & r_23[29] /*9570*/;
  assign _12217_ = _12215_ | _12216_ /*9569*/;
  assign _12218_ = inv_24[30] ^ r_23[30] /*9567*/;
  assign sum_24[30] = _12218_ ^ _12217_ /*9566*/;
  assign _12219_ = _12218_ & _12217_ /*9565*/;
  assign _12220_ = inv_24[30] & r_23[30] /*9564*/;
  assign _12221_ = _12219_ | _12220_ /*9563*/;
  assign _12222_ = inv_24[31] ^ r_23[31] /*9561*/;
  assign sum_24[31] = _12222_ ^ _12221_ /*9560*/;
  assign _12223_ = _12222_ & _12221_ /*9559*/;
  assign _12224_ = inv_24[31] & r_23[31] /*9558*/;
  assign _12225_ = _12223_ | _12224_ /*9557*/;
  assign _12226_ = inv_24[32] ^ r_23[32] /*9555*/;
  assign sum_24[32] = _12226_ ^ _12225_ /*9554*/;
  assign _12227_ = _12226_ & _12225_ /*9553*/;
  assign _12228_ = inv_24[32] & r_23[32] /*9552*/;
  assign _12229_ = _12227_ | _12228_ /*9551*/;
  assign _12230_ = inv_24[33] ^ r_23[33] /*9549*/;
  assign sum_24[33] = _12230_ ^ _12229_ /*9548*/;
  assign _12231_ = _12230_ & _12229_ /*9547*/;
  assign _12232_ = inv_24[33] & r_23[33] /*9546*/;
  assign _12233_ = _12231_ | _12232_ /*9545*/;
  assign _12234_ = inv_24[34] ^ r_23[34] /*9543*/;
  assign sum_24[34] = _12234_ ^ _12233_ /*9542*/;
  assign _12235_ = _12234_ & _12233_ /*9541*/;
  assign _12236_ = inv_24[34] & r_23[34] /*9540*/;
  assign _12237_ = _12235_ | _12236_ /*9539*/;
  assign _12238_ = inv_24[35] ^ r_23[35] /*9537*/;
  assign sum_24[35] = _12238_ ^ _12237_ /*9536*/;
  assign _12239_ = _12238_ & _12237_ /*9535*/;
  assign _12240_ = inv_24[35] & r_23[35] /*9534*/;
  assign _12241_ = _12239_ | _12240_ /*9533*/;
  assign _12242_ = inv_24[36] ^ r_23[36] /*9531*/;
  assign sum_24[36] = _12242_ ^ _12241_ /*9530*/;
  assign _12243_ = _12242_ & _12241_ /*9529*/;
  assign _12244_ = inv_24[36] & r_23[36] /*9528*/;
  assign _12245_ = _12243_ | _12244_ /*9527*/;
  assign _12246_ = inv_24[37] ^ r_23[37] /*9525*/;
  assign sum_24[37] = _12246_ ^ _12245_ /*9524*/;
  assign _12247_ = _12246_ & _12245_ /*9523*/;
  assign _12248_ = inv_24[37] & r_23[37] /*9522*/;
  assign _12249_ = _12247_ | _12248_ /*9521*/;
  assign _12250_ = inv_24[38] ^ r_23[38] /*9519*/;
  assign sum_24[38] = _12250_ ^ _12249_ /*9518*/;
  assign _12251_ = _12250_ & _12249_ /*9517*/;
  assign _12252_ = inv_24[38] & r_23[38] /*9516*/;
  assign _12253_ = _12251_ | _12252_ /*9515*/;
  assign _12254_ = inv_24[39] ^ r_23[39] /*9513*/;
  assign sum_24[39] = _12254_ ^ _12253_ /*9512*/;
  assign _12255_ = _12254_ & _12253_ /*9511*/;
  assign _12256_ = inv_24[39] & r_23[39] /*9510*/;
  assign _12257_ = _12255_ | _12256_ /*9509*/;
  assign _12258_ = inv_24[40] ^ r_23[40] /*9507*/;
  assign sum_24[40] = _12258_ ^ _12257_ /*9506*/;
  assign _12259_ = _12258_ & _12257_ /*9505*/;
  assign _12260_ = inv_24[40] & r_23[40] /*9504*/;
  assign _12261_ = _12259_ | _12260_ /*9503*/;
  assign _12262_ = inv_24[41] ^ r_23[41] /*9501*/;
  assign sum_24[41] = _12262_ ^ _12261_ /*9500*/;
  assign _12263_ = _12262_ & _12261_ /*9499*/;
  assign _12264_ = inv_24[41] & r_23[41] /*9498*/;
  assign _12265_ = _12263_ | _12264_ /*9497*/;
  assign _12266_ = inv_24[42] ^ r_23[42] /*9495*/;
  assign sum_24[42] = _12266_ ^ _12265_ /*9494*/;
  assign _12267_ = _12266_ & _12265_ /*9493*/;
  assign _12268_ = inv_24[42] & r_23[42] /*9492*/;
  assign _12269_ = _12267_ | _12268_ /*9491*/;
  assign _12270_ = inv_24[43] ^ r_23[43] /*9489*/;
  assign sum_24[43] = _12270_ ^ _12269_ /*9488*/;
  assign _12271_ = _12270_ & _12269_ /*9487*/;
  assign _12272_ = inv_24[43] & r_23[43] /*9486*/;
  assign _12273_ = _12271_ | _12272_ /*9485*/;
  assign _12274_ = inv_24[44] ^ r_23[44] /*9483*/;
  assign sum_24[44] = _12274_ ^ _12273_ /*9482*/;
  assign _12275_ = _12274_ & _12273_ /*9481*/;
  assign _12276_ = inv_24[44] & r_23[44] /*9480*/;
  assign _12277_ = _12275_ | _12276_ /*9479*/;
  assign _12278_ = inv_24[45] ^ r_23[45] /*9477*/;
  assign sum_24[45] = _12278_ ^ _12277_ /*9476*/;
  assign _12279_ = _12278_ & _12277_ /*9475*/;
  assign _12280_ = inv_24[45] & r_23[45] /*9474*/;
  assign _12281_ = _12279_ | _12280_ /*9473*/;
  assign _12282_ = inv_24[46] ^ r_23[46] /*9471*/;
  assign sum_24[46] = _12282_ ^ _12281_ /*9470*/;
  assign _12283_ = _12282_ & _12281_ /*9469*/;
  assign _12284_ = inv_24[46] & r_23[46] /*9468*/;
  assign _12285_ = _12283_ | _12284_ /*9467*/;
  assign _12286_ = inv_24[47] ^ r_23[47] /*9465*/;
  assign sum_24[47] = _12286_ ^ _12285_ /*9464*/;
  assign _12287_ = _12286_ & _12285_ /*9463*/;
  assign _12288_ = inv_24[47] & r_23[47] /*9462*/;
  assign _12289_ = _12287_ | _12288_ /*9461*/;
  assign _12290_ = inv_24[48] ^ r_23[48] /*9459*/;
  assign sum_24[48] = _12290_ ^ _12289_ /*9458*/;
  assign _12291_ = _12290_ & _12289_ /*9457*/;
  assign _12292_ = inv_24[48] & r_23[48] /*9456*/;
  assign _12293_ = _12291_ | _12292_ /*9455*/;
  assign _12294_ = inv_24[49] ^ r_23[49] /*9453*/;
  assign sum_24[49] = _12294_ ^ _12293_ /*9452*/;
  assign _12295_ = _12294_ & _12293_ /*9451*/;
  assign _12296_ = inv_24[49] & r_23[49] /*9450*/;
  assign _12297_ = _12295_ | _12296_ /*9449*/;
  assign _12298_ = inv_24[50] ^ r_23[50] /*9447*/;
  assign sum_24[50] = _12298_ ^ _12297_ /*9446*/;
  assign _12299_ = _12298_ & _12297_ /*9445*/;
  assign _12300_ = inv_24[50] & r_23[50] /*9444*/;
  assign _12301_ = _12299_ | _12300_ /*9443*/;
  assign _12302_ = inv_24[51] ^ r_23[51] /*9441*/;
  assign sum_24[51] = _12302_ ^ _12301_ /*9440*/;
  assign _12303_ = _12302_ & _12301_ /*9439*/;
  assign _12304_ = inv_24[51] & r_23[51] /*9438*/;
  assign _12305_ = _12303_ | _12304_ /*9437*/;
  assign _12306_ = inv_24[52] ^ r_23[52] /*9435*/;
  assign sum_24[52] = _12306_ ^ _12305_ /*9434*/;
  assign _12307_ = _12306_ & _12305_ /*9433*/;
  assign _12308_ = inv_24[52] & r_23[52] /*9432*/;
  assign _12309_ = _12307_ | _12308_ /*9431*/;
  assign _12310_ = inv_24[53] ^ r_23[53] /*9429*/;
  assign sum_24[53] = _12310_ ^ _12309_ /*9428*/;
  assign _12311_ = _12310_ & _12309_ /*9427*/;
  assign _12312_ = inv_24[53] & r_23[53] /*9426*/;
  assign _12313_ = _12311_ | _12312_ /*9425*/;
  assign _12314_ = inv_24[54] ^ r_23[54] /*9423*/;
  assign sum_24[54] = _12314_ ^ _12313_ /*9422*/;
  assign _12315_ = _12314_ & _12313_ /*9421*/;
  assign _12316_ = inv_24[54] & r_23[54] /*9420*/;
  assign _12317_ = _12315_ | _12316_ /*9419*/;
  assign _12318_ = inv_24[55] ^ r_23[55] /*9417*/;
  assign sum_24[55] = _12318_ ^ _12317_ /*9416*/;
  assign _12319_ = _12318_ & _12317_ /*9415*/;
  assign _12320_ = inv_24[55] & r_23[55] /*9414*/;
  assign _12321_ = _12319_ | _12320_ /*9413*/;
  assign _12322_ = inv_24[56] ^ r_23[56] /*9411*/;
  assign sum_24[56] = _12322_ ^ _12321_ /*9410*/;
  assign _12323_ = _12322_ & _12321_ /*9409*/;
  assign _12324_ = inv_24[56] & r_23[56] /*9408*/;
  assign _12325_ = _12323_ | _12324_ /*9407*/;
  assign _12326_ = inv_24[57] ^ r_23[57] /*9405*/;
  assign sum_24[57] = _12326_ ^ _12325_ /*9404*/;
  assign _12327_ = _12326_ & _12325_ /*9403*/;
  assign _12328_ = inv_24[57] & r_23[57] /*9402*/;
  assign _12329_ = _12327_ | _12328_ /*9401*/;
  assign _12330_ = inv_24[58] ^ r_23[58] /*9399*/;
  assign sum_24[58] = _12330_ ^ _12329_ /*9398*/;
  assign _12331_ = _12330_ & _12329_ /*9397*/;
  assign _12332_ = inv_24[58] & r_23[58] /*9396*/;
  assign _12333_ = _12331_ | _12332_ /*9395*/;
  assign _12334_ = inv_24[59] ^ r_23[59] /*9393*/;
  assign sum_24[59] = _12334_ ^ _12333_ /*9392*/;
  assign _12335_ = _12334_ & _12333_ /*9391*/;
  assign _12336_ = inv_24[59] & r_23[59] /*9390*/;
  assign _12337_ = _12335_ | _12336_ /*9389*/;
  assign _12338_ = inv_24[60] ^ r_23[60] /*9387*/;
  assign sum_24[60] = _12338_ ^ _12337_ /*9386*/;
  assign _12339_ = _12338_ & _12337_ /*9385*/;
  assign _12340_ = inv_24[60] & r_23[60] /*9384*/;
  assign _12341_ = _12339_ | _12340_ /*9383*/;
  assign _12342_ = inv_24[61] ^ r_23[61] /*9381*/;
  assign sum_24[61] = _12342_ ^ _12341_ /*9380*/;
  assign _12343_ = _12342_ & _12341_ /*9379*/;
  assign _12344_ = inv_24[61] & r_23[61] /*9378*/;
  assign _12345_ = _12343_ | _12344_ /*9377*/;
  assign _12346_ = inv_24[62] ^ r_23[62] /*9375*/;
  assign sum_24[62] = _12346_ ^ _12345_ /*9374*/;
  assign _12347_ = _12346_ & _12345_ /*9373*/;
  assign _12348_ = inv_24[62] & r_23[62] /*9372*/;
  assign _12349_ = _12347_ | _12348_ /*9371*/;
  assign _12350_ = inv_24[63] ^ r_23[63] /*9369*/;
  assign sum_24[63] = _12350_ ^ _12349_ /*9368*/;
  assign _12351_ = _12350_ & _12349_ /*9367*/;
  assign _12352_ = inv_24[63] & r_23[63] /*9366*/;
  assign _12353_ = _12351_ | _12352_ /*9365*/;
  assign _12354_ = inv_24[64] ^ r_23[64] /*9363*/;
  assign sum_24[64] = _12354_ ^ _12353_ /*9362*/;
  assign _12355_ = _12354_ & _12353_ /*9361*/;
  assign _12356_ = inv_24[64] & r_23[64] /*9360*/;
  assign _12357_ = _12355_ | _12356_ /*9359*/;
  assign _12358_ = inv_24[65] ^ r_23[65] /*9357*/;
  assign sum_24[65] = _12358_ ^ _12357_ /*9356*/;
  assign _12359_ = _12358_ & _12357_ /*9355*/;
  assign _12360_ = inv_24[65] & r_23[65] /*9354*/;
  assign _12361_ = _12359_ | _12360_ /*9353*/;
  assign _12362_ = inv_24[66] ^ r_23[66] /*9351*/;
  assign sum_24[66] = _12362_ ^ _12361_ /*9350*/;
  assign _12363_ = _12362_ & _12361_ /*9349*/;
  assign _12364_ = inv_24[66] & r_23[66] /*9348*/;
  assign _12365_ = _12363_ | _12364_ /*9347*/;
  assign _12366_ = inv_24[67] ^ r_23[67] /*9345*/;
  assign sum_24[67] = _12366_ ^ _12365_ /*9344*/;
  assign _12367_ = _12366_ & _12365_ /*9343*/;
  assign _12368_ = inv_24[67] & r_23[67] /*9342*/;
  assign _12369_ = _12367_ | _12368_ /*9341*/;
  assign _12370_ = inv_24[68] ^ r_23[68] /*9339*/;
  assign sum_24[68] = _12370_ ^ _12369_ /*9338*/;
  assign _12371_ = _12370_ & _12369_ /*9337*/;
  assign _12372_ = inv_24[68] & r_23[68] /*9336*/;
  assign _12373_ = _12371_ | _12372_ /*9335*/;
  assign _12374_ = inv_24[69] ^ r_23[69] /*9333*/;
  assign sum_24[69] = _12374_ ^ _12373_ /*9332*/;
  assign _12375_ = _12374_ & _12373_ /*9331*/;
  assign _12376_ = inv_24[69] & r_23[69] /*9330*/;
  assign _12377_ = _12375_ | _12376_ /*9329*/;
  assign _12378_ = inv_24[70] ^ r_23[70] /*9327*/;
  assign sum_24[70] = _12378_ ^ _12377_ /*9326*/;
  assign _12379_ = _12378_ & _12377_ /*9325*/;
  assign _12380_ = inv_24[70] & r_23[70] /*9324*/;
  assign _12381_ = _12379_ | _12380_ /*9323*/;
  assign _12382_ = inv_24[71] ^ r_23[71] /*9321*/;
  assign sum_24[71] = _12382_ ^ _12381_ /*9320*/;
  assign _12383_ = _12382_ & _12381_ /*9319*/;
  assign _12384_ = inv_24[71] & r_23[71] /*9318*/;
  assign _12385_ = _12383_ | _12384_ /*9317*/;
  assign _12386_ = inv_24[72] ^ r_23[72] /*9315*/;
  assign sum_24[72] = _12386_ ^ _12385_ /*9314*/;
  assign _12387_ = _12386_ & _12385_ /*9313*/;
  assign _12388_ = inv_24[72] & r_23[72] /*9312*/;
  assign _12389_ = _12387_ | _12388_ /*9311*/;
  assign _12390_ = inv_24[73] ^ r_23[73] /*9309*/;
  assign sum_24[73] = _12390_ ^ _12389_ /*9308*/;
  assign _12391_ = _12390_ & _12389_ /*9307*/;
  assign _12392_ = inv_24[73] & r_23[73] /*9306*/;
  assign _12393_ = _12391_ | _12392_ /*9305*/;
  assign _12394_ = inv_24[74] ^ r_23[74] /*9303*/;
  assign sum_24[74] = _12394_ ^ _12393_ /*9302*/;
  assign _12395_ = _12394_ & _12393_ /*9301*/;
  assign _12396_ = inv_24[74] & r_23[74] /*9300*/;
  assign _12397_ = _12395_ | _12396_ /*9299*/;
  assign _12398_ = inv_24[75] ^ r_23[75] /*9297*/;
  assign sum_24[75] = _12398_ ^ _12397_ /*9296*/;
  assign _12399_ = _12398_ & _12397_ /*9295*/;
  assign _12400_ = inv_24[75] & r_23[75] /*9294*/;
  assign _12401_ = _12399_ | _12400_ /*9293*/;
  assign _12402_ = inv_24[76] ^ r_23[76] /*9291*/;
  assign sum_24[76] = _12402_ ^ _12401_ /*9290*/;
  assign _12403_ = _12402_ & _12401_ /*9289*/;
  assign _12404_ = inv_24[76] & r_23[76] /*9288*/;
  assign _12405_ = _12403_ | _12404_ /*9287*/;
  assign _12406_ = inv_24[77] ^ r_23[77] /*9285*/;
  assign sum_24[77] = _12406_ ^ _12405_ /*9284*/;
  assign _12407_ = _12406_ & _12405_ /*9283*/;
  assign _12408_ = inv_24[77] & r_23[77] /*9282*/;
  assign _12409_ = _12407_ | _12408_ /*9281*/;
  assign _12410_ = inv_24[78] ^ r_23[78] /*9279*/;
  assign sum_24[78] = _12410_ ^ _12409_ /*9278*/;
  assign _12411_ = _12410_ & _12409_ /*9277*/;
  assign _12412_ = inv_24[78] & r_23[78] /*9276*/;
  assign _12413_ = _12411_ | _12412_ /*9275*/;
  assign _12414_ = inv_24[79] ^ r_23[79] /*9273*/;
  assign sum_24[79] = _12414_ ^ _12413_ /*9272*/;
  assign _12415_ = _12414_ & _12413_ /*9271*/;
  assign _12416_ = inv_24[79] & r_23[79] /*9270*/;
  assign _12417_ = _12415_ | _12416_ /*9269*/;
  assign _12418_ = inv_24[80] ^ r_23[80] /*9267*/;
  assign sum_24[80] = _12418_ ^ _12417_ /*9266*/;
  assign _12419_ = _12418_ & _12417_ /*9265*/;
  assign _12420_ = inv_24[80] & r_23[80] /*9264*/;
  assign _12421_ = _12419_ | _12420_ /*9263*/;
  assign _12422_ = inv_24[81] ^ r_23[81] /*9261*/;
  assign sum_24[81] = _12422_ ^ _12421_ /*9260*/;
  assign _12423_ = _12422_ & _12421_ /*9259*/;
  assign _12424_ = inv_24[81] & r_23[81] /*9258*/;
  assign _12425_ = _12423_ | _12424_ /*9257*/;
  assign _12426_ = inv_24[82] ^ r_23[82] /*9255*/;
  assign sum_24[82] = _12426_ ^ _12425_ /*9254*/;
  assign _12427_ = _12426_ & _12425_ /*9253*/;
  assign _12428_ = inv_24[82] & r_23[82] /*9252*/;
  assign _12429_ = _12427_ | _12428_ /*9251*/;
  assign _12430_ = inv_24[83] ^ r_23[83] /*9249*/;
  assign sum_24[83] = _12430_ ^ _12429_ /*9248*/;
  assign _12431_ = _12430_ & _12429_ /*9247*/;
  assign _12432_ = inv_24[83] & r_23[83] /*9246*/;
  assign _12433_ = _12431_ | _12432_ /*9245*/;
  assign _12434_ = inv_24[84] ^ r_23[84] /*9243*/;
  assign sum_24[84] = _12434_ ^ _12433_ /*9242*/;
  assign _12435_ = _12434_ & _12433_ /*9241*/;
  assign _12436_ = inv_24[84] & r_23[84] /*9240*/;
  assign _12437_ = _12435_ | _12436_ /*9239*/;
  assign _12438_ = inv_24[85] ^ r_23[85] /*9237*/;
  assign sum_24[85] = _12438_ ^ _12437_ /*9236*/;
  assign _12439_ = _12438_ & _12437_ /*9235*/;
  assign _12440_ = inv_24[85] & r_23[85] /*9234*/;
  assign _12441_ = _12439_ | _12440_ /*9233*/;
  assign _12442_ = _12441_ ^ _12437_ /*9232*/;
  assign _12443_ = ~_12442_ /*9231*/;
  assign _12444_ = sum_24[85] & _12443_ /*9230*/;
  assign _12445_ = _12442_ & _12441_ /*9229*/;
  assign sum_24[86] = _12445_ | _12444_ /*9228*/;
  assign q[8] = ~sum_24[86] /*9227*/;
  assign m_24[0] = r_23[0] /*9226*/;
  assign m_24[1] = r_23[1] /*9225*/;
  assign m_24[2] = r_23[2] /*9224*/;
  assign m_24[3] = r_23[3] /*9223*/;
  assign m_24[4] = r_23[4] /*9222*/;
  assign m_24[5] = r_23[5] /*9221*/;
  assign m_24[6] = r_23[6] /*9220*/;
  assign m_24[7] = r_23[7] /*9219*/;
  assign m_24[8] = r_23[8] /*9218*/;
  assign m_24[9] = r_23[9] /*9217*/;
  assign m_24[10] = r_23[10] /*9216*/;
  assign m_24[11] = r_23[11] /*9215*/;
  assign m_24[12] = r_23[12] /*9214*/;
  assign m_24[13] = r_23[13] /*9213*/;
  assign m_24[14] = r_23[14] /*9212*/;
  assign m_24[15] = r_23[15] /*9211*/;
  assign m_24[16] = r_23[16] /*9210*/;
  assign m_24[17] = r_23[17] /*9209*/;
  assign m_24[18] = r_23[18] /*9208*/;
  assign m_24[19] = r_23[19] /*9207*/;
  assign m_24[20] = r_23[20] /*9206*/;
  assign m_24[21] = r_23[21] /*9205*/;
  assign m_24[22] = r_23[22] /*9204*/;
  assign m_24[23] = r_23[23] /*9203*/;
  assign m_24[24] = r_23[24] /*9202*/;
  assign m_24[25] = r_23[25] /*9201*/;
  assign m_24[26] = r_23[26] /*9200*/;
  assign m_24[27] = r_23[27] /*9199*/;
  assign m_24[28] = r_23[28] /*9198*/;
  assign m_24[29] = r_23[29] /*9197*/;
  assign m_24[30] = r_23[30] /*9196*/;
  assign m_24[31] = r_23[31] /*9195*/;
  assign m_24[32] = r_23[32] /*9194*/;
  assign m_24[33] = r_23[33] /*9193*/;
  assign m_24[34] = r_23[34] /*9192*/;
  assign m_24[35] = r_23[35] /*9191*/;
  assign m_24[36] = r_23[36] /*9190*/;
  assign m_24[37] = r_23[37] /*9189*/;
  assign m_24[38] = r_23[38] /*9188*/;
  assign m_24[39] = r_23[39] /*9187*/;
  assign m_24[40] = r_23[40] /*9186*/;
  assign m_24[41] = r_23[41] /*9185*/;
  assign m_24[42] = r_23[42] /*9184*/;
  assign m_24[43] = r_23[43] /*9183*/;
  assign m_24[44] = r_23[44] /*9182*/;
  assign m_24[45] = r_23[45] /*9181*/;
  assign m_24[46] = r_23[46] /*9180*/;
  assign m_24[47] = r_23[47] /*9179*/;
  assign m_24[48] = r_23[48] /*9178*/;
  assign m_24[49] = r_23[49] /*9177*/;
  assign m_24[50] = r_23[50] /*9176*/;
  assign m_24[51] = r_23[51] /*9175*/;
  assign m_24[52] = r_23[52] /*9174*/;
  assign m_24[53] = r_23[53] /*9173*/;
  assign m_24[54] = r_23[54] /*9172*/;
  assign m_24[55] = r_23[55] /*9171*/;
  assign m_24[56] = r_23[56] /*9170*/;
  assign m_24[57] = r_23[57] /*9169*/;
  assign m_24[58] = r_23[58] /*9168*/;
  assign m_24[59] = r_23[59] /*9167*/;
  assign m_24[60] = r_23[60] /*9166*/;
  assign m_24[61] = r_23[61] /*9165*/;
  assign m_24[62] = r_23[62] /*9164*/;
  assign m_24[63] = r_23[63] /*9163*/;
  assign m_24[64] = r_23[64] /*9162*/;
  assign m_24[65] = r_23[65] /*9161*/;
  assign m_24[66] = r_23[66] /*9160*/;
  assign m_24[67] = r_23[67] /*9159*/;
  assign m_24[68] = r_23[68] /*9158*/;
  assign m_24[69] = r_23[69] /*9157*/;
  assign m_24[70] = r_23[70] /*9156*/;
  assign m_24[71] = r_23[71] /*9155*/;
  assign m_24[72] = r_23[72] /*9154*/;
  assign m_24[73] = r_23[73] /*9153*/;
  assign m_24[74] = r_23[74] /*9152*/;
  assign m_24[75] = r_23[75] /*9151*/;
  assign m_24[76] = r_23[76] /*9150*/;
  assign m_24[77] = r_23[77] /*9149*/;
  assign m_24[78] = r_23[78] /*9148*/;
  assign m_24[79] = r_23[79] /*9147*/;
  assign m_24[80] = r_23[80] /*9146*/;
  assign m_24[81] = r_23[81] /*9145*/;
  assign m_24[82] = r_23[82] /*9144*/;
  assign m_24[83] = r_23[83] /*9143*/;
  assign m_24[84] = r_23[84] /*9142*/;
  assign m_24[85] = r_23[85] /*9141*/;
  assign m_24[86] = r_23[85] /*9140*/;
  assign _12447_ = ~q[8] /*9139*/;
  assign _12448_ = sum_24[0] & q[8] /*9138*/;
  assign _12449_ = m_24[0] & _12447_ /*9137*/;
  assign r_24[0] = _12449_ | _12448_ /*9136*/;
  assign _12450_ = ~q[8] /*9135*/;
  assign _12451_ = sum_24[1] & q[8] /*9134*/;
  assign _12452_ = m_24[1] & _12450_ /*9133*/;
  assign r_24[1] = _12452_ | _12451_ /*9132*/;
  assign _12453_ = ~q[8] /*9131*/;
  assign _12454_ = sum_24[2] & q[8] /*9130*/;
  assign _12455_ = m_24[2] & _12453_ /*9129*/;
  assign r_24[2] = _12455_ | _12454_ /*9128*/;
  assign _12456_ = ~q[8] /*9127*/;
  assign _12457_ = sum_24[3] & q[8] /*9126*/;
  assign _12458_ = m_24[3] & _12456_ /*9125*/;
  assign r_24[3] = _12458_ | _12457_ /*9124*/;
  assign _12459_ = ~q[8] /*9123*/;
  assign _12460_ = sum_24[4] & q[8] /*9122*/;
  assign _12461_ = m_24[4] & _12459_ /*9121*/;
  assign r_24[4] = _12461_ | _12460_ /*9120*/;
  assign _12462_ = ~q[8] /*9119*/;
  assign _12463_ = sum_24[5] & q[8] /*9118*/;
  assign _12464_ = m_24[5] & _12462_ /*9117*/;
  assign r_24[5] = _12464_ | _12463_ /*9116*/;
  assign _12465_ = ~q[8] /*9115*/;
  assign _12466_ = sum_24[6] & q[8] /*9114*/;
  assign _12467_ = m_24[6] & _12465_ /*9113*/;
  assign r_24[6] = _12467_ | _12466_ /*9112*/;
  assign _12468_ = ~q[8] /*9111*/;
  assign _12469_ = sum_24[7] & q[8] /*9110*/;
  assign _12470_ = m_24[7] & _12468_ /*9109*/;
  assign r_24[7] = _12470_ | _12469_ /*9108*/;
  assign _12471_ = ~q[8] /*9107*/;
  assign _12472_ = sum_24[8] & q[8] /*9106*/;
  assign _12473_ = m_24[8] & _12471_ /*9105*/;
  assign r_24[8] = _12473_ | _12472_ /*9104*/;
  assign _12474_ = ~q[8] /*9103*/;
  assign _12475_ = sum_24[9] & q[8] /*9102*/;
  assign _12476_ = m_24[9] & _12474_ /*9101*/;
  assign r_24[9] = _12476_ | _12475_ /*9100*/;
  assign _12477_ = ~q[8] /*9099*/;
  assign _12478_ = sum_24[10] & q[8] /*9098*/;
  assign _12479_ = m_24[10] & _12477_ /*9097*/;
  assign r_24[10] = _12479_ | _12478_ /*9096*/;
  assign _12480_ = ~q[8] /*9095*/;
  assign _12481_ = sum_24[11] & q[8] /*9094*/;
  assign _12482_ = m_24[11] & _12480_ /*9093*/;
  assign r_24[11] = _12482_ | _12481_ /*9092*/;
  assign _12483_ = ~q[8] /*9091*/;
  assign _12484_ = sum_24[12] & q[8] /*9090*/;
  assign _12485_ = m_24[12] & _12483_ /*9089*/;
  assign r_24[12] = _12485_ | _12484_ /*9088*/;
  assign _12486_ = ~q[8] /*9087*/;
  assign _12487_ = sum_24[13] & q[8] /*9086*/;
  assign _12488_ = m_24[13] & _12486_ /*9085*/;
  assign r_24[13] = _12488_ | _12487_ /*9084*/;
  assign _12489_ = ~q[8] /*9083*/;
  assign _12490_ = sum_24[14] & q[8] /*9082*/;
  assign _12491_ = m_24[14] & _12489_ /*9081*/;
  assign r_24[14] = _12491_ | _12490_ /*9080*/;
  assign _12492_ = ~q[8] /*9079*/;
  assign _12493_ = sum_24[15] & q[8] /*9078*/;
  assign _12494_ = m_24[15] & _12492_ /*9077*/;
  assign r_24[15] = _12494_ | _12493_ /*9076*/;
  assign _12495_ = ~q[8] /*9075*/;
  assign _12496_ = sum_24[16] & q[8] /*9074*/;
  assign _12497_ = m_24[16] & _12495_ /*9073*/;
  assign r_24[16] = _12497_ | _12496_ /*9072*/;
  assign _12498_ = ~q[8] /*9071*/;
  assign _12499_ = sum_24[17] & q[8] /*9070*/;
  assign _12500_ = m_24[17] & _12498_ /*9069*/;
  assign r_24[17] = _12500_ | _12499_ /*9068*/;
  assign _12501_ = ~q[8] /*9067*/;
  assign _12502_ = sum_24[18] & q[8] /*9066*/;
  assign _12503_ = m_24[18] & _12501_ /*9065*/;
  assign r_24[18] = _12503_ | _12502_ /*9064*/;
  assign _12504_ = ~q[8] /*9063*/;
  assign _12505_ = sum_24[19] & q[8] /*9062*/;
  assign _12506_ = m_24[19] & _12504_ /*9061*/;
  assign r_24[19] = _12506_ | _12505_ /*9060*/;
  assign _12507_ = ~q[8] /*9059*/;
  assign _12508_ = sum_24[20] & q[8] /*9058*/;
  assign _12509_ = m_24[20] & _12507_ /*9057*/;
  assign r_24[20] = _12509_ | _12508_ /*9056*/;
  assign _12510_ = ~q[8] /*9055*/;
  assign _12511_ = sum_24[21] & q[8] /*9054*/;
  assign _12512_ = m_24[21] & _12510_ /*9053*/;
  assign r_24[21] = _12512_ | _12511_ /*9052*/;
  assign _12513_ = ~q[8] /*9051*/;
  assign _12514_ = sum_24[22] & q[8] /*9050*/;
  assign _12515_ = m_24[22] & _12513_ /*9049*/;
  assign r_24[22] = _12515_ | _12514_ /*9048*/;
  assign _12516_ = ~q[8] /*9047*/;
  assign _12517_ = sum_24[23] & q[8] /*9046*/;
  assign _12518_ = m_24[23] & _12516_ /*9045*/;
  assign r_24[23] = _12518_ | _12517_ /*9044*/;
  assign _12519_ = ~q[8] /*9043*/;
  assign _12520_ = sum_24[24] & q[8] /*9042*/;
  assign _12521_ = m_24[24] & _12519_ /*9041*/;
  assign r_24[24] = _12521_ | _12520_ /*9040*/;
  assign _12522_ = ~q[8] /*9039*/;
  assign _12523_ = sum_24[25] & q[8] /*9038*/;
  assign _12524_ = m_24[25] & _12522_ /*9037*/;
  assign r_24[25] = _12524_ | _12523_ /*9036*/;
  assign _12525_ = ~q[8] /*9035*/;
  assign _12526_ = sum_24[26] & q[8] /*9034*/;
  assign _12527_ = m_24[26] & _12525_ /*9033*/;
  assign r_24[26] = _12527_ | _12526_ /*9032*/;
  assign _12528_ = ~q[8] /*9031*/;
  assign _12529_ = sum_24[27] & q[8] /*9030*/;
  assign _12530_ = m_24[27] & _12528_ /*9029*/;
  assign r_24[27] = _12530_ | _12529_ /*9028*/;
  assign _12531_ = ~q[8] /*9027*/;
  assign _12532_ = sum_24[28] & q[8] /*9026*/;
  assign _12533_ = m_24[28] & _12531_ /*9025*/;
  assign r_24[28] = _12533_ | _12532_ /*9024*/;
  assign _12534_ = ~q[8] /*9023*/;
  assign _12535_ = sum_24[29] & q[8] /*9022*/;
  assign _12536_ = m_24[29] & _12534_ /*9021*/;
  assign r_24[29] = _12536_ | _12535_ /*9020*/;
  assign _12537_ = ~q[8] /*9019*/;
  assign _12538_ = sum_24[30] & q[8] /*9018*/;
  assign _12539_ = m_24[30] & _12537_ /*9017*/;
  assign r_24[30] = _12539_ | _12538_ /*9016*/;
  assign _12540_ = ~q[8] /*9015*/;
  assign _12541_ = sum_24[31] & q[8] /*9014*/;
  assign _12542_ = m_24[31] & _12540_ /*9013*/;
  assign r_24[31] = _12542_ | _12541_ /*9012*/;
  assign _12543_ = ~q[8] /*9011*/;
  assign _12544_ = sum_24[32] & q[8] /*9010*/;
  assign _12545_ = m_24[32] & _12543_ /*9009*/;
  assign r_24[32] = _12545_ | _12544_ /*9008*/;
  assign _12546_ = ~q[8] /*9007*/;
  assign _12547_ = sum_24[33] & q[8] /*9006*/;
  assign _12548_ = m_24[33] & _12546_ /*9005*/;
  assign r_24[33] = _12548_ | _12547_ /*9004*/;
  assign _12549_ = ~q[8] /*9003*/;
  assign _12550_ = sum_24[34] & q[8] /*9002*/;
  assign _12551_ = m_24[34] & _12549_ /*9001*/;
  assign r_24[34] = _12551_ | _12550_ /*9000*/;
  assign _12552_ = ~q[8] /*8999*/;
  assign _12553_ = sum_24[35] & q[8] /*8998*/;
  assign _12554_ = m_24[35] & _12552_ /*8997*/;
  assign r_24[35] = _12554_ | _12553_ /*8996*/;
  assign _12555_ = ~q[8] /*8995*/;
  assign _12556_ = sum_24[36] & q[8] /*8994*/;
  assign _12557_ = m_24[36] & _12555_ /*8993*/;
  assign r_24[36] = _12557_ | _12556_ /*8992*/;
  assign _12558_ = ~q[8] /*8991*/;
  assign _12559_ = sum_24[37] & q[8] /*8990*/;
  assign _12560_ = m_24[37] & _12558_ /*8989*/;
  assign r_24[37] = _12560_ | _12559_ /*8988*/;
  assign _12561_ = ~q[8] /*8987*/;
  assign _12562_ = sum_24[38] & q[8] /*8986*/;
  assign _12563_ = m_24[38] & _12561_ /*8985*/;
  assign r_24[38] = _12563_ | _12562_ /*8984*/;
  assign _12564_ = ~q[8] /*8983*/;
  assign _12565_ = sum_24[39] & q[8] /*8982*/;
  assign _12566_ = m_24[39] & _12564_ /*8981*/;
  assign r_24[39] = _12566_ | _12565_ /*8980*/;
  assign _12567_ = ~q[8] /*8979*/;
  assign _12568_ = sum_24[40] & q[8] /*8978*/;
  assign _12569_ = m_24[40] & _12567_ /*8977*/;
  assign r_24[40] = _12569_ | _12568_ /*8976*/;
  assign _12570_ = ~q[8] /*8975*/;
  assign _12571_ = sum_24[41] & q[8] /*8974*/;
  assign _12572_ = m_24[41] & _12570_ /*8973*/;
  assign r_24[41] = _12572_ | _12571_ /*8972*/;
  assign _12573_ = ~q[8] /*8971*/;
  assign _12574_ = sum_24[42] & q[8] /*8970*/;
  assign _12575_ = m_24[42] & _12573_ /*8969*/;
  assign r_24[42] = _12575_ | _12574_ /*8968*/;
  assign _12576_ = ~q[8] /*8967*/;
  assign _12577_ = sum_24[43] & q[8] /*8966*/;
  assign _12578_ = m_24[43] & _12576_ /*8965*/;
  assign r_24[43] = _12578_ | _12577_ /*8964*/;
  assign _12579_ = ~q[8] /*8963*/;
  assign _12580_ = sum_24[44] & q[8] /*8962*/;
  assign _12581_ = m_24[44] & _12579_ /*8961*/;
  assign r_24[44] = _12581_ | _12580_ /*8960*/;
  assign _12582_ = ~q[8] /*8959*/;
  assign _12583_ = sum_24[45] & q[8] /*8958*/;
  assign _12584_ = m_24[45] & _12582_ /*8957*/;
  assign r_24[45] = _12584_ | _12583_ /*8956*/;
  assign _12585_ = ~q[8] /*8955*/;
  assign _12586_ = sum_24[46] & q[8] /*8954*/;
  assign _12587_ = m_24[46] & _12585_ /*8953*/;
  assign r_24[46] = _12587_ | _12586_ /*8952*/;
  assign _12588_ = ~q[8] /*8951*/;
  assign _12589_ = sum_24[47] & q[8] /*8950*/;
  assign _12590_ = m_24[47] & _12588_ /*8949*/;
  assign r_24[47] = _12590_ | _12589_ /*8948*/;
  assign _12591_ = ~q[8] /*8947*/;
  assign _12592_ = sum_24[48] & q[8] /*8946*/;
  assign _12593_ = m_24[48] & _12591_ /*8945*/;
  assign r_24[48] = _12593_ | _12592_ /*8944*/;
  assign _12594_ = ~q[8] /*8943*/;
  assign _12595_ = sum_24[49] & q[8] /*8942*/;
  assign _12596_ = m_24[49] & _12594_ /*8941*/;
  assign r_24[49] = _12596_ | _12595_ /*8940*/;
  assign _12597_ = ~q[8] /*8939*/;
  assign _12598_ = sum_24[50] & q[8] /*8938*/;
  assign _12599_ = m_24[50] & _12597_ /*8937*/;
  assign r_24[50] = _12599_ | _12598_ /*8936*/;
  assign _12600_ = ~q[8] /*8935*/;
  assign _12601_ = sum_24[51] & q[8] /*8934*/;
  assign _12602_ = m_24[51] & _12600_ /*8933*/;
  assign r_24[51] = _12602_ | _12601_ /*8932*/;
  assign _12603_ = ~q[8] /*8931*/;
  assign _12604_ = sum_24[52] & q[8] /*8930*/;
  assign _12605_ = m_24[52] & _12603_ /*8929*/;
  assign r_24[52] = _12605_ | _12604_ /*8928*/;
  assign _12606_ = ~q[8] /*8927*/;
  assign _12607_ = sum_24[53] & q[8] /*8926*/;
  assign _12608_ = m_24[53] & _12606_ /*8925*/;
  assign r_24[53] = _12608_ | _12607_ /*8924*/;
  assign _12609_ = ~q[8] /*8923*/;
  assign _12610_ = sum_24[54] & q[8] /*8922*/;
  assign _12611_ = m_24[54] & _12609_ /*8921*/;
  assign r_24[54] = _12611_ | _12610_ /*8920*/;
  assign _12612_ = ~q[8] /*8919*/;
  assign _12613_ = sum_24[55] & q[8] /*8918*/;
  assign _12614_ = m_24[55] & _12612_ /*8917*/;
  assign r_24[55] = _12614_ | _12613_ /*8916*/;
  assign _12615_ = ~q[8] /*8915*/;
  assign _12616_ = sum_24[56] & q[8] /*8914*/;
  assign _12617_ = m_24[56] & _12615_ /*8913*/;
  assign r_24[56] = _12617_ | _12616_ /*8912*/;
  assign _12618_ = ~q[8] /*8911*/;
  assign _12619_ = sum_24[57] & q[8] /*8910*/;
  assign _12620_ = m_24[57] & _12618_ /*8909*/;
  assign r_24[57] = _12620_ | _12619_ /*8908*/;
  assign _12621_ = ~q[8] /*8907*/;
  assign _12622_ = sum_24[58] & q[8] /*8906*/;
  assign _12623_ = m_24[58] & _12621_ /*8905*/;
  assign r_24[58] = _12623_ | _12622_ /*8904*/;
  assign _12624_ = ~q[8] /*8903*/;
  assign _12625_ = sum_24[59] & q[8] /*8902*/;
  assign _12626_ = m_24[59] & _12624_ /*8901*/;
  assign r_24[59] = _12626_ | _12625_ /*8900*/;
  assign _12627_ = ~q[8] /*8899*/;
  assign _12628_ = sum_24[60] & q[8] /*8898*/;
  assign _12629_ = m_24[60] & _12627_ /*8897*/;
  assign r_24[60] = _12629_ | _12628_ /*8896*/;
  assign _12630_ = ~q[8] /*8895*/;
  assign _12631_ = sum_24[61] & q[8] /*8894*/;
  assign _12632_ = m_24[61] & _12630_ /*8893*/;
  assign r_24[61] = _12632_ | _12631_ /*8892*/;
  assign _12633_ = ~q[8] /*8891*/;
  assign _12634_ = sum_24[62] & q[8] /*8890*/;
  assign _12635_ = m_24[62] & _12633_ /*8889*/;
  assign r_24[62] = _12635_ | _12634_ /*8888*/;
  assign _12636_ = ~q[8] /*8887*/;
  assign _12637_ = sum_24[63] & q[8] /*8886*/;
  assign _12638_ = m_24[63] & _12636_ /*8885*/;
  assign r_24[63] = _12638_ | _12637_ /*8884*/;
  assign _12639_ = ~q[8] /*8883*/;
  assign _12640_ = sum_24[64] & q[8] /*8882*/;
  assign _12641_ = m_24[64] & _12639_ /*8881*/;
  assign r_24[64] = _12641_ | _12640_ /*8880*/;
  assign _12642_ = ~q[8] /*8879*/;
  assign _12643_ = sum_24[65] & q[8] /*8878*/;
  assign _12644_ = m_24[65] & _12642_ /*8877*/;
  assign r_24[65] = _12644_ | _12643_ /*8876*/;
  assign _12645_ = ~q[8] /*8875*/;
  assign _12646_ = sum_24[66] & q[8] /*8874*/;
  assign _12647_ = m_24[66] & _12645_ /*8873*/;
  assign r_24[66] = _12647_ | _12646_ /*8872*/;
  assign _12648_ = ~q[8] /*8871*/;
  assign _12649_ = sum_24[67] & q[8] /*8870*/;
  assign _12650_ = m_24[67] & _12648_ /*8869*/;
  assign r_24[67] = _12650_ | _12649_ /*8868*/;
  assign _12651_ = ~q[8] /*8867*/;
  assign _12652_ = sum_24[68] & q[8] /*8866*/;
  assign _12653_ = m_24[68] & _12651_ /*8865*/;
  assign r_24[68] = _12653_ | _12652_ /*8864*/;
  assign _12654_ = ~q[8] /*8863*/;
  assign _12655_ = sum_24[69] & q[8] /*8862*/;
  assign _12656_ = m_24[69] & _12654_ /*8861*/;
  assign r_24[69] = _12656_ | _12655_ /*8860*/;
  assign _12657_ = ~q[8] /*8859*/;
  assign _12658_ = sum_24[70] & q[8] /*8858*/;
  assign _12659_ = m_24[70] & _12657_ /*8857*/;
  assign r_24[70] = _12659_ | _12658_ /*8856*/;
  assign _12660_ = ~q[8] /*8855*/;
  assign _12661_ = sum_24[71] & q[8] /*8854*/;
  assign _12662_ = m_24[71] & _12660_ /*8853*/;
  assign r_24[71] = _12662_ | _12661_ /*8852*/;
  assign _12663_ = ~q[8] /*8851*/;
  assign _12664_ = sum_24[72] & q[8] /*8850*/;
  assign _12665_ = m_24[72] & _12663_ /*8849*/;
  assign r_24[72] = _12665_ | _12664_ /*8848*/;
  assign _12666_ = ~q[8] /*8847*/;
  assign _12667_ = sum_24[73] & q[8] /*8846*/;
  assign _12668_ = m_24[73] & _12666_ /*8845*/;
  assign r_24[73] = _12668_ | _12667_ /*8844*/;
  assign _12669_ = ~q[8] /*8843*/;
  assign _12670_ = sum_24[74] & q[8] /*8842*/;
  assign _12671_ = m_24[74] & _12669_ /*8841*/;
  assign r_24[74] = _12671_ | _12670_ /*8840*/;
  assign _12672_ = ~q[8] /*8839*/;
  assign _12673_ = sum_24[75] & q[8] /*8838*/;
  assign _12674_ = m_24[75] & _12672_ /*8837*/;
  assign r_24[75] = _12674_ | _12673_ /*8836*/;
  assign _12675_ = ~q[8] /*8835*/;
  assign _12676_ = sum_24[76] & q[8] /*8834*/;
  assign _12677_ = m_24[76] & _12675_ /*8833*/;
  assign r_24[76] = _12677_ | _12676_ /*8832*/;
  assign _12678_ = ~q[8] /*8831*/;
  assign _12679_ = sum_24[77] & q[8] /*8830*/;
  assign _12680_ = m_24[77] & _12678_ /*8829*/;
  assign r_24[77] = _12680_ | _12679_ /*8828*/;
  assign _12681_ = ~q[8] /*8827*/;
  assign _12682_ = sum_24[78] & q[8] /*8826*/;
  assign _12683_ = m_24[78] & _12681_ /*8825*/;
  assign r_24[78] = _12683_ | _12682_ /*8824*/;
  assign _12684_ = ~q[8] /*8823*/;
  assign _12685_ = sum_24[79] & q[8] /*8822*/;
  assign _12686_ = m_24[79] & _12684_ /*8821*/;
  assign r_24[79] = _12686_ | _12685_ /*8820*/;
  assign _12687_ = ~q[8] /*8819*/;
  assign _12688_ = sum_24[80] & q[8] /*8818*/;
  assign _12689_ = m_24[80] & _12687_ /*8817*/;
  assign r_24[80] = _12689_ | _12688_ /*8816*/;
  assign _12690_ = ~q[8] /*8815*/;
  assign _12691_ = sum_24[81] & q[8] /*8814*/;
  assign _12692_ = m_24[81] & _12690_ /*8813*/;
  assign r_24[81] = _12692_ | _12691_ /*8812*/;
  assign _12693_ = ~q[8] /*8811*/;
  assign _12694_ = sum_24[82] & q[8] /*8810*/;
  assign _12695_ = m_24[82] & _12693_ /*8809*/;
  assign r_24[82] = _12695_ | _12694_ /*8808*/;
  assign _12696_ = ~q[8] /*8807*/;
  assign _12697_ = sum_24[83] & q[8] /*8806*/;
  assign _12698_ = m_24[83] & _12696_ /*8805*/;
  assign r_24[83] = _12698_ | _12697_ /*8804*/;
  assign _12699_ = ~q[8] /*8803*/;
  assign _12700_ = sum_24[84] & q[8] /*8802*/;
  assign _12701_ = m_24[84] & _12699_ /*8801*/;
  assign r_24[84] = _12701_ | _12700_ /*8800*/;
  assign _12702_ = ~q[8] /*8799*/;
  assign _12703_ = sum_24[85] & q[8] /*8798*/;
  assign _12704_ = m_24[85] & _12702_ /*8797*/;
  assign r_24[85] = _12704_ | _12703_ /*8796*/;
  assign _12705_ = ~q[8] /*8795*/;
  assign _12706_ = sum_24[86] & q[8] /*8794*/;
  assign _12707_ = m_24[86] & _12705_ /*8793*/;
  assign r_24[86] = _12707_ | _12706_ /*8792*/;
  assign inv_25[0] = oneWire /*8672*/;
  assign inv_25[1] = oneWire /*8666*/;
  assign inv_25[2] = oneWire /*8660*/;
  assign inv_25[3] = oneWire /*8654*/;
  assign inv_25[4] = oneWire /*8648*/;
  assign inv_25[5] = oneWire /*8642*/;
  assign inv_25[6] = oneWire /*8636*/;
  assign inv_25[7] = ~div[0] /*8630*/;
  assign inv_25[8] = ~div[1] /*8624*/;
  assign inv_25[9] = ~div[2] /*8618*/;
  assign inv_25[10] = ~div[3] /*8612*/;
  assign inv_25[11] = ~div[4] /*8606*/;
  assign inv_25[12] = ~div[5] /*8600*/;
  assign inv_25[13] = ~div[6] /*8594*/;
  assign inv_25[14] = ~div[7] /*8588*/;
  assign inv_25[15] = ~div[8] /*8582*/;
  assign inv_25[16] = ~div[9] /*8576*/;
  assign inv_25[17] = ~div[10] /*8570*/;
  assign inv_25[18] = ~div[11] /*8564*/;
  assign inv_25[19] = ~div[12] /*8558*/;
  assign inv_25[20] = ~div[13] /*8552*/;
  assign inv_25[21] = ~div[14] /*8546*/;
  assign inv_25[22] = ~div[15] /*8540*/;
  assign inv_25[23] = ~div[16] /*8534*/;
  assign inv_25[24] = ~div[17] /*8528*/;
  assign inv_25[25] = ~div[18] /*8522*/;
  assign inv_25[26] = ~div[19] /*8516*/;
  assign inv_25[27] = ~div[20] /*8510*/;
  assign inv_25[28] = ~div[21] /*8504*/;
  assign inv_25[29] = ~div[22] /*8498*/;
  assign inv_25[30] = ~div[23] /*8492*/;
  assign inv_25[31] = ~div[24] /*8486*/;
  assign inv_25[32] = ~div[25] /*8480*/;
  assign inv_25[33] = ~div[26] /*8474*/;
  assign inv_25[34] = ~div[27] /*8468*/;
  assign inv_25[35] = ~div[28] /*8462*/;
  assign inv_25[36] = ~div[29] /*8456*/;
  assign inv_25[37] = ~div[30] /*8450*/;
  assign inv_25[38] = oneWire /*8444*/;
  assign inv_25[39] = oneWire /*8438*/;
  assign inv_25[40] = oneWire /*8432*/;
  assign inv_25[41] = oneWire /*8426*/;
  assign inv_25[42] = oneWire /*8420*/;
  assign inv_25[43] = oneWire /*8414*/;
  assign inv_25[44] = oneWire /*8408*/;
  assign inv_25[45] = oneWire /*8402*/;
  assign inv_25[46] = oneWire /*8396*/;
  assign inv_25[47] = oneWire /*8390*/;
  assign inv_25[48] = oneWire /*8384*/;
  assign inv_25[49] = oneWire /*8378*/;
  assign inv_25[50] = oneWire /*8372*/;
  assign inv_25[51] = oneWire /*8366*/;
  assign inv_25[52] = oneWire /*8360*/;
  assign inv_25[53] = oneWire /*8354*/;
  assign inv_25[54] = oneWire /*8348*/;
  assign inv_25[55] = oneWire /*8342*/;
  assign inv_25[56] = oneWire /*8336*/;
  assign inv_25[57] = oneWire /*8330*/;
  assign inv_25[58] = oneWire /*8324*/;
  assign inv_25[59] = oneWire /*8318*/;
  assign inv_25[60] = oneWire /*8312*/;
  assign inv_25[61] = oneWire /*8306*/;
  assign inv_25[62] = oneWire /*8300*/;
  assign inv_25[63] = oneWire /*8294*/;
  assign inv_25[64] = oneWire /*8288*/;
  assign inv_25[65] = oneWire /*8282*/;
  assign inv_25[66] = oneWire /*8276*/;
  assign inv_25[67] = oneWire /*8270*/;
  assign inv_25[68] = oneWire /*8264*/;
  assign inv_25[69] = oneWire /*8258*/;
  assign inv_25[70] = oneWire /*8252*/;
  assign inv_25[71] = oneWire /*8246*/;
  assign inv_25[72] = oneWire /*8240*/;
  assign inv_25[73] = oneWire /*8234*/;
  assign inv_25[74] = oneWire /*8228*/;
  assign inv_25[75] = oneWire /*8222*/;
  assign inv_25[76] = oneWire /*8216*/;
  assign inv_25[77] = oneWire /*8210*/;
  assign inv_25[78] = oneWire /*8204*/;
  assign inv_25[79] = oneWire /*8198*/;
  assign inv_25[80] = oneWire /*8192*/;
  assign inv_25[81] = oneWire /*8186*/;
  assign inv_25[82] = oneWire /*8180*/;
  assign inv_25[83] = oneWire /*8174*/;
  assign inv_25[84] = oneWire /*8168*/;
  assign inv_25[85] = oneWire /*8162*/;
  assign inv_25[86] = oneWire /*8156*/;
  assign _12708_ = inv_25[0] ^ r_24[0] /*8671*/;
  assign sum_25[0] = _12708_ ^ oneWire /*8670*/;
  assign _12709_ = _12708_ & oneWire /*8669*/;
  assign _12710_ = inv_25[0] & r_24[0] /*8668*/;
  assign _12711_ = _12709_ | _12710_ /*8667*/;
  assign _12712_ = inv_25[1] ^ r_24[1] /*8665*/;
  assign sum_25[1] = _12712_ ^ _12711_ /*8664*/;
  assign _12713_ = _12712_ & _12711_ /*8663*/;
  assign _12714_ = inv_25[1] & r_24[1] /*8662*/;
  assign _12715_ = _12713_ | _12714_ /*8661*/;
  assign _12716_ = inv_25[2] ^ r_24[2] /*8659*/;
  assign sum_25[2] = _12716_ ^ _12715_ /*8658*/;
  assign _12717_ = _12716_ & _12715_ /*8657*/;
  assign _12718_ = inv_25[2] & r_24[2] /*8656*/;
  assign _12719_ = _12717_ | _12718_ /*8655*/;
  assign _12720_ = inv_25[3] ^ r_24[3] /*8653*/;
  assign sum_25[3] = _12720_ ^ _12719_ /*8652*/;
  assign _12721_ = _12720_ & _12719_ /*8651*/;
  assign _12722_ = inv_25[3] & r_24[3] /*8650*/;
  assign _12723_ = _12721_ | _12722_ /*8649*/;
  assign _12724_ = inv_25[4] ^ r_24[4] /*8647*/;
  assign sum_25[4] = _12724_ ^ _12723_ /*8646*/;
  assign _12725_ = _12724_ & _12723_ /*8645*/;
  assign _12726_ = inv_25[4] & r_24[4] /*8644*/;
  assign _12727_ = _12725_ | _12726_ /*8643*/;
  assign _12728_ = inv_25[5] ^ r_24[5] /*8641*/;
  assign sum_25[5] = _12728_ ^ _12727_ /*8640*/;
  assign _12729_ = _12728_ & _12727_ /*8639*/;
  assign _12730_ = inv_25[5] & r_24[5] /*8638*/;
  assign _12731_ = _12729_ | _12730_ /*8637*/;
  assign _12732_ = inv_25[6] ^ r_24[6] /*8635*/;
  assign sum_25[6] = _12732_ ^ _12731_ /*8634*/;
  assign _12733_ = _12732_ & _12731_ /*8633*/;
  assign _12734_ = inv_25[6] & r_24[6] /*8632*/;
  assign _12735_ = _12733_ | _12734_ /*8631*/;
  assign _12736_ = inv_25[7] ^ r_24[7] /*8629*/;
  assign sum_25[7] = _12736_ ^ _12735_ /*8628*/;
  assign _12737_ = _12736_ & _12735_ /*8627*/;
  assign _12738_ = inv_25[7] & r_24[7] /*8626*/;
  assign _12739_ = _12737_ | _12738_ /*8625*/;
  assign _12740_ = inv_25[8] ^ r_24[8] /*8623*/;
  assign sum_25[8] = _12740_ ^ _12739_ /*8622*/;
  assign _12741_ = _12740_ & _12739_ /*8621*/;
  assign _12742_ = inv_25[8] & r_24[8] /*8620*/;
  assign _12743_ = _12741_ | _12742_ /*8619*/;
  assign _12744_ = inv_25[9] ^ r_24[9] /*8617*/;
  assign sum_25[9] = _12744_ ^ _12743_ /*8616*/;
  assign _12745_ = _12744_ & _12743_ /*8615*/;
  assign _12746_ = inv_25[9] & r_24[9] /*8614*/;
  assign _12747_ = _12745_ | _12746_ /*8613*/;
  assign _12748_ = inv_25[10] ^ r_24[10] /*8611*/;
  assign sum_25[10] = _12748_ ^ _12747_ /*8610*/;
  assign _12749_ = _12748_ & _12747_ /*8609*/;
  assign _12750_ = inv_25[10] & r_24[10] /*8608*/;
  assign _12751_ = _12749_ | _12750_ /*8607*/;
  assign _12752_ = inv_25[11] ^ r_24[11] /*8605*/;
  assign sum_25[11] = _12752_ ^ _12751_ /*8604*/;
  assign _12753_ = _12752_ & _12751_ /*8603*/;
  assign _12754_ = inv_25[11] & r_24[11] /*8602*/;
  assign _12755_ = _12753_ | _12754_ /*8601*/;
  assign _12756_ = inv_25[12] ^ r_24[12] /*8599*/;
  assign sum_25[12] = _12756_ ^ _12755_ /*8598*/;
  assign _12757_ = _12756_ & _12755_ /*8597*/;
  assign _12758_ = inv_25[12] & r_24[12] /*8596*/;
  assign _12759_ = _12757_ | _12758_ /*8595*/;
  assign _12760_ = inv_25[13] ^ r_24[13] /*8593*/;
  assign sum_25[13] = _12760_ ^ _12759_ /*8592*/;
  assign _12761_ = _12760_ & _12759_ /*8591*/;
  assign _12762_ = inv_25[13] & r_24[13] /*8590*/;
  assign _12763_ = _12761_ | _12762_ /*8589*/;
  assign _12764_ = inv_25[14] ^ r_24[14] /*8587*/;
  assign sum_25[14] = _12764_ ^ _12763_ /*8586*/;
  assign _12765_ = _12764_ & _12763_ /*8585*/;
  assign _12766_ = inv_25[14] & r_24[14] /*8584*/;
  assign _12767_ = _12765_ | _12766_ /*8583*/;
  assign _12768_ = inv_25[15] ^ r_24[15] /*8581*/;
  assign sum_25[15] = _12768_ ^ _12767_ /*8580*/;
  assign _12769_ = _12768_ & _12767_ /*8579*/;
  assign _12770_ = inv_25[15] & r_24[15] /*8578*/;
  assign _12771_ = _12769_ | _12770_ /*8577*/;
  assign _12772_ = inv_25[16] ^ r_24[16] /*8575*/;
  assign sum_25[16] = _12772_ ^ _12771_ /*8574*/;
  assign _12773_ = _12772_ & _12771_ /*8573*/;
  assign _12774_ = inv_25[16] & r_24[16] /*8572*/;
  assign _12775_ = _12773_ | _12774_ /*8571*/;
  assign _12776_ = inv_25[17] ^ r_24[17] /*8569*/;
  assign sum_25[17] = _12776_ ^ _12775_ /*8568*/;
  assign _12777_ = _12776_ & _12775_ /*8567*/;
  assign _12778_ = inv_25[17] & r_24[17] /*8566*/;
  assign _12779_ = _12777_ | _12778_ /*8565*/;
  assign _12780_ = inv_25[18] ^ r_24[18] /*8563*/;
  assign sum_25[18] = _12780_ ^ _12779_ /*8562*/;
  assign _12781_ = _12780_ & _12779_ /*8561*/;
  assign _12782_ = inv_25[18] & r_24[18] /*8560*/;
  assign _12783_ = _12781_ | _12782_ /*8559*/;
  assign _12784_ = inv_25[19] ^ r_24[19] /*8557*/;
  assign sum_25[19] = _12784_ ^ _12783_ /*8556*/;
  assign _12785_ = _12784_ & _12783_ /*8555*/;
  assign _12786_ = inv_25[19] & r_24[19] /*8554*/;
  assign _12787_ = _12785_ | _12786_ /*8553*/;
  assign _12788_ = inv_25[20] ^ r_24[20] /*8551*/;
  assign sum_25[20] = _12788_ ^ _12787_ /*8550*/;
  assign _12789_ = _12788_ & _12787_ /*8549*/;
  assign _12790_ = inv_25[20] & r_24[20] /*8548*/;
  assign _12791_ = _12789_ | _12790_ /*8547*/;
  assign _12792_ = inv_25[21] ^ r_24[21] /*8545*/;
  assign sum_25[21] = _12792_ ^ _12791_ /*8544*/;
  assign _12793_ = _12792_ & _12791_ /*8543*/;
  assign _12794_ = inv_25[21] & r_24[21] /*8542*/;
  assign _12795_ = _12793_ | _12794_ /*8541*/;
  assign _12796_ = inv_25[22] ^ r_24[22] /*8539*/;
  assign sum_25[22] = _12796_ ^ _12795_ /*8538*/;
  assign _12797_ = _12796_ & _12795_ /*8537*/;
  assign _12798_ = inv_25[22] & r_24[22] /*8536*/;
  assign _12799_ = _12797_ | _12798_ /*8535*/;
  assign _12800_ = inv_25[23] ^ r_24[23] /*8533*/;
  assign sum_25[23] = _12800_ ^ _12799_ /*8532*/;
  assign _12801_ = _12800_ & _12799_ /*8531*/;
  assign _12802_ = inv_25[23] & r_24[23] /*8530*/;
  assign _12803_ = _12801_ | _12802_ /*8529*/;
  assign _12804_ = inv_25[24] ^ r_24[24] /*8527*/;
  assign sum_25[24] = _12804_ ^ _12803_ /*8526*/;
  assign _12805_ = _12804_ & _12803_ /*8525*/;
  assign _12806_ = inv_25[24] & r_24[24] /*8524*/;
  assign _12807_ = _12805_ | _12806_ /*8523*/;
  assign _12808_ = inv_25[25] ^ r_24[25] /*8521*/;
  assign sum_25[25] = _12808_ ^ _12807_ /*8520*/;
  assign _12809_ = _12808_ & _12807_ /*8519*/;
  assign _12810_ = inv_25[25] & r_24[25] /*8518*/;
  assign _12811_ = _12809_ | _12810_ /*8517*/;
  assign _12812_ = inv_25[26] ^ r_24[26] /*8515*/;
  assign sum_25[26] = _12812_ ^ _12811_ /*8514*/;
  assign _12813_ = _12812_ & _12811_ /*8513*/;
  assign _12814_ = inv_25[26] & r_24[26] /*8512*/;
  assign _12815_ = _12813_ | _12814_ /*8511*/;
  assign _12816_ = inv_25[27] ^ r_24[27] /*8509*/;
  assign sum_25[27] = _12816_ ^ _12815_ /*8508*/;
  assign _12817_ = _12816_ & _12815_ /*8507*/;
  assign _12818_ = inv_25[27] & r_24[27] /*8506*/;
  assign _12819_ = _12817_ | _12818_ /*8505*/;
  assign _12820_ = inv_25[28] ^ r_24[28] /*8503*/;
  assign sum_25[28] = _12820_ ^ _12819_ /*8502*/;
  assign _12821_ = _12820_ & _12819_ /*8501*/;
  assign _12822_ = inv_25[28] & r_24[28] /*8500*/;
  assign _12823_ = _12821_ | _12822_ /*8499*/;
  assign _12824_ = inv_25[29] ^ r_24[29] /*8497*/;
  assign sum_25[29] = _12824_ ^ _12823_ /*8496*/;
  assign _12825_ = _12824_ & _12823_ /*8495*/;
  assign _12826_ = inv_25[29] & r_24[29] /*8494*/;
  assign _12827_ = _12825_ | _12826_ /*8493*/;
  assign _12828_ = inv_25[30] ^ r_24[30] /*8491*/;
  assign sum_25[30] = _12828_ ^ _12827_ /*8490*/;
  assign _12829_ = _12828_ & _12827_ /*8489*/;
  assign _12830_ = inv_25[30] & r_24[30] /*8488*/;
  assign _12831_ = _12829_ | _12830_ /*8487*/;
  assign _12832_ = inv_25[31] ^ r_24[31] /*8485*/;
  assign sum_25[31] = _12832_ ^ _12831_ /*8484*/;
  assign _12833_ = _12832_ & _12831_ /*8483*/;
  assign _12834_ = inv_25[31] & r_24[31] /*8482*/;
  assign _12835_ = _12833_ | _12834_ /*8481*/;
  assign _12836_ = inv_25[32] ^ r_24[32] /*8479*/;
  assign sum_25[32] = _12836_ ^ _12835_ /*8478*/;
  assign _12837_ = _12836_ & _12835_ /*8477*/;
  assign _12838_ = inv_25[32] & r_24[32] /*8476*/;
  assign _12839_ = _12837_ | _12838_ /*8475*/;
  assign _12840_ = inv_25[33] ^ r_24[33] /*8473*/;
  assign sum_25[33] = _12840_ ^ _12839_ /*8472*/;
  assign _12841_ = _12840_ & _12839_ /*8471*/;
  assign _12842_ = inv_25[33] & r_24[33] /*8470*/;
  assign _12843_ = _12841_ | _12842_ /*8469*/;
  assign _12844_ = inv_25[34] ^ r_24[34] /*8467*/;
  assign sum_25[34] = _12844_ ^ _12843_ /*8466*/;
  assign _12845_ = _12844_ & _12843_ /*8465*/;
  assign _12846_ = inv_25[34] & r_24[34] /*8464*/;
  assign _12847_ = _12845_ | _12846_ /*8463*/;
  assign _12848_ = inv_25[35] ^ r_24[35] /*8461*/;
  assign sum_25[35] = _12848_ ^ _12847_ /*8460*/;
  assign _12849_ = _12848_ & _12847_ /*8459*/;
  assign _12850_ = inv_25[35] & r_24[35] /*8458*/;
  assign _12851_ = _12849_ | _12850_ /*8457*/;
  assign _12852_ = inv_25[36] ^ r_24[36] /*8455*/;
  assign sum_25[36] = _12852_ ^ _12851_ /*8454*/;
  assign _12853_ = _12852_ & _12851_ /*8453*/;
  assign _12854_ = inv_25[36] & r_24[36] /*8452*/;
  assign _12855_ = _12853_ | _12854_ /*8451*/;
  assign _12856_ = inv_25[37] ^ r_24[37] /*8449*/;
  assign sum_25[37] = _12856_ ^ _12855_ /*8448*/;
  assign _12857_ = _12856_ & _12855_ /*8447*/;
  assign _12858_ = inv_25[37] & r_24[37] /*8446*/;
  assign _12859_ = _12857_ | _12858_ /*8445*/;
  assign _12860_ = inv_25[38] ^ r_24[38] /*8443*/;
  assign sum_25[38] = _12860_ ^ _12859_ /*8442*/;
  assign _12861_ = _12860_ & _12859_ /*8441*/;
  assign _12862_ = inv_25[38] & r_24[38] /*8440*/;
  assign _12863_ = _12861_ | _12862_ /*8439*/;
  assign _12864_ = inv_25[39] ^ r_24[39] /*8437*/;
  assign sum_25[39] = _12864_ ^ _12863_ /*8436*/;
  assign _12865_ = _12864_ & _12863_ /*8435*/;
  assign _12866_ = inv_25[39] & r_24[39] /*8434*/;
  assign _12867_ = _12865_ | _12866_ /*8433*/;
  assign _12868_ = inv_25[40] ^ r_24[40] /*8431*/;
  assign sum_25[40] = _12868_ ^ _12867_ /*8430*/;
  assign _12869_ = _12868_ & _12867_ /*8429*/;
  assign _12870_ = inv_25[40] & r_24[40] /*8428*/;
  assign _12871_ = _12869_ | _12870_ /*8427*/;
  assign _12872_ = inv_25[41] ^ r_24[41] /*8425*/;
  assign sum_25[41] = _12872_ ^ _12871_ /*8424*/;
  assign _12873_ = _12872_ & _12871_ /*8423*/;
  assign _12874_ = inv_25[41] & r_24[41] /*8422*/;
  assign _12875_ = _12873_ | _12874_ /*8421*/;
  assign _12876_ = inv_25[42] ^ r_24[42] /*8419*/;
  assign sum_25[42] = _12876_ ^ _12875_ /*8418*/;
  assign _12877_ = _12876_ & _12875_ /*8417*/;
  assign _12878_ = inv_25[42] & r_24[42] /*8416*/;
  assign _12879_ = _12877_ | _12878_ /*8415*/;
  assign _12880_ = inv_25[43] ^ r_24[43] /*8413*/;
  assign sum_25[43] = _12880_ ^ _12879_ /*8412*/;
  assign _12881_ = _12880_ & _12879_ /*8411*/;
  assign _12882_ = inv_25[43] & r_24[43] /*8410*/;
  assign _12883_ = _12881_ | _12882_ /*8409*/;
  assign _12884_ = inv_25[44] ^ r_24[44] /*8407*/;
  assign sum_25[44] = _12884_ ^ _12883_ /*8406*/;
  assign _12885_ = _12884_ & _12883_ /*8405*/;
  assign _12886_ = inv_25[44] & r_24[44] /*8404*/;
  assign _12887_ = _12885_ | _12886_ /*8403*/;
  assign _12888_ = inv_25[45] ^ r_24[45] /*8401*/;
  assign sum_25[45] = _12888_ ^ _12887_ /*8400*/;
  assign _12889_ = _12888_ & _12887_ /*8399*/;
  assign _12890_ = inv_25[45] & r_24[45] /*8398*/;
  assign _12891_ = _12889_ | _12890_ /*8397*/;
  assign _12892_ = inv_25[46] ^ r_24[46] /*8395*/;
  assign sum_25[46] = _12892_ ^ _12891_ /*8394*/;
  assign _12893_ = _12892_ & _12891_ /*8393*/;
  assign _12894_ = inv_25[46] & r_24[46] /*8392*/;
  assign _12895_ = _12893_ | _12894_ /*8391*/;
  assign _12896_ = inv_25[47] ^ r_24[47] /*8389*/;
  assign sum_25[47] = _12896_ ^ _12895_ /*8388*/;
  assign _12897_ = _12896_ & _12895_ /*8387*/;
  assign _12898_ = inv_25[47] & r_24[47] /*8386*/;
  assign _12899_ = _12897_ | _12898_ /*8385*/;
  assign _12900_ = inv_25[48] ^ r_24[48] /*8383*/;
  assign sum_25[48] = _12900_ ^ _12899_ /*8382*/;
  assign _12901_ = _12900_ & _12899_ /*8381*/;
  assign _12902_ = inv_25[48] & r_24[48] /*8380*/;
  assign _12903_ = _12901_ | _12902_ /*8379*/;
  assign _12904_ = inv_25[49] ^ r_24[49] /*8377*/;
  assign sum_25[49] = _12904_ ^ _12903_ /*8376*/;
  assign _12905_ = _12904_ & _12903_ /*8375*/;
  assign _12906_ = inv_25[49] & r_24[49] /*8374*/;
  assign _12907_ = _12905_ | _12906_ /*8373*/;
  assign _12908_ = inv_25[50] ^ r_24[50] /*8371*/;
  assign sum_25[50] = _12908_ ^ _12907_ /*8370*/;
  assign _12909_ = _12908_ & _12907_ /*8369*/;
  assign _12910_ = inv_25[50] & r_24[50] /*8368*/;
  assign _12911_ = _12909_ | _12910_ /*8367*/;
  assign _12912_ = inv_25[51] ^ r_24[51] /*8365*/;
  assign sum_25[51] = _12912_ ^ _12911_ /*8364*/;
  assign _12913_ = _12912_ & _12911_ /*8363*/;
  assign _12914_ = inv_25[51] & r_24[51] /*8362*/;
  assign _12915_ = _12913_ | _12914_ /*8361*/;
  assign _12916_ = inv_25[52] ^ r_24[52] /*8359*/;
  assign sum_25[52] = _12916_ ^ _12915_ /*8358*/;
  assign _12917_ = _12916_ & _12915_ /*8357*/;
  assign _12918_ = inv_25[52] & r_24[52] /*8356*/;
  assign _12919_ = _12917_ | _12918_ /*8355*/;
  assign _12920_ = inv_25[53] ^ r_24[53] /*8353*/;
  assign sum_25[53] = _12920_ ^ _12919_ /*8352*/;
  assign _12921_ = _12920_ & _12919_ /*8351*/;
  assign _12922_ = inv_25[53] & r_24[53] /*8350*/;
  assign _12923_ = _12921_ | _12922_ /*8349*/;
  assign _12924_ = inv_25[54] ^ r_24[54] /*8347*/;
  assign sum_25[54] = _12924_ ^ _12923_ /*8346*/;
  assign _12925_ = _12924_ & _12923_ /*8345*/;
  assign _12926_ = inv_25[54] & r_24[54] /*8344*/;
  assign _12927_ = _12925_ | _12926_ /*8343*/;
  assign _12928_ = inv_25[55] ^ r_24[55] /*8341*/;
  assign sum_25[55] = _12928_ ^ _12927_ /*8340*/;
  assign _12929_ = _12928_ & _12927_ /*8339*/;
  assign _12930_ = inv_25[55] & r_24[55] /*8338*/;
  assign _12931_ = _12929_ | _12930_ /*8337*/;
  assign _12932_ = inv_25[56] ^ r_24[56] /*8335*/;
  assign sum_25[56] = _12932_ ^ _12931_ /*8334*/;
  assign _12933_ = _12932_ & _12931_ /*8333*/;
  assign _12934_ = inv_25[56] & r_24[56] /*8332*/;
  assign _12935_ = _12933_ | _12934_ /*8331*/;
  assign _12936_ = inv_25[57] ^ r_24[57] /*8329*/;
  assign sum_25[57] = _12936_ ^ _12935_ /*8328*/;
  assign _12937_ = _12936_ & _12935_ /*8327*/;
  assign _12938_ = inv_25[57] & r_24[57] /*8326*/;
  assign _12939_ = _12937_ | _12938_ /*8325*/;
  assign _12940_ = inv_25[58] ^ r_24[58] /*8323*/;
  assign sum_25[58] = _12940_ ^ _12939_ /*8322*/;
  assign _12941_ = _12940_ & _12939_ /*8321*/;
  assign _12942_ = inv_25[58] & r_24[58] /*8320*/;
  assign _12943_ = _12941_ | _12942_ /*8319*/;
  assign _12944_ = inv_25[59] ^ r_24[59] /*8317*/;
  assign sum_25[59] = _12944_ ^ _12943_ /*8316*/;
  assign _12945_ = _12944_ & _12943_ /*8315*/;
  assign _12946_ = inv_25[59] & r_24[59] /*8314*/;
  assign _12947_ = _12945_ | _12946_ /*8313*/;
  assign _12948_ = inv_25[60] ^ r_24[60] /*8311*/;
  assign sum_25[60] = _12948_ ^ _12947_ /*8310*/;
  assign _12949_ = _12948_ & _12947_ /*8309*/;
  assign _12950_ = inv_25[60] & r_24[60] /*8308*/;
  assign _12951_ = _12949_ | _12950_ /*8307*/;
  assign _12952_ = inv_25[61] ^ r_24[61] /*8305*/;
  assign sum_25[61] = _12952_ ^ _12951_ /*8304*/;
  assign _12953_ = _12952_ & _12951_ /*8303*/;
  assign _12954_ = inv_25[61] & r_24[61] /*8302*/;
  assign _12955_ = _12953_ | _12954_ /*8301*/;
  assign _12956_ = inv_25[62] ^ r_24[62] /*8299*/;
  assign sum_25[62] = _12956_ ^ _12955_ /*8298*/;
  assign _12957_ = _12956_ & _12955_ /*8297*/;
  assign _12958_ = inv_25[62] & r_24[62] /*8296*/;
  assign _12959_ = _12957_ | _12958_ /*8295*/;
  assign _12960_ = inv_25[63] ^ r_24[63] /*8293*/;
  assign sum_25[63] = _12960_ ^ _12959_ /*8292*/;
  assign _12961_ = _12960_ & _12959_ /*8291*/;
  assign _12962_ = inv_25[63] & r_24[63] /*8290*/;
  assign _12963_ = _12961_ | _12962_ /*8289*/;
  assign _12964_ = inv_25[64] ^ r_24[64] /*8287*/;
  assign sum_25[64] = _12964_ ^ _12963_ /*8286*/;
  assign _12965_ = _12964_ & _12963_ /*8285*/;
  assign _12966_ = inv_25[64] & r_24[64] /*8284*/;
  assign _12967_ = _12965_ | _12966_ /*8283*/;
  assign _12968_ = inv_25[65] ^ r_24[65] /*8281*/;
  assign sum_25[65] = _12968_ ^ _12967_ /*8280*/;
  assign _12969_ = _12968_ & _12967_ /*8279*/;
  assign _12970_ = inv_25[65] & r_24[65] /*8278*/;
  assign _12971_ = _12969_ | _12970_ /*8277*/;
  assign _12972_ = inv_25[66] ^ r_24[66] /*8275*/;
  assign sum_25[66] = _12972_ ^ _12971_ /*8274*/;
  assign _12973_ = _12972_ & _12971_ /*8273*/;
  assign _12974_ = inv_25[66] & r_24[66] /*8272*/;
  assign _12975_ = _12973_ | _12974_ /*8271*/;
  assign _12976_ = inv_25[67] ^ r_24[67] /*8269*/;
  assign sum_25[67] = _12976_ ^ _12975_ /*8268*/;
  assign _12977_ = _12976_ & _12975_ /*8267*/;
  assign _12978_ = inv_25[67] & r_24[67] /*8266*/;
  assign _12979_ = _12977_ | _12978_ /*8265*/;
  assign _12980_ = inv_25[68] ^ r_24[68] /*8263*/;
  assign sum_25[68] = _12980_ ^ _12979_ /*8262*/;
  assign _12981_ = _12980_ & _12979_ /*8261*/;
  assign _12982_ = inv_25[68] & r_24[68] /*8260*/;
  assign _12983_ = _12981_ | _12982_ /*8259*/;
  assign _12984_ = inv_25[69] ^ r_24[69] /*8257*/;
  assign sum_25[69] = _12984_ ^ _12983_ /*8256*/;
  assign _12985_ = _12984_ & _12983_ /*8255*/;
  assign _12986_ = inv_25[69] & r_24[69] /*8254*/;
  assign _12987_ = _12985_ | _12986_ /*8253*/;
  assign _12988_ = inv_25[70] ^ r_24[70] /*8251*/;
  assign sum_25[70] = _12988_ ^ _12987_ /*8250*/;
  assign _12989_ = _12988_ & _12987_ /*8249*/;
  assign _12990_ = inv_25[70] & r_24[70] /*8248*/;
  assign _12991_ = _12989_ | _12990_ /*8247*/;
  assign _12992_ = inv_25[71] ^ r_24[71] /*8245*/;
  assign sum_25[71] = _12992_ ^ _12991_ /*8244*/;
  assign _12993_ = _12992_ & _12991_ /*8243*/;
  assign _12994_ = inv_25[71] & r_24[71] /*8242*/;
  assign _12995_ = _12993_ | _12994_ /*8241*/;
  assign _12996_ = inv_25[72] ^ r_24[72] /*8239*/;
  assign sum_25[72] = _12996_ ^ _12995_ /*8238*/;
  assign _12997_ = _12996_ & _12995_ /*8237*/;
  assign _12998_ = inv_25[72] & r_24[72] /*8236*/;
  assign _12999_ = _12997_ | _12998_ /*8235*/;
  assign _13000_ = inv_25[73] ^ r_24[73] /*8233*/;
  assign sum_25[73] = _13000_ ^ _12999_ /*8232*/;
  assign _13001_ = _13000_ & _12999_ /*8231*/;
  assign _13002_ = inv_25[73] & r_24[73] /*8230*/;
  assign _13003_ = _13001_ | _13002_ /*8229*/;
  assign _13004_ = inv_25[74] ^ r_24[74] /*8227*/;
  assign sum_25[74] = _13004_ ^ _13003_ /*8226*/;
  assign _13005_ = _13004_ & _13003_ /*8225*/;
  assign _13006_ = inv_25[74] & r_24[74] /*8224*/;
  assign _13007_ = _13005_ | _13006_ /*8223*/;
  assign _13008_ = inv_25[75] ^ r_24[75] /*8221*/;
  assign sum_25[75] = _13008_ ^ _13007_ /*8220*/;
  assign _13009_ = _13008_ & _13007_ /*8219*/;
  assign _13010_ = inv_25[75] & r_24[75] /*8218*/;
  assign _13011_ = _13009_ | _13010_ /*8217*/;
  assign _13012_ = inv_25[76] ^ r_24[76] /*8215*/;
  assign sum_25[76] = _13012_ ^ _13011_ /*8214*/;
  assign _13013_ = _13012_ & _13011_ /*8213*/;
  assign _13014_ = inv_25[76] & r_24[76] /*8212*/;
  assign _13015_ = _13013_ | _13014_ /*8211*/;
  assign _13016_ = inv_25[77] ^ r_24[77] /*8209*/;
  assign sum_25[77] = _13016_ ^ _13015_ /*8208*/;
  assign _13017_ = _13016_ & _13015_ /*8207*/;
  assign _13018_ = inv_25[77] & r_24[77] /*8206*/;
  assign _13019_ = _13017_ | _13018_ /*8205*/;
  assign _13020_ = inv_25[78] ^ r_24[78] /*8203*/;
  assign sum_25[78] = _13020_ ^ _13019_ /*8202*/;
  assign _13021_ = _13020_ & _13019_ /*8201*/;
  assign _13022_ = inv_25[78] & r_24[78] /*8200*/;
  assign _13023_ = _13021_ | _13022_ /*8199*/;
  assign _13024_ = inv_25[79] ^ r_24[79] /*8197*/;
  assign sum_25[79] = _13024_ ^ _13023_ /*8196*/;
  assign _13025_ = _13024_ & _13023_ /*8195*/;
  assign _13026_ = inv_25[79] & r_24[79] /*8194*/;
  assign _13027_ = _13025_ | _13026_ /*8193*/;
  assign _13028_ = inv_25[80] ^ r_24[80] /*8191*/;
  assign sum_25[80] = _13028_ ^ _13027_ /*8190*/;
  assign _13029_ = _13028_ & _13027_ /*8189*/;
  assign _13030_ = inv_25[80] & r_24[80] /*8188*/;
  assign _13031_ = _13029_ | _13030_ /*8187*/;
  assign _13032_ = inv_25[81] ^ r_24[81] /*8185*/;
  assign sum_25[81] = _13032_ ^ _13031_ /*8184*/;
  assign _13033_ = _13032_ & _13031_ /*8183*/;
  assign _13034_ = inv_25[81] & r_24[81] /*8182*/;
  assign _13035_ = _13033_ | _13034_ /*8181*/;
  assign _13036_ = inv_25[82] ^ r_24[82] /*8179*/;
  assign sum_25[82] = _13036_ ^ _13035_ /*8178*/;
  assign _13037_ = _13036_ & _13035_ /*8177*/;
  assign _13038_ = inv_25[82] & r_24[82] /*8176*/;
  assign _13039_ = _13037_ | _13038_ /*8175*/;
  assign _13040_ = inv_25[83] ^ r_24[83] /*8173*/;
  assign sum_25[83] = _13040_ ^ _13039_ /*8172*/;
  assign _13041_ = _13040_ & _13039_ /*8171*/;
  assign _13042_ = inv_25[83] & r_24[83] /*8170*/;
  assign _13043_ = _13041_ | _13042_ /*8169*/;
  assign _13044_ = inv_25[84] ^ r_24[84] /*8167*/;
  assign sum_25[84] = _13044_ ^ _13043_ /*8166*/;
  assign _13045_ = _13044_ & _13043_ /*8165*/;
  assign _13046_ = inv_25[84] & r_24[84] /*8164*/;
  assign _13047_ = _13045_ | _13046_ /*8163*/;
  assign _13048_ = inv_25[85] ^ r_24[85] /*8161*/;
  assign sum_25[85] = _13048_ ^ _13047_ /*8160*/;
  assign _13049_ = _13048_ & _13047_ /*8159*/;
  assign _13050_ = inv_25[85] & r_24[85] /*8158*/;
  assign _13051_ = _13049_ | _13050_ /*8157*/;
  assign _13052_ = inv_25[86] ^ r_24[86] /*8155*/;
  assign sum_25[86] = _13052_ ^ _13051_ /*8154*/;
  assign _13053_ = _13052_ & _13051_ /*8153*/;
  assign _13054_ = inv_25[86] & r_24[86] /*8152*/;
  assign _13055_ = _13053_ | _13054_ /*8151*/;
  assign _13056_ = _13055_ ^ _13051_ /*8150*/;
  assign _13057_ = ~_13056_ /*8149*/;
  assign _13058_ = sum_25[86] & _13057_ /*8148*/;
  assign _13059_ = _13056_ & _13055_ /*8147*/;
  assign sum_25[87] = _13059_ | _13058_ /*8146*/;
  assign q[7] = ~sum_25[87] /*8145*/;
  assign m_25[0] = r_24[0] /*8144*/;
  assign m_25[1] = r_24[1] /*8143*/;
  assign m_25[2] = r_24[2] /*8142*/;
  assign m_25[3] = r_24[3] /*8141*/;
  assign m_25[4] = r_24[4] /*8140*/;
  assign m_25[5] = r_24[5] /*8139*/;
  assign m_25[6] = r_24[6] /*8138*/;
  assign m_25[7] = r_24[7] /*8137*/;
  assign m_25[8] = r_24[8] /*8136*/;
  assign m_25[9] = r_24[9] /*8135*/;
  assign m_25[10] = r_24[10] /*8134*/;
  assign m_25[11] = r_24[11] /*8133*/;
  assign m_25[12] = r_24[12] /*8132*/;
  assign m_25[13] = r_24[13] /*8131*/;
  assign m_25[14] = r_24[14] /*8130*/;
  assign m_25[15] = r_24[15] /*8129*/;
  assign m_25[16] = r_24[16] /*8128*/;
  assign m_25[17] = r_24[17] /*8127*/;
  assign m_25[18] = r_24[18] /*8126*/;
  assign m_25[19] = r_24[19] /*8125*/;
  assign m_25[20] = r_24[20] /*8124*/;
  assign m_25[21] = r_24[21] /*8123*/;
  assign m_25[22] = r_24[22] /*8122*/;
  assign m_25[23] = r_24[23] /*8121*/;
  assign m_25[24] = r_24[24] /*8120*/;
  assign m_25[25] = r_24[25] /*8119*/;
  assign m_25[26] = r_24[26] /*8118*/;
  assign m_25[27] = r_24[27] /*8117*/;
  assign m_25[28] = r_24[28] /*8116*/;
  assign m_25[29] = r_24[29] /*8115*/;
  assign m_25[30] = r_24[30] /*8114*/;
  assign m_25[31] = r_24[31] /*8113*/;
  assign m_25[32] = r_24[32] /*8112*/;
  assign m_25[33] = r_24[33] /*8111*/;
  assign m_25[34] = r_24[34] /*8110*/;
  assign m_25[35] = r_24[35] /*8109*/;
  assign m_25[36] = r_24[36] /*8108*/;
  assign m_25[37] = r_24[37] /*8107*/;
  assign m_25[38] = r_24[38] /*8106*/;
  assign m_25[39] = r_24[39] /*8105*/;
  assign m_25[40] = r_24[40] /*8104*/;
  assign m_25[41] = r_24[41] /*8103*/;
  assign m_25[42] = r_24[42] /*8102*/;
  assign m_25[43] = r_24[43] /*8101*/;
  assign m_25[44] = r_24[44] /*8100*/;
  assign m_25[45] = r_24[45] /*8099*/;
  assign m_25[46] = r_24[46] /*8098*/;
  assign m_25[47] = r_24[47] /*8097*/;
  assign m_25[48] = r_24[48] /*8096*/;
  assign m_25[49] = r_24[49] /*8095*/;
  assign m_25[50] = r_24[50] /*8094*/;
  assign m_25[51] = r_24[51] /*8093*/;
  assign m_25[52] = r_24[52] /*8092*/;
  assign m_25[53] = r_24[53] /*8091*/;
  assign m_25[54] = r_24[54] /*8090*/;
  assign m_25[55] = r_24[55] /*8089*/;
  assign m_25[56] = r_24[56] /*8088*/;
  assign m_25[57] = r_24[57] /*8087*/;
  assign m_25[58] = r_24[58] /*8086*/;
  assign m_25[59] = r_24[59] /*8085*/;
  assign m_25[60] = r_24[60] /*8084*/;
  assign m_25[61] = r_24[61] /*8083*/;
  assign m_25[62] = r_24[62] /*8082*/;
  assign m_25[63] = r_24[63] /*8081*/;
  assign m_25[64] = r_24[64] /*8080*/;
  assign m_25[65] = r_24[65] /*8079*/;
  assign m_25[66] = r_24[66] /*8078*/;
  assign m_25[67] = r_24[67] /*8077*/;
  assign m_25[68] = r_24[68] /*8076*/;
  assign m_25[69] = r_24[69] /*8075*/;
  assign m_25[70] = r_24[70] /*8074*/;
  assign m_25[71] = r_24[71] /*8073*/;
  assign m_25[72] = r_24[72] /*8072*/;
  assign m_25[73] = r_24[73] /*8071*/;
  assign m_25[74] = r_24[74] /*8070*/;
  assign m_25[75] = r_24[75] /*8069*/;
  assign m_25[76] = r_24[76] /*8068*/;
  assign m_25[77] = r_24[77] /*8067*/;
  assign m_25[78] = r_24[78] /*8066*/;
  assign m_25[79] = r_24[79] /*8065*/;
  assign m_25[80] = r_24[80] /*8064*/;
  assign m_25[81] = r_24[81] /*8063*/;
  assign m_25[82] = r_24[82] /*8062*/;
  assign m_25[83] = r_24[83] /*8061*/;
  assign m_25[84] = r_24[84] /*8060*/;
  assign m_25[85] = r_24[85] /*8059*/;
  assign m_25[86] = r_24[86] /*8058*/;
  assign m_25[87] = r_24[86] /*8057*/;
  assign _13061_ = ~q[7] /*8056*/;
  assign _13062_ = sum_25[0] & q[7] /*8055*/;
  assign _13063_ = m_25[0] & _13061_ /*8054*/;
  assign r_25[0] = _13063_ | _13062_ /*8053*/;
  assign _13064_ = ~q[7] /*8052*/;
  assign _13065_ = sum_25[1] & q[7] /*8051*/;
  assign _13066_ = m_25[1] & _13064_ /*8050*/;
  assign r_25[1] = _13066_ | _13065_ /*8049*/;
  assign _13067_ = ~q[7] /*8048*/;
  assign _13068_ = sum_25[2] & q[7] /*8047*/;
  assign _13069_ = m_25[2] & _13067_ /*8046*/;
  assign r_25[2] = _13069_ | _13068_ /*8045*/;
  assign _13070_ = ~q[7] /*8044*/;
  assign _13071_ = sum_25[3] & q[7] /*8043*/;
  assign _13072_ = m_25[3] & _13070_ /*8042*/;
  assign r_25[3] = _13072_ | _13071_ /*8041*/;
  assign _13073_ = ~q[7] /*8040*/;
  assign _13074_ = sum_25[4] & q[7] /*8039*/;
  assign _13075_ = m_25[4] & _13073_ /*8038*/;
  assign r_25[4] = _13075_ | _13074_ /*8037*/;
  assign _13076_ = ~q[7] /*8036*/;
  assign _13077_ = sum_25[5] & q[7] /*8035*/;
  assign _13078_ = m_25[5] & _13076_ /*8034*/;
  assign r_25[5] = _13078_ | _13077_ /*8033*/;
  assign _13079_ = ~q[7] /*8032*/;
  assign _13080_ = sum_25[6] & q[7] /*8031*/;
  assign _13081_ = m_25[6] & _13079_ /*8030*/;
  assign r_25[6] = _13081_ | _13080_ /*8029*/;
  assign _13082_ = ~q[7] /*8028*/;
  assign _13083_ = sum_25[7] & q[7] /*8027*/;
  assign _13084_ = m_25[7] & _13082_ /*8026*/;
  assign r_25[7] = _13084_ | _13083_ /*8025*/;
  assign _13085_ = ~q[7] /*8024*/;
  assign _13086_ = sum_25[8] & q[7] /*8023*/;
  assign _13087_ = m_25[8] & _13085_ /*8022*/;
  assign r_25[8] = _13087_ | _13086_ /*8021*/;
  assign _13088_ = ~q[7] /*8020*/;
  assign _13089_ = sum_25[9] & q[7] /*8019*/;
  assign _13090_ = m_25[9] & _13088_ /*8018*/;
  assign r_25[9] = _13090_ | _13089_ /*8017*/;
  assign _13091_ = ~q[7] /*8016*/;
  assign _13092_ = sum_25[10] & q[7] /*8015*/;
  assign _13093_ = m_25[10] & _13091_ /*8014*/;
  assign r_25[10] = _13093_ | _13092_ /*8013*/;
  assign _13094_ = ~q[7] /*8012*/;
  assign _13095_ = sum_25[11] & q[7] /*8011*/;
  assign _13096_ = m_25[11] & _13094_ /*8010*/;
  assign r_25[11] = _13096_ | _13095_ /*8009*/;
  assign _13097_ = ~q[7] /*8008*/;
  assign _13098_ = sum_25[12] & q[7] /*8007*/;
  assign _13099_ = m_25[12] & _13097_ /*8006*/;
  assign r_25[12] = _13099_ | _13098_ /*8005*/;
  assign _13100_ = ~q[7] /*8004*/;
  assign _13101_ = sum_25[13] & q[7] /*8003*/;
  assign _13102_ = m_25[13] & _13100_ /*8002*/;
  assign r_25[13] = _13102_ | _13101_ /*8001*/;
  assign _13103_ = ~q[7] /*8000*/;
  assign _13104_ = sum_25[14] & q[7] /*7999*/;
  assign _13105_ = m_25[14] & _13103_ /*7998*/;
  assign r_25[14] = _13105_ | _13104_ /*7997*/;
  assign _13106_ = ~q[7] /*7996*/;
  assign _13107_ = sum_25[15] & q[7] /*7995*/;
  assign _13108_ = m_25[15] & _13106_ /*7994*/;
  assign r_25[15] = _13108_ | _13107_ /*7993*/;
  assign _13109_ = ~q[7] /*7992*/;
  assign _13110_ = sum_25[16] & q[7] /*7991*/;
  assign _13111_ = m_25[16] & _13109_ /*7990*/;
  assign r_25[16] = _13111_ | _13110_ /*7989*/;
  assign _13112_ = ~q[7] /*7988*/;
  assign _13113_ = sum_25[17] & q[7] /*7987*/;
  assign _13114_ = m_25[17] & _13112_ /*7986*/;
  assign r_25[17] = _13114_ | _13113_ /*7985*/;
  assign _13115_ = ~q[7] /*7984*/;
  assign _13116_ = sum_25[18] & q[7] /*7983*/;
  assign _13117_ = m_25[18] & _13115_ /*7982*/;
  assign r_25[18] = _13117_ | _13116_ /*7981*/;
  assign _13118_ = ~q[7] /*7980*/;
  assign _13119_ = sum_25[19] & q[7] /*7979*/;
  assign _13120_ = m_25[19] & _13118_ /*7978*/;
  assign r_25[19] = _13120_ | _13119_ /*7977*/;
  assign _13121_ = ~q[7] /*7976*/;
  assign _13122_ = sum_25[20] & q[7] /*7975*/;
  assign _13123_ = m_25[20] & _13121_ /*7974*/;
  assign r_25[20] = _13123_ | _13122_ /*7973*/;
  assign _13124_ = ~q[7] /*7972*/;
  assign _13125_ = sum_25[21] & q[7] /*7971*/;
  assign _13126_ = m_25[21] & _13124_ /*7970*/;
  assign r_25[21] = _13126_ | _13125_ /*7969*/;
  assign _13127_ = ~q[7] /*7968*/;
  assign _13128_ = sum_25[22] & q[7] /*7967*/;
  assign _13129_ = m_25[22] & _13127_ /*7966*/;
  assign r_25[22] = _13129_ | _13128_ /*7965*/;
  assign _13130_ = ~q[7] /*7964*/;
  assign _13131_ = sum_25[23] & q[7] /*7963*/;
  assign _13132_ = m_25[23] & _13130_ /*7962*/;
  assign r_25[23] = _13132_ | _13131_ /*7961*/;
  assign _13133_ = ~q[7] /*7960*/;
  assign _13134_ = sum_25[24] & q[7] /*7959*/;
  assign _13135_ = m_25[24] & _13133_ /*7958*/;
  assign r_25[24] = _13135_ | _13134_ /*7957*/;
  assign _13136_ = ~q[7] /*7956*/;
  assign _13137_ = sum_25[25] & q[7] /*7955*/;
  assign _13138_ = m_25[25] & _13136_ /*7954*/;
  assign r_25[25] = _13138_ | _13137_ /*7953*/;
  assign _13139_ = ~q[7] /*7952*/;
  assign _13140_ = sum_25[26] & q[7] /*7951*/;
  assign _13141_ = m_25[26] & _13139_ /*7950*/;
  assign r_25[26] = _13141_ | _13140_ /*7949*/;
  assign _13142_ = ~q[7] /*7948*/;
  assign _13143_ = sum_25[27] & q[7] /*7947*/;
  assign _13144_ = m_25[27] & _13142_ /*7946*/;
  assign r_25[27] = _13144_ | _13143_ /*7945*/;
  assign _13145_ = ~q[7] /*7944*/;
  assign _13146_ = sum_25[28] & q[7] /*7943*/;
  assign _13147_ = m_25[28] & _13145_ /*7942*/;
  assign r_25[28] = _13147_ | _13146_ /*7941*/;
  assign _13148_ = ~q[7] /*7940*/;
  assign _13149_ = sum_25[29] & q[7] /*7939*/;
  assign _13150_ = m_25[29] & _13148_ /*7938*/;
  assign r_25[29] = _13150_ | _13149_ /*7937*/;
  assign _13151_ = ~q[7] /*7936*/;
  assign _13152_ = sum_25[30] & q[7] /*7935*/;
  assign _13153_ = m_25[30] & _13151_ /*7934*/;
  assign r_25[30] = _13153_ | _13152_ /*7933*/;
  assign _13154_ = ~q[7] /*7932*/;
  assign _13155_ = sum_25[31] & q[7] /*7931*/;
  assign _13156_ = m_25[31] & _13154_ /*7930*/;
  assign r_25[31] = _13156_ | _13155_ /*7929*/;
  assign _13157_ = ~q[7] /*7928*/;
  assign _13158_ = sum_25[32] & q[7] /*7927*/;
  assign _13159_ = m_25[32] & _13157_ /*7926*/;
  assign r_25[32] = _13159_ | _13158_ /*7925*/;
  assign _13160_ = ~q[7] /*7924*/;
  assign _13161_ = sum_25[33] & q[7] /*7923*/;
  assign _13162_ = m_25[33] & _13160_ /*7922*/;
  assign r_25[33] = _13162_ | _13161_ /*7921*/;
  assign _13163_ = ~q[7] /*7920*/;
  assign _13164_ = sum_25[34] & q[7] /*7919*/;
  assign _13165_ = m_25[34] & _13163_ /*7918*/;
  assign r_25[34] = _13165_ | _13164_ /*7917*/;
  assign _13166_ = ~q[7] /*7916*/;
  assign _13167_ = sum_25[35] & q[7] /*7915*/;
  assign _13168_ = m_25[35] & _13166_ /*7914*/;
  assign r_25[35] = _13168_ | _13167_ /*7913*/;
  assign _13169_ = ~q[7] /*7912*/;
  assign _13170_ = sum_25[36] & q[7] /*7911*/;
  assign _13171_ = m_25[36] & _13169_ /*7910*/;
  assign r_25[36] = _13171_ | _13170_ /*7909*/;
  assign _13172_ = ~q[7] /*7908*/;
  assign _13173_ = sum_25[37] & q[7] /*7907*/;
  assign _13174_ = m_25[37] & _13172_ /*7906*/;
  assign r_25[37] = _13174_ | _13173_ /*7905*/;
  assign _13175_ = ~q[7] /*7904*/;
  assign _13176_ = sum_25[38] & q[7] /*7903*/;
  assign _13177_ = m_25[38] & _13175_ /*7902*/;
  assign r_25[38] = _13177_ | _13176_ /*7901*/;
  assign _13178_ = ~q[7] /*7900*/;
  assign _13179_ = sum_25[39] & q[7] /*7899*/;
  assign _13180_ = m_25[39] & _13178_ /*7898*/;
  assign r_25[39] = _13180_ | _13179_ /*7897*/;
  assign _13181_ = ~q[7] /*7896*/;
  assign _13182_ = sum_25[40] & q[7] /*7895*/;
  assign _13183_ = m_25[40] & _13181_ /*7894*/;
  assign r_25[40] = _13183_ | _13182_ /*7893*/;
  assign _13184_ = ~q[7] /*7892*/;
  assign _13185_ = sum_25[41] & q[7] /*7891*/;
  assign _13186_ = m_25[41] & _13184_ /*7890*/;
  assign r_25[41] = _13186_ | _13185_ /*7889*/;
  assign _13187_ = ~q[7] /*7888*/;
  assign _13188_ = sum_25[42] & q[7] /*7887*/;
  assign _13189_ = m_25[42] & _13187_ /*7886*/;
  assign r_25[42] = _13189_ | _13188_ /*7885*/;
  assign _13190_ = ~q[7] /*7884*/;
  assign _13191_ = sum_25[43] & q[7] /*7883*/;
  assign _13192_ = m_25[43] & _13190_ /*7882*/;
  assign r_25[43] = _13192_ | _13191_ /*7881*/;
  assign _13193_ = ~q[7] /*7880*/;
  assign _13194_ = sum_25[44] & q[7] /*7879*/;
  assign _13195_ = m_25[44] & _13193_ /*7878*/;
  assign r_25[44] = _13195_ | _13194_ /*7877*/;
  assign _13196_ = ~q[7] /*7876*/;
  assign _13197_ = sum_25[45] & q[7] /*7875*/;
  assign _13198_ = m_25[45] & _13196_ /*7874*/;
  assign r_25[45] = _13198_ | _13197_ /*7873*/;
  assign _13199_ = ~q[7] /*7872*/;
  assign _13200_ = sum_25[46] & q[7] /*7871*/;
  assign _13201_ = m_25[46] & _13199_ /*7870*/;
  assign r_25[46] = _13201_ | _13200_ /*7869*/;
  assign _13202_ = ~q[7] /*7868*/;
  assign _13203_ = sum_25[47] & q[7] /*7867*/;
  assign _13204_ = m_25[47] & _13202_ /*7866*/;
  assign r_25[47] = _13204_ | _13203_ /*7865*/;
  assign _13205_ = ~q[7] /*7864*/;
  assign _13206_ = sum_25[48] & q[7] /*7863*/;
  assign _13207_ = m_25[48] & _13205_ /*7862*/;
  assign r_25[48] = _13207_ | _13206_ /*7861*/;
  assign _13208_ = ~q[7] /*7860*/;
  assign _13209_ = sum_25[49] & q[7] /*7859*/;
  assign _13210_ = m_25[49] & _13208_ /*7858*/;
  assign r_25[49] = _13210_ | _13209_ /*7857*/;
  assign _13211_ = ~q[7] /*7856*/;
  assign _13212_ = sum_25[50] & q[7] /*7855*/;
  assign _13213_ = m_25[50] & _13211_ /*7854*/;
  assign r_25[50] = _13213_ | _13212_ /*7853*/;
  assign _13214_ = ~q[7] /*7852*/;
  assign _13215_ = sum_25[51] & q[7] /*7851*/;
  assign _13216_ = m_25[51] & _13214_ /*7850*/;
  assign r_25[51] = _13216_ | _13215_ /*7849*/;
  assign _13217_ = ~q[7] /*7848*/;
  assign _13218_ = sum_25[52] & q[7] /*7847*/;
  assign _13219_ = m_25[52] & _13217_ /*7846*/;
  assign r_25[52] = _13219_ | _13218_ /*7845*/;
  assign _13220_ = ~q[7] /*7844*/;
  assign _13221_ = sum_25[53] & q[7] /*7843*/;
  assign _13222_ = m_25[53] & _13220_ /*7842*/;
  assign r_25[53] = _13222_ | _13221_ /*7841*/;
  assign _13223_ = ~q[7] /*7840*/;
  assign _13224_ = sum_25[54] & q[7] /*7839*/;
  assign _13225_ = m_25[54] & _13223_ /*7838*/;
  assign r_25[54] = _13225_ | _13224_ /*7837*/;
  assign _13226_ = ~q[7] /*7836*/;
  assign _13227_ = sum_25[55] & q[7] /*7835*/;
  assign _13228_ = m_25[55] & _13226_ /*7834*/;
  assign r_25[55] = _13228_ | _13227_ /*7833*/;
  assign _13229_ = ~q[7] /*7832*/;
  assign _13230_ = sum_25[56] & q[7] /*7831*/;
  assign _13231_ = m_25[56] & _13229_ /*7830*/;
  assign r_25[56] = _13231_ | _13230_ /*7829*/;
  assign _13232_ = ~q[7] /*7828*/;
  assign _13233_ = sum_25[57] & q[7] /*7827*/;
  assign _13234_ = m_25[57] & _13232_ /*7826*/;
  assign r_25[57] = _13234_ | _13233_ /*7825*/;
  assign _13235_ = ~q[7] /*7824*/;
  assign _13236_ = sum_25[58] & q[7] /*7823*/;
  assign _13237_ = m_25[58] & _13235_ /*7822*/;
  assign r_25[58] = _13237_ | _13236_ /*7821*/;
  assign _13238_ = ~q[7] /*7820*/;
  assign _13239_ = sum_25[59] & q[7] /*7819*/;
  assign _13240_ = m_25[59] & _13238_ /*7818*/;
  assign r_25[59] = _13240_ | _13239_ /*7817*/;
  assign _13241_ = ~q[7] /*7816*/;
  assign _13242_ = sum_25[60] & q[7] /*7815*/;
  assign _13243_ = m_25[60] & _13241_ /*7814*/;
  assign r_25[60] = _13243_ | _13242_ /*7813*/;
  assign _13244_ = ~q[7] /*7812*/;
  assign _13245_ = sum_25[61] & q[7] /*7811*/;
  assign _13246_ = m_25[61] & _13244_ /*7810*/;
  assign r_25[61] = _13246_ | _13245_ /*7809*/;
  assign _13247_ = ~q[7] /*7808*/;
  assign _13248_ = sum_25[62] & q[7] /*7807*/;
  assign _13249_ = m_25[62] & _13247_ /*7806*/;
  assign r_25[62] = _13249_ | _13248_ /*7805*/;
  assign _13250_ = ~q[7] /*7804*/;
  assign _13251_ = sum_25[63] & q[7] /*7803*/;
  assign _13252_ = m_25[63] & _13250_ /*7802*/;
  assign r_25[63] = _13252_ | _13251_ /*7801*/;
  assign _13253_ = ~q[7] /*7800*/;
  assign _13254_ = sum_25[64] & q[7] /*7799*/;
  assign _13255_ = m_25[64] & _13253_ /*7798*/;
  assign r_25[64] = _13255_ | _13254_ /*7797*/;
  assign _13256_ = ~q[7] /*7796*/;
  assign _13257_ = sum_25[65] & q[7] /*7795*/;
  assign _13258_ = m_25[65] & _13256_ /*7794*/;
  assign r_25[65] = _13258_ | _13257_ /*7793*/;
  assign _13259_ = ~q[7] /*7792*/;
  assign _13260_ = sum_25[66] & q[7] /*7791*/;
  assign _13261_ = m_25[66] & _13259_ /*7790*/;
  assign r_25[66] = _13261_ | _13260_ /*7789*/;
  assign _13262_ = ~q[7] /*7788*/;
  assign _13263_ = sum_25[67] & q[7] /*7787*/;
  assign _13264_ = m_25[67] & _13262_ /*7786*/;
  assign r_25[67] = _13264_ | _13263_ /*7785*/;
  assign _13265_ = ~q[7] /*7784*/;
  assign _13266_ = sum_25[68] & q[7] /*7783*/;
  assign _13267_ = m_25[68] & _13265_ /*7782*/;
  assign r_25[68] = _13267_ | _13266_ /*7781*/;
  assign _13268_ = ~q[7] /*7780*/;
  assign _13269_ = sum_25[69] & q[7] /*7779*/;
  assign _13270_ = m_25[69] & _13268_ /*7778*/;
  assign r_25[69] = _13270_ | _13269_ /*7777*/;
  assign _13271_ = ~q[7] /*7776*/;
  assign _13272_ = sum_25[70] & q[7] /*7775*/;
  assign _13273_ = m_25[70] & _13271_ /*7774*/;
  assign r_25[70] = _13273_ | _13272_ /*7773*/;
  assign _13274_ = ~q[7] /*7772*/;
  assign _13275_ = sum_25[71] & q[7] /*7771*/;
  assign _13276_ = m_25[71] & _13274_ /*7770*/;
  assign r_25[71] = _13276_ | _13275_ /*7769*/;
  assign _13277_ = ~q[7] /*7768*/;
  assign _13278_ = sum_25[72] & q[7] /*7767*/;
  assign _13279_ = m_25[72] & _13277_ /*7766*/;
  assign r_25[72] = _13279_ | _13278_ /*7765*/;
  assign _13280_ = ~q[7] /*7764*/;
  assign _13281_ = sum_25[73] & q[7] /*7763*/;
  assign _13282_ = m_25[73] & _13280_ /*7762*/;
  assign r_25[73] = _13282_ | _13281_ /*7761*/;
  assign _13283_ = ~q[7] /*7760*/;
  assign _13284_ = sum_25[74] & q[7] /*7759*/;
  assign _13285_ = m_25[74] & _13283_ /*7758*/;
  assign r_25[74] = _13285_ | _13284_ /*7757*/;
  assign _13286_ = ~q[7] /*7756*/;
  assign _13287_ = sum_25[75] & q[7] /*7755*/;
  assign _13288_ = m_25[75] & _13286_ /*7754*/;
  assign r_25[75] = _13288_ | _13287_ /*7753*/;
  assign _13289_ = ~q[7] /*7752*/;
  assign _13290_ = sum_25[76] & q[7] /*7751*/;
  assign _13291_ = m_25[76] & _13289_ /*7750*/;
  assign r_25[76] = _13291_ | _13290_ /*7749*/;
  assign _13292_ = ~q[7] /*7748*/;
  assign _13293_ = sum_25[77] & q[7] /*7747*/;
  assign _13294_ = m_25[77] & _13292_ /*7746*/;
  assign r_25[77] = _13294_ | _13293_ /*7745*/;
  assign _13295_ = ~q[7] /*7744*/;
  assign _13296_ = sum_25[78] & q[7] /*7743*/;
  assign _13297_ = m_25[78] & _13295_ /*7742*/;
  assign r_25[78] = _13297_ | _13296_ /*7741*/;
  assign _13298_ = ~q[7] /*7740*/;
  assign _13299_ = sum_25[79] & q[7] /*7739*/;
  assign _13300_ = m_25[79] & _13298_ /*7738*/;
  assign r_25[79] = _13300_ | _13299_ /*7737*/;
  assign _13301_ = ~q[7] /*7736*/;
  assign _13302_ = sum_25[80] & q[7] /*7735*/;
  assign _13303_ = m_25[80] & _13301_ /*7734*/;
  assign r_25[80] = _13303_ | _13302_ /*7733*/;
  assign _13304_ = ~q[7] /*7732*/;
  assign _13305_ = sum_25[81] & q[7] /*7731*/;
  assign _13306_ = m_25[81] & _13304_ /*7730*/;
  assign r_25[81] = _13306_ | _13305_ /*7729*/;
  assign _13307_ = ~q[7] /*7728*/;
  assign _13308_ = sum_25[82] & q[7] /*7727*/;
  assign _13309_ = m_25[82] & _13307_ /*7726*/;
  assign r_25[82] = _13309_ | _13308_ /*7725*/;
  assign _13310_ = ~q[7] /*7724*/;
  assign _13311_ = sum_25[83] & q[7] /*7723*/;
  assign _13312_ = m_25[83] & _13310_ /*7722*/;
  assign r_25[83] = _13312_ | _13311_ /*7721*/;
  assign _13313_ = ~q[7] /*7720*/;
  assign _13314_ = sum_25[84] & q[7] /*7719*/;
  assign _13315_ = m_25[84] & _13313_ /*7718*/;
  assign r_25[84] = _13315_ | _13314_ /*7717*/;
  assign _13316_ = ~q[7] /*7716*/;
  assign _13317_ = sum_25[85] & q[7] /*7715*/;
  assign _13318_ = m_25[85] & _13316_ /*7714*/;
  assign r_25[85] = _13318_ | _13317_ /*7713*/;
  assign _13319_ = ~q[7] /*7712*/;
  assign _13320_ = sum_25[86] & q[7] /*7711*/;
  assign _13321_ = m_25[86] & _13319_ /*7710*/;
  assign r_25[86] = _13321_ | _13320_ /*7709*/;
  assign _13322_ = ~q[7] /*7708*/;
  assign _13323_ = sum_25[87] & q[7] /*7707*/;
  assign _13324_ = m_25[87] & _13322_ /*7706*/;
  assign r_25[87] = _13324_ | _13323_ /*7705*/;
  assign inv_26[0] = oneWire /*7596*/;
  assign inv_26[1] = oneWire /*7590*/;
  assign inv_26[2] = oneWire /*7584*/;
  assign inv_26[3] = oneWire /*7578*/;
  assign inv_26[4] = oneWire /*7572*/;
  assign inv_26[5] = oneWire /*7566*/;
  assign inv_26[6] = ~div[0] /*7560*/;
  assign inv_26[7] = ~div[1] /*7554*/;
  assign inv_26[8] = ~div[2] /*7548*/;
  assign inv_26[9] = ~div[3] /*7542*/;
  assign inv_26[10] = ~div[4] /*7536*/;
  assign inv_26[11] = ~div[5] /*7530*/;
  assign inv_26[12] = ~div[6] /*7524*/;
  assign inv_26[13] = ~div[7] /*7518*/;
  assign inv_26[14] = ~div[8] /*7512*/;
  assign inv_26[15] = ~div[9] /*7506*/;
  assign inv_26[16] = ~div[10] /*7500*/;
  assign inv_26[17] = ~div[11] /*7494*/;
  assign inv_26[18] = ~div[12] /*7488*/;
  assign inv_26[19] = ~div[13] /*7482*/;
  assign inv_26[20] = ~div[14] /*7476*/;
  assign inv_26[21] = ~div[15] /*7470*/;
  assign inv_26[22] = ~div[16] /*7464*/;
  assign inv_26[23] = ~div[17] /*7458*/;
  assign inv_26[24] = ~div[18] /*7452*/;
  assign inv_26[25] = ~div[19] /*7446*/;
  assign inv_26[26] = ~div[20] /*7440*/;
  assign inv_26[27] = ~div[21] /*7434*/;
  assign inv_26[28] = ~div[22] /*7428*/;
  assign inv_26[29] = ~div[23] /*7422*/;
  assign inv_26[30] = ~div[24] /*7416*/;
  assign inv_26[31] = ~div[25] /*7410*/;
  assign inv_26[32] = ~div[26] /*7404*/;
  assign inv_26[33] = ~div[27] /*7398*/;
  assign inv_26[34] = ~div[28] /*7392*/;
  assign inv_26[35] = ~div[29] /*7386*/;
  assign inv_26[36] = ~div[30] /*7380*/;
  assign inv_26[37] = oneWire /*7374*/;
  assign inv_26[38] = oneWire /*7368*/;
  assign inv_26[39] = oneWire /*7362*/;
  assign inv_26[40] = oneWire /*7356*/;
  assign inv_26[41] = oneWire /*7350*/;
  assign inv_26[42] = oneWire /*7344*/;
  assign inv_26[43] = oneWire /*7338*/;
  assign inv_26[44] = oneWire /*7332*/;
  assign inv_26[45] = oneWire /*7326*/;
  assign inv_26[46] = oneWire /*7320*/;
  assign inv_26[47] = oneWire /*7314*/;
  assign inv_26[48] = oneWire /*7308*/;
  assign inv_26[49] = oneWire /*7302*/;
  assign inv_26[50] = oneWire /*7296*/;
  assign inv_26[51] = oneWire /*7290*/;
  assign inv_26[52] = oneWire /*7284*/;
  assign inv_26[53] = oneWire /*7278*/;
  assign inv_26[54] = oneWire /*7272*/;
  assign inv_26[55] = oneWire /*7266*/;
  assign inv_26[56] = oneWire /*7260*/;
  assign inv_26[57] = oneWire /*7254*/;
  assign inv_26[58] = oneWire /*7248*/;
  assign inv_26[59] = oneWire /*7242*/;
  assign inv_26[60] = oneWire /*7236*/;
  assign inv_26[61] = oneWire /*7230*/;
  assign inv_26[62] = oneWire /*7224*/;
  assign inv_26[63] = oneWire /*7218*/;
  assign inv_26[64] = oneWire /*7212*/;
  assign inv_26[65] = oneWire /*7206*/;
  assign inv_26[66] = oneWire /*7200*/;
  assign inv_26[67] = oneWire /*7194*/;
  assign inv_26[68] = oneWire /*7188*/;
  assign inv_26[69] = oneWire /*7182*/;
  assign inv_26[70] = oneWire /*7176*/;
  assign inv_26[71] = oneWire /*7170*/;
  assign inv_26[72] = oneWire /*7164*/;
  assign inv_26[73] = oneWire /*7158*/;
  assign inv_26[74] = oneWire /*7152*/;
  assign inv_26[75] = oneWire /*7146*/;
  assign inv_26[76] = oneWire /*7140*/;
  assign inv_26[77] = oneWire /*7134*/;
  assign inv_26[78] = oneWire /*7128*/;
  assign inv_26[79] = oneWire /*7122*/;
  assign inv_26[80] = oneWire /*7116*/;
  assign inv_26[81] = oneWire /*7110*/;
  assign inv_26[82] = oneWire /*7104*/;
  assign inv_26[83] = oneWire /*7098*/;
  assign inv_26[84] = oneWire /*7092*/;
  assign inv_26[85] = oneWire /*7086*/;
  assign inv_26[86] = oneWire /*7080*/;
  assign inv_26[87] = oneWire /*7074*/;
  assign _13325_ = inv_26[0] ^ r_25[0] /*7595*/;
  assign sum_26[0] = _13325_ ^ oneWire /*7594*/;
  assign _13326_ = _13325_ & oneWire /*7593*/;
  assign _13327_ = inv_26[0] & r_25[0] /*7592*/;
  assign _13328_ = _13326_ | _13327_ /*7591*/;
  assign _13329_ = inv_26[1] ^ r_25[1] /*7589*/;
  assign sum_26[1] = _13329_ ^ _13328_ /*7588*/;
  assign _13330_ = _13329_ & _13328_ /*7587*/;
  assign _13331_ = inv_26[1] & r_25[1] /*7586*/;
  assign _13332_ = _13330_ | _13331_ /*7585*/;
  assign _13333_ = inv_26[2] ^ r_25[2] /*7583*/;
  assign sum_26[2] = _13333_ ^ _13332_ /*7582*/;
  assign _13334_ = _13333_ & _13332_ /*7581*/;
  assign _13335_ = inv_26[2] & r_25[2] /*7580*/;
  assign _13336_ = _13334_ | _13335_ /*7579*/;
  assign _13337_ = inv_26[3] ^ r_25[3] /*7577*/;
  assign sum_26[3] = _13337_ ^ _13336_ /*7576*/;
  assign _13338_ = _13337_ & _13336_ /*7575*/;
  assign _13339_ = inv_26[3] & r_25[3] /*7574*/;
  assign _13340_ = _13338_ | _13339_ /*7573*/;
  assign _13341_ = inv_26[4] ^ r_25[4] /*7571*/;
  assign sum_26[4] = _13341_ ^ _13340_ /*7570*/;
  assign _13342_ = _13341_ & _13340_ /*7569*/;
  assign _13343_ = inv_26[4] & r_25[4] /*7568*/;
  assign _13344_ = _13342_ | _13343_ /*7567*/;
  assign _13345_ = inv_26[5] ^ r_25[5] /*7565*/;
  assign sum_26[5] = _13345_ ^ _13344_ /*7564*/;
  assign _13346_ = _13345_ & _13344_ /*7563*/;
  assign _13347_ = inv_26[5] & r_25[5] /*7562*/;
  assign _13348_ = _13346_ | _13347_ /*7561*/;
  assign _13349_ = inv_26[6] ^ r_25[6] /*7559*/;
  assign sum_26[6] = _13349_ ^ _13348_ /*7558*/;
  assign _13350_ = _13349_ & _13348_ /*7557*/;
  assign _13351_ = inv_26[6] & r_25[6] /*7556*/;
  assign _13352_ = _13350_ | _13351_ /*7555*/;
  assign _13353_ = inv_26[7] ^ r_25[7] /*7553*/;
  assign sum_26[7] = _13353_ ^ _13352_ /*7552*/;
  assign _13354_ = _13353_ & _13352_ /*7551*/;
  assign _13355_ = inv_26[7] & r_25[7] /*7550*/;
  assign _13356_ = _13354_ | _13355_ /*7549*/;
  assign _13357_ = inv_26[8] ^ r_25[8] /*7547*/;
  assign sum_26[8] = _13357_ ^ _13356_ /*7546*/;
  assign _13358_ = _13357_ & _13356_ /*7545*/;
  assign _13359_ = inv_26[8] & r_25[8] /*7544*/;
  assign _13360_ = _13358_ | _13359_ /*7543*/;
  assign _13361_ = inv_26[9] ^ r_25[9] /*7541*/;
  assign sum_26[9] = _13361_ ^ _13360_ /*7540*/;
  assign _13362_ = _13361_ & _13360_ /*7539*/;
  assign _13363_ = inv_26[9] & r_25[9] /*7538*/;
  assign _13364_ = _13362_ | _13363_ /*7537*/;
  assign _13365_ = inv_26[10] ^ r_25[10] /*7535*/;
  assign sum_26[10] = _13365_ ^ _13364_ /*7534*/;
  assign _13366_ = _13365_ & _13364_ /*7533*/;
  assign _13367_ = inv_26[10] & r_25[10] /*7532*/;
  assign _13368_ = _13366_ | _13367_ /*7531*/;
  assign _13369_ = inv_26[11] ^ r_25[11] /*7529*/;
  assign sum_26[11] = _13369_ ^ _13368_ /*7528*/;
  assign _13370_ = _13369_ & _13368_ /*7527*/;
  assign _13371_ = inv_26[11] & r_25[11] /*7526*/;
  assign _13372_ = _13370_ | _13371_ /*7525*/;
  assign _13373_ = inv_26[12] ^ r_25[12] /*7523*/;
  assign sum_26[12] = _13373_ ^ _13372_ /*7522*/;
  assign _13374_ = _13373_ & _13372_ /*7521*/;
  assign _13375_ = inv_26[12] & r_25[12] /*7520*/;
  assign _13376_ = _13374_ | _13375_ /*7519*/;
  assign _13377_ = inv_26[13] ^ r_25[13] /*7517*/;
  assign sum_26[13] = _13377_ ^ _13376_ /*7516*/;
  assign _13378_ = _13377_ & _13376_ /*7515*/;
  assign _13379_ = inv_26[13] & r_25[13] /*7514*/;
  assign _13380_ = _13378_ | _13379_ /*7513*/;
  assign _13381_ = inv_26[14] ^ r_25[14] /*7511*/;
  assign sum_26[14] = _13381_ ^ _13380_ /*7510*/;
  assign _13382_ = _13381_ & _13380_ /*7509*/;
  assign _13383_ = inv_26[14] & r_25[14] /*7508*/;
  assign _13384_ = _13382_ | _13383_ /*7507*/;
  assign _13385_ = inv_26[15] ^ r_25[15] /*7505*/;
  assign sum_26[15] = _13385_ ^ _13384_ /*7504*/;
  assign _13386_ = _13385_ & _13384_ /*7503*/;
  assign _13387_ = inv_26[15] & r_25[15] /*7502*/;
  assign _13388_ = _13386_ | _13387_ /*7501*/;
  assign _13389_ = inv_26[16] ^ r_25[16] /*7499*/;
  assign sum_26[16] = _13389_ ^ _13388_ /*7498*/;
  assign _13390_ = _13389_ & _13388_ /*7497*/;
  assign _13391_ = inv_26[16] & r_25[16] /*7496*/;
  assign _13392_ = _13390_ | _13391_ /*7495*/;
  assign _13393_ = inv_26[17] ^ r_25[17] /*7493*/;
  assign sum_26[17] = _13393_ ^ _13392_ /*7492*/;
  assign _13394_ = _13393_ & _13392_ /*7491*/;
  assign _13395_ = inv_26[17] & r_25[17] /*7490*/;
  assign _13396_ = _13394_ | _13395_ /*7489*/;
  assign _13397_ = inv_26[18] ^ r_25[18] /*7487*/;
  assign sum_26[18] = _13397_ ^ _13396_ /*7486*/;
  assign _13398_ = _13397_ & _13396_ /*7485*/;
  assign _13399_ = inv_26[18] & r_25[18] /*7484*/;
  assign _13400_ = _13398_ | _13399_ /*7483*/;
  assign _13401_ = inv_26[19] ^ r_25[19] /*7481*/;
  assign sum_26[19] = _13401_ ^ _13400_ /*7480*/;
  assign _13402_ = _13401_ & _13400_ /*7479*/;
  assign _13403_ = inv_26[19] & r_25[19] /*7478*/;
  assign _13404_ = _13402_ | _13403_ /*7477*/;
  assign _13405_ = inv_26[20] ^ r_25[20] /*7475*/;
  assign sum_26[20] = _13405_ ^ _13404_ /*7474*/;
  assign _13406_ = _13405_ & _13404_ /*7473*/;
  assign _13407_ = inv_26[20] & r_25[20] /*7472*/;
  assign _13408_ = _13406_ | _13407_ /*7471*/;
  assign _13409_ = inv_26[21] ^ r_25[21] /*7469*/;
  assign sum_26[21] = _13409_ ^ _13408_ /*7468*/;
  assign _13410_ = _13409_ & _13408_ /*7467*/;
  assign _13411_ = inv_26[21] & r_25[21] /*7466*/;
  assign _13412_ = _13410_ | _13411_ /*7465*/;
  assign _13413_ = inv_26[22] ^ r_25[22] /*7463*/;
  assign sum_26[22] = _13413_ ^ _13412_ /*7462*/;
  assign _13414_ = _13413_ & _13412_ /*7461*/;
  assign _13415_ = inv_26[22] & r_25[22] /*7460*/;
  assign _13416_ = _13414_ | _13415_ /*7459*/;
  assign _13417_ = inv_26[23] ^ r_25[23] /*7457*/;
  assign sum_26[23] = _13417_ ^ _13416_ /*7456*/;
  assign _13418_ = _13417_ & _13416_ /*7455*/;
  assign _13419_ = inv_26[23] & r_25[23] /*7454*/;
  assign _13420_ = _13418_ | _13419_ /*7453*/;
  assign _13421_ = inv_26[24] ^ r_25[24] /*7451*/;
  assign sum_26[24] = _13421_ ^ _13420_ /*7450*/;
  assign _13422_ = _13421_ & _13420_ /*7449*/;
  assign _13423_ = inv_26[24] & r_25[24] /*7448*/;
  assign _13424_ = _13422_ | _13423_ /*7447*/;
  assign _13425_ = inv_26[25] ^ r_25[25] /*7445*/;
  assign sum_26[25] = _13425_ ^ _13424_ /*7444*/;
  assign _13426_ = _13425_ & _13424_ /*7443*/;
  assign _13427_ = inv_26[25] & r_25[25] /*7442*/;
  assign _13428_ = _13426_ | _13427_ /*7441*/;
  assign _13429_ = inv_26[26] ^ r_25[26] /*7439*/;
  assign sum_26[26] = _13429_ ^ _13428_ /*7438*/;
  assign _13430_ = _13429_ & _13428_ /*7437*/;
  assign _13431_ = inv_26[26] & r_25[26] /*7436*/;
  assign _13432_ = _13430_ | _13431_ /*7435*/;
  assign _13433_ = inv_26[27] ^ r_25[27] /*7433*/;
  assign sum_26[27] = _13433_ ^ _13432_ /*7432*/;
  assign _13434_ = _13433_ & _13432_ /*7431*/;
  assign _13435_ = inv_26[27] & r_25[27] /*7430*/;
  assign _13436_ = _13434_ | _13435_ /*7429*/;
  assign _13437_ = inv_26[28] ^ r_25[28] /*7427*/;
  assign sum_26[28] = _13437_ ^ _13436_ /*7426*/;
  assign _13438_ = _13437_ & _13436_ /*7425*/;
  assign _13439_ = inv_26[28] & r_25[28] /*7424*/;
  assign _13440_ = _13438_ | _13439_ /*7423*/;
  assign _13441_ = inv_26[29] ^ r_25[29] /*7421*/;
  assign sum_26[29] = _13441_ ^ _13440_ /*7420*/;
  assign _13442_ = _13441_ & _13440_ /*7419*/;
  assign _13443_ = inv_26[29] & r_25[29] /*7418*/;
  assign _13444_ = _13442_ | _13443_ /*7417*/;
  assign _13445_ = inv_26[30] ^ r_25[30] /*7415*/;
  assign sum_26[30] = _13445_ ^ _13444_ /*7414*/;
  assign _13446_ = _13445_ & _13444_ /*7413*/;
  assign _13447_ = inv_26[30] & r_25[30] /*7412*/;
  assign _13448_ = _13446_ | _13447_ /*7411*/;
  assign _13449_ = inv_26[31] ^ r_25[31] /*7409*/;
  assign sum_26[31] = _13449_ ^ _13448_ /*7408*/;
  assign _13450_ = _13449_ & _13448_ /*7407*/;
  assign _13451_ = inv_26[31] & r_25[31] /*7406*/;
  assign _13452_ = _13450_ | _13451_ /*7405*/;
  assign _13453_ = inv_26[32] ^ r_25[32] /*7403*/;
  assign sum_26[32] = _13453_ ^ _13452_ /*7402*/;
  assign _13454_ = _13453_ & _13452_ /*7401*/;
  assign _13455_ = inv_26[32] & r_25[32] /*7400*/;
  assign _13456_ = _13454_ | _13455_ /*7399*/;
  assign _13457_ = inv_26[33] ^ r_25[33] /*7397*/;
  assign sum_26[33] = _13457_ ^ _13456_ /*7396*/;
  assign _13458_ = _13457_ & _13456_ /*7395*/;
  assign _13459_ = inv_26[33] & r_25[33] /*7394*/;
  assign _13460_ = _13458_ | _13459_ /*7393*/;
  assign _13461_ = inv_26[34] ^ r_25[34] /*7391*/;
  assign sum_26[34] = _13461_ ^ _13460_ /*7390*/;
  assign _13462_ = _13461_ & _13460_ /*7389*/;
  assign _13463_ = inv_26[34] & r_25[34] /*7388*/;
  assign _13464_ = _13462_ | _13463_ /*7387*/;
  assign _13465_ = inv_26[35] ^ r_25[35] /*7385*/;
  assign sum_26[35] = _13465_ ^ _13464_ /*7384*/;
  assign _13466_ = _13465_ & _13464_ /*7383*/;
  assign _13467_ = inv_26[35] & r_25[35] /*7382*/;
  assign _13468_ = _13466_ | _13467_ /*7381*/;
  assign _13469_ = inv_26[36] ^ r_25[36] /*7379*/;
  assign sum_26[36] = _13469_ ^ _13468_ /*7378*/;
  assign _13470_ = _13469_ & _13468_ /*7377*/;
  assign _13471_ = inv_26[36] & r_25[36] /*7376*/;
  assign _13472_ = _13470_ | _13471_ /*7375*/;
  assign _13473_ = inv_26[37] ^ r_25[37] /*7373*/;
  assign sum_26[37] = _13473_ ^ _13472_ /*7372*/;
  assign _13474_ = _13473_ & _13472_ /*7371*/;
  assign _13475_ = inv_26[37] & r_25[37] /*7370*/;
  assign _13476_ = _13474_ | _13475_ /*7369*/;
  assign _13477_ = inv_26[38] ^ r_25[38] /*7367*/;
  assign sum_26[38] = _13477_ ^ _13476_ /*7366*/;
  assign _13478_ = _13477_ & _13476_ /*7365*/;
  assign _13479_ = inv_26[38] & r_25[38] /*7364*/;
  assign _13480_ = _13478_ | _13479_ /*7363*/;
  assign _13481_ = inv_26[39] ^ r_25[39] /*7361*/;
  assign sum_26[39] = _13481_ ^ _13480_ /*7360*/;
  assign _13482_ = _13481_ & _13480_ /*7359*/;
  assign _13483_ = inv_26[39] & r_25[39] /*7358*/;
  assign _13484_ = _13482_ | _13483_ /*7357*/;
  assign _13485_ = inv_26[40] ^ r_25[40] /*7355*/;
  assign sum_26[40] = _13485_ ^ _13484_ /*7354*/;
  assign _13486_ = _13485_ & _13484_ /*7353*/;
  assign _13487_ = inv_26[40] & r_25[40] /*7352*/;
  assign _13488_ = _13486_ | _13487_ /*7351*/;
  assign _13489_ = inv_26[41] ^ r_25[41] /*7349*/;
  assign sum_26[41] = _13489_ ^ _13488_ /*7348*/;
  assign _13490_ = _13489_ & _13488_ /*7347*/;
  assign _13491_ = inv_26[41] & r_25[41] /*7346*/;
  assign _13492_ = _13490_ | _13491_ /*7345*/;
  assign _13493_ = inv_26[42] ^ r_25[42] /*7343*/;
  assign sum_26[42] = _13493_ ^ _13492_ /*7342*/;
  assign _13494_ = _13493_ & _13492_ /*7341*/;
  assign _13495_ = inv_26[42] & r_25[42] /*7340*/;
  assign _13496_ = _13494_ | _13495_ /*7339*/;
  assign _13497_ = inv_26[43] ^ r_25[43] /*7337*/;
  assign sum_26[43] = _13497_ ^ _13496_ /*7336*/;
  assign _13498_ = _13497_ & _13496_ /*7335*/;
  assign _13499_ = inv_26[43] & r_25[43] /*7334*/;
  assign _13500_ = _13498_ | _13499_ /*7333*/;
  assign _13501_ = inv_26[44] ^ r_25[44] /*7331*/;
  assign sum_26[44] = _13501_ ^ _13500_ /*7330*/;
  assign _13502_ = _13501_ & _13500_ /*7329*/;
  assign _13503_ = inv_26[44] & r_25[44] /*7328*/;
  assign _13504_ = _13502_ | _13503_ /*7327*/;
  assign _13505_ = inv_26[45] ^ r_25[45] /*7325*/;
  assign sum_26[45] = _13505_ ^ _13504_ /*7324*/;
  assign _13506_ = _13505_ & _13504_ /*7323*/;
  assign _13507_ = inv_26[45] & r_25[45] /*7322*/;
  assign _13508_ = _13506_ | _13507_ /*7321*/;
  assign _13509_ = inv_26[46] ^ r_25[46] /*7319*/;
  assign sum_26[46] = _13509_ ^ _13508_ /*7318*/;
  assign _13510_ = _13509_ & _13508_ /*7317*/;
  assign _13511_ = inv_26[46] & r_25[46] /*7316*/;
  assign _13512_ = _13510_ | _13511_ /*7315*/;
  assign _13513_ = inv_26[47] ^ r_25[47] /*7313*/;
  assign sum_26[47] = _13513_ ^ _13512_ /*7312*/;
  assign _13514_ = _13513_ & _13512_ /*7311*/;
  assign _13515_ = inv_26[47] & r_25[47] /*7310*/;
  assign _13516_ = _13514_ | _13515_ /*7309*/;
  assign _13517_ = inv_26[48] ^ r_25[48] /*7307*/;
  assign sum_26[48] = _13517_ ^ _13516_ /*7306*/;
  assign _13518_ = _13517_ & _13516_ /*7305*/;
  assign _13519_ = inv_26[48] & r_25[48] /*7304*/;
  assign _13520_ = _13518_ | _13519_ /*7303*/;
  assign _13521_ = inv_26[49] ^ r_25[49] /*7301*/;
  assign sum_26[49] = _13521_ ^ _13520_ /*7300*/;
  assign _13522_ = _13521_ & _13520_ /*7299*/;
  assign _13523_ = inv_26[49] & r_25[49] /*7298*/;
  assign _13524_ = _13522_ | _13523_ /*7297*/;
  assign _13525_ = inv_26[50] ^ r_25[50] /*7295*/;
  assign sum_26[50] = _13525_ ^ _13524_ /*7294*/;
  assign _13526_ = _13525_ & _13524_ /*7293*/;
  assign _13527_ = inv_26[50] & r_25[50] /*7292*/;
  assign _13528_ = _13526_ | _13527_ /*7291*/;
  assign _13529_ = inv_26[51] ^ r_25[51] /*7289*/;
  assign sum_26[51] = _13529_ ^ _13528_ /*7288*/;
  assign _13530_ = _13529_ & _13528_ /*7287*/;
  assign _13531_ = inv_26[51] & r_25[51] /*7286*/;
  assign _13532_ = _13530_ | _13531_ /*7285*/;
  assign _13533_ = inv_26[52] ^ r_25[52] /*7283*/;
  assign sum_26[52] = _13533_ ^ _13532_ /*7282*/;
  assign _13534_ = _13533_ & _13532_ /*7281*/;
  assign _13535_ = inv_26[52] & r_25[52] /*7280*/;
  assign _13536_ = _13534_ | _13535_ /*7279*/;
  assign _13537_ = inv_26[53] ^ r_25[53] /*7277*/;
  assign sum_26[53] = _13537_ ^ _13536_ /*7276*/;
  assign _13538_ = _13537_ & _13536_ /*7275*/;
  assign _13539_ = inv_26[53] & r_25[53] /*7274*/;
  assign _13540_ = _13538_ | _13539_ /*7273*/;
  assign _13541_ = inv_26[54] ^ r_25[54] /*7271*/;
  assign sum_26[54] = _13541_ ^ _13540_ /*7270*/;
  assign _13542_ = _13541_ & _13540_ /*7269*/;
  assign _13543_ = inv_26[54] & r_25[54] /*7268*/;
  assign _13544_ = _13542_ | _13543_ /*7267*/;
  assign _13545_ = inv_26[55] ^ r_25[55] /*7265*/;
  assign sum_26[55] = _13545_ ^ _13544_ /*7264*/;
  assign _13546_ = _13545_ & _13544_ /*7263*/;
  assign _13547_ = inv_26[55] & r_25[55] /*7262*/;
  assign _13548_ = _13546_ | _13547_ /*7261*/;
  assign _13549_ = inv_26[56] ^ r_25[56] /*7259*/;
  assign sum_26[56] = _13549_ ^ _13548_ /*7258*/;
  assign _13550_ = _13549_ & _13548_ /*7257*/;
  assign _13551_ = inv_26[56] & r_25[56] /*7256*/;
  assign _13552_ = _13550_ | _13551_ /*7255*/;
  assign _13553_ = inv_26[57] ^ r_25[57] /*7253*/;
  assign sum_26[57] = _13553_ ^ _13552_ /*7252*/;
  assign _13554_ = _13553_ & _13552_ /*7251*/;
  assign _13555_ = inv_26[57] & r_25[57] /*7250*/;
  assign _13556_ = _13554_ | _13555_ /*7249*/;
  assign _13557_ = inv_26[58] ^ r_25[58] /*7247*/;
  assign sum_26[58] = _13557_ ^ _13556_ /*7246*/;
  assign _13558_ = _13557_ & _13556_ /*7245*/;
  assign _13559_ = inv_26[58] & r_25[58] /*7244*/;
  assign _13560_ = _13558_ | _13559_ /*7243*/;
  assign _13561_ = inv_26[59] ^ r_25[59] /*7241*/;
  assign sum_26[59] = _13561_ ^ _13560_ /*7240*/;
  assign _13562_ = _13561_ & _13560_ /*7239*/;
  assign _13563_ = inv_26[59] & r_25[59] /*7238*/;
  assign _13564_ = _13562_ | _13563_ /*7237*/;
  assign _13565_ = inv_26[60] ^ r_25[60] /*7235*/;
  assign sum_26[60] = _13565_ ^ _13564_ /*7234*/;
  assign _13566_ = _13565_ & _13564_ /*7233*/;
  assign _13567_ = inv_26[60] & r_25[60] /*7232*/;
  assign _13568_ = _13566_ | _13567_ /*7231*/;
  assign _13569_ = inv_26[61] ^ r_25[61] /*7229*/;
  assign sum_26[61] = _13569_ ^ _13568_ /*7228*/;
  assign _13570_ = _13569_ & _13568_ /*7227*/;
  assign _13571_ = inv_26[61] & r_25[61] /*7226*/;
  assign _13572_ = _13570_ | _13571_ /*7225*/;
  assign _13573_ = inv_26[62] ^ r_25[62] /*7223*/;
  assign sum_26[62] = _13573_ ^ _13572_ /*7222*/;
  assign _13574_ = _13573_ & _13572_ /*7221*/;
  assign _13575_ = inv_26[62] & r_25[62] /*7220*/;
  assign _13576_ = _13574_ | _13575_ /*7219*/;
  assign _13577_ = inv_26[63] ^ r_25[63] /*7217*/;
  assign sum_26[63] = _13577_ ^ _13576_ /*7216*/;
  assign _13578_ = _13577_ & _13576_ /*7215*/;
  assign _13579_ = inv_26[63] & r_25[63] /*7214*/;
  assign _13580_ = _13578_ | _13579_ /*7213*/;
  assign _13581_ = inv_26[64] ^ r_25[64] /*7211*/;
  assign sum_26[64] = _13581_ ^ _13580_ /*7210*/;
  assign _13582_ = _13581_ & _13580_ /*7209*/;
  assign _13583_ = inv_26[64] & r_25[64] /*7208*/;
  assign _13584_ = _13582_ | _13583_ /*7207*/;
  assign _13585_ = inv_26[65] ^ r_25[65] /*7205*/;
  assign sum_26[65] = _13585_ ^ _13584_ /*7204*/;
  assign _13586_ = _13585_ & _13584_ /*7203*/;
  assign _13587_ = inv_26[65] & r_25[65] /*7202*/;
  assign _13588_ = _13586_ | _13587_ /*7201*/;
  assign _13589_ = inv_26[66] ^ r_25[66] /*7199*/;
  assign sum_26[66] = _13589_ ^ _13588_ /*7198*/;
  assign _13590_ = _13589_ & _13588_ /*7197*/;
  assign _13591_ = inv_26[66] & r_25[66] /*7196*/;
  assign _13592_ = _13590_ | _13591_ /*7195*/;
  assign _13593_ = inv_26[67] ^ r_25[67] /*7193*/;
  assign sum_26[67] = _13593_ ^ _13592_ /*7192*/;
  assign _13594_ = _13593_ & _13592_ /*7191*/;
  assign _13595_ = inv_26[67] & r_25[67] /*7190*/;
  assign _13596_ = _13594_ | _13595_ /*7189*/;
  assign _13597_ = inv_26[68] ^ r_25[68] /*7187*/;
  assign sum_26[68] = _13597_ ^ _13596_ /*7186*/;
  assign _13598_ = _13597_ & _13596_ /*7185*/;
  assign _13599_ = inv_26[68] & r_25[68] /*7184*/;
  assign _13600_ = _13598_ | _13599_ /*7183*/;
  assign _13601_ = inv_26[69] ^ r_25[69] /*7181*/;
  assign sum_26[69] = _13601_ ^ _13600_ /*7180*/;
  assign _13602_ = _13601_ & _13600_ /*7179*/;
  assign _13603_ = inv_26[69] & r_25[69] /*7178*/;
  assign _13604_ = _13602_ | _13603_ /*7177*/;
  assign _13605_ = inv_26[70] ^ r_25[70] /*7175*/;
  assign sum_26[70] = _13605_ ^ _13604_ /*7174*/;
  assign _13606_ = _13605_ & _13604_ /*7173*/;
  assign _13607_ = inv_26[70] & r_25[70] /*7172*/;
  assign _13608_ = _13606_ | _13607_ /*7171*/;
  assign _13609_ = inv_26[71] ^ r_25[71] /*7169*/;
  assign sum_26[71] = _13609_ ^ _13608_ /*7168*/;
  assign _13610_ = _13609_ & _13608_ /*7167*/;
  assign _13611_ = inv_26[71] & r_25[71] /*7166*/;
  assign _13612_ = _13610_ | _13611_ /*7165*/;
  assign _13613_ = inv_26[72] ^ r_25[72] /*7163*/;
  assign sum_26[72] = _13613_ ^ _13612_ /*7162*/;
  assign _13614_ = _13613_ & _13612_ /*7161*/;
  assign _13615_ = inv_26[72] & r_25[72] /*7160*/;
  assign _13616_ = _13614_ | _13615_ /*7159*/;
  assign _13617_ = inv_26[73] ^ r_25[73] /*7157*/;
  assign sum_26[73] = _13617_ ^ _13616_ /*7156*/;
  assign _13618_ = _13617_ & _13616_ /*7155*/;
  assign _13619_ = inv_26[73] & r_25[73] /*7154*/;
  assign _13620_ = _13618_ | _13619_ /*7153*/;
  assign _13621_ = inv_26[74] ^ r_25[74] /*7151*/;
  assign sum_26[74] = _13621_ ^ _13620_ /*7150*/;
  assign _13622_ = _13621_ & _13620_ /*7149*/;
  assign _13623_ = inv_26[74] & r_25[74] /*7148*/;
  assign _13624_ = _13622_ | _13623_ /*7147*/;
  assign _13625_ = inv_26[75] ^ r_25[75] /*7145*/;
  assign sum_26[75] = _13625_ ^ _13624_ /*7144*/;
  assign _13626_ = _13625_ & _13624_ /*7143*/;
  assign _13627_ = inv_26[75] & r_25[75] /*7142*/;
  assign _13628_ = _13626_ | _13627_ /*7141*/;
  assign _13629_ = inv_26[76] ^ r_25[76] /*7139*/;
  assign sum_26[76] = _13629_ ^ _13628_ /*7138*/;
  assign _13630_ = _13629_ & _13628_ /*7137*/;
  assign _13631_ = inv_26[76] & r_25[76] /*7136*/;
  assign _13632_ = _13630_ | _13631_ /*7135*/;
  assign _13633_ = inv_26[77] ^ r_25[77] /*7133*/;
  assign sum_26[77] = _13633_ ^ _13632_ /*7132*/;
  assign _13634_ = _13633_ & _13632_ /*7131*/;
  assign _13635_ = inv_26[77] & r_25[77] /*7130*/;
  assign _13636_ = _13634_ | _13635_ /*7129*/;
  assign _13637_ = inv_26[78] ^ r_25[78] /*7127*/;
  assign sum_26[78] = _13637_ ^ _13636_ /*7126*/;
  assign _13638_ = _13637_ & _13636_ /*7125*/;
  assign _13639_ = inv_26[78] & r_25[78] /*7124*/;
  assign _13640_ = _13638_ | _13639_ /*7123*/;
  assign _13641_ = inv_26[79] ^ r_25[79] /*7121*/;
  assign sum_26[79] = _13641_ ^ _13640_ /*7120*/;
  assign _13642_ = _13641_ & _13640_ /*7119*/;
  assign _13643_ = inv_26[79] & r_25[79] /*7118*/;
  assign _13644_ = _13642_ | _13643_ /*7117*/;
  assign _13645_ = inv_26[80] ^ r_25[80] /*7115*/;
  assign sum_26[80] = _13645_ ^ _13644_ /*7114*/;
  assign _13646_ = _13645_ & _13644_ /*7113*/;
  assign _13647_ = inv_26[80] & r_25[80] /*7112*/;
  assign _13648_ = _13646_ | _13647_ /*7111*/;
  assign _13649_ = inv_26[81] ^ r_25[81] /*7109*/;
  assign sum_26[81] = _13649_ ^ _13648_ /*7108*/;
  assign _13650_ = _13649_ & _13648_ /*7107*/;
  assign _13651_ = inv_26[81] & r_25[81] /*7106*/;
  assign _13652_ = _13650_ | _13651_ /*7105*/;
  assign _13653_ = inv_26[82] ^ r_25[82] /*7103*/;
  assign sum_26[82] = _13653_ ^ _13652_ /*7102*/;
  assign _13654_ = _13653_ & _13652_ /*7101*/;
  assign _13655_ = inv_26[82] & r_25[82] /*7100*/;
  assign _13656_ = _13654_ | _13655_ /*7099*/;
  assign _13657_ = inv_26[83] ^ r_25[83] /*7097*/;
  assign sum_26[83] = _13657_ ^ _13656_ /*7096*/;
  assign _13658_ = _13657_ & _13656_ /*7095*/;
  assign _13659_ = inv_26[83] & r_25[83] /*7094*/;
  assign _13660_ = _13658_ | _13659_ /*7093*/;
  assign _13661_ = inv_26[84] ^ r_25[84] /*7091*/;
  assign sum_26[84] = _13661_ ^ _13660_ /*7090*/;
  assign _13662_ = _13661_ & _13660_ /*7089*/;
  assign _13663_ = inv_26[84] & r_25[84] /*7088*/;
  assign _13664_ = _13662_ | _13663_ /*7087*/;
  assign _13665_ = inv_26[85] ^ r_25[85] /*7085*/;
  assign sum_26[85] = _13665_ ^ _13664_ /*7084*/;
  assign _13666_ = _13665_ & _13664_ /*7083*/;
  assign _13667_ = inv_26[85] & r_25[85] /*7082*/;
  assign _13668_ = _13666_ | _13667_ /*7081*/;
  assign _13669_ = inv_26[86] ^ r_25[86] /*7079*/;
  assign sum_26[86] = _13669_ ^ _13668_ /*7078*/;
  assign _13670_ = _13669_ & _13668_ /*7077*/;
  assign _13671_ = inv_26[86] & r_25[86] /*7076*/;
  assign _13672_ = _13670_ | _13671_ /*7075*/;
  assign _13673_ = inv_26[87] ^ r_25[87] /*7073*/;
  assign sum_26[87] = _13673_ ^ _13672_ /*7072*/;
  assign _13674_ = _13673_ & _13672_ /*7071*/;
  assign _13675_ = inv_26[87] & r_25[87] /*7070*/;
  assign _13676_ = _13674_ | _13675_ /*7069*/;
  assign _13677_ = _13676_ ^ _13672_ /*7068*/;
  assign _13678_ = ~_13677_ /*7067*/;
  assign _13679_ = sum_26[87] & _13678_ /*7066*/;
  assign _13680_ = _13677_ & _13676_ /*7065*/;
  assign sum_26[88] = _13680_ | _13679_ /*7064*/;
  assign q[6] = ~sum_26[88] /*7063*/;
  assign m_26[0] = r_25[0] /*7062*/;
  assign m_26[1] = r_25[1] /*7061*/;
  assign m_26[2] = r_25[2] /*7060*/;
  assign m_26[3] = r_25[3] /*7059*/;
  assign m_26[4] = r_25[4] /*7058*/;
  assign m_26[5] = r_25[5] /*7057*/;
  assign m_26[6] = r_25[6] /*7056*/;
  assign m_26[7] = r_25[7] /*7055*/;
  assign m_26[8] = r_25[8] /*7054*/;
  assign m_26[9] = r_25[9] /*7053*/;
  assign m_26[10] = r_25[10] /*7052*/;
  assign m_26[11] = r_25[11] /*7051*/;
  assign m_26[12] = r_25[12] /*7050*/;
  assign m_26[13] = r_25[13] /*7049*/;
  assign m_26[14] = r_25[14] /*7048*/;
  assign m_26[15] = r_25[15] /*7047*/;
  assign m_26[16] = r_25[16] /*7046*/;
  assign m_26[17] = r_25[17] /*7045*/;
  assign m_26[18] = r_25[18] /*7044*/;
  assign m_26[19] = r_25[19] /*7043*/;
  assign m_26[20] = r_25[20] /*7042*/;
  assign m_26[21] = r_25[21] /*7041*/;
  assign m_26[22] = r_25[22] /*7040*/;
  assign m_26[23] = r_25[23] /*7039*/;
  assign m_26[24] = r_25[24] /*7038*/;
  assign m_26[25] = r_25[25] /*7037*/;
  assign m_26[26] = r_25[26] /*7036*/;
  assign m_26[27] = r_25[27] /*7035*/;
  assign m_26[28] = r_25[28] /*7034*/;
  assign m_26[29] = r_25[29] /*7033*/;
  assign m_26[30] = r_25[30] /*7032*/;
  assign m_26[31] = r_25[31] /*7031*/;
  assign m_26[32] = r_25[32] /*7030*/;
  assign m_26[33] = r_25[33] /*7029*/;
  assign m_26[34] = r_25[34] /*7028*/;
  assign m_26[35] = r_25[35] /*7027*/;
  assign m_26[36] = r_25[36] /*7026*/;
  assign m_26[37] = r_25[37] /*7025*/;
  assign m_26[38] = r_25[38] /*7024*/;
  assign m_26[39] = r_25[39] /*7023*/;
  assign m_26[40] = r_25[40] /*7022*/;
  assign m_26[41] = r_25[41] /*7021*/;
  assign m_26[42] = r_25[42] /*7020*/;
  assign m_26[43] = r_25[43] /*7019*/;
  assign m_26[44] = r_25[44] /*7018*/;
  assign m_26[45] = r_25[45] /*7017*/;
  assign m_26[46] = r_25[46] /*7016*/;
  assign m_26[47] = r_25[47] /*7015*/;
  assign m_26[48] = r_25[48] /*7014*/;
  assign m_26[49] = r_25[49] /*7013*/;
  assign m_26[50] = r_25[50] /*7012*/;
  assign m_26[51] = r_25[51] /*7011*/;
  assign m_26[52] = r_25[52] /*7010*/;
  assign m_26[53] = r_25[53] /*7009*/;
  assign m_26[54] = r_25[54] /*7008*/;
  assign m_26[55] = r_25[55] /*7007*/;
  assign m_26[56] = r_25[56] /*7006*/;
  assign m_26[57] = r_25[57] /*7005*/;
  assign m_26[58] = r_25[58] /*7004*/;
  assign m_26[59] = r_25[59] /*7003*/;
  assign m_26[60] = r_25[60] /*7002*/;
  assign m_26[61] = r_25[61] /*7001*/;
  assign m_26[62] = r_25[62] /*7000*/;
  assign m_26[63] = r_25[63] /*6999*/;
  assign m_26[64] = r_25[64] /*6998*/;
  assign m_26[65] = r_25[65] /*6997*/;
  assign m_26[66] = r_25[66] /*6996*/;
  assign m_26[67] = r_25[67] /*6995*/;
  assign m_26[68] = r_25[68] /*6994*/;
  assign m_26[69] = r_25[69] /*6993*/;
  assign m_26[70] = r_25[70] /*6992*/;
  assign m_26[71] = r_25[71] /*6991*/;
  assign m_26[72] = r_25[72] /*6990*/;
  assign m_26[73] = r_25[73] /*6989*/;
  assign m_26[74] = r_25[74] /*6988*/;
  assign m_26[75] = r_25[75] /*6987*/;
  assign m_26[76] = r_25[76] /*6986*/;
  assign m_26[77] = r_25[77] /*6985*/;
  assign m_26[78] = r_25[78] /*6984*/;
  assign m_26[79] = r_25[79] /*6983*/;
  assign m_26[80] = r_25[80] /*6982*/;
  assign m_26[81] = r_25[81] /*6981*/;
  assign m_26[82] = r_25[82] /*6980*/;
  assign m_26[83] = r_25[83] /*6979*/;
  assign m_26[84] = r_25[84] /*6978*/;
  assign m_26[85] = r_25[85] /*6977*/;
  assign m_26[86] = r_25[86] /*6976*/;
  assign m_26[87] = r_25[87] /*6975*/;
  assign m_26[88] = r_25[87] /*6974*/;
  assign _13682_ = ~q[6] /*6973*/;
  assign _13683_ = sum_26[0] & q[6] /*6972*/;
  assign _13684_ = m_26[0] & _13682_ /*6971*/;
  assign r_26[0] = _13684_ | _13683_ /*6970*/;
  assign _13685_ = ~q[6] /*6969*/;
  assign _13686_ = sum_26[1] & q[6] /*6968*/;
  assign _13687_ = m_26[1] & _13685_ /*6967*/;
  assign r_26[1] = _13687_ | _13686_ /*6966*/;
  assign _13688_ = ~q[6] /*6965*/;
  assign _13689_ = sum_26[2] & q[6] /*6964*/;
  assign _13690_ = m_26[2] & _13688_ /*6963*/;
  assign r_26[2] = _13690_ | _13689_ /*6962*/;
  assign _13691_ = ~q[6] /*6961*/;
  assign _13692_ = sum_26[3] & q[6] /*6960*/;
  assign _13693_ = m_26[3] & _13691_ /*6959*/;
  assign r_26[3] = _13693_ | _13692_ /*6958*/;
  assign _13694_ = ~q[6] /*6957*/;
  assign _13695_ = sum_26[4] & q[6] /*6956*/;
  assign _13696_ = m_26[4] & _13694_ /*6955*/;
  assign r_26[4] = _13696_ | _13695_ /*6954*/;
  assign _13697_ = ~q[6] /*6953*/;
  assign _13698_ = sum_26[5] & q[6] /*6952*/;
  assign _13699_ = m_26[5] & _13697_ /*6951*/;
  assign r_26[5] = _13699_ | _13698_ /*6950*/;
  assign _13700_ = ~q[6] /*6949*/;
  assign _13701_ = sum_26[6] & q[6] /*6948*/;
  assign _13702_ = m_26[6] & _13700_ /*6947*/;
  assign r_26[6] = _13702_ | _13701_ /*6946*/;
  assign _13703_ = ~q[6] /*6945*/;
  assign _13704_ = sum_26[7] & q[6] /*6944*/;
  assign _13705_ = m_26[7] & _13703_ /*6943*/;
  assign r_26[7] = _13705_ | _13704_ /*6942*/;
  assign _13706_ = ~q[6] /*6941*/;
  assign _13707_ = sum_26[8] & q[6] /*6940*/;
  assign _13708_ = m_26[8] & _13706_ /*6939*/;
  assign r_26[8] = _13708_ | _13707_ /*6938*/;
  assign _13709_ = ~q[6] /*6937*/;
  assign _13710_ = sum_26[9] & q[6] /*6936*/;
  assign _13711_ = m_26[9] & _13709_ /*6935*/;
  assign r_26[9] = _13711_ | _13710_ /*6934*/;
  assign _13712_ = ~q[6] /*6933*/;
  assign _13713_ = sum_26[10] & q[6] /*6932*/;
  assign _13714_ = m_26[10] & _13712_ /*6931*/;
  assign r_26[10] = _13714_ | _13713_ /*6930*/;
  assign _13715_ = ~q[6] /*6929*/;
  assign _13716_ = sum_26[11] & q[6] /*6928*/;
  assign _13717_ = m_26[11] & _13715_ /*6927*/;
  assign r_26[11] = _13717_ | _13716_ /*6926*/;
  assign _13718_ = ~q[6] /*6925*/;
  assign _13719_ = sum_26[12] & q[6] /*6924*/;
  assign _13720_ = m_26[12] & _13718_ /*6923*/;
  assign r_26[12] = _13720_ | _13719_ /*6922*/;
  assign _13721_ = ~q[6] /*6921*/;
  assign _13722_ = sum_26[13] & q[6] /*6920*/;
  assign _13723_ = m_26[13] & _13721_ /*6919*/;
  assign r_26[13] = _13723_ | _13722_ /*6918*/;
  assign _13724_ = ~q[6] /*6917*/;
  assign _13725_ = sum_26[14] & q[6] /*6916*/;
  assign _13726_ = m_26[14] & _13724_ /*6915*/;
  assign r_26[14] = _13726_ | _13725_ /*6914*/;
  assign _13727_ = ~q[6] /*6913*/;
  assign _13728_ = sum_26[15] & q[6] /*6912*/;
  assign _13729_ = m_26[15] & _13727_ /*6911*/;
  assign r_26[15] = _13729_ | _13728_ /*6910*/;
  assign _13730_ = ~q[6] /*6909*/;
  assign _13731_ = sum_26[16] & q[6] /*6908*/;
  assign _13732_ = m_26[16] & _13730_ /*6907*/;
  assign r_26[16] = _13732_ | _13731_ /*6906*/;
  assign _13733_ = ~q[6] /*6905*/;
  assign _13734_ = sum_26[17] & q[6] /*6904*/;
  assign _13735_ = m_26[17] & _13733_ /*6903*/;
  assign r_26[17] = _13735_ | _13734_ /*6902*/;
  assign _13736_ = ~q[6] /*6901*/;
  assign _13737_ = sum_26[18] & q[6] /*6900*/;
  assign _13738_ = m_26[18] & _13736_ /*6899*/;
  assign r_26[18] = _13738_ | _13737_ /*6898*/;
  assign _13739_ = ~q[6] /*6897*/;
  assign _13740_ = sum_26[19] & q[6] /*6896*/;
  assign _13741_ = m_26[19] & _13739_ /*6895*/;
  assign r_26[19] = _13741_ | _13740_ /*6894*/;
  assign _13742_ = ~q[6] /*6893*/;
  assign _13743_ = sum_26[20] & q[6] /*6892*/;
  assign _13744_ = m_26[20] & _13742_ /*6891*/;
  assign r_26[20] = _13744_ | _13743_ /*6890*/;
  assign _13745_ = ~q[6] /*6889*/;
  assign _13746_ = sum_26[21] & q[6] /*6888*/;
  assign _13747_ = m_26[21] & _13745_ /*6887*/;
  assign r_26[21] = _13747_ | _13746_ /*6886*/;
  assign _13748_ = ~q[6] /*6885*/;
  assign _13749_ = sum_26[22] & q[6] /*6884*/;
  assign _13750_ = m_26[22] & _13748_ /*6883*/;
  assign r_26[22] = _13750_ | _13749_ /*6882*/;
  assign _13751_ = ~q[6] /*6881*/;
  assign _13752_ = sum_26[23] & q[6] /*6880*/;
  assign _13753_ = m_26[23] & _13751_ /*6879*/;
  assign r_26[23] = _13753_ | _13752_ /*6878*/;
  assign _13754_ = ~q[6] /*6877*/;
  assign _13755_ = sum_26[24] & q[6] /*6876*/;
  assign _13756_ = m_26[24] & _13754_ /*6875*/;
  assign r_26[24] = _13756_ | _13755_ /*6874*/;
  assign _13757_ = ~q[6] /*6873*/;
  assign _13758_ = sum_26[25] & q[6] /*6872*/;
  assign _13759_ = m_26[25] & _13757_ /*6871*/;
  assign r_26[25] = _13759_ | _13758_ /*6870*/;
  assign _13760_ = ~q[6] /*6869*/;
  assign _13761_ = sum_26[26] & q[6] /*6868*/;
  assign _13762_ = m_26[26] & _13760_ /*6867*/;
  assign r_26[26] = _13762_ | _13761_ /*6866*/;
  assign _13763_ = ~q[6] /*6865*/;
  assign _13764_ = sum_26[27] & q[6] /*6864*/;
  assign _13765_ = m_26[27] & _13763_ /*6863*/;
  assign r_26[27] = _13765_ | _13764_ /*6862*/;
  assign _13766_ = ~q[6] /*6861*/;
  assign _13767_ = sum_26[28] & q[6] /*6860*/;
  assign _13768_ = m_26[28] & _13766_ /*6859*/;
  assign r_26[28] = _13768_ | _13767_ /*6858*/;
  assign _13769_ = ~q[6] /*6857*/;
  assign _13770_ = sum_26[29] & q[6] /*6856*/;
  assign _13771_ = m_26[29] & _13769_ /*6855*/;
  assign r_26[29] = _13771_ | _13770_ /*6854*/;
  assign _13772_ = ~q[6] /*6853*/;
  assign _13773_ = sum_26[30] & q[6] /*6852*/;
  assign _13774_ = m_26[30] & _13772_ /*6851*/;
  assign r_26[30] = _13774_ | _13773_ /*6850*/;
  assign _13775_ = ~q[6] /*6849*/;
  assign _13776_ = sum_26[31] & q[6] /*6848*/;
  assign _13777_ = m_26[31] & _13775_ /*6847*/;
  assign r_26[31] = _13777_ | _13776_ /*6846*/;
  assign _13778_ = ~q[6] /*6845*/;
  assign _13779_ = sum_26[32] & q[6] /*6844*/;
  assign _13780_ = m_26[32] & _13778_ /*6843*/;
  assign r_26[32] = _13780_ | _13779_ /*6842*/;
  assign _13781_ = ~q[6] /*6841*/;
  assign _13782_ = sum_26[33] & q[6] /*6840*/;
  assign _13783_ = m_26[33] & _13781_ /*6839*/;
  assign r_26[33] = _13783_ | _13782_ /*6838*/;
  assign _13784_ = ~q[6] /*6837*/;
  assign _13785_ = sum_26[34] & q[6] /*6836*/;
  assign _13786_ = m_26[34] & _13784_ /*6835*/;
  assign r_26[34] = _13786_ | _13785_ /*6834*/;
  assign _13787_ = ~q[6] /*6833*/;
  assign _13788_ = sum_26[35] & q[6] /*6832*/;
  assign _13789_ = m_26[35] & _13787_ /*6831*/;
  assign r_26[35] = _13789_ | _13788_ /*6830*/;
  assign _13790_ = ~q[6] /*6829*/;
  assign _13791_ = sum_26[36] & q[6] /*6828*/;
  assign _13792_ = m_26[36] & _13790_ /*6827*/;
  assign r_26[36] = _13792_ | _13791_ /*6826*/;
  assign _13793_ = ~q[6] /*6825*/;
  assign _13794_ = sum_26[37] & q[6] /*6824*/;
  assign _13795_ = m_26[37] & _13793_ /*6823*/;
  assign r_26[37] = _13795_ | _13794_ /*6822*/;
  assign _13796_ = ~q[6] /*6821*/;
  assign _13797_ = sum_26[38] & q[6] /*6820*/;
  assign _13798_ = m_26[38] & _13796_ /*6819*/;
  assign r_26[38] = _13798_ | _13797_ /*6818*/;
  assign _13799_ = ~q[6] /*6817*/;
  assign _13800_ = sum_26[39] & q[6] /*6816*/;
  assign _13801_ = m_26[39] & _13799_ /*6815*/;
  assign r_26[39] = _13801_ | _13800_ /*6814*/;
  assign _13802_ = ~q[6] /*6813*/;
  assign _13803_ = sum_26[40] & q[6] /*6812*/;
  assign _13804_ = m_26[40] & _13802_ /*6811*/;
  assign r_26[40] = _13804_ | _13803_ /*6810*/;
  assign _13805_ = ~q[6] /*6809*/;
  assign _13806_ = sum_26[41] & q[6] /*6808*/;
  assign _13807_ = m_26[41] & _13805_ /*6807*/;
  assign r_26[41] = _13807_ | _13806_ /*6806*/;
  assign _13808_ = ~q[6] /*6805*/;
  assign _13809_ = sum_26[42] & q[6] /*6804*/;
  assign _13810_ = m_26[42] & _13808_ /*6803*/;
  assign r_26[42] = _13810_ | _13809_ /*6802*/;
  assign _13811_ = ~q[6] /*6801*/;
  assign _13812_ = sum_26[43] & q[6] /*6800*/;
  assign _13813_ = m_26[43] & _13811_ /*6799*/;
  assign r_26[43] = _13813_ | _13812_ /*6798*/;
  assign _13814_ = ~q[6] /*6797*/;
  assign _13815_ = sum_26[44] & q[6] /*6796*/;
  assign _13816_ = m_26[44] & _13814_ /*6795*/;
  assign r_26[44] = _13816_ | _13815_ /*6794*/;
  assign _13817_ = ~q[6] /*6793*/;
  assign _13818_ = sum_26[45] & q[6] /*6792*/;
  assign _13819_ = m_26[45] & _13817_ /*6791*/;
  assign r_26[45] = _13819_ | _13818_ /*6790*/;
  assign _13820_ = ~q[6] /*6789*/;
  assign _13821_ = sum_26[46] & q[6] /*6788*/;
  assign _13822_ = m_26[46] & _13820_ /*6787*/;
  assign r_26[46] = _13822_ | _13821_ /*6786*/;
  assign _13823_ = ~q[6] /*6785*/;
  assign _13824_ = sum_26[47] & q[6] /*6784*/;
  assign _13825_ = m_26[47] & _13823_ /*6783*/;
  assign r_26[47] = _13825_ | _13824_ /*6782*/;
  assign _13826_ = ~q[6] /*6781*/;
  assign _13827_ = sum_26[48] & q[6] /*6780*/;
  assign _13828_ = m_26[48] & _13826_ /*6779*/;
  assign r_26[48] = _13828_ | _13827_ /*6778*/;
  assign _13829_ = ~q[6] /*6777*/;
  assign _13830_ = sum_26[49] & q[6] /*6776*/;
  assign _13831_ = m_26[49] & _13829_ /*6775*/;
  assign r_26[49] = _13831_ | _13830_ /*6774*/;
  assign _13832_ = ~q[6] /*6773*/;
  assign _13833_ = sum_26[50] & q[6] /*6772*/;
  assign _13834_ = m_26[50] & _13832_ /*6771*/;
  assign r_26[50] = _13834_ | _13833_ /*6770*/;
  assign _13835_ = ~q[6] /*6769*/;
  assign _13836_ = sum_26[51] & q[6] /*6768*/;
  assign _13837_ = m_26[51] & _13835_ /*6767*/;
  assign r_26[51] = _13837_ | _13836_ /*6766*/;
  assign _13838_ = ~q[6] /*6765*/;
  assign _13839_ = sum_26[52] & q[6] /*6764*/;
  assign _13840_ = m_26[52] & _13838_ /*6763*/;
  assign r_26[52] = _13840_ | _13839_ /*6762*/;
  assign _13841_ = ~q[6] /*6761*/;
  assign _13842_ = sum_26[53] & q[6] /*6760*/;
  assign _13843_ = m_26[53] & _13841_ /*6759*/;
  assign r_26[53] = _13843_ | _13842_ /*6758*/;
  assign _13844_ = ~q[6] /*6757*/;
  assign _13845_ = sum_26[54] & q[6] /*6756*/;
  assign _13846_ = m_26[54] & _13844_ /*6755*/;
  assign r_26[54] = _13846_ | _13845_ /*6754*/;
  assign _13847_ = ~q[6] /*6753*/;
  assign _13848_ = sum_26[55] & q[6] /*6752*/;
  assign _13849_ = m_26[55] & _13847_ /*6751*/;
  assign r_26[55] = _13849_ | _13848_ /*6750*/;
  assign _13850_ = ~q[6] /*6749*/;
  assign _13851_ = sum_26[56] & q[6] /*6748*/;
  assign _13852_ = m_26[56] & _13850_ /*6747*/;
  assign r_26[56] = _13852_ | _13851_ /*6746*/;
  assign _13853_ = ~q[6] /*6745*/;
  assign _13854_ = sum_26[57] & q[6] /*6744*/;
  assign _13855_ = m_26[57] & _13853_ /*6743*/;
  assign r_26[57] = _13855_ | _13854_ /*6742*/;
  assign _13856_ = ~q[6] /*6741*/;
  assign _13857_ = sum_26[58] & q[6] /*6740*/;
  assign _13858_ = m_26[58] & _13856_ /*6739*/;
  assign r_26[58] = _13858_ | _13857_ /*6738*/;
  assign _13859_ = ~q[6] /*6737*/;
  assign _13860_ = sum_26[59] & q[6] /*6736*/;
  assign _13861_ = m_26[59] & _13859_ /*6735*/;
  assign r_26[59] = _13861_ | _13860_ /*6734*/;
  assign _13862_ = ~q[6] /*6733*/;
  assign _13863_ = sum_26[60] & q[6] /*6732*/;
  assign _13864_ = m_26[60] & _13862_ /*6731*/;
  assign r_26[60] = _13864_ | _13863_ /*6730*/;
  assign _13865_ = ~q[6] /*6729*/;
  assign _13866_ = sum_26[61] & q[6] /*6728*/;
  assign _13867_ = m_26[61] & _13865_ /*6727*/;
  assign r_26[61] = _13867_ | _13866_ /*6726*/;
  assign _13868_ = ~q[6] /*6725*/;
  assign _13869_ = sum_26[62] & q[6] /*6724*/;
  assign _13870_ = m_26[62] & _13868_ /*6723*/;
  assign r_26[62] = _13870_ | _13869_ /*6722*/;
  assign _13871_ = ~q[6] /*6721*/;
  assign _13872_ = sum_26[63] & q[6] /*6720*/;
  assign _13873_ = m_26[63] & _13871_ /*6719*/;
  assign r_26[63] = _13873_ | _13872_ /*6718*/;
  assign _13874_ = ~q[6] /*6717*/;
  assign _13875_ = sum_26[64] & q[6] /*6716*/;
  assign _13876_ = m_26[64] & _13874_ /*6715*/;
  assign r_26[64] = _13876_ | _13875_ /*6714*/;
  assign _13877_ = ~q[6] /*6713*/;
  assign _13878_ = sum_26[65] & q[6] /*6712*/;
  assign _13879_ = m_26[65] & _13877_ /*6711*/;
  assign r_26[65] = _13879_ | _13878_ /*6710*/;
  assign _13880_ = ~q[6] /*6709*/;
  assign _13881_ = sum_26[66] & q[6] /*6708*/;
  assign _13882_ = m_26[66] & _13880_ /*6707*/;
  assign r_26[66] = _13882_ | _13881_ /*6706*/;
  assign _13883_ = ~q[6] /*6705*/;
  assign _13884_ = sum_26[67] & q[6] /*6704*/;
  assign _13885_ = m_26[67] & _13883_ /*6703*/;
  assign r_26[67] = _13885_ | _13884_ /*6702*/;
  assign _13886_ = ~q[6] /*6701*/;
  assign _13887_ = sum_26[68] & q[6] /*6700*/;
  assign _13888_ = m_26[68] & _13886_ /*6699*/;
  assign r_26[68] = _13888_ | _13887_ /*6698*/;
  assign _13889_ = ~q[6] /*6697*/;
  assign _13890_ = sum_26[69] & q[6] /*6696*/;
  assign _13891_ = m_26[69] & _13889_ /*6695*/;
  assign r_26[69] = _13891_ | _13890_ /*6694*/;
  assign _13892_ = ~q[6] /*6693*/;
  assign _13893_ = sum_26[70] & q[6] /*6692*/;
  assign _13894_ = m_26[70] & _13892_ /*6691*/;
  assign r_26[70] = _13894_ | _13893_ /*6690*/;
  assign _13895_ = ~q[6] /*6689*/;
  assign _13896_ = sum_26[71] & q[6] /*6688*/;
  assign _13897_ = m_26[71] & _13895_ /*6687*/;
  assign r_26[71] = _13897_ | _13896_ /*6686*/;
  assign _13898_ = ~q[6] /*6685*/;
  assign _13899_ = sum_26[72] & q[6] /*6684*/;
  assign _13900_ = m_26[72] & _13898_ /*6683*/;
  assign r_26[72] = _13900_ | _13899_ /*6682*/;
  assign _13901_ = ~q[6] /*6681*/;
  assign _13902_ = sum_26[73] & q[6] /*6680*/;
  assign _13903_ = m_26[73] & _13901_ /*6679*/;
  assign r_26[73] = _13903_ | _13902_ /*6678*/;
  assign _13904_ = ~q[6] /*6677*/;
  assign _13905_ = sum_26[74] & q[6] /*6676*/;
  assign _13906_ = m_26[74] & _13904_ /*6675*/;
  assign r_26[74] = _13906_ | _13905_ /*6674*/;
  assign _13907_ = ~q[6] /*6673*/;
  assign _13908_ = sum_26[75] & q[6] /*6672*/;
  assign _13909_ = m_26[75] & _13907_ /*6671*/;
  assign r_26[75] = _13909_ | _13908_ /*6670*/;
  assign _13910_ = ~q[6] /*6669*/;
  assign _13911_ = sum_26[76] & q[6] /*6668*/;
  assign _13912_ = m_26[76] & _13910_ /*6667*/;
  assign r_26[76] = _13912_ | _13911_ /*6666*/;
  assign _13913_ = ~q[6] /*6665*/;
  assign _13914_ = sum_26[77] & q[6] /*6664*/;
  assign _13915_ = m_26[77] & _13913_ /*6663*/;
  assign r_26[77] = _13915_ | _13914_ /*6662*/;
  assign _13916_ = ~q[6] /*6661*/;
  assign _13917_ = sum_26[78] & q[6] /*6660*/;
  assign _13918_ = m_26[78] & _13916_ /*6659*/;
  assign r_26[78] = _13918_ | _13917_ /*6658*/;
  assign _13919_ = ~q[6] /*6657*/;
  assign _13920_ = sum_26[79] & q[6] /*6656*/;
  assign _13921_ = m_26[79] & _13919_ /*6655*/;
  assign r_26[79] = _13921_ | _13920_ /*6654*/;
  assign _13922_ = ~q[6] /*6653*/;
  assign _13923_ = sum_26[80] & q[6] /*6652*/;
  assign _13924_ = m_26[80] & _13922_ /*6651*/;
  assign r_26[80] = _13924_ | _13923_ /*6650*/;
  assign _13925_ = ~q[6] /*6649*/;
  assign _13926_ = sum_26[81] & q[6] /*6648*/;
  assign _13927_ = m_26[81] & _13925_ /*6647*/;
  assign r_26[81] = _13927_ | _13926_ /*6646*/;
  assign _13928_ = ~q[6] /*6645*/;
  assign _13929_ = sum_26[82] & q[6] /*6644*/;
  assign _13930_ = m_26[82] & _13928_ /*6643*/;
  assign r_26[82] = _13930_ | _13929_ /*6642*/;
  assign _13931_ = ~q[6] /*6641*/;
  assign _13932_ = sum_26[83] & q[6] /*6640*/;
  assign _13933_ = m_26[83] & _13931_ /*6639*/;
  assign r_26[83] = _13933_ | _13932_ /*6638*/;
  assign _13934_ = ~q[6] /*6637*/;
  assign _13935_ = sum_26[84] & q[6] /*6636*/;
  assign _13936_ = m_26[84] & _13934_ /*6635*/;
  assign r_26[84] = _13936_ | _13935_ /*6634*/;
  assign _13937_ = ~q[6] /*6633*/;
  assign _13938_ = sum_26[85] & q[6] /*6632*/;
  assign _13939_ = m_26[85] & _13937_ /*6631*/;
  assign r_26[85] = _13939_ | _13938_ /*6630*/;
  assign _13940_ = ~q[6] /*6629*/;
  assign _13941_ = sum_26[86] & q[6] /*6628*/;
  assign _13942_ = m_26[86] & _13940_ /*6627*/;
  assign r_26[86] = _13942_ | _13941_ /*6626*/;
  assign _13943_ = ~q[6] /*6625*/;
  assign _13944_ = sum_26[87] & q[6] /*6624*/;
  assign _13945_ = m_26[87] & _13943_ /*6623*/;
  assign r_26[87] = _13945_ | _13944_ /*6622*/;
  assign _13946_ = ~q[6] /*6621*/;
  assign _13947_ = sum_26[88] & q[6] /*6620*/;
  assign _13948_ = m_26[88] & _13946_ /*6619*/;
  assign r_26[88] = _13948_ | _13947_ /*6618*/;
  assign inv_27[0] = oneWire /*6520*/;
  assign inv_27[1] = oneWire /*6514*/;
  assign inv_27[2] = oneWire /*6508*/;
  assign inv_27[3] = oneWire /*6502*/;
  assign inv_27[4] = oneWire /*6496*/;
  assign inv_27[5] = ~div[0] /*6490*/;
  assign inv_27[6] = ~div[1] /*6484*/;
  assign inv_27[7] = ~div[2] /*6478*/;
  assign inv_27[8] = ~div[3] /*6472*/;
  assign inv_27[9] = ~div[4] /*6466*/;
  assign inv_27[10] = ~div[5] /*6460*/;
  assign inv_27[11] = ~div[6] /*6454*/;
  assign inv_27[12] = ~div[7] /*6448*/;
  assign inv_27[13] = ~div[8] /*6442*/;
  assign inv_27[14] = ~div[9] /*6436*/;
  assign inv_27[15] = ~div[10] /*6430*/;
  assign inv_27[16] = ~div[11] /*6424*/;
  assign inv_27[17] = ~div[12] /*6418*/;
  assign inv_27[18] = ~div[13] /*6412*/;
  assign inv_27[19] = ~div[14] /*6406*/;
  assign inv_27[20] = ~div[15] /*6400*/;
  assign inv_27[21] = ~div[16] /*6394*/;
  assign inv_27[22] = ~div[17] /*6388*/;
  assign inv_27[23] = ~div[18] /*6382*/;
  assign inv_27[24] = ~div[19] /*6376*/;
  assign inv_27[25] = ~div[20] /*6370*/;
  assign inv_27[26] = ~div[21] /*6364*/;
  assign inv_27[27] = ~div[22] /*6358*/;
  assign inv_27[28] = ~div[23] /*6352*/;
  assign inv_27[29] = ~div[24] /*6346*/;
  assign inv_27[30] = ~div[25] /*6340*/;
  assign inv_27[31] = ~div[26] /*6334*/;
  assign inv_27[32] = ~div[27] /*6328*/;
  assign inv_27[33] = ~div[28] /*6322*/;
  assign inv_27[34] = ~div[29] /*6316*/;
  assign inv_27[35] = ~div[30] /*6310*/;
  assign inv_27[36] = oneWire /*6304*/;
  assign inv_27[37] = oneWire /*6298*/;
  assign inv_27[38] = oneWire /*6292*/;
  assign inv_27[39] = oneWire /*6286*/;
  assign inv_27[40] = oneWire /*6280*/;
  assign inv_27[41] = oneWire /*6274*/;
  assign inv_27[42] = oneWire /*6268*/;
  assign inv_27[43] = oneWire /*6262*/;
  assign inv_27[44] = oneWire /*6256*/;
  assign inv_27[45] = oneWire /*6250*/;
  assign inv_27[46] = oneWire /*6244*/;
  assign inv_27[47] = oneWire /*6238*/;
  assign inv_27[48] = oneWire /*6232*/;
  assign inv_27[49] = oneWire /*6226*/;
  assign inv_27[50] = oneWire /*6220*/;
  assign inv_27[51] = oneWire /*6214*/;
  assign inv_27[52] = oneWire /*6208*/;
  assign inv_27[53] = oneWire /*6202*/;
  assign inv_27[54] = oneWire /*6196*/;
  assign inv_27[55] = oneWire /*6190*/;
  assign inv_27[56] = oneWire /*6184*/;
  assign inv_27[57] = oneWire /*6178*/;
  assign inv_27[58] = oneWire /*6172*/;
  assign inv_27[59] = oneWire /*6166*/;
  assign inv_27[60] = oneWire /*6160*/;
  assign inv_27[61] = oneWire /*6154*/;
  assign inv_27[62] = oneWire /*6148*/;
  assign inv_27[63] = oneWire /*6142*/;
  assign inv_27[64] = oneWire /*6136*/;
  assign inv_27[65] = oneWire /*6130*/;
  assign inv_27[66] = oneWire /*6124*/;
  assign inv_27[67] = oneWire /*6118*/;
  assign inv_27[68] = oneWire /*6112*/;
  assign inv_27[69] = oneWire /*6106*/;
  assign inv_27[70] = oneWire /*6100*/;
  assign inv_27[71] = oneWire /*6094*/;
  assign inv_27[72] = oneWire /*6088*/;
  assign inv_27[73] = oneWire /*6082*/;
  assign inv_27[74] = oneWire /*6076*/;
  assign inv_27[75] = oneWire /*6070*/;
  assign inv_27[76] = oneWire /*6064*/;
  assign inv_27[77] = oneWire /*6058*/;
  assign inv_27[78] = oneWire /*6052*/;
  assign inv_27[79] = oneWire /*6046*/;
  assign inv_27[80] = oneWire /*6040*/;
  assign inv_27[81] = oneWire /*6034*/;
  assign inv_27[82] = oneWire /*6028*/;
  assign inv_27[83] = oneWire /*6022*/;
  assign inv_27[84] = oneWire /*6016*/;
  assign inv_27[85] = oneWire /*6010*/;
  assign inv_27[86] = oneWire /*6004*/;
  assign inv_27[87] = oneWire /*5998*/;
  assign inv_27[88] = oneWire /*5992*/;
  assign _13949_ = inv_27[0] ^ r_26[0] /*6519*/;
  assign sum_27[0] = _13949_ ^ oneWire /*6518*/;
  assign _13950_ = _13949_ & oneWire /*6517*/;
  assign _13951_ = inv_27[0] & r_26[0] /*6516*/;
  assign _13952_ = _13950_ | _13951_ /*6515*/;
  assign _13953_ = inv_27[1] ^ r_26[1] /*6513*/;
  assign sum_27[1] = _13953_ ^ _13952_ /*6512*/;
  assign _13954_ = _13953_ & _13952_ /*6511*/;
  assign _13955_ = inv_27[1] & r_26[1] /*6510*/;
  assign _13956_ = _13954_ | _13955_ /*6509*/;
  assign _13957_ = inv_27[2] ^ r_26[2] /*6507*/;
  assign sum_27[2] = _13957_ ^ _13956_ /*6506*/;
  assign _13958_ = _13957_ & _13956_ /*6505*/;
  assign _13959_ = inv_27[2] & r_26[2] /*6504*/;
  assign _13960_ = _13958_ | _13959_ /*6503*/;
  assign _13961_ = inv_27[3] ^ r_26[3] /*6501*/;
  assign sum_27[3] = _13961_ ^ _13960_ /*6500*/;
  assign _13962_ = _13961_ & _13960_ /*6499*/;
  assign _13963_ = inv_27[3] & r_26[3] /*6498*/;
  assign _13964_ = _13962_ | _13963_ /*6497*/;
  assign _13965_ = inv_27[4] ^ r_26[4] /*6495*/;
  assign sum_27[4] = _13965_ ^ _13964_ /*6494*/;
  assign _13966_ = _13965_ & _13964_ /*6493*/;
  assign _13967_ = inv_27[4] & r_26[4] /*6492*/;
  assign _13968_ = _13966_ | _13967_ /*6491*/;
  assign _13969_ = inv_27[5] ^ r_26[5] /*6489*/;
  assign sum_27[5] = _13969_ ^ _13968_ /*6488*/;
  assign _13970_ = _13969_ & _13968_ /*6487*/;
  assign _13971_ = inv_27[5] & r_26[5] /*6486*/;
  assign _13972_ = _13970_ | _13971_ /*6485*/;
  assign _13973_ = inv_27[6] ^ r_26[6] /*6483*/;
  assign sum_27[6] = _13973_ ^ _13972_ /*6482*/;
  assign _13974_ = _13973_ & _13972_ /*6481*/;
  assign _13975_ = inv_27[6] & r_26[6] /*6480*/;
  assign _13976_ = _13974_ | _13975_ /*6479*/;
  assign _13977_ = inv_27[7] ^ r_26[7] /*6477*/;
  assign sum_27[7] = _13977_ ^ _13976_ /*6476*/;
  assign _13978_ = _13977_ & _13976_ /*6475*/;
  assign _13979_ = inv_27[7] & r_26[7] /*6474*/;
  assign _13980_ = _13978_ | _13979_ /*6473*/;
  assign _13981_ = inv_27[8] ^ r_26[8] /*6471*/;
  assign sum_27[8] = _13981_ ^ _13980_ /*6470*/;
  assign _13982_ = _13981_ & _13980_ /*6469*/;
  assign _13983_ = inv_27[8] & r_26[8] /*6468*/;
  assign _13984_ = _13982_ | _13983_ /*6467*/;
  assign _13985_ = inv_27[9] ^ r_26[9] /*6465*/;
  assign sum_27[9] = _13985_ ^ _13984_ /*6464*/;
  assign _13986_ = _13985_ & _13984_ /*6463*/;
  assign _13987_ = inv_27[9] & r_26[9] /*6462*/;
  assign _13988_ = _13986_ | _13987_ /*6461*/;
  assign _13989_ = inv_27[10] ^ r_26[10] /*6459*/;
  assign sum_27[10] = _13989_ ^ _13988_ /*6458*/;
  assign _13990_ = _13989_ & _13988_ /*6457*/;
  assign _13991_ = inv_27[10] & r_26[10] /*6456*/;
  assign _13992_ = _13990_ | _13991_ /*6455*/;
  assign _13993_ = inv_27[11] ^ r_26[11] /*6453*/;
  assign sum_27[11] = _13993_ ^ _13992_ /*6452*/;
  assign _13994_ = _13993_ & _13992_ /*6451*/;
  assign _13995_ = inv_27[11] & r_26[11] /*6450*/;
  assign _13996_ = _13994_ | _13995_ /*6449*/;
  assign _13997_ = inv_27[12] ^ r_26[12] /*6447*/;
  assign sum_27[12] = _13997_ ^ _13996_ /*6446*/;
  assign _13998_ = _13997_ & _13996_ /*6445*/;
  assign _13999_ = inv_27[12] & r_26[12] /*6444*/;
  assign _14000_ = _13998_ | _13999_ /*6443*/;
  assign _14001_ = inv_27[13] ^ r_26[13] /*6441*/;
  assign sum_27[13] = _14001_ ^ _14000_ /*6440*/;
  assign _14002_ = _14001_ & _14000_ /*6439*/;
  assign _14003_ = inv_27[13] & r_26[13] /*6438*/;
  assign _14004_ = _14002_ | _14003_ /*6437*/;
  assign _14005_ = inv_27[14] ^ r_26[14] /*6435*/;
  assign sum_27[14] = _14005_ ^ _14004_ /*6434*/;
  assign _14006_ = _14005_ & _14004_ /*6433*/;
  assign _14007_ = inv_27[14] & r_26[14] /*6432*/;
  assign _14008_ = _14006_ | _14007_ /*6431*/;
  assign _14009_ = inv_27[15] ^ r_26[15] /*6429*/;
  assign sum_27[15] = _14009_ ^ _14008_ /*6428*/;
  assign _14010_ = _14009_ & _14008_ /*6427*/;
  assign _14011_ = inv_27[15] & r_26[15] /*6426*/;
  assign _14012_ = _14010_ | _14011_ /*6425*/;
  assign _14013_ = inv_27[16] ^ r_26[16] /*6423*/;
  assign sum_27[16] = _14013_ ^ _14012_ /*6422*/;
  assign _14014_ = _14013_ & _14012_ /*6421*/;
  assign _14015_ = inv_27[16] & r_26[16] /*6420*/;
  assign _14016_ = _14014_ | _14015_ /*6419*/;
  assign _14017_ = inv_27[17] ^ r_26[17] /*6417*/;
  assign sum_27[17] = _14017_ ^ _14016_ /*6416*/;
  assign _14018_ = _14017_ & _14016_ /*6415*/;
  assign _14019_ = inv_27[17] & r_26[17] /*6414*/;
  assign _14020_ = _14018_ | _14019_ /*6413*/;
  assign _14021_ = inv_27[18] ^ r_26[18] /*6411*/;
  assign sum_27[18] = _14021_ ^ _14020_ /*6410*/;
  assign _14022_ = _14021_ & _14020_ /*6409*/;
  assign _14023_ = inv_27[18] & r_26[18] /*6408*/;
  assign _14024_ = _14022_ | _14023_ /*6407*/;
  assign _14025_ = inv_27[19] ^ r_26[19] /*6405*/;
  assign sum_27[19] = _14025_ ^ _14024_ /*6404*/;
  assign _14026_ = _14025_ & _14024_ /*6403*/;
  assign _14027_ = inv_27[19] & r_26[19] /*6402*/;
  assign _14028_ = _14026_ | _14027_ /*6401*/;
  assign _14029_ = inv_27[20] ^ r_26[20] /*6399*/;
  assign sum_27[20] = _14029_ ^ _14028_ /*6398*/;
  assign _14030_ = _14029_ & _14028_ /*6397*/;
  assign _14031_ = inv_27[20] & r_26[20] /*6396*/;
  assign _14032_ = _14030_ | _14031_ /*6395*/;
  assign _14033_ = inv_27[21] ^ r_26[21] /*6393*/;
  assign sum_27[21] = _14033_ ^ _14032_ /*6392*/;
  assign _14034_ = _14033_ & _14032_ /*6391*/;
  assign _14035_ = inv_27[21] & r_26[21] /*6390*/;
  assign _14036_ = _14034_ | _14035_ /*6389*/;
  assign _14037_ = inv_27[22] ^ r_26[22] /*6387*/;
  assign sum_27[22] = _14037_ ^ _14036_ /*6386*/;
  assign _14038_ = _14037_ & _14036_ /*6385*/;
  assign _14039_ = inv_27[22] & r_26[22] /*6384*/;
  assign _14040_ = _14038_ | _14039_ /*6383*/;
  assign _14041_ = inv_27[23] ^ r_26[23] /*6381*/;
  assign sum_27[23] = _14041_ ^ _14040_ /*6380*/;
  assign _14042_ = _14041_ & _14040_ /*6379*/;
  assign _14043_ = inv_27[23] & r_26[23] /*6378*/;
  assign _14044_ = _14042_ | _14043_ /*6377*/;
  assign _14045_ = inv_27[24] ^ r_26[24] /*6375*/;
  assign sum_27[24] = _14045_ ^ _14044_ /*6374*/;
  assign _14046_ = _14045_ & _14044_ /*6373*/;
  assign _14047_ = inv_27[24] & r_26[24] /*6372*/;
  assign _14048_ = _14046_ | _14047_ /*6371*/;
  assign _14049_ = inv_27[25] ^ r_26[25] /*6369*/;
  assign sum_27[25] = _14049_ ^ _14048_ /*6368*/;
  assign _14050_ = _14049_ & _14048_ /*6367*/;
  assign _14051_ = inv_27[25] & r_26[25] /*6366*/;
  assign _14052_ = _14050_ | _14051_ /*6365*/;
  assign _14053_ = inv_27[26] ^ r_26[26] /*6363*/;
  assign sum_27[26] = _14053_ ^ _14052_ /*6362*/;
  assign _14054_ = _14053_ & _14052_ /*6361*/;
  assign _14055_ = inv_27[26] & r_26[26] /*6360*/;
  assign _14056_ = _14054_ | _14055_ /*6359*/;
  assign _14057_ = inv_27[27] ^ r_26[27] /*6357*/;
  assign sum_27[27] = _14057_ ^ _14056_ /*6356*/;
  assign _14058_ = _14057_ & _14056_ /*6355*/;
  assign _14059_ = inv_27[27] & r_26[27] /*6354*/;
  assign _14060_ = _14058_ | _14059_ /*6353*/;
  assign _14061_ = inv_27[28] ^ r_26[28] /*6351*/;
  assign sum_27[28] = _14061_ ^ _14060_ /*6350*/;
  assign _14062_ = _14061_ & _14060_ /*6349*/;
  assign _14063_ = inv_27[28] & r_26[28] /*6348*/;
  assign _14064_ = _14062_ | _14063_ /*6347*/;
  assign _14065_ = inv_27[29] ^ r_26[29] /*6345*/;
  assign sum_27[29] = _14065_ ^ _14064_ /*6344*/;
  assign _14066_ = _14065_ & _14064_ /*6343*/;
  assign _14067_ = inv_27[29] & r_26[29] /*6342*/;
  assign _14068_ = _14066_ | _14067_ /*6341*/;
  assign _14069_ = inv_27[30] ^ r_26[30] /*6339*/;
  assign sum_27[30] = _14069_ ^ _14068_ /*6338*/;
  assign _14070_ = _14069_ & _14068_ /*6337*/;
  assign _14071_ = inv_27[30] & r_26[30] /*6336*/;
  assign _14072_ = _14070_ | _14071_ /*6335*/;
  assign _14073_ = inv_27[31] ^ r_26[31] /*6333*/;
  assign sum_27[31] = _14073_ ^ _14072_ /*6332*/;
  assign _14074_ = _14073_ & _14072_ /*6331*/;
  assign _14075_ = inv_27[31] & r_26[31] /*6330*/;
  assign _14076_ = _14074_ | _14075_ /*6329*/;
  assign _14077_ = inv_27[32] ^ r_26[32] /*6327*/;
  assign sum_27[32] = _14077_ ^ _14076_ /*6326*/;
  assign _14078_ = _14077_ & _14076_ /*6325*/;
  assign _14079_ = inv_27[32] & r_26[32] /*6324*/;
  assign _14080_ = _14078_ | _14079_ /*6323*/;
  assign _14081_ = inv_27[33] ^ r_26[33] /*6321*/;
  assign sum_27[33] = _14081_ ^ _14080_ /*6320*/;
  assign _14082_ = _14081_ & _14080_ /*6319*/;
  assign _14083_ = inv_27[33] & r_26[33] /*6318*/;
  assign _14084_ = _14082_ | _14083_ /*6317*/;
  assign _14085_ = inv_27[34] ^ r_26[34] /*6315*/;
  assign sum_27[34] = _14085_ ^ _14084_ /*6314*/;
  assign _14086_ = _14085_ & _14084_ /*6313*/;
  assign _14087_ = inv_27[34] & r_26[34] /*6312*/;
  assign _14088_ = _14086_ | _14087_ /*6311*/;
  assign _14089_ = inv_27[35] ^ r_26[35] /*6309*/;
  assign sum_27[35] = _14089_ ^ _14088_ /*6308*/;
  assign _14090_ = _14089_ & _14088_ /*6307*/;
  assign _14091_ = inv_27[35] & r_26[35] /*6306*/;
  assign _14092_ = _14090_ | _14091_ /*6305*/;
  assign _14093_ = inv_27[36] ^ r_26[36] /*6303*/;
  assign sum_27[36] = _14093_ ^ _14092_ /*6302*/;
  assign _14094_ = _14093_ & _14092_ /*6301*/;
  assign _14095_ = inv_27[36] & r_26[36] /*6300*/;
  assign _14096_ = _14094_ | _14095_ /*6299*/;
  assign _14097_ = inv_27[37] ^ r_26[37] /*6297*/;
  assign sum_27[37] = _14097_ ^ _14096_ /*6296*/;
  assign _14098_ = _14097_ & _14096_ /*6295*/;
  assign _14099_ = inv_27[37] & r_26[37] /*6294*/;
  assign _14100_ = _14098_ | _14099_ /*6293*/;
  assign _14101_ = inv_27[38] ^ r_26[38] /*6291*/;
  assign sum_27[38] = _14101_ ^ _14100_ /*6290*/;
  assign _14102_ = _14101_ & _14100_ /*6289*/;
  assign _14103_ = inv_27[38] & r_26[38] /*6288*/;
  assign _14104_ = _14102_ | _14103_ /*6287*/;
  assign _14105_ = inv_27[39] ^ r_26[39] /*6285*/;
  assign sum_27[39] = _14105_ ^ _14104_ /*6284*/;
  assign _14106_ = _14105_ & _14104_ /*6283*/;
  assign _14107_ = inv_27[39] & r_26[39] /*6282*/;
  assign _14108_ = _14106_ | _14107_ /*6281*/;
  assign _14109_ = inv_27[40] ^ r_26[40] /*6279*/;
  assign sum_27[40] = _14109_ ^ _14108_ /*6278*/;
  assign _14110_ = _14109_ & _14108_ /*6277*/;
  assign _14111_ = inv_27[40] & r_26[40] /*6276*/;
  assign _14112_ = _14110_ | _14111_ /*6275*/;
  assign _14113_ = inv_27[41] ^ r_26[41] /*6273*/;
  assign sum_27[41] = _14113_ ^ _14112_ /*6272*/;
  assign _14114_ = _14113_ & _14112_ /*6271*/;
  assign _14115_ = inv_27[41] & r_26[41] /*6270*/;
  assign _14116_ = _14114_ | _14115_ /*6269*/;
  assign _14117_ = inv_27[42] ^ r_26[42] /*6267*/;
  assign sum_27[42] = _14117_ ^ _14116_ /*6266*/;
  assign _14118_ = _14117_ & _14116_ /*6265*/;
  assign _14119_ = inv_27[42] & r_26[42] /*6264*/;
  assign _14120_ = _14118_ | _14119_ /*6263*/;
  assign _14121_ = inv_27[43] ^ r_26[43] /*6261*/;
  assign sum_27[43] = _14121_ ^ _14120_ /*6260*/;
  assign _14122_ = _14121_ & _14120_ /*6259*/;
  assign _14123_ = inv_27[43] & r_26[43] /*6258*/;
  assign _14124_ = _14122_ | _14123_ /*6257*/;
  assign _14125_ = inv_27[44] ^ r_26[44] /*6255*/;
  assign sum_27[44] = _14125_ ^ _14124_ /*6254*/;
  assign _14126_ = _14125_ & _14124_ /*6253*/;
  assign _14127_ = inv_27[44] & r_26[44] /*6252*/;
  assign _14128_ = _14126_ | _14127_ /*6251*/;
  assign _14129_ = inv_27[45] ^ r_26[45] /*6249*/;
  assign sum_27[45] = _14129_ ^ _14128_ /*6248*/;
  assign _14130_ = _14129_ & _14128_ /*6247*/;
  assign _14131_ = inv_27[45] & r_26[45] /*6246*/;
  assign _14132_ = _14130_ | _14131_ /*6245*/;
  assign _14133_ = inv_27[46] ^ r_26[46] /*6243*/;
  assign sum_27[46] = _14133_ ^ _14132_ /*6242*/;
  assign _14134_ = _14133_ & _14132_ /*6241*/;
  assign _14135_ = inv_27[46] & r_26[46] /*6240*/;
  assign _14136_ = _14134_ | _14135_ /*6239*/;
  assign _14137_ = inv_27[47] ^ r_26[47] /*6237*/;
  assign sum_27[47] = _14137_ ^ _14136_ /*6236*/;
  assign _14138_ = _14137_ & _14136_ /*6235*/;
  assign _14139_ = inv_27[47] & r_26[47] /*6234*/;
  assign _14140_ = _14138_ | _14139_ /*6233*/;
  assign _14141_ = inv_27[48] ^ r_26[48] /*6231*/;
  assign sum_27[48] = _14141_ ^ _14140_ /*6230*/;
  assign _14142_ = _14141_ & _14140_ /*6229*/;
  assign _14143_ = inv_27[48] & r_26[48] /*6228*/;
  assign _14144_ = _14142_ | _14143_ /*6227*/;
  assign _14145_ = inv_27[49] ^ r_26[49] /*6225*/;
  assign sum_27[49] = _14145_ ^ _14144_ /*6224*/;
  assign _14146_ = _14145_ & _14144_ /*6223*/;
  assign _14147_ = inv_27[49] & r_26[49] /*6222*/;
  assign _14148_ = _14146_ | _14147_ /*6221*/;
  assign _14149_ = inv_27[50] ^ r_26[50] /*6219*/;
  assign sum_27[50] = _14149_ ^ _14148_ /*6218*/;
  assign _14150_ = _14149_ & _14148_ /*6217*/;
  assign _14151_ = inv_27[50] & r_26[50] /*6216*/;
  assign _14152_ = _14150_ | _14151_ /*6215*/;
  assign _14153_ = inv_27[51] ^ r_26[51] /*6213*/;
  assign sum_27[51] = _14153_ ^ _14152_ /*6212*/;
  assign _14154_ = _14153_ & _14152_ /*6211*/;
  assign _14155_ = inv_27[51] & r_26[51] /*6210*/;
  assign _14156_ = _14154_ | _14155_ /*6209*/;
  assign _14157_ = inv_27[52] ^ r_26[52] /*6207*/;
  assign sum_27[52] = _14157_ ^ _14156_ /*6206*/;
  assign _14158_ = _14157_ & _14156_ /*6205*/;
  assign _14159_ = inv_27[52] & r_26[52] /*6204*/;
  assign _14160_ = _14158_ | _14159_ /*6203*/;
  assign _14161_ = inv_27[53] ^ r_26[53] /*6201*/;
  assign sum_27[53] = _14161_ ^ _14160_ /*6200*/;
  assign _14162_ = _14161_ & _14160_ /*6199*/;
  assign _14163_ = inv_27[53] & r_26[53] /*6198*/;
  assign _14164_ = _14162_ | _14163_ /*6197*/;
  assign _14165_ = inv_27[54] ^ r_26[54] /*6195*/;
  assign sum_27[54] = _14165_ ^ _14164_ /*6194*/;
  assign _14166_ = _14165_ & _14164_ /*6193*/;
  assign _14167_ = inv_27[54] & r_26[54] /*6192*/;
  assign _14168_ = _14166_ | _14167_ /*6191*/;
  assign _14169_ = inv_27[55] ^ r_26[55] /*6189*/;
  assign sum_27[55] = _14169_ ^ _14168_ /*6188*/;
  assign _14170_ = _14169_ & _14168_ /*6187*/;
  assign _14171_ = inv_27[55] & r_26[55] /*6186*/;
  assign _14172_ = _14170_ | _14171_ /*6185*/;
  assign _14173_ = inv_27[56] ^ r_26[56] /*6183*/;
  assign sum_27[56] = _14173_ ^ _14172_ /*6182*/;
  assign _14174_ = _14173_ & _14172_ /*6181*/;
  assign _14175_ = inv_27[56] & r_26[56] /*6180*/;
  assign _14176_ = _14174_ | _14175_ /*6179*/;
  assign _14177_ = inv_27[57] ^ r_26[57] /*6177*/;
  assign sum_27[57] = _14177_ ^ _14176_ /*6176*/;
  assign _14178_ = _14177_ & _14176_ /*6175*/;
  assign _14179_ = inv_27[57] & r_26[57] /*6174*/;
  assign _14180_ = _14178_ | _14179_ /*6173*/;
  assign _14181_ = inv_27[58] ^ r_26[58] /*6171*/;
  assign sum_27[58] = _14181_ ^ _14180_ /*6170*/;
  assign _14182_ = _14181_ & _14180_ /*6169*/;
  assign _14183_ = inv_27[58] & r_26[58] /*6168*/;
  assign _14184_ = _14182_ | _14183_ /*6167*/;
  assign _14185_ = inv_27[59] ^ r_26[59] /*6165*/;
  assign sum_27[59] = _14185_ ^ _14184_ /*6164*/;
  assign _14186_ = _14185_ & _14184_ /*6163*/;
  assign _14187_ = inv_27[59] & r_26[59] /*6162*/;
  assign _14188_ = _14186_ | _14187_ /*6161*/;
  assign _14189_ = inv_27[60] ^ r_26[60] /*6159*/;
  assign sum_27[60] = _14189_ ^ _14188_ /*6158*/;
  assign _14190_ = _14189_ & _14188_ /*6157*/;
  assign _14191_ = inv_27[60] & r_26[60] /*6156*/;
  assign _14192_ = _14190_ | _14191_ /*6155*/;
  assign _14193_ = inv_27[61] ^ r_26[61] /*6153*/;
  assign sum_27[61] = _14193_ ^ _14192_ /*6152*/;
  assign _14194_ = _14193_ & _14192_ /*6151*/;
  assign _14195_ = inv_27[61] & r_26[61] /*6150*/;
  assign _14196_ = _14194_ | _14195_ /*6149*/;
  assign _14197_ = inv_27[62] ^ r_26[62] /*6147*/;
  assign sum_27[62] = _14197_ ^ _14196_ /*6146*/;
  assign _14198_ = _14197_ & _14196_ /*6145*/;
  assign _14199_ = inv_27[62] & r_26[62] /*6144*/;
  assign _14200_ = _14198_ | _14199_ /*6143*/;
  assign _14201_ = inv_27[63] ^ r_26[63] /*6141*/;
  assign sum_27[63] = _14201_ ^ _14200_ /*6140*/;
  assign _14202_ = _14201_ & _14200_ /*6139*/;
  assign _14203_ = inv_27[63] & r_26[63] /*6138*/;
  assign _14204_ = _14202_ | _14203_ /*6137*/;
  assign _14205_ = inv_27[64] ^ r_26[64] /*6135*/;
  assign sum_27[64] = _14205_ ^ _14204_ /*6134*/;
  assign _14206_ = _14205_ & _14204_ /*6133*/;
  assign _14207_ = inv_27[64] & r_26[64] /*6132*/;
  assign _14208_ = _14206_ | _14207_ /*6131*/;
  assign _14209_ = inv_27[65] ^ r_26[65] /*6129*/;
  assign sum_27[65] = _14209_ ^ _14208_ /*6128*/;
  assign _14210_ = _14209_ & _14208_ /*6127*/;
  assign _14211_ = inv_27[65] & r_26[65] /*6126*/;
  assign _14212_ = _14210_ | _14211_ /*6125*/;
  assign _14213_ = inv_27[66] ^ r_26[66] /*6123*/;
  assign sum_27[66] = _14213_ ^ _14212_ /*6122*/;
  assign _14214_ = _14213_ & _14212_ /*6121*/;
  assign _14215_ = inv_27[66] & r_26[66] /*6120*/;
  assign _14216_ = _14214_ | _14215_ /*6119*/;
  assign _14217_ = inv_27[67] ^ r_26[67] /*6117*/;
  assign sum_27[67] = _14217_ ^ _14216_ /*6116*/;
  assign _14218_ = _14217_ & _14216_ /*6115*/;
  assign _14219_ = inv_27[67] & r_26[67] /*6114*/;
  assign _14220_ = _14218_ | _14219_ /*6113*/;
  assign _14221_ = inv_27[68] ^ r_26[68] /*6111*/;
  assign sum_27[68] = _14221_ ^ _14220_ /*6110*/;
  assign _14222_ = _14221_ & _14220_ /*6109*/;
  assign _14223_ = inv_27[68] & r_26[68] /*6108*/;
  assign _14224_ = _14222_ | _14223_ /*6107*/;
  assign _14225_ = inv_27[69] ^ r_26[69] /*6105*/;
  assign sum_27[69] = _14225_ ^ _14224_ /*6104*/;
  assign _14226_ = _14225_ & _14224_ /*6103*/;
  assign _14227_ = inv_27[69] & r_26[69] /*6102*/;
  assign _14228_ = _14226_ | _14227_ /*6101*/;
  assign _14229_ = inv_27[70] ^ r_26[70] /*6099*/;
  assign sum_27[70] = _14229_ ^ _14228_ /*6098*/;
  assign _14230_ = _14229_ & _14228_ /*6097*/;
  assign _14231_ = inv_27[70] & r_26[70] /*6096*/;
  assign _14232_ = _14230_ | _14231_ /*6095*/;
  assign _14233_ = inv_27[71] ^ r_26[71] /*6093*/;
  assign sum_27[71] = _14233_ ^ _14232_ /*6092*/;
  assign _14234_ = _14233_ & _14232_ /*6091*/;
  assign _14235_ = inv_27[71] & r_26[71] /*6090*/;
  assign _14236_ = _14234_ | _14235_ /*6089*/;
  assign _14237_ = inv_27[72] ^ r_26[72] /*6087*/;
  assign sum_27[72] = _14237_ ^ _14236_ /*6086*/;
  assign _14238_ = _14237_ & _14236_ /*6085*/;
  assign _14239_ = inv_27[72] & r_26[72] /*6084*/;
  assign _14240_ = _14238_ | _14239_ /*6083*/;
  assign _14241_ = inv_27[73] ^ r_26[73] /*6081*/;
  assign sum_27[73] = _14241_ ^ _14240_ /*6080*/;
  assign _14242_ = _14241_ & _14240_ /*6079*/;
  assign _14243_ = inv_27[73] & r_26[73] /*6078*/;
  assign _14244_ = _14242_ | _14243_ /*6077*/;
  assign _14245_ = inv_27[74] ^ r_26[74] /*6075*/;
  assign sum_27[74] = _14245_ ^ _14244_ /*6074*/;
  assign _14246_ = _14245_ & _14244_ /*6073*/;
  assign _14247_ = inv_27[74] & r_26[74] /*6072*/;
  assign _14248_ = _14246_ | _14247_ /*6071*/;
  assign _14249_ = inv_27[75] ^ r_26[75] /*6069*/;
  assign sum_27[75] = _14249_ ^ _14248_ /*6068*/;
  assign _14250_ = _14249_ & _14248_ /*6067*/;
  assign _14251_ = inv_27[75] & r_26[75] /*6066*/;
  assign _14252_ = _14250_ | _14251_ /*6065*/;
  assign _14253_ = inv_27[76] ^ r_26[76] /*6063*/;
  assign sum_27[76] = _14253_ ^ _14252_ /*6062*/;
  assign _14254_ = _14253_ & _14252_ /*6061*/;
  assign _14255_ = inv_27[76] & r_26[76] /*6060*/;
  assign _14256_ = _14254_ | _14255_ /*6059*/;
  assign _14257_ = inv_27[77] ^ r_26[77] /*6057*/;
  assign sum_27[77] = _14257_ ^ _14256_ /*6056*/;
  assign _14258_ = _14257_ & _14256_ /*6055*/;
  assign _14259_ = inv_27[77] & r_26[77] /*6054*/;
  assign _14260_ = _14258_ | _14259_ /*6053*/;
  assign _14261_ = inv_27[78] ^ r_26[78] /*6051*/;
  assign sum_27[78] = _14261_ ^ _14260_ /*6050*/;
  assign _14262_ = _14261_ & _14260_ /*6049*/;
  assign _14263_ = inv_27[78] & r_26[78] /*6048*/;
  assign _14264_ = _14262_ | _14263_ /*6047*/;
  assign _14265_ = inv_27[79] ^ r_26[79] /*6045*/;
  assign sum_27[79] = _14265_ ^ _14264_ /*6044*/;
  assign _14266_ = _14265_ & _14264_ /*6043*/;
  assign _14267_ = inv_27[79] & r_26[79] /*6042*/;
  assign _14268_ = _14266_ | _14267_ /*6041*/;
  assign _14269_ = inv_27[80] ^ r_26[80] /*6039*/;
  assign sum_27[80] = _14269_ ^ _14268_ /*6038*/;
  assign _14270_ = _14269_ & _14268_ /*6037*/;
  assign _14271_ = inv_27[80] & r_26[80] /*6036*/;
  assign _14272_ = _14270_ | _14271_ /*6035*/;
  assign _14273_ = inv_27[81] ^ r_26[81] /*6033*/;
  assign sum_27[81] = _14273_ ^ _14272_ /*6032*/;
  assign _14274_ = _14273_ & _14272_ /*6031*/;
  assign _14275_ = inv_27[81] & r_26[81] /*6030*/;
  assign _14276_ = _14274_ | _14275_ /*6029*/;
  assign _14277_ = inv_27[82] ^ r_26[82] /*6027*/;
  assign sum_27[82] = _14277_ ^ _14276_ /*6026*/;
  assign _14278_ = _14277_ & _14276_ /*6025*/;
  assign _14279_ = inv_27[82] & r_26[82] /*6024*/;
  assign _14280_ = _14278_ | _14279_ /*6023*/;
  assign _14281_ = inv_27[83] ^ r_26[83] /*6021*/;
  assign sum_27[83] = _14281_ ^ _14280_ /*6020*/;
  assign _14282_ = _14281_ & _14280_ /*6019*/;
  assign _14283_ = inv_27[83] & r_26[83] /*6018*/;
  assign _14284_ = _14282_ | _14283_ /*6017*/;
  assign _14285_ = inv_27[84] ^ r_26[84] /*6015*/;
  assign sum_27[84] = _14285_ ^ _14284_ /*6014*/;
  assign _14286_ = _14285_ & _14284_ /*6013*/;
  assign _14287_ = inv_27[84] & r_26[84] /*6012*/;
  assign _14288_ = _14286_ | _14287_ /*6011*/;
  assign _14289_ = inv_27[85] ^ r_26[85] /*6009*/;
  assign sum_27[85] = _14289_ ^ _14288_ /*6008*/;
  assign _14290_ = _14289_ & _14288_ /*6007*/;
  assign _14291_ = inv_27[85] & r_26[85] /*6006*/;
  assign _14292_ = _14290_ | _14291_ /*6005*/;
  assign _14293_ = inv_27[86] ^ r_26[86] /*6003*/;
  assign sum_27[86] = _14293_ ^ _14292_ /*6002*/;
  assign _14294_ = _14293_ & _14292_ /*6001*/;
  assign _14295_ = inv_27[86] & r_26[86] /*6000*/;
  assign _14296_ = _14294_ | _14295_ /*5999*/;
  assign _14297_ = inv_27[87] ^ r_26[87] /*5997*/;
  assign sum_27[87] = _14297_ ^ _14296_ /*5996*/;
  assign _14298_ = _14297_ & _14296_ /*5995*/;
  assign _14299_ = inv_27[87] & r_26[87] /*5994*/;
  assign _14300_ = _14298_ | _14299_ /*5993*/;
  assign _14301_ = inv_27[88] ^ r_26[88] /*5991*/;
  assign sum_27[88] = _14301_ ^ _14300_ /*5990*/;
  assign _14302_ = _14301_ & _14300_ /*5989*/;
  assign _14303_ = inv_27[88] & r_26[88] /*5988*/;
  assign _14304_ = _14302_ | _14303_ /*5987*/;
  assign _14305_ = _14304_ ^ _14300_ /*5986*/;
  assign _14306_ = ~_14305_ /*5985*/;
  assign _14307_ = sum_27[88] & _14306_ /*5984*/;
  assign _14308_ = _14305_ & _14304_ /*5983*/;
  assign sum_27[89] = _14308_ | _14307_ /*5982*/;
  assign q[5] = ~sum_27[89] /*5981*/;
  assign m_27[0] = r_26[0] /*5980*/;
  assign m_27[1] = r_26[1] /*5979*/;
  assign m_27[2] = r_26[2] /*5978*/;
  assign m_27[3] = r_26[3] /*5977*/;
  assign m_27[4] = r_26[4] /*5976*/;
  assign m_27[5] = r_26[5] /*5975*/;
  assign m_27[6] = r_26[6] /*5974*/;
  assign m_27[7] = r_26[7] /*5973*/;
  assign m_27[8] = r_26[8] /*5972*/;
  assign m_27[9] = r_26[9] /*5971*/;
  assign m_27[10] = r_26[10] /*5970*/;
  assign m_27[11] = r_26[11] /*5969*/;
  assign m_27[12] = r_26[12] /*5968*/;
  assign m_27[13] = r_26[13] /*5967*/;
  assign m_27[14] = r_26[14] /*5966*/;
  assign m_27[15] = r_26[15] /*5965*/;
  assign m_27[16] = r_26[16] /*5964*/;
  assign m_27[17] = r_26[17] /*5963*/;
  assign m_27[18] = r_26[18] /*5962*/;
  assign m_27[19] = r_26[19] /*5961*/;
  assign m_27[20] = r_26[20] /*5960*/;
  assign m_27[21] = r_26[21] /*5959*/;
  assign m_27[22] = r_26[22] /*5958*/;
  assign m_27[23] = r_26[23] /*5957*/;
  assign m_27[24] = r_26[24] /*5956*/;
  assign m_27[25] = r_26[25] /*5955*/;
  assign m_27[26] = r_26[26] /*5954*/;
  assign m_27[27] = r_26[27] /*5953*/;
  assign m_27[28] = r_26[28] /*5952*/;
  assign m_27[29] = r_26[29] /*5951*/;
  assign m_27[30] = r_26[30] /*5950*/;
  assign m_27[31] = r_26[31] /*5949*/;
  assign m_27[32] = r_26[32] /*5948*/;
  assign m_27[33] = r_26[33] /*5947*/;
  assign m_27[34] = r_26[34] /*5946*/;
  assign m_27[35] = r_26[35] /*5945*/;
  assign m_27[36] = r_26[36] /*5944*/;
  assign m_27[37] = r_26[37] /*5943*/;
  assign m_27[38] = r_26[38] /*5942*/;
  assign m_27[39] = r_26[39] /*5941*/;
  assign m_27[40] = r_26[40] /*5940*/;
  assign m_27[41] = r_26[41] /*5939*/;
  assign m_27[42] = r_26[42] /*5938*/;
  assign m_27[43] = r_26[43] /*5937*/;
  assign m_27[44] = r_26[44] /*5936*/;
  assign m_27[45] = r_26[45] /*5935*/;
  assign m_27[46] = r_26[46] /*5934*/;
  assign m_27[47] = r_26[47] /*5933*/;
  assign m_27[48] = r_26[48] /*5932*/;
  assign m_27[49] = r_26[49] /*5931*/;
  assign m_27[50] = r_26[50] /*5930*/;
  assign m_27[51] = r_26[51] /*5929*/;
  assign m_27[52] = r_26[52] /*5928*/;
  assign m_27[53] = r_26[53] /*5927*/;
  assign m_27[54] = r_26[54] /*5926*/;
  assign m_27[55] = r_26[55] /*5925*/;
  assign m_27[56] = r_26[56] /*5924*/;
  assign m_27[57] = r_26[57] /*5923*/;
  assign m_27[58] = r_26[58] /*5922*/;
  assign m_27[59] = r_26[59] /*5921*/;
  assign m_27[60] = r_26[60] /*5920*/;
  assign m_27[61] = r_26[61] /*5919*/;
  assign m_27[62] = r_26[62] /*5918*/;
  assign m_27[63] = r_26[63] /*5917*/;
  assign m_27[64] = r_26[64] /*5916*/;
  assign m_27[65] = r_26[65] /*5915*/;
  assign m_27[66] = r_26[66] /*5914*/;
  assign m_27[67] = r_26[67] /*5913*/;
  assign m_27[68] = r_26[68] /*5912*/;
  assign m_27[69] = r_26[69] /*5911*/;
  assign m_27[70] = r_26[70] /*5910*/;
  assign m_27[71] = r_26[71] /*5909*/;
  assign m_27[72] = r_26[72] /*5908*/;
  assign m_27[73] = r_26[73] /*5907*/;
  assign m_27[74] = r_26[74] /*5906*/;
  assign m_27[75] = r_26[75] /*5905*/;
  assign m_27[76] = r_26[76] /*5904*/;
  assign m_27[77] = r_26[77] /*5903*/;
  assign m_27[78] = r_26[78] /*5902*/;
  assign m_27[79] = r_26[79] /*5901*/;
  assign m_27[80] = r_26[80] /*5900*/;
  assign m_27[81] = r_26[81] /*5899*/;
  assign m_27[82] = r_26[82] /*5898*/;
  assign m_27[83] = r_26[83] /*5897*/;
  assign m_27[84] = r_26[84] /*5896*/;
  assign m_27[85] = r_26[85] /*5895*/;
  assign m_27[86] = r_26[86] /*5894*/;
  assign m_27[87] = r_26[87] /*5893*/;
  assign m_27[88] = r_26[88] /*5892*/;
  assign m_27[89] = r_26[88] /*5891*/;
  assign _14310_ = ~q[5] /*5890*/;
  assign _14311_ = sum_27[0] & q[5] /*5889*/;
  assign _14312_ = m_27[0] & _14310_ /*5888*/;
  assign r_27[0] = _14312_ | _14311_ /*5887*/;
  assign _14313_ = ~q[5] /*5886*/;
  assign _14314_ = sum_27[1] & q[5] /*5885*/;
  assign _14315_ = m_27[1] & _14313_ /*5884*/;
  assign r_27[1] = _14315_ | _14314_ /*5883*/;
  assign _14316_ = ~q[5] /*5882*/;
  assign _14317_ = sum_27[2] & q[5] /*5881*/;
  assign _14318_ = m_27[2] & _14316_ /*5880*/;
  assign r_27[2] = _14318_ | _14317_ /*5879*/;
  assign _14319_ = ~q[5] /*5878*/;
  assign _14320_ = sum_27[3] & q[5] /*5877*/;
  assign _14321_ = m_27[3] & _14319_ /*5876*/;
  assign r_27[3] = _14321_ | _14320_ /*5875*/;
  assign _14322_ = ~q[5] /*5874*/;
  assign _14323_ = sum_27[4] & q[5] /*5873*/;
  assign _14324_ = m_27[4] & _14322_ /*5872*/;
  assign r_27[4] = _14324_ | _14323_ /*5871*/;
  assign _14325_ = ~q[5] /*5870*/;
  assign _14326_ = sum_27[5] & q[5] /*5869*/;
  assign _14327_ = m_27[5] & _14325_ /*5868*/;
  assign r_27[5] = _14327_ | _14326_ /*5867*/;
  assign _14328_ = ~q[5] /*5866*/;
  assign _14329_ = sum_27[6] & q[5] /*5865*/;
  assign _14330_ = m_27[6] & _14328_ /*5864*/;
  assign r_27[6] = _14330_ | _14329_ /*5863*/;
  assign _14331_ = ~q[5] /*5862*/;
  assign _14332_ = sum_27[7] & q[5] /*5861*/;
  assign _14333_ = m_27[7] & _14331_ /*5860*/;
  assign r_27[7] = _14333_ | _14332_ /*5859*/;
  assign _14334_ = ~q[5] /*5858*/;
  assign _14335_ = sum_27[8] & q[5] /*5857*/;
  assign _14336_ = m_27[8] & _14334_ /*5856*/;
  assign r_27[8] = _14336_ | _14335_ /*5855*/;
  assign _14337_ = ~q[5] /*5854*/;
  assign _14338_ = sum_27[9] & q[5] /*5853*/;
  assign _14339_ = m_27[9] & _14337_ /*5852*/;
  assign r_27[9] = _14339_ | _14338_ /*5851*/;
  assign _14340_ = ~q[5] /*5850*/;
  assign _14341_ = sum_27[10] & q[5] /*5849*/;
  assign _14342_ = m_27[10] & _14340_ /*5848*/;
  assign r_27[10] = _14342_ | _14341_ /*5847*/;
  assign _14343_ = ~q[5] /*5846*/;
  assign _14344_ = sum_27[11] & q[5] /*5845*/;
  assign _14345_ = m_27[11] & _14343_ /*5844*/;
  assign r_27[11] = _14345_ | _14344_ /*5843*/;
  assign _14346_ = ~q[5] /*5842*/;
  assign _14347_ = sum_27[12] & q[5] /*5841*/;
  assign _14348_ = m_27[12] & _14346_ /*5840*/;
  assign r_27[12] = _14348_ | _14347_ /*5839*/;
  assign _14349_ = ~q[5] /*5838*/;
  assign _14350_ = sum_27[13] & q[5] /*5837*/;
  assign _14351_ = m_27[13] & _14349_ /*5836*/;
  assign r_27[13] = _14351_ | _14350_ /*5835*/;
  assign _14352_ = ~q[5] /*5834*/;
  assign _14353_ = sum_27[14] & q[5] /*5833*/;
  assign _14354_ = m_27[14] & _14352_ /*5832*/;
  assign r_27[14] = _14354_ | _14353_ /*5831*/;
  assign _14355_ = ~q[5] /*5830*/;
  assign _14356_ = sum_27[15] & q[5] /*5829*/;
  assign _14357_ = m_27[15] & _14355_ /*5828*/;
  assign r_27[15] = _14357_ | _14356_ /*5827*/;
  assign _14358_ = ~q[5] /*5826*/;
  assign _14359_ = sum_27[16] & q[5] /*5825*/;
  assign _14360_ = m_27[16] & _14358_ /*5824*/;
  assign r_27[16] = _14360_ | _14359_ /*5823*/;
  assign _14361_ = ~q[5] /*5822*/;
  assign _14362_ = sum_27[17] & q[5] /*5821*/;
  assign _14363_ = m_27[17] & _14361_ /*5820*/;
  assign r_27[17] = _14363_ | _14362_ /*5819*/;
  assign _14364_ = ~q[5] /*5818*/;
  assign _14365_ = sum_27[18] & q[5] /*5817*/;
  assign _14366_ = m_27[18] & _14364_ /*5816*/;
  assign r_27[18] = _14366_ | _14365_ /*5815*/;
  assign _14367_ = ~q[5] /*5814*/;
  assign _14368_ = sum_27[19] & q[5] /*5813*/;
  assign _14369_ = m_27[19] & _14367_ /*5812*/;
  assign r_27[19] = _14369_ | _14368_ /*5811*/;
  assign _14370_ = ~q[5] /*5810*/;
  assign _14371_ = sum_27[20] & q[5] /*5809*/;
  assign _14372_ = m_27[20] & _14370_ /*5808*/;
  assign r_27[20] = _14372_ | _14371_ /*5807*/;
  assign _14373_ = ~q[5] /*5806*/;
  assign _14374_ = sum_27[21] & q[5] /*5805*/;
  assign _14375_ = m_27[21] & _14373_ /*5804*/;
  assign r_27[21] = _14375_ | _14374_ /*5803*/;
  assign _14376_ = ~q[5] /*5802*/;
  assign _14377_ = sum_27[22] & q[5] /*5801*/;
  assign _14378_ = m_27[22] & _14376_ /*5800*/;
  assign r_27[22] = _14378_ | _14377_ /*5799*/;
  assign _14379_ = ~q[5] /*5798*/;
  assign _14380_ = sum_27[23] & q[5] /*5797*/;
  assign _14381_ = m_27[23] & _14379_ /*5796*/;
  assign r_27[23] = _14381_ | _14380_ /*5795*/;
  assign _14382_ = ~q[5] /*5794*/;
  assign _14383_ = sum_27[24] & q[5] /*5793*/;
  assign _14384_ = m_27[24] & _14382_ /*5792*/;
  assign r_27[24] = _14384_ | _14383_ /*5791*/;
  assign _14385_ = ~q[5] /*5790*/;
  assign _14386_ = sum_27[25] & q[5] /*5789*/;
  assign _14387_ = m_27[25] & _14385_ /*5788*/;
  assign r_27[25] = _14387_ | _14386_ /*5787*/;
  assign _14388_ = ~q[5] /*5786*/;
  assign _14389_ = sum_27[26] & q[5] /*5785*/;
  assign _14390_ = m_27[26] & _14388_ /*5784*/;
  assign r_27[26] = _14390_ | _14389_ /*5783*/;
  assign _14391_ = ~q[5] /*5782*/;
  assign _14392_ = sum_27[27] & q[5] /*5781*/;
  assign _14393_ = m_27[27] & _14391_ /*5780*/;
  assign r_27[27] = _14393_ | _14392_ /*5779*/;
  assign _14394_ = ~q[5] /*5778*/;
  assign _14395_ = sum_27[28] & q[5] /*5777*/;
  assign _14396_ = m_27[28] & _14394_ /*5776*/;
  assign r_27[28] = _14396_ | _14395_ /*5775*/;
  assign _14397_ = ~q[5] /*5774*/;
  assign _14398_ = sum_27[29] & q[5] /*5773*/;
  assign _14399_ = m_27[29] & _14397_ /*5772*/;
  assign r_27[29] = _14399_ | _14398_ /*5771*/;
  assign _14400_ = ~q[5] /*5770*/;
  assign _14401_ = sum_27[30] & q[5] /*5769*/;
  assign _14402_ = m_27[30] & _14400_ /*5768*/;
  assign r_27[30] = _14402_ | _14401_ /*5767*/;
  assign _14403_ = ~q[5] /*5766*/;
  assign _14404_ = sum_27[31] & q[5] /*5765*/;
  assign _14405_ = m_27[31] & _14403_ /*5764*/;
  assign r_27[31] = _14405_ | _14404_ /*5763*/;
  assign _14406_ = ~q[5] /*5762*/;
  assign _14407_ = sum_27[32] & q[5] /*5761*/;
  assign _14408_ = m_27[32] & _14406_ /*5760*/;
  assign r_27[32] = _14408_ | _14407_ /*5759*/;
  assign _14409_ = ~q[5] /*5758*/;
  assign _14410_ = sum_27[33] & q[5] /*5757*/;
  assign _14411_ = m_27[33] & _14409_ /*5756*/;
  assign r_27[33] = _14411_ | _14410_ /*5755*/;
  assign _14412_ = ~q[5] /*5754*/;
  assign _14413_ = sum_27[34] & q[5] /*5753*/;
  assign _14414_ = m_27[34] & _14412_ /*5752*/;
  assign r_27[34] = _14414_ | _14413_ /*5751*/;
  assign _14415_ = ~q[5] /*5750*/;
  assign _14416_ = sum_27[35] & q[5] /*5749*/;
  assign _14417_ = m_27[35] & _14415_ /*5748*/;
  assign r_27[35] = _14417_ | _14416_ /*5747*/;
  assign _14418_ = ~q[5] /*5746*/;
  assign _14419_ = sum_27[36] & q[5] /*5745*/;
  assign _14420_ = m_27[36] & _14418_ /*5744*/;
  assign r_27[36] = _14420_ | _14419_ /*5743*/;
  assign _14421_ = ~q[5] /*5742*/;
  assign _14422_ = sum_27[37] & q[5] /*5741*/;
  assign _14423_ = m_27[37] & _14421_ /*5740*/;
  assign r_27[37] = _14423_ | _14422_ /*5739*/;
  assign _14424_ = ~q[5] /*5738*/;
  assign _14425_ = sum_27[38] & q[5] /*5737*/;
  assign _14426_ = m_27[38] & _14424_ /*5736*/;
  assign r_27[38] = _14426_ | _14425_ /*5735*/;
  assign _14427_ = ~q[5] /*5734*/;
  assign _14428_ = sum_27[39] & q[5] /*5733*/;
  assign _14429_ = m_27[39] & _14427_ /*5732*/;
  assign r_27[39] = _14429_ | _14428_ /*5731*/;
  assign _14430_ = ~q[5] /*5730*/;
  assign _14431_ = sum_27[40] & q[5] /*5729*/;
  assign _14432_ = m_27[40] & _14430_ /*5728*/;
  assign r_27[40] = _14432_ | _14431_ /*5727*/;
  assign _14433_ = ~q[5] /*5726*/;
  assign _14434_ = sum_27[41] & q[5] /*5725*/;
  assign _14435_ = m_27[41] & _14433_ /*5724*/;
  assign r_27[41] = _14435_ | _14434_ /*5723*/;
  assign _14436_ = ~q[5] /*5722*/;
  assign _14437_ = sum_27[42] & q[5] /*5721*/;
  assign _14438_ = m_27[42] & _14436_ /*5720*/;
  assign r_27[42] = _14438_ | _14437_ /*5719*/;
  assign _14439_ = ~q[5] /*5718*/;
  assign _14440_ = sum_27[43] & q[5] /*5717*/;
  assign _14441_ = m_27[43] & _14439_ /*5716*/;
  assign r_27[43] = _14441_ | _14440_ /*5715*/;
  assign _14442_ = ~q[5] /*5714*/;
  assign _14443_ = sum_27[44] & q[5] /*5713*/;
  assign _14444_ = m_27[44] & _14442_ /*5712*/;
  assign r_27[44] = _14444_ | _14443_ /*5711*/;
  assign _14445_ = ~q[5] /*5710*/;
  assign _14446_ = sum_27[45] & q[5] /*5709*/;
  assign _14447_ = m_27[45] & _14445_ /*5708*/;
  assign r_27[45] = _14447_ | _14446_ /*5707*/;
  assign _14448_ = ~q[5] /*5706*/;
  assign _14449_ = sum_27[46] & q[5] /*5705*/;
  assign _14450_ = m_27[46] & _14448_ /*5704*/;
  assign r_27[46] = _14450_ | _14449_ /*5703*/;
  assign _14451_ = ~q[5] /*5702*/;
  assign _14452_ = sum_27[47] & q[5] /*5701*/;
  assign _14453_ = m_27[47] & _14451_ /*5700*/;
  assign r_27[47] = _14453_ | _14452_ /*5699*/;
  assign _14454_ = ~q[5] /*5698*/;
  assign _14455_ = sum_27[48] & q[5] /*5697*/;
  assign _14456_ = m_27[48] & _14454_ /*5696*/;
  assign r_27[48] = _14456_ | _14455_ /*5695*/;
  assign _14457_ = ~q[5] /*5694*/;
  assign _14458_ = sum_27[49] & q[5] /*5693*/;
  assign _14459_ = m_27[49] & _14457_ /*5692*/;
  assign r_27[49] = _14459_ | _14458_ /*5691*/;
  assign _14460_ = ~q[5] /*5690*/;
  assign _14461_ = sum_27[50] & q[5] /*5689*/;
  assign _14462_ = m_27[50] & _14460_ /*5688*/;
  assign r_27[50] = _14462_ | _14461_ /*5687*/;
  assign _14463_ = ~q[5] /*5686*/;
  assign _14464_ = sum_27[51] & q[5] /*5685*/;
  assign _14465_ = m_27[51] & _14463_ /*5684*/;
  assign r_27[51] = _14465_ | _14464_ /*5683*/;
  assign _14466_ = ~q[5] /*5682*/;
  assign _14467_ = sum_27[52] & q[5] /*5681*/;
  assign _14468_ = m_27[52] & _14466_ /*5680*/;
  assign r_27[52] = _14468_ | _14467_ /*5679*/;
  assign _14469_ = ~q[5] /*5678*/;
  assign _14470_ = sum_27[53] & q[5] /*5677*/;
  assign _14471_ = m_27[53] & _14469_ /*5676*/;
  assign r_27[53] = _14471_ | _14470_ /*5675*/;
  assign _14472_ = ~q[5] /*5674*/;
  assign _14473_ = sum_27[54] & q[5] /*5673*/;
  assign _14474_ = m_27[54] & _14472_ /*5672*/;
  assign r_27[54] = _14474_ | _14473_ /*5671*/;
  assign _14475_ = ~q[5] /*5670*/;
  assign _14476_ = sum_27[55] & q[5] /*5669*/;
  assign _14477_ = m_27[55] & _14475_ /*5668*/;
  assign r_27[55] = _14477_ | _14476_ /*5667*/;
  assign _14478_ = ~q[5] /*5666*/;
  assign _14479_ = sum_27[56] & q[5] /*5665*/;
  assign _14480_ = m_27[56] & _14478_ /*5664*/;
  assign r_27[56] = _14480_ | _14479_ /*5663*/;
  assign _14481_ = ~q[5] /*5662*/;
  assign _14482_ = sum_27[57] & q[5] /*5661*/;
  assign _14483_ = m_27[57] & _14481_ /*5660*/;
  assign r_27[57] = _14483_ | _14482_ /*5659*/;
  assign _14484_ = ~q[5] /*5658*/;
  assign _14485_ = sum_27[58] & q[5] /*5657*/;
  assign _14486_ = m_27[58] & _14484_ /*5656*/;
  assign r_27[58] = _14486_ | _14485_ /*5655*/;
  assign _14487_ = ~q[5] /*5654*/;
  assign _14488_ = sum_27[59] & q[5] /*5653*/;
  assign _14489_ = m_27[59] & _14487_ /*5652*/;
  assign r_27[59] = _14489_ | _14488_ /*5651*/;
  assign _14490_ = ~q[5] /*5650*/;
  assign _14491_ = sum_27[60] & q[5] /*5649*/;
  assign _14492_ = m_27[60] & _14490_ /*5648*/;
  assign r_27[60] = _14492_ | _14491_ /*5647*/;
  assign _14493_ = ~q[5] /*5646*/;
  assign _14494_ = sum_27[61] & q[5] /*5645*/;
  assign _14495_ = m_27[61] & _14493_ /*5644*/;
  assign r_27[61] = _14495_ | _14494_ /*5643*/;
  assign _14496_ = ~q[5] /*5642*/;
  assign _14497_ = sum_27[62] & q[5] /*5641*/;
  assign _14498_ = m_27[62] & _14496_ /*5640*/;
  assign r_27[62] = _14498_ | _14497_ /*5639*/;
  assign _14499_ = ~q[5] /*5638*/;
  assign _14500_ = sum_27[63] & q[5] /*5637*/;
  assign _14501_ = m_27[63] & _14499_ /*5636*/;
  assign r_27[63] = _14501_ | _14500_ /*5635*/;
  assign _14502_ = ~q[5] /*5634*/;
  assign _14503_ = sum_27[64] & q[5] /*5633*/;
  assign _14504_ = m_27[64] & _14502_ /*5632*/;
  assign r_27[64] = _14504_ | _14503_ /*5631*/;
  assign _14505_ = ~q[5] /*5630*/;
  assign _14506_ = sum_27[65] & q[5] /*5629*/;
  assign _14507_ = m_27[65] & _14505_ /*5628*/;
  assign r_27[65] = _14507_ | _14506_ /*5627*/;
  assign _14508_ = ~q[5] /*5626*/;
  assign _14509_ = sum_27[66] & q[5] /*5625*/;
  assign _14510_ = m_27[66] & _14508_ /*5624*/;
  assign r_27[66] = _14510_ | _14509_ /*5623*/;
  assign _14511_ = ~q[5] /*5622*/;
  assign _14512_ = sum_27[67] & q[5] /*5621*/;
  assign _14513_ = m_27[67] & _14511_ /*5620*/;
  assign r_27[67] = _14513_ | _14512_ /*5619*/;
  assign _14514_ = ~q[5] /*5618*/;
  assign _14515_ = sum_27[68] & q[5] /*5617*/;
  assign _14516_ = m_27[68] & _14514_ /*5616*/;
  assign r_27[68] = _14516_ | _14515_ /*5615*/;
  assign _14517_ = ~q[5] /*5614*/;
  assign _14518_ = sum_27[69] & q[5] /*5613*/;
  assign _14519_ = m_27[69] & _14517_ /*5612*/;
  assign r_27[69] = _14519_ | _14518_ /*5611*/;
  assign _14520_ = ~q[5] /*5610*/;
  assign _14521_ = sum_27[70] & q[5] /*5609*/;
  assign _14522_ = m_27[70] & _14520_ /*5608*/;
  assign r_27[70] = _14522_ | _14521_ /*5607*/;
  assign _14523_ = ~q[5] /*5606*/;
  assign _14524_ = sum_27[71] & q[5] /*5605*/;
  assign _14525_ = m_27[71] & _14523_ /*5604*/;
  assign r_27[71] = _14525_ | _14524_ /*5603*/;
  assign _14526_ = ~q[5] /*5602*/;
  assign _14527_ = sum_27[72] & q[5] /*5601*/;
  assign _14528_ = m_27[72] & _14526_ /*5600*/;
  assign r_27[72] = _14528_ | _14527_ /*5599*/;
  assign _14529_ = ~q[5] /*5598*/;
  assign _14530_ = sum_27[73] & q[5] /*5597*/;
  assign _14531_ = m_27[73] & _14529_ /*5596*/;
  assign r_27[73] = _14531_ | _14530_ /*5595*/;
  assign _14532_ = ~q[5] /*5594*/;
  assign _14533_ = sum_27[74] & q[5] /*5593*/;
  assign _14534_ = m_27[74] & _14532_ /*5592*/;
  assign r_27[74] = _14534_ | _14533_ /*5591*/;
  assign _14535_ = ~q[5] /*5590*/;
  assign _14536_ = sum_27[75] & q[5] /*5589*/;
  assign _14537_ = m_27[75] & _14535_ /*5588*/;
  assign r_27[75] = _14537_ | _14536_ /*5587*/;
  assign _14538_ = ~q[5] /*5586*/;
  assign _14539_ = sum_27[76] & q[5] /*5585*/;
  assign _14540_ = m_27[76] & _14538_ /*5584*/;
  assign r_27[76] = _14540_ | _14539_ /*5583*/;
  assign _14541_ = ~q[5] /*5582*/;
  assign _14542_ = sum_27[77] & q[5] /*5581*/;
  assign _14543_ = m_27[77] & _14541_ /*5580*/;
  assign r_27[77] = _14543_ | _14542_ /*5579*/;
  assign _14544_ = ~q[5] /*5578*/;
  assign _14545_ = sum_27[78] & q[5] /*5577*/;
  assign _14546_ = m_27[78] & _14544_ /*5576*/;
  assign r_27[78] = _14546_ | _14545_ /*5575*/;
  assign _14547_ = ~q[5] /*5574*/;
  assign _14548_ = sum_27[79] & q[5] /*5573*/;
  assign _14549_ = m_27[79] & _14547_ /*5572*/;
  assign r_27[79] = _14549_ | _14548_ /*5571*/;
  assign _14550_ = ~q[5] /*5570*/;
  assign _14551_ = sum_27[80] & q[5] /*5569*/;
  assign _14552_ = m_27[80] & _14550_ /*5568*/;
  assign r_27[80] = _14552_ | _14551_ /*5567*/;
  assign _14553_ = ~q[5] /*5566*/;
  assign _14554_ = sum_27[81] & q[5] /*5565*/;
  assign _14555_ = m_27[81] & _14553_ /*5564*/;
  assign r_27[81] = _14555_ | _14554_ /*5563*/;
  assign _14556_ = ~q[5] /*5562*/;
  assign _14557_ = sum_27[82] & q[5] /*5561*/;
  assign _14558_ = m_27[82] & _14556_ /*5560*/;
  assign r_27[82] = _14558_ | _14557_ /*5559*/;
  assign _14559_ = ~q[5] /*5558*/;
  assign _14560_ = sum_27[83] & q[5] /*5557*/;
  assign _14561_ = m_27[83] & _14559_ /*5556*/;
  assign r_27[83] = _14561_ | _14560_ /*5555*/;
  assign _14562_ = ~q[5] /*5554*/;
  assign _14563_ = sum_27[84] & q[5] /*5553*/;
  assign _14564_ = m_27[84] & _14562_ /*5552*/;
  assign r_27[84] = _14564_ | _14563_ /*5551*/;
  assign _14565_ = ~q[5] /*5550*/;
  assign _14566_ = sum_27[85] & q[5] /*5549*/;
  assign _14567_ = m_27[85] & _14565_ /*5548*/;
  assign r_27[85] = _14567_ | _14566_ /*5547*/;
  assign _14568_ = ~q[5] /*5546*/;
  assign _14569_ = sum_27[86] & q[5] /*5545*/;
  assign _14570_ = m_27[86] & _14568_ /*5544*/;
  assign r_27[86] = _14570_ | _14569_ /*5543*/;
  assign _14571_ = ~q[5] /*5542*/;
  assign _14572_ = sum_27[87] & q[5] /*5541*/;
  assign _14573_ = m_27[87] & _14571_ /*5540*/;
  assign r_27[87] = _14573_ | _14572_ /*5539*/;
  assign _14574_ = ~q[5] /*5538*/;
  assign _14575_ = sum_27[88] & q[5] /*5537*/;
  assign _14576_ = m_27[88] & _14574_ /*5536*/;
  assign r_27[88] = _14576_ | _14575_ /*5535*/;
  assign _14577_ = ~q[5] /*5534*/;
  assign _14578_ = sum_27[89] & q[5] /*5533*/;
  assign _14579_ = m_27[89] & _14577_ /*5532*/;
  assign r_27[89] = _14579_ | _14578_ /*5531*/;
  assign inv_28[0] = oneWire /*5444*/;
  assign inv_28[1] = oneWire /*5438*/;
  assign inv_28[2] = oneWire /*5432*/;
  assign inv_28[3] = oneWire /*5426*/;
  assign inv_28[4] = ~div[0] /*5420*/;
  assign inv_28[5] = ~div[1] /*5414*/;
  assign inv_28[6] = ~div[2] /*5408*/;
  assign inv_28[7] = ~div[3] /*5402*/;
  assign inv_28[8] = ~div[4] /*5396*/;
  assign inv_28[9] = ~div[5] /*5390*/;
  assign inv_28[10] = ~div[6] /*5384*/;
  assign inv_28[11] = ~div[7] /*5378*/;
  assign inv_28[12] = ~div[8] /*5372*/;
  assign inv_28[13] = ~div[9] /*5366*/;
  assign inv_28[14] = ~div[10] /*5360*/;
  assign inv_28[15] = ~div[11] /*5354*/;
  assign inv_28[16] = ~div[12] /*5348*/;
  assign inv_28[17] = ~div[13] /*5342*/;
  assign inv_28[18] = ~div[14] /*5336*/;
  assign inv_28[19] = ~div[15] /*5330*/;
  assign inv_28[20] = ~div[16] /*5324*/;
  assign inv_28[21] = ~div[17] /*5318*/;
  assign inv_28[22] = ~div[18] /*5312*/;
  assign inv_28[23] = ~div[19] /*5306*/;
  assign inv_28[24] = ~div[20] /*5300*/;
  assign inv_28[25] = ~div[21] /*5294*/;
  assign inv_28[26] = ~div[22] /*5288*/;
  assign inv_28[27] = ~div[23] /*5282*/;
  assign inv_28[28] = ~div[24] /*5276*/;
  assign inv_28[29] = ~div[25] /*5270*/;
  assign inv_28[30] = ~div[26] /*5264*/;
  assign inv_28[31] = ~div[27] /*5258*/;
  assign inv_28[32] = ~div[28] /*5252*/;
  assign inv_28[33] = ~div[29] /*5246*/;
  assign inv_28[34] = ~div[30] /*5240*/;
  assign inv_28[35] = oneWire /*5234*/;
  assign inv_28[36] = oneWire /*5228*/;
  assign inv_28[37] = oneWire /*5222*/;
  assign inv_28[38] = oneWire /*5216*/;
  assign inv_28[39] = oneWire /*5210*/;
  assign inv_28[40] = oneWire /*5204*/;
  assign inv_28[41] = oneWire /*5198*/;
  assign inv_28[42] = oneWire /*5192*/;
  assign inv_28[43] = oneWire /*5186*/;
  assign inv_28[44] = oneWire /*5180*/;
  assign inv_28[45] = oneWire /*5174*/;
  assign inv_28[46] = oneWire /*5168*/;
  assign inv_28[47] = oneWire /*5162*/;
  assign inv_28[48] = oneWire /*5156*/;
  assign inv_28[49] = oneWire /*5150*/;
  assign inv_28[50] = oneWire /*5144*/;
  assign inv_28[51] = oneWire /*5138*/;
  assign inv_28[52] = oneWire /*5132*/;
  assign inv_28[53] = oneWire /*5126*/;
  assign inv_28[54] = oneWire /*5120*/;
  assign inv_28[55] = oneWire /*5114*/;
  assign inv_28[56] = oneWire /*5108*/;
  assign inv_28[57] = oneWire /*5102*/;
  assign inv_28[58] = oneWire /*5096*/;
  assign inv_28[59] = oneWire /*5090*/;
  assign inv_28[60] = oneWire /*5084*/;
  assign inv_28[61] = oneWire /*5078*/;
  assign inv_28[62] = oneWire /*5072*/;
  assign inv_28[63] = oneWire /*5066*/;
  assign inv_28[64] = oneWire /*5060*/;
  assign inv_28[65] = oneWire /*5054*/;
  assign inv_28[66] = oneWire /*5048*/;
  assign inv_28[67] = oneWire /*5042*/;
  assign inv_28[68] = oneWire /*5036*/;
  assign inv_28[69] = oneWire /*5030*/;
  assign inv_28[70] = oneWire /*5024*/;
  assign inv_28[71] = oneWire /*5018*/;
  assign inv_28[72] = oneWire /*5012*/;
  assign inv_28[73] = oneWire /*5006*/;
  assign inv_28[74] = oneWire /*5000*/;
  assign inv_28[75] = oneWire /*4994*/;
  assign inv_28[76] = oneWire /*4988*/;
  assign inv_28[77] = oneWire /*4982*/;
  assign inv_28[78] = oneWire /*4976*/;
  assign inv_28[79] = oneWire /*4970*/;
  assign inv_28[80] = oneWire /*4964*/;
  assign inv_28[81] = oneWire /*4958*/;
  assign inv_28[82] = oneWire /*4952*/;
  assign inv_28[83] = oneWire /*4946*/;
  assign inv_28[84] = oneWire /*4940*/;
  assign inv_28[85] = oneWire /*4934*/;
  assign inv_28[86] = oneWire /*4928*/;
  assign inv_28[87] = oneWire /*4922*/;
  assign inv_28[88] = oneWire /*4916*/;
  assign inv_28[89] = oneWire /*4910*/;
  assign _14580_ = inv_28[0] ^ r_27[0] /*5443*/;
  assign sum_28[0] = _14580_ ^ oneWire /*5442*/;
  assign _14581_ = _14580_ & oneWire /*5441*/;
  assign _14582_ = inv_28[0] & r_27[0] /*5440*/;
  assign _14583_ = _14581_ | _14582_ /*5439*/;
  assign _14584_ = inv_28[1] ^ r_27[1] /*5437*/;
  assign sum_28[1] = _14584_ ^ _14583_ /*5436*/;
  assign _14585_ = _14584_ & _14583_ /*5435*/;
  assign _14586_ = inv_28[1] & r_27[1] /*5434*/;
  assign _14587_ = _14585_ | _14586_ /*5433*/;
  assign _14588_ = inv_28[2] ^ r_27[2] /*5431*/;
  assign sum_28[2] = _14588_ ^ _14587_ /*5430*/;
  assign _14589_ = _14588_ & _14587_ /*5429*/;
  assign _14590_ = inv_28[2] & r_27[2] /*5428*/;
  assign _14591_ = _14589_ | _14590_ /*5427*/;
  assign _14592_ = inv_28[3] ^ r_27[3] /*5425*/;
  assign sum_28[3] = _14592_ ^ _14591_ /*5424*/;
  assign _14593_ = _14592_ & _14591_ /*5423*/;
  assign _14594_ = inv_28[3] & r_27[3] /*5422*/;
  assign _14595_ = _14593_ | _14594_ /*5421*/;
  assign _14596_ = inv_28[4] ^ r_27[4] /*5419*/;
  assign sum_28[4] = _14596_ ^ _14595_ /*5418*/;
  assign _14597_ = _14596_ & _14595_ /*5417*/;
  assign _14598_ = inv_28[4] & r_27[4] /*5416*/;
  assign _14599_ = _14597_ | _14598_ /*5415*/;
  assign _14600_ = inv_28[5] ^ r_27[5] /*5413*/;
  assign sum_28[5] = _14600_ ^ _14599_ /*5412*/;
  assign _14601_ = _14600_ & _14599_ /*5411*/;
  assign _14602_ = inv_28[5] & r_27[5] /*5410*/;
  assign _14603_ = _14601_ | _14602_ /*5409*/;
  assign _14604_ = inv_28[6] ^ r_27[6] /*5407*/;
  assign sum_28[6] = _14604_ ^ _14603_ /*5406*/;
  assign _14605_ = _14604_ & _14603_ /*5405*/;
  assign _14606_ = inv_28[6] & r_27[6] /*5404*/;
  assign _14607_ = _14605_ | _14606_ /*5403*/;
  assign _14608_ = inv_28[7] ^ r_27[7] /*5401*/;
  assign sum_28[7] = _14608_ ^ _14607_ /*5400*/;
  assign _14609_ = _14608_ & _14607_ /*5399*/;
  assign _14610_ = inv_28[7] & r_27[7] /*5398*/;
  assign _14611_ = _14609_ | _14610_ /*5397*/;
  assign _14612_ = inv_28[8] ^ r_27[8] /*5395*/;
  assign sum_28[8] = _14612_ ^ _14611_ /*5394*/;
  assign _14613_ = _14612_ & _14611_ /*5393*/;
  assign _14614_ = inv_28[8] & r_27[8] /*5392*/;
  assign _14615_ = _14613_ | _14614_ /*5391*/;
  assign _14616_ = inv_28[9] ^ r_27[9] /*5389*/;
  assign sum_28[9] = _14616_ ^ _14615_ /*5388*/;
  assign _14617_ = _14616_ & _14615_ /*5387*/;
  assign _14618_ = inv_28[9] & r_27[9] /*5386*/;
  assign _14619_ = _14617_ | _14618_ /*5385*/;
  assign _14620_ = inv_28[10] ^ r_27[10] /*5383*/;
  assign sum_28[10] = _14620_ ^ _14619_ /*5382*/;
  assign _14621_ = _14620_ & _14619_ /*5381*/;
  assign _14622_ = inv_28[10] & r_27[10] /*5380*/;
  assign _14623_ = _14621_ | _14622_ /*5379*/;
  assign _14624_ = inv_28[11] ^ r_27[11] /*5377*/;
  assign sum_28[11] = _14624_ ^ _14623_ /*5376*/;
  assign _14625_ = _14624_ & _14623_ /*5375*/;
  assign _14626_ = inv_28[11] & r_27[11] /*5374*/;
  assign _14627_ = _14625_ | _14626_ /*5373*/;
  assign _14628_ = inv_28[12] ^ r_27[12] /*5371*/;
  assign sum_28[12] = _14628_ ^ _14627_ /*5370*/;
  assign _14629_ = _14628_ & _14627_ /*5369*/;
  assign _14630_ = inv_28[12] & r_27[12] /*5368*/;
  assign _14631_ = _14629_ | _14630_ /*5367*/;
  assign _14632_ = inv_28[13] ^ r_27[13] /*5365*/;
  assign sum_28[13] = _14632_ ^ _14631_ /*5364*/;
  assign _14633_ = _14632_ & _14631_ /*5363*/;
  assign _14634_ = inv_28[13] & r_27[13] /*5362*/;
  assign _14635_ = _14633_ | _14634_ /*5361*/;
  assign _14636_ = inv_28[14] ^ r_27[14] /*5359*/;
  assign sum_28[14] = _14636_ ^ _14635_ /*5358*/;
  assign _14637_ = _14636_ & _14635_ /*5357*/;
  assign _14638_ = inv_28[14] & r_27[14] /*5356*/;
  assign _14639_ = _14637_ | _14638_ /*5355*/;
  assign _14640_ = inv_28[15] ^ r_27[15] /*5353*/;
  assign sum_28[15] = _14640_ ^ _14639_ /*5352*/;
  assign _14641_ = _14640_ & _14639_ /*5351*/;
  assign _14642_ = inv_28[15] & r_27[15] /*5350*/;
  assign _14643_ = _14641_ | _14642_ /*5349*/;
  assign _14644_ = inv_28[16] ^ r_27[16] /*5347*/;
  assign sum_28[16] = _14644_ ^ _14643_ /*5346*/;
  assign _14645_ = _14644_ & _14643_ /*5345*/;
  assign _14646_ = inv_28[16] & r_27[16] /*5344*/;
  assign _14647_ = _14645_ | _14646_ /*5343*/;
  assign _14648_ = inv_28[17] ^ r_27[17] /*5341*/;
  assign sum_28[17] = _14648_ ^ _14647_ /*5340*/;
  assign _14649_ = _14648_ & _14647_ /*5339*/;
  assign _14650_ = inv_28[17] & r_27[17] /*5338*/;
  assign _14651_ = _14649_ | _14650_ /*5337*/;
  assign _14652_ = inv_28[18] ^ r_27[18] /*5335*/;
  assign sum_28[18] = _14652_ ^ _14651_ /*5334*/;
  assign _14653_ = _14652_ & _14651_ /*5333*/;
  assign _14654_ = inv_28[18] & r_27[18] /*5332*/;
  assign _14655_ = _14653_ | _14654_ /*5331*/;
  assign _14656_ = inv_28[19] ^ r_27[19] /*5329*/;
  assign sum_28[19] = _14656_ ^ _14655_ /*5328*/;
  assign _14657_ = _14656_ & _14655_ /*5327*/;
  assign _14658_ = inv_28[19] & r_27[19] /*5326*/;
  assign _14659_ = _14657_ | _14658_ /*5325*/;
  assign _14660_ = inv_28[20] ^ r_27[20] /*5323*/;
  assign sum_28[20] = _14660_ ^ _14659_ /*5322*/;
  assign _14661_ = _14660_ & _14659_ /*5321*/;
  assign _14662_ = inv_28[20] & r_27[20] /*5320*/;
  assign _14663_ = _14661_ | _14662_ /*5319*/;
  assign _14664_ = inv_28[21] ^ r_27[21] /*5317*/;
  assign sum_28[21] = _14664_ ^ _14663_ /*5316*/;
  assign _14665_ = _14664_ & _14663_ /*5315*/;
  assign _14666_ = inv_28[21] & r_27[21] /*5314*/;
  assign _14667_ = _14665_ | _14666_ /*5313*/;
  assign _14668_ = inv_28[22] ^ r_27[22] /*5311*/;
  assign sum_28[22] = _14668_ ^ _14667_ /*5310*/;
  assign _14669_ = _14668_ & _14667_ /*5309*/;
  assign _14670_ = inv_28[22] & r_27[22] /*5308*/;
  assign _14671_ = _14669_ | _14670_ /*5307*/;
  assign _14672_ = inv_28[23] ^ r_27[23] /*5305*/;
  assign sum_28[23] = _14672_ ^ _14671_ /*5304*/;
  assign _14673_ = _14672_ & _14671_ /*5303*/;
  assign _14674_ = inv_28[23] & r_27[23] /*5302*/;
  assign _14675_ = _14673_ | _14674_ /*5301*/;
  assign _14676_ = inv_28[24] ^ r_27[24] /*5299*/;
  assign sum_28[24] = _14676_ ^ _14675_ /*5298*/;
  assign _14677_ = _14676_ & _14675_ /*5297*/;
  assign _14678_ = inv_28[24] & r_27[24] /*5296*/;
  assign _14679_ = _14677_ | _14678_ /*5295*/;
  assign _14680_ = inv_28[25] ^ r_27[25] /*5293*/;
  assign sum_28[25] = _14680_ ^ _14679_ /*5292*/;
  assign _14681_ = _14680_ & _14679_ /*5291*/;
  assign _14682_ = inv_28[25] & r_27[25] /*5290*/;
  assign _14683_ = _14681_ | _14682_ /*5289*/;
  assign _14684_ = inv_28[26] ^ r_27[26] /*5287*/;
  assign sum_28[26] = _14684_ ^ _14683_ /*5286*/;
  assign _14685_ = _14684_ & _14683_ /*5285*/;
  assign _14686_ = inv_28[26] & r_27[26] /*5284*/;
  assign _14687_ = _14685_ | _14686_ /*5283*/;
  assign _14688_ = inv_28[27] ^ r_27[27] /*5281*/;
  assign sum_28[27] = _14688_ ^ _14687_ /*5280*/;
  assign _14689_ = _14688_ & _14687_ /*5279*/;
  assign _14690_ = inv_28[27] & r_27[27] /*5278*/;
  assign _14691_ = _14689_ | _14690_ /*5277*/;
  assign _14692_ = inv_28[28] ^ r_27[28] /*5275*/;
  assign sum_28[28] = _14692_ ^ _14691_ /*5274*/;
  assign _14693_ = _14692_ & _14691_ /*5273*/;
  assign _14694_ = inv_28[28] & r_27[28] /*5272*/;
  assign _14695_ = _14693_ | _14694_ /*5271*/;
  assign _14696_ = inv_28[29] ^ r_27[29] /*5269*/;
  assign sum_28[29] = _14696_ ^ _14695_ /*5268*/;
  assign _14697_ = _14696_ & _14695_ /*5267*/;
  assign _14698_ = inv_28[29] & r_27[29] /*5266*/;
  assign _14699_ = _14697_ | _14698_ /*5265*/;
  assign _14700_ = inv_28[30] ^ r_27[30] /*5263*/;
  assign sum_28[30] = _14700_ ^ _14699_ /*5262*/;
  assign _14701_ = _14700_ & _14699_ /*5261*/;
  assign _14702_ = inv_28[30] & r_27[30] /*5260*/;
  assign _14703_ = _14701_ | _14702_ /*5259*/;
  assign _14704_ = inv_28[31] ^ r_27[31] /*5257*/;
  assign sum_28[31] = _14704_ ^ _14703_ /*5256*/;
  assign _14705_ = _14704_ & _14703_ /*5255*/;
  assign _14706_ = inv_28[31] & r_27[31] /*5254*/;
  assign _14707_ = _14705_ | _14706_ /*5253*/;
  assign _14708_ = inv_28[32] ^ r_27[32] /*5251*/;
  assign sum_28[32] = _14708_ ^ _14707_ /*5250*/;
  assign _14709_ = _14708_ & _14707_ /*5249*/;
  assign _14710_ = inv_28[32] & r_27[32] /*5248*/;
  assign _14711_ = _14709_ | _14710_ /*5247*/;
  assign _14712_ = inv_28[33] ^ r_27[33] /*5245*/;
  assign sum_28[33] = _14712_ ^ _14711_ /*5244*/;
  assign _14713_ = _14712_ & _14711_ /*5243*/;
  assign _14714_ = inv_28[33] & r_27[33] /*5242*/;
  assign _14715_ = _14713_ | _14714_ /*5241*/;
  assign _14716_ = inv_28[34] ^ r_27[34] /*5239*/;
  assign sum_28[34] = _14716_ ^ _14715_ /*5238*/;
  assign _14717_ = _14716_ & _14715_ /*5237*/;
  assign _14718_ = inv_28[34] & r_27[34] /*5236*/;
  assign _14719_ = _14717_ | _14718_ /*5235*/;
  assign _14720_ = inv_28[35] ^ r_27[35] /*5233*/;
  assign sum_28[35] = _14720_ ^ _14719_ /*5232*/;
  assign _14721_ = _14720_ & _14719_ /*5231*/;
  assign _14722_ = inv_28[35] & r_27[35] /*5230*/;
  assign _14723_ = _14721_ | _14722_ /*5229*/;
  assign _14724_ = inv_28[36] ^ r_27[36] /*5227*/;
  assign sum_28[36] = _14724_ ^ _14723_ /*5226*/;
  assign _14725_ = _14724_ & _14723_ /*5225*/;
  assign _14726_ = inv_28[36] & r_27[36] /*5224*/;
  assign _14727_ = _14725_ | _14726_ /*5223*/;
  assign _14728_ = inv_28[37] ^ r_27[37] /*5221*/;
  assign sum_28[37] = _14728_ ^ _14727_ /*5220*/;
  assign _14729_ = _14728_ & _14727_ /*5219*/;
  assign _14730_ = inv_28[37] & r_27[37] /*5218*/;
  assign _14731_ = _14729_ | _14730_ /*5217*/;
  assign _14732_ = inv_28[38] ^ r_27[38] /*5215*/;
  assign sum_28[38] = _14732_ ^ _14731_ /*5214*/;
  assign _14733_ = _14732_ & _14731_ /*5213*/;
  assign _14734_ = inv_28[38] & r_27[38] /*5212*/;
  assign _14735_ = _14733_ | _14734_ /*5211*/;
  assign _14736_ = inv_28[39] ^ r_27[39] /*5209*/;
  assign sum_28[39] = _14736_ ^ _14735_ /*5208*/;
  assign _14737_ = _14736_ & _14735_ /*5207*/;
  assign _14738_ = inv_28[39] & r_27[39] /*5206*/;
  assign _14739_ = _14737_ | _14738_ /*5205*/;
  assign _14740_ = inv_28[40] ^ r_27[40] /*5203*/;
  assign sum_28[40] = _14740_ ^ _14739_ /*5202*/;
  assign _14741_ = _14740_ & _14739_ /*5201*/;
  assign _14742_ = inv_28[40] & r_27[40] /*5200*/;
  assign _14743_ = _14741_ | _14742_ /*5199*/;
  assign _14744_ = inv_28[41] ^ r_27[41] /*5197*/;
  assign sum_28[41] = _14744_ ^ _14743_ /*5196*/;
  assign _14745_ = _14744_ & _14743_ /*5195*/;
  assign _14746_ = inv_28[41] & r_27[41] /*5194*/;
  assign _14747_ = _14745_ | _14746_ /*5193*/;
  assign _14748_ = inv_28[42] ^ r_27[42] /*5191*/;
  assign sum_28[42] = _14748_ ^ _14747_ /*5190*/;
  assign _14749_ = _14748_ & _14747_ /*5189*/;
  assign _14750_ = inv_28[42] & r_27[42] /*5188*/;
  assign _14751_ = _14749_ | _14750_ /*5187*/;
  assign _14752_ = inv_28[43] ^ r_27[43] /*5185*/;
  assign sum_28[43] = _14752_ ^ _14751_ /*5184*/;
  assign _14753_ = _14752_ & _14751_ /*5183*/;
  assign _14754_ = inv_28[43] & r_27[43] /*5182*/;
  assign _14755_ = _14753_ | _14754_ /*5181*/;
  assign _14756_ = inv_28[44] ^ r_27[44] /*5179*/;
  assign sum_28[44] = _14756_ ^ _14755_ /*5178*/;
  assign _14757_ = _14756_ & _14755_ /*5177*/;
  assign _14758_ = inv_28[44] & r_27[44] /*5176*/;
  assign _14759_ = _14757_ | _14758_ /*5175*/;
  assign _14760_ = inv_28[45] ^ r_27[45] /*5173*/;
  assign sum_28[45] = _14760_ ^ _14759_ /*5172*/;
  assign _14761_ = _14760_ & _14759_ /*5171*/;
  assign _14762_ = inv_28[45] & r_27[45] /*5170*/;
  assign _14763_ = _14761_ | _14762_ /*5169*/;
  assign _14764_ = inv_28[46] ^ r_27[46] /*5167*/;
  assign sum_28[46] = _14764_ ^ _14763_ /*5166*/;
  assign _14765_ = _14764_ & _14763_ /*5165*/;
  assign _14766_ = inv_28[46] & r_27[46] /*5164*/;
  assign _14767_ = _14765_ | _14766_ /*5163*/;
  assign _14768_ = inv_28[47] ^ r_27[47] /*5161*/;
  assign sum_28[47] = _14768_ ^ _14767_ /*5160*/;
  assign _14769_ = _14768_ & _14767_ /*5159*/;
  assign _14770_ = inv_28[47] & r_27[47] /*5158*/;
  assign _14771_ = _14769_ | _14770_ /*5157*/;
  assign _14772_ = inv_28[48] ^ r_27[48] /*5155*/;
  assign sum_28[48] = _14772_ ^ _14771_ /*5154*/;
  assign _14773_ = _14772_ & _14771_ /*5153*/;
  assign _14774_ = inv_28[48] & r_27[48] /*5152*/;
  assign _14775_ = _14773_ | _14774_ /*5151*/;
  assign _14776_ = inv_28[49] ^ r_27[49] /*5149*/;
  assign sum_28[49] = _14776_ ^ _14775_ /*5148*/;
  assign _14777_ = _14776_ & _14775_ /*5147*/;
  assign _14778_ = inv_28[49] & r_27[49] /*5146*/;
  assign _14779_ = _14777_ | _14778_ /*5145*/;
  assign _14780_ = inv_28[50] ^ r_27[50] /*5143*/;
  assign sum_28[50] = _14780_ ^ _14779_ /*5142*/;
  assign _14781_ = _14780_ & _14779_ /*5141*/;
  assign _14782_ = inv_28[50] & r_27[50] /*5140*/;
  assign _14783_ = _14781_ | _14782_ /*5139*/;
  assign _14784_ = inv_28[51] ^ r_27[51] /*5137*/;
  assign sum_28[51] = _14784_ ^ _14783_ /*5136*/;
  assign _14785_ = _14784_ & _14783_ /*5135*/;
  assign _14786_ = inv_28[51] & r_27[51] /*5134*/;
  assign _14787_ = _14785_ | _14786_ /*5133*/;
  assign _14788_ = inv_28[52] ^ r_27[52] /*5131*/;
  assign sum_28[52] = _14788_ ^ _14787_ /*5130*/;
  assign _14789_ = _14788_ & _14787_ /*5129*/;
  assign _14790_ = inv_28[52] & r_27[52] /*5128*/;
  assign _14791_ = _14789_ | _14790_ /*5127*/;
  assign _14792_ = inv_28[53] ^ r_27[53] /*5125*/;
  assign sum_28[53] = _14792_ ^ _14791_ /*5124*/;
  assign _14793_ = _14792_ & _14791_ /*5123*/;
  assign _14794_ = inv_28[53] & r_27[53] /*5122*/;
  assign _14795_ = _14793_ | _14794_ /*5121*/;
  assign _14796_ = inv_28[54] ^ r_27[54] /*5119*/;
  assign sum_28[54] = _14796_ ^ _14795_ /*5118*/;
  assign _14797_ = _14796_ & _14795_ /*5117*/;
  assign _14798_ = inv_28[54] & r_27[54] /*5116*/;
  assign _14799_ = _14797_ | _14798_ /*5115*/;
  assign _14800_ = inv_28[55] ^ r_27[55] /*5113*/;
  assign sum_28[55] = _14800_ ^ _14799_ /*5112*/;
  assign _14801_ = _14800_ & _14799_ /*5111*/;
  assign _14802_ = inv_28[55] & r_27[55] /*5110*/;
  assign _14803_ = _14801_ | _14802_ /*5109*/;
  assign _14804_ = inv_28[56] ^ r_27[56] /*5107*/;
  assign sum_28[56] = _14804_ ^ _14803_ /*5106*/;
  assign _14805_ = _14804_ & _14803_ /*5105*/;
  assign _14806_ = inv_28[56] & r_27[56] /*5104*/;
  assign _14807_ = _14805_ | _14806_ /*5103*/;
  assign _14808_ = inv_28[57] ^ r_27[57] /*5101*/;
  assign sum_28[57] = _14808_ ^ _14807_ /*5100*/;
  assign _14809_ = _14808_ & _14807_ /*5099*/;
  assign _14810_ = inv_28[57] & r_27[57] /*5098*/;
  assign _14811_ = _14809_ | _14810_ /*5097*/;
  assign _14812_ = inv_28[58] ^ r_27[58] /*5095*/;
  assign sum_28[58] = _14812_ ^ _14811_ /*5094*/;
  assign _14813_ = _14812_ & _14811_ /*5093*/;
  assign _14814_ = inv_28[58] & r_27[58] /*5092*/;
  assign _14815_ = _14813_ | _14814_ /*5091*/;
  assign _14816_ = inv_28[59] ^ r_27[59] /*5089*/;
  assign sum_28[59] = _14816_ ^ _14815_ /*5088*/;
  assign _14817_ = _14816_ & _14815_ /*5087*/;
  assign _14818_ = inv_28[59] & r_27[59] /*5086*/;
  assign _14819_ = _14817_ | _14818_ /*5085*/;
  assign _14820_ = inv_28[60] ^ r_27[60] /*5083*/;
  assign sum_28[60] = _14820_ ^ _14819_ /*5082*/;
  assign _14821_ = _14820_ & _14819_ /*5081*/;
  assign _14822_ = inv_28[60] & r_27[60] /*5080*/;
  assign _14823_ = _14821_ | _14822_ /*5079*/;
  assign _14824_ = inv_28[61] ^ r_27[61] /*5077*/;
  assign sum_28[61] = _14824_ ^ _14823_ /*5076*/;
  assign _14825_ = _14824_ & _14823_ /*5075*/;
  assign _14826_ = inv_28[61] & r_27[61] /*5074*/;
  assign _14827_ = _14825_ | _14826_ /*5073*/;
  assign _14828_ = inv_28[62] ^ r_27[62] /*5071*/;
  assign sum_28[62] = _14828_ ^ _14827_ /*5070*/;
  assign _14829_ = _14828_ & _14827_ /*5069*/;
  assign _14830_ = inv_28[62] & r_27[62] /*5068*/;
  assign _14831_ = _14829_ | _14830_ /*5067*/;
  assign _14832_ = inv_28[63] ^ r_27[63] /*5065*/;
  assign sum_28[63] = _14832_ ^ _14831_ /*5064*/;
  assign _14833_ = _14832_ & _14831_ /*5063*/;
  assign _14834_ = inv_28[63] & r_27[63] /*5062*/;
  assign _14835_ = _14833_ | _14834_ /*5061*/;
  assign _14836_ = inv_28[64] ^ r_27[64] /*5059*/;
  assign sum_28[64] = _14836_ ^ _14835_ /*5058*/;
  assign _14837_ = _14836_ & _14835_ /*5057*/;
  assign _14838_ = inv_28[64] & r_27[64] /*5056*/;
  assign _14839_ = _14837_ | _14838_ /*5055*/;
  assign _14840_ = inv_28[65] ^ r_27[65] /*5053*/;
  assign sum_28[65] = _14840_ ^ _14839_ /*5052*/;
  assign _14841_ = _14840_ & _14839_ /*5051*/;
  assign _14842_ = inv_28[65] & r_27[65] /*5050*/;
  assign _14843_ = _14841_ | _14842_ /*5049*/;
  assign _14844_ = inv_28[66] ^ r_27[66] /*5047*/;
  assign sum_28[66] = _14844_ ^ _14843_ /*5046*/;
  assign _14845_ = _14844_ & _14843_ /*5045*/;
  assign _14846_ = inv_28[66] & r_27[66] /*5044*/;
  assign _14847_ = _14845_ | _14846_ /*5043*/;
  assign _14848_ = inv_28[67] ^ r_27[67] /*5041*/;
  assign sum_28[67] = _14848_ ^ _14847_ /*5040*/;
  assign _14849_ = _14848_ & _14847_ /*5039*/;
  assign _14850_ = inv_28[67] & r_27[67] /*5038*/;
  assign _14851_ = _14849_ | _14850_ /*5037*/;
  assign _14852_ = inv_28[68] ^ r_27[68] /*5035*/;
  assign sum_28[68] = _14852_ ^ _14851_ /*5034*/;
  assign _14853_ = _14852_ & _14851_ /*5033*/;
  assign _14854_ = inv_28[68] & r_27[68] /*5032*/;
  assign _14855_ = _14853_ | _14854_ /*5031*/;
  assign _14856_ = inv_28[69] ^ r_27[69] /*5029*/;
  assign sum_28[69] = _14856_ ^ _14855_ /*5028*/;
  assign _14857_ = _14856_ & _14855_ /*5027*/;
  assign _14858_ = inv_28[69] & r_27[69] /*5026*/;
  assign _14859_ = _14857_ | _14858_ /*5025*/;
  assign _14860_ = inv_28[70] ^ r_27[70] /*5023*/;
  assign sum_28[70] = _14860_ ^ _14859_ /*5022*/;
  assign _14861_ = _14860_ & _14859_ /*5021*/;
  assign _14862_ = inv_28[70] & r_27[70] /*5020*/;
  assign _14863_ = _14861_ | _14862_ /*5019*/;
  assign _14864_ = inv_28[71] ^ r_27[71] /*5017*/;
  assign sum_28[71] = _14864_ ^ _14863_ /*5016*/;
  assign _14865_ = _14864_ & _14863_ /*5015*/;
  assign _14866_ = inv_28[71] & r_27[71] /*5014*/;
  assign _14867_ = _14865_ | _14866_ /*5013*/;
  assign _14868_ = inv_28[72] ^ r_27[72] /*5011*/;
  assign sum_28[72] = _14868_ ^ _14867_ /*5010*/;
  assign _14869_ = _14868_ & _14867_ /*5009*/;
  assign _14870_ = inv_28[72] & r_27[72] /*5008*/;
  assign _14871_ = _14869_ | _14870_ /*5007*/;
  assign _14872_ = inv_28[73] ^ r_27[73] /*5005*/;
  assign sum_28[73] = _14872_ ^ _14871_ /*5004*/;
  assign _14873_ = _14872_ & _14871_ /*5003*/;
  assign _14874_ = inv_28[73] & r_27[73] /*5002*/;
  assign _14875_ = _14873_ | _14874_ /*5001*/;
  assign _14876_ = inv_28[74] ^ r_27[74] /*4999*/;
  assign sum_28[74] = _14876_ ^ _14875_ /*4998*/;
  assign _14877_ = _14876_ & _14875_ /*4997*/;
  assign _14878_ = inv_28[74] & r_27[74] /*4996*/;
  assign _14879_ = _14877_ | _14878_ /*4995*/;
  assign _14880_ = inv_28[75] ^ r_27[75] /*4993*/;
  assign sum_28[75] = _14880_ ^ _14879_ /*4992*/;
  assign _14881_ = _14880_ & _14879_ /*4991*/;
  assign _14882_ = inv_28[75] & r_27[75] /*4990*/;
  assign _14883_ = _14881_ | _14882_ /*4989*/;
  assign _14884_ = inv_28[76] ^ r_27[76] /*4987*/;
  assign sum_28[76] = _14884_ ^ _14883_ /*4986*/;
  assign _14885_ = _14884_ & _14883_ /*4985*/;
  assign _14886_ = inv_28[76] & r_27[76] /*4984*/;
  assign _14887_ = _14885_ | _14886_ /*4983*/;
  assign _14888_ = inv_28[77] ^ r_27[77] /*4981*/;
  assign sum_28[77] = _14888_ ^ _14887_ /*4980*/;
  assign _14889_ = _14888_ & _14887_ /*4979*/;
  assign _14890_ = inv_28[77] & r_27[77] /*4978*/;
  assign _14891_ = _14889_ | _14890_ /*4977*/;
  assign _14892_ = inv_28[78] ^ r_27[78] /*4975*/;
  assign sum_28[78] = _14892_ ^ _14891_ /*4974*/;
  assign _14893_ = _14892_ & _14891_ /*4973*/;
  assign _14894_ = inv_28[78] & r_27[78] /*4972*/;
  assign _14895_ = _14893_ | _14894_ /*4971*/;
  assign _14896_ = inv_28[79] ^ r_27[79] /*4969*/;
  assign sum_28[79] = _14896_ ^ _14895_ /*4968*/;
  assign _14897_ = _14896_ & _14895_ /*4967*/;
  assign _14898_ = inv_28[79] & r_27[79] /*4966*/;
  assign _14899_ = _14897_ | _14898_ /*4965*/;
  assign _14900_ = inv_28[80] ^ r_27[80] /*4963*/;
  assign sum_28[80] = _14900_ ^ _14899_ /*4962*/;
  assign _14901_ = _14900_ & _14899_ /*4961*/;
  assign _14902_ = inv_28[80] & r_27[80] /*4960*/;
  assign _14903_ = _14901_ | _14902_ /*4959*/;
  assign _14904_ = inv_28[81] ^ r_27[81] /*4957*/;
  assign sum_28[81] = _14904_ ^ _14903_ /*4956*/;
  assign _14905_ = _14904_ & _14903_ /*4955*/;
  assign _14906_ = inv_28[81] & r_27[81] /*4954*/;
  assign _14907_ = _14905_ | _14906_ /*4953*/;
  assign _14908_ = inv_28[82] ^ r_27[82] /*4951*/;
  assign sum_28[82] = _14908_ ^ _14907_ /*4950*/;
  assign _14909_ = _14908_ & _14907_ /*4949*/;
  assign _14910_ = inv_28[82] & r_27[82] /*4948*/;
  assign _14911_ = _14909_ | _14910_ /*4947*/;
  assign _14912_ = inv_28[83] ^ r_27[83] /*4945*/;
  assign sum_28[83] = _14912_ ^ _14911_ /*4944*/;
  assign _14913_ = _14912_ & _14911_ /*4943*/;
  assign _14914_ = inv_28[83] & r_27[83] /*4942*/;
  assign _14915_ = _14913_ | _14914_ /*4941*/;
  assign _14916_ = inv_28[84] ^ r_27[84] /*4939*/;
  assign sum_28[84] = _14916_ ^ _14915_ /*4938*/;
  assign _14917_ = _14916_ & _14915_ /*4937*/;
  assign _14918_ = inv_28[84] & r_27[84] /*4936*/;
  assign _14919_ = _14917_ | _14918_ /*4935*/;
  assign _14920_ = inv_28[85] ^ r_27[85] /*4933*/;
  assign sum_28[85] = _14920_ ^ _14919_ /*4932*/;
  assign _14921_ = _14920_ & _14919_ /*4931*/;
  assign _14922_ = inv_28[85] & r_27[85] /*4930*/;
  assign _14923_ = _14921_ | _14922_ /*4929*/;
  assign _14924_ = inv_28[86] ^ r_27[86] /*4927*/;
  assign sum_28[86] = _14924_ ^ _14923_ /*4926*/;
  assign _14925_ = _14924_ & _14923_ /*4925*/;
  assign _14926_ = inv_28[86] & r_27[86] /*4924*/;
  assign _14927_ = _14925_ | _14926_ /*4923*/;
  assign _14928_ = inv_28[87] ^ r_27[87] /*4921*/;
  assign sum_28[87] = _14928_ ^ _14927_ /*4920*/;
  assign _14929_ = _14928_ & _14927_ /*4919*/;
  assign _14930_ = inv_28[87] & r_27[87] /*4918*/;
  assign _14931_ = _14929_ | _14930_ /*4917*/;
  assign _14932_ = inv_28[88] ^ r_27[88] /*4915*/;
  assign sum_28[88] = _14932_ ^ _14931_ /*4914*/;
  assign _14933_ = _14932_ & _14931_ /*4913*/;
  assign _14934_ = inv_28[88] & r_27[88] /*4912*/;
  assign _14935_ = _14933_ | _14934_ /*4911*/;
  assign _14936_ = inv_28[89] ^ r_27[89] /*4909*/;
  assign sum_28[89] = _14936_ ^ _14935_ /*4908*/;
  assign _14937_ = _14936_ & _14935_ /*4907*/;
  assign _14938_ = inv_28[89] & r_27[89] /*4906*/;
  assign _14939_ = _14937_ | _14938_ /*4905*/;
  assign _14940_ = _14939_ ^ _14935_ /*4904*/;
  assign _14941_ = ~_14940_ /*4903*/;
  assign _14942_ = sum_28[89] & _14941_ /*4902*/;
  assign _14943_ = _14940_ & _14939_ /*4901*/;
  assign sum_28[90] = _14943_ | _14942_ /*4900*/;
  assign q[4] = ~sum_28[90] /*4899*/;
  assign m_28[0] = r_27[0] /*4898*/;
  assign m_28[1] = r_27[1] /*4897*/;
  assign m_28[2] = r_27[2] /*4896*/;
  assign m_28[3] = r_27[3] /*4895*/;
  assign m_28[4] = r_27[4] /*4894*/;
  assign m_28[5] = r_27[5] /*4893*/;
  assign m_28[6] = r_27[6] /*4892*/;
  assign m_28[7] = r_27[7] /*4891*/;
  assign m_28[8] = r_27[8] /*4890*/;
  assign m_28[9] = r_27[9] /*4889*/;
  assign m_28[10] = r_27[10] /*4888*/;
  assign m_28[11] = r_27[11] /*4887*/;
  assign m_28[12] = r_27[12] /*4886*/;
  assign m_28[13] = r_27[13] /*4885*/;
  assign m_28[14] = r_27[14] /*4884*/;
  assign m_28[15] = r_27[15] /*4883*/;
  assign m_28[16] = r_27[16] /*4882*/;
  assign m_28[17] = r_27[17] /*4881*/;
  assign m_28[18] = r_27[18] /*4880*/;
  assign m_28[19] = r_27[19] /*4879*/;
  assign m_28[20] = r_27[20] /*4878*/;
  assign m_28[21] = r_27[21] /*4877*/;
  assign m_28[22] = r_27[22] /*4876*/;
  assign m_28[23] = r_27[23] /*4875*/;
  assign m_28[24] = r_27[24] /*4874*/;
  assign m_28[25] = r_27[25] /*4873*/;
  assign m_28[26] = r_27[26] /*4872*/;
  assign m_28[27] = r_27[27] /*4871*/;
  assign m_28[28] = r_27[28] /*4870*/;
  assign m_28[29] = r_27[29] /*4869*/;
  assign m_28[30] = r_27[30] /*4868*/;
  assign m_28[31] = r_27[31] /*4867*/;
  assign m_28[32] = r_27[32] /*4866*/;
  assign m_28[33] = r_27[33] /*4865*/;
  assign m_28[34] = r_27[34] /*4864*/;
  assign m_28[35] = r_27[35] /*4863*/;
  assign m_28[36] = r_27[36] /*4862*/;
  assign m_28[37] = r_27[37] /*4861*/;
  assign m_28[38] = r_27[38] /*4860*/;
  assign m_28[39] = r_27[39] /*4859*/;
  assign m_28[40] = r_27[40] /*4858*/;
  assign m_28[41] = r_27[41] /*4857*/;
  assign m_28[42] = r_27[42] /*4856*/;
  assign m_28[43] = r_27[43] /*4855*/;
  assign m_28[44] = r_27[44] /*4854*/;
  assign m_28[45] = r_27[45] /*4853*/;
  assign m_28[46] = r_27[46] /*4852*/;
  assign m_28[47] = r_27[47] /*4851*/;
  assign m_28[48] = r_27[48] /*4850*/;
  assign m_28[49] = r_27[49] /*4849*/;
  assign m_28[50] = r_27[50] /*4848*/;
  assign m_28[51] = r_27[51] /*4847*/;
  assign m_28[52] = r_27[52] /*4846*/;
  assign m_28[53] = r_27[53] /*4845*/;
  assign m_28[54] = r_27[54] /*4844*/;
  assign m_28[55] = r_27[55] /*4843*/;
  assign m_28[56] = r_27[56] /*4842*/;
  assign m_28[57] = r_27[57] /*4841*/;
  assign m_28[58] = r_27[58] /*4840*/;
  assign m_28[59] = r_27[59] /*4839*/;
  assign m_28[60] = r_27[60] /*4838*/;
  assign m_28[61] = r_27[61] /*4837*/;
  assign m_28[62] = r_27[62] /*4836*/;
  assign m_28[63] = r_27[63] /*4835*/;
  assign m_28[64] = r_27[64] /*4834*/;
  assign m_28[65] = r_27[65] /*4833*/;
  assign m_28[66] = r_27[66] /*4832*/;
  assign m_28[67] = r_27[67] /*4831*/;
  assign m_28[68] = r_27[68] /*4830*/;
  assign m_28[69] = r_27[69] /*4829*/;
  assign m_28[70] = r_27[70] /*4828*/;
  assign m_28[71] = r_27[71] /*4827*/;
  assign m_28[72] = r_27[72] /*4826*/;
  assign m_28[73] = r_27[73] /*4825*/;
  assign m_28[74] = r_27[74] /*4824*/;
  assign m_28[75] = r_27[75] /*4823*/;
  assign m_28[76] = r_27[76] /*4822*/;
  assign m_28[77] = r_27[77] /*4821*/;
  assign m_28[78] = r_27[78] /*4820*/;
  assign m_28[79] = r_27[79] /*4819*/;
  assign m_28[80] = r_27[80] /*4818*/;
  assign m_28[81] = r_27[81] /*4817*/;
  assign m_28[82] = r_27[82] /*4816*/;
  assign m_28[83] = r_27[83] /*4815*/;
  assign m_28[84] = r_27[84] /*4814*/;
  assign m_28[85] = r_27[85] /*4813*/;
  assign m_28[86] = r_27[86] /*4812*/;
  assign m_28[87] = r_27[87] /*4811*/;
  assign m_28[88] = r_27[88] /*4810*/;
  assign m_28[89] = r_27[89] /*4809*/;
  assign m_28[90] = r_27[89] /*4808*/;
  assign _14945_ = ~q[4] /*4807*/;
  assign _14946_ = sum_28[0] & q[4] /*4806*/;
  assign _14947_ = m_28[0] & _14945_ /*4805*/;
  assign r_28[0] = _14947_ | _14946_ /*4804*/;
  assign _14948_ = ~q[4] /*4803*/;
  assign _14949_ = sum_28[1] & q[4] /*4802*/;
  assign _14950_ = m_28[1] & _14948_ /*4801*/;
  assign r_28[1] = _14950_ | _14949_ /*4800*/;
  assign _14951_ = ~q[4] /*4799*/;
  assign _14952_ = sum_28[2] & q[4] /*4798*/;
  assign _14953_ = m_28[2] & _14951_ /*4797*/;
  assign r_28[2] = _14953_ | _14952_ /*4796*/;
  assign _14954_ = ~q[4] /*4795*/;
  assign _14955_ = sum_28[3] & q[4] /*4794*/;
  assign _14956_ = m_28[3] & _14954_ /*4793*/;
  assign r_28[3] = _14956_ | _14955_ /*4792*/;
  assign _14957_ = ~q[4] /*4791*/;
  assign _14958_ = sum_28[4] & q[4] /*4790*/;
  assign _14959_ = m_28[4] & _14957_ /*4789*/;
  assign r_28[4] = _14959_ | _14958_ /*4788*/;
  assign _14960_ = ~q[4] /*4787*/;
  assign _14961_ = sum_28[5] & q[4] /*4786*/;
  assign _14962_ = m_28[5] & _14960_ /*4785*/;
  assign r_28[5] = _14962_ | _14961_ /*4784*/;
  assign _14963_ = ~q[4] /*4783*/;
  assign _14964_ = sum_28[6] & q[4] /*4782*/;
  assign _14965_ = m_28[6] & _14963_ /*4781*/;
  assign r_28[6] = _14965_ | _14964_ /*4780*/;
  assign _14966_ = ~q[4] /*4779*/;
  assign _14967_ = sum_28[7] & q[4] /*4778*/;
  assign _14968_ = m_28[7] & _14966_ /*4777*/;
  assign r_28[7] = _14968_ | _14967_ /*4776*/;
  assign _14969_ = ~q[4] /*4775*/;
  assign _14970_ = sum_28[8] & q[4] /*4774*/;
  assign _14971_ = m_28[8] & _14969_ /*4773*/;
  assign r_28[8] = _14971_ | _14970_ /*4772*/;
  assign _14972_ = ~q[4] /*4771*/;
  assign _14973_ = sum_28[9] & q[4] /*4770*/;
  assign _14974_ = m_28[9] & _14972_ /*4769*/;
  assign r_28[9] = _14974_ | _14973_ /*4768*/;
  assign _14975_ = ~q[4] /*4767*/;
  assign _14976_ = sum_28[10] & q[4] /*4766*/;
  assign _14977_ = m_28[10] & _14975_ /*4765*/;
  assign r_28[10] = _14977_ | _14976_ /*4764*/;
  assign _14978_ = ~q[4] /*4763*/;
  assign _14979_ = sum_28[11] & q[4] /*4762*/;
  assign _14980_ = m_28[11] & _14978_ /*4761*/;
  assign r_28[11] = _14980_ | _14979_ /*4760*/;
  assign _14981_ = ~q[4] /*4759*/;
  assign _14982_ = sum_28[12] & q[4] /*4758*/;
  assign _14983_ = m_28[12] & _14981_ /*4757*/;
  assign r_28[12] = _14983_ | _14982_ /*4756*/;
  assign _14984_ = ~q[4] /*4755*/;
  assign _14985_ = sum_28[13] & q[4] /*4754*/;
  assign _14986_ = m_28[13] & _14984_ /*4753*/;
  assign r_28[13] = _14986_ | _14985_ /*4752*/;
  assign _14987_ = ~q[4] /*4751*/;
  assign _14988_ = sum_28[14] & q[4] /*4750*/;
  assign _14989_ = m_28[14] & _14987_ /*4749*/;
  assign r_28[14] = _14989_ | _14988_ /*4748*/;
  assign _14990_ = ~q[4] /*4747*/;
  assign _14991_ = sum_28[15] & q[4] /*4746*/;
  assign _14992_ = m_28[15] & _14990_ /*4745*/;
  assign r_28[15] = _14992_ | _14991_ /*4744*/;
  assign _14993_ = ~q[4] /*4743*/;
  assign _14994_ = sum_28[16] & q[4] /*4742*/;
  assign _14995_ = m_28[16] & _14993_ /*4741*/;
  assign r_28[16] = _14995_ | _14994_ /*4740*/;
  assign _14996_ = ~q[4] /*4739*/;
  assign _14997_ = sum_28[17] & q[4] /*4738*/;
  assign _14998_ = m_28[17] & _14996_ /*4737*/;
  assign r_28[17] = _14998_ | _14997_ /*4736*/;
  assign _14999_ = ~q[4] /*4735*/;
  assign _15000_ = sum_28[18] & q[4] /*4734*/;
  assign _15001_ = m_28[18] & _14999_ /*4733*/;
  assign r_28[18] = _15001_ | _15000_ /*4732*/;
  assign _15002_ = ~q[4] /*4731*/;
  assign _15003_ = sum_28[19] & q[4] /*4730*/;
  assign _15004_ = m_28[19] & _15002_ /*4729*/;
  assign r_28[19] = _15004_ | _15003_ /*4728*/;
  assign _15005_ = ~q[4] /*4727*/;
  assign _15006_ = sum_28[20] & q[4] /*4726*/;
  assign _15007_ = m_28[20] & _15005_ /*4725*/;
  assign r_28[20] = _15007_ | _15006_ /*4724*/;
  assign _15008_ = ~q[4] /*4723*/;
  assign _15009_ = sum_28[21] & q[4] /*4722*/;
  assign _15010_ = m_28[21] & _15008_ /*4721*/;
  assign r_28[21] = _15010_ | _15009_ /*4720*/;
  assign _15011_ = ~q[4] /*4719*/;
  assign _15012_ = sum_28[22] & q[4] /*4718*/;
  assign _15013_ = m_28[22] & _15011_ /*4717*/;
  assign r_28[22] = _15013_ | _15012_ /*4716*/;
  assign _15014_ = ~q[4] /*4715*/;
  assign _15015_ = sum_28[23] & q[4] /*4714*/;
  assign _15016_ = m_28[23] & _15014_ /*4713*/;
  assign r_28[23] = _15016_ | _15015_ /*4712*/;
  assign _15017_ = ~q[4] /*4711*/;
  assign _15018_ = sum_28[24] & q[4] /*4710*/;
  assign _15019_ = m_28[24] & _15017_ /*4709*/;
  assign r_28[24] = _15019_ | _15018_ /*4708*/;
  assign _15020_ = ~q[4] /*4707*/;
  assign _15021_ = sum_28[25] & q[4] /*4706*/;
  assign _15022_ = m_28[25] & _15020_ /*4705*/;
  assign r_28[25] = _15022_ | _15021_ /*4704*/;
  assign _15023_ = ~q[4] /*4703*/;
  assign _15024_ = sum_28[26] & q[4] /*4702*/;
  assign _15025_ = m_28[26] & _15023_ /*4701*/;
  assign r_28[26] = _15025_ | _15024_ /*4700*/;
  assign _15026_ = ~q[4] /*4699*/;
  assign _15027_ = sum_28[27] & q[4] /*4698*/;
  assign _15028_ = m_28[27] & _15026_ /*4697*/;
  assign r_28[27] = _15028_ | _15027_ /*4696*/;
  assign _15029_ = ~q[4] /*4695*/;
  assign _15030_ = sum_28[28] & q[4] /*4694*/;
  assign _15031_ = m_28[28] & _15029_ /*4693*/;
  assign r_28[28] = _15031_ | _15030_ /*4692*/;
  assign _15032_ = ~q[4] /*4691*/;
  assign _15033_ = sum_28[29] & q[4] /*4690*/;
  assign _15034_ = m_28[29] & _15032_ /*4689*/;
  assign r_28[29] = _15034_ | _15033_ /*4688*/;
  assign _15035_ = ~q[4] /*4687*/;
  assign _15036_ = sum_28[30] & q[4] /*4686*/;
  assign _15037_ = m_28[30] & _15035_ /*4685*/;
  assign r_28[30] = _15037_ | _15036_ /*4684*/;
  assign _15038_ = ~q[4] /*4683*/;
  assign _15039_ = sum_28[31] & q[4] /*4682*/;
  assign _15040_ = m_28[31] & _15038_ /*4681*/;
  assign r_28[31] = _15040_ | _15039_ /*4680*/;
  assign _15041_ = ~q[4] /*4679*/;
  assign _15042_ = sum_28[32] & q[4] /*4678*/;
  assign _15043_ = m_28[32] & _15041_ /*4677*/;
  assign r_28[32] = _15043_ | _15042_ /*4676*/;
  assign _15044_ = ~q[4] /*4675*/;
  assign _15045_ = sum_28[33] & q[4] /*4674*/;
  assign _15046_ = m_28[33] & _15044_ /*4673*/;
  assign r_28[33] = _15046_ | _15045_ /*4672*/;
  assign _15047_ = ~q[4] /*4671*/;
  assign _15048_ = sum_28[34] & q[4] /*4670*/;
  assign _15049_ = m_28[34] & _15047_ /*4669*/;
  assign r_28[34] = _15049_ | _15048_ /*4668*/;
  assign _15050_ = ~q[4] /*4667*/;
  assign _15051_ = sum_28[35] & q[4] /*4666*/;
  assign _15052_ = m_28[35] & _15050_ /*4665*/;
  assign r_28[35] = _15052_ | _15051_ /*4664*/;
  assign _15053_ = ~q[4] /*4663*/;
  assign _15054_ = sum_28[36] & q[4] /*4662*/;
  assign _15055_ = m_28[36] & _15053_ /*4661*/;
  assign r_28[36] = _15055_ | _15054_ /*4660*/;
  assign _15056_ = ~q[4] /*4659*/;
  assign _15057_ = sum_28[37] & q[4] /*4658*/;
  assign _15058_ = m_28[37] & _15056_ /*4657*/;
  assign r_28[37] = _15058_ | _15057_ /*4656*/;
  assign _15059_ = ~q[4] /*4655*/;
  assign _15060_ = sum_28[38] & q[4] /*4654*/;
  assign _15061_ = m_28[38] & _15059_ /*4653*/;
  assign r_28[38] = _15061_ | _15060_ /*4652*/;
  assign _15062_ = ~q[4] /*4651*/;
  assign _15063_ = sum_28[39] & q[4] /*4650*/;
  assign _15064_ = m_28[39] & _15062_ /*4649*/;
  assign r_28[39] = _15064_ | _15063_ /*4648*/;
  assign _15065_ = ~q[4] /*4647*/;
  assign _15066_ = sum_28[40] & q[4] /*4646*/;
  assign _15067_ = m_28[40] & _15065_ /*4645*/;
  assign r_28[40] = _15067_ | _15066_ /*4644*/;
  assign _15068_ = ~q[4] /*4643*/;
  assign _15069_ = sum_28[41] & q[4] /*4642*/;
  assign _15070_ = m_28[41] & _15068_ /*4641*/;
  assign r_28[41] = _15070_ | _15069_ /*4640*/;
  assign _15071_ = ~q[4] /*4639*/;
  assign _15072_ = sum_28[42] & q[4] /*4638*/;
  assign _15073_ = m_28[42] & _15071_ /*4637*/;
  assign r_28[42] = _15073_ | _15072_ /*4636*/;
  assign _15074_ = ~q[4] /*4635*/;
  assign _15075_ = sum_28[43] & q[4] /*4634*/;
  assign _15076_ = m_28[43] & _15074_ /*4633*/;
  assign r_28[43] = _15076_ | _15075_ /*4632*/;
  assign _15077_ = ~q[4] /*4631*/;
  assign _15078_ = sum_28[44] & q[4] /*4630*/;
  assign _15079_ = m_28[44] & _15077_ /*4629*/;
  assign r_28[44] = _15079_ | _15078_ /*4628*/;
  assign _15080_ = ~q[4] /*4627*/;
  assign _15081_ = sum_28[45] & q[4] /*4626*/;
  assign _15082_ = m_28[45] & _15080_ /*4625*/;
  assign r_28[45] = _15082_ | _15081_ /*4624*/;
  assign _15083_ = ~q[4] /*4623*/;
  assign _15084_ = sum_28[46] & q[4] /*4622*/;
  assign _15085_ = m_28[46] & _15083_ /*4621*/;
  assign r_28[46] = _15085_ | _15084_ /*4620*/;
  assign _15086_ = ~q[4] /*4619*/;
  assign _15087_ = sum_28[47] & q[4] /*4618*/;
  assign _15088_ = m_28[47] & _15086_ /*4617*/;
  assign r_28[47] = _15088_ | _15087_ /*4616*/;
  assign _15089_ = ~q[4] /*4615*/;
  assign _15090_ = sum_28[48] & q[4] /*4614*/;
  assign _15091_ = m_28[48] & _15089_ /*4613*/;
  assign r_28[48] = _15091_ | _15090_ /*4612*/;
  assign _15092_ = ~q[4] /*4611*/;
  assign _15093_ = sum_28[49] & q[4] /*4610*/;
  assign _15094_ = m_28[49] & _15092_ /*4609*/;
  assign r_28[49] = _15094_ | _15093_ /*4608*/;
  assign _15095_ = ~q[4] /*4607*/;
  assign _15096_ = sum_28[50] & q[4] /*4606*/;
  assign _15097_ = m_28[50] & _15095_ /*4605*/;
  assign r_28[50] = _15097_ | _15096_ /*4604*/;
  assign _15098_ = ~q[4] /*4603*/;
  assign _15099_ = sum_28[51] & q[4] /*4602*/;
  assign _15100_ = m_28[51] & _15098_ /*4601*/;
  assign r_28[51] = _15100_ | _15099_ /*4600*/;
  assign _15101_ = ~q[4] /*4599*/;
  assign _15102_ = sum_28[52] & q[4] /*4598*/;
  assign _15103_ = m_28[52] & _15101_ /*4597*/;
  assign r_28[52] = _15103_ | _15102_ /*4596*/;
  assign _15104_ = ~q[4] /*4595*/;
  assign _15105_ = sum_28[53] & q[4] /*4594*/;
  assign _15106_ = m_28[53] & _15104_ /*4593*/;
  assign r_28[53] = _15106_ | _15105_ /*4592*/;
  assign _15107_ = ~q[4] /*4591*/;
  assign _15108_ = sum_28[54] & q[4] /*4590*/;
  assign _15109_ = m_28[54] & _15107_ /*4589*/;
  assign r_28[54] = _15109_ | _15108_ /*4588*/;
  assign _15110_ = ~q[4] /*4587*/;
  assign _15111_ = sum_28[55] & q[4] /*4586*/;
  assign _15112_ = m_28[55] & _15110_ /*4585*/;
  assign r_28[55] = _15112_ | _15111_ /*4584*/;
  assign _15113_ = ~q[4] /*4583*/;
  assign _15114_ = sum_28[56] & q[4] /*4582*/;
  assign _15115_ = m_28[56] & _15113_ /*4581*/;
  assign r_28[56] = _15115_ | _15114_ /*4580*/;
  assign _15116_ = ~q[4] /*4579*/;
  assign _15117_ = sum_28[57] & q[4] /*4578*/;
  assign _15118_ = m_28[57] & _15116_ /*4577*/;
  assign r_28[57] = _15118_ | _15117_ /*4576*/;
  assign _15119_ = ~q[4] /*4575*/;
  assign _15120_ = sum_28[58] & q[4] /*4574*/;
  assign _15121_ = m_28[58] & _15119_ /*4573*/;
  assign r_28[58] = _15121_ | _15120_ /*4572*/;
  assign _15122_ = ~q[4] /*4571*/;
  assign _15123_ = sum_28[59] & q[4] /*4570*/;
  assign _15124_ = m_28[59] & _15122_ /*4569*/;
  assign r_28[59] = _15124_ | _15123_ /*4568*/;
  assign _15125_ = ~q[4] /*4567*/;
  assign _15126_ = sum_28[60] & q[4] /*4566*/;
  assign _15127_ = m_28[60] & _15125_ /*4565*/;
  assign r_28[60] = _15127_ | _15126_ /*4564*/;
  assign _15128_ = ~q[4] /*4563*/;
  assign _15129_ = sum_28[61] & q[4] /*4562*/;
  assign _15130_ = m_28[61] & _15128_ /*4561*/;
  assign r_28[61] = _15130_ | _15129_ /*4560*/;
  assign _15131_ = ~q[4] /*4559*/;
  assign _15132_ = sum_28[62] & q[4] /*4558*/;
  assign _15133_ = m_28[62] & _15131_ /*4557*/;
  assign r_28[62] = _15133_ | _15132_ /*4556*/;
  assign _15134_ = ~q[4] /*4555*/;
  assign _15135_ = sum_28[63] & q[4] /*4554*/;
  assign _15136_ = m_28[63] & _15134_ /*4553*/;
  assign r_28[63] = _15136_ | _15135_ /*4552*/;
  assign _15137_ = ~q[4] /*4551*/;
  assign _15138_ = sum_28[64] & q[4] /*4550*/;
  assign _15139_ = m_28[64] & _15137_ /*4549*/;
  assign r_28[64] = _15139_ | _15138_ /*4548*/;
  assign _15140_ = ~q[4] /*4547*/;
  assign _15141_ = sum_28[65] & q[4] /*4546*/;
  assign _15142_ = m_28[65] & _15140_ /*4545*/;
  assign r_28[65] = _15142_ | _15141_ /*4544*/;
  assign _15143_ = ~q[4] /*4543*/;
  assign _15144_ = sum_28[66] & q[4] /*4542*/;
  assign _15145_ = m_28[66] & _15143_ /*4541*/;
  assign r_28[66] = _15145_ | _15144_ /*4540*/;
  assign _15146_ = ~q[4] /*4539*/;
  assign _15147_ = sum_28[67] & q[4] /*4538*/;
  assign _15148_ = m_28[67] & _15146_ /*4537*/;
  assign r_28[67] = _15148_ | _15147_ /*4536*/;
  assign _15149_ = ~q[4] /*4535*/;
  assign _15150_ = sum_28[68] & q[4] /*4534*/;
  assign _15151_ = m_28[68] & _15149_ /*4533*/;
  assign r_28[68] = _15151_ | _15150_ /*4532*/;
  assign _15152_ = ~q[4] /*4531*/;
  assign _15153_ = sum_28[69] & q[4] /*4530*/;
  assign _15154_ = m_28[69] & _15152_ /*4529*/;
  assign r_28[69] = _15154_ | _15153_ /*4528*/;
  assign _15155_ = ~q[4] /*4527*/;
  assign _15156_ = sum_28[70] & q[4] /*4526*/;
  assign _15157_ = m_28[70] & _15155_ /*4525*/;
  assign r_28[70] = _15157_ | _15156_ /*4524*/;
  assign _15158_ = ~q[4] /*4523*/;
  assign _15159_ = sum_28[71] & q[4] /*4522*/;
  assign _15160_ = m_28[71] & _15158_ /*4521*/;
  assign r_28[71] = _15160_ | _15159_ /*4520*/;
  assign _15161_ = ~q[4] /*4519*/;
  assign _15162_ = sum_28[72] & q[4] /*4518*/;
  assign _15163_ = m_28[72] & _15161_ /*4517*/;
  assign r_28[72] = _15163_ | _15162_ /*4516*/;
  assign _15164_ = ~q[4] /*4515*/;
  assign _15165_ = sum_28[73] & q[4] /*4514*/;
  assign _15166_ = m_28[73] & _15164_ /*4513*/;
  assign r_28[73] = _15166_ | _15165_ /*4512*/;
  assign _15167_ = ~q[4] /*4511*/;
  assign _15168_ = sum_28[74] & q[4] /*4510*/;
  assign _15169_ = m_28[74] & _15167_ /*4509*/;
  assign r_28[74] = _15169_ | _15168_ /*4508*/;
  assign _15170_ = ~q[4] /*4507*/;
  assign _15171_ = sum_28[75] & q[4] /*4506*/;
  assign _15172_ = m_28[75] & _15170_ /*4505*/;
  assign r_28[75] = _15172_ | _15171_ /*4504*/;
  assign _15173_ = ~q[4] /*4503*/;
  assign _15174_ = sum_28[76] & q[4] /*4502*/;
  assign _15175_ = m_28[76] & _15173_ /*4501*/;
  assign r_28[76] = _15175_ | _15174_ /*4500*/;
  assign _15176_ = ~q[4] /*4499*/;
  assign _15177_ = sum_28[77] & q[4] /*4498*/;
  assign _15178_ = m_28[77] & _15176_ /*4497*/;
  assign r_28[77] = _15178_ | _15177_ /*4496*/;
  assign _15179_ = ~q[4] /*4495*/;
  assign _15180_ = sum_28[78] & q[4] /*4494*/;
  assign _15181_ = m_28[78] & _15179_ /*4493*/;
  assign r_28[78] = _15181_ | _15180_ /*4492*/;
  assign _15182_ = ~q[4] /*4491*/;
  assign _15183_ = sum_28[79] & q[4] /*4490*/;
  assign _15184_ = m_28[79] & _15182_ /*4489*/;
  assign r_28[79] = _15184_ | _15183_ /*4488*/;
  assign _15185_ = ~q[4] /*4487*/;
  assign _15186_ = sum_28[80] & q[4] /*4486*/;
  assign _15187_ = m_28[80] & _15185_ /*4485*/;
  assign r_28[80] = _15187_ | _15186_ /*4484*/;
  assign _15188_ = ~q[4] /*4483*/;
  assign _15189_ = sum_28[81] & q[4] /*4482*/;
  assign _15190_ = m_28[81] & _15188_ /*4481*/;
  assign r_28[81] = _15190_ | _15189_ /*4480*/;
  assign _15191_ = ~q[4] /*4479*/;
  assign _15192_ = sum_28[82] & q[4] /*4478*/;
  assign _15193_ = m_28[82] & _15191_ /*4477*/;
  assign r_28[82] = _15193_ | _15192_ /*4476*/;
  assign _15194_ = ~q[4] /*4475*/;
  assign _15195_ = sum_28[83] & q[4] /*4474*/;
  assign _15196_ = m_28[83] & _15194_ /*4473*/;
  assign r_28[83] = _15196_ | _15195_ /*4472*/;
  assign _15197_ = ~q[4] /*4471*/;
  assign _15198_ = sum_28[84] & q[4] /*4470*/;
  assign _15199_ = m_28[84] & _15197_ /*4469*/;
  assign r_28[84] = _15199_ | _15198_ /*4468*/;
  assign _15200_ = ~q[4] /*4467*/;
  assign _15201_ = sum_28[85] & q[4] /*4466*/;
  assign _15202_ = m_28[85] & _15200_ /*4465*/;
  assign r_28[85] = _15202_ | _15201_ /*4464*/;
  assign _15203_ = ~q[4] /*4463*/;
  assign _15204_ = sum_28[86] & q[4] /*4462*/;
  assign _15205_ = m_28[86] & _15203_ /*4461*/;
  assign r_28[86] = _15205_ | _15204_ /*4460*/;
  assign _15206_ = ~q[4] /*4459*/;
  assign _15207_ = sum_28[87] & q[4] /*4458*/;
  assign _15208_ = m_28[87] & _15206_ /*4457*/;
  assign r_28[87] = _15208_ | _15207_ /*4456*/;
  assign _15209_ = ~q[4] /*4455*/;
  assign _15210_ = sum_28[88] & q[4] /*4454*/;
  assign _15211_ = m_28[88] & _15209_ /*4453*/;
  assign r_28[88] = _15211_ | _15210_ /*4452*/;
  assign _15212_ = ~q[4] /*4451*/;
  assign _15213_ = sum_28[89] & q[4] /*4450*/;
  assign _15214_ = m_28[89] & _15212_ /*4449*/;
  assign r_28[89] = _15214_ | _15213_ /*4448*/;
  assign _15215_ = ~q[4] /*4447*/;
  assign _15216_ = sum_28[90] & q[4] /*4446*/;
  assign _15217_ = m_28[90] & _15215_ /*4445*/;
  assign r_28[90] = _15217_ | _15216_ /*4444*/;
  assign inv_29[0] = oneWire /*4368*/;
  assign inv_29[1] = oneWire /*4362*/;
  assign inv_29[2] = oneWire /*4356*/;
  assign inv_29[3] = ~div[0] /*4350*/;
  assign inv_29[4] = ~div[1] /*4344*/;
  assign inv_29[5] = ~div[2] /*4338*/;
  assign inv_29[6] = ~div[3] /*4332*/;
  assign inv_29[7] = ~div[4] /*4326*/;
  assign inv_29[8] = ~div[5] /*4320*/;
  assign inv_29[9] = ~div[6] /*4314*/;
  assign inv_29[10] = ~div[7] /*4308*/;
  assign inv_29[11] = ~div[8] /*4302*/;
  assign inv_29[12] = ~div[9] /*4296*/;
  assign inv_29[13] = ~div[10] /*4290*/;
  assign inv_29[14] = ~div[11] /*4284*/;
  assign inv_29[15] = ~div[12] /*4278*/;
  assign inv_29[16] = ~div[13] /*4272*/;
  assign inv_29[17] = ~div[14] /*4266*/;
  assign inv_29[18] = ~div[15] /*4260*/;
  assign inv_29[19] = ~div[16] /*4254*/;
  assign inv_29[20] = ~div[17] /*4248*/;
  assign inv_29[21] = ~div[18] /*4242*/;
  assign inv_29[22] = ~div[19] /*4236*/;
  assign inv_29[23] = ~div[20] /*4230*/;
  assign inv_29[24] = ~div[21] /*4224*/;
  assign inv_29[25] = ~div[22] /*4218*/;
  assign inv_29[26] = ~div[23] /*4212*/;
  assign inv_29[27] = ~div[24] /*4206*/;
  assign inv_29[28] = ~div[25] /*4200*/;
  assign inv_29[29] = ~div[26] /*4194*/;
  assign inv_29[30] = ~div[27] /*4188*/;
  assign inv_29[31] = ~div[28] /*4182*/;
  assign inv_29[32] = ~div[29] /*4176*/;
  assign inv_29[33] = ~div[30] /*4170*/;
  assign inv_29[34] = oneWire /*4164*/;
  assign inv_29[35] = oneWire /*4158*/;
  assign inv_29[36] = oneWire /*4152*/;
  assign inv_29[37] = oneWire /*4146*/;
  assign inv_29[38] = oneWire /*4140*/;
  assign inv_29[39] = oneWire /*4134*/;
  assign inv_29[40] = oneWire /*4128*/;
  assign inv_29[41] = oneWire /*4122*/;
  assign inv_29[42] = oneWire /*4116*/;
  assign inv_29[43] = oneWire /*4110*/;
  assign inv_29[44] = oneWire /*4104*/;
  assign inv_29[45] = oneWire /*4098*/;
  assign inv_29[46] = oneWire /*4092*/;
  assign inv_29[47] = oneWire /*4086*/;
  assign inv_29[48] = oneWire /*4080*/;
  assign inv_29[49] = oneWire /*4074*/;
  assign inv_29[50] = oneWire /*4068*/;
  assign inv_29[51] = oneWire /*4062*/;
  assign inv_29[52] = oneWire /*4056*/;
  assign inv_29[53] = oneWire /*4050*/;
  assign inv_29[54] = oneWire /*4044*/;
  assign inv_29[55] = oneWire /*4038*/;
  assign inv_29[56] = oneWire /*4032*/;
  assign inv_29[57] = oneWire /*4026*/;
  assign inv_29[58] = oneWire /*4020*/;
  assign inv_29[59] = oneWire /*4014*/;
  assign inv_29[60] = oneWire /*4008*/;
  assign inv_29[61] = oneWire /*4002*/;
  assign inv_29[62] = oneWire /*3996*/;
  assign inv_29[63] = oneWire /*3990*/;
  assign inv_29[64] = oneWire /*3984*/;
  assign inv_29[65] = oneWire /*3978*/;
  assign inv_29[66] = oneWire /*3972*/;
  assign inv_29[67] = oneWire /*3966*/;
  assign inv_29[68] = oneWire /*3960*/;
  assign inv_29[69] = oneWire /*3954*/;
  assign inv_29[70] = oneWire /*3948*/;
  assign inv_29[71] = oneWire /*3942*/;
  assign inv_29[72] = oneWire /*3936*/;
  assign inv_29[73] = oneWire /*3930*/;
  assign inv_29[74] = oneWire /*3924*/;
  assign inv_29[75] = oneWire /*3918*/;
  assign inv_29[76] = oneWire /*3912*/;
  assign inv_29[77] = oneWire /*3906*/;
  assign inv_29[78] = oneWire /*3900*/;
  assign inv_29[79] = oneWire /*3894*/;
  assign inv_29[80] = oneWire /*3888*/;
  assign inv_29[81] = oneWire /*3882*/;
  assign inv_29[82] = oneWire /*3876*/;
  assign inv_29[83] = oneWire /*3870*/;
  assign inv_29[84] = oneWire /*3864*/;
  assign inv_29[85] = oneWire /*3858*/;
  assign inv_29[86] = oneWire /*3852*/;
  assign inv_29[87] = oneWire /*3846*/;
  assign inv_29[88] = oneWire /*3840*/;
  assign inv_29[89] = oneWire /*3834*/;
  assign inv_29[90] = oneWire /*3828*/;
  assign _15218_ = inv_29[0] ^ r_28[0] /*4367*/;
  assign sum_29[0] = _15218_ ^ oneWire /*4366*/;
  assign _15219_ = _15218_ & oneWire /*4365*/;
  assign _15220_ = inv_29[0] & r_28[0] /*4364*/;
  assign _15221_ = _15219_ | _15220_ /*4363*/;
  assign _15222_ = inv_29[1] ^ r_28[1] /*4361*/;
  assign sum_29[1] = _15222_ ^ _15221_ /*4360*/;
  assign _15223_ = _15222_ & _15221_ /*4359*/;
  assign _15224_ = inv_29[1] & r_28[1] /*4358*/;
  assign _15225_ = _15223_ | _15224_ /*4357*/;
  assign _15226_ = inv_29[2] ^ r_28[2] /*4355*/;
  assign sum_29[2] = _15226_ ^ _15225_ /*4354*/;
  assign _15227_ = _15226_ & _15225_ /*4353*/;
  assign _15228_ = inv_29[2] & r_28[2] /*4352*/;
  assign _15229_ = _15227_ | _15228_ /*4351*/;
  assign _15230_ = inv_29[3] ^ r_28[3] /*4349*/;
  assign sum_29[3] = _15230_ ^ _15229_ /*4348*/;
  assign _15231_ = _15230_ & _15229_ /*4347*/;
  assign _15232_ = inv_29[3] & r_28[3] /*4346*/;
  assign _15233_ = _15231_ | _15232_ /*4345*/;
  assign _15234_ = inv_29[4] ^ r_28[4] /*4343*/;
  assign sum_29[4] = _15234_ ^ _15233_ /*4342*/;
  assign _15235_ = _15234_ & _15233_ /*4341*/;
  assign _15236_ = inv_29[4] & r_28[4] /*4340*/;
  assign _15237_ = _15235_ | _15236_ /*4339*/;
  assign _15238_ = inv_29[5] ^ r_28[5] /*4337*/;
  assign sum_29[5] = _15238_ ^ _15237_ /*4336*/;
  assign _15239_ = _15238_ & _15237_ /*4335*/;
  assign _15240_ = inv_29[5] & r_28[5] /*4334*/;
  assign _15241_ = _15239_ | _15240_ /*4333*/;
  assign _15242_ = inv_29[6] ^ r_28[6] /*4331*/;
  assign sum_29[6] = _15242_ ^ _15241_ /*4330*/;
  assign _15243_ = _15242_ & _15241_ /*4329*/;
  assign _15244_ = inv_29[6] & r_28[6] /*4328*/;
  assign _15245_ = _15243_ | _15244_ /*4327*/;
  assign _15246_ = inv_29[7] ^ r_28[7] /*4325*/;
  assign sum_29[7] = _15246_ ^ _15245_ /*4324*/;
  assign _15247_ = _15246_ & _15245_ /*4323*/;
  assign _15248_ = inv_29[7] & r_28[7] /*4322*/;
  assign _15249_ = _15247_ | _15248_ /*4321*/;
  assign _15250_ = inv_29[8] ^ r_28[8] /*4319*/;
  assign sum_29[8] = _15250_ ^ _15249_ /*4318*/;
  assign _15251_ = _15250_ & _15249_ /*4317*/;
  assign _15252_ = inv_29[8] & r_28[8] /*4316*/;
  assign _15253_ = _15251_ | _15252_ /*4315*/;
  assign _15254_ = inv_29[9] ^ r_28[9] /*4313*/;
  assign sum_29[9] = _15254_ ^ _15253_ /*4312*/;
  assign _15255_ = _15254_ & _15253_ /*4311*/;
  assign _15256_ = inv_29[9] & r_28[9] /*4310*/;
  assign _15257_ = _15255_ | _15256_ /*4309*/;
  assign _15258_ = inv_29[10] ^ r_28[10] /*4307*/;
  assign sum_29[10] = _15258_ ^ _15257_ /*4306*/;
  assign _15259_ = _15258_ & _15257_ /*4305*/;
  assign _15260_ = inv_29[10] & r_28[10] /*4304*/;
  assign _15261_ = _15259_ | _15260_ /*4303*/;
  assign _15262_ = inv_29[11] ^ r_28[11] /*4301*/;
  assign sum_29[11] = _15262_ ^ _15261_ /*4300*/;
  assign _15263_ = _15262_ & _15261_ /*4299*/;
  assign _15264_ = inv_29[11] & r_28[11] /*4298*/;
  assign _15265_ = _15263_ | _15264_ /*4297*/;
  assign _15266_ = inv_29[12] ^ r_28[12] /*4295*/;
  assign sum_29[12] = _15266_ ^ _15265_ /*4294*/;
  assign _15267_ = _15266_ & _15265_ /*4293*/;
  assign _15268_ = inv_29[12] & r_28[12] /*4292*/;
  assign _15269_ = _15267_ | _15268_ /*4291*/;
  assign _15270_ = inv_29[13] ^ r_28[13] /*4289*/;
  assign sum_29[13] = _15270_ ^ _15269_ /*4288*/;
  assign _15271_ = _15270_ & _15269_ /*4287*/;
  assign _15272_ = inv_29[13] & r_28[13] /*4286*/;
  assign _15273_ = _15271_ | _15272_ /*4285*/;
  assign _15274_ = inv_29[14] ^ r_28[14] /*4283*/;
  assign sum_29[14] = _15274_ ^ _15273_ /*4282*/;
  assign _15275_ = _15274_ & _15273_ /*4281*/;
  assign _15276_ = inv_29[14] & r_28[14] /*4280*/;
  assign _15277_ = _15275_ | _15276_ /*4279*/;
  assign _15278_ = inv_29[15] ^ r_28[15] /*4277*/;
  assign sum_29[15] = _15278_ ^ _15277_ /*4276*/;
  assign _15279_ = _15278_ & _15277_ /*4275*/;
  assign _15280_ = inv_29[15] & r_28[15] /*4274*/;
  assign _15281_ = _15279_ | _15280_ /*4273*/;
  assign _15282_ = inv_29[16] ^ r_28[16] /*4271*/;
  assign sum_29[16] = _15282_ ^ _15281_ /*4270*/;
  assign _15283_ = _15282_ & _15281_ /*4269*/;
  assign _15284_ = inv_29[16] & r_28[16] /*4268*/;
  assign _15285_ = _15283_ | _15284_ /*4267*/;
  assign _15286_ = inv_29[17] ^ r_28[17] /*4265*/;
  assign sum_29[17] = _15286_ ^ _15285_ /*4264*/;
  assign _15287_ = _15286_ & _15285_ /*4263*/;
  assign _15288_ = inv_29[17] & r_28[17] /*4262*/;
  assign _15289_ = _15287_ | _15288_ /*4261*/;
  assign _15290_ = inv_29[18] ^ r_28[18] /*4259*/;
  assign sum_29[18] = _15290_ ^ _15289_ /*4258*/;
  assign _15291_ = _15290_ & _15289_ /*4257*/;
  assign _15292_ = inv_29[18] & r_28[18] /*4256*/;
  assign _15293_ = _15291_ | _15292_ /*4255*/;
  assign _15294_ = inv_29[19] ^ r_28[19] /*4253*/;
  assign sum_29[19] = _15294_ ^ _15293_ /*4252*/;
  assign _15295_ = _15294_ & _15293_ /*4251*/;
  assign _15296_ = inv_29[19] & r_28[19] /*4250*/;
  assign _15297_ = _15295_ | _15296_ /*4249*/;
  assign _15298_ = inv_29[20] ^ r_28[20] /*4247*/;
  assign sum_29[20] = _15298_ ^ _15297_ /*4246*/;
  assign _15299_ = _15298_ & _15297_ /*4245*/;
  assign _15300_ = inv_29[20] & r_28[20] /*4244*/;
  assign _15301_ = _15299_ | _15300_ /*4243*/;
  assign _15302_ = inv_29[21] ^ r_28[21] /*4241*/;
  assign sum_29[21] = _15302_ ^ _15301_ /*4240*/;
  assign _15303_ = _15302_ & _15301_ /*4239*/;
  assign _15304_ = inv_29[21] & r_28[21] /*4238*/;
  assign _15305_ = _15303_ | _15304_ /*4237*/;
  assign _15306_ = inv_29[22] ^ r_28[22] /*4235*/;
  assign sum_29[22] = _15306_ ^ _15305_ /*4234*/;
  assign _15307_ = _15306_ & _15305_ /*4233*/;
  assign _15308_ = inv_29[22] & r_28[22] /*4232*/;
  assign _15309_ = _15307_ | _15308_ /*4231*/;
  assign _15310_ = inv_29[23] ^ r_28[23] /*4229*/;
  assign sum_29[23] = _15310_ ^ _15309_ /*4228*/;
  assign _15311_ = _15310_ & _15309_ /*4227*/;
  assign _15312_ = inv_29[23] & r_28[23] /*4226*/;
  assign _15313_ = _15311_ | _15312_ /*4225*/;
  assign _15314_ = inv_29[24] ^ r_28[24] /*4223*/;
  assign sum_29[24] = _15314_ ^ _15313_ /*4222*/;
  assign _15315_ = _15314_ & _15313_ /*4221*/;
  assign _15316_ = inv_29[24] & r_28[24] /*4220*/;
  assign _15317_ = _15315_ | _15316_ /*4219*/;
  assign _15318_ = inv_29[25] ^ r_28[25] /*4217*/;
  assign sum_29[25] = _15318_ ^ _15317_ /*4216*/;
  assign _15319_ = _15318_ & _15317_ /*4215*/;
  assign _15320_ = inv_29[25] & r_28[25] /*4214*/;
  assign _15321_ = _15319_ | _15320_ /*4213*/;
  assign _15322_ = inv_29[26] ^ r_28[26] /*4211*/;
  assign sum_29[26] = _15322_ ^ _15321_ /*4210*/;
  assign _15323_ = _15322_ & _15321_ /*4209*/;
  assign _15324_ = inv_29[26] & r_28[26] /*4208*/;
  assign _15325_ = _15323_ | _15324_ /*4207*/;
  assign _15326_ = inv_29[27] ^ r_28[27] /*4205*/;
  assign sum_29[27] = _15326_ ^ _15325_ /*4204*/;
  assign _15327_ = _15326_ & _15325_ /*4203*/;
  assign _15328_ = inv_29[27] & r_28[27] /*4202*/;
  assign _15329_ = _15327_ | _15328_ /*4201*/;
  assign _15330_ = inv_29[28] ^ r_28[28] /*4199*/;
  assign sum_29[28] = _15330_ ^ _15329_ /*4198*/;
  assign _15331_ = _15330_ & _15329_ /*4197*/;
  assign _15332_ = inv_29[28] & r_28[28] /*4196*/;
  assign _15333_ = _15331_ | _15332_ /*4195*/;
  assign _15334_ = inv_29[29] ^ r_28[29] /*4193*/;
  assign sum_29[29] = _15334_ ^ _15333_ /*4192*/;
  assign _15335_ = _15334_ & _15333_ /*4191*/;
  assign _15336_ = inv_29[29] & r_28[29] /*4190*/;
  assign _15337_ = _15335_ | _15336_ /*4189*/;
  assign _15338_ = inv_29[30] ^ r_28[30] /*4187*/;
  assign sum_29[30] = _15338_ ^ _15337_ /*4186*/;
  assign _15339_ = _15338_ & _15337_ /*4185*/;
  assign _15340_ = inv_29[30] & r_28[30] /*4184*/;
  assign _15341_ = _15339_ | _15340_ /*4183*/;
  assign _15342_ = inv_29[31] ^ r_28[31] /*4181*/;
  assign sum_29[31] = _15342_ ^ _15341_ /*4180*/;
  assign _15343_ = _15342_ & _15341_ /*4179*/;
  assign _15344_ = inv_29[31] & r_28[31] /*4178*/;
  assign _15345_ = _15343_ | _15344_ /*4177*/;
  assign _15346_ = inv_29[32] ^ r_28[32] /*4175*/;
  assign sum_29[32] = _15346_ ^ _15345_ /*4174*/;
  assign _15347_ = _15346_ & _15345_ /*4173*/;
  assign _15348_ = inv_29[32] & r_28[32] /*4172*/;
  assign _15349_ = _15347_ | _15348_ /*4171*/;
  assign _15350_ = inv_29[33] ^ r_28[33] /*4169*/;
  assign sum_29[33] = _15350_ ^ _15349_ /*4168*/;
  assign _15351_ = _15350_ & _15349_ /*4167*/;
  assign _15352_ = inv_29[33] & r_28[33] /*4166*/;
  assign _15353_ = _15351_ | _15352_ /*4165*/;
  assign _15354_ = inv_29[34] ^ r_28[34] /*4163*/;
  assign sum_29[34] = _15354_ ^ _15353_ /*4162*/;
  assign _15355_ = _15354_ & _15353_ /*4161*/;
  assign _15356_ = inv_29[34] & r_28[34] /*4160*/;
  assign _15357_ = _15355_ | _15356_ /*4159*/;
  assign _15358_ = inv_29[35] ^ r_28[35] /*4157*/;
  assign sum_29[35] = _15358_ ^ _15357_ /*4156*/;
  assign _15359_ = _15358_ & _15357_ /*4155*/;
  assign _15360_ = inv_29[35] & r_28[35] /*4154*/;
  assign _15361_ = _15359_ | _15360_ /*4153*/;
  assign _15362_ = inv_29[36] ^ r_28[36] /*4151*/;
  assign sum_29[36] = _15362_ ^ _15361_ /*4150*/;
  assign _15363_ = _15362_ & _15361_ /*4149*/;
  assign _15364_ = inv_29[36] & r_28[36] /*4148*/;
  assign _15365_ = _15363_ | _15364_ /*4147*/;
  assign _15366_ = inv_29[37] ^ r_28[37] /*4145*/;
  assign sum_29[37] = _15366_ ^ _15365_ /*4144*/;
  assign _15367_ = _15366_ & _15365_ /*4143*/;
  assign _15368_ = inv_29[37] & r_28[37] /*4142*/;
  assign _15369_ = _15367_ | _15368_ /*4141*/;
  assign _15370_ = inv_29[38] ^ r_28[38] /*4139*/;
  assign sum_29[38] = _15370_ ^ _15369_ /*4138*/;
  assign _15371_ = _15370_ & _15369_ /*4137*/;
  assign _15372_ = inv_29[38] & r_28[38] /*4136*/;
  assign _15373_ = _15371_ | _15372_ /*4135*/;
  assign _15374_ = inv_29[39] ^ r_28[39] /*4133*/;
  assign sum_29[39] = _15374_ ^ _15373_ /*4132*/;
  assign _15375_ = _15374_ & _15373_ /*4131*/;
  assign _15376_ = inv_29[39] & r_28[39] /*4130*/;
  assign _15377_ = _15375_ | _15376_ /*4129*/;
  assign _15378_ = inv_29[40] ^ r_28[40] /*4127*/;
  assign sum_29[40] = _15378_ ^ _15377_ /*4126*/;
  assign _15379_ = _15378_ & _15377_ /*4125*/;
  assign _15380_ = inv_29[40] & r_28[40] /*4124*/;
  assign _15381_ = _15379_ | _15380_ /*4123*/;
  assign _15382_ = inv_29[41] ^ r_28[41] /*4121*/;
  assign sum_29[41] = _15382_ ^ _15381_ /*4120*/;
  assign _15383_ = _15382_ & _15381_ /*4119*/;
  assign _15384_ = inv_29[41] & r_28[41] /*4118*/;
  assign _15385_ = _15383_ | _15384_ /*4117*/;
  assign _15386_ = inv_29[42] ^ r_28[42] /*4115*/;
  assign sum_29[42] = _15386_ ^ _15385_ /*4114*/;
  assign _15387_ = _15386_ & _15385_ /*4113*/;
  assign _15388_ = inv_29[42] & r_28[42] /*4112*/;
  assign _15389_ = _15387_ | _15388_ /*4111*/;
  assign _15390_ = inv_29[43] ^ r_28[43] /*4109*/;
  assign sum_29[43] = _15390_ ^ _15389_ /*4108*/;
  assign _15391_ = _15390_ & _15389_ /*4107*/;
  assign _15392_ = inv_29[43] & r_28[43] /*4106*/;
  assign _15393_ = _15391_ | _15392_ /*4105*/;
  assign _15394_ = inv_29[44] ^ r_28[44] /*4103*/;
  assign sum_29[44] = _15394_ ^ _15393_ /*4102*/;
  assign _15395_ = _15394_ & _15393_ /*4101*/;
  assign _15396_ = inv_29[44] & r_28[44] /*4100*/;
  assign _15397_ = _15395_ | _15396_ /*4099*/;
  assign _15398_ = inv_29[45] ^ r_28[45] /*4097*/;
  assign sum_29[45] = _15398_ ^ _15397_ /*4096*/;
  assign _15399_ = _15398_ & _15397_ /*4095*/;
  assign _15400_ = inv_29[45] & r_28[45] /*4094*/;
  assign _15401_ = _15399_ | _15400_ /*4093*/;
  assign _15402_ = inv_29[46] ^ r_28[46] /*4091*/;
  assign sum_29[46] = _15402_ ^ _15401_ /*4090*/;
  assign _15403_ = _15402_ & _15401_ /*4089*/;
  assign _15404_ = inv_29[46] & r_28[46] /*4088*/;
  assign _15405_ = _15403_ | _15404_ /*4087*/;
  assign _15406_ = inv_29[47] ^ r_28[47] /*4085*/;
  assign sum_29[47] = _15406_ ^ _15405_ /*4084*/;
  assign _15407_ = _15406_ & _15405_ /*4083*/;
  assign _15408_ = inv_29[47] & r_28[47] /*4082*/;
  assign _15409_ = _15407_ | _15408_ /*4081*/;
  assign _15410_ = inv_29[48] ^ r_28[48] /*4079*/;
  assign sum_29[48] = _15410_ ^ _15409_ /*4078*/;
  assign _15411_ = _15410_ & _15409_ /*4077*/;
  assign _15412_ = inv_29[48] & r_28[48] /*4076*/;
  assign _15413_ = _15411_ | _15412_ /*4075*/;
  assign _15414_ = inv_29[49] ^ r_28[49] /*4073*/;
  assign sum_29[49] = _15414_ ^ _15413_ /*4072*/;
  assign _15415_ = _15414_ & _15413_ /*4071*/;
  assign _15416_ = inv_29[49] & r_28[49] /*4070*/;
  assign _15417_ = _15415_ | _15416_ /*4069*/;
  assign _15418_ = inv_29[50] ^ r_28[50] /*4067*/;
  assign sum_29[50] = _15418_ ^ _15417_ /*4066*/;
  assign _15419_ = _15418_ & _15417_ /*4065*/;
  assign _15420_ = inv_29[50] & r_28[50] /*4064*/;
  assign _15421_ = _15419_ | _15420_ /*4063*/;
  assign _15422_ = inv_29[51] ^ r_28[51] /*4061*/;
  assign sum_29[51] = _15422_ ^ _15421_ /*4060*/;
  assign _15423_ = _15422_ & _15421_ /*4059*/;
  assign _15424_ = inv_29[51] & r_28[51] /*4058*/;
  assign _15425_ = _15423_ | _15424_ /*4057*/;
  assign _15426_ = inv_29[52] ^ r_28[52] /*4055*/;
  assign sum_29[52] = _15426_ ^ _15425_ /*4054*/;
  assign _15427_ = _15426_ & _15425_ /*4053*/;
  assign _15428_ = inv_29[52] & r_28[52] /*4052*/;
  assign _15429_ = _15427_ | _15428_ /*4051*/;
  assign _15430_ = inv_29[53] ^ r_28[53] /*4049*/;
  assign sum_29[53] = _15430_ ^ _15429_ /*4048*/;
  assign _15431_ = _15430_ & _15429_ /*4047*/;
  assign _15432_ = inv_29[53] & r_28[53] /*4046*/;
  assign _15433_ = _15431_ | _15432_ /*4045*/;
  assign _15434_ = inv_29[54] ^ r_28[54] /*4043*/;
  assign sum_29[54] = _15434_ ^ _15433_ /*4042*/;
  assign _15435_ = _15434_ & _15433_ /*4041*/;
  assign _15436_ = inv_29[54] & r_28[54] /*4040*/;
  assign _15437_ = _15435_ | _15436_ /*4039*/;
  assign _15438_ = inv_29[55] ^ r_28[55] /*4037*/;
  assign sum_29[55] = _15438_ ^ _15437_ /*4036*/;
  assign _15439_ = _15438_ & _15437_ /*4035*/;
  assign _15440_ = inv_29[55] & r_28[55] /*4034*/;
  assign _15441_ = _15439_ | _15440_ /*4033*/;
  assign _15442_ = inv_29[56] ^ r_28[56] /*4031*/;
  assign sum_29[56] = _15442_ ^ _15441_ /*4030*/;
  assign _15443_ = _15442_ & _15441_ /*4029*/;
  assign _15444_ = inv_29[56] & r_28[56] /*4028*/;
  assign _15445_ = _15443_ | _15444_ /*4027*/;
  assign _15446_ = inv_29[57] ^ r_28[57] /*4025*/;
  assign sum_29[57] = _15446_ ^ _15445_ /*4024*/;
  assign _15447_ = _15446_ & _15445_ /*4023*/;
  assign _15448_ = inv_29[57] & r_28[57] /*4022*/;
  assign _15449_ = _15447_ | _15448_ /*4021*/;
  assign _15450_ = inv_29[58] ^ r_28[58] /*4019*/;
  assign sum_29[58] = _15450_ ^ _15449_ /*4018*/;
  assign _15451_ = _15450_ & _15449_ /*4017*/;
  assign _15452_ = inv_29[58] & r_28[58] /*4016*/;
  assign _15453_ = _15451_ | _15452_ /*4015*/;
  assign _15454_ = inv_29[59] ^ r_28[59] /*4013*/;
  assign sum_29[59] = _15454_ ^ _15453_ /*4012*/;
  assign _15455_ = _15454_ & _15453_ /*4011*/;
  assign _15456_ = inv_29[59] & r_28[59] /*4010*/;
  assign _15457_ = _15455_ | _15456_ /*4009*/;
  assign _15458_ = inv_29[60] ^ r_28[60] /*4007*/;
  assign sum_29[60] = _15458_ ^ _15457_ /*4006*/;
  assign _15459_ = _15458_ & _15457_ /*4005*/;
  assign _15460_ = inv_29[60] & r_28[60] /*4004*/;
  assign _15461_ = _15459_ | _15460_ /*4003*/;
  assign _15462_ = inv_29[61] ^ r_28[61] /*4001*/;
  assign sum_29[61] = _15462_ ^ _15461_ /*4000*/;
  assign _15463_ = _15462_ & _15461_ /*3999*/;
  assign _15464_ = inv_29[61] & r_28[61] /*3998*/;
  assign _15465_ = _15463_ | _15464_ /*3997*/;
  assign _15466_ = inv_29[62] ^ r_28[62] /*3995*/;
  assign sum_29[62] = _15466_ ^ _15465_ /*3994*/;
  assign _15467_ = _15466_ & _15465_ /*3993*/;
  assign _15468_ = inv_29[62] & r_28[62] /*3992*/;
  assign _15469_ = _15467_ | _15468_ /*3991*/;
  assign _15470_ = inv_29[63] ^ r_28[63] /*3989*/;
  assign sum_29[63] = _15470_ ^ _15469_ /*3988*/;
  assign _15471_ = _15470_ & _15469_ /*3987*/;
  assign _15472_ = inv_29[63] & r_28[63] /*3986*/;
  assign _15473_ = _15471_ | _15472_ /*3985*/;
  assign _15474_ = inv_29[64] ^ r_28[64] /*3983*/;
  assign sum_29[64] = _15474_ ^ _15473_ /*3982*/;
  assign _15475_ = _15474_ & _15473_ /*3981*/;
  assign _15476_ = inv_29[64] & r_28[64] /*3980*/;
  assign _15477_ = _15475_ | _15476_ /*3979*/;
  assign _15478_ = inv_29[65] ^ r_28[65] /*3977*/;
  assign sum_29[65] = _15478_ ^ _15477_ /*3976*/;
  assign _15479_ = _15478_ & _15477_ /*3975*/;
  assign _15480_ = inv_29[65] & r_28[65] /*3974*/;
  assign _15481_ = _15479_ | _15480_ /*3973*/;
  assign _15482_ = inv_29[66] ^ r_28[66] /*3971*/;
  assign sum_29[66] = _15482_ ^ _15481_ /*3970*/;
  assign _15483_ = _15482_ & _15481_ /*3969*/;
  assign _15484_ = inv_29[66] & r_28[66] /*3968*/;
  assign _15485_ = _15483_ | _15484_ /*3967*/;
  assign _15486_ = inv_29[67] ^ r_28[67] /*3965*/;
  assign sum_29[67] = _15486_ ^ _15485_ /*3964*/;
  assign _15487_ = _15486_ & _15485_ /*3963*/;
  assign _15488_ = inv_29[67] & r_28[67] /*3962*/;
  assign _15489_ = _15487_ | _15488_ /*3961*/;
  assign _15490_ = inv_29[68] ^ r_28[68] /*3959*/;
  assign sum_29[68] = _15490_ ^ _15489_ /*3958*/;
  assign _15491_ = _15490_ & _15489_ /*3957*/;
  assign _15492_ = inv_29[68] & r_28[68] /*3956*/;
  assign _15493_ = _15491_ | _15492_ /*3955*/;
  assign _15494_ = inv_29[69] ^ r_28[69] /*3953*/;
  assign sum_29[69] = _15494_ ^ _15493_ /*3952*/;
  assign _15495_ = _15494_ & _15493_ /*3951*/;
  assign _15496_ = inv_29[69] & r_28[69] /*3950*/;
  assign _15497_ = _15495_ | _15496_ /*3949*/;
  assign _15498_ = inv_29[70] ^ r_28[70] /*3947*/;
  assign sum_29[70] = _15498_ ^ _15497_ /*3946*/;
  assign _15499_ = _15498_ & _15497_ /*3945*/;
  assign _15500_ = inv_29[70] & r_28[70] /*3944*/;
  assign _15501_ = _15499_ | _15500_ /*3943*/;
  assign _15502_ = inv_29[71] ^ r_28[71] /*3941*/;
  assign sum_29[71] = _15502_ ^ _15501_ /*3940*/;
  assign _15503_ = _15502_ & _15501_ /*3939*/;
  assign _15504_ = inv_29[71] & r_28[71] /*3938*/;
  assign _15505_ = _15503_ | _15504_ /*3937*/;
  assign _15506_ = inv_29[72] ^ r_28[72] /*3935*/;
  assign sum_29[72] = _15506_ ^ _15505_ /*3934*/;
  assign _15507_ = _15506_ & _15505_ /*3933*/;
  assign _15508_ = inv_29[72] & r_28[72] /*3932*/;
  assign _15509_ = _15507_ | _15508_ /*3931*/;
  assign _15510_ = inv_29[73] ^ r_28[73] /*3929*/;
  assign sum_29[73] = _15510_ ^ _15509_ /*3928*/;
  assign _15511_ = _15510_ & _15509_ /*3927*/;
  assign _15512_ = inv_29[73] & r_28[73] /*3926*/;
  assign _15513_ = _15511_ | _15512_ /*3925*/;
  assign _15514_ = inv_29[74] ^ r_28[74] /*3923*/;
  assign sum_29[74] = _15514_ ^ _15513_ /*3922*/;
  assign _15515_ = _15514_ & _15513_ /*3921*/;
  assign _15516_ = inv_29[74] & r_28[74] /*3920*/;
  assign _15517_ = _15515_ | _15516_ /*3919*/;
  assign _15518_ = inv_29[75] ^ r_28[75] /*3917*/;
  assign sum_29[75] = _15518_ ^ _15517_ /*3916*/;
  assign _15519_ = _15518_ & _15517_ /*3915*/;
  assign _15520_ = inv_29[75] & r_28[75] /*3914*/;
  assign _15521_ = _15519_ | _15520_ /*3913*/;
  assign _15522_ = inv_29[76] ^ r_28[76] /*3911*/;
  assign sum_29[76] = _15522_ ^ _15521_ /*3910*/;
  assign _15523_ = _15522_ & _15521_ /*3909*/;
  assign _15524_ = inv_29[76] & r_28[76] /*3908*/;
  assign _15525_ = _15523_ | _15524_ /*3907*/;
  assign _15526_ = inv_29[77] ^ r_28[77] /*3905*/;
  assign sum_29[77] = _15526_ ^ _15525_ /*3904*/;
  assign _15527_ = _15526_ & _15525_ /*3903*/;
  assign _15528_ = inv_29[77] & r_28[77] /*3902*/;
  assign _15529_ = _15527_ | _15528_ /*3901*/;
  assign _15530_ = inv_29[78] ^ r_28[78] /*3899*/;
  assign sum_29[78] = _15530_ ^ _15529_ /*3898*/;
  assign _15531_ = _15530_ & _15529_ /*3897*/;
  assign _15532_ = inv_29[78] & r_28[78] /*3896*/;
  assign _15533_ = _15531_ | _15532_ /*3895*/;
  assign _15534_ = inv_29[79] ^ r_28[79] /*3893*/;
  assign sum_29[79] = _15534_ ^ _15533_ /*3892*/;
  assign _15535_ = _15534_ & _15533_ /*3891*/;
  assign _15536_ = inv_29[79] & r_28[79] /*3890*/;
  assign _15537_ = _15535_ | _15536_ /*3889*/;
  assign _15538_ = inv_29[80] ^ r_28[80] /*3887*/;
  assign sum_29[80] = _15538_ ^ _15537_ /*3886*/;
  assign _15539_ = _15538_ & _15537_ /*3885*/;
  assign _15540_ = inv_29[80] & r_28[80] /*3884*/;
  assign _15541_ = _15539_ | _15540_ /*3883*/;
  assign _15542_ = inv_29[81] ^ r_28[81] /*3881*/;
  assign sum_29[81] = _15542_ ^ _15541_ /*3880*/;
  assign _15543_ = _15542_ & _15541_ /*3879*/;
  assign _15544_ = inv_29[81] & r_28[81] /*3878*/;
  assign _15545_ = _15543_ | _15544_ /*3877*/;
  assign _15546_ = inv_29[82] ^ r_28[82] /*3875*/;
  assign sum_29[82] = _15546_ ^ _15545_ /*3874*/;
  assign _15547_ = _15546_ & _15545_ /*3873*/;
  assign _15548_ = inv_29[82] & r_28[82] /*3872*/;
  assign _15549_ = _15547_ | _15548_ /*3871*/;
  assign _15550_ = inv_29[83] ^ r_28[83] /*3869*/;
  assign sum_29[83] = _15550_ ^ _15549_ /*3868*/;
  assign _15551_ = _15550_ & _15549_ /*3867*/;
  assign _15552_ = inv_29[83] & r_28[83] /*3866*/;
  assign _15553_ = _15551_ | _15552_ /*3865*/;
  assign _15554_ = inv_29[84] ^ r_28[84] /*3863*/;
  assign sum_29[84] = _15554_ ^ _15553_ /*3862*/;
  assign _15555_ = _15554_ & _15553_ /*3861*/;
  assign _15556_ = inv_29[84] & r_28[84] /*3860*/;
  assign _15557_ = _15555_ | _15556_ /*3859*/;
  assign _15558_ = inv_29[85] ^ r_28[85] /*3857*/;
  assign sum_29[85] = _15558_ ^ _15557_ /*3856*/;
  assign _15559_ = _15558_ & _15557_ /*3855*/;
  assign _15560_ = inv_29[85] & r_28[85] /*3854*/;
  assign _15561_ = _15559_ | _15560_ /*3853*/;
  assign _15562_ = inv_29[86] ^ r_28[86] /*3851*/;
  assign sum_29[86] = _15562_ ^ _15561_ /*3850*/;
  assign _15563_ = _15562_ & _15561_ /*3849*/;
  assign _15564_ = inv_29[86] & r_28[86] /*3848*/;
  assign _15565_ = _15563_ | _15564_ /*3847*/;
  assign _15566_ = inv_29[87] ^ r_28[87] /*3845*/;
  assign sum_29[87] = _15566_ ^ _15565_ /*3844*/;
  assign _15567_ = _15566_ & _15565_ /*3843*/;
  assign _15568_ = inv_29[87] & r_28[87] /*3842*/;
  assign _15569_ = _15567_ | _15568_ /*3841*/;
  assign _15570_ = inv_29[88] ^ r_28[88] /*3839*/;
  assign sum_29[88] = _15570_ ^ _15569_ /*3838*/;
  assign _15571_ = _15570_ & _15569_ /*3837*/;
  assign _15572_ = inv_29[88] & r_28[88] /*3836*/;
  assign _15573_ = _15571_ | _15572_ /*3835*/;
  assign _15574_ = inv_29[89] ^ r_28[89] /*3833*/;
  assign sum_29[89] = _15574_ ^ _15573_ /*3832*/;
  assign _15575_ = _15574_ & _15573_ /*3831*/;
  assign _15576_ = inv_29[89] & r_28[89] /*3830*/;
  assign _15577_ = _15575_ | _15576_ /*3829*/;
  assign _15578_ = inv_29[90] ^ r_28[90] /*3827*/;
  assign sum_29[90] = _15578_ ^ _15577_ /*3826*/;
  assign _15579_ = _15578_ & _15577_ /*3825*/;
  assign _15580_ = inv_29[90] & r_28[90] /*3824*/;
  assign _15581_ = _15579_ | _15580_ /*3823*/;
  assign _15582_ = _15581_ ^ _15577_ /*3822*/;
  assign _15583_ = ~_15582_ /*3821*/;
  assign _15584_ = sum_29[90] & _15583_ /*3820*/;
  assign _15585_ = _15582_ & _15581_ /*3819*/;
  assign sum_29[91] = _15585_ | _15584_ /*3818*/;
  assign q[3] = ~sum_29[91] /*3817*/;
  assign m_29[0] = r_28[0] /*3816*/;
  assign m_29[1] = r_28[1] /*3815*/;
  assign m_29[2] = r_28[2] /*3814*/;
  assign m_29[3] = r_28[3] /*3813*/;
  assign m_29[4] = r_28[4] /*3812*/;
  assign m_29[5] = r_28[5] /*3811*/;
  assign m_29[6] = r_28[6] /*3810*/;
  assign m_29[7] = r_28[7] /*3809*/;
  assign m_29[8] = r_28[8] /*3808*/;
  assign m_29[9] = r_28[9] /*3807*/;
  assign m_29[10] = r_28[10] /*3806*/;
  assign m_29[11] = r_28[11] /*3805*/;
  assign m_29[12] = r_28[12] /*3804*/;
  assign m_29[13] = r_28[13] /*3803*/;
  assign m_29[14] = r_28[14] /*3802*/;
  assign m_29[15] = r_28[15] /*3801*/;
  assign m_29[16] = r_28[16] /*3800*/;
  assign m_29[17] = r_28[17] /*3799*/;
  assign m_29[18] = r_28[18] /*3798*/;
  assign m_29[19] = r_28[19] /*3797*/;
  assign m_29[20] = r_28[20] /*3796*/;
  assign m_29[21] = r_28[21] /*3795*/;
  assign m_29[22] = r_28[22] /*3794*/;
  assign m_29[23] = r_28[23] /*3793*/;
  assign m_29[24] = r_28[24] /*3792*/;
  assign m_29[25] = r_28[25] /*3791*/;
  assign m_29[26] = r_28[26] /*3790*/;
  assign m_29[27] = r_28[27] /*3789*/;
  assign m_29[28] = r_28[28] /*3788*/;
  assign m_29[29] = r_28[29] /*3787*/;
  assign m_29[30] = r_28[30] /*3786*/;
  assign m_29[31] = r_28[31] /*3785*/;
  assign m_29[32] = r_28[32] /*3784*/;
  assign m_29[33] = r_28[33] /*3783*/;
  assign m_29[34] = r_28[34] /*3782*/;
  assign m_29[35] = r_28[35] /*3781*/;
  assign m_29[36] = r_28[36] /*3780*/;
  assign m_29[37] = r_28[37] /*3779*/;
  assign m_29[38] = r_28[38] /*3778*/;
  assign m_29[39] = r_28[39] /*3777*/;
  assign m_29[40] = r_28[40] /*3776*/;
  assign m_29[41] = r_28[41] /*3775*/;
  assign m_29[42] = r_28[42] /*3774*/;
  assign m_29[43] = r_28[43] /*3773*/;
  assign m_29[44] = r_28[44] /*3772*/;
  assign m_29[45] = r_28[45] /*3771*/;
  assign m_29[46] = r_28[46] /*3770*/;
  assign m_29[47] = r_28[47] /*3769*/;
  assign m_29[48] = r_28[48] /*3768*/;
  assign m_29[49] = r_28[49] /*3767*/;
  assign m_29[50] = r_28[50] /*3766*/;
  assign m_29[51] = r_28[51] /*3765*/;
  assign m_29[52] = r_28[52] /*3764*/;
  assign m_29[53] = r_28[53] /*3763*/;
  assign m_29[54] = r_28[54] /*3762*/;
  assign m_29[55] = r_28[55] /*3761*/;
  assign m_29[56] = r_28[56] /*3760*/;
  assign m_29[57] = r_28[57] /*3759*/;
  assign m_29[58] = r_28[58] /*3758*/;
  assign m_29[59] = r_28[59] /*3757*/;
  assign m_29[60] = r_28[60] /*3756*/;
  assign m_29[61] = r_28[61] /*3755*/;
  assign m_29[62] = r_28[62] /*3754*/;
  assign m_29[63] = r_28[63] /*3753*/;
  assign m_29[64] = r_28[64] /*3752*/;
  assign m_29[65] = r_28[65] /*3751*/;
  assign m_29[66] = r_28[66] /*3750*/;
  assign m_29[67] = r_28[67] /*3749*/;
  assign m_29[68] = r_28[68] /*3748*/;
  assign m_29[69] = r_28[69] /*3747*/;
  assign m_29[70] = r_28[70] /*3746*/;
  assign m_29[71] = r_28[71] /*3745*/;
  assign m_29[72] = r_28[72] /*3744*/;
  assign m_29[73] = r_28[73] /*3743*/;
  assign m_29[74] = r_28[74] /*3742*/;
  assign m_29[75] = r_28[75] /*3741*/;
  assign m_29[76] = r_28[76] /*3740*/;
  assign m_29[77] = r_28[77] /*3739*/;
  assign m_29[78] = r_28[78] /*3738*/;
  assign m_29[79] = r_28[79] /*3737*/;
  assign m_29[80] = r_28[80] /*3736*/;
  assign m_29[81] = r_28[81] /*3735*/;
  assign m_29[82] = r_28[82] /*3734*/;
  assign m_29[83] = r_28[83] /*3733*/;
  assign m_29[84] = r_28[84] /*3732*/;
  assign m_29[85] = r_28[85] /*3731*/;
  assign m_29[86] = r_28[86] /*3730*/;
  assign m_29[87] = r_28[87] /*3729*/;
  assign m_29[88] = r_28[88] /*3728*/;
  assign m_29[89] = r_28[89] /*3727*/;
  assign m_29[90] = r_28[90] /*3726*/;
  assign m_29[91] = r_28[90] /*3725*/;
  assign _15587_ = ~q[3] /*3724*/;
  assign _15588_ = sum_29[0] & q[3] /*3723*/;
  assign _15589_ = m_29[0] & _15587_ /*3722*/;
  assign r_29[0] = _15589_ | _15588_ /*3721*/;
  assign _15590_ = ~q[3] /*3720*/;
  assign _15591_ = sum_29[1] & q[3] /*3719*/;
  assign _15592_ = m_29[1] & _15590_ /*3718*/;
  assign r_29[1] = _15592_ | _15591_ /*3717*/;
  assign _15593_ = ~q[3] /*3716*/;
  assign _15594_ = sum_29[2] & q[3] /*3715*/;
  assign _15595_ = m_29[2] & _15593_ /*3714*/;
  assign r_29[2] = _15595_ | _15594_ /*3713*/;
  assign _15596_ = ~q[3] /*3712*/;
  assign _15597_ = sum_29[3] & q[3] /*3711*/;
  assign _15598_ = m_29[3] & _15596_ /*3710*/;
  assign r_29[3] = _15598_ | _15597_ /*3709*/;
  assign _15599_ = ~q[3] /*3708*/;
  assign _15600_ = sum_29[4] & q[3] /*3707*/;
  assign _15601_ = m_29[4] & _15599_ /*3706*/;
  assign r_29[4] = _15601_ | _15600_ /*3705*/;
  assign _15602_ = ~q[3] /*3704*/;
  assign _15603_ = sum_29[5] & q[3] /*3703*/;
  assign _15604_ = m_29[5] & _15602_ /*3702*/;
  assign r_29[5] = _15604_ | _15603_ /*3701*/;
  assign _15605_ = ~q[3] /*3700*/;
  assign _15606_ = sum_29[6] & q[3] /*3699*/;
  assign _15607_ = m_29[6] & _15605_ /*3698*/;
  assign r_29[6] = _15607_ | _15606_ /*3697*/;
  assign _15608_ = ~q[3] /*3696*/;
  assign _15609_ = sum_29[7] & q[3] /*3695*/;
  assign _15610_ = m_29[7] & _15608_ /*3694*/;
  assign r_29[7] = _15610_ | _15609_ /*3693*/;
  assign _15611_ = ~q[3] /*3692*/;
  assign _15612_ = sum_29[8] & q[3] /*3691*/;
  assign _15613_ = m_29[8] & _15611_ /*3690*/;
  assign r_29[8] = _15613_ | _15612_ /*3689*/;
  assign _15614_ = ~q[3] /*3688*/;
  assign _15615_ = sum_29[9] & q[3] /*3687*/;
  assign _15616_ = m_29[9] & _15614_ /*3686*/;
  assign r_29[9] = _15616_ | _15615_ /*3685*/;
  assign _15617_ = ~q[3] /*3684*/;
  assign _15618_ = sum_29[10] & q[3] /*3683*/;
  assign _15619_ = m_29[10] & _15617_ /*3682*/;
  assign r_29[10] = _15619_ | _15618_ /*3681*/;
  assign _15620_ = ~q[3] /*3680*/;
  assign _15621_ = sum_29[11] & q[3] /*3679*/;
  assign _15622_ = m_29[11] & _15620_ /*3678*/;
  assign r_29[11] = _15622_ | _15621_ /*3677*/;
  assign _15623_ = ~q[3] /*3676*/;
  assign _15624_ = sum_29[12] & q[3] /*3675*/;
  assign _15625_ = m_29[12] & _15623_ /*3674*/;
  assign r_29[12] = _15625_ | _15624_ /*3673*/;
  assign _15626_ = ~q[3] /*3672*/;
  assign _15627_ = sum_29[13] & q[3] /*3671*/;
  assign _15628_ = m_29[13] & _15626_ /*3670*/;
  assign r_29[13] = _15628_ | _15627_ /*3669*/;
  assign _15629_ = ~q[3] /*3668*/;
  assign _15630_ = sum_29[14] & q[3] /*3667*/;
  assign _15631_ = m_29[14] & _15629_ /*3666*/;
  assign r_29[14] = _15631_ | _15630_ /*3665*/;
  assign _15632_ = ~q[3] /*3664*/;
  assign _15633_ = sum_29[15] & q[3] /*3663*/;
  assign _15634_ = m_29[15] & _15632_ /*3662*/;
  assign r_29[15] = _15634_ | _15633_ /*3661*/;
  assign _15635_ = ~q[3] /*3660*/;
  assign _15636_ = sum_29[16] & q[3] /*3659*/;
  assign _15637_ = m_29[16] & _15635_ /*3658*/;
  assign r_29[16] = _15637_ | _15636_ /*3657*/;
  assign _15638_ = ~q[3] /*3656*/;
  assign _15639_ = sum_29[17] & q[3] /*3655*/;
  assign _15640_ = m_29[17] & _15638_ /*3654*/;
  assign r_29[17] = _15640_ | _15639_ /*3653*/;
  assign _15641_ = ~q[3] /*3652*/;
  assign _15642_ = sum_29[18] & q[3] /*3651*/;
  assign _15643_ = m_29[18] & _15641_ /*3650*/;
  assign r_29[18] = _15643_ | _15642_ /*3649*/;
  assign _15644_ = ~q[3] /*3648*/;
  assign _15645_ = sum_29[19] & q[3] /*3647*/;
  assign _15646_ = m_29[19] & _15644_ /*3646*/;
  assign r_29[19] = _15646_ | _15645_ /*3645*/;
  assign _15647_ = ~q[3] /*3644*/;
  assign _15648_ = sum_29[20] & q[3] /*3643*/;
  assign _15649_ = m_29[20] & _15647_ /*3642*/;
  assign r_29[20] = _15649_ | _15648_ /*3641*/;
  assign _15650_ = ~q[3] /*3640*/;
  assign _15651_ = sum_29[21] & q[3] /*3639*/;
  assign _15652_ = m_29[21] & _15650_ /*3638*/;
  assign r_29[21] = _15652_ | _15651_ /*3637*/;
  assign _15653_ = ~q[3] /*3636*/;
  assign _15654_ = sum_29[22] & q[3] /*3635*/;
  assign _15655_ = m_29[22] & _15653_ /*3634*/;
  assign r_29[22] = _15655_ | _15654_ /*3633*/;
  assign _15656_ = ~q[3] /*3632*/;
  assign _15657_ = sum_29[23] & q[3] /*3631*/;
  assign _15658_ = m_29[23] & _15656_ /*3630*/;
  assign r_29[23] = _15658_ | _15657_ /*3629*/;
  assign _15659_ = ~q[3] /*3628*/;
  assign _15660_ = sum_29[24] & q[3] /*3627*/;
  assign _15661_ = m_29[24] & _15659_ /*3626*/;
  assign r_29[24] = _15661_ | _15660_ /*3625*/;
  assign _15662_ = ~q[3] /*3624*/;
  assign _15663_ = sum_29[25] & q[3] /*3623*/;
  assign _15664_ = m_29[25] & _15662_ /*3622*/;
  assign r_29[25] = _15664_ | _15663_ /*3621*/;
  assign _15665_ = ~q[3] /*3620*/;
  assign _15666_ = sum_29[26] & q[3] /*3619*/;
  assign _15667_ = m_29[26] & _15665_ /*3618*/;
  assign r_29[26] = _15667_ | _15666_ /*3617*/;
  assign _15668_ = ~q[3] /*3616*/;
  assign _15669_ = sum_29[27] & q[3] /*3615*/;
  assign _15670_ = m_29[27] & _15668_ /*3614*/;
  assign r_29[27] = _15670_ | _15669_ /*3613*/;
  assign _15671_ = ~q[3] /*3612*/;
  assign _15672_ = sum_29[28] & q[3] /*3611*/;
  assign _15673_ = m_29[28] & _15671_ /*3610*/;
  assign r_29[28] = _15673_ | _15672_ /*3609*/;
  assign _15674_ = ~q[3] /*3608*/;
  assign _15675_ = sum_29[29] & q[3] /*3607*/;
  assign _15676_ = m_29[29] & _15674_ /*3606*/;
  assign r_29[29] = _15676_ | _15675_ /*3605*/;
  assign _15677_ = ~q[3] /*3604*/;
  assign _15678_ = sum_29[30] & q[3] /*3603*/;
  assign _15679_ = m_29[30] & _15677_ /*3602*/;
  assign r_29[30] = _15679_ | _15678_ /*3601*/;
  assign _15680_ = ~q[3] /*3600*/;
  assign _15681_ = sum_29[31] & q[3] /*3599*/;
  assign _15682_ = m_29[31] & _15680_ /*3598*/;
  assign r_29[31] = _15682_ | _15681_ /*3597*/;
  assign _15683_ = ~q[3] /*3596*/;
  assign _15684_ = sum_29[32] & q[3] /*3595*/;
  assign _15685_ = m_29[32] & _15683_ /*3594*/;
  assign r_29[32] = _15685_ | _15684_ /*3593*/;
  assign _15686_ = ~q[3] /*3592*/;
  assign _15687_ = sum_29[33] & q[3] /*3591*/;
  assign _15688_ = m_29[33] & _15686_ /*3590*/;
  assign r_29[33] = _15688_ | _15687_ /*3589*/;
  assign _15689_ = ~q[3] /*3588*/;
  assign _15690_ = sum_29[34] & q[3] /*3587*/;
  assign _15691_ = m_29[34] & _15689_ /*3586*/;
  assign r_29[34] = _15691_ | _15690_ /*3585*/;
  assign _15692_ = ~q[3] /*3584*/;
  assign _15693_ = sum_29[35] & q[3] /*3583*/;
  assign _15694_ = m_29[35] & _15692_ /*3582*/;
  assign r_29[35] = _15694_ | _15693_ /*3581*/;
  assign _15695_ = ~q[3] /*3580*/;
  assign _15696_ = sum_29[36] & q[3] /*3579*/;
  assign _15697_ = m_29[36] & _15695_ /*3578*/;
  assign r_29[36] = _15697_ | _15696_ /*3577*/;
  assign _15698_ = ~q[3] /*3576*/;
  assign _15699_ = sum_29[37] & q[3] /*3575*/;
  assign _15700_ = m_29[37] & _15698_ /*3574*/;
  assign r_29[37] = _15700_ | _15699_ /*3573*/;
  assign _15701_ = ~q[3] /*3572*/;
  assign _15702_ = sum_29[38] & q[3] /*3571*/;
  assign _15703_ = m_29[38] & _15701_ /*3570*/;
  assign r_29[38] = _15703_ | _15702_ /*3569*/;
  assign _15704_ = ~q[3] /*3568*/;
  assign _15705_ = sum_29[39] & q[3] /*3567*/;
  assign _15706_ = m_29[39] & _15704_ /*3566*/;
  assign r_29[39] = _15706_ | _15705_ /*3565*/;
  assign _15707_ = ~q[3] /*3564*/;
  assign _15708_ = sum_29[40] & q[3] /*3563*/;
  assign _15709_ = m_29[40] & _15707_ /*3562*/;
  assign r_29[40] = _15709_ | _15708_ /*3561*/;
  assign _15710_ = ~q[3] /*3560*/;
  assign _15711_ = sum_29[41] & q[3] /*3559*/;
  assign _15712_ = m_29[41] & _15710_ /*3558*/;
  assign r_29[41] = _15712_ | _15711_ /*3557*/;
  assign _15713_ = ~q[3] /*3556*/;
  assign _15714_ = sum_29[42] & q[3] /*3555*/;
  assign _15715_ = m_29[42] & _15713_ /*3554*/;
  assign r_29[42] = _15715_ | _15714_ /*3553*/;
  assign _15716_ = ~q[3] /*3552*/;
  assign _15717_ = sum_29[43] & q[3] /*3551*/;
  assign _15718_ = m_29[43] & _15716_ /*3550*/;
  assign r_29[43] = _15718_ | _15717_ /*3549*/;
  assign _15719_ = ~q[3] /*3548*/;
  assign _15720_ = sum_29[44] & q[3] /*3547*/;
  assign _15721_ = m_29[44] & _15719_ /*3546*/;
  assign r_29[44] = _15721_ | _15720_ /*3545*/;
  assign _15722_ = ~q[3] /*3544*/;
  assign _15723_ = sum_29[45] & q[3] /*3543*/;
  assign _15724_ = m_29[45] & _15722_ /*3542*/;
  assign r_29[45] = _15724_ | _15723_ /*3541*/;
  assign _15725_ = ~q[3] /*3540*/;
  assign _15726_ = sum_29[46] & q[3] /*3539*/;
  assign _15727_ = m_29[46] & _15725_ /*3538*/;
  assign r_29[46] = _15727_ | _15726_ /*3537*/;
  assign _15728_ = ~q[3] /*3536*/;
  assign _15729_ = sum_29[47] & q[3] /*3535*/;
  assign _15730_ = m_29[47] & _15728_ /*3534*/;
  assign r_29[47] = _15730_ | _15729_ /*3533*/;
  assign _15731_ = ~q[3] /*3532*/;
  assign _15732_ = sum_29[48] & q[3] /*3531*/;
  assign _15733_ = m_29[48] & _15731_ /*3530*/;
  assign r_29[48] = _15733_ | _15732_ /*3529*/;
  assign _15734_ = ~q[3] /*3528*/;
  assign _15735_ = sum_29[49] & q[3] /*3527*/;
  assign _15736_ = m_29[49] & _15734_ /*3526*/;
  assign r_29[49] = _15736_ | _15735_ /*3525*/;
  assign _15737_ = ~q[3] /*3524*/;
  assign _15738_ = sum_29[50] & q[3] /*3523*/;
  assign _15739_ = m_29[50] & _15737_ /*3522*/;
  assign r_29[50] = _15739_ | _15738_ /*3521*/;
  assign _15740_ = ~q[3] /*3520*/;
  assign _15741_ = sum_29[51] & q[3] /*3519*/;
  assign _15742_ = m_29[51] & _15740_ /*3518*/;
  assign r_29[51] = _15742_ | _15741_ /*3517*/;
  assign _15743_ = ~q[3] /*3516*/;
  assign _15744_ = sum_29[52] & q[3] /*3515*/;
  assign _15745_ = m_29[52] & _15743_ /*3514*/;
  assign r_29[52] = _15745_ | _15744_ /*3513*/;
  assign _15746_ = ~q[3] /*3512*/;
  assign _15747_ = sum_29[53] & q[3] /*3511*/;
  assign _15748_ = m_29[53] & _15746_ /*3510*/;
  assign r_29[53] = _15748_ | _15747_ /*3509*/;
  assign _15749_ = ~q[3] /*3508*/;
  assign _15750_ = sum_29[54] & q[3] /*3507*/;
  assign _15751_ = m_29[54] & _15749_ /*3506*/;
  assign r_29[54] = _15751_ | _15750_ /*3505*/;
  assign _15752_ = ~q[3] /*3504*/;
  assign _15753_ = sum_29[55] & q[3] /*3503*/;
  assign _15754_ = m_29[55] & _15752_ /*3502*/;
  assign r_29[55] = _15754_ | _15753_ /*3501*/;
  assign _15755_ = ~q[3] /*3500*/;
  assign _15756_ = sum_29[56] & q[3] /*3499*/;
  assign _15757_ = m_29[56] & _15755_ /*3498*/;
  assign r_29[56] = _15757_ | _15756_ /*3497*/;
  assign _15758_ = ~q[3] /*3496*/;
  assign _15759_ = sum_29[57] & q[3] /*3495*/;
  assign _15760_ = m_29[57] & _15758_ /*3494*/;
  assign r_29[57] = _15760_ | _15759_ /*3493*/;
  assign _15761_ = ~q[3] /*3492*/;
  assign _15762_ = sum_29[58] & q[3] /*3491*/;
  assign _15763_ = m_29[58] & _15761_ /*3490*/;
  assign r_29[58] = _15763_ | _15762_ /*3489*/;
  assign _15764_ = ~q[3] /*3488*/;
  assign _15765_ = sum_29[59] & q[3] /*3487*/;
  assign _15766_ = m_29[59] & _15764_ /*3486*/;
  assign r_29[59] = _15766_ | _15765_ /*3485*/;
  assign _15767_ = ~q[3] /*3484*/;
  assign _15768_ = sum_29[60] & q[3] /*3483*/;
  assign _15769_ = m_29[60] & _15767_ /*3482*/;
  assign r_29[60] = _15769_ | _15768_ /*3481*/;
  assign _15770_ = ~q[3] /*3480*/;
  assign _15771_ = sum_29[61] & q[3] /*3479*/;
  assign _15772_ = m_29[61] & _15770_ /*3478*/;
  assign r_29[61] = _15772_ | _15771_ /*3477*/;
  assign _15773_ = ~q[3] /*3476*/;
  assign _15774_ = sum_29[62] & q[3] /*3475*/;
  assign _15775_ = m_29[62] & _15773_ /*3474*/;
  assign r_29[62] = _15775_ | _15774_ /*3473*/;
  assign _15776_ = ~q[3] /*3472*/;
  assign _15777_ = sum_29[63] & q[3] /*3471*/;
  assign _15778_ = m_29[63] & _15776_ /*3470*/;
  assign r_29[63] = _15778_ | _15777_ /*3469*/;
  assign _15779_ = ~q[3] /*3468*/;
  assign _15780_ = sum_29[64] & q[3] /*3467*/;
  assign _15781_ = m_29[64] & _15779_ /*3466*/;
  assign r_29[64] = _15781_ | _15780_ /*3465*/;
  assign _15782_ = ~q[3] /*3464*/;
  assign _15783_ = sum_29[65] & q[3] /*3463*/;
  assign _15784_ = m_29[65] & _15782_ /*3462*/;
  assign r_29[65] = _15784_ | _15783_ /*3461*/;
  assign _15785_ = ~q[3] /*3460*/;
  assign _15786_ = sum_29[66] & q[3] /*3459*/;
  assign _15787_ = m_29[66] & _15785_ /*3458*/;
  assign r_29[66] = _15787_ | _15786_ /*3457*/;
  assign _15788_ = ~q[3] /*3456*/;
  assign _15789_ = sum_29[67] & q[3] /*3455*/;
  assign _15790_ = m_29[67] & _15788_ /*3454*/;
  assign r_29[67] = _15790_ | _15789_ /*3453*/;
  assign _15791_ = ~q[3] /*3452*/;
  assign _15792_ = sum_29[68] & q[3] /*3451*/;
  assign _15793_ = m_29[68] & _15791_ /*3450*/;
  assign r_29[68] = _15793_ | _15792_ /*3449*/;
  assign _15794_ = ~q[3] /*3448*/;
  assign _15795_ = sum_29[69] & q[3] /*3447*/;
  assign _15796_ = m_29[69] & _15794_ /*3446*/;
  assign r_29[69] = _15796_ | _15795_ /*3445*/;
  assign _15797_ = ~q[3] /*3444*/;
  assign _15798_ = sum_29[70] & q[3] /*3443*/;
  assign _15799_ = m_29[70] & _15797_ /*3442*/;
  assign r_29[70] = _15799_ | _15798_ /*3441*/;
  assign _15800_ = ~q[3] /*3440*/;
  assign _15801_ = sum_29[71] & q[3] /*3439*/;
  assign _15802_ = m_29[71] & _15800_ /*3438*/;
  assign r_29[71] = _15802_ | _15801_ /*3437*/;
  assign _15803_ = ~q[3] /*3436*/;
  assign _15804_ = sum_29[72] & q[3] /*3435*/;
  assign _15805_ = m_29[72] & _15803_ /*3434*/;
  assign r_29[72] = _15805_ | _15804_ /*3433*/;
  assign _15806_ = ~q[3] /*3432*/;
  assign _15807_ = sum_29[73] & q[3] /*3431*/;
  assign _15808_ = m_29[73] & _15806_ /*3430*/;
  assign r_29[73] = _15808_ | _15807_ /*3429*/;
  assign _15809_ = ~q[3] /*3428*/;
  assign _15810_ = sum_29[74] & q[3] /*3427*/;
  assign _15811_ = m_29[74] & _15809_ /*3426*/;
  assign r_29[74] = _15811_ | _15810_ /*3425*/;
  assign _15812_ = ~q[3] /*3424*/;
  assign _15813_ = sum_29[75] & q[3] /*3423*/;
  assign _15814_ = m_29[75] & _15812_ /*3422*/;
  assign r_29[75] = _15814_ | _15813_ /*3421*/;
  assign _15815_ = ~q[3] /*3420*/;
  assign _15816_ = sum_29[76] & q[3] /*3419*/;
  assign _15817_ = m_29[76] & _15815_ /*3418*/;
  assign r_29[76] = _15817_ | _15816_ /*3417*/;
  assign _15818_ = ~q[3] /*3416*/;
  assign _15819_ = sum_29[77] & q[3] /*3415*/;
  assign _15820_ = m_29[77] & _15818_ /*3414*/;
  assign r_29[77] = _15820_ | _15819_ /*3413*/;
  assign _15821_ = ~q[3] /*3412*/;
  assign _15822_ = sum_29[78] & q[3] /*3411*/;
  assign _15823_ = m_29[78] & _15821_ /*3410*/;
  assign r_29[78] = _15823_ | _15822_ /*3409*/;
  assign _15824_ = ~q[3] /*3408*/;
  assign _15825_ = sum_29[79] & q[3] /*3407*/;
  assign _15826_ = m_29[79] & _15824_ /*3406*/;
  assign r_29[79] = _15826_ | _15825_ /*3405*/;
  assign _15827_ = ~q[3] /*3404*/;
  assign _15828_ = sum_29[80] & q[3] /*3403*/;
  assign _15829_ = m_29[80] & _15827_ /*3402*/;
  assign r_29[80] = _15829_ | _15828_ /*3401*/;
  assign _15830_ = ~q[3] /*3400*/;
  assign _15831_ = sum_29[81] & q[3] /*3399*/;
  assign _15832_ = m_29[81] & _15830_ /*3398*/;
  assign r_29[81] = _15832_ | _15831_ /*3397*/;
  assign _15833_ = ~q[3] /*3396*/;
  assign _15834_ = sum_29[82] & q[3] /*3395*/;
  assign _15835_ = m_29[82] & _15833_ /*3394*/;
  assign r_29[82] = _15835_ | _15834_ /*3393*/;
  assign _15836_ = ~q[3] /*3392*/;
  assign _15837_ = sum_29[83] & q[3] /*3391*/;
  assign _15838_ = m_29[83] & _15836_ /*3390*/;
  assign r_29[83] = _15838_ | _15837_ /*3389*/;
  assign _15839_ = ~q[3] /*3388*/;
  assign _15840_ = sum_29[84] & q[3] /*3387*/;
  assign _15841_ = m_29[84] & _15839_ /*3386*/;
  assign r_29[84] = _15841_ | _15840_ /*3385*/;
  assign _15842_ = ~q[3] /*3384*/;
  assign _15843_ = sum_29[85] & q[3] /*3383*/;
  assign _15844_ = m_29[85] & _15842_ /*3382*/;
  assign r_29[85] = _15844_ | _15843_ /*3381*/;
  assign _15845_ = ~q[3] /*3380*/;
  assign _15846_ = sum_29[86] & q[3] /*3379*/;
  assign _15847_ = m_29[86] & _15845_ /*3378*/;
  assign r_29[86] = _15847_ | _15846_ /*3377*/;
  assign _15848_ = ~q[3] /*3376*/;
  assign _15849_ = sum_29[87] & q[3] /*3375*/;
  assign _15850_ = m_29[87] & _15848_ /*3374*/;
  assign r_29[87] = _15850_ | _15849_ /*3373*/;
  assign _15851_ = ~q[3] /*3372*/;
  assign _15852_ = sum_29[88] & q[3] /*3371*/;
  assign _15853_ = m_29[88] & _15851_ /*3370*/;
  assign r_29[88] = _15853_ | _15852_ /*3369*/;
  assign _15854_ = ~q[3] /*3368*/;
  assign _15855_ = sum_29[89] & q[3] /*3367*/;
  assign _15856_ = m_29[89] & _15854_ /*3366*/;
  assign r_29[89] = _15856_ | _15855_ /*3365*/;
  assign _15857_ = ~q[3] /*3364*/;
  assign _15858_ = sum_29[90] & q[3] /*3363*/;
  assign _15859_ = m_29[90] & _15857_ /*3362*/;
  assign r_29[90] = _15859_ | _15858_ /*3361*/;
  assign _15860_ = ~q[3] /*3360*/;
  assign _15861_ = sum_29[91] & q[3] /*3359*/;
  assign _15862_ = m_29[91] & _15860_ /*3358*/;
  assign r_29[91] = _15862_ | _15861_ /*3357*/;
  assign inv_30[0] = oneWire /*3292*/;
  assign inv_30[1] = oneWire /*3286*/;
  assign inv_30[2] = ~div[0] /*3280*/;
  assign inv_30[3] = ~div[1] /*3274*/;
  assign inv_30[4] = ~div[2] /*3268*/;
  assign inv_30[5] = ~div[3] /*3262*/;
  assign inv_30[6] = ~div[4] /*3256*/;
  assign inv_30[7] = ~div[5] /*3250*/;
  assign inv_30[8] = ~div[6] /*3244*/;
  assign inv_30[9] = ~div[7] /*3238*/;
  assign inv_30[10] = ~div[8] /*3232*/;
  assign inv_30[11] = ~div[9] /*3226*/;
  assign inv_30[12] = ~div[10] /*3220*/;
  assign inv_30[13] = ~div[11] /*3214*/;
  assign inv_30[14] = ~div[12] /*3208*/;
  assign inv_30[15] = ~div[13] /*3202*/;
  assign inv_30[16] = ~div[14] /*3196*/;
  assign inv_30[17] = ~div[15] /*3190*/;
  assign inv_30[18] = ~div[16] /*3184*/;
  assign inv_30[19] = ~div[17] /*3178*/;
  assign inv_30[20] = ~div[18] /*3172*/;
  assign inv_30[21] = ~div[19] /*3166*/;
  assign inv_30[22] = ~div[20] /*3160*/;
  assign inv_30[23] = ~div[21] /*3154*/;
  assign inv_30[24] = ~div[22] /*3148*/;
  assign inv_30[25] = ~div[23] /*3142*/;
  assign inv_30[26] = ~div[24] /*3136*/;
  assign inv_30[27] = ~div[25] /*3130*/;
  assign inv_30[28] = ~div[26] /*3124*/;
  assign inv_30[29] = ~div[27] /*3118*/;
  assign inv_30[30] = ~div[28] /*3112*/;
  assign inv_30[31] = ~div[29] /*3106*/;
  assign inv_30[32] = ~div[30] /*3100*/;
  assign inv_30[33] = oneWire /*3094*/;
  assign inv_30[34] = oneWire /*3088*/;
  assign inv_30[35] = oneWire /*3082*/;
  assign inv_30[36] = oneWire /*3076*/;
  assign inv_30[37] = oneWire /*3070*/;
  assign inv_30[38] = oneWire /*3064*/;
  assign inv_30[39] = oneWire /*3058*/;
  assign inv_30[40] = oneWire /*3052*/;
  assign inv_30[41] = oneWire /*3046*/;
  assign inv_30[42] = oneWire /*3040*/;
  assign inv_30[43] = oneWire /*3034*/;
  assign inv_30[44] = oneWire /*3028*/;
  assign inv_30[45] = oneWire /*3022*/;
  assign inv_30[46] = oneWire /*3016*/;
  assign inv_30[47] = oneWire /*3010*/;
  assign inv_30[48] = oneWire /*3004*/;
  assign inv_30[49] = oneWire /*2998*/;
  assign inv_30[50] = oneWire /*2992*/;
  assign inv_30[51] = oneWire /*2986*/;
  assign inv_30[52] = oneWire /*2980*/;
  assign inv_30[53] = oneWire /*2974*/;
  assign inv_30[54] = oneWire /*2968*/;
  assign inv_30[55] = oneWire /*2962*/;
  assign inv_30[56] = oneWire /*2956*/;
  assign inv_30[57] = oneWire /*2950*/;
  assign inv_30[58] = oneWire /*2944*/;
  assign inv_30[59] = oneWire /*2938*/;
  assign inv_30[60] = oneWire /*2932*/;
  assign inv_30[61] = oneWire /*2926*/;
  assign inv_30[62] = oneWire /*2920*/;
  assign inv_30[63] = oneWire /*2914*/;
  assign inv_30[64] = oneWire /*2908*/;
  assign inv_30[65] = oneWire /*2902*/;
  assign inv_30[66] = oneWire /*2896*/;
  assign inv_30[67] = oneWire /*2890*/;
  assign inv_30[68] = oneWire /*2884*/;
  assign inv_30[69] = oneWire /*2878*/;
  assign inv_30[70] = oneWire /*2872*/;
  assign inv_30[71] = oneWire /*2866*/;
  assign inv_30[72] = oneWire /*2860*/;
  assign inv_30[73] = oneWire /*2854*/;
  assign inv_30[74] = oneWire /*2848*/;
  assign inv_30[75] = oneWire /*2842*/;
  assign inv_30[76] = oneWire /*2836*/;
  assign inv_30[77] = oneWire /*2830*/;
  assign inv_30[78] = oneWire /*2824*/;
  assign inv_30[79] = oneWire /*2818*/;
  assign inv_30[80] = oneWire /*2812*/;
  assign inv_30[81] = oneWire /*2806*/;
  assign inv_30[82] = oneWire /*2800*/;
  assign inv_30[83] = oneWire /*2794*/;
  assign inv_30[84] = oneWire /*2788*/;
  assign inv_30[85] = oneWire /*2782*/;
  assign inv_30[86] = oneWire /*2776*/;
  assign inv_30[87] = oneWire /*2770*/;
  assign inv_30[88] = oneWire /*2764*/;
  assign inv_30[89] = oneWire /*2758*/;
  assign inv_30[90] = oneWire /*2752*/;
  assign inv_30[91] = oneWire /*2746*/;
  assign _15863_ = inv_30[0] ^ r_29[0] /*3291*/;
  assign sum_30[0] = _15863_ ^ oneWire /*3290*/;
  assign _15864_ = _15863_ & oneWire /*3289*/;
  assign _15865_ = inv_30[0] & r_29[0] /*3288*/;
  assign _15866_ = _15864_ | _15865_ /*3287*/;
  assign _15867_ = inv_30[1] ^ r_29[1] /*3285*/;
  assign sum_30[1] = _15867_ ^ _15866_ /*3284*/;
  assign _15868_ = _15867_ & _15866_ /*3283*/;
  assign _15869_ = inv_30[1] & r_29[1] /*3282*/;
  assign _15870_ = _15868_ | _15869_ /*3281*/;
  assign _15871_ = inv_30[2] ^ r_29[2] /*3279*/;
  assign sum_30[2] = _15871_ ^ _15870_ /*3278*/;
  assign _15872_ = _15871_ & _15870_ /*3277*/;
  assign _15873_ = inv_30[2] & r_29[2] /*3276*/;
  assign _15874_ = _15872_ | _15873_ /*3275*/;
  assign _15875_ = inv_30[3] ^ r_29[3] /*3273*/;
  assign sum_30[3] = _15875_ ^ _15874_ /*3272*/;
  assign _15876_ = _15875_ & _15874_ /*3271*/;
  assign _15877_ = inv_30[3] & r_29[3] /*3270*/;
  assign _15878_ = _15876_ | _15877_ /*3269*/;
  assign _15879_ = inv_30[4] ^ r_29[4] /*3267*/;
  assign sum_30[4] = _15879_ ^ _15878_ /*3266*/;
  assign _15880_ = _15879_ & _15878_ /*3265*/;
  assign _15881_ = inv_30[4] & r_29[4] /*3264*/;
  assign _15882_ = _15880_ | _15881_ /*3263*/;
  assign _15883_ = inv_30[5] ^ r_29[5] /*3261*/;
  assign sum_30[5] = _15883_ ^ _15882_ /*3260*/;
  assign _15884_ = _15883_ & _15882_ /*3259*/;
  assign _15885_ = inv_30[5] & r_29[5] /*3258*/;
  assign _15886_ = _15884_ | _15885_ /*3257*/;
  assign _15887_ = inv_30[6] ^ r_29[6] /*3255*/;
  assign sum_30[6] = _15887_ ^ _15886_ /*3254*/;
  assign _15888_ = _15887_ & _15886_ /*3253*/;
  assign _15889_ = inv_30[6] & r_29[6] /*3252*/;
  assign _15890_ = _15888_ | _15889_ /*3251*/;
  assign _15891_ = inv_30[7] ^ r_29[7] /*3249*/;
  assign sum_30[7] = _15891_ ^ _15890_ /*3248*/;
  assign _15892_ = _15891_ & _15890_ /*3247*/;
  assign _15893_ = inv_30[7] & r_29[7] /*3246*/;
  assign _15894_ = _15892_ | _15893_ /*3245*/;
  assign _15895_ = inv_30[8] ^ r_29[8] /*3243*/;
  assign sum_30[8] = _15895_ ^ _15894_ /*3242*/;
  assign _15896_ = _15895_ & _15894_ /*3241*/;
  assign _15897_ = inv_30[8] & r_29[8] /*3240*/;
  assign _15898_ = _15896_ | _15897_ /*3239*/;
  assign _15899_ = inv_30[9] ^ r_29[9] /*3237*/;
  assign sum_30[9] = _15899_ ^ _15898_ /*3236*/;
  assign _15900_ = _15899_ & _15898_ /*3235*/;
  assign _15901_ = inv_30[9] & r_29[9] /*3234*/;
  assign _15902_ = _15900_ | _15901_ /*3233*/;
  assign _15903_ = inv_30[10] ^ r_29[10] /*3231*/;
  assign sum_30[10] = _15903_ ^ _15902_ /*3230*/;
  assign _15904_ = _15903_ & _15902_ /*3229*/;
  assign _15905_ = inv_30[10] & r_29[10] /*3228*/;
  assign _15906_ = _15904_ | _15905_ /*3227*/;
  assign _15907_ = inv_30[11] ^ r_29[11] /*3225*/;
  assign sum_30[11] = _15907_ ^ _15906_ /*3224*/;
  assign _15908_ = _15907_ & _15906_ /*3223*/;
  assign _15909_ = inv_30[11] & r_29[11] /*3222*/;
  assign _15910_ = _15908_ | _15909_ /*3221*/;
  assign _15911_ = inv_30[12] ^ r_29[12] /*3219*/;
  assign sum_30[12] = _15911_ ^ _15910_ /*3218*/;
  assign _15912_ = _15911_ & _15910_ /*3217*/;
  assign _15913_ = inv_30[12] & r_29[12] /*3216*/;
  assign _15914_ = _15912_ | _15913_ /*3215*/;
  assign _15915_ = inv_30[13] ^ r_29[13] /*3213*/;
  assign sum_30[13] = _15915_ ^ _15914_ /*3212*/;
  assign _15916_ = _15915_ & _15914_ /*3211*/;
  assign _15917_ = inv_30[13] & r_29[13] /*3210*/;
  assign _15918_ = _15916_ | _15917_ /*3209*/;
  assign _15919_ = inv_30[14] ^ r_29[14] /*3207*/;
  assign sum_30[14] = _15919_ ^ _15918_ /*3206*/;
  assign _15920_ = _15919_ & _15918_ /*3205*/;
  assign _15921_ = inv_30[14] & r_29[14] /*3204*/;
  assign _15922_ = _15920_ | _15921_ /*3203*/;
  assign _15923_ = inv_30[15] ^ r_29[15] /*3201*/;
  assign sum_30[15] = _15923_ ^ _15922_ /*3200*/;
  assign _15924_ = _15923_ & _15922_ /*3199*/;
  assign _15925_ = inv_30[15] & r_29[15] /*3198*/;
  assign _15926_ = _15924_ | _15925_ /*3197*/;
  assign _15927_ = inv_30[16] ^ r_29[16] /*3195*/;
  assign sum_30[16] = _15927_ ^ _15926_ /*3194*/;
  assign _15928_ = _15927_ & _15926_ /*3193*/;
  assign _15929_ = inv_30[16] & r_29[16] /*3192*/;
  assign _15930_ = _15928_ | _15929_ /*3191*/;
  assign _15931_ = inv_30[17] ^ r_29[17] /*3189*/;
  assign sum_30[17] = _15931_ ^ _15930_ /*3188*/;
  assign _15932_ = _15931_ & _15930_ /*3187*/;
  assign _15933_ = inv_30[17] & r_29[17] /*3186*/;
  assign _15934_ = _15932_ | _15933_ /*3185*/;
  assign _15935_ = inv_30[18] ^ r_29[18] /*3183*/;
  assign sum_30[18] = _15935_ ^ _15934_ /*3182*/;
  assign _15936_ = _15935_ & _15934_ /*3181*/;
  assign _15937_ = inv_30[18] & r_29[18] /*3180*/;
  assign _15938_ = _15936_ | _15937_ /*3179*/;
  assign _15939_ = inv_30[19] ^ r_29[19] /*3177*/;
  assign sum_30[19] = _15939_ ^ _15938_ /*3176*/;
  assign _15940_ = _15939_ & _15938_ /*3175*/;
  assign _15941_ = inv_30[19] & r_29[19] /*3174*/;
  assign _15942_ = _15940_ | _15941_ /*3173*/;
  assign _15943_ = inv_30[20] ^ r_29[20] /*3171*/;
  assign sum_30[20] = _15943_ ^ _15942_ /*3170*/;
  assign _15944_ = _15943_ & _15942_ /*3169*/;
  assign _15945_ = inv_30[20] & r_29[20] /*3168*/;
  assign _15946_ = _15944_ | _15945_ /*3167*/;
  assign _15947_ = inv_30[21] ^ r_29[21] /*3165*/;
  assign sum_30[21] = _15947_ ^ _15946_ /*3164*/;
  assign _15948_ = _15947_ & _15946_ /*3163*/;
  assign _15949_ = inv_30[21] & r_29[21] /*3162*/;
  assign _15950_ = _15948_ | _15949_ /*3161*/;
  assign _15951_ = inv_30[22] ^ r_29[22] /*3159*/;
  assign sum_30[22] = _15951_ ^ _15950_ /*3158*/;
  assign _15952_ = _15951_ & _15950_ /*3157*/;
  assign _15953_ = inv_30[22] & r_29[22] /*3156*/;
  assign _15954_ = _15952_ | _15953_ /*3155*/;
  assign _15955_ = inv_30[23] ^ r_29[23] /*3153*/;
  assign sum_30[23] = _15955_ ^ _15954_ /*3152*/;
  assign _15956_ = _15955_ & _15954_ /*3151*/;
  assign _15957_ = inv_30[23] & r_29[23] /*3150*/;
  assign _15958_ = _15956_ | _15957_ /*3149*/;
  assign _15959_ = inv_30[24] ^ r_29[24] /*3147*/;
  assign sum_30[24] = _15959_ ^ _15958_ /*3146*/;
  assign _15960_ = _15959_ & _15958_ /*3145*/;
  assign _15961_ = inv_30[24] & r_29[24] /*3144*/;
  assign _15962_ = _15960_ | _15961_ /*3143*/;
  assign _15963_ = inv_30[25] ^ r_29[25] /*3141*/;
  assign sum_30[25] = _15963_ ^ _15962_ /*3140*/;
  assign _15964_ = _15963_ & _15962_ /*3139*/;
  assign _15965_ = inv_30[25] & r_29[25] /*3138*/;
  assign _15966_ = _15964_ | _15965_ /*3137*/;
  assign _15967_ = inv_30[26] ^ r_29[26] /*3135*/;
  assign sum_30[26] = _15967_ ^ _15966_ /*3134*/;
  assign _15968_ = _15967_ & _15966_ /*3133*/;
  assign _15969_ = inv_30[26] & r_29[26] /*3132*/;
  assign _15970_ = _15968_ | _15969_ /*3131*/;
  assign _15971_ = inv_30[27] ^ r_29[27] /*3129*/;
  assign sum_30[27] = _15971_ ^ _15970_ /*3128*/;
  assign _15972_ = _15971_ & _15970_ /*3127*/;
  assign _15973_ = inv_30[27] & r_29[27] /*3126*/;
  assign _15974_ = _15972_ | _15973_ /*3125*/;
  assign _15975_ = inv_30[28] ^ r_29[28] /*3123*/;
  assign sum_30[28] = _15975_ ^ _15974_ /*3122*/;
  assign _15976_ = _15975_ & _15974_ /*3121*/;
  assign _15977_ = inv_30[28] & r_29[28] /*3120*/;
  assign _15978_ = _15976_ | _15977_ /*3119*/;
  assign _15979_ = inv_30[29] ^ r_29[29] /*3117*/;
  assign sum_30[29] = _15979_ ^ _15978_ /*3116*/;
  assign _15980_ = _15979_ & _15978_ /*3115*/;
  assign _15981_ = inv_30[29] & r_29[29] /*3114*/;
  assign _15982_ = _15980_ | _15981_ /*3113*/;
  assign _15983_ = inv_30[30] ^ r_29[30] /*3111*/;
  assign sum_30[30] = _15983_ ^ _15982_ /*3110*/;
  assign _15984_ = _15983_ & _15982_ /*3109*/;
  assign _15985_ = inv_30[30] & r_29[30] /*3108*/;
  assign _15986_ = _15984_ | _15985_ /*3107*/;
  assign _15987_ = inv_30[31] ^ r_29[31] /*3105*/;
  assign sum_30[31] = _15987_ ^ _15986_ /*3104*/;
  assign _15988_ = _15987_ & _15986_ /*3103*/;
  assign _15989_ = inv_30[31] & r_29[31] /*3102*/;
  assign _15990_ = _15988_ | _15989_ /*3101*/;
  assign _15991_ = inv_30[32] ^ r_29[32] /*3099*/;
  assign sum_30[32] = _15991_ ^ _15990_ /*3098*/;
  assign _15992_ = _15991_ & _15990_ /*3097*/;
  assign _15993_ = inv_30[32] & r_29[32] /*3096*/;
  assign _15994_ = _15992_ | _15993_ /*3095*/;
  assign _15995_ = inv_30[33] ^ r_29[33] /*3093*/;
  assign sum_30[33] = _15995_ ^ _15994_ /*3092*/;
  assign _15996_ = _15995_ & _15994_ /*3091*/;
  assign _15997_ = inv_30[33] & r_29[33] /*3090*/;
  assign _15998_ = _15996_ | _15997_ /*3089*/;
  assign _15999_ = inv_30[34] ^ r_29[34] /*3087*/;
  assign sum_30[34] = _15999_ ^ _15998_ /*3086*/;
  assign _16000_ = _15999_ & _15998_ /*3085*/;
  assign _16001_ = inv_30[34] & r_29[34] /*3084*/;
  assign _16002_ = _16000_ | _16001_ /*3083*/;
  assign _16003_ = inv_30[35] ^ r_29[35] /*3081*/;
  assign sum_30[35] = _16003_ ^ _16002_ /*3080*/;
  assign _16004_ = _16003_ & _16002_ /*3079*/;
  assign _16005_ = inv_30[35] & r_29[35] /*3078*/;
  assign _16006_ = _16004_ | _16005_ /*3077*/;
  assign _16007_ = inv_30[36] ^ r_29[36] /*3075*/;
  assign sum_30[36] = _16007_ ^ _16006_ /*3074*/;
  assign _16008_ = _16007_ & _16006_ /*3073*/;
  assign _16009_ = inv_30[36] & r_29[36] /*3072*/;
  assign _16010_ = _16008_ | _16009_ /*3071*/;
  assign _16011_ = inv_30[37] ^ r_29[37] /*3069*/;
  assign sum_30[37] = _16011_ ^ _16010_ /*3068*/;
  assign _16012_ = _16011_ & _16010_ /*3067*/;
  assign _16013_ = inv_30[37] & r_29[37] /*3066*/;
  assign _16014_ = _16012_ | _16013_ /*3065*/;
  assign _16015_ = inv_30[38] ^ r_29[38] /*3063*/;
  assign sum_30[38] = _16015_ ^ _16014_ /*3062*/;
  assign _16016_ = _16015_ & _16014_ /*3061*/;
  assign _16017_ = inv_30[38] & r_29[38] /*3060*/;
  assign _16018_ = _16016_ | _16017_ /*3059*/;
  assign _16019_ = inv_30[39] ^ r_29[39] /*3057*/;
  assign sum_30[39] = _16019_ ^ _16018_ /*3056*/;
  assign _16020_ = _16019_ & _16018_ /*3055*/;
  assign _16021_ = inv_30[39] & r_29[39] /*3054*/;
  assign _16022_ = _16020_ | _16021_ /*3053*/;
  assign _16023_ = inv_30[40] ^ r_29[40] /*3051*/;
  assign sum_30[40] = _16023_ ^ _16022_ /*3050*/;
  assign _16024_ = _16023_ & _16022_ /*3049*/;
  assign _16025_ = inv_30[40] & r_29[40] /*3048*/;
  assign _16026_ = _16024_ | _16025_ /*3047*/;
  assign _16027_ = inv_30[41] ^ r_29[41] /*3045*/;
  assign sum_30[41] = _16027_ ^ _16026_ /*3044*/;
  assign _16028_ = _16027_ & _16026_ /*3043*/;
  assign _16029_ = inv_30[41] & r_29[41] /*3042*/;
  assign _16030_ = _16028_ | _16029_ /*3041*/;
  assign _16031_ = inv_30[42] ^ r_29[42] /*3039*/;
  assign sum_30[42] = _16031_ ^ _16030_ /*3038*/;
  assign _16032_ = _16031_ & _16030_ /*3037*/;
  assign _16033_ = inv_30[42] & r_29[42] /*3036*/;
  assign _16034_ = _16032_ | _16033_ /*3035*/;
  assign _16035_ = inv_30[43] ^ r_29[43] /*3033*/;
  assign sum_30[43] = _16035_ ^ _16034_ /*3032*/;
  assign _16036_ = _16035_ & _16034_ /*3031*/;
  assign _16037_ = inv_30[43] & r_29[43] /*3030*/;
  assign _16038_ = _16036_ | _16037_ /*3029*/;
  assign _16039_ = inv_30[44] ^ r_29[44] /*3027*/;
  assign sum_30[44] = _16039_ ^ _16038_ /*3026*/;
  assign _16040_ = _16039_ & _16038_ /*3025*/;
  assign _16041_ = inv_30[44] & r_29[44] /*3024*/;
  assign _16042_ = _16040_ | _16041_ /*3023*/;
  assign _16043_ = inv_30[45] ^ r_29[45] /*3021*/;
  assign sum_30[45] = _16043_ ^ _16042_ /*3020*/;
  assign _16044_ = _16043_ & _16042_ /*3019*/;
  assign _16045_ = inv_30[45] & r_29[45] /*3018*/;
  assign _16046_ = _16044_ | _16045_ /*3017*/;
  assign _16047_ = inv_30[46] ^ r_29[46] /*3015*/;
  assign sum_30[46] = _16047_ ^ _16046_ /*3014*/;
  assign _16048_ = _16047_ & _16046_ /*3013*/;
  assign _16049_ = inv_30[46] & r_29[46] /*3012*/;
  assign _16050_ = _16048_ | _16049_ /*3011*/;
  assign _16051_ = inv_30[47] ^ r_29[47] /*3009*/;
  assign sum_30[47] = _16051_ ^ _16050_ /*3008*/;
  assign _16052_ = _16051_ & _16050_ /*3007*/;
  assign _16053_ = inv_30[47] & r_29[47] /*3006*/;
  assign _16054_ = _16052_ | _16053_ /*3005*/;
  assign _16055_ = inv_30[48] ^ r_29[48] /*3003*/;
  assign sum_30[48] = _16055_ ^ _16054_ /*3002*/;
  assign _16056_ = _16055_ & _16054_ /*3001*/;
  assign _16057_ = inv_30[48] & r_29[48] /*3000*/;
  assign _16058_ = _16056_ | _16057_ /*2999*/;
  assign _16059_ = inv_30[49] ^ r_29[49] /*2997*/;
  assign sum_30[49] = _16059_ ^ _16058_ /*2996*/;
  assign _16060_ = _16059_ & _16058_ /*2995*/;
  assign _16061_ = inv_30[49] & r_29[49] /*2994*/;
  assign _16062_ = _16060_ | _16061_ /*2993*/;
  assign _16063_ = inv_30[50] ^ r_29[50] /*2991*/;
  assign sum_30[50] = _16063_ ^ _16062_ /*2990*/;
  assign _16064_ = _16063_ & _16062_ /*2989*/;
  assign _16065_ = inv_30[50] & r_29[50] /*2988*/;
  assign _16066_ = _16064_ | _16065_ /*2987*/;
  assign _16067_ = inv_30[51] ^ r_29[51] /*2985*/;
  assign sum_30[51] = _16067_ ^ _16066_ /*2984*/;
  assign _16068_ = _16067_ & _16066_ /*2983*/;
  assign _16069_ = inv_30[51] & r_29[51] /*2982*/;
  assign _16070_ = _16068_ | _16069_ /*2981*/;
  assign _16071_ = inv_30[52] ^ r_29[52] /*2979*/;
  assign sum_30[52] = _16071_ ^ _16070_ /*2978*/;
  assign _16072_ = _16071_ & _16070_ /*2977*/;
  assign _16073_ = inv_30[52] & r_29[52] /*2976*/;
  assign _16074_ = _16072_ | _16073_ /*2975*/;
  assign _16075_ = inv_30[53] ^ r_29[53] /*2973*/;
  assign sum_30[53] = _16075_ ^ _16074_ /*2972*/;
  assign _16076_ = _16075_ & _16074_ /*2971*/;
  assign _16077_ = inv_30[53] & r_29[53] /*2970*/;
  assign _16078_ = _16076_ | _16077_ /*2969*/;
  assign _16079_ = inv_30[54] ^ r_29[54] /*2967*/;
  assign sum_30[54] = _16079_ ^ _16078_ /*2966*/;
  assign _16080_ = _16079_ & _16078_ /*2965*/;
  assign _16081_ = inv_30[54] & r_29[54] /*2964*/;
  assign _16082_ = _16080_ | _16081_ /*2963*/;
  assign _16083_ = inv_30[55] ^ r_29[55] /*2961*/;
  assign sum_30[55] = _16083_ ^ _16082_ /*2960*/;
  assign _16084_ = _16083_ & _16082_ /*2959*/;
  assign _16085_ = inv_30[55] & r_29[55] /*2958*/;
  assign _16086_ = _16084_ | _16085_ /*2957*/;
  assign _16087_ = inv_30[56] ^ r_29[56] /*2955*/;
  assign sum_30[56] = _16087_ ^ _16086_ /*2954*/;
  assign _16088_ = _16087_ & _16086_ /*2953*/;
  assign _16089_ = inv_30[56] & r_29[56] /*2952*/;
  assign _16090_ = _16088_ | _16089_ /*2951*/;
  assign _16091_ = inv_30[57] ^ r_29[57] /*2949*/;
  assign sum_30[57] = _16091_ ^ _16090_ /*2948*/;
  assign _16092_ = _16091_ & _16090_ /*2947*/;
  assign _16093_ = inv_30[57] & r_29[57] /*2946*/;
  assign _16094_ = _16092_ | _16093_ /*2945*/;
  assign _16095_ = inv_30[58] ^ r_29[58] /*2943*/;
  assign sum_30[58] = _16095_ ^ _16094_ /*2942*/;
  assign _16096_ = _16095_ & _16094_ /*2941*/;
  assign _16097_ = inv_30[58] & r_29[58] /*2940*/;
  assign _16098_ = _16096_ | _16097_ /*2939*/;
  assign _16099_ = inv_30[59] ^ r_29[59] /*2937*/;
  assign sum_30[59] = _16099_ ^ _16098_ /*2936*/;
  assign _16100_ = _16099_ & _16098_ /*2935*/;
  assign _16101_ = inv_30[59] & r_29[59] /*2934*/;
  assign _16102_ = _16100_ | _16101_ /*2933*/;
  assign _16103_ = inv_30[60] ^ r_29[60] /*2931*/;
  assign sum_30[60] = _16103_ ^ _16102_ /*2930*/;
  assign _16104_ = _16103_ & _16102_ /*2929*/;
  assign _16105_ = inv_30[60] & r_29[60] /*2928*/;
  assign _16106_ = _16104_ | _16105_ /*2927*/;
  assign _16107_ = inv_30[61] ^ r_29[61] /*2925*/;
  assign sum_30[61] = _16107_ ^ _16106_ /*2924*/;
  assign _16108_ = _16107_ & _16106_ /*2923*/;
  assign _16109_ = inv_30[61] & r_29[61] /*2922*/;
  assign _16110_ = _16108_ | _16109_ /*2921*/;
  assign _16111_ = inv_30[62] ^ r_29[62] /*2919*/;
  assign sum_30[62] = _16111_ ^ _16110_ /*2918*/;
  assign _16112_ = _16111_ & _16110_ /*2917*/;
  assign _16113_ = inv_30[62] & r_29[62] /*2916*/;
  assign _16114_ = _16112_ | _16113_ /*2915*/;
  assign _16115_ = inv_30[63] ^ r_29[63] /*2913*/;
  assign sum_30[63] = _16115_ ^ _16114_ /*2912*/;
  assign _16116_ = _16115_ & _16114_ /*2911*/;
  assign _16117_ = inv_30[63] & r_29[63] /*2910*/;
  assign _16118_ = _16116_ | _16117_ /*2909*/;
  assign _16119_ = inv_30[64] ^ r_29[64] /*2907*/;
  assign sum_30[64] = _16119_ ^ _16118_ /*2906*/;
  assign _16120_ = _16119_ & _16118_ /*2905*/;
  assign _16121_ = inv_30[64] & r_29[64] /*2904*/;
  assign _16122_ = _16120_ | _16121_ /*2903*/;
  assign _16123_ = inv_30[65] ^ r_29[65] /*2901*/;
  assign sum_30[65] = _16123_ ^ _16122_ /*2900*/;
  assign _16124_ = _16123_ & _16122_ /*2899*/;
  assign _16125_ = inv_30[65] & r_29[65] /*2898*/;
  assign _16126_ = _16124_ | _16125_ /*2897*/;
  assign _16127_ = inv_30[66] ^ r_29[66] /*2895*/;
  assign sum_30[66] = _16127_ ^ _16126_ /*2894*/;
  assign _16128_ = _16127_ & _16126_ /*2893*/;
  assign _16129_ = inv_30[66] & r_29[66] /*2892*/;
  assign _16130_ = _16128_ | _16129_ /*2891*/;
  assign _16131_ = inv_30[67] ^ r_29[67] /*2889*/;
  assign sum_30[67] = _16131_ ^ _16130_ /*2888*/;
  assign _16132_ = _16131_ & _16130_ /*2887*/;
  assign _16133_ = inv_30[67] & r_29[67] /*2886*/;
  assign _16134_ = _16132_ | _16133_ /*2885*/;
  assign _16135_ = inv_30[68] ^ r_29[68] /*2883*/;
  assign sum_30[68] = _16135_ ^ _16134_ /*2882*/;
  assign _16136_ = _16135_ & _16134_ /*2881*/;
  assign _16137_ = inv_30[68] & r_29[68] /*2880*/;
  assign _16138_ = _16136_ | _16137_ /*2879*/;
  assign _16139_ = inv_30[69] ^ r_29[69] /*2877*/;
  assign sum_30[69] = _16139_ ^ _16138_ /*2876*/;
  assign _16140_ = _16139_ & _16138_ /*2875*/;
  assign _16141_ = inv_30[69] & r_29[69] /*2874*/;
  assign _16142_ = _16140_ | _16141_ /*2873*/;
  assign _16143_ = inv_30[70] ^ r_29[70] /*2871*/;
  assign sum_30[70] = _16143_ ^ _16142_ /*2870*/;
  assign _16144_ = _16143_ & _16142_ /*2869*/;
  assign _16145_ = inv_30[70] & r_29[70] /*2868*/;
  assign _16146_ = _16144_ | _16145_ /*2867*/;
  assign _16147_ = inv_30[71] ^ r_29[71] /*2865*/;
  assign sum_30[71] = _16147_ ^ _16146_ /*2864*/;
  assign _16148_ = _16147_ & _16146_ /*2863*/;
  assign _16149_ = inv_30[71] & r_29[71] /*2862*/;
  assign _16150_ = _16148_ | _16149_ /*2861*/;
  assign _16151_ = inv_30[72] ^ r_29[72] /*2859*/;
  assign sum_30[72] = _16151_ ^ _16150_ /*2858*/;
  assign _16152_ = _16151_ & _16150_ /*2857*/;
  assign _16153_ = inv_30[72] & r_29[72] /*2856*/;
  assign _16154_ = _16152_ | _16153_ /*2855*/;
  assign _16155_ = inv_30[73] ^ r_29[73] /*2853*/;
  assign sum_30[73] = _16155_ ^ _16154_ /*2852*/;
  assign _16156_ = _16155_ & _16154_ /*2851*/;
  assign _16157_ = inv_30[73] & r_29[73] /*2850*/;
  assign _16158_ = _16156_ | _16157_ /*2849*/;
  assign _16159_ = inv_30[74] ^ r_29[74] /*2847*/;
  assign sum_30[74] = _16159_ ^ _16158_ /*2846*/;
  assign _16160_ = _16159_ & _16158_ /*2845*/;
  assign _16161_ = inv_30[74] & r_29[74] /*2844*/;
  assign _16162_ = _16160_ | _16161_ /*2843*/;
  assign _16163_ = inv_30[75] ^ r_29[75] /*2841*/;
  assign sum_30[75] = _16163_ ^ _16162_ /*2840*/;
  assign _16164_ = _16163_ & _16162_ /*2839*/;
  assign _16165_ = inv_30[75] & r_29[75] /*2838*/;
  assign _16166_ = _16164_ | _16165_ /*2837*/;
  assign _16167_ = inv_30[76] ^ r_29[76] /*2835*/;
  assign sum_30[76] = _16167_ ^ _16166_ /*2834*/;
  assign _16168_ = _16167_ & _16166_ /*2833*/;
  assign _16169_ = inv_30[76] & r_29[76] /*2832*/;
  assign _16170_ = _16168_ | _16169_ /*2831*/;
  assign _16171_ = inv_30[77] ^ r_29[77] /*2829*/;
  assign sum_30[77] = _16171_ ^ _16170_ /*2828*/;
  assign _16172_ = _16171_ & _16170_ /*2827*/;
  assign _16173_ = inv_30[77] & r_29[77] /*2826*/;
  assign _16174_ = _16172_ | _16173_ /*2825*/;
  assign _16175_ = inv_30[78] ^ r_29[78] /*2823*/;
  assign sum_30[78] = _16175_ ^ _16174_ /*2822*/;
  assign _16176_ = _16175_ & _16174_ /*2821*/;
  assign _16177_ = inv_30[78] & r_29[78] /*2820*/;
  assign _16178_ = _16176_ | _16177_ /*2819*/;
  assign _16179_ = inv_30[79] ^ r_29[79] /*2817*/;
  assign sum_30[79] = _16179_ ^ _16178_ /*2816*/;
  assign _16180_ = _16179_ & _16178_ /*2815*/;
  assign _16181_ = inv_30[79] & r_29[79] /*2814*/;
  assign _16182_ = _16180_ | _16181_ /*2813*/;
  assign _16183_ = inv_30[80] ^ r_29[80] /*2811*/;
  assign sum_30[80] = _16183_ ^ _16182_ /*2810*/;
  assign _16184_ = _16183_ & _16182_ /*2809*/;
  assign _16185_ = inv_30[80] & r_29[80] /*2808*/;
  assign _16186_ = _16184_ | _16185_ /*2807*/;
  assign _16187_ = inv_30[81] ^ r_29[81] /*2805*/;
  assign sum_30[81] = _16187_ ^ _16186_ /*2804*/;
  assign _16188_ = _16187_ & _16186_ /*2803*/;
  assign _16189_ = inv_30[81] & r_29[81] /*2802*/;
  assign _16190_ = _16188_ | _16189_ /*2801*/;
  assign _16191_ = inv_30[82] ^ r_29[82] /*2799*/;
  assign sum_30[82] = _16191_ ^ _16190_ /*2798*/;
  assign _16192_ = _16191_ & _16190_ /*2797*/;
  assign _16193_ = inv_30[82] & r_29[82] /*2796*/;
  assign _16194_ = _16192_ | _16193_ /*2795*/;
  assign _16195_ = inv_30[83] ^ r_29[83] /*2793*/;
  assign sum_30[83] = _16195_ ^ _16194_ /*2792*/;
  assign _16196_ = _16195_ & _16194_ /*2791*/;
  assign _16197_ = inv_30[83] & r_29[83] /*2790*/;
  assign _16198_ = _16196_ | _16197_ /*2789*/;
  assign _16199_ = inv_30[84] ^ r_29[84] /*2787*/;
  assign sum_30[84] = _16199_ ^ _16198_ /*2786*/;
  assign _16200_ = _16199_ & _16198_ /*2785*/;
  assign _16201_ = inv_30[84] & r_29[84] /*2784*/;
  assign _16202_ = _16200_ | _16201_ /*2783*/;
  assign _16203_ = inv_30[85] ^ r_29[85] /*2781*/;
  assign sum_30[85] = _16203_ ^ _16202_ /*2780*/;
  assign _16204_ = _16203_ & _16202_ /*2779*/;
  assign _16205_ = inv_30[85] & r_29[85] /*2778*/;
  assign _16206_ = _16204_ | _16205_ /*2777*/;
  assign _16207_ = inv_30[86] ^ r_29[86] /*2775*/;
  assign sum_30[86] = _16207_ ^ _16206_ /*2774*/;
  assign _16208_ = _16207_ & _16206_ /*2773*/;
  assign _16209_ = inv_30[86] & r_29[86] /*2772*/;
  assign _16210_ = _16208_ | _16209_ /*2771*/;
  assign _16211_ = inv_30[87] ^ r_29[87] /*2769*/;
  assign sum_30[87] = _16211_ ^ _16210_ /*2768*/;
  assign _16212_ = _16211_ & _16210_ /*2767*/;
  assign _16213_ = inv_30[87] & r_29[87] /*2766*/;
  assign _16214_ = _16212_ | _16213_ /*2765*/;
  assign _16215_ = inv_30[88] ^ r_29[88] /*2763*/;
  assign sum_30[88] = _16215_ ^ _16214_ /*2762*/;
  assign _16216_ = _16215_ & _16214_ /*2761*/;
  assign _16217_ = inv_30[88] & r_29[88] /*2760*/;
  assign _16218_ = _16216_ | _16217_ /*2759*/;
  assign _16219_ = inv_30[89] ^ r_29[89] /*2757*/;
  assign sum_30[89] = _16219_ ^ _16218_ /*2756*/;
  assign _16220_ = _16219_ & _16218_ /*2755*/;
  assign _16221_ = inv_30[89] & r_29[89] /*2754*/;
  assign _16222_ = _16220_ | _16221_ /*2753*/;
  assign _16223_ = inv_30[90] ^ r_29[90] /*2751*/;
  assign sum_30[90] = _16223_ ^ _16222_ /*2750*/;
  assign _16224_ = _16223_ & _16222_ /*2749*/;
  assign _16225_ = inv_30[90] & r_29[90] /*2748*/;
  assign _16226_ = _16224_ | _16225_ /*2747*/;
  assign _16227_ = inv_30[91] ^ r_29[91] /*2745*/;
  assign sum_30[91] = _16227_ ^ _16226_ /*2744*/;
  assign _16228_ = _16227_ & _16226_ /*2743*/;
  assign _16229_ = inv_30[91] & r_29[91] /*2742*/;
  assign _16230_ = _16228_ | _16229_ /*2741*/;
  assign _16231_ = _16230_ ^ _16226_ /*2740*/;
  assign _16232_ = ~_16231_ /*2739*/;
  assign _16233_ = sum_30[91] & _16232_ /*2738*/;
  assign _16234_ = _16231_ & _16230_ /*2737*/;
  assign sum_30[92] = _16234_ | _16233_ /*2736*/;
  assign q[2] = ~sum_30[92] /*2735*/;
  assign m_30[0] = r_29[0] /*2734*/;
  assign m_30[1] = r_29[1] /*2733*/;
  assign m_30[2] = r_29[2] /*2732*/;
  assign m_30[3] = r_29[3] /*2731*/;
  assign m_30[4] = r_29[4] /*2730*/;
  assign m_30[5] = r_29[5] /*2729*/;
  assign m_30[6] = r_29[6] /*2728*/;
  assign m_30[7] = r_29[7] /*2727*/;
  assign m_30[8] = r_29[8] /*2726*/;
  assign m_30[9] = r_29[9] /*2725*/;
  assign m_30[10] = r_29[10] /*2724*/;
  assign m_30[11] = r_29[11] /*2723*/;
  assign m_30[12] = r_29[12] /*2722*/;
  assign m_30[13] = r_29[13] /*2721*/;
  assign m_30[14] = r_29[14] /*2720*/;
  assign m_30[15] = r_29[15] /*2719*/;
  assign m_30[16] = r_29[16] /*2718*/;
  assign m_30[17] = r_29[17] /*2717*/;
  assign m_30[18] = r_29[18] /*2716*/;
  assign m_30[19] = r_29[19] /*2715*/;
  assign m_30[20] = r_29[20] /*2714*/;
  assign m_30[21] = r_29[21] /*2713*/;
  assign m_30[22] = r_29[22] /*2712*/;
  assign m_30[23] = r_29[23] /*2711*/;
  assign m_30[24] = r_29[24] /*2710*/;
  assign m_30[25] = r_29[25] /*2709*/;
  assign m_30[26] = r_29[26] /*2708*/;
  assign m_30[27] = r_29[27] /*2707*/;
  assign m_30[28] = r_29[28] /*2706*/;
  assign m_30[29] = r_29[29] /*2705*/;
  assign m_30[30] = r_29[30] /*2704*/;
  assign m_30[31] = r_29[31] /*2703*/;
  assign m_30[32] = r_29[32] /*2702*/;
  assign m_30[33] = r_29[33] /*2701*/;
  assign m_30[34] = r_29[34] /*2700*/;
  assign m_30[35] = r_29[35] /*2699*/;
  assign m_30[36] = r_29[36] /*2698*/;
  assign m_30[37] = r_29[37] /*2697*/;
  assign m_30[38] = r_29[38] /*2696*/;
  assign m_30[39] = r_29[39] /*2695*/;
  assign m_30[40] = r_29[40] /*2694*/;
  assign m_30[41] = r_29[41] /*2693*/;
  assign m_30[42] = r_29[42] /*2692*/;
  assign m_30[43] = r_29[43] /*2691*/;
  assign m_30[44] = r_29[44] /*2690*/;
  assign m_30[45] = r_29[45] /*2689*/;
  assign m_30[46] = r_29[46] /*2688*/;
  assign m_30[47] = r_29[47] /*2687*/;
  assign m_30[48] = r_29[48] /*2686*/;
  assign m_30[49] = r_29[49] /*2685*/;
  assign m_30[50] = r_29[50] /*2684*/;
  assign m_30[51] = r_29[51] /*2683*/;
  assign m_30[52] = r_29[52] /*2682*/;
  assign m_30[53] = r_29[53] /*2681*/;
  assign m_30[54] = r_29[54] /*2680*/;
  assign m_30[55] = r_29[55] /*2679*/;
  assign m_30[56] = r_29[56] /*2678*/;
  assign m_30[57] = r_29[57] /*2677*/;
  assign m_30[58] = r_29[58] /*2676*/;
  assign m_30[59] = r_29[59] /*2675*/;
  assign m_30[60] = r_29[60] /*2674*/;
  assign m_30[61] = r_29[61] /*2673*/;
  assign m_30[62] = r_29[62] /*2672*/;
  assign m_30[63] = r_29[63] /*2671*/;
  assign m_30[64] = r_29[64] /*2670*/;
  assign m_30[65] = r_29[65] /*2669*/;
  assign m_30[66] = r_29[66] /*2668*/;
  assign m_30[67] = r_29[67] /*2667*/;
  assign m_30[68] = r_29[68] /*2666*/;
  assign m_30[69] = r_29[69] /*2665*/;
  assign m_30[70] = r_29[70] /*2664*/;
  assign m_30[71] = r_29[71] /*2663*/;
  assign m_30[72] = r_29[72] /*2662*/;
  assign m_30[73] = r_29[73] /*2661*/;
  assign m_30[74] = r_29[74] /*2660*/;
  assign m_30[75] = r_29[75] /*2659*/;
  assign m_30[76] = r_29[76] /*2658*/;
  assign m_30[77] = r_29[77] /*2657*/;
  assign m_30[78] = r_29[78] /*2656*/;
  assign m_30[79] = r_29[79] /*2655*/;
  assign m_30[80] = r_29[80] /*2654*/;
  assign m_30[81] = r_29[81] /*2653*/;
  assign m_30[82] = r_29[82] /*2652*/;
  assign m_30[83] = r_29[83] /*2651*/;
  assign m_30[84] = r_29[84] /*2650*/;
  assign m_30[85] = r_29[85] /*2649*/;
  assign m_30[86] = r_29[86] /*2648*/;
  assign m_30[87] = r_29[87] /*2647*/;
  assign m_30[88] = r_29[88] /*2646*/;
  assign m_30[89] = r_29[89] /*2645*/;
  assign m_30[90] = r_29[90] /*2644*/;
  assign m_30[91] = r_29[91] /*2643*/;
  assign m_30[92] = r_29[91] /*2642*/;
  assign _16236_ = ~q[2] /*2641*/;
  assign _16237_ = sum_30[0] & q[2] /*2640*/;
  assign _16238_ = m_30[0] & _16236_ /*2639*/;
  assign r_30[0] = _16238_ | _16237_ /*2638*/;
  assign _16239_ = ~q[2] /*2637*/;
  assign _16240_ = sum_30[1] & q[2] /*2636*/;
  assign _16241_ = m_30[1] & _16239_ /*2635*/;
  assign r_30[1] = _16241_ | _16240_ /*2634*/;
  assign _16242_ = ~q[2] /*2633*/;
  assign _16243_ = sum_30[2] & q[2] /*2632*/;
  assign _16244_ = m_30[2] & _16242_ /*2631*/;
  assign r_30[2] = _16244_ | _16243_ /*2630*/;
  assign _16245_ = ~q[2] /*2629*/;
  assign _16246_ = sum_30[3] & q[2] /*2628*/;
  assign _16247_ = m_30[3] & _16245_ /*2627*/;
  assign r_30[3] = _16247_ | _16246_ /*2626*/;
  assign _16248_ = ~q[2] /*2625*/;
  assign _16249_ = sum_30[4] & q[2] /*2624*/;
  assign _16250_ = m_30[4] & _16248_ /*2623*/;
  assign r_30[4] = _16250_ | _16249_ /*2622*/;
  assign _16251_ = ~q[2] /*2621*/;
  assign _16252_ = sum_30[5] & q[2] /*2620*/;
  assign _16253_ = m_30[5] & _16251_ /*2619*/;
  assign r_30[5] = _16253_ | _16252_ /*2618*/;
  assign _16254_ = ~q[2] /*2617*/;
  assign _16255_ = sum_30[6] & q[2] /*2616*/;
  assign _16256_ = m_30[6] & _16254_ /*2615*/;
  assign r_30[6] = _16256_ | _16255_ /*2614*/;
  assign _16257_ = ~q[2] /*2613*/;
  assign _16258_ = sum_30[7] & q[2] /*2612*/;
  assign _16259_ = m_30[7] & _16257_ /*2611*/;
  assign r_30[7] = _16259_ | _16258_ /*2610*/;
  assign _16260_ = ~q[2] /*2609*/;
  assign _16261_ = sum_30[8] & q[2] /*2608*/;
  assign _16262_ = m_30[8] & _16260_ /*2607*/;
  assign r_30[8] = _16262_ | _16261_ /*2606*/;
  assign _16263_ = ~q[2] /*2605*/;
  assign _16264_ = sum_30[9] & q[2] /*2604*/;
  assign _16265_ = m_30[9] & _16263_ /*2603*/;
  assign r_30[9] = _16265_ | _16264_ /*2602*/;
  assign _16266_ = ~q[2] /*2601*/;
  assign _16267_ = sum_30[10] & q[2] /*2600*/;
  assign _16268_ = m_30[10] & _16266_ /*2599*/;
  assign r_30[10] = _16268_ | _16267_ /*2598*/;
  assign _16269_ = ~q[2] /*2597*/;
  assign _16270_ = sum_30[11] & q[2] /*2596*/;
  assign _16271_ = m_30[11] & _16269_ /*2595*/;
  assign r_30[11] = _16271_ | _16270_ /*2594*/;
  assign _16272_ = ~q[2] /*2593*/;
  assign _16273_ = sum_30[12] & q[2] /*2592*/;
  assign _16274_ = m_30[12] & _16272_ /*2591*/;
  assign r_30[12] = _16274_ | _16273_ /*2590*/;
  assign _16275_ = ~q[2] /*2589*/;
  assign _16276_ = sum_30[13] & q[2] /*2588*/;
  assign _16277_ = m_30[13] & _16275_ /*2587*/;
  assign r_30[13] = _16277_ | _16276_ /*2586*/;
  assign _16278_ = ~q[2] /*2585*/;
  assign _16279_ = sum_30[14] & q[2] /*2584*/;
  assign _16280_ = m_30[14] & _16278_ /*2583*/;
  assign r_30[14] = _16280_ | _16279_ /*2582*/;
  assign _16281_ = ~q[2] /*2581*/;
  assign _16282_ = sum_30[15] & q[2] /*2580*/;
  assign _16283_ = m_30[15] & _16281_ /*2579*/;
  assign r_30[15] = _16283_ | _16282_ /*2578*/;
  assign _16284_ = ~q[2] /*2577*/;
  assign _16285_ = sum_30[16] & q[2] /*2576*/;
  assign _16286_ = m_30[16] & _16284_ /*2575*/;
  assign r_30[16] = _16286_ | _16285_ /*2574*/;
  assign _16287_ = ~q[2] /*2573*/;
  assign _16288_ = sum_30[17] & q[2] /*2572*/;
  assign _16289_ = m_30[17] & _16287_ /*2571*/;
  assign r_30[17] = _16289_ | _16288_ /*2570*/;
  assign _16290_ = ~q[2] /*2569*/;
  assign _16291_ = sum_30[18] & q[2] /*2568*/;
  assign _16292_ = m_30[18] & _16290_ /*2567*/;
  assign r_30[18] = _16292_ | _16291_ /*2566*/;
  assign _16293_ = ~q[2] /*2565*/;
  assign _16294_ = sum_30[19] & q[2] /*2564*/;
  assign _16295_ = m_30[19] & _16293_ /*2563*/;
  assign r_30[19] = _16295_ | _16294_ /*2562*/;
  assign _16296_ = ~q[2] /*2561*/;
  assign _16297_ = sum_30[20] & q[2] /*2560*/;
  assign _16298_ = m_30[20] & _16296_ /*2559*/;
  assign r_30[20] = _16298_ | _16297_ /*2558*/;
  assign _16299_ = ~q[2] /*2557*/;
  assign _16300_ = sum_30[21] & q[2] /*2556*/;
  assign _16301_ = m_30[21] & _16299_ /*2555*/;
  assign r_30[21] = _16301_ | _16300_ /*2554*/;
  assign _16302_ = ~q[2] /*2553*/;
  assign _16303_ = sum_30[22] & q[2] /*2552*/;
  assign _16304_ = m_30[22] & _16302_ /*2551*/;
  assign r_30[22] = _16304_ | _16303_ /*2550*/;
  assign _16305_ = ~q[2] /*2549*/;
  assign _16306_ = sum_30[23] & q[2] /*2548*/;
  assign _16307_ = m_30[23] & _16305_ /*2547*/;
  assign r_30[23] = _16307_ | _16306_ /*2546*/;
  assign _16308_ = ~q[2] /*2545*/;
  assign _16309_ = sum_30[24] & q[2] /*2544*/;
  assign _16310_ = m_30[24] & _16308_ /*2543*/;
  assign r_30[24] = _16310_ | _16309_ /*2542*/;
  assign _16311_ = ~q[2] /*2541*/;
  assign _16312_ = sum_30[25] & q[2] /*2540*/;
  assign _16313_ = m_30[25] & _16311_ /*2539*/;
  assign r_30[25] = _16313_ | _16312_ /*2538*/;
  assign _16314_ = ~q[2] /*2537*/;
  assign _16315_ = sum_30[26] & q[2] /*2536*/;
  assign _16316_ = m_30[26] & _16314_ /*2535*/;
  assign r_30[26] = _16316_ | _16315_ /*2534*/;
  assign _16317_ = ~q[2] /*2533*/;
  assign _16318_ = sum_30[27] & q[2] /*2532*/;
  assign _16319_ = m_30[27] & _16317_ /*2531*/;
  assign r_30[27] = _16319_ | _16318_ /*2530*/;
  assign _16320_ = ~q[2] /*2529*/;
  assign _16321_ = sum_30[28] & q[2] /*2528*/;
  assign _16322_ = m_30[28] & _16320_ /*2527*/;
  assign r_30[28] = _16322_ | _16321_ /*2526*/;
  assign _16323_ = ~q[2] /*2525*/;
  assign _16324_ = sum_30[29] & q[2] /*2524*/;
  assign _16325_ = m_30[29] & _16323_ /*2523*/;
  assign r_30[29] = _16325_ | _16324_ /*2522*/;
  assign _16326_ = ~q[2] /*2521*/;
  assign _16327_ = sum_30[30] & q[2] /*2520*/;
  assign _16328_ = m_30[30] & _16326_ /*2519*/;
  assign r_30[30] = _16328_ | _16327_ /*2518*/;
  assign _16329_ = ~q[2] /*2517*/;
  assign _16330_ = sum_30[31] & q[2] /*2516*/;
  assign _16331_ = m_30[31] & _16329_ /*2515*/;
  assign r_30[31] = _16331_ | _16330_ /*2514*/;
  assign _16332_ = ~q[2] /*2513*/;
  assign _16333_ = sum_30[32] & q[2] /*2512*/;
  assign _16334_ = m_30[32] & _16332_ /*2511*/;
  assign r_30[32] = _16334_ | _16333_ /*2510*/;
  assign _16335_ = ~q[2] /*2509*/;
  assign _16336_ = sum_30[33] & q[2] /*2508*/;
  assign _16337_ = m_30[33] & _16335_ /*2507*/;
  assign r_30[33] = _16337_ | _16336_ /*2506*/;
  assign _16338_ = ~q[2] /*2505*/;
  assign _16339_ = sum_30[34] & q[2] /*2504*/;
  assign _16340_ = m_30[34] & _16338_ /*2503*/;
  assign r_30[34] = _16340_ | _16339_ /*2502*/;
  assign _16341_ = ~q[2] /*2501*/;
  assign _16342_ = sum_30[35] & q[2] /*2500*/;
  assign _16343_ = m_30[35] & _16341_ /*2499*/;
  assign r_30[35] = _16343_ | _16342_ /*2498*/;
  assign _16344_ = ~q[2] /*2497*/;
  assign _16345_ = sum_30[36] & q[2] /*2496*/;
  assign _16346_ = m_30[36] & _16344_ /*2495*/;
  assign r_30[36] = _16346_ | _16345_ /*2494*/;
  assign _16347_ = ~q[2] /*2493*/;
  assign _16348_ = sum_30[37] & q[2] /*2492*/;
  assign _16349_ = m_30[37] & _16347_ /*2491*/;
  assign r_30[37] = _16349_ | _16348_ /*2490*/;
  assign _16350_ = ~q[2] /*2489*/;
  assign _16351_ = sum_30[38] & q[2] /*2488*/;
  assign _16352_ = m_30[38] & _16350_ /*2487*/;
  assign r_30[38] = _16352_ | _16351_ /*2486*/;
  assign _16353_ = ~q[2] /*2485*/;
  assign _16354_ = sum_30[39] & q[2] /*2484*/;
  assign _16355_ = m_30[39] & _16353_ /*2483*/;
  assign r_30[39] = _16355_ | _16354_ /*2482*/;
  assign _16356_ = ~q[2] /*2481*/;
  assign _16357_ = sum_30[40] & q[2] /*2480*/;
  assign _16358_ = m_30[40] & _16356_ /*2479*/;
  assign r_30[40] = _16358_ | _16357_ /*2478*/;
  assign _16359_ = ~q[2] /*2477*/;
  assign _16360_ = sum_30[41] & q[2] /*2476*/;
  assign _16361_ = m_30[41] & _16359_ /*2475*/;
  assign r_30[41] = _16361_ | _16360_ /*2474*/;
  assign _16362_ = ~q[2] /*2473*/;
  assign _16363_ = sum_30[42] & q[2] /*2472*/;
  assign _16364_ = m_30[42] & _16362_ /*2471*/;
  assign r_30[42] = _16364_ | _16363_ /*2470*/;
  assign _16365_ = ~q[2] /*2469*/;
  assign _16366_ = sum_30[43] & q[2] /*2468*/;
  assign _16367_ = m_30[43] & _16365_ /*2467*/;
  assign r_30[43] = _16367_ | _16366_ /*2466*/;
  assign _16368_ = ~q[2] /*2465*/;
  assign _16369_ = sum_30[44] & q[2] /*2464*/;
  assign _16370_ = m_30[44] & _16368_ /*2463*/;
  assign r_30[44] = _16370_ | _16369_ /*2462*/;
  assign _16371_ = ~q[2] /*2461*/;
  assign _16372_ = sum_30[45] & q[2] /*2460*/;
  assign _16373_ = m_30[45] & _16371_ /*2459*/;
  assign r_30[45] = _16373_ | _16372_ /*2458*/;
  assign _16374_ = ~q[2] /*2457*/;
  assign _16375_ = sum_30[46] & q[2] /*2456*/;
  assign _16376_ = m_30[46] & _16374_ /*2455*/;
  assign r_30[46] = _16376_ | _16375_ /*2454*/;
  assign _16377_ = ~q[2] /*2453*/;
  assign _16378_ = sum_30[47] & q[2] /*2452*/;
  assign _16379_ = m_30[47] & _16377_ /*2451*/;
  assign r_30[47] = _16379_ | _16378_ /*2450*/;
  assign _16380_ = ~q[2] /*2449*/;
  assign _16381_ = sum_30[48] & q[2] /*2448*/;
  assign _16382_ = m_30[48] & _16380_ /*2447*/;
  assign r_30[48] = _16382_ | _16381_ /*2446*/;
  assign _16383_ = ~q[2] /*2445*/;
  assign _16384_ = sum_30[49] & q[2] /*2444*/;
  assign _16385_ = m_30[49] & _16383_ /*2443*/;
  assign r_30[49] = _16385_ | _16384_ /*2442*/;
  assign _16386_ = ~q[2] /*2441*/;
  assign _16387_ = sum_30[50] & q[2] /*2440*/;
  assign _16388_ = m_30[50] & _16386_ /*2439*/;
  assign r_30[50] = _16388_ | _16387_ /*2438*/;
  assign _16389_ = ~q[2] /*2437*/;
  assign _16390_ = sum_30[51] & q[2] /*2436*/;
  assign _16391_ = m_30[51] & _16389_ /*2435*/;
  assign r_30[51] = _16391_ | _16390_ /*2434*/;
  assign _16392_ = ~q[2] /*2433*/;
  assign _16393_ = sum_30[52] & q[2] /*2432*/;
  assign _16394_ = m_30[52] & _16392_ /*2431*/;
  assign r_30[52] = _16394_ | _16393_ /*2430*/;
  assign _16395_ = ~q[2] /*2429*/;
  assign _16396_ = sum_30[53] & q[2] /*2428*/;
  assign _16397_ = m_30[53] & _16395_ /*2427*/;
  assign r_30[53] = _16397_ | _16396_ /*2426*/;
  assign _16398_ = ~q[2] /*2425*/;
  assign _16399_ = sum_30[54] & q[2] /*2424*/;
  assign _16400_ = m_30[54] & _16398_ /*2423*/;
  assign r_30[54] = _16400_ | _16399_ /*2422*/;
  assign _16401_ = ~q[2] /*2421*/;
  assign _16402_ = sum_30[55] & q[2] /*2420*/;
  assign _16403_ = m_30[55] & _16401_ /*2419*/;
  assign r_30[55] = _16403_ | _16402_ /*2418*/;
  assign _16404_ = ~q[2] /*2417*/;
  assign _16405_ = sum_30[56] & q[2] /*2416*/;
  assign _16406_ = m_30[56] & _16404_ /*2415*/;
  assign r_30[56] = _16406_ | _16405_ /*2414*/;
  assign _16407_ = ~q[2] /*2413*/;
  assign _16408_ = sum_30[57] & q[2] /*2412*/;
  assign _16409_ = m_30[57] & _16407_ /*2411*/;
  assign r_30[57] = _16409_ | _16408_ /*2410*/;
  assign _16410_ = ~q[2] /*2409*/;
  assign _16411_ = sum_30[58] & q[2] /*2408*/;
  assign _16412_ = m_30[58] & _16410_ /*2407*/;
  assign r_30[58] = _16412_ | _16411_ /*2406*/;
  assign _16413_ = ~q[2] /*2405*/;
  assign _16414_ = sum_30[59] & q[2] /*2404*/;
  assign _16415_ = m_30[59] & _16413_ /*2403*/;
  assign r_30[59] = _16415_ | _16414_ /*2402*/;
  assign _16416_ = ~q[2] /*2401*/;
  assign _16417_ = sum_30[60] & q[2] /*2400*/;
  assign _16418_ = m_30[60] & _16416_ /*2399*/;
  assign r_30[60] = _16418_ | _16417_ /*2398*/;
  assign _16419_ = ~q[2] /*2397*/;
  assign _16420_ = sum_30[61] & q[2] /*2396*/;
  assign _16421_ = m_30[61] & _16419_ /*2395*/;
  assign r_30[61] = _16421_ | _16420_ /*2394*/;
  assign _16422_ = ~q[2] /*2393*/;
  assign _16423_ = sum_30[62] & q[2] /*2392*/;
  assign _16424_ = m_30[62] & _16422_ /*2391*/;
  assign r_30[62] = _16424_ | _16423_ /*2390*/;
  assign _16425_ = ~q[2] /*2389*/;
  assign _16426_ = sum_30[63] & q[2] /*2388*/;
  assign _16427_ = m_30[63] & _16425_ /*2387*/;
  assign r_30[63] = _16427_ | _16426_ /*2386*/;
  assign _16428_ = ~q[2] /*2385*/;
  assign _16429_ = sum_30[64] & q[2] /*2384*/;
  assign _16430_ = m_30[64] & _16428_ /*2383*/;
  assign r_30[64] = _16430_ | _16429_ /*2382*/;
  assign _16431_ = ~q[2] /*2381*/;
  assign _16432_ = sum_30[65] & q[2] /*2380*/;
  assign _16433_ = m_30[65] & _16431_ /*2379*/;
  assign r_30[65] = _16433_ | _16432_ /*2378*/;
  assign _16434_ = ~q[2] /*2377*/;
  assign _16435_ = sum_30[66] & q[2] /*2376*/;
  assign _16436_ = m_30[66] & _16434_ /*2375*/;
  assign r_30[66] = _16436_ | _16435_ /*2374*/;
  assign _16437_ = ~q[2] /*2373*/;
  assign _16438_ = sum_30[67] & q[2] /*2372*/;
  assign _16439_ = m_30[67] & _16437_ /*2371*/;
  assign r_30[67] = _16439_ | _16438_ /*2370*/;
  assign _16440_ = ~q[2] /*2369*/;
  assign _16441_ = sum_30[68] & q[2] /*2368*/;
  assign _16442_ = m_30[68] & _16440_ /*2367*/;
  assign r_30[68] = _16442_ | _16441_ /*2366*/;
  assign _16443_ = ~q[2] /*2365*/;
  assign _16444_ = sum_30[69] & q[2] /*2364*/;
  assign _16445_ = m_30[69] & _16443_ /*2363*/;
  assign r_30[69] = _16445_ | _16444_ /*2362*/;
  assign _16446_ = ~q[2] /*2361*/;
  assign _16447_ = sum_30[70] & q[2] /*2360*/;
  assign _16448_ = m_30[70] & _16446_ /*2359*/;
  assign r_30[70] = _16448_ | _16447_ /*2358*/;
  assign _16449_ = ~q[2] /*2357*/;
  assign _16450_ = sum_30[71] & q[2] /*2356*/;
  assign _16451_ = m_30[71] & _16449_ /*2355*/;
  assign r_30[71] = _16451_ | _16450_ /*2354*/;
  assign _16452_ = ~q[2] /*2353*/;
  assign _16453_ = sum_30[72] & q[2] /*2352*/;
  assign _16454_ = m_30[72] & _16452_ /*2351*/;
  assign r_30[72] = _16454_ | _16453_ /*2350*/;
  assign _16455_ = ~q[2] /*2349*/;
  assign _16456_ = sum_30[73] & q[2] /*2348*/;
  assign _16457_ = m_30[73] & _16455_ /*2347*/;
  assign r_30[73] = _16457_ | _16456_ /*2346*/;
  assign _16458_ = ~q[2] /*2345*/;
  assign _16459_ = sum_30[74] & q[2] /*2344*/;
  assign _16460_ = m_30[74] & _16458_ /*2343*/;
  assign r_30[74] = _16460_ | _16459_ /*2342*/;
  assign _16461_ = ~q[2] /*2341*/;
  assign _16462_ = sum_30[75] & q[2] /*2340*/;
  assign _16463_ = m_30[75] & _16461_ /*2339*/;
  assign r_30[75] = _16463_ | _16462_ /*2338*/;
  assign _16464_ = ~q[2] /*2337*/;
  assign _16465_ = sum_30[76] & q[2] /*2336*/;
  assign _16466_ = m_30[76] & _16464_ /*2335*/;
  assign r_30[76] = _16466_ | _16465_ /*2334*/;
  assign _16467_ = ~q[2] /*2333*/;
  assign _16468_ = sum_30[77] & q[2] /*2332*/;
  assign _16469_ = m_30[77] & _16467_ /*2331*/;
  assign r_30[77] = _16469_ | _16468_ /*2330*/;
  assign _16470_ = ~q[2] /*2329*/;
  assign _16471_ = sum_30[78] & q[2] /*2328*/;
  assign _16472_ = m_30[78] & _16470_ /*2327*/;
  assign r_30[78] = _16472_ | _16471_ /*2326*/;
  assign _16473_ = ~q[2] /*2325*/;
  assign _16474_ = sum_30[79] & q[2] /*2324*/;
  assign _16475_ = m_30[79] & _16473_ /*2323*/;
  assign r_30[79] = _16475_ | _16474_ /*2322*/;
  assign _16476_ = ~q[2] /*2321*/;
  assign _16477_ = sum_30[80] & q[2] /*2320*/;
  assign _16478_ = m_30[80] & _16476_ /*2319*/;
  assign r_30[80] = _16478_ | _16477_ /*2318*/;
  assign _16479_ = ~q[2] /*2317*/;
  assign _16480_ = sum_30[81] & q[2] /*2316*/;
  assign _16481_ = m_30[81] & _16479_ /*2315*/;
  assign r_30[81] = _16481_ | _16480_ /*2314*/;
  assign _16482_ = ~q[2] /*2313*/;
  assign _16483_ = sum_30[82] & q[2] /*2312*/;
  assign _16484_ = m_30[82] & _16482_ /*2311*/;
  assign r_30[82] = _16484_ | _16483_ /*2310*/;
  assign _16485_ = ~q[2] /*2309*/;
  assign _16486_ = sum_30[83] & q[2] /*2308*/;
  assign _16487_ = m_30[83] & _16485_ /*2307*/;
  assign r_30[83] = _16487_ | _16486_ /*2306*/;
  assign _16488_ = ~q[2] /*2305*/;
  assign _16489_ = sum_30[84] & q[2] /*2304*/;
  assign _16490_ = m_30[84] & _16488_ /*2303*/;
  assign r_30[84] = _16490_ | _16489_ /*2302*/;
  assign _16491_ = ~q[2] /*2301*/;
  assign _16492_ = sum_30[85] & q[2] /*2300*/;
  assign _16493_ = m_30[85] & _16491_ /*2299*/;
  assign r_30[85] = _16493_ | _16492_ /*2298*/;
  assign _16494_ = ~q[2] /*2297*/;
  assign _16495_ = sum_30[86] & q[2] /*2296*/;
  assign _16496_ = m_30[86] & _16494_ /*2295*/;
  assign r_30[86] = _16496_ | _16495_ /*2294*/;
  assign _16497_ = ~q[2] /*2293*/;
  assign _16498_ = sum_30[87] & q[2] /*2292*/;
  assign _16499_ = m_30[87] & _16497_ /*2291*/;
  assign r_30[87] = _16499_ | _16498_ /*2290*/;
  assign _16500_ = ~q[2] /*2289*/;
  assign _16501_ = sum_30[88] & q[2] /*2288*/;
  assign _16502_ = m_30[88] & _16500_ /*2287*/;
  assign r_30[88] = _16502_ | _16501_ /*2286*/;
  assign _16503_ = ~q[2] /*2285*/;
  assign _16504_ = sum_30[89] & q[2] /*2284*/;
  assign _16505_ = m_30[89] & _16503_ /*2283*/;
  assign r_30[89] = _16505_ | _16504_ /*2282*/;
  assign _16506_ = ~q[2] /*2281*/;
  assign _16507_ = sum_30[90] & q[2] /*2280*/;
  assign _16508_ = m_30[90] & _16506_ /*2279*/;
  assign r_30[90] = _16508_ | _16507_ /*2278*/;
  assign _16509_ = ~q[2] /*2277*/;
  assign _16510_ = sum_30[91] & q[2] /*2276*/;
  assign _16511_ = m_30[91] & _16509_ /*2275*/;
  assign r_30[91] = _16511_ | _16510_ /*2274*/;
  assign _16512_ = ~q[2] /*2273*/;
  assign _16513_ = sum_30[92] & q[2] /*2272*/;
  assign _16514_ = m_30[92] & _16512_ /*2271*/;
  assign r_30[92] = _16514_ | _16513_ /*2270*/;
  assign inv_31[0] = oneWire /*2216*/;
  assign inv_31[1] = ~div[0] /*2210*/;
  assign inv_31[2] = ~div[1] /*2204*/;
  assign inv_31[3] = ~div[2] /*2198*/;
  assign inv_31[4] = ~div[3] /*2192*/;
  assign inv_31[5] = ~div[4] /*2186*/;
  assign inv_31[6] = ~div[5] /*2180*/;
  assign inv_31[7] = ~div[6] /*2174*/;
  assign inv_31[8] = ~div[7] /*2168*/;
  assign inv_31[9] = ~div[8] /*2162*/;
  assign inv_31[10] = ~div[9] /*2156*/;
  assign inv_31[11] = ~div[10] /*2150*/;
  assign inv_31[12] = ~div[11] /*2144*/;
  assign inv_31[13] = ~div[12] /*2138*/;
  assign inv_31[14] = ~div[13] /*2132*/;
  assign inv_31[15] = ~div[14] /*2126*/;
  assign inv_31[16] = ~div[15] /*2120*/;
  assign inv_31[17] = ~div[16] /*2114*/;
  assign inv_31[18] = ~div[17] /*2108*/;
  assign inv_31[19] = ~div[18] /*2102*/;
  assign inv_31[20] = ~div[19] /*2096*/;
  assign inv_31[21] = ~div[20] /*2090*/;
  assign inv_31[22] = ~div[21] /*2084*/;
  assign inv_31[23] = ~div[22] /*2078*/;
  assign inv_31[24] = ~div[23] /*2072*/;
  assign inv_31[25] = ~div[24] /*2066*/;
  assign inv_31[26] = ~div[25] /*2060*/;
  assign inv_31[27] = ~div[26] /*2054*/;
  assign inv_31[28] = ~div[27] /*2048*/;
  assign inv_31[29] = ~div[28] /*2042*/;
  assign inv_31[30] = ~div[29] /*2036*/;
  assign inv_31[31] = ~div[30] /*2030*/;
  assign inv_31[32] = oneWire /*2024*/;
  assign inv_31[33] = oneWire /*2018*/;
  assign inv_31[34] = oneWire /*2012*/;
  assign inv_31[35] = oneWire /*2006*/;
  assign inv_31[36] = oneWire /*2000*/;
  assign inv_31[37] = oneWire /*1994*/;
  assign inv_31[38] = oneWire /*1988*/;
  assign inv_31[39] = oneWire /*1982*/;
  assign inv_31[40] = oneWire /*1976*/;
  assign inv_31[41] = oneWire /*1970*/;
  assign inv_31[42] = oneWire /*1964*/;
  assign inv_31[43] = oneWire /*1958*/;
  assign inv_31[44] = oneWire /*1952*/;
  assign inv_31[45] = oneWire /*1946*/;
  assign inv_31[46] = oneWire /*1940*/;
  assign inv_31[47] = oneWire /*1934*/;
  assign inv_31[48] = oneWire /*1928*/;
  assign inv_31[49] = oneWire /*1922*/;
  assign inv_31[50] = oneWire /*1916*/;
  assign inv_31[51] = oneWire /*1910*/;
  assign inv_31[52] = oneWire /*1904*/;
  assign inv_31[53] = oneWire /*1898*/;
  assign inv_31[54] = oneWire /*1892*/;
  assign inv_31[55] = oneWire /*1886*/;
  assign inv_31[56] = oneWire /*1880*/;
  assign inv_31[57] = oneWire /*1874*/;
  assign inv_31[58] = oneWire /*1868*/;
  assign inv_31[59] = oneWire /*1862*/;
  assign inv_31[60] = oneWire /*1856*/;
  assign inv_31[61] = oneWire /*1850*/;
  assign inv_31[62] = oneWire /*1844*/;
  assign inv_31[63] = oneWire /*1838*/;
  assign inv_31[64] = oneWire /*1832*/;
  assign inv_31[65] = oneWire /*1826*/;
  assign inv_31[66] = oneWire /*1820*/;
  assign inv_31[67] = oneWire /*1814*/;
  assign inv_31[68] = oneWire /*1808*/;
  assign inv_31[69] = oneWire /*1802*/;
  assign inv_31[70] = oneWire /*1796*/;
  assign inv_31[71] = oneWire /*1790*/;
  assign inv_31[72] = oneWire /*1784*/;
  assign inv_31[73] = oneWire /*1778*/;
  assign inv_31[74] = oneWire /*1772*/;
  assign inv_31[75] = oneWire /*1766*/;
  assign inv_31[76] = oneWire /*1760*/;
  assign inv_31[77] = oneWire /*1754*/;
  assign inv_31[78] = oneWire /*1748*/;
  assign inv_31[79] = oneWire /*1742*/;
  assign inv_31[80] = oneWire /*1736*/;
  assign inv_31[81] = oneWire /*1730*/;
  assign inv_31[82] = oneWire /*1724*/;
  assign inv_31[83] = oneWire /*1718*/;
  assign inv_31[84] = oneWire /*1712*/;
  assign inv_31[85] = oneWire /*1706*/;
  assign inv_31[86] = oneWire /*1700*/;
  assign inv_31[87] = oneWire /*1694*/;
  assign inv_31[88] = oneWire /*1688*/;
  assign inv_31[89] = oneWire /*1682*/;
  assign inv_31[90] = oneWire /*1676*/;
  assign inv_31[91] = oneWire /*1670*/;
  assign inv_31[92] = oneWire /*1664*/;
  assign _16515_ = inv_31[0] ^ r_30[0] /*2215*/;
  assign sum_31[0] = _16515_ ^ oneWire /*2214*/;
  assign _16516_ = _16515_ & oneWire /*2213*/;
  assign _16517_ = inv_31[0] & r_30[0] /*2212*/;
  assign _16518_ = _16516_ | _16517_ /*2211*/;
  assign _16519_ = inv_31[1] ^ r_30[1] /*2209*/;
  assign sum_31[1] = _16519_ ^ _16518_ /*2208*/;
  assign _16520_ = _16519_ & _16518_ /*2207*/;
  assign _16521_ = inv_31[1] & r_30[1] /*2206*/;
  assign _16522_ = _16520_ | _16521_ /*2205*/;
  assign _16523_ = inv_31[2] ^ r_30[2] /*2203*/;
  assign sum_31[2] = _16523_ ^ _16522_ /*2202*/;
  assign _16524_ = _16523_ & _16522_ /*2201*/;
  assign _16525_ = inv_31[2] & r_30[2] /*2200*/;
  assign _16526_ = _16524_ | _16525_ /*2199*/;
  assign _16527_ = inv_31[3] ^ r_30[3] /*2197*/;
  assign sum_31[3] = _16527_ ^ _16526_ /*2196*/;
  assign _16528_ = _16527_ & _16526_ /*2195*/;
  assign _16529_ = inv_31[3] & r_30[3] /*2194*/;
  assign _16530_ = _16528_ | _16529_ /*2193*/;
  assign _16531_ = inv_31[4] ^ r_30[4] /*2191*/;
  assign sum_31[4] = _16531_ ^ _16530_ /*2190*/;
  assign _16532_ = _16531_ & _16530_ /*2189*/;
  assign _16533_ = inv_31[4] & r_30[4] /*2188*/;
  assign _16534_ = _16532_ | _16533_ /*2187*/;
  assign _16535_ = inv_31[5] ^ r_30[5] /*2185*/;
  assign sum_31[5] = _16535_ ^ _16534_ /*2184*/;
  assign _16536_ = _16535_ & _16534_ /*2183*/;
  assign _16537_ = inv_31[5] & r_30[5] /*2182*/;
  assign _16538_ = _16536_ | _16537_ /*2181*/;
  assign _16539_ = inv_31[6] ^ r_30[6] /*2179*/;
  assign sum_31[6] = _16539_ ^ _16538_ /*2178*/;
  assign _16540_ = _16539_ & _16538_ /*2177*/;
  assign _16541_ = inv_31[6] & r_30[6] /*2176*/;
  assign _16542_ = _16540_ | _16541_ /*2175*/;
  assign _16543_ = inv_31[7] ^ r_30[7] /*2173*/;
  assign sum_31[7] = _16543_ ^ _16542_ /*2172*/;
  assign _16544_ = _16543_ & _16542_ /*2171*/;
  assign _16545_ = inv_31[7] & r_30[7] /*2170*/;
  assign _16546_ = _16544_ | _16545_ /*2169*/;
  assign _16547_ = inv_31[8] ^ r_30[8] /*2167*/;
  assign sum_31[8] = _16547_ ^ _16546_ /*2166*/;
  assign _16548_ = _16547_ & _16546_ /*2165*/;
  assign _16549_ = inv_31[8] & r_30[8] /*2164*/;
  assign _16550_ = _16548_ | _16549_ /*2163*/;
  assign _16551_ = inv_31[9] ^ r_30[9] /*2161*/;
  assign sum_31[9] = _16551_ ^ _16550_ /*2160*/;
  assign _16552_ = _16551_ & _16550_ /*2159*/;
  assign _16553_ = inv_31[9] & r_30[9] /*2158*/;
  assign _16554_ = _16552_ | _16553_ /*2157*/;
  assign _16555_ = inv_31[10] ^ r_30[10] /*2155*/;
  assign sum_31[10] = _16555_ ^ _16554_ /*2154*/;
  assign _16556_ = _16555_ & _16554_ /*2153*/;
  assign _16557_ = inv_31[10] & r_30[10] /*2152*/;
  assign _16558_ = _16556_ | _16557_ /*2151*/;
  assign _16559_ = inv_31[11] ^ r_30[11] /*2149*/;
  assign sum_31[11] = _16559_ ^ _16558_ /*2148*/;
  assign _16560_ = _16559_ & _16558_ /*2147*/;
  assign _16561_ = inv_31[11] & r_30[11] /*2146*/;
  assign _16562_ = _16560_ | _16561_ /*2145*/;
  assign _16563_ = inv_31[12] ^ r_30[12] /*2143*/;
  assign sum_31[12] = _16563_ ^ _16562_ /*2142*/;
  assign _16564_ = _16563_ & _16562_ /*2141*/;
  assign _16565_ = inv_31[12] & r_30[12] /*2140*/;
  assign _16566_ = _16564_ | _16565_ /*2139*/;
  assign _16567_ = inv_31[13] ^ r_30[13] /*2137*/;
  assign sum_31[13] = _16567_ ^ _16566_ /*2136*/;
  assign _16568_ = _16567_ & _16566_ /*2135*/;
  assign _16569_ = inv_31[13] & r_30[13] /*2134*/;
  assign _16570_ = _16568_ | _16569_ /*2133*/;
  assign _16571_ = inv_31[14] ^ r_30[14] /*2131*/;
  assign sum_31[14] = _16571_ ^ _16570_ /*2130*/;
  assign _16572_ = _16571_ & _16570_ /*2129*/;
  assign _16573_ = inv_31[14] & r_30[14] /*2128*/;
  assign _16574_ = _16572_ | _16573_ /*2127*/;
  assign _16575_ = inv_31[15] ^ r_30[15] /*2125*/;
  assign sum_31[15] = _16575_ ^ _16574_ /*2124*/;
  assign _16576_ = _16575_ & _16574_ /*2123*/;
  assign _16577_ = inv_31[15] & r_30[15] /*2122*/;
  assign _16578_ = _16576_ | _16577_ /*2121*/;
  assign _16579_ = inv_31[16] ^ r_30[16] /*2119*/;
  assign sum_31[16] = _16579_ ^ _16578_ /*2118*/;
  assign _16580_ = _16579_ & _16578_ /*2117*/;
  assign _16581_ = inv_31[16] & r_30[16] /*2116*/;
  assign _16582_ = _16580_ | _16581_ /*2115*/;
  assign _16583_ = inv_31[17] ^ r_30[17] /*2113*/;
  assign sum_31[17] = _16583_ ^ _16582_ /*2112*/;
  assign _16584_ = _16583_ & _16582_ /*2111*/;
  assign _16585_ = inv_31[17] & r_30[17] /*2110*/;
  assign _16586_ = _16584_ | _16585_ /*2109*/;
  assign _16587_ = inv_31[18] ^ r_30[18] /*2107*/;
  assign sum_31[18] = _16587_ ^ _16586_ /*2106*/;
  assign _16588_ = _16587_ & _16586_ /*2105*/;
  assign _16589_ = inv_31[18] & r_30[18] /*2104*/;
  assign _16590_ = _16588_ | _16589_ /*2103*/;
  assign _16591_ = inv_31[19] ^ r_30[19] /*2101*/;
  assign sum_31[19] = _16591_ ^ _16590_ /*2100*/;
  assign _16592_ = _16591_ & _16590_ /*2099*/;
  assign _16593_ = inv_31[19] & r_30[19] /*2098*/;
  assign _16594_ = _16592_ | _16593_ /*2097*/;
  assign _16595_ = inv_31[20] ^ r_30[20] /*2095*/;
  assign sum_31[20] = _16595_ ^ _16594_ /*2094*/;
  assign _16596_ = _16595_ & _16594_ /*2093*/;
  assign _16597_ = inv_31[20] & r_30[20] /*2092*/;
  assign _16598_ = _16596_ | _16597_ /*2091*/;
  assign _16599_ = inv_31[21] ^ r_30[21] /*2089*/;
  assign sum_31[21] = _16599_ ^ _16598_ /*2088*/;
  assign _16600_ = _16599_ & _16598_ /*2087*/;
  assign _16601_ = inv_31[21] & r_30[21] /*2086*/;
  assign _16602_ = _16600_ | _16601_ /*2085*/;
  assign _16603_ = inv_31[22] ^ r_30[22] /*2083*/;
  assign sum_31[22] = _16603_ ^ _16602_ /*2082*/;
  assign _16604_ = _16603_ & _16602_ /*2081*/;
  assign _16605_ = inv_31[22] & r_30[22] /*2080*/;
  assign _16606_ = _16604_ | _16605_ /*2079*/;
  assign _16607_ = inv_31[23] ^ r_30[23] /*2077*/;
  assign sum_31[23] = _16607_ ^ _16606_ /*2076*/;
  assign _16608_ = _16607_ & _16606_ /*2075*/;
  assign _16609_ = inv_31[23] & r_30[23] /*2074*/;
  assign _16610_ = _16608_ | _16609_ /*2073*/;
  assign _16611_ = inv_31[24] ^ r_30[24] /*2071*/;
  assign sum_31[24] = _16611_ ^ _16610_ /*2070*/;
  assign _16612_ = _16611_ & _16610_ /*2069*/;
  assign _16613_ = inv_31[24] & r_30[24] /*2068*/;
  assign _16614_ = _16612_ | _16613_ /*2067*/;
  assign _16615_ = inv_31[25] ^ r_30[25] /*2065*/;
  assign sum_31[25] = _16615_ ^ _16614_ /*2064*/;
  assign _16616_ = _16615_ & _16614_ /*2063*/;
  assign _16617_ = inv_31[25] & r_30[25] /*2062*/;
  assign _16618_ = _16616_ | _16617_ /*2061*/;
  assign _16619_ = inv_31[26] ^ r_30[26] /*2059*/;
  assign sum_31[26] = _16619_ ^ _16618_ /*2058*/;
  assign _16620_ = _16619_ & _16618_ /*2057*/;
  assign _16621_ = inv_31[26] & r_30[26] /*2056*/;
  assign _16622_ = _16620_ | _16621_ /*2055*/;
  assign _16623_ = inv_31[27] ^ r_30[27] /*2053*/;
  assign sum_31[27] = _16623_ ^ _16622_ /*2052*/;
  assign _16624_ = _16623_ & _16622_ /*2051*/;
  assign _16625_ = inv_31[27] & r_30[27] /*2050*/;
  assign _16626_ = _16624_ | _16625_ /*2049*/;
  assign _16627_ = inv_31[28] ^ r_30[28] /*2047*/;
  assign sum_31[28] = _16627_ ^ _16626_ /*2046*/;
  assign _16628_ = _16627_ & _16626_ /*2045*/;
  assign _16629_ = inv_31[28] & r_30[28] /*2044*/;
  assign _16630_ = _16628_ | _16629_ /*2043*/;
  assign _16631_ = inv_31[29] ^ r_30[29] /*2041*/;
  assign sum_31[29] = _16631_ ^ _16630_ /*2040*/;
  assign _16632_ = _16631_ & _16630_ /*2039*/;
  assign _16633_ = inv_31[29] & r_30[29] /*2038*/;
  assign _16634_ = _16632_ | _16633_ /*2037*/;
  assign _16635_ = inv_31[30] ^ r_30[30] /*2035*/;
  assign sum_31[30] = _16635_ ^ _16634_ /*2034*/;
  assign _16636_ = _16635_ & _16634_ /*2033*/;
  assign _16637_ = inv_31[30] & r_30[30] /*2032*/;
  assign _16638_ = _16636_ | _16637_ /*2031*/;
  assign _16639_ = inv_31[31] ^ r_30[31] /*2029*/;
  assign sum_31[31] = _16639_ ^ _16638_ /*2028*/;
  assign _16640_ = _16639_ & _16638_ /*2027*/;
  assign _16641_ = inv_31[31] & r_30[31] /*2026*/;
  assign _16642_ = _16640_ | _16641_ /*2025*/;
  assign _16643_ = inv_31[32] ^ r_30[32] /*2023*/;
  assign sum_31[32] = _16643_ ^ _16642_ /*2022*/;
  assign _16644_ = _16643_ & _16642_ /*2021*/;
  assign _16645_ = inv_31[32] & r_30[32] /*2020*/;
  assign _16646_ = _16644_ | _16645_ /*2019*/;
  assign _16647_ = inv_31[33] ^ r_30[33] /*2017*/;
  assign sum_31[33] = _16647_ ^ _16646_ /*2016*/;
  assign _16648_ = _16647_ & _16646_ /*2015*/;
  assign _16649_ = inv_31[33] & r_30[33] /*2014*/;
  assign _16650_ = _16648_ | _16649_ /*2013*/;
  assign _16651_ = inv_31[34] ^ r_30[34] /*2011*/;
  assign sum_31[34] = _16651_ ^ _16650_ /*2010*/;
  assign _16652_ = _16651_ & _16650_ /*2009*/;
  assign _16653_ = inv_31[34] & r_30[34] /*2008*/;
  assign _16654_ = _16652_ | _16653_ /*2007*/;
  assign _16655_ = inv_31[35] ^ r_30[35] /*2005*/;
  assign sum_31[35] = _16655_ ^ _16654_ /*2004*/;
  assign _16656_ = _16655_ & _16654_ /*2003*/;
  assign _16657_ = inv_31[35] & r_30[35] /*2002*/;
  assign _16658_ = _16656_ | _16657_ /*2001*/;
  assign _16659_ = inv_31[36] ^ r_30[36] /*1999*/;
  assign sum_31[36] = _16659_ ^ _16658_ /*1998*/;
  assign _16660_ = _16659_ & _16658_ /*1997*/;
  assign _16661_ = inv_31[36] & r_30[36] /*1996*/;
  assign _16662_ = _16660_ | _16661_ /*1995*/;
  assign _16663_ = inv_31[37] ^ r_30[37] /*1993*/;
  assign sum_31[37] = _16663_ ^ _16662_ /*1992*/;
  assign _16664_ = _16663_ & _16662_ /*1991*/;
  assign _16665_ = inv_31[37] & r_30[37] /*1990*/;
  assign _16666_ = _16664_ | _16665_ /*1989*/;
  assign _16667_ = inv_31[38] ^ r_30[38] /*1987*/;
  assign sum_31[38] = _16667_ ^ _16666_ /*1986*/;
  assign _16668_ = _16667_ & _16666_ /*1985*/;
  assign _16669_ = inv_31[38] & r_30[38] /*1984*/;
  assign _16670_ = _16668_ | _16669_ /*1983*/;
  assign _16671_ = inv_31[39] ^ r_30[39] /*1981*/;
  assign sum_31[39] = _16671_ ^ _16670_ /*1980*/;
  assign _16672_ = _16671_ & _16670_ /*1979*/;
  assign _16673_ = inv_31[39] & r_30[39] /*1978*/;
  assign _16674_ = _16672_ | _16673_ /*1977*/;
  assign _16675_ = inv_31[40] ^ r_30[40] /*1975*/;
  assign sum_31[40] = _16675_ ^ _16674_ /*1974*/;
  assign _16676_ = _16675_ & _16674_ /*1973*/;
  assign _16677_ = inv_31[40] & r_30[40] /*1972*/;
  assign _16678_ = _16676_ | _16677_ /*1971*/;
  assign _16679_ = inv_31[41] ^ r_30[41] /*1969*/;
  assign sum_31[41] = _16679_ ^ _16678_ /*1968*/;
  assign _16680_ = _16679_ & _16678_ /*1967*/;
  assign _16681_ = inv_31[41] & r_30[41] /*1966*/;
  assign _16682_ = _16680_ | _16681_ /*1965*/;
  assign _16683_ = inv_31[42] ^ r_30[42] /*1963*/;
  assign sum_31[42] = _16683_ ^ _16682_ /*1962*/;
  assign _16684_ = _16683_ & _16682_ /*1961*/;
  assign _16685_ = inv_31[42] & r_30[42] /*1960*/;
  assign _16686_ = _16684_ | _16685_ /*1959*/;
  assign _16687_ = inv_31[43] ^ r_30[43] /*1957*/;
  assign sum_31[43] = _16687_ ^ _16686_ /*1956*/;
  assign _16688_ = _16687_ & _16686_ /*1955*/;
  assign _16689_ = inv_31[43] & r_30[43] /*1954*/;
  assign _16690_ = _16688_ | _16689_ /*1953*/;
  assign _16691_ = inv_31[44] ^ r_30[44] /*1951*/;
  assign sum_31[44] = _16691_ ^ _16690_ /*1950*/;
  assign _16692_ = _16691_ & _16690_ /*1949*/;
  assign _16693_ = inv_31[44] & r_30[44] /*1948*/;
  assign _16694_ = _16692_ | _16693_ /*1947*/;
  assign _16695_ = inv_31[45] ^ r_30[45] /*1945*/;
  assign sum_31[45] = _16695_ ^ _16694_ /*1944*/;
  assign _16696_ = _16695_ & _16694_ /*1943*/;
  assign _16697_ = inv_31[45] & r_30[45] /*1942*/;
  assign _16698_ = _16696_ | _16697_ /*1941*/;
  assign _16699_ = inv_31[46] ^ r_30[46] /*1939*/;
  assign sum_31[46] = _16699_ ^ _16698_ /*1938*/;
  assign _16700_ = _16699_ & _16698_ /*1937*/;
  assign _16701_ = inv_31[46] & r_30[46] /*1936*/;
  assign _16702_ = _16700_ | _16701_ /*1935*/;
  assign _16703_ = inv_31[47] ^ r_30[47] /*1933*/;
  assign sum_31[47] = _16703_ ^ _16702_ /*1932*/;
  assign _16704_ = _16703_ & _16702_ /*1931*/;
  assign _16705_ = inv_31[47] & r_30[47] /*1930*/;
  assign _16706_ = _16704_ | _16705_ /*1929*/;
  assign _16707_ = inv_31[48] ^ r_30[48] /*1927*/;
  assign sum_31[48] = _16707_ ^ _16706_ /*1926*/;
  assign _16708_ = _16707_ & _16706_ /*1925*/;
  assign _16709_ = inv_31[48] & r_30[48] /*1924*/;
  assign _16710_ = _16708_ | _16709_ /*1923*/;
  assign _16711_ = inv_31[49] ^ r_30[49] /*1921*/;
  assign sum_31[49] = _16711_ ^ _16710_ /*1920*/;
  assign _16712_ = _16711_ & _16710_ /*1919*/;
  assign _16713_ = inv_31[49] & r_30[49] /*1918*/;
  assign _16714_ = _16712_ | _16713_ /*1917*/;
  assign _16715_ = inv_31[50] ^ r_30[50] /*1915*/;
  assign sum_31[50] = _16715_ ^ _16714_ /*1914*/;
  assign _16716_ = _16715_ & _16714_ /*1913*/;
  assign _16717_ = inv_31[50] & r_30[50] /*1912*/;
  assign _16718_ = _16716_ | _16717_ /*1911*/;
  assign _16719_ = inv_31[51] ^ r_30[51] /*1909*/;
  assign sum_31[51] = _16719_ ^ _16718_ /*1908*/;
  assign _16720_ = _16719_ & _16718_ /*1907*/;
  assign _16721_ = inv_31[51] & r_30[51] /*1906*/;
  assign _16722_ = _16720_ | _16721_ /*1905*/;
  assign _16723_ = inv_31[52] ^ r_30[52] /*1903*/;
  assign sum_31[52] = _16723_ ^ _16722_ /*1902*/;
  assign _16724_ = _16723_ & _16722_ /*1901*/;
  assign _16725_ = inv_31[52] & r_30[52] /*1900*/;
  assign _16726_ = _16724_ | _16725_ /*1899*/;
  assign _16727_ = inv_31[53] ^ r_30[53] /*1897*/;
  assign sum_31[53] = _16727_ ^ _16726_ /*1896*/;
  assign _16728_ = _16727_ & _16726_ /*1895*/;
  assign _16729_ = inv_31[53] & r_30[53] /*1894*/;
  assign _16730_ = _16728_ | _16729_ /*1893*/;
  assign _16731_ = inv_31[54] ^ r_30[54] /*1891*/;
  assign sum_31[54] = _16731_ ^ _16730_ /*1890*/;
  assign _16732_ = _16731_ & _16730_ /*1889*/;
  assign _16733_ = inv_31[54] & r_30[54] /*1888*/;
  assign _16734_ = _16732_ | _16733_ /*1887*/;
  assign _16735_ = inv_31[55] ^ r_30[55] /*1885*/;
  assign sum_31[55] = _16735_ ^ _16734_ /*1884*/;
  assign _16736_ = _16735_ & _16734_ /*1883*/;
  assign _16737_ = inv_31[55] & r_30[55] /*1882*/;
  assign _16738_ = _16736_ | _16737_ /*1881*/;
  assign _16739_ = inv_31[56] ^ r_30[56] /*1879*/;
  assign sum_31[56] = _16739_ ^ _16738_ /*1878*/;
  assign _16740_ = _16739_ & _16738_ /*1877*/;
  assign _16741_ = inv_31[56] & r_30[56] /*1876*/;
  assign _16742_ = _16740_ | _16741_ /*1875*/;
  assign _16743_ = inv_31[57] ^ r_30[57] /*1873*/;
  assign sum_31[57] = _16743_ ^ _16742_ /*1872*/;
  assign _16744_ = _16743_ & _16742_ /*1871*/;
  assign _16745_ = inv_31[57] & r_30[57] /*1870*/;
  assign _16746_ = _16744_ | _16745_ /*1869*/;
  assign _16747_ = inv_31[58] ^ r_30[58] /*1867*/;
  assign sum_31[58] = _16747_ ^ _16746_ /*1866*/;
  assign _16748_ = _16747_ & _16746_ /*1865*/;
  assign _16749_ = inv_31[58] & r_30[58] /*1864*/;
  assign _16750_ = _16748_ | _16749_ /*1863*/;
  assign _16751_ = inv_31[59] ^ r_30[59] /*1861*/;
  assign sum_31[59] = _16751_ ^ _16750_ /*1860*/;
  assign _16752_ = _16751_ & _16750_ /*1859*/;
  assign _16753_ = inv_31[59] & r_30[59] /*1858*/;
  assign _16754_ = _16752_ | _16753_ /*1857*/;
  assign _16755_ = inv_31[60] ^ r_30[60] /*1855*/;
  assign sum_31[60] = _16755_ ^ _16754_ /*1854*/;
  assign _16756_ = _16755_ & _16754_ /*1853*/;
  assign _16757_ = inv_31[60] & r_30[60] /*1852*/;
  assign _16758_ = _16756_ | _16757_ /*1851*/;
  assign _16759_ = inv_31[61] ^ r_30[61] /*1849*/;
  assign sum_31[61] = _16759_ ^ _16758_ /*1848*/;
  assign _16760_ = _16759_ & _16758_ /*1847*/;
  assign _16761_ = inv_31[61] & r_30[61] /*1846*/;
  assign _16762_ = _16760_ | _16761_ /*1845*/;
  assign _16763_ = inv_31[62] ^ r_30[62] /*1843*/;
  assign sum_31[62] = _16763_ ^ _16762_ /*1842*/;
  assign _16764_ = _16763_ & _16762_ /*1841*/;
  assign _16765_ = inv_31[62] & r_30[62] /*1840*/;
  assign _16766_ = _16764_ | _16765_ /*1839*/;
  assign _16767_ = inv_31[63] ^ r_30[63] /*1837*/;
  assign sum_31[63] = _16767_ ^ _16766_ /*1836*/;
  assign _16768_ = _16767_ & _16766_ /*1835*/;
  assign _16769_ = inv_31[63] & r_30[63] /*1834*/;
  assign _16770_ = _16768_ | _16769_ /*1833*/;
  assign _16771_ = inv_31[64] ^ r_30[64] /*1831*/;
  assign sum_31[64] = _16771_ ^ _16770_ /*1830*/;
  assign _16772_ = _16771_ & _16770_ /*1829*/;
  assign _16773_ = inv_31[64] & r_30[64] /*1828*/;
  assign _16774_ = _16772_ | _16773_ /*1827*/;
  assign _16775_ = inv_31[65] ^ r_30[65] /*1825*/;
  assign sum_31[65] = _16775_ ^ _16774_ /*1824*/;
  assign _16776_ = _16775_ & _16774_ /*1823*/;
  assign _16777_ = inv_31[65] & r_30[65] /*1822*/;
  assign _16778_ = _16776_ | _16777_ /*1821*/;
  assign _16779_ = inv_31[66] ^ r_30[66] /*1819*/;
  assign sum_31[66] = _16779_ ^ _16778_ /*1818*/;
  assign _16780_ = _16779_ & _16778_ /*1817*/;
  assign _16781_ = inv_31[66] & r_30[66] /*1816*/;
  assign _16782_ = _16780_ | _16781_ /*1815*/;
  assign _16783_ = inv_31[67] ^ r_30[67] /*1813*/;
  assign sum_31[67] = _16783_ ^ _16782_ /*1812*/;
  assign _16784_ = _16783_ & _16782_ /*1811*/;
  assign _16785_ = inv_31[67] & r_30[67] /*1810*/;
  assign _16786_ = _16784_ | _16785_ /*1809*/;
  assign _16787_ = inv_31[68] ^ r_30[68] /*1807*/;
  assign sum_31[68] = _16787_ ^ _16786_ /*1806*/;
  assign _16788_ = _16787_ & _16786_ /*1805*/;
  assign _16789_ = inv_31[68] & r_30[68] /*1804*/;
  assign _16790_ = _16788_ | _16789_ /*1803*/;
  assign _16791_ = inv_31[69] ^ r_30[69] /*1801*/;
  assign sum_31[69] = _16791_ ^ _16790_ /*1800*/;
  assign _16792_ = _16791_ & _16790_ /*1799*/;
  assign _16793_ = inv_31[69] & r_30[69] /*1798*/;
  assign _16794_ = _16792_ | _16793_ /*1797*/;
  assign _16795_ = inv_31[70] ^ r_30[70] /*1795*/;
  assign sum_31[70] = _16795_ ^ _16794_ /*1794*/;
  assign _16796_ = _16795_ & _16794_ /*1793*/;
  assign _16797_ = inv_31[70] & r_30[70] /*1792*/;
  assign _16798_ = _16796_ | _16797_ /*1791*/;
  assign _16799_ = inv_31[71] ^ r_30[71] /*1789*/;
  assign sum_31[71] = _16799_ ^ _16798_ /*1788*/;
  assign _16800_ = _16799_ & _16798_ /*1787*/;
  assign _16801_ = inv_31[71] & r_30[71] /*1786*/;
  assign _16802_ = _16800_ | _16801_ /*1785*/;
  assign _16803_ = inv_31[72] ^ r_30[72] /*1783*/;
  assign sum_31[72] = _16803_ ^ _16802_ /*1782*/;
  assign _16804_ = _16803_ & _16802_ /*1781*/;
  assign _16805_ = inv_31[72] & r_30[72] /*1780*/;
  assign _16806_ = _16804_ | _16805_ /*1779*/;
  assign _16807_ = inv_31[73] ^ r_30[73] /*1777*/;
  assign sum_31[73] = _16807_ ^ _16806_ /*1776*/;
  assign _16808_ = _16807_ & _16806_ /*1775*/;
  assign _16809_ = inv_31[73] & r_30[73] /*1774*/;
  assign _16810_ = _16808_ | _16809_ /*1773*/;
  assign _16811_ = inv_31[74] ^ r_30[74] /*1771*/;
  assign sum_31[74] = _16811_ ^ _16810_ /*1770*/;
  assign _16812_ = _16811_ & _16810_ /*1769*/;
  assign _16813_ = inv_31[74] & r_30[74] /*1768*/;
  assign _16814_ = _16812_ | _16813_ /*1767*/;
  assign _16815_ = inv_31[75] ^ r_30[75] /*1765*/;
  assign sum_31[75] = _16815_ ^ _16814_ /*1764*/;
  assign _16816_ = _16815_ & _16814_ /*1763*/;
  assign _16817_ = inv_31[75] & r_30[75] /*1762*/;
  assign _16818_ = _16816_ | _16817_ /*1761*/;
  assign _16819_ = inv_31[76] ^ r_30[76] /*1759*/;
  assign sum_31[76] = _16819_ ^ _16818_ /*1758*/;
  assign _16820_ = _16819_ & _16818_ /*1757*/;
  assign _16821_ = inv_31[76] & r_30[76] /*1756*/;
  assign _16822_ = _16820_ | _16821_ /*1755*/;
  assign _16823_ = inv_31[77] ^ r_30[77] /*1753*/;
  assign sum_31[77] = _16823_ ^ _16822_ /*1752*/;
  assign _16824_ = _16823_ & _16822_ /*1751*/;
  assign _16825_ = inv_31[77] & r_30[77] /*1750*/;
  assign _16826_ = _16824_ | _16825_ /*1749*/;
  assign _16827_ = inv_31[78] ^ r_30[78] /*1747*/;
  assign sum_31[78] = _16827_ ^ _16826_ /*1746*/;
  assign _16828_ = _16827_ & _16826_ /*1745*/;
  assign _16829_ = inv_31[78] & r_30[78] /*1744*/;
  assign _16830_ = _16828_ | _16829_ /*1743*/;
  assign _16831_ = inv_31[79] ^ r_30[79] /*1741*/;
  assign sum_31[79] = _16831_ ^ _16830_ /*1740*/;
  assign _16832_ = _16831_ & _16830_ /*1739*/;
  assign _16833_ = inv_31[79] & r_30[79] /*1738*/;
  assign _16834_ = _16832_ | _16833_ /*1737*/;
  assign _16835_ = inv_31[80] ^ r_30[80] /*1735*/;
  assign sum_31[80] = _16835_ ^ _16834_ /*1734*/;
  assign _16836_ = _16835_ & _16834_ /*1733*/;
  assign _16837_ = inv_31[80] & r_30[80] /*1732*/;
  assign _16838_ = _16836_ | _16837_ /*1731*/;
  assign _16839_ = inv_31[81] ^ r_30[81] /*1729*/;
  assign sum_31[81] = _16839_ ^ _16838_ /*1728*/;
  assign _16840_ = _16839_ & _16838_ /*1727*/;
  assign _16841_ = inv_31[81] & r_30[81] /*1726*/;
  assign _16842_ = _16840_ | _16841_ /*1725*/;
  assign _16843_ = inv_31[82] ^ r_30[82] /*1723*/;
  assign sum_31[82] = _16843_ ^ _16842_ /*1722*/;
  assign _16844_ = _16843_ & _16842_ /*1721*/;
  assign _16845_ = inv_31[82] & r_30[82] /*1720*/;
  assign _16846_ = _16844_ | _16845_ /*1719*/;
  assign _16847_ = inv_31[83] ^ r_30[83] /*1717*/;
  assign sum_31[83] = _16847_ ^ _16846_ /*1716*/;
  assign _16848_ = _16847_ & _16846_ /*1715*/;
  assign _16849_ = inv_31[83] & r_30[83] /*1714*/;
  assign _16850_ = _16848_ | _16849_ /*1713*/;
  assign _16851_ = inv_31[84] ^ r_30[84] /*1711*/;
  assign sum_31[84] = _16851_ ^ _16850_ /*1710*/;
  assign _16852_ = _16851_ & _16850_ /*1709*/;
  assign _16853_ = inv_31[84] & r_30[84] /*1708*/;
  assign _16854_ = _16852_ | _16853_ /*1707*/;
  assign _16855_ = inv_31[85] ^ r_30[85] /*1705*/;
  assign sum_31[85] = _16855_ ^ _16854_ /*1704*/;
  assign _16856_ = _16855_ & _16854_ /*1703*/;
  assign _16857_ = inv_31[85] & r_30[85] /*1702*/;
  assign _16858_ = _16856_ | _16857_ /*1701*/;
  assign _16859_ = inv_31[86] ^ r_30[86] /*1699*/;
  assign sum_31[86] = _16859_ ^ _16858_ /*1698*/;
  assign _16860_ = _16859_ & _16858_ /*1697*/;
  assign _16861_ = inv_31[86] & r_30[86] /*1696*/;
  assign _16862_ = _16860_ | _16861_ /*1695*/;
  assign _16863_ = inv_31[87] ^ r_30[87] /*1693*/;
  assign sum_31[87] = _16863_ ^ _16862_ /*1692*/;
  assign _16864_ = _16863_ & _16862_ /*1691*/;
  assign _16865_ = inv_31[87] & r_30[87] /*1690*/;
  assign _16866_ = _16864_ | _16865_ /*1689*/;
  assign _16867_ = inv_31[88] ^ r_30[88] /*1687*/;
  assign sum_31[88] = _16867_ ^ _16866_ /*1686*/;
  assign _16868_ = _16867_ & _16866_ /*1685*/;
  assign _16869_ = inv_31[88] & r_30[88] /*1684*/;
  assign _16870_ = _16868_ | _16869_ /*1683*/;
  assign _16871_ = inv_31[89] ^ r_30[89] /*1681*/;
  assign sum_31[89] = _16871_ ^ _16870_ /*1680*/;
  assign _16872_ = _16871_ & _16870_ /*1679*/;
  assign _16873_ = inv_31[89] & r_30[89] /*1678*/;
  assign _16874_ = _16872_ | _16873_ /*1677*/;
  assign _16875_ = inv_31[90] ^ r_30[90] /*1675*/;
  assign sum_31[90] = _16875_ ^ _16874_ /*1674*/;
  assign _16876_ = _16875_ & _16874_ /*1673*/;
  assign _16877_ = inv_31[90] & r_30[90] /*1672*/;
  assign _16878_ = _16876_ | _16877_ /*1671*/;
  assign _16879_ = inv_31[91] ^ r_30[91] /*1669*/;
  assign sum_31[91] = _16879_ ^ _16878_ /*1668*/;
  assign _16880_ = _16879_ & _16878_ /*1667*/;
  assign _16881_ = inv_31[91] & r_30[91] /*1666*/;
  assign _16882_ = _16880_ | _16881_ /*1665*/;
  assign _16883_ = inv_31[92] ^ r_30[92] /*1663*/;
  assign sum_31[92] = _16883_ ^ _16882_ /*1662*/;
  assign _16884_ = _16883_ & _16882_ /*1661*/;
  assign _16885_ = inv_31[92] & r_30[92] /*1660*/;
  assign _16886_ = _16884_ | _16885_ /*1659*/;
  assign _16887_ = _16886_ ^ _16882_ /*1658*/;
  assign _16888_ = ~_16887_ /*1657*/;
  assign _16889_ = sum_31[92] & _16888_ /*1656*/;
  assign _16890_ = _16887_ & _16886_ /*1655*/;
  assign sum_31[93] = _16890_ | _16889_ /*1654*/;
  assign q[1] = ~sum_31[93] /*1653*/;
  assign m_31[0] = r_30[0] /*1652*/;
  assign m_31[1] = r_30[1] /*1651*/;
  assign m_31[2] = r_30[2] /*1650*/;
  assign m_31[3] = r_30[3] /*1649*/;
  assign m_31[4] = r_30[4] /*1648*/;
  assign m_31[5] = r_30[5] /*1647*/;
  assign m_31[6] = r_30[6] /*1646*/;
  assign m_31[7] = r_30[7] /*1645*/;
  assign m_31[8] = r_30[8] /*1644*/;
  assign m_31[9] = r_30[9] /*1643*/;
  assign m_31[10] = r_30[10] /*1642*/;
  assign m_31[11] = r_30[11] /*1641*/;
  assign m_31[12] = r_30[12] /*1640*/;
  assign m_31[13] = r_30[13] /*1639*/;
  assign m_31[14] = r_30[14] /*1638*/;
  assign m_31[15] = r_30[15] /*1637*/;
  assign m_31[16] = r_30[16] /*1636*/;
  assign m_31[17] = r_30[17] /*1635*/;
  assign m_31[18] = r_30[18] /*1634*/;
  assign m_31[19] = r_30[19] /*1633*/;
  assign m_31[20] = r_30[20] /*1632*/;
  assign m_31[21] = r_30[21] /*1631*/;
  assign m_31[22] = r_30[22] /*1630*/;
  assign m_31[23] = r_30[23] /*1629*/;
  assign m_31[24] = r_30[24] /*1628*/;
  assign m_31[25] = r_30[25] /*1627*/;
  assign m_31[26] = r_30[26] /*1626*/;
  assign m_31[27] = r_30[27] /*1625*/;
  assign m_31[28] = r_30[28] /*1624*/;
  assign m_31[29] = r_30[29] /*1623*/;
  assign m_31[30] = r_30[30] /*1622*/;
  assign m_31[31] = r_30[31] /*1621*/;
  assign m_31[32] = r_30[32] /*1620*/;
  assign m_31[33] = r_30[33] /*1619*/;
  assign m_31[34] = r_30[34] /*1618*/;
  assign m_31[35] = r_30[35] /*1617*/;
  assign m_31[36] = r_30[36] /*1616*/;
  assign m_31[37] = r_30[37] /*1615*/;
  assign m_31[38] = r_30[38] /*1614*/;
  assign m_31[39] = r_30[39] /*1613*/;
  assign m_31[40] = r_30[40] /*1612*/;
  assign m_31[41] = r_30[41] /*1611*/;
  assign m_31[42] = r_30[42] /*1610*/;
  assign m_31[43] = r_30[43] /*1609*/;
  assign m_31[44] = r_30[44] /*1608*/;
  assign m_31[45] = r_30[45] /*1607*/;
  assign m_31[46] = r_30[46] /*1606*/;
  assign m_31[47] = r_30[47] /*1605*/;
  assign m_31[48] = r_30[48] /*1604*/;
  assign m_31[49] = r_30[49] /*1603*/;
  assign m_31[50] = r_30[50] /*1602*/;
  assign m_31[51] = r_30[51] /*1601*/;
  assign m_31[52] = r_30[52] /*1600*/;
  assign m_31[53] = r_30[53] /*1599*/;
  assign m_31[54] = r_30[54] /*1598*/;
  assign m_31[55] = r_30[55] /*1597*/;
  assign m_31[56] = r_30[56] /*1596*/;
  assign m_31[57] = r_30[57] /*1595*/;
  assign m_31[58] = r_30[58] /*1594*/;
  assign m_31[59] = r_30[59] /*1593*/;
  assign m_31[60] = r_30[60] /*1592*/;
  assign m_31[61] = r_30[61] /*1591*/;
  assign m_31[62] = r_30[62] /*1590*/;
  assign m_31[63] = r_30[63] /*1589*/;
  assign m_31[64] = r_30[64] /*1588*/;
  assign m_31[65] = r_30[65] /*1587*/;
  assign m_31[66] = r_30[66] /*1586*/;
  assign m_31[67] = r_30[67] /*1585*/;
  assign m_31[68] = r_30[68] /*1584*/;
  assign m_31[69] = r_30[69] /*1583*/;
  assign m_31[70] = r_30[70] /*1582*/;
  assign m_31[71] = r_30[71] /*1581*/;
  assign m_31[72] = r_30[72] /*1580*/;
  assign m_31[73] = r_30[73] /*1579*/;
  assign m_31[74] = r_30[74] /*1578*/;
  assign m_31[75] = r_30[75] /*1577*/;
  assign m_31[76] = r_30[76] /*1576*/;
  assign m_31[77] = r_30[77] /*1575*/;
  assign m_31[78] = r_30[78] /*1574*/;
  assign m_31[79] = r_30[79] /*1573*/;
  assign m_31[80] = r_30[80] /*1572*/;
  assign m_31[81] = r_30[81] /*1571*/;
  assign m_31[82] = r_30[82] /*1570*/;
  assign m_31[83] = r_30[83] /*1569*/;
  assign m_31[84] = r_30[84] /*1568*/;
  assign m_31[85] = r_30[85] /*1567*/;
  assign m_31[86] = r_30[86] /*1566*/;
  assign m_31[87] = r_30[87] /*1565*/;
  assign m_31[88] = r_30[88] /*1564*/;
  assign m_31[89] = r_30[89] /*1563*/;
  assign m_31[90] = r_30[90] /*1562*/;
  assign m_31[91] = r_30[91] /*1561*/;
  assign m_31[92] = r_30[92] /*1560*/;
  assign m_31[93] = r_30[92] /*1559*/;
  assign _16892_ = ~q[1] /*1558*/;
  assign _16893_ = sum_31[0] & q[1] /*1557*/;
  assign _16894_ = m_31[0] & _16892_ /*1556*/;
  assign r_31[0] = _16894_ | _16893_ /*1555*/;
  assign _16895_ = ~q[1] /*1554*/;
  assign _16896_ = sum_31[1] & q[1] /*1553*/;
  assign _16897_ = m_31[1] & _16895_ /*1552*/;
  assign r_31[1] = _16897_ | _16896_ /*1551*/;
  assign _16898_ = ~q[1] /*1550*/;
  assign _16899_ = sum_31[2] & q[1] /*1549*/;
  assign _16900_ = m_31[2] & _16898_ /*1548*/;
  assign r_31[2] = _16900_ | _16899_ /*1547*/;
  assign _16901_ = ~q[1] /*1546*/;
  assign _16902_ = sum_31[3] & q[1] /*1545*/;
  assign _16903_ = m_31[3] & _16901_ /*1544*/;
  assign r_31[3] = _16903_ | _16902_ /*1543*/;
  assign _16904_ = ~q[1] /*1542*/;
  assign _16905_ = sum_31[4] & q[1] /*1541*/;
  assign _16906_ = m_31[4] & _16904_ /*1540*/;
  assign r_31[4] = _16906_ | _16905_ /*1539*/;
  assign _16907_ = ~q[1] /*1538*/;
  assign _16908_ = sum_31[5] & q[1] /*1537*/;
  assign _16909_ = m_31[5] & _16907_ /*1536*/;
  assign r_31[5] = _16909_ | _16908_ /*1535*/;
  assign _16910_ = ~q[1] /*1534*/;
  assign _16911_ = sum_31[6] & q[1] /*1533*/;
  assign _16912_ = m_31[6] & _16910_ /*1532*/;
  assign r_31[6] = _16912_ | _16911_ /*1531*/;
  assign _16913_ = ~q[1] /*1530*/;
  assign _16914_ = sum_31[7] & q[1] /*1529*/;
  assign _16915_ = m_31[7] & _16913_ /*1528*/;
  assign r_31[7] = _16915_ | _16914_ /*1527*/;
  assign _16916_ = ~q[1] /*1526*/;
  assign _16917_ = sum_31[8] & q[1] /*1525*/;
  assign _16918_ = m_31[8] & _16916_ /*1524*/;
  assign r_31[8] = _16918_ | _16917_ /*1523*/;
  assign _16919_ = ~q[1] /*1522*/;
  assign _16920_ = sum_31[9] & q[1] /*1521*/;
  assign _16921_ = m_31[9] & _16919_ /*1520*/;
  assign r_31[9] = _16921_ | _16920_ /*1519*/;
  assign _16922_ = ~q[1] /*1518*/;
  assign _16923_ = sum_31[10] & q[1] /*1517*/;
  assign _16924_ = m_31[10] & _16922_ /*1516*/;
  assign r_31[10] = _16924_ | _16923_ /*1515*/;
  assign _16925_ = ~q[1] /*1514*/;
  assign _16926_ = sum_31[11] & q[1] /*1513*/;
  assign _16927_ = m_31[11] & _16925_ /*1512*/;
  assign r_31[11] = _16927_ | _16926_ /*1511*/;
  assign _16928_ = ~q[1] /*1510*/;
  assign _16929_ = sum_31[12] & q[1] /*1509*/;
  assign _16930_ = m_31[12] & _16928_ /*1508*/;
  assign r_31[12] = _16930_ | _16929_ /*1507*/;
  assign _16931_ = ~q[1] /*1506*/;
  assign _16932_ = sum_31[13] & q[1] /*1505*/;
  assign _16933_ = m_31[13] & _16931_ /*1504*/;
  assign r_31[13] = _16933_ | _16932_ /*1503*/;
  assign _16934_ = ~q[1] /*1502*/;
  assign _16935_ = sum_31[14] & q[1] /*1501*/;
  assign _16936_ = m_31[14] & _16934_ /*1500*/;
  assign r_31[14] = _16936_ | _16935_ /*1499*/;
  assign _16937_ = ~q[1] /*1498*/;
  assign _16938_ = sum_31[15] & q[1] /*1497*/;
  assign _16939_ = m_31[15] & _16937_ /*1496*/;
  assign r_31[15] = _16939_ | _16938_ /*1495*/;
  assign _16940_ = ~q[1] /*1494*/;
  assign _16941_ = sum_31[16] & q[1] /*1493*/;
  assign _16942_ = m_31[16] & _16940_ /*1492*/;
  assign r_31[16] = _16942_ | _16941_ /*1491*/;
  assign _16943_ = ~q[1] /*1490*/;
  assign _16944_ = sum_31[17] & q[1] /*1489*/;
  assign _16945_ = m_31[17] & _16943_ /*1488*/;
  assign r_31[17] = _16945_ | _16944_ /*1487*/;
  assign _16946_ = ~q[1] /*1486*/;
  assign _16947_ = sum_31[18] & q[1] /*1485*/;
  assign _16948_ = m_31[18] & _16946_ /*1484*/;
  assign r_31[18] = _16948_ | _16947_ /*1483*/;
  assign _16949_ = ~q[1] /*1482*/;
  assign _16950_ = sum_31[19] & q[1] /*1481*/;
  assign _16951_ = m_31[19] & _16949_ /*1480*/;
  assign r_31[19] = _16951_ | _16950_ /*1479*/;
  assign _16952_ = ~q[1] /*1478*/;
  assign _16953_ = sum_31[20] & q[1] /*1477*/;
  assign _16954_ = m_31[20] & _16952_ /*1476*/;
  assign r_31[20] = _16954_ | _16953_ /*1475*/;
  assign _16955_ = ~q[1] /*1474*/;
  assign _16956_ = sum_31[21] & q[1] /*1473*/;
  assign _16957_ = m_31[21] & _16955_ /*1472*/;
  assign r_31[21] = _16957_ | _16956_ /*1471*/;
  assign _16958_ = ~q[1] /*1470*/;
  assign _16959_ = sum_31[22] & q[1] /*1469*/;
  assign _16960_ = m_31[22] & _16958_ /*1468*/;
  assign r_31[22] = _16960_ | _16959_ /*1467*/;
  assign _16961_ = ~q[1] /*1466*/;
  assign _16962_ = sum_31[23] & q[1] /*1465*/;
  assign _16963_ = m_31[23] & _16961_ /*1464*/;
  assign r_31[23] = _16963_ | _16962_ /*1463*/;
  assign _16964_ = ~q[1] /*1462*/;
  assign _16965_ = sum_31[24] & q[1] /*1461*/;
  assign _16966_ = m_31[24] & _16964_ /*1460*/;
  assign r_31[24] = _16966_ | _16965_ /*1459*/;
  assign _16967_ = ~q[1] /*1458*/;
  assign _16968_ = sum_31[25] & q[1] /*1457*/;
  assign _16969_ = m_31[25] & _16967_ /*1456*/;
  assign r_31[25] = _16969_ | _16968_ /*1455*/;
  assign _16970_ = ~q[1] /*1454*/;
  assign _16971_ = sum_31[26] & q[1] /*1453*/;
  assign _16972_ = m_31[26] & _16970_ /*1452*/;
  assign r_31[26] = _16972_ | _16971_ /*1451*/;
  assign _16973_ = ~q[1] /*1450*/;
  assign _16974_ = sum_31[27] & q[1] /*1449*/;
  assign _16975_ = m_31[27] & _16973_ /*1448*/;
  assign r_31[27] = _16975_ | _16974_ /*1447*/;
  assign _16976_ = ~q[1] /*1446*/;
  assign _16977_ = sum_31[28] & q[1] /*1445*/;
  assign _16978_ = m_31[28] & _16976_ /*1444*/;
  assign r_31[28] = _16978_ | _16977_ /*1443*/;
  assign _16979_ = ~q[1] /*1442*/;
  assign _16980_ = sum_31[29] & q[1] /*1441*/;
  assign _16981_ = m_31[29] & _16979_ /*1440*/;
  assign r_31[29] = _16981_ | _16980_ /*1439*/;
  assign _16982_ = ~q[1] /*1438*/;
  assign _16983_ = sum_31[30] & q[1] /*1437*/;
  assign _16984_ = m_31[30] & _16982_ /*1436*/;
  assign r_31[30] = _16984_ | _16983_ /*1435*/;
  assign _16985_ = ~q[1] /*1434*/;
  assign _16986_ = sum_31[31] & q[1] /*1433*/;
  assign _16987_ = m_31[31] & _16985_ /*1432*/;
  assign r_31[31] = _16987_ | _16986_ /*1431*/;
  assign _16988_ = ~q[1] /*1430*/;
  assign _16989_ = sum_31[32] & q[1] /*1429*/;
  assign _16990_ = m_31[32] & _16988_ /*1428*/;
  assign r_31[32] = _16990_ | _16989_ /*1427*/;
  assign _16991_ = ~q[1] /*1426*/;
  assign _16992_ = sum_31[33] & q[1] /*1425*/;
  assign _16993_ = m_31[33] & _16991_ /*1424*/;
  assign r_31[33] = _16993_ | _16992_ /*1423*/;
  assign _16994_ = ~q[1] /*1422*/;
  assign _16995_ = sum_31[34] & q[1] /*1421*/;
  assign _16996_ = m_31[34] & _16994_ /*1420*/;
  assign r_31[34] = _16996_ | _16995_ /*1419*/;
  assign _16997_ = ~q[1] /*1418*/;
  assign _16998_ = sum_31[35] & q[1] /*1417*/;
  assign _16999_ = m_31[35] & _16997_ /*1416*/;
  assign r_31[35] = _16999_ | _16998_ /*1415*/;
  assign _17000_ = ~q[1] /*1414*/;
  assign _17001_ = sum_31[36] & q[1] /*1413*/;
  assign _17002_ = m_31[36] & _17000_ /*1412*/;
  assign r_31[36] = _17002_ | _17001_ /*1411*/;
  assign _17003_ = ~q[1] /*1410*/;
  assign _17004_ = sum_31[37] & q[1] /*1409*/;
  assign _17005_ = m_31[37] & _17003_ /*1408*/;
  assign r_31[37] = _17005_ | _17004_ /*1407*/;
  assign _17006_ = ~q[1] /*1406*/;
  assign _17007_ = sum_31[38] & q[1] /*1405*/;
  assign _17008_ = m_31[38] & _17006_ /*1404*/;
  assign r_31[38] = _17008_ | _17007_ /*1403*/;
  assign _17009_ = ~q[1] /*1402*/;
  assign _17010_ = sum_31[39] & q[1] /*1401*/;
  assign _17011_ = m_31[39] & _17009_ /*1400*/;
  assign r_31[39] = _17011_ | _17010_ /*1399*/;
  assign _17012_ = ~q[1] /*1398*/;
  assign _17013_ = sum_31[40] & q[1] /*1397*/;
  assign _17014_ = m_31[40] & _17012_ /*1396*/;
  assign r_31[40] = _17014_ | _17013_ /*1395*/;
  assign _17015_ = ~q[1] /*1394*/;
  assign _17016_ = sum_31[41] & q[1] /*1393*/;
  assign _17017_ = m_31[41] & _17015_ /*1392*/;
  assign r_31[41] = _17017_ | _17016_ /*1391*/;
  assign _17018_ = ~q[1] /*1390*/;
  assign _17019_ = sum_31[42] & q[1] /*1389*/;
  assign _17020_ = m_31[42] & _17018_ /*1388*/;
  assign r_31[42] = _17020_ | _17019_ /*1387*/;
  assign _17021_ = ~q[1] /*1386*/;
  assign _17022_ = sum_31[43] & q[1] /*1385*/;
  assign _17023_ = m_31[43] & _17021_ /*1384*/;
  assign r_31[43] = _17023_ | _17022_ /*1383*/;
  assign _17024_ = ~q[1] /*1382*/;
  assign _17025_ = sum_31[44] & q[1] /*1381*/;
  assign _17026_ = m_31[44] & _17024_ /*1380*/;
  assign r_31[44] = _17026_ | _17025_ /*1379*/;
  assign _17027_ = ~q[1] /*1378*/;
  assign _17028_ = sum_31[45] & q[1] /*1377*/;
  assign _17029_ = m_31[45] & _17027_ /*1376*/;
  assign r_31[45] = _17029_ | _17028_ /*1375*/;
  assign _17030_ = ~q[1] /*1374*/;
  assign _17031_ = sum_31[46] & q[1] /*1373*/;
  assign _17032_ = m_31[46] & _17030_ /*1372*/;
  assign r_31[46] = _17032_ | _17031_ /*1371*/;
  assign _17033_ = ~q[1] /*1370*/;
  assign _17034_ = sum_31[47] & q[1] /*1369*/;
  assign _17035_ = m_31[47] & _17033_ /*1368*/;
  assign r_31[47] = _17035_ | _17034_ /*1367*/;
  assign _17036_ = ~q[1] /*1366*/;
  assign _17037_ = sum_31[48] & q[1] /*1365*/;
  assign _17038_ = m_31[48] & _17036_ /*1364*/;
  assign r_31[48] = _17038_ | _17037_ /*1363*/;
  assign _17039_ = ~q[1] /*1362*/;
  assign _17040_ = sum_31[49] & q[1] /*1361*/;
  assign _17041_ = m_31[49] & _17039_ /*1360*/;
  assign r_31[49] = _17041_ | _17040_ /*1359*/;
  assign _17042_ = ~q[1] /*1358*/;
  assign _17043_ = sum_31[50] & q[1] /*1357*/;
  assign _17044_ = m_31[50] & _17042_ /*1356*/;
  assign r_31[50] = _17044_ | _17043_ /*1355*/;
  assign _17045_ = ~q[1] /*1354*/;
  assign _17046_ = sum_31[51] & q[1] /*1353*/;
  assign _17047_ = m_31[51] & _17045_ /*1352*/;
  assign r_31[51] = _17047_ | _17046_ /*1351*/;
  assign _17048_ = ~q[1] /*1350*/;
  assign _17049_ = sum_31[52] & q[1] /*1349*/;
  assign _17050_ = m_31[52] & _17048_ /*1348*/;
  assign r_31[52] = _17050_ | _17049_ /*1347*/;
  assign _17051_ = ~q[1] /*1346*/;
  assign _17052_ = sum_31[53] & q[1] /*1345*/;
  assign _17053_ = m_31[53] & _17051_ /*1344*/;
  assign r_31[53] = _17053_ | _17052_ /*1343*/;
  assign _17054_ = ~q[1] /*1342*/;
  assign _17055_ = sum_31[54] & q[1] /*1341*/;
  assign _17056_ = m_31[54] & _17054_ /*1340*/;
  assign r_31[54] = _17056_ | _17055_ /*1339*/;
  assign _17057_ = ~q[1] /*1338*/;
  assign _17058_ = sum_31[55] & q[1] /*1337*/;
  assign _17059_ = m_31[55] & _17057_ /*1336*/;
  assign r_31[55] = _17059_ | _17058_ /*1335*/;
  assign _17060_ = ~q[1] /*1334*/;
  assign _17061_ = sum_31[56] & q[1] /*1333*/;
  assign _17062_ = m_31[56] & _17060_ /*1332*/;
  assign r_31[56] = _17062_ | _17061_ /*1331*/;
  assign _17063_ = ~q[1] /*1330*/;
  assign _17064_ = sum_31[57] & q[1] /*1329*/;
  assign _17065_ = m_31[57] & _17063_ /*1328*/;
  assign r_31[57] = _17065_ | _17064_ /*1327*/;
  assign _17066_ = ~q[1] /*1326*/;
  assign _17067_ = sum_31[58] & q[1] /*1325*/;
  assign _17068_ = m_31[58] & _17066_ /*1324*/;
  assign r_31[58] = _17068_ | _17067_ /*1323*/;
  assign _17069_ = ~q[1] /*1322*/;
  assign _17070_ = sum_31[59] & q[1] /*1321*/;
  assign _17071_ = m_31[59] & _17069_ /*1320*/;
  assign r_31[59] = _17071_ | _17070_ /*1319*/;
  assign _17072_ = ~q[1] /*1318*/;
  assign _17073_ = sum_31[60] & q[1] /*1317*/;
  assign _17074_ = m_31[60] & _17072_ /*1316*/;
  assign r_31[60] = _17074_ | _17073_ /*1315*/;
  assign _17075_ = ~q[1] /*1314*/;
  assign _17076_ = sum_31[61] & q[1] /*1313*/;
  assign _17077_ = m_31[61] & _17075_ /*1312*/;
  assign r_31[61] = _17077_ | _17076_ /*1311*/;
  assign _17078_ = ~q[1] /*1310*/;
  assign _17079_ = sum_31[62] & q[1] /*1309*/;
  assign _17080_ = m_31[62] & _17078_ /*1308*/;
  assign r_31[62] = _17080_ | _17079_ /*1307*/;
  assign _17081_ = ~q[1] /*1306*/;
  assign _17082_ = sum_31[63] & q[1] /*1305*/;
  assign _17083_ = m_31[63] & _17081_ /*1304*/;
  assign r_31[63] = _17083_ | _17082_ /*1303*/;
  assign _17084_ = ~q[1] /*1302*/;
  assign _17085_ = sum_31[64] & q[1] /*1301*/;
  assign _17086_ = m_31[64] & _17084_ /*1300*/;
  assign r_31[64] = _17086_ | _17085_ /*1299*/;
  assign _17087_ = ~q[1] /*1298*/;
  assign _17088_ = sum_31[65] & q[1] /*1297*/;
  assign _17089_ = m_31[65] & _17087_ /*1296*/;
  assign r_31[65] = _17089_ | _17088_ /*1295*/;
  assign _17090_ = ~q[1] /*1294*/;
  assign _17091_ = sum_31[66] & q[1] /*1293*/;
  assign _17092_ = m_31[66] & _17090_ /*1292*/;
  assign r_31[66] = _17092_ | _17091_ /*1291*/;
  assign _17093_ = ~q[1] /*1290*/;
  assign _17094_ = sum_31[67] & q[1] /*1289*/;
  assign _17095_ = m_31[67] & _17093_ /*1288*/;
  assign r_31[67] = _17095_ | _17094_ /*1287*/;
  assign _17096_ = ~q[1] /*1286*/;
  assign _17097_ = sum_31[68] & q[1] /*1285*/;
  assign _17098_ = m_31[68] & _17096_ /*1284*/;
  assign r_31[68] = _17098_ | _17097_ /*1283*/;
  assign _17099_ = ~q[1] /*1282*/;
  assign _17100_ = sum_31[69] & q[1] /*1281*/;
  assign _17101_ = m_31[69] & _17099_ /*1280*/;
  assign r_31[69] = _17101_ | _17100_ /*1279*/;
  assign _17102_ = ~q[1] /*1278*/;
  assign _17103_ = sum_31[70] & q[1] /*1277*/;
  assign _17104_ = m_31[70] & _17102_ /*1276*/;
  assign r_31[70] = _17104_ | _17103_ /*1275*/;
  assign _17105_ = ~q[1] /*1274*/;
  assign _17106_ = sum_31[71] & q[1] /*1273*/;
  assign _17107_ = m_31[71] & _17105_ /*1272*/;
  assign r_31[71] = _17107_ | _17106_ /*1271*/;
  assign _17108_ = ~q[1] /*1270*/;
  assign _17109_ = sum_31[72] & q[1] /*1269*/;
  assign _17110_ = m_31[72] & _17108_ /*1268*/;
  assign r_31[72] = _17110_ | _17109_ /*1267*/;
  assign _17111_ = ~q[1] /*1266*/;
  assign _17112_ = sum_31[73] & q[1] /*1265*/;
  assign _17113_ = m_31[73] & _17111_ /*1264*/;
  assign r_31[73] = _17113_ | _17112_ /*1263*/;
  assign _17114_ = ~q[1] /*1262*/;
  assign _17115_ = sum_31[74] & q[1] /*1261*/;
  assign _17116_ = m_31[74] & _17114_ /*1260*/;
  assign r_31[74] = _17116_ | _17115_ /*1259*/;
  assign _17117_ = ~q[1] /*1258*/;
  assign _17118_ = sum_31[75] & q[1] /*1257*/;
  assign _17119_ = m_31[75] & _17117_ /*1256*/;
  assign r_31[75] = _17119_ | _17118_ /*1255*/;
  assign _17120_ = ~q[1] /*1254*/;
  assign _17121_ = sum_31[76] & q[1] /*1253*/;
  assign _17122_ = m_31[76] & _17120_ /*1252*/;
  assign r_31[76] = _17122_ | _17121_ /*1251*/;
  assign _17123_ = ~q[1] /*1250*/;
  assign _17124_ = sum_31[77] & q[1] /*1249*/;
  assign _17125_ = m_31[77] & _17123_ /*1248*/;
  assign r_31[77] = _17125_ | _17124_ /*1247*/;
  assign _17126_ = ~q[1] /*1246*/;
  assign _17127_ = sum_31[78] & q[1] /*1245*/;
  assign _17128_ = m_31[78] & _17126_ /*1244*/;
  assign r_31[78] = _17128_ | _17127_ /*1243*/;
  assign _17129_ = ~q[1] /*1242*/;
  assign _17130_ = sum_31[79] & q[1] /*1241*/;
  assign _17131_ = m_31[79] & _17129_ /*1240*/;
  assign r_31[79] = _17131_ | _17130_ /*1239*/;
  assign _17132_ = ~q[1] /*1238*/;
  assign _17133_ = sum_31[80] & q[1] /*1237*/;
  assign _17134_ = m_31[80] & _17132_ /*1236*/;
  assign r_31[80] = _17134_ | _17133_ /*1235*/;
  assign _17135_ = ~q[1] /*1234*/;
  assign _17136_ = sum_31[81] & q[1] /*1233*/;
  assign _17137_ = m_31[81] & _17135_ /*1232*/;
  assign r_31[81] = _17137_ | _17136_ /*1231*/;
  assign _17138_ = ~q[1] /*1230*/;
  assign _17139_ = sum_31[82] & q[1] /*1229*/;
  assign _17140_ = m_31[82] & _17138_ /*1228*/;
  assign r_31[82] = _17140_ | _17139_ /*1227*/;
  assign _17141_ = ~q[1] /*1226*/;
  assign _17142_ = sum_31[83] & q[1] /*1225*/;
  assign _17143_ = m_31[83] & _17141_ /*1224*/;
  assign r_31[83] = _17143_ | _17142_ /*1223*/;
  assign _17144_ = ~q[1] /*1222*/;
  assign _17145_ = sum_31[84] & q[1] /*1221*/;
  assign _17146_ = m_31[84] & _17144_ /*1220*/;
  assign r_31[84] = _17146_ | _17145_ /*1219*/;
  assign _17147_ = ~q[1] /*1218*/;
  assign _17148_ = sum_31[85] & q[1] /*1217*/;
  assign _17149_ = m_31[85] & _17147_ /*1216*/;
  assign r_31[85] = _17149_ | _17148_ /*1215*/;
  assign _17150_ = ~q[1] /*1214*/;
  assign _17151_ = sum_31[86] & q[1] /*1213*/;
  assign _17152_ = m_31[86] & _17150_ /*1212*/;
  assign r_31[86] = _17152_ | _17151_ /*1211*/;
  assign _17153_ = ~q[1] /*1210*/;
  assign _17154_ = sum_31[87] & q[1] /*1209*/;
  assign _17155_ = m_31[87] & _17153_ /*1208*/;
  assign r_31[87] = _17155_ | _17154_ /*1207*/;
  assign _17156_ = ~q[1] /*1206*/;
  assign _17157_ = sum_31[88] & q[1] /*1205*/;
  assign _17158_ = m_31[88] & _17156_ /*1204*/;
  assign r_31[88] = _17158_ | _17157_ /*1203*/;
  assign _17159_ = ~q[1] /*1202*/;
  assign _17160_ = sum_31[89] & q[1] /*1201*/;
  assign _17161_ = m_31[89] & _17159_ /*1200*/;
  assign r_31[89] = _17161_ | _17160_ /*1199*/;
  assign _17162_ = ~q[1] /*1198*/;
  assign _17163_ = sum_31[90] & q[1] /*1197*/;
  assign _17164_ = m_31[90] & _17162_ /*1196*/;
  assign r_31[90] = _17164_ | _17163_ /*1195*/;
  assign _17165_ = ~q[1] /*1194*/;
  assign _17166_ = sum_31[91] & q[1] /*1193*/;
  assign _17167_ = m_31[91] & _17165_ /*1192*/;
  assign r_31[91] = _17167_ | _17166_ /*1191*/;
  assign _17168_ = ~q[1] /*1190*/;
  assign _17169_ = sum_31[92] & q[1] /*1189*/;
  assign _17170_ = m_31[92] & _17168_ /*1188*/;
  assign r_31[92] = _17170_ | _17169_ /*1187*/;
  assign _17171_ = ~q[1] /*1186*/;
  assign _17172_ = sum_31[93] & q[1] /*1185*/;
  assign _17173_ = m_31[93] & _17171_ /*1184*/;
  assign r_31[93] = _17173_ | _17172_ /*1183*/;
  assign inv_32[0] = ~div[0] /*1140*/;
  assign inv_32[1] = ~div[1] /*1134*/;
  assign inv_32[2] = ~div[2] /*1128*/;
  assign inv_32[3] = ~div[3] /*1122*/;
  assign inv_32[4] = ~div[4] /*1116*/;
  assign inv_32[5] = ~div[5] /*1110*/;
  assign inv_32[6] = ~div[6] /*1104*/;
  assign inv_32[7] = ~div[7] /*1098*/;
  assign inv_32[8] = ~div[8] /*1092*/;
  assign inv_32[9] = ~div[9] /*1086*/;
  assign inv_32[10] = ~div[10] /*1080*/;
  assign inv_32[11] = ~div[11] /*1074*/;
  assign inv_32[12] = ~div[12] /*1068*/;
  assign inv_32[13] = ~div[13] /*1062*/;
  assign inv_32[14] = ~div[14] /*1056*/;
  assign inv_32[15] = ~div[15] /*1050*/;
  assign inv_32[16] = ~div[16] /*1044*/;
  assign inv_32[17] = ~div[17] /*1038*/;
  assign inv_32[18] = ~div[18] /*1032*/;
  assign inv_32[19] = ~div[19] /*1026*/;
  assign inv_32[20] = ~div[20] /*1020*/;
  assign inv_32[21] = ~div[21] /*1014*/;
  assign inv_32[22] = ~div[22] /*1008*/;
  assign inv_32[23] = ~div[23] /*1002*/;
  assign inv_32[24] = ~div[24] /*996*/;
  assign inv_32[25] = ~div[25] /*990*/;
  assign inv_32[26] = ~div[26] /*984*/;
  assign inv_32[27] = ~div[27] /*978*/;
  assign inv_32[28] = ~div[28] /*972*/;
  assign inv_32[29] = ~div[29] /*966*/;
  assign inv_32[30] = ~div[30] /*960*/;
  assign inv_32[31] = oneWire /*954*/;
  assign inv_32[32] = oneWire /*948*/;
  assign inv_32[33] = oneWire /*942*/;
  assign inv_32[34] = oneWire /*936*/;
  assign inv_32[35] = oneWire /*930*/;
  assign inv_32[36] = oneWire /*924*/;
  assign inv_32[37] = oneWire /*918*/;
  assign inv_32[38] = oneWire /*912*/;
  assign inv_32[39] = oneWire /*906*/;
  assign inv_32[40] = oneWire /*900*/;
  assign inv_32[41] = oneWire /*894*/;
  assign inv_32[42] = oneWire /*888*/;
  assign inv_32[43] = oneWire /*882*/;
  assign inv_32[44] = oneWire /*876*/;
  assign inv_32[45] = oneWire /*870*/;
  assign inv_32[46] = oneWire /*864*/;
  assign inv_32[47] = oneWire /*858*/;
  assign inv_32[48] = oneWire /*852*/;
  assign inv_32[49] = oneWire /*846*/;
  assign inv_32[50] = oneWire /*840*/;
  assign inv_32[51] = oneWire /*834*/;
  assign inv_32[52] = oneWire /*828*/;
  assign inv_32[53] = oneWire /*822*/;
  assign inv_32[54] = oneWire /*816*/;
  assign inv_32[55] = oneWire /*810*/;
  assign inv_32[56] = oneWire /*804*/;
  assign inv_32[57] = oneWire /*798*/;
  assign inv_32[58] = oneWire /*792*/;
  assign inv_32[59] = oneWire /*786*/;
  assign inv_32[60] = oneWire /*780*/;
  assign inv_32[61] = oneWire /*774*/;
  assign inv_32[62] = oneWire /*768*/;
  assign inv_32[63] = oneWire /*762*/;
  assign inv_32[64] = oneWire /*756*/;
  assign inv_32[65] = oneWire /*750*/;
  assign inv_32[66] = oneWire /*744*/;
  assign inv_32[67] = oneWire /*738*/;
  assign inv_32[68] = oneWire /*732*/;
  assign inv_32[69] = oneWire /*726*/;
  assign inv_32[70] = oneWire /*720*/;
  assign inv_32[71] = oneWire /*714*/;
  assign inv_32[72] = oneWire /*708*/;
  assign inv_32[73] = oneWire /*702*/;
  assign inv_32[74] = oneWire /*696*/;
  assign inv_32[75] = oneWire /*690*/;
  assign inv_32[76] = oneWire /*684*/;
  assign inv_32[77] = oneWire /*678*/;
  assign inv_32[78] = oneWire /*672*/;
  assign inv_32[79] = oneWire /*666*/;
  assign inv_32[80] = oneWire /*660*/;
  assign inv_32[81] = oneWire /*654*/;
  assign inv_32[82] = oneWire /*648*/;
  assign inv_32[83] = oneWire /*642*/;
  assign inv_32[84] = oneWire /*636*/;
  assign inv_32[85] = oneWire /*630*/;
  assign inv_32[86] = oneWire /*624*/;
  assign inv_32[87] = oneWire /*618*/;
  assign inv_32[88] = oneWire /*612*/;
  assign inv_32[89] = oneWire /*606*/;
  assign inv_32[90] = oneWire /*600*/;
  assign inv_32[91] = oneWire /*594*/;
  assign inv_32[92] = oneWire /*588*/;
  assign inv_32[93] = oneWire /*582*/;
  assign _17174_ = inv_32[0] ^ r_31[0] /*1139*/;
  assign sum_32[0] = _17174_ ^ oneWire /*1138*/;
  assign _17175_ = _17174_ & oneWire /*1137*/;
  assign _17176_ = inv_32[0] & r_31[0] /*1136*/;
  assign _17177_ = _17175_ | _17176_ /*1135*/;
  assign _17178_ = inv_32[1] ^ r_31[1] /*1133*/;
  assign sum_32[1] = _17178_ ^ _17177_ /*1132*/;
  assign _17179_ = _17178_ & _17177_ /*1131*/;
  assign _17180_ = inv_32[1] & r_31[1] /*1130*/;
  assign _17181_ = _17179_ | _17180_ /*1129*/;
  assign _17182_ = inv_32[2] ^ r_31[2] /*1127*/;
  assign sum_32[2] = _17182_ ^ _17181_ /*1126*/;
  assign _17183_ = _17182_ & _17181_ /*1125*/;
  assign _17184_ = inv_32[2] & r_31[2] /*1124*/;
  assign _17185_ = _17183_ | _17184_ /*1123*/;
  assign _17186_ = inv_32[3] ^ r_31[3] /*1121*/;
  assign sum_32[3] = _17186_ ^ _17185_ /*1120*/;
  assign _17187_ = _17186_ & _17185_ /*1119*/;
  assign _17188_ = inv_32[3] & r_31[3] /*1118*/;
  assign _17189_ = _17187_ | _17188_ /*1117*/;
  assign _17190_ = inv_32[4] ^ r_31[4] /*1115*/;
  assign sum_32[4] = _17190_ ^ _17189_ /*1114*/;
  assign _17191_ = _17190_ & _17189_ /*1113*/;
  assign _17192_ = inv_32[4] & r_31[4] /*1112*/;
  assign _17193_ = _17191_ | _17192_ /*1111*/;
  assign _17194_ = inv_32[5] ^ r_31[5] /*1109*/;
  assign sum_32[5] = _17194_ ^ _17193_ /*1108*/;
  assign _17195_ = _17194_ & _17193_ /*1107*/;
  assign _17196_ = inv_32[5] & r_31[5] /*1106*/;
  assign _17197_ = _17195_ | _17196_ /*1105*/;
  assign _17198_ = inv_32[6] ^ r_31[6] /*1103*/;
  assign sum_32[6] = _17198_ ^ _17197_ /*1102*/;
  assign _17199_ = _17198_ & _17197_ /*1101*/;
  assign _17200_ = inv_32[6] & r_31[6] /*1100*/;
  assign _17201_ = _17199_ | _17200_ /*1099*/;
  assign _17202_ = inv_32[7] ^ r_31[7] /*1097*/;
  assign sum_32[7] = _17202_ ^ _17201_ /*1096*/;
  assign _17203_ = _17202_ & _17201_ /*1095*/;
  assign _17204_ = inv_32[7] & r_31[7] /*1094*/;
  assign _17205_ = _17203_ | _17204_ /*1093*/;
  assign _17206_ = inv_32[8] ^ r_31[8] /*1091*/;
  assign sum_32[8] = _17206_ ^ _17205_ /*1090*/;
  assign _17207_ = _17206_ & _17205_ /*1089*/;
  assign _17208_ = inv_32[8] & r_31[8] /*1088*/;
  assign _17209_ = _17207_ | _17208_ /*1087*/;
  assign _17210_ = inv_32[9] ^ r_31[9] /*1085*/;
  assign sum_32[9] = _17210_ ^ _17209_ /*1084*/;
  assign _17211_ = _17210_ & _17209_ /*1083*/;
  assign _17212_ = inv_32[9] & r_31[9] /*1082*/;
  assign _17213_ = _17211_ | _17212_ /*1081*/;
  assign _17214_ = inv_32[10] ^ r_31[10] /*1079*/;
  assign sum_32[10] = _17214_ ^ _17213_ /*1078*/;
  assign _17215_ = _17214_ & _17213_ /*1077*/;
  assign _17216_ = inv_32[10] & r_31[10] /*1076*/;
  assign _17217_ = _17215_ | _17216_ /*1075*/;
  assign _17218_ = inv_32[11] ^ r_31[11] /*1073*/;
  assign sum_32[11] = _17218_ ^ _17217_ /*1072*/;
  assign _17219_ = _17218_ & _17217_ /*1071*/;
  assign _17220_ = inv_32[11] & r_31[11] /*1070*/;
  assign _17221_ = _17219_ | _17220_ /*1069*/;
  assign _17222_ = inv_32[12] ^ r_31[12] /*1067*/;
  assign sum_32[12] = _17222_ ^ _17221_ /*1066*/;
  assign _17223_ = _17222_ & _17221_ /*1065*/;
  assign _17224_ = inv_32[12] & r_31[12] /*1064*/;
  assign _17225_ = _17223_ | _17224_ /*1063*/;
  assign _17226_ = inv_32[13] ^ r_31[13] /*1061*/;
  assign sum_32[13] = _17226_ ^ _17225_ /*1060*/;
  assign _17227_ = _17226_ & _17225_ /*1059*/;
  assign _17228_ = inv_32[13] & r_31[13] /*1058*/;
  assign _17229_ = _17227_ | _17228_ /*1057*/;
  assign _17230_ = inv_32[14] ^ r_31[14] /*1055*/;
  assign sum_32[14] = _17230_ ^ _17229_ /*1054*/;
  assign _17231_ = _17230_ & _17229_ /*1053*/;
  assign _17232_ = inv_32[14] & r_31[14] /*1052*/;
  assign _17233_ = _17231_ | _17232_ /*1051*/;
  assign _17234_ = inv_32[15] ^ r_31[15] /*1049*/;
  assign sum_32[15] = _17234_ ^ _17233_ /*1048*/;
  assign _17235_ = _17234_ & _17233_ /*1047*/;
  assign _17236_ = inv_32[15] & r_31[15] /*1046*/;
  assign _17237_ = _17235_ | _17236_ /*1045*/;
  assign _17238_ = inv_32[16] ^ r_31[16] /*1043*/;
  assign sum_32[16] = _17238_ ^ _17237_ /*1042*/;
  assign _17239_ = _17238_ & _17237_ /*1041*/;
  assign _17240_ = inv_32[16] & r_31[16] /*1040*/;
  assign _17241_ = _17239_ | _17240_ /*1039*/;
  assign _17242_ = inv_32[17] ^ r_31[17] /*1037*/;
  assign sum_32[17] = _17242_ ^ _17241_ /*1036*/;
  assign _17243_ = _17242_ & _17241_ /*1035*/;
  assign _17244_ = inv_32[17] & r_31[17] /*1034*/;
  assign _17245_ = _17243_ | _17244_ /*1033*/;
  assign _17246_ = inv_32[18] ^ r_31[18] /*1031*/;
  assign sum_32[18] = _17246_ ^ _17245_ /*1030*/;
  assign _17247_ = _17246_ & _17245_ /*1029*/;
  assign _17248_ = inv_32[18] & r_31[18] /*1028*/;
  assign _17249_ = _17247_ | _17248_ /*1027*/;
  assign _17250_ = inv_32[19] ^ r_31[19] /*1025*/;
  assign sum_32[19] = _17250_ ^ _17249_ /*1024*/;
  assign _17251_ = _17250_ & _17249_ /*1023*/;
  assign _17252_ = inv_32[19] & r_31[19] /*1022*/;
  assign _17253_ = _17251_ | _17252_ /*1021*/;
  assign _17254_ = inv_32[20] ^ r_31[20] /*1019*/;
  assign sum_32[20] = _17254_ ^ _17253_ /*1018*/;
  assign _17255_ = _17254_ & _17253_ /*1017*/;
  assign _17256_ = inv_32[20] & r_31[20] /*1016*/;
  assign _17257_ = _17255_ | _17256_ /*1015*/;
  assign _17258_ = inv_32[21] ^ r_31[21] /*1013*/;
  assign sum_32[21] = _17258_ ^ _17257_ /*1012*/;
  assign _17259_ = _17258_ & _17257_ /*1011*/;
  assign _17260_ = inv_32[21] & r_31[21] /*1010*/;
  assign _17261_ = _17259_ | _17260_ /*1009*/;
  assign _17262_ = inv_32[22] ^ r_31[22] /*1007*/;
  assign sum_32[22] = _17262_ ^ _17261_ /*1006*/;
  assign _17263_ = _17262_ & _17261_ /*1005*/;
  assign _17264_ = inv_32[22] & r_31[22] /*1004*/;
  assign _17265_ = _17263_ | _17264_ /*1003*/;
  assign _17266_ = inv_32[23] ^ r_31[23] /*1001*/;
  assign sum_32[23] = _17266_ ^ _17265_ /*1000*/;
  assign _17267_ = _17266_ & _17265_ /*999*/;
  assign _17268_ = inv_32[23] & r_31[23] /*998*/;
  assign _17269_ = _17267_ | _17268_ /*997*/;
  assign _17270_ = inv_32[24] ^ r_31[24] /*995*/;
  assign sum_32[24] = _17270_ ^ _17269_ /*994*/;
  assign _17271_ = _17270_ & _17269_ /*993*/;
  assign _17272_ = inv_32[24] & r_31[24] /*992*/;
  assign _17273_ = _17271_ | _17272_ /*991*/;
  assign _17274_ = inv_32[25] ^ r_31[25] /*989*/;
  assign sum_32[25] = _17274_ ^ _17273_ /*988*/;
  assign _17275_ = _17274_ & _17273_ /*987*/;
  assign _17276_ = inv_32[25] & r_31[25] /*986*/;
  assign _17277_ = _17275_ | _17276_ /*985*/;
  assign _17278_ = inv_32[26] ^ r_31[26] /*983*/;
  assign sum_32[26] = _17278_ ^ _17277_ /*982*/;
  assign _17279_ = _17278_ & _17277_ /*981*/;
  assign _17280_ = inv_32[26] & r_31[26] /*980*/;
  assign _17281_ = _17279_ | _17280_ /*979*/;
  assign _17282_ = inv_32[27] ^ r_31[27] /*977*/;
  assign sum_32[27] = _17282_ ^ _17281_ /*976*/;
  assign _17283_ = _17282_ & _17281_ /*975*/;
  assign _17284_ = inv_32[27] & r_31[27] /*974*/;
  assign _17285_ = _17283_ | _17284_ /*973*/;
  assign _17286_ = inv_32[28] ^ r_31[28] /*971*/;
  assign sum_32[28] = _17286_ ^ _17285_ /*970*/;
  assign _17287_ = _17286_ & _17285_ /*969*/;
  assign _17288_ = inv_32[28] & r_31[28] /*968*/;
  assign _17289_ = _17287_ | _17288_ /*967*/;
  assign _17290_ = inv_32[29] ^ r_31[29] /*965*/;
  assign sum_32[29] = _17290_ ^ _17289_ /*964*/;
  assign _17291_ = _17290_ & _17289_ /*963*/;
  assign _17292_ = inv_32[29] & r_31[29] /*962*/;
  assign _17293_ = _17291_ | _17292_ /*961*/;
  assign _17294_ = inv_32[30] ^ r_31[30] /*959*/;
  assign sum_32[30] = _17294_ ^ _17293_ /*958*/;
  assign _17295_ = _17294_ & _17293_ /*957*/;
  assign _17296_ = inv_32[30] & r_31[30] /*956*/;
  assign _17297_ = _17295_ | _17296_ /*955*/;
  assign _17298_ = inv_32[31] ^ r_31[31] /*953*/;
  assign sum_32[31] = _17298_ ^ _17297_ /*952*/;
  assign _17299_ = _17298_ & _17297_ /*951*/;
  assign _17300_ = inv_32[31] & r_31[31] /*950*/;
  assign _17301_ = _17299_ | _17300_ /*949*/;
  assign _17302_ = inv_32[32] ^ r_31[32] /*947*/;
  assign sum_32[32] = _17302_ ^ _17301_ /*946*/;
  assign _17303_ = _17302_ & _17301_ /*945*/;
  assign _17304_ = inv_32[32] & r_31[32] /*944*/;
  assign _17305_ = _17303_ | _17304_ /*943*/;
  assign _17306_ = inv_32[33] ^ r_31[33] /*941*/;
  assign sum_32[33] = _17306_ ^ _17305_ /*940*/;
  assign _17307_ = _17306_ & _17305_ /*939*/;
  assign _17308_ = inv_32[33] & r_31[33] /*938*/;
  assign _17309_ = _17307_ | _17308_ /*937*/;
  assign _17310_ = inv_32[34] ^ r_31[34] /*935*/;
  assign sum_32[34] = _17310_ ^ _17309_ /*934*/;
  assign _17311_ = _17310_ & _17309_ /*933*/;
  assign _17312_ = inv_32[34] & r_31[34] /*932*/;
  assign _17313_ = _17311_ | _17312_ /*931*/;
  assign _17314_ = inv_32[35] ^ r_31[35] /*929*/;
  assign sum_32[35] = _17314_ ^ _17313_ /*928*/;
  assign _17315_ = _17314_ & _17313_ /*927*/;
  assign _17316_ = inv_32[35] & r_31[35] /*926*/;
  assign _17317_ = _17315_ | _17316_ /*925*/;
  assign _17318_ = inv_32[36] ^ r_31[36] /*923*/;
  assign sum_32[36] = _17318_ ^ _17317_ /*922*/;
  assign _17319_ = _17318_ & _17317_ /*921*/;
  assign _17320_ = inv_32[36] & r_31[36] /*920*/;
  assign _17321_ = _17319_ | _17320_ /*919*/;
  assign _17322_ = inv_32[37] ^ r_31[37] /*917*/;
  assign sum_32[37] = _17322_ ^ _17321_ /*916*/;
  assign _17323_ = _17322_ & _17321_ /*915*/;
  assign _17324_ = inv_32[37] & r_31[37] /*914*/;
  assign _17325_ = _17323_ | _17324_ /*913*/;
  assign _17326_ = inv_32[38] ^ r_31[38] /*911*/;
  assign sum_32[38] = _17326_ ^ _17325_ /*910*/;
  assign _17327_ = _17326_ & _17325_ /*909*/;
  assign _17328_ = inv_32[38] & r_31[38] /*908*/;
  assign _17329_ = _17327_ | _17328_ /*907*/;
  assign _17330_ = inv_32[39] ^ r_31[39] /*905*/;
  assign sum_32[39] = _17330_ ^ _17329_ /*904*/;
  assign _17331_ = _17330_ & _17329_ /*903*/;
  assign _17332_ = inv_32[39] & r_31[39] /*902*/;
  assign _17333_ = _17331_ | _17332_ /*901*/;
  assign _17334_ = inv_32[40] ^ r_31[40] /*899*/;
  assign sum_32[40] = _17334_ ^ _17333_ /*898*/;
  assign _17335_ = _17334_ & _17333_ /*897*/;
  assign _17336_ = inv_32[40] & r_31[40] /*896*/;
  assign _17337_ = _17335_ | _17336_ /*895*/;
  assign _17338_ = inv_32[41] ^ r_31[41] /*893*/;
  assign sum_32[41] = _17338_ ^ _17337_ /*892*/;
  assign _17339_ = _17338_ & _17337_ /*891*/;
  assign _17340_ = inv_32[41] & r_31[41] /*890*/;
  assign _17341_ = _17339_ | _17340_ /*889*/;
  assign _17342_ = inv_32[42] ^ r_31[42] /*887*/;
  assign sum_32[42] = _17342_ ^ _17341_ /*886*/;
  assign _17343_ = _17342_ & _17341_ /*885*/;
  assign _17344_ = inv_32[42] & r_31[42] /*884*/;
  assign _17345_ = _17343_ | _17344_ /*883*/;
  assign _17346_ = inv_32[43] ^ r_31[43] /*881*/;
  assign sum_32[43] = _17346_ ^ _17345_ /*880*/;
  assign _17347_ = _17346_ & _17345_ /*879*/;
  assign _17348_ = inv_32[43] & r_31[43] /*878*/;
  assign _17349_ = _17347_ | _17348_ /*877*/;
  assign _17350_ = inv_32[44] ^ r_31[44] /*875*/;
  assign sum_32[44] = _17350_ ^ _17349_ /*874*/;
  assign _17351_ = _17350_ & _17349_ /*873*/;
  assign _17352_ = inv_32[44] & r_31[44] /*872*/;
  assign _17353_ = _17351_ | _17352_ /*871*/;
  assign _17354_ = inv_32[45] ^ r_31[45] /*869*/;
  assign sum_32[45] = _17354_ ^ _17353_ /*868*/;
  assign _17355_ = _17354_ & _17353_ /*867*/;
  assign _17356_ = inv_32[45] & r_31[45] /*866*/;
  assign _17357_ = _17355_ | _17356_ /*865*/;
  assign _17358_ = inv_32[46] ^ r_31[46] /*863*/;
  assign sum_32[46] = _17358_ ^ _17357_ /*862*/;
  assign _17359_ = _17358_ & _17357_ /*861*/;
  assign _17360_ = inv_32[46] & r_31[46] /*860*/;
  assign _17361_ = _17359_ | _17360_ /*859*/;
  assign _17362_ = inv_32[47] ^ r_31[47] /*857*/;
  assign sum_32[47] = _17362_ ^ _17361_ /*856*/;
  assign _17363_ = _17362_ & _17361_ /*855*/;
  assign _17364_ = inv_32[47] & r_31[47] /*854*/;
  assign _17365_ = _17363_ | _17364_ /*853*/;
  assign _17366_ = inv_32[48] ^ r_31[48] /*851*/;
  assign sum_32[48] = _17366_ ^ _17365_ /*850*/;
  assign _17367_ = _17366_ & _17365_ /*849*/;
  assign _17368_ = inv_32[48] & r_31[48] /*848*/;
  assign _17369_ = _17367_ | _17368_ /*847*/;
  assign _17370_ = inv_32[49] ^ r_31[49] /*845*/;
  assign sum_32[49] = _17370_ ^ _17369_ /*844*/;
  assign _17371_ = _17370_ & _17369_ /*843*/;
  assign _17372_ = inv_32[49] & r_31[49] /*842*/;
  assign _17373_ = _17371_ | _17372_ /*841*/;
  assign _17374_ = inv_32[50] ^ r_31[50] /*839*/;
  assign sum_32[50] = _17374_ ^ _17373_ /*838*/;
  assign _17375_ = _17374_ & _17373_ /*837*/;
  assign _17376_ = inv_32[50] & r_31[50] /*836*/;
  assign _17377_ = _17375_ | _17376_ /*835*/;
  assign _17378_ = inv_32[51] ^ r_31[51] /*833*/;
  assign sum_32[51] = _17378_ ^ _17377_ /*832*/;
  assign _17379_ = _17378_ & _17377_ /*831*/;
  assign _17380_ = inv_32[51] & r_31[51] /*830*/;
  assign _17381_ = _17379_ | _17380_ /*829*/;
  assign _17382_ = inv_32[52] ^ r_31[52] /*827*/;
  assign sum_32[52] = _17382_ ^ _17381_ /*826*/;
  assign _17383_ = _17382_ & _17381_ /*825*/;
  assign _17384_ = inv_32[52] & r_31[52] /*824*/;
  assign _17385_ = _17383_ | _17384_ /*823*/;
  assign _17386_ = inv_32[53] ^ r_31[53] /*821*/;
  assign sum_32[53] = _17386_ ^ _17385_ /*820*/;
  assign _17387_ = _17386_ & _17385_ /*819*/;
  assign _17388_ = inv_32[53] & r_31[53] /*818*/;
  assign _17389_ = _17387_ | _17388_ /*817*/;
  assign _17390_ = inv_32[54] ^ r_31[54] /*815*/;
  assign sum_32[54] = _17390_ ^ _17389_ /*814*/;
  assign _17391_ = _17390_ & _17389_ /*813*/;
  assign _17392_ = inv_32[54] & r_31[54] /*812*/;
  assign _17393_ = _17391_ | _17392_ /*811*/;
  assign _17394_ = inv_32[55] ^ r_31[55] /*809*/;
  assign sum_32[55] = _17394_ ^ _17393_ /*808*/;
  assign _17395_ = _17394_ & _17393_ /*807*/;
  assign _17396_ = inv_32[55] & r_31[55] /*806*/;
  assign _17397_ = _17395_ | _17396_ /*805*/;
  assign _17398_ = inv_32[56] ^ r_31[56] /*803*/;
  assign sum_32[56] = _17398_ ^ _17397_ /*802*/;
  assign _17399_ = _17398_ & _17397_ /*801*/;
  assign _17400_ = inv_32[56] & r_31[56] /*800*/;
  assign _17401_ = _17399_ | _17400_ /*799*/;
  assign _17402_ = inv_32[57] ^ r_31[57] /*797*/;
  assign sum_32[57] = _17402_ ^ _17401_ /*796*/;
  assign _17403_ = _17402_ & _17401_ /*795*/;
  assign _17404_ = inv_32[57] & r_31[57] /*794*/;
  assign _17405_ = _17403_ | _17404_ /*793*/;
  assign _17406_ = inv_32[58] ^ r_31[58] /*791*/;
  assign sum_32[58] = _17406_ ^ _17405_ /*790*/;
  assign _17407_ = _17406_ & _17405_ /*789*/;
  assign _17408_ = inv_32[58] & r_31[58] /*788*/;
  assign _17409_ = _17407_ | _17408_ /*787*/;
  assign _17410_ = inv_32[59] ^ r_31[59] /*785*/;
  assign sum_32[59] = _17410_ ^ _17409_ /*784*/;
  assign _17411_ = _17410_ & _17409_ /*783*/;
  assign _17412_ = inv_32[59] & r_31[59] /*782*/;
  assign _17413_ = _17411_ | _17412_ /*781*/;
  assign _17414_ = inv_32[60] ^ r_31[60] /*779*/;
  assign sum_32[60] = _17414_ ^ _17413_ /*778*/;
  assign _17415_ = _17414_ & _17413_ /*777*/;
  assign _17416_ = inv_32[60] & r_31[60] /*776*/;
  assign _17417_ = _17415_ | _17416_ /*775*/;
  assign _17418_ = inv_32[61] ^ r_31[61] /*773*/;
  assign sum_32[61] = _17418_ ^ _17417_ /*772*/;
  assign _17419_ = _17418_ & _17417_ /*771*/;
  assign _17420_ = inv_32[61] & r_31[61] /*770*/;
  assign _17421_ = _17419_ | _17420_ /*769*/;
  assign _17422_ = inv_32[62] ^ r_31[62] /*767*/;
  assign sum_32[62] = _17422_ ^ _17421_ /*766*/;
  assign _17423_ = _17422_ & _17421_ /*765*/;
  assign _17424_ = inv_32[62] & r_31[62] /*764*/;
  assign _17425_ = _17423_ | _17424_ /*763*/;
  assign _17426_ = inv_32[63] ^ r_31[63] /*761*/;
  assign sum_32[63] = _17426_ ^ _17425_ /*760*/;
  assign _17427_ = _17426_ & _17425_ /*759*/;
  assign _17428_ = inv_32[63] & r_31[63] /*758*/;
  assign _17429_ = _17427_ | _17428_ /*757*/;
  assign _17430_ = inv_32[64] ^ r_31[64] /*755*/;
  assign sum_32[64] = _17430_ ^ _17429_ /*754*/;
  assign _17431_ = _17430_ & _17429_ /*753*/;
  assign _17432_ = inv_32[64] & r_31[64] /*752*/;
  assign _17433_ = _17431_ | _17432_ /*751*/;
  assign _17434_ = inv_32[65] ^ r_31[65] /*749*/;
  assign sum_32[65] = _17434_ ^ _17433_ /*748*/;
  assign _17435_ = _17434_ & _17433_ /*747*/;
  assign _17436_ = inv_32[65] & r_31[65] /*746*/;
  assign _17437_ = _17435_ | _17436_ /*745*/;
  assign _17438_ = inv_32[66] ^ r_31[66] /*743*/;
  assign sum_32[66] = _17438_ ^ _17437_ /*742*/;
  assign _17439_ = _17438_ & _17437_ /*741*/;
  assign _17440_ = inv_32[66] & r_31[66] /*740*/;
  assign _17441_ = _17439_ | _17440_ /*739*/;
  assign _17442_ = inv_32[67] ^ r_31[67] /*737*/;
  assign sum_32[67] = _17442_ ^ _17441_ /*736*/;
  assign _17443_ = _17442_ & _17441_ /*735*/;
  assign _17444_ = inv_32[67] & r_31[67] /*734*/;
  assign _17445_ = _17443_ | _17444_ /*733*/;
  assign _17446_ = inv_32[68] ^ r_31[68] /*731*/;
  assign sum_32[68] = _17446_ ^ _17445_ /*730*/;
  assign _17447_ = _17446_ & _17445_ /*729*/;
  assign _17448_ = inv_32[68] & r_31[68] /*728*/;
  assign _17449_ = _17447_ | _17448_ /*727*/;
  assign _17450_ = inv_32[69] ^ r_31[69] /*725*/;
  assign sum_32[69] = _17450_ ^ _17449_ /*724*/;
  assign _17451_ = _17450_ & _17449_ /*723*/;
  assign _17452_ = inv_32[69] & r_31[69] /*722*/;
  assign _17453_ = _17451_ | _17452_ /*721*/;
  assign _17454_ = inv_32[70] ^ r_31[70] /*719*/;
  assign sum_32[70] = _17454_ ^ _17453_ /*718*/;
  assign _17455_ = _17454_ & _17453_ /*717*/;
  assign _17456_ = inv_32[70] & r_31[70] /*716*/;
  assign _17457_ = _17455_ | _17456_ /*715*/;
  assign _17458_ = inv_32[71] ^ r_31[71] /*713*/;
  assign sum_32[71] = _17458_ ^ _17457_ /*712*/;
  assign _17459_ = _17458_ & _17457_ /*711*/;
  assign _17460_ = inv_32[71] & r_31[71] /*710*/;
  assign _17461_ = _17459_ | _17460_ /*709*/;
  assign _17462_ = inv_32[72] ^ r_31[72] /*707*/;
  assign sum_32[72] = _17462_ ^ _17461_ /*706*/;
  assign _17463_ = _17462_ & _17461_ /*705*/;
  assign _17464_ = inv_32[72] & r_31[72] /*704*/;
  assign _17465_ = _17463_ | _17464_ /*703*/;
  assign _17466_ = inv_32[73] ^ r_31[73] /*701*/;
  assign sum_32[73] = _17466_ ^ _17465_ /*700*/;
  assign _17467_ = _17466_ & _17465_ /*699*/;
  assign _17468_ = inv_32[73] & r_31[73] /*698*/;
  assign _17469_ = _17467_ | _17468_ /*697*/;
  assign _17470_ = inv_32[74] ^ r_31[74] /*695*/;
  assign sum_32[74] = _17470_ ^ _17469_ /*694*/;
  assign _17471_ = _17470_ & _17469_ /*693*/;
  assign _17472_ = inv_32[74] & r_31[74] /*692*/;
  assign _17473_ = _17471_ | _17472_ /*691*/;
  assign _17474_ = inv_32[75] ^ r_31[75] /*689*/;
  assign sum_32[75] = _17474_ ^ _17473_ /*688*/;
  assign _17475_ = _17474_ & _17473_ /*687*/;
  assign _17476_ = inv_32[75] & r_31[75] /*686*/;
  assign _17477_ = _17475_ | _17476_ /*685*/;
  assign _17478_ = inv_32[76] ^ r_31[76] /*683*/;
  assign sum_32[76] = _17478_ ^ _17477_ /*682*/;
  assign _17479_ = _17478_ & _17477_ /*681*/;
  assign _17480_ = inv_32[76] & r_31[76] /*680*/;
  assign _17481_ = _17479_ | _17480_ /*679*/;
  assign _17482_ = inv_32[77] ^ r_31[77] /*677*/;
  assign sum_32[77] = _17482_ ^ _17481_ /*676*/;
  assign _17483_ = _17482_ & _17481_ /*675*/;
  assign _17484_ = inv_32[77] & r_31[77] /*674*/;
  assign _17485_ = _17483_ | _17484_ /*673*/;
  assign _17486_ = inv_32[78] ^ r_31[78] /*671*/;
  assign sum_32[78] = _17486_ ^ _17485_ /*670*/;
  assign _17487_ = _17486_ & _17485_ /*669*/;
  assign _17488_ = inv_32[78] & r_31[78] /*668*/;
  assign _17489_ = _17487_ | _17488_ /*667*/;
  assign _17490_ = inv_32[79] ^ r_31[79] /*665*/;
  assign sum_32[79] = _17490_ ^ _17489_ /*664*/;
  assign _17491_ = _17490_ & _17489_ /*663*/;
  assign _17492_ = inv_32[79] & r_31[79] /*662*/;
  assign _17493_ = _17491_ | _17492_ /*661*/;
  assign _17494_ = inv_32[80] ^ r_31[80] /*659*/;
  assign sum_32[80] = _17494_ ^ _17493_ /*658*/;
  assign _17495_ = _17494_ & _17493_ /*657*/;
  assign _17496_ = inv_32[80] & r_31[80] /*656*/;
  assign _17497_ = _17495_ | _17496_ /*655*/;
  assign _17498_ = inv_32[81] ^ r_31[81] /*653*/;
  assign sum_32[81] = _17498_ ^ _17497_ /*652*/;
  assign _17499_ = _17498_ & _17497_ /*651*/;
  assign _17500_ = inv_32[81] & r_31[81] /*650*/;
  assign _17501_ = _17499_ | _17500_ /*649*/;
  assign _17502_ = inv_32[82] ^ r_31[82] /*647*/;
  assign sum_32[82] = _17502_ ^ _17501_ /*646*/;
  assign _17503_ = _17502_ & _17501_ /*645*/;
  assign _17504_ = inv_32[82] & r_31[82] /*644*/;
  assign _17505_ = _17503_ | _17504_ /*643*/;
  assign _17506_ = inv_32[83] ^ r_31[83] /*641*/;
  assign sum_32[83] = _17506_ ^ _17505_ /*640*/;
  assign _17507_ = _17506_ & _17505_ /*639*/;
  assign _17508_ = inv_32[83] & r_31[83] /*638*/;
  assign _17509_ = _17507_ | _17508_ /*637*/;
  assign _17510_ = inv_32[84] ^ r_31[84] /*635*/;
  assign sum_32[84] = _17510_ ^ _17509_ /*634*/;
  assign _17511_ = _17510_ & _17509_ /*633*/;
  assign _17512_ = inv_32[84] & r_31[84] /*632*/;
  assign _17513_ = _17511_ | _17512_ /*631*/;
  assign _17514_ = inv_32[85] ^ r_31[85] /*629*/;
  assign sum_32[85] = _17514_ ^ _17513_ /*628*/;
  assign _17515_ = _17514_ & _17513_ /*627*/;
  assign _17516_ = inv_32[85] & r_31[85] /*626*/;
  assign _17517_ = _17515_ | _17516_ /*625*/;
  assign _17518_ = inv_32[86] ^ r_31[86] /*623*/;
  assign sum_32[86] = _17518_ ^ _17517_ /*622*/;
  assign _17519_ = _17518_ & _17517_ /*621*/;
  assign _17520_ = inv_32[86] & r_31[86] /*620*/;
  assign _17521_ = _17519_ | _17520_ /*619*/;
  assign _17522_ = inv_32[87] ^ r_31[87] /*617*/;
  assign sum_32[87] = _17522_ ^ _17521_ /*616*/;
  assign _17523_ = _17522_ & _17521_ /*615*/;
  assign _17524_ = inv_32[87] & r_31[87] /*614*/;
  assign _17525_ = _17523_ | _17524_ /*613*/;
  assign _17526_ = inv_32[88] ^ r_31[88] /*611*/;
  assign sum_32[88] = _17526_ ^ _17525_ /*610*/;
  assign _17527_ = _17526_ & _17525_ /*609*/;
  assign _17528_ = inv_32[88] & r_31[88] /*608*/;
  assign _17529_ = _17527_ | _17528_ /*607*/;
  assign _17530_ = inv_32[89] ^ r_31[89] /*605*/;
  assign sum_32[89] = _17530_ ^ _17529_ /*604*/;
  assign _17531_ = _17530_ & _17529_ /*603*/;
  assign _17532_ = inv_32[89] & r_31[89] /*602*/;
  assign _17533_ = _17531_ | _17532_ /*601*/;
  assign _17534_ = inv_32[90] ^ r_31[90] /*599*/;
  assign sum_32[90] = _17534_ ^ _17533_ /*598*/;
  assign _17535_ = _17534_ & _17533_ /*597*/;
  assign _17536_ = inv_32[90] & r_31[90] /*596*/;
  assign _17537_ = _17535_ | _17536_ /*595*/;
  assign _17538_ = inv_32[91] ^ r_31[91] /*593*/;
  assign sum_32[91] = _17538_ ^ _17537_ /*592*/;
  assign _17539_ = _17538_ & _17537_ /*591*/;
  assign _17540_ = inv_32[91] & r_31[91] /*590*/;
  assign _17541_ = _17539_ | _17540_ /*589*/;
  assign _17542_ = inv_32[92] ^ r_31[92] /*587*/;
  assign sum_32[92] = _17542_ ^ _17541_ /*586*/;
  assign _17543_ = _17542_ & _17541_ /*585*/;
  assign _17544_ = inv_32[92] & r_31[92] /*584*/;
  assign _17545_ = _17543_ | _17544_ /*583*/;
  assign _17546_ = inv_32[93] ^ r_31[93] /*581*/;
  assign sum_32[93] = _17546_ ^ _17545_ /*580*/;
  assign _17547_ = _17546_ & _17545_ /*579*/;
  assign _17548_ = inv_32[93] & r_31[93] /*578*/;
  assign _17549_ = _17547_ | _17548_ /*577*/;
  assign _17550_ = _17549_ ^ _17545_ /*576*/;
  assign _17551_ = ~_17550_ /*575*/;
  assign _17552_ = sum_32[93] & _17551_ /*574*/;
  assign _17553_ = _17550_ & _17549_ /*573*/;
  assign sum_32[94] = _17553_ | _17552_ /*572*/;
  assign q[0] = ~sum_32[94] /*571*/;
  assign m_32[0] = r_31[0] /*570*/;
  assign m_32[1] = r_31[1] /*569*/;
  assign m_32[2] = r_31[2] /*568*/;
  assign m_32[3] = r_31[3] /*567*/;
  assign m_32[4] = r_31[4] /*566*/;
  assign m_32[5] = r_31[5] /*565*/;
  assign m_32[6] = r_31[6] /*564*/;
  assign m_32[7] = r_31[7] /*563*/;
  assign m_32[8] = r_31[8] /*562*/;
  assign m_32[9] = r_31[9] /*561*/;
  assign m_32[10] = r_31[10] /*560*/;
  assign m_32[11] = r_31[11] /*559*/;
  assign m_32[12] = r_31[12] /*558*/;
  assign m_32[13] = r_31[13] /*557*/;
  assign m_32[14] = r_31[14] /*556*/;
  assign m_32[15] = r_31[15] /*555*/;
  assign m_32[16] = r_31[16] /*554*/;
  assign m_32[17] = r_31[17] /*553*/;
  assign m_32[18] = r_31[18] /*552*/;
  assign m_32[19] = r_31[19] /*551*/;
  assign m_32[20] = r_31[20] /*550*/;
  assign m_32[21] = r_31[21] /*549*/;
  assign m_32[22] = r_31[22] /*548*/;
  assign m_32[23] = r_31[23] /*547*/;
  assign m_32[24] = r_31[24] /*546*/;
  assign m_32[25] = r_31[25] /*545*/;
  assign m_32[26] = r_31[26] /*544*/;
  assign m_32[27] = r_31[27] /*543*/;
  assign m_32[28] = r_31[28] /*542*/;
  assign m_32[29] = r_31[29] /*541*/;
  assign m_32[30] = r_31[30] /*540*/;
  assign m_32[31] = r_31[31] /*539*/;
  assign m_32[32] = r_31[32] /*538*/;
  assign m_32[33] = r_31[33] /*537*/;
  assign m_32[34] = r_31[34] /*536*/;
  assign m_32[35] = r_31[35] /*535*/;
  assign m_32[36] = r_31[36] /*534*/;
  assign m_32[37] = r_31[37] /*533*/;
  assign m_32[38] = r_31[38] /*532*/;
  assign m_32[39] = r_31[39] /*531*/;
  assign m_32[40] = r_31[40] /*530*/;
  assign m_32[41] = r_31[41] /*529*/;
  assign m_32[42] = r_31[42] /*528*/;
  assign m_32[43] = r_31[43] /*527*/;
  assign m_32[44] = r_31[44] /*526*/;
  assign m_32[45] = r_31[45] /*525*/;
  assign m_32[46] = r_31[46] /*524*/;
  assign m_32[47] = r_31[47] /*523*/;
  assign m_32[48] = r_31[48] /*522*/;
  assign m_32[49] = r_31[49] /*521*/;
  assign m_32[50] = r_31[50] /*520*/;
  assign m_32[51] = r_31[51] /*519*/;
  assign m_32[52] = r_31[52] /*518*/;
  assign m_32[53] = r_31[53] /*517*/;
  assign m_32[54] = r_31[54] /*516*/;
  assign m_32[55] = r_31[55] /*515*/;
  assign m_32[56] = r_31[56] /*514*/;
  assign m_32[57] = r_31[57] /*513*/;
  assign m_32[58] = r_31[58] /*512*/;
  assign m_32[59] = r_31[59] /*511*/;
  assign m_32[60] = r_31[60] /*510*/;
  assign m_32[61] = r_31[61] /*509*/;
  assign m_32[62] = r_31[62] /*508*/;
  assign m_32[63] = r_31[63] /*507*/;
  assign m_32[64] = r_31[64] /*506*/;
  assign m_32[65] = r_31[65] /*505*/;
  assign m_32[66] = r_31[66] /*504*/;
  assign m_32[67] = r_31[67] /*503*/;
  assign m_32[68] = r_31[68] /*502*/;
  assign m_32[69] = r_31[69] /*501*/;
  assign m_32[70] = r_31[70] /*500*/;
  assign m_32[71] = r_31[71] /*499*/;
  assign m_32[72] = r_31[72] /*498*/;
  assign m_32[73] = r_31[73] /*497*/;
  assign m_32[74] = r_31[74] /*496*/;
  assign m_32[75] = r_31[75] /*495*/;
  assign m_32[76] = r_31[76] /*494*/;
  assign m_32[77] = r_31[77] /*493*/;
  assign m_32[78] = r_31[78] /*492*/;
  assign m_32[79] = r_31[79] /*491*/;
  assign m_32[80] = r_31[80] /*490*/;
  assign m_32[81] = r_31[81] /*489*/;
  assign m_32[82] = r_31[82] /*488*/;
  assign m_32[83] = r_31[83] /*487*/;
  assign m_32[84] = r_31[84] /*486*/;
  assign m_32[85] = r_31[85] /*485*/;
  assign m_32[86] = r_31[86] /*484*/;
  assign m_32[87] = r_31[87] /*483*/;
  assign m_32[88] = r_31[88] /*482*/;
  assign m_32[89] = r_31[89] /*481*/;
  assign m_32[90] = r_31[90] /*480*/;
  assign m_32[91] = r_31[91] /*479*/;
  assign m_32[92] = r_31[92] /*478*/;
  assign m_32[93] = r_31[93] /*477*/;
  assign m_32[94] = r_31[93] /*476*/;
  assign _17555_ = ~q[0] /*475*/;
  assign _17556_ = sum_32[0] & q[0] /*474*/;
  assign _17557_ = m_32[0] & _17555_ /*473*/;
  assign r_32[0] = _17557_ | _17556_ /*472*/;
  assign _17558_ = ~q[0] /*471*/;
  assign _17559_ = sum_32[1] & q[0] /*470*/;
  assign _17560_ = m_32[1] & _17558_ /*469*/;
  assign r_32[1] = _17560_ | _17559_ /*468*/;
  assign _17561_ = ~q[0] /*467*/;
  assign _17562_ = sum_32[2] & q[0] /*466*/;
  assign _17563_ = m_32[2] & _17561_ /*465*/;
  assign r_32[2] = _17563_ | _17562_ /*464*/;
  assign _17564_ = ~q[0] /*463*/;
  assign _17565_ = sum_32[3] & q[0] /*462*/;
  assign _17566_ = m_32[3] & _17564_ /*461*/;
  assign r_32[3] = _17566_ | _17565_ /*460*/;
  assign _17567_ = ~q[0] /*459*/;
  assign _17568_ = sum_32[4] & q[0] /*458*/;
  assign _17569_ = m_32[4] & _17567_ /*457*/;
  assign r_32[4] = _17569_ | _17568_ /*456*/;
  assign _17570_ = ~q[0] /*455*/;
  assign _17571_ = sum_32[5] & q[0] /*454*/;
  assign _17572_ = m_32[5] & _17570_ /*453*/;
  assign r_32[5] = _17572_ | _17571_ /*452*/;
  assign _17573_ = ~q[0] /*451*/;
  assign _17574_ = sum_32[6] & q[0] /*450*/;
  assign _17575_ = m_32[6] & _17573_ /*449*/;
  assign r_32[6] = _17575_ | _17574_ /*448*/;
  assign _17576_ = ~q[0] /*447*/;
  assign _17577_ = sum_32[7] & q[0] /*446*/;
  assign _17578_ = m_32[7] & _17576_ /*445*/;
  assign r_32[7] = _17578_ | _17577_ /*444*/;
  assign _17579_ = ~q[0] /*443*/;
  assign _17580_ = sum_32[8] & q[0] /*442*/;
  assign _17581_ = m_32[8] & _17579_ /*441*/;
  assign r_32[8] = _17581_ | _17580_ /*440*/;
  assign _17582_ = ~q[0] /*439*/;
  assign _17583_ = sum_32[9] & q[0] /*438*/;
  assign _17584_ = m_32[9] & _17582_ /*437*/;
  assign r_32[9] = _17584_ | _17583_ /*436*/;
  assign _17585_ = ~q[0] /*435*/;
  assign _17586_ = sum_32[10] & q[0] /*434*/;
  assign _17587_ = m_32[10] & _17585_ /*433*/;
  assign r_32[10] = _17587_ | _17586_ /*432*/;
  assign _17588_ = ~q[0] /*431*/;
  assign _17589_ = sum_32[11] & q[0] /*430*/;
  assign _17590_ = m_32[11] & _17588_ /*429*/;
  assign r_32[11] = _17590_ | _17589_ /*428*/;
  assign _17591_ = ~q[0] /*427*/;
  assign _17592_ = sum_32[12] & q[0] /*426*/;
  assign _17593_ = m_32[12] & _17591_ /*425*/;
  assign r_32[12] = _17593_ | _17592_ /*424*/;
  assign _17594_ = ~q[0] /*423*/;
  assign _17595_ = sum_32[13] & q[0] /*422*/;
  assign _17596_ = m_32[13] & _17594_ /*421*/;
  assign r_32[13] = _17596_ | _17595_ /*420*/;
  assign _17597_ = ~q[0] /*419*/;
  assign _17598_ = sum_32[14] & q[0] /*418*/;
  assign _17599_ = m_32[14] & _17597_ /*417*/;
  assign r_32[14] = _17599_ | _17598_ /*416*/;
  assign _17600_ = ~q[0] /*415*/;
  assign _17601_ = sum_32[15] & q[0] /*414*/;
  assign _17602_ = m_32[15] & _17600_ /*413*/;
  assign r_32[15] = _17602_ | _17601_ /*412*/;
  assign _17603_ = ~q[0] /*411*/;
  assign _17604_ = sum_32[16] & q[0] /*410*/;
  assign _17605_ = m_32[16] & _17603_ /*409*/;
  assign r_32[16] = _17605_ | _17604_ /*408*/;
  assign _17606_ = ~q[0] /*407*/;
  assign _17607_ = sum_32[17] & q[0] /*406*/;
  assign _17608_ = m_32[17] & _17606_ /*405*/;
  assign r_32[17] = _17608_ | _17607_ /*404*/;
  assign _17609_ = ~q[0] /*403*/;
  assign _17610_ = sum_32[18] & q[0] /*402*/;
  assign _17611_ = m_32[18] & _17609_ /*401*/;
  assign r_32[18] = _17611_ | _17610_ /*400*/;
  assign _17612_ = ~q[0] /*399*/;
  assign _17613_ = sum_32[19] & q[0] /*398*/;
  assign _17614_ = m_32[19] & _17612_ /*397*/;
  assign r_32[19] = _17614_ | _17613_ /*396*/;
  assign _17615_ = ~q[0] /*395*/;
  assign _17616_ = sum_32[20] & q[0] /*394*/;
  assign _17617_ = m_32[20] & _17615_ /*393*/;
  assign r_32[20] = _17617_ | _17616_ /*392*/;
  assign _17618_ = ~q[0] /*391*/;
  assign _17619_ = sum_32[21] & q[0] /*390*/;
  assign _17620_ = m_32[21] & _17618_ /*389*/;
  assign r_32[21] = _17620_ | _17619_ /*388*/;
  assign _17621_ = ~q[0] /*387*/;
  assign _17622_ = sum_32[22] & q[0] /*386*/;
  assign _17623_ = m_32[22] & _17621_ /*385*/;
  assign r_32[22] = _17623_ | _17622_ /*384*/;
  assign _17624_ = ~q[0] /*383*/;
  assign _17625_ = sum_32[23] & q[0] /*382*/;
  assign _17626_ = m_32[23] & _17624_ /*381*/;
  assign r_32[23] = _17626_ | _17625_ /*380*/;
  assign _17627_ = ~q[0] /*379*/;
  assign _17628_ = sum_32[24] & q[0] /*378*/;
  assign _17629_ = m_32[24] & _17627_ /*377*/;
  assign r_32[24] = _17629_ | _17628_ /*376*/;
  assign _17630_ = ~q[0] /*375*/;
  assign _17631_ = sum_32[25] & q[0] /*374*/;
  assign _17632_ = m_32[25] & _17630_ /*373*/;
  assign r_32[25] = _17632_ | _17631_ /*372*/;
  assign _17633_ = ~q[0] /*371*/;
  assign _17634_ = sum_32[26] & q[0] /*370*/;
  assign _17635_ = m_32[26] & _17633_ /*369*/;
  assign r_32[26] = _17635_ | _17634_ /*368*/;
  assign _17636_ = ~q[0] /*367*/;
  assign _17637_ = sum_32[27] & q[0] /*366*/;
  assign _17638_ = m_32[27] & _17636_ /*365*/;
  assign r_32[27] = _17638_ | _17637_ /*364*/;
  assign _17639_ = ~q[0] /*363*/;
  assign _17640_ = sum_32[28] & q[0] /*362*/;
  assign _17641_ = m_32[28] & _17639_ /*361*/;
  assign r_32[28] = _17641_ | _17640_ /*360*/;
  assign _17642_ = ~q[0] /*359*/;
  assign _17643_ = sum_32[29] & q[0] /*358*/;
  assign _17644_ = m_32[29] & _17642_ /*357*/;
  assign r_32[29] = _17644_ | _17643_ /*356*/;
  assign _17645_ = ~q[0] /*355*/;
  assign _17646_ = sum_32[30] & q[0] /*354*/;
  assign _17647_ = m_32[30] & _17645_ /*353*/;
  assign r_32[30] = _17647_ | _17646_ /*352*/;
  assign _17648_ = ~q[0] /*351*/;
  assign _17649_ = sum_32[31] & q[0] /*350*/;
  assign _17650_ = m_32[31] & _17648_ /*349*/;
  assign r_32[31] = _17650_ | _17649_ /*348*/;
  assign _17651_ = ~q[0] /*347*/;
  assign _17652_ = sum_32[32] & q[0] /*346*/;
  assign _17653_ = m_32[32] & _17651_ /*345*/;
  assign r_32[32] = _17653_ | _17652_ /*344*/;
  assign _17654_ = ~q[0] /*343*/;
  assign _17655_ = sum_32[33] & q[0] /*342*/;
  assign _17656_ = m_32[33] & _17654_ /*341*/;
  assign r_32[33] = _17656_ | _17655_ /*340*/;
  assign _17657_ = ~q[0] /*339*/;
  assign _17658_ = sum_32[34] & q[0] /*338*/;
  assign _17659_ = m_32[34] & _17657_ /*337*/;
  assign r_32[34] = _17659_ | _17658_ /*336*/;
  assign _17660_ = ~q[0] /*335*/;
  assign _17661_ = sum_32[35] & q[0] /*334*/;
  assign _17662_ = m_32[35] & _17660_ /*333*/;
  assign r_32[35] = _17662_ | _17661_ /*332*/;
  assign _17663_ = ~q[0] /*331*/;
  assign _17664_ = sum_32[36] & q[0] /*330*/;
  assign _17665_ = m_32[36] & _17663_ /*329*/;
  assign r_32[36] = _17665_ | _17664_ /*328*/;
  assign _17666_ = ~q[0] /*327*/;
  assign _17667_ = sum_32[37] & q[0] /*326*/;
  assign _17668_ = m_32[37] & _17666_ /*325*/;
  assign r_32[37] = _17668_ | _17667_ /*324*/;
  assign _17669_ = ~q[0] /*323*/;
  assign _17670_ = sum_32[38] & q[0] /*322*/;
  assign _17671_ = m_32[38] & _17669_ /*321*/;
  assign r_32[38] = _17671_ | _17670_ /*320*/;
  assign _17672_ = ~q[0] /*319*/;
  assign _17673_ = sum_32[39] & q[0] /*318*/;
  assign _17674_ = m_32[39] & _17672_ /*317*/;
  assign r_32[39] = _17674_ | _17673_ /*316*/;
  assign _17675_ = ~q[0] /*315*/;
  assign _17676_ = sum_32[40] & q[0] /*314*/;
  assign _17677_ = m_32[40] & _17675_ /*313*/;
  assign r_32[40] = _17677_ | _17676_ /*312*/;
  assign _17678_ = ~q[0] /*311*/;
  assign _17679_ = sum_32[41] & q[0] /*310*/;
  assign _17680_ = m_32[41] & _17678_ /*309*/;
  assign r_32[41] = _17680_ | _17679_ /*308*/;
  assign _17681_ = ~q[0] /*307*/;
  assign _17682_ = sum_32[42] & q[0] /*306*/;
  assign _17683_ = m_32[42] & _17681_ /*305*/;
  assign r_32[42] = _17683_ | _17682_ /*304*/;
  assign _17684_ = ~q[0] /*303*/;
  assign _17685_ = sum_32[43] & q[0] /*302*/;
  assign _17686_ = m_32[43] & _17684_ /*301*/;
  assign r_32[43] = _17686_ | _17685_ /*300*/;
  assign _17687_ = ~q[0] /*299*/;
  assign _17688_ = sum_32[44] & q[0] /*298*/;
  assign _17689_ = m_32[44] & _17687_ /*297*/;
  assign r_32[44] = _17689_ | _17688_ /*296*/;
  assign _17690_ = ~q[0] /*295*/;
  assign _17691_ = sum_32[45] & q[0] /*294*/;
  assign _17692_ = m_32[45] & _17690_ /*293*/;
  assign r_32[45] = _17692_ | _17691_ /*292*/;
  assign _17693_ = ~q[0] /*291*/;
  assign _17694_ = sum_32[46] & q[0] /*290*/;
  assign _17695_ = m_32[46] & _17693_ /*289*/;
  assign r_32[46] = _17695_ | _17694_ /*288*/;
  assign _17696_ = ~q[0] /*287*/;
  assign _17697_ = sum_32[47] & q[0] /*286*/;
  assign _17698_ = m_32[47] & _17696_ /*285*/;
  assign r_32[47] = _17698_ | _17697_ /*284*/;
  assign _17699_ = ~q[0] /*283*/;
  assign _17700_ = sum_32[48] & q[0] /*282*/;
  assign _17701_ = m_32[48] & _17699_ /*281*/;
  assign r_32[48] = _17701_ | _17700_ /*280*/;
  assign _17702_ = ~q[0] /*279*/;
  assign _17703_ = sum_32[49] & q[0] /*278*/;
  assign _17704_ = m_32[49] & _17702_ /*277*/;
  assign r_32[49] = _17704_ | _17703_ /*276*/;
  assign _17705_ = ~q[0] /*275*/;
  assign _17706_ = sum_32[50] & q[0] /*274*/;
  assign _17707_ = m_32[50] & _17705_ /*273*/;
  assign r_32[50] = _17707_ | _17706_ /*272*/;
  assign _17708_ = ~q[0] /*271*/;
  assign _17709_ = sum_32[51] & q[0] /*270*/;
  assign _17710_ = m_32[51] & _17708_ /*269*/;
  assign r_32[51] = _17710_ | _17709_ /*268*/;
  assign _17711_ = ~q[0] /*267*/;
  assign _17712_ = sum_32[52] & q[0] /*266*/;
  assign _17713_ = m_32[52] & _17711_ /*265*/;
  assign r_32[52] = _17713_ | _17712_ /*264*/;
  assign _17714_ = ~q[0] /*263*/;
  assign _17715_ = sum_32[53] & q[0] /*262*/;
  assign _17716_ = m_32[53] & _17714_ /*261*/;
  assign r_32[53] = _17716_ | _17715_ /*260*/;
  assign _17717_ = ~q[0] /*259*/;
  assign _17718_ = sum_32[54] & q[0] /*258*/;
  assign _17719_ = m_32[54] & _17717_ /*257*/;
  assign r_32[54] = _17719_ | _17718_ /*256*/;
  assign _17720_ = ~q[0] /*255*/;
  assign _17721_ = sum_32[55] & q[0] /*254*/;
  assign _17722_ = m_32[55] & _17720_ /*253*/;
  assign r_32[55] = _17722_ | _17721_ /*252*/;
  assign _17723_ = ~q[0] /*251*/;
  assign _17724_ = sum_32[56] & q[0] /*250*/;
  assign _17725_ = m_32[56] & _17723_ /*249*/;
  assign r_32[56] = _17725_ | _17724_ /*248*/;
  assign _17726_ = ~q[0] /*247*/;
  assign _17727_ = sum_32[57] & q[0] /*246*/;
  assign _17728_ = m_32[57] & _17726_ /*245*/;
  assign r_32[57] = _17728_ | _17727_ /*244*/;
  assign _17729_ = ~q[0] /*243*/;
  assign _17730_ = sum_32[58] & q[0] /*242*/;
  assign _17731_ = m_32[58] & _17729_ /*241*/;
  assign r_32[58] = _17731_ | _17730_ /*240*/;
  assign _17732_ = ~q[0] /*239*/;
  assign _17733_ = sum_32[59] & q[0] /*238*/;
  assign _17734_ = m_32[59] & _17732_ /*237*/;
  assign r_32[59] = _17734_ | _17733_ /*236*/;
  assign _17735_ = ~q[0] /*235*/;
  assign _17736_ = sum_32[60] & q[0] /*234*/;
  assign _17737_ = m_32[60] & _17735_ /*233*/;
  assign r_32[60] = _17737_ | _17736_ /*232*/;
  assign _17738_ = ~q[0] /*231*/;
  assign _17739_ = sum_32[61] & q[0] /*230*/;
  assign _17740_ = m_32[61] & _17738_ /*229*/;
  assign r_32[61] = _17740_ | _17739_ /*228*/;
  assign _17741_ = ~q[0] /*227*/;
  assign _17742_ = sum_32[62] & q[0] /*226*/;
  assign _17743_ = m_32[62] & _17741_ /*225*/;
  assign r_32[62] = _17743_ | _17742_ /*224*/;
  assign _17744_ = ~q[0] /*223*/;
  assign _17745_ = sum_32[63] & q[0] /*222*/;
  assign _17746_ = m_32[63] & _17744_ /*221*/;
  assign r_32[63] = _17746_ | _17745_ /*220*/;
  assign _17747_ = ~q[0] /*219*/;
  assign _17748_ = sum_32[64] & q[0] /*218*/;
  assign _17749_ = m_32[64] & _17747_ /*217*/;
  assign r_32[64] = _17749_ | _17748_ /*216*/;
  assign _17750_ = ~q[0] /*215*/;
  assign _17751_ = sum_32[65] & q[0] /*214*/;
  assign _17752_ = m_32[65] & _17750_ /*213*/;
  assign r_32[65] = _17752_ | _17751_ /*212*/;
  assign _17753_ = ~q[0] /*211*/;
  assign _17754_ = sum_32[66] & q[0] /*210*/;
  assign _17755_ = m_32[66] & _17753_ /*209*/;
  assign r_32[66] = _17755_ | _17754_ /*208*/;
  assign _17756_ = ~q[0] /*207*/;
  assign _17757_ = sum_32[67] & q[0] /*206*/;
  assign _17758_ = m_32[67] & _17756_ /*205*/;
  assign r_32[67] = _17758_ | _17757_ /*204*/;
  assign _17759_ = ~q[0] /*203*/;
  assign _17760_ = sum_32[68] & q[0] /*202*/;
  assign _17761_ = m_32[68] & _17759_ /*201*/;
  assign r_32[68] = _17761_ | _17760_ /*200*/;
  assign _17762_ = ~q[0] /*199*/;
  assign _17763_ = sum_32[69] & q[0] /*198*/;
  assign _17764_ = m_32[69] & _17762_ /*197*/;
  assign r_32[69] = _17764_ | _17763_ /*196*/;
  assign _17765_ = ~q[0] /*195*/;
  assign _17766_ = sum_32[70] & q[0] /*194*/;
  assign _17767_ = m_32[70] & _17765_ /*193*/;
  assign r_32[70] = _17767_ | _17766_ /*192*/;
  assign _17768_ = ~q[0] /*191*/;
  assign _17769_ = sum_32[71] & q[0] /*190*/;
  assign _17770_ = m_32[71] & _17768_ /*189*/;
  assign r_32[71] = _17770_ | _17769_ /*188*/;
  assign _17771_ = ~q[0] /*187*/;
  assign _17772_ = sum_32[72] & q[0] /*186*/;
  assign _17773_ = m_32[72] & _17771_ /*185*/;
  assign r_32[72] = _17773_ | _17772_ /*184*/;
  assign _17774_ = ~q[0] /*183*/;
  assign _17775_ = sum_32[73] & q[0] /*182*/;
  assign _17776_ = m_32[73] & _17774_ /*181*/;
  assign r_32[73] = _17776_ | _17775_ /*180*/;
  assign _17777_ = ~q[0] /*179*/;
  assign _17778_ = sum_32[74] & q[0] /*178*/;
  assign _17779_ = m_32[74] & _17777_ /*177*/;
  assign r_32[74] = _17779_ | _17778_ /*176*/;
  assign _17780_ = ~q[0] /*175*/;
  assign _17781_ = sum_32[75] & q[0] /*174*/;
  assign _17782_ = m_32[75] & _17780_ /*173*/;
  assign r_32[75] = _17782_ | _17781_ /*172*/;
  assign _17783_ = ~q[0] /*171*/;
  assign _17784_ = sum_32[76] & q[0] /*170*/;
  assign _17785_ = m_32[76] & _17783_ /*169*/;
  assign r_32[76] = _17785_ | _17784_ /*168*/;
  assign _17786_ = ~q[0] /*167*/;
  assign _17787_ = sum_32[77] & q[0] /*166*/;
  assign _17788_ = m_32[77] & _17786_ /*165*/;
  assign r_32[77] = _17788_ | _17787_ /*164*/;
  assign _17789_ = ~q[0] /*163*/;
  assign _17790_ = sum_32[78] & q[0] /*162*/;
  assign _17791_ = m_32[78] & _17789_ /*161*/;
  assign r_32[78] = _17791_ | _17790_ /*160*/;
  assign _17792_ = ~q[0] /*159*/;
  assign _17793_ = sum_32[79] & q[0] /*158*/;
  assign _17794_ = m_32[79] & _17792_ /*157*/;
  assign r_32[79] = _17794_ | _17793_ /*156*/;
  assign _17795_ = ~q[0] /*155*/;
  assign _17796_ = sum_32[80] & q[0] /*154*/;
  assign _17797_ = m_32[80] & _17795_ /*153*/;
  assign r_32[80] = _17797_ | _17796_ /*152*/;
  assign _17798_ = ~q[0] /*151*/;
  assign _17799_ = sum_32[81] & q[0] /*150*/;
  assign _17800_ = m_32[81] & _17798_ /*149*/;
  assign r_32[81] = _17800_ | _17799_ /*148*/;
  assign _17801_ = ~q[0] /*147*/;
  assign _17802_ = sum_32[82] & q[0] /*146*/;
  assign _17803_ = m_32[82] & _17801_ /*145*/;
  assign r_32[82] = _17803_ | _17802_ /*144*/;
  assign _17804_ = ~q[0] /*143*/;
  assign _17805_ = sum_32[83] & q[0] /*142*/;
  assign _17806_ = m_32[83] & _17804_ /*141*/;
  assign r_32[83] = _17806_ | _17805_ /*140*/;
  assign _17807_ = ~q[0] /*139*/;
  assign _17808_ = sum_32[84] & q[0] /*138*/;
  assign _17809_ = m_32[84] & _17807_ /*137*/;
  assign r_32[84] = _17809_ | _17808_ /*136*/;
  assign _17810_ = ~q[0] /*135*/;
  assign _17811_ = sum_32[85] & q[0] /*134*/;
  assign _17812_ = m_32[85] & _17810_ /*133*/;
  assign r_32[85] = _17812_ | _17811_ /*132*/;
  assign _17813_ = ~q[0] /*131*/;
  assign _17814_ = sum_32[86] & q[0] /*130*/;
  assign _17815_ = m_32[86] & _17813_ /*129*/;
  assign r_32[86] = _17815_ | _17814_ /*128*/;
  assign _17816_ = ~q[0] /*127*/;
  assign _17817_ = sum_32[87] & q[0] /*126*/;
  assign _17818_ = m_32[87] & _17816_ /*125*/;
  assign r_32[87] = _17818_ | _17817_ /*124*/;
  assign _17819_ = ~q[0] /*123*/;
  assign _17820_ = sum_32[88] & q[0] /*122*/;
  assign _17821_ = m_32[88] & _17819_ /*121*/;
  assign r_32[88] = _17821_ | _17820_ /*120*/;
  assign _17822_ = ~q[0] /*119*/;
  assign _17823_ = sum_32[89] & q[0] /*118*/;
  assign _17824_ = m_32[89] & _17822_ /*117*/;
  assign r_32[89] = _17824_ | _17823_ /*116*/;
  assign _17825_ = ~q[0] /*115*/;
  assign _17826_ = sum_32[90] & q[0] /*114*/;
  assign _17827_ = m_32[90] & _17825_ /*113*/;
  assign r_32[90] = _17827_ | _17826_ /*112*/;
  assign _17828_ = ~q[0] /*111*/;
  assign _17829_ = sum_32[91] & q[0] /*110*/;
  assign _17830_ = m_32[91] & _17828_ /*109*/;
  assign r_32[91] = _17830_ | _17829_ /*108*/;
  assign _17831_ = ~q[0] /*107*/;
  assign _17832_ = sum_32[92] & q[0] /*106*/;
  assign _17833_ = m_32[92] & _17831_ /*105*/;
  assign r_32[92] = _17833_ | _17832_ /*104*/;
  assign _17834_ = ~q[0] /*103*/;
  assign _17835_ = sum_32[93] & q[0] /*102*/;
  assign _17836_ = m_32[93] & _17834_ /*101*/;
  assign r_32[93] = _17836_ | _17835_ /*100*/;
  assign _17837_ = ~q[0] /*99*/;
  assign _17838_ = sum_32[94] & q[0] /*98*/;
  assign _17839_ = m_32[94] & _17837_ /*97*/;
  assign r_32[94] = _17839_ | _17838_ /*96*/;
  assign rout[0] = r_32[0] /*0*/;
  assign rout[1] = r_32[1] /*1*/;
  assign rout[2] = r_32[2] /*2*/;
  assign rout[3] = r_32[3] /*3*/;
  assign rout[4] = r_32[4] /*4*/;
  assign rout[5] = r_32[5] /*5*/;
  assign rout[6] = r_32[6] /*6*/;
  assign rout[7] = r_32[7] /*7*/;
  assign rout[8] = r_32[8] /*8*/;
  assign rout[9] = r_32[9] /*9*/;
  assign rout[10] = r_32[10] /*10*/;
  assign rout[11] = r_32[11] /*11*/;
  assign rout[12] = r_32[12] /*12*/;
  assign rout[13] = r_32[13] /*13*/;
  assign rout[14] = r_32[14] /*14*/;
  assign rout[15] = r_32[15] /*15*/;
  assign rout[16] = r_32[16] /*16*/;
  assign rout[17] = r_32[17] /*17*/;
  assign rout[18] = r_32[18] /*18*/;
  assign rout[19] = r_32[19] /*19*/;
  assign rout[20] = r_32[20] /*20*/;
  assign rout[21] = r_32[21] /*21*/;
  assign rout[22] = r_32[22] /*22*/;
  assign rout[23] = r_32[23] /*23*/;
  assign rout[24] = r_32[24] /*24*/;
  assign rout[25] = r_32[25] /*25*/;
  assign rout[26] = r_32[26] /*26*/;
  assign rout[27] = r_32[27] /*27*/;
  assign rout[28] = r_32[28] /*28*/;
  assign rout[29] = r_32[29] /*29*/;
  assign rout[30] = r_32[30] /*30*/;
  assign rout[31] = r_32[31] /*31*/;
  assign rout[32] = r_32[32] /*32*/;
  assign rout[33] = r_32[33] /*33*/;
  assign rout[34] = r_32[34] /*34*/;
  assign rout[35] = r_32[35] /*35*/;
  assign rout[36] = r_32[36] /*36*/;
  assign rout[37] = r_32[37] /*37*/;
  assign rout[38] = r_32[38] /*38*/;
  assign rout[39] = r_32[39] /*39*/;
  assign rout[40] = r_32[40] /*40*/;
  assign rout[41] = r_32[41] /*41*/;
  assign rout[42] = r_32[42] /*42*/;
  assign rout[43] = r_32[43] /*43*/;
  assign rout[44] = r_32[44] /*44*/;
  assign rout[45] = r_32[45] /*45*/;
  assign rout[46] = r_32[46] /*46*/;
  assign rout[47] = r_32[47] /*47*/;
  assign rout[48] = r_32[48] /*48*/;
  assign rout[49] = r_32[49] /*49*/;
  assign rout[50] = r_32[50] /*50*/;
  assign rout[51] = r_32[51] /*51*/;
  assign rout[52] = r_32[52] /*52*/;
  assign rout[53] = r_32[53] /*53*/;
  assign rout[54] = r_32[54] /*54*/;
  assign rout[55] = r_32[55] /*55*/;
  assign rout[56] = r_32[56] /*56*/;
  assign rout[57] = r_32[57] /*57*/;
  assign rout[58] = r_32[58] /*58*/;
  assign rout[59] = r_32[59] /*59*/;
  assign rout[60] = r_32[60] /*60*/;
  assign rout[61] = r_32[61] /*61*/;
  assign rout[62] = r_32[62] /*62*/;
  assign rout[63] = r_32[63] /*63*/;
  assign rout[64] = r_32[64] /*64*/;
  assign rout[65] = r_32[65] /*65*/;
  assign rout[66] = r_32[66] /*66*/;
  assign rout[67] = r_32[67] /*67*/;
  assign rout[68] = r_32[68] /*68*/;
  assign rout[69] = r_32[69] /*69*/;
  assign rout[70] = r_32[70] /*70*/;
  assign rout[71] = r_32[71] /*71*/;
  assign rout[72] = r_32[72] /*72*/;
  assign rout[73] = r_32[73] /*73*/;
  assign rout[74] = r_32[74] /*74*/;
  assign rout[75] = r_32[75] /*75*/;
  assign rout[76] = r_32[76] /*76*/;
  assign rout[77] = r_32[77] /*77*/;
  assign rout[78] = r_32[78] /*78*/;
  assign rout[79] = r_32[79] /*79*/;
  assign rout[80] = r_32[80] /*80*/;
  assign rout[81] = r_32[81] /*81*/;
  assign rout[82] = r_32[82] /*82*/;
  assign rout[83] = r_32[83] /*83*/;
  assign rout[84] = r_32[84] /*84*/;
  assign rout[85] = r_32[85] /*85*/;
  assign rout[86] = r_32[86] /*86*/;
  assign rout[87] = r_32[87] /*87*/;
  assign rout[88] = r_32[88] /*88*/;
  assign rout[89] = r_32[89] /*89*/;
  assign rout[90] = r_32[90] /*90*/;
  assign rout[91] = r_32[91] /*91*/;
  assign rout[92] = r_32[92] /*92*/;
  assign rout[93] = r_32[93] /*93*/;
  assign rout[94] = r_32[94] /*94*/;
endmodule