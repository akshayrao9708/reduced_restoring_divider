module nonresdivReduced(R_0, D, Q, R_n1);
input [5:0] R_0;
input [2:0] D;
output [3:0] Q;
output [2:0] R_n1;
wire _0_;
wire _1_;
wire _2_;
wire _3_;
wire _4_;
wire _5_;
wire _6_;
wire _7_;
wire _8_;
wire _9_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire _30_;
wire _31_;
wire _32_;
wire _33_;
wire _34_;
wire _35_;
wire _36_;
wire _37_;
wire _38_;
wire _39_;
wire _40_;
wire _41_;
wire _42_;
wire _43_;
wire _44_;
wire _45_;
wire _46_;
wire _47_;
wire _48_;
wire _49_;
wire _50_;
wire _51_;
wire _52_;
wire _53_;
wire _54_;
wire _55_;
wire _56_;
wire _57_;
wire _58_;
wire _59_;
wire _60_;
wire _61_;
wire _62_;
wire _63_;
wire _64_;
wire _65_;
wire _66_;
wire _67_;
wire _68_;
wire _69_;
wire _70_;
wire _71_;
wire _72_;
wire _73_;
wire _74_;
wire _75_;
wire _76_;
wire _77_;
wire _78_;
wire _79_;
wire _80_;
wire _81_;
wire _82_;
wire _83_;
wire _84_;
wire _85_;
wire _86_;
wire _87_;
wire _88_;
wire _89_;
wire _90_;
wire _91_;
wire _92_;
wire _93_;
wire _94_;
wire _95_;
wire _96_;
wire _97_;
wire _98_;
wire _99_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire zeroWire;
wire oneWire;
assign zeroWire = 1'b0 /*255*/;
assign oneWire = 1'b1 /*255*/;
assign _9_ = ~D[0] /*229*/;
assign _6_ = R_0[3] & _9_ /*225*/;
assign _7_ = R_0[3] ^ _9_ /*228*/;
assign _8_ = oneWire & _7_ /*226*/;
assign _0_ = oneWire ^ _7_ /*227*/;
assign _5_ = _6_ | _8_ /*224*/;
assign _14_ = ~D[1] /*223*/;
assign _11_ = R_0[4] & _14_ /*219*/;
assign _12_ = R_0[4] ^ _14_ /*222*/;
assign _13_ = _5_ & _12_ /*220*/;
assign _1_ = _5_ ^ _12_ /*221*/;
assign _10_ = _11_ | _13_ /*218*/;
assign _19_ = ~D[2] /*217*/;
assign _16_ = R_0[5] & _19_ /*213*/;
assign _17_ = R_0[5] ^ _19_ /*216*/;
assign _18_ = _10_ & _17_ /*214*/;
assign _2_ = _10_ ^ _17_ /*215*/;
assign _15_ = _16_ | _18_ /*212*/;
assign _20_ = zeroWire & oneWire /*207*/;
assign _21_ = zeroWire ^ oneWire /*210*/;
assign _22_ = _15_ & _21_ /*208*/;
assign _3_ = _15_ ^ _21_ /*209*/;
assign Q[3] = _20_ | _22_ /*206*/;
assign _34_ = D[0] ^ Q[3] /*182*/;
assign _31_ = R_0[2] & _34_ /*178*/;
assign _32_ = R_0[2] ^ _34_ /*181*/;
assign _33_ = Q[3] & _32_ /*179*/;
assign _25_ = Q[3] ^ _32_ /*180*/;
assign _30_ = _31_ | _33_ /*177*/;
assign _39_ = D[1] ^ Q[3] /*176*/;
assign _36_ = _0_ & _39_ /*172*/;
assign _37_ = _0_ ^ _39_ /*175*/;
assign _38_ = _30_ & _37_ /*173*/;
assign _26_ = _30_ ^ _37_ /*174*/;
assign _35_ = _36_ | _38_ /*171*/;
assign _44_ = D[2] ^ Q[3] /*170*/;
assign _41_ = _1_ & _44_ /*166*/;
assign _42_ = _1_ ^ _44_ /*169*/;
assign _43_ = _35_ & _42_ /*167*/;
assign _27_ = _35_ ^ _42_ /*168*/;
assign _40_ = _41_ | _43_ /*165*/;
assign _48_ = zeroWire ^ Q[3] /*164*/;
assign _45_ = _2_ & _48_ /*160*/;
assign _46_ = _2_ ^ _48_ /*163*/;
assign _47_ = _40_ & _46_ /*161*/;
assign _28_ = _40_ ^ _46_ /*162*/;
assign Q[2] = _45_ | _47_ /*159*/;
assign _59_ = D[0] ^ Q[2] /*133*/;
assign _56_ = R_0[1] & _59_ /*129*/;
assign _57_ = R_0[1] ^ _59_ /*132*/;
assign _58_ = Q[2] & _57_ /*130*/;
assign _50_ = Q[2] ^ _57_ /*131*/;
assign _55_ = _56_ | _58_ /*128*/;
assign _64_ = D[1] ^ Q[2] /*127*/;
assign _61_ = _25_ & _64_ /*123*/;
assign _62_ = _25_ ^ _64_ /*126*/;
assign _63_ = _55_ & _62_ /*124*/;
assign _51_ = _55_ ^ _62_ /*125*/;
assign _60_ = _61_ | _63_ /*122*/;
assign _69_ = D[2] ^ Q[2] /*121*/;
assign _66_ = _26_ & _69_ /*117*/;
assign _67_ = _26_ ^ _69_ /*120*/;
assign _68_ = _60_ & _67_ /*118*/;
assign _52_ = _60_ ^ _67_ /*119*/;
assign _65_ = _66_ | _68_ /*116*/;
assign _73_ = zeroWire ^ Q[2] /*115*/;
assign _70_ = _27_ & _73_ /*111*/;
assign _71_ = _27_ ^ _73_ /*114*/;
assign _72_ = _65_ & _71_ /*112*/;
assign _53_ = _65_ ^ _71_ /*113*/;
assign Q[1] = _70_ | _72_ /*110*/;
assign _84_ = D[0] ^ Q[1] /*84*/;
assign _81_ = R_0[0] & _84_ /*80*/;
assign _82_ = R_0[0] ^ _84_ /*83*/;
assign _83_ = Q[1] & _82_ /*81*/;
assign _75_ = Q[1] ^ _82_ /*82*/;
assign _80_ = _81_ | _83_ /*79*/;
assign _89_ = D[1] ^ Q[1] /*78*/;
assign _86_ = _50_ & _89_ /*74*/;
assign _87_ = _50_ ^ _89_ /*77*/;
assign _88_ = _80_ & _87_ /*75*/;
assign _76_ = _80_ ^ _87_ /*76*/;
assign _85_ = _86_ | _88_ /*73*/;
assign _94_ = D[2] ^ Q[1] /*72*/;
assign _91_ = _51_ & _94_ /*68*/;
assign _92_ = _51_ ^ _94_ /*71*/;
assign _93_ = _85_ & _92_ /*69*/;
assign _77_ = _85_ ^ _92_ /*70*/;
assign _90_ = _91_ | _93_ /*67*/;
assign _98_ = zeroWire ^ Q[1] /*66*/;
assign _95_ = _52_ & _98_ /*62*/;
assign _96_ = _52_ ^ _98_ /*65*/;
assign _97_ = _90_ & _96_ /*63*/;
assign _78_ = _90_ ^ _96_ /*64*/;
assign Q[0] = _95_ | _97_ /*61*/;
assign _102_ = ~Q[0] /*34*/;
assign _101_ = _102_ & D[0] /*33*/;
assign _104_ = _75_ & _101_ /*28*/;
assign _105_ = _75_ ^ _101_ /*31*/;
assign _106_ = zeroWire & _105_ /*29*/;
assign R_n1[0] = zeroWire ^ _105_ /*30*/;
assign _103_ = _104_ | _106_ /*27*/;
assign _108_ = ~Q[0] /*26*/;
assign _107_ = _108_ & D[1] /*25*/;
assign _110_ = _76_ & _107_ /*20*/;
assign _111_ = _76_ ^ _107_ /*23*/;
assign _112_ = _103_ & _111_ /*21*/;
assign R_n1[1] = _103_ ^ _111_ /*22*/;
assign _109_ = _110_ | _112_ /*19*/;
assign _114_ = ~Q[0] /*18*/;
assign _113_ = _114_ & D[2] /*17*/;
assign _116_ = _77_ & _113_ /*12*/;
assign _117_ = _77_ ^ _113_ /*15*/;
assign _118_ = _109_ & _117_ /*13*/;
assign R_n1[2] = _109_ ^ _117_ /*14*/;
assign _115_ = _116_ | _118_ /*11*/;
endmodule
