module divider(q, rout, rin, div);
  wire _0_;
  wire _1_;
  wire _2_;
  wire _3_;
  wire _4_;
  wire _5_;
  wire _6_;
  wire _7_;
  wire _8_;
  wire _9_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  wire _38_;
  wire _39_;
  wire _40_;
  wire _41_;
  wire _42_;
  wire _43_;
  wire _44_;
  wire _45_;
  wire _46_;
  wire _47_;
  wire _48_;
  wire _49_;
  wire _50_;
  wire _51_;
  wire _52_;
  wire _53_;
  wire _54_;
  wire _55_;
  wire _56_;
  wire _57_;
  wire _58_;
  wire _59_;
  wire _60_;
  wire _61_;
  wire _62_;
  wire _63_;
  wire _64_;
  wire _65_;
  wire _66_;
  wire _67_;
  wire _68_;
  wire _69_;
  wire _70_;
  wire _71_;
  wire _72_;
  wire _73_;
  wire _74_;
  wire _75_;
  wire _76_;
  wire _77_;
  wire _78_;
  wire _79_;
  wire _80_;
  wire _81_;
  wire _82_;
  wire _83_;
  wire _84_;
  wire _85_;
  wire _86_;
  wire _87_;
  wire _88_;
  wire _89_;
  wire _90_;
  wire _91_;
  wire _92_;
  wire _93_;
  wire _94_;
  wire _95_;
  wire _96_;
  wire _97_;
  wire _98_;
  wire _99_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire _304_;
  wire _305_;
  wire _306_;
  wire _307_;
  wire _308_;
  wire _309_;
  wire _310_;
  wire _311_;
  wire _312_;
  wire _313_;
  wire _314_;
  wire _315_;
  wire _316_;
  wire _317_;
  wire _318_;
  wire _319_;
  wire _320_;
  wire _321_;
  wire _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire _326_;
  wire _327_;
  wire _328_;
  wire _329_;
  wire _330_;
  wire _331_;
  wire _332_;
  wire _333_;
  wire _334_;
  wire _335_;
  wire _336_;
  wire _337_;
  wire _338_;
  wire _339_;
  wire _340_;
  wire _341_;
  wire _342_;
  wire _343_;
  wire _344_;
  wire _345_;
  wire _346_;
  wire _347_;
  wire _348_;
  wire _349_;
  wire _350_;
  wire _351_;
  wire _352_;
  wire _353_;
  wire _354_;
  wire _355_;
  wire _356_;
  wire _357_;
  wire _358_;
  wire _359_;
  wire _360_;
  wire _361_;
  wire _362_;
  wire _363_;
  wire _364_;
  wire _365_;
  wire _366_;
  wire _367_;
  wire _368_;
  wire _369_;
  wire _370_;
  wire _371_;
  wire _372_;
  wire _373_;
  wire _374_;
  wire _375_;
  wire _376_;
  wire _377_;
  wire _378_;
  wire _379_;
  wire _380_;
  wire _381_;
  wire _382_;
  wire _383_;
  wire _384_;
  wire _385_;
  wire _386_;
  wire _387_;
  wire _388_;
  wire _389_;
  wire _390_;
  wire _391_;
  wire _392_;
  wire _393_;
  wire _394_;
  wire _395_;
  wire _396_;
  wire _397_;
  wire _398_;
  wire _399_;
  wire _400_;
  wire _401_;
  wire _402_;
  wire _403_;
  wire _404_;
  wire _405_;
  wire _406_;
  wire _407_;
  wire _408_;
  wire _409_;
  wire _410_;
  wire _411_;
  wire _412_;
  wire _413_;
  wire _414_;
  wire _415_;
  wire _416_;
  wire _417_;
  wire _418_;
  wire _419_;
  wire _420_;
  wire _421_;
  wire _422_;
  wire _423_;
  wire _424_;
  wire _425_;
  wire _426_;
  wire _427_;
  wire _428_;
  wire _429_;
  wire _430_;
  wire _431_;
  wire _432_;
  wire _433_;
  wire _434_;
  wire _435_;
  wire _436_;
  wire _437_;
  wire _438_;
  wire _439_;
  wire _440_;
  wire _441_;
  wire _442_;
  wire _443_;
  wire _444_;
  wire _445_;
  wire _446_;
  wire _447_;
  wire _448_;
  wire _449_;
  wire _450_;
  wire _451_;
  wire _452_;
  wire _453_;
  wire _454_;
  wire _455_;
  wire _456_;
  wire _457_;
  wire _458_;
  wire _459_;
  wire _460_;
  wire _461_;
  wire _462_;
  wire _463_;
  wire _464_;
  wire _465_;
  wire _466_;
  wire _467_;
  wire _468_;
  wire _469_;
  wire _470_;
  wire _471_;
  wire _472_;
  wire _473_;
  wire _474_;
  wire _475_;
  wire _476_;
  wire _477_;
  wire _478_;
  wire _479_;
  wire _480_;
  wire _481_;
  wire _482_;
  wire _483_;
  wire _484_;
  wire _485_;
  wire _486_;
  wire _487_;
  wire _488_;
  wire _489_;
  wire _490_;
  wire _491_;
  wire _492_;
  wire _493_;
  wire _494_;
  wire _495_;
  wire _496_;
  wire _497_;
  wire _498_;
  wire _499_;
  wire _500_;
  wire _501_;
  wire _502_;
  wire _503_;
  wire _504_;
  wire _505_;
  wire _506_;
  wire _507_;
  wire _508_;
  wire _509_;
  wire _510_;
  wire _511_;
  wire _512_;
  wire _513_;
  wire _514_;
  wire _515_;
  wire _516_;
  wire _517_;
  wire _518_;
  wire _519_;
  wire _520_;
  wire _521_;
  wire _522_;
  wire _523_;
  wire _524_;
  wire _525_;
  wire _526_;
  wire _527_;
  wire _528_;
  wire _529_;
  wire _530_;
  wire _531_;
  wire _532_;
  wire _533_;
  wire _534_;
  wire _535_;
  wire _536_;
  wire _537_;
  wire _538_;
  wire _539_;
  wire _540_;
  wire _541_;
  wire _542_;
  wire _543_;
  wire _544_;
  wire _545_;
  wire _546_;
  wire _547_;
  wire _548_;
  wire _549_;
  wire _550_;
  wire _551_;
  wire _552_;
  wire _553_;
  wire _554_;
  wire _555_;
  wire _556_;
  wire _557_;
  wire _558_;
  wire _559_;
  wire _560_;
  wire _561_;
  wire _562_;
  wire _563_;
  wire _564_;
  wire _565_;
  wire _566_;
  wire _567_;
  wire _568_;
  wire _569_;
  wire _570_;
  wire _571_;
  wire _572_;
  wire _573_;
  wire _574_;
  wire _575_;
  wire _576_;
  wire _577_;
  wire _578_;
  wire _579_;
  wire _580_;
  wire _581_;
  wire _582_;
  wire _583_;
  wire _584_;
  wire _585_;
  wire _586_;
  wire _587_;
  wire _588_;
  wire _589_;
  wire _590_;
  wire _591_;
  wire _592_;
  wire _593_;
  wire _594_;
  wire _595_;
  wire _596_;
  wire _597_;
  wire _598_;
  wire _599_;
  wire _600_;
  wire _601_;
  wire _602_;
  wire _603_;
  wire _604_;
  wire _605_;
  wire _606_;
  wire _607_;
  wire _608_;
  wire _609_;
  wire _610_;
  wire _611_;
  wire _612_;
  wire _613_;
  wire _614_;
  wire _615_;
  wire _616_;
  wire _617_;
  wire _618_;
  wire _619_;
  wire _620_;
  wire _621_;
  wire _622_;
  wire _623_;
  wire _624_;
  wire _625_;
  wire _626_;
  wire _627_;
  wire _628_;
  wire _629_;
  wire _630_;
  wire _631_;
  wire _632_;
  wire _633_;
  wire _634_;
  wire _635_;
  wire _636_;
  wire _637_;
  wire _638_;
  wire _639_;
  wire _640_;
  wire _641_;
  wire _642_;
  wire _643_;
  wire _644_;
  wire _645_;
  wire _646_;
  wire _647_;
  wire _648_;
  wire _649_;
  wire _650_;
  wire _651_;
  wire _652_;
  wire _653_;
  wire _654_;
  wire _655_;
  wire _656_;
  wire _657_;
  wire _658_;
  wire _659_;
  wire _660_;
  wire _661_;
  wire _662_;
  wire _663_;
  wire _664_;
  wire _665_;
  wire _666_;
  wire _667_;
  wire _668_;
  wire _669_;
  wire _670_;
  wire _671_;
  wire _672_;
  wire _673_;
  wire _674_;
  wire _675_;
  wire _676_;
  wire _677_;
  wire _678_;
  wire _679_;
  wire _680_;
  wire _681_;
  wire _682_;
  wire _683_;
  wire _684_;
  wire _685_;
  wire _686_;
  wire _687_;
  wire _688_;
  wire _689_;
  wire _690_;
  wire _691_;
  wire _692_;
  wire _693_;
  wire _694_;
  wire _695_;
  wire _696_;
  wire _697_;
  wire _698_;
  wire _699_;
  wire _700_;
  wire _701_;
  wire _702_;
  wire _703_;
  wire _704_;
  wire _705_;
  wire _706_;
  wire _707_;
  wire _708_;
  wire _709_;
  wire _710_;
  wire _711_;
  wire _712_;
  wire _713_;
  wire _714_;
  wire _715_;
  wire _716_;
  wire _717_;
  wire _718_;
  wire _719_;
  wire _720_;
  wire _721_;
  wire _722_;
  wire _723_;
  wire _724_;
  wire _725_;
  wire _726_;
  wire _727_;
  wire _728_;
  wire _729_;
  wire _730_;
  wire _731_;
  wire _732_;
  wire _733_;
  wire _734_;
  wire _735_;
  wire _736_;
  wire _737_;
  wire _738_;
  wire _739_;
  wire _740_;
  wire _741_;
  wire _742_;
  wire _743_;
  wire _744_;
  wire _745_;
  wire _746_;
  wire _747_;
  wire _748_;
  wire _749_;
  wire _750_;
  wire _751_;
  wire _752_;
  wire _753_;
  wire _754_;
  wire _755_;
  wire _756_;
  wire _757_;
  wire _758_;
  wire _759_;
  wire _760_;
  wire _761_;
  wire _762_;
  wire _763_;
  wire _764_;
  wire _765_;
  wire _766_;
  wire _767_;
  wire _768_;
  wire _769_;
  wire _770_;
  wire _771_;
  wire _772_;
  wire _773_;
  wire _774_;
  wire _775_;
  wire _776_;
  wire _777_;
  wire _778_;
  wire _779_;
  wire _780_;
  wire _781_;
  wire _782_;
  wire _783_;
  wire _784_;
  wire _785_;
  wire _786_;
  wire _787_;
  wire _788_;
  wire _789_;
  wire _790_;
  wire _791_;
  wire _792_;
  wire _793_;
  wire _794_;
  wire _795_;
  wire _796_;
  wire _797_;
  wire _798_;
  wire _799_;
  wire _800_;
  wire _801_;
  wire _802_;
  wire _803_;
  wire _804_;
  wire _805_;
  wire _806_;
  wire _807_;
  wire _808_;
  wire _809_;
  wire _810_;
  wire _811_;
  wire _812_;
  wire _813_;
  wire _814_;
  wire _815_;
  wire _816_;
  wire _817_;
  wire _818_;
  wire _819_;
  wire _820_;
  wire _821_;
  wire _822_;
  wire _823_;
  wire _824_;
  wire _825_;
  wire _826_;
  wire _827_;
  wire _828_;
  wire _829_;
  wire _830_;
  wire _831_;
  wire _832_;
  wire _833_;
  wire _834_;
  wire _835_;
  wire _836_;
  wire _837_;
  wire _838_;
  wire _839_;
  wire _840_;
  wire _841_;
  wire _842_;
  wire _843_;
  wire _844_;
  wire _845_;
  wire _846_;
  wire _847_;
  wire _848_;
  wire _849_;
  wire _850_;
  wire _851_;
  wire _852_;
  wire _853_;
  wire _854_;
  wire _855_;
  wire _856_;
  wire _857_;
  wire _858_;
  wire _859_;
  wire _860_;
  wire _861_;
  wire _862_;
  wire _863_;
  wire _864_;
  wire _865_;
  wire _866_;
  wire _867_;
  wire _868_;
  wire _869_;
  wire _870_;
  wire _871_;
  wire _872_;
  wire _873_;
  wire _874_;
  wire _875_;
  wire _876_;
  wire _877_;
  wire _878_;
  wire _879_;
  wire _880_;
  wire _881_;
  wire _882_;
  wire _883_;
  wire _884_;
  wire _885_;
  wire _886_;
  wire _887_;
  wire _888_;
  wire _889_;
  wire _890_;
  wire _891_;
  wire _892_;
  wire _893_;
  wire _894_;
  wire _895_;
  wire _896_;
  wire _897_;
  wire _898_;
  wire _899_;
  wire _900_;
  wire _901_;
  wire _902_;
  wire _903_;
  wire _904_;
  wire _905_;
  wire _906_;
  wire _907_;
  wire _908_;
  wire _909_;
  wire _910_;
  wire _911_;
  wire _912_;
  wire _913_;
  wire _914_;
  wire _915_;
  wire _916_;
  wire _917_;
  wire _918_;
  wire _919_;
  wire _920_;
  wire _921_;
  wire _922_;
  wire _923_;
  wire _924_;
  wire _925_;
  wire _926_;
  wire _927_;
  wire _928_;
  wire _929_;
  wire _930_;
  wire _931_;
  wire _932_;
  wire _933_;
  wire _934_;
  wire _935_;
  wire _936_;
  wire _937_;
  wire _938_;
  wire _939_;
  wire _940_;
  wire _941_;
  wire _942_;
  wire _943_;
  wire _944_;
  wire _945_;
  wire _946_;
  wire _947_;
  wire _948_;
  wire _949_;
  wire _950_;
  wire _951_;
  wire _952_;
  wire _953_;
  wire _954_;
  wire _955_;
  wire _956_;
  wire _957_;
  wire _958_;
  wire _959_;
  wire _960_;
  wire _961_;
  wire _962_;
  wire _963_;
  wire _964_;
  wire _965_;
  wire _966_;
  wire _967_;
  wire _968_;
  wire _969_;
  wire _970_;
  wire _971_;
  wire _972_;
  wire _973_;
  wire _974_;
  wire _975_;
  wire _976_;
  wire _977_;
  wire _978_;
  wire _979_;
  wire _980_;
  wire _981_;
  wire _982_;
  wire _983_;
  wire _984_;
  wire _985_;
  wire _986_;
  wire _987_;
  wire _988_;
  wire _989_;
  wire _990_;
  wire _991_;
  wire _992_;
  wire _993_;
  wire _994_;
  wire _995_;
  wire _996_;
  wire _997_;
  wire _998_;
  wire _999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire _1601_;
  wire _1602_;
  wire _1603_;
  wire _1604_;
  wire _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire _1611_;
  wire _1612_;
  wire _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire _1629_;
  wire _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire _1720_;
  wire _1721_;
  wire _1722_;
  wire _1723_;
  wire _1724_;
  wire _1725_;
  wire _1726_;
  wire _1727_;
  wire _1728_;
  wire _1729_;
  wire _1730_;
  wire _1731_;
  wire _1732_;
  wire _1733_;
  wire _1734_;
  wire _1735_;
  wire _1736_;
  wire _1737_;
  wire _1738_;
  wire _1739_;
  wire _1740_;
  wire _1741_;
  wire _1742_;
  wire _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire _1751_;
  wire _1752_;
  wire _1753_;
  wire _1754_;
  wire _1755_;
  wire _1756_;
  wire _1757_;
  wire _1758_;
  wire _1759_;
  wire _1760_;
  wire _1761_;
  wire _1762_;
  wire _1763_;
  wire _1764_;
  wire _1765_;
  wire _1766_;
  wire _1767_;
  wire _1768_;
  wire _1769_;
  wire _1770_;
  wire _1771_;
  wire _1772_;
  wire _1773_;
  wire _1774_;
  wire _1775_;
  wire _1776_;
  wire _1777_;
  wire _1778_;
  wire _1779_;
  wire _1780_;
  wire _1781_;
  wire _1782_;
  wire _1783_;
  wire _1784_;
  wire _1785_;
  wire _1786_;
  wire _1787_;
  wire _1788_;
  wire _1789_;
  wire _1790_;
  wire _1791_;
  wire _1792_;
  wire _1793_;
  wire _1794_;
  wire _1795_;
  wire _1796_;
  wire _1797_;
  wire _1798_;
  wire _1799_;
  wire _1800_;
  wire _1801_;
  wire _1802_;
  wire _1803_;
  wire _1804_;
  wire _1805_;
  wire _1806_;
  wire _1807_;
  wire _1808_;
  wire _1809_;
  wire _1810_;
  wire _1811_;
  wire _1812_;
  wire _1813_;
  wire _1814_;
  wire _1815_;
  wire _1816_;
  wire _1817_;
  wire _1818_;
  wire _1819_;
  wire _1820_;
  wire _1821_;
  wire _1822_;
  wire _1823_;
  wire _1824_;
  wire _1825_;
  wire _1826_;
  wire _1827_;
  wire _1828_;
  wire _1829_;
  wire _1830_;
  wire _1831_;
  wire _1832_;
  wire _1833_;
  wire _1834_;
  wire _1835_;
  wire _1836_;
  wire _1837_;
  wire _1838_;
  wire _1839_;
  wire _1840_;
  wire _1841_;
  wire _1842_;
  wire _1843_;
  wire _1844_;
  wire _1845_;
  wire _1846_;
  wire _1847_;
  wire _1848_;
  wire _1849_;
  wire _1850_;
  wire _1851_;
  wire _1852_;
  wire _1853_;
  wire _1854_;
  wire _1855_;
  wire _1856_;
  wire _1857_;
  wire _1858_;
  wire _1859_;
  wire _1860_;
  wire _1861_;
  wire _1862_;
  wire _1863_;
  wire _1864_;
  wire _1865_;
  wire _1866_;
  wire _1867_;
  wire _1868_;
  wire _1869_;
  wire _1870_;
  wire _1871_;
  wire _1872_;
  wire _1873_;
  wire _1874_;
  wire _1875_;
  wire _1876_;
  wire _1877_;
  wire _1878_;
  wire _1879_;
  wire _1880_;
  wire _1881_;
  wire _1882_;
  wire _1883_;
  wire _1884_;
  wire _1885_;
  wire _1886_;
  wire _1887_;
  wire _1888_;
  wire _1889_;
  wire _1890_;
  wire _1891_;
  wire _1892_;
  wire _1893_;
  wire _1894_;
  wire _1895_;
  wire _1896_;
  wire _1897_;
  wire _1898_;
  wire _1899_;
  wire _1900_;
  wire _1901_;
  wire _1902_;
  wire _1903_;
  wire _1904_;
  wire _1905_;
  wire _1906_;
  wire _1907_;
  wire _1908_;
  wire _1909_;
  wire _1910_;
  wire _1911_;
  wire _1912_;
  wire _1913_;
  wire _1914_;
  wire _1915_;
  wire _1916_;
  wire _1917_;
  wire _1918_;
  wire _1919_;
  wire _1920_;
  wire _1921_;
  wire _1922_;
  wire _1923_;
  wire _1924_;
  wire _1925_;
  wire _1926_;
  wire _1927_;
  wire _1928_;
  wire _1929_;
  wire _1930_;
  wire _1931_;
  wire _1932_;
  wire _1933_;
  wire _1934_;
  wire _1935_;
  wire _1936_;
  wire _1937_;
  wire _1938_;
  wire _1939_;
  wire _1940_;
  wire _1941_;
  wire _1942_;
  wire _1943_;
  wire _1944_;
  wire _1945_;
  wire _1946_;
  wire _1947_;
  wire _1948_;
  wire _1949_;
  wire _1950_;
  wire _1951_;
  wire _1952_;
  wire _1953_;
  wire _1954_;
  wire _1955_;
  wire _1956_;
  wire _1957_;
  wire _1958_;
  wire _1959_;
  wire _1960_;
  wire _1961_;
  wire _1962_;
  wire _1963_;
  wire _1964_;
  wire _1965_;
  wire _1966_;
  wire _1967_;
  wire _1968_;
  wire _1969_;
  wire _1970_;
  wire _1971_;
  wire _1972_;
  wire _1973_;
  wire _1974_;
  wire _1975_;
  wire _1976_;
  wire _1977_;
  wire _1978_;
  wire _1979_;
  wire _1980_;
  wire _1981_;
  wire _1982_;
  wire _1983_;
  wire _1984_;
  wire _1985_;
  wire _1986_;
  wire _1987_;
  wire _1988_;
  wire _1989_;
  wire _1990_;
  wire _1991_;
  wire _1992_;
  wire _1993_;
  wire _1994_;
  wire _1995_;
  wire _1996_;
  wire _1997_;
  wire _1998_;
  wire _1999_;
  wire _2000_;
  wire _2001_;
  wire _2002_;
  wire _2003_;
  wire _2004_;
  wire _2005_;
  wire _2006_;
  wire _2007_;
  wire _2008_;
  wire _2009_;
  wire _2010_;
  wire _2011_;
  wire _2012_;
  wire _2013_;
  wire _2014_;
  wire _2015_;
  wire _2016_;
  wire _2017_;
  wire _2018_;
  wire _2019_;
  wire _2020_;
  wire _2021_;
  wire _2022_;
  wire _2023_;
  wire _2024_;
  wire _2025_;
  wire _2026_;
  wire _2027_;
  wire _2028_;
  wire _2029_;
  wire _2030_;
  wire _2031_;
  wire _2032_;
  wire _2033_;
  wire _2034_;
  wire _2035_;
  wire _2036_;
  wire _2037_;
  wire _2038_;
  wire _2039_;
  wire _2040_;
  wire _2041_;
  wire _2042_;
  wire _2043_;
  wire _2044_;
  wire _2045_;
  wire _2046_;
  wire _2047_;
  wire _2048_;
  wire _2049_;
  wire _2050_;
  wire _2051_;
  wire _2052_;
  wire _2053_;
  wire _2054_;
  wire _2055_;
  wire _2056_;
  wire _2057_;
  wire _2058_;
  wire _2059_;
  wire _2060_;
  wire _2061_;
  wire _2062_;
  wire _2063_;
  wire _2064_;
  wire _2065_;
  wire _2066_;
  wire _2067_;
  wire _2068_;
  wire _2069_;
  wire _2070_;
  wire _2071_;
  wire _2072_;
  wire _2073_;
  wire _2074_;
  wire _2075_;
  wire _2076_;
  wire _2077_;
  wire _2078_;
  wire _2079_;
  wire _2080_;
  wire _2081_;
  wire _2082_;
  wire _2083_;
  wire _2084_;
  wire _2085_;
  wire _2086_;
  wire _2087_;
  wire _2088_;
  wire _2089_;
  wire _2090_;
  wire _2091_;
  wire _2092_;
  wire _2093_;
  wire _2094_;
  wire _2095_;
  wire _2096_;
  wire _2097_;
  wire _2098_;
  wire _2099_;
  wire _2100_;
  wire _2101_;
  wire _2102_;
  wire _2103_;
  wire _2104_;
  wire _2105_;
  wire _2106_;
  wire _2107_;
  wire _2108_;
  wire _2109_;
  wire _2110_;
  wire _2111_;
  wire _2112_;
  wire _2113_;
  wire _2114_;
  wire _2115_;
  wire _2116_;
  wire _2117_;
  wire _2118_;
  wire _2119_;
  wire _2120_;
  wire _2121_;
  wire _2122_;
  wire _2123_;
  wire _2124_;
  wire _2125_;
  wire _2126_;
  wire _2127_;
  wire _2128_;
  wire _2129_;
  wire _2130_;
  wire _2131_;
  wire _2132_;
  wire _2133_;
  wire _2134_;
  wire _2135_;
  wire _2136_;
  wire _2137_;
  wire _2138_;
  wire _2139_;
  wire _2140_;
  wire _2141_;
  wire _2142_;
  wire _2143_;
  wire _2144_;
  wire _2145_;
  wire _2146_;
  wire _2147_;
  wire _2148_;
  wire _2149_;
  wire _2150_;
  wire _2151_;
  wire _2152_;
  wire _2153_;
  wire _2154_;
  wire _2155_;
  wire _2156_;
  wire _2157_;
  wire _2158_;
  wire _2159_;
  wire _2160_;
  wire _2161_;
  wire _2162_;
  wire _2163_;
  wire _2164_;
  wire _2165_;
  wire _2166_;
  wire _2167_;
  wire _2168_;
  wire _2169_;
  wire _2170_;
  wire _2171_;
  wire _2172_;
  wire _2173_;
  wire _2174_;
  wire _2175_;
  wire _2176_;
  wire _2177_;
  wire _2178_;
  wire _2179_;
  wire _2180_;
  wire _2181_;
  wire _2182_;
  wire _2183_;
  wire _2184_;
  wire _2185_;
  wire _2186_;
  wire _2187_;
  wire _2188_;
  wire _2189_;
  wire _2190_;
  wire _2191_;
  wire _2192_;
  wire _2193_;
  wire _2194_;
  wire _2195_;
  wire _2196_;
  wire _2197_;
  wire _2198_;
  wire _2199_;
  wire _2200_;
  wire _2201_;
  wire _2202_;
  wire _2203_;
  wire _2204_;
  wire _2205_;
  wire _2206_;
  wire _2207_;
  wire _2208_;
  wire _2209_;
  wire _2210_;
  wire _2211_;
  wire _2212_;
  wire _2213_;
  wire _2214_;
  wire _2215_;
  wire _2216_;
  wire _2217_;
  wire _2218_;
  wire _2219_;
  wire _2220_;
  wire _2221_;
  wire _2222_;
  wire _2223_;
  wire _2224_;
  wire _2225_;
  wire _2226_;
  wire _2227_;
  wire _2228_;
  wire _2229_;
  wire _2230_;
  wire _2231_;
  wire _2232_;
  wire _2233_;
  wire _2234_;
  wire _2235_;
  wire _2236_;
  wire _2237_;
  wire _2238_;
  wire _2239_;
  wire _2240_;
  wire _2241_;
  wire _2242_;
  wire _2243_;
  wire _2244_;
  wire _2245_;
  wire _2246_;
  wire _2247_;
  wire _2248_;
  wire _2249_;
  wire _2250_;
  wire _2251_;
  wire _2252_;
  wire _2253_;
  wire _2254_;
  wire _2255_;
  wire _2256_;
  wire _2257_;
  wire _2258_;
  wire _2259_;
  wire _2260_;
  wire _2261_;
  wire _2262_;
  wire _2263_;
  wire _2264_;
  wire _2265_;
  wire _2266_;
  wire _2267_;
  wire _2268_;
  wire _2269_;
  wire _2270_;
  wire _2271_;
  wire _2272_;
  wire _2273_;
  wire _2274_;
  wire _2275_;
  wire _2276_;
  wire _2277_;
  wire _2278_;
  wire _2279_;
  wire _2280_;
  wire _2281_;
  wire _2282_;
  wire _2283_;
  wire _2284_;
  wire _2285_;
  wire _2286_;
  wire _2287_;
  wire _2288_;
  wire _2289_;
  wire _2290_;
  wire _2291_;
  wire _2292_;
  wire _2293_;
  wire _2294_;
  wire _2295_;
  wire _2296_;
  wire _2297_;
  wire _2298_;
  wire _2299_;
  wire _2300_;
  wire _2301_;
  wire _2302_;
  wire _2303_;
  wire _2304_;
  wire _2305_;
  wire _2306_;
  wire _2307_;
  wire _2308_;
  wire _2309_;
  wire _2310_;
  wire _2311_;
  wire _2312_;
  wire _2313_;
  wire _2314_;
  wire _2315_;
  wire _2316_;
  wire _2317_;
  wire _2318_;
  wire _2319_;
  wire _2320_;
  wire _2321_;
  wire _2322_;
  wire _2323_;
  wire _2324_;
  wire _2325_;
  wire _2326_;
  wire _2327_;
  wire _2328_;
  wire _2329_;
  wire _2330_;
  wire _2331_;
  wire _2332_;
  wire _2333_;
  wire _2334_;
  wire _2335_;
  wire _2336_;
  wire _2337_;
  wire _2338_;
  wire _2339_;
  wire _2340_;
  wire _2341_;
  wire _2342_;
  wire _2343_;
  wire _2344_;
  wire _2345_;
  wire _2346_;
  wire _2347_;
  wire _2348_;
  wire _2349_;
  wire _2350_;
  wire _2351_;
  wire _2352_;
  wire _2353_;
  wire _2354_;
  wire _2355_;
  wire _2356_;
  wire _2357_;
  wire _2358_;
  wire _2359_;
  wire _2360_;
  wire _2361_;
  wire _2362_;
  wire _2363_;
  wire _2364_;
  wire _2365_;
  wire _2366_;
  wire _2367_;
  wire _2368_;
  wire _2369_;
  wire _2370_;
  wire _2371_;
  wire _2372_;
  wire _2373_;
  wire _2374_;
  wire _2375_;
  wire _2376_;
  wire _2377_;
  wire _2378_;
  wire _2379_;
  wire _2380_;
  wire _2381_;
  wire _2382_;
  wire _2383_;
  wire _2384_;
  wire _2385_;
  wire _2386_;
  wire _2387_;
  wire _2388_;
  wire _2389_;
  wire _2390_;
  wire _2391_;
  wire _2392_;
  wire _2393_;
  wire _2394_;
  wire _2395_;
  wire _2396_;
  wire _2397_;
  wire _2398_;
  wire _2399_;
  wire _2400_;
  wire _2401_;
  wire _2402_;
  wire _2403_;
  wire _2404_;
  wire _2405_;
  wire _2406_;
  wire _2407_;
  wire _2408_;
  wire _2409_;
  wire _2410_;
  wire _2411_;
  wire _2412_;
  wire _2413_;
  wire _2414_;
  wire _2415_;
  wire _2416_;
  wire _2417_;
  wire _2418_;
  wire _2419_;
  wire _2420_;
  wire _2421_;
  wire _2422_;
  wire _2423_;
  wire _2424_;
  wire _2425_;
  wire _2426_;
  wire _2427_;
  wire _2428_;
  wire _2429_;
  wire _2430_;
  wire _2431_;
  wire _2432_;
  wire _2433_;
  wire _2434_;
  wire _2435_;
  wire _2436_;
  wire _2437_;
  wire _2438_;
  wire _2439_;
  wire _2440_;
  wire _2441_;
  wire _2442_;
  wire _2443_;
  wire _2444_;
  wire _2445_;
  wire _2446_;
  wire _2447_;
  wire _2448_;
  wire _2449_;
  wire _2450_;
  wire _2451_;
  wire _2452_;
  wire _2453_;
  wire _2454_;
  wire _2455_;
  wire _2456_;
  wire _2457_;
  wire _2458_;
  wire _2459_;
  wire _2460_;
  wire _2461_;
  wire _2462_;
  wire _2463_;
  wire _2464_;
  wire _2465_;
  wire _2466_;
  wire _2467_;
  wire _2468_;
  wire _2469_;
  wire _2470_;
  wire _2471_;
  wire _2472_;
  wire _2473_;
  wire _2474_;
  wire _2475_;
  wire _2476_;
  wire _2477_;
  wire _2478_;
  wire _2479_;
  wire _2480_;
  wire _2481_;
  wire _2482_;
  wire _2483_;
  wire _2484_;
  wire _2485_;
  wire _2486_;
  wire _2487_;
  wire _2488_;
  wire _2489_;
  wire _2490_;
  wire _2491_;
  wire _2492_;
  wire _2493_;
  wire _2494_;
  wire _2495_;
  wire _2496_;
  wire _2497_;
  wire _2498_;
  wire _2499_;
  wire _2500_;
  wire _2501_;
  wire _2502_;
  wire _2503_;
  wire _2504_;
  wire _2505_;
  wire _2506_;
  wire _2507_;
  wire _2508_;
  wire _2509_;
  wire _2510_;
  wire _2511_;
  wire _2512_;
  wire _2513_;
  wire _2514_;
  wire _2515_;
  wire _2516_;
  wire _2517_;
  wire _2518_;
  wire _2519_;
  wire _2520_;
  wire _2521_;
  wire _2522_;
  wire _2523_;
  wire _2524_;
  wire _2525_;
  wire _2526_;
  wire _2527_;
  wire _2528_;
  wire _2529_;
  wire _2530_;
  wire _2531_;
  wire _2532_;
  wire _2533_;
  wire _2534_;
  wire _2535_;
  wire _2536_;
  wire _2537_;
  wire _2538_;
  wire _2539_;
  wire _2540_;
  wire _2541_;
  wire _2542_;
  wire _2543_;
  wire _2544_;
  wire _2545_;
  wire _2546_;
  wire _2547_;
  wire _2548_;
  wire _2549_;
  wire _2550_;
  wire _2551_;
  wire _2552_;
  wire _2553_;
  wire _2554_;
  wire _2555_;
  wire _2556_;
  wire _2557_;
  wire _2558_;
  wire _2559_;
  wire _2560_;
  wire _2561_;
  wire _2562_;
  wire _2563_;
  wire _2564_;
  wire _2565_;
  wire _2566_;
  wire _2567_;
  wire _2568_;
  wire _2569_;
  wire _2570_;
  wire _2571_;
  wire _2572_;
  wire _2573_;
  wire _2574_;
  wire _2575_;
  wire _2576_;
  wire _2577_;
  wire _2578_;
  wire _2579_;
  wire _2580_;
  wire _2581_;
  wire _2582_;
  wire _2583_;
  wire _2584_;
  wire _2585_;
  wire _2586_;
  wire _2587_;
  wire _2588_;
  wire _2589_;
  wire _2590_;
  wire _2591_;
  wire _2592_;
  wire _2593_;
  wire _2594_;
  wire _2595_;
  wire _2596_;
  wire _2597_;
  wire _2598_;
  wire _2599_;
  wire _2600_;
  wire _2601_;
  wire _2602_;
  wire _2603_;
  wire _2604_;
  wire _2605_;
  wire _2606_;
  wire _2607_;
  wire _2608_;
  wire _2609_;
  wire _2610_;
  wire _2611_;
  wire _2612_;
  wire _2613_;
  wire _2614_;
  wire _2615_;
  wire _2616_;
  wire _2617_;
  wire _2618_;
  wire _2619_;
  wire _2620_;
  wire _2621_;
  wire _2622_;
  wire _2623_;
  wire _2624_;
  wire _2625_;
  wire _2626_;
  wire _2627_;
  wire _2628_;
  wire _2629_;
  wire _2630_;
  wire _2631_;
  wire _2632_;
  wire _2633_;
  wire _2634_;
  wire _2635_;
  wire _2636_;
  wire _2637_;
  wire _2638_;
  wire _2639_;
  wire _2640_;
  wire _2641_;
  wire _2642_;
  wire _2643_;
  wire _2644_;
  wire _2645_;
  wire _2646_;
  wire _2647_;
  wire _2648_;
  wire _2649_;
  wire _2650_;
  wire _2651_;
  wire _2652_;
  wire _2653_;
  wire _2654_;
  wire _2655_;
  wire _2656_;
  wire _2657_;
  wire _2658_;
  wire _2659_;
  wire _2660_;
  wire _2661_;
  wire _2662_;
  wire _2663_;
  wire _2664_;
  wire _2665_;
  wire _2666_;
  wire _2667_;
  wire _2668_;
  wire _2669_;
  wire _2670_;
  wire _2671_;
  wire _2672_;
  wire _2673_;
  wire _2674_;
  wire _2675_;
  wire _2676_;
  wire _2677_;
  wire _2678_;
  wire _2679_;
  wire _2680_;
  wire _2681_;
  wire _2682_;
  wire _2683_;
  wire _2684_;
  wire _2685_;
  wire _2686_;
  wire _2687_;
  wire _2688_;
  wire _2689_;
  wire _2690_;
  wire _2691_;
  wire _2692_;
  wire _2693_;
  wire _2694_;
  wire _2695_;
  wire _2696_;
  wire _2697_;
  wire _2698_;
  wire _2699_;
  wire _2700_;
  wire _2701_;
  wire _2702_;
  wire _2703_;
  wire _2704_;
  wire _2705_;
  wire _2706_;
  wire _2707_;
  wire _2708_;
  wire _2709_;
  wire _2710_;
  wire _2711_;
  wire _2712_;
  wire _2713_;
  wire _2714_;
  wire _2715_;
  wire _2716_;
  wire _2717_;
  wire _2718_;
  wire _2719_;
  wire _2720_;
  wire _2721_;
  wire _2722_;
  wire _2723_;
  wire _2724_;
  wire _2725_;
  wire _2726_;
  wire _2727_;
  wire _2728_;
  wire _2729_;
  wire _2730_;
  wire _2731_;
  wire _2732_;
  wire _2733_;
  wire _2734_;
  wire _2735_;
  wire _2736_;
  wire _2737_;
  wire _2738_;
  wire _2739_;
  wire _2740_;
  wire _2741_;
  wire _2742_;
  wire _2743_;
  wire _2744_;
  wire _2745_;
  wire _2746_;
  wire _2747_;
  wire _2748_;
  wire _2749_;
  wire _2750_;
  wire _2751_;
  wire _2752_;
  wire _2753_;
  wire _2754_;
  wire _2755_;
  wire _2756_;
  wire _2757_;
  wire _2758_;
  wire _2759_;
  wire _2760_;
  wire _2761_;
  wire _2762_;
  wire _2763_;
  wire _2764_;
  wire _2765_;
  wire _2766_;
  wire _2767_;
  wire _2768_;
  wire _2769_;
  wire _2770_;
  wire _2771_;
  wire _2772_;
  wire _2773_;
  wire _2774_;
  wire _2775_;
  wire _2776_;
  wire _2777_;
  wire _2778_;
  wire _2779_;
  wire _2780_;
  wire _2781_;
  wire _2782_;
  wire _2783_;
  wire _2784_;
  wire _2785_;
  wire _2786_;
  wire _2787_;
  wire _2788_;
  wire _2789_;
  wire _2790_;
  wire _2791_;
  wire _2792_;
  wire _2793_;
  wire _2794_;
  wire _2795_;
  wire _2796_;
  wire _2797_;
  wire _2798_;
  wire _2799_;
  wire _2800_;
  wire _2801_;
  wire _2802_;
  wire _2803_;
  wire _2804_;
  wire _2805_;
  wire _2806_;
  wire _2807_;
  wire _2808_;
  wire _2809_;
  wire _2810_;
  wire _2811_;
  wire _2812_;
  wire _2813_;
  wire _2814_;
  wire _2815_;
  wire _2816_;
  wire _2817_;
  wire _2818_;
  wire _2819_;
  wire _2820_;
  wire _2821_;
  wire _2822_;
  wire _2823_;
  wire _2824_;
  wire _2825_;
  wire _2826_;
  wire _2827_;
  wire _2828_;
  wire _2829_;
  wire _2830_;
  wire _2831_;
  wire _2832_;
  wire _2833_;
  wire _2834_;
  wire _2835_;
  wire _2836_;
  wire _2837_;
  wire _2838_;
  wire _2839_;
  wire _2840_;
  wire _2841_;
  wire _2842_;
  wire _2843_;
  wire _2844_;
  wire _2845_;
  wire _2846_;
  wire _2847_;
  wire _2848_;
  wire _2849_;
  wire _2850_;
  wire _2851_;
  wire _2852_;
  wire _2853_;
  wire _2854_;
  wire _2855_;
  wire _2856_;
  wire _2857_;
  wire _2858_;
  wire _2859_;
  wire _2860_;
  wire _2861_;
  wire _2862_;
  wire _2863_;
  wire _2864_;
  wire _2865_;
  wire _2866_;
  wire _2867_;
  wire _2868_;
  wire _2869_;
  wire _2870_;
  wire _2871_;
  wire _2872_;
  wire _2873_;
  wire _2874_;
  wire _2875_;
  wire _2876_;
  wire _2877_;
  wire _2878_;
  wire _2879_;
  wire _2880_;
  wire _2881_;
  wire _2882_;
  wire _2883_;
  wire _2884_;
  wire _2885_;
  wire _2886_;
  wire _2887_;
  wire _2888_;
  wire _2889_;
  wire _2890_;
  wire _2891_;
  wire _2892_;
  wire _2893_;
  wire _2894_;
  wire _2895_;
  wire _2896_;
  wire _2897_;
  wire _2898_;
  wire _2899_;
  wire _2900_;
  wire _2901_;
  wire _2902_;
  wire _2903_;
  wire _2904_;
  wire _2905_;
  wire _2906_;
  wire _2907_;
  wire _2908_;
  wire _2909_;
  wire _2910_;
  wire _2911_;
  wire _2912_;
  wire _2913_;
  wire _2914_;
  wire _2915_;
  wire _2916_;
  wire _2917_;
  wire _2918_;
  wire _2919_;
  wire _2920_;
  wire _2921_;
  wire _2922_;
  wire _2923_;
  wire _2924_;
  wire _2925_;
  wire _2926_;
  wire _2927_;
  wire _2928_;
  wire _2929_;
  wire _2930_;
  wire _2931_;
  wire _2932_;
  wire _2933_;
  wire _2934_;
  wire _2935_;
  wire _2936_;
  wire _2937_;
  wire _2938_;
  wire _2939_;
  wire _2940_;
  wire _2941_;
  wire _2942_;
  wire _2943_;
  wire _2944_;
  wire _2945_;
  wire _2946_;
  wire _2947_;
  wire _2948_;
  wire _2949_;
  wire _2950_;
  wire _2951_;
  wire _2952_;
  wire _2953_;
  wire _2954_;
  wire _2955_;
  wire _2956_;
  wire _2957_;
  wire _2958_;
  wire _2959_;
  wire _2960_;
  wire _2961_;
  wire _2962_;
  wire _2963_;
  wire _2964_;
  wire _2965_;
  wire _2966_;
  wire _2967_;
  wire _2968_;
  wire _2969_;
  wire _2970_;
  wire _2971_;
  wire _2972_;
  wire _2973_;
  wire _2974_;
  wire _2975_;
  wire _2976_;
  wire _2977_;
  wire _2978_;
  wire _2979_;
  wire _2980_;
  wire _2981_;
  wire _2982_;
  wire _2983_;
  wire _2984_;
  wire _2985_;
  wire _2986_;
  wire _2987_;
  wire _2988_;
  wire _2989_;
  wire _2990_;
  wire _2991_;
  wire _2992_;
  wire _2993_;
  wire _2994_;
  wire _2995_;
  wire _2996_;
  wire _2997_;
  wire _2998_;
  wire _2999_;
  wire _3000_;
  wire _3001_;
  wire _3002_;
  wire _3003_;
  wire _3004_;
  wire _3005_;
  wire _3006_;
  wire _3007_;
  wire _3008_;
  wire _3009_;
  wire _3010_;
  wire _3011_;
  wire _3012_;
  wire _3013_;
  wire _3014_;
  wire _3015_;
  wire _3016_;
  wire _3017_;
  wire _3018_;
  wire _3019_;
  wire _3020_;
  wire _3021_;
  wire _3022_;
  wire _3023_;
  wire _3024_;
  wire _3025_;
  wire _3026_;
  wire _3027_;
  wire _3028_;
  wire _3029_;
  wire _3030_;
  wire _3031_;
  wire _3032_;
  wire _3033_;
  wire _3034_;
  wire _3035_;
  wire _3036_;
  wire _3037_;
  wire _3038_;
  wire _3039_;
  wire _3040_;
  wire _3041_;
  wire _3042_;
  wire _3043_;
  wire _3044_;
  wire _3045_;
  wire _3046_;
  wire _3047_;
  wire _3048_;
  wire _3049_;
  wire _3050_;
  wire _3051_;
  wire _3052_;
  wire _3053_;
  wire _3054_;
  wire _3055_;
  wire _3056_;
  wire _3057_;
  wire _3058_;
  wire _3059_;
  wire _3060_;
  wire _3061_;
  wire _3062_;
  wire _3063_;
  wire _3064_;
  wire _3065_;
  wire _3066_;
  wire _3067_;
  wire _3068_;
  wire _3069_;
  wire _3070_;
  wire _3071_;
  wire _3072_;
  wire _3073_;
  wire _3074_;
  wire _3075_;
  wire _3076_;
  wire _3077_;
  wire _3078_;
  wire _3079_;
  wire _3080_;
  wire _3081_;
  wire _3082_;
  wire _3083_;
  wire _3084_;
  wire _3085_;
  wire _3086_;
  wire _3087_;
  wire _3088_;
  wire _3089_;
  wire _3090_;
  wire _3091_;
  wire _3092_;
  wire _3093_;
  wire _3094_;
  wire _3095_;
  wire _3096_;
  wire _3097_;
  wire _3098_;
  wire _3099_;
  wire _3100_;
  wire _3101_;
  wire _3102_;
  wire _3103_;
  wire _3104_;
  wire _3105_;
  wire _3106_;
  wire _3107_;
  wire _3108_;
  wire _3109_;
  wire _3110_;
  wire _3111_;
  wire _3112_;
  wire _3113_;
  wire _3114_;
  wire _3115_;
  wire _3116_;
  wire _3117_;
  wire _3118_;
  wire _3119_;
  wire _3120_;
  wire _3121_;
  wire _3122_;
  wire _3123_;
  wire _3124_;
  wire _3125_;
  wire _3126_;
  wire _3127_;
  wire _3128_;
  wire _3129_;
  wire _3130_;
  wire _3131_;
  wire _3132_;
  wire _3133_;
  wire _3134_;
  wire _3135_;
  wire _3136_;
  wire _3137_;
  wire _3138_;
  wire _3139_;
  wire _3140_;
  wire _3141_;
  wire _3142_;
  wire _3143_;
  wire _3144_;
  wire _3145_;
  wire _3146_;
  wire _3147_;
  wire _3148_;
  wire _3149_;
  wire _3150_;
  wire _3151_;
  wire _3152_;
  wire _3153_;
  wire _3154_;
  wire _3155_;
  wire _3156_;
  wire _3157_;
  wire _3158_;
  wire _3159_;
  wire _3160_;
  wire _3161_;
  wire _3162_;
  wire _3163_;
  wire _3164_;
  wire _3165_;
  wire _3166_;
  wire _3167_;
  wire _3168_;
  wire _3169_;
  wire _3170_;
  wire _3171_;
  wire _3172_;
  wire _3173_;
  wire _3174_;
  wire _3175_;
  wire _3176_;
  wire _3177_;
  wire _3178_;
  wire _3179_;
  wire _3180_;
  wire _3181_;
  wire _3182_;
  wire _3183_;
  wire _3184_;
  wire _3185_;
  wire _3186_;
  wire _3187_;
  wire _3188_;
  wire _3189_;
  wire _3190_;
  wire _3191_;
  wire _3192_;
  wire _3193_;
  wire _3194_;
  wire _3195_;
  wire _3196_;
  wire _3197_;
  wire _3198_;
  wire _3199_;
  wire _3200_;
  wire _3201_;
  wire _3202_;
  wire _3203_;
  wire _3204_;
  wire _3205_;
  wire _3206_;
  wire _3207_;
  wire _3208_;
  wire _3209_;
  wire _3210_;
  wire _3211_;
  wire _3212_;
  wire _3213_;
  wire _3214_;
  wire _3215_;
  wire _3216_;
  wire _3217_;
  wire _3218_;
  wire _3219_;
  wire _3220_;
  wire _3221_;
  wire _3222_;
  wire _3223_;
  wire _3224_;
  wire _3225_;
  wire _3226_;
  wire _3227_;
  wire _3228_;
  wire _3229_;
  wire _3230_;
  wire _3231_;
  wire _3232_;
  wire _3233_;
  wire _3234_;
  wire _3235_;
  wire _3236_;
  wire _3237_;
  wire _3238_;
  wire _3239_;
  wire _3240_;
  wire _3241_;
  wire _3242_;
  wire _3243_;
  wire _3244_;
  wire _3245_;
  wire _3246_;
  wire _3247_;
  wire _3248_;
  wire _3249_;
  wire _3250_;
  wire _3251_;
  wire _3252_;
  wire _3253_;
  wire _3254_;
  wire _3255_;
  wire _3256_;
  wire _3257_;
  wire _3258_;
  wire _3259_;
  wire _3260_;
  wire _3261_;
  wire _3262_;
  wire _3263_;
  wire _3264_;
  wire _3265_;
  wire _3266_;
  wire _3267_;
  wire _3268_;
  wire _3269_;
  wire _3270_;
  wire _3271_;
  wire _3272_;
  wire _3273_;
  wire _3274_;
  wire _3275_;
  wire _3276_;
  wire _3277_;
  wire _3278_;
  wire _3279_;
  wire _3280_;
  wire _3281_;
  wire _3282_;
  wire _3283_;
  wire _3284_;
  wire _3285_;
  wire _3286_;
  wire _3287_;
  wire _3288_;
  wire _3289_;
  wire _3290_;
  wire _3291_;
  wire _3292_;
  wire _3293_;
  wire _3294_;
  wire _3295_;
  wire _3296_;
  wire _3297_;
  wire _3298_;
  wire _3299_;
  wire _3300_;
  wire _3301_;
  wire _3302_;
  wire _3303_;
  wire _3304_;
  wire _3305_;
  wire _3306_;
  wire _3307_;
  wire _3308_;
  wire _3309_;
  wire _3310_;
  wire _3311_;
  wire _3312_;
  wire _3313_;
  wire _3314_;
  wire _3315_;
  wire _3316_;
  wire _3317_;
  wire _3318_;
  wire _3319_;
  wire _3320_;
  wire _3321_;
  wire _3322_;
  wire _3323_;
  wire _3324_;
  wire _3325_;
  wire _3326_;
  wire _3327_;
  wire _3328_;
  wire _3329_;
  wire _3330_;
  wire _3331_;
  wire _3332_;
  wire _3333_;
  wire _3334_;
  wire _3335_;
  wire _3336_;
  wire _3337_;
  wire _3338_;
  wire _3339_;
  wire _3340_;
  wire _3341_;
  wire _3342_;
  wire _3343_;
  wire _3344_;
  wire _3345_;
  wire _3346_;
  wire _3347_;
  wire _3348_;
  wire _3349_;
  wire _3350_;
  wire _3351_;
  wire _3352_;
  wire _3353_;
  wire _3354_;
  wire _3355_;
  wire _3356_;
  wire _3357_;
  wire _3358_;
  wire _3359_;
  wire _3360_;
  wire _3361_;
  wire _3362_;
  wire _3363_;
  wire _3364_;
  wire _3365_;
  wire _3366_;
  wire _3367_;
  wire _3368_;
  wire _3369_;
  wire _3370_;
  wire _3371_;
  wire _3372_;
  wire _3373_;
  wire _3374_;
  wire _3375_;
  wire _3376_;
  wire _3377_;
  wire _3378_;
  wire _3379_;
  wire _3380_;
  wire _3381_;
  wire _3382_;
  wire _3383_;
  wire _3384_;
  wire _3385_;
  wire _3386_;
  wire _3387_;
  wire _3388_;
  wire _3389_;
  wire _3390_;
  wire _3391_;
  wire _3392_;
  wire _3393_;
  wire _3394_;
  wire _3395_;
  wire _3396_;
  wire _3397_;
  wire _3398_;
  wire _3399_;
  wire _3400_;
  wire _3401_;
  wire _3402_;
  wire _3403_;
  wire _3404_;
  wire _3405_;
  wire _3406_;
  wire _3407_;
  wire _3408_;
  wire _3409_;
  wire _3410_;
  wire _3411_;
  wire _3412_;
  wire _3413_;
  wire _3414_;
  wire _3415_;
  wire _3416_;
  wire _3417_;
  wire _3418_;
  wire _3419_;
  wire _3420_;
  wire _3421_;
  wire _3422_;
  wire _3423_;
  wire _3424_;
  wire _3425_;
  wire _3426_;
  wire _3427_;
  wire _3428_;
  wire _3429_;
  wire _3430_;
  wire _3431_;
  wire _3432_;
  wire _3433_;
  wire _3434_;
  wire _3435_;
  wire _3436_;
  wire _3437_;
  wire _3438_;
  wire _3439_;
  wire _3440_;
  wire _3441_;
  wire _3442_;
  wire _3443_;
  wire _3444_;
  wire _3445_;
  wire _3446_;
  wire _3447_;
  wire _3448_;
  wire _3449_;
  wire _3450_;
  wire _3451_;
  wire _3452_;
  wire _3453_;
  wire _3454_;
  wire _3455_;
  wire _3456_;
  wire _3457_;
  wire _3458_;
  wire _3459_;
  wire _3460_;
  wire _3461_;
  wire _3462_;
  wire _3463_;
  wire _3464_;
  wire _3465_;
  wire _3466_;
  wire _3467_;
  wire _3468_;
  wire _3469_;
  wire _3470_;
  wire _3471_;
  wire _3472_;
  wire _3473_;
  wire _3474_;
  wire _3475_;
  wire _3476_;
  wire _3477_;
  wire _3478_;
  wire _3479_;
  wire _3480_;
  wire _3481_;
  wire _3482_;
  wire _3483_;
  wire _3484_;
  wire _3485_;
  wire _3486_;
  wire _3487_;
  wire _3488_;
  wire _3489_;
  wire _3490_;
  wire _3491_;
  wire _3492_;
  wire _3493_;
  wire _3494_;
  wire _3495_;
  wire _3496_;
  wire _3497_;
  wire _3498_;
  wire _3499_;
  wire _3500_;
  wire _3501_;
  wire _3502_;
  wire _3503_;
  wire _3504_;
  wire _3505_;
  wire _3506_;
  wire _3507_;
  wire _3508_;
  wire _3509_;
  wire _3510_;
  wire _3511_;
  wire _3512_;
  wire _3513_;
  wire _3514_;
  wire _3515_;
  wire _3516_;
  wire _3517_;
  wire _3518_;
  wire _3519_;
  wire _3520_;
  wire _3521_;
  wire _3522_;
  wire _3523_;
  wire _3524_;
  wire _3525_;
  wire _3526_;
  wire _3527_;
  wire _3528_;
  wire _3529_;
  wire _3530_;
  wire _3531_;
  wire _3532_;
  wire _3533_;
  wire _3534_;
  wire _3535_;
  wire _3536_;
  wire _3537_;
  wire _3538_;
  wire _3539_;
  wire _3540_;
  wire _3541_;
  wire _3542_;
  wire _3543_;
  wire _3544_;
  wire _3545_;
  wire _3546_;
  wire _3547_;
  wire _3548_;
  wire _3549_;
  wire _3550_;
  wire _3551_;
  wire _3552_;
  wire _3553_;
  wire _3554_;
  wire _3555_;
  wire _3556_;
  wire _3557_;
  wire _3558_;
  wire _3559_;
  wire _3560_;
  wire _3561_;
  wire _3562_;
  wire _3563_;
  wire _3564_;
  wire _3565_;
  wire _3566_;
  wire _3567_;
  wire _3568_;
  wire _3569_;
  wire _3570_;
  wire _3571_;
  wire _3572_;
  wire _3573_;
  wire _3574_;
  wire _3575_;
  wire _3576_;
  wire _3577_;
  wire _3578_;
  wire _3579_;
  wire _3580_;
  wire _3581_;
  wire _3582_;
  wire _3583_;
  wire _3584_;
  wire _3585_;
  wire _3586_;
  wire _3587_;
  wire _3588_;
  wire _3589_;
  wire _3590_;
  wire _3591_;
  wire _3592_;
  wire _3593_;
  wire _3594_;
  wire _3595_;
  wire _3596_;
  wire _3597_;
  wire _3598_;
  wire _3599_;
  wire _3600_;
  wire _3601_;
  wire _3602_;
  wire _3603_;
  wire _3604_;
  wire _3605_;
  wire _3606_;
  wire _3607_;
  wire _3608_;
  wire _3609_;
  wire _3610_;
  wire _3611_;
  wire _3612_;
  wire _3613_;
  wire _3614_;
  wire _3615_;
  wire _3616_;
  wire _3617_;
  wire _3618_;
  wire _3619_;
  wire _3620_;
  wire _3621_;
  wire _3622_;
  wire _3623_;
  wire _3624_;
  wire _3625_;
  wire _3626_;
  wire _3627_;
  wire _3628_;
  wire _3629_;
  wire _3630_;
  wire _3631_;
  wire _3632_;
  wire _3633_;
  wire _3634_;
  wire _3635_;
  wire _3636_;
  wire _3637_;
  wire _3638_;
  wire _3639_;
  wire _3640_;
  wire _3641_;
  wire _3642_;
  wire _3643_;
  wire _3644_;
  wire _3645_;
  wire _3646_;
  wire _3647_;
  wire _3648_;
  wire _3649_;
  wire _3650_;
  wire _3651_;
  wire _3652_;
  wire _3653_;
  wire _3654_;
  wire _3655_;
  wire _3656_;
  wire _3657_;
  wire _3658_;
  wire _3659_;
  wire _3660_;
  wire _3661_;
  wire _3662_;
  wire _3663_;
  wire _3664_;
  wire _3665_;
  wire _3666_;
  wire _3667_;
  wire _3668_;
  wire _3669_;
  wire _3670_;
  wire _3671_;
  wire _3672_;
  wire _3673_;
  wire _3674_;
  wire _3675_;
  wire _3676_;
  wire _3677_;
  wire _3678_;
  wire _3679_;
  wire _3680_;
  wire _3681_;
  wire _3682_;
  wire _3683_;
  wire _3684_;
  wire _3685_;
  wire _3686_;
  wire _3687_;
  wire _3688_;
  wire _3689_;
  wire _3690_;
  wire _3691_;
  wire _3692_;
  wire _3693_;
  wire _3694_;
  wire _3695_;
  wire _3696_;
  wire _3697_;
  wire _3698_;
  wire _3699_;
  wire _3700_;
  wire _3701_;
  wire _3702_;
  wire _3703_;
  wire _3704_;
  wire _3705_;
  wire _3706_;
  wire _3707_;
  wire _3708_;
  wire _3709_;
  wire _3710_;
  wire _3711_;
  wire _3712_;
  wire _3713_;
  wire _3714_;
  wire _3715_;
  wire _3716_;
  wire _3717_;
  wire _3718_;
  wire _3719_;
  wire _3720_;
  wire _3721_;
  wire _3722_;
  wire _3723_;
  wire _3724_;
  wire _3725_;
  wire _3726_;
  wire _3727_;
  wire _3728_;
  wire _3729_;
  wire _3730_;
  wire _3731_;
  wire _3732_;
  wire _3733_;
  wire _3734_;
  wire _3735_;
  wire _3736_;
  wire _3737_;
  wire _3738_;
  wire _3739_;
  wire _3740_;
  wire _3741_;
  wire _3742_;
  wire _3743_;
  wire _3744_;
  wire _3745_;
  wire _3746_;
  wire _3747_;
  wire _3748_;
  wire _3749_;
  wire _3750_;
  wire _3751_;
  wire _3752_;
  wire _3753_;
  wire _3754_;
  wire _3755_;
  wire _3756_;
  wire _3757_;
  wire _3758_;
  wire _3759_;
  wire _3760_;
  wire _3761_;
  wire _3762_;
  wire _3763_;
  wire _3764_;
  wire _3765_;
  wire _3766_;
  wire _3767_;
  wire _3768_;
  wire _3769_;
  wire _3770_;
  wire _3771_;
  wire _3772_;
  wire _3773_;
  wire _3774_;
  wire _3775_;
  wire _3776_;
  wire _3777_;
  wire _3778_;
  wire _3779_;
  wire _3780_;
  wire _3781_;
  wire _3782_;
  wire _3783_;
  wire _3784_;
  wire _3785_;
  wire _3786_;
  wire _3787_;
  wire _3788_;
  wire _3789_;
  wire _3790_;
  wire _3791_;
  wire _3792_;
  wire _3793_;
  wire _3794_;
  wire _3795_;
  wire _3796_;
  wire _3797_;
  wire _3798_;
  wire _3799_;
  wire _3800_;
  wire _3801_;
  wire _3802_;
  wire _3803_;
  wire _3804_;
  wire _3805_;
  wire _3806_;
  wire _3807_;
  wire _3808_;
  wire _3809_;
  wire _3810_;
  wire _3811_;
  wire _3812_;
  wire _3813_;
  wire _3814_;
  wire _3815_;
  wire _3816_;
  wire _3817_;
  wire _3818_;
  wire _3819_;
  wire _3820_;
  wire _3821_;
  wire _3822_;
  wire _3823_;
  wire _3824_;
  wire _3825_;
  wire _3826_;
  wire _3827_;
  wire _3828_;
  wire _3829_;
  wire _3830_;
  wire _3831_;
  wire _3832_;
  wire _3833_;
  wire _3834_;
  wire _3835_;
  wire _3836_;
  wire _3837_;
  wire _3838_;
  wire _3839_;
  wire _3840_;
  wire _3841_;
  wire _3842_;
  wire _3843_;
  wire _3844_;
  wire _3845_;
  wire _3846_;
  wire _3847_;
  wire _3848_;
  wire _3849_;
  wire _3850_;
  wire _3851_;
  wire _3852_;
  wire _3853_;
  wire _3854_;
  wire _3855_;
  wire _3856_;
  wire _3857_;
  wire _3858_;
  wire _3859_;
  wire _3860_;
  wire _3861_;
  wire _3862_;
  wire _3863_;
  wire _3864_;
  wire _3865_;
  wire _3866_;
  wire _3867_;
  wire _3868_;
  wire _3869_;
  wire _3870_;
  wire _3871_;
  wire _3872_;
  wire _3873_;
  wire _3874_;
  wire _3875_;
  wire _3876_;
  wire _3877_;
  wire _3878_;
  wire _3879_;
  wire _3880_;
  wire _3881_;
  wire _3882_;
  wire _3883_;
  wire _3884_;
  wire _3885_;
  wire _3886_;
  wire _3887_;
  wire _3888_;
  wire _3889_;
  wire _3890_;
  wire _3891_;
  wire _3892_;
  wire _3893_;
  wire _3894_;
  wire _3895_;
  wire _3896_;
  wire _3897_;
  wire _3898_;
  wire _3899_;
  wire _3900_;
  wire _3901_;
  wire _3902_;
  wire _3903_;
  wire _3904_;
  wire _3905_;
  wire _3906_;
  wire _3907_;
  wire _3908_;
  wire _3909_;
  wire _3910_;
  wire _3911_;
  wire _3912_;
  wire _3913_;
  wire _3914_;
  wire _3915_;
  wire _3916_;
  wire _3917_;
  wire _3918_;
  wire _3919_;
  wire _3920_;
  wire _3921_;
  wire _3922_;
  wire _3923_;
  wire _3924_;
  wire _3925_;
  wire _3926_;
  wire _3927_;
  wire _3928_;
  wire _3929_;
  wire _3930_;
  wire _3931_;
  wire _3932_;
  wire _3933_;
  wire _3934_;
  wire _3935_;
  wire _3936_;
  wire _3937_;
  wire _3938_;
  wire _3939_;
  wire _3940_;
  wire _3941_;
  wire _3942_;
  wire _3943_;
  wire _3944_;
  wire _3945_;
  wire _3946_;
  wire _3947_;
  wire _3948_;
  wire _3949_;
  wire _3950_;
  wire _3951_;
  wire _3952_;
  wire _3953_;
  wire _3954_;
  wire _3955_;
  wire _3956_;
  wire _3957_;
  wire _3958_;
  wire _3959_;
  wire _3960_;
  wire _3961_;
  wire _3962_;
  wire _3963_;
  wire _3964_;
  wire _3965_;
  wire _3966_;
  wire _3967_;
  wire _3968_;
  wire _3969_;
  wire _3970_;
  wire _3971_;
  wire _3972_;
  wire _3973_;
  wire _3974_;
  wire _3975_;
  wire _3976_;
  wire _3977_;
  wire _3978_;
  wire _3979_;
  wire _3980_;
  wire _3981_;
  wire _3982_;
  wire _3983_;
  wire _3984_;
  wire _3985_;
  wire _3986_;
  wire _3987_;
  wire _3988_;
  wire _3989_;
  wire _3990_;
  wire _3991_;
  wire _3992_;
  wire _3993_;
  wire _3994_;
  wire _3995_;
  wire _3996_;
  wire _3997_;
  wire _3998_;
  wire _3999_;
  wire _4000_;
  wire _4001_;
  wire _4002_;
  wire _4003_;
  wire _4004_;
  wire _4005_;
  wire _4006_;
  wire _4007_;
  wire _4008_;
  wire _4009_;
  wire _4010_;
  wire _4011_;
  wire _4012_;
  wire _4013_;
  wire _4014_;
  wire _4015_;
  wire _4016_;
  wire _4017_;
  wire _4018_;
  wire _4019_;
  wire _4020_;
  wire _4021_;
  wire _4022_;
  wire _4023_;
  wire _4024_;
  wire _4025_;
  wire _4026_;
  wire _4027_;
  wire _4028_;
  wire _4029_;
  wire _4030_;
  wire _4031_;
  wire _4032_;
  wire _4033_;
  wire _4034_;
  wire _4035_;
  wire _4036_;
  wire _4037_;
  wire _4038_;
  wire _4039_;
  wire _4040_;
  wire _4041_;
  wire _4042_;
  wire _4043_;
  wire _4044_;
  wire _4045_;
  wire _4046_;
  wire _4047_;
  wire _4048_;
  wire _4049_;
  wire _4050_;
  wire _4051_;
  wire _4052_;
  wire _4053_;
  wire _4054_;
  wire _4055_;
  wire _4056_;
  wire _4057_;
  wire _4058_;
  wire _4059_;
  wire _4060_;
  wire _4061_;
  wire _4062_;
  wire _4063_;
  wire _4064_;
  wire _4065_;
  wire _4066_;
  wire _4067_;
  wire _4068_;
  wire _4069_;
  wire _4070_;
  wire _4071_;
  wire _4072_;
  wire _4073_;
  wire _4074_;
  wire _4075_;
  wire _4076_;
  wire _4077_;
  wire _4078_;
  wire _4079_;
  wire _4080_;
  wire _4081_;
  wire _4082_;
  wire _4083_;
  wire _4084_;
  wire _4085_;
  wire _4086_;
  wire _4087_;
  wire _4088_;
  wire _4089_;
  wire _4090_;
  wire _4091_;
  wire _4092_;
  wire _4093_;
  wire _4094_;
  wire _4095_;
  wire _4096_;
  wire _4097_;
  wire _4098_;
  wire _4099_;
  wire _4100_;
  wire _4101_;
  wire _4102_;
  wire _4103_;
  wire _4104_;
  wire _4105_;
  wire _4106_;
  wire _4107_;
  wire _4108_;
  wire _4109_;
  wire _4110_;
  wire _4111_;
  wire _4112_;
  wire _4113_;
  wire _4114_;
  wire _4115_;
  wire _4116_;
  wire _4117_;
  wire _4118_;
  wire _4119_;
  wire _4120_;
  wire _4121_;
  wire _4122_;
  wire _4123_;
  wire _4124_;
  wire _4125_;
  wire _4126_;
  wire _4127_;
  wire _4128_;
  wire _4129_;
  wire _4130_;
  wire _4131_;
  wire _4132_;
  wire _4133_;
  wire _4134_;
  wire _4135_;
  wire _4136_;
  wire _4137_;
  wire _4138_;
  wire _4139_;
  wire _4140_;
  wire _4141_;
  wire _4142_;
  wire _4143_;
  wire _4144_;
  wire _4145_;
  wire _4146_;
  wire _4147_;
  wire _4148_;
  wire _4149_;
  wire _4150_;
  wire _4151_;
  wire _4152_;
  wire _4153_;
  wire _4154_;
  wire _4155_;
  wire _4156_;
  wire _4157_;
  wire _4158_;
  wire _4159_;
  wire _4160_;
  wire _4161_;
  wire _4162_;
  wire _4163_;
  wire _4164_;
  wire _4165_;
  wire _4166_;
  wire _4167_;
  wire _4168_;
  wire _4169_;
  wire _4170_;
  wire _4171_;
  wire _4172_;
  wire _4173_;
  wire _4174_;
  wire _4175_;
  wire _4176_;
  wire _4177_;
  wire _4178_;
  wire _4179_;
  wire _4180_;
  wire _4181_;
  wire _4182_;
  wire _4183_;
  wire _4184_;
  wire _4185_;
  wire _4186_;
  wire _4187_;
  wire _4188_;
  wire _4189_;
  wire _4190_;
  wire _4191_;
  wire _4192_;
  wire _4193_;
  wire _4194_;
  wire _4195_;
  wire _4196_;
  wire _4197_;
  wire _4198_;
  wire _4199_;
  wire _4200_;
  wire _4201_;
  wire _4202_;
  wire _4203_;
  wire _4204_;
  wire _4205_;
  wire _4206_;
  wire _4207_;
  wire _4208_;
  wire _4209_;
  wire _4210_;
  wire _4211_;
  wire _4212_;
  wire _4213_;
  wire _4214_;
  wire _4215_;
  wire _4216_;
  wire _4217_;
  wire _4218_;
  wire _4219_;
  wire _4220_;
  wire _4221_;
  wire _4222_;
  wire _4223_;
  wire _4224_;
  wire _4225_;
  wire _4226_;
  wire _4227_;
  wire _4228_;
  wire _4229_;
  wire _4230_;
  wire _4231_;
  wire _4232_;
  wire _4233_;
  wire _4234_;
  wire _4235_;
  wire _4236_;
  wire _4237_;
  wire _4238_;
  wire _4239_;
  wire _4240_;
  wire _4241_;
  wire _4242_;
  wire _4243_;
  wire _4244_;
  wire _4245_;
  wire _4246_;
  wire _4247_;
  wire _4248_;
  wire _4249_;
  wire _4250_;
  wire _4251_;
  wire _4252_;
  wire _4253_;
  wire _4254_;
  wire _4255_;
  wire _4256_;
  wire _4257_;
  wire _4258_;
  wire _4259_;
  wire _4260_;
  wire _4261_;
  wire _4262_;
  wire _4263_;
  wire _4264_;
  wire _4265_;
  wire _4266_;
  wire _4267_;
  wire _4268_;
  wire _4269_;
  wire _4270_;
  wire _4271_;
  wire _4272_;
  wire _4273_;
  wire _4274_;
  wire _4275_;
  wire _4276_;
  wire _4277_;
  wire _4278_;
  wire _4279_;
  wire _4280_;
  wire _4281_;
  wire _4282_;
  wire _4283_;
  wire _4284_;
  wire _4285_;
  wire _4286_;
  wire _4287_;
  wire _4288_;
  wire _4289_;
  wire _4290_;
  wire _4291_;
  wire _4292_;
  wire _4293_;
  wire _4294_;
  wire _4295_;
  wire _4296_;
  wire _4297_;
  wire _4298_;
  wire _4299_;
  wire _4300_;
  wire _4301_;
  wire _4302_;
  wire _4303_;
  wire _4304_;
  wire _4305_;
  wire _4306_;
  wire _4307_;
  wire _4308_;
  wire _4309_;
  wire _4310_;
  wire _4311_;
  wire _4312_;
  wire _4313_;
  wire _4314_;
  wire _4315_;
  wire _4316_;
  wire _4317_;
  wire _4318_;
  wire _4319_;
  wire _4320_;
  wire _4321_;
  wire _4322_;
  wire _4323_;
  wire _4324_;
  wire _4325_;
  wire _4326_;
  wire _4327_;
  wire _4328_;
  wire _4329_;
  wire _4330_;
  wire _4331_;
  wire _4332_;
  wire _4333_;
  wire _4334_;
  wire _4335_;
  wire _4336_;
  wire _4337_;
  wire _4338_;
  wire _4339_;
  wire _4340_;
  wire _4341_;
  wire _4342_;
  wire _4343_;
  wire _4344_;
  wire _4345_;
  wire _4346_;
  wire _4347_;
  wire _4348_;
  wire _4349_;
  wire _4350_;
  wire _4351_;
  wire _4352_;
  wire _4353_;
  wire _4354_;
  wire _4355_;
  wire _4356_;
  wire _4357_;
  wire _4358_;
  wire _4359_;
  wire _4360_;
  wire _4361_;
  wire _4362_;
  wire _4363_;
  wire _4364_;
  wire _4365_;
  wire _4366_;
  wire _4367_;
  wire _4368_;
  wire _4369_;
  wire _4370_;
  wire _4371_;
  wire _4372_;
  wire _4373_;
  wire _4374_;
  wire _4375_;
  wire _4376_;
  wire _4377_;
  wire _4378_;
  wire _4379_;
  wire _4380_;
  wire _4381_;
  wire _4382_;
  wire _4383_;
  wire _4384_;
  wire _4385_;
  wire _4386_;
  wire _4387_;
  wire _4388_;
  wire _4389_;
  wire _4390_;
  wire _4391_;
  wire _4392_;
  wire _4393_;
  wire _4394_;
  wire _4395_;
  wire _4396_;
  wire _4397_;
  wire _4398_;
  wire _4399_;
  wire _4400_;
  wire _4401_;
  wire _4402_;
  wire _4403_;
  wire _4404_;
  wire _4405_;
  wire _4406_;
  wire _4407_;
  wire _4408_;
  wire _4409_;
  wire _4410_;
  wire _4411_;
  wire _4412_;
  wire _4413_;
  wire _4414_;
  wire _4415_;
  wire _4416_;
  wire _4417_;
  wire _4418_;
  wire _4419_;
  wire _4420_;
  wire _4421_;
  wire _4422_;
  wire _4423_;
  wire _4424_;
  wire _4425_;
  wire _4426_;
  wire _4427_;
  wire _4428_;
  wire _4429_;
  wire _4430_;
  wire _4431_;
  wire _4432_;
  wire _4433_;
  wire _4434_;
  wire _4435_;
  wire _4436_;
  wire _4437_;
  wire _4438_;
  wire _4439_;
  wire _4440_;
  wire _4441_;
  wire _4442_;
  wire _4443_;
  wire _4444_;
  wire _4445_;
  wire _4446_;
  wire _4447_;
  wire _4448_;
  wire _4449_;
  wire _4450_;
  wire _4451_;
  wire _4452_;
  wire _4453_;
  wire _4454_;
  wire _4455_;
  wire _4456_;
  wire _4457_;
  wire _4458_;
  wire _4459_;
  wire _4460_;
  wire _4461_;
  wire _4462_;
  wire _4463_;
  wire _4464_;
  wire _4465_;
  wire _4466_;
  wire _4467_;
  wire _4468_;
  wire _4469_;
  wire _4470_;
  wire _4471_;
  wire _4472_;
  wire _4473_;
  wire _4474_;
  wire _4475_;
  wire _4476_;
  wire _4477_;
  wire _4478_;
  wire _4479_;
  wire _4480_;
  wire _4481_;
  wire _4482_;
  wire _4483_;
  wire _4484_;
  wire _4485_;
  wire _4486_;
  wire _4487_;
  wire _4488_;
  wire _4489_;
  wire _4490_;
  wire _4491_;
  wire _4492_;
  wire _4493_;
  wire _4494_;
  wire _4495_;
  wire _4496_;
  wire _4497_;
  wire _4498_;
  wire _4499_;
  wire _4500_;
  wire _4501_;
  wire _4502_;
  wire _4503_;
  wire _4504_;
  wire _4505_;
  wire _4506_;
  wire _4507_;
  wire _4508_;
  wire _4509_;
  wire _4510_;
  wire _4511_;
  wire _4512_;
  wire _4513_;
  wire _4514_;
  wire _4515_;
  wire _4516_;
  wire _4517_;
  wire _4518_;
  wire _4519_;
  wire _4520_;
  wire _4521_;
  wire _4522_;
  wire _4523_;
  wire _4524_;
  wire _4525_;
  wire _4526_;
  wire _4527_;
  wire _4528_;
  wire _4529_;
  wire _4530_;
  wire _4531_;
  wire _4532_;
  wire _4533_;
  wire _4534_;
  wire _4535_;
  wire _4536_;
  wire _4537_;
  wire _4538_;
  wire _4539_;
  wire _4540_;
  wire _4541_;
  wire _4542_;
  wire _4543_;
  wire _4544_;
  wire _4545_;
  wire _4546_;
  wire _4547_;
  wire _4548_;
  wire _4549_;
  wire _4550_;
  wire _4551_;
  wire _4552_;
  wire _4553_;
  wire _4554_;
  wire _4555_;
  wire _4556_;
  wire _4557_;
  wire _4558_;
  wire _4559_;
  wire _4560_;
  wire _4561_;
  wire _4562_;
  wire _4563_;
  wire _4564_;
  wire _4565_;
  wire _4566_;
  wire _4567_;
  wire _4568_;
  wire _4569_;
  wire _4570_;
  wire _4571_;
  wire _4572_;
  wire _4573_;
  wire _4574_;
  wire _4575_;
  wire _4576_;
  wire _4577_;
  wire _4578_;
  wire _4579_;
  wire _4580_;
  wire _4581_;
  wire _4582_;
  wire _4583_;
  wire _4584_;
  wire _4585_;
  wire _4586_;
  wire _4587_;
  wire _4588_;
  wire _4589_;
  wire _4590_;
  wire _4591_;
  wire _4592_;
  wire _4593_;
  wire _4594_;
  wire _4595_;
  wire _4596_;
  wire _4597_;
  wire _4598_;
  wire _4599_;
  wire _4600_;
  wire _4601_;
  wire _4602_;
  wire _4603_;
  wire _4604_;
  wire _4605_;
  wire _4606_;
  wire _4607_;
  wire _4608_;
  wire _4609_;
  wire _4610_;
  wire _4611_;
  wire _4612_;
  wire _4613_;
  wire _4614_;
  wire _4615_;
  wire _4616_;
  wire _4617_;
  wire _4618_;
  wire _4619_;
  wire _4620_;
  wire _4621_;
  wire _4622_;
  wire _4623_;
  wire _4624_;
  wire _4625_;
  wire _4626_;
  wire _4627_;
  wire _4628_;
  wire _4629_;
  wire _4630_;
  wire _4631_;
  wire _4632_;
  wire _4633_;
  wire _4634_;
  wire _4635_;
  wire _4636_;
  wire _4637_;
  wire _4638_;
  wire _4639_;
  wire _4640_;
  wire _4641_;
  wire _4642_;
  wire _4643_;
  wire _4644_;
  wire _4645_;
  wire _4646_;
  wire _4647_;
  wire _4648_;
  wire _4649_;
  wire _4650_;
  wire _4651_;
  wire _4652_;
  wire _4653_;
  wire _4654_;
  wire _4655_;
  wire _4656_;
  wire _4657_;
  wire _4658_;
  wire _4659_;
  wire _4660_;
  wire _4661_;
  wire _4662_;
  wire _4663_;
  wire _4664_;
  wire _4665_;
  wire _4666_;
  wire _4667_;
  wire _4668_;
  wire _4669_;
  wire _4670_;
  wire _4671_;
  wire _4672_;
  wire _4673_;
  wire _4674_;
  wire _4675_;
  wire _4676_;
  wire _4677_;
  wire _4678_;
  wire _4679_;
  wire _4680_;
  wire _4681_;
  wire _4682_;
  wire _4683_;
  wire _4684_;
  wire _4685_;
  wire _4686_;
  wire _4687_;
  wire _4688_;
  wire _4689_;
  wire _4690_;
  wire _4691_;
  wire _4692_;
  wire _4693_;
  wire _4694_;
  wire _4695_;
  wire _4696_;
  wire _4697_;
  wire _4698_;
  wire _4699_;
  wire _4700_;
  wire _4701_;
  wire _4702_;
  wire _4703_;
  wire _4704_;
  wire _4705_;
  wire _4706_;
  wire _4707_;
  wire _4708_;
  wire _4709_;
  wire _4710_;
  wire _4711_;
  wire _4712_;
  wire _4713_;
  wire _4714_;
  wire _4715_;
  wire _4716_;
  wire _4717_;
  wire _4718_;
  wire _4719_;
  wire _4720_;
  wire _4721_;
  wire _4722_;
  wire _4723_;
  wire _4724_;
  wire _4725_;
  wire _4726_;
  wire _4727_;
  wire _4728_;
  wire _4729_;
  wire _4730_;
  wire _4731_;
  wire _4732_;
  wire _4733_;
  wire _4734_;
  wire _4735_;
  wire _4736_;
  wire _4737_;
  wire _4738_;
  wire _4739_;
  wire _4740_;
  wire _4741_;
  wire _4742_;
  wire _4743_;
  wire _4744_;
  wire _4745_;
  wire _4746_;
  wire _4747_;
  wire _4748_;
  wire _4749_;
  wire _4750_;
  wire _4751_;
  wire _4752_;
  wire _4753_;
  wire _4754_;
  wire _4755_;
  wire _4756_;
  wire _4757_;
  wire _4758_;
  wire _4759_;
  wire _4760_;
  wire _4761_;
  wire _4762_;
  wire _4763_;
  wire _4764_;
  wire _4765_;
  wire _4766_;
  wire _4767_;
  wire _4768_;
  wire _4769_;
  wire _4770_;
  wire _4771_;
  wire _4772_;
  wire _4773_;
  wire _4774_;
  wire _4775_;
  wire _4776_;
  wire _4777_;
  wire _4778_;
  wire _4779_;
  wire _4780_;
  wire _4781_;
  wire _4782_;
  wire _4783_;
  wire _4784_;
  wire _4785_;
  wire _4786_;
  wire _4787_;
  wire _4788_;
  wire _4789_;
  wire _4790_;
  wire _4791_;
  wire _4792_;
  wire _4793_;
  wire _4794_;
  wire _4795_;
  wire _4796_;
  wire _4797_;
  wire _4798_;
  wire _4799_;
  wire _4800_;
  wire _4801_;
  wire _4802_;
  wire _4803_;
  wire _4804_;
  wire _4805_;
  wire _4806_;
  wire _4807_;
  wire _4808_;
  wire _4809_;
  wire _4810_;
  wire _4811_;
  wire _4812_;
  wire _4813_;
  wire _4814_;
  wire _4815_;
  wire _4816_;
  wire _4817_;
  wire _4818_;
  wire _4819_;
  wire _4820_;
  wire _4821_;
  wire _4822_;
  wire _4823_;
  wire _4824_;
  wire _4825_;
  wire _4826_;
  wire _4827_;
  wire _4828_;
  wire _4829_;
  wire _4830_;
  wire _4831_;
  wire _4832_;
  wire _4833_;
  wire _4834_;
  wire _4835_;
  wire _4836_;
  wire _4837_;
  wire _4838_;
  wire _4839_;
  wire _4840_;
  wire _4841_;
  wire _4842_;
  wire _4843_;
  wire _4844_;
  wire _4845_;
  wire _4846_;
  wire _4847_;
  wire _4848_;
  wire _4849_;
  wire _4850_;
  wire _4851_;
  wire _4852_;
  wire _4853_;
  wire _4854_;
  wire _4855_;
  wire _4856_;
  wire _4857_;
  wire _4858_;
  wire _4859_;
  wire _4860_;
  wire _4861_;
  wire _4862_;
  wire _4863_;
  wire _4864_;
  wire _4865_;
  wire _4866_;
  wire _4867_;
  wire _4868_;
  wire _4869_;
  wire _4870_;
  wire _4871_;
  wire _4872_;
  wire _4873_;
  wire _4874_;
  wire _4875_;
  wire _4876_;
  wire _4877_;
  wire _4878_;
  wire _4879_;
  wire _4880_;
  wire _4881_;
  wire _4882_;
  wire _4883_;
  wire _4884_;
  wire _4885_;
  wire _4886_;
  wire _4887_;
  wire _4888_;
  wire _4889_;
  wire _4890_;
  wire _4891_;
  wire _4892_;
  wire _4893_;
  wire _4894_;
  wire _4895_;
  wire _4896_;
  wire _4897_;
  wire _4898_;
  wire _4899_;
  wire _4900_;
  wire _4901_;
  wire _4902_;
  wire _4903_;
  wire _4904_;
  wire _4905_;
  wire _4906_;
  wire _4907_;
  wire _4908_;
  wire _4909_;
  wire _4910_;
  wire _4911_;
  wire _4912_;
  wire _4913_;
  wire _4914_;
  wire _4915_;
  wire _4916_;
  wire _4917_;
  wire _4918_;
  wire _4919_;
  wire _4920_;
  wire _4921_;
  wire _4922_;
  wire _4923_;
  wire _4924_;
  wire _4925_;
  wire _4926_;
  wire _4927_;
  wire _4928_;
  wire _4929_;
  wire _4930_;
  wire _4931_;
  wire _4932_;
  wire _4933_;
  wire _4934_;
  wire _4935_;
  wire _4936_;
  wire _4937_;
  wire _4938_;
  wire _4939_;
  wire _4940_;
  wire _4941_;
  wire _4942_;
  wire _4943_;
  wire _4944_;
  wire _4945_;
  wire _4946_;
  wire _4947_;
  wire _4948_;
  wire _4949_;
  wire _4950_;
  wire _4951_;
  wire _4952_;
  wire _4953_;
  wire _4954_;
  wire _4955_;
  wire _4956_;
  wire _4957_;
  wire _4958_;
  wire _4959_;
  wire _4960_;
  wire _4961_;
  wire _4962_;
  wire _4963_;
  wire _4964_;
  wire _4965_;
  wire _4966_;
  wire _4967_;
  wire _4968_;
  wire _4969_;
  wire _4970_;
  wire _4971_;
  wire _4972_;
  wire _4973_;
  wire _4974_;
  wire _4975_;
  wire _4976_;
  wire _4977_;
  wire _4978_;
  wire _4979_;
  wire _4980_;
  wire _4981_;
  wire _4982_;
  wire _4983_;
  wire _4984_;
  wire _4985_;
  wire _4986_;
  wire _4987_;
  wire _4988_;
  wire _4989_;
  wire _4990_;
  wire _4991_;
  wire _4992_;
  wire _4993_;
  wire _4994_;
  wire _4995_;
  wire _4996_;
  wire _4997_;
  wire _4998_;
  wire _4999_;
  wire _5000_;
  wire _5001_;
  wire _5002_;
  wire _5003_;
  wire _5004_;
  wire _5005_;
  wire _5006_;
  wire _5007_;
  wire _5008_;
  wire _5009_;
  wire _5010_;
  wire _5011_;
  wire _5012_;
  wire _5013_;
  wire _5014_;
  wire _5015_;
  wire _5016_;
  wire _5017_;
  wire _5018_;
  wire _5019_;
  wire _5020_;
  wire _5021_;
  wire _5022_;
  wire _5023_;
  wire _5024_;
  wire _5025_;
  wire _5026_;
  wire _5027_;
  wire _5028_;
  wire _5029_;
  wire _5030_;
  wire _5031_;
  wire _5032_;
  wire _5033_;
  wire _5034_;
  wire _5035_;
  wire _5036_;
  wire _5037_;
  wire _5038_;
  wire _5039_;
  wire _5040_;
  wire _5041_;
  wire _5042_;
  wire _5043_;
  wire _5044_;
  wire _5045_;
  wire _5046_;
  wire _5047_;
  wire _5048_;
  wire _5049_;
  wire _5050_;
  wire _5051_;
  wire _5052_;
  wire _5053_;
  wire _5054_;
  wire _5055_;
  wire _5056_;
  wire _5057_;
  wire _5058_;
  wire _5059_;
  wire _5060_;
  wire _5061_;
  wire _5062_;
  wire _5063_;
  wire _5064_;
  wire _5065_;
  wire _5066_;
  wire _5067_;
  wire _5068_;
  wire _5069_;
  wire _5070_;
  wire _5071_;
  wire _5072_;
  wire _5073_;
  wire _5074_;
  wire _5075_;
  wire _5076_;
  wire _5077_;
  wire _5078_;
  wire _5079_;
  wire _5080_;
  wire _5081_;
  wire _5082_;
  wire _5083_;
  wire _5084_;
  wire _5085_;
  wire _5086_;
  wire _5087_;
  wire _5088_;
  wire _5089_;
  wire _5090_;
  wire _5091_;
  wire _5092_;
  wire _5093_;
  wire _5094_;
  wire _5095_;
  wire _5096_;
  wire _5097_;
  wire _5098_;
  wire _5099_;
  wire _5100_;
  wire _5101_;
  wire _5102_;
  wire _5103_;
  wire _5104_;
  wire _5105_;
  wire _5106_;
  wire _5107_;
  wire _5108_;
  wire _5109_;
  wire _5110_;
  wire _5111_;
  wire _5112_;
  wire _5113_;
  wire _5114_;
  wire _5115_;
  wire _5116_;
  wire _5117_;
  wire _5118_;
  wire _5119_;
  wire _5120_;
  wire _5121_;
  wire _5122_;
  wire _5123_;
  wire _5124_;
  wire _5125_;
  wire _5126_;
  wire _5127_;
  wire _5128_;
  wire _5129_;
  wire _5130_;
  wire _5131_;
  wire _5132_;
  wire _5133_;
  wire _5134_;
  wire _5135_;
  wire _5136_;
  wire _5137_;
  wire _5138_;
  wire _5139_;
  wire _5140_;
  wire _5141_;
  wire _5142_;
  wire _5143_;
  wire _5144_;
  wire _5145_;
  wire _5146_;
  wire _5147_;
  wire _5148_;
  wire _5149_;
  wire _5150_;
  wire _5151_;
  wire _5152_;
  wire _5153_;
  wire _5154_;
  wire _5155_;
  wire _5156_;
  wire _5157_;
  wire _5158_;
  wire _5159_;
  wire _5160_;
  wire _5161_;
  wire _5162_;
  wire _5163_;
  wire _5164_;
  wire _5165_;
  wire _5166_;
  wire _5167_;
  wire _5168_;
  wire _5169_;
  wire _5170_;
  wire _5171_;
  wire _5172_;
  wire _5173_;
  wire _5174_;
  wire _5175_;
  wire _5176_;
  wire _5177_;
  wire _5178_;
  wire _5179_;
  wire _5180_;
  wire _5181_;
  wire _5182_;
  wire _5183_;
  wire _5184_;
  wire _5185_;
  wire _5186_;
  wire _5187_;
  wire _5188_;
  wire _5189_;
  wire _5190_;
  wire _5191_;
  wire _5192_;
  wire _5193_;
  wire _5194_;
  wire _5195_;
  wire _5196_;
  wire _5197_;
  wire _5198_;
  wire _5199_;
  wire _5200_;
  wire _5201_;
  wire _5202_;
  wire _5203_;
  wire _5204_;
  wire _5205_;
  wire _5206_;
  wire _5207_;
  wire _5208_;
  wire _5209_;
  wire _5210_;
  wire _5211_;
  wire _5212_;
  wire _5213_;
  wire _5214_;
  wire _5215_;
  wire _5216_;
  wire _5217_;
  wire _5218_;
  wire _5219_;
  wire _5220_;
  wire _5221_;
  wire _5222_;
  wire _5223_;
  wire _5224_;
  wire _5225_;
  wire _5226_;
  wire _5227_;
  wire _5228_;
  wire _5229_;
  wire _5230_;
  wire _5231_;
  wire _5232_;
  wire _5233_;
  wire _5234_;
  wire _5235_;
  wire _5236_;
  wire _5237_;
  wire _5238_;
  wire _5239_;
  wire _5240_;
  wire _5241_;
  wire _5242_;
  wire _5243_;
  wire _5244_;
  wire _5245_;
  wire _5246_;
  wire _5247_;
  wire _5248_;
  wire _5249_;
  wire _5250_;
  wire _5251_;
  wire _5252_;
  wire _5253_;
  wire _5254_;
  wire _5255_;
  wire _5256_;
  wire _5257_;
  wire _5258_;
  wire _5259_;
  wire _5260_;
  wire _5261_;
  wire _5262_;
  wire _5263_;
  wire _5264_;
  wire _5265_;
  wire _5266_;
  wire _5267_;
  wire _5268_;
  wire _5269_;
  wire _5270_;
  wire _5271_;
  wire _5272_;
  wire _5273_;
  wire _5274_;
  wire _5275_;
  wire _5276_;
  wire _5277_;
  wire _5278_;
  wire _5279_;
  wire _5280_;
  wire _5281_;
  wire _5282_;
  wire _5283_;
  wire _5284_;
  wire _5285_;
  wire _5286_;
  wire _5287_;
  wire _5288_;
  wire _5289_;
  wire _5290_;
  wire _5291_;
  wire _5292_;
  wire _5293_;
  wire _5294_;
  wire _5295_;
  wire _5296_;
  wire _5297_;
  wire _5298_;
  wire _5299_;
  wire _5300_;
  wire _5301_;
  wire _5302_;
  wire _5303_;
  wire _5304_;
  wire _5305_;
  wire _5306_;
  wire _5307_;
  wire _5308_;
  wire _5309_;
  wire _5310_;
  wire _5311_;
  wire _5312_;
  wire _5313_;
  wire _5314_;
  wire _5315_;
  wire _5316_;
  wire _5317_;
  wire _5318_;
  wire _5319_;
  wire _5320_;
  wire _5321_;
  wire _5322_;
  wire _5323_;
  wire _5324_;
  wire _5325_;
  wire _5326_;
  wire _5327_;
  wire _5328_;
  wire _5329_;
  wire _5330_;
  wire _5331_;
  wire _5332_;
  wire _5333_;
  wire _5334_;
  wire _5335_;
  wire _5336_;
  wire _5337_;
  wire _5338_;
  wire _5339_;
  wire _5340_;
  wire _5341_;
  wire _5342_;
  wire _5343_;
  wire _5344_;
  wire _5345_;
  wire _5346_;
  wire _5347_;
  wire _5348_;
  wire _5349_;
  wire _5350_;
  wire _5351_;
  wire _5352_;
  wire _5353_;
  wire _5354_;
  wire _5355_;
  wire _5356_;
  wire _5357_;
  wire _5358_;
  wire _5359_;
  wire _5360_;
  wire _5361_;
  wire _5362_;
  wire _5363_;
  wire _5364_;
  wire _5365_;
  wire _5366_;
  wire _5367_;
  wire _5368_;
  wire _5369_;
  wire _5370_;
  wire _5371_;
  wire _5372_;
  wire _5373_;
  wire _5374_;
  wire _5375_;
  wire _5376_;
  wire _5377_;
  wire _5378_;
  wire _5379_;
  wire _5380_;
  wire _5381_;
  wire _5382_;
  wire _5383_;
  wire _5384_;
  wire _5385_;
  wire _5386_;
  wire _5387_;
  wire _5388_;
  wire _5389_;
  wire _5390_;
  wire _5391_;
  wire _5392_;
  wire _5393_;
  wire _5394_;
  wire _5395_;
  wire _5396_;
  wire _5397_;
  wire _5398_;
  wire _5399_;
  wire _5400_;
  wire _5401_;
  wire _5402_;
  wire _5403_;
  wire _5404_;
  wire _5405_;
  wire _5406_;
  wire _5407_;
  wire _5408_;
  wire _5409_;
  wire _5410_;
  wire _5411_;
  wire _5412_;
  wire _5413_;
  wire _5414_;
  wire _5415_;
  wire _5416_;
  wire _5417_;
  wire _5418_;
  wire _5419_;
  wire _5420_;
  wire _5421_;
  wire _5422_;
  wire _5423_;
  wire _5424_;
  wire _5425_;
  wire _5426_;
  wire _5427_;
  wire _5428_;
  wire _5429_;
  wire _5430_;
  wire _5431_;
  wire _5432_;
  wire _5433_;
  wire _5434_;
  wire _5435_;
  wire _5436_;
  wire _5437_;
  wire _5438_;
  wire _5439_;
  wire _5440_;
  wire _5441_;
  wire _5442_;
  wire _5443_;
  wire _5444_;
  wire _5445_;
  wire _5446_;
  wire _5447_;
  wire _5448_;
  wire _5449_;
  wire _5450_;
  wire _5451_;
  wire _5452_;
  wire _5453_;
  wire _5454_;
  wire _5455_;
  wire _5456_;
  wire _5457_;
  wire _5458_;
  wire _5459_;
  wire _5460_;
  wire _5461_;
  wire _5462_;
  wire _5463_;
  wire _5464_;
  wire _5465_;
  wire _5466_;
  wire _5467_;
  wire _5468_;
  wire _5469_;
  wire _5470_;
  wire _5471_;
  wire _5472_;
  wire _5473_;
  wire _5474_;
  wire _5475_;
  wire _5476_;
  wire _5477_;
  wire _5478_;
  wire _5479_;
  wire _5480_;
  wire _5481_;
  wire _5482_;
  wire _5483_;
  wire _5484_;
  wire _5485_;
  wire _5486_;
  wire _5487_;
  wire _5488_;
  wire _5489_;
  wire _5490_;
  wire _5491_;
  wire _5492_;
  wire _5493_;
  wire _5494_;
  wire _5495_;
  wire _5496_;
  wire _5497_;
  wire _5498_;
  wire _5499_;
  wire _5500_;
  wire _5501_;
  wire _5502_;
  wire _5503_;
  wire _5504_;
  wire _5505_;
  wire _5506_;
  wire _5507_;
  wire _5508_;
  wire _5509_;
  wire _5510_;
  wire _5511_;
  wire _5512_;
  wire _5513_;
  wire _5514_;
  wire _5515_;
  wire _5516_;
  wire _5517_;
  wire _5518_;
  wire _5519_;
  wire _5520_;
  wire _5521_;
  wire _5522_;
  wire _5523_;
  wire _5524_;
  wire _5525_;
  wire _5526_;
  wire _5527_;
  wire _5528_;
  wire _5529_;
  wire _5530_;
  wire _5531_;
  wire _5532_;
  wire _5533_;
  wire _5534_;
  wire _5535_;
  wire _5536_;
  wire _5537_;
  wire _5538_;
  wire _5539_;
  wire _5540_;
  wire _5541_;
  wire _5542_;
  wire _5543_;
  wire _5544_;
  wire _5545_;
  wire _5546_;
  wire _5547_;
  wire _5548_;
  wire _5549_;
  wire _5550_;
  wire _5551_;
  wire _5552_;
  wire _5553_;
  wire _5554_;
  wire _5555_;
  wire _5556_;
  wire _5557_;
  wire _5558_;
  wire _5559_;
  wire _5560_;
  wire _5561_;
  wire _5562_;
  wire _5563_;
  wire _5564_;
  wire _5565_;
  wire _5566_;
  wire _5567_;
  wire _5568_;
  wire _5569_;
  wire _5570_;
  wire _5571_;
  wire _5572_;
  wire _5573_;
  wire _5574_;
  wire _5575_;
  wire _5576_;
  wire _5577_;
  wire _5578_;
  wire _5579_;
  wire _5580_;
  wire _5581_;
  wire _5582_;
  wire _5583_;
  wire _5584_;
  wire _5585_;
  wire _5586_;
  wire _5587_;
  wire _5588_;
  wire _5589_;
  wire _5590_;
  wire _5591_;
  wire _5592_;
  wire _5593_;
  wire _5594_;
  wire _5595_;
  wire _5596_;
  wire _5597_;
  wire _5598_;
  wire _5599_;
  wire _5600_;
  wire _5601_;
  wire _5602_;
  wire _5603_;
  wire _5604_;
  wire _5605_;
  wire _5606_;
  wire _5607_;
  wire _5608_;
  wire _5609_;
  wire _5610_;
  wire _5611_;
  wire _5612_;
  wire _5613_;
  wire _5614_;
  wire _5615_;
  wire _5616_;
  wire _5617_;
  wire _5618_;
  wire _5619_;
  wire _5620_;
  wire _5621_;
  wire _5622_;
  wire _5623_;
  wire _5624_;
  wire _5625_;
  wire _5626_;
  wire _5627_;
  wire _5628_;
  wire _5629_;
  wire _5630_;
  wire _5631_;
  wire _5632_;
  wire _5633_;
  wire _5634_;
  wire _5635_;
  wire _5636_;
  wire _5637_;
  wire _5638_;
  wire _5639_;
  wire _5640_;
  wire _5641_;
  wire _5642_;
  wire _5643_;
  wire _5644_;
  wire _5645_;
  wire _5646_;
  wire _5647_;
  wire _5648_;
  wire _5649_;
  wire _5650_;
  wire _5651_;
  wire _5652_;
  wire _5653_;
  wire _5654_;
  wire _5655_;
  wire _5656_;
  wire _5657_;
  wire _5658_;
  wire _5659_;
  wire _5660_;
  wire _5661_;
  wire _5662_;
  wire _5663_;
  wire _5664_;
  wire _5665_;
  wire _5666_;
  wire _5667_;
  wire _5668_;
  wire _5669_;
  wire _5670_;
  wire _5671_;
  wire _5672_;
  wire _5673_;
  wire _5674_;
  wire _5675_;
  wire _5676_;
  wire _5677_;
  wire _5678_;
  wire _5679_;
  wire _5680_;
  wire _5681_;
  wire _5682_;
  wire _5683_;
  wire _5684_;
  wire _5685_;
  wire _5686_;
  wire _5687_;
  wire _5688_;
  wire _5689_;
  wire _5690_;
  wire _5691_;
  wire _5692_;
  wire _5693_;
  wire _5694_;
  wire _5695_;
  wire _5696_;
  wire _5697_;
  wire _5698_;
  wire _5699_;
  wire _5700_;
  wire _5701_;
  wire _5702_;
  wire _5703_;
  wire _5704_;
  wire _5705_;
  wire _5706_;
  wire _5707_;
  wire _5708_;
  wire _5709_;
  wire _5710_;
  wire _5711_;
  wire _5712_;
  wire _5713_;
  wire _5714_;
  wire _5715_;
  wire _5716_;
  wire _5717_;
  wire _5718_;
  wire _5719_;
  wire _5720_;
  wire _5721_;
  wire _5722_;
  wire _5723_;
  wire _5724_;
  wire _5725_;
  wire _5726_;
  wire _5727_;
  wire _5728_;
  wire _5729_;
  wire _5730_;
  wire _5731_;
  wire _5732_;
  wire _5733_;
  wire _5734_;
  wire _5735_;
  wire _5736_;
  wire _5737_;
  wire _5738_;
  wire _5739_;
  wire _5740_;
  wire _5741_;
  wire _5742_;
  wire _5743_;
  wire _5744_;
  wire _5745_;
  wire _5746_;
  wire _5747_;
  wire _5748_;
  wire _5749_;
  wire _5750_;
  wire _5751_;
  wire _5752_;
  wire _5753_;
  wire _5754_;
  wire _5755_;
  wire _5756_;
  wire _5757_;
  wire _5758_;
  wire _5759_;
  wire _5760_;
  wire _5761_;
  wire _5762_;
  wire _5763_;
  wire _5764_;
  wire _5765_;
  wire _5766_;
  wire _5767_;
  wire _5768_;
  wire _5769_;
  wire _5770_;
  wire _5771_;
  wire _5772_;
  wire _5773_;
  wire _5774_;
  wire _5775_;
  wire _5776_;
  wire _5777_;
  wire _5778_;
  wire _5779_;
  wire _5780_;
  wire _5781_;
  wire _5782_;
  wire _5783_;
  wire _5784_;
  wire _5785_;
  wire _5786_;
  wire _5787_;
  wire _5788_;
  wire _5789_;
  wire _5790_;
  wire _5791_;
  wire _5792_;
  wire _5793_;
  wire _5794_;
  wire _5795_;
  wire _5796_;
  wire _5797_;
  wire _5798_;
  wire _5799_;
  wire _5800_;
  wire _5801_;
  wire _5802_;
  wire _5803_;
  wire _5804_;
  wire _5805_;
  wire _5806_;
  wire _5807_;
  wire _5808_;
  wire _5809_;
  wire _5810_;
  wire _5811_;
  wire _5812_;
  wire _5813_;
  wire _5814_;
  wire _5815_;
  wire _5816_;
  wire _5817_;
  wire _5818_;
  wire _5819_;
  wire _5820_;
  wire _5821_;
  wire _5822_;
  wire _5823_;
  wire _5824_;
  wire _5825_;
  wire _5826_;
  wire _5827_;
  wire _5828_;
  wire _5829_;
  wire _5830_;
  wire _5831_;
  wire _5832_;
  wire _5833_;
  wire _5834_;
  wire _5835_;
  wire _5836_;
  wire _5837_;
  wire _5838_;
  wire _5839_;
  wire _5840_;
  wire _5841_;
  wire _5842_;
  wire _5843_;
  wire _5844_;
  wire _5845_;
  wire _5846_;
  wire _5847_;
  wire _5848_;
  wire _5849_;
  wire _5850_;
  wire _5851_;
  wire _5852_;
  wire _5853_;
  wire _5854_;
  wire _5855_;
  wire _5856_;
  wire _5857_;
  wire _5858_;
  wire _5859_;
  wire _5860_;
  wire _5861_;
  wire _5862_;
  wire _5863_;
  wire _5864_;
  wire _5865_;
  wire _5866_;
  wire _5867_;
  wire _5868_;
  wire _5869_;
  wire _5870_;
  wire _5871_;
  wire _5872_;
  wire _5873_;
  wire _5874_;
  wire _5875_;
  wire _5876_;
  wire _5877_;
  wire _5878_;
  wire _5879_;
  wire _5880_;
  wire _5881_;
  wire _5882_;
  wire _5883_;
  wire _5884_;
  wire _5885_;
  wire _5886_;
  wire _5887_;
  wire _5888_;
  wire _5889_;
  wire _5890_;
  wire _5891_;
  wire _5892_;
  wire _5893_;
  wire _5894_;
  wire _5895_;
  wire _5896_;
  wire _5897_;
  wire _5898_;
  wire _5899_;
  wire _5900_;
  wire _5901_;
  wire _5902_;
  wire _5903_;
  wire _5904_;
  wire _5905_;
  wire _5906_;
  wire _5907_;
  wire _5908_;
  wire _5909_;
  wire _5910_;
  wire _5911_;
  wire _5912_;
  wire _5913_;
  wire _5914_;
  wire _5915_;
  wire _5916_;
  wire _5917_;
  wire _5918_;
  wire _5919_;
  wire _5920_;
  wire _5921_;
  wire _5922_;
  wire _5923_;
  wire _5924_;
  wire _5925_;
  wire _5926_;
  wire _5927_;
  wire _5928_;
  wire _5929_;
  wire _5930_;
  wire _5931_;
  wire _5932_;
  wire _5933_;
  wire _5934_;
  wire _5935_;
  wire _5936_;
  wire _5937_;
  wire _5938_;
  wire _5939_;
  wire _5940_;
  wire _5941_;
  wire _5942_;
  wire _5943_;
  wire _5944_;
  wire _5945_;
  wire _5946_;
  wire _5947_;
  wire _5948_;
  wire _5949_;
  wire _5950_;
  wire _5951_;
  wire _5952_;
  wire _5953_;
  wire _5954_;
  wire _5955_;
  wire _5956_;
  wire _5957_;
  wire _5958_;
  wire _5959_;
  wire _5960_;
  wire _5961_;
  wire _5962_;
  wire _5963_;
  wire _5964_;
  wire _5965_;
  wire _5966_;
  wire _5967_;
  wire _5968_;
  wire _5969_;
  wire _5970_;
  wire _5971_;
  wire _5972_;
  wire _5973_;
  wire _5974_;
  wire _5975_;
  wire _5976_;
  wire _5977_;
  wire _5978_;
  wire _5979_;
  wire _5980_;
  wire _5981_;
  wire _5982_;
  wire _5983_;
  wire _5984_;
  wire _5985_;
  wire _5986_;
  wire _5987_;
  wire _5988_;
  wire _5989_;
  wire _5990_;
  wire _5991_;
  wire _5992_;
  wire _5993_;
  wire _5994_;
  wire _5995_;
  wire _5996_;
  wire _5997_;
  wire _5998_;
  wire _5999_;
  wire _6000_;
  wire _6001_;
  wire _6002_;
  wire _6003_;
  wire _6004_;
  wire _6005_;
  wire _6006_;
  wire _6007_;
  wire _6008_;
  wire _6009_;
  wire _6010_;
  wire _6011_;
  wire _6012_;
  wire _6013_;
  wire _6014_;
  wire _6015_;
  wire _6016_;
  wire _6017_;
  wire _6018_;
  wire _6019_;
  wire _6020_;
  wire _6021_;
  wire _6022_;
  wire _6023_;
  wire _6024_;
  wire _6025_;
  wire _6026_;
  wire _6027_;
  wire _6028_;
  wire _6029_;
  wire _6030_;
  wire _6031_;
  wire _6032_;
  wire _6033_;
  wire _6034_;
  wire _6035_;
  wire _6036_;
  wire _6037_;
  wire _6038_;
  wire _6039_;
  wire _6040_;
  wire _6041_;
  wire _6042_;
  wire _6043_;
  wire _6044_;
  wire _6045_;
  wire _6046_;
  wire _6047_;
  wire _6048_;
  wire _6049_;
  wire _6050_;
  wire _6051_;
  wire _6052_;
  wire _6053_;
  wire _6054_;
  wire _6055_;
  wire _6056_;
  wire _6057_;
  wire _6058_;
  wire _6059_;
  wire _6060_;
  wire _6061_;
  wire _6062_;
  wire _6063_;
  wire _6064_;
  wire _6065_;
  wire _6066_;
  wire _6067_;
  wire _6068_;
  wire _6069_;
  wire _6070_;
  wire _6071_;
  wire _6072_;
  wire _6073_;
  wire _6074_;
  wire _6075_;
  wire _6076_;
  wire _6077_;
  wire _6078_;
  wire _6079_;
  wire _6080_;
  wire _6081_;
  wire _6082_;
  wire _6083_;
  wire _6084_;
  wire _6085_;
  wire _6086_;
  wire _6087_;
  wire _6088_;
  wire _6089_;
  wire _6090_;
  wire _6091_;
  wire _6092_;
  wire _6093_;
  wire _6094_;
  wire _6095_;
  wire _6096_;
  wire _6097_;
  wire _6098_;
  wire _6099_;
  wire _6100_;
  wire _6101_;
  wire _6102_;
  wire _6103_;
  wire _6104_;
  wire _6105_;
  wire _6106_;
  wire _6107_;
  wire _6108_;
  wire _6109_;
  wire _6110_;
  wire _6111_;
  wire _6112_;
  wire _6113_;
  wire _6114_;
  wire _6115_;
  wire _6116_;
  wire _6117_;
  wire _6118_;
  wire _6119_;
  wire _6120_;
  wire _6121_;
  wire _6122_;
  wire _6123_;
  wire _6124_;
  wire _6125_;
  wire _6126_;
  wire _6127_;
  wire _6128_;
  wire _6129_;
  wire _6130_;
  wire _6131_;
  wire _6132_;
  wire _6133_;
  wire _6134_;
  wire _6135_;
  wire _6136_;
  wire _6137_;
  wire _6138_;
  wire _6139_;
  wire _6140_;
  wire _6141_;
  wire _6142_;
  wire _6143_;
  wire _6144_;
  wire _6145_;
  wire _6146_;
  wire _6147_;
  wire _6148_;
  wire _6149_;
  wire _6150_;
  wire _6151_;
  wire _6152_;
  wire _6153_;
  wire _6154_;
  wire _6155_;
  wire _6156_;
  wire _6157_;
  wire _6158_;
  wire _6159_;
  wire _6160_;
  wire _6161_;
  wire _6162_;
  wire _6163_;
  wire _6164_;
  wire _6165_;
  wire _6166_;
  wire _6167_;
  wire _6168_;
  wire _6169_;
  wire _6170_;
  wire _6171_;
  wire _6172_;
  wire _6173_;
  wire _6174_;
  wire _6175_;
  wire _6176_;
  wire _6177_;
  wire _6178_;
  wire _6179_;
  wire _6180_;
  wire _6181_;
  wire _6182_;
  wire _6183_;
  wire _6184_;
  wire _6185_;
  wire _6186_;
  wire _6187_;
  wire _6188_;
  wire _6189_;
  wire _6190_;
  wire _6191_;
  wire _6192_;
  wire _6193_;
  wire _6194_;
  wire _6195_;
  wire _6196_;
  wire _6197_;
  wire _6198_;
  wire _6199_;
  wire _6200_;
  wire _6201_;
  wire _6202_;
  wire _6203_;
  wire _6204_;
  wire _6205_;
  wire _6206_;
  wire _6207_;
  wire _6208_;
  wire _6209_;
  wire _6210_;
  wire _6211_;
  wire _6212_;
  wire _6213_;
  wire _6214_;
  wire _6215_;
  wire _6216_;
  wire _6217_;
  wire _6218_;
  wire _6219_;
  wire _6220_;
  wire _6221_;
  wire _6222_;
  wire _6223_;
  wire _6224_;
  wire _6225_;
  wire _6226_;
  wire _6227_;
  wire _6228_;
  wire _6229_;
  wire _6230_;
  wire _6231_;
  wire _6232_;
  wire _6233_;
  wire _6234_;
  wire _6235_;
  wire _6236_;
  wire _6237_;
  wire _6238_;
  wire _6239_;
  wire _6240_;
  wire _6241_;
  wire _6242_;
  wire _6243_;
  wire _6244_;
  wire _6245_;
  wire _6246_;
  wire _6247_;
  wire _6248_;
  wire _6249_;
  wire _6250_;
  wire _6251_;
  wire _6252_;
  wire _6253_;
  wire _6254_;
  wire _6255_;
  wire _6256_;
  wire _6257_;
  wire _6258_;
  wire _6259_;
  wire _6260_;
  wire _6261_;
  wire _6262_;
  wire _6263_;
  wire _6264_;
  wire _6265_;
  wire _6266_;
  wire _6267_;
  wire _6268_;
  wire _6269_;
  wire _6270_;
  wire _6271_;
  wire _6272_;
  wire _6273_;
  wire _6274_;
  wire _6275_;
  wire _6276_;
  wire _6277_;
  wire _6278_;
  wire _6279_;
  wire _6280_;
  wire _6281_;
  wire _6282_;
  wire _6283_;
  wire _6284_;
  wire _6285_;
  wire _6286_;
  wire _6287_;
  wire _6288_;
  wire _6289_;
  wire _6290_;
  wire _6291_;
  wire _6292_;
  wire _6293_;
  wire _6294_;
  wire _6295_;
  wire _6296_;
  wire _6297_;
  wire _6298_;
  wire _6299_;
  wire _6300_;
  wire _6301_;
  wire _6302_;
  wire _6303_;
  wire _6304_;
  wire _6305_;
  wire _6306_;
  wire _6307_;
  wire _6308_;
  wire _6309_;
  wire _6310_;
  wire _6311_;
  wire _6312_;
  wire _6313_;
  wire _6314_;
  wire _6315_;
  wire _6316_;
  wire _6317_;
  wire _6318_;
  wire _6319_;
  wire _6320_;
  wire _6321_;
  wire _6322_;
  wire _6323_;
  wire _6324_;
  wire _6325_;
  wire _6326_;
  wire _6327_;
  wire _6328_;
  wire _6329_;
  wire _6330_;
  wire _6331_;
  wire _6332_;
  wire _6333_;
  wire _6334_;
  wire _6335_;
  wire _6336_;
  wire _6337_;
  wire _6338_;
  wire _6339_;
  wire _6340_;
  wire _6341_;
  wire _6342_;
  wire _6343_;
  wire _6344_;
  wire _6345_;
  wire _6346_;
  wire _6347_;
  wire _6348_;
  wire _6349_;
  wire _6350_;
  wire _6351_;
  wire _6352_;
  wire _6353_;
  wire _6354_;
  wire _6355_;
  wire _6356_;
  wire _6357_;
  wire _6358_;
  wire _6359_;
  wire _6360_;
  wire _6361_;
  wire _6362_;
  wire _6363_;
  wire _6364_;
  wire _6365_;
  wire _6366_;
  wire _6367_;
  wire _6368_;
  wire _6369_;
  wire _6370_;
  wire _6371_;
  wire _6372_;
  wire _6373_;
  wire _6374_;
  wire _6375_;
  wire _6376_;
  wire _6377_;
  wire _6378_;
  wire _6379_;
  wire _6380_;
  wire _6381_;
  wire _6382_;
  wire _6383_;
  wire _6384_;
  wire _6385_;
  wire _6386_;
  wire _6387_;
  wire _6388_;
  wire _6389_;
  wire _6390_;
  wire _6391_;
  wire _6392_;
  wire _6393_;
  wire _6394_;
  wire _6395_;
  wire _6396_;
  wire _6397_;
  wire _6398_;
  wire _6399_;
  wire _6400_;
  wire _6401_;
  wire _6402_;
  wire _6403_;
  wire _6404_;
  wire _6405_;
  wire _6406_;
  wire _6407_;
  wire _6408_;
  wire _6409_;
  wire _6410_;
  wire _6411_;
  wire _6412_;
  wire _6413_;
  wire _6414_;
  wire _6415_;
  wire _6416_;
  wire _6417_;
  wire _6418_;
  wire _6419_;
  wire _6420_;
  wire _6421_;
  wire _6422_;
  wire _6423_;
  wire _6424_;
  wire _6425_;
  wire _6426_;
  wire _6427_;
  wire _6428_;
  wire _6429_;
  wire _6430_;
  wire _6431_;
  wire _6432_;
  wire _6433_;
  wire _6434_;
  wire _6435_;
  wire _6436_;
  wire _6437_;
  wire _6438_;
  wire _6439_;
  wire _6440_;
  wire _6441_;
  wire _6442_;
  wire _6443_;
  wire _6444_;
  wire _6445_;
  wire _6446_;
  wire _6447_;
  wire _6448_;
  wire _6449_;
  wire _6450_;
  wire _6451_;
  wire _6452_;
  wire _6453_;
  wire _6454_;
  wire _6455_;
  wire _6456_;
  wire _6457_;
  wire _6458_;
  wire _6459_;
  wire _6460_;
  wire _6461_;
  wire _6462_;
  wire _6463_;
  wire _6464_;
  wire _6465_;
  wire _6466_;
  wire _6467_;
  wire _6468_;
  wire _6469_;
  wire _6470_;
  wire _6471_;
  wire _6472_;
  wire _6473_;
  wire _6474_;
  wire _6475_;
  wire _6476_;
  wire _6477_;
  wire _6478_;
  wire _6479_;
  wire _6480_;
  wire _6481_;
  wire _6482_;
  wire _6483_;
  wire _6484_;
  wire _6485_;
  wire _6486_;
  wire _6487_;
  wire _6488_;
  wire _6489_;
  wire _6490_;
  wire _6491_;
  wire _6492_;
  wire _6493_;
  wire _6494_;
  wire _6495_;
  wire _6496_;
  wire _6497_;
  wire _6498_;
  wire _6499_;
  wire _6500_;
  wire _6501_;
  wire _6502_;
  wire _6503_;
  wire _6504_;
  wire _6505_;
  wire _6506_;
  wire _6507_;
  wire _6508_;
  wire _6509_;
  wire _6510_;
  wire _6511_;
  wire _6512_;
  wire _6513_;
  wire _6514_;
  wire _6515_;
  wire _6516_;
  wire _6517_;
  wire _6518_;
  wire _6519_;
  wire _6520_;
  wire _6521_;
  wire _6522_;
  wire _6523_;
  wire _6524_;
  wire _6525_;
  wire _6526_;
  wire _6527_;
  wire _6528_;
  wire _6529_;
  wire _6530_;
  wire _6531_;
  wire _6532_;
  wire _6533_;
  wire _6534_;
  wire _6535_;
  wire _6536_;
  wire _6537_;
  wire _6538_;
  wire _6539_;
  wire _6540_;
  wire _6541_;
  wire _6542_;
  wire _6543_;
  wire _6544_;
  wire _6545_;
  wire _6546_;
  wire _6547_;
  wire _6548_;
  wire _6549_;
  wire _6550_;
  wire _6551_;
  wire _6552_;
  wire _6553_;
  wire _6554_;
  wire _6555_;
  wire _6556_;
  wire _6557_;
  wire _6558_;
  wire _6559_;
  wire _6560_;
  wire _6561_;
  wire _6562_;
  wire _6563_;
  wire _6564_;
  wire _6565_;
  wire _6566_;
  wire _6567_;
  wire _6568_;
  wire _6569_;
  wire _6570_;
  wire _6571_;
  wire _6572_;
  wire _6573_;
  wire _6574_;
  wire _6575_;
  wire _6576_;
  wire _6577_;
  wire _6578_;
  wire _6579_;
  wire _6580_;
  wire _6581_;
  wire _6582_;
  wire _6583_;
  wire _6584_;
  wire _6585_;
  wire _6586_;
  wire _6587_;
  wire _6588_;
  wire _6589_;
  wire _6590_;
  wire _6591_;
  wire _6592_;
  wire _6593_;
  wire _6594_;
  wire _6595_;
  wire _6596_;
  wire _6597_;
  wire _6598_;
  wire _6599_;
  wire _6600_;
  wire _6601_;
  wire _6602_;
  wire _6603_;
  wire _6604_;
  wire _6605_;
  wire _6606_;
  wire _6607_;
  wire _6608_;
  wire _6609_;
  wire _6610_;
  wire _6611_;
  wire _6612_;
  wire _6613_;
  wire _6614_;
  wire _6615_;
  wire _6616_;
  wire _6617_;
  wire _6618_;
  wire _6619_;
  wire _6620_;
  wire _6621_;
  wire _6622_;
  wire _6623_;
  wire _6624_;
  wire _6625_;
  wire _6626_;
  wire _6627_;
  wire _6628_;
  wire _6629_;
  wire _6630_;
  wire _6631_;
  wire _6632_;
  wire _6633_;
  wire _6634_;
  wire _6635_;
  wire _6636_;
  wire _6637_;
  wire _6638_;
  wire _6639_;
  wire _6640_;
  wire _6641_;
  wire _6642_;
  wire _6643_;
  wire _6644_;
  wire _6645_;
  wire _6646_;
  wire _6647_;
  wire _6648_;
  wire _6649_;
  wire _6650_;
  wire _6651_;
  wire _6652_;
  wire _6653_;
  wire _6654_;
  wire _6655_;
  wire _6656_;
  wire _6657_;
  wire _6658_;
  wire _6659_;
  wire _6660_;
  wire _6661_;
  wire _6662_;
  wire _6663_;
  wire _6664_;
  wire _6665_;
  wire _6666_;
  wire _6667_;
  wire _6668_;
  wire _6669_;
  wire _6670_;
  wire _6671_;
  wire _6672_;
  wire _6673_;
  wire _6674_;
  wire _6675_;
  wire _6676_;
  wire _6677_;
  wire _6678_;
  wire _6679_;
  wire _6680_;
  wire _6681_;
  wire _6682_;
  wire _6683_;
  wire _6684_;
  wire _6685_;
  wire _6686_;
  wire _6687_;
  wire _6688_;
  wire _6689_;
  wire _6690_;
  wire _6691_;
  wire _6692_;
  wire _6693_;
  wire _6694_;
  wire _6695_;
  wire _6696_;
  wire _6697_;
  wire _6698_;
  wire _6699_;
  wire _6700_;
  wire _6701_;
  wire _6702_;
  wire _6703_;
  wire _6704_;
  wire _6705_;
  wire _6706_;
  wire _6707_;
  wire _6708_;
  wire _6709_;
  wire _6710_;
  wire _6711_;
  wire _6712_;
  wire _6713_;
  wire _6714_;
  wire _6715_;
  wire _6716_;
  wire _6717_;
  wire _6718_;
  wire _6719_;
  wire _6720_;
  wire _6721_;
  wire _6722_;
  wire _6723_;
  wire _6724_;
  wire _6725_;
  wire _6726_;
  wire _6727_;
  wire _6728_;
  wire _6729_;
  wire _6730_;
  wire _6731_;
  wire _6732_;
  wire _6733_;
  wire _6734_;
  wire _6735_;
  wire _6736_;
  wire _6737_;
  wire _6738_;
  wire _6739_;
  wire _6740_;
  wire _6741_;
  wire _6742_;
  wire _6743_;
  wire _6744_;
  wire _6745_;
  wire _6746_;
  wire _6747_;
  wire _6748_;
  wire _6749_;
  wire _6750_;
  wire _6751_;
  wire _6752_;
  wire _6753_;
  wire _6754_;
  wire _6755_;
  wire _6756_;
  wire _6757_;
  wire _6758_;
  wire _6759_;
  wire _6760_;
  wire _6761_;
  wire _6762_;
  wire _6763_;
  wire _6764_;
  wire _6765_;
  wire _6766_;
  wire _6767_;
  wire _6768_;
  wire _6769_;
  wire _6770_;
  wire _6771_;
  wire _6772_;
  wire _6773_;
  wire _6774_;
  wire _6775_;
  wire _6776_;
  wire _6777_;
  wire _6778_;
  wire _6779_;
  wire _6780_;
  wire _6781_;
  wire _6782_;
  wire _6783_;
  wire _6784_;
  wire _6785_;
  wire _6786_;
  wire _6787_;
  wire _6788_;
  wire _6789_;
  wire _6790_;
  wire _6791_;
  wire _6792_;
  wire _6793_;
  wire _6794_;
  wire _6795_;
  wire _6796_;
  wire _6797_;
  wire _6798_;
  wire _6799_;
  wire _6800_;
  wire _6801_;
  wire _6802_;
  wire _6803_;
  wire _6804_;
  wire _6805_;
  wire _6806_;
  wire _6807_;
  wire _6808_;
  wire _6809_;
  wire _6810_;
  wire _6811_;
  wire _6812_;
  wire _6813_;
  wire _6814_;
  wire _6815_;
  wire _6816_;
  wire _6817_;
  wire _6818_;
  wire _6819_;
  wire _6820_;
  wire _6821_;
  wire _6822_;
  wire _6823_;
  wire _6824_;
  wire _6825_;
  wire _6826_;
  wire _6827_;
  wire _6828_;
  wire _6829_;
  wire _6830_;
  wire _6831_;
  wire _6832_;
  wire _6833_;
  wire _6834_;
  wire _6835_;
  wire _6836_;
  wire _6837_;
  wire _6838_;
  wire _6839_;
  wire _6840_;
  wire _6841_;
  wire _6842_;
  wire _6843_;
  wire _6844_;
  wire _6845_;
  wire _6846_;
  wire _6847_;
  wire _6848_;
  wire _6849_;
  wire _6850_;
  wire _6851_;
  wire _6852_;
  wire _6853_;
  wire _6854_;
  wire _6855_;
  wire _6856_;
  wire _6857_;
  wire _6858_;
  wire _6859_;
  wire _6860_;
  wire _6861_;
  wire _6862_;
  wire _6863_;
  wire _6864_;
  wire _6865_;
  wire _6866_;
  wire _6867_;
  wire _6868_;
  wire _6869_;
  wire _6870_;
  wire _6871_;
  wire _6872_;
  wire _6873_;
  wire _6874_;
  wire _6875_;
  wire _6876_;
  wire _6877_;
  wire _6878_;
  wire _6879_;
  wire _6880_;
  wire _6881_;
  wire _6882_;
  wire _6883_;
  wire _6884_;
  wire _6885_;
  wire _6886_;
  wire _6887_;
  wire _6888_;
  wire _6889_;
  wire _6890_;
  wire _6891_;
  wire _6892_;
  wire _6893_;
  wire _6894_;
  wire _6895_;
  wire _6896_;
  wire _6897_;
  wire _6898_;
  wire _6899_;
  wire _6900_;
  wire _6901_;
  wire _6902_;
  wire _6903_;
  wire _6904_;
  wire _6905_;
  wire _6906_;
  wire _6907_;
  wire _6908_;
  wire _6909_;
  wire _6910_;
  wire _6911_;
  wire _6912_;
  wire _6913_;
  wire _6914_;
  wire _6915_;
  wire _6916_;
  wire _6917_;
  wire _6918_;
  wire _6919_;
  wire _6920_;
  wire _6921_;
  wire _6922_;
  wire _6923_;
  wire _6924_;
  wire _6925_;
  wire _6926_;
  wire _6927_;
  wire _6928_;
  wire _6929_;
  wire _6930_;
  wire _6931_;
  wire _6932_;
  wire _6933_;
  wire _6934_;
  wire _6935_;
  wire _6936_;
  wire _6937_;
  wire _6938_;
  wire _6939_;
  wire _6940_;
  wire _6941_;
  wire _6942_;
  wire _6943_;
  wire _6944_;
  wire _6945_;
  wire _6946_;
  wire _6947_;
  wire _6948_;
  wire _6949_;
  wire _6950_;
  wire _6951_;
  wire _6952_;
  wire _6953_;
  wire _6954_;
  wire _6955_;
  wire _6956_;
  wire _6957_;
  wire _6958_;
  wire _6959_;
  wire _6960_;
  wire _6961_;
  wire _6962_;
  wire _6963_;
  wire _6964_;
  wire _6965_;
  wire _6966_;
  wire _6967_;
  wire _6968_;
  wire _6969_;
  wire _6970_;
  wire _6971_;
  wire _6972_;
  wire _6973_;
  wire _6974_;
  wire _6975_;
  wire _6976_;
  wire _6977_;
  wire _6978_;
  wire _6979_;
  wire _6980_;
  wire _6981_;
  wire _6982_;
  wire _6983_;
  wire _6984_;
  wire _6985_;
  wire _6986_;
  wire _6987_;
  wire _6988_;
  wire _6989_;
  wire _6990_;
  wire _6991_;
  wire _6992_;
  wire _6993_;
  wire _6994_;
  wire _6995_;
  wire _6996_;
  wire _6997_;
  wire _6998_;
  wire _6999_;
  wire _7000_;
  wire _7001_;
  wire _7002_;
  wire _7003_;
  wire _7004_;
  wire _7005_;
  wire _7006_;
  wire _7007_;
  wire _7008_;
  wire _7009_;
  wire _7010_;
  wire _7011_;
  wire _7012_;
  wire _7013_;
  wire _7014_;
  wire _7015_;
  wire _7016_;
  wire _7017_;
  wire _7018_;
  wire _7019_;
  wire _7020_;
  wire _7021_;
  wire _7022_;
  wire _7023_;
  wire _7024_;
  wire _7025_;
  wire _7026_;
  wire _7027_;
  wire _7028_;
  wire _7029_;
  wire _7030_;
  wire _7031_;
  wire _7032_;
  wire _7033_;
  wire _7034_;
  wire _7035_;
  wire _7036_;
  wire _7037_;
  wire _7038_;
  wire _7039_;
  wire _7040_;
  wire _7041_;
  wire _7042_;
  wire _7043_;
  wire _7044_;
  wire _7045_;
  wire _7046_;
  wire _7047_;
  wire _7048_;
  wire _7049_;
  wire _7050_;
  wire _7051_;
  wire _7052_;
  wire _7053_;
  wire _7054_;
  wire _7055_;
  wire _7056_;
  wire _7057_;
  wire _7058_;
  wire _7059_;
  wire _7060_;
  wire _7061_;
  wire _7062_;
  wire _7063_;
  wire _7064_;
  wire _7065_;
  wire _7066_;
  wire _7067_;
  wire _7068_;
  wire _7069_;
  wire _7070_;
  wire _7071_;
  wire _7072_;
  wire _7073_;
  wire _7074_;
  wire _7075_;
  wire _7076_;
  wire _7077_;
  wire _7078_;
  wire _7079_;
  wire _7080_;
  wire _7081_;
  wire _7082_;
  wire _7083_;
  wire _7084_;
  wire _7085_;
  wire _7086_;
  wire _7087_;
  wire _7088_;
  wire _7089_;
  wire _7090_;
  wire _7091_;
  wire _7092_;
  wire _7093_;
  wire _7094_;
  wire _7095_;
  wire _7096_;
  wire _7097_;
  wire _7098_;
  wire _7099_;
  wire _7100_;
  wire _7101_;
  wire _7102_;
  wire _7103_;
  wire _7104_;
  wire _7105_;
  wire _7106_;
  wire _7107_;
  wire _7108_;
  wire _7109_;
  wire _7110_;
  wire _7111_;
  wire _7112_;
  wire _7113_;
  wire _7114_;
  wire _7115_;
  wire _7116_;
  wire _7117_;
  wire _7118_;
  wire _7119_;
  wire _7120_;
  wire _7121_;
  wire _7122_;
  wire _7123_;
  wire _7124_;
  wire _7125_;
  wire _7126_;
  wire _7127_;
  wire _7128_;
  wire _7129_;
  wire _7130_;
  wire _7131_;
  wire _7132_;
  wire _7133_;
  wire _7134_;
  wire _7135_;
  wire _7136_;
  wire _7137_;
  wire _7138_;
  wire _7139_;
  wire _7140_;
  wire _7141_;
  wire _7142_;
  wire _7143_;
  wire _7144_;
  wire _7145_;
  wire _7146_;
  wire _7147_;
  wire _7148_;
  wire _7149_;
  wire _7150_;
  wire _7151_;
  wire _7152_;
  wire _7153_;
  wire _7154_;
  wire _7155_;
  wire _7156_;
  wire _7157_;
  wire _7158_;
  wire _7159_;
  wire _7160_;
  wire _7161_;
  wire _7162_;
  wire _7163_;
  wire _7164_;
  wire _7165_;
  wire _7166_;
  wire _7167_;
  wire [62:0] r_0;
  wire [62:0] r_1;
  wire [31:0] m_1;
  wire [31:0] sum_1;
  wire [31:0] inv_1;
  wire [61:0] r_2;
  wire [31:0] m_2;
  wire [31:0] sum_2;
  wire [31:0] inv_2;
  wire [60:0] r_3;
  wire [31:0] m_3;
  wire [31:0] sum_3;
  wire [31:0] inv_3;
  wire [59:0] r_4;
  wire [31:0] m_4;
  wire [31:0] sum_4;
  wire [31:0] inv_4;
  wire [58:0] r_5;
  wire [31:0] m_5;
  wire [31:0] sum_5;
  wire [31:0] inv_5;
  wire [57:0] r_6;
  wire [31:0] m_6;
  wire [31:0] sum_6;
  wire [31:0] inv_6;
  wire [56:0] r_7;
  wire [31:0] m_7;
  wire [31:0] sum_7;
  wire [31:0] inv_7;
  wire [55:0] r_8;
  wire [31:0] m_8;
  wire [31:0] sum_8;
  wire [31:0] inv_8;
  wire [54:0] r_9;
  wire [31:0] m_9;
  wire [31:0] sum_9;
  wire [31:0] inv_9;
  wire [53:0] r_10;
  wire [31:0] m_10;
  wire [31:0] sum_10;
  wire [31:0] inv_10;
  wire [52:0] r_11;
  wire [31:0] m_11;
  wire [31:0] sum_11;
  wire [31:0] inv_11;
  wire [51:0] r_12;
  wire [31:0] m_12;
  wire [31:0] sum_12;
  wire [31:0] inv_12;
  wire [50:0] r_13;
  wire [31:0] m_13;
  wire [31:0] sum_13;
  wire [31:0] inv_13;
  wire [49:0] r_14;
  wire [31:0] m_14;
  wire [31:0] sum_14;
  wire [31:0] inv_14;
  wire [48:0] r_15;
  wire [31:0] m_15;
  wire [31:0] sum_15;
  wire [31:0] inv_15;
  wire [47:0] r_16;
  wire [31:0] m_16;
  wire [31:0] sum_16;
  wire [31:0] inv_16;
  wire [46:0] r_17;
  wire [31:0] m_17;
  wire [31:0] sum_17;
  wire [31:0] inv_17;
  wire [45:0] r_18;
  wire [31:0] m_18;
  wire [31:0] sum_18;
  wire [31:0] inv_18;
  wire [44:0] r_19;
  wire [31:0] m_19;
  wire [31:0] sum_19;
  wire [31:0] inv_19;
  wire [43:0] r_20;
  wire [31:0] m_20;
  wire [31:0] sum_20;
  wire [31:0] inv_20;
  wire [42:0] r_21;
  wire [31:0] m_21;
  wire [31:0] sum_21;
  wire [31:0] inv_21;
  wire [41:0] r_22;
  wire [31:0] m_22;
  wire [31:0] sum_22;
  wire [31:0] inv_22;
  wire [40:0] r_23;
  wire [31:0] m_23;
  wire [31:0] sum_23;
  wire [31:0] inv_23;
  wire [39:0] r_24;
  wire [31:0] m_24;
  wire [31:0] sum_24;
  wire [31:0] inv_24;
  wire [38:0] r_25;
  wire [31:0] m_25;
  wire [31:0] sum_25;
  wire [31:0] inv_25;
  wire [37:0] r_26;
  wire [31:0] m_26;
  wire [31:0] sum_26;
  wire [31:0] inv_26;
  wire [36:0] r_27;
  wire [31:0] m_27;
  wire [31:0] sum_27;
  wire [31:0] inv_27;
  wire [35:0] r_28;
  wire [31:0] m_28;
  wire [31:0] sum_28;
  wire [31:0] inv_28;
  wire [34:0] r_29;
  wire [31:0] m_29;
  wire [31:0] sum_29;
  wire [31:0] inv_29;
  wire [33:0] r_30;
  wire [31:0] m_30;
  wire [31:0] sum_30;
  wire [31:0] inv_30;
  wire [32:0] r_31;
  wire [31:0] m_31;
  wire [31:0] sum_31;
  wire [31:0] inv_31;
  wire [31:0] r_32;
  wire [31:0] m_32;
  wire [31:0] sum_32;
  wire [31:0] inv_32;
  wire zeroWire;
  wire oneWire;
  input [61:0] rin;
  input [30:0] div;
  output [31:0] q;
  output [31:0] rout;
  assign zeroWire = 1'b0 /*0*/;
  assign oneWire = 1'b1 /*0*/;
  assign r_0[0] = rin[0] /*41735*/;
  assign r_0[1] = rin[1] /*41734*/;
  assign r_0[2] = rin[2] /*41733*/;
  assign r_0[3] = rin[3] /*41732*/;
  assign r_0[4] = rin[4] /*41731*/;
  assign r_0[5] = rin[5] /*41730*/;
  assign r_0[6] = rin[6] /*41729*/;
  assign r_0[7] = rin[7] /*41728*/;
  assign r_0[8] = rin[8] /*41727*/;
  assign r_0[9] = rin[9] /*41726*/;
  assign r_0[10] = rin[10] /*41725*/;
  assign r_0[11] = rin[11] /*41724*/;
  assign r_0[12] = rin[12] /*41723*/;
  assign r_0[13] = rin[13] /*41722*/;
  assign r_0[14] = rin[14] /*41721*/;
  assign r_0[15] = rin[15] /*41720*/;
  assign r_0[16] = rin[16] /*41719*/;
  assign r_0[17] = rin[17] /*41718*/;
  assign r_0[18] = rin[18] /*41717*/;
  assign r_0[19] = rin[19] /*41716*/;
  assign r_0[20] = rin[20] /*41715*/;
  assign r_0[21] = rin[21] /*41714*/;
  assign r_0[22] = rin[22] /*41713*/;
  assign r_0[23] = rin[23] /*41712*/;
  assign r_0[24] = rin[24] /*41711*/;
  assign r_0[25] = rin[25] /*41710*/;
  assign r_0[26] = rin[26] /*41709*/;
  assign r_0[27] = rin[27] /*41708*/;
  assign r_0[28] = rin[28] /*41707*/;
  assign r_0[29] = rin[29] /*41706*/;
  assign r_0[30] = rin[30] /*41705*/;
  assign r_0[31] = rin[31] /*41704*/;
  assign r_0[32] = rin[32] /*41703*/;
  assign r_0[33] = rin[33] /*41702*/;
  assign r_0[34] = rin[34] /*41701*/;
  assign r_0[35] = rin[35] /*41700*/;
  assign r_0[36] = rin[36] /*41699*/;
  assign r_0[37] = rin[37] /*41698*/;
  assign r_0[38] = rin[38] /*41697*/;
  assign r_0[39] = rin[39] /*41696*/;
  assign r_0[40] = rin[40] /*41695*/;
  assign r_0[41] = rin[41] /*41694*/;
  assign r_0[42] = rin[42] /*41693*/;
  assign r_0[43] = rin[43] /*41692*/;
  assign r_0[44] = rin[44] /*41691*/;
  assign r_0[45] = rin[45] /*41690*/;
  assign r_0[46] = rin[46] /*41689*/;
  assign r_0[47] = rin[47] /*41688*/;
  assign r_0[48] = rin[48] /*41687*/;
  assign r_0[49] = rin[49] /*41686*/;
  assign r_0[50] = rin[50] /*41685*/;
  assign r_0[51] = rin[51] /*41684*/;
  assign r_0[52] = rin[52] /*41683*/;
  assign r_0[53] = rin[53] /*41682*/;
  assign r_0[54] = rin[54] /*41681*/;
  assign r_0[55] = rin[55] /*41680*/;
  assign r_0[56] = rin[56] /*41679*/;
  assign r_0[57] = rin[57] /*41678*/;
  assign r_0[58] = rin[58] /*41677*/;
  assign r_0[59] = rin[59] /*41676*/;
  assign r_0[60] = rin[60] /*41675*/;
  assign r_0[61] = rin[61] /*41674*/;
  assign r_0[62] = zeroWire /*41673*/;
  assign inv_1[0] = ~div[0] /*41672*/;
  assign inv_1[1] = ~div[1] /*41671*/;
  assign inv_1[2] = ~div[2] /*41670*/;
  assign inv_1[3] = ~div[3] /*41669*/;
  assign inv_1[4] = ~div[4] /*41668*/;
  assign inv_1[5] = ~div[5] /*41667*/;
  assign inv_1[6] = ~div[6] /*41666*/;
  assign inv_1[7] = ~div[7] /*41665*/;
  assign inv_1[8] = ~div[8] /*41664*/;
  assign inv_1[9] = ~div[9] /*41663*/;
  assign inv_1[10] = ~div[10] /*41662*/;
  assign inv_1[11] = ~div[11] /*41661*/;
  assign inv_1[12] = ~div[12] /*41660*/;
  assign inv_1[13] = ~div[13] /*41659*/;
  assign inv_1[14] = ~div[14] /*41658*/;
  assign inv_1[15] = ~div[15] /*41657*/;
  assign inv_1[16] = ~div[16] /*41656*/;
  assign inv_1[17] = ~div[17] /*41655*/;
  assign inv_1[18] = ~div[18] /*41654*/;
  assign inv_1[19] = ~div[19] /*41653*/;
  assign inv_1[20] = ~div[20] /*41652*/;
  assign inv_1[21] = ~div[21] /*41651*/;
  assign inv_1[22] = ~div[22] /*41650*/;
  assign inv_1[23] = ~div[23] /*41649*/;
  assign inv_1[24] = ~div[24] /*41648*/;
  assign inv_1[25] = ~div[25] /*41647*/;
  assign inv_1[26] = ~div[26] /*41646*/;
  assign inv_1[27] = ~div[27] /*41645*/;
  assign inv_1[28] = ~div[28] /*41644*/;
  assign inv_1[29] = ~div[29] /*41643*/;
  assign inv_1[30] = ~div[30] /*41642*/;
assign inv_1[31] = oneWire /*41641*/;
  assign _0_ = inv_1[0] ^ r_0[31] /*41639*/;
  assign sum_1[0] = _0_ ^ oneWire /*41638*/;
  assign _1_ = _0_ & oneWire /*41637*/;
  assign _2_ = inv_1[0] & r_0[31] /*41636*/;
  assign _3_ = _1_ | _2_ /*41635*/;
  assign _4_ = inv_1[1] ^ r_0[32] /*41634*/;
  assign sum_1[1] = _4_ ^ _3_ /*41633*/;
  assign _5_ = _4_ & _3_ /*41632*/;
  assign _6_ = inv_1[1] & r_0[32] /*41631*/;
  assign _7_ = _5_ | _6_ /*41630*/;
  assign _8_ = inv_1[2] ^ r_0[33] /*41628*/;
  assign sum_1[2] = _8_ ^ _7_ /*41627*/;
  assign _9_ = _8_ & _7_ /*41626*/;
  assign _10_ = inv_1[2] & r_0[33] /*41625*/;
  assign _11_ = _9_ | _10_ /*41624*/;
  assign _12_ = inv_1[3] ^ r_0[34] /*41622*/;
  assign sum_1[3] = _12_ ^ _11_ /*41621*/;
  assign _13_ = _12_ & _11_ /*41620*/;
  assign _14_ = inv_1[3] & r_0[34] /*41619*/;
  assign _15_ = _13_ | _14_ /*41618*/;
  assign _16_ = inv_1[4] ^ r_0[35] /*41616*/;
  assign sum_1[4] = _16_ ^ _15_ /*41615*/;
  assign _17_ = _16_ & _15_ /*41614*/;
  assign _18_ = inv_1[4] & r_0[35] /*41613*/;
  assign _19_ = _17_ | _18_ /*41612*/;
  assign _20_ = inv_1[5] ^ r_0[36] /*41610*/;
  assign sum_1[5] = _20_ ^ _19_ /*41609*/;
  assign _21_ = _20_ & _19_ /*41608*/;
  assign _22_ = inv_1[5] & r_0[36] /*41607*/;
  assign _23_ = _21_ | _22_ /*41606*/;
  assign _24_ = inv_1[6] ^ r_0[37] /*41604*/;
  assign sum_1[6] = _24_ ^ _23_ /*41603*/;
  assign _25_ = _24_ & _23_ /*41602*/;
  assign _26_ = inv_1[6] & r_0[37] /*41601*/;
  assign _27_ = _25_ | _26_ /*41600*/;
  assign _28_ = inv_1[7] ^ r_0[38] /*41598*/;
  assign sum_1[7] = _28_ ^ _27_ /*41597*/;
  assign _29_ = _28_ & _27_ /*41596*/;
  assign _30_ = inv_1[7] & r_0[38] /*41595*/;
  assign _31_ = _29_ | _30_ /*41594*/;
  assign _32_ = inv_1[8] ^ r_0[39] /*41592*/;
  assign sum_1[8] = _32_ ^ _31_ /*41591*/;
  assign _33_ = _32_ & _31_ /*41590*/;
  assign _34_ = inv_1[8] & r_0[39] /*41589*/;
  assign _35_ = _33_ | _34_ /*41588*/;
  assign _36_ = inv_1[9] ^ r_0[40] /*41586*/;
  assign sum_1[9] = _36_ ^ _35_ /*41585*/;
  assign _37_ = _36_ & _35_ /*41584*/;
  assign _38_ = inv_1[9] & r_0[40] /*41583*/;
  assign _39_ = _37_ | _38_ /*41582*/;
  assign _40_ = inv_1[10] ^ r_0[41] /*41580*/;
  assign sum_1[10] = _40_ ^ _39_ /*41579*/;
  assign _41_ = _40_ & _39_ /*41578*/;
  assign _42_ = inv_1[10] & r_0[41] /*41577*/;
  assign _43_ = _41_ | _42_ /*41576*/;
  assign _44_ = inv_1[11] ^ r_0[42] /*41574*/;
  assign sum_1[11] = _44_ ^ _43_ /*41573*/;
  assign _45_ = _44_ & _43_ /*41572*/;
  assign _46_ = inv_1[11] & r_0[42] /*41571*/;
  assign _47_ = _45_ | _46_ /*41570*/;
  assign _48_ = inv_1[12] ^ r_0[43] /*41568*/;
  assign sum_1[12] = _48_ ^ _47_ /*41567*/;
  assign _49_ = _48_ & _47_ /*41566*/;
  assign _50_ = inv_1[12] & r_0[43] /*41565*/;
  assign _51_ = _49_ | _50_ /*41564*/;
  assign _52_ = inv_1[13] ^ r_0[44] /*41562*/;
  assign sum_1[13] = _52_ ^ _51_ /*41561*/;
  assign _53_ = _52_ & _51_ /*41560*/;
  assign _54_ = inv_1[13] & r_0[44] /*41559*/;
  assign _55_ = _53_ | _54_ /*41558*/;
  assign _56_ = inv_1[14] ^ r_0[45] /*41556*/;
  assign sum_1[14] = _56_ ^ _55_ /*41555*/;
  assign _57_ = _56_ & _55_ /*41554*/;
  assign _58_ = inv_1[14] & r_0[45] /*41553*/;
  assign _59_ = _57_ | _58_ /*41552*/;
  assign _60_ = inv_1[15] ^ r_0[46] /*41550*/;
  assign sum_1[15] = _60_ ^ _59_ /*41549*/;
  assign _61_ = _60_ & _59_ /*41548*/;
  assign _62_ = inv_1[15] & r_0[46] /*41547*/;
  assign _63_ = _61_ | _62_ /*41546*/;
  assign _64_ = inv_1[16] ^ r_0[47] /*41544*/;
  assign sum_1[16] = _64_ ^ _63_ /*41543*/;
  assign _65_ = _64_ & _63_ /*41542*/;
  assign _66_ = inv_1[16] & r_0[47] /*41541*/;
  assign _67_ = _65_ | _66_ /*41540*/;
  assign _68_ = inv_1[17] ^ r_0[48] /*41538*/;
  assign sum_1[17] = _68_ ^ _67_ /*41537*/;
  assign _69_ = _68_ & _67_ /*41536*/;
  assign _70_ = inv_1[17] & r_0[48] /*41535*/;
  assign _71_ = _69_ | _70_ /*41534*/;
  assign _72_ = inv_1[18] ^ r_0[49] /*41532*/;
  assign sum_1[18] = _72_ ^ _71_ /*41531*/;
  assign _73_ = _72_ & _71_ /*41530*/;
  assign _74_ = inv_1[18] & r_0[49] /*41529*/;
  assign _75_ = _73_ | _74_ /*41528*/;
  assign _76_ = inv_1[19] ^ r_0[50] /*41526*/;
  assign sum_1[19] = _76_ ^ _75_ /*41525*/;
  assign _77_ = _76_ & _75_ /*41524*/;
  assign _78_ = inv_1[19] & r_0[50] /*41523*/;
  assign _79_ = _77_ | _78_ /*41522*/;
  assign _80_ = inv_1[20] ^ r_0[51] /*41520*/;
  assign sum_1[20] = _80_ ^ _79_ /*41519*/;
  assign _81_ = _80_ & _79_ /*41518*/;
  assign _82_ = inv_1[20] & r_0[51] /*41517*/;
  assign _83_ = _81_ | _82_ /*41516*/;
  assign _84_ = inv_1[21] ^ r_0[52] /*41514*/;
  assign sum_1[21] = _84_ ^ _83_ /*41513*/;
  assign _85_ = _84_ & _83_ /*41512*/;
  assign _86_ = inv_1[21] & r_0[52] /*41511*/;
  assign _87_ = _85_ | _86_ /*41510*/;
  assign _88_ = inv_1[22] ^ r_0[53] /*41508*/;
  assign sum_1[22] = _88_ ^ _87_ /*41507*/;
  assign _89_ = _88_ & _87_ /*41506*/;
  assign _90_ = inv_1[22] & r_0[53] /*41505*/;
  assign _91_ = _89_ | _90_ /*41504*/;
  assign _92_ = inv_1[23] ^ r_0[54] /*41502*/;
  assign sum_1[23] = _92_ ^ _91_ /*41501*/;
  assign _93_ = _92_ & _91_ /*41500*/;
  assign _94_ = inv_1[23] & r_0[54] /*41499*/;
  assign _95_ = _93_ | _94_ /*41498*/;
  assign _96_ = inv_1[24] ^ r_0[55] /*41496*/;
  assign sum_1[24] = _96_ ^ _95_ /*41495*/;
  assign _97_ = _96_ & _95_ /*41494*/;
  assign _98_ = inv_1[24] & r_0[55] /*41493*/;
  assign _99_ = _97_ | _98_ /*41492*/;
  assign _100_ = inv_1[25] ^ r_0[56] /*41490*/;
  assign sum_1[25] = _100_ ^ _99_ /*41489*/;
  assign _101_ = _100_ & _99_ /*41488*/;
  assign _102_ = inv_1[25] & r_0[56] /*41487*/;
  assign _103_ = _101_ | _102_ /*41486*/;
  assign _104_ = inv_1[26] ^ r_0[57] /*41484*/;
  assign sum_1[26] = _104_ ^ _103_ /*41483*/;
  assign _105_ = _104_ & _103_ /*41482*/;
  assign _106_ = inv_1[26] & r_0[57] /*41481*/;
  assign _107_ = _105_ | _106_ /*41480*/;
  assign _108_ = inv_1[27] ^ r_0[58] /*41478*/;
  assign sum_1[27] = _108_ ^ _107_ /*41477*/;
  assign _109_ = _108_ & _107_ /*41476*/;
  assign _110_ = inv_1[27] & r_0[58] /*41475*/;
  assign _111_ = _109_ | _110_ /*41474*/;
  assign _112_ = inv_1[28] ^ r_0[59] /*41472*/;
  assign sum_1[28] = _112_ ^ _111_ /*41471*/;
  assign _113_ = _112_ & _111_ /*41470*/;
  assign _114_ = inv_1[28] & r_0[59] /*41469*/;
  assign _115_ = _113_ | _114_ /*41468*/;
  assign _116_ = inv_1[29] ^ r_0[60] /*41466*/;
  assign sum_1[29] = _116_ ^ _115_ /*41465*/;
  assign _117_ = _116_ & _115_ /*41464*/;
  assign _118_ = inv_1[29] & r_0[60] /*41463*/;
  assign _119_ = _117_ | _118_ /*41462*/;
  assign _120_ = inv_1[30] ^ r_0[61] /*41460*/;
  assign sum_1[30] = _120_ ^ _119_ /*41459*/;
  assign _121_ = _120_ & _119_ /*41458*/;
  assign _122_ = inv_1[30] & r_0[61] /*41457*/;
  assign _123_ = _121_ | _122_ /*41456*/;
  assign _124_ = inv_1[31] ^ r_0[62] /*41454*/;
  assign sum_1[31] = _124_ ^ _123_ /*41453*/;
  assign _125_ = _124_ & _123_ /*41452*/;
  assign _126_ = inv_1[31] & r_0[62] /*41451*/;
  assign _127_ = _125_ | _126_ /*41450*/;
  assign q[31] = ~sum_1[31] /*41477*/;
  assign m_1[0] = r_0[31] /*41476*/;
  assign m_1[1] = r_0[32] /*41475*/;
  assign m_1[2] = r_0[33] /*41474*/;
  assign m_1[3] = r_0[34] /*41473*/;
  assign m_1[4] = r_0[35] /*41472*/;
  assign m_1[5] = r_0[36] /*41471*/;
  assign m_1[6] = r_0[37] /*41470*/;
  assign m_1[7] = r_0[38] /*41469*/;
  assign m_1[8] = r_0[39] /*41468*/;
  assign m_1[9] = r_0[40] /*41467*/;
  assign m_1[10] = r_0[41] /*41466*/;
  assign m_1[11] = r_0[42] /*41465*/;
  assign m_1[12] = r_0[43] /*41464*/;
  assign m_1[13] = r_0[44] /*41463*/;
  assign m_1[14] = r_0[45] /*41462*/;
  assign m_1[15] = r_0[46] /*41461*/;
  assign m_1[16] = r_0[47] /*41460*/;
  assign m_1[17] = r_0[48] /*41459*/;
  assign m_1[18] = r_0[49] /*41458*/;
  assign m_1[19] = r_0[50] /*41457*/;
  assign m_1[20] = r_0[51] /*41456*/;
  assign m_1[21] = r_0[52] /*41455*/;
  assign m_1[22] = r_0[53] /*41454*/;
  assign m_1[23] = r_0[54] /*41453*/;
  assign m_1[24] = r_0[55] /*41452*/;
  assign m_1[25] = r_0[56] /*41451*/;
  assign m_1[26] = r_0[57] /*41450*/;
  assign m_1[27] = r_0[58] /*41449*/;
  assign m_1[28] = r_0[59] /*41448*/;
  assign m_1[29] = r_0[60] /*41447*/;
  assign m_1[30] = r_0[61] /*41446*/;
  assign m_1[31] = r_0[62] /*41445*/;
  assign _128_ = ~q[31] /*41443*/;
  assign _129_ = sum_1[0] & q[31] /*41442*/;
  assign _130_ = m_1[0] & _128_ /*41441*/;
  assign r_1[31] = _130_ | _129_ /*41440*/;
  assign _131_ = ~q[31] /*41439*/;
  assign _132_ = sum_1[1] & q[31] /*41438*/;
  assign _133_ = m_1[1] & _131_ /*41437*/;
  assign r_1[32] = _133_ | _132_ /*41436*/;
  assign _134_ = ~q[31] /*41435*/;
  assign _135_ = sum_1[2] & q[31] /*41434*/;
  assign _136_ = m_1[2] & _134_ /*41433*/;
  assign r_1[33] = _136_ | _135_ /*41432*/;
  assign _137_ = ~q[31] /*41431*/;
  assign _138_ = sum_1[3] & q[31] /*41430*/;
  assign _139_ = m_1[3] & _137_ /*41429*/;
  assign r_1[34] = _139_ | _138_ /*41428*/;
  assign _140_ = ~q[31] /*41427*/;
  assign _141_ = sum_1[4] & q[31] /*41426*/;
  assign _142_ = m_1[4] & _140_ /*41425*/;
  assign r_1[35] = _142_ | _141_ /*41424*/;
  assign _143_ = ~q[31] /*41423*/;
  assign _144_ = sum_1[5] & q[31] /*41422*/;
  assign _145_ = m_1[5] & _143_ /*41421*/;
  assign r_1[36] = _145_ | _144_ /*41420*/;
  assign _146_ = ~q[31] /*41419*/;
  assign _147_ = sum_1[6] & q[31] /*41418*/;
  assign _148_ = m_1[6] & _146_ /*41417*/;
  assign r_1[37] = _148_ | _147_ /*41416*/;
  assign _149_ = ~q[31] /*41415*/;
  assign _150_ = sum_1[7] & q[31] /*41414*/;
  assign _151_ = m_1[7] & _149_ /*41413*/;
  assign r_1[38] = _151_ | _150_ /*41412*/;
  assign _152_ = ~q[31] /*41411*/;
  assign _153_ = sum_1[8] & q[31] /*41410*/;
  assign _154_ = m_1[8] & _152_ /*41409*/;
  assign r_1[39] = _154_ | _153_ /*41408*/;
  assign _155_ = ~q[31] /*41407*/;
  assign _156_ = sum_1[9] & q[31] /*41406*/;
  assign _157_ = m_1[9] & _155_ /*41405*/;
  assign r_1[40] = _157_ | _156_ /*41404*/;
  assign _158_ = ~q[31] /*41403*/;
  assign _159_ = sum_1[10] & q[31] /*41402*/;
  assign _160_ = m_1[10] & _158_ /*41401*/;
  assign r_1[41] = _160_ | _159_ /*41400*/;
  assign _161_ = ~q[31] /*41399*/;
  assign _162_ = sum_1[11] & q[31] /*41398*/;
  assign _163_ = m_1[11] & _161_ /*41397*/;
  assign r_1[42] = _163_ | _162_ /*41396*/;
  assign _164_ = ~q[31] /*41395*/;
  assign _165_ = sum_1[12] & q[31] /*41394*/;
  assign _166_ = m_1[12] & _164_ /*41393*/;
  assign r_1[43] = _166_ | _165_ /*41392*/;
  assign _167_ = ~q[31] /*41391*/;
  assign _168_ = sum_1[13] & q[31] /*41390*/;
  assign _169_ = m_1[13] & _167_ /*41389*/;
  assign r_1[44] = _169_ | _168_ /*41388*/;
  assign _170_ = ~q[31] /*41387*/;
  assign _171_ = sum_1[14] & q[31] /*41386*/;
  assign _172_ = m_1[14] & _170_ /*41385*/;
  assign r_1[45] = _172_ | _171_ /*41384*/;
  assign _173_ = ~q[31] /*41383*/;
  assign _174_ = sum_1[15] & q[31] /*41382*/;
  assign _175_ = m_1[15] & _173_ /*41381*/;
  assign r_1[46] = _175_ | _174_ /*41380*/;
  assign _176_ = ~q[31] /*41379*/;
  assign _177_ = sum_1[16] & q[31] /*41378*/;
  assign _178_ = m_1[16] & _176_ /*41377*/;
  assign r_1[47] = _178_ | _177_ /*41376*/;
  assign _179_ = ~q[31] /*41375*/;
  assign _180_ = sum_1[17] & q[31] /*41374*/;
  assign _181_ = m_1[17] & _179_ /*41373*/;
  assign r_1[48] = _181_ | _180_ /*41372*/;
  assign _182_ = ~q[31] /*41371*/;
  assign _183_ = sum_1[18] & q[31] /*41370*/;
  assign _184_ = m_1[18] & _182_ /*41369*/;
  assign r_1[49] = _184_ | _183_ /*41368*/;
  assign _185_ = ~q[31] /*41367*/;
  assign _186_ = sum_1[19] & q[31] /*41366*/;
  assign _187_ = m_1[19] & _185_ /*41365*/;
  assign r_1[50] = _187_ | _186_ /*41364*/;
  assign _188_ = ~q[31] /*41363*/;
  assign _189_ = sum_1[20] & q[31] /*41362*/;
  assign _190_ = m_1[20] & _188_ /*41361*/;
  assign r_1[51] = _190_ | _189_ /*41360*/;
  assign _191_ = ~q[31] /*41359*/;
  assign _192_ = sum_1[21] & q[31] /*41358*/;
  assign _193_ = m_1[21] & _191_ /*41357*/;
  assign r_1[52] = _193_ | _192_ /*41356*/;
  assign _194_ = ~q[31] /*41355*/;
  assign _195_ = sum_1[22] & q[31] /*41354*/;
  assign _196_ = m_1[22] & _194_ /*41353*/;
  assign r_1[53] = _196_ | _195_ /*41352*/;
  assign _197_ = ~q[31] /*41351*/;
  assign _198_ = sum_1[23] & q[31] /*41350*/;
  assign _199_ = m_1[23] & _197_ /*41349*/;
  assign r_1[54] = _199_ | _198_ /*41348*/;
  assign _200_ = ~q[31] /*41347*/;
  assign _201_ = sum_1[24] & q[31] /*41346*/;
  assign _202_ = m_1[24] & _200_ /*41345*/;
  assign r_1[55] = _202_ | _201_ /*41344*/;
  assign _203_ = ~q[31] /*41343*/;
  assign _204_ = sum_1[25] & q[31] /*41342*/;
  assign _205_ = m_1[25] & _203_ /*41341*/;
  assign r_1[56] = _205_ | _204_ /*41340*/;
  assign _206_ = ~q[31] /*41339*/;
  assign _207_ = sum_1[26] & q[31] /*41338*/;
  assign _208_ = m_1[26] & _206_ /*41337*/;
  assign r_1[57] = _208_ | _207_ /*41336*/;
  assign _209_ = ~q[31] /*41335*/;
  assign _210_ = sum_1[27] & q[31] /*41334*/;
  assign _211_ = m_1[27] & _209_ /*41333*/;
  assign r_1[58] = _211_ | _210_ /*41332*/;
  assign _212_ = ~q[31] /*41331*/;
  assign _213_ = sum_1[28] & q[31] /*41330*/;
  assign _214_ = m_1[28] & _212_ /*41329*/;
  assign r_1[59] = _214_ | _213_ /*41328*/;
  assign _215_ = ~q[31] /*41327*/;
  assign _216_ = sum_1[29] & q[31] /*41326*/;
  assign _217_ = m_1[29] & _215_ /*41325*/;
  assign r_1[60] = _217_ | _216_ /*41324*/;
  assign _218_ = ~q[31] /*41323*/;
  assign _219_ = sum_1[30] & q[31] /*41322*/;
  assign _220_ = m_1[30] & _218_ /*41321*/;
  assign r_1[61] = _220_ | _219_ /*41320*/;
  assign _221_ = ~q[31] /*41319*/;
  assign _222_ = sum_1[31] & q[31] /*41318*/;
  assign _223_ = m_1[31] & _221_ /*41317*/;
  assign r_1[62] = _223_ | _222_ /*41316*/;
assign r_1[0]= r_0[0] /*41315*/;
assign r_1[1]= r_0[1] /*41314*/;
assign r_1[2]= r_0[2] /*41313*/;
assign r_1[3]= r_0[3] /*41312*/;
assign r_1[4]= r_0[4] /*41311*/;
assign r_1[5]= r_0[5] /*41310*/;
assign r_1[6]= r_0[6] /*41309*/;
assign r_1[7]= r_0[7] /*41308*/;
assign r_1[8]= r_0[8] /*41307*/;
assign r_1[9]= r_0[9] /*41306*/;
assign r_1[10]= r_0[10] /*41305*/;
assign r_1[11]= r_0[11] /*41304*/;
assign r_1[12]= r_0[12] /*41303*/;
assign r_1[13]= r_0[13] /*41302*/;
assign r_1[14]= r_0[14] /*41301*/;
assign r_1[15]= r_0[15] /*41300*/;
assign r_1[16]= r_0[16] /*41299*/;
assign r_1[17]= r_0[17] /*41298*/;
assign r_1[18]= r_0[18] /*41297*/;
assign r_1[19]= r_0[19] /*41296*/;
assign r_1[20]= r_0[20] /*41295*/;
assign r_1[21]= r_0[21] /*41294*/;
assign r_1[22]= r_0[22] /*41293*/;
assign r_1[23]= r_0[23] /*41292*/;
assign r_1[24]= r_0[24] /*41291*/;
assign r_1[25]= r_0[25] /*41290*/;
assign r_1[26]= r_0[26] /*41289*/;
assign r_1[27]= r_0[27] /*41288*/;
assign r_1[28]= r_0[28] /*41287*/;
assign r_1[29]= r_0[29] /*41286*/;
assign r_1[30]= r_0[30] /*41285*/;
  assign inv_2[0] = ~div[0] /*41224*/;
  assign inv_2[1] = ~div[1] /*41223*/;
  assign inv_2[2] = ~div[2] /*41222*/;
  assign inv_2[3] = ~div[3] /*41221*/;
  assign inv_2[4] = ~div[4] /*41220*/;
  assign inv_2[5] = ~div[5] /*41219*/;
  assign inv_2[6] = ~div[6] /*41218*/;
  assign inv_2[7] = ~div[7] /*41217*/;
  assign inv_2[8] = ~div[8] /*41216*/;
  assign inv_2[9] = ~div[9] /*41215*/;
  assign inv_2[10] = ~div[10] /*41214*/;
  assign inv_2[11] = ~div[11] /*41213*/;
  assign inv_2[12] = ~div[12] /*41212*/;
  assign inv_2[13] = ~div[13] /*41211*/;
  assign inv_2[14] = ~div[14] /*41210*/;
  assign inv_2[15] = ~div[15] /*41209*/;
  assign inv_2[16] = ~div[16] /*41208*/;
  assign inv_2[17] = ~div[17] /*41207*/;
  assign inv_2[18] = ~div[18] /*41206*/;
  assign inv_2[19] = ~div[19] /*41205*/;
  assign inv_2[20] = ~div[20] /*41204*/;
  assign inv_2[21] = ~div[21] /*41203*/;
  assign inv_2[22] = ~div[22] /*41202*/;
  assign inv_2[23] = ~div[23] /*41201*/;
  assign inv_2[24] = ~div[24] /*41200*/;
  assign inv_2[25] = ~div[25] /*41199*/;
  assign inv_2[26] = ~div[26] /*41198*/;
  assign inv_2[27] = ~div[27] /*41197*/;
  assign inv_2[28] = ~div[28] /*41196*/;
  assign inv_2[29] = ~div[29] /*41195*/;
  assign inv_2[30] = ~div[30] /*41194*/;
assign inv_2[31] = oneWire /*41193*/;
  assign _224_ = inv_2[0] ^ r_1[30] /*41191*/;
  assign sum_2[0] = _224_ ^ oneWire /*41190*/;
  assign _225_ = _224_ & oneWire /*41189*/;
  assign _226_ = inv_2[0] & r_1[30] /*41188*/;
  assign _227_ = _225_ | _226_ /*41187*/;
  assign _228_ = inv_2[1] ^ r_1[31] /*41186*/;
  assign sum_2[1] = _228_ ^ _227_ /*41185*/;
  assign _229_ = _228_ & _227_ /*41184*/;
  assign _230_ = inv_2[1] & r_1[31] /*41183*/;
  assign _231_ = _229_ | _230_ /*41182*/;
  assign _232_ = inv_2[2] ^ r_1[32] /*41180*/;
  assign sum_2[2] = _232_ ^ _231_ /*41179*/;
  assign _233_ = _232_ & _231_ /*41178*/;
  assign _234_ = inv_2[2] & r_1[32] /*41177*/;
  assign _235_ = _233_ | _234_ /*41176*/;
  assign _236_ = inv_2[3] ^ r_1[33] /*41174*/;
  assign sum_2[3] = _236_ ^ _235_ /*41173*/;
  assign _237_ = _236_ & _235_ /*41172*/;
  assign _238_ = inv_2[3] & r_1[33] /*41171*/;
  assign _239_ = _237_ | _238_ /*41170*/;
  assign _240_ = inv_2[4] ^ r_1[34] /*41168*/;
  assign sum_2[4] = _240_ ^ _239_ /*41167*/;
  assign _241_ = _240_ & _239_ /*41166*/;
  assign _242_ = inv_2[4] & r_1[34] /*41165*/;
  assign _243_ = _241_ | _242_ /*41164*/;
  assign _244_ = inv_2[5] ^ r_1[35] /*41162*/;
  assign sum_2[5] = _244_ ^ _243_ /*41161*/;
  assign _245_ = _244_ & _243_ /*41160*/;
  assign _246_ = inv_2[5] & r_1[35] /*41159*/;
  assign _247_ = _245_ | _246_ /*41158*/;
  assign _248_ = inv_2[6] ^ r_1[36] /*41156*/;
  assign sum_2[6] = _248_ ^ _247_ /*41155*/;
  assign _249_ = _248_ & _247_ /*41154*/;
  assign _250_ = inv_2[6] & r_1[36] /*41153*/;
  assign _251_ = _249_ | _250_ /*41152*/;
  assign _252_ = inv_2[7] ^ r_1[37] /*41150*/;
  assign sum_2[7] = _252_ ^ _251_ /*41149*/;
  assign _253_ = _252_ & _251_ /*41148*/;
  assign _254_ = inv_2[7] & r_1[37] /*41147*/;
  assign _255_ = _253_ | _254_ /*41146*/;
  assign _256_ = inv_2[8] ^ r_1[38] /*41144*/;
  assign sum_2[8] = _256_ ^ _255_ /*41143*/;
  assign _257_ = _256_ & _255_ /*41142*/;
  assign _258_ = inv_2[8] & r_1[38] /*41141*/;
  assign _259_ = _257_ | _258_ /*41140*/;
  assign _260_ = inv_2[9] ^ r_1[39] /*41138*/;
  assign sum_2[9] = _260_ ^ _259_ /*41137*/;
  assign _261_ = _260_ & _259_ /*41136*/;
  assign _262_ = inv_2[9] & r_1[39] /*41135*/;
  assign _263_ = _261_ | _262_ /*41134*/;
  assign _264_ = inv_2[10] ^ r_1[40] /*41132*/;
  assign sum_2[10] = _264_ ^ _263_ /*41131*/;
  assign _265_ = _264_ & _263_ /*41130*/;
  assign _266_ = inv_2[10] & r_1[40] /*41129*/;
  assign _267_ = _265_ | _266_ /*41128*/;
  assign _268_ = inv_2[11] ^ r_1[41] /*41126*/;
  assign sum_2[11] = _268_ ^ _267_ /*41125*/;
  assign _269_ = _268_ & _267_ /*41124*/;
  assign _270_ = inv_2[11] & r_1[41] /*41123*/;
  assign _271_ = _269_ | _270_ /*41122*/;
  assign _272_ = inv_2[12] ^ r_1[42] /*41120*/;
  assign sum_2[12] = _272_ ^ _271_ /*41119*/;
  assign _273_ = _272_ & _271_ /*41118*/;
  assign _274_ = inv_2[12] & r_1[42] /*41117*/;
  assign _275_ = _273_ | _274_ /*41116*/;
  assign _276_ = inv_2[13] ^ r_1[43] /*41114*/;
  assign sum_2[13] = _276_ ^ _275_ /*41113*/;
  assign _277_ = _276_ & _275_ /*41112*/;
  assign _278_ = inv_2[13] & r_1[43] /*41111*/;
  assign _279_ = _277_ | _278_ /*41110*/;
  assign _280_ = inv_2[14] ^ r_1[44] /*41108*/;
  assign sum_2[14] = _280_ ^ _279_ /*41107*/;
  assign _281_ = _280_ & _279_ /*41106*/;
  assign _282_ = inv_2[14] & r_1[44] /*41105*/;
  assign _283_ = _281_ | _282_ /*41104*/;
  assign _284_ = inv_2[15] ^ r_1[45] /*41102*/;
  assign sum_2[15] = _284_ ^ _283_ /*41101*/;
  assign _285_ = _284_ & _283_ /*41100*/;
  assign _286_ = inv_2[15] & r_1[45] /*41099*/;
  assign _287_ = _285_ | _286_ /*41098*/;
  assign _288_ = inv_2[16] ^ r_1[46] /*41096*/;
  assign sum_2[16] = _288_ ^ _287_ /*41095*/;
  assign _289_ = _288_ & _287_ /*41094*/;
  assign _290_ = inv_2[16] & r_1[46] /*41093*/;
  assign _291_ = _289_ | _290_ /*41092*/;
  assign _292_ = inv_2[17] ^ r_1[47] /*41090*/;
  assign sum_2[17] = _292_ ^ _291_ /*41089*/;
  assign _293_ = _292_ & _291_ /*41088*/;
  assign _294_ = inv_2[17] & r_1[47] /*41087*/;
  assign _295_ = _293_ | _294_ /*41086*/;
  assign _296_ = inv_2[18] ^ r_1[48] /*41084*/;
  assign sum_2[18] = _296_ ^ _295_ /*41083*/;
  assign _297_ = _296_ & _295_ /*41082*/;
  assign _298_ = inv_2[18] & r_1[48] /*41081*/;
  assign _299_ = _297_ | _298_ /*41080*/;
  assign _300_ = inv_2[19] ^ r_1[49] /*41078*/;
  assign sum_2[19] = _300_ ^ _299_ /*41077*/;
  assign _301_ = _300_ & _299_ /*41076*/;
  assign _302_ = inv_2[19] & r_1[49] /*41075*/;
  assign _303_ = _301_ | _302_ /*41074*/;
  assign _304_ = inv_2[20] ^ r_1[50] /*41072*/;
  assign sum_2[20] = _304_ ^ _303_ /*41071*/;
  assign _305_ = _304_ & _303_ /*41070*/;
  assign _306_ = inv_2[20] & r_1[50] /*41069*/;
  assign _307_ = _305_ | _306_ /*41068*/;
  assign _308_ = inv_2[21] ^ r_1[51] /*41066*/;
  assign sum_2[21] = _308_ ^ _307_ /*41065*/;
  assign _309_ = _308_ & _307_ /*41064*/;
  assign _310_ = inv_2[21] & r_1[51] /*41063*/;
  assign _311_ = _309_ | _310_ /*41062*/;
  assign _312_ = inv_2[22] ^ r_1[52] /*41060*/;
  assign sum_2[22] = _312_ ^ _311_ /*41059*/;
  assign _313_ = _312_ & _311_ /*41058*/;
  assign _314_ = inv_2[22] & r_1[52] /*41057*/;
  assign _315_ = _313_ | _314_ /*41056*/;
  assign _316_ = inv_2[23] ^ r_1[53] /*41054*/;
  assign sum_2[23] = _316_ ^ _315_ /*41053*/;
  assign _317_ = _316_ & _315_ /*41052*/;
  assign _318_ = inv_2[23] & r_1[53] /*41051*/;
  assign _319_ = _317_ | _318_ /*41050*/;
  assign _320_ = inv_2[24] ^ r_1[54] /*41048*/;
  assign sum_2[24] = _320_ ^ _319_ /*41047*/;
  assign _321_ = _320_ & _319_ /*41046*/;
  assign _322_ = inv_2[24] & r_1[54] /*41045*/;
  assign _323_ = _321_ | _322_ /*41044*/;
  assign _324_ = inv_2[25] ^ r_1[55] /*41042*/;
  assign sum_2[25] = _324_ ^ _323_ /*41041*/;
  assign _325_ = _324_ & _323_ /*41040*/;
  assign _326_ = inv_2[25] & r_1[55] /*41039*/;
  assign _327_ = _325_ | _326_ /*41038*/;
  assign _328_ = inv_2[26] ^ r_1[56] /*41036*/;
  assign sum_2[26] = _328_ ^ _327_ /*41035*/;
  assign _329_ = _328_ & _327_ /*41034*/;
  assign _330_ = inv_2[26] & r_1[56] /*41033*/;
  assign _331_ = _329_ | _330_ /*41032*/;
  assign _332_ = inv_2[27] ^ r_1[57] /*41030*/;
  assign sum_2[27] = _332_ ^ _331_ /*41029*/;
  assign _333_ = _332_ & _331_ /*41028*/;
  assign _334_ = inv_2[27] & r_1[57] /*41027*/;
  assign _335_ = _333_ | _334_ /*41026*/;
  assign _336_ = inv_2[28] ^ r_1[58] /*41024*/;
  assign sum_2[28] = _336_ ^ _335_ /*41023*/;
  assign _337_ = _336_ & _335_ /*41022*/;
  assign _338_ = inv_2[28] & r_1[58] /*41021*/;
  assign _339_ = _337_ | _338_ /*41020*/;
  assign _340_ = inv_2[29] ^ r_1[59] /*41018*/;
  assign sum_2[29] = _340_ ^ _339_ /*41017*/;
  assign _341_ = _340_ & _339_ /*41016*/;
  assign _342_ = inv_2[29] & r_1[59] /*41015*/;
  assign _343_ = _341_ | _342_ /*41014*/;
  assign _344_ = inv_2[30] ^ r_1[60] /*41012*/;
  assign sum_2[30] = _344_ ^ _343_ /*41011*/;
  assign _345_ = _344_ & _343_ /*41010*/;
  assign _346_ = inv_2[30] & r_1[60] /*41009*/;
  assign _347_ = _345_ | _346_ /*41008*/;
  assign _348_ = inv_2[31] ^ r_1[61] /*41006*/;
  assign sum_2[31] = _348_ ^ _347_ /*41005*/;
  assign _349_ = _348_ & _347_ /*41004*/;
  assign _350_ = inv_2[31] & r_1[61] /*41003*/;
  assign _351_ = _349_ | _350_ /*41002*/;
  assign q[30] = ~sum_2[31] /*41029*/;
  assign m_2[0] = r_1[30] /*41028*/;
  assign m_2[1] = r_1[31] /*41027*/;
  assign m_2[2] = r_1[32] /*41026*/;
  assign m_2[3] = r_1[33] /*41025*/;
  assign m_2[4] = r_1[34] /*41024*/;
  assign m_2[5] = r_1[35] /*41023*/;
  assign m_2[6] = r_1[36] /*41022*/;
  assign m_2[7] = r_1[37] /*41021*/;
  assign m_2[8] = r_1[38] /*41020*/;
  assign m_2[9] = r_1[39] /*41019*/;
  assign m_2[10] = r_1[40] /*41018*/;
  assign m_2[11] = r_1[41] /*41017*/;
  assign m_2[12] = r_1[42] /*41016*/;
  assign m_2[13] = r_1[43] /*41015*/;
  assign m_2[14] = r_1[44] /*41014*/;
  assign m_2[15] = r_1[45] /*41013*/;
  assign m_2[16] = r_1[46] /*41012*/;
  assign m_2[17] = r_1[47] /*41011*/;
  assign m_2[18] = r_1[48] /*41010*/;
  assign m_2[19] = r_1[49] /*41009*/;
  assign m_2[20] = r_1[50] /*41008*/;
  assign m_2[21] = r_1[51] /*41007*/;
  assign m_2[22] = r_1[52] /*41006*/;
  assign m_2[23] = r_1[53] /*41005*/;
  assign m_2[24] = r_1[54] /*41004*/;
  assign m_2[25] = r_1[55] /*41003*/;
  assign m_2[26] = r_1[56] /*41002*/;
  assign m_2[27] = r_1[57] /*41001*/;
  assign m_2[28] = r_1[58] /*41000*/;
  assign m_2[29] = r_1[59] /*40999*/;
  assign m_2[30] = r_1[60] /*40998*/;
  assign m_2[31] = r_1[61] /*40997*/;
  assign _352_ = ~q[30] /*40995*/;
  assign _353_ = sum_2[0] & q[30] /*40994*/;
  assign _354_ = m_2[0] & _352_ /*40993*/;
  assign r_2[30] = _354_ | _353_ /*40992*/;
  assign _355_ = ~q[30] /*40991*/;
  assign _356_ = sum_2[1] & q[30] /*40990*/;
  assign _357_ = m_2[1] & _355_ /*40989*/;
  assign r_2[31] = _357_ | _356_ /*40988*/;
  assign _358_ = ~q[30] /*40987*/;
  assign _359_ = sum_2[2] & q[30] /*40986*/;
  assign _360_ = m_2[2] & _358_ /*40985*/;
  assign r_2[32] = _360_ | _359_ /*40984*/;
  assign _361_ = ~q[30] /*40983*/;
  assign _362_ = sum_2[3] & q[30] /*40982*/;
  assign _363_ = m_2[3] & _361_ /*40981*/;
  assign r_2[33] = _363_ | _362_ /*40980*/;
  assign _364_ = ~q[30] /*40979*/;
  assign _365_ = sum_2[4] & q[30] /*40978*/;
  assign _366_ = m_2[4] & _364_ /*40977*/;
  assign r_2[34] = _366_ | _365_ /*40976*/;
  assign _367_ = ~q[30] /*40975*/;
  assign _368_ = sum_2[5] & q[30] /*40974*/;
  assign _369_ = m_2[5] & _367_ /*40973*/;
  assign r_2[35] = _369_ | _368_ /*40972*/;
  assign _370_ = ~q[30] /*40971*/;
  assign _371_ = sum_2[6] & q[30] /*40970*/;
  assign _372_ = m_2[6] & _370_ /*40969*/;
  assign r_2[36] = _372_ | _371_ /*40968*/;
  assign _373_ = ~q[30] /*40967*/;
  assign _374_ = sum_2[7] & q[30] /*40966*/;
  assign _375_ = m_2[7] & _373_ /*40965*/;
  assign r_2[37] = _375_ | _374_ /*40964*/;
  assign _376_ = ~q[30] /*40963*/;
  assign _377_ = sum_2[8] & q[30] /*40962*/;
  assign _378_ = m_2[8] & _376_ /*40961*/;
  assign r_2[38] = _378_ | _377_ /*40960*/;
  assign _379_ = ~q[30] /*40959*/;
  assign _380_ = sum_2[9] & q[30] /*40958*/;
  assign _381_ = m_2[9] & _379_ /*40957*/;
  assign r_2[39] = _381_ | _380_ /*40956*/;
  assign _382_ = ~q[30] /*40955*/;
  assign _383_ = sum_2[10] & q[30] /*40954*/;
  assign _384_ = m_2[10] & _382_ /*40953*/;
  assign r_2[40] = _384_ | _383_ /*40952*/;
  assign _385_ = ~q[30] /*40951*/;
  assign _386_ = sum_2[11] & q[30] /*40950*/;
  assign _387_ = m_2[11] & _385_ /*40949*/;
  assign r_2[41] = _387_ | _386_ /*40948*/;
  assign _388_ = ~q[30] /*40947*/;
  assign _389_ = sum_2[12] & q[30] /*40946*/;
  assign _390_ = m_2[12] & _388_ /*40945*/;
  assign r_2[42] = _390_ | _389_ /*40944*/;
  assign _391_ = ~q[30] /*40943*/;
  assign _392_ = sum_2[13] & q[30] /*40942*/;
  assign _393_ = m_2[13] & _391_ /*40941*/;
  assign r_2[43] = _393_ | _392_ /*40940*/;
  assign _394_ = ~q[30] /*40939*/;
  assign _395_ = sum_2[14] & q[30] /*40938*/;
  assign _396_ = m_2[14] & _394_ /*40937*/;
  assign r_2[44] = _396_ | _395_ /*40936*/;
  assign _397_ = ~q[30] /*40935*/;
  assign _398_ = sum_2[15] & q[30] /*40934*/;
  assign _399_ = m_2[15] & _397_ /*40933*/;
  assign r_2[45] = _399_ | _398_ /*40932*/;
  assign _400_ = ~q[30] /*40931*/;
  assign _401_ = sum_2[16] & q[30] /*40930*/;
  assign _402_ = m_2[16] & _400_ /*40929*/;
  assign r_2[46] = _402_ | _401_ /*40928*/;
  assign _403_ = ~q[30] /*40927*/;
  assign _404_ = sum_2[17] & q[30] /*40926*/;
  assign _405_ = m_2[17] & _403_ /*40925*/;
  assign r_2[47] = _405_ | _404_ /*40924*/;
  assign _406_ = ~q[30] /*40923*/;
  assign _407_ = sum_2[18] & q[30] /*40922*/;
  assign _408_ = m_2[18] & _406_ /*40921*/;
  assign r_2[48] = _408_ | _407_ /*40920*/;
  assign _409_ = ~q[30] /*40919*/;
  assign _410_ = sum_2[19] & q[30] /*40918*/;
  assign _411_ = m_2[19] & _409_ /*40917*/;
  assign r_2[49] = _411_ | _410_ /*40916*/;
  assign _412_ = ~q[30] /*40915*/;
  assign _413_ = sum_2[20] & q[30] /*40914*/;
  assign _414_ = m_2[20] & _412_ /*40913*/;
  assign r_2[50] = _414_ | _413_ /*40912*/;
  assign _415_ = ~q[30] /*40911*/;
  assign _416_ = sum_2[21] & q[30] /*40910*/;
  assign _417_ = m_2[21] & _415_ /*40909*/;
  assign r_2[51] = _417_ | _416_ /*40908*/;
  assign _418_ = ~q[30] /*40907*/;
  assign _419_ = sum_2[22] & q[30] /*40906*/;
  assign _420_ = m_2[22] & _418_ /*40905*/;
  assign r_2[52] = _420_ | _419_ /*40904*/;
  assign _421_ = ~q[30] /*40903*/;
  assign _422_ = sum_2[23] & q[30] /*40902*/;
  assign _423_ = m_2[23] & _421_ /*40901*/;
  assign r_2[53] = _423_ | _422_ /*40900*/;
  assign _424_ = ~q[30] /*40899*/;
  assign _425_ = sum_2[24] & q[30] /*40898*/;
  assign _426_ = m_2[24] & _424_ /*40897*/;
  assign r_2[54] = _426_ | _425_ /*40896*/;
  assign _427_ = ~q[30] /*40895*/;
  assign _428_ = sum_2[25] & q[30] /*40894*/;
  assign _429_ = m_2[25] & _427_ /*40893*/;
  assign r_2[55] = _429_ | _428_ /*40892*/;
  assign _430_ = ~q[30] /*40891*/;
  assign _431_ = sum_2[26] & q[30] /*40890*/;
  assign _432_ = m_2[26] & _430_ /*40889*/;
  assign r_2[56] = _432_ | _431_ /*40888*/;
  assign _433_ = ~q[30] /*40887*/;
  assign _434_ = sum_2[27] & q[30] /*40886*/;
  assign _435_ = m_2[27] & _433_ /*40885*/;
  assign r_2[57] = _435_ | _434_ /*40884*/;
  assign _436_ = ~q[30] /*40883*/;
  assign _437_ = sum_2[28] & q[30] /*40882*/;
  assign _438_ = m_2[28] & _436_ /*40881*/;
  assign r_2[58] = _438_ | _437_ /*40880*/;
  assign _439_ = ~q[30] /*40879*/;
  assign _440_ = sum_2[29] & q[30] /*40878*/;
  assign _441_ = m_2[29] & _439_ /*40877*/;
  assign r_2[59] = _441_ | _440_ /*40876*/;
  assign _442_ = ~q[30] /*40875*/;
  assign _443_ = sum_2[30] & q[30] /*40874*/;
  assign _444_ = m_2[30] & _442_ /*40873*/;
  assign r_2[60] = _444_ | _443_ /*40872*/;
  assign _445_ = ~q[30] /*40871*/;
  assign _446_ = sum_2[31] & q[30] /*40870*/;
  assign _447_ = m_2[31] & _445_ /*40869*/;
  assign r_2[61] = _447_ | _446_ /*40868*/;
assign r_2[0]= r_1[0] /*40867*/;
assign r_2[1]= r_1[1] /*40866*/;
assign r_2[2]= r_1[2] /*40865*/;
assign r_2[3]= r_1[3] /*40864*/;
assign r_2[4]= r_1[4] /*40863*/;
assign r_2[5]= r_1[5] /*40862*/;
assign r_2[6]= r_1[6] /*40861*/;
assign r_2[7]= r_1[7] /*40860*/;
assign r_2[8]= r_1[8] /*40859*/;
assign r_2[9]= r_1[9] /*40858*/;
assign r_2[10]= r_1[10] /*40857*/;
assign r_2[11]= r_1[11] /*40856*/;
assign r_2[12]= r_1[12] /*40855*/;
assign r_2[13]= r_1[13] /*40854*/;
assign r_2[14]= r_1[14] /*40853*/;
assign r_2[15]= r_1[15] /*40852*/;
assign r_2[16]= r_1[16] /*40851*/;
assign r_2[17]= r_1[17] /*40850*/;
assign r_2[18]= r_1[18] /*40849*/;
assign r_2[19]= r_1[19] /*40848*/;
assign r_2[20]= r_1[20] /*40847*/;
assign r_2[21]= r_1[21] /*40846*/;
assign r_2[22]= r_1[22] /*40845*/;
assign r_2[23]= r_1[23] /*40844*/;
assign r_2[24]= r_1[24] /*40843*/;
assign r_2[25]= r_1[25] /*40842*/;
assign r_2[26]= r_1[26] /*40841*/;
assign r_2[27]= r_1[27] /*40840*/;
assign r_2[28]= r_1[28] /*40839*/;
assign r_2[29]= r_1[29] /*40838*/;
  assign inv_3[0] = ~div[0] /*40776*/;
  assign inv_3[1] = ~div[1] /*40775*/;
  assign inv_3[2] = ~div[2] /*40774*/;
  assign inv_3[3] = ~div[3] /*40773*/;
  assign inv_3[4] = ~div[4] /*40772*/;
  assign inv_3[5] = ~div[5] /*40771*/;
  assign inv_3[6] = ~div[6] /*40770*/;
  assign inv_3[7] = ~div[7] /*40769*/;
  assign inv_3[8] = ~div[8] /*40768*/;
  assign inv_3[9] = ~div[9] /*40767*/;
  assign inv_3[10] = ~div[10] /*40766*/;
  assign inv_3[11] = ~div[11] /*40765*/;
  assign inv_3[12] = ~div[12] /*40764*/;
  assign inv_3[13] = ~div[13] /*40763*/;
  assign inv_3[14] = ~div[14] /*40762*/;
  assign inv_3[15] = ~div[15] /*40761*/;
  assign inv_3[16] = ~div[16] /*40760*/;
  assign inv_3[17] = ~div[17] /*40759*/;
  assign inv_3[18] = ~div[18] /*40758*/;
  assign inv_3[19] = ~div[19] /*40757*/;
  assign inv_3[20] = ~div[20] /*40756*/;
  assign inv_3[21] = ~div[21] /*40755*/;
  assign inv_3[22] = ~div[22] /*40754*/;
  assign inv_3[23] = ~div[23] /*40753*/;
  assign inv_3[24] = ~div[24] /*40752*/;
  assign inv_3[25] = ~div[25] /*40751*/;
  assign inv_3[26] = ~div[26] /*40750*/;
  assign inv_3[27] = ~div[27] /*40749*/;
  assign inv_3[28] = ~div[28] /*40748*/;
  assign inv_3[29] = ~div[29] /*40747*/;
  assign inv_3[30] = ~div[30] /*40746*/;
assign inv_3[31] = oneWire /*40745*/;
  assign _448_ = inv_3[0] ^ r_2[29] /*40743*/;
  assign sum_3[0] = _448_ ^ oneWire /*40742*/;
  assign _449_ = _448_ & oneWire /*40741*/;
  assign _450_ = inv_3[0] & r_2[29] /*40740*/;
  assign _451_ = _449_ | _450_ /*40739*/;
  assign _452_ = inv_3[1] ^ r_2[30] /*40738*/;
  assign sum_3[1] = _452_ ^ _451_ /*40737*/;
  assign _453_ = _452_ & _451_ /*40736*/;
  assign _454_ = inv_3[1] & r_2[30] /*40735*/;
  assign _455_ = _453_ | _454_ /*40734*/;
  assign _456_ = inv_3[2] ^ r_2[31] /*40732*/;
  assign sum_3[2] = _456_ ^ _455_ /*40731*/;
  assign _457_ = _456_ & _455_ /*40730*/;
  assign _458_ = inv_3[2] & r_2[31] /*40729*/;
  assign _459_ = _457_ | _458_ /*40728*/;
  assign _460_ = inv_3[3] ^ r_2[32] /*40726*/;
  assign sum_3[3] = _460_ ^ _459_ /*40725*/;
  assign _461_ = _460_ & _459_ /*40724*/;
  assign _462_ = inv_3[3] & r_2[32] /*40723*/;
  assign _463_ = _461_ | _462_ /*40722*/;
  assign _464_ = inv_3[4] ^ r_2[33] /*40720*/;
  assign sum_3[4] = _464_ ^ _463_ /*40719*/;
  assign _465_ = _464_ & _463_ /*40718*/;
  assign _466_ = inv_3[4] & r_2[33] /*40717*/;
  assign _467_ = _465_ | _466_ /*40716*/;
  assign _468_ = inv_3[5] ^ r_2[34] /*40714*/;
  assign sum_3[5] = _468_ ^ _467_ /*40713*/;
  assign _469_ = _468_ & _467_ /*40712*/;
  assign _470_ = inv_3[5] & r_2[34] /*40711*/;
  assign _471_ = _469_ | _470_ /*40710*/;
  assign _472_ = inv_3[6] ^ r_2[35] /*40708*/;
  assign sum_3[6] = _472_ ^ _471_ /*40707*/;
  assign _473_ = _472_ & _471_ /*40706*/;
  assign _474_ = inv_3[6] & r_2[35] /*40705*/;
  assign _475_ = _473_ | _474_ /*40704*/;
  assign _476_ = inv_3[7] ^ r_2[36] /*40702*/;
  assign sum_3[7] = _476_ ^ _475_ /*40701*/;
  assign _477_ = _476_ & _475_ /*40700*/;
  assign _478_ = inv_3[7] & r_2[36] /*40699*/;
  assign _479_ = _477_ | _478_ /*40698*/;
  assign _480_ = inv_3[8] ^ r_2[37] /*40696*/;
  assign sum_3[8] = _480_ ^ _479_ /*40695*/;
  assign _481_ = _480_ & _479_ /*40694*/;
  assign _482_ = inv_3[8] & r_2[37] /*40693*/;
  assign _483_ = _481_ | _482_ /*40692*/;
  assign _484_ = inv_3[9] ^ r_2[38] /*40690*/;
  assign sum_3[9] = _484_ ^ _483_ /*40689*/;
  assign _485_ = _484_ & _483_ /*40688*/;
  assign _486_ = inv_3[9] & r_2[38] /*40687*/;
  assign _487_ = _485_ | _486_ /*40686*/;
  assign _488_ = inv_3[10] ^ r_2[39] /*40684*/;
  assign sum_3[10] = _488_ ^ _487_ /*40683*/;
  assign _489_ = _488_ & _487_ /*40682*/;
  assign _490_ = inv_3[10] & r_2[39] /*40681*/;
  assign _491_ = _489_ | _490_ /*40680*/;
  assign _492_ = inv_3[11] ^ r_2[40] /*40678*/;
  assign sum_3[11] = _492_ ^ _491_ /*40677*/;
  assign _493_ = _492_ & _491_ /*40676*/;
  assign _494_ = inv_3[11] & r_2[40] /*40675*/;
  assign _495_ = _493_ | _494_ /*40674*/;
  assign _496_ = inv_3[12] ^ r_2[41] /*40672*/;
  assign sum_3[12] = _496_ ^ _495_ /*40671*/;
  assign _497_ = _496_ & _495_ /*40670*/;
  assign _498_ = inv_3[12] & r_2[41] /*40669*/;
  assign _499_ = _497_ | _498_ /*40668*/;
  assign _500_ = inv_3[13] ^ r_2[42] /*40666*/;
  assign sum_3[13] = _500_ ^ _499_ /*40665*/;
  assign _501_ = _500_ & _499_ /*40664*/;
  assign _502_ = inv_3[13] & r_2[42] /*40663*/;
  assign _503_ = _501_ | _502_ /*40662*/;
  assign _504_ = inv_3[14] ^ r_2[43] /*40660*/;
  assign sum_3[14] = _504_ ^ _503_ /*40659*/;
  assign _505_ = _504_ & _503_ /*40658*/;
  assign _506_ = inv_3[14] & r_2[43] /*40657*/;
  assign _507_ = _505_ | _506_ /*40656*/;
  assign _508_ = inv_3[15] ^ r_2[44] /*40654*/;
  assign sum_3[15] = _508_ ^ _507_ /*40653*/;
  assign _509_ = _508_ & _507_ /*40652*/;
  assign _510_ = inv_3[15] & r_2[44] /*40651*/;
  assign _511_ = _509_ | _510_ /*40650*/;
  assign _512_ = inv_3[16] ^ r_2[45] /*40648*/;
  assign sum_3[16] = _512_ ^ _511_ /*40647*/;
  assign _513_ = _512_ & _511_ /*40646*/;
  assign _514_ = inv_3[16] & r_2[45] /*40645*/;
  assign _515_ = _513_ | _514_ /*40644*/;
  assign _516_ = inv_3[17] ^ r_2[46] /*40642*/;
  assign sum_3[17] = _516_ ^ _515_ /*40641*/;
  assign _517_ = _516_ & _515_ /*40640*/;
  assign _518_ = inv_3[17] & r_2[46] /*40639*/;
  assign _519_ = _517_ | _518_ /*40638*/;
  assign _520_ = inv_3[18] ^ r_2[47] /*40636*/;
  assign sum_3[18] = _520_ ^ _519_ /*40635*/;
  assign _521_ = _520_ & _519_ /*40634*/;
  assign _522_ = inv_3[18] & r_2[47] /*40633*/;
  assign _523_ = _521_ | _522_ /*40632*/;
  assign _524_ = inv_3[19] ^ r_2[48] /*40630*/;
  assign sum_3[19] = _524_ ^ _523_ /*40629*/;
  assign _525_ = _524_ & _523_ /*40628*/;
  assign _526_ = inv_3[19] & r_2[48] /*40627*/;
  assign _527_ = _525_ | _526_ /*40626*/;
  assign _528_ = inv_3[20] ^ r_2[49] /*40624*/;
  assign sum_3[20] = _528_ ^ _527_ /*40623*/;
  assign _529_ = _528_ & _527_ /*40622*/;
  assign _530_ = inv_3[20] & r_2[49] /*40621*/;
  assign _531_ = _529_ | _530_ /*40620*/;
  assign _532_ = inv_3[21] ^ r_2[50] /*40618*/;
  assign sum_3[21] = _532_ ^ _531_ /*40617*/;
  assign _533_ = _532_ & _531_ /*40616*/;
  assign _534_ = inv_3[21] & r_2[50] /*40615*/;
  assign _535_ = _533_ | _534_ /*40614*/;
  assign _536_ = inv_3[22] ^ r_2[51] /*40612*/;
  assign sum_3[22] = _536_ ^ _535_ /*40611*/;
  assign _537_ = _536_ & _535_ /*40610*/;
  assign _538_ = inv_3[22] & r_2[51] /*40609*/;
  assign _539_ = _537_ | _538_ /*40608*/;
  assign _540_ = inv_3[23] ^ r_2[52] /*40606*/;
  assign sum_3[23] = _540_ ^ _539_ /*40605*/;
  assign _541_ = _540_ & _539_ /*40604*/;
  assign _542_ = inv_3[23] & r_2[52] /*40603*/;
  assign _543_ = _541_ | _542_ /*40602*/;
  assign _544_ = inv_3[24] ^ r_2[53] /*40600*/;
  assign sum_3[24] = _544_ ^ _543_ /*40599*/;
  assign _545_ = _544_ & _543_ /*40598*/;
  assign _546_ = inv_3[24] & r_2[53] /*40597*/;
  assign _547_ = _545_ | _546_ /*40596*/;
  assign _548_ = inv_3[25] ^ r_2[54] /*40594*/;
  assign sum_3[25] = _548_ ^ _547_ /*40593*/;
  assign _549_ = _548_ & _547_ /*40592*/;
  assign _550_ = inv_3[25] & r_2[54] /*40591*/;
  assign _551_ = _549_ | _550_ /*40590*/;
  assign _552_ = inv_3[26] ^ r_2[55] /*40588*/;
  assign sum_3[26] = _552_ ^ _551_ /*40587*/;
  assign _553_ = _552_ & _551_ /*40586*/;
  assign _554_ = inv_3[26] & r_2[55] /*40585*/;
  assign _555_ = _553_ | _554_ /*40584*/;
  assign _556_ = inv_3[27] ^ r_2[56] /*40582*/;
  assign sum_3[27] = _556_ ^ _555_ /*40581*/;
  assign _557_ = _556_ & _555_ /*40580*/;
  assign _558_ = inv_3[27] & r_2[56] /*40579*/;
  assign _559_ = _557_ | _558_ /*40578*/;
  assign _560_ = inv_3[28] ^ r_2[57] /*40576*/;
  assign sum_3[28] = _560_ ^ _559_ /*40575*/;
  assign _561_ = _560_ & _559_ /*40574*/;
  assign _562_ = inv_3[28] & r_2[57] /*40573*/;
  assign _563_ = _561_ | _562_ /*40572*/;
  assign _564_ = inv_3[29] ^ r_2[58] /*40570*/;
  assign sum_3[29] = _564_ ^ _563_ /*40569*/;
  assign _565_ = _564_ & _563_ /*40568*/;
  assign _566_ = inv_3[29] & r_2[58] /*40567*/;
  assign _567_ = _565_ | _566_ /*40566*/;
  assign _568_ = inv_3[30] ^ r_2[59] /*40564*/;
  assign sum_3[30] = _568_ ^ _567_ /*40563*/;
  assign _569_ = _568_ & _567_ /*40562*/;
  assign _570_ = inv_3[30] & r_2[59] /*40561*/;
  assign _571_ = _569_ | _570_ /*40560*/;
  assign _572_ = inv_3[31] ^ r_2[60] /*40558*/;
  assign sum_3[31] = _572_ ^ _571_ /*40557*/;
  assign _573_ = _572_ & _571_ /*40556*/;
  assign _574_ = inv_3[31] & r_2[60] /*40555*/;
  assign _575_ = _573_ | _574_ /*40554*/;
  assign q[29] = ~sum_3[31] /*40581*/;
  assign m_3[0] = r_2[29] /*40580*/;
  assign m_3[1] = r_2[30] /*40579*/;
  assign m_3[2] = r_2[31] /*40578*/;
  assign m_3[3] = r_2[32] /*40577*/;
  assign m_3[4] = r_2[33] /*40576*/;
  assign m_3[5] = r_2[34] /*40575*/;
  assign m_3[6] = r_2[35] /*40574*/;
  assign m_3[7] = r_2[36] /*40573*/;
  assign m_3[8] = r_2[37] /*40572*/;
  assign m_3[9] = r_2[38] /*40571*/;
  assign m_3[10] = r_2[39] /*40570*/;
  assign m_3[11] = r_2[40] /*40569*/;
  assign m_3[12] = r_2[41] /*40568*/;
  assign m_3[13] = r_2[42] /*40567*/;
  assign m_3[14] = r_2[43] /*40566*/;
  assign m_3[15] = r_2[44] /*40565*/;
  assign m_3[16] = r_2[45] /*40564*/;
  assign m_3[17] = r_2[46] /*40563*/;
  assign m_3[18] = r_2[47] /*40562*/;
  assign m_3[19] = r_2[48] /*40561*/;
  assign m_3[20] = r_2[49] /*40560*/;
  assign m_3[21] = r_2[50] /*40559*/;
  assign m_3[22] = r_2[51] /*40558*/;
  assign m_3[23] = r_2[52] /*40557*/;
  assign m_3[24] = r_2[53] /*40556*/;
  assign m_3[25] = r_2[54] /*40555*/;
  assign m_3[26] = r_2[55] /*40554*/;
  assign m_3[27] = r_2[56] /*40553*/;
  assign m_3[28] = r_2[57] /*40552*/;
  assign m_3[29] = r_2[58] /*40551*/;
  assign m_3[30] = r_2[59] /*40550*/;
  assign m_3[31] = r_2[60] /*40549*/;
  assign _576_ = ~q[29] /*40547*/;
  assign _577_ = sum_3[0] & q[29] /*40546*/;
  assign _578_ = m_3[0] & _576_ /*40545*/;
  assign r_3[29] = _578_ | _577_ /*40544*/;
  assign _579_ = ~q[29] /*40543*/;
  assign _580_ = sum_3[1] & q[29] /*40542*/;
  assign _581_ = m_3[1] & _579_ /*40541*/;
  assign r_3[30] = _581_ | _580_ /*40540*/;
  assign _582_ = ~q[29] /*40539*/;
  assign _583_ = sum_3[2] & q[29] /*40538*/;
  assign _584_ = m_3[2] & _582_ /*40537*/;
  assign r_3[31] = _584_ | _583_ /*40536*/;
  assign _585_ = ~q[29] /*40535*/;
  assign _586_ = sum_3[3] & q[29] /*40534*/;
  assign _587_ = m_3[3] & _585_ /*40533*/;
  assign r_3[32] = _587_ | _586_ /*40532*/;
  assign _588_ = ~q[29] /*40531*/;
  assign _589_ = sum_3[4] & q[29] /*40530*/;
  assign _590_ = m_3[4] & _588_ /*40529*/;
  assign r_3[33] = _590_ | _589_ /*40528*/;
  assign _591_ = ~q[29] /*40527*/;
  assign _592_ = sum_3[5] & q[29] /*40526*/;
  assign _593_ = m_3[5] & _591_ /*40525*/;
  assign r_3[34] = _593_ | _592_ /*40524*/;
  assign _594_ = ~q[29] /*40523*/;
  assign _595_ = sum_3[6] & q[29] /*40522*/;
  assign _596_ = m_3[6] & _594_ /*40521*/;
  assign r_3[35] = _596_ | _595_ /*40520*/;
  assign _597_ = ~q[29] /*40519*/;
  assign _598_ = sum_3[7] & q[29] /*40518*/;
  assign _599_ = m_3[7] & _597_ /*40517*/;
  assign r_3[36] = _599_ | _598_ /*40516*/;
  assign _600_ = ~q[29] /*40515*/;
  assign _601_ = sum_3[8] & q[29] /*40514*/;
  assign _602_ = m_3[8] & _600_ /*40513*/;
  assign r_3[37] = _602_ | _601_ /*40512*/;
  assign _603_ = ~q[29] /*40511*/;
  assign _604_ = sum_3[9] & q[29] /*40510*/;
  assign _605_ = m_3[9] & _603_ /*40509*/;
  assign r_3[38] = _605_ | _604_ /*40508*/;
  assign _606_ = ~q[29] /*40507*/;
  assign _607_ = sum_3[10] & q[29] /*40506*/;
  assign _608_ = m_3[10] & _606_ /*40505*/;
  assign r_3[39] = _608_ | _607_ /*40504*/;
  assign _609_ = ~q[29] /*40503*/;
  assign _610_ = sum_3[11] & q[29] /*40502*/;
  assign _611_ = m_3[11] & _609_ /*40501*/;
  assign r_3[40] = _611_ | _610_ /*40500*/;
  assign _612_ = ~q[29] /*40499*/;
  assign _613_ = sum_3[12] & q[29] /*40498*/;
  assign _614_ = m_3[12] & _612_ /*40497*/;
  assign r_3[41] = _614_ | _613_ /*40496*/;
  assign _615_ = ~q[29] /*40495*/;
  assign _616_ = sum_3[13] & q[29] /*40494*/;
  assign _617_ = m_3[13] & _615_ /*40493*/;
  assign r_3[42] = _617_ | _616_ /*40492*/;
  assign _618_ = ~q[29] /*40491*/;
  assign _619_ = sum_3[14] & q[29] /*40490*/;
  assign _620_ = m_3[14] & _618_ /*40489*/;
  assign r_3[43] = _620_ | _619_ /*40488*/;
  assign _621_ = ~q[29] /*40487*/;
  assign _622_ = sum_3[15] & q[29] /*40486*/;
  assign _623_ = m_3[15] & _621_ /*40485*/;
  assign r_3[44] = _623_ | _622_ /*40484*/;
  assign _624_ = ~q[29] /*40483*/;
  assign _625_ = sum_3[16] & q[29] /*40482*/;
  assign _626_ = m_3[16] & _624_ /*40481*/;
  assign r_3[45] = _626_ | _625_ /*40480*/;
  assign _627_ = ~q[29] /*40479*/;
  assign _628_ = sum_3[17] & q[29] /*40478*/;
  assign _629_ = m_3[17] & _627_ /*40477*/;
  assign r_3[46] = _629_ | _628_ /*40476*/;
  assign _630_ = ~q[29] /*40475*/;
  assign _631_ = sum_3[18] & q[29] /*40474*/;
  assign _632_ = m_3[18] & _630_ /*40473*/;
  assign r_3[47] = _632_ | _631_ /*40472*/;
  assign _633_ = ~q[29] /*40471*/;
  assign _634_ = sum_3[19] & q[29] /*40470*/;
  assign _635_ = m_3[19] & _633_ /*40469*/;
  assign r_3[48] = _635_ | _634_ /*40468*/;
  assign _636_ = ~q[29] /*40467*/;
  assign _637_ = sum_3[20] & q[29] /*40466*/;
  assign _638_ = m_3[20] & _636_ /*40465*/;
  assign r_3[49] = _638_ | _637_ /*40464*/;
  assign _639_ = ~q[29] /*40463*/;
  assign _640_ = sum_3[21] & q[29] /*40462*/;
  assign _641_ = m_3[21] & _639_ /*40461*/;
  assign r_3[50] = _641_ | _640_ /*40460*/;
  assign _642_ = ~q[29] /*40459*/;
  assign _643_ = sum_3[22] & q[29] /*40458*/;
  assign _644_ = m_3[22] & _642_ /*40457*/;
  assign r_3[51] = _644_ | _643_ /*40456*/;
  assign _645_ = ~q[29] /*40455*/;
  assign _646_ = sum_3[23] & q[29] /*40454*/;
  assign _647_ = m_3[23] & _645_ /*40453*/;
  assign r_3[52] = _647_ | _646_ /*40452*/;
  assign _648_ = ~q[29] /*40451*/;
  assign _649_ = sum_3[24] & q[29] /*40450*/;
  assign _650_ = m_3[24] & _648_ /*40449*/;
  assign r_3[53] = _650_ | _649_ /*40448*/;
  assign _651_ = ~q[29] /*40447*/;
  assign _652_ = sum_3[25] & q[29] /*40446*/;
  assign _653_ = m_3[25] & _651_ /*40445*/;
  assign r_3[54] = _653_ | _652_ /*40444*/;
  assign _654_ = ~q[29] /*40443*/;
  assign _655_ = sum_3[26] & q[29] /*40442*/;
  assign _656_ = m_3[26] & _654_ /*40441*/;
  assign r_3[55] = _656_ | _655_ /*40440*/;
  assign _657_ = ~q[29] /*40439*/;
  assign _658_ = sum_3[27] & q[29] /*40438*/;
  assign _659_ = m_3[27] & _657_ /*40437*/;
  assign r_3[56] = _659_ | _658_ /*40436*/;
  assign _660_ = ~q[29] /*40435*/;
  assign _661_ = sum_3[28] & q[29] /*40434*/;
  assign _662_ = m_3[28] & _660_ /*40433*/;
  assign r_3[57] = _662_ | _661_ /*40432*/;
  assign _663_ = ~q[29] /*40431*/;
  assign _664_ = sum_3[29] & q[29] /*40430*/;
  assign _665_ = m_3[29] & _663_ /*40429*/;
  assign r_3[58] = _665_ | _664_ /*40428*/;
  assign _666_ = ~q[29] /*40427*/;
  assign _667_ = sum_3[30] & q[29] /*40426*/;
  assign _668_ = m_3[30] & _666_ /*40425*/;
  assign r_3[59] = _668_ | _667_ /*40424*/;
  assign _669_ = ~q[29] /*40423*/;
  assign _670_ = sum_3[31] & q[29] /*40422*/;
  assign _671_ = m_3[31] & _669_ /*40421*/;
  assign r_3[60] = _671_ | _670_ /*40420*/;
assign r_3[0]= r_2[0] /*40419*/;
assign r_3[1]= r_2[1] /*40418*/;
assign r_3[2]= r_2[2] /*40417*/;
assign r_3[3]= r_2[3] /*40416*/;
assign r_3[4]= r_2[4] /*40415*/;
assign r_3[5]= r_2[5] /*40414*/;
assign r_3[6]= r_2[6] /*40413*/;
assign r_3[7]= r_2[7] /*40412*/;
assign r_3[8]= r_2[8] /*40411*/;
assign r_3[9]= r_2[9] /*40410*/;
assign r_3[10]= r_2[10] /*40409*/;
assign r_3[11]= r_2[11] /*40408*/;
assign r_3[12]= r_2[12] /*40407*/;
assign r_3[13]= r_2[13] /*40406*/;
assign r_3[14]= r_2[14] /*40405*/;
assign r_3[15]= r_2[15] /*40404*/;
assign r_3[16]= r_2[16] /*40403*/;
assign r_3[17]= r_2[17] /*40402*/;
assign r_3[18]= r_2[18] /*40401*/;
assign r_3[19]= r_2[19] /*40400*/;
assign r_3[20]= r_2[20] /*40399*/;
assign r_3[21]= r_2[21] /*40398*/;
assign r_3[22]= r_2[22] /*40397*/;
assign r_3[23]= r_2[23] /*40396*/;
assign r_3[24]= r_2[24] /*40395*/;
assign r_3[25]= r_2[25] /*40394*/;
assign r_3[26]= r_2[26] /*40393*/;
assign r_3[27]= r_2[27] /*40392*/;
assign r_3[28]= r_2[28] /*40391*/;
  assign inv_4[0] = ~div[0] /*40328*/;
  assign inv_4[1] = ~div[1] /*40327*/;
  assign inv_4[2] = ~div[2] /*40326*/;
  assign inv_4[3] = ~div[3] /*40325*/;
  assign inv_4[4] = ~div[4] /*40324*/;
  assign inv_4[5] = ~div[5] /*40323*/;
  assign inv_4[6] = ~div[6] /*40322*/;
  assign inv_4[7] = ~div[7] /*40321*/;
  assign inv_4[8] = ~div[8] /*40320*/;
  assign inv_4[9] = ~div[9] /*40319*/;
  assign inv_4[10] = ~div[10] /*40318*/;
  assign inv_4[11] = ~div[11] /*40317*/;
  assign inv_4[12] = ~div[12] /*40316*/;
  assign inv_4[13] = ~div[13] /*40315*/;
  assign inv_4[14] = ~div[14] /*40314*/;
  assign inv_4[15] = ~div[15] /*40313*/;
  assign inv_4[16] = ~div[16] /*40312*/;
  assign inv_4[17] = ~div[17] /*40311*/;
  assign inv_4[18] = ~div[18] /*40310*/;
  assign inv_4[19] = ~div[19] /*40309*/;
  assign inv_4[20] = ~div[20] /*40308*/;
  assign inv_4[21] = ~div[21] /*40307*/;
  assign inv_4[22] = ~div[22] /*40306*/;
  assign inv_4[23] = ~div[23] /*40305*/;
  assign inv_4[24] = ~div[24] /*40304*/;
  assign inv_4[25] = ~div[25] /*40303*/;
  assign inv_4[26] = ~div[26] /*40302*/;
  assign inv_4[27] = ~div[27] /*40301*/;
  assign inv_4[28] = ~div[28] /*40300*/;
  assign inv_4[29] = ~div[29] /*40299*/;
  assign inv_4[30] = ~div[30] /*40298*/;
assign inv_4[31] = oneWire /*40297*/;
  assign _672_ = inv_4[0] ^ r_3[28] /*40295*/;
  assign sum_4[0] = _672_ ^ oneWire /*40294*/;
  assign _673_ = _672_ & oneWire /*40293*/;
  assign _674_ = inv_4[0] & r_3[28] /*40292*/;
  assign _675_ = _673_ | _674_ /*40291*/;
  assign _676_ = inv_4[1] ^ r_3[29] /*40290*/;
  assign sum_4[1] = _676_ ^ _675_ /*40289*/;
  assign _677_ = _676_ & _675_ /*40288*/;
  assign _678_ = inv_4[1] & r_3[29] /*40287*/;
  assign _679_ = _677_ | _678_ /*40286*/;
  assign _680_ = inv_4[2] ^ r_3[30] /*40284*/;
  assign sum_4[2] = _680_ ^ _679_ /*40283*/;
  assign _681_ = _680_ & _679_ /*40282*/;
  assign _682_ = inv_4[2] & r_3[30] /*40281*/;
  assign _683_ = _681_ | _682_ /*40280*/;
  assign _684_ = inv_4[3] ^ r_3[31] /*40278*/;
  assign sum_4[3] = _684_ ^ _683_ /*40277*/;
  assign _685_ = _684_ & _683_ /*40276*/;
  assign _686_ = inv_4[3] & r_3[31] /*40275*/;
  assign _687_ = _685_ | _686_ /*40274*/;
  assign _688_ = inv_4[4] ^ r_3[32] /*40272*/;
  assign sum_4[4] = _688_ ^ _687_ /*40271*/;
  assign _689_ = _688_ & _687_ /*40270*/;
  assign _690_ = inv_4[4] & r_3[32] /*40269*/;
  assign _691_ = _689_ | _690_ /*40268*/;
  assign _692_ = inv_4[5] ^ r_3[33] /*40266*/;
  assign sum_4[5] = _692_ ^ _691_ /*40265*/;
  assign _693_ = _692_ & _691_ /*40264*/;
  assign _694_ = inv_4[5] & r_3[33] /*40263*/;
  assign _695_ = _693_ | _694_ /*40262*/;
  assign _696_ = inv_4[6] ^ r_3[34] /*40260*/;
  assign sum_4[6] = _696_ ^ _695_ /*40259*/;
  assign _697_ = _696_ & _695_ /*40258*/;
  assign _698_ = inv_4[6] & r_3[34] /*40257*/;
  assign _699_ = _697_ | _698_ /*40256*/;
  assign _700_ = inv_4[7] ^ r_3[35] /*40254*/;
  assign sum_4[7] = _700_ ^ _699_ /*40253*/;
  assign _701_ = _700_ & _699_ /*40252*/;
  assign _702_ = inv_4[7] & r_3[35] /*40251*/;
  assign _703_ = _701_ | _702_ /*40250*/;
  assign _704_ = inv_4[8] ^ r_3[36] /*40248*/;
  assign sum_4[8] = _704_ ^ _703_ /*40247*/;
  assign _705_ = _704_ & _703_ /*40246*/;
  assign _706_ = inv_4[8] & r_3[36] /*40245*/;
  assign _707_ = _705_ | _706_ /*40244*/;
  assign _708_ = inv_4[9] ^ r_3[37] /*40242*/;
  assign sum_4[9] = _708_ ^ _707_ /*40241*/;
  assign _709_ = _708_ & _707_ /*40240*/;
  assign _710_ = inv_4[9] & r_3[37] /*40239*/;
  assign _711_ = _709_ | _710_ /*40238*/;
  assign _712_ = inv_4[10] ^ r_3[38] /*40236*/;
  assign sum_4[10] = _712_ ^ _711_ /*40235*/;
  assign _713_ = _712_ & _711_ /*40234*/;
  assign _714_ = inv_4[10] & r_3[38] /*40233*/;
  assign _715_ = _713_ | _714_ /*40232*/;
  assign _716_ = inv_4[11] ^ r_3[39] /*40230*/;
  assign sum_4[11] = _716_ ^ _715_ /*40229*/;
  assign _717_ = _716_ & _715_ /*40228*/;
  assign _718_ = inv_4[11] & r_3[39] /*40227*/;
  assign _719_ = _717_ | _718_ /*40226*/;
  assign _720_ = inv_4[12] ^ r_3[40] /*40224*/;
  assign sum_4[12] = _720_ ^ _719_ /*40223*/;
  assign _721_ = _720_ & _719_ /*40222*/;
  assign _722_ = inv_4[12] & r_3[40] /*40221*/;
  assign _723_ = _721_ | _722_ /*40220*/;
  assign _724_ = inv_4[13] ^ r_3[41] /*40218*/;
  assign sum_4[13] = _724_ ^ _723_ /*40217*/;
  assign _725_ = _724_ & _723_ /*40216*/;
  assign _726_ = inv_4[13] & r_3[41] /*40215*/;
  assign _727_ = _725_ | _726_ /*40214*/;
  assign _728_ = inv_4[14] ^ r_3[42] /*40212*/;
  assign sum_4[14] = _728_ ^ _727_ /*40211*/;
  assign _729_ = _728_ & _727_ /*40210*/;
  assign _730_ = inv_4[14] & r_3[42] /*40209*/;
  assign _731_ = _729_ | _730_ /*40208*/;
  assign _732_ = inv_4[15] ^ r_3[43] /*40206*/;
  assign sum_4[15] = _732_ ^ _731_ /*40205*/;
  assign _733_ = _732_ & _731_ /*40204*/;
  assign _734_ = inv_4[15] & r_3[43] /*40203*/;
  assign _735_ = _733_ | _734_ /*40202*/;
  assign _736_ = inv_4[16] ^ r_3[44] /*40200*/;
  assign sum_4[16] = _736_ ^ _735_ /*40199*/;
  assign _737_ = _736_ & _735_ /*40198*/;
  assign _738_ = inv_4[16] & r_3[44] /*40197*/;
  assign _739_ = _737_ | _738_ /*40196*/;
  assign _740_ = inv_4[17] ^ r_3[45] /*40194*/;
  assign sum_4[17] = _740_ ^ _739_ /*40193*/;
  assign _741_ = _740_ & _739_ /*40192*/;
  assign _742_ = inv_4[17] & r_3[45] /*40191*/;
  assign _743_ = _741_ | _742_ /*40190*/;
  assign _744_ = inv_4[18] ^ r_3[46] /*40188*/;
  assign sum_4[18] = _744_ ^ _743_ /*40187*/;
  assign _745_ = _744_ & _743_ /*40186*/;
  assign _746_ = inv_4[18] & r_3[46] /*40185*/;
  assign _747_ = _745_ | _746_ /*40184*/;
  assign _748_ = inv_4[19] ^ r_3[47] /*40182*/;
  assign sum_4[19] = _748_ ^ _747_ /*40181*/;
  assign _749_ = _748_ & _747_ /*40180*/;
  assign _750_ = inv_4[19] & r_3[47] /*40179*/;
  assign _751_ = _749_ | _750_ /*40178*/;
  assign _752_ = inv_4[20] ^ r_3[48] /*40176*/;
  assign sum_4[20] = _752_ ^ _751_ /*40175*/;
  assign _753_ = _752_ & _751_ /*40174*/;
  assign _754_ = inv_4[20] & r_3[48] /*40173*/;
  assign _755_ = _753_ | _754_ /*40172*/;
  assign _756_ = inv_4[21] ^ r_3[49] /*40170*/;
  assign sum_4[21] = _756_ ^ _755_ /*40169*/;
  assign _757_ = _756_ & _755_ /*40168*/;
  assign _758_ = inv_4[21] & r_3[49] /*40167*/;
  assign _759_ = _757_ | _758_ /*40166*/;
  assign _760_ = inv_4[22] ^ r_3[50] /*40164*/;
  assign sum_4[22] = _760_ ^ _759_ /*40163*/;
  assign _761_ = _760_ & _759_ /*40162*/;
  assign _762_ = inv_4[22] & r_3[50] /*40161*/;
  assign _763_ = _761_ | _762_ /*40160*/;
  assign _764_ = inv_4[23] ^ r_3[51] /*40158*/;
  assign sum_4[23] = _764_ ^ _763_ /*40157*/;
  assign _765_ = _764_ & _763_ /*40156*/;
  assign _766_ = inv_4[23] & r_3[51] /*40155*/;
  assign _767_ = _765_ | _766_ /*40154*/;
  assign _768_ = inv_4[24] ^ r_3[52] /*40152*/;
  assign sum_4[24] = _768_ ^ _767_ /*40151*/;
  assign _769_ = _768_ & _767_ /*40150*/;
  assign _770_ = inv_4[24] & r_3[52] /*40149*/;
  assign _771_ = _769_ | _770_ /*40148*/;
  assign _772_ = inv_4[25] ^ r_3[53] /*40146*/;
  assign sum_4[25] = _772_ ^ _771_ /*40145*/;
  assign _773_ = _772_ & _771_ /*40144*/;
  assign _774_ = inv_4[25] & r_3[53] /*40143*/;
  assign _775_ = _773_ | _774_ /*40142*/;
  assign _776_ = inv_4[26] ^ r_3[54] /*40140*/;
  assign sum_4[26] = _776_ ^ _775_ /*40139*/;
  assign _777_ = _776_ & _775_ /*40138*/;
  assign _778_ = inv_4[26] & r_3[54] /*40137*/;
  assign _779_ = _777_ | _778_ /*40136*/;
  assign _780_ = inv_4[27] ^ r_3[55] /*40134*/;
  assign sum_4[27] = _780_ ^ _779_ /*40133*/;
  assign _781_ = _780_ & _779_ /*40132*/;
  assign _782_ = inv_4[27] & r_3[55] /*40131*/;
  assign _783_ = _781_ | _782_ /*40130*/;
  assign _784_ = inv_4[28] ^ r_3[56] /*40128*/;
  assign sum_4[28] = _784_ ^ _783_ /*40127*/;
  assign _785_ = _784_ & _783_ /*40126*/;
  assign _786_ = inv_4[28] & r_3[56] /*40125*/;
  assign _787_ = _785_ | _786_ /*40124*/;
  assign _788_ = inv_4[29] ^ r_3[57] /*40122*/;
  assign sum_4[29] = _788_ ^ _787_ /*40121*/;
  assign _789_ = _788_ & _787_ /*40120*/;
  assign _790_ = inv_4[29] & r_3[57] /*40119*/;
  assign _791_ = _789_ | _790_ /*40118*/;
  assign _792_ = inv_4[30] ^ r_3[58] /*40116*/;
  assign sum_4[30] = _792_ ^ _791_ /*40115*/;
  assign _793_ = _792_ & _791_ /*40114*/;
  assign _794_ = inv_4[30] & r_3[58] /*40113*/;
  assign _795_ = _793_ | _794_ /*40112*/;
  assign _796_ = inv_4[31] ^ r_3[59] /*40110*/;
  assign sum_4[31] = _796_ ^ _795_ /*40109*/;
  assign _797_ = _796_ & _795_ /*40108*/;
  assign _798_ = inv_4[31] & r_3[59] /*40107*/;
  assign _799_ = _797_ | _798_ /*40106*/;
  assign q[28] = ~sum_4[31] /*40133*/;
  assign m_4[0] = r_3[28] /*40132*/;
  assign m_4[1] = r_3[29] /*40131*/;
  assign m_4[2] = r_3[30] /*40130*/;
  assign m_4[3] = r_3[31] /*40129*/;
  assign m_4[4] = r_3[32] /*40128*/;
  assign m_4[5] = r_3[33] /*40127*/;
  assign m_4[6] = r_3[34] /*40126*/;
  assign m_4[7] = r_3[35] /*40125*/;
  assign m_4[8] = r_3[36] /*40124*/;
  assign m_4[9] = r_3[37] /*40123*/;
  assign m_4[10] = r_3[38] /*40122*/;
  assign m_4[11] = r_3[39] /*40121*/;
  assign m_4[12] = r_3[40] /*40120*/;
  assign m_4[13] = r_3[41] /*40119*/;
  assign m_4[14] = r_3[42] /*40118*/;
  assign m_4[15] = r_3[43] /*40117*/;
  assign m_4[16] = r_3[44] /*40116*/;
  assign m_4[17] = r_3[45] /*40115*/;
  assign m_4[18] = r_3[46] /*40114*/;
  assign m_4[19] = r_3[47] /*40113*/;
  assign m_4[20] = r_3[48] /*40112*/;
  assign m_4[21] = r_3[49] /*40111*/;
  assign m_4[22] = r_3[50] /*40110*/;
  assign m_4[23] = r_3[51] /*40109*/;
  assign m_4[24] = r_3[52] /*40108*/;
  assign m_4[25] = r_3[53] /*40107*/;
  assign m_4[26] = r_3[54] /*40106*/;
  assign m_4[27] = r_3[55] /*40105*/;
  assign m_4[28] = r_3[56] /*40104*/;
  assign m_4[29] = r_3[57] /*40103*/;
  assign m_4[30] = r_3[58] /*40102*/;
  assign m_4[31] = r_3[59] /*40101*/;
  assign _800_ = ~q[28] /*40099*/;
  assign _801_ = sum_4[0] & q[28] /*40098*/;
  assign _802_ = m_4[0] & _800_ /*40097*/;
  assign r_4[28] = _802_ | _801_ /*40096*/;
  assign _803_ = ~q[28] /*40095*/;
  assign _804_ = sum_4[1] & q[28] /*40094*/;
  assign _805_ = m_4[1] & _803_ /*40093*/;
  assign r_4[29] = _805_ | _804_ /*40092*/;
  assign _806_ = ~q[28] /*40091*/;
  assign _807_ = sum_4[2] & q[28] /*40090*/;
  assign _808_ = m_4[2] & _806_ /*40089*/;
  assign r_4[30] = _808_ | _807_ /*40088*/;
  assign _809_ = ~q[28] /*40087*/;
  assign _810_ = sum_4[3] & q[28] /*40086*/;
  assign _811_ = m_4[3] & _809_ /*40085*/;
  assign r_4[31] = _811_ | _810_ /*40084*/;
  assign _812_ = ~q[28] /*40083*/;
  assign _813_ = sum_4[4] & q[28] /*40082*/;
  assign _814_ = m_4[4] & _812_ /*40081*/;
  assign r_4[32] = _814_ | _813_ /*40080*/;
  assign _815_ = ~q[28] /*40079*/;
  assign _816_ = sum_4[5] & q[28] /*40078*/;
  assign _817_ = m_4[5] & _815_ /*40077*/;
  assign r_4[33] = _817_ | _816_ /*40076*/;
  assign _818_ = ~q[28] /*40075*/;
  assign _819_ = sum_4[6] & q[28] /*40074*/;
  assign _820_ = m_4[6] & _818_ /*40073*/;
  assign r_4[34] = _820_ | _819_ /*40072*/;
  assign _821_ = ~q[28] /*40071*/;
  assign _822_ = sum_4[7] & q[28] /*40070*/;
  assign _823_ = m_4[7] & _821_ /*40069*/;
  assign r_4[35] = _823_ | _822_ /*40068*/;
  assign _824_ = ~q[28] /*40067*/;
  assign _825_ = sum_4[8] & q[28] /*40066*/;
  assign _826_ = m_4[8] & _824_ /*40065*/;
  assign r_4[36] = _826_ | _825_ /*40064*/;
  assign _827_ = ~q[28] /*40063*/;
  assign _828_ = sum_4[9] & q[28] /*40062*/;
  assign _829_ = m_4[9] & _827_ /*40061*/;
  assign r_4[37] = _829_ | _828_ /*40060*/;
  assign _830_ = ~q[28] /*40059*/;
  assign _831_ = sum_4[10] & q[28] /*40058*/;
  assign _832_ = m_4[10] & _830_ /*40057*/;
  assign r_4[38] = _832_ | _831_ /*40056*/;
  assign _833_ = ~q[28] /*40055*/;
  assign _834_ = sum_4[11] & q[28] /*40054*/;
  assign _835_ = m_4[11] & _833_ /*40053*/;
  assign r_4[39] = _835_ | _834_ /*40052*/;
  assign _836_ = ~q[28] /*40051*/;
  assign _837_ = sum_4[12] & q[28] /*40050*/;
  assign _838_ = m_4[12] & _836_ /*40049*/;
  assign r_4[40] = _838_ | _837_ /*40048*/;
  assign _839_ = ~q[28] /*40047*/;
  assign _840_ = sum_4[13] & q[28] /*40046*/;
  assign _841_ = m_4[13] & _839_ /*40045*/;
  assign r_4[41] = _841_ | _840_ /*40044*/;
  assign _842_ = ~q[28] /*40043*/;
  assign _843_ = sum_4[14] & q[28] /*40042*/;
  assign _844_ = m_4[14] & _842_ /*40041*/;
  assign r_4[42] = _844_ | _843_ /*40040*/;
  assign _845_ = ~q[28] /*40039*/;
  assign _846_ = sum_4[15] & q[28] /*40038*/;
  assign _847_ = m_4[15] & _845_ /*40037*/;
  assign r_4[43] = _847_ | _846_ /*40036*/;
  assign _848_ = ~q[28] /*40035*/;
  assign _849_ = sum_4[16] & q[28] /*40034*/;
  assign _850_ = m_4[16] & _848_ /*40033*/;
  assign r_4[44] = _850_ | _849_ /*40032*/;
  assign _851_ = ~q[28] /*40031*/;
  assign _852_ = sum_4[17] & q[28] /*40030*/;
  assign _853_ = m_4[17] & _851_ /*40029*/;
  assign r_4[45] = _853_ | _852_ /*40028*/;
  assign _854_ = ~q[28] /*40027*/;
  assign _855_ = sum_4[18] & q[28] /*40026*/;
  assign _856_ = m_4[18] & _854_ /*40025*/;
  assign r_4[46] = _856_ | _855_ /*40024*/;
  assign _857_ = ~q[28] /*40023*/;
  assign _858_ = sum_4[19] & q[28] /*40022*/;
  assign _859_ = m_4[19] & _857_ /*40021*/;
  assign r_4[47] = _859_ | _858_ /*40020*/;
  assign _860_ = ~q[28] /*40019*/;
  assign _861_ = sum_4[20] & q[28] /*40018*/;
  assign _862_ = m_4[20] & _860_ /*40017*/;
  assign r_4[48] = _862_ | _861_ /*40016*/;
  assign _863_ = ~q[28] /*40015*/;
  assign _864_ = sum_4[21] & q[28] /*40014*/;
  assign _865_ = m_4[21] & _863_ /*40013*/;
  assign r_4[49] = _865_ | _864_ /*40012*/;
  assign _866_ = ~q[28] /*40011*/;
  assign _867_ = sum_4[22] & q[28] /*40010*/;
  assign _868_ = m_4[22] & _866_ /*40009*/;
  assign r_4[50] = _868_ | _867_ /*40008*/;
  assign _869_ = ~q[28] /*40007*/;
  assign _870_ = sum_4[23] & q[28] /*40006*/;
  assign _871_ = m_4[23] & _869_ /*40005*/;
  assign r_4[51] = _871_ | _870_ /*40004*/;
  assign _872_ = ~q[28] /*40003*/;
  assign _873_ = sum_4[24] & q[28] /*40002*/;
  assign _874_ = m_4[24] & _872_ /*40001*/;
  assign r_4[52] = _874_ | _873_ /*40000*/;
  assign _875_ = ~q[28] /*39999*/;
  assign _876_ = sum_4[25] & q[28] /*39998*/;
  assign _877_ = m_4[25] & _875_ /*39997*/;
  assign r_4[53] = _877_ | _876_ /*39996*/;
  assign _878_ = ~q[28] /*39995*/;
  assign _879_ = sum_4[26] & q[28] /*39994*/;
  assign _880_ = m_4[26] & _878_ /*39993*/;
  assign r_4[54] = _880_ | _879_ /*39992*/;
  assign _881_ = ~q[28] /*39991*/;
  assign _882_ = sum_4[27] & q[28] /*39990*/;
  assign _883_ = m_4[27] & _881_ /*39989*/;
  assign r_4[55] = _883_ | _882_ /*39988*/;
  assign _884_ = ~q[28] /*39987*/;
  assign _885_ = sum_4[28] & q[28] /*39986*/;
  assign _886_ = m_4[28] & _884_ /*39985*/;
  assign r_4[56] = _886_ | _885_ /*39984*/;
  assign _887_ = ~q[28] /*39983*/;
  assign _888_ = sum_4[29] & q[28] /*39982*/;
  assign _889_ = m_4[29] & _887_ /*39981*/;
  assign r_4[57] = _889_ | _888_ /*39980*/;
  assign _890_ = ~q[28] /*39979*/;
  assign _891_ = sum_4[30] & q[28] /*39978*/;
  assign _892_ = m_4[30] & _890_ /*39977*/;
  assign r_4[58] = _892_ | _891_ /*39976*/;
  assign _893_ = ~q[28] /*39975*/;
  assign _894_ = sum_4[31] & q[28] /*39974*/;
  assign _895_ = m_4[31] & _893_ /*39973*/;
  assign r_4[59] = _895_ | _894_ /*39972*/;
assign r_4[0]= r_3[0] /*39971*/;
assign r_4[1]= r_3[1] /*39970*/;
assign r_4[2]= r_3[2] /*39969*/;
assign r_4[3]= r_3[3] /*39968*/;
assign r_4[4]= r_3[4] /*39967*/;
assign r_4[5]= r_3[5] /*39966*/;
assign r_4[6]= r_3[6] /*39965*/;
assign r_4[7]= r_3[7] /*39964*/;
assign r_4[8]= r_3[8] /*39963*/;
assign r_4[9]= r_3[9] /*39962*/;
assign r_4[10]= r_3[10] /*39961*/;
assign r_4[11]= r_3[11] /*39960*/;
assign r_4[12]= r_3[12] /*39959*/;
assign r_4[13]= r_3[13] /*39958*/;
assign r_4[14]= r_3[14] /*39957*/;
assign r_4[15]= r_3[15] /*39956*/;
assign r_4[16]= r_3[16] /*39955*/;
assign r_4[17]= r_3[17] /*39954*/;
assign r_4[18]= r_3[18] /*39953*/;
assign r_4[19]= r_3[19] /*39952*/;
assign r_4[20]= r_3[20] /*39951*/;
assign r_4[21]= r_3[21] /*39950*/;
assign r_4[22]= r_3[22] /*39949*/;
assign r_4[23]= r_3[23] /*39948*/;
assign r_4[24]= r_3[24] /*39947*/;
assign r_4[25]= r_3[25] /*39946*/;
assign r_4[26]= r_3[26] /*39945*/;
assign r_4[27]= r_3[27] /*39944*/;
  assign inv_5[0] = ~div[0] /*39880*/;
  assign inv_5[1] = ~div[1] /*39879*/;
  assign inv_5[2] = ~div[2] /*39878*/;
  assign inv_5[3] = ~div[3] /*39877*/;
  assign inv_5[4] = ~div[4] /*39876*/;
  assign inv_5[5] = ~div[5] /*39875*/;
  assign inv_5[6] = ~div[6] /*39874*/;
  assign inv_5[7] = ~div[7] /*39873*/;
  assign inv_5[8] = ~div[8] /*39872*/;
  assign inv_5[9] = ~div[9] /*39871*/;
  assign inv_5[10] = ~div[10] /*39870*/;
  assign inv_5[11] = ~div[11] /*39869*/;
  assign inv_5[12] = ~div[12] /*39868*/;
  assign inv_5[13] = ~div[13] /*39867*/;
  assign inv_5[14] = ~div[14] /*39866*/;
  assign inv_5[15] = ~div[15] /*39865*/;
  assign inv_5[16] = ~div[16] /*39864*/;
  assign inv_5[17] = ~div[17] /*39863*/;
  assign inv_5[18] = ~div[18] /*39862*/;
  assign inv_5[19] = ~div[19] /*39861*/;
  assign inv_5[20] = ~div[20] /*39860*/;
  assign inv_5[21] = ~div[21] /*39859*/;
  assign inv_5[22] = ~div[22] /*39858*/;
  assign inv_5[23] = ~div[23] /*39857*/;
  assign inv_5[24] = ~div[24] /*39856*/;
  assign inv_5[25] = ~div[25] /*39855*/;
  assign inv_5[26] = ~div[26] /*39854*/;
  assign inv_5[27] = ~div[27] /*39853*/;
  assign inv_5[28] = ~div[28] /*39852*/;
  assign inv_5[29] = ~div[29] /*39851*/;
  assign inv_5[30] = ~div[30] /*39850*/;
assign inv_5[31] = oneWire /*39849*/;
  assign _896_ = inv_5[0] ^ r_4[27] /*39847*/;
  assign sum_5[0] = _896_ ^ oneWire /*39846*/;
  assign _897_ = _896_ & oneWire /*39845*/;
  assign _898_ = inv_5[0] & r_4[27] /*39844*/;
  assign _899_ = _897_ | _898_ /*39843*/;
  assign _900_ = inv_5[1] ^ r_4[28] /*39842*/;
  assign sum_5[1] = _900_ ^ _899_ /*39841*/;
  assign _901_ = _900_ & _899_ /*39840*/;
  assign _902_ = inv_5[1] & r_4[28] /*39839*/;
  assign _903_ = _901_ | _902_ /*39838*/;
  assign _904_ = inv_5[2] ^ r_4[29] /*39836*/;
  assign sum_5[2] = _904_ ^ _903_ /*39835*/;
  assign _905_ = _904_ & _903_ /*39834*/;
  assign _906_ = inv_5[2] & r_4[29] /*39833*/;
  assign _907_ = _905_ | _906_ /*39832*/;
  assign _908_ = inv_5[3] ^ r_4[30] /*39830*/;
  assign sum_5[3] = _908_ ^ _907_ /*39829*/;
  assign _909_ = _908_ & _907_ /*39828*/;
  assign _910_ = inv_5[3] & r_4[30] /*39827*/;
  assign _911_ = _909_ | _910_ /*39826*/;
  assign _912_ = inv_5[4] ^ r_4[31] /*39824*/;
  assign sum_5[4] = _912_ ^ _911_ /*39823*/;
  assign _913_ = _912_ & _911_ /*39822*/;
  assign _914_ = inv_5[4] & r_4[31] /*39821*/;
  assign _915_ = _913_ | _914_ /*39820*/;
  assign _916_ = inv_5[5] ^ r_4[32] /*39818*/;
  assign sum_5[5] = _916_ ^ _915_ /*39817*/;
  assign _917_ = _916_ & _915_ /*39816*/;
  assign _918_ = inv_5[5] & r_4[32] /*39815*/;
  assign _919_ = _917_ | _918_ /*39814*/;
  assign _920_ = inv_5[6] ^ r_4[33] /*39812*/;
  assign sum_5[6] = _920_ ^ _919_ /*39811*/;
  assign _921_ = _920_ & _919_ /*39810*/;
  assign _922_ = inv_5[6] & r_4[33] /*39809*/;
  assign _923_ = _921_ | _922_ /*39808*/;
  assign _924_ = inv_5[7] ^ r_4[34] /*39806*/;
  assign sum_5[7] = _924_ ^ _923_ /*39805*/;
  assign _925_ = _924_ & _923_ /*39804*/;
  assign _926_ = inv_5[7] & r_4[34] /*39803*/;
  assign _927_ = _925_ | _926_ /*39802*/;
  assign _928_ = inv_5[8] ^ r_4[35] /*39800*/;
  assign sum_5[8] = _928_ ^ _927_ /*39799*/;
  assign _929_ = _928_ & _927_ /*39798*/;
  assign _930_ = inv_5[8] & r_4[35] /*39797*/;
  assign _931_ = _929_ | _930_ /*39796*/;
  assign _932_ = inv_5[9] ^ r_4[36] /*39794*/;
  assign sum_5[9] = _932_ ^ _931_ /*39793*/;
  assign _933_ = _932_ & _931_ /*39792*/;
  assign _934_ = inv_5[9] & r_4[36] /*39791*/;
  assign _935_ = _933_ | _934_ /*39790*/;
  assign _936_ = inv_5[10] ^ r_4[37] /*39788*/;
  assign sum_5[10] = _936_ ^ _935_ /*39787*/;
  assign _937_ = _936_ & _935_ /*39786*/;
  assign _938_ = inv_5[10] & r_4[37] /*39785*/;
  assign _939_ = _937_ | _938_ /*39784*/;
  assign _940_ = inv_5[11] ^ r_4[38] /*39782*/;
  assign sum_5[11] = _940_ ^ _939_ /*39781*/;
  assign _941_ = _940_ & _939_ /*39780*/;
  assign _942_ = inv_5[11] & r_4[38] /*39779*/;
  assign _943_ = _941_ | _942_ /*39778*/;
  assign _944_ = inv_5[12] ^ r_4[39] /*39776*/;
  assign sum_5[12] = _944_ ^ _943_ /*39775*/;
  assign _945_ = _944_ & _943_ /*39774*/;
  assign _946_ = inv_5[12] & r_4[39] /*39773*/;
  assign _947_ = _945_ | _946_ /*39772*/;
  assign _948_ = inv_5[13] ^ r_4[40] /*39770*/;
  assign sum_5[13] = _948_ ^ _947_ /*39769*/;
  assign _949_ = _948_ & _947_ /*39768*/;
  assign _950_ = inv_5[13] & r_4[40] /*39767*/;
  assign _951_ = _949_ | _950_ /*39766*/;
  assign _952_ = inv_5[14] ^ r_4[41] /*39764*/;
  assign sum_5[14] = _952_ ^ _951_ /*39763*/;
  assign _953_ = _952_ & _951_ /*39762*/;
  assign _954_ = inv_5[14] & r_4[41] /*39761*/;
  assign _955_ = _953_ | _954_ /*39760*/;
  assign _956_ = inv_5[15] ^ r_4[42] /*39758*/;
  assign sum_5[15] = _956_ ^ _955_ /*39757*/;
  assign _957_ = _956_ & _955_ /*39756*/;
  assign _958_ = inv_5[15] & r_4[42] /*39755*/;
  assign _959_ = _957_ | _958_ /*39754*/;
  assign _960_ = inv_5[16] ^ r_4[43] /*39752*/;
  assign sum_5[16] = _960_ ^ _959_ /*39751*/;
  assign _961_ = _960_ & _959_ /*39750*/;
  assign _962_ = inv_5[16] & r_4[43] /*39749*/;
  assign _963_ = _961_ | _962_ /*39748*/;
  assign _964_ = inv_5[17] ^ r_4[44] /*39746*/;
  assign sum_5[17] = _964_ ^ _963_ /*39745*/;
  assign _965_ = _964_ & _963_ /*39744*/;
  assign _966_ = inv_5[17] & r_4[44] /*39743*/;
  assign _967_ = _965_ | _966_ /*39742*/;
  assign _968_ = inv_5[18] ^ r_4[45] /*39740*/;
  assign sum_5[18] = _968_ ^ _967_ /*39739*/;
  assign _969_ = _968_ & _967_ /*39738*/;
  assign _970_ = inv_5[18] & r_4[45] /*39737*/;
  assign _971_ = _969_ | _970_ /*39736*/;
  assign _972_ = inv_5[19] ^ r_4[46] /*39734*/;
  assign sum_5[19] = _972_ ^ _971_ /*39733*/;
  assign _973_ = _972_ & _971_ /*39732*/;
  assign _974_ = inv_5[19] & r_4[46] /*39731*/;
  assign _975_ = _973_ | _974_ /*39730*/;
  assign _976_ = inv_5[20] ^ r_4[47] /*39728*/;
  assign sum_5[20] = _976_ ^ _975_ /*39727*/;
  assign _977_ = _976_ & _975_ /*39726*/;
  assign _978_ = inv_5[20] & r_4[47] /*39725*/;
  assign _979_ = _977_ | _978_ /*39724*/;
  assign _980_ = inv_5[21] ^ r_4[48] /*39722*/;
  assign sum_5[21] = _980_ ^ _979_ /*39721*/;
  assign _981_ = _980_ & _979_ /*39720*/;
  assign _982_ = inv_5[21] & r_4[48] /*39719*/;
  assign _983_ = _981_ | _982_ /*39718*/;
  assign _984_ = inv_5[22] ^ r_4[49] /*39716*/;
  assign sum_5[22] = _984_ ^ _983_ /*39715*/;
  assign _985_ = _984_ & _983_ /*39714*/;
  assign _986_ = inv_5[22] & r_4[49] /*39713*/;
  assign _987_ = _985_ | _986_ /*39712*/;
  assign _988_ = inv_5[23] ^ r_4[50] /*39710*/;
  assign sum_5[23] = _988_ ^ _987_ /*39709*/;
  assign _989_ = _988_ & _987_ /*39708*/;
  assign _990_ = inv_5[23] & r_4[50] /*39707*/;
  assign _991_ = _989_ | _990_ /*39706*/;
  assign _992_ = inv_5[24] ^ r_4[51] /*39704*/;
  assign sum_5[24] = _992_ ^ _991_ /*39703*/;
  assign _993_ = _992_ & _991_ /*39702*/;
  assign _994_ = inv_5[24] & r_4[51] /*39701*/;
  assign _995_ = _993_ | _994_ /*39700*/;
  assign _996_ = inv_5[25] ^ r_4[52] /*39698*/;
  assign sum_5[25] = _996_ ^ _995_ /*39697*/;
  assign _997_ = _996_ & _995_ /*39696*/;
  assign _998_ = inv_5[25] & r_4[52] /*39695*/;
  assign _999_ = _997_ | _998_ /*39694*/;
  assign _1000_ = inv_5[26] ^ r_4[53] /*39692*/;
  assign sum_5[26] = _1000_ ^ _999_ /*39691*/;
  assign _1001_ = _1000_ & _999_ /*39690*/;
  assign _1002_ = inv_5[26] & r_4[53] /*39689*/;
  assign _1003_ = _1001_ | _1002_ /*39688*/;
  assign _1004_ = inv_5[27] ^ r_4[54] /*39686*/;
  assign sum_5[27] = _1004_ ^ _1003_ /*39685*/;
  assign _1005_ = _1004_ & _1003_ /*39684*/;
  assign _1006_ = inv_5[27] & r_4[54] /*39683*/;
  assign _1007_ = _1005_ | _1006_ /*39682*/;
  assign _1008_ = inv_5[28] ^ r_4[55] /*39680*/;
  assign sum_5[28] = _1008_ ^ _1007_ /*39679*/;
  assign _1009_ = _1008_ & _1007_ /*39678*/;
  assign _1010_ = inv_5[28] & r_4[55] /*39677*/;
  assign _1011_ = _1009_ | _1010_ /*39676*/;
  assign _1012_ = inv_5[29] ^ r_4[56] /*39674*/;
  assign sum_5[29] = _1012_ ^ _1011_ /*39673*/;
  assign _1013_ = _1012_ & _1011_ /*39672*/;
  assign _1014_ = inv_5[29] & r_4[56] /*39671*/;
  assign _1015_ = _1013_ | _1014_ /*39670*/;
  assign _1016_ = inv_5[30] ^ r_4[57] /*39668*/;
  assign sum_5[30] = _1016_ ^ _1015_ /*39667*/;
  assign _1017_ = _1016_ & _1015_ /*39666*/;
  assign _1018_ = inv_5[30] & r_4[57] /*39665*/;
  assign _1019_ = _1017_ | _1018_ /*39664*/;
  assign _1020_ = inv_5[31] ^ r_4[58] /*39662*/;
  assign sum_5[31] = _1020_ ^ _1019_ /*39661*/;
  assign _1021_ = _1020_ & _1019_ /*39660*/;
  assign _1022_ = inv_5[31] & r_4[58] /*39659*/;
  assign _1023_ = _1021_ | _1022_ /*39658*/;
  assign q[27] = ~sum_5[31] /*39685*/;
  assign m_5[0] = r_4[27] /*39684*/;
  assign m_5[1] = r_4[28] /*39683*/;
  assign m_5[2] = r_4[29] /*39682*/;
  assign m_5[3] = r_4[30] /*39681*/;
  assign m_5[4] = r_4[31] /*39680*/;
  assign m_5[5] = r_4[32] /*39679*/;
  assign m_5[6] = r_4[33] /*39678*/;
  assign m_5[7] = r_4[34] /*39677*/;
  assign m_5[8] = r_4[35] /*39676*/;
  assign m_5[9] = r_4[36] /*39675*/;
  assign m_5[10] = r_4[37] /*39674*/;
  assign m_5[11] = r_4[38] /*39673*/;
  assign m_5[12] = r_4[39] /*39672*/;
  assign m_5[13] = r_4[40] /*39671*/;
  assign m_5[14] = r_4[41] /*39670*/;
  assign m_5[15] = r_4[42] /*39669*/;
  assign m_5[16] = r_4[43] /*39668*/;
  assign m_5[17] = r_4[44] /*39667*/;
  assign m_5[18] = r_4[45] /*39666*/;
  assign m_5[19] = r_4[46] /*39665*/;
  assign m_5[20] = r_4[47] /*39664*/;
  assign m_5[21] = r_4[48] /*39663*/;
  assign m_5[22] = r_4[49] /*39662*/;
  assign m_5[23] = r_4[50] /*39661*/;
  assign m_5[24] = r_4[51] /*39660*/;
  assign m_5[25] = r_4[52] /*39659*/;
  assign m_5[26] = r_4[53] /*39658*/;
  assign m_5[27] = r_4[54] /*39657*/;
  assign m_5[28] = r_4[55] /*39656*/;
  assign m_5[29] = r_4[56] /*39655*/;
  assign m_5[30] = r_4[57] /*39654*/;
  assign m_5[31] = r_4[58] /*39653*/;
  assign _1024_ = ~q[27] /*39651*/;
  assign _1025_ = sum_5[0] & q[27] /*39650*/;
  assign _1026_ = m_5[0] & _1024_ /*39649*/;
  assign r_5[27] = _1026_ | _1025_ /*39648*/;
  assign _1027_ = ~q[27] /*39647*/;
  assign _1028_ = sum_5[1] & q[27] /*39646*/;
  assign _1029_ = m_5[1] & _1027_ /*39645*/;
  assign r_5[28] = _1029_ | _1028_ /*39644*/;
  assign _1030_ = ~q[27] /*39643*/;
  assign _1031_ = sum_5[2] & q[27] /*39642*/;
  assign _1032_ = m_5[2] & _1030_ /*39641*/;
  assign r_5[29] = _1032_ | _1031_ /*39640*/;
  assign _1033_ = ~q[27] /*39639*/;
  assign _1034_ = sum_5[3] & q[27] /*39638*/;
  assign _1035_ = m_5[3] & _1033_ /*39637*/;
  assign r_5[30] = _1035_ | _1034_ /*39636*/;
  assign _1036_ = ~q[27] /*39635*/;
  assign _1037_ = sum_5[4] & q[27] /*39634*/;
  assign _1038_ = m_5[4] & _1036_ /*39633*/;
  assign r_5[31] = _1038_ | _1037_ /*39632*/;
  assign _1039_ = ~q[27] /*39631*/;
  assign _1040_ = sum_5[5] & q[27] /*39630*/;
  assign _1041_ = m_5[5] & _1039_ /*39629*/;
  assign r_5[32] = _1041_ | _1040_ /*39628*/;
  assign _1042_ = ~q[27] /*39627*/;
  assign _1043_ = sum_5[6] & q[27] /*39626*/;
  assign _1044_ = m_5[6] & _1042_ /*39625*/;
  assign r_5[33] = _1044_ | _1043_ /*39624*/;
  assign _1045_ = ~q[27] /*39623*/;
  assign _1046_ = sum_5[7] & q[27] /*39622*/;
  assign _1047_ = m_5[7] & _1045_ /*39621*/;
  assign r_5[34] = _1047_ | _1046_ /*39620*/;
  assign _1048_ = ~q[27] /*39619*/;
  assign _1049_ = sum_5[8] & q[27] /*39618*/;
  assign _1050_ = m_5[8] & _1048_ /*39617*/;
  assign r_5[35] = _1050_ | _1049_ /*39616*/;
  assign _1051_ = ~q[27] /*39615*/;
  assign _1052_ = sum_5[9] & q[27] /*39614*/;
  assign _1053_ = m_5[9] & _1051_ /*39613*/;
  assign r_5[36] = _1053_ | _1052_ /*39612*/;
  assign _1054_ = ~q[27] /*39611*/;
  assign _1055_ = sum_5[10] & q[27] /*39610*/;
  assign _1056_ = m_5[10] & _1054_ /*39609*/;
  assign r_5[37] = _1056_ | _1055_ /*39608*/;
  assign _1057_ = ~q[27] /*39607*/;
  assign _1058_ = sum_5[11] & q[27] /*39606*/;
  assign _1059_ = m_5[11] & _1057_ /*39605*/;
  assign r_5[38] = _1059_ | _1058_ /*39604*/;
  assign _1060_ = ~q[27] /*39603*/;
  assign _1061_ = sum_5[12] & q[27] /*39602*/;
  assign _1062_ = m_5[12] & _1060_ /*39601*/;
  assign r_5[39] = _1062_ | _1061_ /*39600*/;
  assign _1063_ = ~q[27] /*39599*/;
  assign _1064_ = sum_5[13] & q[27] /*39598*/;
  assign _1065_ = m_5[13] & _1063_ /*39597*/;
  assign r_5[40] = _1065_ | _1064_ /*39596*/;
  assign _1066_ = ~q[27] /*39595*/;
  assign _1067_ = sum_5[14] & q[27] /*39594*/;
  assign _1068_ = m_5[14] & _1066_ /*39593*/;
  assign r_5[41] = _1068_ | _1067_ /*39592*/;
  assign _1069_ = ~q[27] /*39591*/;
  assign _1070_ = sum_5[15] & q[27] /*39590*/;
  assign _1071_ = m_5[15] & _1069_ /*39589*/;
  assign r_5[42] = _1071_ | _1070_ /*39588*/;
  assign _1072_ = ~q[27] /*39587*/;
  assign _1073_ = sum_5[16] & q[27] /*39586*/;
  assign _1074_ = m_5[16] & _1072_ /*39585*/;
  assign r_5[43] = _1074_ | _1073_ /*39584*/;
  assign _1075_ = ~q[27] /*39583*/;
  assign _1076_ = sum_5[17] & q[27] /*39582*/;
  assign _1077_ = m_5[17] & _1075_ /*39581*/;
  assign r_5[44] = _1077_ | _1076_ /*39580*/;
  assign _1078_ = ~q[27] /*39579*/;
  assign _1079_ = sum_5[18] & q[27] /*39578*/;
  assign _1080_ = m_5[18] & _1078_ /*39577*/;
  assign r_5[45] = _1080_ | _1079_ /*39576*/;
  assign _1081_ = ~q[27] /*39575*/;
  assign _1082_ = sum_5[19] & q[27] /*39574*/;
  assign _1083_ = m_5[19] & _1081_ /*39573*/;
  assign r_5[46] = _1083_ | _1082_ /*39572*/;
  assign _1084_ = ~q[27] /*39571*/;
  assign _1085_ = sum_5[20] & q[27] /*39570*/;
  assign _1086_ = m_5[20] & _1084_ /*39569*/;
  assign r_5[47] = _1086_ | _1085_ /*39568*/;
  assign _1087_ = ~q[27] /*39567*/;
  assign _1088_ = sum_5[21] & q[27] /*39566*/;
  assign _1089_ = m_5[21] & _1087_ /*39565*/;
  assign r_5[48] = _1089_ | _1088_ /*39564*/;
  assign _1090_ = ~q[27] /*39563*/;
  assign _1091_ = sum_5[22] & q[27] /*39562*/;
  assign _1092_ = m_5[22] & _1090_ /*39561*/;
  assign r_5[49] = _1092_ | _1091_ /*39560*/;
  assign _1093_ = ~q[27] /*39559*/;
  assign _1094_ = sum_5[23] & q[27] /*39558*/;
  assign _1095_ = m_5[23] & _1093_ /*39557*/;
  assign r_5[50] = _1095_ | _1094_ /*39556*/;
  assign _1096_ = ~q[27] /*39555*/;
  assign _1097_ = sum_5[24] & q[27] /*39554*/;
  assign _1098_ = m_5[24] & _1096_ /*39553*/;
  assign r_5[51] = _1098_ | _1097_ /*39552*/;
  assign _1099_ = ~q[27] /*39551*/;
  assign _1100_ = sum_5[25] & q[27] /*39550*/;
  assign _1101_ = m_5[25] & _1099_ /*39549*/;
  assign r_5[52] = _1101_ | _1100_ /*39548*/;
  assign _1102_ = ~q[27] /*39547*/;
  assign _1103_ = sum_5[26] & q[27] /*39546*/;
  assign _1104_ = m_5[26] & _1102_ /*39545*/;
  assign r_5[53] = _1104_ | _1103_ /*39544*/;
  assign _1105_ = ~q[27] /*39543*/;
  assign _1106_ = sum_5[27] & q[27] /*39542*/;
  assign _1107_ = m_5[27] & _1105_ /*39541*/;
  assign r_5[54] = _1107_ | _1106_ /*39540*/;
  assign _1108_ = ~q[27] /*39539*/;
  assign _1109_ = sum_5[28] & q[27] /*39538*/;
  assign _1110_ = m_5[28] & _1108_ /*39537*/;
  assign r_5[55] = _1110_ | _1109_ /*39536*/;
  assign _1111_ = ~q[27] /*39535*/;
  assign _1112_ = sum_5[29] & q[27] /*39534*/;
  assign _1113_ = m_5[29] & _1111_ /*39533*/;
  assign r_5[56] = _1113_ | _1112_ /*39532*/;
  assign _1114_ = ~q[27] /*39531*/;
  assign _1115_ = sum_5[30] & q[27] /*39530*/;
  assign _1116_ = m_5[30] & _1114_ /*39529*/;
  assign r_5[57] = _1116_ | _1115_ /*39528*/;
  assign _1117_ = ~q[27] /*39527*/;
  assign _1118_ = sum_5[31] & q[27] /*39526*/;
  assign _1119_ = m_5[31] & _1117_ /*39525*/;
  assign r_5[58] = _1119_ | _1118_ /*39524*/;
assign r_5[0]= r_4[0] /*39523*/;
assign r_5[1]= r_4[1] /*39522*/;
assign r_5[2]= r_4[2] /*39521*/;
assign r_5[3]= r_4[3] /*39520*/;
assign r_5[4]= r_4[4] /*39519*/;
assign r_5[5]= r_4[5] /*39518*/;
assign r_5[6]= r_4[6] /*39517*/;
assign r_5[7]= r_4[7] /*39516*/;
assign r_5[8]= r_4[8] /*39515*/;
assign r_5[9]= r_4[9] /*39514*/;
assign r_5[10]= r_4[10] /*39513*/;
assign r_5[11]= r_4[11] /*39512*/;
assign r_5[12]= r_4[12] /*39511*/;
assign r_5[13]= r_4[13] /*39510*/;
assign r_5[14]= r_4[14] /*39509*/;
assign r_5[15]= r_4[15] /*39508*/;
assign r_5[16]= r_4[16] /*39507*/;
assign r_5[17]= r_4[17] /*39506*/;
assign r_5[18]= r_4[18] /*39505*/;
assign r_5[19]= r_4[19] /*39504*/;
assign r_5[20]= r_4[20] /*39503*/;
assign r_5[21]= r_4[21] /*39502*/;
assign r_5[22]= r_4[22] /*39501*/;
assign r_5[23]= r_4[23] /*39500*/;
assign r_5[24]= r_4[24] /*39499*/;
assign r_5[25]= r_4[25] /*39498*/;
assign r_5[26]= r_4[26] /*39497*/;
  assign inv_6[0] = ~div[0] /*39432*/;
  assign inv_6[1] = ~div[1] /*39431*/;
  assign inv_6[2] = ~div[2] /*39430*/;
  assign inv_6[3] = ~div[3] /*39429*/;
  assign inv_6[4] = ~div[4] /*39428*/;
  assign inv_6[5] = ~div[5] /*39427*/;
  assign inv_6[6] = ~div[6] /*39426*/;
  assign inv_6[7] = ~div[7] /*39425*/;
  assign inv_6[8] = ~div[8] /*39424*/;
  assign inv_6[9] = ~div[9] /*39423*/;
  assign inv_6[10] = ~div[10] /*39422*/;
  assign inv_6[11] = ~div[11] /*39421*/;
  assign inv_6[12] = ~div[12] /*39420*/;
  assign inv_6[13] = ~div[13] /*39419*/;
  assign inv_6[14] = ~div[14] /*39418*/;
  assign inv_6[15] = ~div[15] /*39417*/;
  assign inv_6[16] = ~div[16] /*39416*/;
  assign inv_6[17] = ~div[17] /*39415*/;
  assign inv_6[18] = ~div[18] /*39414*/;
  assign inv_6[19] = ~div[19] /*39413*/;
  assign inv_6[20] = ~div[20] /*39412*/;
  assign inv_6[21] = ~div[21] /*39411*/;
  assign inv_6[22] = ~div[22] /*39410*/;
  assign inv_6[23] = ~div[23] /*39409*/;
  assign inv_6[24] = ~div[24] /*39408*/;
  assign inv_6[25] = ~div[25] /*39407*/;
  assign inv_6[26] = ~div[26] /*39406*/;
  assign inv_6[27] = ~div[27] /*39405*/;
  assign inv_6[28] = ~div[28] /*39404*/;
  assign inv_6[29] = ~div[29] /*39403*/;
  assign inv_6[30] = ~div[30] /*39402*/;
assign inv_6[31] = oneWire /*39401*/;
  assign _1120_ = inv_6[0] ^ r_5[26] /*39399*/;
  assign sum_6[0] = _1120_ ^ oneWire /*39398*/;
  assign _1121_ = _1120_ & oneWire /*39397*/;
  assign _1122_ = inv_6[0] & r_5[26] /*39396*/;
  assign _1123_ = _1121_ | _1122_ /*39395*/;
  assign _1124_ = inv_6[1] ^ r_5[27] /*39394*/;
  assign sum_6[1] = _1124_ ^ _1123_ /*39393*/;
  assign _1125_ = _1124_ & _1123_ /*39392*/;
  assign _1126_ = inv_6[1] & r_5[27] /*39391*/;
  assign _1127_ = _1125_ | _1126_ /*39390*/;
  assign _1128_ = inv_6[2] ^ r_5[28] /*39388*/;
  assign sum_6[2] = _1128_ ^ _1127_ /*39387*/;
  assign _1129_ = _1128_ & _1127_ /*39386*/;
  assign _1130_ = inv_6[2] & r_5[28] /*39385*/;
  assign _1131_ = _1129_ | _1130_ /*39384*/;
  assign _1132_ = inv_6[3] ^ r_5[29] /*39382*/;
  assign sum_6[3] = _1132_ ^ _1131_ /*39381*/;
  assign _1133_ = _1132_ & _1131_ /*39380*/;
  assign _1134_ = inv_6[3] & r_5[29] /*39379*/;
  assign _1135_ = _1133_ | _1134_ /*39378*/;
  assign _1136_ = inv_6[4] ^ r_5[30] /*39376*/;
  assign sum_6[4] = _1136_ ^ _1135_ /*39375*/;
  assign _1137_ = _1136_ & _1135_ /*39374*/;
  assign _1138_ = inv_6[4] & r_5[30] /*39373*/;
  assign _1139_ = _1137_ | _1138_ /*39372*/;
  assign _1140_ = inv_6[5] ^ r_5[31] /*39370*/;
  assign sum_6[5] = _1140_ ^ _1139_ /*39369*/;
  assign _1141_ = _1140_ & _1139_ /*39368*/;
  assign _1142_ = inv_6[5] & r_5[31] /*39367*/;
  assign _1143_ = _1141_ | _1142_ /*39366*/;
  assign _1144_ = inv_6[6] ^ r_5[32] /*39364*/;
  assign sum_6[6] = _1144_ ^ _1143_ /*39363*/;
  assign _1145_ = _1144_ & _1143_ /*39362*/;
  assign _1146_ = inv_6[6] & r_5[32] /*39361*/;
  assign _1147_ = _1145_ | _1146_ /*39360*/;
  assign _1148_ = inv_6[7] ^ r_5[33] /*39358*/;
  assign sum_6[7] = _1148_ ^ _1147_ /*39357*/;
  assign _1149_ = _1148_ & _1147_ /*39356*/;
  assign _1150_ = inv_6[7] & r_5[33] /*39355*/;
  assign _1151_ = _1149_ | _1150_ /*39354*/;
  assign _1152_ = inv_6[8] ^ r_5[34] /*39352*/;
  assign sum_6[8] = _1152_ ^ _1151_ /*39351*/;
  assign _1153_ = _1152_ & _1151_ /*39350*/;
  assign _1154_ = inv_6[8] & r_5[34] /*39349*/;
  assign _1155_ = _1153_ | _1154_ /*39348*/;
  assign _1156_ = inv_6[9] ^ r_5[35] /*39346*/;
  assign sum_6[9] = _1156_ ^ _1155_ /*39345*/;
  assign _1157_ = _1156_ & _1155_ /*39344*/;
  assign _1158_ = inv_6[9] & r_5[35] /*39343*/;
  assign _1159_ = _1157_ | _1158_ /*39342*/;
  assign _1160_ = inv_6[10] ^ r_5[36] /*39340*/;
  assign sum_6[10] = _1160_ ^ _1159_ /*39339*/;
  assign _1161_ = _1160_ & _1159_ /*39338*/;
  assign _1162_ = inv_6[10] & r_5[36] /*39337*/;
  assign _1163_ = _1161_ | _1162_ /*39336*/;
  assign _1164_ = inv_6[11] ^ r_5[37] /*39334*/;
  assign sum_6[11] = _1164_ ^ _1163_ /*39333*/;
  assign _1165_ = _1164_ & _1163_ /*39332*/;
  assign _1166_ = inv_6[11] & r_5[37] /*39331*/;
  assign _1167_ = _1165_ | _1166_ /*39330*/;
  assign _1168_ = inv_6[12] ^ r_5[38] /*39328*/;
  assign sum_6[12] = _1168_ ^ _1167_ /*39327*/;
  assign _1169_ = _1168_ & _1167_ /*39326*/;
  assign _1170_ = inv_6[12] & r_5[38] /*39325*/;
  assign _1171_ = _1169_ | _1170_ /*39324*/;
  assign _1172_ = inv_6[13] ^ r_5[39] /*39322*/;
  assign sum_6[13] = _1172_ ^ _1171_ /*39321*/;
  assign _1173_ = _1172_ & _1171_ /*39320*/;
  assign _1174_ = inv_6[13] & r_5[39] /*39319*/;
  assign _1175_ = _1173_ | _1174_ /*39318*/;
  assign _1176_ = inv_6[14] ^ r_5[40] /*39316*/;
  assign sum_6[14] = _1176_ ^ _1175_ /*39315*/;
  assign _1177_ = _1176_ & _1175_ /*39314*/;
  assign _1178_ = inv_6[14] & r_5[40] /*39313*/;
  assign _1179_ = _1177_ | _1178_ /*39312*/;
  assign _1180_ = inv_6[15] ^ r_5[41] /*39310*/;
  assign sum_6[15] = _1180_ ^ _1179_ /*39309*/;
  assign _1181_ = _1180_ & _1179_ /*39308*/;
  assign _1182_ = inv_6[15] & r_5[41] /*39307*/;
  assign _1183_ = _1181_ | _1182_ /*39306*/;
  assign _1184_ = inv_6[16] ^ r_5[42] /*39304*/;
  assign sum_6[16] = _1184_ ^ _1183_ /*39303*/;
  assign _1185_ = _1184_ & _1183_ /*39302*/;
  assign _1186_ = inv_6[16] & r_5[42] /*39301*/;
  assign _1187_ = _1185_ | _1186_ /*39300*/;
  assign _1188_ = inv_6[17] ^ r_5[43] /*39298*/;
  assign sum_6[17] = _1188_ ^ _1187_ /*39297*/;
  assign _1189_ = _1188_ & _1187_ /*39296*/;
  assign _1190_ = inv_6[17] & r_5[43] /*39295*/;
  assign _1191_ = _1189_ | _1190_ /*39294*/;
  assign _1192_ = inv_6[18] ^ r_5[44] /*39292*/;
  assign sum_6[18] = _1192_ ^ _1191_ /*39291*/;
  assign _1193_ = _1192_ & _1191_ /*39290*/;
  assign _1194_ = inv_6[18] & r_5[44] /*39289*/;
  assign _1195_ = _1193_ | _1194_ /*39288*/;
  assign _1196_ = inv_6[19] ^ r_5[45] /*39286*/;
  assign sum_6[19] = _1196_ ^ _1195_ /*39285*/;
  assign _1197_ = _1196_ & _1195_ /*39284*/;
  assign _1198_ = inv_6[19] & r_5[45] /*39283*/;
  assign _1199_ = _1197_ | _1198_ /*39282*/;
  assign _1200_ = inv_6[20] ^ r_5[46] /*39280*/;
  assign sum_6[20] = _1200_ ^ _1199_ /*39279*/;
  assign _1201_ = _1200_ & _1199_ /*39278*/;
  assign _1202_ = inv_6[20] & r_5[46] /*39277*/;
  assign _1203_ = _1201_ | _1202_ /*39276*/;
  assign _1204_ = inv_6[21] ^ r_5[47] /*39274*/;
  assign sum_6[21] = _1204_ ^ _1203_ /*39273*/;
  assign _1205_ = _1204_ & _1203_ /*39272*/;
  assign _1206_ = inv_6[21] & r_5[47] /*39271*/;
  assign _1207_ = _1205_ | _1206_ /*39270*/;
  assign _1208_ = inv_6[22] ^ r_5[48] /*39268*/;
  assign sum_6[22] = _1208_ ^ _1207_ /*39267*/;
  assign _1209_ = _1208_ & _1207_ /*39266*/;
  assign _1210_ = inv_6[22] & r_5[48] /*39265*/;
  assign _1211_ = _1209_ | _1210_ /*39264*/;
  assign _1212_ = inv_6[23] ^ r_5[49] /*39262*/;
  assign sum_6[23] = _1212_ ^ _1211_ /*39261*/;
  assign _1213_ = _1212_ & _1211_ /*39260*/;
  assign _1214_ = inv_6[23] & r_5[49] /*39259*/;
  assign _1215_ = _1213_ | _1214_ /*39258*/;
  assign _1216_ = inv_6[24] ^ r_5[50] /*39256*/;
  assign sum_6[24] = _1216_ ^ _1215_ /*39255*/;
  assign _1217_ = _1216_ & _1215_ /*39254*/;
  assign _1218_ = inv_6[24] & r_5[50] /*39253*/;
  assign _1219_ = _1217_ | _1218_ /*39252*/;
  assign _1220_ = inv_6[25] ^ r_5[51] /*39250*/;
  assign sum_6[25] = _1220_ ^ _1219_ /*39249*/;
  assign _1221_ = _1220_ & _1219_ /*39248*/;
  assign _1222_ = inv_6[25] & r_5[51] /*39247*/;
  assign _1223_ = _1221_ | _1222_ /*39246*/;
  assign _1224_ = inv_6[26] ^ r_5[52] /*39244*/;
  assign sum_6[26] = _1224_ ^ _1223_ /*39243*/;
  assign _1225_ = _1224_ & _1223_ /*39242*/;
  assign _1226_ = inv_6[26] & r_5[52] /*39241*/;
  assign _1227_ = _1225_ | _1226_ /*39240*/;
  assign _1228_ = inv_6[27] ^ r_5[53] /*39238*/;
  assign sum_6[27] = _1228_ ^ _1227_ /*39237*/;
  assign _1229_ = _1228_ & _1227_ /*39236*/;
  assign _1230_ = inv_6[27] & r_5[53] /*39235*/;
  assign _1231_ = _1229_ | _1230_ /*39234*/;
  assign _1232_ = inv_6[28] ^ r_5[54] /*39232*/;
  assign sum_6[28] = _1232_ ^ _1231_ /*39231*/;
  assign _1233_ = _1232_ & _1231_ /*39230*/;
  assign _1234_ = inv_6[28] & r_5[54] /*39229*/;
  assign _1235_ = _1233_ | _1234_ /*39228*/;
  assign _1236_ = inv_6[29] ^ r_5[55] /*39226*/;
  assign sum_6[29] = _1236_ ^ _1235_ /*39225*/;
  assign _1237_ = _1236_ & _1235_ /*39224*/;
  assign _1238_ = inv_6[29] & r_5[55] /*39223*/;
  assign _1239_ = _1237_ | _1238_ /*39222*/;
  assign _1240_ = inv_6[30] ^ r_5[56] /*39220*/;
  assign sum_6[30] = _1240_ ^ _1239_ /*39219*/;
  assign _1241_ = _1240_ & _1239_ /*39218*/;
  assign _1242_ = inv_6[30] & r_5[56] /*39217*/;
  assign _1243_ = _1241_ | _1242_ /*39216*/;
  assign _1244_ = inv_6[31] ^ r_5[57] /*39214*/;
  assign sum_6[31] = _1244_ ^ _1243_ /*39213*/;
  assign _1245_ = _1244_ & _1243_ /*39212*/;
  assign _1246_ = inv_6[31] & r_5[57] /*39211*/;
  assign _1247_ = _1245_ | _1246_ /*39210*/;
  assign q[26] = ~sum_6[31] /*39237*/;
  assign m_6[0] = r_5[26] /*39236*/;
  assign m_6[1] = r_5[27] /*39235*/;
  assign m_6[2] = r_5[28] /*39234*/;
  assign m_6[3] = r_5[29] /*39233*/;
  assign m_6[4] = r_5[30] /*39232*/;
  assign m_6[5] = r_5[31] /*39231*/;
  assign m_6[6] = r_5[32] /*39230*/;
  assign m_6[7] = r_5[33] /*39229*/;
  assign m_6[8] = r_5[34] /*39228*/;
  assign m_6[9] = r_5[35] /*39227*/;
  assign m_6[10] = r_5[36] /*39226*/;
  assign m_6[11] = r_5[37] /*39225*/;
  assign m_6[12] = r_5[38] /*39224*/;
  assign m_6[13] = r_5[39] /*39223*/;
  assign m_6[14] = r_5[40] /*39222*/;
  assign m_6[15] = r_5[41] /*39221*/;
  assign m_6[16] = r_5[42] /*39220*/;
  assign m_6[17] = r_5[43] /*39219*/;
  assign m_6[18] = r_5[44] /*39218*/;
  assign m_6[19] = r_5[45] /*39217*/;
  assign m_6[20] = r_5[46] /*39216*/;
  assign m_6[21] = r_5[47] /*39215*/;
  assign m_6[22] = r_5[48] /*39214*/;
  assign m_6[23] = r_5[49] /*39213*/;
  assign m_6[24] = r_5[50] /*39212*/;
  assign m_6[25] = r_5[51] /*39211*/;
  assign m_6[26] = r_5[52] /*39210*/;
  assign m_6[27] = r_5[53] /*39209*/;
  assign m_6[28] = r_5[54] /*39208*/;
  assign m_6[29] = r_5[55] /*39207*/;
  assign m_6[30] = r_5[56] /*39206*/;
  assign m_6[31] = r_5[57] /*39205*/;
  assign _1248_ = ~q[26] /*39203*/;
  assign _1249_ = sum_6[0] & q[26] /*39202*/;
  assign _1250_ = m_6[0] & _1248_ /*39201*/;
  assign r_6[26] = _1250_ | _1249_ /*39200*/;
  assign _1251_ = ~q[26] /*39199*/;
  assign _1252_ = sum_6[1] & q[26] /*39198*/;
  assign _1253_ = m_6[1] & _1251_ /*39197*/;
  assign r_6[27] = _1253_ | _1252_ /*39196*/;
  assign _1254_ = ~q[26] /*39195*/;
  assign _1255_ = sum_6[2] & q[26] /*39194*/;
  assign _1256_ = m_6[2] & _1254_ /*39193*/;
  assign r_6[28] = _1256_ | _1255_ /*39192*/;
  assign _1257_ = ~q[26] /*39191*/;
  assign _1258_ = sum_6[3] & q[26] /*39190*/;
  assign _1259_ = m_6[3] & _1257_ /*39189*/;
  assign r_6[29] = _1259_ | _1258_ /*39188*/;
  assign _1260_ = ~q[26] /*39187*/;
  assign _1261_ = sum_6[4] & q[26] /*39186*/;
  assign _1262_ = m_6[4] & _1260_ /*39185*/;
  assign r_6[30] = _1262_ | _1261_ /*39184*/;
  assign _1263_ = ~q[26] /*39183*/;
  assign _1264_ = sum_6[5] & q[26] /*39182*/;
  assign _1265_ = m_6[5] & _1263_ /*39181*/;
  assign r_6[31] = _1265_ | _1264_ /*39180*/;
  assign _1266_ = ~q[26] /*39179*/;
  assign _1267_ = sum_6[6] & q[26] /*39178*/;
  assign _1268_ = m_6[6] & _1266_ /*39177*/;
  assign r_6[32] = _1268_ | _1267_ /*39176*/;
  assign _1269_ = ~q[26] /*39175*/;
  assign _1270_ = sum_6[7] & q[26] /*39174*/;
  assign _1271_ = m_6[7] & _1269_ /*39173*/;
  assign r_6[33] = _1271_ | _1270_ /*39172*/;
  assign _1272_ = ~q[26] /*39171*/;
  assign _1273_ = sum_6[8] & q[26] /*39170*/;
  assign _1274_ = m_6[8] & _1272_ /*39169*/;
  assign r_6[34] = _1274_ | _1273_ /*39168*/;
  assign _1275_ = ~q[26] /*39167*/;
  assign _1276_ = sum_6[9] & q[26] /*39166*/;
  assign _1277_ = m_6[9] & _1275_ /*39165*/;
  assign r_6[35] = _1277_ | _1276_ /*39164*/;
  assign _1278_ = ~q[26] /*39163*/;
  assign _1279_ = sum_6[10] & q[26] /*39162*/;
  assign _1280_ = m_6[10] & _1278_ /*39161*/;
  assign r_6[36] = _1280_ | _1279_ /*39160*/;
  assign _1281_ = ~q[26] /*39159*/;
  assign _1282_ = sum_6[11] & q[26] /*39158*/;
  assign _1283_ = m_6[11] & _1281_ /*39157*/;
  assign r_6[37] = _1283_ | _1282_ /*39156*/;
  assign _1284_ = ~q[26] /*39155*/;
  assign _1285_ = sum_6[12] & q[26] /*39154*/;
  assign _1286_ = m_6[12] & _1284_ /*39153*/;
  assign r_6[38] = _1286_ | _1285_ /*39152*/;
  assign _1287_ = ~q[26] /*39151*/;
  assign _1288_ = sum_6[13] & q[26] /*39150*/;
  assign _1289_ = m_6[13] & _1287_ /*39149*/;
  assign r_6[39] = _1289_ | _1288_ /*39148*/;
  assign _1290_ = ~q[26] /*39147*/;
  assign _1291_ = sum_6[14] & q[26] /*39146*/;
  assign _1292_ = m_6[14] & _1290_ /*39145*/;
  assign r_6[40] = _1292_ | _1291_ /*39144*/;
  assign _1293_ = ~q[26] /*39143*/;
  assign _1294_ = sum_6[15] & q[26] /*39142*/;
  assign _1295_ = m_6[15] & _1293_ /*39141*/;
  assign r_6[41] = _1295_ | _1294_ /*39140*/;
  assign _1296_ = ~q[26] /*39139*/;
  assign _1297_ = sum_6[16] & q[26] /*39138*/;
  assign _1298_ = m_6[16] & _1296_ /*39137*/;
  assign r_6[42] = _1298_ | _1297_ /*39136*/;
  assign _1299_ = ~q[26] /*39135*/;
  assign _1300_ = sum_6[17] & q[26] /*39134*/;
  assign _1301_ = m_6[17] & _1299_ /*39133*/;
  assign r_6[43] = _1301_ | _1300_ /*39132*/;
  assign _1302_ = ~q[26] /*39131*/;
  assign _1303_ = sum_6[18] & q[26] /*39130*/;
  assign _1304_ = m_6[18] & _1302_ /*39129*/;
  assign r_6[44] = _1304_ | _1303_ /*39128*/;
  assign _1305_ = ~q[26] /*39127*/;
  assign _1306_ = sum_6[19] & q[26] /*39126*/;
  assign _1307_ = m_6[19] & _1305_ /*39125*/;
  assign r_6[45] = _1307_ | _1306_ /*39124*/;
  assign _1308_ = ~q[26] /*39123*/;
  assign _1309_ = sum_6[20] & q[26] /*39122*/;
  assign _1310_ = m_6[20] & _1308_ /*39121*/;
  assign r_6[46] = _1310_ | _1309_ /*39120*/;
  assign _1311_ = ~q[26] /*39119*/;
  assign _1312_ = sum_6[21] & q[26] /*39118*/;
  assign _1313_ = m_6[21] & _1311_ /*39117*/;
  assign r_6[47] = _1313_ | _1312_ /*39116*/;
  assign _1314_ = ~q[26] /*39115*/;
  assign _1315_ = sum_6[22] & q[26] /*39114*/;
  assign _1316_ = m_6[22] & _1314_ /*39113*/;
  assign r_6[48] = _1316_ | _1315_ /*39112*/;
  assign _1317_ = ~q[26] /*39111*/;
  assign _1318_ = sum_6[23] & q[26] /*39110*/;
  assign _1319_ = m_6[23] & _1317_ /*39109*/;
  assign r_6[49] = _1319_ | _1318_ /*39108*/;
  assign _1320_ = ~q[26] /*39107*/;
  assign _1321_ = sum_6[24] & q[26] /*39106*/;
  assign _1322_ = m_6[24] & _1320_ /*39105*/;
  assign r_6[50] = _1322_ | _1321_ /*39104*/;
  assign _1323_ = ~q[26] /*39103*/;
  assign _1324_ = sum_6[25] & q[26] /*39102*/;
  assign _1325_ = m_6[25] & _1323_ /*39101*/;
  assign r_6[51] = _1325_ | _1324_ /*39100*/;
  assign _1326_ = ~q[26] /*39099*/;
  assign _1327_ = sum_6[26] & q[26] /*39098*/;
  assign _1328_ = m_6[26] & _1326_ /*39097*/;
  assign r_6[52] = _1328_ | _1327_ /*39096*/;
  assign _1329_ = ~q[26] /*39095*/;
  assign _1330_ = sum_6[27] & q[26] /*39094*/;
  assign _1331_ = m_6[27] & _1329_ /*39093*/;
  assign r_6[53] = _1331_ | _1330_ /*39092*/;
  assign _1332_ = ~q[26] /*39091*/;
  assign _1333_ = sum_6[28] & q[26] /*39090*/;
  assign _1334_ = m_6[28] & _1332_ /*39089*/;
  assign r_6[54] = _1334_ | _1333_ /*39088*/;
  assign _1335_ = ~q[26] /*39087*/;
  assign _1336_ = sum_6[29] & q[26] /*39086*/;
  assign _1337_ = m_6[29] & _1335_ /*39085*/;
  assign r_6[55] = _1337_ | _1336_ /*39084*/;
  assign _1338_ = ~q[26] /*39083*/;
  assign _1339_ = sum_6[30] & q[26] /*39082*/;
  assign _1340_ = m_6[30] & _1338_ /*39081*/;
  assign r_6[56] = _1340_ | _1339_ /*39080*/;
  assign _1341_ = ~q[26] /*39079*/;
  assign _1342_ = sum_6[31] & q[26] /*39078*/;
  assign _1343_ = m_6[31] & _1341_ /*39077*/;
  assign r_6[57] = _1343_ | _1342_ /*39076*/;
assign r_6[0]= r_5[0] /*39075*/;
assign r_6[1]= r_5[1] /*39074*/;
assign r_6[2]= r_5[2] /*39073*/;
assign r_6[3]= r_5[3] /*39072*/;
assign r_6[4]= r_5[4] /*39071*/;
assign r_6[5]= r_5[5] /*39070*/;
assign r_6[6]= r_5[6] /*39069*/;
assign r_6[7]= r_5[7] /*39068*/;
assign r_6[8]= r_5[8] /*39067*/;
assign r_6[9]= r_5[9] /*39066*/;
assign r_6[10]= r_5[10] /*39065*/;
assign r_6[11]= r_5[11] /*39064*/;
assign r_6[12]= r_5[12] /*39063*/;
assign r_6[13]= r_5[13] /*39062*/;
assign r_6[14]= r_5[14] /*39061*/;
assign r_6[15]= r_5[15] /*39060*/;
assign r_6[16]= r_5[16] /*39059*/;
assign r_6[17]= r_5[17] /*39058*/;
assign r_6[18]= r_5[18] /*39057*/;
assign r_6[19]= r_5[19] /*39056*/;
assign r_6[20]= r_5[20] /*39055*/;
assign r_6[21]= r_5[21] /*39054*/;
assign r_6[22]= r_5[22] /*39053*/;
assign r_6[23]= r_5[23] /*39052*/;
assign r_6[24]= r_5[24] /*39051*/;
assign r_6[25]= r_5[25] /*39050*/;
  assign inv_7[0] = ~div[0] /*38984*/;
  assign inv_7[1] = ~div[1] /*38983*/;
  assign inv_7[2] = ~div[2] /*38982*/;
  assign inv_7[3] = ~div[3] /*38981*/;
  assign inv_7[4] = ~div[4] /*38980*/;
  assign inv_7[5] = ~div[5] /*38979*/;
  assign inv_7[6] = ~div[6] /*38978*/;
  assign inv_7[7] = ~div[7] /*38977*/;
  assign inv_7[8] = ~div[8] /*38976*/;
  assign inv_7[9] = ~div[9] /*38975*/;
  assign inv_7[10] = ~div[10] /*38974*/;
  assign inv_7[11] = ~div[11] /*38973*/;
  assign inv_7[12] = ~div[12] /*38972*/;
  assign inv_7[13] = ~div[13] /*38971*/;
  assign inv_7[14] = ~div[14] /*38970*/;
  assign inv_7[15] = ~div[15] /*38969*/;
  assign inv_7[16] = ~div[16] /*38968*/;
  assign inv_7[17] = ~div[17] /*38967*/;
  assign inv_7[18] = ~div[18] /*38966*/;
  assign inv_7[19] = ~div[19] /*38965*/;
  assign inv_7[20] = ~div[20] /*38964*/;
  assign inv_7[21] = ~div[21] /*38963*/;
  assign inv_7[22] = ~div[22] /*38962*/;
  assign inv_7[23] = ~div[23] /*38961*/;
  assign inv_7[24] = ~div[24] /*38960*/;
  assign inv_7[25] = ~div[25] /*38959*/;
  assign inv_7[26] = ~div[26] /*38958*/;
  assign inv_7[27] = ~div[27] /*38957*/;
  assign inv_7[28] = ~div[28] /*38956*/;
  assign inv_7[29] = ~div[29] /*38955*/;
  assign inv_7[30] = ~div[30] /*38954*/;
assign inv_7[31] = oneWire /*38953*/;
  assign _1344_ = inv_7[0] ^ r_6[25] /*38951*/;
  assign sum_7[0] = _1344_ ^ oneWire /*38950*/;
  assign _1345_ = _1344_ & oneWire /*38949*/;
  assign _1346_ = inv_7[0] & r_6[25] /*38948*/;
  assign _1347_ = _1345_ | _1346_ /*38947*/;
  assign _1348_ = inv_7[1] ^ r_6[26] /*38946*/;
  assign sum_7[1] = _1348_ ^ _1347_ /*38945*/;
  assign _1349_ = _1348_ & _1347_ /*38944*/;
  assign _1350_ = inv_7[1] & r_6[26] /*38943*/;
  assign _1351_ = _1349_ | _1350_ /*38942*/;
  assign _1352_ = inv_7[2] ^ r_6[27] /*38940*/;
  assign sum_7[2] = _1352_ ^ _1351_ /*38939*/;
  assign _1353_ = _1352_ & _1351_ /*38938*/;
  assign _1354_ = inv_7[2] & r_6[27] /*38937*/;
  assign _1355_ = _1353_ | _1354_ /*38936*/;
  assign _1356_ = inv_7[3] ^ r_6[28] /*38934*/;
  assign sum_7[3] = _1356_ ^ _1355_ /*38933*/;
  assign _1357_ = _1356_ & _1355_ /*38932*/;
  assign _1358_ = inv_7[3] & r_6[28] /*38931*/;
  assign _1359_ = _1357_ | _1358_ /*38930*/;
  assign _1360_ = inv_7[4] ^ r_6[29] /*38928*/;
  assign sum_7[4] = _1360_ ^ _1359_ /*38927*/;
  assign _1361_ = _1360_ & _1359_ /*38926*/;
  assign _1362_ = inv_7[4] & r_6[29] /*38925*/;
  assign _1363_ = _1361_ | _1362_ /*38924*/;
  assign _1364_ = inv_7[5] ^ r_6[30] /*38922*/;
  assign sum_7[5] = _1364_ ^ _1363_ /*38921*/;
  assign _1365_ = _1364_ & _1363_ /*38920*/;
  assign _1366_ = inv_7[5] & r_6[30] /*38919*/;
  assign _1367_ = _1365_ | _1366_ /*38918*/;
  assign _1368_ = inv_7[6] ^ r_6[31] /*38916*/;
  assign sum_7[6] = _1368_ ^ _1367_ /*38915*/;
  assign _1369_ = _1368_ & _1367_ /*38914*/;
  assign _1370_ = inv_7[6] & r_6[31] /*38913*/;
  assign _1371_ = _1369_ | _1370_ /*38912*/;
  assign _1372_ = inv_7[7] ^ r_6[32] /*38910*/;
  assign sum_7[7] = _1372_ ^ _1371_ /*38909*/;
  assign _1373_ = _1372_ & _1371_ /*38908*/;
  assign _1374_ = inv_7[7] & r_6[32] /*38907*/;
  assign _1375_ = _1373_ | _1374_ /*38906*/;
  assign _1376_ = inv_7[8] ^ r_6[33] /*38904*/;
  assign sum_7[8] = _1376_ ^ _1375_ /*38903*/;
  assign _1377_ = _1376_ & _1375_ /*38902*/;
  assign _1378_ = inv_7[8] & r_6[33] /*38901*/;
  assign _1379_ = _1377_ | _1378_ /*38900*/;
  assign _1380_ = inv_7[9] ^ r_6[34] /*38898*/;
  assign sum_7[9] = _1380_ ^ _1379_ /*38897*/;
  assign _1381_ = _1380_ & _1379_ /*38896*/;
  assign _1382_ = inv_7[9] & r_6[34] /*38895*/;
  assign _1383_ = _1381_ | _1382_ /*38894*/;
  assign _1384_ = inv_7[10] ^ r_6[35] /*38892*/;
  assign sum_7[10] = _1384_ ^ _1383_ /*38891*/;
  assign _1385_ = _1384_ & _1383_ /*38890*/;
  assign _1386_ = inv_7[10] & r_6[35] /*38889*/;
  assign _1387_ = _1385_ | _1386_ /*38888*/;
  assign _1388_ = inv_7[11] ^ r_6[36] /*38886*/;
  assign sum_7[11] = _1388_ ^ _1387_ /*38885*/;
  assign _1389_ = _1388_ & _1387_ /*38884*/;
  assign _1390_ = inv_7[11] & r_6[36] /*38883*/;
  assign _1391_ = _1389_ | _1390_ /*38882*/;
  assign _1392_ = inv_7[12] ^ r_6[37] /*38880*/;
  assign sum_7[12] = _1392_ ^ _1391_ /*38879*/;
  assign _1393_ = _1392_ & _1391_ /*38878*/;
  assign _1394_ = inv_7[12] & r_6[37] /*38877*/;
  assign _1395_ = _1393_ | _1394_ /*38876*/;
  assign _1396_ = inv_7[13] ^ r_6[38] /*38874*/;
  assign sum_7[13] = _1396_ ^ _1395_ /*38873*/;
  assign _1397_ = _1396_ & _1395_ /*38872*/;
  assign _1398_ = inv_7[13] & r_6[38] /*38871*/;
  assign _1399_ = _1397_ | _1398_ /*38870*/;
  assign _1400_ = inv_7[14] ^ r_6[39] /*38868*/;
  assign sum_7[14] = _1400_ ^ _1399_ /*38867*/;
  assign _1401_ = _1400_ & _1399_ /*38866*/;
  assign _1402_ = inv_7[14] & r_6[39] /*38865*/;
  assign _1403_ = _1401_ | _1402_ /*38864*/;
  assign _1404_ = inv_7[15] ^ r_6[40] /*38862*/;
  assign sum_7[15] = _1404_ ^ _1403_ /*38861*/;
  assign _1405_ = _1404_ & _1403_ /*38860*/;
  assign _1406_ = inv_7[15] & r_6[40] /*38859*/;
  assign _1407_ = _1405_ | _1406_ /*38858*/;
  assign _1408_ = inv_7[16] ^ r_6[41] /*38856*/;
  assign sum_7[16] = _1408_ ^ _1407_ /*38855*/;
  assign _1409_ = _1408_ & _1407_ /*38854*/;
  assign _1410_ = inv_7[16] & r_6[41] /*38853*/;
  assign _1411_ = _1409_ | _1410_ /*38852*/;
  assign _1412_ = inv_7[17] ^ r_6[42] /*38850*/;
  assign sum_7[17] = _1412_ ^ _1411_ /*38849*/;
  assign _1413_ = _1412_ & _1411_ /*38848*/;
  assign _1414_ = inv_7[17] & r_6[42] /*38847*/;
  assign _1415_ = _1413_ | _1414_ /*38846*/;
  assign _1416_ = inv_7[18] ^ r_6[43] /*38844*/;
  assign sum_7[18] = _1416_ ^ _1415_ /*38843*/;
  assign _1417_ = _1416_ & _1415_ /*38842*/;
  assign _1418_ = inv_7[18] & r_6[43] /*38841*/;
  assign _1419_ = _1417_ | _1418_ /*38840*/;
  assign _1420_ = inv_7[19] ^ r_6[44] /*38838*/;
  assign sum_7[19] = _1420_ ^ _1419_ /*38837*/;
  assign _1421_ = _1420_ & _1419_ /*38836*/;
  assign _1422_ = inv_7[19] & r_6[44] /*38835*/;
  assign _1423_ = _1421_ | _1422_ /*38834*/;
  assign _1424_ = inv_7[20] ^ r_6[45] /*38832*/;
  assign sum_7[20] = _1424_ ^ _1423_ /*38831*/;
  assign _1425_ = _1424_ & _1423_ /*38830*/;
  assign _1426_ = inv_7[20] & r_6[45] /*38829*/;
  assign _1427_ = _1425_ | _1426_ /*38828*/;
  assign _1428_ = inv_7[21] ^ r_6[46] /*38826*/;
  assign sum_7[21] = _1428_ ^ _1427_ /*38825*/;
  assign _1429_ = _1428_ & _1427_ /*38824*/;
  assign _1430_ = inv_7[21] & r_6[46] /*38823*/;
  assign _1431_ = _1429_ | _1430_ /*38822*/;
  assign _1432_ = inv_7[22] ^ r_6[47] /*38820*/;
  assign sum_7[22] = _1432_ ^ _1431_ /*38819*/;
  assign _1433_ = _1432_ & _1431_ /*38818*/;
  assign _1434_ = inv_7[22] & r_6[47] /*38817*/;
  assign _1435_ = _1433_ | _1434_ /*38816*/;
  assign _1436_ = inv_7[23] ^ r_6[48] /*38814*/;
  assign sum_7[23] = _1436_ ^ _1435_ /*38813*/;
  assign _1437_ = _1436_ & _1435_ /*38812*/;
  assign _1438_ = inv_7[23] & r_6[48] /*38811*/;
  assign _1439_ = _1437_ | _1438_ /*38810*/;
  assign _1440_ = inv_7[24] ^ r_6[49] /*38808*/;
  assign sum_7[24] = _1440_ ^ _1439_ /*38807*/;
  assign _1441_ = _1440_ & _1439_ /*38806*/;
  assign _1442_ = inv_7[24] & r_6[49] /*38805*/;
  assign _1443_ = _1441_ | _1442_ /*38804*/;
  assign _1444_ = inv_7[25] ^ r_6[50] /*38802*/;
  assign sum_7[25] = _1444_ ^ _1443_ /*38801*/;
  assign _1445_ = _1444_ & _1443_ /*38800*/;
  assign _1446_ = inv_7[25] & r_6[50] /*38799*/;
  assign _1447_ = _1445_ | _1446_ /*38798*/;
  assign _1448_ = inv_7[26] ^ r_6[51] /*38796*/;
  assign sum_7[26] = _1448_ ^ _1447_ /*38795*/;
  assign _1449_ = _1448_ & _1447_ /*38794*/;
  assign _1450_ = inv_7[26] & r_6[51] /*38793*/;
  assign _1451_ = _1449_ | _1450_ /*38792*/;
  assign _1452_ = inv_7[27] ^ r_6[52] /*38790*/;
  assign sum_7[27] = _1452_ ^ _1451_ /*38789*/;
  assign _1453_ = _1452_ & _1451_ /*38788*/;
  assign _1454_ = inv_7[27] & r_6[52] /*38787*/;
  assign _1455_ = _1453_ | _1454_ /*38786*/;
  assign _1456_ = inv_7[28] ^ r_6[53] /*38784*/;
  assign sum_7[28] = _1456_ ^ _1455_ /*38783*/;
  assign _1457_ = _1456_ & _1455_ /*38782*/;
  assign _1458_ = inv_7[28] & r_6[53] /*38781*/;
  assign _1459_ = _1457_ | _1458_ /*38780*/;
  assign _1460_ = inv_7[29] ^ r_6[54] /*38778*/;
  assign sum_7[29] = _1460_ ^ _1459_ /*38777*/;
  assign _1461_ = _1460_ & _1459_ /*38776*/;
  assign _1462_ = inv_7[29] & r_6[54] /*38775*/;
  assign _1463_ = _1461_ | _1462_ /*38774*/;
  assign _1464_ = inv_7[30] ^ r_6[55] /*38772*/;
  assign sum_7[30] = _1464_ ^ _1463_ /*38771*/;
  assign _1465_ = _1464_ & _1463_ /*38770*/;
  assign _1466_ = inv_7[30] & r_6[55] /*38769*/;
  assign _1467_ = _1465_ | _1466_ /*38768*/;
  assign _1468_ = inv_7[31] ^ r_6[56] /*38766*/;
  assign sum_7[31] = _1468_ ^ _1467_ /*38765*/;
  assign _1469_ = _1468_ & _1467_ /*38764*/;
  assign _1470_ = inv_7[31] & r_6[56] /*38763*/;
  assign _1471_ = _1469_ | _1470_ /*38762*/;
  assign q[25] = ~sum_7[31] /*38789*/;
  assign m_7[0] = r_6[25] /*38788*/;
  assign m_7[1] = r_6[26] /*38787*/;
  assign m_7[2] = r_6[27] /*38786*/;
  assign m_7[3] = r_6[28] /*38785*/;
  assign m_7[4] = r_6[29] /*38784*/;
  assign m_7[5] = r_6[30] /*38783*/;
  assign m_7[6] = r_6[31] /*38782*/;
  assign m_7[7] = r_6[32] /*38781*/;
  assign m_7[8] = r_6[33] /*38780*/;
  assign m_7[9] = r_6[34] /*38779*/;
  assign m_7[10] = r_6[35] /*38778*/;
  assign m_7[11] = r_6[36] /*38777*/;
  assign m_7[12] = r_6[37] /*38776*/;
  assign m_7[13] = r_6[38] /*38775*/;
  assign m_7[14] = r_6[39] /*38774*/;
  assign m_7[15] = r_6[40] /*38773*/;
  assign m_7[16] = r_6[41] /*38772*/;
  assign m_7[17] = r_6[42] /*38771*/;
  assign m_7[18] = r_6[43] /*38770*/;
  assign m_7[19] = r_6[44] /*38769*/;
  assign m_7[20] = r_6[45] /*38768*/;
  assign m_7[21] = r_6[46] /*38767*/;
  assign m_7[22] = r_6[47] /*38766*/;
  assign m_7[23] = r_6[48] /*38765*/;
  assign m_7[24] = r_6[49] /*38764*/;
  assign m_7[25] = r_6[50] /*38763*/;
  assign m_7[26] = r_6[51] /*38762*/;
  assign m_7[27] = r_6[52] /*38761*/;
  assign m_7[28] = r_6[53] /*38760*/;
  assign m_7[29] = r_6[54] /*38759*/;
  assign m_7[30] = r_6[55] /*38758*/;
  assign m_7[31] = r_6[56] /*38757*/;
  assign _1472_ = ~q[25] /*38755*/;
  assign _1473_ = sum_7[0] & q[25] /*38754*/;
  assign _1474_ = m_7[0] & _1472_ /*38753*/;
  assign r_7[25] = _1474_ | _1473_ /*38752*/;
  assign _1475_ = ~q[25] /*38751*/;
  assign _1476_ = sum_7[1] & q[25] /*38750*/;
  assign _1477_ = m_7[1] & _1475_ /*38749*/;
  assign r_7[26] = _1477_ | _1476_ /*38748*/;
  assign _1478_ = ~q[25] /*38747*/;
  assign _1479_ = sum_7[2] & q[25] /*38746*/;
  assign _1480_ = m_7[2] & _1478_ /*38745*/;
  assign r_7[27] = _1480_ | _1479_ /*38744*/;
  assign _1481_ = ~q[25] /*38743*/;
  assign _1482_ = sum_7[3] & q[25] /*38742*/;
  assign _1483_ = m_7[3] & _1481_ /*38741*/;
  assign r_7[28] = _1483_ | _1482_ /*38740*/;
  assign _1484_ = ~q[25] /*38739*/;
  assign _1485_ = sum_7[4] & q[25] /*38738*/;
  assign _1486_ = m_7[4] & _1484_ /*38737*/;
  assign r_7[29] = _1486_ | _1485_ /*38736*/;
  assign _1487_ = ~q[25] /*38735*/;
  assign _1488_ = sum_7[5] & q[25] /*38734*/;
  assign _1489_ = m_7[5] & _1487_ /*38733*/;
  assign r_7[30] = _1489_ | _1488_ /*38732*/;
  assign _1490_ = ~q[25] /*38731*/;
  assign _1491_ = sum_7[6] & q[25] /*38730*/;
  assign _1492_ = m_7[6] & _1490_ /*38729*/;
  assign r_7[31] = _1492_ | _1491_ /*38728*/;
  assign _1493_ = ~q[25] /*38727*/;
  assign _1494_ = sum_7[7] & q[25] /*38726*/;
  assign _1495_ = m_7[7] & _1493_ /*38725*/;
  assign r_7[32] = _1495_ | _1494_ /*38724*/;
  assign _1496_ = ~q[25] /*38723*/;
  assign _1497_ = sum_7[8] & q[25] /*38722*/;
  assign _1498_ = m_7[8] & _1496_ /*38721*/;
  assign r_7[33] = _1498_ | _1497_ /*38720*/;
  assign _1499_ = ~q[25] /*38719*/;
  assign _1500_ = sum_7[9] & q[25] /*38718*/;
  assign _1501_ = m_7[9] & _1499_ /*38717*/;
  assign r_7[34] = _1501_ | _1500_ /*38716*/;
  assign _1502_ = ~q[25] /*38715*/;
  assign _1503_ = sum_7[10] & q[25] /*38714*/;
  assign _1504_ = m_7[10] & _1502_ /*38713*/;
  assign r_7[35] = _1504_ | _1503_ /*38712*/;
  assign _1505_ = ~q[25] /*38711*/;
  assign _1506_ = sum_7[11] & q[25] /*38710*/;
  assign _1507_ = m_7[11] & _1505_ /*38709*/;
  assign r_7[36] = _1507_ | _1506_ /*38708*/;
  assign _1508_ = ~q[25] /*38707*/;
  assign _1509_ = sum_7[12] & q[25] /*38706*/;
  assign _1510_ = m_7[12] & _1508_ /*38705*/;
  assign r_7[37] = _1510_ | _1509_ /*38704*/;
  assign _1511_ = ~q[25] /*38703*/;
  assign _1512_ = sum_7[13] & q[25] /*38702*/;
  assign _1513_ = m_7[13] & _1511_ /*38701*/;
  assign r_7[38] = _1513_ | _1512_ /*38700*/;
  assign _1514_ = ~q[25] /*38699*/;
  assign _1515_ = sum_7[14] & q[25] /*38698*/;
  assign _1516_ = m_7[14] & _1514_ /*38697*/;
  assign r_7[39] = _1516_ | _1515_ /*38696*/;
  assign _1517_ = ~q[25] /*38695*/;
  assign _1518_ = sum_7[15] & q[25] /*38694*/;
  assign _1519_ = m_7[15] & _1517_ /*38693*/;
  assign r_7[40] = _1519_ | _1518_ /*38692*/;
  assign _1520_ = ~q[25] /*38691*/;
  assign _1521_ = sum_7[16] & q[25] /*38690*/;
  assign _1522_ = m_7[16] & _1520_ /*38689*/;
  assign r_7[41] = _1522_ | _1521_ /*38688*/;
  assign _1523_ = ~q[25] /*38687*/;
  assign _1524_ = sum_7[17] & q[25] /*38686*/;
  assign _1525_ = m_7[17] & _1523_ /*38685*/;
  assign r_7[42] = _1525_ | _1524_ /*38684*/;
  assign _1526_ = ~q[25] /*38683*/;
  assign _1527_ = sum_7[18] & q[25] /*38682*/;
  assign _1528_ = m_7[18] & _1526_ /*38681*/;
  assign r_7[43] = _1528_ | _1527_ /*38680*/;
  assign _1529_ = ~q[25] /*38679*/;
  assign _1530_ = sum_7[19] & q[25] /*38678*/;
  assign _1531_ = m_7[19] & _1529_ /*38677*/;
  assign r_7[44] = _1531_ | _1530_ /*38676*/;
  assign _1532_ = ~q[25] /*38675*/;
  assign _1533_ = sum_7[20] & q[25] /*38674*/;
  assign _1534_ = m_7[20] & _1532_ /*38673*/;
  assign r_7[45] = _1534_ | _1533_ /*38672*/;
  assign _1535_ = ~q[25] /*38671*/;
  assign _1536_ = sum_7[21] & q[25] /*38670*/;
  assign _1537_ = m_7[21] & _1535_ /*38669*/;
  assign r_7[46] = _1537_ | _1536_ /*38668*/;
  assign _1538_ = ~q[25] /*38667*/;
  assign _1539_ = sum_7[22] & q[25] /*38666*/;
  assign _1540_ = m_7[22] & _1538_ /*38665*/;
  assign r_7[47] = _1540_ | _1539_ /*38664*/;
  assign _1541_ = ~q[25] /*38663*/;
  assign _1542_ = sum_7[23] & q[25] /*38662*/;
  assign _1543_ = m_7[23] & _1541_ /*38661*/;
  assign r_7[48] = _1543_ | _1542_ /*38660*/;
  assign _1544_ = ~q[25] /*38659*/;
  assign _1545_ = sum_7[24] & q[25] /*38658*/;
  assign _1546_ = m_7[24] & _1544_ /*38657*/;
  assign r_7[49] = _1546_ | _1545_ /*38656*/;
  assign _1547_ = ~q[25] /*38655*/;
  assign _1548_ = sum_7[25] & q[25] /*38654*/;
  assign _1549_ = m_7[25] & _1547_ /*38653*/;
  assign r_7[50] = _1549_ | _1548_ /*38652*/;
  assign _1550_ = ~q[25] /*38651*/;
  assign _1551_ = sum_7[26] & q[25] /*38650*/;
  assign _1552_ = m_7[26] & _1550_ /*38649*/;
  assign r_7[51] = _1552_ | _1551_ /*38648*/;
  assign _1553_ = ~q[25] /*38647*/;
  assign _1554_ = sum_7[27] & q[25] /*38646*/;
  assign _1555_ = m_7[27] & _1553_ /*38645*/;
  assign r_7[52] = _1555_ | _1554_ /*38644*/;
  assign _1556_ = ~q[25] /*38643*/;
  assign _1557_ = sum_7[28] & q[25] /*38642*/;
  assign _1558_ = m_7[28] & _1556_ /*38641*/;
  assign r_7[53] = _1558_ | _1557_ /*38640*/;
  assign _1559_ = ~q[25] /*38639*/;
  assign _1560_ = sum_7[29] & q[25] /*38638*/;
  assign _1561_ = m_7[29] & _1559_ /*38637*/;
  assign r_7[54] = _1561_ | _1560_ /*38636*/;
  assign _1562_ = ~q[25] /*38635*/;
  assign _1563_ = sum_7[30] & q[25] /*38634*/;
  assign _1564_ = m_7[30] & _1562_ /*38633*/;
  assign r_7[55] = _1564_ | _1563_ /*38632*/;
  assign _1565_ = ~q[25] /*38631*/;
  assign _1566_ = sum_7[31] & q[25] /*38630*/;
  assign _1567_ = m_7[31] & _1565_ /*38629*/;
  assign r_7[56] = _1567_ | _1566_ /*38628*/;
assign r_7[0]= r_6[0] /*38627*/;
assign r_7[1]= r_6[1] /*38626*/;
assign r_7[2]= r_6[2] /*38625*/;
assign r_7[3]= r_6[3] /*38624*/;
assign r_7[4]= r_6[4] /*38623*/;
assign r_7[5]= r_6[5] /*38622*/;
assign r_7[6]= r_6[6] /*38621*/;
assign r_7[7]= r_6[7] /*38620*/;
assign r_7[8]= r_6[8] /*38619*/;
assign r_7[9]= r_6[9] /*38618*/;
assign r_7[10]= r_6[10] /*38617*/;
assign r_7[11]= r_6[11] /*38616*/;
assign r_7[12]= r_6[12] /*38615*/;
assign r_7[13]= r_6[13] /*38614*/;
assign r_7[14]= r_6[14] /*38613*/;
assign r_7[15]= r_6[15] /*38612*/;
assign r_7[16]= r_6[16] /*38611*/;
assign r_7[17]= r_6[17] /*38610*/;
assign r_7[18]= r_6[18] /*38609*/;
assign r_7[19]= r_6[19] /*38608*/;
assign r_7[20]= r_6[20] /*38607*/;
assign r_7[21]= r_6[21] /*38606*/;
assign r_7[22]= r_6[22] /*38605*/;
assign r_7[23]= r_6[23] /*38604*/;
assign r_7[24]= r_6[24] /*38603*/;
  assign inv_8[0] = ~div[0] /*38536*/;
  assign inv_8[1] = ~div[1] /*38535*/;
  assign inv_8[2] = ~div[2] /*38534*/;
  assign inv_8[3] = ~div[3] /*38533*/;
  assign inv_8[4] = ~div[4] /*38532*/;
  assign inv_8[5] = ~div[5] /*38531*/;
  assign inv_8[6] = ~div[6] /*38530*/;
  assign inv_8[7] = ~div[7] /*38529*/;
  assign inv_8[8] = ~div[8] /*38528*/;
  assign inv_8[9] = ~div[9] /*38527*/;
  assign inv_8[10] = ~div[10] /*38526*/;
  assign inv_8[11] = ~div[11] /*38525*/;
  assign inv_8[12] = ~div[12] /*38524*/;
  assign inv_8[13] = ~div[13] /*38523*/;
  assign inv_8[14] = ~div[14] /*38522*/;
  assign inv_8[15] = ~div[15] /*38521*/;
  assign inv_8[16] = ~div[16] /*38520*/;
  assign inv_8[17] = ~div[17] /*38519*/;
  assign inv_8[18] = ~div[18] /*38518*/;
  assign inv_8[19] = ~div[19] /*38517*/;
  assign inv_8[20] = ~div[20] /*38516*/;
  assign inv_8[21] = ~div[21] /*38515*/;
  assign inv_8[22] = ~div[22] /*38514*/;
  assign inv_8[23] = ~div[23] /*38513*/;
  assign inv_8[24] = ~div[24] /*38512*/;
  assign inv_8[25] = ~div[25] /*38511*/;
  assign inv_8[26] = ~div[26] /*38510*/;
  assign inv_8[27] = ~div[27] /*38509*/;
  assign inv_8[28] = ~div[28] /*38508*/;
  assign inv_8[29] = ~div[29] /*38507*/;
  assign inv_8[30] = ~div[30] /*38506*/;
assign inv_8[31] = oneWire /*38505*/;
  assign _1568_ = inv_8[0] ^ r_7[24] /*38503*/;
  assign sum_8[0] = _1568_ ^ oneWire /*38502*/;
  assign _1569_ = _1568_ & oneWire /*38501*/;
  assign _1570_ = inv_8[0] & r_7[24] /*38500*/;
  assign _1571_ = _1569_ | _1570_ /*38499*/;
  assign _1572_ = inv_8[1] ^ r_7[25] /*38498*/;
  assign sum_8[1] = _1572_ ^ _1571_ /*38497*/;
  assign _1573_ = _1572_ & _1571_ /*38496*/;
  assign _1574_ = inv_8[1] & r_7[25] /*38495*/;
  assign _1575_ = _1573_ | _1574_ /*38494*/;
  assign _1576_ = inv_8[2] ^ r_7[26] /*38492*/;
  assign sum_8[2] = _1576_ ^ _1575_ /*38491*/;
  assign _1577_ = _1576_ & _1575_ /*38490*/;
  assign _1578_ = inv_8[2] & r_7[26] /*38489*/;
  assign _1579_ = _1577_ | _1578_ /*38488*/;
  assign _1580_ = inv_8[3] ^ r_7[27] /*38486*/;
  assign sum_8[3] = _1580_ ^ _1579_ /*38485*/;
  assign _1581_ = _1580_ & _1579_ /*38484*/;
  assign _1582_ = inv_8[3] & r_7[27] /*38483*/;
  assign _1583_ = _1581_ | _1582_ /*38482*/;
  assign _1584_ = inv_8[4] ^ r_7[28] /*38480*/;
  assign sum_8[4] = _1584_ ^ _1583_ /*38479*/;
  assign _1585_ = _1584_ & _1583_ /*38478*/;
  assign _1586_ = inv_8[4] & r_7[28] /*38477*/;
  assign _1587_ = _1585_ | _1586_ /*38476*/;
  assign _1588_ = inv_8[5] ^ r_7[29] /*38474*/;
  assign sum_8[5] = _1588_ ^ _1587_ /*38473*/;
  assign _1589_ = _1588_ & _1587_ /*38472*/;
  assign _1590_ = inv_8[5] & r_7[29] /*38471*/;
  assign _1591_ = _1589_ | _1590_ /*38470*/;
  assign _1592_ = inv_8[6] ^ r_7[30] /*38468*/;
  assign sum_8[6] = _1592_ ^ _1591_ /*38467*/;
  assign _1593_ = _1592_ & _1591_ /*38466*/;
  assign _1594_ = inv_8[6] & r_7[30] /*38465*/;
  assign _1595_ = _1593_ | _1594_ /*38464*/;
  assign _1596_ = inv_8[7] ^ r_7[31] /*38462*/;
  assign sum_8[7] = _1596_ ^ _1595_ /*38461*/;
  assign _1597_ = _1596_ & _1595_ /*38460*/;
  assign _1598_ = inv_8[7] & r_7[31] /*38459*/;
  assign _1599_ = _1597_ | _1598_ /*38458*/;
  assign _1600_ = inv_8[8] ^ r_7[32] /*38456*/;
  assign sum_8[8] = _1600_ ^ _1599_ /*38455*/;
  assign _1601_ = _1600_ & _1599_ /*38454*/;
  assign _1602_ = inv_8[8] & r_7[32] /*38453*/;
  assign _1603_ = _1601_ | _1602_ /*38452*/;
  assign _1604_ = inv_8[9] ^ r_7[33] /*38450*/;
  assign sum_8[9] = _1604_ ^ _1603_ /*38449*/;
  assign _1605_ = _1604_ & _1603_ /*38448*/;
  assign _1606_ = inv_8[9] & r_7[33] /*38447*/;
  assign _1607_ = _1605_ | _1606_ /*38446*/;
  assign _1608_ = inv_8[10] ^ r_7[34] /*38444*/;
  assign sum_8[10] = _1608_ ^ _1607_ /*38443*/;
  assign _1609_ = _1608_ & _1607_ /*38442*/;
  assign _1610_ = inv_8[10] & r_7[34] /*38441*/;
  assign _1611_ = _1609_ | _1610_ /*38440*/;
  assign _1612_ = inv_8[11] ^ r_7[35] /*38438*/;
  assign sum_8[11] = _1612_ ^ _1611_ /*38437*/;
  assign _1613_ = _1612_ & _1611_ /*38436*/;
  assign _1614_ = inv_8[11] & r_7[35] /*38435*/;
  assign _1615_ = _1613_ | _1614_ /*38434*/;
  assign _1616_ = inv_8[12] ^ r_7[36] /*38432*/;
  assign sum_8[12] = _1616_ ^ _1615_ /*38431*/;
  assign _1617_ = _1616_ & _1615_ /*38430*/;
  assign _1618_ = inv_8[12] & r_7[36] /*38429*/;
  assign _1619_ = _1617_ | _1618_ /*38428*/;
  assign _1620_ = inv_8[13] ^ r_7[37] /*38426*/;
  assign sum_8[13] = _1620_ ^ _1619_ /*38425*/;
  assign _1621_ = _1620_ & _1619_ /*38424*/;
  assign _1622_ = inv_8[13] & r_7[37] /*38423*/;
  assign _1623_ = _1621_ | _1622_ /*38422*/;
  assign _1624_ = inv_8[14] ^ r_7[38] /*38420*/;
  assign sum_8[14] = _1624_ ^ _1623_ /*38419*/;
  assign _1625_ = _1624_ & _1623_ /*38418*/;
  assign _1626_ = inv_8[14] & r_7[38] /*38417*/;
  assign _1627_ = _1625_ | _1626_ /*38416*/;
  assign _1628_ = inv_8[15] ^ r_7[39] /*38414*/;
  assign sum_8[15] = _1628_ ^ _1627_ /*38413*/;
  assign _1629_ = _1628_ & _1627_ /*38412*/;
  assign _1630_ = inv_8[15] & r_7[39] /*38411*/;
  assign _1631_ = _1629_ | _1630_ /*38410*/;
  assign _1632_ = inv_8[16] ^ r_7[40] /*38408*/;
  assign sum_8[16] = _1632_ ^ _1631_ /*38407*/;
  assign _1633_ = _1632_ & _1631_ /*38406*/;
  assign _1634_ = inv_8[16] & r_7[40] /*38405*/;
  assign _1635_ = _1633_ | _1634_ /*38404*/;
  assign _1636_ = inv_8[17] ^ r_7[41] /*38402*/;
  assign sum_8[17] = _1636_ ^ _1635_ /*38401*/;
  assign _1637_ = _1636_ & _1635_ /*38400*/;
  assign _1638_ = inv_8[17] & r_7[41] /*38399*/;
  assign _1639_ = _1637_ | _1638_ /*38398*/;
  assign _1640_ = inv_8[18] ^ r_7[42] /*38396*/;
  assign sum_8[18] = _1640_ ^ _1639_ /*38395*/;
  assign _1641_ = _1640_ & _1639_ /*38394*/;
  assign _1642_ = inv_8[18] & r_7[42] /*38393*/;
  assign _1643_ = _1641_ | _1642_ /*38392*/;
  assign _1644_ = inv_8[19] ^ r_7[43] /*38390*/;
  assign sum_8[19] = _1644_ ^ _1643_ /*38389*/;
  assign _1645_ = _1644_ & _1643_ /*38388*/;
  assign _1646_ = inv_8[19] & r_7[43] /*38387*/;
  assign _1647_ = _1645_ | _1646_ /*38386*/;
  assign _1648_ = inv_8[20] ^ r_7[44] /*38384*/;
  assign sum_8[20] = _1648_ ^ _1647_ /*38383*/;
  assign _1649_ = _1648_ & _1647_ /*38382*/;
  assign _1650_ = inv_8[20] & r_7[44] /*38381*/;
  assign _1651_ = _1649_ | _1650_ /*38380*/;
  assign _1652_ = inv_8[21] ^ r_7[45] /*38378*/;
  assign sum_8[21] = _1652_ ^ _1651_ /*38377*/;
  assign _1653_ = _1652_ & _1651_ /*38376*/;
  assign _1654_ = inv_8[21] & r_7[45] /*38375*/;
  assign _1655_ = _1653_ | _1654_ /*38374*/;
  assign _1656_ = inv_8[22] ^ r_7[46] /*38372*/;
  assign sum_8[22] = _1656_ ^ _1655_ /*38371*/;
  assign _1657_ = _1656_ & _1655_ /*38370*/;
  assign _1658_ = inv_8[22] & r_7[46] /*38369*/;
  assign _1659_ = _1657_ | _1658_ /*38368*/;
  assign _1660_ = inv_8[23] ^ r_7[47] /*38366*/;
  assign sum_8[23] = _1660_ ^ _1659_ /*38365*/;
  assign _1661_ = _1660_ & _1659_ /*38364*/;
  assign _1662_ = inv_8[23] & r_7[47] /*38363*/;
  assign _1663_ = _1661_ | _1662_ /*38362*/;
  assign _1664_ = inv_8[24] ^ r_7[48] /*38360*/;
  assign sum_8[24] = _1664_ ^ _1663_ /*38359*/;
  assign _1665_ = _1664_ & _1663_ /*38358*/;
  assign _1666_ = inv_8[24] & r_7[48] /*38357*/;
  assign _1667_ = _1665_ | _1666_ /*38356*/;
  assign _1668_ = inv_8[25] ^ r_7[49] /*38354*/;
  assign sum_8[25] = _1668_ ^ _1667_ /*38353*/;
  assign _1669_ = _1668_ & _1667_ /*38352*/;
  assign _1670_ = inv_8[25] & r_7[49] /*38351*/;
  assign _1671_ = _1669_ | _1670_ /*38350*/;
  assign _1672_ = inv_8[26] ^ r_7[50] /*38348*/;
  assign sum_8[26] = _1672_ ^ _1671_ /*38347*/;
  assign _1673_ = _1672_ & _1671_ /*38346*/;
  assign _1674_ = inv_8[26] & r_7[50] /*38345*/;
  assign _1675_ = _1673_ | _1674_ /*38344*/;
  assign _1676_ = inv_8[27] ^ r_7[51] /*38342*/;
  assign sum_8[27] = _1676_ ^ _1675_ /*38341*/;
  assign _1677_ = _1676_ & _1675_ /*38340*/;
  assign _1678_ = inv_8[27] & r_7[51] /*38339*/;
  assign _1679_ = _1677_ | _1678_ /*38338*/;
  assign _1680_ = inv_8[28] ^ r_7[52] /*38336*/;
  assign sum_8[28] = _1680_ ^ _1679_ /*38335*/;
  assign _1681_ = _1680_ & _1679_ /*38334*/;
  assign _1682_ = inv_8[28] & r_7[52] /*38333*/;
  assign _1683_ = _1681_ | _1682_ /*38332*/;
  assign _1684_ = inv_8[29] ^ r_7[53] /*38330*/;
  assign sum_8[29] = _1684_ ^ _1683_ /*38329*/;
  assign _1685_ = _1684_ & _1683_ /*38328*/;
  assign _1686_ = inv_8[29] & r_7[53] /*38327*/;
  assign _1687_ = _1685_ | _1686_ /*38326*/;
  assign _1688_ = inv_8[30] ^ r_7[54] /*38324*/;
  assign sum_8[30] = _1688_ ^ _1687_ /*38323*/;
  assign _1689_ = _1688_ & _1687_ /*38322*/;
  assign _1690_ = inv_8[30] & r_7[54] /*38321*/;
  assign _1691_ = _1689_ | _1690_ /*38320*/;
  assign _1692_ = inv_8[31] ^ r_7[55] /*38318*/;
  assign sum_8[31] = _1692_ ^ _1691_ /*38317*/;
  assign _1693_ = _1692_ & _1691_ /*38316*/;
  assign _1694_ = inv_8[31] & r_7[55] /*38315*/;
  assign _1695_ = _1693_ | _1694_ /*38314*/;
  assign q[24] = ~sum_8[31] /*38341*/;
  assign m_8[0] = r_7[24] /*38340*/;
  assign m_8[1] = r_7[25] /*38339*/;
  assign m_8[2] = r_7[26] /*38338*/;
  assign m_8[3] = r_7[27] /*38337*/;
  assign m_8[4] = r_7[28] /*38336*/;
  assign m_8[5] = r_7[29] /*38335*/;
  assign m_8[6] = r_7[30] /*38334*/;
  assign m_8[7] = r_7[31] /*38333*/;
  assign m_8[8] = r_7[32] /*38332*/;
  assign m_8[9] = r_7[33] /*38331*/;
  assign m_8[10] = r_7[34] /*38330*/;
  assign m_8[11] = r_7[35] /*38329*/;
  assign m_8[12] = r_7[36] /*38328*/;
  assign m_8[13] = r_7[37] /*38327*/;
  assign m_8[14] = r_7[38] /*38326*/;
  assign m_8[15] = r_7[39] /*38325*/;
  assign m_8[16] = r_7[40] /*38324*/;
  assign m_8[17] = r_7[41] /*38323*/;
  assign m_8[18] = r_7[42] /*38322*/;
  assign m_8[19] = r_7[43] /*38321*/;
  assign m_8[20] = r_7[44] /*38320*/;
  assign m_8[21] = r_7[45] /*38319*/;
  assign m_8[22] = r_7[46] /*38318*/;
  assign m_8[23] = r_7[47] /*38317*/;
  assign m_8[24] = r_7[48] /*38316*/;
  assign m_8[25] = r_7[49] /*38315*/;
  assign m_8[26] = r_7[50] /*38314*/;
  assign m_8[27] = r_7[51] /*38313*/;
  assign m_8[28] = r_7[52] /*38312*/;
  assign m_8[29] = r_7[53] /*38311*/;
  assign m_8[30] = r_7[54] /*38310*/;
  assign m_8[31] = r_7[55] /*38309*/;
  assign _1696_ = ~q[24] /*38307*/;
  assign _1697_ = sum_8[0] & q[24] /*38306*/;
  assign _1698_ = m_8[0] & _1696_ /*38305*/;
  assign r_8[24] = _1698_ | _1697_ /*38304*/;
  assign _1699_ = ~q[24] /*38303*/;
  assign _1700_ = sum_8[1] & q[24] /*38302*/;
  assign _1701_ = m_8[1] & _1699_ /*38301*/;
  assign r_8[25] = _1701_ | _1700_ /*38300*/;
  assign _1702_ = ~q[24] /*38299*/;
  assign _1703_ = sum_8[2] & q[24] /*38298*/;
  assign _1704_ = m_8[2] & _1702_ /*38297*/;
  assign r_8[26] = _1704_ | _1703_ /*38296*/;
  assign _1705_ = ~q[24] /*38295*/;
  assign _1706_ = sum_8[3] & q[24] /*38294*/;
  assign _1707_ = m_8[3] & _1705_ /*38293*/;
  assign r_8[27] = _1707_ | _1706_ /*38292*/;
  assign _1708_ = ~q[24] /*38291*/;
  assign _1709_ = sum_8[4] & q[24] /*38290*/;
  assign _1710_ = m_8[4] & _1708_ /*38289*/;
  assign r_8[28] = _1710_ | _1709_ /*38288*/;
  assign _1711_ = ~q[24] /*38287*/;
  assign _1712_ = sum_8[5] & q[24] /*38286*/;
  assign _1713_ = m_8[5] & _1711_ /*38285*/;
  assign r_8[29] = _1713_ | _1712_ /*38284*/;
  assign _1714_ = ~q[24] /*38283*/;
  assign _1715_ = sum_8[6] & q[24] /*38282*/;
  assign _1716_ = m_8[6] & _1714_ /*38281*/;
  assign r_8[30] = _1716_ | _1715_ /*38280*/;
  assign _1717_ = ~q[24] /*38279*/;
  assign _1718_ = sum_8[7] & q[24] /*38278*/;
  assign _1719_ = m_8[7] & _1717_ /*38277*/;
  assign r_8[31] = _1719_ | _1718_ /*38276*/;
  assign _1720_ = ~q[24] /*38275*/;
  assign _1721_ = sum_8[8] & q[24] /*38274*/;
  assign _1722_ = m_8[8] & _1720_ /*38273*/;
  assign r_8[32] = _1722_ | _1721_ /*38272*/;
  assign _1723_ = ~q[24] /*38271*/;
  assign _1724_ = sum_8[9] & q[24] /*38270*/;
  assign _1725_ = m_8[9] & _1723_ /*38269*/;
  assign r_8[33] = _1725_ | _1724_ /*38268*/;
  assign _1726_ = ~q[24] /*38267*/;
  assign _1727_ = sum_8[10] & q[24] /*38266*/;
  assign _1728_ = m_8[10] & _1726_ /*38265*/;
  assign r_8[34] = _1728_ | _1727_ /*38264*/;
  assign _1729_ = ~q[24] /*38263*/;
  assign _1730_ = sum_8[11] & q[24] /*38262*/;
  assign _1731_ = m_8[11] & _1729_ /*38261*/;
  assign r_8[35] = _1731_ | _1730_ /*38260*/;
  assign _1732_ = ~q[24] /*38259*/;
  assign _1733_ = sum_8[12] & q[24] /*38258*/;
  assign _1734_ = m_8[12] & _1732_ /*38257*/;
  assign r_8[36] = _1734_ | _1733_ /*38256*/;
  assign _1735_ = ~q[24] /*38255*/;
  assign _1736_ = sum_8[13] & q[24] /*38254*/;
  assign _1737_ = m_8[13] & _1735_ /*38253*/;
  assign r_8[37] = _1737_ | _1736_ /*38252*/;
  assign _1738_ = ~q[24] /*38251*/;
  assign _1739_ = sum_8[14] & q[24] /*38250*/;
  assign _1740_ = m_8[14] & _1738_ /*38249*/;
  assign r_8[38] = _1740_ | _1739_ /*38248*/;
  assign _1741_ = ~q[24] /*38247*/;
  assign _1742_ = sum_8[15] & q[24] /*38246*/;
  assign _1743_ = m_8[15] & _1741_ /*38245*/;
  assign r_8[39] = _1743_ | _1742_ /*38244*/;
  assign _1744_ = ~q[24] /*38243*/;
  assign _1745_ = sum_8[16] & q[24] /*38242*/;
  assign _1746_ = m_8[16] & _1744_ /*38241*/;
  assign r_8[40] = _1746_ | _1745_ /*38240*/;
  assign _1747_ = ~q[24] /*38239*/;
  assign _1748_ = sum_8[17] & q[24] /*38238*/;
  assign _1749_ = m_8[17] & _1747_ /*38237*/;
  assign r_8[41] = _1749_ | _1748_ /*38236*/;
  assign _1750_ = ~q[24] /*38235*/;
  assign _1751_ = sum_8[18] & q[24] /*38234*/;
  assign _1752_ = m_8[18] & _1750_ /*38233*/;
  assign r_8[42] = _1752_ | _1751_ /*38232*/;
  assign _1753_ = ~q[24] /*38231*/;
  assign _1754_ = sum_8[19] & q[24] /*38230*/;
  assign _1755_ = m_8[19] & _1753_ /*38229*/;
  assign r_8[43] = _1755_ | _1754_ /*38228*/;
  assign _1756_ = ~q[24] /*38227*/;
  assign _1757_ = sum_8[20] & q[24] /*38226*/;
  assign _1758_ = m_8[20] & _1756_ /*38225*/;
  assign r_8[44] = _1758_ | _1757_ /*38224*/;
  assign _1759_ = ~q[24] /*38223*/;
  assign _1760_ = sum_8[21] & q[24] /*38222*/;
  assign _1761_ = m_8[21] & _1759_ /*38221*/;
  assign r_8[45] = _1761_ | _1760_ /*38220*/;
  assign _1762_ = ~q[24] /*38219*/;
  assign _1763_ = sum_8[22] & q[24] /*38218*/;
  assign _1764_ = m_8[22] & _1762_ /*38217*/;
  assign r_8[46] = _1764_ | _1763_ /*38216*/;
  assign _1765_ = ~q[24] /*38215*/;
  assign _1766_ = sum_8[23] & q[24] /*38214*/;
  assign _1767_ = m_8[23] & _1765_ /*38213*/;
  assign r_8[47] = _1767_ | _1766_ /*38212*/;
  assign _1768_ = ~q[24] /*38211*/;
  assign _1769_ = sum_8[24] & q[24] /*38210*/;
  assign _1770_ = m_8[24] & _1768_ /*38209*/;
  assign r_8[48] = _1770_ | _1769_ /*38208*/;
  assign _1771_ = ~q[24] /*38207*/;
  assign _1772_ = sum_8[25] & q[24] /*38206*/;
  assign _1773_ = m_8[25] & _1771_ /*38205*/;
  assign r_8[49] = _1773_ | _1772_ /*38204*/;
  assign _1774_ = ~q[24] /*38203*/;
  assign _1775_ = sum_8[26] & q[24] /*38202*/;
  assign _1776_ = m_8[26] & _1774_ /*38201*/;
  assign r_8[50] = _1776_ | _1775_ /*38200*/;
  assign _1777_ = ~q[24] /*38199*/;
  assign _1778_ = sum_8[27] & q[24] /*38198*/;
  assign _1779_ = m_8[27] & _1777_ /*38197*/;
  assign r_8[51] = _1779_ | _1778_ /*38196*/;
  assign _1780_ = ~q[24] /*38195*/;
  assign _1781_ = sum_8[28] & q[24] /*38194*/;
  assign _1782_ = m_8[28] & _1780_ /*38193*/;
  assign r_8[52] = _1782_ | _1781_ /*38192*/;
  assign _1783_ = ~q[24] /*38191*/;
  assign _1784_ = sum_8[29] & q[24] /*38190*/;
  assign _1785_ = m_8[29] & _1783_ /*38189*/;
  assign r_8[53] = _1785_ | _1784_ /*38188*/;
  assign _1786_ = ~q[24] /*38187*/;
  assign _1787_ = sum_8[30] & q[24] /*38186*/;
  assign _1788_ = m_8[30] & _1786_ /*38185*/;
  assign r_8[54] = _1788_ | _1787_ /*38184*/;
  assign _1789_ = ~q[24] /*38183*/;
  assign _1790_ = sum_8[31] & q[24] /*38182*/;
  assign _1791_ = m_8[31] & _1789_ /*38181*/;
  assign r_8[55] = _1791_ | _1790_ /*38180*/;
assign r_8[0]= r_7[0] /*38179*/;
assign r_8[1]= r_7[1] /*38178*/;
assign r_8[2]= r_7[2] /*38177*/;
assign r_8[3]= r_7[3] /*38176*/;
assign r_8[4]= r_7[4] /*38175*/;
assign r_8[5]= r_7[5] /*38174*/;
assign r_8[6]= r_7[6] /*38173*/;
assign r_8[7]= r_7[7] /*38172*/;
assign r_8[8]= r_7[8] /*38171*/;
assign r_8[9]= r_7[9] /*38170*/;
assign r_8[10]= r_7[10] /*38169*/;
assign r_8[11]= r_7[11] /*38168*/;
assign r_8[12]= r_7[12] /*38167*/;
assign r_8[13]= r_7[13] /*38166*/;
assign r_8[14]= r_7[14] /*38165*/;
assign r_8[15]= r_7[15] /*38164*/;
assign r_8[16]= r_7[16] /*38163*/;
assign r_8[17]= r_7[17] /*38162*/;
assign r_8[18]= r_7[18] /*38161*/;
assign r_8[19]= r_7[19] /*38160*/;
assign r_8[20]= r_7[20] /*38159*/;
assign r_8[21]= r_7[21] /*38158*/;
assign r_8[22]= r_7[22] /*38157*/;
assign r_8[23]= r_7[23] /*38156*/;
  assign inv_9[0] = ~div[0] /*38088*/;
  assign inv_9[1] = ~div[1] /*38087*/;
  assign inv_9[2] = ~div[2] /*38086*/;
  assign inv_9[3] = ~div[3] /*38085*/;
  assign inv_9[4] = ~div[4] /*38084*/;
  assign inv_9[5] = ~div[5] /*38083*/;
  assign inv_9[6] = ~div[6] /*38082*/;
  assign inv_9[7] = ~div[7] /*38081*/;
  assign inv_9[8] = ~div[8] /*38080*/;
  assign inv_9[9] = ~div[9] /*38079*/;
  assign inv_9[10] = ~div[10] /*38078*/;
  assign inv_9[11] = ~div[11] /*38077*/;
  assign inv_9[12] = ~div[12] /*38076*/;
  assign inv_9[13] = ~div[13] /*38075*/;
  assign inv_9[14] = ~div[14] /*38074*/;
  assign inv_9[15] = ~div[15] /*38073*/;
  assign inv_9[16] = ~div[16] /*38072*/;
  assign inv_9[17] = ~div[17] /*38071*/;
  assign inv_9[18] = ~div[18] /*38070*/;
  assign inv_9[19] = ~div[19] /*38069*/;
  assign inv_9[20] = ~div[20] /*38068*/;
  assign inv_9[21] = ~div[21] /*38067*/;
  assign inv_9[22] = ~div[22] /*38066*/;
  assign inv_9[23] = ~div[23] /*38065*/;
  assign inv_9[24] = ~div[24] /*38064*/;
  assign inv_9[25] = ~div[25] /*38063*/;
  assign inv_9[26] = ~div[26] /*38062*/;
  assign inv_9[27] = ~div[27] /*38061*/;
  assign inv_9[28] = ~div[28] /*38060*/;
  assign inv_9[29] = ~div[29] /*38059*/;
  assign inv_9[30] = ~div[30] /*38058*/;
assign inv_9[31] = oneWire /*38057*/;
  assign _1792_ = inv_9[0] ^ r_8[23] /*38055*/;
  assign sum_9[0] = _1792_ ^ oneWire /*38054*/;
  assign _1793_ = _1792_ & oneWire /*38053*/;
  assign _1794_ = inv_9[0] & r_8[23] /*38052*/;
  assign _1795_ = _1793_ | _1794_ /*38051*/;
  assign _1796_ = inv_9[1] ^ r_8[24] /*38050*/;
  assign sum_9[1] = _1796_ ^ _1795_ /*38049*/;
  assign _1797_ = _1796_ & _1795_ /*38048*/;
  assign _1798_ = inv_9[1] & r_8[24] /*38047*/;
  assign _1799_ = _1797_ | _1798_ /*38046*/;
  assign _1800_ = inv_9[2] ^ r_8[25] /*38044*/;
  assign sum_9[2] = _1800_ ^ _1799_ /*38043*/;
  assign _1801_ = _1800_ & _1799_ /*38042*/;
  assign _1802_ = inv_9[2] & r_8[25] /*38041*/;
  assign _1803_ = _1801_ | _1802_ /*38040*/;
  assign _1804_ = inv_9[3] ^ r_8[26] /*38038*/;
  assign sum_9[3] = _1804_ ^ _1803_ /*38037*/;
  assign _1805_ = _1804_ & _1803_ /*38036*/;
  assign _1806_ = inv_9[3] & r_8[26] /*38035*/;
  assign _1807_ = _1805_ | _1806_ /*38034*/;
  assign _1808_ = inv_9[4] ^ r_8[27] /*38032*/;
  assign sum_9[4] = _1808_ ^ _1807_ /*38031*/;
  assign _1809_ = _1808_ & _1807_ /*38030*/;
  assign _1810_ = inv_9[4] & r_8[27] /*38029*/;
  assign _1811_ = _1809_ | _1810_ /*38028*/;
  assign _1812_ = inv_9[5] ^ r_8[28] /*38026*/;
  assign sum_9[5] = _1812_ ^ _1811_ /*38025*/;
  assign _1813_ = _1812_ & _1811_ /*38024*/;
  assign _1814_ = inv_9[5] & r_8[28] /*38023*/;
  assign _1815_ = _1813_ | _1814_ /*38022*/;
  assign _1816_ = inv_9[6] ^ r_8[29] /*38020*/;
  assign sum_9[6] = _1816_ ^ _1815_ /*38019*/;
  assign _1817_ = _1816_ & _1815_ /*38018*/;
  assign _1818_ = inv_9[6] & r_8[29] /*38017*/;
  assign _1819_ = _1817_ | _1818_ /*38016*/;
  assign _1820_ = inv_9[7] ^ r_8[30] /*38014*/;
  assign sum_9[7] = _1820_ ^ _1819_ /*38013*/;
  assign _1821_ = _1820_ & _1819_ /*38012*/;
  assign _1822_ = inv_9[7] & r_8[30] /*38011*/;
  assign _1823_ = _1821_ | _1822_ /*38010*/;
  assign _1824_ = inv_9[8] ^ r_8[31] /*38008*/;
  assign sum_9[8] = _1824_ ^ _1823_ /*38007*/;
  assign _1825_ = _1824_ & _1823_ /*38006*/;
  assign _1826_ = inv_9[8] & r_8[31] /*38005*/;
  assign _1827_ = _1825_ | _1826_ /*38004*/;
  assign _1828_ = inv_9[9] ^ r_8[32] /*38002*/;
  assign sum_9[9] = _1828_ ^ _1827_ /*38001*/;
  assign _1829_ = _1828_ & _1827_ /*38000*/;
  assign _1830_ = inv_9[9] & r_8[32] /*37999*/;
  assign _1831_ = _1829_ | _1830_ /*37998*/;
  assign _1832_ = inv_9[10] ^ r_8[33] /*37996*/;
  assign sum_9[10] = _1832_ ^ _1831_ /*37995*/;
  assign _1833_ = _1832_ & _1831_ /*37994*/;
  assign _1834_ = inv_9[10] & r_8[33] /*37993*/;
  assign _1835_ = _1833_ | _1834_ /*37992*/;
  assign _1836_ = inv_9[11] ^ r_8[34] /*37990*/;
  assign sum_9[11] = _1836_ ^ _1835_ /*37989*/;
  assign _1837_ = _1836_ & _1835_ /*37988*/;
  assign _1838_ = inv_9[11] & r_8[34] /*37987*/;
  assign _1839_ = _1837_ | _1838_ /*37986*/;
  assign _1840_ = inv_9[12] ^ r_8[35] /*37984*/;
  assign sum_9[12] = _1840_ ^ _1839_ /*37983*/;
  assign _1841_ = _1840_ & _1839_ /*37982*/;
  assign _1842_ = inv_9[12] & r_8[35] /*37981*/;
  assign _1843_ = _1841_ | _1842_ /*37980*/;
  assign _1844_ = inv_9[13] ^ r_8[36] /*37978*/;
  assign sum_9[13] = _1844_ ^ _1843_ /*37977*/;
  assign _1845_ = _1844_ & _1843_ /*37976*/;
  assign _1846_ = inv_9[13] & r_8[36] /*37975*/;
  assign _1847_ = _1845_ | _1846_ /*37974*/;
  assign _1848_ = inv_9[14] ^ r_8[37] /*37972*/;
  assign sum_9[14] = _1848_ ^ _1847_ /*37971*/;
  assign _1849_ = _1848_ & _1847_ /*37970*/;
  assign _1850_ = inv_9[14] & r_8[37] /*37969*/;
  assign _1851_ = _1849_ | _1850_ /*37968*/;
  assign _1852_ = inv_9[15] ^ r_8[38] /*37966*/;
  assign sum_9[15] = _1852_ ^ _1851_ /*37965*/;
  assign _1853_ = _1852_ & _1851_ /*37964*/;
  assign _1854_ = inv_9[15] & r_8[38] /*37963*/;
  assign _1855_ = _1853_ | _1854_ /*37962*/;
  assign _1856_ = inv_9[16] ^ r_8[39] /*37960*/;
  assign sum_9[16] = _1856_ ^ _1855_ /*37959*/;
  assign _1857_ = _1856_ & _1855_ /*37958*/;
  assign _1858_ = inv_9[16] & r_8[39] /*37957*/;
  assign _1859_ = _1857_ | _1858_ /*37956*/;
  assign _1860_ = inv_9[17] ^ r_8[40] /*37954*/;
  assign sum_9[17] = _1860_ ^ _1859_ /*37953*/;
  assign _1861_ = _1860_ & _1859_ /*37952*/;
  assign _1862_ = inv_9[17] & r_8[40] /*37951*/;
  assign _1863_ = _1861_ | _1862_ /*37950*/;
  assign _1864_ = inv_9[18] ^ r_8[41] /*37948*/;
  assign sum_9[18] = _1864_ ^ _1863_ /*37947*/;
  assign _1865_ = _1864_ & _1863_ /*37946*/;
  assign _1866_ = inv_9[18] & r_8[41] /*37945*/;
  assign _1867_ = _1865_ | _1866_ /*37944*/;
  assign _1868_ = inv_9[19] ^ r_8[42] /*37942*/;
  assign sum_9[19] = _1868_ ^ _1867_ /*37941*/;
  assign _1869_ = _1868_ & _1867_ /*37940*/;
  assign _1870_ = inv_9[19] & r_8[42] /*37939*/;
  assign _1871_ = _1869_ | _1870_ /*37938*/;
  assign _1872_ = inv_9[20] ^ r_8[43] /*37936*/;
  assign sum_9[20] = _1872_ ^ _1871_ /*37935*/;
  assign _1873_ = _1872_ & _1871_ /*37934*/;
  assign _1874_ = inv_9[20] & r_8[43] /*37933*/;
  assign _1875_ = _1873_ | _1874_ /*37932*/;
  assign _1876_ = inv_9[21] ^ r_8[44] /*37930*/;
  assign sum_9[21] = _1876_ ^ _1875_ /*37929*/;
  assign _1877_ = _1876_ & _1875_ /*37928*/;
  assign _1878_ = inv_9[21] & r_8[44] /*37927*/;
  assign _1879_ = _1877_ | _1878_ /*37926*/;
  assign _1880_ = inv_9[22] ^ r_8[45] /*37924*/;
  assign sum_9[22] = _1880_ ^ _1879_ /*37923*/;
  assign _1881_ = _1880_ & _1879_ /*37922*/;
  assign _1882_ = inv_9[22] & r_8[45] /*37921*/;
  assign _1883_ = _1881_ | _1882_ /*37920*/;
  assign _1884_ = inv_9[23] ^ r_8[46] /*37918*/;
  assign sum_9[23] = _1884_ ^ _1883_ /*37917*/;
  assign _1885_ = _1884_ & _1883_ /*37916*/;
  assign _1886_ = inv_9[23] & r_8[46] /*37915*/;
  assign _1887_ = _1885_ | _1886_ /*37914*/;
  assign _1888_ = inv_9[24] ^ r_8[47] /*37912*/;
  assign sum_9[24] = _1888_ ^ _1887_ /*37911*/;
  assign _1889_ = _1888_ & _1887_ /*37910*/;
  assign _1890_ = inv_9[24] & r_8[47] /*37909*/;
  assign _1891_ = _1889_ | _1890_ /*37908*/;
  assign _1892_ = inv_9[25] ^ r_8[48] /*37906*/;
  assign sum_9[25] = _1892_ ^ _1891_ /*37905*/;
  assign _1893_ = _1892_ & _1891_ /*37904*/;
  assign _1894_ = inv_9[25] & r_8[48] /*37903*/;
  assign _1895_ = _1893_ | _1894_ /*37902*/;
  assign _1896_ = inv_9[26] ^ r_8[49] /*37900*/;
  assign sum_9[26] = _1896_ ^ _1895_ /*37899*/;
  assign _1897_ = _1896_ & _1895_ /*37898*/;
  assign _1898_ = inv_9[26] & r_8[49] /*37897*/;
  assign _1899_ = _1897_ | _1898_ /*37896*/;
  assign _1900_ = inv_9[27] ^ r_8[50] /*37894*/;
  assign sum_9[27] = _1900_ ^ _1899_ /*37893*/;
  assign _1901_ = _1900_ & _1899_ /*37892*/;
  assign _1902_ = inv_9[27] & r_8[50] /*37891*/;
  assign _1903_ = _1901_ | _1902_ /*37890*/;
  assign _1904_ = inv_9[28] ^ r_8[51] /*37888*/;
  assign sum_9[28] = _1904_ ^ _1903_ /*37887*/;
  assign _1905_ = _1904_ & _1903_ /*37886*/;
  assign _1906_ = inv_9[28] & r_8[51] /*37885*/;
  assign _1907_ = _1905_ | _1906_ /*37884*/;
  assign _1908_ = inv_9[29] ^ r_8[52] /*37882*/;
  assign sum_9[29] = _1908_ ^ _1907_ /*37881*/;
  assign _1909_ = _1908_ & _1907_ /*37880*/;
  assign _1910_ = inv_9[29] & r_8[52] /*37879*/;
  assign _1911_ = _1909_ | _1910_ /*37878*/;
  assign _1912_ = inv_9[30] ^ r_8[53] /*37876*/;
  assign sum_9[30] = _1912_ ^ _1911_ /*37875*/;
  assign _1913_ = _1912_ & _1911_ /*37874*/;
  assign _1914_ = inv_9[30] & r_8[53] /*37873*/;
  assign _1915_ = _1913_ | _1914_ /*37872*/;
  assign _1916_ = inv_9[31] ^ r_8[54] /*37870*/;
  assign sum_9[31] = _1916_ ^ _1915_ /*37869*/;
  assign _1917_ = _1916_ & _1915_ /*37868*/;
  assign _1918_ = inv_9[31] & r_8[54] /*37867*/;
  assign _1919_ = _1917_ | _1918_ /*37866*/;
  assign q[23] = ~sum_9[31] /*37893*/;
  assign m_9[0] = r_8[23] /*37892*/;
  assign m_9[1] = r_8[24] /*37891*/;
  assign m_9[2] = r_8[25] /*37890*/;
  assign m_9[3] = r_8[26] /*37889*/;
  assign m_9[4] = r_8[27] /*37888*/;
  assign m_9[5] = r_8[28] /*37887*/;
  assign m_9[6] = r_8[29] /*37886*/;
  assign m_9[7] = r_8[30] /*37885*/;
  assign m_9[8] = r_8[31] /*37884*/;
  assign m_9[9] = r_8[32] /*37883*/;
  assign m_9[10] = r_8[33] /*37882*/;
  assign m_9[11] = r_8[34] /*37881*/;
  assign m_9[12] = r_8[35] /*37880*/;
  assign m_9[13] = r_8[36] /*37879*/;
  assign m_9[14] = r_8[37] /*37878*/;
  assign m_9[15] = r_8[38] /*37877*/;
  assign m_9[16] = r_8[39] /*37876*/;
  assign m_9[17] = r_8[40] /*37875*/;
  assign m_9[18] = r_8[41] /*37874*/;
  assign m_9[19] = r_8[42] /*37873*/;
  assign m_9[20] = r_8[43] /*37872*/;
  assign m_9[21] = r_8[44] /*37871*/;
  assign m_9[22] = r_8[45] /*37870*/;
  assign m_9[23] = r_8[46] /*37869*/;
  assign m_9[24] = r_8[47] /*37868*/;
  assign m_9[25] = r_8[48] /*37867*/;
  assign m_9[26] = r_8[49] /*37866*/;
  assign m_9[27] = r_8[50] /*37865*/;
  assign m_9[28] = r_8[51] /*37864*/;
  assign m_9[29] = r_8[52] /*37863*/;
  assign m_9[30] = r_8[53] /*37862*/;
  assign m_9[31] = r_8[54] /*37861*/;
  assign _1920_ = ~q[23] /*37859*/;
  assign _1921_ = sum_9[0] & q[23] /*37858*/;
  assign _1922_ = m_9[0] & _1920_ /*37857*/;
  assign r_9[23] = _1922_ | _1921_ /*37856*/;
  assign _1923_ = ~q[23] /*37855*/;
  assign _1924_ = sum_9[1] & q[23] /*37854*/;
  assign _1925_ = m_9[1] & _1923_ /*37853*/;
  assign r_9[24] = _1925_ | _1924_ /*37852*/;
  assign _1926_ = ~q[23] /*37851*/;
  assign _1927_ = sum_9[2] & q[23] /*37850*/;
  assign _1928_ = m_9[2] & _1926_ /*37849*/;
  assign r_9[25] = _1928_ | _1927_ /*37848*/;
  assign _1929_ = ~q[23] /*37847*/;
  assign _1930_ = sum_9[3] & q[23] /*37846*/;
  assign _1931_ = m_9[3] & _1929_ /*37845*/;
  assign r_9[26] = _1931_ | _1930_ /*37844*/;
  assign _1932_ = ~q[23] /*37843*/;
  assign _1933_ = sum_9[4] & q[23] /*37842*/;
  assign _1934_ = m_9[4] & _1932_ /*37841*/;
  assign r_9[27] = _1934_ | _1933_ /*37840*/;
  assign _1935_ = ~q[23] /*37839*/;
  assign _1936_ = sum_9[5] & q[23] /*37838*/;
  assign _1937_ = m_9[5] & _1935_ /*37837*/;
  assign r_9[28] = _1937_ | _1936_ /*37836*/;
  assign _1938_ = ~q[23] /*37835*/;
  assign _1939_ = sum_9[6] & q[23] /*37834*/;
  assign _1940_ = m_9[6] & _1938_ /*37833*/;
  assign r_9[29] = _1940_ | _1939_ /*37832*/;
  assign _1941_ = ~q[23] /*37831*/;
  assign _1942_ = sum_9[7] & q[23] /*37830*/;
  assign _1943_ = m_9[7] & _1941_ /*37829*/;
  assign r_9[30] = _1943_ | _1942_ /*37828*/;
  assign _1944_ = ~q[23] /*37827*/;
  assign _1945_ = sum_9[8] & q[23] /*37826*/;
  assign _1946_ = m_9[8] & _1944_ /*37825*/;
  assign r_9[31] = _1946_ | _1945_ /*37824*/;
  assign _1947_ = ~q[23] /*37823*/;
  assign _1948_ = sum_9[9] & q[23] /*37822*/;
  assign _1949_ = m_9[9] & _1947_ /*37821*/;
  assign r_9[32] = _1949_ | _1948_ /*37820*/;
  assign _1950_ = ~q[23] /*37819*/;
  assign _1951_ = sum_9[10] & q[23] /*37818*/;
  assign _1952_ = m_9[10] & _1950_ /*37817*/;
  assign r_9[33] = _1952_ | _1951_ /*37816*/;
  assign _1953_ = ~q[23] /*37815*/;
  assign _1954_ = sum_9[11] & q[23] /*37814*/;
  assign _1955_ = m_9[11] & _1953_ /*37813*/;
  assign r_9[34] = _1955_ | _1954_ /*37812*/;
  assign _1956_ = ~q[23] /*37811*/;
  assign _1957_ = sum_9[12] & q[23] /*37810*/;
  assign _1958_ = m_9[12] & _1956_ /*37809*/;
  assign r_9[35] = _1958_ | _1957_ /*37808*/;
  assign _1959_ = ~q[23] /*37807*/;
  assign _1960_ = sum_9[13] & q[23] /*37806*/;
  assign _1961_ = m_9[13] & _1959_ /*37805*/;
  assign r_9[36] = _1961_ | _1960_ /*37804*/;
  assign _1962_ = ~q[23] /*37803*/;
  assign _1963_ = sum_9[14] & q[23] /*37802*/;
  assign _1964_ = m_9[14] & _1962_ /*37801*/;
  assign r_9[37] = _1964_ | _1963_ /*37800*/;
  assign _1965_ = ~q[23] /*37799*/;
  assign _1966_ = sum_9[15] & q[23] /*37798*/;
  assign _1967_ = m_9[15] & _1965_ /*37797*/;
  assign r_9[38] = _1967_ | _1966_ /*37796*/;
  assign _1968_ = ~q[23] /*37795*/;
  assign _1969_ = sum_9[16] & q[23] /*37794*/;
  assign _1970_ = m_9[16] & _1968_ /*37793*/;
  assign r_9[39] = _1970_ | _1969_ /*37792*/;
  assign _1971_ = ~q[23] /*37791*/;
  assign _1972_ = sum_9[17] & q[23] /*37790*/;
  assign _1973_ = m_9[17] & _1971_ /*37789*/;
  assign r_9[40] = _1973_ | _1972_ /*37788*/;
  assign _1974_ = ~q[23] /*37787*/;
  assign _1975_ = sum_9[18] & q[23] /*37786*/;
  assign _1976_ = m_9[18] & _1974_ /*37785*/;
  assign r_9[41] = _1976_ | _1975_ /*37784*/;
  assign _1977_ = ~q[23] /*37783*/;
  assign _1978_ = sum_9[19] & q[23] /*37782*/;
  assign _1979_ = m_9[19] & _1977_ /*37781*/;
  assign r_9[42] = _1979_ | _1978_ /*37780*/;
  assign _1980_ = ~q[23] /*37779*/;
  assign _1981_ = sum_9[20] & q[23] /*37778*/;
  assign _1982_ = m_9[20] & _1980_ /*37777*/;
  assign r_9[43] = _1982_ | _1981_ /*37776*/;
  assign _1983_ = ~q[23] /*37775*/;
  assign _1984_ = sum_9[21] & q[23] /*37774*/;
  assign _1985_ = m_9[21] & _1983_ /*37773*/;
  assign r_9[44] = _1985_ | _1984_ /*37772*/;
  assign _1986_ = ~q[23] /*37771*/;
  assign _1987_ = sum_9[22] & q[23] /*37770*/;
  assign _1988_ = m_9[22] & _1986_ /*37769*/;
  assign r_9[45] = _1988_ | _1987_ /*37768*/;
  assign _1989_ = ~q[23] /*37767*/;
  assign _1990_ = sum_9[23] & q[23] /*37766*/;
  assign _1991_ = m_9[23] & _1989_ /*37765*/;
  assign r_9[46] = _1991_ | _1990_ /*37764*/;
  assign _1992_ = ~q[23] /*37763*/;
  assign _1993_ = sum_9[24] & q[23] /*37762*/;
  assign _1994_ = m_9[24] & _1992_ /*37761*/;
  assign r_9[47] = _1994_ | _1993_ /*37760*/;
  assign _1995_ = ~q[23] /*37759*/;
  assign _1996_ = sum_9[25] & q[23] /*37758*/;
  assign _1997_ = m_9[25] & _1995_ /*37757*/;
  assign r_9[48] = _1997_ | _1996_ /*37756*/;
  assign _1998_ = ~q[23] /*37755*/;
  assign _1999_ = sum_9[26] & q[23] /*37754*/;
  assign _2000_ = m_9[26] & _1998_ /*37753*/;
  assign r_9[49] = _2000_ | _1999_ /*37752*/;
  assign _2001_ = ~q[23] /*37751*/;
  assign _2002_ = sum_9[27] & q[23] /*37750*/;
  assign _2003_ = m_9[27] & _2001_ /*37749*/;
  assign r_9[50] = _2003_ | _2002_ /*37748*/;
  assign _2004_ = ~q[23] /*37747*/;
  assign _2005_ = sum_9[28] & q[23] /*37746*/;
  assign _2006_ = m_9[28] & _2004_ /*37745*/;
  assign r_9[51] = _2006_ | _2005_ /*37744*/;
  assign _2007_ = ~q[23] /*37743*/;
  assign _2008_ = sum_9[29] & q[23] /*37742*/;
  assign _2009_ = m_9[29] & _2007_ /*37741*/;
  assign r_9[52] = _2009_ | _2008_ /*37740*/;
  assign _2010_ = ~q[23] /*37739*/;
  assign _2011_ = sum_9[30] & q[23] /*37738*/;
  assign _2012_ = m_9[30] & _2010_ /*37737*/;
  assign r_9[53] = _2012_ | _2011_ /*37736*/;
  assign _2013_ = ~q[23] /*37735*/;
  assign _2014_ = sum_9[31] & q[23] /*37734*/;
  assign _2015_ = m_9[31] & _2013_ /*37733*/;
  assign r_9[54] = _2015_ | _2014_ /*37732*/;
assign r_9[0]= r_8[0] /*37731*/;
assign r_9[1]= r_8[1] /*37730*/;
assign r_9[2]= r_8[2] /*37729*/;
assign r_9[3]= r_8[3] /*37728*/;
assign r_9[4]= r_8[4] /*37727*/;
assign r_9[5]= r_8[5] /*37726*/;
assign r_9[6]= r_8[6] /*37725*/;
assign r_9[7]= r_8[7] /*37724*/;
assign r_9[8]= r_8[8] /*37723*/;
assign r_9[9]= r_8[9] /*37722*/;
assign r_9[10]= r_8[10] /*37721*/;
assign r_9[11]= r_8[11] /*37720*/;
assign r_9[12]= r_8[12] /*37719*/;
assign r_9[13]= r_8[13] /*37718*/;
assign r_9[14]= r_8[14] /*37717*/;
assign r_9[15]= r_8[15] /*37716*/;
assign r_9[16]= r_8[16] /*37715*/;
assign r_9[17]= r_8[17] /*37714*/;
assign r_9[18]= r_8[18] /*37713*/;
assign r_9[19]= r_8[19] /*37712*/;
assign r_9[20]= r_8[20] /*37711*/;
assign r_9[21]= r_8[21] /*37710*/;
assign r_9[22]= r_8[22] /*37709*/;
  assign inv_10[0] = ~div[0] /*37640*/;
  assign inv_10[1] = ~div[1] /*37639*/;
  assign inv_10[2] = ~div[2] /*37638*/;
  assign inv_10[3] = ~div[3] /*37637*/;
  assign inv_10[4] = ~div[4] /*37636*/;
  assign inv_10[5] = ~div[5] /*37635*/;
  assign inv_10[6] = ~div[6] /*37634*/;
  assign inv_10[7] = ~div[7] /*37633*/;
  assign inv_10[8] = ~div[8] /*37632*/;
  assign inv_10[9] = ~div[9] /*37631*/;
  assign inv_10[10] = ~div[10] /*37630*/;
  assign inv_10[11] = ~div[11] /*37629*/;
  assign inv_10[12] = ~div[12] /*37628*/;
  assign inv_10[13] = ~div[13] /*37627*/;
  assign inv_10[14] = ~div[14] /*37626*/;
  assign inv_10[15] = ~div[15] /*37625*/;
  assign inv_10[16] = ~div[16] /*37624*/;
  assign inv_10[17] = ~div[17] /*37623*/;
  assign inv_10[18] = ~div[18] /*37622*/;
  assign inv_10[19] = ~div[19] /*37621*/;
  assign inv_10[20] = ~div[20] /*37620*/;
  assign inv_10[21] = ~div[21] /*37619*/;
  assign inv_10[22] = ~div[22] /*37618*/;
  assign inv_10[23] = ~div[23] /*37617*/;
  assign inv_10[24] = ~div[24] /*37616*/;
  assign inv_10[25] = ~div[25] /*37615*/;
  assign inv_10[26] = ~div[26] /*37614*/;
  assign inv_10[27] = ~div[27] /*37613*/;
  assign inv_10[28] = ~div[28] /*37612*/;
  assign inv_10[29] = ~div[29] /*37611*/;
  assign inv_10[30] = ~div[30] /*37610*/;
assign inv_10[31] = oneWire /*37609*/;
  assign _2016_ = inv_10[0] ^ r_9[22] /*37607*/;
  assign sum_10[0] = _2016_ ^ oneWire /*37606*/;
  assign _2017_ = _2016_ & oneWire /*37605*/;
  assign _2018_ = inv_10[0] & r_9[22] /*37604*/;
  assign _2019_ = _2017_ | _2018_ /*37603*/;
  assign _2020_ = inv_10[1] ^ r_9[23] /*37602*/;
  assign sum_10[1] = _2020_ ^ _2019_ /*37601*/;
  assign _2021_ = _2020_ & _2019_ /*37600*/;
  assign _2022_ = inv_10[1] & r_9[23] /*37599*/;
  assign _2023_ = _2021_ | _2022_ /*37598*/;
  assign _2024_ = inv_10[2] ^ r_9[24] /*37596*/;
  assign sum_10[2] = _2024_ ^ _2023_ /*37595*/;
  assign _2025_ = _2024_ & _2023_ /*37594*/;
  assign _2026_ = inv_10[2] & r_9[24] /*37593*/;
  assign _2027_ = _2025_ | _2026_ /*37592*/;
  assign _2028_ = inv_10[3] ^ r_9[25] /*37590*/;
  assign sum_10[3] = _2028_ ^ _2027_ /*37589*/;
  assign _2029_ = _2028_ & _2027_ /*37588*/;
  assign _2030_ = inv_10[3] & r_9[25] /*37587*/;
  assign _2031_ = _2029_ | _2030_ /*37586*/;
  assign _2032_ = inv_10[4] ^ r_9[26] /*37584*/;
  assign sum_10[4] = _2032_ ^ _2031_ /*37583*/;
  assign _2033_ = _2032_ & _2031_ /*37582*/;
  assign _2034_ = inv_10[4] & r_9[26] /*37581*/;
  assign _2035_ = _2033_ | _2034_ /*37580*/;
  assign _2036_ = inv_10[5] ^ r_9[27] /*37578*/;
  assign sum_10[5] = _2036_ ^ _2035_ /*37577*/;
  assign _2037_ = _2036_ & _2035_ /*37576*/;
  assign _2038_ = inv_10[5] & r_9[27] /*37575*/;
  assign _2039_ = _2037_ | _2038_ /*37574*/;
  assign _2040_ = inv_10[6] ^ r_9[28] /*37572*/;
  assign sum_10[6] = _2040_ ^ _2039_ /*37571*/;
  assign _2041_ = _2040_ & _2039_ /*37570*/;
  assign _2042_ = inv_10[6] & r_9[28] /*37569*/;
  assign _2043_ = _2041_ | _2042_ /*37568*/;
  assign _2044_ = inv_10[7] ^ r_9[29] /*37566*/;
  assign sum_10[7] = _2044_ ^ _2043_ /*37565*/;
  assign _2045_ = _2044_ & _2043_ /*37564*/;
  assign _2046_ = inv_10[7] & r_9[29] /*37563*/;
  assign _2047_ = _2045_ | _2046_ /*37562*/;
  assign _2048_ = inv_10[8] ^ r_9[30] /*37560*/;
  assign sum_10[8] = _2048_ ^ _2047_ /*37559*/;
  assign _2049_ = _2048_ & _2047_ /*37558*/;
  assign _2050_ = inv_10[8] & r_9[30] /*37557*/;
  assign _2051_ = _2049_ | _2050_ /*37556*/;
  assign _2052_ = inv_10[9] ^ r_9[31] /*37554*/;
  assign sum_10[9] = _2052_ ^ _2051_ /*37553*/;
  assign _2053_ = _2052_ & _2051_ /*37552*/;
  assign _2054_ = inv_10[9] & r_9[31] /*37551*/;
  assign _2055_ = _2053_ | _2054_ /*37550*/;
  assign _2056_ = inv_10[10] ^ r_9[32] /*37548*/;
  assign sum_10[10] = _2056_ ^ _2055_ /*37547*/;
  assign _2057_ = _2056_ & _2055_ /*37546*/;
  assign _2058_ = inv_10[10] & r_9[32] /*37545*/;
  assign _2059_ = _2057_ | _2058_ /*37544*/;
  assign _2060_ = inv_10[11] ^ r_9[33] /*37542*/;
  assign sum_10[11] = _2060_ ^ _2059_ /*37541*/;
  assign _2061_ = _2060_ & _2059_ /*37540*/;
  assign _2062_ = inv_10[11] & r_9[33] /*37539*/;
  assign _2063_ = _2061_ | _2062_ /*37538*/;
  assign _2064_ = inv_10[12] ^ r_9[34] /*37536*/;
  assign sum_10[12] = _2064_ ^ _2063_ /*37535*/;
  assign _2065_ = _2064_ & _2063_ /*37534*/;
  assign _2066_ = inv_10[12] & r_9[34] /*37533*/;
  assign _2067_ = _2065_ | _2066_ /*37532*/;
  assign _2068_ = inv_10[13] ^ r_9[35] /*37530*/;
  assign sum_10[13] = _2068_ ^ _2067_ /*37529*/;
  assign _2069_ = _2068_ & _2067_ /*37528*/;
  assign _2070_ = inv_10[13] & r_9[35] /*37527*/;
  assign _2071_ = _2069_ | _2070_ /*37526*/;
  assign _2072_ = inv_10[14] ^ r_9[36] /*37524*/;
  assign sum_10[14] = _2072_ ^ _2071_ /*37523*/;
  assign _2073_ = _2072_ & _2071_ /*37522*/;
  assign _2074_ = inv_10[14] & r_9[36] /*37521*/;
  assign _2075_ = _2073_ | _2074_ /*37520*/;
  assign _2076_ = inv_10[15] ^ r_9[37] /*37518*/;
  assign sum_10[15] = _2076_ ^ _2075_ /*37517*/;
  assign _2077_ = _2076_ & _2075_ /*37516*/;
  assign _2078_ = inv_10[15] & r_9[37] /*37515*/;
  assign _2079_ = _2077_ | _2078_ /*37514*/;
  assign _2080_ = inv_10[16] ^ r_9[38] /*37512*/;
  assign sum_10[16] = _2080_ ^ _2079_ /*37511*/;
  assign _2081_ = _2080_ & _2079_ /*37510*/;
  assign _2082_ = inv_10[16] & r_9[38] /*37509*/;
  assign _2083_ = _2081_ | _2082_ /*37508*/;
  assign _2084_ = inv_10[17] ^ r_9[39] /*37506*/;
  assign sum_10[17] = _2084_ ^ _2083_ /*37505*/;
  assign _2085_ = _2084_ & _2083_ /*37504*/;
  assign _2086_ = inv_10[17] & r_9[39] /*37503*/;
  assign _2087_ = _2085_ | _2086_ /*37502*/;
  assign _2088_ = inv_10[18] ^ r_9[40] /*37500*/;
  assign sum_10[18] = _2088_ ^ _2087_ /*37499*/;
  assign _2089_ = _2088_ & _2087_ /*37498*/;
  assign _2090_ = inv_10[18] & r_9[40] /*37497*/;
  assign _2091_ = _2089_ | _2090_ /*37496*/;
  assign _2092_ = inv_10[19] ^ r_9[41] /*37494*/;
  assign sum_10[19] = _2092_ ^ _2091_ /*37493*/;
  assign _2093_ = _2092_ & _2091_ /*37492*/;
  assign _2094_ = inv_10[19] & r_9[41] /*37491*/;
  assign _2095_ = _2093_ | _2094_ /*37490*/;
  assign _2096_ = inv_10[20] ^ r_9[42] /*37488*/;
  assign sum_10[20] = _2096_ ^ _2095_ /*37487*/;
  assign _2097_ = _2096_ & _2095_ /*37486*/;
  assign _2098_ = inv_10[20] & r_9[42] /*37485*/;
  assign _2099_ = _2097_ | _2098_ /*37484*/;
  assign _2100_ = inv_10[21] ^ r_9[43] /*37482*/;
  assign sum_10[21] = _2100_ ^ _2099_ /*37481*/;
  assign _2101_ = _2100_ & _2099_ /*37480*/;
  assign _2102_ = inv_10[21] & r_9[43] /*37479*/;
  assign _2103_ = _2101_ | _2102_ /*37478*/;
  assign _2104_ = inv_10[22] ^ r_9[44] /*37476*/;
  assign sum_10[22] = _2104_ ^ _2103_ /*37475*/;
  assign _2105_ = _2104_ & _2103_ /*37474*/;
  assign _2106_ = inv_10[22] & r_9[44] /*37473*/;
  assign _2107_ = _2105_ | _2106_ /*37472*/;
  assign _2108_ = inv_10[23] ^ r_9[45] /*37470*/;
  assign sum_10[23] = _2108_ ^ _2107_ /*37469*/;
  assign _2109_ = _2108_ & _2107_ /*37468*/;
  assign _2110_ = inv_10[23] & r_9[45] /*37467*/;
  assign _2111_ = _2109_ | _2110_ /*37466*/;
  assign _2112_ = inv_10[24] ^ r_9[46] /*37464*/;
  assign sum_10[24] = _2112_ ^ _2111_ /*37463*/;
  assign _2113_ = _2112_ & _2111_ /*37462*/;
  assign _2114_ = inv_10[24] & r_9[46] /*37461*/;
  assign _2115_ = _2113_ | _2114_ /*37460*/;
  assign _2116_ = inv_10[25] ^ r_9[47] /*37458*/;
  assign sum_10[25] = _2116_ ^ _2115_ /*37457*/;
  assign _2117_ = _2116_ & _2115_ /*37456*/;
  assign _2118_ = inv_10[25] & r_9[47] /*37455*/;
  assign _2119_ = _2117_ | _2118_ /*37454*/;
  assign _2120_ = inv_10[26] ^ r_9[48] /*37452*/;
  assign sum_10[26] = _2120_ ^ _2119_ /*37451*/;
  assign _2121_ = _2120_ & _2119_ /*37450*/;
  assign _2122_ = inv_10[26] & r_9[48] /*37449*/;
  assign _2123_ = _2121_ | _2122_ /*37448*/;
  assign _2124_ = inv_10[27] ^ r_9[49] /*37446*/;
  assign sum_10[27] = _2124_ ^ _2123_ /*37445*/;
  assign _2125_ = _2124_ & _2123_ /*37444*/;
  assign _2126_ = inv_10[27] & r_9[49] /*37443*/;
  assign _2127_ = _2125_ | _2126_ /*37442*/;
  assign _2128_ = inv_10[28] ^ r_9[50] /*37440*/;
  assign sum_10[28] = _2128_ ^ _2127_ /*37439*/;
  assign _2129_ = _2128_ & _2127_ /*37438*/;
  assign _2130_ = inv_10[28] & r_9[50] /*37437*/;
  assign _2131_ = _2129_ | _2130_ /*37436*/;
  assign _2132_ = inv_10[29] ^ r_9[51] /*37434*/;
  assign sum_10[29] = _2132_ ^ _2131_ /*37433*/;
  assign _2133_ = _2132_ & _2131_ /*37432*/;
  assign _2134_ = inv_10[29] & r_9[51] /*37431*/;
  assign _2135_ = _2133_ | _2134_ /*37430*/;
  assign _2136_ = inv_10[30] ^ r_9[52] /*37428*/;
  assign sum_10[30] = _2136_ ^ _2135_ /*37427*/;
  assign _2137_ = _2136_ & _2135_ /*37426*/;
  assign _2138_ = inv_10[30] & r_9[52] /*37425*/;
  assign _2139_ = _2137_ | _2138_ /*37424*/;
  assign _2140_ = inv_10[31] ^ r_9[53] /*37422*/;
  assign sum_10[31] = _2140_ ^ _2139_ /*37421*/;
  assign _2141_ = _2140_ & _2139_ /*37420*/;
  assign _2142_ = inv_10[31] & r_9[53] /*37419*/;
  assign _2143_ = _2141_ | _2142_ /*37418*/;
  assign q[22] = ~sum_10[31] /*37445*/;
  assign m_10[0] = r_9[22] /*37444*/;
  assign m_10[1] = r_9[23] /*37443*/;
  assign m_10[2] = r_9[24] /*37442*/;
  assign m_10[3] = r_9[25] /*37441*/;
  assign m_10[4] = r_9[26] /*37440*/;
  assign m_10[5] = r_9[27] /*37439*/;
  assign m_10[6] = r_9[28] /*37438*/;
  assign m_10[7] = r_9[29] /*37437*/;
  assign m_10[8] = r_9[30] /*37436*/;
  assign m_10[9] = r_9[31] /*37435*/;
  assign m_10[10] = r_9[32] /*37434*/;
  assign m_10[11] = r_9[33] /*37433*/;
  assign m_10[12] = r_9[34] /*37432*/;
  assign m_10[13] = r_9[35] /*37431*/;
  assign m_10[14] = r_9[36] /*37430*/;
  assign m_10[15] = r_9[37] /*37429*/;
  assign m_10[16] = r_9[38] /*37428*/;
  assign m_10[17] = r_9[39] /*37427*/;
  assign m_10[18] = r_9[40] /*37426*/;
  assign m_10[19] = r_9[41] /*37425*/;
  assign m_10[20] = r_9[42] /*37424*/;
  assign m_10[21] = r_9[43] /*37423*/;
  assign m_10[22] = r_9[44] /*37422*/;
  assign m_10[23] = r_9[45] /*37421*/;
  assign m_10[24] = r_9[46] /*37420*/;
  assign m_10[25] = r_9[47] /*37419*/;
  assign m_10[26] = r_9[48] /*37418*/;
  assign m_10[27] = r_9[49] /*37417*/;
  assign m_10[28] = r_9[50] /*37416*/;
  assign m_10[29] = r_9[51] /*37415*/;
  assign m_10[30] = r_9[52] /*37414*/;
  assign m_10[31] = r_9[53] /*37413*/;
  assign _2144_ = ~q[22] /*37411*/;
  assign _2145_ = sum_10[0] & q[22] /*37410*/;
  assign _2146_ = m_10[0] & _2144_ /*37409*/;
  assign r_10[22] = _2146_ | _2145_ /*37408*/;
  assign _2147_ = ~q[22] /*37407*/;
  assign _2148_ = sum_10[1] & q[22] /*37406*/;
  assign _2149_ = m_10[1] & _2147_ /*37405*/;
  assign r_10[23] = _2149_ | _2148_ /*37404*/;
  assign _2150_ = ~q[22] /*37403*/;
  assign _2151_ = sum_10[2] & q[22] /*37402*/;
  assign _2152_ = m_10[2] & _2150_ /*37401*/;
  assign r_10[24] = _2152_ | _2151_ /*37400*/;
  assign _2153_ = ~q[22] /*37399*/;
  assign _2154_ = sum_10[3] & q[22] /*37398*/;
  assign _2155_ = m_10[3] & _2153_ /*37397*/;
  assign r_10[25] = _2155_ | _2154_ /*37396*/;
  assign _2156_ = ~q[22] /*37395*/;
  assign _2157_ = sum_10[4] & q[22] /*37394*/;
  assign _2158_ = m_10[4] & _2156_ /*37393*/;
  assign r_10[26] = _2158_ | _2157_ /*37392*/;
  assign _2159_ = ~q[22] /*37391*/;
  assign _2160_ = sum_10[5] & q[22] /*37390*/;
  assign _2161_ = m_10[5] & _2159_ /*37389*/;
  assign r_10[27] = _2161_ | _2160_ /*37388*/;
  assign _2162_ = ~q[22] /*37387*/;
  assign _2163_ = sum_10[6] & q[22] /*37386*/;
  assign _2164_ = m_10[6] & _2162_ /*37385*/;
  assign r_10[28] = _2164_ | _2163_ /*37384*/;
  assign _2165_ = ~q[22] /*37383*/;
  assign _2166_ = sum_10[7] & q[22] /*37382*/;
  assign _2167_ = m_10[7] & _2165_ /*37381*/;
  assign r_10[29] = _2167_ | _2166_ /*37380*/;
  assign _2168_ = ~q[22] /*37379*/;
  assign _2169_ = sum_10[8] & q[22] /*37378*/;
  assign _2170_ = m_10[8] & _2168_ /*37377*/;
  assign r_10[30] = _2170_ | _2169_ /*37376*/;
  assign _2171_ = ~q[22] /*37375*/;
  assign _2172_ = sum_10[9] & q[22] /*37374*/;
  assign _2173_ = m_10[9] & _2171_ /*37373*/;
  assign r_10[31] = _2173_ | _2172_ /*37372*/;
  assign _2174_ = ~q[22] /*37371*/;
  assign _2175_ = sum_10[10] & q[22] /*37370*/;
  assign _2176_ = m_10[10] & _2174_ /*37369*/;
  assign r_10[32] = _2176_ | _2175_ /*37368*/;
  assign _2177_ = ~q[22] /*37367*/;
  assign _2178_ = sum_10[11] & q[22] /*37366*/;
  assign _2179_ = m_10[11] & _2177_ /*37365*/;
  assign r_10[33] = _2179_ | _2178_ /*37364*/;
  assign _2180_ = ~q[22] /*37363*/;
  assign _2181_ = sum_10[12] & q[22] /*37362*/;
  assign _2182_ = m_10[12] & _2180_ /*37361*/;
  assign r_10[34] = _2182_ | _2181_ /*37360*/;
  assign _2183_ = ~q[22] /*37359*/;
  assign _2184_ = sum_10[13] & q[22] /*37358*/;
  assign _2185_ = m_10[13] & _2183_ /*37357*/;
  assign r_10[35] = _2185_ | _2184_ /*37356*/;
  assign _2186_ = ~q[22] /*37355*/;
  assign _2187_ = sum_10[14] & q[22] /*37354*/;
  assign _2188_ = m_10[14] & _2186_ /*37353*/;
  assign r_10[36] = _2188_ | _2187_ /*37352*/;
  assign _2189_ = ~q[22] /*37351*/;
  assign _2190_ = sum_10[15] & q[22] /*37350*/;
  assign _2191_ = m_10[15] & _2189_ /*37349*/;
  assign r_10[37] = _2191_ | _2190_ /*37348*/;
  assign _2192_ = ~q[22] /*37347*/;
  assign _2193_ = sum_10[16] & q[22] /*37346*/;
  assign _2194_ = m_10[16] & _2192_ /*37345*/;
  assign r_10[38] = _2194_ | _2193_ /*37344*/;
  assign _2195_ = ~q[22] /*37343*/;
  assign _2196_ = sum_10[17] & q[22] /*37342*/;
  assign _2197_ = m_10[17] & _2195_ /*37341*/;
  assign r_10[39] = _2197_ | _2196_ /*37340*/;
  assign _2198_ = ~q[22] /*37339*/;
  assign _2199_ = sum_10[18] & q[22] /*37338*/;
  assign _2200_ = m_10[18] & _2198_ /*37337*/;
  assign r_10[40] = _2200_ | _2199_ /*37336*/;
  assign _2201_ = ~q[22] /*37335*/;
  assign _2202_ = sum_10[19] & q[22] /*37334*/;
  assign _2203_ = m_10[19] & _2201_ /*37333*/;
  assign r_10[41] = _2203_ | _2202_ /*37332*/;
  assign _2204_ = ~q[22] /*37331*/;
  assign _2205_ = sum_10[20] & q[22] /*37330*/;
  assign _2206_ = m_10[20] & _2204_ /*37329*/;
  assign r_10[42] = _2206_ | _2205_ /*37328*/;
  assign _2207_ = ~q[22] /*37327*/;
  assign _2208_ = sum_10[21] & q[22] /*37326*/;
  assign _2209_ = m_10[21] & _2207_ /*37325*/;
  assign r_10[43] = _2209_ | _2208_ /*37324*/;
  assign _2210_ = ~q[22] /*37323*/;
  assign _2211_ = sum_10[22] & q[22] /*37322*/;
  assign _2212_ = m_10[22] & _2210_ /*37321*/;
  assign r_10[44] = _2212_ | _2211_ /*37320*/;
  assign _2213_ = ~q[22] /*37319*/;
  assign _2214_ = sum_10[23] & q[22] /*37318*/;
  assign _2215_ = m_10[23] & _2213_ /*37317*/;
  assign r_10[45] = _2215_ | _2214_ /*37316*/;
  assign _2216_ = ~q[22] /*37315*/;
  assign _2217_ = sum_10[24] & q[22] /*37314*/;
  assign _2218_ = m_10[24] & _2216_ /*37313*/;
  assign r_10[46] = _2218_ | _2217_ /*37312*/;
  assign _2219_ = ~q[22] /*37311*/;
  assign _2220_ = sum_10[25] & q[22] /*37310*/;
  assign _2221_ = m_10[25] & _2219_ /*37309*/;
  assign r_10[47] = _2221_ | _2220_ /*37308*/;
  assign _2222_ = ~q[22] /*37307*/;
  assign _2223_ = sum_10[26] & q[22] /*37306*/;
  assign _2224_ = m_10[26] & _2222_ /*37305*/;
  assign r_10[48] = _2224_ | _2223_ /*37304*/;
  assign _2225_ = ~q[22] /*37303*/;
  assign _2226_ = sum_10[27] & q[22] /*37302*/;
  assign _2227_ = m_10[27] & _2225_ /*37301*/;
  assign r_10[49] = _2227_ | _2226_ /*37300*/;
  assign _2228_ = ~q[22] /*37299*/;
  assign _2229_ = sum_10[28] & q[22] /*37298*/;
  assign _2230_ = m_10[28] & _2228_ /*37297*/;
  assign r_10[50] = _2230_ | _2229_ /*37296*/;
  assign _2231_ = ~q[22] /*37295*/;
  assign _2232_ = sum_10[29] & q[22] /*37294*/;
  assign _2233_ = m_10[29] & _2231_ /*37293*/;
  assign r_10[51] = _2233_ | _2232_ /*37292*/;
  assign _2234_ = ~q[22] /*37291*/;
  assign _2235_ = sum_10[30] & q[22] /*37290*/;
  assign _2236_ = m_10[30] & _2234_ /*37289*/;
  assign r_10[52] = _2236_ | _2235_ /*37288*/;
  assign _2237_ = ~q[22] /*37287*/;
  assign _2238_ = sum_10[31] & q[22] /*37286*/;
  assign _2239_ = m_10[31] & _2237_ /*37285*/;
  assign r_10[53] = _2239_ | _2238_ /*37284*/;
assign r_10[0]= r_9[0] /*37283*/;
assign r_10[1]= r_9[1] /*37282*/;
assign r_10[2]= r_9[2] /*37281*/;
assign r_10[3]= r_9[3] /*37280*/;
assign r_10[4]= r_9[4] /*37279*/;
assign r_10[5]= r_9[5] /*37278*/;
assign r_10[6]= r_9[6] /*37277*/;
assign r_10[7]= r_9[7] /*37276*/;
assign r_10[8]= r_9[8] /*37275*/;
assign r_10[9]= r_9[9] /*37274*/;
assign r_10[10]= r_9[10] /*37273*/;
assign r_10[11]= r_9[11] /*37272*/;
assign r_10[12]= r_9[12] /*37271*/;
assign r_10[13]= r_9[13] /*37270*/;
assign r_10[14]= r_9[14] /*37269*/;
assign r_10[15]= r_9[15] /*37268*/;
assign r_10[16]= r_9[16] /*37267*/;
assign r_10[17]= r_9[17] /*37266*/;
assign r_10[18]= r_9[18] /*37265*/;
assign r_10[19]= r_9[19] /*37264*/;
assign r_10[20]= r_9[20] /*37263*/;
assign r_10[21]= r_9[21] /*37262*/;
  assign inv_11[0] = ~div[0] /*37192*/;
  assign inv_11[1] = ~div[1] /*37191*/;
  assign inv_11[2] = ~div[2] /*37190*/;
  assign inv_11[3] = ~div[3] /*37189*/;
  assign inv_11[4] = ~div[4] /*37188*/;
  assign inv_11[5] = ~div[5] /*37187*/;
  assign inv_11[6] = ~div[6] /*37186*/;
  assign inv_11[7] = ~div[7] /*37185*/;
  assign inv_11[8] = ~div[8] /*37184*/;
  assign inv_11[9] = ~div[9] /*37183*/;
  assign inv_11[10] = ~div[10] /*37182*/;
  assign inv_11[11] = ~div[11] /*37181*/;
  assign inv_11[12] = ~div[12] /*37180*/;
  assign inv_11[13] = ~div[13] /*37179*/;
  assign inv_11[14] = ~div[14] /*37178*/;
  assign inv_11[15] = ~div[15] /*37177*/;
  assign inv_11[16] = ~div[16] /*37176*/;
  assign inv_11[17] = ~div[17] /*37175*/;
  assign inv_11[18] = ~div[18] /*37174*/;
  assign inv_11[19] = ~div[19] /*37173*/;
  assign inv_11[20] = ~div[20] /*37172*/;
  assign inv_11[21] = ~div[21] /*37171*/;
  assign inv_11[22] = ~div[22] /*37170*/;
  assign inv_11[23] = ~div[23] /*37169*/;
  assign inv_11[24] = ~div[24] /*37168*/;
  assign inv_11[25] = ~div[25] /*37167*/;
  assign inv_11[26] = ~div[26] /*37166*/;
  assign inv_11[27] = ~div[27] /*37165*/;
  assign inv_11[28] = ~div[28] /*37164*/;
  assign inv_11[29] = ~div[29] /*37163*/;
  assign inv_11[30] = ~div[30] /*37162*/;
assign inv_11[31] = oneWire /*37161*/;
  assign _2240_ = inv_11[0] ^ r_10[21] /*37159*/;
  assign sum_11[0] = _2240_ ^ oneWire /*37158*/;
  assign _2241_ = _2240_ & oneWire /*37157*/;
  assign _2242_ = inv_11[0] & r_10[21] /*37156*/;
  assign _2243_ = _2241_ | _2242_ /*37155*/;
  assign _2244_ = inv_11[1] ^ r_10[22] /*37154*/;
  assign sum_11[1] = _2244_ ^ _2243_ /*37153*/;
  assign _2245_ = _2244_ & _2243_ /*37152*/;
  assign _2246_ = inv_11[1] & r_10[22] /*37151*/;
  assign _2247_ = _2245_ | _2246_ /*37150*/;
  assign _2248_ = inv_11[2] ^ r_10[23] /*37148*/;
  assign sum_11[2] = _2248_ ^ _2247_ /*37147*/;
  assign _2249_ = _2248_ & _2247_ /*37146*/;
  assign _2250_ = inv_11[2] & r_10[23] /*37145*/;
  assign _2251_ = _2249_ | _2250_ /*37144*/;
  assign _2252_ = inv_11[3] ^ r_10[24] /*37142*/;
  assign sum_11[3] = _2252_ ^ _2251_ /*37141*/;
  assign _2253_ = _2252_ & _2251_ /*37140*/;
  assign _2254_ = inv_11[3] & r_10[24] /*37139*/;
  assign _2255_ = _2253_ | _2254_ /*37138*/;
  assign _2256_ = inv_11[4] ^ r_10[25] /*37136*/;
  assign sum_11[4] = _2256_ ^ _2255_ /*37135*/;
  assign _2257_ = _2256_ & _2255_ /*37134*/;
  assign _2258_ = inv_11[4] & r_10[25] /*37133*/;
  assign _2259_ = _2257_ | _2258_ /*37132*/;
  assign _2260_ = inv_11[5] ^ r_10[26] /*37130*/;
  assign sum_11[5] = _2260_ ^ _2259_ /*37129*/;
  assign _2261_ = _2260_ & _2259_ /*37128*/;
  assign _2262_ = inv_11[5] & r_10[26] /*37127*/;
  assign _2263_ = _2261_ | _2262_ /*37126*/;
  assign _2264_ = inv_11[6] ^ r_10[27] /*37124*/;
  assign sum_11[6] = _2264_ ^ _2263_ /*37123*/;
  assign _2265_ = _2264_ & _2263_ /*37122*/;
  assign _2266_ = inv_11[6] & r_10[27] /*37121*/;
  assign _2267_ = _2265_ | _2266_ /*37120*/;
  assign _2268_ = inv_11[7] ^ r_10[28] /*37118*/;
  assign sum_11[7] = _2268_ ^ _2267_ /*37117*/;
  assign _2269_ = _2268_ & _2267_ /*37116*/;
  assign _2270_ = inv_11[7] & r_10[28] /*37115*/;
  assign _2271_ = _2269_ | _2270_ /*37114*/;
  assign _2272_ = inv_11[8] ^ r_10[29] /*37112*/;
  assign sum_11[8] = _2272_ ^ _2271_ /*37111*/;
  assign _2273_ = _2272_ & _2271_ /*37110*/;
  assign _2274_ = inv_11[8] & r_10[29] /*37109*/;
  assign _2275_ = _2273_ | _2274_ /*37108*/;
  assign _2276_ = inv_11[9] ^ r_10[30] /*37106*/;
  assign sum_11[9] = _2276_ ^ _2275_ /*37105*/;
  assign _2277_ = _2276_ & _2275_ /*37104*/;
  assign _2278_ = inv_11[9] & r_10[30] /*37103*/;
  assign _2279_ = _2277_ | _2278_ /*37102*/;
  assign _2280_ = inv_11[10] ^ r_10[31] /*37100*/;
  assign sum_11[10] = _2280_ ^ _2279_ /*37099*/;
  assign _2281_ = _2280_ & _2279_ /*37098*/;
  assign _2282_ = inv_11[10] & r_10[31] /*37097*/;
  assign _2283_ = _2281_ | _2282_ /*37096*/;
  assign _2284_ = inv_11[11] ^ r_10[32] /*37094*/;
  assign sum_11[11] = _2284_ ^ _2283_ /*37093*/;
  assign _2285_ = _2284_ & _2283_ /*37092*/;
  assign _2286_ = inv_11[11] & r_10[32] /*37091*/;
  assign _2287_ = _2285_ | _2286_ /*37090*/;
  assign _2288_ = inv_11[12] ^ r_10[33] /*37088*/;
  assign sum_11[12] = _2288_ ^ _2287_ /*37087*/;
  assign _2289_ = _2288_ & _2287_ /*37086*/;
  assign _2290_ = inv_11[12] & r_10[33] /*37085*/;
  assign _2291_ = _2289_ | _2290_ /*37084*/;
  assign _2292_ = inv_11[13] ^ r_10[34] /*37082*/;
  assign sum_11[13] = _2292_ ^ _2291_ /*37081*/;
  assign _2293_ = _2292_ & _2291_ /*37080*/;
  assign _2294_ = inv_11[13] & r_10[34] /*37079*/;
  assign _2295_ = _2293_ | _2294_ /*37078*/;
  assign _2296_ = inv_11[14] ^ r_10[35] /*37076*/;
  assign sum_11[14] = _2296_ ^ _2295_ /*37075*/;
  assign _2297_ = _2296_ & _2295_ /*37074*/;
  assign _2298_ = inv_11[14] & r_10[35] /*37073*/;
  assign _2299_ = _2297_ | _2298_ /*37072*/;
  assign _2300_ = inv_11[15] ^ r_10[36] /*37070*/;
  assign sum_11[15] = _2300_ ^ _2299_ /*37069*/;
  assign _2301_ = _2300_ & _2299_ /*37068*/;
  assign _2302_ = inv_11[15] & r_10[36] /*37067*/;
  assign _2303_ = _2301_ | _2302_ /*37066*/;
  assign _2304_ = inv_11[16] ^ r_10[37] /*37064*/;
  assign sum_11[16] = _2304_ ^ _2303_ /*37063*/;
  assign _2305_ = _2304_ & _2303_ /*37062*/;
  assign _2306_ = inv_11[16] & r_10[37] /*37061*/;
  assign _2307_ = _2305_ | _2306_ /*37060*/;
  assign _2308_ = inv_11[17] ^ r_10[38] /*37058*/;
  assign sum_11[17] = _2308_ ^ _2307_ /*37057*/;
  assign _2309_ = _2308_ & _2307_ /*37056*/;
  assign _2310_ = inv_11[17] & r_10[38] /*37055*/;
  assign _2311_ = _2309_ | _2310_ /*37054*/;
  assign _2312_ = inv_11[18] ^ r_10[39] /*37052*/;
  assign sum_11[18] = _2312_ ^ _2311_ /*37051*/;
  assign _2313_ = _2312_ & _2311_ /*37050*/;
  assign _2314_ = inv_11[18] & r_10[39] /*37049*/;
  assign _2315_ = _2313_ | _2314_ /*37048*/;
  assign _2316_ = inv_11[19] ^ r_10[40] /*37046*/;
  assign sum_11[19] = _2316_ ^ _2315_ /*37045*/;
  assign _2317_ = _2316_ & _2315_ /*37044*/;
  assign _2318_ = inv_11[19] & r_10[40] /*37043*/;
  assign _2319_ = _2317_ | _2318_ /*37042*/;
  assign _2320_ = inv_11[20] ^ r_10[41] /*37040*/;
  assign sum_11[20] = _2320_ ^ _2319_ /*37039*/;
  assign _2321_ = _2320_ & _2319_ /*37038*/;
  assign _2322_ = inv_11[20] & r_10[41] /*37037*/;
  assign _2323_ = _2321_ | _2322_ /*37036*/;
  assign _2324_ = inv_11[21] ^ r_10[42] /*37034*/;
  assign sum_11[21] = _2324_ ^ _2323_ /*37033*/;
  assign _2325_ = _2324_ & _2323_ /*37032*/;
  assign _2326_ = inv_11[21] & r_10[42] /*37031*/;
  assign _2327_ = _2325_ | _2326_ /*37030*/;
  assign _2328_ = inv_11[22] ^ r_10[43] /*37028*/;
  assign sum_11[22] = _2328_ ^ _2327_ /*37027*/;
  assign _2329_ = _2328_ & _2327_ /*37026*/;
  assign _2330_ = inv_11[22] & r_10[43] /*37025*/;
  assign _2331_ = _2329_ | _2330_ /*37024*/;
  assign _2332_ = inv_11[23] ^ r_10[44] /*37022*/;
  assign sum_11[23] = _2332_ ^ _2331_ /*37021*/;
  assign _2333_ = _2332_ & _2331_ /*37020*/;
  assign _2334_ = inv_11[23] & r_10[44] /*37019*/;
  assign _2335_ = _2333_ | _2334_ /*37018*/;
  assign _2336_ = inv_11[24] ^ r_10[45] /*37016*/;
  assign sum_11[24] = _2336_ ^ _2335_ /*37015*/;
  assign _2337_ = _2336_ & _2335_ /*37014*/;
  assign _2338_ = inv_11[24] & r_10[45] /*37013*/;
  assign _2339_ = _2337_ | _2338_ /*37012*/;
  assign _2340_ = inv_11[25] ^ r_10[46] /*37010*/;
  assign sum_11[25] = _2340_ ^ _2339_ /*37009*/;
  assign _2341_ = _2340_ & _2339_ /*37008*/;
  assign _2342_ = inv_11[25] & r_10[46] /*37007*/;
  assign _2343_ = _2341_ | _2342_ /*37006*/;
  assign _2344_ = inv_11[26] ^ r_10[47] /*37004*/;
  assign sum_11[26] = _2344_ ^ _2343_ /*37003*/;
  assign _2345_ = _2344_ & _2343_ /*37002*/;
  assign _2346_ = inv_11[26] & r_10[47] /*37001*/;
  assign _2347_ = _2345_ | _2346_ /*37000*/;
  assign _2348_ = inv_11[27] ^ r_10[48] /*36998*/;
  assign sum_11[27] = _2348_ ^ _2347_ /*36997*/;
  assign _2349_ = _2348_ & _2347_ /*36996*/;
  assign _2350_ = inv_11[27] & r_10[48] /*36995*/;
  assign _2351_ = _2349_ | _2350_ /*36994*/;
  assign _2352_ = inv_11[28] ^ r_10[49] /*36992*/;
  assign sum_11[28] = _2352_ ^ _2351_ /*36991*/;
  assign _2353_ = _2352_ & _2351_ /*36990*/;
  assign _2354_ = inv_11[28] & r_10[49] /*36989*/;
  assign _2355_ = _2353_ | _2354_ /*36988*/;
  assign _2356_ = inv_11[29] ^ r_10[50] /*36986*/;
  assign sum_11[29] = _2356_ ^ _2355_ /*36985*/;
  assign _2357_ = _2356_ & _2355_ /*36984*/;
  assign _2358_ = inv_11[29] & r_10[50] /*36983*/;
  assign _2359_ = _2357_ | _2358_ /*36982*/;
  assign _2360_ = inv_11[30] ^ r_10[51] /*36980*/;
  assign sum_11[30] = _2360_ ^ _2359_ /*36979*/;
  assign _2361_ = _2360_ & _2359_ /*36978*/;
  assign _2362_ = inv_11[30] & r_10[51] /*36977*/;
  assign _2363_ = _2361_ | _2362_ /*36976*/;
  assign _2364_ = inv_11[31] ^ r_10[52] /*36974*/;
  assign sum_11[31] = _2364_ ^ _2363_ /*36973*/;
  assign _2365_ = _2364_ & _2363_ /*36972*/;
  assign _2366_ = inv_11[31] & r_10[52] /*36971*/;
  assign _2367_ = _2365_ | _2366_ /*36970*/;
  assign q[21] = ~sum_11[31] /*36997*/;
  assign m_11[0] = r_10[21] /*36996*/;
  assign m_11[1] = r_10[22] /*36995*/;
  assign m_11[2] = r_10[23] /*36994*/;
  assign m_11[3] = r_10[24] /*36993*/;
  assign m_11[4] = r_10[25] /*36992*/;
  assign m_11[5] = r_10[26] /*36991*/;
  assign m_11[6] = r_10[27] /*36990*/;
  assign m_11[7] = r_10[28] /*36989*/;
  assign m_11[8] = r_10[29] /*36988*/;
  assign m_11[9] = r_10[30] /*36987*/;
  assign m_11[10] = r_10[31] /*36986*/;
  assign m_11[11] = r_10[32] /*36985*/;
  assign m_11[12] = r_10[33] /*36984*/;
  assign m_11[13] = r_10[34] /*36983*/;
  assign m_11[14] = r_10[35] /*36982*/;
  assign m_11[15] = r_10[36] /*36981*/;
  assign m_11[16] = r_10[37] /*36980*/;
  assign m_11[17] = r_10[38] /*36979*/;
  assign m_11[18] = r_10[39] /*36978*/;
  assign m_11[19] = r_10[40] /*36977*/;
  assign m_11[20] = r_10[41] /*36976*/;
  assign m_11[21] = r_10[42] /*36975*/;
  assign m_11[22] = r_10[43] /*36974*/;
  assign m_11[23] = r_10[44] /*36973*/;
  assign m_11[24] = r_10[45] /*36972*/;
  assign m_11[25] = r_10[46] /*36971*/;
  assign m_11[26] = r_10[47] /*36970*/;
  assign m_11[27] = r_10[48] /*36969*/;
  assign m_11[28] = r_10[49] /*36968*/;
  assign m_11[29] = r_10[50] /*36967*/;
  assign m_11[30] = r_10[51] /*36966*/;
  assign m_11[31] = r_10[52] /*36965*/;
  assign _2368_ = ~q[21] /*36963*/;
  assign _2369_ = sum_11[0] & q[21] /*36962*/;
  assign _2370_ = m_11[0] & _2368_ /*36961*/;
  assign r_11[21] = _2370_ | _2369_ /*36960*/;
  assign _2371_ = ~q[21] /*36959*/;
  assign _2372_ = sum_11[1] & q[21] /*36958*/;
  assign _2373_ = m_11[1] & _2371_ /*36957*/;
  assign r_11[22] = _2373_ | _2372_ /*36956*/;
  assign _2374_ = ~q[21] /*36955*/;
  assign _2375_ = sum_11[2] & q[21] /*36954*/;
  assign _2376_ = m_11[2] & _2374_ /*36953*/;
  assign r_11[23] = _2376_ | _2375_ /*36952*/;
  assign _2377_ = ~q[21] /*36951*/;
  assign _2378_ = sum_11[3] & q[21] /*36950*/;
  assign _2379_ = m_11[3] & _2377_ /*36949*/;
  assign r_11[24] = _2379_ | _2378_ /*36948*/;
  assign _2380_ = ~q[21] /*36947*/;
  assign _2381_ = sum_11[4] & q[21] /*36946*/;
  assign _2382_ = m_11[4] & _2380_ /*36945*/;
  assign r_11[25] = _2382_ | _2381_ /*36944*/;
  assign _2383_ = ~q[21] /*36943*/;
  assign _2384_ = sum_11[5] & q[21] /*36942*/;
  assign _2385_ = m_11[5] & _2383_ /*36941*/;
  assign r_11[26] = _2385_ | _2384_ /*36940*/;
  assign _2386_ = ~q[21] /*36939*/;
  assign _2387_ = sum_11[6] & q[21] /*36938*/;
  assign _2388_ = m_11[6] & _2386_ /*36937*/;
  assign r_11[27] = _2388_ | _2387_ /*36936*/;
  assign _2389_ = ~q[21] /*36935*/;
  assign _2390_ = sum_11[7] & q[21] /*36934*/;
  assign _2391_ = m_11[7] & _2389_ /*36933*/;
  assign r_11[28] = _2391_ | _2390_ /*36932*/;
  assign _2392_ = ~q[21] /*36931*/;
  assign _2393_ = sum_11[8] & q[21] /*36930*/;
  assign _2394_ = m_11[8] & _2392_ /*36929*/;
  assign r_11[29] = _2394_ | _2393_ /*36928*/;
  assign _2395_ = ~q[21] /*36927*/;
  assign _2396_ = sum_11[9] & q[21] /*36926*/;
  assign _2397_ = m_11[9] & _2395_ /*36925*/;
  assign r_11[30] = _2397_ | _2396_ /*36924*/;
  assign _2398_ = ~q[21] /*36923*/;
  assign _2399_ = sum_11[10] & q[21] /*36922*/;
  assign _2400_ = m_11[10] & _2398_ /*36921*/;
  assign r_11[31] = _2400_ | _2399_ /*36920*/;
  assign _2401_ = ~q[21] /*36919*/;
  assign _2402_ = sum_11[11] & q[21] /*36918*/;
  assign _2403_ = m_11[11] & _2401_ /*36917*/;
  assign r_11[32] = _2403_ | _2402_ /*36916*/;
  assign _2404_ = ~q[21] /*36915*/;
  assign _2405_ = sum_11[12] & q[21] /*36914*/;
  assign _2406_ = m_11[12] & _2404_ /*36913*/;
  assign r_11[33] = _2406_ | _2405_ /*36912*/;
  assign _2407_ = ~q[21] /*36911*/;
  assign _2408_ = sum_11[13] & q[21] /*36910*/;
  assign _2409_ = m_11[13] & _2407_ /*36909*/;
  assign r_11[34] = _2409_ | _2408_ /*36908*/;
  assign _2410_ = ~q[21] /*36907*/;
  assign _2411_ = sum_11[14] & q[21] /*36906*/;
  assign _2412_ = m_11[14] & _2410_ /*36905*/;
  assign r_11[35] = _2412_ | _2411_ /*36904*/;
  assign _2413_ = ~q[21] /*36903*/;
  assign _2414_ = sum_11[15] & q[21] /*36902*/;
  assign _2415_ = m_11[15] & _2413_ /*36901*/;
  assign r_11[36] = _2415_ | _2414_ /*36900*/;
  assign _2416_ = ~q[21] /*36899*/;
  assign _2417_ = sum_11[16] & q[21] /*36898*/;
  assign _2418_ = m_11[16] & _2416_ /*36897*/;
  assign r_11[37] = _2418_ | _2417_ /*36896*/;
  assign _2419_ = ~q[21] /*36895*/;
  assign _2420_ = sum_11[17] & q[21] /*36894*/;
  assign _2421_ = m_11[17] & _2419_ /*36893*/;
  assign r_11[38] = _2421_ | _2420_ /*36892*/;
  assign _2422_ = ~q[21] /*36891*/;
  assign _2423_ = sum_11[18] & q[21] /*36890*/;
  assign _2424_ = m_11[18] & _2422_ /*36889*/;
  assign r_11[39] = _2424_ | _2423_ /*36888*/;
  assign _2425_ = ~q[21] /*36887*/;
  assign _2426_ = sum_11[19] & q[21] /*36886*/;
  assign _2427_ = m_11[19] & _2425_ /*36885*/;
  assign r_11[40] = _2427_ | _2426_ /*36884*/;
  assign _2428_ = ~q[21] /*36883*/;
  assign _2429_ = sum_11[20] & q[21] /*36882*/;
  assign _2430_ = m_11[20] & _2428_ /*36881*/;
  assign r_11[41] = _2430_ | _2429_ /*36880*/;
  assign _2431_ = ~q[21] /*36879*/;
  assign _2432_ = sum_11[21] & q[21] /*36878*/;
  assign _2433_ = m_11[21] & _2431_ /*36877*/;
  assign r_11[42] = _2433_ | _2432_ /*36876*/;
  assign _2434_ = ~q[21] /*36875*/;
  assign _2435_ = sum_11[22] & q[21] /*36874*/;
  assign _2436_ = m_11[22] & _2434_ /*36873*/;
  assign r_11[43] = _2436_ | _2435_ /*36872*/;
  assign _2437_ = ~q[21] /*36871*/;
  assign _2438_ = sum_11[23] & q[21] /*36870*/;
  assign _2439_ = m_11[23] & _2437_ /*36869*/;
  assign r_11[44] = _2439_ | _2438_ /*36868*/;
  assign _2440_ = ~q[21] /*36867*/;
  assign _2441_ = sum_11[24] & q[21] /*36866*/;
  assign _2442_ = m_11[24] & _2440_ /*36865*/;
  assign r_11[45] = _2442_ | _2441_ /*36864*/;
  assign _2443_ = ~q[21] /*36863*/;
  assign _2444_ = sum_11[25] & q[21] /*36862*/;
  assign _2445_ = m_11[25] & _2443_ /*36861*/;
  assign r_11[46] = _2445_ | _2444_ /*36860*/;
  assign _2446_ = ~q[21] /*36859*/;
  assign _2447_ = sum_11[26] & q[21] /*36858*/;
  assign _2448_ = m_11[26] & _2446_ /*36857*/;
  assign r_11[47] = _2448_ | _2447_ /*36856*/;
  assign _2449_ = ~q[21] /*36855*/;
  assign _2450_ = sum_11[27] & q[21] /*36854*/;
  assign _2451_ = m_11[27] & _2449_ /*36853*/;
  assign r_11[48] = _2451_ | _2450_ /*36852*/;
  assign _2452_ = ~q[21] /*36851*/;
  assign _2453_ = sum_11[28] & q[21] /*36850*/;
  assign _2454_ = m_11[28] & _2452_ /*36849*/;
  assign r_11[49] = _2454_ | _2453_ /*36848*/;
  assign _2455_ = ~q[21] /*36847*/;
  assign _2456_ = sum_11[29] & q[21] /*36846*/;
  assign _2457_ = m_11[29] & _2455_ /*36845*/;
  assign r_11[50] = _2457_ | _2456_ /*36844*/;
  assign _2458_ = ~q[21] /*36843*/;
  assign _2459_ = sum_11[30] & q[21] /*36842*/;
  assign _2460_ = m_11[30] & _2458_ /*36841*/;
  assign r_11[51] = _2460_ | _2459_ /*36840*/;
  assign _2461_ = ~q[21] /*36839*/;
  assign _2462_ = sum_11[31] & q[21] /*36838*/;
  assign _2463_ = m_11[31] & _2461_ /*36837*/;
  assign r_11[52] = _2463_ | _2462_ /*36836*/;
assign r_11[0]= r_10[0] /*36835*/;
assign r_11[1]= r_10[1] /*36834*/;
assign r_11[2]= r_10[2] /*36833*/;
assign r_11[3]= r_10[3] /*36832*/;
assign r_11[4]= r_10[4] /*36831*/;
assign r_11[5]= r_10[5] /*36830*/;
assign r_11[6]= r_10[6] /*36829*/;
assign r_11[7]= r_10[7] /*36828*/;
assign r_11[8]= r_10[8] /*36827*/;
assign r_11[9]= r_10[9] /*36826*/;
assign r_11[10]= r_10[10] /*36825*/;
assign r_11[11]= r_10[11] /*36824*/;
assign r_11[12]= r_10[12] /*36823*/;
assign r_11[13]= r_10[13] /*36822*/;
assign r_11[14]= r_10[14] /*36821*/;
assign r_11[15]= r_10[15] /*36820*/;
assign r_11[16]= r_10[16] /*36819*/;
assign r_11[17]= r_10[17] /*36818*/;
assign r_11[18]= r_10[18] /*36817*/;
assign r_11[19]= r_10[19] /*36816*/;
assign r_11[20]= r_10[20] /*36815*/;
  assign inv_12[0] = ~div[0] /*36744*/;
  assign inv_12[1] = ~div[1] /*36743*/;
  assign inv_12[2] = ~div[2] /*36742*/;
  assign inv_12[3] = ~div[3] /*36741*/;
  assign inv_12[4] = ~div[4] /*36740*/;
  assign inv_12[5] = ~div[5] /*36739*/;
  assign inv_12[6] = ~div[6] /*36738*/;
  assign inv_12[7] = ~div[7] /*36737*/;
  assign inv_12[8] = ~div[8] /*36736*/;
  assign inv_12[9] = ~div[9] /*36735*/;
  assign inv_12[10] = ~div[10] /*36734*/;
  assign inv_12[11] = ~div[11] /*36733*/;
  assign inv_12[12] = ~div[12] /*36732*/;
  assign inv_12[13] = ~div[13] /*36731*/;
  assign inv_12[14] = ~div[14] /*36730*/;
  assign inv_12[15] = ~div[15] /*36729*/;
  assign inv_12[16] = ~div[16] /*36728*/;
  assign inv_12[17] = ~div[17] /*36727*/;
  assign inv_12[18] = ~div[18] /*36726*/;
  assign inv_12[19] = ~div[19] /*36725*/;
  assign inv_12[20] = ~div[20] /*36724*/;
  assign inv_12[21] = ~div[21] /*36723*/;
  assign inv_12[22] = ~div[22] /*36722*/;
  assign inv_12[23] = ~div[23] /*36721*/;
  assign inv_12[24] = ~div[24] /*36720*/;
  assign inv_12[25] = ~div[25] /*36719*/;
  assign inv_12[26] = ~div[26] /*36718*/;
  assign inv_12[27] = ~div[27] /*36717*/;
  assign inv_12[28] = ~div[28] /*36716*/;
  assign inv_12[29] = ~div[29] /*36715*/;
  assign inv_12[30] = ~div[30] /*36714*/;
assign inv_12[31] = oneWire /*36713*/;
  assign _2464_ = inv_12[0] ^ r_11[20] /*36711*/;
  assign sum_12[0] = _2464_ ^ oneWire /*36710*/;
  assign _2465_ = _2464_ & oneWire /*36709*/;
  assign _2466_ = inv_12[0] & r_11[20] /*36708*/;
  assign _2467_ = _2465_ | _2466_ /*36707*/;
  assign _2468_ = inv_12[1] ^ r_11[21] /*36706*/;
  assign sum_12[1] = _2468_ ^ _2467_ /*36705*/;
  assign _2469_ = _2468_ & _2467_ /*36704*/;
  assign _2470_ = inv_12[1] & r_11[21] /*36703*/;
  assign _2471_ = _2469_ | _2470_ /*36702*/;
  assign _2472_ = inv_12[2] ^ r_11[22] /*36700*/;
  assign sum_12[2] = _2472_ ^ _2471_ /*36699*/;
  assign _2473_ = _2472_ & _2471_ /*36698*/;
  assign _2474_ = inv_12[2] & r_11[22] /*36697*/;
  assign _2475_ = _2473_ | _2474_ /*36696*/;
  assign _2476_ = inv_12[3] ^ r_11[23] /*36694*/;
  assign sum_12[3] = _2476_ ^ _2475_ /*36693*/;
  assign _2477_ = _2476_ & _2475_ /*36692*/;
  assign _2478_ = inv_12[3] & r_11[23] /*36691*/;
  assign _2479_ = _2477_ | _2478_ /*36690*/;
  assign _2480_ = inv_12[4] ^ r_11[24] /*36688*/;
  assign sum_12[4] = _2480_ ^ _2479_ /*36687*/;
  assign _2481_ = _2480_ & _2479_ /*36686*/;
  assign _2482_ = inv_12[4] & r_11[24] /*36685*/;
  assign _2483_ = _2481_ | _2482_ /*36684*/;
  assign _2484_ = inv_12[5] ^ r_11[25] /*36682*/;
  assign sum_12[5] = _2484_ ^ _2483_ /*36681*/;
  assign _2485_ = _2484_ & _2483_ /*36680*/;
  assign _2486_ = inv_12[5] & r_11[25] /*36679*/;
  assign _2487_ = _2485_ | _2486_ /*36678*/;
  assign _2488_ = inv_12[6] ^ r_11[26] /*36676*/;
  assign sum_12[6] = _2488_ ^ _2487_ /*36675*/;
  assign _2489_ = _2488_ & _2487_ /*36674*/;
  assign _2490_ = inv_12[6] & r_11[26] /*36673*/;
  assign _2491_ = _2489_ | _2490_ /*36672*/;
  assign _2492_ = inv_12[7] ^ r_11[27] /*36670*/;
  assign sum_12[7] = _2492_ ^ _2491_ /*36669*/;
  assign _2493_ = _2492_ & _2491_ /*36668*/;
  assign _2494_ = inv_12[7] & r_11[27] /*36667*/;
  assign _2495_ = _2493_ | _2494_ /*36666*/;
  assign _2496_ = inv_12[8] ^ r_11[28] /*36664*/;
  assign sum_12[8] = _2496_ ^ _2495_ /*36663*/;
  assign _2497_ = _2496_ & _2495_ /*36662*/;
  assign _2498_ = inv_12[8] & r_11[28] /*36661*/;
  assign _2499_ = _2497_ | _2498_ /*36660*/;
  assign _2500_ = inv_12[9] ^ r_11[29] /*36658*/;
  assign sum_12[9] = _2500_ ^ _2499_ /*36657*/;
  assign _2501_ = _2500_ & _2499_ /*36656*/;
  assign _2502_ = inv_12[9] & r_11[29] /*36655*/;
  assign _2503_ = _2501_ | _2502_ /*36654*/;
  assign _2504_ = inv_12[10] ^ r_11[30] /*36652*/;
  assign sum_12[10] = _2504_ ^ _2503_ /*36651*/;
  assign _2505_ = _2504_ & _2503_ /*36650*/;
  assign _2506_ = inv_12[10] & r_11[30] /*36649*/;
  assign _2507_ = _2505_ | _2506_ /*36648*/;
  assign _2508_ = inv_12[11] ^ r_11[31] /*36646*/;
  assign sum_12[11] = _2508_ ^ _2507_ /*36645*/;
  assign _2509_ = _2508_ & _2507_ /*36644*/;
  assign _2510_ = inv_12[11] & r_11[31] /*36643*/;
  assign _2511_ = _2509_ | _2510_ /*36642*/;
  assign _2512_ = inv_12[12] ^ r_11[32] /*36640*/;
  assign sum_12[12] = _2512_ ^ _2511_ /*36639*/;
  assign _2513_ = _2512_ & _2511_ /*36638*/;
  assign _2514_ = inv_12[12] & r_11[32] /*36637*/;
  assign _2515_ = _2513_ | _2514_ /*36636*/;
  assign _2516_ = inv_12[13] ^ r_11[33] /*36634*/;
  assign sum_12[13] = _2516_ ^ _2515_ /*36633*/;
  assign _2517_ = _2516_ & _2515_ /*36632*/;
  assign _2518_ = inv_12[13] & r_11[33] /*36631*/;
  assign _2519_ = _2517_ | _2518_ /*36630*/;
  assign _2520_ = inv_12[14] ^ r_11[34] /*36628*/;
  assign sum_12[14] = _2520_ ^ _2519_ /*36627*/;
  assign _2521_ = _2520_ & _2519_ /*36626*/;
  assign _2522_ = inv_12[14] & r_11[34] /*36625*/;
  assign _2523_ = _2521_ | _2522_ /*36624*/;
  assign _2524_ = inv_12[15] ^ r_11[35] /*36622*/;
  assign sum_12[15] = _2524_ ^ _2523_ /*36621*/;
  assign _2525_ = _2524_ & _2523_ /*36620*/;
  assign _2526_ = inv_12[15] & r_11[35] /*36619*/;
  assign _2527_ = _2525_ | _2526_ /*36618*/;
  assign _2528_ = inv_12[16] ^ r_11[36] /*36616*/;
  assign sum_12[16] = _2528_ ^ _2527_ /*36615*/;
  assign _2529_ = _2528_ & _2527_ /*36614*/;
  assign _2530_ = inv_12[16] & r_11[36] /*36613*/;
  assign _2531_ = _2529_ | _2530_ /*36612*/;
  assign _2532_ = inv_12[17] ^ r_11[37] /*36610*/;
  assign sum_12[17] = _2532_ ^ _2531_ /*36609*/;
  assign _2533_ = _2532_ & _2531_ /*36608*/;
  assign _2534_ = inv_12[17] & r_11[37] /*36607*/;
  assign _2535_ = _2533_ | _2534_ /*36606*/;
  assign _2536_ = inv_12[18] ^ r_11[38] /*36604*/;
  assign sum_12[18] = _2536_ ^ _2535_ /*36603*/;
  assign _2537_ = _2536_ & _2535_ /*36602*/;
  assign _2538_ = inv_12[18] & r_11[38] /*36601*/;
  assign _2539_ = _2537_ | _2538_ /*36600*/;
  assign _2540_ = inv_12[19] ^ r_11[39] /*36598*/;
  assign sum_12[19] = _2540_ ^ _2539_ /*36597*/;
  assign _2541_ = _2540_ & _2539_ /*36596*/;
  assign _2542_ = inv_12[19] & r_11[39] /*36595*/;
  assign _2543_ = _2541_ | _2542_ /*36594*/;
  assign _2544_ = inv_12[20] ^ r_11[40] /*36592*/;
  assign sum_12[20] = _2544_ ^ _2543_ /*36591*/;
  assign _2545_ = _2544_ & _2543_ /*36590*/;
  assign _2546_ = inv_12[20] & r_11[40] /*36589*/;
  assign _2547_ = _2545_ | _2546_ /*36588*/;
  assign _2548_ = inv_12[21] ^ r_11[41] /*36586*/;
  assign sum_12[21] = _2548_ ^ _2547_ /*36585*/;
  assign _2549_ = _2548_ & _2547_ /*36584*/;
  assign _2550_ = inv_12[21] & r_11[41] /*36583*/;
  assign _2551_ = _2549_ | _2550_ /*36582*/;
  assign _2552_ = inv_12[22] ^ r_11[42] /*36580*/;
  assign sum_12[22] = _2552_ ^ _2551_ /*36579*/;
  assign _2553_ = _2552_ & _2551_ /*36578*/;
  assign _2554_ = inv_12[22] & r_11[42] /*36577*/;
  assign _2555_ = _2553_ | _2554_ /*36576*/;
  assign _2556_ = inv_12[23] ^ r_11[43] /*36574*/;
  assign sum_12[23] = _2556_ ^ _2555_ /*36573*/;
  assign _2557_ = _2556_ & _2555_ /*36572*/;
  assign _2558_ = inv_12[23] & r_11[43] /*36571*/;
  assign _2559_ = _2557_ | _2558_ /*36570*/;
  assign _2560_ = inv_12[24] ^ r_11[44] /*36568*/;
  assign sum_12[24] = _2560_ ^ _2559_ /*36567*/;
  assign _2561_ = _2560_ & _2559_ /*36566*/;
  assign _2562_ = inv_12[24] & r_11[44] /*36565*/;
  assign _2563_ = _2561_ | _2562_ /*36564*/;
  assign _2564_ = inv_12[25] ^ r_11[45] /*36562*/;
  assign sum_12[25] = _2564_ ^ _2563_ /*36561*/;
  assign _2565_ = _2564_ & _2563_ /*36560*/;
  assign _2566_ = inv_12[25] & r_11[45] /*36559*/;
  assign _2567_ = _2565_ | _2566_ /*36558*/;
  assign _2568_ = inv_12[26] ^ r_11[46] /*36556*/;
  assign sum_12[26] = _2568_ ^ _2567_ /*36555*/;
  assign _2569_ = _2568_ & _2567_ /*36554*/;
  assign _2570_ = inv_12[26] & r_11[46] /*36553*/;
  assign _2571_ = _2569_ | _2570_ /*36552*/;
  assign _2572_ = inv_12[27] ^ r_11[47] /*36550*/;
  assign sum_12[27] = _2572_ ^ _2571_ /*36549*/;
  assign _2573_ = _2572_ & _2571_ /*36548*/;
  assign _2574_ = inv_12[27] & r_11[47] /*36547*/;
  assign _2575_ = _2573_ | _2574_ /*36546*/;
  assign _2576_ = inv_12[28] ^ r_11[48] /*36544*/;
  assign sum_12[28] = _2576_ ^ _2575_ /*36543*/;
  assign _2577_ = _2576_ & _2575_ /*36542*/;
  assign _2578_ = inv_12[28] & r_11[48] /*36541*/;
  assign _2579_ = _2577_ | _2578_ /*36540*/;
  assign _2580_ = inv_12[29] ^ r_11[49] /*36538*/;
  assign sum_12[29] = _2580_ ^ _2579_ /*36537*/;
  assign _2581_ = _2580_ & _2579_ /*36536*/;
  assign _2582_ = inv_12[29] & r_11[49] /*36535*/;
  assign _2583_ = _2581_ | _2582_ /*36534*/;
  assign _2584_ = inv_12[30] ^ r_11[50] /*36532*/;
  assign sum_12[30] = _2584_ ^ _2583_ /*36531*/;
  assign _2585_ = _2584_ & _2583_ /*36530*/;
  assign _2586_ = inv_12[30] & r_11[50] /*36529*/;
  assign _2587_ = _2585_ | _2586_ /*36528*/;
  assign _2588_ = inv_12[31] ^ r_11[51] /*36526*/;
  assign sum_12[31] = _2588_ ^ _2587_ /*36525*/;
  assign _2589_ = _2588_ & _2587_ /*36524*/;
  assign _2590_ = inv_12[31] & r_11[51] /*36523*/;
  assign _2591_ = _2589_ | _2590_ /*36522*/;
  assign q[20] = ~sum_12[31] /*36549*/;
  assign m_12[0] = r_11[20] /*36548*/;
  assign m_12[1] = r_11[21] /*36547*/;
  assign m_12[2] = r_11[22] /*36546*/;
  assign m_12[3] = r_11[23] /*36545*/;
  assign m_12[4] = r_11[24] /*36544*/;
  assign m_12[5] = r_11[25] /*36543*/;
  assign m_12[6] = r_11[26] /*36542*/;
  assign m_12[7] = r_11[27] /*36541*/;
  assign m_12[8] = r_11[28] /*36540*/;
  assign m_12[9] = r_11[29] /*36539*/;
  assign m_12[10] = r_11[30] /*36538*/;
  assign m_12[11] = r_11[31] /*36537*/;
  assign m_12[12] = r_11[32] /*36536*/;
  assign m_12[13] = r_11[33] /*36535*/;
  assign m_12[14] = r_11[34] /*36534*/;
  assign m_12[15] = r_11[35] /*36533*/;
  assign m_12[16] = r_11[36] /*36532*/;
  assign m_12[17] = r_11[37] /*36531*/;
  assign m_12[18] = r_11[38] /*36530*/;
  assign m_12[19] = r_11[39] /*36529*/;
  assign m_12[20] = r_11[40] /*36528*/;
  assign m_12[21] = r_11[41] /*36527*/;
  assign m_12[22] = r_11[42] /*36526*/;
  assign m_12[23] = r_11[43] /*36525*/;
  assign m_12[24] = r_11[44] /*36524*/;
  assign m_12[25] = r_11[45] /*36523*/;
  assign m_12[26] = r_11[46] /*36522*/;
  assign m_12[27] = r_11[47] /*36521*/;
  assign m_12[28] = r_11[48] /*36520*/;
  assign m_12[29] = r_11[49] /*36519*/;
  assign m_12[30] = r_11[50] /*36518*/;
  assign m_12[31] = r_11[51] /*36517*/;
  assign _2592_ = ~q[20] /*36515*/;
  assign _2593_ = sum_12[0] & q[20] /*36514*/;
  assign _2594_ = m_12[0] & _2592_ /*36513*/;
  assign r_12[20] = _2594_ | _2593_ /*36512*/;
  assign _2595_ = ~q[20] /*36511*/;
  assign _2596_ = sum_12[1] & q[20] /*36510*/;
  assign _2597_ = m_12[1] & _2595_ /*36509*/;
  assign r_12[21] = _2597_ | _2596_ /*36508*/;
  assign _2598_ = ~q[20] /*36507*/;
  assign _2599_ = sum_12[2] & q[20] /*36506*/;
  assign _2600_ = m_12[2] & _2598_ /*36505*/;
  assign r_12[22] = _2600_ | _2599_ /*36504*/;
  assign _2601_ = ~q[20] /*36503*/;
  assign _2602_ = sum_12[3] & q[20] /*36502*/;
  assign _2603_ = m_12[3] & _2601_ /*36501*/;
  assign r_12[23] = _2603_ | _2602_ /*36500*/;
  assign _2604_ = ~q[20] /*36499*/;
  assign _2605_ = sum_12[4] & q[20] /*36498*/;
  assign _2606_ = m_12[4] & _2604_ /*36497*/;
  assign r_12[24] = _2606_ | _2605_ /*36496*/;
  assign _2607_ = ~q[20] /*36495*/;
  assign _2608_ = sum_12[5] & q[20] /*36494*/;
  assign _2609_ = m_12[5] & _2607_ /*36493*/;
  assign r_12[25] = _2609_ | _2608_ /*36492*/;
  assign _2610_ = ~q[20] /*36491*/;
  assign _2611_ = sum_12[6] & q[20] /*36490*/;
  assign _2612_ = m_12[6] & _2610_ /*36489*/;
  assign r_12[26] = _2612_ | _2611_ /*36488*/;
  assign _2613_ = ~q[20] /*36487*/;
  assign _2614_ = sum_12[7] & q[20] /*36486*/;
  assign _2615_ = m_12[7] & _2613_ /*36485*/;
  assign r_12[27] = _2615_ | _2614_ /*36484*/;
  assign _2616_ = ~q[20] /*36483*/;
  assign _2617_ = sum_12[8] & q[20] /*36482*/;
  assign _2618_ = m_12[8] & _2616_ /*36481*/;
  assign r_12[28] = _2618_ | _2617_ /*36480*/;
  assign _2619_ = ~q[20] /*36479*/;
  assign _2620_ = sum_12[9] & q[20] /*36478*/;
  assign _2621_ = m_12[9] & _2619_ /*36477*/;
  assign r_12[29] = _2621_ | _2620_ /*36476*/;
  assign _2622_ = ~q[20] /*36475*/;
  assign _2623_ = sum_12[10] & q[20] /*36474*/;
  assign _2624_ = m_12[10] & _2622_ /*36473*/;
  assign r_12[30] = _2624_ | _2623_ /*36472*/;
  assign _2625_ = ~q[20] /*36471*/;
  assign _2626_ = sum_12[11] & q[20] /*36470*/;
  assign _2627_ = m_12[11] & _2625_ /*36469*/;
  assign r_12[31] = _2627_ | _2626_ /*36468*/;
  assign _2628_ = ~q[20] /*36467*/;
  assign _2629_ = sum_12[12] & q[20] /*36466*/;
  assign _2630_ = m_12[12] & _2628_ /*36465*/;
  assign r_12[32] = _2630_ | _2629_ /*36464*/;
  assign _2631_ = ~q[20] /*36463*/;
  assign _2632_ = sum_12[13] & q[20] /*36462*/;
  assign _2633_ = m_12[13] & _2631_ /*36461*/;
  assign r_12[33] = _2633_ | _2632_ /*36460*/;
  assign _2634_ = ~q[20] /*36459*/;
  assign _2635_ = sum_12[14] & q[20] /*36458*/;
  assign _2636_ = m_12[14] & _2634_ /*36457*/;
  assign r_12[34] = _2636_ | _2635_ /*36456*/;
  assign _2637_ = ~q[20] /*36455*/;
  assign _2638_ = sum_12[15] & q[20] /*36454*/;
  assign _2639_ = m_12[15] & _2637_ /*36453*/;
  assign r_12[35] = _2639_ | _2638_ /*36452*/;
  assign _2640_ = ~q[20] /*36451*/;
  assign _2641_ = sum_12[16] & q[20] /*36450*/;
  assign _2642_ = m_12[16] & _2640_ /*36449*/;
  assign r_12[36] = _2642_ | _2641_ /*36448*/;
  assign _2643_ = ~q[20] /*36447*/;
  assign _2644_ = sum_12[17] & q[20] /*36446*/;
  assign _2645_ = m_12[17] & _2643_ /*36445*/;
  assign r_12[37] = _2645_ | _2644_ /*36444*/;
  assign _2646_ = ~q[20] /*36443*/;
  assign _2647_ = sum_12[18] & q[20] /*36442*/;
  assign _2648_ = m_12[18] & _2646_ /*36441*/;
  assign r_12[38] = _2648_ | _2647_ /*36440*/;
  assign _2649_ = ~q[20] /*36439*/;
  assign _2650_ = sum_12[19] & q[20] /*36438*/;
  assign _2651_ = m_12[19] & _2649_ /*36437*/;
  assign r_12[39] = _2651_ | _2650_ /*36436*/;
  assign _2652_ = ~q[20] /*36435*/;
  assign _2653_ = sum_12[20] & q[20] /*36434*/;
  assign _2654_ = m_12[20] & _2652_ /*36433*/;
  assign r_12[40] = _2654_ | _2653_ /*36432*/;
  assign _2655_ = ~q[20] /*36431*/;
  assign _2656_ = sum_12[21] & q[20] /*36430*/;
  assign _2657_ = m_12[21] & _2655_ /*36429*/;
  assign r_12[41] = _2657_ | _2656_ /*36428*/;
  assign _2658_ = ~q[20] /*36427*/;
  assign _2659_ = sum_12[22] & q[20] /*36426*/;
  assign _2660_ = m_12[22] & _2658_ /*36425*/;
  assign r_12[42] = _2660_ | _2659_ /*36424*/;
  assign _2661_ = ~q[20] /*36423*/;
  assign _2662_ = sum_12[23] & q[20] /*36422*/;
  assign _2663_ = m_12[23] & _2661_ /*36421*/;
  assign r_12[43] = _2663_ | _2662_ /*36420*/;
  assign _2664_ = ~q[20] /*36419*/;
  assign _2665_ = sum_12[24] & q[20] /*36418*/;
  assign _2666_ = m_12[24] & _2664_ /*36417*/;
  assign r_12[44] = _2666_ | _2665_ /*36416*/;
  assign _2667_ = ~q[20] /*36415*/;
  assign _2668_ = sum_12[25] & q[20] /*36414*/;
  assign _2669_ = m_12[25] & _2667_ /*36413*/;
  assign r_12[45] = _2669_ | _2668_ /*36412*/;
  assign _2670_ = ~q[20] /*36411*/;
  assign _2671_ = sum_12[26] & q[20] /*36410*/;
  assign _2672_ = m_12[26] & _2670_ /*36409*/;
  assign r_12[46] = _2672_ | _2671_ /*36408*/;
  assign _2673_ = ~q[20] /*36407*/;
  assign _2674_ = sum_12[27] & q[20] /*36406*/;
  assign _2675_ = m_12[27] & _2673_ /*36405*/;
  assign r_12[47] = _2675_ | _2674_ /*36404*/;
  assign _2676_ = ~q[20] /*36403*/;
  assign _2677_ = sum_12[28] & q[20] /*36402*/;
  assign _2678_ = m_12[28] & _2676_ /*36401*/;
  assign r_12[48] = _2678_ | _2677_ /*36400*/;
  assign _2679_ = ~q[20] /*36399*/;
  assign _2680_ = sum_12[29] & q[20] /*36398*/;
  assign _2681_ = m_12[29] & _2679_ /*36397*/;
  assign r_12[49] = _2681_ | _2680_ /*36396*/;
  assign _2682_ = ~q[20] /*36395*/;
  assign _2683_ = sum_12[30] & q[20] /*36394*/;
  assign _2684_ = m_12[30] & _2682_ /*36393*/;
  assign r_12[50] = _2684_ | _2683_ /*36392*/;
  assign _2685_ = ~q[20] /*36391*/;
  assign _2686_ = sum_12[31] & q[20] /*36390*/;
  assign _2687_ = m_12[31] & _2685_ /*36389*/;
  assign r_12[51] = _2687_ | _2686_ /*36388*/;
assign r_12[0]= r_11[0] /*36387*/;
assign r_12[1]= r_11[1] /*36386*/;
assign r_12[2]= r_11[2] /*36385*/;
assign r_12[3]= r_11[3] /*36384*/;
assign r_12[4]= r_11[4] /*36383*/;
assign r_12[5]= r_11[5] /*36382*/;
assign r_12[6]= r_11[6] /*36381*/;
assign r_12[7]= r_11[7] /*36380*/;
assign r_12[8]= r_11[8] /*36379*/;
assign r_12[9]= r_11[9] /*36378*/;
assign r_12[10]= r_11[10] /*36377*/;
assign r_12[11]= r_11[11] /*36376*/;
assign r_12[12]= r_11[12] /*36375*/;
assign r_12[13]= r_11[13] /*36374*/;
assign r_12[14]= r_11[14] /*36373*/;
assign r_12[15]= r_11[15] /*36372*/;
assign r_12[16]= r_11[16] /*36371*/;
assign r_12[17]= r_11[17] /*36370*/;
assign r_12[18]= r_11[18] /*36369*/;
assign r_12[19]= r_11[19] /*36368*/;
  assign inv_13[0] = ~div[0] /*36296*/;
  assign inv_13[1] = ~div[1] /*36295*/;
  assign inv_13[2] = ~div[2] /*36294*/;
  assign inv_13[3] = ~div[3] /*36293*/;
  assign inv_13[4] = ~div[4] /*36292*/;
  assign inv_13[5] = ~div[5] /*36291*/;
  assign inv_13[6] = ~div[6] /*36290*/;
  assign inv_13[7] = ~div[7] /*36289*/;
  assign inv_13[8] = ~div[8] /*36288*/;
  assign inv_13[9] = ~div[9] /*36287*/;
  assign inv_13[10] = ~div[10] /*36286*/;
  assign inv_13[11] = ~div[11] /*36285*/;
  assign inv_13[12] = ~div[12] /*36284*/;
  assign inv_13[13] = ~div[13] /*36283*/;
  assign inv_13[14] = ~div[14] /*36282*/;
  assign inv_13[15] = ~div[15] /*36281*/;
  assign inv_13[16] = ~div[16] /*36280*/;
  assign inv_13[17] = ~div[17] /*36279*/;
  assign inv_13[18] = ~div[18] /*36278*/;
  assign inv_13[19] = ~div[19] /*36277*/;
  assign inv_13[20] = ~div[20] /*36276*/;
  assign inv_13[21] = ~div[21] /*36275*/;
  assign inv_13[22] = ~div[22] /*36274*/;
  assign inv_13[23] = ~div[23] /*36273*/;
  assign inv_13[24] = ~div[24] /*36272*/;
  assign inv_13[25] = ~div[25] /*36271*/;
  assign inv_13[26] = ~div[26] /*36270*/;
  assign inv_13[27] = ~div[27] /*36269*/;
  assign inv_13[28] = ~div[28] /*36268*/;
  assign inv_13[29] = ~div[29] /*36267*/;
  assign inv_13[30] = ~div[30] /*36266*/;
assign inv_13[31] = oneWire /*36265*/;
  assign _2688_ = inv_13[0] ^ r_12[19] /*36263*/;
  assign sum_13[0] = _2688_ ^ oneWire /*36262*/;
  assign _2689_ = _2688_ & oneWire /*36261*/;
  assign _2690_ = inv_13[0] & r_12[19] /*36260*/;
  assign _2691_ = _2689_ | _2690_ /*36259*/;
  assign _2692_ = inv_13[1] ^ r_12[20] /*36258*/;
  assign sum_13[1] = _2692_ ^ _2691_ /*36257*/;
  assign _2693_ = _2692_ & _2691_ /*36256*/;
  assign _2694_ = inv_13[1] & r_12[20] /*36255*/;
  assign _2695_ = _2693_ | _2694_ /*36254*/;
  assign _2696_ = inv_13[2] ^ r_12[21] /*36252*/;
  assign sum_13[2] = _2696_ ^ _2695_ /*36251*/;
  assign _2697_ = _2696_ & _2695_ /*36250*/;
  assign _2698_ = inv_13[2] & r_12[21] /*36249*/;
  assign _2699_ = _2697_ | _2698_ /*36248*/;
  assign _2700_ = inv_13[3] ^ r_12[22] /*36246*/;
  assign sum_13[3] = _2700_ ^ _2699_ /*36245*/;
  assign _2701_ = _2700_ & _2699_ /*36244*/;
  assign _2702_ = inv_13[3] & r_12[22] /*36243*/;
  assign _2703_ = _2701_ | _2702_ /*36242*/;
  assign _2704_ = inv_13[4] ^ r_12[23] /*36240*/;
  assign sum_13[4] = _2704_ ^ _2703_ /*36239*/;
  assign _2705_ = _2704_ & _2703_ /*36238*/;
  assign _2706_ = inv_13[4] & r_12[23] /*36237*/;
  assign _2707_ = _2705_ | _2706_ /*36236*/;
  assign _2708_ = inv_13[5] ^ r_12[24] /*36234*/;
  assign sum_13[5] = _2708_ ^ _2707_ /*36233*/;
  assign _2709_ = _2708_ & _2707_ /*36232*/;
  assign _2710_ = inv_13[5] & r_12[24] /*36231*/;
  assign _2711_ = _2709_ | _2710_ /*36230*/;
  assign _2712_ = inv_13[6] ^ r_12[25] /*36228*/;
  assign sum_13[6] = _2712_ ^ _2711_ /*36227*/;
  assign _2713_ = _2712_ & _2711_ /*36226*/;
  assign _2714_ = inv_13[6] & r_12[25] /*36225*/;
  assign _2715_ = _2713_ | _2714_ /*36224*/;
  assign _2716_ = inv_13[7] ^ r_12[26] /*36222*/;
  assign sum_13[7] = _2716_ ^ _2715_ /*36221*/;
  assign _2717_ = _2716_ & _2715_ /*36220*/;
  assign _2718_ = inv_13[7] & r_12[26] /*36219*/;
  assign _2719_ = _2717_ | _2718_ /*36218*/;
  assign _2720_ = inv_13[8] ^ r_12[27] /*36216*/;
  assign sum_13[8] = _2720_ ^ _2719_ /*36215*/;
  assign _2721_ = _2720_ & _2719_ /*36214*/;
  assign _2722_ = inv_13[8] & r_12[27] /*36213*/;
  assign _2723_ = _2721_ | _2722_ /*36212*/;
  assign _2724_ = inv_13[9] ^ r_12[28] /*36210*/;
  assign sum_13[9] = _2724_ ^ _2723_ /*36209*/;
  assign _2725_ = _2724_ & _2723_ /*36208*/;
  assign _2726_ = inv_13[9] & r_12[28] /*36207*/;
  assign _2727_ = _2725_ | _2726_ /*36206*/;
  assign _2728_ = inv_13[10] ^ r_12[29] /*36204*/;
  assign sum_13[10] = _2728_ ^ _2727_ /*36203*/;
  assign _2729_ = _2728_ & _2727_ /*36202*/;
  assign _2730_ = inv_13[10] & r_12[29] /*36201*/;
  assign _2731_ = _2729_ | _2730_ /*36200*/;
  assign _2732_ = inv_13[11] ^ r_12[30] /*36198*/;
  assign sum_13[11] = _2732_ ^ _2731_ /*36197*/;
  assign _2733_ = _2732_ & _2731_ /*36196*/;
  assign _2734_ = inv_13[11] & r_12[30] /*36195*/;
  assign _2735_ = _2733_ | _2734_ /*36194*/;
  assign _2736_ = inv_13[12] ^ r_12[31] /*36192*/;
  assign sum_13[12] = _2736_ ^ _2735_ /*36191*/;
  assign _2737_ = _2736_ & _2735_ /*36190*/;
  assign _2738_ = inv_13[12] & r_12[31] /*36189*/;
  assign _2739_ = _2737_ | _2738_ /*36188*/;
  assign _2740_ = inv_13[13] ^ r_12[32] /*36186*/;
  assign sum_13[13] = _2740_ ^ _2739_ /*36185*/;
  assign _2741_ = _2740_ & _2739_ /*36184*/;
  assign _2742_ = inv_13[13] & r_12[32] /*36183*/;
  assign _2743_ = _2741_ | _2742_ /*36182*/;
  assign _2744_ = inv_13[14] ^ r_12[33] /*36180*/;
  assign sum_13[14] = _2744_ ^ _2743_ /*36179*/;
  assign _2745_ = _2744_ & _2743_ /*36178*/;
  assign _2746_ = inv_13[14] & r_12[33] /*36177*/;
  assign _2747_ = _2745_ | _2746_ /*36176*/;
  assign _2748_ = inv_13[15] ^ r_12[34] /*36174*/;
  assign sum_13[15] = _2748_ ^ _2747_ /*36173*/;
  assign _2749_ = _2748_ & _2747_ /*36172*/;
  assign _2750_ = inv_13[15] & r_12[34] /*36171*/;
  assign _2751_ = _2749_ | _2750_ /*36170*/;
  assign _2752_ = inv_13[16] ^ r_12[35] /*36168*/;
  assign sum_13[16] = _2752_ ^ _2751_ /*36167*/;
  assign _2753_ = _2752_ & _2751_ /*36166*/;
  assign _2754_ = inv_13[16] & r_12[35] /*36165*/;
  assign _2755_ = _2753_ | _2754_ /*36164*/;
  assign _2756_ = inv_13[17] ^ r_12[36] /*36162*/;
  assign sum_13[17] = _2756_ ^ _2755_ /*36161*/;
  assign _2757_ = _2756_ & _2755_ /*36160*/;
  assign _2758_ = inv_13[17] & r_12[36] /*36159*/;
  assign _2759_ = _2757_ | _2758_ /*36158*/;
  assign _2760_ = inv_13[18] ^ r_12[37] /*36156*/;
  assign sum_13[18] = _2760_ ^ _2759_ /*36155*/;
  assign _2761_ = _2760_ & _2759_ /*36154*/;
  assign _2762_ = inv_13[18] & r_12[37] /*36153*/;
  assign _2763_ = _2761_ | _2762_ /*36152*/;
  assign _2764_ = inv_13[19] ^ r_12[38] /*36150*/;
  assign sum_13[19] = _2764_ ^ _2763_ /*36149*/;
  assign _2765_ = _2764_ & _2763_ /*36148*/;
  assign _2766_ = inv_13[19] & r_12[38] /*36147*/;
  assign _2767_ = _2765_ | _2766_ /*36146*/;
  assign _2768_ = inv_13[20] ^ r_12[39] /*36144*/;
  assign sum_13[20] = _2768_ ^ _2767_ /*36143*/;
  assign _2769_ = _2768_ & _2767_ /*36142*/;
  assign _2770_ = inv_13[20] & r_12[39] /*36141*/;
  assign _2771_ = _2769_ | _2770_ /*36140*/;
  assign _2772_ = inv_13[21] ^ r_12[40] /*36138*/;
  assign sum_13[21] = _2772_ ^ _2771_ /*36137*/;
  assign _2773_ = _2772_ & _2771_ /*36136*/;
  assign _2774_ = inv_13[21] & r_12[40] /*36135*/;
  assign _2775_ = _2773_ | _2774_ /*36134*/;
  assign _2776_ = inv_13[22] ^ r_12[41] /*36132*/;
  assign sum_13[22] = _2776_ ^ _2775_ /*36131*/;
  assign _2777_ = _2776_ & _2775_ /*36130*/;
  assign _2778_ = inv_13[22] & r_12[41] /*36129*/;
  assign _2779_ = _2777_ | _2778_ /*36128*/;
  assign _2780_ = inv_13[23] ^ r_12[42] /*36126*/;
  assign sum_13[23] = _2780_ ^ _2779_ /*36125*/;
  assign _2781_ = _2780_ & _2779_ /*36124*/;
  assign _2782_ = inv_13[23] & r_12[42] /*36123*/;
  assign _2783_ = _2781_ | _2782_ /*36122*/;
  assign _2784_ = inv_13[24] ^ r_12[43] /*36120*/;
  assign sum_13[24] = _2784_ ^ _2783_ /*36119*/;
  assign _2785_ = _2784_ & _2783_ /*36118*/;
  assign _2786_ = inv_13[24] & r_12[43] /*36117*/;
  assign _2787_ = _2785_ | _2786_ /*36116*/;
  assign _2788_ = inv_13[25] ^ r_12[44] /*36114*/;
  assign sum_13[25] = _2788_ ^ _2787_ /*36113*/;
  assign _2789_ = _2788_ & _2787_ /*36112*/;
  assign _2790_ = inv_13[25] & r_12[44] /*36111*/;
  assign _2791_ = _2789_ | _2790_ /*36110*/;
  assign _2792_ = inv_13[26] ^ r_12[45] /*36108*/;
  assign sum_13[26] = _2792_ ^ _2791_ /*36107*/;
  assign _2793_ = _2792_ & _2791_ /*36106*/;
  assign _2794_ = inv_13[26] & r_12[45] /*36105*/;
  assign _2795_ = _2793_ | _2794_ /*36104*/;
  assign _2796_ = inv_13[27] ^ r_12[46] /*36102*/;
  assign sum_13[27] = _2796_ ^ _2795_ /*36101*/;
  assign _2797_ = _2796_ & _2795_ /*36100*/;
  assign _2798_ = inv_13[27] & r_12[46] /*36099*/;
  assign _2799_ = _2797_ | _2798_ /*36098*/;
  assign _2800_ = inv_13[28] ^ r_12[47] /*36096*/;
  assign sum_13[28] = _2800_ ^ _2799_ /*36095*/;
  assign _2801_ = _2800_ & _2799_ /*36094*/;
  assign _2802_ = inv_13[28] & r_12[47] /*36093*/;
  assign _2803_ = _2801_ | _2802_ /*36092*/;
  assign _2804_ = inv_13[29] ^ r_12[48] /*36090*/;
  assign sum_13[29] = _2804_ ^ _2803_ /*36089*/;
  assign _2805_ = _2804_ & _2803_ /*36088*/;
  assign _2806_ = inv_13[29] & r_12[48] /*36087*/;
  assign _2807_ = _2805_ | _2806_ /*36086*/;
  assign _2808_ = inv_13[30] ^ r_12[49] /*36084*/;
  assign sum_13[30] = _2808_ ^ _2807_ /*36083*/;
  assign _2809_ = _2808_ & _2807_ /*36082*/;
  assign _2810_ = inv_13[30] & r_12[49] /*36081*/;
  assign _2811_ = _2809_ | _2810_ /*36080*/;
  assign _2812_ = inv_13[31] ^ r_12[50] /*36078*/;
  assign sum_13[31] = _2812_ ^ _2811_ /*36077*/;
  assign _2813_ = _2812_ & _2811_ /*36076*/;
  assign _2814_ = inv_13[31] & r_12[50] /*36075*/;
  assign _2815_ = _2813_ | _2814_ /*36074*/;
  assign q[19] = ~sum_13[31] /*36101*/;
  assign m_13[0] = r_12[19] /*36100*/;
  assign m_13[1] = r_12[20] /*36099*/;
  assign m_13[2] = r_12[21] /*36098*/;
  assign m_13[3] = r_12[22] /*36097*/;
  assign m_13[4] = r_12[23] /*36096*/;
  assign m_13[5] = r_12[24] /*36095*/;
  assign m_13[6] = r_12[25] /*36094*/;
  assign m_13[7] = r_12[26] /*36093*/;
  assign m_13[8] = r_12[27] /*36092*/;
  assign m_13[9] = r_12[28] /*36091*/;
  assign m_13[10] = r_12[29] /*36090*/;
  assign m_13[11] = r_12[30] /*36089*/;
  assign m_13[12] = r_12[31] /*36088*/;
  assign m_13[13] = r_12[32] /*36087*/;
  assign m_13[14] = r_12[33] /*36086*/;
  assign m_13[15] = r_12[34] /*36085*/;
  assign m_13[16] = r_12[35] /*36084*/;
  assign m_13[17] = r_12[36] /*36083*/;
  assign m_13[18] = r_12[37] /*36082*/;
  assign m_13[19] = r_12[38] /*36081*/;
  assign m_13[20] = r_12[39] /*36080*/;
  assign m_13[21] = r_12[40] /*36079*/;
  assign m_13[22] = r_12[41] /*36078*/;
  assign m_13[23] = r_12[42] /*36077*/;
  assign m_13[24] = r_12[43] /*36076*/;
  assign m_13[25] = r_12[44] /*36075*/;
  assign m_13[26] = r_12[45] /*36074*/;
  assign m_13[27] = r_12[46] /*36073*/;
  assign m_13[28] = r_12[47] /*36072*/;
  assign m_13[29] = r_12[48] /*36071*/;
  assign m_13[30] = r_12[49] /*36070*/;
  assign m_13[31] = r_12[50] /*36069*/;
  assign _2816_ = ~q[19] /*36067*/;
  assign _2817_ = sum_13[0] & q[19] /*36066*/;
  assign _2818_ = m_13[0] & _2816_ /*36065*/;
  assign r_13[19] = _2818_ | _2817_ /*36064*/;
  assign _2819_ = ~q[19] /*36063*/;
  assign _2820_ = sum_13[1] & q[19] /*36062*/;
  assign _2821_ = m_13[1] & _2819_ /*36061*/;
  assign r_13[20] = _2821_ | _2820_ /*36060*/;
  assign _2822_ = ~q[19] /*36059*/;
  assign _2823_ = sum_13[2] & q[19] /*36058*/;
  assign _2824_ = m_13[2] & _2822_ /*36057*/;
  assign r_13[21] = _2824_ | _2823_ /*36056*/;
  assign _2825_ = ~q[19] /*36055*/;
  assign _2826_ = sum_13[3] & q[19] /*36054*/;
  assign _2827_ = m_13[3] & _2825_ /*36053*/;
  assign r_13[22] = _2827_ | _2826_ /*36052*/;
  assign _2828_ = ~q[19] /*36051*/;
  assign _2829_ = sum_13[4] & q[19] /*36050*/;
  assign _2830_ = m_13[4] & _2828_ /*36049*/;
  assign r_13[23] = _2830_ | _2829_ /*36048*/;
  assign _2831_ = ~q[19] /*36047*/;
  assign _2832_ = sum_13[5] & q[19] /*36046*/;
  assign _2833_ = m_13[5] & _2831_ /*36045*/;
  assign r_13[24] = _2833_ | _2832_ /*36044*/;
  assign _2834_ = ~q[19] /*36043*/;
  assign _2835_ = sum_13[6] & q[19] /*36042*/;
  assign _2836_ = m_13[6] & _2834_ /*36041*/;
  assign r_13[25] = _2836_ | _2835_ /*36040*/;
  assign _2837_ = ~q[19] /*36039*/;
  assign _2838_ = sum_13[7] & q[19] /*36038*/;
  assign _2839_ = m_13[7] & _2837_ /*36037*/;
  assign r_13[26] = _2839_ | _2838_ /*36036*/;
  assign _2840_ = ~q[19] /*36035*/;
  assign _2841_ = sum_13[8] & q[19] /*36034*/;
  assign _2842_ = m_13[8] & _2840_ /*36033*/;
  assign r_13[27] = _2842_ | _2841_ /*36032*/;
  assign _2843_ = ~q[19] /*36031*/;
  assign _2844_ = sum_13[9] & q[19] /*36030*/;
  assign _2845_ = m_13[9] & _2843_ /*36029*/;
  assign r_13[28] = _2845_ | _2844_ /*36028*/;
  assign _2846_ = ~q[19] /*36027*/;
  assign _2847_ = sum_13[10] & q[19] /*36026*/;
  assign _2848_ = m_13[10] & _2846_ /*36025*/;
  assign r_13[29] = _2848_ | _2847_ /*36024*/;
  assign _2849_ = ~q[19] /*36023*/;
  assign _2850_ = sum_13[11] & q[19] /*36022*/;
  assign _2851_ = m_13[11] & _2849_ /*36021*/;
  assign r_13[30] = _2851_ | _2850_ /*36020*/;
  assign _2852_ = ~q[19] /*36019*/;
  assign _2853_ = sum_13[12] & q[19] /*36018*/;
  assign _2854_ = m_13[12] & _2852_ /*36017*/;
  assign r_13[31] = _2854_ | _2853_ /*36016*/;
  assign _2855_ = ~q[19] /*36015*/;
  assign _2856_ = sum_13[13] & q[19] /*36014*/;
  assign _2857_ = m_13[13] & _2855_ /*36013*/;
  assign r_13[32] = _2857_ | _2856_ /*36012*/;
  assign _2858_ = ~q[19] /*36011*/;
  assign _2859_ = sum_13[14] & q[19] /*36010*/;
  assign _2860_ = m_13[14] & _2858_ /*36009*/;
  assign r_13[33] = _2860_ | _2859_ /*36008*/;
  assign _2861_ = ~q[19] /*36007*/;
  assign _2862_ = sum_13[15] & q[19] /*36006*/;
  assign _2863_ = m_13[15] & _2861_ /*36005*/;
  assign r_13[34] = _2863_ | _2862_ /*36004*/;
  assign _2864_ = ~q[19] /*36003*/;
  assign _2865_ = sum_13[16] & q[19] /*36002*/;
  assign _2866_ = m_13[16] & _2864_ /*36001*/;
  assign r_13[35] = _2866_ | _2865_ /*36000*/;
  assign _2867_ = ~q[19] /*35999*/;
  assign _2868_ = sum_13[17] & q[19] /*35998*/;
  assign _2869_ = m_13[17] & _2867_ /*35997*/;
  assign r_13[36] = _2869_ | _2868_ /*35996*/;
  assign _2870_ = ~q[19] /*35995*/;
  assign _2871_ = sum_13[18] & q[19] /*35994*/;
  assign _2872_ = m_13[18] & _2870_ /*35993*/;
  assign r_13[37] = _2872_ | _2871_ /*35992*/;
  assign _2873_ = ~q[19] /*35991*/;
  assign _2874_ = sum_13[19] & q[19] /*35990*/;
  assign _2875_ = m_13[19] & _2873_ /*35989*/;
  assign r_13[38] = _2875_ | _2874_ /*35988*/;
  assign _2876_ = ~q[19] /*35987*/;
  assign _2877_ = sum_13[20] & q[19] /*35986*/;
  assign _2878_ = m_13[20] & _2876_ /*35985*/;
  assign r_13[39] = _2878_ | _2877_ /*35984*/;
  assign _2879_ = ~q[19] /*35983*/;
  assign _2880_ = sum_13[21] & q[19] /*35982*/;
  assign _2881_ = m_13[21] & _2879_ /*35981*/;
  assign r_13[40] = _2881_ | _2880_ /*35980*/;
  assign _2882_ = ~q[19] /*35979*/;
  assign _2883_ = sum_13[22] & q[19] /*35978*/;
  assign _2884_ = m_13[22] & _2882_ /*35977*/;
  assign r_13[41] = _2884_ | _2883_ /*35976*/;
  assign _2885_ = ~q[19] /*35975*/;
  assign _2886_ = sum_13[23] & q[19] /*35974*/;
  assign _2887_ = m_13[23] & _2885_ /*35973*/;
  assign r_13[42] = _2887_ | _2886_ /*35972*/;
  assign _2888_ = ~q[19] /*35971*/;
  assign _2889_ = sum_13[24] & q[19] /*35970*/;
  assign _2890_ = m_13[24] & _2888_ /*35969*/;
  assign r_13[43] = _2890_ | _2889_ /*35968*/;
  assign _2891_ = ~q[19] /*35967*/;
  assign _2892_ = sum_13[25] & q[19] /*35966*/;
  assign _2893_ = m_13[25] & _2891_ /*35965*/;
  assign r_13[44] = _2893_ | _2892_ /*35964*/;
  assign _2894_ = ~q[19] /*35963*/;
  assign _2895_ = sum_13[26] & q[19] /*35962*/;
  assign _2896_ = m_13[26] & _2894_ /*35961*/;
  assign r_13[45] = _2896_ | _2895_ /*35960*/;
  assign _2897_ = ~q[19] /*35959*/;
  assign _2898_ = sum_13[27] & q[19] /*35958*/;
  assign _2899_ = m_13[27] & _2897_ /*35957*/;
  assign r_13[46] = _2899_ | _2898_ /*35956*/;
  assign _2900_ = ~q[19] /*35955*/;
  assign _2901_ = sum_13[28] & q[19] /*35954*/;
  assign _2902_ = m_13[28] & _2900_ /*35953*/;
  assign r_13[47] = _2902_ | _2901_ /*35952*/;
  assign _2903_ = ~q[19] /*35951*/;
  assign _2904_ = sum_13[29] & q[19] /*35950*/;
  assign _2905_ = m_13[29] & _2903_ /*35949*/;
  assign r_13[48] = _2905_ | _2904_ /*35948*/;
  assign _2906_ = ~q[19] /*35947*/;
  assign _2907_ = sum_13[30] & q[19] /*35946*/;
  assign _2908_ = m_13[30] & _2906_ /*35945*/;
  assign r_13[49] = _2908_ | _2907_ /*35944*/;
  assign _2909_ = ~q[19] /*35943*/;
  assign _2910_ = sum_13[31] & q[19] /*35942*/;
  assign _2911_ = m_13[31] & _2909_ /*35941*/;
  assign r_13[50] = _2911_ | _2910_ /*35940*/;
assign r_13[0]= r_12[0] /*35939*/;
assign r_13[1]= r_12[1] /*35938*/;
assign r_13[2]= r_12[2] /*35937*/;
assign r_13[3]= r_12[3] /*35936*/;
assign r_13[4]= r_12[4] /*35935*/;
assign r_13[5]= r_12[5] /*35934*/;
assign r_13[6]= r_12[6] /*35933*/;
assign r_13[7]= r_12[7] /*35932*/;
assign r_13[8]= r_12[8] /*35931*/;
assign r_13[9]= r_12[9] /*35930*/;
assign r_13[10]= r_12[10] /*35929*/;
assign r_13[11]= r_12[11] /*35928*/;
assign r_13[12]= r_12[12] /*35927*/;
assign r_13[13]= r_12[13] /*35926*/;
assign r_13[14]= r_12[14] /*35925*/;
assign r_13[15]= r_12[15] /*35924*/;
assign r_13[16]= r_12[16] /*35923*/;
assign r_13[17]= r_12[17] /*35922*/;
assign r_13[18]= r_12[18] /*35921*/;
  assign inv_14[0] = ~div[0] /*35848*/;
  assign inv_14[1] = ~div[1] /*35847*/;
  assign inv_14[2] = ~div[2] /*35846*/;
  assign inv_14[3] = ~div[3] /*35845*/;
  assign inv_14[4] = ~div[4] /*35844*/;
  assign inv_14[5] = ~div[5] /*35843*/;
  assign inv_14[6] = ~div[6] /*35842*/;
  assign inv_14[7] = ~div[7] /*35841*/;
  assign inv_14[8] = ~div[8] /*35840*/;
  assign inv_14[9] = ~div[9] /*35839*/;
  assign inv_14[10] = ~div[10] /*35838*/;
  assign inv_14[11] = ~div[11] /*35837*/;
  assign inv_14[12] = ~div[12] /*35836*/;
  assign inv_14[13] = ~div[13] /*35835*/;
  assign inv_14[14] = ~div[14] /*35834*/;
  assign inv_14[15] = ~div[15] /*35833*/;
  assign inv_14[16] = ~div[16] /*35832*/;
  assign inv_14[17] = ~div[17] /*35831*/;
  assign inv_14[18] = ~div[18] /*35830*/;
  assign inv_14[19] = ~div[19] /*35829*/;
  assign inv_14[20] = ~div[20] /*35828*/;
  assign inv_14[21] = ~div[21] /*35827*/;
  assign inv_14[22] = ~div[22] /*35826*/;
  assign inv_14[23] = ~div[23] /*35825*/;
  assign inv_14[24] = ~div[24] /*35824*/;
  assign inv_14[25] = ~div[25] /*35823*/;
  assign inv_14[26] = ~div[26] /*35822*/;
  assign inv_14[27] = ~div[27] /*35821*/;
  assign inv_14[28] = ~div[28] /*35820*/;
  assign inv_14[29] = ~div[29] /*35819*/;
  assign inv_14[30] = ~div[30] /*35818*/;
assign inv_14[31] = oneWire /*35817*/;
  assign _2912_ = inv_14[0] ^ r_13[18] /*35815*/;
  assign sum_14[0] = _2912_ ^ oneWire /*35814*/;
  assign _2913_ = _2912_ & oneWire /*35813*/;
  assign _2914_ = inv_14[0] & r_13[18] /*35812*/;
  assign _2915_ = _2913_ | _2914_ /*35811*/;
  assign _2916_ = inv_14[1] ^ r_13[19] /*35810*/;
  assign sum_14[1] = _2916_ ^ _2915_ /*35809*/;
  assign _2917_ = _2916_ & _2915_ /*35808*/;
  assign _2918_ = inv_14[1] & r_13[19] /*35807*/;
  assign _2919_ = _2917_ | _2918_ /*35806*/;
  assign _2920_ = inv_14[2] ^ r_13[20] /*35804*/;
  assign sum_14[2] = _2920_ ^ _2919_ /*35803*/;
  assign _2921_ = _2920_ & _2919_ /*35802*/;
  assign _2922_ = inv_14[2] & r_13[20] /*35801*/;
  assign _2923_ = _2921_ | _2922_ /*35800*/;
  assign _2924_ = inv_14[3] ^ r_13[21] /*35798*/;
  assign sum_14[3] = _2924_ ^ _2923_ /*35797*/;
  assign _2925_ = _2924_ & _2923_ /*35796*/;
  assign _2926_ = inv_14[3] & r_13[21] /*35795*/;
  assign _2927_ = _2925_ | _2926_ /*35794*/;
  assign _2928_ = inv_14[4] ^ r_13[22] /*35792*/;
  assign sum_14[4] = _2928_ ^ _2927_ /*35791*/;
  assign _2929_ = _2928_ & _2927_ /*35790*/;
  assign _2930_ = inv_14[4] & r_13[22] /*35789*/;
  assign _2931_ = _2929_ | _2930_ /*35788*/;
  assign _2932_ = inv_14[5] ^ r_13[23] /*35786*/;
  assign sum_14[5] = _2932_ ^ _2931_ /*35785*/;
  assign _2933_ = _2932_ & _2931_ /*35784*/;
  assign _2934_ = inv_14[5] & r_13[23] /*35783*/;
  assign _2935_ = _2933_ | _2934_ /*35782*/;
  assign _2936_ = inv_14[6] ^ r_13[24] /*35780*/;
  assign sum_14[6] = _2936_ ^ _2935_ /*35779*/;
  assign _2937_ = _2936_ & _2935_ /*35778*/;
  assign _2938_ = inv_14[6] & r_13[24] /*35777*/;
  assign _2939_ = _2937_ | _2938_ /*35776*/;
  assign _2940_ = inv_14[7] ^ r_13[25] /*35774*/;
  assign sum_14[7] = _2940_ ^ _2939_ /*35773*/;
  assign _2941_ = _2940_ & _2939_ /*35772*/;
  assign _2942_ = inv_14[7] & r_13[25] /*35771*/;
  assign _2943_ = _2941_ | _2942_ /*35770*/;
  assign _2944_ = inv_14[8] ^ r_13[26] /*35768*/;
  assign sum_14[8] = _2944_ ^ _2943_ /*35767*/;
  assign _2945_ = _2944_ & _2943_ /*35766*/;
  assign _2946_ = inv_14[8] & r_13[26] /*35765*/;
  assign _2947_ = _2945_ | _2946_ /*35764*/;
  assign _2948_ = inv_14[9] ^ r_13[27] /*35762*/;
  assign sum_14[9] = _2948_ ^ _2947_ /*35761*/;
  assign _2949_ = _2948_ & _2947_ /*35760*/;
  assign _2950_ = inv_14[9] & r_13[27] /*35759*/;
  assign _2951_ = _2949_ | _2950_ /*35758*/;
  assign _2952_ = inv_14[10] ^ r_13[28] /*35756*/;
  assign sum_14[10] = _2952_ ^ _2951_ /*35755*/;
  assign _2953_ = _2952_ & _2951_ /*35754*/;
  assign _2954_ = inv_14[10] & r_13[28] /*35753*/;
  assign _2955_ = _2953_ | _2954_ /*35752*/;
  assign _2956_ = inv_14[11] ^ r_13[29] /*35750*/;
  assign sum_14[11] = _2956_ ^ _2955_ /*35749*/;
  assign _2957_ = _2956_ & _2955_ /*35748*/;
  assign _2958_ = inv_14[11] & r_13[29] /*35747*/;
  assign _2959_ = _2957_ | _2958_ /*35746*/;
  assign _2960_ = inv_14[12] ^ r_13[30] /*35744*/;
  assign sum_14[12] = _2960_ ^ _2959_ /*35743*/;
  assign _2961_ = _2960_ & _2959_ /*35742*/;
  assign _2962_ = inv_14[12] & r_13[30] /*35741*/;
  assign _2963_ = _2961_ | _2962_ /*35740*/;
  assign _2964_ = inv_14[13] ^ r_13[31] /*35738*/;
  assign sum_14[13] = _2964_ ^ _2963_ /*35737*/;
  assign _2965_ = _2964_ & _2963_ /*35736*/;
  assign _2966_ = inv_14[13] & r_13[31] /*35735*/;
  assign _2967_ = _2965_ | _2966_ /*35734*/;
  assign _2968_ = inv_14[14] ^ r_13[32] /*35732*/;
  assign sum_14[14] = _2968_ ^ _2967_ /*35731*/;
  assign _2969_ = _2968_ & _2967_ /*35730*/;
  assign _2970_ = inv_14[14] & r_13[32] /*35729*/;
  assign _2971_ = _2969_ | _2970_ /*35728*/;
  assign _2972_ = inv_14[15] ^ r_13[33] /*35726*/;
  assign sum_14[15] = _2972_ ^ _2971_ /*35725*/;
  assign _2973_ = _2972_ & _2971_ /*35724*/;
  assign _2974_ = inv_14[15] & r_13[33] /*35723*/;
  assign _2975_ = _2973_ | _2974_ /*35722*/;
  assign _2976_ = inv_14[16] ^ r_13[34] /*35720*/;
  assign sum_14[16] = _2976_ ^ _2975_ /*35719*/;
  assign _2977_ = _2976_ & _2975_ /*35718*/;
  assign _2978_ = inv_14[16] & r_13[34] /*35717*/;
  assign _2979_ = _2977_ | _2978_ /*35716*/;
  assign _2980_ = inv_14[17] ^ r_13[35] /*35714*/;
  assign sum_14[17] = _2980_ ^ _2979_ /*35713*/;
  assign _2981_ = _2980_ & _2979_ /*35712*/;
  assign _2982_ = inv_14[17] & r_13[35] /*35711*/;
  assign _2983_ = _2981_ | _2982_ /*35710*/;
  assign _2984_ = inv_14[18] ^ r_13[36] /*35708*/;
  assign sum_14[18] = _2984_ ^ _2983_ /*35707*/;
  assign _2985_ = _2984_ & _2983_ /*35706*/;
  assign _2986_ = inv_14[18] & r_13[36] /*35705*/;
  assign _2987_ = _2985_ | _2986_ /*35704*/;
  assign _2988_ = inv_14[19] ^ r_13[37] /*35702*/;
  assign sum_14[19] = _2988_ ^ _2987_ /*35701*/;
  assign _2989_ = _2988_ & _2987_ /*35700*/;
  assign _2990_ = inv_14[19] & r_13[37] /*35699*/;
  assign _2991_ = _2989_ | _2990_ /*35698*/;
  assign _2992_ = inv_14[20] ^ r_13[38] /*35696*/;
  assign sum_14[20] = _2992_ ^ _2991_ /*35695*/;
  assign _2993_ = _2992_ & _2991_ /*35694*/;
  assign _2994_ = inv_14[20] & r_13[38] /*35693*/;
  assign _2995_ = _2993_ | _2994_ /*35692*/;
  assign _2996_ = inv_14[21] ^ r_13[39] /*35690*/;
  assign sum_14[21] = _2996_ ^ _2995_ /*35689*/;
  assign _2997_ = _2996_ & _2995_ /*35688*/;
  assign _2998_ = inv_14[21] & r_13[39] /*35687*/;
  assign _2999_ = _2997_ | _2998_ /*35686*/;
  assign _3000_ = inv_14[22] ^ r_13[40] /*35684*/;
  assign sum_14[22] = _3000_ ^ _2999_ /*35683*/;
  assign _3001_ = _3000_ & _2999_ /*35682*/;
  assign _3002_ = inv_14[22] & r_13[40] /*35681*/;
  assign _3003_ = _3001_ | _3002_ /*35680*/;
  assign _3004_ = inv_14[23] ^ r_13[41] /*35678*/;
  assign sum_14[23] = _3004_ ^ _3003_ /*35677*/;
  assign _3005_ = _3004_ & _3003_ /*35676*/;
  assign _3006_ = inv_14[23] & r_13[41] /*35675*/;
  assign _3007_ = _3005_ | _3006_ /*35674*/;
  assign _3008_ = inv_14[24] ^ r_13[42] /*35672*/;
  assign sum_14[24] = _3008_ ^ _3007_ /*35671*/;
  assign _3009_ = _3008_ & _3007_ /*35670*/;
  assign _3010_ = inv_14[24] & r_13[42] /*35669*/;
  assign _3011_ = _3009_ | _3010_ /*35668*/;
  assign _3012_ = inv_14[25] ^ r_13[43] /*35666*/;
  assign sum_14[25] = _3012_ ^ _3011_ /*35665*/;
  assign _3013_ = _3012_ & _3011_ /*35664*/;
  assign _3014_ = inv_14[25] & r_13[43] /*35663*/;
  assign _3015_ = _3013_ | _3014_ /*35662*/;
  assign _3016_ = inv_14[26] ^ r_13[44] /*35660*/;
  assign sum_14[26] = _3016_ ^ _3015_ /*35659*/;
  assign _3017_ = _3016_ & _3015_ /*35658*/;
  assign _3018_ = inv_14[26] & r_13[44] /*35657*/;
  assign _3019_ = _3017_ | _3018_ /*35656*/;
  assign _3020_ = inv_14[27] ^ r_13[45] /*35654*/;
  assign sum_14[27] = _3020_ ^ _3019_ /*35653*/;
  assign _3021_ = _3020_ & _3019_ /*35652*/;
  assign _3022_ = inv_14[27] & r_13[45] /*35651*/;
  assign _3023_ = _3021_ | _3022_ /*35650*/;
  assign _3024_ = inv_14[28] ^ r_13[46] /*35648*/;
  assign sum_14[28] = _3024_ ^ _3023_ /*35647*/;
  assign _3025_ = _3024_ & _3023_ /*35646*/;
  assign _3026_ = inv_14[28] & r_13[46] /*35645*/;
  assign _3027_ = _3025_ | _3026_ /*35644*/;
  assign _3028_ = inv_14[29] ^ r_13[47] /*35642*/;
  assign sum_14[29] = _3028_ ^ _3027_ /*35641*/;
  assign _3029_ = _3028_ & _3027_ /*35640*/;
  assign _3030_ = inv_14[29] & r_13[47] /*35639*/;
  assign _3031_ = _3029_ | _3030_ /*35638*/;
  assign _3032_ = inv_14[30] ^ r_13[48] /*35636*/;
  assign sum_14[30] = _3032_ ^ _3031_ /*35635*/;
  assign _3033_ = _3032_ & _3031_ /*35634*/;
  assign _3034_ = inv_14[30] & r_13[48] /*35633*/;
  assign _3035_ = _3033_ | _3034_ /*35632*/;
  assign _3036_ = inv_14[31] ^ r_13[49] /*35630*/;
  assign sum_14[31] = _3036_ ^ _3035_ /*35629*/;
  assign _3037_ = _3036_ & _3035_ /*35628*/;
  assign _3038_ = inv_14[31] & r_13[49] /*35627*/;
  assign _3039_ = _3037_ | _3038_ /*35626*/;
  assign q[18] = ~sum_14[31] /*35653*/;
  assign m_14[0] = r_13[18] /*35652*/;
  assign m_14[1] = r_13[19] /*35651*/;
  assign m_14[2] = r_13[20] /*35650*/;
  assign m_14[3] = r_13[21] /*35649*/;
  assign m_14[4] = r_13[22] /*35648*/;
  assign m_14[5] = r_13[23] /*35647*/;
  assign m_14[6] = r_13[24] /*35646*/;
  assign m_14[7] = r_13[25] /*35645*/;
  assign m_14[8] = r_13[26] /*35644*/;
  assign m_14[9] = r_13[27] /*35643*/;
  assign m_14[10] = r_13[28] /*35642*/;
  assign m_14[11] = r_13[29] /*35641*/;
  assign m_14[12] = r_13[30] /*35640*/;
  assign m_14[13] = r_13[31] /*35639*/;
  assign m_14[14] = r_13[32] /*35638*/;
  assign m_14[15] = r_13[33] /*35637*/;
  assign m_14[16] = r_13[34] /*35636*/;
  assign m_14[17] = r_13[35] /*35635*/;
  assign m_14[18] = r_13[36] /*35634*/;
  assign m_14[19] = r_13[37] /*35633*/;
  assign m_14[20] = r_13[38] /*35632*/;
  assign m_14[21] = r_13[39] /*35631*/;
  assign m_14[22] = r_13[40] /*35630*/;
  assign m_14[23] = r_13[41] /*35629*/;
  assign m_14[24] = r_13[42] /*35628*/;
  assign m_14[25] = r_13[43] /*35627*/;
  assign m_14[26] = r_13[44] /*35626*/;
  assign m_14[27] = r_13[45] /*35625*/;
  assign m_14[28] = r_13[46] /*35624*/;
  assign m_14[29] = r_13[47] /*35623*/;
  assign m_14[30] = r_13[48] /*35622*/;
  assign m_14[31] = r_13[49] /*35621*/;
  assign _3040_ = ~q[18] /*35619*/;
  assign _3041_ = sum_14[0] & q[18] /*35618*/;
  assign _3042_ = m_14[0] & _3040_ /*35617*/;
  assign r_14[18] = _3042_ | _3041_ /*35616*/;
  assign _3043_ = ~q[18] /*35615*/;
  assign _3044_ = sum_14[1] & q[18] /*35614*/;
  assign _3045_ = m_14[1] & _3043_ /*35613*/;
  assign r_14[19] = _3045_ | _3044_ /*35612*/;
  assign _3046_ = ~q[18] /*35611*/;
  assign _3047_ = sum_14[2] & q[18] /*35610*/;
  assign _3048_ = m_14[2] & _3046_ /*35609*/;
  assign r_14[20] = _3048_ | _3047_ /*35608*/;
  assign _3049_ = ~q[18] /*35607*/;
  assign _3050_ = sum_14[3] & q[18] /*35606*/;
  assign _3051_ = m_14[3] & _3049_ /*35605*/;
  assign r_14[21] = _3051_ | _3050_ /*35604*/;
  assign _3052_ = ~q[18] /*35603*/;
  assign _3053_ = sum_14[4] & q[18] /*35602*/;
  assign _3054_ = m_14[4] & _3052_ /*35601*/;
  assign r_14[22] = _3054_ | _3053_ /*35600*/;
  assign _3055_ = ~q[18] /*35599*/;
  assign _3056_ = sum_14[5] & q[18] /*35598*/;
  assign _3057_ = m_14[5] & _3055_ /*35597*/;
  assign r_14[23] = _3057_ | _3056_ /*35596*/;
  assign _3058_ = ~q[18] /*35595*/;
  assign _3059_ = sum_14[6] & q[18] /*35594*/;
  assign _3060_ = m_14[6] & _3058_ /*35593*/;
  assign r_14[24] = _3060_ | _3059_ /*35592*/;
  assign _3061_ = ~q[18] /*35591*/;
  assign _3062_ = sum_14[7] & q[18] /*35590*/;
  assign _3063_ = m_14[7] & _3061_ /*35589*/;
  assign r_14[25] = _3063_ | _3062_ /*35588*/;
  assign _3064_ = ~q[18] /*35587*/;
  assign _3065_ = sum_14[8] & q[18] /*35586*/;
  assign _3066_ = m_14[8] & _3064_ /*35585*/;
  assign r_14[26] = _3066_ | _3065_ /*35584*/;
  assign _3067_ = ~q[18] /*35583*/;
  assign _3068_ = sum_14[9] & q[18] /*35582*/;
  assign _3069_ = m_14[9] & _3067_ /*35581*/;
  assign r_14[27] = _3069_ | _3068_ /*35580*/;
  assign _3070_ = ~q[18] /*35579*/;
  assign _3071_ = sum_14[10] & q[18] /*35578*/;
  assign _3072_ = m_14[10] & _3070_ /*35577*/;
  assign r_14[28] = _3072_ | _3071_ /*35576*/;
  assign _3073_ = ~q[18] /*35575*/;
  assign _3074_ = sum_14[11] & q[18] /*35574*/;
  assign _3075_ = m_14[11] & _3073_ /*35573*/;
  assign r_14[29] = _3075_ | _3074_ /*35572*/;
  assign _3076_ = ~q[18] /*35571*/;
  assign _3077_ = sum_14[12] & q[18] /*35570*/;
  assign _3078_ = m_14[12] & _3076_ /*35569*/;
  assign r_14[30] = _3078_ | _3077_ /*35568*/;
  assign _3079_ = ~q[18] /*35567*/;
  assign _3080_ = sum_14[13] & q[18] /*35566*/;
  assign _3081_ = m_14[13] & _3079_ /*35565*/;
  assign r_14[31] = _3081_ | _3080_ /*35564*/;
  assign _3082_ = ~q[18] /*35563*/;
  assign _3083_ = sum_14[14] & q[18] /*35562*/;
  assign _3084_ = m_14[14] & _3082_ /*35561*/;
  assign r_14[32] = _3084_ | _3083_ /*35560*/;
  assign _3085_ = ~q[18] /*35559*/;
  assign _3086_ = sum_14[15] & q[18] /*35558*/;
  assign _3087_ = m_14[15] & _3085_ /*35557*/;
  assign r_14[33] = _3087_ | _3086_ /*35556*/;
  assign _3088_ = ~q[18] /*35555*/;
  assign _3089_ = sum_14[16] & q[18] /*35554*/;
  assign _3090_ = m_14[16] & _3088_ /*35553*/;
  assign r_14[34] = _3090_ | _3089_ /*35552*/;
  assign _3091_ = ~q[18] /*35551*/;
  assign _3092_ = sum_14[17] & q[18] /*35550*/;
  assign _3093_ = m_14[17] & _3091_ /*35549*/;
  assign r_14[35] = _3093_ | _3092_ /*35548*/;
  assign _3094_ = ~q[18] /*35547*/;
  assign _3095_ = sum_14[18] & q[18] /*35546*/;
  assign _3096_ = m_14[18] & _3094_ /*35545*/;
  assign r_14[36] = _3096_ | _3095_ /*35544*/;
  assign _3097_ = ~q[18] /*35543*/;
  assign _3098_ = sum_14[19] & q[18] /*35542*/;
  assign _3099_ = m_14[19] & _3097_ /*35541*/;
  assign r_14[37] = _3099_ | _3098_ /*35540*/;
  assign _3100_ = ~q[18] /*35539*/;
  assign _3101_ = sum_14[20] & q[18] /*35538*/;
  assign _3102_ = m_14[20] & _3100_ /*35537*/;
  assign r_14[38] = _3102_ | _3101_ /*35536*/;
  assign _3103_ = ~q[18] /*35535*/;
  assign _3104_ = sum_14[21] & q[18] /*35534*/;
  assign _3105_ = m_14[21] & _3103_ /*35533*/;
  assign r_14[39] = _3105_ | _3104_ /*35532*/;
  assign _3106_ = ~q[18] /*35531*/;
  assign _3107_ = sum_14[22] & q[18] /*35530*/;
  assign _3108_ = m_14[22] & _3106_ /*35529*/;
  assign r_14[40] = _3108_ | _3107_ /*35528*/;
  assign _3109_ = ~q[18] /*35527*/;
  assign _3110_ = sum_14[23] & q[18] /*35526*/;
  assign _3111_ = m_14[23] & _3109_ /*35525*/;
  assign r_14[41] = _3111_ | _3110_ /*35524*/;
  assign _3112_ = ~q[18] /*35523*/;
  assign _3113_ = sum_14[24] & q[18] /*35522*/;
  assign _3114_ = m_14[24] & _3112_ /*35521*/;
  assign r_14[42] = _3114_ | _3113_ /*35520*/;
  assign _3115_ = ~q[18] /*35519*/;
  assign _3116_ = sum_14[25] & q[18] /*35518*/;
  assign _3117_ = m_14[25] & _3115_ /*35517*/;
  assign r_14[43] = _3117_ | _3116_ /*35516*/;
  assign _3118_ = ~q[18] /*35515*/;
  assign _3119_ = sum_14[26] & q[18] /*35514*/;
  assign _3120_ = m_14[26] & _3118_ /*35513*/;
  assign r_14[44] = _3120_ | _3119_ /*35512*/;
  assign _3121_ = ~q[18] /*35511*/;
  assign _3122_ = sum_14[27] & q[18] /*35510*/;
  assign _3123_ = m_14[27] & _3121_ /*35509*/;
  assign r_14[45] = _3123_ | _3122_ /*35508*/;
  assign _3124_ = ~q[18] /*35507*/;
  assign _3125_ = sum_14[28] & q[18] /*35506*/;
  assign _3126_ = m_14[28] & _3124_ /*35505*/;
  assign r_14[46] = _3126_ | _3125_ /*35504*/;
  assign _3127_ = ~q[18] /*35503*/;
  assign _3128_ = sum_14[29] & q[18] /*35502*/;
  assign _3129_ = m_14[29] & _3127_ /*35501*/;
  assign r_14[47] = _3129_ | _3128_ /*35500*/;
  assign _3130_ = ~q[18] /*35499*/;
  assign _3131_ = sum_14[30] & q[18] /*35498*/;
  assign _3132_ = m_14[30] & _3130_ /*35497*/;
  assign r_14[48] = _3132_ | _3131_ /*35496*/;
  assign _3133_ = ~q[18] /*35495*/;
  assign _3134_ = sum_14[31] & q[18] /*35494*/;
  assign _3135_ = m_14[31] & _3133_ /*35493*/;
  assign r_14[49] = _3135_ | _3134_ /*35492*/;
assign r_14[0]= r_13[0] /*35491*/;
assign r_14[1]= r_13[1] /*35490*/;
assign r_14[2]= r_13[2] /*35489*/;
assign r_14[3]= r_13[3] /*35488*/;
assign r_14[4]= r_13[4] /*35487*/;
assign r_14[5]= r_13[5] /*35486*/;
assign r_14[6]= r_13[6] /*35485*/;
assign r_14[7]= r_13[7] /*35484*/;
assign r_14[8]= r_13[8] /*35483*/;
assign r_14[9]= r_13[9] /*35482*/;
assign r_14[10]= r_13[10] /*35481*/;
assign r_14[11]= r_13[11] /*35480*/;
assign r_14[12]= r_13[12] /*35479*/;
assign r_14[13]= r_13[13] /*35478*/;
assign r_14[14]= r_13[14] /*35477*/;
assign r_14[15]= r_13[15] /*35476*/;
assign r_14[16]= r_13[16] /*35475*/;
assign r_14[17]= r_13[17] /*35474*/;
  assign inv_15[0] = ~div[0] /*35400*/;
  assign inv_15[1] = ~div[1] /*35399*/;
  assign inv_15[2] = ~div[2] /*35398*/;
  assign inv_15[3] = ~div[3] /*35397*/;
  assign inv_15[4] = ~div[4] /*35396*/;
  assign inv_15[5] = ~div[5] /*35395*/;
  assign inv_15[6] = ~div[6] /*35394*/;
  assign inv_15[7] = ~div[7] /*35393*/;
  assign inv_15[8] = ~div[8] /*35392*/;
  assign inv_15[9] = ~div[9] /*35391*/;
  assign inv_15[10] = ~div[10] /*35390*/;
  assign inv_15[11] = ~div[11] /*35389*/;
  assign inv_15[12] = ~div[12] /*35388*/;
  assign inv_15[13] = ~div[13] /*35387*/;
  assign inv_15[14] = ~div[14] /*35386*/;
  assign inv_15[15] = ~div[15] /*35385*/;
  assign inv_15[16] = ~div[16] /*35384*/;
  assign inv_15[17] = ~div[17] /*35383*/;
  assign inv_15[18] = ~div[18] /*35382*/;
  assign inv_15[19] = ~div[19] /*35381*/;
  assign inv_15[20] = ~div[20] /*35380*/;
  assign inv_15[21] = ~div[21] /*35379*/;
  assign inv_15[22] = ~div[22] /*35378*/;
  assign inv_15[23] = ~div[23] /*35377*/;
  assign inv_15[24] = ~div[24] /*35376*/;
  assign inv_15[25] = ~div[25] /*35375*/;
  assign inv_15[26] = ~div[26] /*35374*/;
  assign inv_15[27] = ~div[27] /*35373*/;
  assign inv_15[28] = ~div[28] /*35372*/;
  assign inv_15[29] = ~div[29] /*35371*/;
  assign inv_15[30] = ~div[30] /*35370*/;
assign inv_15[31] = oneWire /*35369*/;
  assign _3136_ = inv_15[0] ^ r_14[17] /*35367*/;
  assign sum_15[0] = _3136_ ^ oneWire /*35366*/;
  assign _3137_ = _3136_ & oneWire /*35365*/;
  assign _3138_ = inv_15[0] & r_14[17] /*35364*/;
  assign _3139_ = _3137_ | _3138_ /*35363*/;
  assign _3140_ = inv_15[1] ^ r_14[18] /*35362*/;
  assign sum_15[1] = _3140_ ^ _3139_ /*35361*/;
  assign _3141_ = _3140_ & _3139_ /*35360*/;
  assign _3142_ = inv_15[1] & r_14[18] /*35359*/;
  assign _3143_ = _3141_ | _3142_ /*35358*/;
  assign _3144_ = inv_15[2] ^ r_14[19] /*35356*/;
  assign sum_15[2] = _3144_ ^ _3143_ /*35355*/;
  assign _3145_ = _3144_ & _3143_ /*35354*/;
  assign _3146_ = inv_15[2] & r_14[19] /*35353*/;
  assign _3147_ = _3145_ | _3146_ /*35352*/;
  assign _3148_ = inv_15[3] ^ r_14[20] /*35350*/;
  assign sum_15[3] = _3148_ ^ _3147_ /*35349*/;
  assign _3149_ = _3148_ & _3147_ /*35348*/;
  assign _3150_ = inv_15[3] & r_14[20] /*35347*/;
  assign _3151_ = _3149_ | _3150_ /*35346*/;
  assign _3152_ = inv_15[4] ^ r_14[21] /*35344*/;
  assign sum_15[4] = _3152_ ^ _3151_ /*35343*/;
  assign _3153_ = _3152_ & _3151_ /*35342*/;
  assign _3154_ = inv_15[4] & r_14[21] /*35341*/;
  assign _3155_ = _3153_ | _3154_ /*35340*/;
  assign _3156_ = inv_15[5] ^ r_14[22] /*35338*/;
  assign sum_15[5] = _3156_ ^ _3155_ /*35337*/;
  assign _3157_ = _3156_ & _3155_ /*35336*/;
  assign _3158_ = inv_15[5] & r_14[22] /*35335*/;
  assign _3159_ = _3157_ | _3158_ /*35334*/;
  assign _3160_ = inv_15[6] ^ r_14[23] /*35332*/;
  assign sum_15[6] = _3160_ ^ _3159_ /*35331*/;
  assign _3161_ = _3160_ & _3159_ /*35330*/;
  assign _3162_ = inv_15[6] & r_14[23] /*35329*/;
  assign _3163_ = _3161_ | _3162_ /*35328*/;
  assign _3164_ = inv_15[7] ^ r_14[24] /*35326*/;
  assign sum_15[7] = _3164_ ^ _3163_ /*35325*/;
  assign _3165_ = _3164_ & _3163_ /*35324*/;
  assign _3166_ = inv_15[7] & r_14[24] /*35323*/;
  assign _3167_ = _3165_ | _3166_ /*35322*/;
  assign _3168_ = inv_15[8] ^ r_14[25] /*35320*/;
  assign sum_15[8] = _3168_ ^ _3167_ /*35319*/;
  assign _3169_ = _3168_ & _3167_ /*35318*/;
  assign _3170_ = inv_15[8] & r_14[25] /*35317*/;
  assign _3171_ = _3169_ | _3170_ /*35316*/;
  assign _3172_ = inv_15[9] ^ r_14[26] /*35314*/;
  assign sum_15[9] = _3172_ ^ _3171_ /*35313*/;
  assign _3173_ = _3172_ & _3171_ /*35312*/;
  assign _3174_ = inv_15[9] & r_14[26] /*35311*/;
  assign _3175_ = _3173_ | _3174_ /*35310*/;
  assign _3176_ = inv_15[10] ^ r_14[27] /*35308*/;
  assign sum_15[10] = _3176_ ^ _3175_ /*35307*/;
  assign _3177_ = _3176_ & _3175_ /*35306*/;
  assign _3178_ = inv_15[10] & r_14[27] /*35305*/;
  assign _3179_ = _3177_ | _3178_ /*35304*/;
  assign _3180_ = inv_15[11] ^ r_14[28] /*35302*/;
  assign sum_15[11] = _3180_ ^ _3179_ /*35301*/;
  assign _3181_ = _3180_ & _3179_ /*35300*/;
  assign _3182_ = inv_15[11] & r_14[28] /*35299*/;
  assign _3183_ = _3181_ | _3182_ /*35298*/;
  assign _3184_ = inv_15[12] ^ r_14[29] /*35296*/;
  assign sum_15[12] = _3184_ ^ _3183_ /*35295*/;
  assign _3185_ = _3184_ & _3183_ /*35294*/;
  assign _3186_ = inv_15[12] & r_14[29] /*35293*/;
  assign _3187_ = _3185_ | _3186_ /*35292*/;
  assign _3188_ = inv_15[13] ^ r_14[30] /*35290*/;
  assign sum_15[13] = _3188_ ^ _3187_ /*35289*/;
  assign _3189_ = _3188_ & _3187_ /*35288*/;
  assign _3190_ = inv_15[13] & r_14[30] /*35287*/;
  assign _3191_ = _3189_ | _3190_ /*35286*/;
  assign _3192_ = inv_15[14] ^ r_14[31] /*35284*/;
  assign sum_15[14] = _3192_ ^ _3191_ /*35283*/;
  assign _3193_ = _3192_ & _3191_ /*35282*/;
  assign _3194_ = inv_15[14] & r_14[31] /*35281*/;
  assign _3195_ = _3193_ | _3194_ /*35280*/;
  assign _3196_ = inv_15[15] ^ r_14[32] /*35278*/;
  assign sum_15[15] = _3196_ ^ _3195_ /*35277*/;
  assign _3197_ = _3196_ & _3195_ /*35276*/;
  assign _3198_ = inv_15[15] & r_14[32] /*35275*/;
  assign _3199_ = _3197_ | _3198_ /*35274*/;
  assign _3200_ = inv_15[16] ^ r_14[33] /*35272*/;
  assign sum_15[16] = _3200_ ^ _3199_ /*35271*/;
  assign _3201_ = _3200_ & _3199_ /*35270*/;
  assign _3202_ = inv_15[16] & r_14[33] /*35269*/;
  assign _3203_ = _3201_ | _3202_ /*35268*/;
  assign _3204_ = inv_15[17] ^ r_14[34] /*35266*/;
  assign sum_15[17] = _3204_ ^ _3203_ /*35265*/;
  assign _3205_ = _3204_ & _3203_ /*35264*/;
  assign _3206_ = inv_15[17] & r_14[34] /*35263*/;
  assign _3207_ = _3205_ | _3206_ /*35262*/;
  assign _3208_ = inv_15[18] ^ r_14[35] /*35260*/;
  assign sum_15[18] = _3208_ ^ _3207_ /*35259*/;
  assign _3209_ = _3208_ & _3207_ /*35258*/;
  assign _3210_ = inv_15[18] & r_14[35] /*35257*/;
  assign _3211_ = _3209_ | _3210_ /*35256*/;
  assign _3212_ = inv_15[19] ^ r_14[36] /*35254*/;
  assign sum_15[19] = _3212_ ^ _3211_ /*35253*/;
  assign _3213_ = _3212_ & _3211_ /*35252*/;
  assign _3214_ = inv_15[19] & r_14[36] /*35251*/;
  assign _3215_ = _3213_ | _3214_ /*35250*/;
  assign _3216_ = inv_15[20] ^ r_14[37] /*35248*/;
  assign sum_15[20] = _3216_ ^ _3215_ /*35247*/;
  assign _3217_ = _3216_ & _3215_ /*35246*/;
  assign _3218_ = inv_15[20] & r_14[37] /*35245*/;
  assign _3219_ = _3217_ | _3218_ /*35244*/;
  assign _3220_ = inv_15[21] ^ r_14[38] /*35242*/;
  assign sum_15[21] = _3220_ ^ _3219_ /*35241*/;
  assign _3221_ = _3220_ & _3219_ /*35240*/;
  assign _3222_ = inv_15[21] & r_14[38] /*35239*/;
  assign _3223_ = _3221_ | _3222_ /*35238*/;
  assign _3224_ = inv_15[22] ^ r_14[39] /*35236*/;
  assign sum_15[22] = _3224_ ^ _3223_ /*35235*/;
  assign _3225_ = _3224_ & _3223_ /*35234*/;
  assign _3226_ = inv_15[22] & r_14[39] /*35233*/;
  assign _3227_ = _3225_ | _3226_ /*35232*/;
  assign _3228_ = inv_15[23] ^ r_14[40] /*35230*/;
  assign sum_15[23] = _3228_ ^ _3227_ /*35229*/;
  assign _3229_ = _3228_ & _3227_ /*35228*/;
  assign _3230_ = inv_15[23] & r_14[40] /*35227*/;
  assign _3231_ = _3229_ | _3230_ /*35226*/;
  assign _3232_ = inv_15[24] ^ r_14[41] /*35224*/;
  assign sum_15[24] = _3232_ ^ _3231_ /*35223*/;
  assign _3233_ = _3232_ & _3231_ /*35222*/;
  assign _3234_ = inv_15[24] & r_14[41] /*35221*/;
  assign _3235_ = _3233_ | _3234_ /*35220*/;
  assign _3236_ = inv_15[25] ^ r_14[42] /*35218*/;
  assign sum_15[25] = _3236_ ^ _3235_ /*35217*/;
  assign _3237_ = _3236_ & _3235_ /*35216*/;
  assign _3238_ = inv_15[25] & r_14[42] /*35215*/;
  assign _3239_ = _3237_ | _3238_ /*35214*/;
  assign _3240_ = inv_15[26] ^ r_14[43] /*35212*/;
  assign sum_15[26] = _3240_ ^ _3239_ /*35211*/;
  assign _3241_ = _3240_ & _3239_ /*35210*/;
  assign _3242_ = inv_15[26] & r_14[43] /*35209*/;
  assign _3243_ = _3241_ | _3242_ /*35208*/;
  assign _3244_ = inv_15[27] ^ r_14[44] /*35206*/;
  assign sum_15[27] = _3244_ ^ _3243_ /*35205*/;
  assign _3245_ = _3244_ & _3243_ /*35204*/;
  assign _3246_ = inv_15[27] & r_14[44] /*35203*/;
  assign _3247_ = _3245_ | _3246_ /*35202*/;
  assign _3248_ = inv_15[28] ^ r_14[45] /*35200*/;
  assign sum_15[28] = _3248_ ^ _3247_ /*35199*/;
  assign _3249_ = _3248_ & _3247_ /*35198*/;
  assign _3250_ = inv_15[28] & r_14[45] /*35197*/;
  assign _3251_ = _3249_ | _3250_ /*35196*/;
  assign _3252_ = inv_15[29] ^ r_14[46] /*35194*/;
  assign sum_15[29] = _3252_ ^ _3251_ /*35193*/;
  assign _3253_ = _3252_ & _3251_ /*35192*/;
  assign _3254_ = inv_15[29] & r_14[46] /*35191*/;
  assign _3255_ = _3253_ | _3254_ /*35190*/;
  assign _3256_ = inv_15[30] ^ r_14[47] /*35188*/;
  assign sum_15[30] = _3256_ ^ _3255_ /*35187*/;
  assign _3257_ = _3256_ & _3255_ /*35186*/;
  assign _3258_ = inv_15[30] & r_14[47] /*35185*/;
  assign _3259_ = _3257_ | _3258_ /*35184*/;
  assign _3260_ = inv_15[31] ^ r_14[48] /*35182*/;
  assign sum_15[31] = _3260_ ^ _3259_ /*35181*/;
  assign _3261_ = _3260_ & _3259_ /*35180*/;
  assign _3262_ = inv_15[31] & r_14[48] /*35179*/;
  assign _3263_ = _3261_ | _3262_ /*35178*/;
  assign q[17] = ~sum_15[31] /*35205*/;
  assign m_15[0] = r_14[17] /*35204*/;
  assign m_15[1] = r_14[18] /*35203*/;
  assign m_15[2] = r_14[19] /*35202*/;
  assign m_15[3] = r_14[20] /*35201*/;
  assign m_15[4] = r_14[21] /*35200*/;
  assign m_15[5] = r_14[22] /*35199*/;
  assign m_15[6] = r_14[23] /*35198*/;
  assign m_15[7] = r_14[24] /*35197*/;
  assign m_15[8] = r_14[25] /*35196*/;
  assign m_15[9] = r_14[26] /*35195*/;
  assign m_15[10] = r_14[27] /*35194*/;
  assign m_15[11] = r_14[28] /*35193*/;
  assign m_15[12] = r_14[29] /*35192*/;
  assign m_15[13] = r_14[30] /*35191*/;
  assign m_15[14] = r_14[31] /*35190*/;
  assign m_15[15] = r_14[32] /*35189*/;
  assign m_15[16] = r_14[33] /*35188*/;
  assign m_15[17] = r_14[34] /*35187*/;
  assign m_15[18] = r_14[35] /*35186*/;
  assign m_15[19] = r_14[36] /*35185*/;
  assign m_15[20] = r_14[37] /*35184*/;
  assign m_15[21] = r_14[38] /*35183*/;
  assign m_15[22] = r_14[39] /*35182*/;
  assign m_15[23] = r_14[40] /*35181*/;
  assign m_15[24] = r_14[41] /*35180*/;
  assign m_15[25] = r_14[42] /*35179*/;
  assign m_15[26] = r_14[43] /*35178*/;
  assign m_15[27] = r_14[44] /*35177*/;
  assign m_15[28] = r_14[45] /*35176*/;
  assign m_15[29] = r_14[46] /*35175*/;
  assign m_15[30] = r_14[47] /*35174*/;
  assign m_15[31] = r_14[48] /*35173*/;
  assign _3264_ = ~q[17] /*35171*/;
  assign _3265_ = sum_15[0] & q[17] /*35170*/;
  assign _3266_ = m_15[0] & _3264_ /*35169*/;
  assign r_15[17] = _3266_ | _3265_ /*35168*/;
  assign _3267_ = ~q[17] /*35167*/;
  assign _3268_ = sum_15[1] & q[17] /*35166*/;
  assign _3269_ = m_15[1] & _3267_ /*35165*/;
  assign r_15[18] = _3269_ | _3268_ /*35164*/;
  assign _3270_ = ~q[17] /*35163*/;
  assign _3271_ = sum_15[2] & q[17] /*35162*/;
  assign _3272_ = m_15[2] & _3270_ /*35161*/;
  assign r_15[19] = _3272_ | _3271_ /*35160*/;
  assign _3273_ = ~q[17] /*35159*/;
  assign _3274_ = sum_15[3] & q[17] /*35158*/;
  assign _3275_ = m_15[3] & _3273_ /*35157*/;
  assign r_15[20] = _3275_ | _3274_ /*35156*/;
  assign _3276_ = ~q[17] /*35155*/;
  assign _3277_ = sum_15[4] & q[17] /*35154*/;
  assign _3278_ = m_15[4] & _3276_ /*35153*/;
  assign r_15[21] = _3278_ | _3277_ /*35152*/;
  assign _3279_ = ~q[17] /*35151*/;
  assign _3280_ = sum_15[5] & q[17] /*35150*/;
  assign _3281_ = m_15[5] & _3279_ /*35149*/;
  assign r_15[22] = _3281_ | _3280_ /*35148*/;
  assign _3282_ = ~q[17] /*35147*/;
  assign _3283_ = sum_15[6] & q[17] /*35146*/;
  assign _3284_ = m_15[6] & _3282_ /*35145*/;
  assign r_15[23] = _3284_ | _3283_ /*35144*/;
  assign _3285_ = ~q[17] /*35143*/;
  assign _3286_ = sum_15[7] & q[17] /*35142*/;
  assign _3287_ = m_15[7] & _3285_ /*35141*/;
  assign r_15[24] = _3287_ | _3286_ /*35140*/;
  assign _3288_ = ~q[17] /*35139*/;
  assign _3289_ = sum_15[8] & q[17] /*35138*/;
  assign _3290_ = m_15[8] & _3288_ /*35137*/;
  assign r_15[25] = _3290_ | _3289_ /*35136*/;
  assign _3291_ = ~q[17] /*35135*/;
  assign _3292_ = sum_15[9] & q[17] /*35134*/;
  assign _3293_ = m_15[9] & _3291_ /*35133*/;
  assign r_15[26] = _3293_ | _3292_ /*35132*/;
  assign _3294_ = ~q[17] /*35131*/;
  assign _3295_ = sum_15[10] & q[17] /*35130*/;
  assign _3296_ = m_15[10] & _3294_ /*35129*/;
  assign r_15[27] = _3296_ | _3295_ /*35128*/;
  assign _3297_ = ~q[17] /*35127*/;
  assign _3298_ = sum_15[11] & q[17] /*35126*/;
  assign _3299_ = m_15[11] & _3297_ /*35125*/;
  assign r_15[28] = _3299_ | _3298_ /*35124*/;
  assign _3300_ = ~q[17] /*35123*/;
  assign _3301_ = sum_15[12] & q[17] /*35122*/;
  assign _3302_ = m_15[12] & _3300_ /*35121*/;
  assign r_15[29] = _3302_ | _3301_ /*35120*/;
  assign _3303_ = ~q[17] /*35119*/;
  assign _3304_ = sum_15[13] & q[17] /*35118*/;
  assign _3305_ = m_15[13] & _3303_ /*35117*/;
  assign r_15[30] = _3305_ | _3304_ /*35116*/;
  assign _3306_ = ~q[17] /*35115*/;
  assign _3307_ = sum_15[14] & q[17] /*35114*/;
  assign _3308_ = m_15[14] & _3306_ /*35113*/;
  assign r_15[31] = _3308_ | _3307_ /*35112*/;
  assign _3309_ = ~q[17] /*35111*/;
  assign _3310_ = sum_15[15] & q[17] /*35110*/;
  assign _3311_ = m_15[15] & _3309_ /*35109*/;
  assign r_15[32] = _3311_ | _3310_ /*35108*/;
  assign _3312_ = ~q[17] /*35107*/;
  assign _3313_ = sum_15[16] & q[17] /*35106*/;
  assign _3314_ = m_15[16] & _3312_ /*35105*/;
  assign r_15[33] = _3314_ | _3313_ /*35104*/;
  assign _3315_ = ~q[17] /*35103*/;
  assign _3316_ = sum_15[17] & q[17] /*35102*/;
  assign _3317_ = m_15[17] & _3315_ /*35101*/;
  assign r_15[34] = _3317_ | _3316_ /*35100*/;
  assign _3318_ = ~q[17] /*35099*/;
  assign _3319_ = sum_15[18] & q[17] /*35098*/;
  assign _3320_ = m_15[18] & _3318_ /*35097*/;
  assign r_15[35] = _3320_ | _3319_ /*35096*/;
  assign _3321_ = ~q[17] /*35095*/;
  assign _3322_ = sum_15[19] & q[17] /*35094*/;
  assign _3323_ = m_15[19] & _3321_ /*35093*/;
  assign r_15[36] = _3323_ | _3322_ /*35092*/;
  assign _3324_ = ~q[17] /*35091*/;
  assign _3325_ = sum_15[20] & q[17] /*35090*/;
  assign _3326_ = m_15[20] & _3324_ /*35089*/;
  assign r_15[37] = _3326_ | _3325_ /*35088*/;
  assign _3327_ = ~q[17] /*35087*/;
  assign _3328_ = sum_15[21] & q[17] /*35086*/;
  assign _3329_ = m_15[21] & _3327_ /*35085*/;
  assign r_15[38] = _3329_ | _3328_ /*35084*/;
  assign _3330_ = ~q[17] /*35083*/;
  assign _3331_ = sum_15[22] & q[17] /*35082*/;
  assign _3332_ = m_15[22] & _3330_ /*35081*/;
  assign r_15[39] = _3332_ | _3331_ /*35080*/;
  assign _3333_ = ~q[17] /*35079*/;
  assign _3334_ = sum_15[23] & q[17] /*35078*/;
  assign _3335_ = m_15[23] & _3333_ /*35077*/;
  assign r_15[40] = _3335_ | _3334_ /*35076*/;
  assign _3336_ = ~q[17] /*35075*/;
  assign _3337_ = sum_15[24] & q[17] /*35074*/;
  assign _3338_ = m_15[24] & _3336_ /*35073*/;
  assign r_15[41] = _3338_ | _3337_ /*35072*/;
  assign _3339_ = ~q[17] /*35071*/;
  assign _3340_ = sum_15[25] & q[17] /*35070*/;
  assign _3341_ = m_15[25] & _3339_ /*35069*/;
  assign r_15[42] = _3341_ | _3340_ /*35068*/;
  assign _3342_ = ~q[17] /*35067*/;
  assign _3343_ = sum_15[26] & q[17] /*35066*/;
  assign _3344_ = m_15[26] & _3342_ /*35065*/;
  assign r_15[43] = _3344_ | _3343_ /*35064*/;
  assign _3345_ = ~q[17] /*35063*/;
  assign _3346_ = sum_15[27] & q[17] /*35062*/;
  assign _3347_ = m_15[27] & _3345_ /*35061*/;
  assign r_15[44] = _3347_ | _3346_ /*35060*/;
  assign _3348_ = ~q[17] /*35059*/;
  assign _3349_ = sum_15[28] & q[17] /*35058*/;
  assign _3350_ = m_15[28] & _3348_ /*35057*/;
  assign r_15[45] = _3350_ | _3349_ /*35056*/;
  assign _3351_ = ~q[17] /*35055*/;
  assign _3352_ = sum_15[29] & q[17] /*35054*/;
  assign _3353_ = m_15[29] & _3351_ /*35053*/;
  assign r_15[46] = _3353_ | _3352_ /*35052*/;
  assign _3354_ = ~q[17] /*35051*/;
  assign _3355_ = sum_15[30] & q[17] /*35050*/;
  assign _3356_ = m_15[30] & _3354_ /*35049*/;
  assign r_15[47] = _3356_ | _3355_ /*35048*/;
  assign _3357_ = ~q[17] /*35047*/;
  assign _3358_ = sum_15[31] & q[17] /*35046*/;
  assign _3359_ = m_15[31] & _3357_ /*35045*/;
  assign r_15[48] = _3359_ | _3358_ /*35044*/;
assign r_15[0]= r_14[0] /*35043*/;
assign r_15[1]= r_14[1] /*35042*/;
assign r_15[2]= r_14[2] /*35041*/;
assign r_15[3]= r_14[3] /*35040*/;
assign r_15[4]= r_14[4] /*35039*/;
assign r_15[5]= r_14[5] /*35038*/;
assign r_15[6]= r_14[6] /*35037*/;
assign r_15[7]= r_14[7] /*35036*/;
assign r_15[8]= r_14[8] /*35035*/;
assign r_15[9]= r_14[9] /*35034*/;
assign r_15[10]= r_14[10] /*35033*/;
assign r_15[11]= r_14[11] /*35032*/;
assign r_15[12]= r_14[12] /*35031*/;
assign r_15[13]= r_14[13] /*35030*/;
assign r_15[14]= r_14[14] /*35029*/;
assign r_15[15]= r_14[15] /*35028*/;
assign r_15[16]= r_14[16] /*35027*/;
  assign inv_16[0] = ~div[0] /*34952*/;
  assign inv_16[1] = ~div[1] /*34951*/;
  assign inv_16[2] = ~div[2] /*34950*/;
  assign inv_16[3] = ~div[3] /*34949*/;
  assign inv_16[4] = ~div[4] /*34948*/;
  assign inv_16[5] = ~div[5] /*34947*/;
  assign inv_16[6] = ~div[6] /*34946*/;
  assign inv_16[7] = ~div[7] /*34945*/;
  assign inv_16[8] = ~div[8] /*34944*/;
  assign inv_16[9] = ~div[9] /*34943*/;
  assign inv_16[10] = ~div[10] /*34942*/;
  assign inv_16[11] = ~div[11] /*34941*/;
  assign inv_16[12] = ~div[12] /*34940*/;
  assign inv_16[13] = ~div[13] /*34939*/;
  assign inv_16[14] = ~div[14] /*34938*/;
  assign inv_16[15] = ~div[15] /*34937*/;
  assign inv_16[16] = ~div[16] /*34936*/;
  assign inv_16[17] = ~div[17] /*34935*/;
  assign inv_16[18] = ~div[18] /*34934*/;
  assign inv_16[19] = ~div[19] /*34933*/;
  assign inv_16[20] = ~div[20] /*34932*/;
  assign inv_16[21] = ~div[21] /*34931*/;
  assign inv_16[22] = ~div[22] /*34930*/;
  assign inv_16[23] = ~div[23] /*34929*/;
  assign inv_16[24] = ~div[24] /*34928*/;
  assign inv_16[25] = ~div[25] /*34927*/;
  assign inv_16[26] = ~div[26] /*34926*/;
  assign inv_16[27] = ~div[27] /*34925*/;
  assign inv_16[28] = ~div[28] /*34924*/;
  assign inv_16[29] = ~div[29] /*34923*/;
  assign inv_16[30] = ~div[30] /*34922*/;
assign inv_16[31] = oneWire /*34921*/;
  assign _3360_ = inv_16[0] ^ r_15[16] /*34919*/;
  assign sum_16[0] = _3360_ ^ oneWire /*34918*/;
  assign _3361_ = _3360_ & oneWire /*34917*/;
  assign _3362_ = inv_16[0] & r_15[16] /*34916*/;
  assign _3363_ = _3361_ | _3362_ /*34915*/;
  assign _3364_ = inv_16[1] ^ r_15[17] /*34914*/;
  assign sum_16[1] = _3364_ ^ _3363_ /*34913*/;
  assign _3365_ = _3364_ & _3363_ /*34912*/;
  assign _3366_ = inv_16[1] & r_15[17] /*34911*/;
  assign _3367_ = _3365_ | _3366_ /*34910*/;
  assign _3368_ = inv_16[2] ^ r_15[18] /*34908*/;
  assign sum_16[2] = _3368_ ^ _3367_ /*34907*/;
  assign _3369_ = _3368_ & _3367_ /*34906*/;
  assign _3370_ = inv_16[2] & r_15[18] /*34905*/;
  assign _3371_ = _3369_ | _3370_ /*34904*/;
  assign _3372_ = inv_16[3] ^ r_15[19] /*34902*/;
  assign sum_16[3] = _3372_ ^ _3371_ /*34901*/;
  assign _3373_ = _3372_ & _3371_ /*34900*/;
  assign _3374_ = inv_16[3] & r_15[19] /*34899*/;
  assign _3375_ = _3373_ | _3374_ /*34898*/;
  assign _3376_ = inv_16[4] ^ r_15[20] /*34896*/;
  assign sum_16[4] = _3376_ ^ _3375_ /*34895*/;
  assign _3377_ = _3376_ & _3375_ /*34894*/;
  assign _3378_ = inv_16[4] & r_15[20] /*34893*/;
  assign _3379_ = _3377_ | _3378_ /*34892*/;
  assign _3380_ = inv_16[5] ^ r_15[21] /*34890*/;
  assign sum_16[5] = _3380_ ^ _3379_ /*34889*/;
  assign _3381_ = _3380_ & _3379_ /*34888*/;
  assign _3382_ = inv_16[5] & r_15[21] /*34887*/;
  assign _3383_ = _3381_ | _3382_ /*34886*/;
  assign _3384_ = inv_16[6] ^ r_15[22] /*34884*/;
  assign sum_16[6] = _3384_ ^ _3383_ /*34883*/;
  assign _3385_ = _3384_ & _3383_ /*34882*/;
  assign _3386_ = inv_16[6] & r_15[22] /*34881*/;
  assign _3387_ = _3385_ | _3386_ /*34880*/;
  assign _3388_ = inv_16[7] ^ r_15[23] /*34878*/;
  assign sum_16[7] = _3388_ ^ _3387_ /*34877*/;
  assign _3389_ = _3388_ & _3387_ /*34876*/;
  assign _3390_ = inv_16[7] & r_15[23] /*34875*/;
  assign _3391_ = _3389_ | _3390_ /*34874*/;
  assign _3392_ = inv_16[8] ^ r_15[24] /*34872*/;
  assign sum_16[8] = _3392_ ^ _3391_ /*34871*/;
  assign _3393_ = _3392_ & _3391_ /*34870*/;
  assign _3394_ = inv_16[8] & r_15[24] /*34869*/;
  assign _3395_ = _3393_ | _3394_ /*34868*/;
  assign _3396_ = inv_16[9] ^ r_15[25] /*34866*/;
  assign sum_16[9] = _3396_ ^ _3395_ /*34865*/;
  assign _3397_ = _3396_ & _3395_ /*34864*/;
  assign _3398_ = inv_16[9] & r_15[25] /*34863*/;
  assign _3399_ = _3397_ | _3398_ /*34862*/;
  assign _3400_ = inv_16[10] ^ r_15[26] /*34860*/;
  assign sum_16[10] = _3400_ ^ _3399_ /*34859*/;
  assign _3401_ = _3400_ & _3399_ /*34858*/;
  assign _3402_ = inv_16[10] & r_15[26] /*34857*/;
  assign _3403_ = _3401_ | _3402_ /*34856*/;
  assign _3404_ = inv_16[11] ^ r_15[27] /*34854*/;
  assign sum_16[11] = _3404_ ^ _3403_ /*34853*/;
  assign _3405_ = _3404_ & _3403_ /*34852*/;
  assign _3406_ = inv_16[11] & r_15[27] /*34851*/;
  assign _3407_ = _3405_ | _3406_ /*34850*/;
  assign _3408_ = inv_16[12] ^ r_15[28] /*34848*/;
  assign sum_16[12] = _3408_ ^ _3407_ /*34847*/;
  assign _3409_ = _3408_ & _3407_ /*34846*/;
  assign _3410_ = inv_16[12] & r_15[28] /*34845*/;
  assign _3411_ = _3409_ | _3410_ /*34844*/;
  assign _3412_ = inv_16[13] ^ r_15[29] /*34842*/;
  assign sum_16[13] = _3412_ ^ _3411_ /*34841*/;
  assign _3413_ = _3412_ & _3411_ /*34840*/;
  assign _3414_ = inv_16[13] & r_15[29] /*34839*/;
  assign _3415_ = _3413_ | _3414_ /*34838*/;
  assign _3416_ = inv_16[14] ^ r_15[30] /*34836*/;
  assign sum_16[14] = _3416_ ^ _3415_ /*34835*/;
  assign _3417_ = _3416_ & _3415_ /*34834*/;
  assign _3418_ = inv_16[14] & r_15[30] /*34833*/;
  assign _3419_ = _3417_ | _3418_ /*34832*/;
  assign _3420_ = inv_16[15] ^ r_15[31] /*34830*/;
  assign sum_16[15] = _3420_ ^ _3419_ /*34829*/;
  assign _3421_ = _3420_ & _3419_ /*34828*/;
  assign _3422_ = inv_16[15] & r_15[31] /*34827*/;
  assign _3423_ = _3421_ | _3422_ /*34826*/;
  assign _3424_ = inv_16[16] ^ r_15[32] /*34824*/;
  assign sum_16[16] = _3424_ ^ _3423_ /*34823*/;
  assign _3425_ = _3424_ & _3423_ /*34822*/;
  assign _3426_ = inv_16[16] & r_15[32] /*34821*/;
  assign _3427_ = _3425_ | _3426_ /*34820*/;
  assign _3428_ = inv_16[17] ^ r_15[33] /*34818*/;
  assign sum_16[17] = _3428_ ^ _3427_ /*34817*/;
  assign _3429_ = _3428_ & _3427_ /*34816*/;
  assign _3430_ = inv_16[17] & r_15[33] /*34815*/;
  assign _3431_ = _3429_ | _3430_ /*34814*/;
  assign _3432_ = inv_16[18] ^ r_15[34] /*34812*/;
  assign sum_16[18] = _3432_ ^ _3431_ /*34811*/;
  assign _3433_ = _3432_ & _3431_ /*34810*/;
  assign _3434_ = inv_16[18] & r_15[34] /*34809*/;
  assign _3435_ = _3433_ | _3434_ /*34808*/;
  assign _3436_ = inv_16[19] ^ r_15[35] /*34806*/;
  assign sum_16[19] = _3436_ ^ _3435_ /*34805*/;
  assign _3437_ = _3436_ & _3435_ /*34804*/;
  assign _3438_ = inv_16[19] & r_15[35] /*34803*/;
  assign _3439_ = _3437_ | _3438_ /*34802*/;
  assign _3440_ = inv_16[20] ^ r_15[36] /*34800*/;
  assign sum_16[20] = _3440_ ^ _3439_ /*34799*/;
  assign _3441_ = _3440_ & _3439_ /*34798*/;
  assign _3442_ = inv_16[20] & r_15[36] /*34797*/;
  assign _3443_ = _3441_ | _3442_ /*34796*/;
  assign _3444_ = inv_16[21] ^ r_15[37] /*34794*/;
  assign sum_16[21] = _3444_ ^ _3443_ /*34793*/;
  assign _3445_ = _3444_ & _3443_ /*34792*/;
  assign _3446_ = inv_16[21] & r_15[37] /*34791*/;
  assign _3447_ = _3445_ | _3446_ /*34790*/;
  assign _3448_ = inv_16[22] ^ r_15[38] /*34788*/;
  assign sum_16[22] = _3448_ ^ _3447_ /*34787*/;
  assign _3449_ = _3448_ & _3447_ /*34786*/;
  assign _3450_ = inv_16[22] & r_15[38] /*34785*/;
  assign _3451_ = _3449_ | _3450_ /*34784*/;
  assign _3452_ = inv_16[23] ^ r_15[39] /*34782*/;
  assign sum_16[23] = _3452_ ^ _3451_ /*34781*/;
  assign _3453_ = _3452_ & _3451_ /*34780*/;
  assign _3454_ = inv_16[23] & r_15[39] /*34779*/;
  assign _3455_ = _3453_ | _3454_ /*34778*/;
  assign _3456_ = inv_16[24] ^ r_15[40] /*34776*/;
  assign sum_16[24] = _3456_ ^ _3455_ /*34775*/;
  assign _3457_ = _3456_ & _3455_ /*34774*/;
  assign _3458_ = inv_16[24] & r_15[40] /*34773*/;
  assign _3459_ = _3457_ | _3458_ /*34772*/;
  assign _3460_ = inv_16[25] ^ r_15[41] /*34770*/;
  assign sum_16[25] = _3460_ ^ _3459_ /*34769*/;
  assign _3461_ = _3460_ & _3459_ /*34768*/;
  assign _3462_ = inv_16[25] & r_15[41] /*34767*/;
  assign _3463_ = _3461_ | _3462_ /*34766*/;
  assign _3464_ = inv_16[26] ^ r_15[42] /*34764*/;
  assign sum_16[26] = _3464_ ^ _3463_ /*34763*/;
  assign _3465_ = _3464_ & _3463_ /*34762*/;
  assign _3466_ = inv_16[26] & r_15[42] /*34761*/;
  assign _3467_ = _3465_ | _3466_ /*34760*/;
  assign _3468_ = inv_16[27] ^ r_15[43] /*34758*/;
  assign sum_16[27] = _3468_ ^ _3467_ /*34757*/;
  assign _3469_ = _3468_ & _3467_ /*34756*/;
  assign _3470_ = inv_16[27] & r_15[43] /*34755*/;
  assign _3471_ = _3469_ | _3470_ /*34754*/;
  assign _3472_ = inv_16[28] ^ r_15[44] /*34752*/;
  assign sum_16[28] = _3472_ ^ _3471_ /*34751*/;
  assign _3473_ = _3472_ & _3471_ /*34750*/;
  assign _3474_ = inv_16[28] & r_15[44] /*34749*/;
  assign _3475_ = _3473_ | _3474_ /*34748*/;
  assign _3476_ = inv_16[29] ^ r_15[45] /*34746*/;
  assign sum_16[29] = _3476_ ^ _3475_ /*34745*/;
  assign _3477_ = _3476_ & _3475_ /*34744*/;
  assign _3478_ = inv_16[29] & r_15[45] /*34743*/;
  assign _3479_ = _3477_ | _3478_ /*34742*/;
  assign _3480_ = inv_16[30] ^ r_15[46] /*34740*/;
  assign sum_16[30] = _3480_ ^ _3479_ /*34739*/;
  assign _3481_ = _3480_ & _3479_ /*34738*/;
  assign _3482_ = inv_16[30] & r_15[46] /*34737*/;
  assign _3483_ = _3481_ | _3482_ /*34736*/;
  assign _3484_ = inv_16[31] ^ r_15[47] /*34734*/;
  assign sum_16[31] = _3484_ ^ _3483_ /*34733*/;
  assign _3485_ = _3484_ & _3483_ /*34732*/;
  assign _3486_ = inv_16[31] & r_15[47] /*34731*/;
  assign _3487_ = _3485_ | _3486_ /*34730*/;
  assign q[16] = ~sum_16[31] /*34757*/;
  assign m_16[0] = r_15[16] /*34756*/;
  assign m_16[1] = r_15[17] /*34755*/;
  assign m_16[2] = r_15[18] /*34754*/;
  assign m_16[3] = r_15[19] /*34753*/;
  assign m_16[4] = r_15[20] /*34752*/;
  assign m_16[5] = r_15[21] /*34751*/;
  assign m_16[6] = r_15[22] /*34750*/;
  assign m_16[7] = r_15[23] /*34749*/;
  assign m_16[8] = r_15[24] /*34748*/;
  assign m_16[9] = r_15[25] /*34747*/;
  assign m_16[10] = r_15[26] /*34746*/;
  assign m_16[11] = r_15[27] /*34745*/;
  assign m_16[12] = r_15[28] /*34744*/;
  assign m_16[13] = r_15[29] /*34743*/;
  assign m_16[14] = r_15[30] /*34742*/;
  assign m_16[15] = r_15[31] /*34741*/;
  assign m_16[16] = r_15[32] /*34740*/;
  assign m_16[17] = r_15[33] /*34739*/;
  assign m_16[18] = r_15[34] /*34738*/;
  assign m_16[19] = r_15[35] /*34737*/;
  assign m_16[20] = r_15[36] /*34736*/;
  assign m_16[21] = r_15[37] /*34735*/;
  assign m_16[22] = r_15[38] /*34734*/;
  assign m_16[23] = r_15[39] /*34733*/;
  assign m_16[24] = r_15[40] /*34732*/;
  assign m_16[25] = r_15[41] /*34731*/;
  assign m_16[26] = r_15[42] /*34730*/;
  assign m_16[27] = r_15[43] /*34729*/;
  assign m_16[28] = r_15[44] /*34728*/;
  assign m_16[29] = r_15[45] /*34727*/;
  assign m_16[30] = r_15[46] /*34726*/;
  assign m_16[31] = r_15[47] /*34725*/;
  assign _3488_ = ~q[16] /*34723*/;
  assign _3489_ = sum_16[0] & q[16] /*34722*/;
  assign _3490_ = m_16[0] & _3488_ /*34721*/;
  assign r_16[16] = _3490_ | _3489_ /*34720*/;
  assign _3491_ = ~q[16] /*34719*/;
  assign _3492_ = sum_16[1] & q[16] /*34718*/;
  assign _3493_ = m_16[1] & _3491_ /*34717*/;
  assign r_16[17] = _3493_ | _3492_ /*34716*/;
  assign _3494_ = ~q[16] /*34715*/;
  assign _3495_ = sum_16[2] & q[16] /*34714*/;
  assign _3496_ = m_16[2] & _3494_ /*34713*/;
  assign r_16[18] = _3496_ | _3495_ /*34712*/;
  assign _3497_ = ~q[16] /*34711*/;
  assign _3498_ = sum_16[3] & q[16] /*34710*/;
  assign _3499_ = m_16[3] & _3497_ /*34709*/;
  assign r_16[19] = _3499_ | _3498_ /*34708*/;
  assign _3500_ = ~q[16] /*34707*/;
  assign _3501_ = sum_16[4] & q[16] /*34706*/;
  assign _3502_ = m_16[4] & _3500_ /*34705*/;
  assign r_16[20] = _3502_ | _3501_ /*34704*/;
  assign _3503_ = ~q[16] /*34703*/;
  assign _3504_ = sum_16[5] & q[16] /*34702*/;
  assign _3505_ = m_16[5] & _3503_ /*34701*/;
  assign r_16[21] = _3505_ | _3504_ /*34700*/;
  assign _3506_ = ~q[16] /*34699*/;
  assign _3507_ = sum_16[6] & q[16] /*34698*/;
  assign _3508_ = m_16[6] & _3506_ /*34697*/;
  assign r_16[22] = _3508_ | _3507_ /*34696*/;
  assign _3509_ = ~q[16] /*34695*/;
  assign _3510_ = sum_16[7] & q[16] /*34694*/;
  assign _3511_ = m_16[7] & _3509_ /*34693*/;
  assign r_16[23] = _3511_ | _3510_ /*34692*/;
  assign _3512_ = ~q[16] /*34691*/;
  assign _3513_ = sum_16[8] & q[16] /*34690*/;
  assign _3514_ = m_16[8] & _3512_ /*34689*/;
  assign r_16[24] = _3514_ | _3513_ /*34688*/;
  assign _3515_ = ~q[16] /*34687*/;
  assign _3516_ = sum_16[9] & q[16] /*34686*/;
  assign _3517_ = m_16[9] & _3515_ /*34685*/;
  assign r_16[25] = _3517_ | _3516_ /*34684*/;
  assign _3518_ = ~q[16] /*34683*/;
  assign _3519_ = sum_16[10] & q[16] /*34682*/;
  assign _3520_ = m_16[10] & _3518_ /*34681*/;
  assign r_16[26] = _3520_ | _3519_ /*34680*/;
  assign _3521_ = ~q[16] /*34679*/;
  assign _3522_ = sum_16[11] & q[16] /*34678*/;
  assign _3523_ = m_16[11] & _3521_ /*34677*/;
  assign r_16[27] = _3523_ | _3522_ /*34676*/;
  assign _3524_ = ~q[16] /*34675*/;
  assign _3525_ = sum_16[12] & q[16] /*34674*/;
  assign _3526_ = m_16[12] & _3524_ /*34673*/;
  assign r_16[28] = _3526_ | _3525_ /*34672*/;
  assign _3527_ = ~q[16] /*34671*/;
  assign _3528_ = sum_16[13] & q[16] /*34670*/;
  assign _3529_ = m_16[13] & _3527_ /*34669*/;
  assign r_16[29] = _3529_ | _3528_ /*34668*/;
  assign _3530_ = ~q[16] /*34667*/;
  assign _3531_ = sum_16[14] & q[16] /*34666*/;
  assign _3532_ = m_16[14] & _3530_ /*34665*/;
  assign r_16[30] = _3532_ | _3531_ /*34664*/;
  assign _3533_ = ~q[16] /*34663*/;
  assign _3534_ = sum_16[15] & q[16] /*34662*/;
  assign _3535_ = m_16[15] & _3533_ /*34661*/;
  assign r_16[31] = _3535_ | _3534_ /*34660*/;
  assign _3536_ = ~q[16] /*34659*/;
  assign _3537_ = sum_16[16] & q[16] /*34658*/;
  assign _3538_ = m_16[16] & _3536_ /*34657*/;
  assign r_16[32] = _3538_ | _3537_ /*34656*/;
  assign _3539_ = ~q[16] /*34655*/;
  assign _3540_ = sum_16[17] & q[16] /*34654*/;
  assign _3541_ = m_16[17] & _3539_ /*34653*/;
  assign r_16[33] = _3541_ | _3540_ /*34652*/;
  assign _3542_ = ~q[16] /*34651*/;
  assign _3543_ = sum_16[18] & q[16] /*34650*/;
  assign _3544_ = m_16[18] & _3542_ /*34649*/;
  assign r_16[34] = _3544_ | _3543_ /*34648*/;
  assign _3545_ = ~q[16] /*34647*/;
  assign _3546_ = sum_16[19] & q[16] /*34646*/;
  assign _3547_ = m_16[19] & _3545_ /*34645*/;
  assign r_16[35] = _3547_ | _3546_ /*34644*/;
  assign _3548_ = ~q[16] /*34643*/;
  assign _3549_ = sum_16[20] & q[16] /*34642*/;
  assign _3550_ = m_16[20] & _3548_ /*34641*/;
  assign r_16[36] = _3550_ | _3549_ /*34640*/;
  assign _3551_ = ~q[16] /*34639*/;
  assign _3552_ = sum_16[21] & q[16] /*34638*/;
  assign _3553_ = m_16[21] & _3551_ /*34637*/;
  assign r_16[37] = _3553_ | _3552_ /*34636*/;
  assign _3554_ = ~q[16] /*34635*/;
  assign _3555_ = sum_16[22] & q[16] /*34634*/;
  assign _3556_ = m_16[22] & _3554_ /*34633*/;
  assign r_16[38] = _3556_ | _3555_ /*34632*/;
  assign _3557_ = ~q[16] /*34631*/;
  assign _3558_ = sum_16[23] & q[16] /*34630*/;
  assign _3559_ = m_16[23] & _3557_ /*34629*/;
  assign r_16[39] = _3559_ | _3558_ /*34628*/;
  assign _3560_ = ~q[16] /*34627*/;
  assign _3561_ = sum_16[24] & q[16] /*34626*/;
  assign _3562_ = m_16[24] & _3560_ /*34625*/;
  assign r_16[40] = _3562_ | _3561_ /*34624*/;
  assign _3563_ = ~q[16] /*34623*/;
  assign _3564_ = sum_16[25] & q[16] /*34622*/;
  assign _3565_ = m_16[25] & _3563_ /*34621*/;
  assign r_16[41] = _3565_ | _3564_ /*34620*/;
  assign _3566_ = ~q[16] /*34619*/;
  assign _3567_ = sum_16[26] & q[16] /*34618*/;
  assign _3568_ = m_16[26] & _3566_ /*34617*/;
  assign r_16[42] = _3568_ | _3567_ /*34616*/;
  assign _3569_ = ~q[16] /*34615*/;
  assign _3570_ = sum_16[27] & q[16] /*34614*/;
  assign _3571_ = m_16[27] & _3569_ /*34613*/;
  assign r_16[43] = _3571_ | _3570_ /*34612*/;
  assign _3572_ = ~q[16] /*34611*/;
  assign _3573_ = sum_16[28] & q[16] /*34610*/;
  assign _3574_ = m_16[28] & _3572_ /*34609*/;
  assign r_16[44] = _3574_ | _3573_ /*34608*/;
  assign _3575_ = ~q[16] /*34607*/;
  assign _3576_ = sum_16[29] & q[16] /*34606*/;
  assign _3577_ = m_16[29] & _3575_ /*34605*/;
  assign r_16[45] = _3577_ | _3576_ /*34604*/;
  assign _3578_ = ~q[16] /*34603*/;
  assign _3579_ = sum_16[30] & q[16] /*34602*/;
  assign _3580_ = m_16[30] & _3578_ /*34601*/;
  assign r_16[46] = _3580_ | _3579_ /*34600*/;
  assign _3581_ = ~q[16] /*34599*/;
  assign _3582_ = sum_16[31] & q[16] /*34598*/;
  assign _3583_ = m_16[31] & _3581_ /*34597*/;
  assign r_16[47] = _3583_ | _3582_ /*34596*/;
assign r_16[0]= r_15[0] /*34595*/;
assign r_16[1]= r_15[1] /*34594*/;
assign r_16[2]= r_15[2] /*34593*/;
assign r_16[3]= r_15[3] /*34592*/;
assign r_16[4]= r_15[4] /*34591*/;
assign r_16[5]= r_15[5] /*34590*/;
assign r_16[6]= r_15[6] /*34589*/;
assign r_16[7]= r_15[7] /*34588*/;
assign r_16[8]= r_15[8] /*34587*/;
assign r_16[9]= r_15[9] /*34586*/;
assign r_16[10]= r_15[10] /*34585*/;
assign r_16[11]= r_15[11] /*34584*/;
assign r_16[12]= r_15[12] /*34583*/;
assign r_16[13]= r_15[13] /*34582*/;
assign r_16[14]= r_15[14] /*34581*/;
assign r_16[15]= r_15[15] /*34580*/;
  assign inv_17[0] = ~div[0] /*34504*/;
  assign inv_17[1] = ~div[1] /*34503*/;
  assign inv_17[2] = ~div[2] /*34502*/;
  assign inv_17[3] = ~div[3] /*34501*/;
  assign inv_17[4] = ~div[4] /*34500*/;
  assign inv_17[5] = ~div[5] /*34499*/;
  assign inv_17[6] = ~div[6] /*34498*/;
  assign inv_17[7] = ~div[7] /*34497*/;
  assign inv_17[8] = ~div[8] /*34496*/;
  assign inv_17[9] = ~div[9] /*34495*/;
  assign inv_17[10] = ~div[10] /*34494*/;
  assign inv_17[11] = ~div[11] /*34493*/;
  assign inv_17[12] = ~div[12] /*34492*/;
  assign inv_17[13] = ~div[13] /*34491*/;
  assign inv_17[14] = ~div[14] /*34490*/;
  assign inv_17[15] = ~div[15] /*34489*/;
  assign inv_17[16] = ~div[16] /*34488*/;
  assign inv_17[17] = ~div[17] /*34487*/;
  assign inv_17[18] = ~div[18] /*34486*/;
  assign inv_17[19] = ~div[19] /*34485*/;
  assign inv_17[20] = ~div[20] /*34484*/;
  assign inv_17[21] = ~div[21] /*34483*/;
  assign inv_17[22] = ~div[22] /*34482*/;
  assign inv_17[23] = ~div[23] /*34481*/;
  assign inv_17[24] = ~div[24] /*34480*/;
  assign inv_17[25] = ~div[25] /*34479*/;
  assign inv_17[26] = ~div[26] /*34478*/;
  assign inv_17[27] = ~div[27] /*34477*/;
  assign inv_17[28] = ~div[28] /*34476*/;
  assign inv_17[29] = ~div[29] /*34475*/;
  assign inv_17[30] = ~div[30] /*34474*/;
assign inv_17[31] = oneWire /*34473*/;
  assign _3584_ = inv_17[0] ^ r_16[15] /*34471*/;
  assign sum_17[0] = _3584_ ^ oneWire /*34470*/;
  assign _3585_ = _3584_ & oneWire /*34469*/;
  assign _3586_ = inv_17[0] & r_16[15] /*34468*/;
  assign _3587_ = _3585_ | _3586_ /*34467*/;
  assign _3588_ = inv_17[1] ^ r_16[16] /*34466*/;
  assign sum_17[1] = _3588_ ^ _3587_ /*34465*/;
  assign _3589_ = _3588_ & _3587_ /*34464*/;
  assign _3590_ = inv_17[1] & r_16[16] /*34463*/;
  assign _3591_ = _3589_ | _3590_ /*34462*/;
  assign _3592_ = inv_17[2] ^ r_16[17] /*34460*/;
  assign sum_17[2] = _3592_ ^ _3591_ /*34459*/;
  assign _3593_ = _3592_ & _3591_ /*34458*/;
  assign _3594_ = inv_17[2] & r_16[17] /*34457*/;
  assign _3595_ = _3593_ | _3594_ /*34456*/;
  assign _3596_ = inv_17[3] ^ r_16[18] /*34454*/;
  assign sum_17[3] = _3596_ ^ _3595_ /*34453*/;
  assign _3597_ = _3596_ & _3595_ /*34452*/;
  assign _3598_ = inv_17[3] & r_16[18] /*34451*/;
  assign _3599_ = _3597_ | _3598_ /*34450*/;
  assign _3600_ = inv_17[4] ^ r_16[19] /*34448*/;
  assign sum_17[4] = _3600_ ^ _3599_ /*34447*/;
  assign _3601_ = _3600_ & _3599_ /*34446*/;
  assign _3602_ = inv_17[4] & r_16[19] /*34445*/;
  assign _3603_ = _3601_ | _3602_ /*34444*/;
  assign _3604_ = inv_17[5] ^ r_16[20] /*34442*/;
  assign sum_17[5] = _3604_ ^ _3603_ /*34441*/;
  assign _3605_ = _3604_ & _3603_ /*34440*/;
  assign _3606_ = inv_17[5] & r_16[20] /*34439*/;
  assign _3607_ = _3605_ | _3606_ /*34438*/;
  assign _3608_ = inv_17[6] ^ r_16[21] /*34436*/;
  assign sum_17[6] = _3608_ ^ _3607_ /*34435*/;
  assign _3609_ = _3608_ & _3607_ /*34434*/;
  assign _3610_ = inv_17[6] & r_16[21] /*34433*/;
  assign _3611_ = _3609_ | _3610_ /*34432*/;
  assign _3612_ = inv_17[7] ^ r_16[22] /*34430*/;
  assign sum_17[7] = _3612_ ^ _3611_ /*34429*/;
  assign _3613_ = _3612_ & _3611_ /*34428*/;
  assign _3614_ = inv_17[7] & r_16[22] /*34427*/;
  assign _3615_ = _3613_ | _3614_ /*34426*/;
  assign _3616_ = inv_17[8] ^ r_16[23] /*34424*/;
  assign sum_17[8] = _3616_ ^ _3615_ /*34423*/;
  assign _3617_ = _3616_ & _3615_ /*34422*/;
  assign _3618_ = inv_17[8] & r_16[23] /*34421*/;
  assign _3619_ = _3617_ | _3618_ /*34420*/;
  assign _3620_ = inv_17[9] ^ r_16[24] /*34418*/;
  assign sum_17[9] = _3620_ ^ _3619_ /*34417*/;
  assign _3621_ = _3620_ & _3619_ /*34416*/;
  assign _3622_ = inv_17[9] & r_16[24] /*34415*/;
  assign _3623_ = _3621_ | _3622_ /*34414*/;
  assign _3624_ = inv_17[10] ^ r_16[25] /*34412*/;
  assign sum_17[10] = _3624_ ^ _3623_ /*34411*/;
  assign _3625_ = _3624_ & _3623_ /*34410*/;
  assign _3626_ = inv_17[10] & r_16[25] /*34409*/;
  assign _3627_ = _3625_ | _3626_ /*34408*/;
  assign _3628_ = inv_17[11] ^ r_16[26] /*34406*/;
  assign sum_17[11] = _3628_ ^ _3627_ /*34405*/;
  assign _3629_ = _3628_ & _3627_ /*34404*/;
  assign _3630_ = inv_17[11] & r_16[26] /*34403*/;
  assign _3631_ = _3629_ | _3630_ /*34402*/;
  assign _3632_ = inv_17[12] ^ r_16[27] /*34400*/;
  assign sum_17[12] = _3632_ ^ _3631_ /*34399*/;
  assign _3633_ = _3632_ & _3631_ /*34398*/;
  assign _3634_ = inv_17[12] & r_16[27] /*34397*/;
  assign _3635_ = _3633_ | _3634_ /*34396*/;
  assign _3636_ = inv_17[13] ^ r_16[28] /*34394*/;
  assign sum_17[13] = _3636_ ^ _3635_ /*34393*/;
  assign _3637_ = _3636_ & _3635_ /*34392*/;
  assign _3638_ = inv_17[13] & r_16[28] /*34391*/;
  assign _3639_ = _3637_ | _3638_ /*34390*/;
  assign _3640_ = inv_17[14] ^ r_16[29] /*34388*/;
  assign sum_17[14] = _3640_ ^ _3639_ /*34387*/;
  assign _3641_ = _3640_ & _3639_ /*34386*/;
  assign _3642_ = inv_17[14] & r_16[29] /*34385*/;
  assign _3643_ = _3641_ | _3642_ /*34384*/;
  assign _3644_ = inv_17[15] ^ r_16[30] /*34382*/;
  assign sum_17[15] = _3644_ ^ _3643_ /*34381*/;
  assign _3645_ = _3644_ & _3643_ /*34380*/;
  assign _3646_ = inv_17[15] & r_16[30] /*34379*/;
  assign _3647_ = _3645_ | _3646_ /*34378*/;
  assign _3648_ = inv_17[16] ^ r_16[31] /*34376*/;
  assign sum_17[16] = _3648_ ^ _3647_ /*34375*/;
  assign _3649_ = _3648_ & _3647_ /*34374*/;
  assign _3650_ = inv_17[16] & r_16[31] /*34373*/;
  assign _3651_ = _3649_ | _3650_ /*34372*/;
  assign _3652_ = inv_17[17] ^ r_16[32] /*34370*/;
  assign sum_17[17] = _3652_ ^ _3651_ /*34369*/;
  assign _3653_ = _3652_ & _3651_ /*34368*/;
  assign _3654_ = inv_17[17] & r_16[32] /*34367*/;
  assign _3655_ = _3653_ | _3654_ /*34366*/;
  assign _3656_ = inv_17[18] ^ r_16[33] /*34364*/;
  assign sum_17[18] = _3656_ ^ _3655_ /*34363*/;
  assign _3657_ = _3656_ & _3655_ /*34362*/;
  assign _3658_ = inv_17[18] & r_16[33] /*34361*/;
  assign _3659_ = _3657_ | _3658_ /*34360*/;
  assign _3660_ = inv_17[19] ^ r_16[34] /*34358*/;
  assign sum_17[19] = _3660_ ^ _3659_ /*34357*/;
  assign _3661_ = _3660_ & _3659_ /*34356*/;
  assign _3662_ = inv_17[19] & r_16[34] /*34355*/;
  assign _3663_ = _3661_ | _3662_ /*34354*/;
  assign _3664_ = inv_17[20] ^ r_16[35] /*34352*/;
  assign sum_17[20] = _3664_ ^ _3663_ /*34351*/;
  assign _3665_ = _3664_ & _3663_ /*34350*/;
  assign _3666_ = inv_17[20] & r_16[35] /*34349*/;
  assign _3667_ = _3665_ | _3666_ /*34348*/;
  assign _3668_ = inv_17[21] ^ r_16[36] /*34346*/;
  assign sum_17[21] = _3668_ ^ _3667_ /*34345*/;
  assign _3669_ = _3668_ & _3667_ /*34344*/;
  assign _3670_ = inv_17[21] & r_16[36] /*34343*/;
  assign _3671_ = _3669_ | _3670_ /*34342*/;
  assign _3672_ = inv_17[22] ^ r_16[37] /*34340*/;
  assign sum_17[22] = _3672_ ^ _3671_ /*34339*/;
  assign _3673_ = _3672_ & _3671_ /*34338*/;
  assign _3674_ = inv_17[22] & r_16[37] /*34337*/;
  assign _3675_ = _3673_ | _3674_ /*34336*/;
  assign _3676_ = inv_17[23] ^ r_16[38] /*34334*/;
  assign sum_17[23] = _3676_ ^ _3675_ /*34333*/;
  assign _3677_ = _3676_ & _3675_ /*34332*/;
  assign _3678_ = inv_17[23] & r_16[38] /*34331*/;
  assign _3679_ = _3677_ | _3678_ /*34330*/;
  assign _3680_ = inv_17[24] ^ r_16[39] /*34328*/;
  assign sum_17[24] = _3680_ ^ _3679_ /*34327*/;
  assign _3681_ = _3680_ & _3679_ /*34326*/;
  assign _3682_ = inv_17[24] & r_16[39] /*34325*/;
  assign _3683_ = _3681_ | _3682_ /*34324*/;
  assign _3684_ = inv_17[25] ^ r_16[40] /*34322*/;
  assign sum_17[25] = _3684_ ^ _3683_ /*34321*/;
  assign _3685_ = _3684_ & _3683_ /*34320*/;
  assign _3686_ = inv_17[25] & r_16[40] /*34319*/;
  assign _3687_ = _3685_ | _3686_ /*34318*/;
  assign _3688_ = inv_17[26] ^ r_16[41] /*34316*/;
  assign sum_17[26] = _3688_ ^ _3687_ /*34315*/;
  assign _3689_ = _3688_ & _3687_ /*34314*/;
  assign _3690_ = inv_17[26] & r_16[41] /*34313*/;
  assign _3691_ = _3689_ | _3690_ /*34312*/;
  assign _3692_ = inv_17[27] ^ r_16[42] /*34310*/;
  assign sum_17[27] = _3692_ ^ _3691_ /*34309*/;
  assign _3693_ = _3692_ & _3691_ /*34308*/;
  assign _3694_ = inv_17[27] & r_16[42] /*34307*/;
  assign _3695_ = _3693_ | _3694_ /*34306*/;
  assign _3696_ = inv_17[28] ^ r_16[43] /*34304*/;
  assign sum_17[28] = _3696_ ^ _3695_ /*34303*/;
  assign _3697_ = _3696_ & _3695_ /*34302*/;
  assign _3698_ = inv_17[28] & r_16[43] /*34301*/;
  assign _3699_ = _3697_ | _3698_ /*34300*/;
  assign _3700_ = inv_17[29] ^ r_16[44] /*34298*/;
  assign sum_17[29] = _3700_ ^ _3699_ /*34297*/;
  assign _3701_ = _3700_ & _3699_ /*34296*/;
  assign _3702_ = inv_17[29] & r_16[44] /*34295*/;
  assign _3703_ = _3701_ | _3702_ /*34294*/;
  assign _3704_ = inv_17[30] ^ r_16[45] /*34292*/;
  assign sum_17[30] = _3704_ ^ _3703_ /*34291*/;
  assign _3705_ = _3704_ & _3703_ /*34290*/;
  assign _3706_ = inv_17[30] & r_16[45] /*34289*/;
  assign _3707_ = _3705_ | _3706_ /*34288*/;
  assign _3708_ = inv_17[31] ^ r_16[46] /*34286*/;
  assign sum_17[31] = _3708_ ^ _3707_ /*34285*/;
  assign _3709_ = _3708_ & _3707_ /*34284*/;
  assign _3710_ = inv_17[31] & r_16[46] /*34283*/;
  assign _3711_ = _3709_ | _3710_ /*34282*/;
  assign q[15] = ~sum_17[31] /*34309*/;
  assign m_17[0] = r_16[15] /*34308*/;
  assign m_17[1] = r_16[16] /*34307*/;
  assign m_17[2] = r_16[17] /*34306*/;
  assign m_17[3] = r_16[18] /*34305*/;
  assign m_17[4] = r_16[19] /*34304*/;
  assign m_17[5] = r_16[20] /*34303*/;
  assign m_17[6] = r_16[21] /*34302*/;
  assign m_17[7] = r_16[22] /*34301*/;
  assign m_17[8] = r_16[23] /*34300*/;
  assign m_17[9] = r_16[24] /*34299*/;
  assign m_17[10] = r_16[25] /*34298*/;
  assign m_17[11] = r_16[26] /*34297*/;
  assign m_17[12] = r_16[27] /*34296*/;
  assign m_17[13] = r_16[28] /*34295*/;
  assign m_17[14] = r_16[29] /*34294*/;
  assign m_17[15] = r_16[30] /*34293*/;
  assign m_17[16] = r_16[31] /*34292*/;
  assign m_17[17] = r_16[32] /*34291*/;
  assign m_17[18] = r_16[33] /*34290*/;
  assign m_17[19] = r_16[34] /*34289*/;
  assign m_17[20] = r_16[35] /*34288*/;
  assign m_17[21] = r_16[36] /*34287*/;
  assign m_17[22] = r_16[37] /*34286*/;
  assign m_17[23] = r_16[38] /*34285*/;
  assign m_17[24] = r_16[39] /*34284*/;
  assign m_17[25] = r_16[40] /*34283*/;
  assign m_17[26] = r_16[41] /*34282*/;
  assign m_17[27] = r_16[42] /*34281*/;
  assign m_17[28] = r_16[43] /*34280*/;
  assign m_17[29] = r_16[44] /*34279*/;
  assign m_17[30] = r_16[45] /*34278*/;
  assign m_17[31] = r_16[46] /*34277*/;
  assign _3712_ = ~q[15] /*34275*/;
  assign _3713_ = sum_17[0] & q[15] /*34274*/;
  assign _3714_ = m_17[0] & _3712_ /*34273*/;
  assign r_17[15] = _3714_ | _3713_ /*34272*/;
  assign _3715_ = ~q[15] /*34271*/;
  assign _3716_ = sum_17[1] & q[15] /*34270*/;
  assign _3717_ = m_17[1] & _3715_ /*34269*/;
  assign r_17[16] = _3717_ | _3716_ /*34268*/;
  assign _3718_ = ~q[15] /*34267*/;
  assign _3719_ = sum_17[2] & q[15] /*34266*/;
  assign _3720_ = m_17[2] & _3718_ /*34265*/;
  assign r_17[17] = _3720_ | _3719_ /*34264*/;
  assign _3721_ = ~q[15] /*34263*/;
  assign _3722_ = sum_17[3] & q[15] /*34262*/;
  assign _3723_ = m_17[3] & _3721_ /*34261*/;
  assign r_17[18] = _3723_ | _3722_ /*34260*/;
  assign _3724_ = ~q[15] /*34259*/;
  assign _3725_ = sum_17[4] & q[15] /*34258*/;
  assign _3726_ = m_17[4] & _3724_ /*34257*/;
  assign r_17[19] = _3726_ | _3725_ /*34256*/;
  assign _3727_ = ~q[15] /*34255*/;
  assign _3728_ = sum_17[5] & q[15] /*34254*/;
  assign _3729_ = m_17[5] & _3727_ /*34253*/;
  assign r_17[20] = _3729_ | _3728_ /*34252*/;
  assign _3730_ = ~q[15] /*34251*/;
  assign _3731_ = sum_17[6] & q[15] /*34250*/;
  assign _3732_ = m_17[6] & _3730_ /*34249*/;
  assign r_17[21] = _3732_ | _3731_ /*34248*/;
  assign _3733_ = ~q[15] /*34247*/;
  assign _3734_ = sum_17[7] & q[15] /*34246*/;
  assign _3735_ = m_17[7] & _3733_ /*34245*/;
  assign r_17[22] = _3735_ | _3734_ /*34244*/;
  assign _3736_ = ~q[15] /*34243*/;
  assign _3737_ = sum_17[8] & q[15] /*34242*/;
  assign _3738_ = m_17[8] & _3736_ /*34241*/;
  assign r_17[23] = _3738_ | _3737_ /*34240*/;
  assign _3739_ = ~q[15] /*34239*/;
  assign _3740_ = sum_17[9] & q[15] /*34238*/;
  assign _3741_ = m_17[9] & _3739_ /*34237*/;
  assign r_17[24] = _3741_ | _3740_ /*34236*/;
  assign _3742_ = ~q[15] /*34235*/;
  assign _3743_ = sum_17[10] & q[15] /*34234*/;
  assign _3744_ = m_17[10] & _3742_ /*34233*/;
  assign r_17[25] = _3744_ | _3743_ /*34232*/;
  assign _3745_ = ~q[15] /*34231*/;
  assign _3746_ = sum_17[11] & q[15] /*34230*/;
  assign _3747_ = m_17[11] & _3745_ /*34229*/;
  assign r_17[26] = _3747_ | _3746_ /*34228*/;
  assign _3748_ = ~q[15] /*34227*/;
  assign _3749_ = sum_17[12] & q[15] /*34226*/;
  assign _3750_ = m_17[12] & _3748_ /*34225*/;
  assign r_17[27] = _3750_ | _3749_ /*34224*/;
  assign _3751_ = ~q[15] /*34223*/;
  assign _3752_ = sum_17[13] & q[15] /*34222*/;
  assign _3753_ = m_17[13] & _3751_ /*34221*/;
  assign r_17[28] = _3753_ | _3752_ /*34220*/;
  assign _3754_ = ~q[15] /*34219*/;
  assign _3755_ = sum_17[14] & q[15] /*34218*/;
  assign _3756_ = m_17[14] & _3754_ /*34217*/;
  assign r_17[29] = _3756_ | _3755_ /*34216*/;
  assign _3757_ = ~q[15] /*34215*/;
  assign _3758_ = sum_17[15] & q[15] /*34214*/;
  assign _3759_ = m_17[15] & _3757_ /*34213*/;
  assign r_17[30] = _3759_ | _3758_ /*34212*/;
  assign _3760_ = ~q[15] /*34211*/;
  assign _3761_ = sum_17[16] & q[15] /*34210*/;
  assign _3762_ = m_17[16] & _3760_ /*34209*/;
  assign r_17[31] = _3762_ | _3761_ /*34208*/;
  assign _3763_ = ~q[15] /*34207*/;
  assign _3764_ = sum_17[17] & q[15] /*34206*/;
  assign _3765_ = m_17[17] & _3763_ /*34205*/;
  assign r_17[32] = _3765_ | _3764_ /*34204*/;
  assign _3766_ = ~q[15] /*34203*/;
  assign _3767_ = sum_17[18] & q[15] /*34202*/;
  assign _3768_ = m_17[18] & _3766_ /*34201*/;
  assign r_17[33] = _3768_ | _3767_ /*34200*/;
  assign _3769_ = ~q[15] /*34199*/;
  assign _3770_ = sum_17[19] & q[15] /*34198*/;
  assign _3771_ = m_17[19] & _3769_ /*34197*/;
  assign r_17[34] = _3771_ | _3770_ /*34196*/;
  assign _3772_ = ~q[15] /*34195*/;
  assign _3773_ = sum_17[20] & q[15] /*34194*/;
  assign _3774_ = m_17[20] & _3772_ /*34193*/;
  assign r_17[35] = _3774_ | _3773_ /*34192*/;
  assign _3775_ = ~q[15] /*34191*/;
  assign _3776_ = sum_17[21] & q[15] /*34190*/;
  assign _3777_ = m_17[21] & _3775_ /*34189*/;
  assign r_17[36] = _3777_ | _3776_ /*34188*/;
  assign _3778_ = ~q[15] /*34187*/;
  assign _3779_ = sum_17[22] & q[15] /*34186*/;
  assign _3780_ = m_17[22] & _3778_ /*34185*/;
  assign r_17[37] = _3780_ | _3779_ /*34184*/;
  assign _3781_ = ~q[15] /*34183*/;
  assign _3782_ = sum_17[23] & q[15] /*34182*/;
  assign _3783_ = m_17[23] & _3781_ /*34181*/;
  assign r_17[38] = _3783_ | _3782_ /*34180*/;
  assign _3784_ = ~q[15] /*34179*/;
  assign _3785_ = sum_17[24] & q[15] /*34178*/;
  assign _3786_ = m_17[24] & _3784_ /*34177*/;
  assign r_17[39] = _3786_ | _3785_ /*34176*/;
  assign _3787_ = ~q[15] /*34175*/;
  assign _3788_ = sum_17[25] & q[15] /*34174*/;
  assign _3789_ = m_17[25] & _3787_ /*34173*/;
  assign r_17[40] = _3789_ | _3788_ /*34172*/;
  assign _3790_ = ~q[15] /*34171*/;
  assign _3791_ = sum_17[26] & q[15] /*34170*/;
  assign _3792_ = m_17[26] & _3790_ /*34169*/;
  assign r_17[41] = _3792_ | _3791_ /*34168*/;
  assign _3793_ = ~q[15] /*34167*/;
  assign _3794_ = sum_17[27] & q[15] /*34166*/;
  assign _3795_ = m_17[27] & _3793_ /*34165*/;
  assign r_17[42] = _3795_ | _3794_ /*34164*/;
  assign _3796_ = ~q[15] /*34163*/;
  assign _3797_ = sum_17[28] & q[15] /*34162*/;
  assign _3798_ = m_17[28] & _3796_ /*34161*/;
  assign r_17[43] = _3798_ | _3797_ /*34160*/;
  assign _3799_ = ~q[15] /*34159*/;
  assign _3800_ = sum_17[29] & q[15] /*34158*/;
  assign _3801_ = m_17[29] & _3799_ /*34157*/;
  assign r_17[44] = _3801_ | _3800_ /*34156*/;
  assign _3802_ = ~q[15] /*34155*/;
  assign _3803_ = sum_17[30] & q[15] /*34154*/;
  assign _3804_ = m_17[30] & _3802_ /*34153*/;
  assign r_17[45] = _3804_ | _3803_ /*34152*/;
  assign _3805_ = ~q[15] /*34151*/;
  assign _3806_ = sum_17[31] & q[15] /*34150*/;
  assign _3807_ = m_17[31] & _3805_ /*34149*/;
  assign r_17[46] = _3807_ | _3806_ /*34148*/;
assign r_17[0]= r_16[0] /*34147*/;
assign r_17[1]= r_16[1] /*34146*/;
assign r_17[2]= r_16[2] /*34145*/;
assign r_17[3]= r_16[3] /*34144*/;
assign r_17[4]= r_16[4] /*34143*/;
assign r_17[5]= r_16[5] /*34142*/;
assign r_17[6]= r_16[6] /*34141*/;
assign r_17[7]= r_16[7] /*34140*/;
assign r_17[8]= r_16[8] /*34139*/;
assign r_17[9]= r_16[9] /*34138*/;
assign r_17[10]= r_16[10] /*34137*/;
assign r_17[11]= r_16[11] /*34136*/;
assign r_17[12]= r_16[12] /*34135*/;
assign r_17[13]= r_16[13] /*34134*/;
assign r_17[14]= r_16[14] /*34133*/;
  assign inv_18[0] = ~div[0] /*34056*/;
  assign inv_18[1] = ~div[1] /*34055*/;
  assign inv_18[2] = ~div[2] /*34054*/;
  assign inv_18[3] = ~div[3] /*34053*/;
  assign inv_18[4] = ~div[4] /*34052*/;
  assign inv_18[5] = ~div[5] /*34051*/;
  assign inv_18[6] = ~div[6] /*34050*/;
  assign inv_18[7] = ~div[7] /*34049*/;
  assign inv_18[8] = ~div[8] /*34048*/;
  assign inv_18[9] = ~div[9] /*34047*/;
  assign inv_18[10] = ~div[10] /*34046*/;
  assign inv_18[11] = ~div[11] /*34045*/;
  assign inv_18[12] = ~div[12] /*34044*/;
  assign inv_18[13] = ~div[13] /*34043*/;
  assign inv_18[14] = ~div[14] /*34042*/;
  assign inv_18[15] = ~div[15] /*34041*/;
  assign inv_18[16] = ~div[16] /*34040*/;
  assign inv_18[17] = ~div[17] /*34039*/;
  assign inv_18[18] = ~div[18] /*34038*/;
  assign inv_18[19] = ~div[19] /*34037*/;
  assign inv_18[20] = ~div[20] /*34036*/;
  assign inv_18[21] = ~div[21] /*34035*/;
  assign inv_18[22] = ~div[22] /*34034*/;
  assign inv_18[23] = ~div[23] /*34033*/;
  assign inv_18[24] = ~div[24] /*34032*/;
  assign inv_18[25] = ~div[25] /*34031*/;
  assign inv_18[26] = ~div[26] /*34030*/;
  assign inv_18[27] = ~div[27] /*34029*/;
  assign inv_18[28] = ~div[28] /*34028*/;
  assign inv_18[29] = ~div[29] /*34027*/;
  assign inv_18[30] = ~div[30] /*34026*/;
assign inv_18[31] = oneWire /*34025*/;
  assign _3808_ = inv_18[0] ^ r_17[14] /*34023*/;
  assign sum_18[0] = _3808_ ^ oneWire /*34022*/;
  assign _3809_ = _3808_ & oneWire /*34021*/;
  assign _3810_ = inv_18[0] & r_17[14] /*34020*/;
  assign _3811_ = _3809_ | _3810_ /*34019*/;
  assign _3812_ = inv_18[1] ^ r_17[15] /*34018*/;
  assign sum_18[1] = _3812_ ^ _3811_ /*34017*/;
  assign _3813_ = _3812_ & _3811_ /*34016*/;
  assign _3814_ = inv_18[1] & r_17[15] /*34015*/;
  assign _3815_ = _3813_ | _3814_ /*34014*/;
  assign _3816_ = inv_18[2] ^ r_17[16] /*34012*/;
  assign sum_18[2] = _3816_ ^ _3815_ /*34011*/;
  assign _3817_ = _3816_ & _3815_ /*34010*/;
  assign _3818_ = inv_18[2] & r_17[16] /*34009*/;
  assign _3819_ = _3817_ | _3818_ /*34008*/;
  assign _3820_ = inv_18[3] ^ r_17[17] /*34006*/;
  assign sum_18[3] = _3820_ ^ _3819_ /*34005*/;
  assign _3821_ = _3820_ & _3819_ /*34004*/;
  assign _3822_ = inv_18[3] & r_17[17] /*34003*/;
  assign _3823_ = _3821_ | _3822_ /*34002*/;
  assign _3824_ = inv_18[4] ^ r_17[18] /*34000*/;
  assign sum_18[4] = _3824_ ^ _3823_ /*33999*/;
  assign _3825_ = _3824_ & _3823_ /*33998*/;
  assign _3826_ = inv_18[4] & r_17[18] /*33997*/;
  assign _3827_ = _3825_ | _3826_ /*33996*/;
  assign _3828_ = inv_18[5] ^ r_17[19] /*33994*/;
  assign sum_18[5] = _3828_ ^ _3827_ /*33993*/;
  assign _3829_ = _3828_ & _3827_ /*33992*/;
  assign _3830_ = inv_18[5] & r_17[19] /*33991*/;
  assign _3831_ = _3829_ | _3830_ /*33990*/;
  assign _3832_ = inv_18[6] ^ r_17[20] /*33988*/;
  assign sum_18[6] = _3832_ ^ _3831_ /*33987*/;
  assign _3833_ = _3832_ & _3831_ /*33986*/;
  assign _3834_ = inv_18[6] & r_17[20] /*33985*/;
  assign _3835_ = _3833_ | _3834_ /*33984*/;
  assign _3836_ = inv_18[7] ^ r_17[21] /*33982*/;
  assign sum_18[7] = _3836_ ^ _3835_ /*33981*/;
  assign _3837_ = _3836_ & _3835_ /*33980*/;
  assign _3838_ = inv_18[7] & r_17[21] /*33979*/;
  assign _3839_ = _3837_ | _3838_ /*33978*/;
  assign _3840_ = inv_18[8] ^ r_17[22] /*33976*/;
  assign sum_18[8] = _3840_ ^ _3839_ /*33975*/;
  assign _3841_ = _3840_ & _3839_ /*33974*/;
  assign _3842_ = inv_18[8] & r_17[22] /*33973*/;
  assign _3843_ = _3841_ | _3842_ /*33972*/;
  assign _3844_ = inv_18[9] ^ r_17[23] /*33970*/;
  assign sum_18[9] = _3844_ ^ _3843_ /*33969*/;
  assign _3845_ = _3844_ & _3843_ /*33968*/;
  assign _3846_ = inv_18[9] & r_17[23] /*33967*/;
  assign _3847_ = _3845_ | _3846_ /*33966*/;
  assign _3848_ = inv_18[10] ^ r_17[24] /*33964*/;
  assign sum_18[10] = _3848_ ^ _3847_ /*33963*/;
  assign _3849_ = _3848_ & _3847_ /*33962*/;
  assign _3850_ = inv_18[10] & r_17[24] /*33961*/;
  assign _3851_ = _3849_ | _3850_ /*33960*/;
  assign _3852_ = inv_18[11] ^ r_17[25] /*33958*/;
  assign sum_18[11] = _3852_ ^ _3851_ /*33957*/;
  assign _3853_ = _3852_ & _3851_ /*33956*/;
  assign _3854_ = inv_18[11] & r_17[25] /*33955*/;
  assign _3855_ = _3853_ | _3854_ /*33954*/;
  assign _3856_ = inv_18[12] ^ r_17[26] /*33952*/;
  assign sum_18[12] = _3856_ ^ _3855_ /*33951*/;
  assign _3857_ = _3856_ & _3855_ /*33950*/;
  assign _3858_ = inv_18[12] & r_17[26] /*33949*/;
  assign _3859_ = _3857_ | _3858_ /*33948*/;
  assign _3860_ = inv_18[13] ^ r_17[27] /*33946*/;
  assign sum_18[13] = _3860_ ^ _3859_ /*33945*/;
  assign _3861_ = _3860_ & _3859_ /*33944*/;
  assign _3862_ = inv_18[13] & r_17[27] /*33943*/;
  assign _3863_ = _3861_ | _3862_ /*33942*/;
  assign _3864_ = inv_18[14] ^ r_17[28] /*33940*/;
  assign sum_18[14] = _3864_ ^ _3863_ /*33939*/;
  assign _3865_ = _3864_ & _3863_ /*33938*/;
  assign _3866_ = inv_18[14] & r_17[28] /*33937*/;
  assign _3867_ = _3865_ | _3866_ /*33936*/;
  assign _3868_ = inv_18[15] ^ r_17[29] /*33934*/;
  assign sum_18[15] = _3868_ ^ _3867_ /*33933*/;
  assign _3869_ = _3868_ & _3867_ /*33932*/;
  assign _3870_ = inv_18[15] & r_17[29] /*33931*/;
  assign _3871_ = _3869_ | _3870_ /*33930*/;
  assign _3872_ = inv_18[16] ^ r_17[30] /*33928*/;
  assign sum_18[16] = _3872_ ^ _3871_ /*33927*/;
  assign _3873_ = _3872_ & _3871_ /*33926*/;
  assign _3874_ = inv_18[16] & r_17[30] /*33925*/;
  assign _3875_ = _3873_ | _3874_ /*33924*/;
  assign _3876_ = inv_18[17] ^ r_17[31] /*33922*/;
  assign sum_18[17] = _3876_ ^ _3875_ /*33921*/;
  assign _3877_ = _3876_ & _3875_ /*33920*/;
  assign _3878_ = inv_18[17] & r_17[31] /*33919*/;
  assign _3879_ = _3877_ | _3878_ /*33918*/;
  assign _3880_ = inv_18[18] ^ r_17[32] /*33916*/;
  assign sum_18[18] = _3880_ ^ _3879_ /*33915*/;
  assign _3881_ = _3880_ & _3879_ /*33914*/;
  assign _3882_ = inv_18[18] & r_17[32] /*33913*/;
  assign _3883_ = _3881_ | _3882_ /*33912*/;
  assign _3884_ = inv_18[19] ^ r_17[33] /*33910*/;
  assign sum_18[19] = _3884_ ^ _3883_ /*33909*/;
  assign _3885_ = _3884_ & _3883_ /*33908*/;
  assign _3886_ = inv_18[19] & r_17[33] /*33907*/;
  assign _3887_ = _3885_ | _3886_ /*33906*/;
  assign _3888_ = inv_18[20] ^ r_17[34] /*33904*/;
  assign sum_18[20] = _3888_ ^ _3887_ /*33903*/;
  assign _3889_ = _3888_ & _3887_ /*33902*/;
  assign _3890_ = inv_18[20] & r_17[34] /*33901*/;
  assign _3891_ = _3889_ | _3890_ /*33900*/;
  assign _3892_ = inv_18[21] ^ r_17[35] /*33898*/;
  assign sum_18[21] = _3892_ ^ _3891_ /*33897*/;
  assign _3893_ = _3892_ & _3891_ /*33896*/;
  assign _3894_ = inv_18[21] & r_17[35] /*33895*/;
  assign _3895_ = _3893_ | _3894_ /*33894*/;
  assign _3896_ = inv_18[22] ^ r_17[36] /*33892*/;
  assign sum_18[22] = _3896_ ^ _3895_ /*33891*/;
  assign _3897_ = _3896_ & _3895_ /*33890*/;
  assign _3898_ = inv_18[22] & r_17[36] /*33889*/;
  assign _3899_ = _3897_ | _3898_ /*33888*/;
  assign _3900_ = inv_18[23] ^ r_17[37] /*33886*/;
  assign sum_18[23] = _3900_ ^ _3899_ /*33885*/;
  assign _3901_ = _3900_ & _3899_ /*33884*/;
  assign _3902_ = inv_18[23] & r_17[37] /*33883*/;
  assign _3903_ = _3901_ | _3902_ /*33882*/;
  assign _3904_ = inv_18[24] ^ r_17[38] /*33880*/;
  assign sum_18[24] = _3904_ ^ _3903_ /*33879*/;
  assign _3905_ = _3904_ & _3903_ /*33878*/;
  assign _3906_ = inv_18[24] & r_17[38] /*33877*/;
  assign _3907_ = _3905_ | _3906_ /*33876*/;
  assign _3908_ = inv_18[25] ^ r_17[39] /*33874*/;
  assign sum_18[25] = _3908_ ^ _3907_ /*33873*/;
  assign _3909_ = _3908_ & _3907_ /*33872*/;
  assign _3910_ = inv_18[25] & r_17[39] /*33871*/;
  assign _3911_ = _3909_ | _3910_ /*33870*/;
  assign _3912_ = inv_18[26] ^ r_17[40] /*33868*/;
  assign sum_18[26] = _3912_ ^ _3911_ /*33867*/;
  assign _3913_ = _3912_ & _3911_ /*33866*/;
  assign _3914_ = inv_18[26] & r_17[40] /*33865*/;
  assign _3915_ = _3913_ | _3914_ /*33864*/;
  assign _3916_ = inv_18[27] ^ r_17[41] /*33862*/;
  assign sum_18[27] = _3916_ ^ _3915_ /*33861*/;
  assign _3917_ = _3916_ & _3915_ /*33860*/;
  assign _3918_ = inv_18[27] & r_17[41] /*33859*/;
  assign _3919_ = _3917_ | _3918_ /*33858*/;
  assign _3920_ = inv_18[28] ^ r_17[42] /*33856*/;
  assign sum_18[28] = _3920_ ^ _3919_ /*33855*/;
  assign _3921_ = _3920_ & _3919_ /*33854*/;
  assign _3922_ = inv_18[28] & r_17[42] /*33853*/;
  assign _3923_ = _3921_ | _3922_ /*33852*/;
  assign _3924_ = inv_18[29] ^ r_17[43] /*33850*/;
  assign sum_18[29] = _3924_ ^ _3923_ /*33849*/;
  assign _3925_ = _3924_ & _3923_ /*33848*/;
  assign _3926_ = inv_18[29] & r_17[43] /*33847*/;
  assign _3927_ = _3925_ | _3926_ /*33846*/;
  assign _3928_ = inv_18[30] ^ r_17[44] /*33844*/;
  assign sum_18[30] = _3928_ ^ _3927_ /*33843*/;
  assign _3929_ = _3928_ & _3927_ /*33842*/;
  assign _3930_ = inv_18[30] & r_17[44] /*33841*/;
  assign _3931_ = _3929_ | _3930_ /*33840*/;
  assign _3932_ = inv_18[31] ^ r_17[45] /*33838*/;
  assign sum_18[31] = _3932_ ^ _3931_ /*33837*/;
  assign _3933_ = _3932_ & _3931_ /*33836*/;
  assign _3934_ = inv_18[31] & r_17[45] /*33835*/;
  assign _3935_ = _3933_ | _3934_ /*33834*/;
  assign q[14] = ~sum_18[31] /*33861*/;
  assign m_18[0] = r_17[14] /*33860*/;
  assign m_18[1] = r_17[15] /*33859*/;
  assign m_18[2] = r_17[16] /*33858*/;
  assign m_18[3] = r_17[17] /*33857*/;
  assign m_18[4] = r_17[18] /*33856*/;
  assign m_18[5] = r_17[19] /*33855*/;
  assign m_18[6] = r_17[20] /*33854*/;
  assign m_18[7] = r_17[21] /*33853*/;
  assign m_18[8] = r_17[22] /*33852*/;
  assign m_18[9] = r_17[23] /*33851*/;
  assign m_18[10] = r_17[24] /*33850*/;
  assign m_18[11] = r_17[25] /*33849*/;
  assign m_18[12] = r_17[26] /*33848*/;
  assign m_18[13] = r_17[27] /*33847*/;
  assign m_18[14] = r_17[28] /*33846*/;
  assign m_18[15] = r_17[29] /*33845*/;
  assign m_18[16] = r_17[30] /*33844*/;
  assign m_18[17] = r_17[31] /*33843*/;
  assign m_18[18] = r_17[32] /*33842*/;
  assign m_18[19] = r_17[33] /*33841*/;
  assign m_18[20] = r_17[34] /*33840*/;
  assign m_18[21] = r_17[35] /*33839*/;
  assign m_18[22] = r_17[36] /*33838*/;
  assign m_18[23] = r_17[37] /*33837*/;
  assign m_18[24] = r_17[38] /*33836*/;
  assign m_18[25] = r_17[39] /*33835*/;
  assign m_18[26] = r_17[40] /*33834*/;
  assign m_18[27] = r_17[41] /*33833*/;
  assign m_18[28] = r_17[42] /*33832*/;
  assign m_18[29] = r_17[43] /*33831*/;
  assign m_18[30] = r_17[44] /*33830*/;
  assign m_18[31] = r_17[45] /*33829*/;
  assign _3936_ = ~q[14] /*33827*/;
  assign _3937_ = sum_18[0] & q[14] /*33826*/;
  assign _3938_ = m_18[0] & _3936_ /*33825*/;
  assign r_18[14] = _3938_ | _3937_ /*33824*/;
  assign _3939_ = ~q[14] /*33823*/;
  assign _3940_ = sum_18[1] & q[14] /*33822*/;
  assign _3941_ = m_18[1] & _3939_ /*33821*/;
  assign r_18[15] = _3941_ | _3940_ /*33820*/;
  assign _3942_ = ~q[14] /*33819*/;
  assign _3943_ = sum_18[2] & q[14] /*33818*/;
  assign _3944_ = m_18[2] & _3942_ /*33817*/;
  assign r_18[16] = _3944_ | _3943_ /*33816*/;
  assign _3945_ = ~q[14] /*33815*/;
  assign _3946_ = sum_18[3] & q[14] /*33814*/;
  assign _3947_ = m_18[3] & _3945_ /*33813*/;
  assign r_18[17] = _3947_ | _3946_ /*33812*/;
  assign _3948_ = ~q[14] /*33811*/;
  assign _3949_ = sum_18[4] & q[14] /*33810*/;
  assign _3950_ = m_18[4] & _3948_ /*33809*/;
  assign r_18[18] = _3950_ | _3949_ /*33808*/;
  assign _3951_ = ~q[14] /*33807*/;
  assign _3952_ = sum_18[5] & q[14] /*33806*/;
  assign _3953_ = m_18[5] & _3951_ /*33805*/;
  assign r_18[19] = _3953_ | _3952_ /*33804*/;
  assign _3954_ = ~q[14] /*33803*/;
  assign _3955_ = sum_18[6] & q[14] /*33802*/;
  assign _3956_ = m_18[6] & _3954_ /*33801*/;
  assign r_18[20] = _3956_ | _3955_ /*33800*/;
  assign _3957_ = ~q[14] /*33799*/;
  assign _3958_ = sum_18[7] & q[14] /*33798*/;
  assign _3959_ = m_18[7] & _3957_ /*33797*/;
  assign r_18[21] = _3959_ | _3958_ /*33796*/;
  assign _3960_ = ~q[14] /*33795*/;
  assign _3961_ = sum_18[8] & q[14] /*33794*/;
  assign _3962_ = m_18[8] & _3960_ /*33793*/;
  assign r_18[22] = _3962_ | _3961_ /*33792*/;
  assign _3963_ = ~q[14] /*33791*/;
  assign _3964_ = sum_18[9] & q[14] /*33790*/;
  assign _3965_ = m_18[9] & _3963_ /*33789*/;
  assign r_18[23] = _3965_ | _3964_ /*33788*/;
  assign _3966_ = ~q[14] /*33787*/;
  assign _3967_ = sum_18[10] & q[14] /*33786*/;
  assign _3968_ = m_18[10] & _3966_ /*33785*/;
  assign r_18[24] = _3968_ | _3967_ /*33784*/;
  assign _3969_ = ~q[14] /*33783*/;
  assign _3970_ = sum_18[11] & q[14] /*33782*/;
  assign _3971_ = m_18[11] & _3969_ /*33781*/;
  assign r_18[25] = _3971_ | _3970_ /*33780*/;
  assign _3972_ = ~q[14] /*33779*/;
  assign _3973_ = sum_18[12] & q[14] /*33778*/;
  assign _3974_ = m_18[12] & _3972_ /*33777*/;
  assign r_18[26] = _3974_ | _3973_ /*33776*/;
  assign _3975_ = ~q[14] /*33775*/;
  assign _3976_ = sum_18[13] & q[14] /*33774*/;
  assign _3977_ = m_18[13] & _3975_ /*33773*/;
  assign r_18[27] = _3977_ | _3976_ /*33772*/;
  assign _3978_ = ~q[14] /*33771*/;
  assign _3979_ = sum_18[14] & q[14] /*33770*/;
  assign _3980_ = m_18[14] & _3978_ /*33769*/;
  assign r_18[28] = _3980_ | _3979_ /*33768*/;
  assign _3981_ = ~q[14] /*33767*/;
  assign _3982_ = sum_18[15] & q[14] /*33766*/;
  assign _3983_ = m_18[15] & _3981_ /*33765*/;
  assign r_18[29] = _3983_ | _3982_ /*33764*/;
  assign _3984_ = ~q[14] /*33763*/;
  assign _3985_ = sum_18[16] & q[14] /*33762*/;
  assign _3986_ = m_18[16] & _3984_ /*33761*/;
  assign r_18[30] = _3986_ | _3985_ /*33760*/;
  assign _3987_ = ~q[14] /*33759*/;
  assign _3988_ = sum_18[17] & q[14] /*33758*/;
  assign _3989_ = m_18[17] & _3987_ /*33757*/;
  assign r_18[31] = _3989_ | _3988_ /*33756*/;
  assign _3990_ = ~q[14] /*33755*/;
  assign _3991_ = sum_18[18] & q[14] /*33754*/;
  assign _3992_ = m_18[18] & _3990_ /*33753*/;
  assign r_18[32] = _3992_ | _3991_ /*33752*/;
  assign _3993_ = ~q[14] /*33751*/;
  assign _3994_ = sum_18[19] & q[14] /*33750*/;
  assign _3995_ = m_18[19] & _3993_ /*33749*/;
  assign r_18[33] = _3995_ | _3994_ /*33748*/;
  assign _3996_ = ~q[14] /*33747*/;
  assign _3997_ = sum_18[20] & q[14] /*33746*/;
  assign _3998_ = m_18[20] & _3996_ /*33745*/;
  assign r_18[34] = _3998_ | _3997_ /*33744*/;
  assign _3999_ = ~q[14] /*33743*/;
  assign _4000_ = sum_18[21] & q[14] /*33742*/;
  assign _4001_ = m_18[21] & _3999_ /*33741*/;
  assign r_18[35] = _4001_ | _4000_ /*33740*/;
  assign _4002_ = ~q[14] /*33739*/;
  assign _4003_ = sum_18[22] & q[14] /*33738*/;
  assign _4004_ = m_18[22] & _4002_ /*33737*/;
  assign r_18[36] = _4004_ | _4003_ /*33736*/;
  assign _4005_ = ~q[14] /*33735*/;
  assign _4006_ = sum_18[23] & q[14] /*33734*/;
  assign _4007_ = m_18[23] & _4005_ /*33733*/;
  assign r_18[37] = _4007_ | _4006_ /*33732*/;
  assign _4008_ = ~q[14] /*33731*/;
  assign _4009_ = sum_18[24] & q[14] /*33730*/;
  assign _4010_ = m_18[24] & _4008_ /*33729*/;
  assign r_18[38] = _4010_ | _4009_ /*33728*/;
  assign _4011_ = ~q[14] /*33727*/;
  assign _4012_ = sum_18[25] & q[14] /*33726*/;
  assign _4013_ = m_18[25] & _4011_ /*33725*/;
  assign r_18[39] = _4013_ | _4012_ /*33724*/;
  assign _4014_ = ~q[14] /*33723*/;
  assign _4015_ = sum_18[26] & q[14] /*33722*/;
  assign _4016_ = m_18[26] & _4014_ /*33721*/;
  assign r_18[40] = _4016_ | _4015_ /*33720*/;
  assign _4017_ = ~q[14] /*33719*/;
  assign _4018_ = sum_18[27] & q[14] /*33718*/;
  assign _4019_ = m_18[27] & _4017_ /*33717*/;
  assign r_18[41] = _4019_ | _4018_ /*33716*/;
  assign _4020_ = ~q[14] /*33715*/;
  assign _4021_ = sum_18[28] & q[14] /*33714*/;
  assign _4022_ = m_18[28] & _4020_ /*33713*/;
  assign r_18[42] = _4022_ | _4021_ /*33712*/;
  assign _4023_ = ~q[14] /*33711*/;
  assign _4024_ = sum_18[29] & q[14] /*33710*/;
  assign _4025_ = m_18[29] & _4023_ /*33709*/;
  assign r_18[43] = _4025_ | _4024_ /*33708*/;
  assign _4026_ = ~q[14] /*33707*/;
  assign _4027_ = sum_18[30] & q[14] /*33706*/;
  assign _4028_ = m_18[30] & _4026_ /*33705*/;
  assign r_18[44] = _4028_ | _4027_ /*33704*/;
  assign _4029_ = ~q[14] /*33703*/;
  assign _4030_ = sum_18[31] & q[14] /*33702*/;
  assign _4031_ = m_18[31] & _4029_ /*33701*/;
  assign r_18[45] = _4031_ | _4030_ /*33700*/;
assign r_18[0]= r_17[0] /*33699*/;
assign r_18[1]= r_17[1] /*33698*/;
assign r_18[2]= r_17[2] /*33697*/;
assign r_18[3]= r_17[3] /*33696*/;
assign r_18[4]= r_17[4] /*33695*/;
assign r_18[5]= r_17[5] /*33694*/;
assign r_18[6]= r_17[6] /*33693*/;
assign r_18[7]= r_17[7] /*33692*/;
assign r_18[8]= r_17[8] /*33691*/;
assign r_18[9]= r_17[9] /*33690*/;
assign r_18[10]= r_17[10] /*33689*/;
assign r_18[11]= r_17[11] /*33688*/;
assign r_18[12]= r_17[12] /*33687*/;
assign r_18[13]= r_17[13] /*33686*/;
  assign inv_19[0] = ~div[0] /*33608*/;
  assign inv_19[1] = ~div[1] /*33607*/;
  assign inv_19[2] = ~div[2] /*33606*/;
  assign inv_19[3] = ~div[3] /*33605*/;
  assign inv_19[4] = ~div[4] /*33604*/;
  assign inv_19[5] = ~div[5] /*33603*/;
  assign inv_19[6] = ~div[6] /*33602*/;
  assign inv_19[7] = ~div[7] /*33601*/;
  assign inv_19[8] = ~div[8] /*33600*/;
  assign inv_19[9] = ~div[9] /*33599*/;
  assign inv_19[10] = ~div[10] /*33598*/;
  assign inv_19[11] = ~div[11] /*33597*/;
  assign inv_19[12] = ~div[12] /*33596*/;
  assign inv_19[13] = ~div[13] /*33595*/;
  assign inv_19[14] = ~div[14] /*33594*/;
  assign inv_19[15] = ~div[15] /*33593*/;
  assign inv_19[16] = ~div[16] /*33592*/;
  assign inv_19[17] = ~div[17] /*33591*/;
  assign inv_19[18] = ~div[18] /*33590*/;
  assign inv_19[19] = ~div[19] /*33589*/;
  assign inv_19[20] = ~div[20] /*33588*/;
  assign inv_19[21] = ~div[21] /*33587*/;
  assign inv_19[22] = ~div[22] /*33586*/;
  assign inv_19[23] = ~div[23] /*33585*/;
  assign inv_19[24] = ~div[24] /*33584*/;
  assign inv_19[25] = ~div[25] /*33583*/;
  assign inv_19[26] = ~div[26] /*33582*/;
  assign inv_19[27] = ~div[27] /*33581*/;
  assign inv_19[28] = ~div[28] /*33580*/;
  assign inv_19[29] = ~div[29] /*33579*/;
  assign inv_19[30] = ~div[30] /*33578*/;
assign inv_19[31] = oneWire /*33577*/;
  assign _4032_ = inv_19[0] ^ r_18[13] /*33575*/;
  assign sum_19[0] = _4032_ ^ oneWire /*33574*/;
  assign _4033_ = _4032_ & oneWire /*33573*/;
  assign _4034_ = inv_19[0] & r_18[13] /*33572*/;
  assign _4035_ = _4033_ | _4034_ /*33571*/;
  assign _4036_ = inv_19[1] ^ r_18[14] /*33570*/;
  assign sum_19[1] = _4036_ ^ _4035_ /*33569*/;
  assign _4037_ = _4036_ & _4035_ /*33568*/;
  assign _4038_ = inv_19[1] & r_18[14] /*33567*/;
  assign _4039_ = _4037_ | _4038_ /*33566*/;
  assign _4040_ = inv_19[2] ^ r_18[15] /*33564*/;
  assign sum_19[2] = _4040_ ^ _4039_ /*33563*/;
  assign _4041_ = _4040_ & _4039_ /*33562*/;
  assign _4042_ = inv_19[2] & r_18[15] /*33561*/;
  assign _4043_ = _4041_ | _4042_ /*33560*/;
  assign _4044_ = inv_19[3] ^ r_18[16] /*33558*/;
  assign sum_19[3] = _4044_ ^ _4043_ /*33557*/;
  assign _4045_ = _4044_ & _4043_ /*33556*/;
  assign _4046_ = inv_19[3] & r_18[16] /*33555*/;
  assign _4047_ = _4045_ | _4046_ /*33554*/;
  assign _4048_ = inv_19[4] ^ r_18[17] /*33552*/;
  assign sum_19[4] = _4048_ ^ _4047_ /*33551*/;
  assign _4049_ = _4048_ & _4047_ /*33550*/;
  assign _4050_ = inv_19[4] & r_18[17] /*33549*/;
  assign _4051_ = _4049_ | _4050_ /*33548*/;
  assign _4052_ = inv_19[5] ^ r_18[18] /*33546*/;
  assign sum_19[5] = _4052_ ^ _4051_ /*33545*/;
  assign _4053_ = _4052_ & _4051_ /*33544*/;
  assign _4054_ = inv_19[5] & r_18[18] /*33543*/;
  assign _4055_ = _4053_ | _4054_ /*33542*/;
  assign _4056_ = inv_19[6] ^ r_18[19] /*33540*/;
  assign sum_19[6] = _4056_ ^ _4055_ /*33539*/;
  assign _4057_ = _4056_ & _4055_ /*33538*/;
  assign _4058_ = inv_19[6] & r_18[19] /*33537*/;
  assign _4059_ = _4057_ | _4058_ /*33536*/;
  assign _4060_ = inv_19[7] ^ r_18[20] /*33534*/;
  assign sum_19[7] = _4060_ ^ _4059_ /*33533*/;
  assign _4061_ = _4060_ & _4059_ /*33532*/;
  assign _4062_ = inv_19[7] & r_18[20] /*33531*/;
  assign _4063_ = _4061_ | _4062_ /*33530*/;
  assign _4064_ = inv_19[8] ^ r_18[21] /*33528*/;
  assign sum_19[8] = _4064_ ^ _4063_ /*33527*/;
  assign _4065_ = _4064_ & _4063_ /*33526*/;
  assign _4066_ = inv_19[8] & r_18[21] /*33525*/;
  assign _4067_ = _4065_ | _4066_ /*33524*/;
  assign _4068_ = inv_19[9] ^ r_18[22] /*33522*/;
  assign sum_19[9] = _4068_ ^ _4067_ /*33521*/;
  assign _4069_ = _4068_ & _4067_ /*33520*/;
  assign _4070_ = inv_19[9] & r_18[22] /*33519*/;
  assign _4071_ = _4069_ | _4070_ /*33518*/;
  assign _4072_ = inv_19[10] ^ r_18[23] /*33516*/;
  assign sum_19[10] = _4072_ ^ _4071_ /*33515*/;
  assign _4073_ = _4072_ & _4071_ /*33514*/;
  assign _4074_ = inv_19[10] & r_18[23] /*33513*/;
  assign _4075_ = _4073_ | _4074_ /*33512*/;
  assign _4076_ = inv_19[11] ^ r_18[24] /*33510*/;
  assign sum_19[11] = _4076_ ^ _4075_ /*33509*/;
  assign _4077_ = _4076_ & _4075_ /*33508*/;
  assign _4078_ = inv_19[11] & r_18[24] /*33507*/;
  assign _4079_ = _4077_ | _4078_ /*33506*/;
  assign _4080_ = inv_19[12] ^ r_18[25] /*33504*/;
  assign sum_19[12] = _4080_ ^ _4079_ /*33503*/;
  assign _4081_ = _4080_ & _4079_ /*33502*/;
  assign _4082_ = inv_19[12] & r_18[25] /*33501*/;
  assign _4083_ = _4081_ | _4082_ /*33500*/;
  assign _4084_ = inv_19[13] ^ r_18[26] /*33498*/;
  assign sum_19[13] = _4084_ ^ _4083_ /*33497*/;
  assign _4085_ = _4084_ & _4083_ /*33496*/;
  assign _4086_ = inv_19[13] & r_18[26] /*33495*/;
  assign _4087_ = _4085_ | _4086_ /*33494*/;
  assign _4088_ = inv_19[14] ^ r_18[27] /*33492*/;
  assign sum_19[14] = _4088_ ^ _4087_ /*33491*/;
  assign _4089_ = _4088_ & _4087_ /*33490*/;
  assign _4090_ = inv_19[14] & r_18[27] /*33489*/;
  assign _4091_ = _4089_ | _4090_ /*33488*/;
  assign _4092_ = inv_19[15] ^ r_18[28] /*33486*/;
  assign sum_19[15] = _4092_ ^ _4091_ /*33485*/;
  assign _4093_ = _4092_ & _4091_ /*33484*/;
  assign _4094_ = inv_19[15] & r_18[28] /*33483*/;
  assign _4095_ = _4093_ | _4094_ /*33482*/;
  assign _4096_ = inv_19[16] ^ r_18[29] /*33480*/;
  assign sum_19[16] = _4096_ ^ _4095_ /*33479*/;
  assign _4097_ = _4096_ & _4095_ /*33478*/;
  assign _4098_ = inv_19[16] & r_18[29] /*33477*/;
  assign _4099_ = _4097_ | _4098_ /*33476*/;
  assign _4100_ = inv_19[17] ^ r_18[30] /*33474*/;
  assign sum_19[17] = _4100_ ^ _4099_ /*33473*/;
  assign _4101_ = _4100_ & _4099_ /*33472*/;
  assign _4102_ = inv_19[17] & r_18[30] /*33471*/;
  assign _4103_ = _4101_ | _4102_ /*33470*/;
  assign _4104_ = inv_19[18] ^ r_18[31] /*33468*/;
  assign sum_19[18] = _4104_ ^ _4103_ /*33467*/;
  assign _4105_ = _4104_ & _4103_ /*33466*/;
  assign _4106_ = inv_19[18] & r_18[31] /*33465*/;
  assign _4107_ = _4105_ | _4106_ /*33464*/;
  assign _4108_ = inv_19[19] ^ r_18[32] /*33462*/;
  assign sum_19[19] = _4108_ ^ _4107_ /*33461*/;
  assign _4109_ = _4108_ & _4107_ /*33460*/;
  assign _4110_ = inv_19[19] & r_18[32] /*33459*/;
  assign _4111_ = _4109_ | _4110_ /*33458*/;
  assign _4112_ = inv_19[20] ^ r_18[33] /*33456*/;
  assign sum_19[20] = _4112_ ^ _4111_ /*33455*/;
  assign _4113_ = _4112_ & _4111_ /*33454*/;
  assign _4114_ = inv_19[20] & r_18[33] /*33453*/;
  assign _4115_ = _4113_ | _4114_ /*33452*/;
  assign _4116_ = inv_19[21] ^ r_18[34] /*33450*/;
  assign sum_19[21] = _4116_ ^ _4115_ /*33449*/;
  assign _4117_ = _4116_ & _4115_ /*33448*/;
  assign _4118_ = inv_19[21] & r_18[34] /*33447*/;
  assign _4119_ = _4117_ | _4118_ /*33446*/;
  assign _4120_ = inv_19[22] ^ r_18[35] /*33444*/;
  assign sum_19[22] = _4120_ ^ _4119_ /*33443*/;
  assign _4121_ = _4120_ & _4119_ /*33442*/;
  assign _4122_ = inv_19[22] & r_18[35] /*33441*/;
  assign _4123_ = _4121_ | _4122_ /*33440*/;
  assign _4124_ = inv_19[23] ^ r_18[36] /*33438*/;
  assign sum_19[23] = _4124_ ^ _4123_ /*33437*/;
  assign _4125_ = _4124_ & _4123_ /*33436*/;
  assign _4126_ = inv_19[23] & r_18[36] /*33435*/;
  assign _4127_ = _4125_ | _4126_ /*33434*/;
  assign _4128_ = inv_19[24] ^ r_18[37] /*33432*/;
  assign sum_19[24] = _4128_ ^ _4127_ /*33431*/;
  assign _4129_ = _4128_ & _4127_ /*33430*/;
  assign _4130_ = inv_19[24] & r_18[37] /*33429*/;
  assign _4131_ = _4129_ | _4130_ /*33428*/;
  assign _4132_ = inv_19[25] ^ r_18[38] /*33426*/;
  assign sum_19[25] = _4132_ ^ _4131_ /*33425*/;
  assign _4133_ = _4132_ & _4131_ /*33424*/;
  assign _4134_ = inv_19[25] & r_18[38] /*33423*/;
  assign _4135_ = _4133_ | _4134_ /*33422*/;
  assign _4136_ = inv_19[26] ^ r_18[39] /*33420*/;
  assign sum_19[26] = _4136_ ^ _4135_ /*33419*/;
  assign _4137_ = _4136_ & _4135_ /*33418*/;
  assign _4138_ = inv_19[26] & r_18[39] /*33417*/;
  assign _4139_ = _4137_ | _4138_ /*33416*/;
  assign _4140_ = inv_19[27] ^ r_18[40] /*33414*/;
  assign sum_19[27] = _4140_ ^ _4139_ /*33413*/;
  assign _4141_ = _4140_ & _4139_ /*33412*/;
  assign _4142_ = inv_19[27] & r_18[40] /*33411*/;
  assign _4143_ = _4141_ | _4142_ /*33410*/;
  assign _4144_ = inv_19[28] ^ r_18[41] /*33408*/;
  assign sum_19[28] = _4144_ ^ _4143_ /*33407*/;
  assign _4145_ = _4144_ & _4143_ /*33406*/;
  assign _4146_ = inv_19[28] & r_18[41] /*33405*/;
  assign _4147_ = _4145_ | _4146_ /*33404*/;
  assign _4148_ = inv_19[29] ^ r_18[42] /*33402*/;
  assign sum_19[29] = _4148_ ^ _4147_ /*33401*/;
  assign _4149_ = _4148_ & _4147_ /*33400*/;
  assign _4150_ = inv_19[29] & r_18[42] /*33399*/;
  assign _4151_ = _4149_ | _4150_ /*33398*/;
  assign _4152_ = inv_19[30] ^ r_18[43] /*33396*/;
  assign sum_19[30] = _4152_ ^ _4151_ /*33395*/;
  assign _4153_ = _4152_ & _4151_ /*33394*/;
  assign _4154_ = inv_19[30] & r_18[43] /*33393*/;
  assign _4155_ = _4153_ | _4154_ /*33392*/;
  assign _4156_ = inv_19[31] ^ r_18[44] /*33390*/;
  assign sum_19[31] = _4156_ ^ _4155_ /*33389*/;
  assign _4157_ = _4156_ & _4155_ /*33388*/;
  assign _4158_ = inv_19[31] & r_18[44] /*33387*/;
  assign _4159_ = _4157_ | _4158_ /*33386*/;
  assign q[13] = ~sum_19[31] /*33413*/;
  assign m_19[0] = r_18[13] /*33412*/;
  assign m_19[1] = r_18[14] /*33411*/;
  assign m_19[2] = r_18[15] /*33410*/;
  assign m_19[3] = r_18[16] /*33409*/;
  assign m_19[4] = r_18[17] /*33408*/;
  assign m_19[5] = r_18[18] /*33407*/;
  assign m_19[6] = r_18[19] /*33406*/;
  assign m_19[7] = r_18[20] /*33405*/;
  assign m_19[8] = r_18[21] /*33404*/;
  assign m_19[9] = r_18[22] /*33403*/;
  assign m_19[10] = r_18[23] /*33402*/;
  assign m_19[11] = r_18[24] /*33401*/;
  assign m_19[12] = r_18[25] /*33400*/;
  assign m_19[13] = r_18[26] /*33399*/;
  assign m_19[14] = r_18[27] /*33398*/;
  assign m_19[15] = r_18[28] /*33397*/;
  assign m_19[16] = r_18[29] /*33396*/;
  assign m_19[17] = r_18[30] /*33395*/;
  assign m_19[18] = r_18[31] /*33394*/;
  assign m_19[19] = r_18[32] /*33393*/;
  assign m_19[20] = r_18[33] /*33392*/;
  assign m_19[21] = r_18[34] /*33391*/;
  assign m_19[22] = r_18[35] /*33390*/;
  assign m_19[23] = r_18[36] /*33389*/;
  assign m_19[24] = r_18[37] /*33388*/;
  assign m_19[25] = r_18[38] /*33387*/;
  assign m_19[26] = r_18[39] /*33386*/;
  assign m_19[27] = r_18[40] /*33385*/;
  assign m_19[28] = r_18[41] /*33384*/;
  assign m_19[29] = r_18[42] /*33383*/;
  assign m_19[30] = r_18[43] /*33382*/;
  assign m_19[31] = r_18[44] /*33381*/;
  assign _4160_ = ~q[13] /*33379*/;
  assign _4161_ = sum_19[0] & q[13] /*33378*/;
  assign _4162_ = m_19[0] & _4160_ /*33377*/;
  assign r_19[13] = _4162_ | _4161_ /*33376*/;
  assign _4163_ = ~q[13] /*33375*/;
  assign _4164_ = sum_19[1] & q[13] /*33374*/;
  assign _4165_ = m_19[1] & _4163_ /*33373*/;
  assign r_19[14] = _4165_ | _4164_ /*33372*/;
  assign _4166_ = ~q[13] /*33371*/;
  assign _4167_ = sum_19[2] & q[13] /*33370*/;
  assign _4168_ = m_19[2] & _4166_ /*33369*/;
  assign r_19[15] = _4168_ | _4167_ /*33368*/;
  assign _4169_ = ~q[13] /*33367*/;
  assign _4170_ = sum_19[3] & q[13] /*33366*/;
  assign _4171_ = m_19[3] & _4169_ /*33365*/;
  assign r_19[16] = _4171_ | _4170_ /*33364*/;
  assign _4172_ = ~q[13] /*33363*/;
  assign _4173_ = sum_19[4] & q[13] /*33362*/;
  assign _4174_ = m_19[4] & _4172_ /*33361*/;
  assign r_19[17] = _4174_ | _4173_ /*33360*/;
  assign _4175_ = ~q[13] /*33359*/;
  assign _4176_ = sum_19[5] & q[13] /*33358*/;
  assign _4177_ = m_19[5] & _4175_ /*33357*/;
  assign r_19[18] = _4177_ | _4176_ /*33356*/;
  assign _4178_ = ~q[13] /*33355*/;
  assign _4179_ = sum_19[6] & q[13] /*33354*/;
  assign _4180_ = m_19[6] & _4178_ /*33353*/;
  assign r_19[19] = _4180_ | _4179_ /*33352*/;
  assign _4181_ = ~q[13] /*33351*/;
  assign _4182_ = sum_19[7] & q[13] /*33350*/;
  assign _4183_ = m_19[7] & _4181_ /*33349*/;
  assign r_19[20] = _4183_ | _4182_ /*33348*/;
  assign _4184_ = ~q[13] /*33347*/;
  assign _4185_ = sum_19[8] & q[13] /*33346*/;
  assign _4186_ = m_19[8] & _4184_ /*33345*/;
  assign r_19[21] = _4186_ | _4185_ /*33344*/;
  assign _4187_ = ~q[13] /*33343*/;
  assign _4188_ = sum_19[9] & q[13] /*33342*/;
  assign _4189_ = m_19[9] & _4187_ /*33341*/;
  assign r_19[22] = _4189_ | _4188_ /*33340*/;
  assign _4190_ = ~q[13] /*33339*/;
  assign _4191_ = sum_19[10] & q[13] /*33338*/;
  assign _4192_ = m_19[10] & _4190_ /*33337*/;
  assign r_19[23] = _4192_ | _4191_ /*33336*/;
  assign _4193_ = ~q[13] /*33335*/;
  assign _4194_ = sum_19[11] & q[13] /*33334*/;
  assign _4195_ = m_19[11] & _4193_ /*33333*/;
  assign r_19[24] = _4195_ | _4194_ /*33332*/;
  assign _4196_ = ~q[13] /*33331*/;
  assign _4197_ = sum_19[12] & q[13] /*33330*/;
  assign _4198_ = m_19[12] & _4196_ /*33329*/;
  assign r_19[25] = _4198_ | _4197_ /*33328*/;
  assign _4199_ = ~q[13] /*33327*/;
  assign _4200_ = sum_19[13] & q[13] /*33326*/;
  assign _4201_ = m_19[13] & _4199_ /*33325*/;
  assign r_19[26] = _4201_ | _4200_ /*33324*/;
  assign _4202_ = ~q[13] /*33323*/;
  assign _4203_ = sum_19[14] & q[13] /*33322*/;
  assign _4204_ = m_19[14] & _4202_ /*33321*/;
  assign r_19[27] = _4204_ | _4203_ /*33320*/;
  assign _4205_ = ~q[13] /*33319*/;
  assign _4206_ = sum_19[15] & q[13] /*33318*/;
  assign _4207_ = m_19[15] & _4205_ /*33317*/;
  assign r_19[28] = _4207_ | _4206_ /*33316*/;
  assign _4208_ = ~q[13] /*33315*/;
  assign _4209_ = sum_19[16] & q[13] /*33314*/;
  assign _4210_ = m_19[16] & _4208_ /*33313*/;
  assign r_19[29] = _4210_ | _4209_ /*33312*/;
  assign _4211_ = ~q[13] /*33311*/;
  assign _4212_ = sum_19[17] & q[13] /*33310*/;
  assign _4213_ = m_19[17] & _4211_ /*33309*/;
  assign r_19[30] = _4213_ | _4212_ /*33308*/;
  assign _4214_ = ~q[13] /*33307*/;
  assign _4215_ = sum_19[18] & q[13] /*33306*/;
  assign _4216_ = m_19[18] & _4214_ /*33305*/;
  assign r_19[31] = _4216_ | _4215_ /*33304*/;
  assign _4217_ = ~q[13] /*33303*/;
  assign _4218_ = sum_19[19] & q[13] /*33302*/;
  assign _4219_ = m_19[19] & _4217_ /*33301*/;
  assign r_19[32] = _4219_ | _4218_ /*33300*/;
  assign _4220_ = ~q[13] /*33299*/;
  assign _4221_ = sum_19[20] & q[13] /*33298*/;
  assign _4222_ = m_19[20] & _4220_ /*33297*/;
  assign r_19[33] = _4222_ | _4221_ /*33296*/;
  assign _4223_ = ~q[13] /*33295*/;
  assign _4224_ = sum_19[21] & q[13] /*33294*/;
  assign _4225_ = m_19[21] & _4223_ /*33293*/;
  assign r_19[34] = _4225_ | _4224_ /*33292*/;
  assign _4226_ = ~q[13] /*33291*/;
  assign _4227_ = sum_19[22] & q[13] /*33290*/;
  assign _4228_ = m_19[22] & _4226_ /*33289*/;
  assign r_19[35] = _4228_ | _4227_ /*33288*/;
  assign _4229_ = ~q[13] /*33287*/;
  assign _4230_ = sum_19[23] & q[13] /*33286*/;
  assign _4231_ = m_19[23] & _4229_ /*33285*/;
  assign r_19[36] = _4231_ | _4230_ /*33284*/;
  assign _4232_ = ~q[13] /*33283*/;
  assign _4233_ = sum_19[24] & q[13] /*33282*/;
  assign _4234_ = m_19[24] & _4232_ /*33281*/;
  assign r_19[37] = _4234_ | _4233_ /*33280*/;
  assign _4235_ = ~q[13] /*33279*/;
  assign _4236_ = sum_19[25] & q[13] /*33278*/;
  assign _4237_ = m_19[25] & _4235_ /*33277*/;
  assign r_19[38] = _4237_ | _4236_ /*33276*/;
  assign _4238_ = ~q[13] /*33275*/;
  assign _4239_ = sum_19[26] & q[13] /*33274*/;
  assign _4240_ = m_19[26] & _4238_ /*33273*/;
  assign r_19[39] = _4240_ | _4239_ /*33272*/;
  assign _4241_ = ~q[13] /*33271*/;
  assign _4242_ = sum_19[27] & q[13] /*33270*/;
  assign _4243_ = m_19[27] & _4241_ /*33269*/;
  assign r_19[40] = _4243_ | _4242_ /*33268*/;
  assign _4244_ = ~q[13] /*33267*/;
  assign _4245_ = sum_19[28] & q[13] /*33266*/;
  assign _4246_ = m_19[28] & _4244_ /*33265*/;
  assign r_19[41] = _4246_ | _4245_ /*33264*/;
  assign _4247_ = ~q[13] /*33263*/;
  assign _4248_ = sum_19[29] & q[13] /*33262*/;
  assign _4249_ = m_19[29] & _4247_ /*33261*/;
  assign r_19[42] = _4249_ | _4248_ /*33260*/;
  assign _4250_ = ~q[13] /*33259*/;
  assign _4251_ = sum_19[30] & q[13] /*33258*/;
  assign _4252_ = m_19[30] & _4250_ /*33257*/;
  assign r_19[43] = _4252_ | _4251_ /*33256*/;
  assign _4253_ = ~q[13] /*33255*/;
  assign _4254_ = sum_19[31] & q[13] /*33254*/;
  assign _4255_ = m_19[31] & _4253_ /*33253*/;
  assign r_19[44] = _4255_ | _4254_ /*33252*/;
assign r_19[0]= r_18[0] /*33251*/;
assign r_19[1]= r_18[1] /*33250*/;
assign r_19[2]= r_18[2] /*33249*/;
assign r_19[3]= r_18[3] /*33248*/;
assign r_19[4]= r_18[4] /*33247*/;
assign r_19[5]= r_18[5] /*33246*/;
assign r_19[6]= r_18[6] /*33245*/;
assign r_19[7]= r_18[7] /*33244*/;
assign r_19[8]= r_18[8] /*33243*/;
assign r_19[9]= r_18[9] /*33242*/;
assign r_19[10]= r_18[10] /*33241*/;
assign r_19[11]= r_18[11] /*33240*/;
assign r_19[12]= r_18[12] /*33239*/;
  assign inv_20[0] = ~div[0] /*33160*/;
  assign inv_20[1] = ~div[1] /*33159*/;
  assign inv_20[2] = ~div[2] /*33158*/;
  assign inv_20[3] = ~div[3] /*33157*/;
  assign inv_20[4] = ~div[4] /*33156*/;
  assign inv_20[5] = ~div[5] /*33155*/;
  assign inv_20[6] = ~div[6] /*33154*/;
  assign inv_20[7] = ~div[7] /*33153*/;
  assign inv_20[8] = ~div[8] /*33152*/;
  assign inv_20[9] = ~div[9] /*33151*/;
  assign inv_20[10] = ~div[10] /*33150*/;
  assign inv_20[11] = ~div[11] /*33149*/;
  assign inv_20[12] = ~div[12] /*33148*/;
  assign inv_20[13] = ~div[13] /*33147*/;
  assign inv_20[14] = ~div[14] /*33146*/;
  assign inv_20[15] = ~div[15] /*33145*/;
  assign inv_20[16] = ~div[16] /*33144*/;
  assign inv_20[17] = ~div[17] /*33143*/;
  assign inv_20[18] = ~div[18] /*33142*/;
  assign inv_20[19] = ~div[19] /*33141*/;
  assign inv_20[20] = ~div[20] /*33140*/;
  assign inv_20[21] = ~div[21] /*33139*/;
  assign inv_20[22] = ~div[22] /*33138*/;
  assign inv_20[23] = ~div[23] /*33137*/;
  assign inv_20[24] = ~div[24] /*33136*/;
  assign inv_20[25] = ~div[25] /*33135*/;
  assign inv_20[26] = ~div[26] /*33134*/;
  assign inv_20[27] = ~div[27] /*33133*/;
  assign inv_20[28] = ~div[28] /*33132*/;
  assign inv_20[29] = ~div[29] /*33131*/;
  assign inv_20[30] = ~div[30] /*33130*/;
assign inv_20[31] = oneWire /*33129*/;
  assign _4256_ = inv_20[0] ^ r_19[12] /*33127*/;
  assign sum_20[0] = _4256_ ^ oneWire /*33126*/;
  assign _4257_ = _4256_ & oneWire /*33125*/;
  assign _4258_ = inv_20[0] & r_19[12] /*33124*/;
  assign _4259_ = _4257_ | _4258_ /*33123*/;
  assign _4260_ = inv_20[1] ^ r_19[13] /*33122*/;
  assign sum_20[1] = _4260_ ^ _4259_ /*33121*/;
  assign _4261_ = _4260_ & _4259_ /*33120*/;
  assign _4262_ = inv_20[1] & r_19[13] /*33119*/;
  assign _4263_ = _4261_ | _4262_ /*33118*/;
  assign _4264_ = inv_20[2] ^ r_19[14] /*33116*/;
  assign sum_20[2] = _4264_ ^ _4263_ /*33115*/;
  assign _4265_ = _4264_ & _4263_ /*33114*/;
  assign _4266_ = inv_20[2] & r_19[14] /*33113*/;
  assign _4267_ = _4265_ | _4266_ /*33112*/;
  assign _4268_ = inv_20[3] ^ r_19[15] /*33110*/;
  assign sum_20[3] = _4268_ ^ _4267_ /*33109*/;
  assign _4269_ = _4268_ & _4267_ /*33108*/;
  assign _4270_ = inv_20[3] & r_19[15] /*33107*/;
  assign _4271_ = _4269_ | _4270_ /*33106*/;
  assign _4272_ = inv_20[4] ^ r_19[16] /*33104*/;
  assign sum_20[4] = _4272_ ^ _4271_ /*33103*/;
  assign _4273_ = _4272_ & _4271_ /*33102*/;
  assign _4274_ = inv_20[4] & r_19[16] /*33101*/;
  assign _4275_ = _4273_ | _4274_ /*33100*/;
  assign _4276_ = inv_20[5] ^ r_19[17] /*33098*/;
  assign sum_20[5] = _4276_ ^ _4275_ /*33097*/;
  assign _4277_ = _4276_ & _4275_ /*33096*/;
  assign _4278_ = inv_20[5] & r_19[17] /*33095*/;
  assign _4279_ = _4277_ | _4278_ /*33094*/;
  assign _4280_ = inv_20[6] ^ r_19[18] /*33092*/;
  assign sum_20[6] = _4280_ ^ _4279_ /*33091*/;
  assign _4281_ = _4280_ & _4279_ /*33090*/;
  assign _4282_ = inv_20[6] & r_19[18] /*33089*/;
  assign _4283_ = _4281_ | _4282_ /*33088*/;
  assign _4284_ = inv_20[7] ^ r_19[19] /*33086*/;
  assign sum_20[7] = _4284_ ^ _4283_ /*33085*/;
  assign _4285_ = _4284_ & _4283_ /*33084*/;
  assign _4286_ = inv_20[7] & r_19[19] /*33083*/;
  assign _4287_ = _4285_ | _4286_ /*33082*/;
  assign _4288_ = inv_20[8] ^ r_19[20] /*33080*/;
  assign sum_20[8] = _4288_ ^ _4287_ /*33079*/;
  assign _4289_ = _4288_ & _4287_ /*33078*/;
  assign _4290_ = inv_20[8] & r_19[20] /*33077*/;
  assign _4291_ = _4289_ | _4290_ /*33076*/;
  assign _4292_ = inv_20[9] ^ r_19[21] /*33074*/;
  assign sum_20[9] = _4292_ ^ _4291_ /*33073*/;
  assign _4293_ = _4292_ & _4291_ /*33072*/;
  assign _4294_ = inv_20[9] & r_19[21] /*33071*/;
  assign _4295_ = _4293_ | _4294_ /*33070*/;
  assign _4296_ = inv_20[10] ^ r_19[22] /*33068*/;
  assign sum_20[10] = _4296_ ^ _4295_ /*33067*/;
  assign _4297_ = _4296_ & _4295_ /*33066*/;
  assign _4298_ = inv_20[10] & r_19[22] /*33065*/;
  assign _4299_ = _4297_ | _4298_ /*33064*/;
  assign _4300_ = inv_20[11] ^ r_19[23] /*33062*/;
  assign sum_20[11] = _4300_ ^ _4299_ /*33061*/;
  assign _4301_ = _4300_ & _4299_ /*33060*/;
  assign _4302_ = inv_20[11] & r_19[23] /*33059*/;
  assign _4303_ = _4301_ | _4302_ /*33058*/;
  assign _4304_ = inv_20[12] ^ r_19[24] /*33056*/;
  assign sum_20[12] = _4304_ ^ _4303_ /*33055*/;
  assign _4305_ = _4304_ & _4303_ /*33054*/;
  assign _4306_ = inv_20[12] & r_19[24] /*33053*/;
  assign _4307_ = _4305_ | _4306_ /*33052*/;
  assign _4308_ = inv_20[13] ^ r_19[25] /*33050*/;
  assign sum_20[13] = _4308_ ^ _4307_ /*33049*/;
  assign _4309_ = _4308_ & _4307_ /*33048*/;
  assign _4310_ = inv_20[13] & r_19[25] /*33047*/;
  assign _4311_ = _4309_ | _4310_ /*33046*/;
  assign _4312_ = inv_20[14] ^ r_19[26] /*33044*/;
  assign sum_20[14] = _4312_ ^ _4311_ /*33043*/;
  assign _4313_ = _4312_ & _4311_ /*33042*/;
  assign _4314_ = inv_20[14] & r_19[26] /*33041*/;
  assign _4315_ = _4313_ | _4314_ /*33040*/;
  assign _4316_ = inv_20[15] ^ r_19[27] /*33038*/;
  assign sum_20[15] = _4316_ ^ _4315_ /*33037*/;
  assign _4317_ = _4316_ & _4315_ /*33036*/;
  assign _4318_ = inv_20[15] & r_19[27] /*33035*/;
  assign _4319_ = _4317_ | _4318_ /*33034*/;
  assign _4320_ = inv_20[16] ^ r_19[28] /*33032*/;
  assign sum_20[16] = _4320_ ^ _4319_ /*33031*/;
  assign _4321_ = _4320_ & _4319_ /*33030*/;
  assign _4322_ = inv_20[16] & r_19[28] /*33029*/;
  assign _4323_ = _4321_ | _4322_ /*33028*/;
  assign _4324_ = inv_20[17] ^ r_19[29] /*33026*/;
  assign sum_20[17] = _4324_ ^ _4323_ /*33025*/;
  assign _4325_ = _4324_ & _4323_ /*33024*/;
  assign _4326_ = inv_20[17] & r_19[29] /*33023*/;
  assign _4327_ = _4325_ | _4326_ /*33022*/;
  assign _4328_ = inv_20[18] ^ r_19[30] /*33020*/;
  assign sum_20[18] = _4328_ ^ _4327_ /*33019*/;
  assign _4329_ = _4328_ & _4327_ /*33018*/;
  assign _4330_ = inv_20[18] & r_19[30] /*33017*/;
  assign _4331_ = _4329_ | _4330_ /*33016*/;
  assign _4332_ = inv_20[19] ^ r_19[31] /*33014*/;
  assign sum_20[19] = _4332_ ^ _4331_ /*33013*/;
  assign _4333_ = _4332_ & _4331_ /*33012*/;
  assign _4334_ = inv_20[19] & r_19[31] /*33011*/;
  assign _4335_ = _4333_ | _4334_ /*33010*/;
  assign _4336_ = inv_20[20] ^ r_19[32] /*33008*/;
  assign sum_20[20] = _4336_ ^ _4335_ /*33007*/;
  assign _4337_ = _4336_ & _4335_ /*33006*/;
  assign _4338_ = inv_20[20] & r_19[32] /*33005*/;
  assign _4339_ = _4337_ | _4338_ /*33004*/;
  assign _4340_ = inv_20[21] ^ r_19[33] /*33002*/;
  assign sum_20[21] = _4340_ ^ _4339_ /*33001*/;
  assign _4341_ = _4340_ & _4339_ /*33000*/;
  assign _4342_ = inv_20[21] & r_19[33] /*32999*/;
  assign _4343_ = _4341_ | _4342_ /*32998*/;
  assign _4344_ = inv_20[22] ^ r_19[34] /*32996*/;
  assign sum_20[22] = _4344_ ^ _4343_ /*32995*/;
  assign _4345_ = _4344_ & _4343_ /*32994*/;
  assign _4346_ = inv_20[22] & r_19[34] /*32993*/;
  assign _4347_ = _4345_ | _4346_ /*32992*/;
  assign _4348_ = inv_20[23] ^ r_19[35] /*32990*/;
  assign sum_20[23] = _4348_ ^ _4347_ /*32989*/;
  assign _4349_ = _4348_ & _4347_ /*32988*/;
  assign _4350_ = inv_20[23] & r_19[35] /*32987*/;
  assign _4351_ = _4349_ | _4350_ /*32986*/;
  assign _4352_ = inv_20[24] ^ r_19[36] /*32984*/;
  assign sum_20[24] = _4352_ ^ _4351_ /*32983*/;
  assign _4353_ = _4352_ & _4351_ /*32982*/;
  assign _4354_ = inv_20[24] & r_19[36] /*32981*/;
  assign _4355_ = _4353_ | _4354_ /*32980*/;
  assign _4356_ = inv_20[25] ^ r_19[37] /*32978*/;
  assign sum_20[25] = _4356_ ^ _4355_ /*32977*/;
  assign _4357_ = _4356_ & _4355_ /*32976*/;
  assign _4358_ = inv_20[25] & r_19[37] /*32975*/;
  assign _4359_ = _4357_ | _4358_ /*32974*/;
  assign _4360_ = inv_20[26] ^ r_19[38] /*32972*/;
  assign sum_20[26] = _4360_ ^ _4359_ /*32971*/;
  assign _4361_ = _4360_ & _4359_ /*32970*/;
  assign _4362_ = inv_20[26] & r_19[38] /*32969*/;
  assign _4363_ = _4361_ | _4362_ /*32968*/;
  assign _4364_ = inv_20[27] ^ r_19[39] /*32966*/;
  assign sum_20[27] = _4364_ ^ _4363_ /*32965*/;
  assign _4365_ = _4364_ & _4363_ /*32964*/;
  assign _4366_ = inv_20[27] & r_19[39] /*32963*/;
  assign _4367_ = _4365_ | _4366_ /*32962*/;
  assign _4368_ = inv_20[28] ^ r_19[40] /*32960*/;
  assign sum_20[28] = _4368_ ^ _4367_ /*32959*/;
  assign _4369_ = _4368_ & _4367_ /*32958*/;
  assign _4370_ = inv_20[28] & r_19[40] /*32957*/;
  assign _4371_ = _4369_ | _4370_ /*32956*/;
  assign _4372_ = inv_20[29] ^ r_19[41] /*32954*/;
  assign sum_20[29] = _4372_ ^ _4371_ /*32953*/;
  assign _4373_ = _4372_ & _4371_ /*32952*/;
  assign _4374_ = inv_20[29] & r_19[41] /*32951*/;
  assign _4375_ = _4373_ | _4374_ /*32950*/;
  assign _4376_ = inv_20[30] ^ r_19[42] /*32948*/;
  assign sum_20[30] = _4376_ ^ _4375_ /*32947*/;
  assign _4377_ = _4376_ & _4375_ /*32946*/;
  assign _4378_ = inv_20[30] & r_19[42] /*32945*/;
  assign _4379_ = _4377_ | _4378_ /*32944*/;
  assign _4380_ = inv_20[31] ^ r_19[43] /*32942*/;
  assign sum_20[31] = _4380_ ^ _4379_ /*32941*/;
  assign _4381_ = _4380_ & _4379_ /*32940*/;
  assign _4382_ = inv_20[31] & r_19[43] /*32939*/;
  assign _4383_ = _4381_ | _4382_ /*32938*/;
  assign q[12] = ~sum_20[31] /*32965*/;
  assign m_20[0] = r_19[12] /*32964*/;
  assign m_20[1] = r_19[13] /*32963*/;
  assign m_20[2] = r_19[14] /*32962*/;
  assign m_20[3] = r_19[15] /*32961*/;
  assign m_20[4] = r_19[16] /*32960*/;
  assign m_20[5] = r_19[17] /*32959*/;
  assign m_20[6] = r_19[18] /*32958*/;
  assign m_20[7] = r_19[19] /*32957*/;
  assign m_20[8] = r_19[20] /*32956*/;
  assign m_20[9] = r_19[21] /*32955*/;
  assign m_20[10] = r_19[22] /*32954*/;
  assign m_20[11] = r_19[23] /*32953*/;
  assign m_20[12] = r_19[24] /*32952*/;
  assign m_20[13] = r_19[25] /*32951*/;
  assign m_20[14] = r_19[26] /*32950*/;
  assign m_20[15] = r_19[27] /*32949*/;
  assign m_20[16] = r_19[28] /*32948*/;
  assign m_20[17] = r_19[29] /*32947*/;
  assign m_20[18] = r_19[30] /*32946*/;
  assign m_20[19] = r_19[31] /*32945*/;
  assign m_20[20] = r_19[32] /*32944*/;
  assign m_20[21] = r_19[33] /*32943*/;
  assign m_20[22] = r_19[34] /*32942*/;
  assign m_20[23] = r_19[35] /*32941*/;
  assign m_20[24] = r_19[36] /*32940*/;
  assign m_20[25] = r_19[37] /*32939*/;
  assign m_20[26] = r_19[38] /*32938*/;
  assign m_20[27] = r_19[39] /*32937*/;
  assign m_20[28] = r_19[40] /*32936*/;
  assign m_20[29] = r_19[41] /*32935*/;
  assign m_20[30] = r_19[42] /*32934*/;
  assign m_20[31] = r_19[43] /*32933*/;
  assign _4384_ = ~q[12] /*32931*/;
  assign _4385_ = sum_20[0] & q[12] /*32930*/;
  assign _4386_ = m_20[0] & _4384_ /*32929*/;
  assign r_20[12] = _4386_ | _4385_ /*32928*/;
  assign _4387_ = ~q[12] /*32927*/;
  assign _4388_ = sum_20[1] & q[12] /*32926*/;
  assign _4389_ = m_20[1] & _4387_ /*32925*/;
  assign r_20[13] = _4389_ | _4388_ /*32924*/;
  assign _4390_ = ~q[12] /*32923*/;
  assign _4391_ = sum_20[2] & q[12] /*32922*/;
  assign _4392_ = m_20[2] & _4390_ /*32921*/;
  assign r_20[14] = _4392_ | _4391_ /*32920*/;
  assign _4393_ = ~q[12] /*32919*/;
  assign _4394_ = sum_20[3] & q[12] /*32918*/;
  assign _4395_ = m_20[3] & _4393_ /*32917*/;
  assign r_20[15] = _4395_ | _4394_ /*32916*/;
  assign _4396_ = ~q[12] /*32915*/;
  assign _4397_ = sum_20[4] & q[12] /*32914*/;
  assign _4398_ = m_20[4] & _4396_ /*32913*/;
  assign r_20[16] = _4398_ | _4397_ /*32912*/;
  assign _4399_ = ~q[12] /*32911*/;
  assign _4400_ = sum_20[5] & q[12] /*32910*/;
  assign _4401_ = m_20[5] & _4399_ /*32909*/;
  assign r_20[17] = _4401_ | _4400_ /*32908*/;
  assign _4402_ = ~q[12] /*32907*/;
  assign _4403_ = sum_20[6] & q[12] /*32906*/;
  assign _4404_ = m_20[6] & _4402_ /*32905*/;
  assign r_20[18] = _4404_ | _4403_ /*32904*/;
  assign _4405_ = ~q[12] /*32903*/;
  assign _4406_ = sum_20[7] & q[12] /*32902*/;
  assign _4407_ = m_20[7] & _4405_ /*32901*/;
  assign r_20[19] = _4407_ | _4406_ /*32900*/;
  assign _4408_ = ~q[12] /*32899*/;
  assign _4409_ = sum_20[8] & q[12] /*32898*/;
  assign _4410_ = m_20[8] & _4408_ /*32897*/;
  assign r_20[20] = _4410_ | _4409_ /*32896*/;
  assign _4411_ = ~q[12] /*32895*/;
  assign _4412_ = sum_20[9] & q[12] /*32894*/;
  assign _4413_ = m_20[9] & _4411_ /*32893*/;
  assign r_20[21] = _4413_ | _4412_ /*32892*/;
  assign _4414_ = ~q[12] /*32891*/;
  assign _4415_ = sum_20[10] & q[12] /*32890*/;
  assign _4416_ = m_20[10] & _4414_ /*32889*/;
  assign r_20[22] = _4416_ | _4415_ /*32888*/;
  assign _4417_ = ~q[12] /*32887*/;
  assign _4418_ = sum_20[11] & q[12] /*32886*/;
  assign _4419_ = m_20[11] & _4417_ /*32885*/;
  assign r_20[23] = _4419_ | _4418_ /*32884*/;
  assign _4420_ = ~q[12] /*32883*/;
  assign _4421_ = sum_20[12] & q[12] /*32882*/;
  assign _4422_ = m_20[12] & _4420_ /*32881*/;
  assign r_20[24] = _4422_ | _4421_ /*32880*/;
  assign _4423_ = ~q[12] /*32879*/;
  assign _4424_ = sum_20[13] & q[12] /*32878*/;
  assign _4425_ = m_20[13] & _4423_ /*32877*/;
  assign r_20[25] = _4425_ | _4424_ /*32876*/;
  assign _4426_ = ~q[12] /*32875*/;
  assign _4427_ = sum_20[14] & q[12] /*32874*/;
  assign _4428_ = m_20[14] & _4426_ /*32873*/;
  assign r_20[26] = _4428_ | _4427_ /*32872*/;
  assign _4429_ = ~q[12] /*32871*/;
  assign _4430_ = sum_20[15] & q[12] /*32870*/;
  assign _4431_ = m_20[15] & _4429_ /*32869*/;
  assign r_20[27] = _4431_ | _4430_ /*32868*/;
  assign _4432_ = ~q[12] /*32867*/;
  assign _4433_ = sum_20[16] & q[12] /*32866*/;
  assign _4434_ = m_20[16] & _4432_ /*32865*/;
  assign r_20[28] = _4434_ | _4433_ /*32864*/;
  assign _4435_ = ~q[12] /*32863*/;
  assign _4436_ = sum_20[17] & q[12] /*32862*/;
  assign _4437_ = m_20[17] & _4435_ /*32861*/;
  assign r_20[29] = _4437_ | _4436_ /*32860*/;
  assign _4438_ = ~q[12] /*32859*/;
  assign _4439_ = sum_20[18] & q[12] /*32858*/;
  assign _4440_ = m_20[18] & _4438_ /*32857*/;
  assign r_20[30] = _4440_ | _4439_ /*32856*/;
  assign _4441_ = ~q[12] /*32855*/;
  assign _4442_ = sum_20[19] & q[12] /*32854*/;
  assign _4443_ = m_20[19] & _4441_ /*32853*/;
  assign r_20[31] = _4443_ | _4442_ /*32852*/;
  assign _4444_ = ~q[12] /*32851*/;
  assign _4445_ = sum_20[20] & q[12] /*32850*/;
  assign _4446_ = m_20[20] & _4444_ /*32849*/;
  assign r_20[32] = _4446_ | _4445_ /*32848*/;
  assign _4447_ = ~q[12] /*32847*/;
  assign _4448_ = sum_20[21] & q[12] /*32846*/;
  assign _4449_ = m_20[21] & _4447_ /*32845*/;
  assign r_20[33] = _4449_ | _4448_ /*32844*/;
  assign _4450_ = ~q[12] /*32843*/;
  assign _4451_ = sum_20[22] & q[12] /*32842*/;
  assign _4452_ = m_20[22] & _4450_ /*32841*/;
  assign r_20[34] = _4452_ | _4451_ /*32840*/;
  assign _4453_ = ~q[12] /*32839*/;
  assign _4454_ = sum_20[23] & q[12] /*32838*/;
  assign _4455_ = m_20[23] & _4453_ /*32837*/;
  assign r_20[35] = _4455_ | _4454_ /*32836*/;
  assign _4456_ = ~q[12] /*32835*/;
  assign _4457_ = sum_20[24] & q[12] /*32834*/;
  assign _4458_ = m_20[24] & _4456_ /*32833*/;
  assign r_20[36] = _4458_ | _4457_ /*32832*/;
  assign _4459_ = ~q[12] /*32831*/;
  assign _4460_ = sum_20[25] & q[12] /*32830*/;
  assign _4461_ = m_20[25] & _4459_ /*32829*/;
  assign r_20[37] = _4461_ | _4460_ /*32828*/;
  assign _4462_ = ~q[12] /*32827*/;
  assign _4463_ = sum_20[26] & q[12] /*32826*/;
  assign _4464_ = m_20[26] & _4462_ /*32825*/;
  assign r_20[38] = _4464_ | _4463_ /*32824*/;
  assign _4465_ = ~q[12] /*32823*/;
  assign _4466_ = sum_20[27] & q[12] /*32822*/;
  assign _4467_ = m_20[27] & _4465_ /*32821*/;
  assign r_20[39] = _4467_ | _4466_ /*32820*/;
  assign _4468_ = ~q[12] /*32819*/;
  assign _4469_ = sum_20[28] & q[12] /*32818*/;
  assign _4470_ = m_20[28] & _4468_ /*32817*/;
  assign r_20[40] = _4470_ | _4469_ /*32816*/;
  assign _4471_ = ~q[12] /*32815*/;
  assign _4472_ = sum_20[29] & q[12] /*32814*/;
  assign _4473_ = m_20[29] & _4471_ /*32813*/;
  assign r_20[41] = _4473_ | _4472_ /*32812*/;
  assign _4474_ = ~q[12] /*32811*/;
  assign _4475_ = sum_20[30] & q[12] /*32810*/;
  assign _4476_ = m_20[30] & _4474_ /*32809*/;
  assign r_20[42] = _4476_ | _4475_ /*32808*/;
  assign _4477_ = ~q[12] /*32807*/;
  assign _4478_ = sum_20[31] & q[12] /*32806*/;
  assign _4479_ = m_20[31] & _4477_ /*32805*/;
  assign r_20[43] = _4479_ | _4478_ /*32804*/;
assign r_20[0]= r_19[0] /*32803*/;
assign r_20[1]= r_19[1] /*32802*/;
assign r_20[2]= r_19[2] /*32801*/;
assign r_20[3]= r_19[3] /*32800*/;
assign r_20[4]= r_19[4] /*32799*/;
assign r_20[5]= r_19[5] /*32798*/;
assign r_20[6]= r_19[6] /*32797*/;
assign r_20[7]= r_19[7] /*32796*/;
assign r_20[8]= r_19[8] /*32795*/;
assign r_20[9]= r_19[9] /*32794*/;
assign r_20[10]= r_19[10] /*32793*/;
assign r_20[11]= r_19[11] /*32792*/;
  assign inv_21[0] = ~div[0] /*32712*/;
  assign inv_21[1] = ~div[1] /*32711*/;
  assign inv_21[2] = ~div[2] /*32710*/;
  assign inv_21[3] = ~div[3] /*32709*/;
  assign inv_21[4] = ~div[4] /*32708*/;
  assign inv_21[5] = ~div[5] /*32707*/;
  assign inv_21[6] = ~div[6] /*32706*/;
  assign inv_21[7] = ~div[7] /*32705*/;
  assign inv_21[8] = ~div[8] /*32704*/;
  assign inv_21[9] = ~div[9] /*32703*/;
  assign inv_21[10] = ~div[10] /*32702*/;
  assign inv_21[11] = ~div[11] /*32701*/;
  assign inv_21[12] = ~div[12] /*32700*/;
  assign inv_21[13] = ~div[13] /*32699*/;
  assign inv_21[14] = ~div[14] /*32698*/;
  assign inv_21[15] = ~div[15] /*32697*/;
  assign inv_21[16] = ~div[16] /*32696*/;
  assign inv_21[17] = ~div[17] /*32695*/;
  assign inv_21[18] = ~div[18] /*32694*/;
  assign inv_21[19] = ~div[19] /*32693*/;
  assign inv_21[20] = ~div[20] /*32692*/;
  assign inv_21[21] = ~div[21] /*32691*/;
  assign inv_21[22] = ~div[22] /*32690*/;
  assign inv_21[23] = ~div[23] /*32689*/;
  assign inv_21[24] = ~div[24] /*32688*/;
  assign inv_21[25] = ~div[25] /*32687*/;
  assign inv_21[26] = ~div[26] /*32686*/;
  assign inv_21[27] = ~div[27] /*32685*/;
  assign inv_21[28] = ~div[28] /*32684*/;
  assign inv_21[29] = ~div[29] /*32683*/;
  assign inv_21[30] = ~div[30] /*32682*/;
assign inv_21[31] = oneWire /*32681*/;
  assign _4480_ = inv_21[0] ^ r_20[11] /*32679*/;
  assign sum_21[0] = _4480_ ^ oneWire /*32678*/;
  assign _4481_ = _4480_ & oneWire /*32677*/;
  assign _4482_ = inv_21[0] & r_20[11] /*32676*/;
  assign _4483_ = _4481_ | _4482_ /*32675*/;
  assign _4484_ = inv_21[1] ^ r_20[12] /*32674*/;
  assign sum_21[1] = _4484_ ^ _4483_ /*32673*/;
  assign _4485_ = _4484_ & _4483_ /*32672*/;
  assign _4486_ = inv_21[1] & r_20[12] /*32671*/;
  assign _4487_ = _4485_ | _4486_ /*32670*/;
  assign _4488_ = inv_21[2] ^ r_20[13] /*32668*/;
  assign sum_21[2] = _4488_ ^ _4487_ /*32667*/;
  assign _4489_ = _4488_ & _4487_ /*32666*/;
  assign _4490_ = inv_21[2] & r_20[13] /*32665*/;
  assign _4491_ = _4489_ | _4490_ /*32664*/;
  assign _4492_ = inv_21[3] ^ r_20[14] /*32662*/;
  assign sum_21[3] = _4492_ ^ _4491_ /*32661*/;
  assign _4493_ = _4492_ & _4491_ /*32660*/;
  assign _4494_ = inv_21[3] & r_20[14] /*32659*/;
  assign _4495_ = _4493_ | _4494_ /*32658*/;
  assign _4496_ = inv_21[4] ^ r_20[15] /*32656*/;
  assign sum_21[4] = _4496_ ^ _4495_ /*32655*/;
  assign _4497_ = _4496_ & _4495_ /*32654*/;
  assign _4498_ = inv_21[4] & r_20[15] /*32653*/;
  assign _4499_ = _4497_ | _4498_ /*32652*/;
  assign _4500_ = inv_21[5] ^ r_20[16] /*32650*/;
  assign sum_21[5] = _4500_ ^ _4499_ /*32649*/;
  assign _4501_ = _4500_ & _4499_ /*32648*/;
  assign _4502_ = inv_21[5] & r_20[16] /*32647*/;
  assign _4503_ = _4501_ | _4502_ /*32646*/;
  assign _4504_ = inv_21[6] ^ r_20[17] /*32644*/;
  assign sum_21[6] = _4504_ ^ _4503_ /*32643*/;
  assign _4505_ = _4504_ & _4503_ /*32642*/;
  assign _4506_ = inv_21[6] & r_20[17] /*32641*/;
  assign _4507_ = _4505_ | _4506_ /*32640*/;
  assign _4508_ = inv_21[7] ^ r_20[18] /*32638*/;
  assign sum_21[7] = _4508_ ^ _4507_ /*32637*/;
  assign _4509_ = _4508_ & _4507_ /*32636*/;
  assign _4510_ = inv_21[7] & r_20[18] /*32635*/;
  assign _4511_ = _4509_ | _4510_ /*32634*/;
  assign _4512_ = inv_21[8] ^ r_20[19] /*32632*/;
  assign sum_21[8] = _4512_ ^ _4511_ /*32631*/;
  assign _4513_ = _4512_ & _4511_ /*32630*/;
  assign _4514_ = inv_21[8] & r_20[19] /*32629*/;
  assign _4515_ = _4513_ | _4514_ /*32628*/;
  assign _4516_ = inv_21[9] ^ r_20[20] /*32626*/;
  assign sum_21[9] = _4516_ ^ _4515_ /*32625*/;
  assign _4517_ = _4516_ & _4515_ /*32624*/;
  assign _4518_ = inv_21[9] & r_20[20] /*32623*/;
  assign _4519_ = _4517_ | _4518_ /*32622*/;
  assign _4520_ = inv_21[10] ^ r_20[21] /*32620*/;
  assign sum_21[10] = _4520_ ^ _4519_ /*32619*/;
  assign _4521_ = _4520_ & _4519_ /*32618*/;
  assign _4522_ = inv_21[10] & r_20[21] /*32617*/;
  assign _4523_ = _4521_ | _4522_ /*32616*/;
  assign _4524_ = inv_21[11] ^ r_20[22] /*32614*/;
  assign sum_21[11] = _4524_ ^ _4523_ /*32613*/;
  assign _4525_ = _4524_ & _4523_ /*32612*/;
  assign _4526_ = inv_21[11] & r_20[22] /*32611*/;
  assign _4527_ = _4525_ | _4526_ /*32610*/;
  assign _4528_ = inv_21[12] ^ r_20[23] /*32608*/;
  assign sum_21[12] = _4528_ ^ _4527_ /*32607*/;
  assign _4529_ = _4528_ & _4527_ /*32606*/;
  assign _4530_ = inv_21[12] & r_20[23] /*32605*/;
  assign _4531_ = _4529_ | _4530_ /*32604*/;
  assign _4532_ = inv_21[13] ^ r_20[24] /*32602*/;
  assign sum_21[13] = _4532_ ^ _4531_ /*32601*/;
  assign _4533_ = _4532_ & _4531_ /*32600*/;
  assign _4534_ = inv_21[13] & r_20[24] /*32599*/;
  assign _4535_ = _4533_ | _4534_ /*32598*/;
  assign _4536_ = inv_21[14] ^ r_20[25] /*32596*/;
  assign sum_21[14] = _4536_ ^ _4535_ /*32595*/;
  assign _4537_ = _4536_ & _4535_ /*32594*/;
  assign _4538_ = inv_21[14] & r_20[25] /*32593*/;
  assign _4539_ = _4537_ | _4538_ /*32592*/;
  assign _4540_ = inv_21[15] ^ r_20[26] /*32590*/;
  assign sum_21[15] = _4540_ ^ _4539_ /*32589*/;
  assign _4541_ = _4540_ & _4539_ /*32588*/;
  assign _4542_ = inv_21[15] & r_20[26] /*32587*/;
  assign _4543_ = _4541_ | _4542_ /*32586*/;
  assign _4544_ = inv_21[16] ^ r_20[27] /*32584*/;
  assign sum_21[16] = _4544_ ^ _4543_ /*32583*/;
  assign _4545_ = _4544_ & _4543_ /*32582*/;
  assign _4546_ = inv_21[16] & r_20[27] /*32581*/;
  assign _4547_ = _4545_ | _4546_ /*32580*/;
  assign _4548_ = inv_21[17] ^ r_20[28] /*32578*/;
  assign sum_21[17] = _4548_ ^ _4547_ /*32577*/;
  assign _4549_ = _4548_ & _4547_ /*32576*/;
  assign _4550_ = inv_21[17] & r_20[28] /*32575*/;
  assign _4551_ = _4549_ | _4550_ /*32574*/;
  assign _4552_ = inv_21[18] ^ r_20[29] /*32572*/;
  assign sum_21[18] = _4552_ ^ _4551_ /*32571*/;
  assign _4553_ = _4552_ & _4551_ /*32570*/;
  assign _4554_ = inv_21[18] & r_20[29] /*32569*/;
  assign _4555_ = _4553_ | _4554_ /*32568*/;
  assign _4556_ = inv_21[19] ^ r_20[30] /*32566*/;
  assign sum_21[19] = _4556_ ^ _4555_ /*32565*/;
  assign _4557_ = _4556_ & _4555_ /*32564*/;
  assign _4558_ = inv_21[19] & r_20[30] /*32563*/;
  assign _4559_ = _4557_ | _4558_ /*32562*/;
  assign _4560_ = inv_21[20] ^ r_20[31] /*32560*/;
  assign sum_21[20] = _4560_ ^ _4559_ /*32559*/;
  assign _4561_ = _4560_ & _4559_ /*32558*/;
  assign _4562_ = inv_21[20] & r_20[31] /*32557*/;
  assign _4563_ = _4561_ | _4562_ /*32556*/;
  assign _4564_ = inv_21[21] ^ r_20[32] /*32554*/;
  assign sum_21[21] = _4564_ ^ _4563_ /*32553*/;
  assign _4565_ = _4564_ & _4563_ /*32552*/;
  assign _4566_ = inv_21[21] & r_20[32] /*32551*/;
  assign _4567_ = _4565_ | _4566_ /*32550*/;
  assign _4568_ = inv_21[22] ^ r_20[33] /*32548*/;
  assign sum_21[22] = _4568_ ^ _4567_ /*32547*/;
  assign _4569_ = _4568_ & _4567_ /*32546*/;
  assign _4570_ = inv_21[22] & r_20[33] /*32545*/;
  assign _4571_ = _4569_ | _4570_ /*32544*/;
  assign _4572_ = inv_21[23] ^ r_20[34] /*32542*/;
  assign sum_21[23] = _4572_ ^ _4571_ /*32541*/;
  assign _4573_ = _4572_ & _4571_ /*32540*/;
  assign _4574_ = inv_21[23] & r_20[34] /*32539*/;
  assign _4575_ = _4573_ | _4574_ /*32538*/;
  assign _4576_ = inv_21[24] ^ r_20[35] /*32536*/;
  assign sum_21[24] = _4576_ ^ _4575_ /*32535*/;
  assign _4577_ = _4576_ & _4575_ /*32534*/;
  assign _4578_ = inv_21[24] & r_20[35] /*32533*/;
  assign _4579_ = _4577_ | _4578_ /*32532*/;
  assign _4580_ = inv_21[25] ^ r_20[36] /*32530*/;
  assign sum_21[25] = _4580_ ^ _4579_ /*32529*/;
  assign _4581_ = _4580_ & _4579_ /*32528*/;
  assign _4582_ = inv_21[25] & r_20[36] /*32527*/;
  assign _4583_ = _4581_ | _4582_ /*32526*/;
  assign _4584_ = inv_21[26] ^ r_20[37] /*32524*/;
  assign sum_21[26] = _4584_ ^ _4583_ /*32523*/;
  assign _4585_ = _4584_ & _4583_ /*32522*/;
  assign _4586_ = inv_21[26] & r_20[37] /*32521*/;
  assign _4587_ = _4585_ | _4586_ /*32520*/;
  assign _4588_ = inv_21[27] ^ r_20[38] /*32518*/;
  assign sum_21[27] = _4588_ ^ _4587_ /*32517*/;
  assign _4589_ = _4588_ & _4587_ /*32516*/;
  assign _4590_ = inv_21[27] & r_20[38] /*32515*/;
  assign _4591_ = _4589_ | _4590_ /*32514*/;
  assign _4592_ = inv_21[28] ^ r_20[39] /*32512*/;
  assign sum_21[28] = _4592_ ^ _4591_ /*32511*/;
  assign _4593_ = _4592_ & _4591_ /*32510*/;
  assign _4594_ = inv_21[28] & r_20[39] /*32509*/;
  assign _4595_ = _4593_ | _4594_ /*32508*/;
  assign _4596_ = inv_21[29] ^ r_20[40] /*32506*/;
  assign sum_21[29] = _4596_ ^ _4595_ /*32505*/;
  assign _4597_ = _4596_ & _4595_ /*32504*/;
  assign _4598_ = inv_21[29] & r_20[40] /*32503*/;
  assign _4599_ = _4597_ | _4598_ /*32502*/;
  assign _4600_ = inv_21[30] ^ r_20[41] /*32500*/;
  assign sum_21[30] = _4600_ ^ _4599_ /*32499*/;
  assign _4601_ = _4600_ & _4599_ /*32498*/;
  assign _4602_ = inv_21[30] & r_20[41] /*32497*/;
  assign _4603_ = _4601_ | _4602_ /*32496*/;
  assign _4604_ = inv_21[31] ^ r_20[42] /*32494*/;
  assign sum_21[31] = _4604_ ^ _4603_ /*32493*/;
  assign _4605_ = _4604_ & _4603_ /*32492*/;
  assign _4606_ = inv_21[31] & r_20[42] /*32491*/;
  assign _4607_ = _4605_ | _4606_ /*32490*/;
  assign q[11] = ~sum_21[31] /*32517*/;
  assign m_21[0] = r_20[11] /*32516*/;
  assign m_21[1] = r_20[12] /*32515*/;
  assign m_21[2] = r_20[13] /*32514*/;
  assign m_21[3] = r_20[14] /*32513*/;
  assign m_21[4] = r_20[15] /*32512*/;
  assign m_21[5] = r_20[16] /*32511*/;
  assign m_21[6] = r_20[17] /*32510*/;
  assign m_21[7] = r_20[18] /*32509*/;
  assign m_21[8] = r_20[19] /*32508*/;
  assign m_21[9] = r_20[20] /*32507*/;
  assign m_21[10] = r_20[21] /*32506*/;
  assign m_21[11] = r_20[22] /*32505*/;
  assign m_21[12] = r_20[23] /*32504*/;
  assign m_21[13] = r_20[24] /*32503*/;
  assign m_21[14] = r_20[25] /*32502*/;
  assign m_21[15] = r_20[26] /*32501*/;
  assign m_21[16] = r_20[27] /*32500*/;
  assign m_21[17] = r_20[28] /*32499*/;
  assign m_21[18] = r_20[29] /*32498*/;
  assign m_21[19] = r_20[30] /*32497*/;
  assign m_21[20] = r_20[31] /*32496*/;
  assign m_21[21] = r_20[32] /*32495*/;
  assign m_21[22] = r_20[33] /*32494*/;
  assign m_21[23] = r_20[34] /*32493*/;
  assign m_21[24] = r_20[35] /*32492*/;
  assign m_21[25] = r_20[36] /*32491*/;
  assign m_21[26] = r_20[37] /*32490*/;
  assign m_21[27] = r_20[38] /*32489*/;
  assign m_21[28] = r_20[39] /*32488*/;
  assign m_21[29] = r_20[40] /*32487*/;
  assign m_21[30] = r_20[41] /*32486*/;
  assign m_21[31] = r_20[42] /*32485*/;
  assign _4608_ = ~q[11] /*32483*/;
  assign _4609_ = sum_21[0] & q[11] /*32482*/;
  assign _4610_ = m_21[0] & _4608_ /*32481*/;
  assign r_21[11] = _4610_ | _4609_ /*32480*/;
  assign _4611_ = ~q[11] /*32479*/;
  assign _4612_ = sum_21[1] & q[11] /*32478*/;
  assign _4613_ = m_21[1] & _4611_ /*32477*/;
  assign r_21[12] = _4613_ | _4612_ /*32476*/;
  assign _4614_ = ~q[11] /*32475*/;
  assign _4615_ = sum_21[2] & q[11] /*32474*/;
  assign _4616_ = m_21[2] & _4614_ /*32473*/;
  assign r_21[13] = _4616_ | _4615_ /*32472*/;
  assign _4617_ = ~q[11] /*32471*/;
  assign _4618_ = sum_21[3] & q[11] /*32470*/;
  assign _4619_ = m_21[3] & _4617_ /*32469*/;
  assign r_21[14] = _4619_ | _4618_ /*32468*/;
  assign _4620_ = ~q[11] /*32467*/;
  assign _4621_ = sum_21[4] & q[11] /*32466*/;
  assign _4622_ = m_21[4] & _4620_ /*32465*/;
  assign r_21[15] = _4622_ | _4621_ /*32464*/;
  assign _4623_ = ~q[11] /*32463*/;
  assign _4624_ = sum_21[5] & q[11] /*32462*/;
  assign _4625_ = m_21[5] & _4623_ /*32461*/;
  assign r_21[16] = _4625_ | _4624_ /*32460*/;
  assign _4626_ = ~q[11] /*32459*/;
  assign _4627_ = sum_21[6] & q[11] /*32458*/;
  assign _4628_ = m_21[6] & _4626_ /*32457*/;
  assign r_21[17] = _4628_ | _4627_ /*32456*/;
  assign _4629_ = ~q[11] /*32455*/;
  assign _4630_ = sum_21[7] & q[11] /*32454*/;
  assign _4631_ = m_21[7] & _4629_ /*32453*/;
  assign r_21[18] = _4631_ | _4630_ /*32452*/;
  assign _4632_ = ~q[11] /*32451*/;
  assign _4633_ = sum_21[8] & q[11] /*32450*/;
  assign _4634_ = m_21[8] & _4632_ /*32449*/;
  assign r_21[19] = _4634_ | _4633_ /*32448*/;
  assign _4635_ = ~q[11] /*32447*/;
  assign _4636_ = sum_21[9] & q[11] /*32446*/;
  assign _4637_ = m_21[9] & _4635_ /*32445*/;
  assign r_21[20] = _4637_ | _4636_ /*32444*/;
  assign _4638_ = ~q[11] /*32443*/;
  assign _4639_ = sum_21[10] & q[11] /*32442*/;
  assign _4640_ = m_21[10] & _4638_ /*32441*/;
  assign r_21[21] = _4640_ | _4639_ /*32440*/;
  assign _4641_ = ~q[11] /*32439*/;
  assign _4642_ = sum_21[11] & q[11] /*32438*/;
  assign _4643_ = m_21[11] & _4641_ /*32437*/;
  assign r_21[22] = _4643_ | _4642_ /*32436*/;
  assign _4644_ = ~q[11] /*32435*/;
  assign _4645_ = sum_21[12] & q[11] /*32434*/;
  assign _4646_ = m_21[12] & _4644_ /*32433*/;
  assign r_21[23] = _4646_ | _4645_ /*32432*/;
  assign _4647_ = ~q[11] /*32431*/;
  assign _4648_ = sum_21[13] & q[11] /*32430*/;
  assign _4649_ = m_21[13] & _4647_ /*32429*/;
  assign r_21[24] = _4649_ | _4648_ /*32428*/;
  assign _4650_ = ~q[11] /*32427*/;
  assign _4651_ = sum_21[14] & q[11] /*32426*/;
  assign _4652_ = m_21[14] & _4650_ /*32425*/;
  assign r_21[25] = _4652_ | _4651_ /*32424*/;
  assign _4653_ = ~q[11] /*32423*/;
  assign _4654_ = sum_21[15] & q[11] /*32422*/;
  assign _4655_ = m_21[15] & _4653_ /*32421*/;
  assign r_21[26] = _4655_ | _4654_ /*32420*/;
  assign _4656_ = ~q[11] /*32419*/;
  assign _4657_ = sum_21[16] & q[11] /*32418*/;
  assign _4658_ = m_21[16] & _4656_ /*32417*/;
  assign r_21[27] = _4658_ | _4657_ /*32416*/;
  assign _4659_ = ~q[11] /*32415*/;
  assign _4660_ = sum_21[17] & q[11] /*32414*/;
  assign _4661_ = m_21[17] & _4659_ /*32413*/;
  assign r_21[28] = _4661_ | _4660_ /*32412*/;
  assign _4662_ = ~q[11] /*32411*/;
  assign _4663_ = sum_21[18] & q[11] /*32410*/;
  assign _4664_ = m_21[18] & _4662_ /*32409*/;
  assign r_21[29] = _4664_ | _4663_ /*32408*/;
  assign _4665_ = ~q[11] /*32407*/;
  assign _4666_ = sum_21[19] & q[11] /*32406*/;
  assign _4667_ = m_21[19] & _4665_ /*32405*/;
  assign r_21[30] = _4667_ | _4666_ /*32404*/;
  assign _4668_ = ~q[11] /*32403*/;
  assign _4669_ = sum_21[20] & q[11] /*32402*/;
  assign _4670_ = m_21[20] & _4668_ /*32401*/;
  assign r_21[31] = _4670_ | _4669_ /*32400*/;
  assign _4671_ = ~q[11] /*32399*/;
  assign _4672_ = sum_21[21] & q[11] /*32398*/;
  assign _4673_ = m_21[21] & _4671_ /*32397*/;
  assign r_21[32] = _4673_ | _4672_ /*32396*/;
  assign _4674_ = ~q[11] /*32395*/;
  assign _4675_ = sum_21[22] & q[11] /*32394*/;
  assign _4676_ = m_21[22] & _4674_ /*32393*/;
  assign r_21[33] = _4676_ | _4675_ /*32392*/;
  assign _4677_ = ~q[11] /*32391*/;
  assign _4678_ = sum_21[23] & q[11] /*32390*/;
  assign _4679_ = m_21[23] & _4677_ /*32389*/;
  assign r_21[34] = _4679_ | _4678_ /*32388*/;
  assign _4680_ = ~q[11] /*32387*/;
  assign _4681_ = sum_21[24] & q[11] /*32386*/;
  assign _4682_ = m_21[24] & _4680_ /*32385*/;
  assign r_21[35] = _4682_ | _4681_ /*32384*/;
  assign _4683_ = ~q[11] /*32383*/;
  assign _4684_ = sum_21[25] & q[11] /*32382*/;
  assign _4685_ = m_21[25] & _4683_ /*32381*/;
  assign r_21[36] = _4685_ | _4684_ /*32380*/;
  assign _4686_ = ~q[11] /*32379*/;
  assign _4687_ = sum_21[26] & q[11] /*32378*/;
  assign _4688_ = m_21[26] & _4686_ /*32377*/;
  assign r_21[37] = _4688_ | _4687_ /*32376*/;
  assign _4689_ = ~q[11] /*32375*/;
  assign _4690_ = sum_21[27] & q[11] /*32374*/;
  assign _4691_ = m_21[27] & _4689_ /*32373*/;
  assign r_21[38] = _4691_ | _4690_ /*32372*/;
  assign _4692_ = ~q[11] /*32371*/;
  assign _4693_ = sum_21[28] & q[11] /*32370*/;
  assign _4694_ = m_21[28] & _4692_ /*32369*/;
  assign r_21[39] = _4694_ | _4693_ /*32368*/;
  assign _4695_ = ~q[11] /*32367*/;
  assign _4696_ = sum_21[29] & q[11] /*32366*/;
  assign _4697_ = m_21[29] & _4695_ /*32365*/;
  assign r_21[40] = _4697_ | _4696_ /*32364*/;
  assign _4698_ = ~q[11] /*32363*/;
  assign _4699_ = sum_21[30] & q[11] /*32362*/;
  assign _4700_ = m_21[30] & _4698_ /*32361*/;
  assign r_21[41] = _4700_ | _4699_ /*32360*/;
  assign _4701_ = ~q[11] /*32359*/;
  assign _4702_ = sum_21[31] & q[11] /*32358*/;
  assign _4703_ = m_21[31] & _4701_ /*32357*/;
  assign r_21[42] = _4703_ | _4702_ /*32356*/;
assign r_21[0]= r_20[0] /*32355*/;
assign r_21[1]= r_20[1] /*32354*/;
assign r_21[2]= r_20[2] /*32353*/;
assign r_21[3]= r_20[3] /*32352*/;
assign r_21[4]= r_20[4] /*32351*/;
assign r_21[5]= r_20[5] /*32350*/;
assign r_21[6]= r_20[6] /*32349*/;
assign r_21[7]= r_20[7] /*32348*/;
assign r_21[8]= r_20[8] /*32347*/;
assign r_21[9]= r_20[9] /*32346*/;
assign r_21[10]= r_20[10] /*32345*/;
  assign inv_22[0] = ~div[0] /*32264*/;
  assign inv_22[1] = ~div[1] /*32263*/;
  assign inv_22[2] = ~div[2] /*32262*/;
  assign inv_22[3] = ~div[3] /*32261*/;
  assign inv_22[4] = ~div[4] /*32260*/;
  assign inv_22[5] = ~div[5] /*32259*/;
  assign inv_22[6] = ~div[6] /*32258*/;
  assign inv_22[7] = ~div[7] /*32257*/;
  assign inv_22[8] = ~div[8] /*32256*/;
  assign inv_22[9] = ~div[9] /*32255*/;
  assign inv_22[10] = ~div[10] /*32254*/;
  assign inv_22[11] = ~div[11] /*32253*/;
  assign inv_22[12] = ~div[12] /*32252*/;
  assign inv_22[13] = ~div[13] /*32251*/;
  assign inv_22[14] = ~div[14] /*32250*/;
  assign inv_22[15] = ~div[15] /*32249*/;
  assign inv_22[16] = ~div[16] /*32248*/;
  assign inv_22[17] = ~div[17] /*32247*/;
  assign inv_22[18] = ~div[18] /*32246*/;
  assign inv_22[19] = ~div[19] /*32245*/;
  assign inv_22[20] = ~div[20] /*32244*/;
  assign inv_22[21] = ~div[21] /*32243*/;
  assign inv_22[22] = ~div[22] /*32242*/;
  assign inv_22[23] = ~div[23] /*32241*/;
  assign inv_22[24] = ~div[24] /*32240*/;
  assign inv_22[25] = ~div[25] /*32239*/;
  assign inv_22[26] = ~div[26] /*32238*/;
  assign inv_22[27] = ~div[27] /*32237*/;
  assign inv_22[28] = ~div[28] /*32236*/;
  assign inv_22[29] = ~div[29] /*32235*/;
  assign inv_22[30] = ~div[30] /*32234*/;
assign inv_22[31] = oneWire /*32233*/;
  assign _4704_ = inv_22[0] ^ r_21[10] /*32231*/;
  assign sum_22[0] = _4704_ ^ oneWire /*32230*/;
  assign _4705_ = _4704_ & oneWire /*32229*/;
  assign _4706_ = inv_22[0] & r_21[10] /*32228*/;
  assign _4707_ = _4705_ | _4706_ /*32227*/;
  assign _4708_ = inv_22[1] ^ r_21[11] /*32226*/;
  assign sum_22[1] = _4708_ ^ _4707_ /*32225*/;
  assign _4709_ = _4708_ & _4707_ /*32224*/;
  assign _4710_ = inv_22[1] & r_21[11] /*32223*/;
  assign _4711_ = _4709_ | _4710_ /*32222*/;
  assign _4712_ = inv_22[2] ^ r_21[12] /*32220*/;
  assign sum_22[2] = _4712_ ^ _4711_ /*32219*/;
  assign _4713_ = _4712_ & _4711_ /*32218*/;
  assign _4714_ = inv_22[2] & r_21[12] /*32217*/;
  assign _4715_ = _4713_ | _4714_ /*32216*/;
  assign _4716_ = inv_22[3] ^ r_21[13] /*32214*/;
  assign sum_22[3] = _4716_ ^ _4715_ /*32213*/;
  assign _4717_ = _4716_ & _4715_ /*32212*/;
  assign _4718_ = inv_22[3] & r_21[13] /*32211*/;
  assign _4719_ = _4717_ | _4718_ /*32210*/;
  assign _4720_ = inv_22[4] ^ r_21[14] /*32208*/;
  assign sum_22[4] = _4720_ ^ _4719_ /*32207*/;
  assign _4721_ = _4720_ & _4719_ /*32206*/;
  assign _4722_ = inv_22[4] & r_21[14] /*32205*/;
  assign _4723_ = _4721_ | _4722_ /*32204*/;
  assign _4724_ = inv_22[5] ^ r_21[15] /*32202*/;
  assign sum_22[5] = _4724_ ^ _4723_ /*32201*/;
  assign _4725_ = _4724_ & _4723_ /*32200*/;
  assign _4726_ = inv_22[5] & r_21[15] /*32199*/;
  assign _4727_ = _4725_ | _4726_ /*32198*/;
  assign _4728_ = inv_22[6] ^ r_21[16] /*32196*/;
  assign sum_22[6] = _4728_ ^ _4727_ /*32195*/;
  assign _4729_ = _4728_ & _4727_ /*32194*/;
  assign _4730_ = inv_22[6] & r_21[16] /*32193*/;
  assign _4731_ = _4729_ | _4730_ /*32192*/;
  assign _4732_ = inv_22[7] ^ r_21[17] /*32190*/;
  assign sum_22[7] = _4732_ ^ _4731_ /*32189*/;
  assign _4733_ = _4732_ & _4731_ /*32188*/;
  assign _4734_ = inv_22[7] & r_21[17] /*32187*/;
  assign _4735_ = _4733_ | _4734_ /*32186*/;
  assign _4736_ = inv_22[8] ^ r_21[18] /*32184*/;
  assign sum_22[8] = _4736_ ^ _4735_ /*32183*/;
  assign _4737_ = _4736_ & _4735_ /*32182*/;
  assign _4738_ = inv_22[8] & r_21[18] /*32181*/;
  assign _4739_ = _4737_ | _4738_ /*32180*/;
  assign _4740_ = inv_22[9] ^ r_21[19] /*32178*/;
  assign sum_22[9] = _4740_ ^ _4739_ /*32177*/;
  assign _4741_ = _4740_ & _4739_ /*32176*/;
  assign _4742_ = inv_22[9] & r_21[19] /*32175*/;
  assign _4743_ = _4741_ | _4742_ /*32174*/;
  assign _4744_ = inv_22[10] ^ r_21[20] /*32172*/;
  assign sum_22[10] = _4744_ ^ _4743_ /*32171*/;
  assign _4745_ = _4744_ & _4743_ /*32170*/;
  assign _4746_ = inv_22[10] & r_21[20] /*32169*/;
  assign _4747_ = _4745_ | _4746_ /*32168*/;
  assign _4748_ = inv_22[11] ^ r_21[21] /*32166*/;
  assign sum_22[11] = _4748_ ^ _4747_ /*32165*/;
  assign _4749_ = _4748_ & _4747_ /*32164*/;
  assign _4750_ = inv_22[11] & r_21[21] /*32163*/;
  assign _4751_ = _4749_ | _4750_ /*32162*/;
  assign _4752_ = inv_22[12] ^ r_21[22] /*32160*/;
  assign sum_22[12] = _4752_ ^ _4751_ /*32159*/;
  assign _4753_ = _4752_ & _4751_ /*32158*/;
  assign _4754_ = inv_22[12] & r_21[22] /*32157*/;
  assign _4755_ = _4753_ | _4754_ /*32156*/;
  assign _4756_ = inv_22[13] ^ r_21[23] /*32154*/;
  assign sum_22[13] = _4756_ ^ _4755_ /*32153*/;
  assign _4757_ = _4756_ & _4755_ /*32152*/;
  assign _4758_ = inv_22[13] & r_21[23] /*32151*/;
  assign _4759_ = _4757_ | _4758_ /*32150*/;
  assign _4760_ = inv_22[14] ^ r_21[24] /*32148*/;
  assign sum_22[14] = _4760_ ^ _4759_ /*32147*/;
  assign _4761_ = _4760_ & _4759_ /*32146*/;
  assign _4762_ = inv_22[14] & r_21[24] /*32145*/;
  assign _4763_ = _4761_ | _4762_ /*32144*/;
  assign _4764_ = inv_22[15] ^ r_21[25] /*32142*/;
  assign sum_22[15] = _4764_ ^ _4763_ /*32141*/;
  assign _4765_ = _4764_ & _4763_ /*32140*/;
  assign _4766_ = inv_22[15] & r_21[25] /*32139*/;
  assign _4767_ = _4765_ | _4766_ /*32138*/;
  assign _4768_ = inv_22[16] ^ r_21[26] /*32136*/;
  assign sum_22[16] = _4768_ ^ _4767_ /*32135*/;
  assign _4769_ = _4768_ & _4767_ /*32134*/;
  assign _4770_ = inv_22[16] & r_21[26] /*32133*/;
  assign _4771_ = _4769_ | _4770_ /*32132*/;
  assign _4772_ = inv_22[17] ^ r_21[27] /*32130*/;
  assign sum_22[17] = _4772_ ^ _4771_ /*32129*/;
  assign _4773_ = _4772_ & _4771_ /*32128*/;
  assign _4774_ = inv_22[17] & r_21[27] /*32127*/;
  assign _4775_ = _4773_ | _4774_ /*32126*/;
  assign _4776_ = inv_22[18] ^ r_21[28] /*32124*/;
  assign sum_22[18] = _4776_ ^ _4775_ /*32123*/;
  assign _4777_ = _4776_ & _4775_ /*32122*/;
  assign _4778_ = inv_22[18] & r_21[28] /*32121*/;
  assign _4779_ = _4777_ | _4778_ /*32120*/;
  assign _4780_ = inv_22[19] ^ r_21[29] /*32118*/;
  assign sum_22[19] = _4780_ ^ _4779_ /*32117*/;
  assign _4781_ = _4780_ & _4779_ /*32116*/;
  assign _4782_ = inv_22[19] & r_21[29] /*32115*/;
  assign _4783_ = _4781_ | _4782_ /*32114*/;
  assign _4784_ = inv_22[20] ^ r_21[30] /*32112*/;
  assign sum_22[20] = _4784_ ^ _4783_ /*32111*/;
  assign _4785_ = _4784_ & _4783_ /*32110*/;
  assign _4786_ = inv_22[20] & r_21[30] /*32109*/;
  assign _4787_ = _4785_ | _4786_ /*32108*/;
  assign _4788_ = inv_22[21] ^ r_21[31] /*32106*/;
  assign sum_22[21] = _4788_ ^ _4787_ /*32105*/;
  assign _4789_ = _4788_ & _4787_ /*32104*/;
  assign _4790_ = inv_22[21] & r_21[31] /*32103*/;
  assign _4791_ = _4789_ | _4790_ /*32102*/;
  assign _4792_ = inv_22[22] ^ r_21[32] /*32100*/;
  assign sum_22[22] = _4792_ ^ _4791_ /*32099*/;
  assign _4793_ = _4792_ & _4791_ /*32098*/;
  assign _4794_ = inv_22[22] & r_21[32] /*32097*/;
  assign _4795_ = _4793_ | _4794_ /*32096*/;
  assign _4796_ = inv_22[23] ^ r_21[33] /*32094*/;
  assign sum_22[23] = _4796_ ^ _4795_ /*32093*/;
  assign _4797_ = _4796_ & _4795_ /*32092*/;
  assign _4798_ = inv_22[23] & r_21[33] /*32091*/;
  assign _4799_ = _4797_ | _4798_ /*32090*/;
  assign _4800_ = inv_22[24] ^ r_21[34] /*32088*/;
  assign sum_22[24] = _4800_ ^ _4799_ /*32087*/;
  assign _4801_ = _4800_ & _4799_ /*32086*/;
  assign _4802_ = inv_22[24] & r_21[34] /*32085*/;
  assign _4803_ = _4801_ | _4802_ /*32084*/;
  assign _4804_ = inv_22[25] ^ r_21[35] /*32082*/;
  assign sum_22[25] = _4804_ ^ _4803_ /*32081*/;
  assign _4805_ = _4804_ & _4803_ /*32080*/;
  assign _4806_ = inv_22[25] & r_21[35] /*32079*/;
  assign _4807_ = _4805_ | _4806_ /*32078*/;
  assign _4808_ = inv_22[26] ^ r_21[36] /*32076*/;
  assign sum_22[26] = _4808_ ^ _4807_ /*32075*/;
  assign _4809_ = _4808_ & _4807_ /*32074*/;
  assign _4810_ = inv_22[26] & r_21[36] /*32073*/;
  assign _4811_ = _4809_ | _4810_ /*32072*/;
  assign _4812_ = inv_22[27] ^ r_21[37] /*32070*/;
  assign sum_22[27] = _4812_ ^ _4811_ /*32069*/;
  assign _4813_ = _4812_ & _4811_ /*32068*/;
  assign _4814_ = inv_22[27] & r_21[37] /*32067*/;
  assign _4815_ = _4813_ | _4814_ /*32066*/;
  assign _4816_ = inv_22[28] ^ r_21[38] /*32064*/;
  assign sum_22[28] = _4816_ ^ _4815_ /*32063*/;
  assign _4817_ = _4816_ & _4815_ /*32062*/;
  assign _4818_ = inv_22[28] & r_21[38] /*32061*/;
  assign _4819_ = _4817_ | _4818_ /*32060*/;
  assign _4820_ = inv_22[29] ^ r_21[39] /*32058*/;
  assign sum_22[29] = _4820_ ^ _4819_ /*32057*/;
  assign _4821_ = _4820_ & _4819_ /*32056*/;
  assign _4822_ = inv_22[29] & r_21[39] /*32055*/;
  assign _4823_ = _4821_ | _4822_ /*32054*/;
  assign _4824_ = inv_22[30] ^ r_21[40] /*32052*/;
  assign sum_22[30] = _4824_ ^ _4823_ /*32051*/;
  assign _4825_ = _4824_ & _4823_ /*32050*/;
  assign _4826_ = inv_22[30] & r_21[40] /*32049*/;
  assign _4827_ = _4825_ | _4826_ /*32048*/;
  assign _4828_ = inv_22[31] ^ r_21[41] /*32046*/;
  assign sum_22[31] = _4828_ ^ _4827_ /*32045*/;
  assign _4829_ = _4828_ & _4827_ /*32044*/;
  assign _4830_ = inv_22[31] & r_21[41] /*32043*/;
  assign _4831_ = _4829_ | _4830_ /*32042*/;
  assign q[10] = ~sum_22[31] /*32069*/;
  assign m_22[0] = r_21[10] /*32068*/;
  assign m_22[1] = r_21[11] /*32067*/;
  assign m_22[2] = r_21[12] /*32066*/;
  assign m_22[3] = r_21[13] /*32065*/;
  assign m_22[4] = r_21[14] /*32064*/;
  assign m_22[5] = r_21[15] /*32063*/;
  assign m_22[6] = r_21[16] /*32062*/;
  assign m_22[7] = r_21[17] /*32061*/;
  assign m_22[8] = r_21[18] /*32060*/;
  assign m_22[9] = r_21[19] /*32059*/;
  assign m_22[10] = r_21[20] /*32058*/;
  assign m_22[11] = r_21[21] /*32057*/;
  assign m_22[12] = r_21[22] /*32056*/;
  assign m_22[13] = r_21[23] /*32055*/;
  assign m_22[14] = r_21[24] /*32054*/;
  assign m_22[15] = r_21[25] /*32053*/;
  assign m_22[16] = r_21[26] /*32052*/;
  assign m_22[17] = r_21[27] /*32051*/;
  assign m_22[18] = r_21[28] /*32050*/;
  assign m_22[19] = r_21[29] /*32049*/;
  assign m_22[20] = r_21[30] /*32048*/;
  assign m_22[21] = r_21[31] /*32047*/;
  assign m_22[22] = r_21[32] /*32046*/;
  assign m_22[23] = r_21[33] /*32045*/;
  assign m_22[24] = r_21[34] /*32044*/;
  assign m_22[25] = r_21[35] /*32043*/;
  assign m_22[26] = r_21[36] /*32042*/;
  assign m_22[27] = r_21[37] /*32041*/;
  assign m_22[28] = r_21[38] /*32040*/;
  assign m_22[29] = r_21[39] /*32039*/;
  assign m_22[30] = r_21[40] /*32038*/;
  assign m_22[31] = r_21[41] /*32037*/;
  assign _4832_ = ~q[10] /*32035*/;
  assign _4833_ = sum_22[0] & q[10] /*32034*/;
  assign _4834_ = m_22[0] & _4832_ /*32033*/;
  assign r_22[10] = _4834_ | _4833_ /*32032*/;
  assign _4835_ = ~q[10] /*32031*/;
  assign _4836_ = sum_22[1] & q[10] /*32030*/;
  assign _4837_ = m_22[1] & _4835_ /*32029*/;
  assign r_22[11] = _4837_ | _4836_ /*32028*/;
  assign _4838_ = ~q[10] /*32027*/;
  assign _4839_ = sum_22[2] & q[10] /*32026*/;
  assign _4840_ = m_22[2] & _4838_ /*32025*/;
  assign r_22[12] = _4840_ | _4839_ /*32024*/;
  assign _4841_ = ~q[10] /*32023*/;
  assign _4842_ = sum_22[3] & q[10] /*32022*/;
  assign _4843_ = m_22[3] & _4841_ /*32021*/;
  assign r_22[13] = _4843_ | _4842_ /*32020*/;
  assign _4844_ = ~q[10] /*32019*/;
  assign _4845_ = sum_22[4] & q[10] /*32018*/;
  assign _4846_ = m_22[4] & _4844_ /*32017*/;
  assign r_22[14] = _4846_ | _4845_ /*32016*/;
  assign _4847_ = ~q[10] /*32015*/;
  assign _4848_ = sum_22[5] & q[10] /*32014*/;
  assign _4849_ = m_22[5] & _4847_ /*32013*/;
  assign r_22[15] = _4849_ | _4848_ /*32012*/;
  assign _4850_ = ~q[10] /*32011*/;
  assign _4851_ = sum_22[6] & q[10] /*32010*/;
  assign _4852_ = m_22[6] & _4850_ /*32009*/;
  assign r_22[16] = _4852_ | _4851_ /*32008*/;
  assign _4853_ = ~q[10] /*32007*/;
  assign _4854_ = sum_22[7] & q[10] /*32006*/;
  assign _4855_ = m_22[7] & _4853_ /*32005*/;
  assign r_22[17] = _4855_ | _4854_ /*32004*/;
  assign _4856_ = ~q[10] /*32003*/;
  assign _4857_ = sum_22[8] & q[10] /*32002*/;
  assign _4858_ = m_22[8] & _4856_ /*32001*/;
  assign r_22[18] = _4858_ | _4857_ /*32000*/;
  assign _4859_ = ~q[10] /*31999*/;
  assign _4860_ = sum_22[9] & q[10] /*31998*/;
  assign _4861_ = m_22[9] & _4859_ /*31997*/;
  assign r_22[19] = _4861_ | _4860_ /*31996*/;
  assign _4862_ = ~q[10] /*31995*/;
  assign _4863_ = sum_22[10] & q[10] /*31994*/;
  assign _4864_ = m_22[10] & _4862_ /*31993*/;
  assign r_22[20] = _4864_ | _4863_ /*31992*/;
  assign _4865_ = ~q[10] /*31991*/;
  assign _4866_ = sum_22[11] & q[10] /*31990*/;
  assign _4867_ = m_22[11] & _4865_ /*31989*/;
  assign r_22[21] = _4867_ | _4866_ /*31988*/;
  assign _4868_ = ~q[10] /*31987*/;
  assign _4869_ = sum_22[12] & q[10] /*31986*/;
  assign _4870_ = m_22[12] & _4868_ /*31985*/;
  assign r_22[22] = _4870_ | _4869_ /*31984*/;
  assign _4871_ = ~q[10] /*31983*/;
  assign _4872_ = sum_22[13] & q[10] /*31982*/;
  assign _4873_ = m_22[13] & _4871_ /*31981*/;
  assign r_22[23] = _4873_ | _4872_ /*31980*/;
  assign _4874_ = ~q[10] /*31979*/;
  assign _4875_ = sum_22[14] & q[10] /*31978*/;
  assign _4876_ = m_22[14] & _4874_ /*31977*/;
  assign r_22[24] = _4876_ | _4875_ /*31976*/;
  assign _4877_ = ~q[10] /*31975*/;
  assign _4878_ = sum_22[15] & q[10] /*31974*/;
  assign _4879_ = m_22[15] & _4877_ /*31973*/;
  assign r_22[25] = _4879_ | _4878_ /*31972*/;
  assign _4880_ = ~q[10] /*31971*/;
  assign _4881_ = sum_22[16] & q[10] /*31970*/;
  assign _4882_ = m_22[16] & _4880_ /*31969*/;
  assign r_22[26] = _4882_ | _4881_ /*31968*/;
  assign _4883_ = ~q[10] /*31967*/;
  assign _4884_ = sum_22[17] & q[10] /*31966*/;
  assign _4885_ = m_22[17] & _4883_ /*31965*/;
  assign r_22[27] = _4885_ | _4884_ /*31964*/;
  assign _4886_ = ~q[10] /*31963*/;
  assign _4887_ = sum_22[18] & q[10] /*31962*/;
  assign _4888_ = m_22[18] & _4886_ /*31961*/;
  assign r_22[28] = _4888_ | _4887_ /*31960*/;
  assign _4889_ = ~q[10] /*31959*/;
  assign _4890_ = sum_22[19] & q[10] /*31958*/;
  assign _4891_ = m_22[19] & _4889_ /*31957*/;
  assign r_22[29] = _4891_ | _4890_ /*31956*/;
  assign _4892_ = ~q[10] /*31955*/;
  assign _4893_ = sum_22[20] & q[10] /*31954*/;
  assign _4894_ = m_22[20] & _4892_ /*31953*/;
  assign r_22[30] = _4894_ | _4893_ /*31952*/;
  assign _4895_ = ~q[10] /*31951*/;
  assign _4896_ = sum_22[21] & q[10] /*31950*/;
  assign _4897_ = m_22[21] & _4895_ /*31949*/;
  assign r_22[31] = _4897_ | _4896_ /*31948*/;
  assign _4898_ = ~q[10] /*31947*/;
  assign _4899_ = sum_22[22] & q[10] /*31946*/;
  assign _4900_ = m_22[22] & _4898_ /*31945*/;
  assign r_22[32] = _4900_ | _4899_ /*31944*/;
  assign _4901_ = ~q[10] /*31943*/;
  assign _4902_ = sum_22[23] & q[10] /*31942*/;
  assign _4903_ = m_22[23] & _4901_ /*31941*/;
  assign r_22[33] = _4903_ | _4902_ /*31940*/;
  assign _4904_ = ~q[10] /*31939*/;
  assign _4905_ = sum_22[24] & q[10] /*31938*/;
  assign _4906_ = m_22[24] & _4904_ /*31937*/;
  assign r_22[34] = _4906_ | _4905_ /*31936*/;
  assign _4907_ = ~q[10] /*31935*/;
  assign _4908_ = sum_22[25] & q[10] /*31934*/;
  assign _4909_ = m_22[25] & _4907_ /*31933*/;
  assign r_22[35] = _4909_ | _4908_ /*31932*/;
  assign _4910_ = ~q[10] /*31931*/;
  assign _4911_ = sum_22[26] & q[10] /*31930*/;
  assign _4912_ = m_22[26] & _4910_ /*31929*/;
  assign r_22[36] = _4912_ | _4911_ /*31928*/;
  assign _4913_ = ~q[10] /*31927*/;
  assign _4914_ = sum_22[27] & q[10] /*31926*/;
  assign _4915_ = m_22[27] & _4913_ /*31925*/;
  assign r_22[37] = _4915_ | _4914_ /*31924*/;
  assign _4916_ = ~q[10] /*31923*/;
  assign _4917_ = sum_22[28] & q[10] /*31922*/;
  assign _4918_ = m_22[28] & _4916_ /*31921*/;
  assign r_22[38] = _4918_ | _4917_ /*31920*/;
  assign _4919_ = ~q[10] /*31919*/;
  assign _4920_ = sum_22[29] & q[10] /*31918*/;
  assign _4921_ = m_22[29] & _4919_ /*31917*/;
  assign r_22[39] = _4921_ | _4920_ /*31916*/;
  assign _4922_ = ~q[10] /*31915*/;
  assign _4923_ = sum_22[30] & q[10] /*31914*/;
  assign _4924_ = m_22[30] & _4922_ /*31913*/;
  assign r_22[40] = _4924_ | _4923_ /*31912*/;
  assign _4925_ = ~q[10] /*31911*/;
  assign _4926_ = sum_22[31] & q[10] /*31910*/;
  assign _4927_ = m_22[31] & _4925_ /*31909*/;
  assign r_22[41] = _4927_ | _4926_ /*31908*/;
assign r_22[0]= r_21[0] /*31907*/;
assign r_22[1]= r_21[1] /*31906*/;
assign r_22[2]= r_21[2] /*31905*/;
assign r_22[3]= r_21[3] /*31904*/;
assign r_22[4]= r_21[4] /*31903*/;
assign r_22[5]= r_21[5] /*31902*/;
assign r_22[6]= r_21[6] /*31901*/;
assign r_22[7]= r_21[7] /*31900*/;
assign r_22[8]= r_21[8] /*31899*/;
assign r_22[9]= r_21[9] /*31898*/;
  assign inv_23[0] = ~div[0] /*31816*/;
  assign inv_23[1] = ~div[1] /*31815*/;
  assign inv_23[2] = ~div[2] /*31814*/;
  assign inv_23[3] = ~div[3] /*31813*/;
  assign inv_23[4] = ~div[4] /*31812*/;
  assign inv_23[5] = ~div[5] /*31811*/;
  assign inv_23[6] = ~div[6] /*31810*/;
  assign inv_23[7] = ~div[7] /*31809*/;
  assign inv_23[8] = ~div[8] /*31808*/;
  assign inv_23[9] = ~div[9] /*31807*/;
  assign inv_23[10] = ~div[10] /*31806*/;
  assign inv_23[11] = ~div[11] /*31805*/;
  assign inv_23[12] = ~div[12] /*31804*/;
  assign inv_23[13] = ~div[13] /*31803*/;
  assign inv_23[14] = ~div[14] /*31802*/;
  assign inv_23[15] = ~div[15] /*31801*/;
  assign inv_23[16] = ~div[16] /*31800*/;
  assign inv_23[17] = ~div[17] /*31799*/;
  assign inv_23[18] = ~div[18] /*31798*/;
  assign inv_23[19] = ~div[19] /*31797*/;
  assign inv_23[20] = ~div[20] /*31796*/;
  assign inv_23[21] = ~div[21] /*31795*/;
  assign inv_23[22] = ~div[22] /*31794*/;
  assign inv_23[23] = ~div[23] /*31793*/;
  assign inv_23[24] = ~div[24] /*31792*/;
  assign inv_23[25] = ~div[25] /*31791*/;
  assign inv_23[26] = ~div[26] /*31790*/;
  assign inv_23[27] = ~div[27] /*31789*/;
  assign inv_23[28] = ~div[28] /*31788*/;
  assign inv_23[29] = ~div[29] /*31787*/;
  assign inv_23[30] = ~div[30] /*31786*/;
assign inv_23[31] = oneWire /*31785*/;
  assign _4928_ = inv_23[0] ^ r_22[9] /*31783*/;
  assign sum_23[0] = _4928_ ^ oneWire /*31782*/;
  assign _4929_ = _4928_ & oneWire /*31781*/;
  assign _4930_ = inv_23[0] & r_22[9] /*31780*/;
  assign _4931_ = _4929_ | _4930_ /*31779*/;
  assign _4932_ = inv_23[1] ^ r_22[10] /*31778*/;
  assign sum_23[1] = _4932_ ^ _4931_ /*31777*/;
  assign _4933_ = _4932_ & _4931_ /*31776*/;
  assign _4934_ = inv_23[1] & r_22[10] /*31775*/;
  assign _4935_ = _4933_ | _4934_ /*31774*/;
  assign _4936_ = inv_23[2] ^ r_22[11] /*31772*/;
  assign sum_23[2] = _4936_ ^ _4935_ /*31771*/;
  assign _4937_ = _4936_ & _4935_ /*31770*/;
  assign _4938_ = inv_23[2] & r_22[11] /*31769*/;
  assign _4939_ = _4937_ | _4938_ /*31768*/;
  assign _4940_ = inv_23[3] ^ r_22[12] /*31766*/;
  assign sum_23[3] = _4940_ ^ _4939_ /*31765*/;
  assign _4941_ = _4940_ & _4939_ /*31764*/;
  assign _4942_ = inv_23[3] & r_22[12] /*31763*/;
  assign _4943_ = _4941_ | _4942_ /*31762*/;
  assign _4944_ = inv_23[4] ^ r_22[13] /*31760*/;
  assign sum_23[4] = _4944_ ^ _4943_ /*31759*/;
  assign _4945_ = _4944_ & _4943_ /*31758*/;
  assign _4946_ = inv_23[4] & r_22[13] /*31757*/;
  assign _4947_ = _4945_ | _4946_ /*31756*/;
  assign _4948_ = inv_23[5] ^ r_22[14] /*31754*/;
  assign sum_23[5] = _4948_ ^ _4947_ /*31753*/;
  assign _4949_ = _4948_ & _4947_ /*31752*/;
  assign _4950_ = inv_23[5] & r_22[14] /*31751*/;
  assign _4951_ = _4949_ | _4950_ /*31750*/;
  assign _4952_ = inv_23[6] ^ r_22[15] /*31748*/;
  assign sum_23[6] = _4952_ ^ _4951_ /*31747*/;
  assign _4953_ = _4952_ & _4951_ /*31746*/;
  assign _4954_ = inv_23[6] & r_22[15] /*31745*/;
  assign _4955_ = _4953_ | _4954_ /*31744*/;
  assign _4956_ = inv_23[7] ^ r_22[16] /*31742*/;
  assign sum_23[7] = _4956_ ^ _4955_ /*31741*/;
  assign _4957_ = _4956_ & _4955_ /*31740*/;
  assign _4958_ = inv_23[7] & r_22[16] /*31739*/;
  assign _4959_ = _4957_ | _4958_ /*31738*/;
  assign _4960_ = inv_23[8] ^ r_22[17] /*31736*/;
  assign sum_23[8] = _4960_ ^ _4959_ /*31735*/;
  assign _4961_ = _4960_ & _4959_ /*31734*/;
  assign _4962_ = inv_23[8] & r_22[17] /*31733*/;
  assign _4963_ = _4961_ | _4962_ /*31732*/;
  assign _4964_ = inv_23[9] ^ r_22[18] /*31730*/;
  assign sum_23[9] = _4964_ ^ _4963_ /*31729*/;
  assign _4965_ = _4964_ & _4963_ /*31728*/;
  assign _4966_ = inv_23[9] & r_22[18] /*31727*/;
  assign _4967_ = _4965_ | _4966_ /*31726*/;
  assign _4968_ = inv_23[10] ^ r_22[19] /*31724*/;
  assign sum_23[10] = _4968_ ^ _4967_ /*31723*/;
  assign _4969_ = _4968_ & _4967_ /*31722*/;
  assign _4970_ = inv_23[10] & r_22[19] /*31721*/;
  assign _4971_ = _4969_ | _4970_ /*31720*/;
  assign _4972_ = inv_23[11] ^ r_22[20] /*31718*/;
  assign sum_23[11] = _4972_ ^ _4971_ /*31717*/;
  assign _4973_ = _4972_ & _4971_ /*31716*/;
  assign _4974_ = inv_23[11] & r_22[20] /*31715*/;
  assign _4975_ = _4973_ | _4974_ /*31714*/;
  assign _4976_ = inv_23[12] ^ r_22[21] /*31712*/;
  assign sum_23[12] = _4976_ ^ _4975_ /*31711*/;
  assign _4977_ = _4976_ & _4975_ /*31710*/;
  assign _4978_ = inv_23[12] & r_22[21] /*31709*/;
  assign _4979_ = _4977_ | _4978_ /*31708*/;
  assign _4980_ = inv_23[13] ^ r_22[22] /*31706*/;
  assign sum_23[13] = _4980_ ^ _4979_ /*31705*/;
  assign _4981_ = _4980_ & _4979_ /*31704*/;
  assign _4982_ = inv_23[13] & r_22[22] /*31703*/;
  assign _4983_ = _4981_ | _4982_ /*31702*/;
  assign _4984_ = inv_23[14] ^ r_22[23] /*31700*/;
  assign sum_23[14] = _4984_ ^ _4983_ /*31699*/;
  assign _4985_ = _4984_ & _4983_ /*31698*/;
  assign _4986_ = inv_23[14] & r_22[23] /*31697*/;
  assign _4987_ = _4985_ | _4986_ /*31696*/;
  assign _4988_ = inv_23[15] ^ r_22[24] /*31694*/;
  assign sum_23[15] = _4988_ ^ _4987_ /*31693*/;
  assign _4989_ = _4988_ & _4987_ /*31692*/;
  assign _4990_ = inv_23[15] & r_22[24] /*31691*/;
  assign _4991_ = _4989_ | _4990_ /*31690*/;
  assign _4992_ = inv_23[16] ^ r_22[25] /*31688*/;
  assign sum_23[16] = _4992_ ^ _4991_ /*31687*/;
  assign _4993_ = _4992_ & _4991_ /*31686*/;
  assign _4994_ = inv_23[16] & r_22[25] /*31685*/;
  assign _4995_ = _4993_ | _4994_ /*31684*/;
  assign _4996_ = inv_23[17] ^ r_22[26] /*31682*/;
  assign sum_23[17] = _4996_ ^ _4995_ /*31681*/;
  assign _4997_ = _4996_ & _4995_ /*31680*/;
  assign _4998_ = inv_23[17] & r_22[26] /*31679*/;
  assign _4999_ = _4997_ | _4998_ /*31678*/;
  assign _5000_ = inv_23[18] ^ r_22[27] /*31676*/;
  assign sum_23[18] = _5000_ ^ _4999_ /*31675*/;
  assign _5001_ = _5000_ & _4999_ /*31674*/;
  assign _5002_ = inv_23[18] & r_22[27] /*31673*/;
  assign _5003_ = _5001_ | _5002_ /*31672*/;
  assign _5004_ = inv_23[19] ^ r_22[28] /*31670*/;
  assign sum_23[19] = _5004_ ^ _5003_ /*31669*/;
  assign _5005_ = _5004_ & _5003_ /*31668*/;
  assign _5006_ = inv_23[19] & r_22[28] /*31667*/;
  assign _5007_ = _5005_ | _5006_ /*31666*/;
  assign _5008_ = inv_23[20] ^ r_22[29] /*31664*/;
  assign sum_23[20] = _5008_ ^ _5007_ /*31663*/;
  assign _5009_ = _5008_ & _5007_ /*31662*/;
  assign _5010_ = inv_23[20] & r_22[29] /*31661*/;
  assign _5011_ = _5009_ | _5010_ /*31660*/;
  assign _5012_ = inv_23[21] ^ r_22[30] /*31658*/;
  assign sum_23[21] = _5012_ ^ _5011_ /*31657*/;
  assign _5013_ = _5012_ & _5011_ /*31656*/;
  assign _5014_ = inv_23[21] & r_22[30] /*31655*/;
  assign _5015_ = _5013_ | _5014_ /*31654*/;
  assign _5016_ = inv_23[22] ^ r_22[31] /*31652*/;
  assign sum_23[22] = _5016_ ^ _5015_ /*31651*/;
  assign _5017_ = _5016_ & _5015_ /*31650*/;
  assign _5018_ = inv_23[22] & r_22[31] /*31649*/;
  assign _5019_ = _5017_ | _5018_ /*31648*/;
  assign _5020_ = inv_23[23] ^ r_22[32] /*31646*/;
  assign sum_23[23] = _5020_ ^ _5019_ /*31645*/;
  assign _5021_ = _5020_ & _5019_ /*31644*/;
  assign _5022_ = inv_23[23] & r_22[32] /*31643*/;
  assign _5023_ = _5021_ | _5022_ /*31642*/;
  assign _5024_ = inv_23[24] ^ r_22[33] /*31640*/;
  assign sum_23[24] = _5024_ ^ _5023_ /*31639*/;
  assign _5025_ = _5024_ & _5023_ /*31638*/;
  assign _5026_ = inv_23[24] & r_22[33] /*31637*/;
  assign _5027_ = _5025_ | _5026_ /*31636*/;
  assign _5028_ = inv_23[25] ^ r_22[34] /*31634*/;
  assign sum_23[25] = _5028_ ^ _5027_ /*31633*/;
  assign _5029_ = _5028_ & _5027_ /*31632*/;
  assign _5030_ = inv_23[25] & r_22[34] /*31631*/;
  assign _5031_ = _5029_ | _5030_ /*31630*/;
  assign _5032_ = inv_23[26] ^ r_22[35] /*31628*/;
  assign sum_23[26] = _5032_ ^ _5031_ /*31627*/;
  assign _5033_ = _5032_ & _5031_ /*31626*/;
  assign _5034_ = inv_23[26] & r_22[35] /*31625*/;
  assign _5035_ = _5033_ | _5034_ /*31624*/;
  assign _5036_ = inv_23[27] ^ r_22[36] /*31622*/;
  assign sum_23[27] = _5036_ ^ _5035_ /*31621*/;
  assign _5037_ = _5036_ & _5035_ /*31620*/;
  assign _5038_ = inv_23[27] & r_22[36] /*31619*/;
  assign _5039_ = _5037_ | _5038_ /*31618*/;
  assign _5040_ = inv_23[28] ^ r_22[37] /*31616*/;
  assign sum_23[28] = _5040_ ^ _5039_ /*31615*/;
  assign _5041_ = _5040_ & _5039_ /*31614*/;
  assign _5042_ = inv_23[28] & r_22[37] /*31613*/;
  assign _5043_ = _5041_ | _5042_ /*31612*/;
  assign _5044_ = inv_23[29] ^ r_22[38] /*31610*/;
  assign sum_23[29] = _5044_ ^ _5043_ /*31609*/;
  assign _5045_ = _5044_ & _5043_ /*31608*/;
  assign _5046_ = inv_23[29] & r_22[38] /*31607*/;
  assign _5047_ = _5045_ | _5046_ /*31606*/;
  assign _5048_ = inv_23[30] ^ r_22[39] /*31604*/;
  assign sum_23[30] = _5048_ ^ _5047_ /*31603*/;
  assign _5049_ = _5048_ & _5047_ /*31602*/;
  assign _5050_ = inv_23[30] & r_22[39] /*31601*/;
  assign _5051_ = _5049_ | _5050_ /*31600*/;
  assign _5052_ = inv_23[31] ^ r_22[40] /*31598*/;
  assign sum_23[31] = _5052_ ^ _5051_ /*31597*/;
  assign _5053_ = _5052_ & _5051_ /*31596*/;
  assign _5054_ = inv_23[31] & r_22[40] /*31595*/;
  assign _5055_ = _5053_ | _5054_ /*31594*/;
  assign q[9] = ~sum_23[31] /*31621*/;
  assign m_23[0] = r_22[9] /*31620*/;
  assign m_23[1] = r_22[10] /*31619*/;
  assign m_23[2] = r_22[11] /*31618*/;
  assign m_23[3] = r_22[12] /*31617*/;
  assign m_23[4] = r_22[13] /*31616*/;
  assign m_23[5] = r_22[14] /*31615*/;
  assign m_23[6] = r_22[15] /*31614*/;
  assign m_23[7] = r_22[16] /*31613*/;
  assign m_23[8] = r_22[17] /*31612*/;
  assign m_23[9] = r_22[18] /*31611*/;
  assign m_23[10] = r_22[19] /*31610*/;
  assign m_23[11] = r_22[20] /*31609*/;
  assign m_23[12] = r_22[21] /*31608*/;
  assign m_23[13] = r_22[22] /*31607*/;
  assign m_23[14] = r_22[23] /*31606*/;
  assign m_23[15] = r_22[24] /*31605*/;
  assign m_23[16] = r_22[25] /*31604*/;
  assign m_23[17] = r_22[26] /*31603*/;
  assign m_23[18] = r_22[27] /*31602*/;
  assign m_23[19] = r_22[28] /*31601*/;
  assign m_23[20] = r_22[29] /*31600*/;
  assign m_23[21] = r_22[30] /*31599*/;
  assign m_23[22] = r_22[31] /*31598*/;
  assign m_23[23] = r_22[32] /*31597*/;
  assign m_23[24] = r_22[33] /*31596*/;
  assign m_23[25] = r_22[34] /*31595*/;
  assign m_23[26] = r_22[35] /*31594*/;
  assign m_23[27] = r_22[36] /*31593*/;
  assign m_23[28] = r_22[37] /*31592*/;
  assign m_23[29] = r_22[38] /*31591*/;
  assign m_23[30] = r_22[39] /*31590*/;
  assign m_23[31] = r_22[40] /*31589*/;
  assign _5056_ = ~q[9] /*31587*/;
  assign _5057_ = sum_23[0] & q[9] /*31586*/;
  assign _5058_ = m_23[0] & _5056_ /*31585*/;
  assign r_23[9] = _5058_ | _5057_ /*31584*/;
  assign _5059_ = ~q[9] /*31583*/;
  assign _5060_ = sum_23[1] & q[9] /*31582*/;
  assign _5061_ = m_23[1] & _5059_ /*31581*/;
  assign r_23[10] = _5061_ | _5060_ /*31580*/;
  assign _5062_ = ~q[9] /*31579*/;
  assign _5063_ = sum_23[2] & q[9] /*31578*/;
  assign _5064_ = m_23[2] & _5062_ /*31577*/;
  assign r_23[11] = _5064_ | _5063_ /*31576*/;
  assign _5065_ = ~q[9] /*31575*/;
  assign _5066_ = sum_23[3] & q[9] /*31574*/;
  assign _5067_ = m_23[3] & _5065_ /*31573*/;
  assign r_23[12] = _5067_ | _5066_ /*31572*/;
  assign _5068_ = ~q[9] /*31571*/;
  assign _5069_ = sum_23[4] & q[9] /*31570*/;
  assign _5070_ = m_23[4] & _5068_ /*31569*/;
  assign r_23[13] = _5070_ | _5069_ /*31568*/;
  assign _5071_ = ~q[9] /*31567*/;
  assign _5072_ = sum_23[5] & q[9] /*31566*/;
  assign _5073_ = m_23[5] & _5071_ /*31565*/;
  assign r_23[14] = _5073_ | _5072_ /*31564*/;
  assign _5074_ = ~q[9] /*31563*/;
  assign _5075_ = sum_23[6] & q[9] /*31562*/;
  assign _5076_ = m_23[6] & _5074_ /*31561*/;
  assign r_23[15] = _5076_ | _5075_ /*31560*/;
  assign _5077_ = ~q[9] /*31559*/;
  assign _5078_ = sum_23[7] & q[9] /*31558*/;
  assign _5079_ = m_23[7] & _5077_ /*31557*/;
  assign r_23[16] = _5079_ | _5078_ /*31556*/;
  assign _5080_ = ~q[9] /*31555*/;
  assign _5081_ = sum_23[8] & q[9] /*31554*/;
  assign _5082_ = m_23[8] & _5080_ /*31553*/;
  assign r_23[17] = _5082_ | _5081_ /*31552*/;
  assign _5083_ = ~q[9] /*31551*/;
  assign _5084_ = sum_23[9] & q[9] /*31550*/;
  assign _5085_ = m_23[9] & _5083_ /*31549*/;
  assign r_23[18] = _5085_ | _5084_ /*31548*/;
  assign _5086_ = ~q[9] /*31547*/;
  assign _5087_ = sum_23[10] & q[9] /*31546*/;
  assign _5088_ = m_23[10] & _5086_ /*31545*/;
  assign r_23[19] = _5088_ | _5087_ /*31544*/;
  assign _5089_ = ~q[9] /*31543*/;
  assign _5090_ = sum_23[11] & q[9] /*31542*/;
  assign _5091_ = m_23[11] & _5089_ /*31541*/;
  assign r_23[20] = _5091_ | _5090_ /*31540*/;
  assign _5092_ = ~q[9] /*31539*/;
  assign _5093_ = sum_23[12] & q[9] /*31538*/;
  assign _5094_ = m_23[12] & _5092_ /*31537*/;
  assign r_23[21] = _5094_ | _5093_ /*31536*/;
  assign _5095_ = ~q[9] /*31535*/;
  assign _5096_ = sum_23[13] & q[9] /*31534*/;
  assign _5097_ = m_23[13] & _5095_ /*31533*/;
  assign r_23[22] = _5097_ | _5096_ /*31532*/;
  assign _5098_ = ~q[9] /*31531*/;
  assign _5099_ = sum_23[14] & q[9] /*31530*/;
  assign _5100_ = m_23[14] & _5098_ /*31529*/;
  assign r_23[23] = _5100_ | _5099_ /*31528*/;
  assign _5101_ = ~q[9] /*31527*/;
  assign _5102_ = sum_23[15] & q[9] /*31526*/;
  assign _5103_ = m_23[15] & _5101_ /*31525*/;
  assign r_23[24] = _5103_ | _5102_ /*31524*/;
  assign _5104_ = ~q[9] /*31523*/;
  assign _5105_ = sum_23[16] & q[9] /*31522*/;
  assign _5106_ = m_23[16] & _5104_ /*31521*/;
  assign r_23[25] = _5106_ | _5105_ /*31520*/;
  assign _5107_ = ~q[9] /*31519*/;
  assign _5108_ = sum_23[17] & q[9] /*31518*/;
  assign _5109_ = m_23[17] & _5107_ /*31517*/;
  assign r_23[26] = _5109_ | _5108_ /*31516*/;
  assign _5110_ = ~q[9] /*31515*/;
  assign _5111_ = sum_23[18] & q[9] /*31514*/;
  assign _5112_ = m_23[18] & _5110_ /*31513*/;
  assign r_23[27] = _5112_ | _5111_ /*31512*/;
  assign _5113_ = ~q[9] /*31511*/;
  assign _5114_ = sum_23[19] & q[9] /*31510*/;
  assign _5115_ = m_23[19] & _5113_ /*31509*/;
  assign r_23[28] = _5115_ | _5114_ /*31508*/;
  assign _5116_ = ~q[9] /*31507*/;
  assign _5117_ = sum_23[20] & q[9] /*31506*/;
  assign _5118_ = m_23[20] & _5116_ /*31505*/;
  assign r_23[29] = _5118_ | _5117_ /*31504*/;
  assign _5119_ = ~q[9] /*31503*/;
  assign _5120_ = sum_23[21] & q[9] /*31502*/;
  assign _5121_ = m_23[21] & _5119_ /*31501*/;
  assign r_23[30] = _5121_ | _5120_ /*31500*/;
  assign _5122_ = ~q[9] /*31499*/;
  assign _5123_ = sum_23[22] & q[9] /*31498*/;
  assign _5124_ = m_23[22] & _5122_ /*31497*/;
  assign r_23[31] = _5124_ | _5123_ /*31496*/;
  assign _5125_ = ~q[9] /*31495*/;
  assign _5126_ = sum_23[23] & q[9] /*31494*/;
  assign _5127_ = m_23[23] & _5125_ /*31493*/;
  assign r_23[32] = _5127_ | _5126_ /*31492*/;
  assign _5128_ = ~q[9] /*31491*/;
  assign _5129_ = sum_23[24] & q[9] /*31490*/;
  assign _5130_ = m_23[24] & _5128_ /*31489*/;
  assign r_23[33] = _5130_ | _5129_ /*31488*/;
  assign _5131_ = ~q[9] /*31487*/;
  assign _5132_ = sum_23[25] & q[9] /*31486*/;
  assign _5133_ = m_23[25] & _5131_ /*31485*/;
  assign r_23[34] = _5133_ | _5132_ /*31484*/;
  assign _5134_ = ~q[9] /*31483*/;
  assign _5135_ = sum_23[26] & q[9] /*31482*/;
  assign _5136_ = m_23[26] & _5134_ /*31481*/;
  assign r_23[35] = _5136_ | _5135_ /*31480*/;
  assign _5137_ = ~q[9] /*31479*/;
  assign _5138_ = sum_23[27] & q[9] /*31478*/;
  assign _5139_ = m_23[27] & _5137_ /*31477*/;
  assign r_23[36] = _5139_ | _5138_ /*31476*/;
  assign _5140_ = ~q[9] /*31475*/;
  assign _5141_ = sum_23[28] & q[9] /*31474*/;
  assign _5142_ = m_23[28] & _5140_ /*31473*/;
  assign r_23[37] = _5142_ | _5141_ /*31472*/;
  assign _5143_ = ~q[9] /*31471*/;
  assign _5144_ = sum_23[29] & q[9] /*31470*/;
  assign _5145_ = m_23[29] & _5143_ /*31469*/;
  assign r_23[38] = _5145_ | _5144_ /*31468*/;
  assign _5146_ = ~q[9] /*31467*/;
  assign _5147_ = sum_23[30] & q[9] /*31466*/;
  assign _5148_ = m_23[30] & _5146_ /*31465*/;
  assign r_23[39] = _5148_ | _5147_ /*31464*/;
  assign _5149_ = ~q[9] /*31463*/;
  assign _5150_ = sum_23[31] & q[9] /*31462*/;
  assign _5151_ = m_23[31] & _5149_ /*31461*/;
  assign r_23[40] = _5151_ | _5150_ /*31460*/;
assign r_23[0]= r_22[0] /*31459*/;
assign r_23[1]= r_22[1] /*31458*/;
assign r_23[2]= r_22[2] /*31457*/;
assign r_23[3]= r_22[3] /*31456*/;
assign r_23[4]= r_22[4] /*31455*/;
assign r_23[5]= r_22[5] /*31454*/;
assign r_23[6]= r_22[6] /*31453*/;
assign r_23[7]= r_22[7] /*31452*/;
assign r_23[8]= r_22[8] /*31451*/;
  assign inv_24[0] = ~div[0] /*31368*/;
  assign inv_24[1] = ~div[1] /*31367*/;
  assign inv_24[2] = ~div[2] /*31366*/;
  assign inv_24[3] = ~div[3] /*31365*/;
  assign inv_24[4] = ~div[4] /*31364*/;
  assign inv_24[5] = ~div[5] /*31363*/;
  assign inv_24[6] = ~div[6] /*31362*/;
  assign inv_24[7] = ~div[7] /*31361*/;
  assign inv_24[8] = ~div[8] /*31360*/;
  assign inv_24[9] = ~div[9] /*31359*/;
  assign inv_24[10] = ~div[10] /*31358*/;
  assign inv_24[11] = ~div[11] /*31357*/;
  assign inv_24[12] = ~div[12] /*31356*/;
  assign inv_24[13] = ~div[13] /*31355*/;
  assign inv_24[14] = ~div[14] /*31354*/;
  assign inv_24[15] = ~div[15] /*31353*/;
  assign inv_24[16] = ~div[16] /*31352*/;
  assign inv_24[17] = ~div[17] /*31351*/;
  assign inv_24[18] = ~div[18] /*31350*/;
  assign inv_24[19] = ~div[19] /*31349*/;
  assign inv_24[20] = ~div[20] /*31348*/;
  assign inv_24[21] = ~div[21] /*31347*/;
  assign inv_24[22] = ~div[22] /*31346*/;
  assign inv_24[23] = ~div[23] /*31345*/;
  assign inv_24[24] = ~div[24] /*31344*/;
  assign inv_24[25] = ~div[25] /*31343*/;
  assign inv_24[26] = ~div[26] /*31342*/;
  assign inv_24[27] = ~div[27] /*31341*/;
  assign inv_24[28] = ~div[28] /*31340*/;
  assign inv_24[29] = ~div[29] /*31339*/;
  assign inv_24[30] = ~div[30] /*31338*/;
assign inv_24[31] = oneWire /*31337*/;
  assign _5152_ = inv_24[0] ^ r_23[8] /*31335*/;
  assign sum_24[0] = _5152_ ^ oneWire /*31334*/;
  assign _5153_ = _5152_ & oneWire /*31333*/;
  assign _5154_ = inv_24[0] & r_23[8] /*31332*/;
  assign _5155_ = _5153_ | _5154_ /*31331*/;
  assign _5156_ = inv_24[1] ^ r_23[9] /*31330*/;
  assign sum_24[1] = _5156_ ^ _5155_ /*31329*/;
  assign _5157_ = _5156_ & _5155_ /*31328*/;
  assign _5158_ = inv_24[1] & r_23[9] /*31327*/;
  assign _5159_ = _5157_ | _5158_ /*31326*/;
  assign _5160_ = inv_24[2] ^ r_23[10] /*31324*/;
  assign sum_24[2] = _5160_ ^ _5159_ /*31323*/;
  assign _5161_ = _5160_ & _5159_ /*31322*/;
  assign _5162_ = inv_24[2] & r_23[10] /*31321*/;
  assign _5163_ = _5161_ | _5162_ /*31320*/;
  assign _5164_ = inv_24[3] ^ r_23[11] /*31318*/;
  assign sum_24[3] = _5164_ ^ _5163_ /*31317*/;
  assign _5165_ = _5164_ & _5163_ /*31316*/;
  assign _5166_ = inv_24[3] & r_23[11] /*31315*/;
  assign _5167_ = _5165_ | _5166_ /*31314*/;
  assign _5168_ = inv_24[4] ^ r_23[12] /*31312*/;
  assign sum_24[4] = _5168_ ^ _5167_ /*31311*/;
  assign _5169_ = _5168_ & _5167_ /*31310*/;
  assign _5170_ = inv_24[4] & r_23[12] /*31309*/;
  assign _5171_ = _5169_ | _5170_ /*31308*/;
  assign _5172_ = inv_24[5] ^ r_23[13] /*31306*/;
  assign sum_24[5] = _5172_ ^ _5171_ /*31305*/;
  assign _5173_ = _5172_ & _5171_ /*31304*/;
  assign _5174_ = inv_24[5] & r_23[13] /*31303*/;
  assign _5175_ = _5173_ | _5174_ /*31302*/;
  assign _5176_ = inv_24[6] ^ r_23[14] /*31300*/;
  assign sum_24[6] = _5176_ ^ _5175_ /*31299*/;
  assign _5177_ = _5176_ & _5175_ /*31298*/;
  assign _5178_ = inv_24[6] & r_23[14] /*31297*/;
  assign _5179_ = _5177_ | _5178_ /*31296*/;
  assign _5180_ = inv_24[7] ^ r_23[15] /*31294*/;
  assign sum_24[7] = _5180_ ^ _5179_ /*31293*/;
  assign _5181_ = _5180_ & _5179_ /*31292*/;
  assign _5182_ = inv_24[7] & r_23[15] /*31291*/;
  assign _5183_ = _5181_ | _5182_ /*31290*/;
  assign _5184_ = inv_24[8] ^ r_23[16] /*31288*/;
  assign sum_24[8] = _5184_ ^ _5183_ /*31287*/;
  assign _5185_ = _5184_ & _5183_ /*31286*/;
  assign _5186_ = inv_24[8] & r_23[16] /*31285*/;
  assign _5187_ = _5185_ | _5186_ /*31284*/;
  assign _5188_ = inv_24[9] ^ r_23[17] /*31282*/;
  assign sum_24[9] = _5188_ ^ _5187_ /*31281*/;
  assign _5189_ = _5188_ & _5187_ /*31280*/;
  assign _5190_ = inv_24[9] & r_23[17] /*31279*/;
  assign _5191_ = _5189_ | _5190_ /*31278*/;
  assign _5192_ = inv_24[10] ^ r_23[18] /*31276*/;
  assign sum_24[10] = _5192_ ^ _5191_ /*31275*/;
  assign _5193_ = _5192_ & _5191_ /*31274*/;
  assign _5194_ = inv_24[10] & r_23[18] /*31273*/;
  assign _5195_ = _5193_ | _5194_ /*31272*/;
  assign _5196_ = inv_24[11] ^ r_23[19] /*31270*/;
  assign sum_24[11] = _5196_ ^ _5195_ /*31269*/;
  assign _5197_ = _5196_ & _5195_ /*31268*/;
  assign _5198_ = inv_24[11] & r_23[19] /*31267*/;
  assign _5199_ = _5197_ | _5198_ /*31266*/;
  assign _5200_ = inv_24[12] ^ r_23[20] /*31264*/;
  assign sum_24[12] = _5200_ ^ _5199_ /*31263*/;
  assign _5201_ = _5200_ & _5199_ /*31262*/;
  assign _5202_ = inv_24[12] & r_23[20] /*31261*/;
  assign _5203_ = _5201_ | _5202_ /*31260*/;
  assign _5204_ = inv_24[13] ^ r_23[21] /*31258*/;
  assign sum_24[13] = _5204_ ^ _5203_ /*31257*/;
  assign _5205_ = _5204_ & _5203_ /*31256*/;
  assign _5206_ = inv_24[13] & r_23[21] /*31255*/;
  assign _5207_ = _5205_ | _5206_ /*31254*/;
  assign _5208_ = inv_24[14] ^ r_23[22] /*31252*/;
  assign sum_24[14] = _5208_ ^ _5207_ /*31251*/;
  assign _5209_ = _5208_ & _5207_ /*31250*/;
  assign _5210_ = inv_24[14] & r_23[22] /*31249*/;
  assign _5211_ = _5209_ | _5210_ /*31248*/;
  assign _5212_ = inv_24[15] ^ r_23[23] /*31246*/;
  assign sum_24[15] = _5212_ ^ _5211_ /*31245*/;
  assign _5213_ = _5212_ & _5211_ /*31244*/;
  assign _5214_ = inv_24[15] & r_23[23] /*31243*/;
  assign _5215_ = _5213_ | _5214_ /*31242*/;
  assign _5216_ = inv_24[16] ^ r_23[24] /*31240*/;
  assign sum_24[16] = _5216_ ^ _5215_ /*31239*/;
  assign _5217_ = _5216_ & _5215_ /*31238*/;
  assign _5218_ = inv_24[16] & r_23[24] /*31237*/;
  assign _5219_ = _5217_ | _5218_ /*31236*/;
  assign _5220_ = inv_24[17] ^ r_23[25] /*31234*/;
  assign sum_24[17] = _5220_ ^ _5219_ /*31233*/;
  assign _5221_ = _5220_ & _5219_ /*31232*/;
  assign _5222_ = inv_24[17] & r_23[25] /*31231*/;
  assign _5223_ = _5221_ | _5222_ /*31230*/;
  assign _5224_ = inv_24[18] ^ r_23[26] /*31228*/;
  assign sum_24[18] = _5224_ ^ _5223_ /*31227*/;
  assign _5225_ = _5224_ & _5223_ /*31226*/;
  assign _5226_ = inv_24[18] & r_23[26] /*31225*/;
  assign _5227_ = _5225_ | _5226_ /*31224*/;
  assign _5228_ = inv_24[19] ^ r_23[27] /*31222*/;
  assign sum_24[19] = _5228_ ^ _5227_ /*31221*/;
  assign _5229_ = _5228_ & _5227_ /*31220*/;
  assign _5230_ = inv_24[19] & r_23[27] /*31219*/;
  assign _5231_ = _5229_ | _5230_ /*31218*/;
  assign _5232_ = inv_24[20] ^ r_23[28] /*31216*/;
  assign sum_24[20] = _5232_ ^ _5231_ /*31215*/;
  assign _5233_ = _5232_ & _5231_ /*31214*/;
  assign _5234_ = inv_24[20] & r_23[28] /*31213*/;
  assign _5235_ = _5233_ | _5234_ /*31212*/;
  assign _5236_ = inv_24[21] ^ r_23[29] /*31210*/;
  assign sum_24[21] = _5236_ ^ _5235_ /*31209*/;
  assign _5237_ = _5236_ & _5235_ /*31208*/;
  assign _5238_ = inv_24[21] & r_23[29] /*31207*/;
  assign _5239_ = _5237_ | _5238_ /*31206*/;
  assign _5240_ = inv_24[22] ^ r_23[30] /*31204*/;
  assign sum_24[22] = _5240_ ^ _5239_ /*31203*/;
  assign _5241_ = _5240_ & _5239_ /*31202*/;
  assign _5242_ = inv_24[22] & r_23[30] /*31201*/;
  assign _5243_ = _5241_ | _5242_ /*31200*/;
  assign _5244_ = inv_24[23] ^ r_23[31] /*31198*/;
  assign sum_24[23] = _5244_ ^ _5243_ /*31197*/;
  assign _5245_ = _5244_ & _5243_ /*31196*/;
  assign _5246_ = inv_24[23] & r_23[31] /*31195*/;
  assign _5247_ = _5245_ | _5246_ /*31194*/;
  assign _5248_ = inv_24[24] ^ r_23[32] /*31192*/;
  assign sum_24[24] = _5248_ ^ _5247_ /*31191*/;
  assign _5249_ = _5248_ & _5247_ /*31190*/;
  assign _5250_ = inv_24[24] & r_23[32] /*31189*/;
  assign _5251_ = _5249_ | _5250_ /*31188*/;
  assign _5252_ = inv_24[25] ^ r_23[33] /*31186*/;
  assign sum_24[25] = _5252_ ^ _5251_ /*31185*/;
  assign _5253_ = _5252_ & _5251_ /*31184*/;
  assign _5254_ = inv_24[25] & r_23[33] /*31183*/;
  assign _5255_ = _5253_ | _5254_ /*31182*/;
  assign _5256_ = inv_24[26] ^ r_23[34] /*31180*/;
  assign sum_24[26] = _5256_ ^ _5255_ /*31179*/;
  assign _5257_ = _5256_ & _5255_ /*31178*/;
  assign _5258_ = inv_24[26] & r_23[34] /*31177*/;
  assign _5259_ = _5257_ | _5258_ /*31176*/;
  assign _5260_ = inv_24[27] ^ r_23[35] /*31174*/;
  assign sum_24[27] = _5260_ ^ _5259_ /*31173*/;
  assign _5261_ = _5260_ & _5259_ /*31172*/;
  assign _5262_ = inv_24[27] & r_23[35] /*31171*/;
  assign _5263_ = _5261_ | _5262_ /*31170*/;
  assign _5264_ = inv_24[28] ^ r_23[36] /*31168*/;
  assign sum_24[28] = _5264_ ^ _5263_ /*31167*/;
  assign _5265_ = _5264_ & _5263_ /*31166*/;
  assign _5266_ = inv_24[28] & r_23[36] /*31165*/;
  assign _5267_ = _5265_ | _5266_ /*31164*/;
  assign _5268_ = inv_24[29] ^ r_23[37] /*31162*/;
  assign sum_24[29] = _5268_ ^ _5267_ /*31161*/;
  assign _5269_ = _5268_ & _5267_ /*31160*/;
  assign _5270_ = inv_24[29] & r_23[37] /*31159*/;
  assign _5271_ = _5269_ | _5270_ /*31158*/;
  assign _5272_ = inv_24[30] ^ r_23[38] /*31156*/;
  assign sum_24[30] = _5272_ ^ _5271_ /*31155*/;
  assign _5273_ = _5272_ & _5271_ /*31154*/;
  assign _5274_ = inv_24[30] & r_23[38] /*31153*/;
  assign _5275_ = _5273_ | _5274_ /*31152*/;
  assign _5276_ = inv_24[31] ^ r_23[39] /*31150*/;
  assign sum_24[31] = _5276_ ^ _5275_ /*31149*/;
  assign _5277_ = _5276_ & _5275_ /*31148*/;
  assign _5278_ = inv_24[31] & r_23[39] /*31147*/;
  assign _5279_ = _5277_ | _5278_ /*31146*/;
  assign q[8] = ~sum_24[31] /*31173*/;
  assign m_24[0] = r_23[8] /*31172*/;
  assign m_24[1] = r_23[9] /*31171*/;
  assign m_24[2] = r_23[10] /*31170*/;
  assign m_24[3] = r_23[11] /*31169*/;
  assign m_24[4] = r_23[12] /*31168*/;
  assign m_24[5] = r_23[13] /*31167*/;
  assign m_24[6] = r_23[14] /*31166*/;
  assign m_24[7] = r_23[15] /*31165*/;
  assign m_24[8] = r_23[16] /*31164*/;
  assign m_24[9] = r_23[17] /*31163*/;
  assign m_24[10] = r_23[18] /*31162*/;
  assign m_24[11] = r_23[19] /*31161*/;
  assign m_24[12] = r_23[20] /*31160*/;
  assign m_24[13] = r_23[21] /*31159*/;
  assign m_24[14] = r_23[22] /*31158*/;
  assign m_24[15] = r_23[23] /*31157*/;
  assign m_24[16] = r_23[24] /*31156*/;
  assign m_24[17] = r_23[25] /*31155*/;
  assign m_24[18] = r_23[26] /*31154*/;
  assign m_24[19] = r_23[27] /*31153*/;
  assign m_24[20] = r_23[28] /*31152*/;
  assign m_24[21] = r_23[29] /*31151*/;
  assign m_24[22] = r_23[30] /*31150*/;
  assign m_24[23] = r_23[31] /*31149*/;
  assign m_24[24] = r_23[32] /*31148*/;
  assign m_24[25] = r_23[33] /*31147*/;
  assign m_24[26] = r_23[34] /*31146*/;
  assign m_24[27] = r_23[35] /*31145*/;
  assign m_24[28] = r_23[36] /*31144*/;
  assign m_24[29] = r_23[37] /*31143*/;
  assign m_24[30] = r_23[38] /*31142*/;
  assign m_24[31] = r_23[39] /*31141*/;
  assign _5280_ = ~q[8] /*31139*/;
  assign _5281_ = sum_24[0] & q[8] /*31138*/;
  assign _5282_ = m_24[0] & _5280_ /*31137*/;
  assign r_24[8] = _5282_ | _5281_ /*31136*/;
  assign _5283_ = ~q[8] /*31135*/;
  assign _5284_ = sum_24[1] & q[8] /*31134*/;
  assign _5285_ = m_24[1] & _5283_ /*31133*/;
  assign r_24[9] = _5285_ | _5284_ /*31132*/;
  assign _5286_ = ~q[8] /*31131*/;
  assign _5287_ = sum_24[2] & q[8] /*31130*/;
  assign _5288_ = m_24[2] & _5286_ /*31129*/;
  assign r_24[10] = _5288_ | _5287_ /*31128*/;
  assign _5289_ = ~q[8] /*31127*/;
  assign _5290_ = sum_24[3] & q[8] /*31126*/;
  assign _5291_ = m_24[3] & _5289_ /*31125*/;
  assign r_24[11] = _5291_ | _5290_ /*31124*/;
  assign _5292_ = ~q[8] /*31123*/;
  assign _5293_ = sum_24[4] & q[8] /*31122*/;
  assign _5294_ = m_24[4] & _5292_ /*31121*/;
  assign r_24[12] = _5294_ | _5293_ /*31120*/;
  assign _5295_ = ~q[8] /*31119*/;
  assign _5296_ = sum_24[5] & q[8] /*31118*/;
  assign _5297_ = m_24[5] & _5295_ /*31117*/;
  assign r_24[13] = _5297_ | _5296_ /*31116*/;
  assign _5298_ = ~q[8] /*31115*/;
  assign _5299_ = sum_24[6] & q[8] /*31114*/;
  assign _5300_ = m_24[6] & _5298_ /*31113*/;
  assign r_24[14] = _5300_ | _5299_ /*31112*/;
  assign _5301_ = ~q[8] /*31111*/;
  assign _5302_ = sum_24[7] & q[8] /*31110*/;
  assign _5303_ = m_24[7] & _5301_ /*31109*/;
  assign r_24[15] = _5303_ | _5302_ /*31108*/;
  assign _5304_ = ~q[8] /*31107*/;
  assign _5305_ = sum_24[8] & q[8] /*31106*/;
  assign _5306_ = m_24[8] & _5304_ /*31105*/;
  assign r_24[16] = _5306_ | _5305_ /*31104*/;
  assign _5307_ = ~q[8] /*31103*/;
  assign _5308_ = sum_24[9] & q[8] /*31102*/;
  assign _5309_ = m_24[9] & _5307_ /*31101*/;
  assign r_24[17] = _5309_ | _5308_ /*31100*/;
  assign _5310_ = ~q[8] /*31099*/;
  assign _5311_ = sum_24[10] & q[8] /*31098*/;
  assign _5312_ = m_24[10] & _5310_ /*31097*/;
  assign r_24[18] = _5312_ | _5311_ /*31096*/;
  assign _5313_ = ~q[8] /*31095*/;
  assign _5314_ = sum_24[11] & q[8] /*31094*/;
  assign _5315_ = m_24[11] & _5313_ /*31093*/;
  assign r_24[19] = _5315_ | _5314_ /*31092*/;
  assign _5316_ = ~q[8] /*31091*/;
  assign _5317_ = sum_24[12] & q[8] /*31090*/;
  assign _5318_ = m_24[12] & _5316_ /*31089*/;
  assign r_24[20] = _5318_ | _5317_ /*31088*/;
  assign _5319_ = ~q[8] /*31087*/;
  assign _5320_ = sum_24[13] & q[8] /*31086*/;
  assign _5321_ = m_24[13] & _5319_ /*31085*/;
  assign r_24[21] = _5321_ | _5320_ /*31084*/;
  assign _5322_ = ~q[8] /*31083*/;
  assign _5323_ = sum_24[14] & q[8] /*31082*/;
  assign _5324_ = m_24[14] & _5322_ /*31081*/;
  assign r_24[22] = _5324_ | _5323_ /*31080*/;
  assign _5325_ = ~q[8] /*31079*/;
  assign _5326_ = sum_24[15] & q[8] /*31078*/;
  assign _5327_ = m_24[15] & _5325_ /*31077*/;
  assign r_24[23] = _5327_ | _5326_ /*31076*/;
  assign _5328_ = ~q[8] /*31075*/;
  assign _5329_ = sum_24[16] & q[8] /*31074*/;
  assign _5330_ = m_24[16] & _5328_ /*31073*/;
  assign r_24[24] = _5330_ | _5329_ /*31072*/;
  assign _5331_ = ~q[8] /*31071*/;
  assign _5332_ = sum_24[17] & q[8] /*31070*/;
  assign _5333_ = m_24[17] & _5331_ /*31069*/;
  assign r_24[25] = _5333_ | _5332_ /*31068*/;
  assign _5334_ = ~q[8] /*31067*/;
  assign _5335_ = sum_24[18] & q[8] /*31066*/;
  assign _5336_ = m_24[18] & _5334_ /*31065*/;
  assign r_24[26] = _5336_ | _5335_ /*31064*/;
  assign _5337_ = ~q[8] /*31063*/;
  assign _5338_ = sum_24[19] & q[8] /*31062*/;
  assign _5339_ = m_24[19] & _5337_ /*31061*/;
  assign r_24[27] = _5339_ | _5338_ /*31060*/;
  assign _5340_ = ~q[8] /*31059*/;
  assign _5341_ = sum_24[20] & q[8] /*31058*/;
  assign _5342_ = m_24[20] & _5340_ /*31057*/;
  assign r_24[28] = _5342_ | _5341_ /*31056*/;
  assign _5343_ = ~q[8] /*31055*/;
  assign _5344_ = sum_24[21] & q[8] /*31054*/;
  assign _5345_ = m_24[21] & _5343_ /*31053*/;
  assign r_24[29] = _5345_ | _5344_ /*31052*/;
  assign _5346_ = ~q[8] /*31051*/;
  assign _5347_ = sum_24[22] & q[8] /*31050*/;
  assign _5348_ = m_24[22] & _5346_ /*31049*/;
  assign r_24[30] = _5348_ | _5347_ /*31048*/;
  assign _5349_ = ~q[8] /*31047*/;
  assign _5350_ = sum_24[23] & q[8] /*31046*/;
  assign _5351_ = m_24[23] & _5349_ /*31045*/;
  assign r_24[31] = _5351_ | _5350_ /*31044*/;
  assign _5352_ = ~q[8] /*31043*/;
  assign _5353_ = sum_24[24] & q[8] /*31042*/;
  assign _5354_ = m_24[24] & _5352_ /*31041*/;
  assign r_24[32] = _5354_ | _5353_ /*31040*/;
  assign _5355_ = ~q[8] /*31039*/;
  assign _5356_ = sum_24[25] & q[8] /*31038*/;
  assign _5357_ = m_24[25] & _5355_ /*31037*/;
  assign r_24[33] = _5357_ | _5356_ /*31036*/;
  assign _5358_ = ~q[8] /*31035*/;
  assign _5359_ = sum_24[26] & q[8] /*31034*/;
  assign _5360_ = m_24[26] & _5358_ /*31033*/;
  assign r_24[34] = _5360_ | _5359_ /*31032*/;
  assign _5361_ = ~q[8] /*31031*/;
  assign _5362_ = sum_24[27] & q[8] /*31030*/;
  assign _5363_ = m_24[27] & _5361_ /*31029*/;
  assign r_24[35] = _5363_ | _5362_ /*31028*/;
  assign _5364_ = ~q[8] /*31027*/;
  assign _5365_ = sum_24[28] & q[8] /*31026*/;
  assign _5366_ = m_24[28] & _5364_ /*31025*/;
  assign r_24[36] = _5366_ | _5365_ /*31024*/;
  assign _5367_ = ~q[8] /*31023*/;
  assign _5368_ = sum_24[29] & q[8] /*31022*/;
  assign _5369_ = m_24[29] & _5367_ /*31021*/;
  assign r_24[37] = _5369_ | _5368_ /*31020*/;
  assign _5370_ = ~q[8] /*31019*/;
  assign _5371_ = sum_24[30] & q[8] /*31018*/;
  assign _5372_ = m_24[30] & _5370_ /*31017*/;
  assign r_24[38] = _5372_ | _5371_ /*31016*/;
  assign _5373_ = ~q[8] /*31015*/;
  assign _5374_ = sum_24[31] & q[8] /*31014*/;
  assign _5375_ = m_24[31] & _5373_ /*31013*/;
  assign r_24[39] = _5375_ | _5374_ /*31012*/;
assign r_24[0]= r_23[0] /*31011*/;
assign r_24[1]= r_23[1] /*31010*/;
assign r_24[2]= r_23[2] /*31009*/;
assign r_24[3]= r_23[3] /*31008*/;
assign r_24[4]= r_23[4] /*31007*/;
assign r_24[5]= r_23[5] /*31006*/;
assign r_24[6]= r_23[6] /*31005*/;
assign r_24[7]= r_23[7] /*31004*/;
  assign inv_25[0] = ~div[0] /*30920*/;
  assign inv_25[1] = ~div[1] /*30919*/;
  assign inv_25[2] = ~div[2] /*30918*/;
  assign inv_25[3] = ~div[3] /*30917*/;
  assign inv_25[4] = ~div[4] /*30916*/;
  assign inv_25[5] = ~div[5] /*30915*/;
  assign inv_25[6] = ~div[6] /*30914*/;
  assign inv_25[7] = ~div[7] /*30913*/;
  assign inv_25[8] = ~div[8] /*30912*/;
  assign inv_25[9] = ~div[9] /*30911*/;
  assign inv_25[10] = ~div[10] /*30910*/;
  assign inv_25[11] = ~div[11] /*30909*/;
  assign inv_25[12] = ~div[12] /*30908*/;
  assign inv_25[13] = ~div[13] /*30907*/;
  assign inv_25[14] = ~div[14] /*30906*/;
  assign inv_25[15] = ~div[15] /*30905*/;
  assign inv_25[16] = ~div[16] /*30904*/;
  assign inv_25[17] = ~div[17] /*30903*/;
  assign inv_25[18] = ~div[18] /*30902*/;
  assign inv_25[19] = ~div[19] /*30901*/;
  assign inv_25[20] = ~div[20] /*30900*/;
  assign inv_25[21] = ~div[21] /*30899*/;
  assign inv_25[22] = ~div[22] /*30898*/;
  assign inv_25[23] = ~div[23] /*30897*/;
  assign inv_25[24] = ~div[24] /*30896*/;
  assign inv_25[25] = ~div[25] /*30895*/;
  assign inv_25[26] = ~div[26] /*30894*/;
  assign inv_25[27] = ~div[27] /*30893*/;
  assign inv_25[28] = ~div[28] /*30892*/;
  assign inv_25[29] = ~div[29] /*30891*/;
  assign inv_25[30] = ~div[30] /*30890*/;
assign inv_25[31] = oneWire /*30889*/;
  assign _5376_ = inv_25[0] ^ r_24[7] /*30887*/;
  assign sum_25[0] = _5376_ ^ oneWire /*30886*/;
  assign _5377_ = _5376_ & oneWire /*30885*/;
  assign _5378_ = inv_25[0] & r_24[7] /*30884*/;
  assign _5379_ = _5377_ | _5378_ /*30883*/;
  assign _5380_ = inv_25[1] ^ r_24[8] /*30882*/;
  assign sum_25[1] = _5380_ ^ _5379_ /*30881*/;
  assign _5381_ = _5380_ & _5379_ /*30880*/;
  assign _5382_ = inv_25[1] & r_24[8] /*30879*/;
  assign _5383_ = _5381_ | _5382_ /*30878*/;
  assign _5384_ = inv_25[2] ^ r_24[9] /*30876*/;
  assign sum_25[2] = _5384_ ^ _5383_ /*30875*/;
  assign _5385_ = _5384_ & _5383_ /*30874*/;
  assign _5386_ = inv_25[2] & r_24[9] /*30873*/;
  assign _5387_ = _5385_ | _5386_ /*30872*/;
  assign _5388_ = inv_25[3] ^ r_24[10] /*30870*/;
  assign sum_25[3] = _5388_ ^ _5387_ /*30869*/;
  assign _5389_ = _5388_ & _5387_ /*30868*/;
  assign _5390_ = inv_25[3] & r_24[10] /*30867*/;
  assign _5391_ = _5389_ | _5390_ /*30866*/;
  assign _5392_ = inv_25[4] ^ r_24[11] /*30864*/;
  assign sum_25[4] = _5392_ ^ _5391_ /*30863*/;
  assign _5393_ = _5392_ & _5391_ /*30862*/;
  assign _5394_ = inv_25[4] & r_24[11] /*30861*/;
  assign _5395_ = _5393_ | _5394_ /*30860*/;
  assign _5396_ = inv_25[5] ^ r_24[12] /*30858*/;
  assign sum_25[5] = _5396_ ^ _5395_ /*30857*/;
  assign _5397_ = _5396_ & _5395_ /*30856*/;
  assign _5398_ = inv_25[5] & r_24[12] /*30855*/;
  assign _5399_ = _5397_ | _5398_ /*30854*/;
  assign _5400_ = inv_25[6] ^ r_24[13] /*30852*/;
  assign sum_25[6] = _5400_ ^ _5399_ /*30851*/;
  assign _5401_ = _5400_ & _5399_ /*30850*/;
  assign _5402_ = inv_25[6] & r_24[13] /*30849*/;
  assign _5403_ = _5401_ | _5402_ /*30848*/;
  assign _5404_ = inv_25[7] ^ r_24[14] /*30846*/;
  assign sum_25[7] = _5404_ ^ _5403_ /*30845*/;
  assign _5405_ = _5404_ & _5403_ /*30844*/;
  assign _5406_ = inv_25[7] & r_24[14] /*30843*/;
  assign _5407_ = _5405_ | _5406_ /*30842*/;
  assign _5408_ = inv_25[8] ^ r_24[15] /*30840*/;
  assign sum_25[8] = _5408_ ^ _5407_ /*30839*/;
  assign _5409_ = _5408_ & _5407_ /*30838*/;
  assign _5410_ = inv_25[8] & r_24[15] /*30837*/;
  assign _5411_ = _5409_ | _5410_ /*30836*/;
  assign _5412_ = inv_25[9] ^ r_24[16] /*30834*/;
  assign sum_25[9] = _5412_ ^ _5411_ /*30833*/;
  assign _5413_ = _5412_ & _5411_ /*30832*/;
  assign _5414_ = inv_25[9] & r_24[16] /*30831*/;
  assign _5415_ = _5413_ | _5414_ /*30830*/;
  assign _5416_ = inv_25[10] ^ r_24[17] /*30828*/;
  assign sum_25[10] = _5416_ ^ _5415_ /*30827*/;
  assign _5417_ = _5416_ & _5415_ /*30826*/;
  assign _5418_ = inv_25[10] & r_24[17] /*30825*/;
  assign _5419_ = _5417_ | _5418_ /*30824*/;
  assign _5420_ = inv_25[11] ^ r_24[18] /*30822*/;
  assign sum_25[11] = _5420_ ^ _5419_ /*30821*/;
  assign _5421_ = _5420_ & _5419_ /*30820*/;
  assign _5422_ = inv_25[11] & r_24[18] /*30819*/;
  assign _5423_ = _5421_ | _5422_ /*30818*/;
  assign _5424_ = inv_25[12] ^ r_24[19] /*30816*/;
  assign sum_25[12] = _5424_ ^ _5423_ /*30815*/;
  assign _5425_ = _5424_ & _5423_ /*30814*/;
  assign _5426_ = inv_25[12] & r_24[19] /*30813*/;
  assign _5427_ = _5425_ | _5426_ /*30812*/;
  assign _5428_ = inv_25[13] ^ r_24[20] /*30810*/;
  assign sum_25[13] = _5428_ ^ _5427_ /*30809*/;
  assign _5429_ = _5428_ & _5427_ /*30808*/;
  assign _5430_ = inv_25[13] & r_24[20] /*30807*/;
  assign _5431_ = _5429_ | _5430_ /*30806*/;
  assign _5432_ = inv_25[14] ^ r_24[21] /*30804*/;
  assign sum_25[14] = _5432_ ^ _5431_ /*30803*/;
  assign _5433_ = _5432_ & _5431_ /*30802*/;
  assign _5434_ = inv_25[14] & r_24[21] /*30801*/;
  assign _5435_ = _5433_ | _5434_ /*30800*/;
  assign _5436_ = inv_25[15] ^ r_24[22] /*30798*/;
  assign sum_25[15] = _5436_ ^ _5435_ /*30797*/;
  assign _5437_ = _5436_ & _5435_ /*30796*/;
  assign _5438_ = inv_25[15] & r_24[22] /*30795*/;
  assign _5439_ = _5437_ | _5438_ /*30794*/;
  assign _5440_ = inv_25[16] ^ r_24[23] /*30792*/;
  assign sum_25[16] = _5440_ ^ _5439_ /*30791*/;
  assign _5441_ = _5440_ & _5439_ /*30790*/;
  assign _5442_ = inv_25[16] & r_24[23] /*30789*/;
  assign _5443_ = _5441_ | _5442_ /*30788*/;
  assign _5444_ = inv_25[17] ^ r_24[24] /*30786*/;
  assign sum_25[17] = _5444_ ^ _5443_ /*30785*/;
  assign _5445_ = _5444_ & _5443_ /*30784*/;
  assign _5446_ = inv_25[17] & r_24[24] /*30783*/;
  assign _5447_ = _5445_ | _5446_ /*30782*/;
  assign _5448_ = inv_25[18] ^ r_24[25] /*30780*/;
  assign sum_25[18] = _5448_ ^ _5447_ /*30779*/;
  assign _5449_ = _5448_ & _5447_ /*30778*/;
  assign _5450_ = inv_25[18] & r_24[25] /*30777*/;
  assign _5451_ = _5449_ | _5450_ /*30776*/;
  assign _5452_ = inv_25[19] ^ r_24[26] /*30774*/;
  assign sum_25[19] = _5452_ ^ _5451_ /*30773*/;
  assign _5453_ = _5452_ & _5451_ /*30772*/;
  assign _5454_ = inv_25[19] & r_24[26] /*30771*/;
  assign _5455_ = _5453_ | _5454_ /*30770*/;
  assign _5456_ = inv_25[20] ^ r_24[27] /*30768*/;
  assign sum_25[20] = _5456_ ^ _5455_ /*30767*/;
  assign _5457_ = _5456_ & _5455_ /*30766*/;
  assign _5458_ = inv_25[20] & r_24[27] /*30765*/;
  assign _5459_ = _5457_ | _5458_ /*30764*/;
  assign _5460_ = inv_25[21] ^ r_24[28] /*30762*/;
  assign sum_25[21] = _5460_ ^ _5459_ /*30761*/;
  assign _5461_ = _5460_ & _5459_ /*30760*/;
  assign _5462_ = inv_25[21] & r_24[28] /*30759*/;
  assign _5463_ = _5461_ | _5462_ /*30758*/;
  assign _5464_ = inv_25[22] ^ r_24[29] /*30756*/;
  assign sum_25[22] = _5464_ ^ _5463_ /*30755*/;
  assign _5465_ = _5464_ & _5463_ /*30754*/;
  assign _5466_ = inv_25[22] & r_24[29] /*30753*/;
  assign _5467_ = _5465_ | _5466_ /*30752*/;
  assign _5468_ = inv_25[23] ^ r_24[30] /*30750*/;
  assign sum_25[23] = _5468_ ^ _5467_ /*30749*/;
  assign _5469_ = _5468_ & _5467_ /*30748*/;
  assign _5470_ = inv_25[23] & r_24[30] /*30747*/;
  assign _5471_ = _5469_ | _5470_ /*30746*/;
  assign _5472_ = inv_25[24] ^ r_24[31] /*30744*/;
  assign sum_25[24] = _5472_ ^ _5471_ /*30743*/;
  assign _5473_ = _5472_ & _5471_ /*30742*/;
  assign _5474_ = inv_25[24] & r_24[31] /*30741*/;
  assign _5475_ = _5473_ | _5474_ /*30740*/;
  assign _5476_ = inv_25[25] ^ r_24[32] /*30738*/;
  assign sum_25[25] = _5476_ ^ _5475_ /*30737*/;
  assign _5477_ = _5476_ & _5475_ /*30736*/;
  assign _5478_ = inv_25[25] & r_24[32] /*30735*/;
  assign _5479_ = _5477_ | _5478_ /*30734*/;
  assign _5480_ = inv_25[26] ^ r_24[33] /*30732*/;
  assign sum_25[26] = _5480_ ^ _5479_ /*30731*/;
  assign _5481_ = _5480_ & _5479_ /*30730*/;
  assign _5482_ = inv_25[26] & r_24[33] /*30729*/;
  assign _5483_ = _5481_ | _5482_ /*30728*/;
  assign _5484_ = inv_25[27] ^ r_24[34] /*30726*/;
  assign sum_25[27] = _5484_ ^ _5483_ /*30725*/;
  assign _5485_ = _5484_ & _5483_ /*30724*/;
  assign _5486_ = inv_25[27] & r_24[34] /*30723*/;
  assign _5487_ = _5485_ | _5486_ /*30722*/;
  assign _5488_ = inv_25[28] ^ r_24[35] /*30720*/;
  assign sum_25[28] = _5488_ ^ _5487_ /*30719*/;
  assign _5489_ = _5488_ & _5487_ /*30718*/;
  assign _5490_ = inv_25[28] & r_24[35] /*30717*/;
  assign _5491_ = _5489_ | _5490_ /*30716*/;
  assign _5492_ = inv_25[29] ^ r_24[36] /*30714*/;
  assign sum_25[29] = _5492_ ^ _5491_ /*30713*/;
  assign _5493_ = _5492_ & _5491_ /*30712*/;
  assign _5494_ = inv_25[29] & r_24[36] /*30711*/;
  assign _5495_ = _5493_ | _5494_ /*30710*/;
  assign _5496_ = inv_25[30] ^ r_24[37] /*30708*/;
  assign sum_25[30] = _5496_ ^ _5495_ /*30707*/;
  assign _5497_ = _5496_ & _5495_ /*30706*/;
  assign _5498_ = inv_25[30] & r_24[37] /*30705*/;
  assign _5499_ = _5497_ | _5498_ /*30704*/;
  assign _5500_ = inv_25[31] ^ r_24[38] /*30702*/;
  assign sum_25[31] = _5500_ ^ _5499_ /*30701*/;
  assign _5501_ = _5500_ & _5499_ /*30700*/;
  assign _5502_ = inv_25[31] & r_24[38] /*30699*/;
  assign _5503_ = _5501_ | _5502_ /*30698*/;
  assign q[7] = ~sum_25[31] /*30725*/;
  assign m_25[0] = r_24[7] /*30724*/;
  assign m_25[1] = r_24[8] /*30723*/;
  assign m_25[2] = r_24[9] /*30722*/;
  assign m_25[3] = r_24[10] /*30721*/;
  assign m_25[4] = r_24[11] /*30720*/;
  assign m_25[5] = r_24[12] /*30719*/;
  assign m_25[6] = r_24[13] /*30718*/;
  assign m_25[7] = r_24[14] /*30717*/;
  assign m_25[8] = r_24[15] /*30716*/;
  assign m_25[9] = r_24[16] /*30715*/;
  assign m_25[10] = r_24[17] /*30714*/;
  assign m_25[11] = r_24[18] /*30713*/;
  assign m_25[12] = r_24[19] /*30712*/;
  assign m_25[13] = r_24[20] /*30711*/;
  assign m_25[14] = r_24[21] /*30710*/;
  assign m_25[15] = r_24[22] /*30709*/;
  assign m_25[16] = r_24[23] /*30708*/;
  assign m_25[17] = r_24[24] /*30707*/;
  assign m_25[18] = r_24[25] /*30706*/;
  assign m_25[19] = r_24[26] /*30705*/;
  assign m_25[20] = r_24[27] /*30704*/;
  assign m_25[21] = r_24[28] /*30703*/;
  assign m_25[22] = r_24[29] /*30702*/;
  assign m_25[23] = r_24[30] /*30701*/;
  assign m_25[24] = r_24[31] /*30700*/;
  assign m_25[25] = r_24[32] /*30699*/;
  assign m_25[26] = r_24[33] /*30698*/;
  assign m_25[27] = r_24[34] /*30697*/;
  assign m_25[28] = r_24[35] /*30696*/;
  assign m_25[29] = r_24[36] /*30695*/;
  assign m_25[30] = r_24[37] /*30694*/;
  assign m_25[31] = r_24[38] /*30693*/;
  assign _5504_ = ~q[7] /*30691*/;
  assign _5505_ = sum_25[0] & q[7] /*30690*/;
  assign _5506_ = m_25[0] & _5504_ /*30689*/;
  assign r_25[7] = _5506_ | _5505_ /*30688*/;
  assign _5507_ = ~q[7] /*30687*/;
  assign _5508_ = sum_25[1] & q[7] /*30686*/;
  assign _5509_ = m_25[1] & _5507_ /*30685*/;
  assign r_25[8] = _5509_ | _5508_ /*30684*/;
  assign _5510_ = ~q[7] /*30683*/;
  assign _5511_ = sum_25[2] & q[7] /*30682*/;
  assign _5512_ = m_25[2] & _5510_ /*30681*/;
  assign r_25[9] = _5512_ | _5511_ /*30680*/;
  assign _5513_ = ~q[7] /*30679*/;
  assign _5514_ = sum_25[3] & q[7] /*30678*/;
  assign _5515_ = m_25[3] & _5513_ /*30677*/;
  assign r_25[10] = _5515_ | _5514_ /*30676*/;
  assign _5516_ = ~q[7] /*30675*/;
  assign _5517_ = sum_25[4] & q[7] /*30674*/;
  assign _5518_ = m_25[4] & _5516_ /*30673*/;
  assign r_25[11] = _5518_ | _5517_ /*30672*/;
  assign _5519_ = ~q[7] /*30671*/;
  assign _5520_ = sum_25[5] & q[7] /*30670*/;
  assign _5521_ = m_25[5] & _5519_ /*30669*/;
  assign r_25[12] = _5521_ | _5520_ /*30668*/;
  assign _5522_ = ~q[7] /*30667*/;
  assign _5523_ = sum_25[6] & q[7] /*30666*/;
  assign _5524_ = m_25[6] & _5522_ /*30665*/;
  assign r_25[13] = _5524_ | _5523_ /*30664*/;
  assign _5525_ = ~q[7] /*30663*/;
  assign _5526_ = sum_25[7] & q[7] /*30662*/;
  assign _5527_ = m_25[7] & _5525_ /*30661*/;
  assign r_25[14] = _5527_ | _5526_ /*30660*/;
  assign _5528_ = ~q[7] /*30659*/;
  assign _5529_ = sum_25[8] & q[7] /*30658*/;
  assign _5530_ = m_25[8] & _5528_ /*30657*/;
  assign r_25[15] = _5530_ | _5529_ /*30656*/;
  assign _5531_ = ~q[7] /*30655*/;
  assign _5532_ = sum_25[9] & q[7] /*30654*/;
  assign _5533_ = m_25[9] & _5531_ /*30653*/;
  assign r_25[16] = _5533_ | _5532_ /*30652*/;
  assign _5534_ = ~q[7] /*30651*/;
  assign _5535_ = sum_25[10] & q[7] /*30650*/;
  assign _5536_ = m_25[10] & _5534_ /*30649*/;
  assign r_25[17] = _5536_ | _5535_ /*30648*/;
  assign _5537_ = ~q[7] /*30647*/;
  assign _5538_ = sum_25[11] & q[7] /*30646*/;
  assign _5539_ = m_25[11] & _5537_ /*30645*/;
  assign r_25[18] = _5539_ | _5538_ /*30644*/;
  assign _5540_ = ~q[7] /*30643*/;
  assign _5541_ = sum_25[12] & q[7] /*30642*/;
  assign _5542_ = m_25[12] & _5540_ /*30641*/;
  assign r_25[19] = _5542_ | _5541_ /*30640*/;
  assign _5543_ = ~q[7] /*30639*/;
  assign _5544_ = sum_25[13] & q[7] /*30638*/;
  assign _5545_ = m_25[13] & _5543_ /*30637*/;
  assign r_25[20] = _5545_ | _5544_ /*30636*/;
  assign _5546_ = ~q[7] /*30635*/;
  assign _5547_ = sum_25[14] & q[7] /*30634*/;
  assign _5548_ = m_25[14] & _5546_ /*30633*/;
  assign r_25[21] = _5548_ | _5547_ /*30632*/;
  assign _5549_ = ~q[7] /*30631*/;
  assign _5550_ = sum_25[15] & q[7] /*30630*/;
  assign _5551_ = m_25[15] & _5549_ /*30629*/;
  assign r_25[22] = _5551_ | _5550_ /*30628*/;
  assign _5552_ = ~q[7] /*30627*/;
  assign _5553_ = sum_25[16] & q[7] /*30626*/;
  assign _5554_ = m_25[16] & _5552_ /*30625*/;
  assign r_25[23] = _5554_ | _5553_ /*30624*/;
  assign _5555_ = ~q[7] /*30623*/;
  assign _5556_ = sum_25[17] & q[7] /*30622*/;
  assign _5557_ = m_25[17] & _5555_ /*30621*/;
  assign r_25[24] = _5557_ | _5556_ /*30620*/;
  assign _5558_ = ~q[7] /*30619*/;
  assign _5559_ = sum_25[18] & q[7] /*30618*/;
  assign _5560_ = m_25[18] & _5558_ /*30617*/;
  assign r_25[25] = _5560_ | _5559_ /*30616*/;
  assign _5561_ = ~q[7] /*30615*/;
  assign _5562_ = sum_25[19] & q[7] /*30614*/;
  assign _5563_ = m_25[19] & _5561_ /*30613*/;
  assign r_25[26] = _5563_ | _5562_ /*30612*/;
  assign _5564_ = ~q[7] /*30611*/;
  assign _5565_ = sum_25[20] & q[7] /*30610*/;
  assign _5566_ = m_25[20] & _5564_ /*30609*/;
  assign r_25[27] = _5566_ | _5565_ /*30608*/;
  assign _5567_ = ~q[7] /*30607*/;
  assign _5568_ = sum_25[21] & q[7] /*30606*/;
  assign _5569_ = m_25[21] & _5567_ /*30605*/;
  assign r_25[28] = _5569_ | _5568_ /*30604*/;
  assign _5570_ = ~q[7] /*30603*/;
  assign _5571_ = sum_25[22] & q[7] /*30602*/;
  assign _5572_ = m_25[22] & _5570_ /*30601*/;
  assign r_25[29] = _5572_ | _5571_ /*30600*/;
  assign _5573_ = ~q[7] /*30599*/;
  assign _5574_ = sum_25[23] & q[7] /*30598*/;
  assign _5575_ = m_25[23] & _5573_ /*30597*/;
  assign r_25[30] = _5575_ | _5574_ /*30596*/;
  assign _5576_ = ~q[7] /*30595*/;
  assign _5577_ = sum_25[24] & q[7] /*30594*/;
  assign _5578_ = m_25[24] & _5576_ /*30593*/;
  assign r_25[31] = _5578_ | _5577_ /*30592*/;
  assign _5579_ = ~q[7] /*30591*/;
  assign _5580_ = sum_25[25] & q[7] /*30590*/;
  assign _5581_ = m_25[25] & _5579_ /*30589*/;
  assign r_25[32] = _5581_ | _5580_ /*30588*/;
  assign _5582_ = ~q[7] /*30587*/;
  assign _5583_ = sum_25[26] & q[7] /*30586*/;
  assign _5584_ = m_25[26] & _5582_ /*30585*/;
  assign r_25[33] = _5584_ | _5583_ /*30584*/;
  assign _5585_ = ~q[7] /*30583*/;
  assign _5586_ = sum_25[27] & q[7] /*30582*/;
  assign _5587_ = m_25[27] & _5585_ /*30581*/;
  assign r_25[34] = _5587_ | _5586_ /*30580*/;
  assign _5588_ = ~q[7] /*30579*/;
  assign _5589_ = sum_25[28] & q[7] /*30578*/;
  assign _5590_ = m_25[28] & _5588_ /*30577*/;
  assign r_25[35] = _5590_ | _5589_ /*30576*/;
  assign _5591_ = ~q[7] /*30575*/;
  assign _5592_ = sum_25[29] & q[7] /*30574*/;
  assign _5593_ = m_25[29] & _5591_ /*30573*/;
  assign r_25[36] = _5593_ | _5592_ /*30572*/;
  assign _5594_ = ~q[7] /*30571*/;
  assign _5595_ = sum_25[30] & q[7] /*30570*/;
  assign _5596_ = m_25[30] & _5594_ /*30569*/;
  assign r_25[37] = _5596_ | _5595_ /*30568*/;
  assign _5597_ = ~q[7] /*30567*/;
  assign _5598_ = sum_25[31] & q[7] /*30566*/;
  assign _5599_ = m_25[31] & _5597_ /*30565*/;
  assign r_25[38] = _5599_ | _5598_ /*30564*/;
assign r_25[0]= r_24[0] /*30563*/;
assign r_25[1]= r_24[1] /*30562*/;
assign r_25[2]= r_24[2] /*30561*/;
assign r_25[3]= r_24[3] /*30560*/;
assign r_25[4]= r_24[4] /*30559*/;
assign r_25[5]= r_24[5] /*30558*/;
assign r_25[6]= r_24[6] /*30557*/;
  assign inv_26[0] = ~div[0] /*30472*/;
  assign inv_26[1] = ~div[1] /*30471*/;
  assign inv_26[2] = ~div[2] /*30470*/;
  assign inv_26[3] = ~div[3] /*30469*/;
  assign inv_26[4] = ~div[4] /*30468*/;
  assign inv_26[5] = ~div[5] /*30467*/;
  assign inv_26[6] = ~div[6] /*30466*/;
  assign inv_26[7] = ~div[7] /*30465*/;
  assign inv_26[8] = ~div[8] /*30464*/;
  assign inv_26[9] = ~div[9] /*30463*/;
  assign inv_26[10] = ~div[10] /*30462*/;
  assign inv_26[11] = ~div[11] /*30461*/;
  assign inv_26[12] = ~div[12] /*30460*/;
  assign inv_26[13] = ~div[13] /*30459*/;
  assign inv_26[14] = ~div[14] /*30458*/;
  assign inv_26[15] = ~div[15] /*30457*/;
  assign inv_26[16] = ~div[16] /*30456*/;
  assign inv_26[17] = ~div[17] /*30455*/;
  assign inv_26[18] = ~div[18] /*30454*/;
  assign inv_26[19] = ~div[19] /*30453*/;
  assign inv_26[20] = ~div[20] /*30452*/;
  assign inv_26[21] = ~div[21] /*30451*/;
  assign inv_26[22] = ~div[22] /*30450*/;
  assign inv_26[23] = ~div[23] /*30449*/;
  assign inv_26[24] = ~div[24] /*30448*/;
  assign inv_26[25] = ~div[25] /*30447*/;
  assign inv_26[26] = ~div[26] /*30446*/;
  assign inv_26[27] = ~div[27] /*30445*/;
  assign inv_26[28] = ~div[28] /*30444*/;
  assign inv_26[29] = ~div[29] /*30443*/;
  assign inv_26[30] = ~div[30] /*30442*/;
assign inv_26[31] = oneWire /*30441*/;
  assign _5600_ = inv_26[0] ^ r_25[6] /*30439*/;
  assign sum_26[0] = _5600_ ^ oneWire /*30438*/;
  assign _5601_ = _5600_ & oneWire /*30437*/;
  assign _5602_ = inv_26[0] & r_25[6] /*30436*/;
  assign _5603_ = _5601_ | _5602_ /*30435*/;
  assign _5604_ = inv_26[1] ^ r_25[7] /*30434*/;
  assign sum_26[1] = _5604_ ^ _5603_ /*30433*/;
  assign _5605_ = _5604_ & _5603_ /*30432*/;
  assign _5606_ = inv_26[1] & r_25[7] /*30431*/;
  assign _5607_ = _5605_ | _5606_ /*30430*/;
  assign _5608_ = inv_26[2] ^ r_25[8] /*30428*/;
  assign sum_26[2] = _5608_ ^ _5607_ /*30427*/;
  assign _5609_ = _5608_ & _5607_ /*30426*/;
  assign _5610_ = inv_26[2] & r_25[8] /*30425*/;
  assign _5611_ = _5609_ | _5610_ /*30424*/;
  assign _5612_ = inv_26[3] ^ r_25[9] /*30422*/;
  assign sum_26[3] = _5612_ ^ _5611_ /*30421*/;
  assign _5613_ = _5612_ & _5611_ /*30420*/;
  assign _5614_ = inv_26[3] & r_25[9] /*30419*/;
  assign _5615_ = _5613_ | _5614_ /*30418*/;
  assign _5616_ = inv_26[4] ^ r_25[10] /*30416*/;
  assign sum_26[4] = _5616_ ^ _5615_ /*30415*/;
  assign _5617_ = _5616_ & _5615_ /*30414*/;
  assign _5618_ = inv_26[4] & r_25[10] /*30413*/;
  assign _5619_ = _5617_ | _5618_ /*30412*/;
  assign _5620_ = inv_26[5] ^ r_25[11] /*30410*/;
  assign sum_26[5] = _5620_ ^ _5619_ /*30409*/;
  assign _5621_ = _5620_ & _5619_ /*30408*/;
  assign _5622_ = inv_26[5] & r_25[11] /*30407*/;
  assign _5623_ = _5621_ | _5622_ /*30406*/;
  assign _5624_ = inv_26[6] ^ r_25[12] /*30404*/;
  assign sum_26[6] = _5624_ ^ _5623_ /*30403*/;
  assign _5625_ = _5624_ & _5623_ /*30402*/;
  assign _5626_ = inv_26[6] & r_25[12] /*30401*/;
  assign _5627_ = _5625_ | _5626_ /*30400*/;
  assign _5628_ = inv_26[7] ^ r_25[13] /*30398*/;
  assign sum_26[7] = _5628_ ^ _5627_ /*30397*/;
  assign _5629_ = _5628_ & _5627_ /*30396*/;
  assign _5630_ = inv_26[7] & r_25[13] /*30395*/;
  assign _5631_ = _5629_ | _5630_ /*30394*/;
  assign _5632_ = inv_26[8] ^ r_25[14] /*30392*/;
  assign sum_26[8] = _5632_ ^ _5631_ /*30391*/;
  assign _5633_ = _5632_ & _5631_ /*30390*/;
  assign _5634_ = inv_26[8] & r_25[14] /*30389*/;
  assign _5635_ = _5633_ | _5634_ /*30388*/;
  assign _5636_ = inv_26[9] ^ r_25[15] /*30386*/;
  assign sum_26[9] = _5636_ ^ _5635_ /*30385*/;
  assign _5637_ = _5636_ & _5635_ /*30384*/;
  assign _5638_ = inv_26[9] & r_25[15] /*30383*/;
  assign _5639_ = _5637_ | _5638_ /*30382*/;
  assign _5640_ = inv_26[10] ^ r_25[16] /*30380*/;
  assign sum_26[10] = _5640_ ^ _5639_ /*30379*/;
  assign _5641_ = _5640_ & _5639_ /*30378*/;
  assign _5642_ = inv_26[10] & r_25[16] /*30377*/;
  assign _5643_ = _5641_ | _5642_ /*30376*/;
  assign _5644_ = inv_26[11] ^ r_25[17] /*30374*/;
  assign sum_26[11] = _5644_ ^ _5643_ /*30373*/;
  assign _5645_ = _5644_ & _5643_ /*30372*/;
  assign _5646_ = inv_26[11] & r_25[17] /*30371*/;
  assign _5647_ = _5645_ | _5646_ /*30370*/;
  assign _5648_ = inv_26[12] ^ r_25[18] /*30368*/;
  assign sum_26[12] = _5648_ ^ _5647_ /*30367*/;
  assign _5649_ = _5648_ & _5647_ /*30366*/;
  assign _5650_ = inv_26[12] & r_25[18] /*30365*/;
  assign _5651_ = _5649_ | _5650_ /*30364*/;
  assign _5652_ = inv_26[13] ^ r_25[19] /*30362*/;
  assign sum_26[13] = _5652_ ^ _5651_ /*30361*/;
  assign _5653_ = _5652_ & _5651_ /*30360*/;
  assign _5654_ = inv_26[13] & r_25[19] /*30359*/;
  assign _5655_ = _5653_ | _5654_ /*30358*/;
  assign _5656_ = inv_26[14] ^ r_25[20] /*30356*/;
  assign sum_26[14] = _5656_ ^ _5655_ /*30355*/;
  assign _5657_ = _5656_ & _5655_ /*30354*/;
  assign _5658_ = inv_26[14] & r_25[20] /*30353*/;
  assign _5659_ = _5657_ | _5658_ /*30352*/;
  assign _5660_ = inv_26[15] ^ r_25[21] /*30350*/;
  assign sum_26[15] = _5660_ ^ _5659_ /*30349*/;
  assign _5661_ = _5660_ & _5659_ /*30348*/;
  assign _5662_ = inv_26[15] & r_25[21] /*30347*/;
  assign _5663_ = _5661_ | _5662_ /*30346*/;
  assign _5664_ = inv_26[16] ^ r_25[22] /*30344*/;
  assign sum_26[16] = _5664_ ^ _5663_ /*30343*/;
  assign _5665_ = _5664_ & _5663_ /*30342*/;
  assign _5666_ = inv_26[16] & r_25[22] /*30341*/;
  assign _5667_ = _5665_ | _5666_ /*30340*/;
  assign _5668_ = inv_26[17] ^ r_25[23] /*30338*/;
  assign sum_26[17] = _5668_ ^ _5667_ /*30337*/;
  assign _5669_ = _5668_ & _5667_ /*30336*/;
  assign _5670_ = inv_26[17] & r_25[23] /*30335*/;
  assign _5671_ = _5669_ | _5670_ /*30334*/;
  assign _5672_ = inv_26[18] ^ r_25[24] /*30332*/;
  assign sum_26[18] = _5672_ ^ _5671_ /*30331*/;
  assign _5673_ = _5672_ & _5671_ /*30330*/;
  assign _5674_ = inv_26[18] & r_25[24] /*30329*/;
  assign _5675_ = _5673_ | _5674_ /*30328*/;
  assign _5676_ = inv_26[19] ^ r_25[25] /*30326*/;
  assign sum_26[19] = _5676_ ^ _5675_ /*30325*/;
  assign _5677_ = _5676_ & _5675_ /*30324*/;
  assign _5678_ = inv_26[19] & r_25[25] /*30323*/;
  assign _5679_ = _5677_ | _5678_ /*30322*/;
  assign _5680_ = inv_26[20] ^ r_25[26] /*30320*/;
  assign sum_26[20] = _5680_ ^ _5679_ /*30319*/;
  assign _5681_ = _5680_ & _5679_ /*30318*/;
  assign _5682_ = inv_26[20] & r_25[26] /*30317*/;
  assign _5683_ = _5681_ | _5682_ /*30316*/;
  assign _5684_ = inv_26[21] ^ r_25[27] /*30314*/;
  assign sum_26[21] = _5684_ ^ _5683_ /*30313*/;
  assign _5685_ = _5684_ & _5683_ /*30312*/;
  assign _5686_ = inv_26[21] & r_25[27] /*30311*/;
  assign _5687_ = _5685_ | _5686_ /*30310*/;
  assign _5688_ = inv_26[22] ^ r_25[28] /*30308*/;
  assign sum_26[22] = _5688_ ^ _5687_ /*30307*/;
  assign _5689_ = _5688_ & _5687_ /*30306*/;
  assign _5690_ = inv_26[22] & r_25[28] /*30305*/;
  assign _5691_ = _5689_ | _5690_ /*30304*/;
  assign _5692_ = inv_26[23] ^ r_25[29] /*30302*/;
  assign sum_26[23] = _5692_ ^ _5691_ /*30301*/;
  assign _5693_ = _5692_ & _5691_ /*30300*/;
  assign _5694_ = inv_26[23] & r_25[29] /*30299*/;
  assign _5695_ = _5693_ | _5694_ /*30298*/;
  assign _5696_ = inv_26[24] ^ r_25[30] /*30296*/;
  assign sum_26[24] = _5696_ ^ _5695_ /*30295*/;
  assign _5697_ = _5696_ & _5695_ /*30294*/;
  assign _5698_ = inv_26[24] & r_25[30] /*30293*/;
  assign _5699_ = _5697_ | _5698_ /*30292*/;
  assign _5700_ = inv_26[25] ^ r_25[31] /*30290*/;
  assign sum_26[25] = _5700_ ^ _5699_ /*30289*/;
  assign _5701_ = _5700_ & _5699_ /*30288*/;
  assign _5702_ = inv_26[25] & r_25[31] /*30287*/;
  assign _5703_ = _5701_ | _5702_ /*30286*/;
  assign _5704_ = inv_26[26] ^ r_25[32] /*30284*/;
  assign sum_26[26] = _5704_ ^ _5703_ /*30283*/;
  assign _5705_ = _5704_ & _5703_ /*30282*/;
  assign _5706_ = inv_26[26] & r_25[32] /*30281*/;
  assign _5707_ = _5705_ | _5706_ /*30280*/;
  assign _5708_ = inv_26[27] ^ r_25[33] /*30278*/;
  assign sum_26[27] = _5708_ ^ _5707_ /*30277*/;
  assign _5709_ = _5708_ & _5707_ /*30276*/;
  assign _5710_ = inv_26[27] & r_25[33] /*30275*/;
  assign _5711_ = _5709_ | _5710_ /*30274*/;
  assign _5712_ = inv_26[28] ^ r_25[34] /*30272*/;
  assign sum_26[28] = _5712_ ^ _5711_ /*30271*/;
  assign _5713_ = _5712_ & _5711_ /*30270*/;
  assign _5714_ = inv_26[28] & r_25[34] /*30269*/;
  assign _5715_ = _5713_ | _5714_ /*30268*/;
  assign _5716_ = inv_26[29] ^ r_25[35] /*30266*/;
  assign sum_26[29] = _5716_ ^ _5715_ /*30265*/;
  assign _5717_ = _5716_ & _5715_ /*30264*/;
  assign _5718_ = inv_26[29] & r_25[35] /*30263*/;
  assign _5719_ = _5717_ | _5718_ /*30262*/;
  assign _5720_ = inv_26[30] ^ r_25[36] /*30260*/;
  assign sum_26[30] = _5720_ ^ _5719_ /*30259*/;
  assign _5721_ = _5720_ & _5719_ /*30258*/;
  assign _5722_ = inv_26[30] & r_25[36] /*30257*/;
  assign _5723_ = _5721_ | _5722_ /*30256*/;
  assign _5724_ = inv_26[31] ^ r_25[37] /*30254*/;
  assign sum_26[31] = _5724_ ^ _5723_ /*30253*/;
  assign _5725_ = _5724_ & _5723_ /*30252*/;
  assign _5726_ = inv_26[31] & r_25[37] /*30251*/;
  assign _5727_ = _5725_ | _5726_ /*30250*/;
  assign q[6] = ~sum_26[31] /*30277*/;
  assign m_26[0] = r_25[6] /*30276*/;
  assign m_26[1] = r_25[7] /*30275*/;
  assign m_26[2] = r_25[8] /*30274*/;
  assign m_26[3] = r_25[9] /*30273*/;
  assign m_26[4] = r_25[10] /*30272*/;
  assign m_26[5] = r_25[11] /*30271*/;
  assign m_26[6] = r_25[12] /*30270*/;
  assign m_26[7] = r_25[13] /*30269*/;
  assign m_26[8] = r_25[14] /*30268*/;
  assign m_26[9] = r_25[15] /*30267*/;
  assign m_26[10] = r_25[16] /*30266*/;
  assign m_26[11] = r_25[17] /*30265*/;
  assign m_26[12] = r_25[18] /*30264*/;
  assign m_26[13] = r_25[19] /*30263*/;
  assign m_26[14] = r_25[20] /*30262*/;
  assign m_26[15] = r_25[21] /*30261*/;
  assign m_26[16] = r_25[22] /*30260*/;
  assign m_26[17] = r_25[23] /*30259*/;
  assign m_26[18] = r_25[24] /*30258*/;
  assign m_26[19] = r_25[25] /*30257*/;
  assign m_26[20] = r_25[26] /*30256*/;
  assign m_26[21] = r_25[27] /*30255*/;
  assign m_26[22] = r_25[28] /*30254*/;
  assign m_26[23] = r_25[29] /*30253*/;
  assign m_26[24] = r_25[30] /*30252*/;
  assign m_26[25] = r_25[31] /*30251*/;
  assign m_26[26] = r_25[32] /*30250*/;
  assign m_26[27] = r_25[33] /*30249*/;
  assign m_26[28] = r_25[34] /*30248*/;
  assign m_26[29] = r_25[35] /*30247*/;
  assign m_26[30] = r_25[36] /*30246*/;
  assign m_26[31] = r_25[37] /*30245*/;
  assign _5728_ = ~q[6] /*30243*/;
  assign _5729_ = sum_26[0] & q[6] /*30242*/;
  assign _5730_ = m_26[0] & _5728_ /*30241*/;
  assign r_26[6] = _5730_ | _5729_ /*30240*/;
  assign _5731_ = ~q[6] /*30239*/;
  assign _5732_ = sum_26[1] & q[6] /*30238*/;
  assign _5733_ = m_26[1] & _5731_ /*30237*/;
  assign r_26[7] = _5733_ | _5732_ /*30236*/;
  assign _5734_ = ~q[6] /*30235*/;
  assign _5735_ = sum_26[2] & q[6] /*30234*/;
  assign _5736_ = m_26[2] & _5734_ /*30233*/;
  assign r_26[8] = _5736_ | _5735_ /*30232*/;
  assign _5737_ = ~q[6] /*30231*/;
  assign _5738_ = sum_26[3] & q[6] /*30230*/;
  assign _5739_ = m_26[3] & _5737_ /*30229*/;
  assign r_26[9] = _5739_ | _5738_ /*30228*/;
  assign _5740_ = ~q[6] /*30227*/;
  assign _5741_ = sum_26[4] & q[6] /*30226*/;
  assign _5742_ = m_26[4] & _5740_ /*30225*/;
  assign r_26[10] = _5742_ | _5741_ /*30224*/;
  assign _5743_ = ~q[6] /*30223*/;
  assign _5744_ = sum_26[5] & q[6] /*30222*/;
  assign _5745_ = m_26[5] & _5743_ /*30221*/;
  assign r_26[11] = _5745_ | _5744_ /*30220*/;
  assign _5746_ = ~q[6] /*30219*/;
  assign _5747_ = sum_26[6] & q[6] /*30218*/;
  assign _5748_ = m_26[6] & _5746_ /*30217*/;
  assign r_26[12] = _5748_ | _5747_ /*30216*/;
  assign _5749_ = ~q[6] /*30215*/;
  assign _5750_ = sum_26[7] & q[6] /*30214*/;
  assign _5751_ = m_26[7] & _5749_ /*30213*/;
  assign r_26[13] = _5751_ | _5750_ /*30212*/;
  assign _5752_ = ~q[6] /*30211*/;
  assign _5753_ = sum_26[8] & q[6] /*30210*/;
  assign _5754_ = m_26[8] & _5752_ /*30209*/;
  assign r_26[14] = _5754_ | _5753_ /*30208*/;
  assign _5755_ = ~q[6] /*30207*/;
  assign _5756_ = sum_26[9] & q[6] /*30206*/;
  assign _5757_ = m_26[9] & _5755_ /*30205*/;
  assign r_26[15] = _5757_ | _5756_ /*30204*/;
  assign _5758_ = ~q[6] /*30203*/;
  assign _5759_ = sum_26[10] & q[6] /*30202*/;
  assign _5760_ = m_26[10] & _5758_ /*30201*/;
  assign r_26[16] = _5760_ | _5759_ /*30200*/;
  assign _5761_ = ~q[6] /*30199*/;
  assign _5762_ = sum_26[11] & q[6] /*30198*/;
  assign _5763_ = m_26[11] & _5761_ /*30197*/;
  assign r_26[17] = _5763_ | _5762_ /*30196*/;
  assign _5764_ = ~q[6] /*30195*/;
  assign _5765_ = sum_26[12] & q[6] /*30194*/;
  assign _5766_ = m_26[12] & _5764_ /*30193*/;
  assign r_26[18] = _5766_ | _5765_ /*30192*/;
  assign _5767_ = ~q[6] /*30191*/;
  assign _5768_ = sum_26[13] & q[6] /*30190*/;
  assign _5769_ = m_26[13] & _5767_ /*30189*/;
  assign r_26[19] = _5769_ | _5768_ /*30188*/;
  assign _5770_ = ~q[6] /*30187*/;
  assign _5771_ = sum_26[14] & q[6] /*30186*/;
  assign _5772_ = m_26[14] & _5770_ /*30185*/;
  assign r_26[20] = _5772_ | _5771_ /*30184*/;
  assign _5773_ = ~q[6] /*30183*/;
  assign _5774_ = sum_26[15] & q[6] /*30182*/;
  assign _5775_ = m_26[15] & _5773_ /*30181*/;
  assign r_26[21] = _5775_ | _5774_ /*30180*/;
  assign _5776_ = ~q[6] /*30179*/;
  assign _5777_ = sum_26[16] & q[6] /*30178*/;
  assign _5778_ = m_26[16] & _5776_ /*30177*/;
  assign r_26[22] = _5778_ | _5777_ /*30176*/;
  assign _5779_ = ~q[6] /*30175*/;
  assign _5780_ = sum_26[17] & q[6] /*30174*/;
  assign _5781_ = m_26[17] & _5779_ /*30173*/;
  assign r_26[23] = _5781_ | _5780_ /*30172*/;
  assign _5782_ = ~q[6] /*30171*/;
  assign _5783_ = sum_26[18] & q[6] /*30170*/;
  assign _5784_ = m_26[18] & _5782_ /*30169*/;
  assign r_26[24] = _5784_ | _5783_ /*30168*/;
  assign _5785_ = ~q[6] /*30167*/;
  assign _5786_ = sum_26[19] & q[6] /*30166*/;
  assign _5787_ = m_26[19] & _5785_ /*30165*/;
  assign r_26[25] = _5787_ | _5786_ /*30164*/;
  assign _5788_ = ~q[6] /*30163*/;
  assign _5789_ = sum_26[20] & q[6] /*30162*/;
  assign _5790_ = m_26[20] & _5788_ /*30161*/;
  assign r_26[26] = _5790_ | _5789_ /*30160*/;
  assign _5791_ = ~q[6] /*30159*/;
  assign _5792_ = sum_26[21] & q[6] /*30158*/;
  assign _5793_ = m_26[21] & _5791_ /*30157*/;
  assign r_26[27] = _5793_ | _5792_ /*30156*/;
  assign _5794_ = ~q[6] /*30155*/;
  assign _5795_ = sum_26[22] & q[6] /*30154*/;
  assign _5796_ = m_26[22] & _5794_ /*30153*/;
  assign r_26[28] = _5796_ | _5795_ /*30152*/;
  assign _5797_ = ~q[6] /*30151*/;
  assign _5798_ = sum_26[23] & q[6] /*30150*/;
  assign _5799_ = m_26[23] & _5797_ /*30149*/;
  assign r_26[29] = _5799_ | _5798_ /*30148*/;
  assign _5800_ = ~q[6] /*30147*/;
  assign _5801_ = sum_26[24] & q[6] /*30146*/;
  assign _5802_ = m_26[24] & _5800_ /*30145*/;
  assign r_26[30] = _5802_ | _5801_ /*30144*/;
  assign _5803_ = ~q[6] /*30143*/;
  assign _5804_ = sum_26[25] & q[6] /*30142*/;
  assign _5805_ = m_26[25] & _5803_ /*30141*/;
  assign r_26[31] = _5805_ | _5804_ /*30140*/;
  assign _5806_ = ~q[6] /*30139*/;
  assign _5807_ = sum_26[26] & q[6] /*30138*/;
  assign _5808_ = m_26[26] & _5806_ /*30137*/;
  assign r_26[32] = _5808_ | _5807_ /*30136*/;
  assign _5809_ = ~q[6] /*30135*/;
  assign _5810_ = sum_26[27] & q[6] /*30134*/;
  assign _5811_ = m_26[27] & _5809_ /*30133*/;
  assign r_26[33] = _5811_ | _5810_ /*30132*/;
  assign _5812_ = ~q[6] /*30131*/;
  assign _5813_ = sum_26[28] & q[6] /*30130*/;
  assign _5814_ = m_26[28] & _5812_ /*30129*/;
  assign r_26[34] = _5814_ | _5813_ /*30128*/;
  assign _5815_ = ~q[6] /*30127*/;
  assign _5816_ = sum_26[29] & q[6] /*30126*/;
  assign _5817_ = m_26[29] & _5815_ /*30125*/;
  assign r_26[35] = _5817_ | _5816_ /*30124*/;
  assign _5818_ = ~q[6] /*30123*/;
  assign _5819_ = sum_26[30] & q[6] /*30122*/;
  assign _5820_ = m_26[30] & _5818_ /*30121*/;
  assign r_26[36] = _5820_ | _5819_ /*30120*/;
  assign _5821_ = ~q[6] /*30119*/;
  assign _5822_ = sum_26[31] & q[6] /*30118*/;
  assign _5823_ = m_26[31] & _5821_ /*30117*/;
  assign r_26[37] = _5823_ | _5822_ /*30116*/;
assign r_26[0]= r_25[0] /*30115*/;
assign r_26[1]= r_25[1] /*30114*/;
assign r_26[2]= r_25[2] /*30113*/;
assign r_26[3]= r_25[3] /*30112*/;
assign r_26[4]= r_25[4] /*30111*/;
assign r_26[5]= r_25[5] /*30110*/;
  assign inv_27[0] = ~div[0] /*30024*/;
  assign inv_27[1] = ~div[1] /*30023*/;
  assign inv_27[2] = ~div[2] /*30022*/;
  assign inv_27[3] = ~div[3] /*30021*/;
  assign inv_27[4] = ~div[4] /*30020*/;
  assign inv_27[5] = ~div[5] /*30019*/;
  assign inv_27[6] = ~div[6] /*30018*/;
  assign inv_27[7] = ~div[7] /*30017*/;
  assign inv_27[8] = ~div[8] /*30016*/;
  assign inv_27[9] = ~div[9] /*30015*/;
  assign inv_27[10] = ~div[10] /*30014*/;
  assign inv_27[11] = ~div[11] /*30013*/;
  assign inv_27[12] = ~div[12] /*30012*/;
  assign inv_27[13] = ~div[13] /*30011*/;
  assign inv_27[14] = ~div[14] /*30010*/;
  assign inv_27[15] = ~div[15] /*30009*/;
  assign inv_27[16] = ~div[16] /*30008*/;
  assign inv_27[17] = ~div[17] /*30007*/;
  assign inv_27[18] = ~div[18] /*30006*/;
  assign inv_27[19] = ~div[19] /*30005*/;
  assign inv_27[20] = ~div[20] /*30004*/;
  assign inv_27[21] = ~div[21] /*30003*/;
  assign inv_27[22] = ~div[22] /*30002*/;
  assign inv_27[23] = ~div[23] /*30001*/;
  assign inv_27[24] = ~div[24] /*30000*/;
  assign inv_27[25] = ~div[25] /*29999*/;
  assign inv_27[26] = ~div[26] /*29998*/;
  assign inv_27[27] = ~div[27] /*29997*/;
  assign inv_27[28] = ~div[28] /*29996*/;
  assign inv_27[29] = ~div[29] /*29995*/;
  assign inv_27[30] = ~div[30] /*29994*/;
assign inv_27[31] = oneWire /*29993*/;
  assign _5824_ = inv_27[0] ^ r_26[5] /*29991*/;
  assign sum_27[0] = _5824_ ^ oneWire /*29990*/;
  assign _5825_ = _5824_ & oneWire /*29989*/;
  assign _5826_ = inv_27[0] & r_26[5] /*29988*/;
  assign _5827_ = _5825_ | _5826_ /*29987*/;
  assign _5828_ = inv_27[1] ^ r_26[6] /*29986*/;
  assign sum_27[1] = _5828_ ^ _5827_ /*29985*/;
  assign _5829_ = _5828_ & _5827_ /*29984*/;
  assign _5830_ = inv_27[1] & r_26[6] /*29983*/;
  assign _5831_ = _5829_ | _5830_ /*29982*/;
  assign _5832_ = inv_27[2] ^ r_26[7] /*29980*/;
  assign sum_27[2] = _5832_ ^ _5831_ /*29979*/;
  assign _5833_ = _5832_ & _5831_ /*29978*/;
  assign _5834_ = inv_27[2] & r_26[7] /*29977*/;
  assign _5835_ = _5833_ | _5834_ /*29976*/;
  assign _5836_ = inv_27[3] ^ r_26[8] /*29974*/;
  assign sum_27[3] = _5836_ ^ _5835_ /*29973*/;
  assign _5837_ = _5836_ & _5835_ /*29972*/;
  assign _5838_ = inv_27[3] & r_26[8] /*29971*/;
  assign _5839_ = _5837_ | _5838_ /*29970*/;
  assign _5840_ = inv_27[4] ^ r_26[9] /*29968*/;
  assign sum_27[4] = _5840_ ^ _5839_ /*29967*/;
  assign _5841_ = _5840_ & _5839_ /*29966*/;
  assign _5842_ = inv_27[4] & r_26[9] /*29965*/;
  assign _5843_ = _5841_ | _5842_ /*29964*/;
  assign _5844_ = inv_27[5] ^ r_26[10] /*29962*/;
  assign sum_27[5] = _5844_ ^ _5843_ /*29961*/;
  assign _5845_ = _5844_ & _5843_ /*29960*/;
  assign _5846_ = inv_27[5] & r_26[10] /*29959*/;
  assign _5847_ = _5845_ | _5846_ /*29958*/;
  assign _5848_ = inv_27[6] ^ r_26[11] /*29956*/;
  assign sum_27[6] = _5848_ ^ _5847_ /*29955*/;
  assign _5849_ = _5848_ & _5847_ /*29954*/;
  assign _5850_ = inv_27[6] & r_26[11] /*29953*/;
  assign _5851_ = _5849_ | _5850_ /*29952*/;
  assign _5852_ = inv_27[7] ^ r_26[12] /*29950*/;
  assign sum_27[7] = _5852_ ^ _5851_ /*29949*/;
  assign _5853_ = _5852_ & _5851_ /*29948*/;
  assign _5854_ = inv_27[7] & r_26[12] /*29947*/;
  assign _5855_ = _5853_ | _5854_ /*29946*/;
  assign _5856_ = inv_27[8] ^ r_26[13] /*29944*/;
  assign sum_27[8] = _5856_ ^ _5855_ /*29943*/;
  assign _5857_ = _5856_ & _5855_ /*29942*/;
  assign _5858_ = inv_27[8] & r_26[13] /*29941*/;
  assign _5859_ = _5857_ | _5858_ /*29940*/;
  assign _5860_ = inv_27[9] ^ r_26[14] /*29938*/;
  assign sum_27[9] = _5860_ ^ _5859_ /*29937*/;
  assign _5861_ = _5860_ & _5859_ /*29936*/;
  assign _5862_ = inv_27[9] & r_26[14] /*29935*/;
  assign _5863_ = _5861_ | _5862_ /*29934*/;
  assign _5864_ = inv_27[10] ^ r_26[15] /*29932*/;
  assign sum_27[10] = _5864_ ^ _5863_ /*29931*/;
  assign _5865_ = _5864_ & _5863_ /*29930*/;
  assign _5866_ = inv_27[10] & r_26[15] /*29929*/;
  assign _5867_ = _5865_ | _5866_ /*29928*/;
  assign _5868_ = inv_27[11] ^ r_26[16] /*29926*/;
  assign sum_27[11] = _5868_ ^ _5867_ /*29925*/;
  assign _5869_ = _5868_ & _5867_ /*29924*/;
  assign _5870_ = inv_27[11] & r_26[16] /*29923*/;
  assign _5871_ = _5869_ | _5870_ /*29922*/;
  assign _5872_ = inv_27[12] ^ r_26[17] /*29920*/;
  assign sum_27[12] = _5872_ ^ _5871_ /*29919*/;
  assign _5873_ = _5872_ & _5871_ /*29918*/;
  assign _5874_ = inv_27[12] & r_26[17] /*29917*/;
  assign _5875_ = _5873_ | _5874_ /*29916*/;
  assign _5876_ = inv_27[13] ^ r_26[18] /*29914*/;
  assign sum_27[13] = _5876_ ^ _5875_ /*29913*/;
  assign _5877_ = _5876_ & _5875_ /*29912*/;
  assign _5878_ = inv_27[13] & r_26[18] /*29911*/;
  assign _5879_ = _5877_ | _5878_ /*29910*/;
  assign _5880_ = inv_27[14] ^ r_26[19] /*29908*/;
  assign sum_27[14] = _5880_ ^ _5879_ /*29907*/;
  assign _5881_ = _5880_ & _5879_ /*29906*/;
  assign _5882_ = inv_27[14] & r_26[19] /*29905*/;
  assign _5883_ = _5881_ | _5882_ /*29904*/;
  assign _5884_ = inv_27[15] ^ r_26[20] /*29902*/;
  assign sum_27[15] = _5884_ ^ _5883_ /*29901*/;
  assign _5885_ = _5884_ & _5883_ /*29900*/;
  assign _5886_ = inv_27[15] & r_26[20] /*29899*/;
  assign _5887_ = _5885_ | _5886_ /*29898*/;
  assign _5888_ = inv_27[16] ^ r_26[21] /*29896*/;
  assign sum_27[16] = _5888_ ^ _5887_ /*29895*/;
  assign _5889_ = _5888_ & _5887_ /*29894*/;
  assign _5890_ = inv_27[16] & r_26[21] /*29893*/;
  assign _5891_ = _5889_ | _5890_ /*29892*/;
  assign _5892_ = inv_27[17] ^ r_26[22] /*29890*/;
  assign sum_27[17] = _5892_ ^ _5891_ /*29889*/;
  assign _5893_ = _5892_ & _5891_ /*29888*/;
  assign _5894_ = inv_27[17] & r_26[22] /*29887*/;
  assign _5895_ = _5893_ | _5894_ /*29886*/;
  assign _5896_ = inv_27[18] ^ r_26[23] /*29884*/;
  assign sum_27[18] = _5896_ ^ _5895_ /*29883*/;
  assign _5897_ = _5896_ & _5895_ /*29882*/;
  assign _5898_ = inv_27[18] & r_26[23] /*29881*/;
  assign _5899_ = _5897_ | _5898_ /*29880*/;
  assign _5900_ = inv_27[19] ^ r_26[24] /*29878*/;
  assign sum_27[19] = _5900_ ^ _5899_ /*29877*/;
  assign _5901_ = _5900_ & _5899_ /*29876*/;
  assign _5902_ = inv_27[19] & r_26[24] /*29875*/;
  assign _5903_ = _5901_ | _5902_ /*29874*/;
  assign _5904_ = inv_27[20] ^ r_26[25] /*29872*/;
  assign sum_27[20] = _5904_ ^ _5903_ /*29871*/;
  assign _5905_ = _5904_ & _5903_ /*29870*/;
  assign _5906_ = inv_27[20] & r_26[25] /*29869*/;
  assign _5907_ = _5905_ | _5906_ /*29868*/;
  assign _5908_ = inv_27[21] ^ r_26[26] /*29866*/;
  assign sum_27[21] = _5908_ ^ _5907_ /*29865*/;
  assign _5909_ = _5908_ & _5907_ /*29864*/;
  assign _5910_ = inv_27[21] & r_26[26] /*29863*/;
  assign _5911_ = _5909_ | _5910_ /*29862*/;
  assign _5912_ = inv_27[22] ^ r_26[27] /*29860*/;
  assign sum_27[22] = _5912_ ^ _5911_ /*29859*/;
  assign _5913_ = _5912_ & _5911_ /*29858*/;
  assign _5914_ = inv_27[22] & r_26[27] /*29857*/;
  assign _5915_ = _5913_ | _5914_ /*29856*/;
  assign _5916_ = inv_27[23] ^ r_26[28] /*29854*/;
  assign sum_27[23] = _5916_ ^ _5915_ /*29853*/;
  assign _5917_ = _5916_ & _5915_ /*29852*/;
  assign _5918_ = inv_27[23] & r_26[28] /*29851*/;
  assign _5919_ = _5917_ | _5918_ /*29850*/;
  assign _5920_ = inv_27[24] ^ r_26[29] /*29848*/;
  assign sum_27[24] = _5920_ ^ _5919_ /*29847*/;
  assign _5921_ = _5920_ & _5919_ /*29846*/;
  assign _5922_ = inv_27[24] & r_26[29] /*29845*/;
  assign _5923_ = _5921_ | _5922_ /*29844*/;
  assign _5924_ = inv_27[25] ^ r_26[30] /*29842*/;
  assign sum_27[25] = _5924_ ^ _5923_ /*29841*/;
  assign _5925_ = _5924_ & _5923_ /*29840*/;
  assign _5926_ = inv_27[25] & r_26[30] /*29839*/;
  assign _5927_ = _5925_ | _5926_ /*29838*/;
  assign _5928_ = inv_27[26] ^ r_26[31] /*29836*/;
  assign sum_27[26] = _5928_ ^ _5927_ /*29835*/;
  assign _5929_ = _5928_ & _5927_ /*29834*/;
  assign _5930_ = inv_27[26] & r_26[31] /*29833*/;
  assign _5931_ = _5929_ | _5930_ /*29832*/;
  assign _5932_ = inv_27[27] ^ r_26[32] /*29830*/;
  assign sum_27[27] = _5932_ ^ _5931_ /*29829*/;
  assign _5933_ = _5932_ & _5931_ /*29828*/;
  assign _5934_ = inv_27[27] & r_26[32] /*29827*/;
  assign _5935_ = _5933_ | _5934_ /*29826*/;
  assign _5936_ = inv_27[28] ^ r_26[33] /*29824*/;
  assign sum_27[28] = _5936_ ^ _5935_ /*29823*/;
  assign _5937_ = _5936_ & _5935_ /*29822*/;
  assign _5938_ = inv_27[28] & r_26[33] /*29821*/;
  assign _5939_ = _5937_ | _5938_ /*29820*/;
  assign _5940_ = inv_27[29] ^ r_26[34] /*29818*/;
  assign sum_27[29] = _5940_ ^ _5939_ /*29817*/;
  assign _5941_ = _5940_ & _5939_ /*29816*/;
  assign _5942_ = inv_27[29] & r_26[34] /*29815*/;
  assign _5943_ = _5941_ | _5942_ /*29814*/;
  assign _5944_ = inv_27[30] ^ r_26[35] /*29812*/;
  assign sum_27[30] = _5944_ ^ _5943_ /*29811*/;
  assign _5945_ = _5944_ & _5943_ /*29810*/;
  assign _5946_ = inv_27[30] & r_26[35] /*29809*/;
  assign _5947_ = _5945_ | _5946_ /*29808*/;
  assign _5948_ = inv_27[31] ^ r_26[36] /*29806*/;
  assign sum_27[31] = _5948_ ^ _5947_ /*29805*/;
  assign _5949_ = _5948_ & _5947_ /*29804*/;
  assign _5950_ = inv_27[31] & r_26[36] /*29803*/;
  assign _5951_ = _5949_ | _5950_ /*29802*/;
  assign q[5] = ~sum_27[31] /*29829*/;
  assign m_27[0] = r_26[5] /*29828*/;
  assign m_27[1] = r_26[6] /*29827*/;
  assign m_27[2] = r_26[7] /*29826*/;
  assign m_27[3] = r_26[8] /*29825*/;
  assign m_27[4] = r_26[9] /*29824*/;
  assign m_27[5] = r_26[10] /*29823*/;
  assign m_27[6] = r_26[11] /*29822*/;
  assign m_27[7] = r_26[12] /*29821*/;
  assign m_27[8] = r_26[13] /*29820*/;
  assign m_27[9] = r_26[14] /*29819*/;
  assign m_27[10] = r_26[15] /*29818*/;
  assign m_27[11] = r_26[16] /*29817*/;
  assign m_27[12] = r_26[17] /*29816*/;
  assign m_27[13] = r_26[18] /*29815*/;
  assign m_27[14] = r_26[19] /*29814*/;
  assign m_27[15] = r_26[20] /*29813*/;
  assign m_27[16] = r_26[21] /*29812*/;
  assign m_27[17] = r_26[22] /*29811*/;
  assign m_27[18] = r_26[23] /*29810*/;
  assign m_27[19] = r_26[24] /*29809*/;
  assign m_27[20] = r_26[25] /*29808*/;
  assign m_27[21] = r_26[26] /*29807*/;
  assign m_27[22] = r_26[27] /*29806*/;
  assign m_27[23] = r_26[28] /*29805*/;
  assign m_27[24] = r_26[29] /*29804*/;
  assign m_27[25] = r_26[30] /*29803*/;
  assign m_27[26] = r_26[31] /*29802*/;
  assign m_27[27] = r_26[32] /*29801*/;
  assign m_27[28] = r_26[33] /*29800*/;
  assign m_27[29] = r_26[34] /*29799*/;
  assign m_27[30] = r_26[35] /*29798*/;
  assign m_27[31] = r_26[36] /*29797*/;
  assign _5952_ = ~q[5] /*29795*/;
  assign _5953_ = sum_27[0] & q[5] /*29794*/;
  assign _5954_ = m_27[0] & _5952_ /*29793*/;
  assign r_27[5] = _5954_ | _5953_ /*29792*/;
  assign _5955_ = ~q[5] /*29791*/;
  assign _5956_ = sum_27[1] & q[5] /*29790*/;
  assign _5957_ = m_27[1] & _5955_ /*29789*/;
  assign r_27[6] = _5957_ | _5956_ /*29788*/;
  assign _5958_ = ~q[5] /*29787*/;
  assign _5959_ = sum_27[2] & q[5] /*29786*/;
  assign _5960_ = m_27[2] & _5958_ /*29785*/;
  assign r_27[7] = _5960_ | _5959_ /*29784*/;
  assign _5961_ = ~q[5] /*29783*/;
  assign _5962_ = sum_27[3] & q[5] /*29782*/;
  assign _5963_ = m_27[3] & _5961_ /*29781*/;
  assign r_27[8] = _5963_ | _5962_ /*29780*/;
  assign _5964_ = ~q[5] /*29779*/;
  assign _5965_ = sum_27[4] & q[5] /*29778*/;
  assign _5966_ = m_27[4] & _5964_ /*29777*/;
  assign r_27[9] = _5966_ | _5965_ /*29776*/;
  assign _5967_ = ~q[5] /*29775*/;
  assign _5968_ = sum_27[5] & q[5] /*29774*/;
  assign _5969_ = m_27[5] & _5967_ /*29773*/;
  assign r_27[10] = _5969_ | _5968_ /*29772*/;
  assign _5970_ = ~q[5] /*29771*/;
  assign _5971_ = sum_27[6] & q[5] /*29770*/;
  assign _5972_ = m_27[6] & _5970_ /*29769*/;
  assign r_27[11] = _5972_ | _5971_ /*29768*/;
  assign _5973_ = ~q[5] /*29767*/;
  assign _5974_ = sum_27[7] & q[5] /*29766*/;
  assign _5975_ = m_27[7] & _5973_ /*29765*/;
  assign r_27[12] = _5975_ | _5974_ /*29764*/;
  assign _5976_ = ~q[5] /*29763*/;
  assign _5977_ = sum_27[8] & q[5] /*29762*/;
  assign _5978_ = m_27[8] & _5976_ /*29761*/;
  assign r_27[13] = _5978_ | _5977_ /*29760*/;
  assign _5979_ = ~q[5] /*29759*/;
  assign _5980_ = sum_27[9] & q[5] /*29758*/;
  assign _5981_ = m_27[9] & _5979_ /*29757*/;
  assign r_27[14] = _5981_ | _5980_ /*29756*/;
  assign _5982_ = ~q[5] /*29755*/;
  assign _5983_ = sum_27[10] & q[5] /*29754*/;
  assign _5984_ = m_27[10] & _5982_ /*29753*/;
  assign r_27[15] = _5984_ | _5983_ /*29752*/;
  assign _5985_ = ~q[5] /*29751*/;
  assign _5986_ = sum_27[11] & q[5] /*29750*/;
  assign _5987_ = m_27[11] & _5985_ /*29749*/;
  assign r_27[16] = _5987_ | _5986_ /*29748*/;
  assign _5988_ = ~q[5] /*29747*/;
  assign _5989_ = sum_27[12] & q[5] /*29746*/;
  assign _5990_ = m_27[12] & _5988_ /*29745*/;
  assign r_27[17] = _5990_ | _5989_ /*29744*/;
  assign _5991_ = ~q[5] /*29743*/;
  assign _5992_ = sum_27[13] & q[5] /*29742*/;
  assign _5993_ = m_27[13] & _5991_ /*29741*/;
  assign r_27[18] = _5993_ | _5992_ /*29740*/;
  assign _5994_ = ~q[5] /*29739*/;
  assign _5995_ = sum_27[14] & q[5] /*29738*/;
  assign _5996_ = m_27[14] & _5994_ /*29737*/;
  assign r_27[19] = _5996_ | _5995_ /*29736*/;
  assign _5997_ = ~q[5] /*29735*/;
  assign _5998_ = sum_27[15] & q[5] /*29734*/;
  assign _5999_ = m_27[15] & _5997_ /*29733*/;
  assign r_27[20] = _5999_ | _5998_ /*29732*/;
  assign _6000_ = ~q[5] /*29731*/;
  assign _6001_ = sum_27[16] & q[5] /*29730*/;
  assign _6002_ = m_27[16] & _6000_ /*29729*/;
  assign r_27[21] = _6002_ | _6001_ /*29728*/;
  assign _6003_ = ~q[5] /*29727*/;
  assign _6004_ = sum_27[17] & q[5] /*29726*/;
  assign _6005_ = m_27[17] & _6003_ /*29725*/;
  assign r_27[22] = _6005_ | _6004_ /*29724*/;
  assign _6006_ = ~q[5] /*29723*/;
  assign _6007_ = sum_27[18] & q[5] /*29722*/;
  assign _6008_ = m_27[18] & _6006_ /*29721*/;
  assign r_27[23] = _6008_ | _6007_ /*29720*/;
  assign _6009_ = ~q[5] /*29719*/;
  assign _6010_ = sum_27[19] & q[5] /*29718*/;
  assign _6011_ = m_27[19] & _6009_ /*29717*/;
  assign r_27[24] = _6011_ | _6010_ /*29716*/;
  assign _6012_ = ~q[5] /*29715*/;
  assign _6013_ = sum_27[20] & q[5] /*29714*/;
  assign _6014_ = m_27[20] & _6012_ /*29713*/;
  assign r_27[25] = _6014_ | _6013_ /*29712*/;
  assign _6015_ = ~q[5] /*29711*/;
  assign _6016_ = sum_27[21] & q[5] /*29710*/;
  assign _6017_ = m_27[21] & _6015_ /*29709*/;
  assign r_27[26] = _6017_ | _6016_ /*29708*/;
  assign _6018_ = ~q[5] /*29707*/;
  assign _6019_ = sum_27[22] & q[5] /*29706*/;
  assign _6020_ = m_27[22] & _6018_ /*29705*/;
  assign r_27[27] = _6020_ | _6019_ /*29704*/;
  assign _6021_ = ~q[5] /*29703*/;
  assign _6022_ = sum_27[23] & q[5] /*29702*/;
  assign _6023_ = m_27[23] & _6021_ /*29701*/;
  assign r_27[28] = _6023_ | _6022_ /*29700*/;
  assign _6024_ = ~q[5] /*29699*/;
  assign _6025_ = sum_27[24] & q[5] /*29698*/;
  assign _6026_ = m_27[24] & _6024_ /*29697*/;
  assign r_27[29] = _6026_ | _6025_ /*29696*/;
  assign _6027_ = ~q[5] /*29695*/;
  assign _6028_ = sum_27[25] & q[5] /*29694*/;
  assign _6029_ = m_27[25] & _6027_ /*29693*/;
  assign r_27[30] = _6029_ | _6028_ /*29692*/;
  assign _6030_ = ~q[5] /*29691*/;
  assign _6031_ = sum_27[26] & q[5] /*29690*/;
  assign _6032_ = m_27[26] & _6030_ /*29689*/;
  assign r_27[31] = _6032_ | _6031_ /*29688*/;
  assign _6033_ = ~q[5] /*29687*/;
  assign _6034_ = sum_27[27] & q[5] /*29686*/;
  assign _6035_ = m_27[27] & _6033_ /*29685*/;
  assign r_27[32] = _6035_ | _6034_ /*29684*/;
  assign _6036_ = ~q[5] /*29683*/;
  assign _6037_ = sum_27[28] & q[5] /*29682*/;
  assign _6038_ = m_27[28] & _6036_ /*29681*/;
  assign r_27[33] = _6038_ | _6037_ /*29680*/;
  assign _6039_ = ~q[5] /*29679*/;
  assign _6040_ = sum_27[29] & q[5] /*29678*/;
  assign _6041_ = m_27[29] & _6039_ /*29677*/;
  assign r_27[34] = _6041_ | _6040_ /*29676*/;
  assign _6042_ = ~q[5] /*29675*/;
  assign _6043_ = sum_27[30] & q[5] /*29674*/;
  assign _6044_ = m_27[30] & _6042_ /*29673*/;
  assign r_27[35] = _6044_ | _6043_ /*29672*/;
  assign _6045_ = ~q[5] /*29671*/;
  assign _6046_ = sum_27[31] & q[5] /*29670*/;
  assign _6047_ = m_27[31] & _6045_ /*29669*/;
  assign r_27[36] = _6047_ | _6046_ /*29668*/;
assign r_27[0]= r_26[0] /*29667*/;
assign r_27[1]= r_26[1] /*29666*/;
assign r_27[2]= r_26[2] /*29665*/;
assign r_27[3]= r_26[3] /*29664*/;
assign r_27[4]= r_26[4] /*29663*/;
  assign inv_28[0] = ~div[0] /*29576*/;
  assign inv_28[1] = ~div[1] /*29575*/;
  assign inv_28[2] = ~div[2] /*29574*/;
  assign inv_28[3] = ~div[3] /*29573*/;
  assign inv_28[4] = ~div[4] /*29572*/;
  assign inv_28[5] = ~div[5] /*29571*/;
  assign inv_28[6] = ~div[6] /*29570*/;
  assign inv_28[7] = ~div[7] /*29569*/;
  assign inv_28[8] = ~div[8] /*29568*/;
  assign inv_28[9] = ~div[9] /*29567*/;
  assign inv_28[10] = ~div[10] /*29566*/;
  assign inv_28[11] = ~div[11] /*29565*/;
  assign inv_28[12] = ~div[12] /*29564*/;
  assign inv_28[13] = ~div[13] /*29563*/;
  assign inv_28[14] = ~div[14] /*29562*/;
  assign inv_28[15] = ~div[15] /*29561*/;
  assign inv_28[16] = ~div[16] /*29560*/;
  assign inv_28[17] = ~div[17] /*29559*/;
  assign inv_28[18] = ~div[18] /*29558*/;
  assign inv_28[19] = ~div[19] /*29557*/;
  assign inv_28[20] = ~div[20] /*29556*/;
  assign inv_28[21] = ~div[21] /*29555*/;
  assign inv_28[22] = ~div[22] /*29554*/;
  assign inv_28[23] = ~div[23] /*29553*/;
  assign inv_28[24] = ~div[24] /*29552*/;
  assign inv_28[25] = ~div[25] /*29551*/;
  assign inv_28[26] = ~div[26] /*29550*/;
  assign inv_28[27] = ~div[27] /*29549*/;
  assign inv_28[28] = ~div[28] /*29548*/;
  assign inv_28[29] = ~div[29] /*29547*/;
  assign inv_28[30] = ~div[30] /*29546*/;
assign inv_28[31] = oneWire /*29545*/;
  assign _6048_ = inv_28[0] ^ r_27[4] /*29543*/;
  assign sum_28[0] = _6048_ ^ oneWire /*29542*/;
  assign _6049_ = _6048_ & oneWire /*29541*/;
  assign _6050_ = inv_28[0] & r_27[4] /*29540*/;
  assign _6051_ = _6049_ | _6050_ /*29539*/;
  assign _6052_ = inv_28[1] ^ r_27[5] /*29538*/;
  assign sum_28[1] = _6052_ ^ _6051_ /*29537*/;
  assign _6053_ = _6052_ & _6051_ /*29536*/;
  assign _6054_ = inv_28[1] & r_27[5] /*29535*/;
  assign _6055_ = _6053_ | _6054_ /*29534*/;
  assign _6056_ = inv_28[2] ^ r_27[6] /*29532*/;
  assign sum_28[2] = _6056_ ^ _6055_ /*29531*/;
  assign _6057_ = _6056_ & _6055_ /*29530*/;
  assign _6058_ = inv_28[2] & r_27[6] /*29529*/;
  assign _6059_ = _6057_ | _6058_ /*29528*/;
  assign _6060_ = inv_28[3] ^ r_27[7] /*29526*/;
  assign sum_28[3] = _6060_ ^ _6059_ /*29525*/;
  assign _6061_ = _6060_ & _6059_ /*29524*/;
  assign _6062_ = inv_28[3] & r_27[7] /*29523*/;
  assign _6063_ = _6061_ | _6062_ /*29522*/;
  assign _6064_ = inv_28[4] ^ r_27[8] /*29520*/;
  assign sum_28[4] = _6064_ ^ _6063_ /*29519*/;
  assign _6065_ = _6064_ & _6063_ /*29518*/;
  assign _6066_ = inv_28[4] & r_27[8] /*29517*/;
  assign _6067_ = _6065_ | _6066_ /*29516*/;
  assign _6068_ = inv_28[5] ^ r_27[9] /*29514*/;
  assign sum_28[5] = _6068_ ^ _6067_ /*29513*/;
  assign _6069_ = _6068_ & _6067_ /*29512*/;
  assign _6070_ = inv_28[5] & r_27[9] /*29511*/;
  assign _6071_ = _6069_ | _6070_ /*29510*/;
  assign _6072_ = inv_28[6] ^ r_27[10] /*29508*/;
  assign sum_28[6] = _6072_ ^ _6071_ /*29507*/;
  assign _6073_ = _6072_ & _6071_ /*29506*/;
  assign _6074_ = inv_28[6] & r_27[10] /*29505*/;
  assign _6075_ = _6073_ | _6074_ /*29504*/;
  assign _6076_ = inv_28[7] ^ r_27[11] /*29502*/;
  assign sum_28[7] = _6076_ ^ _6075_ /*29501*/;
  assign _6077_ = _6076_ & _6075_ /*29500*/;
  assign _6078_ = inv_28[7] & r_27[11] /*29499*/;
  assign _6079_ = _6077_ | _6078_ /*29498*/;
  assign _6080_ = inv_28[8] ^ r_27[12] /*29496*/;
  assign sum_28[8] = _6080_ ^ _6079_ /*29495*/;
  assign _6081_ = _6080_ & _6079_ /*29494*/;
  assign _6082_ = inv_28[8] & r_27[12] /*29493*/;
  assign _6083_ = _6081_ | _6082_ /*29492*/;
  assign _6084_ = inv_28[9] ^ r_27[13] /*29490*/;
  assign sum_28[9] = _6084_ ^ _6083_ /*29489*/;
  assign _6085_ = _6084_ & _6083_ /*29488*/;
  assign _6086_ = inv_28[9] & r_27[13] /*29487*/;
  assign _6087_ = _6085_ | _6086_ /*29486*/;
  assign _6088_ = inv_28[10] ^ r_27[14] /*29484*/;
  assign sum_28[10] = _6088_ ^ _6087_ /*29483*/;
  assign _6089_ = _6088_ & _6087_ /*29482*/;
  assign _6090_ = inv_28[10] & r_27[14] /*29481*/;
  assign _6091_ = _6089_ | _6090_ /*29480*/;
  assign _6092_ = inv_28[11] ^ r_27[15] /*29478*/;
  assign sum_28[11] = _6092_ ^ _6091_ /*29477*/;
  assign _6093_ = _6092_ & _6091_ /*29476*/;
  assign _6094_ = inv_28[11] & r_27[15] /*29475*/;
  assign _6095_ = _6093_ | _6094_ /*29474*/;
  assign _6096_ = inv_28[12] ^ r_27[16] /*29472*/;
  assign sum_28[12] = _6096_ ^ _6095_ /*29471*/;
  assign _6097_ = _6096_ & _6095_ /*29470*/;
  assign _6098_ = inv_28[12] & r_27[16] /*29469*/;
  assign _6099_ = _6097_ | _6098_ /*29468*/;
  assign _6100_ = inv_28[13] ^ r_27[17] /*29466*/;
  assign sum_28[13] = _6100_ ^ _6099_ /*29465*/;
  assign _6101_ = _6100_ & _6099_ /*29464*/;
  assign _6102_ = inv_28[13] & r_27[17] /*29463*/;
  assign _6103_ = _6101_ | _6102_ /*29462*/;
  assign _6104_ = inv_28[14] ^ r_27[18] /*29460*/;
  assign sum_28[14] = _6104_ ^ _6103_ /*29459*/;
  assign _6105_ = _6104_ & _6103_ /*29458*/;
  assign _6106_ = inv_28[14] & r_27[18] /*29457*/;
  assign _6107_ = _6105_ | _6106_ /*29456*/;
  assign _6108_ = inv_28[15] ^ r_27[19] /*29454*/;
  assign sum_28[15] = _6108_ ^ _6107_ /*29453*/;
  assign _6109_ = _6108_ & _6107_ /*29452*/;
  assign _6110_ = inv_28[15] & r_27[19] /*29451*/;
  assign _6111_ = _6109_ | _6110_ /*29450*/;
  assign _6112_ = inv_28[16] ^ r_27[20] /*29448*/;
  assign sum_28[16] = _6112_ ^ _6111_ /*29447*/;
  assign _6113_ = _6112_ & _6111_ /*29446*/;
  assign _6114_ = inv_28[16] & r_27[20] /*29445*/;
  assign _6115_ = _6113_ | _6114_ /*29444*/;
  assign _6116_ = inv_28[17] ^ r_27[21] /*29442*/;
  assign sum_28[17] = _6116_ ^ _6115_ /*29441*/;
  assign _6117_ = _6116_ & _6115_ /*29440*/;
  assign _6118_ = inv_28[17] & r_27[21] /*29439*/;
  assign _6119_ = _6117_ | _6118_ /*29438*/;
  assign _6120_ = inv_28[18] ^ r_27[22] /*29436*/;
  assign sum_28[18] = _6120_ ^ _6119_ /*29435*/;
  assign _6121_ = _6120_ & _6119_ /*29434*/;
  assign _6122_ = inv_28[18] & r_27[22] /*29433*/;
  assign _6123_ = _6121_ | _6122_ /*29432*/;
  assign _6124_ = inv_28[19] ^ r_27[23] /*29430*/;
  assign sum_28[19] = _6124_ ^ _6123_ /*29429*/;
  assign _6125_ = _6124_ & _6123_ /*29428*/;
  assign _6126_ = inv_28[19] & r_27[23] /*29427*/;
  assign _6127_ = _6125_ | _6126_ /*29426*/;
  assign _6128_ = inv_28[20] ^ r_27[24] /*29424*/;
  assign sum_28[20] = _6128_ ^ _6127_ /*29423*/;
  assign _6129_ = _6128_ & _6127_ /*29422*/;
  assign _6130_ = inv_28[20] & r_27[24] /*29421*/;
  assign _6131_ = _6129_ | _6130_ /*29420*/;
  assign _6132_ = inv_28[21] ^ r_27[25] /*29418*/;
  assign sum_28[21] = _6132_ ^ _6131_ /*29417*/;
  assign _6133_ = _6132_ & _6131_ /*29416*/;
  assign _6134_ = inv_28[21] & r_27[25] /*29415*/;
  assign _6135_ = _6133_ | _6134_ /*29414*/;
  assign _6136_ = inv_28[22] ^ r_27[26] /*29412*/;
  assign sum_28[22] = _6136_ ^ _6135_ /*29411*/;
  assign _6137_ = _6136_ & _6135_ /*29410*/;
  assign _6138_ = inv_28[22] & r_27[26] /*29409*/;
  assign _6139_ = _6137_ | _6138_ /*29408*/;
  assign _6140_ = inv_28[23] ^ r_27[27] /*29406*/;
  assign sum_28[23] = _6140_ ^ _6139_ /*29405*/;
  assign _6141_ = _6140_ & _6139_ /*29404*/;
  assign _6142_ = inv_28[23] & r_27[27] /*29403*/;
  assign _6143_ = _6141_ | _6142_ /*29402*/;
  assign _6144_ = inv_28[24] ^ r_27[28] /*29400*/;
  assign sum_28[24] = _6144_ ^ _6143_ /*29399*/;
  assign _6145_ = _6144_ & _6143_ /*29398*/;
  assign _6146_ = inv_28[24] & r_27[28] /*29397*/;
  assign _6147_ = _6145_ | _6146_ /*29396*/;
  assign _6148_ = inv_28[25] ^ r_27[29] /*29394*/;
  assign sum_28[25] = _6148_ ^ _6147_ /*29393*/;
  assign _6149_ = _6148_ & _6147_ /*29392*/;
  assign _6150_ = inv_28[25] & r_27[29] /*29391*/;
  assign _6151_ = _6149_ | _6150_ /*29390*/;
  assign _6152_ = inv_28[26] ^ r_27[30] /*29388*/;
  assign sum_28[26] = _6152_ ^ _6151_ /*29387*/;
  assign _6153_ = _6152_ & _6151_ /*29386*/;
  assign _6154_ = inv_28[26] & r_27[30] /*29385*/;
  assign _6155_ = _6153_ | _6154_ /*29384*/;
  assign _6156_ = inv_28[27] ^ r_27[31] /*29382*/;
  assign sum_28[27] = _6156_ ^ _6155_ /*29381*/;
  assign _6157_ = _6156_ & _6155_ /*29380*/;
  assign _6158_ = inv_28[27] & r_27[31] /*29379*/;
  assign _6159_ = _6157_ | _6158_ /*29378*/;
  assign _6160_ = inv_28[28] ^ r_27[32] /*29376*/;
  assign sum_28[28] = _6160_ ^ _6159_ /*29375*/;
  assign _6161_ = _6160_ & _6159_ /*29374*/;
  assign _6162_ = inv_28[28] & r_27[32] /*29373*/;
  assign _6163_ = _6161_ | _6162_ /*29372*/;
  assign _6164_ = inv_28[29] ^ r_27[33] /*29370*/;
  assign sum_28[29] = _6164_ ^ _6163_ /*29369*/;
  assign _6165_ = _6164_ & _6163_ /*29368*/;
  assign _6166_ = inv_28[29] & r_27[33] /*29367*/;
  assign _6167_ = _6165_ | _6166_ /*29366*/;
  assign _6168_ = inv_28[30] ^ r_27[34] /*29364*/;
  assign sum_28[30] = _6168_ ^ _6167_ /*29363*/;
  assign _6169_ = _6168_ & _6167_ /*29362*/;
  assign _6170_ = inv_28[30] & r_27[34] /*29361*/;
  assign _6171_ = _6169_ | _6170_ /*29360*/;
  assign _6172_ = inv_28[31] ^ r_27[35] /*29358*/;
  assign sum_28[31] = _6172_ ^ _6171_ /*29357*/;
  assign _6173_ = _6172_ & _6171_ /*29356*/;
  assign _6174_ = inv_28[31] & r_27[35] /*29355*/;
  assign _6175_ = _6173_ | _6174_ /*29354*/;
  assign q[4] = ~sum_28[31] /*29381*/;
  assign m_28[0] = r_27[4] /*29380*/;
  assign m_28[1] = r_27[5] /*29379*/;
  assign m_28[2] = r_27[6] /*29378*/;
  assign m_28[3] = r_27[7] /*29377*/;
  assign m_28[4] = r_27[8] /*29376*/;
  assign m_28[5] = r_27[9] /*29375*/;
  assign m_28[6] = r_27[10] /*29374*/;
  assign m_28[7] = r_27[11] /*29373*/;
  assign m_28[8] = r_27[12] /*29372*/;
  assign m_28[9] = r_27[13] /*29371*/;
  assign m_28[10] = r_27[14] /*29370*/;
  assign m_28[11] = r_27[15] /*29369*/;
  assign m_28[12] = r_27[16] /*29368*/;
  assign m_28[13] = r_27[17] /*29367*/;
  assign m_28[14] = r_27[18] /*29366*/;
  assign m_28[15] = r_27[19] /*29365*/;
  assign m_28[16] = r_27[20] /*29364*/;
  assign m_28[17] = r_27[21] /*29363*/;
  assign m_28[18] = r_27[22] /*29362*/;
  assign m_28[19] = r_27[23] /*29361*/;
  assign m_28[20] = r_27[24] /*29360*/;
  assign m_28[21] = r_27[25] /*29359*/;
  assign m_28[22] = r_27[26] /*29358*/;
  assign m_28[23] = r_27[27] /*29357*/;
  assign m_28[24] = r_27[28] /*29356*/;
  assign m_28[25] = r_27[29] /*29355*/;
  assign m_28[26] = r_27[30] /*29354*/;
  assign m_28[27] = r_27[31] /*29353*/;
  assign m_28[28] = r_27[32] /*29352*/;
  assign m_28[29] = r_27[33] /*29351*/;
  assign m_28[30] = r_27[34] /*29350*/;
  assign m_28[31] = r_27[35] /*29349*/;
  assign _6176_ = ~q[4] /*29347*/;
  assign _6177_ = sum_28[0] & q[4] /*29346*/;
  assign _6178_ = m_28[0] & _6176_ /*29345*/;
  assign r_28[4] = _6178_ | _6177_ /*29344*/;
  assign _6179_ = ~q[4] /*29343*/;
  assign _6180_ = sum_28[1] & q[4] /*29342*/;
  assign _6181_ = m_28[1] & _6179_ /*29341*/;
  assign r_28[5] = _6181_ | _6180_ /*29340*/;
  assign _6182_ = ~q[4] /*29339*/;
  assign _6183_ = sum_28[2] & q[4] /*29338*/;
  assign _6184_ = m_28[2] & _6182_ /*29337*/;
  assign r_28[6] = _6184_ | _6183_ /*29336*/;
  assign _6185_ = ~q[4] /*29335*/;
  assign _6186_ = sum_28[3] & q[4] /*29334*/;
  assign _6187_ = m_28[3] & _6185_ /*29333*/;
  assign r_28[7] = _6187_ | _6186_ /*29332*/;
  assign _6188_ = ~q[4] /*29331*/;
  assign _6189_ = sum_28[4] & q[4] /*29330*/;
  assign _6190_ = m_28[4] & _6188_ /*29329*/;
  assign r_28[8] = _6190_ | _6189_ /*29328*/;
  assign _6191_ = ~q[4] /*29327*/;
  assign _6192_ = sum_28[5] & q[4] /*29326*/;
  assign _6193_ = m_28[5] & _6191_ /*29325*/;
  assign r_28[9] = _6193_ | _6192_ /*29324*/;
  assign _6194_ = ~q[4] /*29323*/;
  assign _6195_ = sum_28[6] & q[4] /*29322*/;
  assign _6196_ = m_28[6] & _6194_ /*29321*/;
  assign r_28[10] = _6196_ | _6195_ /*29320*/;
  assign _6197_ = ~q[4] /*29319*/;
  assign _6198_ = sum_28[7] & q[4] /*29318*/;
  assign _6199_ = m_28[7] & _6197_ /*29317*/;
  assign r_28[11] = _6199_ | _6198_ /*29316*/;
  assign _6200_ = ~q[4] /*29315*/;
  assign _6201_ = sum_28[8] & q[4] /*29314*/;
  assign _6202_ = m_28[8] & _6200_ /*29313*/;
  assign r_28[12] = _6202_ | _6201_ /*29312*/;
  assign _6203_ = ~q[4] /*29311*/;
  assign _6204_ = sum_28[9] & q[4] /*29310*/;
  assign _6205_ = m_28[9] & _6203_ /*29309*/;
  assign r_28[13] = _6205_ | _6204_ /*29308*/;
  assign _6206_ = ~q[4] /*29307*/;
  assign _6207_ = sum_28[10] & q[4] /*29306*/;
  assign _6208_ = m_28[10] & _6206_ /*29305*/;
  assign r_28[14] = _6208_ | _6207_ /*29304*/;
  assign _6209_ = ~q[4] /*29303*/;
  assign _6210_ = sum_28[11] & q[4] /*29302*/;
  assign _6211_ = m_28[11] & _6209_ /*29301*/;
  assign r_28[15] = _6211_ | _6210_ /*29300*/;
  assign _6212_ = ~q[4] /*29299*/;
  assign _6213_ = sum_28[12] & q[4] /*29298*/;
  assign _6214_ = m_28[12] & _6212_ /*29297*/;
  assign r_28[16] = _6214_ | _6213_ /*29296*/;
  assign _6215_ = ~q[4] /*29295*/;
  assign _6216_ = sum_28[13] & q[4] /*29294*/;
  assign _6217_ = m_28[13] & _6215_ /*29293*/;
  assign r_28[17] = _6217_ | _6216_ /*29292*/;
  assign _6218_ = ~q[4] /*29291*/;
  assign _6219_ = sum_28[14] & q[4] /*29290*/;
  assign _6220_ = m_28[14] & _6218_ /*29289*/;
  assign r_28[18] = _6220_ | _6219_ /*29288*/;
  assign _6221_ = ~q[4] /*29287*/;
  assign _6222_ = sum_28[15] & q[4] /*29286*/;
  assign _6223_ = m_28[15] & _6221_ /*29285*/;
  assign r_28[19] = _6223_ | _6222_ /*29284*/;
  assign _6224_ = ~q[4] /*29283*/;
  assign _6225_ = sum_28[16] & q[4] /*29282*/;
  assign _6226_ = m_28[16] & _6224_ /*29281*/;
  assign r_28[20] = _6226_ | _6225_ /*29280*/;
  assign _6227_ = ~q[4] /*29279*/;
  assign _6228_ = sum_28[17] & q[4] /*29278*/;
  assign _6229_ = m_28[17] & _6227_ /*29277*/;
  assign r_28[21] = _6229_ | _6228_ /*29276*/;
  assign _6230_ = ~q[4] /*29275*/;
  assign _6231_ = sum_28[18] & q[4] /*29274*/;
  assign _6232_ = m_28[18] & _6230_ /*29273*/;
  assign r_28[22] = _6232_ | _6231_ /*29272*/;
  assign _6233_ = ~q[4] /*29271*/;
  assign _6234_ = sum_28[19] & q[4] /*29270*/;
  assign _6235_ = m_28[19] & _6233_ /*29269*/;
  assign r_28[23] = _6235_ | _6234_ /*29268*/;
  assign _6236_ = ~q[4] /*29267*/;
  assign _6237_ = sum_28[20] & q[4] /*29266*/;
  assign _6238_ = m_28[20] & _6236_ /*29265*/;
  assign r_28[24] = _6238_ | _6237_ /*29264*/;
  assign _6239_ = ~q[4] /*29263*/;
  assign _6240_ = sum_28[21] & q[4] /*29262*/;
  assign _6241_ = m_28[21] & _6239_ /*29261*/;
  assign r_28[25] = _6241_ | _6240_ /*29260*/;
  assign _6242_ = ~q[4] /*29259*/;
  assign _6243_ = sum_28[22] & q[4] /*29258*/;
  assign _6244_ = m_28[22] & _6242_ /*29257*/;
  assign r_28[26] = _6244_ | _6243_ /*29256*/;
  assign _6245_ = ~q[4] /*29255*/;
  assign _6246_ = sum_28[23] & q[4] /*29254*/;
  assign _6247_ = m_28[23] & _6245_ /*29253*/;
  assign r_28[27] = _6247_ | _6246_ /*29252*/;
  assign _6248_ = ~q[4] /*29251*/;
  assign _6249_ = sum_28[24] & q[4] /*29250*/;
  assign _6250_ = m_28[24] & _6248_ /*29249*/;
  assign r_28[28] = _6250_ | _6249_ /*29248*/;
  assign _6251_ = ~q[4] /*29247*/;
  assign _6252_ = sum_28[25] & q[4] /*29246*/;
  assign _6253_ = m_28[25] & _6251_ /*29245*/;
  assign r_28[29] = _6253_ | _6252_ /*29244*/;
  assign _6254_ = ~q[4] /*29243*/;
  assign _6255_ = sum_28[26] & q[4] /*29242*/;
  assign _6256_ = m_28[26] & _6254_ /*29241*/;
  assign r_28[30] = _6256_ | _6255_ /*29240*/;
  assign _6257_ = ~q[4] /*29239*/;
  assign _6258_ = sum_28[27] & q[4] /*29238*/;
  assign _6259_ = m_28[27] & _6257_ /*29237*/;
  assign r_28[31] = _6259_ | _6258_ /*29236*/;
  assign _6260_ = ~q[4] /*29235*/;
  assign _6261_ = sum_28[28] & q[4] /*29234*/;
  assign _6262_ = m_28[28] & _6260_ /*29233*/;
  assign r_28[32] = _6262_ | _6261_ /*29232*/;
  assign _6263_ = ~q[4] /*29231*/;
  assign _6264_ = sum_28[29] & q[4] /*29230*/;
  assign _6265_ = m_28[29] & _6263_ /*29229*/;
  assign r_28[33] = _6265_ | _6264_ /*29228*/;
  assign _6266_ = ~q[4] /*29227*/;
  assign _6267_ = sum_28[30] & q[4] /*29226*/;
  assign _6268_ = m_28[30] & _6266_ /*29225*/;
  assign r_28[34] = _6268_ | _6267_ /*29224*/;
  assign _6269_ = ~q[4] /*29223*/;
  assign _6270_ = sum_28[31] & q[4] /*29222*/;
  assign _6271_ = m_28[31] & _6269_ /*29221*/;
  assign r_28[35] = _6271_ | _6270_ /*29220*/;
assign r_28[0]= r_27[0] /*29219*/;
assign r_28[1]= r_27[1] /*29218*/;
assign r_28[2]= r_27[2] /*29217*/;
assign r_28[3]= r_27[3] /*29216*/;
  assign inv_29[0] = ~div[0] /*29128*/;
  assign inv_29[1] = ~div[1] /*29127*/;
  assign inv_29[2] = ~div[2] /*29126*/;
  assign inv_29[3] = ~div[3] /*29125*/;
  assign inv_29[4] = ~div[4] /*29124*/;
  assign inv_29[5] = ~div[5] /*29123*/;
  assign inv_29[6] = ~div[6] /*29122*/;
  assign inv_29[7] = ~div[7] /*29121*/;
  assign inv_29[8] = ~div[8] /*29120*/;
  assign inv_29[9] = ~div[9] /*29119*/;
  assign inv_29[10] = ~div[10] /*29118*/;
  assign inv_29[11] = ~div[11] /*29117*/;
  assign inv_29[12] = ~div[12] /*29116*/;
  assign inv_29[13] = ~div[13] /*29115*/;
  assign inv_29[14] = ~div[14] /*29114*/;
  assign inv_29[15] = ~div[15] /*29113*/;
  assign inv_29[16] = ~div[16] /*29112*/;
  assign inv_29[17] = ~div[17] /*29111*/;
  assign inv_29[18] = ~div[18] /*29110*/;
  assign inv_29[19] = ~div[19] /*29109*/;
  assign inv_29[20] = ~div[20] /*29108*/;
  assign inv_29[21] = ~div[21] /*29107*/;
  assign inv_29[22] = ~div[22] /*29106*/;
  assign inv_29[23] = ~div[23] /*29105*/;
  assign inv_29[24] = ~div[24] /*29104*/;
  assign inv_29[25] = ~div[25] /*29103*/;
  assign inv_29[26] = ~div[26] /*29102*/;
  assign inv_29[27] = ~div[27] /*29101*/;
  assign inv_29[28] = ~div[28] /*29100*/;
  assign inv_29[29] = ~div[29] /*29099*/;
  assign inv_29[30] = ~div[30] /*29098*/;
assign inv_29[31] = oneWire /*29097*/;
  assign _6272_ = inv_29[0] ^ r_28[3] /*29095*/;
  assign sum_29[0] = _6272_ ^ oneWire /*29094*/;
  assign _6273_ = _6272_ & oneWire /*29093*/;
  assign _6274_ = inv_29[0] & r_28[3] /*29092*/;
  assign _6275_ = _6273_ | _6274_ /*29091*/;
  assign _6276_ = inv_29[1] ^ r_28[4] /*29090*/;
  assign sum_29[1] = _6276_ ^ _6275_ /*29089*/;
  assign _6277_ = _6276_ & _6275_ /*29088*/;
  assign _6278_ = inv_29[1] & r_28[4] /*29087*/;
  assign _6279_ = _6277_ | _6278_ /*29086*/;
  assign _6280_ = inv_29[2] ^ r_28[5] /*29084*/;
  assign sum_29[2] = _6280_ ^ _6279_ /*29083*/;
  assign _6281_ = _6280_ & _6279_ /*29082*/;
  assign _6282_ = inv_29[2] & r_28[5] /*29081*/;
  assign _6283_ = _6281_ | _6282_ /*29080*/;
  assign _6284_ = inv_29[3] ^ r_28[6] /*29078*/;
  assign sum_29[3] = _6284_ ^ _6283_ /*29077*/;
  assign _6285_ = _6284_ & _6283_ /*29076*/;
  assign _6286_ = inv_29[3] & r_28[6] /*29075*/;
  assign _6287_ = _6285_ | _6286_ /*29074*/;
  assign _6288_ = inv_29[4] ^ r_28[7] /*29072*/;
  assign sum_29[4] = _6288_ ^ _6287_ /*29071*/;
  assign _6289_ = _6288_ & _6287_ /*29070*/;
  assign _6290_ = inv_29[4] & r_28[7] /*29069*/;
  assign _6291_ = _6289_ | _6290_ /*29068*/;
  assign _6292_ = inv_29[5] ^ r_28[8] /*29066*/;
  assign sum_29[5] = _6292_ ^ _6291_ /*29065*/;
  assign _6293_ = _6292_ & _6291_ /*29064*/;
  assign _6294_ = inv_29[5] & r_28[8] /*29063*/;
  assign _6295_ = _6293_ | _6294_ /*29062*/;
  assign _6296_ = inv_29[6] ^ r_28[9] /*29060*/;
  assign sum_29[6] = _6296_ ^ _6295_ /*29059*/;
  assign _6297_ = _6296_ & _6295_ /*29058*/;
  assign _6298_ = inv_29[6] & r_28[9] /*29057*/;
  assign _6299_ = _6297_ | _6298_ /*29056*/;
  assign _6300_ = inv_29[7] ^ r_28[10] /*29054*/;
  assign sum_29[7] = _6300_ ^ _6299_ /*29053*/;
  assign _6301_ = _6300_ & _6299_ /*29052*/;
  assign _6302_ = inv_29[7] & r_28[10] /*29051*/;
  assign _6303_ = _6301_ | _6302_ /*29050*/;
  assign _6304_ = inv_29[8] ^ r_28[11] /*29048*/;
  assign sum_29[8] = _6304_ ^ _6303_ /*29047*/;
  assign _6305_ = _6304_ & _6303_ /*29046*/;
  assign _6306_ = inv_29[8] & r_28[11] /*29045*/;
  assign _6307_ = _6305_ | _6306_ /*29044*/;
  assign _6308_ = inv_29[9] ^ r_28[12] /*29042*/;
  assign sum_29[9] = _6308_ ^ _6307_ /*29041*/;
  assign _6309_ = _6308_ & _6307_ /*29040*/;
  assign _6310_ = inv_29[9] & r_28[12] /*29039*/;
  assign _6311_ = _6309_ | _6310_ /*29038*/;
  assign _6312_ = inv_29[10] ^ r_28[13] /*29036*/;
  assign sum_29[10] = _6312_ ^ _6311_ /*29035*/;
  assign _6313_ = _6312_ & _6311_ /*29034*/;
  assign _6314_ = inv_29[10] & r_28[13] /*29033*/;
  assign _6315_ = _6313_ | _6314_ /*29032*/;
  assign _6316_ = inv_29[11] ^ r_28[14] /*29030*/;
  assign sum_29[11] = _6316_ ^ _6315_ /*29029*/;
  assign _6317_ = _6316_ & _6315_ /*29028*/;
  assign _6318_ = inv_29[11] & r_28[14] /*29027*/;
  assign _6319_ = _6317_ | _6318_ /*29026*/;
  assign _6320_ = inv_29[12] ^ r_28[15] /*29024*/;
  assign sum_29[12] = _6320_ ^ _6319_ /*29023*/;
  assign _6321_ = _6320_ & _6319_ /*29022*/;
  assign _6322_ = inv_29[12] & r_28[15] /*29021*/;
  assign _6323_ = _6321_ | _6322_ /*29020*/;
  assign _6324_ = inv_29[13] ^ r_28[16] /*29018*/;
  assign sum_29[13] = _6324_ ^ _6323_ /*29017*/;
  assign _6325_ = _6324_ & _6323_ /*29016*/;
  assign _6326_ = inv_29[13] & r_28[16] /*29015*/;
  assign _6327_ = _6325_ | _6326_ /*29014*/;
  assign _6328_ = inv_29[14] ^ r_28[17] /*29012*/;
  assign sum_29[14] = _6328_ ^ _6327_ /*29011*/;
  assign _6329_ = _6328_ & _6327_ /*29010*/;
  assign _6330_ = inv_29[14] & r_28[17] /*29009*/;
  assign _6331_ = _6329_ | _6330_ /*29008*/;
  assign _6332_ = inv_29[15] ^ r_28[18] /*29006*/;
  assign sum_29[15] = _6332_ ^ _6331_ /*29005*/;
  assign _6333_ = _6332_ & _6331_ /*29004*/;
  assign _6334_ = inv_29[15] & r_28[18] /*29003*/;
  assign _6335_ = _6333_ | _6334_ /*29002*/;
  assign _6336_ = inv_29[16] ^ r_28[19] /*29000*/;
  assign sum_29[16] = _6336_ ^ _6335_ /*28999*/;
  assign _6337_ = _6336_ & _6335_ /*28998*/;
  assign _6338_ = inv_29[16] & r_28[19] /*28997*/;
  assign _6339_ = _6337_ | _6338_ /*28996*/;
  assign _6340_ = inv_29[17] ^ r_28[20] /*28994*/;
  assign sum_29[17] = _6340_ ^ _6339_ /*28993*/;
  assign _6341_ = _6340_ & _6339_ /*28992*/;
  assign _6342_ = inv_29[17] & r_28[20] /*28991*/;
  assign _6343_ = _6341_ | _6342_ /*28990*/;
  assign _6344_ = inv_29[18] ^ r_28[21] /*28988*/;
  assign sum_29[18] = _6344_ ^ _6343_ /*28987*/;
  assign _6345_ = _6344_ & _6343_ /*28986*/;
  assign _6346_ = inv_29[18] & r_28[21] /*28985*/;
  assign _6347_ = _6345_ | _6346_ /*28984*/;
  assign _6348_ = inv_29[19] ^ r_28[22] /*28982*/;
  assign sum_29[19] = _6348_ ^ _6347_ /*28981*/;
  assign _6349_ = _6348_ & _6347_ /*28980*/;
  assign _6350_ = inv_29[19] & r_28[22] /*28979*/;
  assign _6351_ = _6349_ | _6350_ /*28978*/;
  assign _6352_ = inv_29[20] ^ r_28[23] /*28976*/;
  assign sum_29[20] = _6352_ ^ _6351_ /*28975*/;
  assign _6353_ = _6352_ & _6351_ /*28974*/;
  assign _6354_ = inv_29[20] & r_28[23] /*28973*/;
  assign _6355_ = _6353_ | _6354_ /*28972*/;
  assign _6356_ = inv_29[21] ^ r_28[24] /*28970*/;
  assign sum_29[21] = _6356_ ^ _6355_ /*28969*/;
  assign _6357_ = _6356_ & _6355_ /*28968*/;
  assign _6358_ = inv_29[21] & r_28[24] /*28967*/;
  assign _6359_ = _6357_ | _6358_ /*28966*/;
  assign _6360_ = inv_29[22] ^ r_28[25] /*28964*/;
  assign sum_29[22] = _6360_ ^ _6359_ /*28963*/;
  assign _6361_ = _6360_ & _6359_ /*28962*/;
  assign _6362_ = inv_29[22] & r_28[25] /*28961*/;
  assign _6363_ = _6361_ | _6362_ /*28960*/;
  assign _6364_ = inv_29[23] ^ r_28[26] /*28958*/;
  assign sum_29[23] = _6364_ ^ _6363_ /*28957*/;
  assign _6365_ = _6364_ & _6363_ /*28956*/;
  assign _6366_ = inv_29[23] & r_28[26] /*28955*/;
  assign _6367_ = _6365_ | _6366_ /*28954*/;
  assign _6368_ = inv_29[24] ^ r_28[27] /*28952*/;
  assign sum_29[24] = _6368_ ^ _6367_ /*28951*/;
  assign _6369_ = _6368_ & _6367_ /*28950*/;
  assign _6370_ = inv_29[24] & r_28[27] /*28949*/;
  assign _6371_ = _6369_ | _6370_ /*28948*/;
  assign _6372_ = inv_29[25] ^ r_28[28] /*28946*/;
  assign sum_29[25] = _6372_ ^ _6371_ /*28945*/;
  assign _6373_ = _6372_ & _6371_ /*28944*/;
  assign _6374_ = inv_29[25] & r_28[28] /*28943*/;
  assign _6375_ = _6373_ | _6374_ /*28942*/;
  assign _6376_ = inv_29[26] ^ r_28[29] /*28940*/;
  assign sum_29[26] = _6376_ ^ _6375_ /*28939*/;
  assign _6377_ = _6376_ & _6375_ /*28938*/;
  assign _6378_ = inv_29[26] & r_28[29] /*28937*/;
  assign _6379_ = _6377_ | _6378_ /*28936*/;
  assign _6380_ = inv_29[27] ^ r_28[30] /*28934*/;
  assign sum_29[27] = _6380_ ^ _6379_ /*28933*/;
  assign _6381_ = _6380_ & _6379_ /*28932*/;
  assign _6382_ = inv_29[27] & r_28[30] /*28931*/;
  assign _6383_ = _6381_ | _6382_ /*28930*/;
  assign _6384_ = inv_29[28] ^ r_28[31] /*28928*/;
  assign sum_29[28] = _6384_ ^ _6383_ /*28927*/;
  assign _6385_ = _6384_ & _6383_ /*28926*/;
  assign _6386_ = inv_29[28] & r_28[31] /*28925*/;
  assign _6387_ = _6385_ | _6386_ /*28924*/;
  assign _6388_ = inv_29[29] ^ r_28[32] /*28922*/;
  assign sum_29[29] = _6388_ ^ _6387_ /*28921*/;
  assign _6389_ = _6388_ & _6387_ /*28920*/;
  assign _6390_ = inv_29[29] & r_28[32] /*28919*/;
  assign _6391_ = _6389_ | _6390_ /*28918*/;
  assign _6392_ = inv_29[30] ^ r_28[33] /*28916*/;
  assign sum_29[30] = _6392_ ^ _6391_ /*28915*/;
  assign _6393_ = _6392_ & _6391_ /*28914*/;
  assign _6394_ = inv_29[30] & r_28[33] /*28913*/;
  assign _6395_ = _6393_ | _6394_ /*28912*/;
  assign _6396_ = inv_29[31] ^ r_28[34] /*28910*/;
  assign sum_29[31] = _6396_ ^ _6395_ /*28909*/;
  assign _6397_ = _6396_ & _6395_ /*28908*/;
  assign _6398_ = inv_29[31] & r_28[34] /*28907*/;
  assign _6399_ = _6397_ | _6398_ /*28906*/;
  assign q[3] = ~sum_29[31] /*28933*/;
  assign m_29[0] = r_28[3] /*28932*/;
  assign m_29[1] = r_28[4] /*28931*/;
  assign m_29[2] = r_28[5] /*28930*/;
  assign m_29[3] = r_28[6] /*28929*/;
  assign m_29[4] = r_28[7] /*28928*/;
  assign m_29[5] = r_28[8] /*28927*/;
  assign m_29[6] = r_28[9] /*28926*/;
  assign m_29[7] = r_28[10] /*28925*/;
  assign m_29[8] = r_28[11] /*28924*/;
  assign m_29[9] = r_28[12] /*28923*/;
  assign m_29[10] = r_28[13] /*28922*/;
  assign m_29[11] = r_28[14] /*28921*/;
  assign m_29[12] = r_28[15] /*28920*/;
  assign m_29[13] = r_28[16] /*28919*/;
  assign m_29[14] = r_28[17] /*28918*/;
  assign m_29[15] = r_28[18] /*28917*/;
  assign m_29[16] = r_28[19] /*28916*/;
  assign m_29[17] = r_28[20] /*28915*/;
  assign m_29[18] = r_28[21] /*28914*/;
  assign m_29[19] = r_28[22] /*28913*/;
  assign m_29[20] = r_28[23] /*28912*/;
  assign m_29[21] = r_28[24] /*28911*/;
  assign m_29[22] = r_28[25] /*28910*/;
  assign m_29[23] = r_28[26] /*28909*/;
  assign m_29[24] = r_28[27] /*28908*/;
  assign m_29[25] = r_28[28] /*28907*/;
  assign m_29[26] = r_28[29] /*28906*/;
  assign m_29[27] = r_28[30] /*28905*/;
  assign m_29[28] = r_28[31] /*28904*/;
  assign m_29[29] = r_28[32] /*28903*/;
  assign m_29[30] = r_28[33] /*28902*/;
  assign m_29[31] = r_28[34] /*28901*/;
  assign _6400_ = ~q[3] /*28899*/;
  assign _6401_ = sum_29[0] & q[3] /*28898*/;
  assign _6402_ = m_29[0] & _6400_ /*28897*/;
  assign r_29[3] = _6402_ | _6401_ /*28896*/;
  assign _6403_ = ~q[3] /*28895*/;
  assign _6404_ = sum_29[1] & q[3] /*28894*/;
  assign _6405_ = m_29[1] & _6403_ /*28893*/;
  assign r_29[4] = _6405_ | _6404_ /*28892*/;
  assign _6406_ = ~q[3] /*28891*/;
  assign _6407_ = sum_29[2] & q[3] /*28890*/;
  assign _6408_ = m_29[2] & _6406_ /*28889*/;
  assign r_29[5] = _6408_ | _6407_ /*28888*/;
  assign _6409_ = ~q[3] /*28887*/;
  assign _6410_ = sum_29[3] & q[3] /*28886*/;
  assign _6411_ = m_29[3] & _6409_ /*28885*/;
  assign r_29[6] = _6411_ | _6410_ /*28884*/;
  assign _6412_ = ~q[3] /*28883*/;
  assign _6413_ = sum_29[4] & q[3] /*28882*/;
  assign _6414_ = m_29[4] & _6412_ /*28881*/;
  assign r_29[7] = _6414_ | _6413_ /*28880*/;
  assign _6415_ = ~q[3] /*28879*/;
  assign _6416_ = sum_29[5] & q[3] /*28878*/;
  assign _6417_ = m_29[5] & _6415_ /*28877*/;
  assign r_29[8] = _6417_ | _6416_ /*28876*/;
  assign _6418_ = ~q[3] /*28875*/;
  assign _6419_ = sum_29[6] & q[3] /*28874*/;
  assign _6420_ = m_29[6] & _6418_ /*28873*/;
  assign r_29[9] = _6420_ | _6419_ /*28872*/;
  assign _6421_ = ~q[3] /*28871*/;
  assign _6422_ = sum_29[7] & q[3] /*28870*/;
  assign _6423_ = m_29[7] & _6421_ /*28869*/;
  assign r_29[10] = _6423_ | _6422_ /*28868*/;
  assign _6424_ = ~q[3] /*28867*/;
  assign _6425_ = sum_29[8] & q[3] /*28866*/;
  assign _6426_ = m_29[8] & _6424_ /*28865*/;
  assign r_29[11] = _6426_ | _6425_ /*28864*/;
  assign _6427_ = ~q[3] /*28863*/;
  assign _6428_ = sum_29[9] & q[3] /*28862*/;
  assign _6429_ = m_29[9] & _6427_ /*28861*/;
  assign r_29[12] = _6429_ | _6428_ /*28860*/;
  assign _6430_ = ~q[3] /*28859*/;
  assign _6431_ = sum_29[10] & q[3] /*28858*/;
  assign _6432_ = m_29[10] & _6430_ /*28857*/;
  assign r_29[13] = _6432_ | _6431_ /*28856*/;
  assign _6433_ = ~q[3] /*28855*/;
  assign _6434_ = sum_29[11] & q[3] /*28854*/;
  assign _6435_ = m_29[11] & _6433_ /*28853*/;
  assign r_29[14] = _6435_ | _6434_ /*28852*/;
  assign _6436_ = ~q[3] /*28851*/;
  assign _6437_ = sum_29[12] & q[3] /*28850*/;
  assign _6438_ = m_29[12] & _6436_ /*28849*/;
  assign r_29[15] = _6438_ | _6437_ /*28848*/;
  assign _6439_ = ~q[3] /*28847*/;
  assign _6440_ = sum_29[13] & q[3] /*28846*/;
  assign _6441_ = m_29[13] & _6439_ /*28845*/;
  assign r_29[16] = _6441_ | _6440_ /*28844*/;
  assign _6442_ = ~q[3] /*28843*/;
  assign _6443_ = sum_29[14] & q[3] /*28842*/;
  assign _6444_ = m_29[14] & _6442_ /*28841*/;
  assign r_29[17] = _6444_ | _6443_ /*28840*/;
  assign _6445_ = ~q[3] /*28839*/;
  assign _6446_ = sum_29[15] & q[3] /*28838*/;
  assign _6447_ = m_29[15] & _6445_ /*28837*/;
  assign r_29[18] = _6447_ | _6446_ /*28836*/;
  assign _6448_ = ~q[3] /*28835*/;
  assign _6449_ = sum_29[16] & q[3] /*28834*/;
  assign _6450_ = m_29[16] & _6448_ /*28833*/;
  assign r_29[19] = _6450_ | _6449_ /*28832*/;
  assign _6451_ = ~q[3] /*28831*/;
  assign _6452_ = sum_29[17] & q[3] /*28830*/;
  assign _6453_ = m_29[17] & _6451_ /*28829*/;
  assign r_29[20] = _6453_ | _6452_ /*28828*/;
  assign _6454_ = ~q[3] /*28827*/;
  assign _6455_ = sum_29[18] & q[3] /*28826*/;
  assign _6456_ = m_29[18] & _6454_ /*28825*/;
  assign r_29[21] = _6456_ | _6455_ /*28824*/;
  assign _6457_ = ~q[3] /*28823*/;
  assign _6458_ = sum_29[19] & q[3] /*28822*/;
  assign _6459_ = m_29[19] & _6457_ /*28821*/;
  assign r_29[22] = _6459_ | _6458_ /*28820*/;
  assign _6460_ = ~q[3] /*28819*/;
  assign _6461_ = sum_29[20] & q[3] /*28818*/;
  assign _6462_ = m_29[20] & _6460_ /*28817*/;
  assign r_29[23] = _6462_ | _6461_ /*28816*/;
  assign _6463_ = ~q[3] /*28815*/;
  assign _6464_ = sum_29[21] & q[3] /*28814*/;
  assign _6465_ = m_29[21] & _6463_ /*28813*/;
  assign r_29[24] = _6465_ | _6464_ /*28812*/;
  assign _6466_ = ~q[3] /*28811*/;
  assign _6467_ = sum_29[22] & q[3] /*28810*/;
  assign _6468_ = m_29[22] & _6466_ /*28809*/;
  assign r_29[25] = _6468_ | _6467_ /*28808*/;
  assign _6469_ = ~q[3] /*28807*/;
  assign _6470_ = sum_29[23] & q[3] /*28806*/;
  assign _6471_ = m_29[23] & _6469_ /*28805*/;
  assign r_29[26] = _6471_ | _6470_ /*28804*/;
  assign _6472_ = ~q[3] /*28803*/;
  assign _6473_ = sum_29[24] & q[3] /*28802*/;
  assign _6474_ = m_29[24] & _6472_ /*28801*/;
  assign r_29[27] = _6474_ | _6473_ /*28800*/;
  assign _6475_ = ~q[3] /*28799*/;
  assign _6476_ = sum_29[25] & q[3] /*28798*/;
  assign _6477_ = m_29[25] & _6475_ /*28797*/;
  assign r_29[28] = _6477_ | _6476_ /*28796*/;
  assign _6478_ = ~q[3] /*28795*/;
  assign _6479_ = sum_29[26] & q[3] /*28794*/;
  assign _6480_ = m_29[26] & _6478_ /*28793*/;
  assign r_29[29] = _6480_ | _6479_ /*28792*/;
  assign _6481_ = ~q[3] /*28791*/;
  assign _6482_ = sum_29[27] & q[3] /*28790*/;
  assign _6483_ = m_29[27] & _6481_ /*28789*/;
  assign r_29[30] = _6483_ | _6482_ /*28788*/;
  assign _6484_ = ~q[3] /*28787*/;
  assign _6485_ = sum_29[28] & q[3] /*28786*/;
  assign _6486_ = m_29[28] & _6484_ /*28785*/;
  assign r_29[31] = _6486_ | _6485_ /*28784*/;
  assign _6487_ = ~q[3] /*28783*/;
  assign _6488_ = sum_29[29] & q[3] /*28782*/;
  assign _6489_ = m_29[29] & _6487_ /*28781*/;
  assign r_29[32] = _6489_ | _6488_ /*28780*/;
  assign _6490_ = ~q[3] /*28779*/;
  assign _6491_ = sum_29[30] & q[3] /*28778*/;
  assign _6492_ = m_29[30] & _6490_ /*28777*/;
  assign r_29[33] = _6492_ | _6491_ /*28776*/;
  assign _6493_ = ~q[3] /*28775*/;
  assign _6494_ = sum_29[31] & q[3] /*28774*/;
  assign _6495_ = m_29[31] & _6493_ /*28773*/;
  assign r_29[34] = _6495_ | _6494_ /*28772*/;
assign r_29[0]= r_28[0] /*28771*/;
assign r_29[1]= r_28[1] /*28770*/;
assign r_29[2]= r_28[2] /*28769*/;
  assign inv_30[0] = ~div[0] /*28680*/;
  assign inv_30[1] = ~div[1] /*28679*/;
  assign inv_30[2] = ~div[2] /*28678*/;
  assign inv_30[3] = ~div[3] /*28677*/;
  assign inv_30[4] = ~div[4] /*28676*/;
  assign inv_30[5] = ~div[5] /*28675*/;
  assign inv_30[6] = ~div[6] /*28674*/;
  assign inv_30[7] = ~div[7] /*28673*/;
  assign inv_30[8] = ~div[8] /*28672*/;
  assign inv_30[9] = ~div[9] /*28671*/;
  assign inv_30[10] = ~div[10] /*28670*/;
  assign inv_30[11] = ~div[11] /*28669*/;
  assign inv_30[12] = ~div[12] /*28668*/;
  assign inv_30[13] = ~div[13] /*28667*/;
  assign inv_30[14] = ~div[14] /*28666*/;
  assign inv_30[15] = ~div[15] /*28665*/;
  assign inv_30[16] = ~div[16] /*28664*/;
  assign inv_30[17] = ~div[17] /*28663*/;
  assign inv_30[18] = ~div[18] /*28662*/;
  assign inv_30[19] = ~div[19] /*28661*/;
  assign inv_30[20] = ~div[20] /*28660*/;
  assign inv_30[21] = ~div[21] /*28659*/;
  assign inv_30[22] = ~div[22] /*28658*/;
  assign inv_30[23] = ~div[23] /*28657*/;
  assign inv_30[24] = ~div[24] /*28656*/;
  assign inv_30[25] = ~div[25] /*28655*/;
  assign inv_30[26] = ~div[26] /*28654*/;
  assign inv_30[27] = ~div[27] /*28653*/;
  assign inv_30[28] = ~div[28] /*28652*/;
  assign inv_30[29] = ~div[29] /*28651*/;
  assign inv_30[30] = ~div[30] /*28650*/;
assign inv_30[31] = oneWire /*28649*/;
  assign _6496_ = inv_30[0] ^ r_29[2] /*28647*/;
  assign sum_30[0] = _6496_ ^ oneWire /*28646*/;
  assign _6497_ = _6496_ & oneWire /*28645*/;
  assign _6498_ = inv_30[0] & r_29[2] /*28644*/;
  assign _6499_ = _6497_ | _6498_ /*28643*/;
  assign _6500_ = inv_30[1] ^ r_29[3] /*28642*/;
  assign sum_30[1] = _6500_ ^ _6499_ /*28641*/;
  assign _6501_ = _6500_ & _6499_ /*28640*/;
  assign _6502_ = inv_30[1] & r_29[3] /*28639*/;
  assign _6503_ = _6501_ | _6502_ /*28638*/;
  assign _6504_ = inv_30[2] ^ r_29[4] /*28636*/;
  assign sum_30[2] = _6504_ ^ _6503_ /*28635*/;
  assign _6505_ = _6504_ & _6503_ /*28634*/;
  assign _6506_ = inv_30[2] & r_29[4] /*28633*/;
  assign _6507_ = _6505_ | _6506_ /*28632*/;
  assign _6508_ = inv_30[3] ^ r_29[5] /*28630*/;
  assign sum_30[3] = _6508_ ^ _6507_ /*28629*/;
  assign _6509_ = _6508_ & _6507_ /*28628*/;
  assign _6510_ = inv_30[3] & r_29[5] /*28627*/;
  assign _6511_ = _6509_ | _6510_ /*28626*/;
  assign _6512_ = inv_30[4] ^ r_29[6] /*28624*/;
  assign sum_30[4] = _6512_ ^ _6511_ /*28623*/;
  assign _6513_ = _6512_ & _6511_ /*28622*/;
  assign _6514_ = inv_30[4] & r_29[6] /*28621*/;
  assign _6515_ = _6513_ | _6514_ /*28620*/;
  assign _6516_ = inv_30[5] ^ r_29[7] /*28618*/;
  assign sum_30[5] = _6516_ ^ _6515_ /*28617*/;
  assign _6517_ = _6516_ & _6515_ /*28616*/;
  assign _6518_ = inv_30[5] & r_29[7] /*28615*/;
  assign _6519_ = _6517_ | _6518_ /*28614*/;
  assign _6520_ = inv_30[6] ^ r_29[8] /*28612*/;
  assign sum_30[6] = _6520_ ^ _6519_ /*28611*/;
  assign _6521_ = _6520_ & _6519_ /*28610*/;
  assign _6522_ = inv_30[6] & r_29[8] /*28609*/;
  assign _6523_ = _6521_ | _6522_ /*28608*/;
  assign _6524_ = inv_30[7] ^ r_29[9] /*28606*/;
  assign sum_30[7] = _6524_ ^ _6523_ /*28605*/;
  assign _6525_ = _6524_ & _6523_ /*28604*/;
  assign _6526_ = inv_30[7] & r_29[9] /*28603*/;
  assign _6527_ = _6525_ | _6526_ /*28602*/;
  assign _6528_ = inv_30[8] ^ r_29[10] /*28600*/;
  assign sum_30[8] = _6528_ ^ _6527_ /*28599*/;
  assign _6529_ = _6528_ & _6527_ /*28598*/;
  assign _6530_ = inv_30[8] & r_29[10] /*28597*/;
  assign _6531_ = _6529_ | _6530_ /*28596*/;
  assign _6532_ = inv_30[9] ^ r_29[11] /*28594*/;
  assign sum_30[9] = _6532_ ^ _6531_ /*28593*/;
  assign _6533_ = _6532_ & _6531_ /*28592*/;
  assign _6534_ = inv_30[9] & r_29[11] /*28591*/;
  assign _6535_ = _6533_ | _6534_ /*28590*/;
  assign _6536_ = inv_30[10] ^ r_29[12] /*28588*/;
  assign sum_30[10] = _6536_ ^ _6535_ /*28587*/;
  assign _6537_ = _6536_ & _6535_ /*28586*/;
  assign _6538_ = inv_30[10] & r_29[12] /*28585*/;
  assign _6539_ = _6537_ | _6538_ /*28584*/;
  assign _6540_ = inv_30[11] ^ r_29[13] /*28582*/;
  assign sum_30[11] = _6540_ ^ _6539_ /*28581*/;
  assign _6541_ = _6540_ & _6539_ /*28580*/;
  assign _6542_ = inv_30[11] & r_29[13] /*28579*/;
  assign _6543_ = _6541_ | _6542_ /*28578*/;
  assign _6544_ = inv_30[12] ^ r_29[14] /*28576*/;
  assign sum_30[12] = _6544_ ^ _6543_ /*28575*/;
  assign _6545_ = _6544_ & _6543_ /*28574*/;
  assign _6546_ = inv_30[12] & r_29[14] /*28573*/;
  assign _6547_ = _6545_ | _6546_ /*28572*/;
  assign _6548_ = inv_30[13] ^ r_29[15] /*28570*/;
  assign sum_30[13] = _6548_ ^ _6547_ /*28569*/;
  assign _6549_ = _6548_ & _6547_ /*28568*/;
  assign _6550_ = inv_30[13] & r_29[15] /*28567*/;
  assign _6551_ = _6549_ | _6550_ /*28566*/;
  assign _6552_ = inv_30[14] ^ r_29[16] /*28564*/;
  assign sum_30[14] = _6552_ ^ _6551_ /*28563*/;
  assign _6553_ = _6552_ & _6551_ /*28562*/;
  assign _6554_ = inv_30[14] & r_29[16] /*28561*/;
  assign _6555_ = _6553_ | _6554_ /*28560*/;
  assign _6556_ = inv_30[15] ^ r_29[17] /*28558*/;
  assign sum_30[15] = _6556_ ^ _6555_ /*28557*/;
  assign _6557_ = _6556_ & _6555_ /*28556*/;
  assign _6558_ = inv_30[15] & r_29[17] /*28555*/;
  assign _6559_ = _6557_ | _6558_ /*28554*/;
  assign _6560_ = inv_30[16] ^ r_29[18] /*28552*/;
  assign sum_30[16] = _6560_ ^ _6559_ /*28551*/;
  assign _6561_ = _6560_ & _6559_ /*28550*/;
  assign _6562_ = inv_30[16] & r_29[18] /*28549*/;
  assign _6563_ = _6561_ | _6562_ /*28548*/;
  assign _6564_ = inv_30[17] ^ r_29[19] /*28546*/;
  assign sum_30[17] = _6564_ ^ _6563_ /*28545*/;
  assign _6565_ = _6564_ & _6563_ /*28544*/;
  assign _6566_ = inv_30[17] & r_29[19] /*28543*/;
  assign _6567_ = _6565_ | _6566_ /*28542*/;
  assign _6568_ = inv_30[18] ^ r_29[20] /*28540*/;
  assign sum_30[18] = _6568_ ^ _6567_ /*28539*/;
  assign _6569_ = _6568_ & _6567_ /*28538*/;
  assign _6570_ = inv_30[18] & r_29[20] /*28537*/;
  assign _6571_ = _6569_ | _6570_ /*28536*/;
  assign _6572_ = inv_30[19] ^ r_29[21] /*28534*/;
  assign sum_30[19] = _6572_ ^ _6571_ /*28533*/;
  assign _6573_ = _6572_ & _6571_ /*28532*/;
  assign _6574_ = inv_30[19] & r_29[21] /*28531*/;
  assign _6575_ = _6573_ | _6574_ /*28530*/;
  assign _6576_ = inv_30[20] ^ r_29[22] /*28528*/;
  assign sum_30[20] = _6576_ ^ _6575_ /*28527*/;
  assign _6577_ = _6576_ & _6575_ /*28526*/;
  assign _6578_ = inv_30[20] & r_29[22] /*28525*/;
  assign _6579_ = _6577_ | _6578_ /*28524*/;
  assign _6580_ = inv_30[21] ^ r_29[23] /*28522*/;
  assign sum_30[21] = _6580_ ^ _6579_ /*28521*/;
  assign _6581_ = _6580_ & _6579_ /*28520*/;
  assign _6582_ = inv_30[21] & r_29[23] /*28519*/;
  assign _6583_ = _6581_ | _6582_ /*28518*/;
  assign _6584_ = inv_30[22] ^ r_29[24] /*28516*/;
  assign sum_30[22] = _6584_ ^ _6583_ /*28515*/;
  assign _6585_ = _6584_ & _6583_ /*28514*/;
  assign _6586_ = inv_30[22] & r_29[24] /*28513*/;
  assign _6587_ = _6585_ | _6586_ /*28512*/;
  assign _6588_ = inv_30[23] ^ r_29[25] /*28510*/;
  assign sum_30[23] = _6588_ ^ _6587_ /*28509*/;
  assign _6589_ = _6588_ & _6587_ /*28508*/;
  assign _6590_ = inv_30[23] & r_29[25] /*28507*/;
  assign _6591_ = _6589_ | _6590_ /*28506*/;
  assign _6592_ = inv_30[24] ^ r_29[26] /*28504*/;
  assign sum_30[24] = _6592_ ^ _6591_ /*28503*/;
  assign _6593_ = _6592_ & _6591_ /*28502*/;
  assign _6594_ = inv_30[24] & r_29[26] /*28501*/;
  assign _6595_ = _6593_ | _6594_ /*28500*/;
  assign _6596_ = inv_30[25] ^ r_29[27] /*28498*/;
  assign sum_30[25] = _6596_ ^ _6595_ /*28497*/;
  assign _6597_ = _6596_ & _6595_ /*28496*/;
  assign _6598_ = inv_30[25] & r_29[27] /*28495*/;
  assign _6599_ = _6597_ | _6598_ /*28494*/;
  assign _6600_ = inv_30[26] ^ r_29[28] /*28492*/;
  assign sum_30[26] = _6600_ ^ _6599_ /*28491*/;
  assign _6601_ = _6600_ & _6599_ /*28490*/;
  assign _6602_ = inv_30[26] & r_29[28] /*28489*/;
  assign _6603_ = _6601_ | _6602_ /*28488*/;
  assign _6604_ = inv_30[27] ^ r_29[29] /*28486*/;
  assign sum_30[27] = _6604_ ^ _6603_ /*28485*/;
  assign _6605_ = _6604_ & _6603_ /*28484*/;
  assign _6606_ = inv_30[27] & r_29[29] /*28483*/;
  assign _6607_ = _6605_ | _6606_ /*28482*/;
  assign _6608_ = inv_30[28] ^ r_29[30] /*28480*/;
  assign sum_30[28] = _6608_ ^ _6607_ /*28479*/;
  assign _6609_ = _6608_ & _6607_ /*28478*/;
  assign _6610_ = inv_30[28] & r_29[30] /*28477*/;
  assign _6611_ = _6609_ | _6610_ /*28476*/;
  assign _6612_ = inv_30[29] ^ r_29[31] /*28474*/;
  assign sum_30[29] = _6612_ ^ _6611_ /*28473*/;
  assign _6613_ = _6612_ & _6611_ /*28472*/;
  assign _6614_ = inv_30[29] & r_29[31] /*28471*/;
  assign _6615_ = _6613_ | _6614_ /*28470*/;
  assign _6616_ = inv_30[30] ^ r_29[32] /*28468*/;
  assign sum_30[30] = _6616_ ^ _6615_ /*28467*/;
  assign _6617_ = _6616_ & _6615_ /*28466*/;
  assign _6618_ = inv_30[30] & r_29[32] /*28465*/;
  assign _6619_ = _6617_ | _6618_ /*28464*/;
  assign _6620_ = inv_30[31] ^ r_29[33] /*28462*/;
  assign sum_30[31] = _6620_ ^ _6619_ /*28461*/;
  assign _6621_ = _6620_ & _6619_ /*28460*/;
  assign _6622_ = inv_30[31] & r_29[33] /*28459*/;
  assign _6623_ = _6621_ | _6622_ /*28458*/;
  assign q[2] = ~sum_30[31] /*28485*/;
  assign m_30[0] = r_29[2] /*28484*/;
  assign m_30[1] = r_29[3] /*28483*/;
  assign m_30[2] = r_29[4] /*28482*/;
  assign m_30[3] = r_29[5] /*28481*/;
  assign m_30[4] = r_29[6] /*28480*/;
  assign m_30[5] = r_29[7] /*28479*/;
  assign m_30[6] = r_29[8] /*28478*/;
  assign m_30[7] = r_29[9] /*28477*/;
  assign m_30[8] = r_29[10] /*28476*/;
  assign m_30[9] = r_29[11] /*28475*/;
  assign m_30[10] = r_29[12] /*28474*/;
  assign m_30[11] = r_29[13] /*28473*/;
  assign m_30[12] = r_29[14] /*28472*/;
  assign m_30[13] = r_29[15] /*28471*/;
  assign m_30[14] = r_29[16] /*28470*/;
  assign m_30[15] = r_29[17] /*28469*/;
  assign m_30[16] = r_29[18] /*28468*/;
  assign m_30[17] = r_29[19] /*28467*/;
  assign m_30[18] = r_29[20] /*28466*/;
  assign m_30[19] = r_29[21] /*28465*/;
  assign m_30[20] = r_29[22] /*28464*/;
  assign m_30[21] = r_29[23] /*28463*/;
  assign m_30[22] = r_29[24] /*28462*/;
  assign m_30[23] = r_29[25] /*28461*/;
  assign m_30[24] = r_29[26] /*28460*/;
  assign m_30[25] = r_29[27] /*28459*/;
  assign m_30[26] = r_29[28] /*28458*/;
  assign m_30[27] = r_29[29] /*28457*/;
  assign m_30[28] = r_29[30] /*28456*/;
  assign m_30[29] = r_29[31] /*28455*/;
  assign m_30[30] = r_29[32] /*28454*/;
  assign m_30[31] = r_29[33] /*28453*/;
  assign _6624_ = ~q[2] /*28451*/;
  assign _6625_ = sum_30[0] & q[2] /*28450*/;
  assign _6626_ = m_30[0] & _6624_ /*28449*/;
  assign r_30[2] = _6626_ | _6625_ /*28448*/;
  assign _6627_ = ~q[2] /*28447*/;
  assign _6628_ = sum_30[1] & q[2] /*28446*/;
  assign _6629_ = m_30[1] & _6627_ /*28445*/;
  assign r_30[3] = _6629_ | _6628_ /*28444*/;
  assign _6630_ = ~q[2] /*28443*/;
  assign _6631_ = sum_30[2] & q[2] /*28442*/;
  assign _6632_ = m_30[2] & _6630_ /*28441*/;
  assign r_30[4] = _6632_ | _6631_ /*28440*/;
  assign _6633_ = ~q[2] /*28439*/;
  assign _6634_ = sum_30[3] & q[2] /*28438*/;
  assign _6635_ = m_30[3] & _6633_ /*28437*/;
  assign r_30[5] = _6635_ | _6634_ /*28436*/;
  assign _6636_ = ~q[2] /*28435*/;
  assign _6637_ = sum_30[4] & q[2] /*28434*/;
  assign _6638_ = m_30[4] & _6636_ /*28433*/;
  assign r_30[6] = _6638_ | _6637_ /*28432*/;
  assign _6639_ = ~q[2] /*28431*/;
  assign _6640_ = sum_30[5] & q[2] /*28430*/;
  assign _6641_ = m_30[5] & _6639_ /*28429*/;
  assign r_30[7] = _6641_ | _6640_ /*28428*/;
  assign _6642_ = ~q[2] /*28427*/;
  assign _6643_ = sum_30[6] & q[2] /*28426*/;
  assign _6644_ = m_30[6] & _6642_ /*28425*/;
  assign r_30[8] = _6644_ | _6643_ /*28424*/;
  assign _6645_ = ~q[2] /*28423*/;
  assign _6646_ = sum_30[7] & q[2] /*28422*/;
  assign _6647_ = m_30[7] & _6645_ /*28421*/;
  assign r_30[9] = _6647_ | _6646_ /*28420*/;
  assign _6648_ = ~q[2] /*28419*/;
  assign _6649_ = sum_30[8] & q[2] /*28418*/;
  assign _6650_ = m_30[8] & _6648_ /*28417*/;
  assign r_30[10] = _6650_ | _6649_ /*28416*/;
  assign _6651_ = ~q[2] /*28415*/;
  assign _6652_ = sum_30[9] & q[2] /*28414*/;
  assign _6653_ = m_30[9] & _6651_ /*28413*/;
  assign r_30[11] = _6653_ | _6652_ /*28412*/;
  assign _6654_ = ~q[2] /*28411*/;
  assign _6655_ = sum_30[10] & q[2] /*28410*/;
  assign _6656_ = m_30[10] & _6654_ /*28409*/;
  assign r_30[12] = _6656_ | _6655_ /*28408*/;
  assign _6657_ = ~q[2] /*28407*/;
  assign _6658_ = sum_30[11] & q[2] /*28406*/;
  assign _6659_ = m_30[11] & _6657_ /*28405*/;
  assign r_30[13] = _6659_ | _6658_ /*28404*/;
  assign _6660_ = ~q[2] /*28403*/;
  assign _6661_ = sum_30[12] & q[2] /*28402*/;
  assign _6662_ = m_30[12] & _6660_ /*28401*/;
  assign r_30[14] = _6662_ | _6661_ /*28400*/;
  assign _6663_ = ~q[2] /*28399*/;
  assign _6664_ = sum_30[13] & q[2] /*28398*/;
  assign _6665_ = m_30[13] & _6663_ /*28397*/;
  assign r_30[15] = _6665_ | _6664_ /*28396*/;
  assign _6666_ = ~q[2] /*28395*/;
  assign _6667_ = sum_30[14] & q[2] /*28394*/;
  assign _6668_ = m_30[14] & _6666_ /*28393*/;
  assign r_30[16] = _6668_ | _6667_ /*28392*/;
  assign _6669_ = ~q[2] /*28391*/;
  assign _6670_ = sum_30[15] & q[2] /*28390*/;
  assign _6671_ = m_30[15] & _6669_ /*28389*/;
  assign r_30[17] = _6671_ | _6670_ /*28388*/;
  assign _6672_ = ~q[2] /*28387*/;
  assign _6673_ = sum_30[16] & q[2] /*28386*/;
  assign _6674_ = m_30[16] & _6672_ /*28385*/;
  assign r_30[18] = _6674_ | _6673_ /*28384*/;
  assign _6675_ = ~q[2] /*28383*/;
  assign _6676_ = sum_30[17] & q[2] /*28382*/;
  assign _6677_ = m_30[17] & _6675_ /*28381*/;
  assign r_30[19] = _6677_ | _6676_ /*28380*/;
  assign _6678_ = ~q[2] /*28379*/;
  assign _6679_ = sum_30[18] & q[2] /*28378*/;
  assign _6680_ = m_30[18] & _6678_ /*28377*/;
  assign r_30[20] = _6680_ | _6679_ /*28376*/;
  assign _6681_ = ~q[2] /*28375*/;
  assign _6682_ = sum_30[19] & q[2] /*28374*/;
  assign _6683_ = m_30[19] & _6681_ /*28373*/;
  assign r_30[21] = _6683_ | _6682_ /*28372*/;
  assign _6684_ = ~q[2] /*28371*/;
  assign _6685_ = sum_30[20] & q[2] /*28370*/;
  assign _6686_ = m_30[20] & _6684_ /*28369*/;
  assign r_30[22] = _6686_ | _6685_ /*28368*/;
  assign _6687_ = ~q[2] /*28367*/;
  assign _6688_ = sum_30[21] & q[2] /*28366*/;
  assign _6689_ = m_30[21] & _6687_ /*28365*/;
  assign r_30[23] = _6689_ | _6688_ /*28364*/;
  assign _6690_ = ~q[2] /*28363*/;
  assign _6691_ = sum_30[22] & q[2] /*28362*/;
  assign _6692_ = m_30[22] & _6690_ /*28361*/;
  assign r_30[24] = _6692_ | _6691_ /*28360*/;
  assign _6693_ = ~q[2] /*28359*/;
  assign _6694_ = sum_30[23] & q[2] /*28358*/;
  assign _6695_ = m_30[23] & _6693_ /*28357*/;
  assign r_30[25] = _6695_ | _6694_ /*28356*/;
  assign _6696_ = ~q[2] /*28355*/;
  assign _6697_ = sum_30[24] & q[2] /*28354*/;
  assign _6698_ = m_30[24] & _6696_ /*28353*/;
  assign r_30[26] = _6698_ | _6697_ /*28352*/;
  assign _6699_ = ~q[2] /*28351*/;
  assign _6700_ = sum_30[25] & q[2] /*28350*/;
  assign _6701_ = m_30[25] & _6699_ /*28349*/;
  assign r_30[27] = _6701_ | _6700_ /*28348*/;
  assign _6702_ = ~q[2] /*28347*/;
  assign _6703_ = sum_30[26] & q[2] /*28346*/;
  assign _6704_ = m_30[26] & _6702_ /*28345*/;
  assign r_30[28] = _6704_ | _6703_ /*28344*/;
  assign _6705_ = ~q[2] /*28343*/;
  assign _6706_ = sum_30[27] & q[2] /*28342*/;
  assign _6707_ = m_30[27] & _6705_ /*28341*/;
  assign r_30[29] = _6707_ | _6706_ /*28340*/;
  assign _6708_ = ~q[2] /*28339*/;
  assign _6709_ = sum_30[28] & q[2] /*28338*/;
  assign _6710_ = m_30[28] & _6708_ /*28337*/;
  assign r_30[30] = _6710_ | _6709_ /*28336*/;
  assign _6711_ = ~q[2] /*28335*/;
  assign _6712_ = sum_30[29] & q[2] /*28334*/;
  assign _6713_ = m_30[29] & _6711_ /*28333*/;
  assign r_30[31] = _6713_ | _6712_ /*28332*/;
  assign _6714_ = ~q[2] /*28331*/;
  assign _6715_ = sum_30[30] & q[2] /*28330*/;
  assign _6716_ = m_30[30] & _6714_ /*28329*/;
  assign r_30[32] = _6716_ | _6715_ /*28328*/;
  assign _6717_ = ~q[2] /*28327*/;
  assign _6718_ = sum_30[31] & q[2] /*28326*/;
  assign _6719_ = m_30[31] & _6717_ /*28325*/;
  assign r_30[33] = _6719_ | _6718_ /*28324*/;
assign r_30[0]= r_29[0] /*28323*/;
assign r_30[1]= r_29[1] /*28322*/;
  assign inv_31[0] = ~div[0] /*28232*/;
  assign inv_31[1] = ~div[1] /*28231*/;
  assign inv_31[2] = ~div[2] /*28230*/;
  assign inv_31[3] = ~div[3] /*28229*/;
  assign inv_31[4] = ~div[4] /*28228*/;
  assign inv_31[5] = ~div[5] /*28227*/;
  assign inv_31[6] = ~div[6] /*28226*/;
  assign inv_31[7] = ~div[7] /*28225*/;
  assign inv_31[8] = ~div[8] /*28224*/;
  assign inv_31[9] = ~div[9] /*28223*/;
  assign inv_31[10] = ~div[10] /*28222*/;
  assign inv_31[11] = ~div[11] /*28221*/;
  assign inv_31[12] = ~div[12] /*28220*/;
  assign inv_31[13] = ~div[13] /*28219*/;
  assign inv_31[14] = ~div[14] /*28218*/;
  assign inv_31[15] = ~div[15] /*28217*/;
  assign inv_31[16] = ~div[16] /*28216*/;
  assign inv_31[17] = ~div[17] /*28215*/;
  assign inv_31[18] = ~div[18] /*28214*/;
  assign inv_31[19] = ~div[19] /*28213*/;
  assign inv_31[20] = ~div[20] /*28212*/;
  assign inv_31[21] = ~div[21] /*28211*/;
  assign inv_31[22] = ~div[22] /*28210*/;
  assign inv_31[23] = ~div[23] /*28209*/;
  assign inv_31[24] = ~div[24] /*28208*/;
  assign inv_31[25] = ~div[25] /*28207*/;
  assign inv_31[26] = ~div[26] /*28206*/;
  assign inv_31[27] = ~div[27] /*28205*/;
  assign inv_31[28] = ~div[28] /*28204*/;
  assign inv_31[29] = ~div[29] /*28203*/;
  assign inv_31[30] = ~div[30] /*28202*/;
assign inv_31[31] = oneWire /*28201*/;
  assign _6720_ = inv_31[0] ^ r_30[1] /*28199*/;
  assign sum_31[0] = _6720_ ^ oneWire /*28198*/;
  assign _6721_ = _6720_ & oneWire /*28197*/;
  assign _6722_ = inv_31[0] & r_30[1] /*28196*/;
  assign _6723_ = _6721_ | _6722_ /*28195*/;
  assign _6724_ = inv_31[1] ^ r_30[2] /*28194*/;
  assign sum_31[1] = _6724_ ^ _6723_ /*28193*/;
  assign _6725_ = _6724_ & _6723_ /*28192*/;
  assign _6726_ = inv_31[1] & r_30[2] /*28191*/;
  assign _6727_ = _6725_ | _6726_ /*28190*/;
  assign _6728_ = inv_31[2] ^ r_30[3] /*28188*/;
  assign sum_31[2] = _6728_ ^ _6727_ /*28187*/;
  assign _6729_ = _6728_ & _6727_ /*28186*/;
  assign _6730_ = inv_31[2] & r_30[3] /*28185*/;
  assign _6731_ = _6729_ | _6730_ /*28184*/;
  assign _6732_ = inv_31[3] ^ r_30[4] /*28182*/;
  assign sum_31[3] = _6732_ ^ _6731_ /*28181*/;
  assign _6733_ = _6732_ & _6731_ /*28180*/;
  assign _6734_ = inv_31[3] & r_30[4] /*28179*/;
  assign _6735_ = _6733_ | _6734_ /*28178*/;
  assign _6736_ = inv_31[4] ^ r_30[5] /*28176*/;
  assign sum_31[4] = _6736_ ^ _6735_ /*28175*/;
  assign _6737_ = _6736_ & _6735_ /*28174*/;
  assign _6738_ = inv_31[4] & r_30[5] /*28173*/;
  assign _6739_ = _6737_ | _6738_ /*28172*/;
  assign _6740_ = inv_31[5] ^ r_30[6] /*28170*/;
  assign sum_31[5] = _6740_ ^ _6739_ /*28169*/;
  assign _6741_ = _6740_ & _6739_ /*28168*/;
  assign _6742_ = inv_31[5] & r_30[6] /*28167*/;
  assign _6743_ = _6741_ | _6742_ /*28166*/;
  assign _6744_ = inv_31[6] ^ r_30[7] /*28164*/;
  assign sum_31[6] = _6744_ ^ _6743_ /*28163*/;
  assign _6745_ = _6744_ & _6743_ /*28162*/;
  assign _6746_ = inv_31[6] & r_30[7] /*28161*/;
  assign _6747_ = _6745_ | _6746_ /*28160*/;
  assign _6748_ = inv_31[7] ^ r_30[8] /*28158*/;
  assign sum_31[7] = _6748_ ^ _6747_ /*28157*/;
  assign _6749_ = _6748_ & _6747_ /*28156*/;
  assign _6750_ = inv_31[7] & r_30[8] /*28155*/;
  assign _6751_ = _6749_ | _6750_ /*28154*/;
  assign _6752_ = inv_31[8] ^ r_30[9] /*28152*/;
  assign sum_31[8] = _6752_ ^ _6751_ /*28151*/;
  assign _6753_ = _6752_ & _6751_ /*28150*/;
  assign _6754_ = inv_31[8] & r_30[9] /*28149*/;
  assign _6755_ = _6753_ | _6754_ /*28148*/;
  assign _6756_ = inv_31[9] ^ r_30[10] /*28146*/;
  assign sum_31[9] = _6756_ ^ _6755_ /*28145*/;
  assign _6757_ = _6756_ & _6755_ /*28144*/;
  assign _6758_ = inv_31[9] & r_30[10] /*28143*/;
  assign _6759_ = _6757_ | _6758_ /*28142*/;
  assign _6760_ = inv_31[10] ^ r_30[11] /*28140*/;
  assign sum_31[10] = _6760_ ^ _6759_ /*28139*/;
  assign _6761_ = _6760_ & _6759_ /*28138*/;
  assign _6762_ = inv_31[10] & r_30[11] /*28137*/;
  assign _6763_ = _6761_ | _6762_ /*28136*/;
  assign _6764_ = inv_31[11] ^ r_30[12] /*28134*/;
  assign sum_31[11] = _6764_ ^ _6763_ /*28133*/;
  assign _6765_ = _6764_ & _6763_ /*28132*/;
  assign _6766_ = inv_31[11] & r_30[12] /*28131*/;
  assign _6767_ = _6765_ | _6766_ /*28130*/;
  assign _6768_ = inv_31[12] ^ r_30[13] /*28128*/;
  assign sum_31[12] = _6768_ ^ _6767_ /*28127*/;
  assign _6769_ = _6768_ & _6767_ /*28126*/;
  assign _6770_ = inv_31[12] & r_30[13] /*28125*/;
  assign _6771_ = _6769_ | _6770_ /*28124*/;
  assign _6772_ = inv_31[13] ^ r_30[14] /*28122*/;
  assign sum_31[13] = _6772_ ^ _6771_ /*28121*/;
  assign _6773_ = _6772_ & _6771_ /*28120*/;
  assign _6774_ = inv_31[13] & r_30[14] /*28119*/;
  assign _6775_ = _6773_ | _6774_ /*28118*/;
  assign _6776_ = inv_31[14] ^ r_30[15] /*28116*/;
  assign sum_31[14] = _6776_ ^ _6775_ /*28115*/;
  assign _6777_ = _6776_ & _6775_ /*28114*/;
  assign _6778_ = inv_31[14] & r_30[15] /*28113*/;
  assign _6779_ = _6777_ | _6778_ /*28112*/;
  assign _6780_ = inv_31[15] ^ r_30[16] /*28110*/;
  assign sum_31[15] = _6780_ ^ _6779_ /*28109*/;
  assign _6781_ = _6780_ & _6779_ /*28108*/;
  assign _6782_ = inv_31[15] & r_30[16] /*28107*/;
  assign _6783_ = _6781_ | _6782_ /*28106*/;
  assign _6784_ = inv_31[16] ^ r_30[17] /*28104*/;
  assign sum_31[16] = _6784_ ^ _6783_ /*28103*/;
  assign _6785_ = _6784_ & _6783_ /*28102*/;
  assign _6786_ = inv_31[16] & r_30[17] /*28101*/;
  assign _6787_ = _6785_ | _6786_ /*28100*/;
  assign _6788_ = inv_31[17] ^ r_30[18] /*28098*/;
  assign sum_31[17] = _6788_ ^ _6787_ /*28097*/;
  assign _6789_ = _6788_ & _6787_ /*28096*/;
  assign _6790_ = inv_31[17] & r_30[18] /*28095*/;
  assign _6791_ = _6789_ | _6790_ /*28094*/;
  assign _6792_ = inv_31[18] ^ r_30[19] /*28092*/;
  assign sum_31[18] = _6792_ ^ _6791_ /*28091*/;
  assign _6793_ = _6792_ & _6791_ /*28090*/;
  assign _6794_ = inv_31[18] & r_30[19] /*28089*/;
  assign _6795_ = _6793_ | _6794_ /*28088*/;
  assign _6796_ = inv_31[19] ^ r_30[20] /*28086*/;
  assign sum_31[19] = _6796_ ^ _6795_ /*28085*/;
  assign _6797_ = _6796_ & _6795_ /*28084*/;
  assign _6798_ = inv_31[19] & r_30[20] /*28083*/;
  assign _6799_ = _6797_ | _6798_ /*28082*/;
  assign _6800_ = inv_31[20] ^ r_30[21] /*28080*/;
  assign sum_31[20] = _6800_ ^ _6799_ /*28079*/;
  assign _6801_ = _6800_ & _6799_ /*28078*/;
  assign _6802_ = inv_31[20] & r_30[21] /*28077*/;
  assign _6803_ = _6801_ | _6802_ /*28076*/;
  assign _6804_ = inv_31[21] ^ r_30[22] /*28074*/;
  assign sum_31[21] = _6804_ ^ _6803_ /*28073*/;
  assign _6805_ = _6804_ & _6803_ /*28072*/;
  assign _6806_ = inv_31[21] & r_30[22] /*28071*/;
  assign _6807_ = _6805_ | _6806_ /*28070*/;
  assign _6808_ = inv_31[22] ^ r_30[23] /*28068*/;
  assign sum_31[22] = _6808_ ^ _6807_ /*28067*/;
  assign _6809_ = _6808_ & _6807_ /*28066*/;
  assign _6810_ = inv_31[22] & r_30[23] /*28065*/;
  assign _6811_ = _6809_ | _6810_ /*28064*/;
  assign _6812_ = inv_31[23] ^ r_30[24] /*28062*/;
  assign sum_31[23] = _6812_ ^ _6811_ /*28061*/;
  assign _6813_ = _6812_ & _6811_ /*28060*/;
  assign _6814_ = inv_31[23] & r_30[24] /*28059*/;
  assign _6815_ = _6813_ | _6814_ /*28058*/;
  assign _6816_ = inv_31[24] ^ r_30[25] /*28056*/;
  assign sum_31[24] = _6816_ ^ _6815_ /*28055*/;
  assign _6817_ = _6816_ & _6815_ /*28054*/;
  assign _6818_ = inv_31[24] & r_30[25] /*28053*/;
  assign _6819_ = _6817_ | _6818_ /*28052*/;
  assign _6820_ = inv_31[25] ^ r_30[26] /*28050*/;
  assign sum_31[25] = _6820_ ^ _6819_ /*28049*/;
  assign _6821_ = _6820_ & _6819_ /*28048*/;
  assign _6822_ = inv_31[25] & r_30[26] /*28047*/;
  assign _6823_ = _6821_ | _6822_ /*28046*/;
  assign _6824_ = inv_31[26] ^ r_30[27] /*28044*/;
  assign sum_31[26] = _6824_ ^ _6823_ /*28043*/;
  assign _6825_ = _6824_ & _6823_ /*28042*/;
  assign _6826_ = inv_31[26] & r_30[27] /*28041*/;
  assign _6827_ = _6825_ | _6826_ /*28040*/;
  assign _6828_ = inv_31[27] ^ r_30[28] /*28038*/;
  assign sum_31[27] = _6828_ ^ _6827_ /*28037*/;
  assign _6829_ = _6828_ & _6827_ /*28036*/;
  assign _6830_ = inv_31[27] & r_30[28] /*28035*/;
  assign _6831_ = _6829_ | _6830_ /*28034*/;
  assign _6832_ = inv_31[28] ^ r_30[29] /*28032*/;
  assign sum_31[28] = _6832_ ^ _6831_ /*28031*/;
  assign _6833_ = _6832_ & _6831_ /*28030*/;
  assign _6834_ = inv_31[28] & r_30[29] /*28029*/;
  assign _6835_ = _6833_ | _6834_ /*28028*/;
  assign _6836_ = inv_31[29] ^ r_30[30] /*28026*/;
  assign sum_31[29] = _6836_ ^ _6835_ /*28025*/;
  assign _6837_ = _6836_ & _6835_ /*28024*/;
  assign _6838_ = inv_31[29] & r_30[30] /*28023*/;
  assign _6839_ = _6837_ | _6838_ /*28022*/;
  assign _6840_ = inv_31[30] ^ r_30[31] /*28020*/;
  assign sum_31[30] = _6840_ ^ _6839_ /*28019*/;
  assign _6841_ = _6840_ & _6839_ /*28018*/;
  assign _6842_ = inv_31[30] & r_30[31] /*28017*/;
  assign _6843_ = _6841_ | _6842_ /*28016*/;
  assign _6844_ = inv_31[31] ^ r_30[32] /*28014*/;
  assign sum_31[31] = _6844_ ^ _6843_ /*28013*/;
  assign _6845_ = _6844_ & _6843_ /*28012*/;
  assign _6846_ = inv_31[31] & r_30[32] /*28011*/;
  assign _6847_ = _6845_ | _6846_ /*28010*/;
  assign q[1] = ~sum_31[31] /*28037*/;
  assign m_31[0] = r_30[1] /*28036*/;
  assign m_31[1] = r_30[2] /*28035*/;
  assign m_31[2] = r_30[3] /*28034*/;
  assign m_31[3] = r_30[4] /*28033*/;
  assign m_31[4] = r_30[5] /*28032*/;
  assign m_31[5] = r_30[6] /*28031*/;
  assign m_31[6] = r_30[7] /*28030*/;
  assign m_31[7] = r_30[8] /*28029*/;
  assign m_31[8] = r_30[9] /*28028*/;
  assign m_31[9] = r_30[10] /*28027*/;
  assign m_31[10] = r_30[11] /*28026*/;
  assign m_31[11] = r_30[12] /*28025*/;
  assign m_31[12] = r_30[13] /*28024*/;
  assign m_31[13] = r_30[14] /*28023*/;
  assign m_31[14] = r_30[15] /*28022*/;
  assign m_31[15] = r_30[16] /*28021*/;
  assign m_31[16] = r_30[17] /*28020*/;
  assign m_31[17] = r_30[18] /*28019*/;
  assign m_31[18] = r_30[19] /*28018*/;
  assign m_31[19] = r_30[20] /*28017*/;
  assign m_31[20] = r_30[21] /*28016*/;
  assign m_31[21] = r_30[22] /*28015*/;
  assign m_31[22] = r_30[23] /*28014*/;
  assign m_31[23] = r_30[24] /*28013*/;
  assign m_31[24] = r_30[25] /*28012*/;
  assign m_31[25] = r_30[26] /*28011*/;
  assign m_31[26] = r_30[27] /*28010*/;
  assign m_31[27] = r_30[28] /*28009*/;
  assign m_31[28] = r_30[29] /*28008*/;
  assign m_31[29] = r_30[30] /*28007*/;
  assign m_31[30] = r_30[31] /*28006*/;
  assign m_31[31] = r_30[32] /*28005*/;
  assign _6848_ = ~q[1] /*28003*/;
  assign _6849_ = sum_31[0] & q[1] /*28002*/;
  assign _6850_ = m_31[0] & _6848_ /*28001*/;
  assign r_31[1] = _6850_ | _6849_ /*28000*/;
  assign _6851_ = ~q[1] /*27999*/;
  assign _6852_ = sum_31[1] & q[1] /*27998*/;
  assign _6853_ = m_31[1] & _6851_ /*27997*/;
  assign r_31[2] = _6853_ | _6852_ /*27996*/;
  assign _6854_ = ~q[1] /*27995*/;
  assign _6855_ = sum_31[2] & q[1] /*27994*/;
  assign _6856_ = m_31[2] & _6854_ /*27993*/;
  assign r_31[3] = _6856_ | _6855_ /*27992*/;
  assign _6857_ = ~q[1] /*27991*/;
  assign _6858_ = sum_31[3] & q[1] /*27990*/;
  assign _6859_ = m_31[3] & _6857_ /*27989*/;
  assign r_31[4] = _6859_ | _6858_ /*27988*/;
  assign _6860_ = ~q[1] /*27987*/;
  assign _6861_ = sum_31[4] & q[1] /*27986*/;
  assign _6862_ = m_31[4] & _6860_ /*27985*/;
  assign r_31[5] = _6862_ | _6861_ /*27984*/;
  assign _6863_ = ~q[1] /*27983*/;
  assign _6864_ = sum_31[5] & q[1] /*27982*/;
  assign _6865_ = m_31[5] & _6863_ /*27981*/;
  assign r_31[6] = _6865_ | _6864_ /*27980*/;
  assign _6866_ = ~q[1] /*27979*/;
  assign _6867_ = sum_31[6] & q[1] /*27978*/;
  assign _6868_ = m_31[6] & _6866_ /*27977*/;
  assign r_31[7] = _6868_ | _6867_ /*27976*/;
  assign _6869_ = ~q[1] /*27975*/;
  assign _6870_ = sum_31[7] & q[1] /*27974*/;
  assign _6871_ = m_31[7] & _6869_ /*27973*/;
  assign r_31[8] = _6871_ | _6870_ /*27972*/;
  assign _6872_ = ~q[1] /*27971*/;
  assign _6873_ = sum_31[8] & q[1] /*27970*/;
  assign _6874_ = m_31[8] & _6872_ /*27969*/;
  assign r_31[9] = _6874_ | _6873_ /*27968*/;
  assign _6875_ = ~q[1] /*27967*/;
  assign _6876_ = sum_31[9] & q[1] /*27966*/;
  assign _6877_ = m_31[9] & _6875_ /*27965*/;
  assign r_31[10] = _6877_ | _6876_ /*27964*/;
  assign _6878_ = ~q[1] /*27963*/;
  assign _6879_ = sum_31[10] & q[1] /*27962*/;
  assign _6880_ = m_31[10] & _6878_ /*27961*/;
  assign r_31[11] = _6880_ | _6879_ /*27960*/;
  assign _6881_ = ~q[1] /*27959*/;
  assign _6882_ = sum_31[11] & q[1] /*27958*/;
  assign _6883_ = m_31[11] & _6881_ /*27957*/;
  assign r_31[12] = _6883_ | _6882_ /*27956*/;
  assign _6884_ = ~q[1] /*27955*/;
  assign _6885_ = sum_31[12] & q[1] /*27954*/;
  assign _6886_ = m_31[12] & _6884_ /*27953*/;
  assign r_31[13] = _6886_ | _6885_ /*27952*/;
  assign _6887_ = ~q[1] /*27951*/;
  assign _6888_ = sum_31[13] & q[1] /*27950*/;
  assign _6889_ = m_31[13] & _6887_ /*27949*/;
  assign r_31[14] = _6889_ | _6888_ /*27948*/;
  assign _6890_ = ~q[1] /*27947*/;
  assign _6891_ = sum_31[14] & q[1] /*27946*/;
  assign _6892_ = m_31[14] & _6890_ /*27945*/;
  assign r_31[15] = _6892_ | _6891_ /*27944*/;
  assign _6893_ = ~q[1] /*27943*/;
  assign _6894_ = sum_31[15] & q[1] /*27942*/;
  assign _6895_ = m_31[15] & _6893_ /*27941*/;
  assign r_31[16] = _6895_ | _6894_ /*27940*/;
  assign _6896_ = ~q[1] /*27939*/;
  assign _6897_ = sum_31[16] & q[1] /*27938*/;
  assign _6898_ = m_31[16] & _6896_ /*27937*/;
  assign r_31[17] = _6898_ | _6897_ /*27936*/;
  assign _6899_ = ~q[1] /*27935*/;
  assign _6900_ = sum_31[17] & q[1] /*27934*/;
  assign _6901_ = m_31[17] & _6899_ /*27933*/;
  assign r_31[18] = _6901_ | _6900_ /*27932*/;
  assign _6902_ = ~q[1] /*27931*/;
  assign _6903_ = sum_31[18] & q[1] /*27930*/;
  assign _6904_ = m_31[18] & _6902_ /*27929*/;
  assign r_31[19] = _6904_ | _6903_ /*27928*/;
  assign _6905_ = ~q[1] /*27927*/;
  assign _6906_ = sum_31[19] & q[1] /*27926*/;
  assign _6907_ = m_31[19] & _6905_ /*27925*/;
  assign r_31[20] = _6907_ | _6906_ /*27924*/;
  assign _6908_ = ~q[1] /*27923*/;
  assign _6909_ = sum_31[20] & q[1] /*27922*/;
  assign _6910_ = m_31[20] & _6908_ /*27921*/;
  assign r_31[21] = _6910_ | _6909_ /*27920*/;
  assign _6911_ = ~q[1] /*27919*/;
  assign _6912_ = sum_31[21] & q[1] /*27918*/;
  assign _6913_ = m_31[21] & _6911_ /*27917*/;
  assign r_31[22] = _6913_ | _6912_ /*27916*/;
  assign _6914_ = ~q[1] /*27915*/;
  assign _6915_ = sum_31[22] & q[1] /*27914*/;
  assign _6916_ = m_31[22] & _6914_ /*27913*/;
  assign r_31[23] = _6916_ | _6915_ /*27912*/;
  assign _6917_ = ~q[1] /*27911*/;
  assign _6918_ = sum_31[23] & q[1] /*27910*/;
  assign _6919_ = m_31[23] & _6917_ /*27909*/;
  assign r_31[24] = _6919_ | _6918_ /*27908*/;
  assign _6920_ = ~q[1] /*27907*/;
  assign _6921_ = sum_31[24] & q[1] /*27906*/;
  assign _6922_ = m_31[24] & _6920_ /*27905*/;
  assign r_31[25] = _6922_ | _6921_ /*27904*/;
  assign _6923_ = ~q[1] /*27903*/;
  assign _6924_ = sum_31[25] & q[1] /*27902*/;
  assign _6925_ = m_31[25] & _6923_ /*27901*/;
  assign r_31[26] = _6925_ | _6924_ /*27900*/;
  assign _6926_ = ~q[1] /*27899*/;
  assign _6927_ = sum_31[26] & q[1] /*27898*/;
  assign _6928_ = m_31[26] & _6926_ /*27897*/;
  assign r_31[27] = _6928_ | _6927_ /*27896*/;
  assign _6929_ = ~q[1] /*27895*/;
  assign _6930_ = sum_31[27] & q[1] /*27894*/;
  assign _6931_ = m_31[27] & _6929_ /*27893*/;
  assign r_31[28] = _6931_ | _6930_ /*27892*/;
  assign _6932_ = ~q[1] /*27891*/;
  assign _6933_ = sum_31[28] & q[1] /*27890*/;
  assign _6934_ = m_31[28] & _6932_ /*27889*/;
  assign r_31[29] = _6934_ | _6933_ /*27888*/;
  assign _6935_ = ~q[1] /*27887*/;
  assign _6936_ = sum_31[29] & q[1] /*27886*/;
  assign _6937_ = m_31[29] & _6935_ /*27885*/;
  assign r_31[30] = _6937_ | _6936_ /*27884*/;
  assign _6938_ = ~q[1] /*27883*/;
  assign _6939_ = sum_31[30] & q[1] /*27882*/;
  assign _6940_ = m_31[30] & _6938_ /*27881*/;
  assign r_31[31] = _6940_ | _6939_ /*27880*/;
  assign _6941_ = ~q[1] /*27879*/;
  assign _6942_ = sum_31[31] & q[1] /*27878*/;
  assign _6943_ = m_31[31] & _6941_ /*27877*/;
  assign r_31[32] = _6943_ | _6942_ /*27876*/;
assign r_31[0]= r_30[0] /*27875*/;
  assign inv_32[0] = ~div[0] /*27784*/;
  assign inv_32[1] = ~div[1] /*27783*/;
  assign inv_32[2] = ~div[2] /*27782*/;
  assign inv_32[3] = ~div[3] /*27781*/;
  assign inv_32[4] = ~div[4] /*27780*/;
  assign inv_32[5] = ~div[5] /*27779*/;
  assign inv_32[6] = ~div[6] /*27778*/;
  assign inv_32[7] = ~div[7] /*27777*/;
  assign inv_32[8] = ~div[8] /*27776*/;
  assign inv_32[9] = ~div[9] /*27775*/;
  assign inv_32[10] = ~div[10] /*27774*/;
  assign inv_32[11] = ~div[11] /*27773*/;
  assign inv_32[12] = ~div[12] /*27772*/;
  assign inv_32[13] = ~div[13] /*27771*/;
  assign inv_32[14] = ~div[14] /*27770*/;
  assign inv_32[15] = ~div[15] /*27769*/;
  assign inv_32[16] = ~div[16] /*27768*/;
  assign inv_32[17] = ~div[17] /*27767*/;
  assign inv_32[18] = ~div[18] /*27766*/;
  assign inv_32[19] = ~div[19] /*27765*/;
  assign inv_32[20] = ~div[20] /*27764*/;
  assign inv_32[21] = ~div[21] /*27763*/;
  assign inv_32[22] = ~div[22] /*27762*/;
  assign inv_32[23] = ~div[23] /*27761*/;
  assign inv_32[24] = ~div[24] /*27760*/;
  assign inv_32[25] = ~div[25] /*27759*/;
  assign inv_32[26] = ~div[26] /*27758*/;
  assign inv_32[27] = ~div[27] /*27757*/;
  assign inv_32[28] = ~div[28] /*27756*/;
  assign inv_32[29] = ~div[29] /*27755*/;
  assign inv_32[30] = ~div[30] /*27754*/;
assign inv_32[31] = oneWire /*27753*/;
  assign _6944_ = inv_32[0] ^ r_31[0] /*27751*/;
  assign sum_32[0] = _6944_ ^ oneWire /*27750*/;
  assign _6945_ = _6944_ & oneWire /*27749*/;
  assign _6946_ = inv_32[0] & r_31[0] /*27748*/;
  assign _6947_ = _6945_ | _6946_ /*27747*/;
  assign _6948_ = inv_32[1] ^ r_31[1] /*27746*/;
  assign sum_32[1] = _6948_ ^ _6947_ /*27745*/;
  assign _6949_ = _6948_ & _6947_ /*27744*/;
  assign _6950_ = inv_32[1] & r_31[1] /*27743*/;
  assign _6951_ = _6949_ | _6950_ /*27742*/;
  assign _6952_ = inv_32[2] ^ r_31[2] /*27740*/;
  assign sum_32[2] = _6952_ ^ _6951_ /*27739*/;
  assign _6953_ = _6952_ & _6951_ /*27738*/;
  assign _6954_ = inv_32[2] & r_31[2] /*27737*/;
  assign _6955_ = _6953_ | _6954_ /*27736*/;
  assign _6956_ = inv_32[3] ^ r_31[3] /*27734*/;
  assign sum_32[3] = _6956_ ^ _6955_ /*27733*/;
  assign _6957_ = _6956_ & _6955_ /*27732*/;
  assign _6958_ = inv_32[3] & r_31[3] /*27731*/;
  assign _6959_ = _6957_ | _6958_ /*27730*/;
  assign _6960_ = inv_32[4] ^ r_31[4] /*27728*/;
  assign sum_32[4] = _6960_ ^ _6959_ /*27727*/;
  assign _6961_ = _6960_ & _6959_ /*27726*/;
  assign _6962_ = inv_32[4] & r_31[4] /*27725*/;
  assign _6963_ = _6961_ | _6962_ /*27724*/;
  assign _6964_ = inv_32[5] ^ r_31[5] /*27722*/;
  assign sum_32[5] = _6964_ ^ _6963_ /*27721*/;
  assign _6965_ = _6964_ & _6963_ /*27720*/;
  assign _6966_ = inv_32[5] & r_31[5] /*27719*/;
  assign _6967_ = _6965_ | _6966_ /*27718*/;
  assign _6968_ = inv_32[6] ^ r_31[6] /*27716*/;
  assign sum_32[6] = _6968_ ^ _6967_ /*27715*/;
  assign _6969_ = _6968_ & _6967_ /*27714*/;
  assign _6970_ = inv_32[6] & r_31[6] /*27713*/;
  assign _6971_ = _6969_ | _6970_ /*27712*/;
  assign _6972_ = inv_32[7] ^ r_31[7] /*27710*/;
  assign sum_32[7] = _6972_ ^ _6971_ /*27709*/;
  assign _6973_ = _6972_ & _6971_ /*27708*/;
  assign _6974_ = inv_32[7] & r_31[7] /*27707*/;
  assign _6975_ = _6973_ | _6974_ /*27706*/;
  assign _6976_ = inv_32[8] ^ r_31[8] /*27704*/;
  assign sum_32[8] = _6976_ ^ _6975_ /*27703*/;
  assign _6977_ = _6976_ & _6975_ /*27702*/;
  assign _6978_ = inv_32[8] & r_31[8] /*27701*/;
  assign _6979_ = _6977_ | _6978_ /*27700*/;
  assign _6980_ = inv_32[9] ^ r_31[9] /*27698*/;
  assign sum_32[9] = _6980_ ^ _6979_ /*27697*/;
  assign _6981_ = _6980_ & _6979_ /*27696*/;
  assign _6982_ = inv_32[9] & r_31[9] /*27695*/;
  assign _6983_ = _6981_ | _6982_ /*27694*/;
  assign _6984_ = inv_32[10] ^ r_31[10] /*27692*/;
  assign sum_32[10] = _6984_ ^ _6983_ /*27691*/;
  assign _6985_ = _6984_ & _6983_ /*27690*/;
  assign _6986_ = inv_32[10] & r_31[10] /*27689*/;
  assign _6987_ = _6985_ | _6986_ /*27688*/;
  assign _6988_ = inv_32[11] ^ r_31[11] /*27686*/;
  assign sum_32[11] = _6988_ ^ _6987_ /*27685*/;
  assign _6989_ = _6988_ & _6987_ /*27684*/;
  assign _6990_ = inv_32[11] & r_31[11] /*27683*/;
  assign _6991_ = _6989_ | _6990_ /*27682*/;
  assign _6992_ = inv_32[12] ^ r_31[12] /*27680*/;
  assign sum_32[12] = _6992_ ^ _6991_ /*27679*/;
  assign _6993_ = _6992_ & _6991_ /*27678*/;
  assign _6994_ = inv_32[12] & r_31[12] /*27677*/;
  assign _6995_ = _6993_ | _6994_ /*27676*/;
  assign _6996_ = inv_32[13] ^ r_31[13] /*27674*/;
  assign sum_32[13] = _6996_ ^ _6995_ /*27673*/;
  assign _6997_ = _6996_ & _6995_ /*27672*/;
  assign _6998_ = inv_32[13] & r_31[13] /*27671*/;
  assign _6999_ = _6997_ | _6998_ /*27670*/;
  assign _7000_ = inv_32[14] ^ r_31[14] /*27668*/;
  assign sum_32[14] = _7000_ ^ _6999_ /*27667*/;
  assign _7001_ = _7000_ & _6999_ /*27666*/;
  assign _7002_ = inv_32[14] & r_31[14] /*27665*/;
  assign _7003_ = _7001_ | _7002_ /*27664*/;
  assign _7004_ = inv_32[15] ^ r_31[15] /*27662*/;
  assign sum_32[15] = _7004_ ^ _7003_ /*27661*/;
  assign _7005_ = _7004_ & _7003_ /*27660*/;
  assign _7006_ = inv_32[15] & r_31[15] /*27659*/;
  assign _7007_ = _7005_ | _7006_ /*27658*/;
  assign _7008_ = inv_32[16] ^ r_31[16] /*27656*/;
  assign sum_32[16] = _7008_ ^ _7007_ /*27655*/;
  assign _7009_ = _7008_ & _7007_ /*27654*/;
  assign _7010_ = inv_32[16] & r_31[16] /*27653*/;
  assign _7011_ = _7009_ | _7010_ /*27652*/;
  assign _7012_ = inv_32[17] ^ r_31[17] /*27650*/;
  assign sum_32[17] = _7012_ ^ _7011_ /*27649*/;
  assign _7013_ = _7012_ & _7011_ /*27648*/;
  assign _7014_ = inv_32[17] & r_31[17] /*27647*/;
  assign _7015_ = _7013_ | _7014_ /*27646*/;
  assign _7016_ = inv_32[18] ^ r_31[18] /*27644*/;
  assign sum_32[18] = _7016_ ^ _7015_ /*27643*/;
  assign _7017_ = _7016_ & _7015_ /*27642*/;
  assign _7018_ = inv_32[18] & r_31[18] /*27641*/;
  assign _7019_ = _7017_ | _7018_ /*27640*/;
  assign _7020_ = inv_32[19] ^ r_31[19] /*27638*/;
  assign sum_32[19] = _7020_ ^ _7019_ /*27637*/;
  assign _7021_ = _7020_ & _7019_ /*27636*/;
  assign _7022_ = inv_32[19] & r_31[19] /*27635*/;
  assign _7023_ = _7021_ | _7022_ /*27634*/;
  assign _7024_ = inv_32[20] ^ r_31[20] /*27632*/;
  assign sum_32[20] = _7024_ ^ _7023_ /*27631*/;
  assign _7025_ = _7024_ & _7023_ /*27630*/;
  assign _7026_ = inv_32[20] & r_31[20] /*27629*/;
  assign _7027_ = _7025_ | _7026_ /*27628*/;
  assign _7028_ = inv_32[21] ^ r_31[21] /*27626*/;
  assign sum_32[21] = _7028_ ^ _7027_ /*27625*/;
  assign _7029_ = _7028_ & _7027_ /*27624*/;
  assign _7030_ = inv_32[21] & r_31[21] /*27623*/;
  assign _7031_ = _7029_ | _7030_ /*27622*/;
  assign _7032_ = inv_32[22] ^ r_31[22] /*27620*/;
  assign sum_32[22] = _7032_ ^ _7031_ /*27619*/;
  assign _7033_ = _7032_ & _7031_ /*27618*/;
  assign _7034_ = inv_32[22] & r_31[22] /*27617*/;
  assign _7035_ = _7033_ | _7034_ /*27616*/;
  assign _7036_ = inv_32[23] ^ r_31[23] /*27614*/;
  assign sum_32[23] = _7036_ ^ _7035_ /*27613*/;
  assign _7037_ = _7036_ & _7035_ /*27612*/;
  assign _7038_ = inv_32[23] & r_31[23] /*27611*/;
  assign _7039_ = _7037_ | _7038_ /*27610*/;
  assign _7040_ = inv_32[24] ^ r_31[24] /*27608*/;
  assign sum_32[24] = _7040_ ^ _7039_ /*27607*/;
  assign _7041_ = _7040_ & _7039_ /*27606*/;
  assign _7042_ = inv_32[24] & r_31[24] /*27605*/;
  assign _7043_ = _7041_ | _7042_ /*27604*/;
  assign _7044_ = inv_32[25] ^ r_31[25] /*27602*/;
  assign sum_32[25] = _7044_ ^ _7043_ /*27601*/;
  assign _7045_ = _7044_ & _7043_ /*27600*/;
  assign _7046_ = inv_32[25] & r_31[25] /*27599*/;
  assign _7047_ = _7045_ | _7046_ /*27598*/;
  assign _7048_ = inv_32[26] ^ r_31[26] /*27596*/;
  assign sum_32[26] = _7048_ ^ _7047_ /*27595*/;
  assign _7049_ = _7048_ & _7047_ /*27594*/;
  assign _7050_ = inv_32[26] & r_31[26] /*27593*/;
  assign _7051_ = _7049_ | _7050_ /*27592*/;
  assign _7052_ = inv_32[27] ^ r_31[27] /*27590*/;
  assign sum_32[27] = _7052_ ^ _7051_ /*27589*/;
  assign _7053_ = _7052_ & _7051_ /*27588*/;
  assign _7054_ = inv_32[27] & r_31[27] /*27587*/;
  assign _7055_ = _7053_ | _7054_ /*27586*/;
  assign _7056_ = inv_32[28] ^ r_31[28] /*27584*/;
  assign sum_32[28] = _7056_ ^ _7055_ /*27583*/;
  assign _7057_ = _7056_ & _7055_ /*27582*/;
  assign _7058_ = inv_32[28] & r_31[28] /*27581*/;
  assign _7059_ = _7057_ | _7058_ /*27580*/;
  assign _7060_ = inv_32[29] ^ r_31[29] /*27578*/;
  assign sum_32[29] = _7060_ ^ _7059_ /*27577*/;
  assign _7061_ = _7060_ & _7059_ /*27576*/;
  assign _7062_ = inv_32[29] & r_31[29] /*27575*/;
  assign _7063_ = _7061_ | _7062_ /*27574*/;
  assign _7064_ = inv_32[30] ^ r_31[30] /*27572*/;
  assign sum_32[30] = _7064_ ^ _7063_ /*27571*/;
  assign _7065_ = _7064_ & _7063_ /*27570*/;
  assign _7066_ = inv_32[30] & r_31[30] /*27569*/;
  assign _7067_ = _7065_ | _7066_ /*27568*/;
  assign _7068_ = inv_32[31] ^ r_31[31] /*27566*/;
  assign sum_32[31] = _7068_ ^ _7067_ /*27565*/;
  assign _7069_ = _7068_ & _7067_ /*27564*/;
  assign _7070_ = inv_32[31] & r_31[31] /*27563*/;
  assign _7071_ = _7069_ | _7070_ /*27562*/;
  assign q[0] = ~sum_32[31] /*27589*/;
  assign m_32[0] = r_31[0] /*27588*/;
  assign m_32[1] = r_31[1] /*27587*/;
  assign m_32[2] = r_31[2] /*27586*/;
  assign m_32[3] = r_31[3] /*27585*/;
  assign m_32[4] = r_31[4] /*27584*/;
  assign m_32[5] = r_31[5] /*27583*/;
  assign m_32[6] = r_31[6] /*27582*/;
  assign m_32[7] = r_31[7] /*27581*/;
  assign m_32[8] = r_31[8] /*27580*/;
  assign m_32[9] = r_31[9] /*27579*/;
  assign m_32[10] = r_31[10] /*27578*/;
  assign m_32[11] = r_31[11] /*27577*/;
  assign m_32[12] = r_31[12] /*27576*/;
  assign m_32[13] = r_31[13] /*27575*/;
  assign m_32[14] = r_31[14] /*27574*/;
  assign m_32[15] = r_31[15] /*27573*/;
  assign m_32[16] = r_31[16] /*27572*/;
  assign m_32[17] = r_31[17] /*27571*/;
  assign m_32[18] = r_31[18] /*27570*/;
  assign m_32[19] = r_31[19] /*27569*/;
  assign m_32[20] = r_31[20] /*27568*/;
  assign m_32[21] = r_31[21] /*27567*/;
  assign m_32[22] = r_31[22] /*27566*/;
  assign m_32[23] = r_31[23] /*27565*/;
  assign m_32[24] = r_31[24] /*27564*/;
  assign m_32[25] = r_31[25] /*27563*/;
  assign m_32[26] = r_31[26] /*27562*/;
  assign m_32[27] = r_31[27] /*27561*/;
  assign m_32[28] = r_31[28] /*27560*/;
  assign m_32[29] = r_31[29] /*27559*/;
  assign m_32[30] = r_31[30] /*27558*/;
  assign m_32[31] = r_31[31] /*27557*/;
  assign _7072_ = ~q[0] /*27555*/;
  assign _7073_ = sum_32[0] & q[0] /*27554*/;
  assign _7074_ = m_32[0] & _7072_ /*27553*/;
  assign r_32[0] = _7074_ | _7073_ /*27552*/;
  assign _7075_ = ~q[0] /*27551*/;
  assign _7076_ = sum_32[1] & q[0] /*27550*/;
  assign _7077_ = m_32[1] & _7075_ /*27549*/;
  assign r_32[1] = _7077_ | _7076_ /*27548*/;
  assign _7078_ = ~q[0] /*27547*/;
  assign _7079_ = sum_32[2] & q[0] /*27546*/;
  assign _7080_ = m_32[2] & _7078_ /*27545*/;
  assign r_32[2] = _7080_ | _7079_ /*27544*/;
  assign _7081_ = ~q[0] /*27543*/;
  assign _7082_ = sum_32[3] & q[0] /*27542*/;
  assign _7083_ = m_32[3] & _7081_ /*27541*/;
  assign r_32[3] = _7083_ | _7082_ /*27540*/;
  assign _7084_ = ~q[0] /*27539*/;
  assign _7085_ = sum_32[4] & q[0] /*27538*/;
  assign _7086_ = m_32[4] & _7084_ /*27537*/;
  assign r_32[4] = _7086_ | _7085_ /*27536*/;
  assign _7087_ = ~q[0] /*27535*/;
  assign _7088_ = sum_32[5] & q[0] /*27534*/;
  assign _7089_ = m_32[5] & _7087_ /*27533*/;
  assign r_32[5] = _7089_ | _7088_ /*27532*/;
  assign _7090_ = ~q[0] /*27531*/;
  assign _7091_ = sum_32[6] & q[0] /*27530*/;
  assign _7092_ = m_32[6] & _7090_ /*27529*/;
  assign r_32[6] = _7092_ | _7091_ /*27528*/;
  assign _7093_ = ~q[0] /*27527*/;
  assign _7094_ = sum_32[7] & q[0] /*27526*/;
  assign _7095_ = m_32[7] & _7093_ /*27525*/;
  assign r_32[7] = _7095_ | _7094_ /*27524*/;
  assign _7096_ = ~q[0] /*27523*/;
  assign _7097_ = sum_32[8] & q[0] /*27522*/;
  assign _7098_ = m_32[8] & _7096_ /*27521*/;
  assign r_32[8] = _7098_ | _7097_ /*27520*/;
  assign _7099_ = ~q[0] /*27519*/;
  assign _7100_ = sum_32[9] & q[0] /*27518*/;
  assign _7101_ = m_32[9] & _7099_ /*27517*/;
  assign r_32[9] = _7101_ | _7100_ /*27516*/;
  assign _7102_ = ~q[0] /*27515*/;
  assign _7103_ = sum_32[10] & q[0] /*27514*/;
  assign _7104_ = m_32[10] & _7102_ /*27513*/;
  assign r_32[10] = _7104_ | _7103_ /*27512*/;
  assign _7105_ = ~q[0] /*27511*/;
  assign _7106_ = sum_32[11] & q[0] /*27510*/;
  assign _7107_ = m_32[11] & _7105_ /*27509*/;
  assign r_32[11] = _7107_ | _7106_ /*27508*/;
  assign _7108_ = ~q[0] /*27507*/;
  assign _7109_ = sum_32[12] & q[0] /*27506*/;
  assign _7110_ = m_32[12] & _7108_ /*27505*/;
  assign r_32[12] = _7110_ | _7109_ /*27504*/;
  assign _7111_ = ~q[0] /*27503*/;
  assign _7112_ = sum_32[13] & q[0] /*27502*/;
  assign _7113_ = m_32[13] & _7111_ /*27501*/;
  assign r_32[13] = _7113_ | _7112_ /*27500*/;
  assign _7114_ = ~q[0] /*27499*/;
  assign _7115_ = sum_32[14] & q[0] /*27498*/;
  assign _7116_ = m_32[14] & _7114_ /*27497*/;
  assign r_32[14] = _7116_ | _7115_ /*27496*/;
  assign _7117_ = ~q[0] /*27495*/;
  assign _7118_ = sum_32[15] & q[0] /*27494*/;
  assign _7119_ = m_32[15] & _7117_ /*27493*/;
  assign r_32[15] = _7119_ | _7118_ /*27492*/;
  assign _7120_ = ~q[0] /*27491*/;
  assign _7121_ = sum_32[16] & q[0] /*27490*/;
  assign _7122_ = m_32[16] & _7120_ /*27489*/;
  assign r_32[16] = _7122_ | _7121_ /*27488*/;
  assign _7123_ = ~q[0] /*27487*/;
  assign _7124_ = sum_32[17] & q[0] /*27486*/;
  assign _7125_ = m_32[17] & _7123_ /*27485*/;
  assign r_32[17] = _7125_ | _7124_ /*27484*/;
  assign _7126_ = ~q[0] /*27483*/;
  assign _7127_ = sum_32[18] & q[0] /*27482*/;
  assign _7128_ = m_32[18] & _7126_ /*27481*/;
  assign r_32[18] = _7128_ | _7127_ /*27480*/;
  assign _7129_ = ~q[0] /*27479*/;
  assign _7130_ = sum_32[19] & q[0] /*27478*/;
  assign _7131_ = m_32[19] & _7129_ /*27477*/;
  assign r_32[19] = _7131_ | _7130_ /*27476*/;
  assign _7132_ = ~q[0] /*27475*/;
  assign _7133_ = sum_32[20] & q[0] /*27474*/;
  assign _7134_ = m_32[20] & _7132_ /*27473*/;
  assign r_32[20] = _7134_ | _7133_ /*27472*/;
  assign _7135_ = ~q[0] /*27471*/;
  assign _7136_ = sum_32[21] & q[0] /*27470*/;
  assign _7137_ = m_32[21] & _7135_ /*27469*/;
  assign r_32[21] = _7137_ | _7136_ /*27468*/;
  assign _7138_ = ~q[0] /*27467*/;
  assign _7139_ = sum_32[22] & q[0] /*27466*/;
  assign _7140_ = m_32[22] & _7138_ /*27465*/;
  assign r_32[22] = _7140_ | _7139_ /*27464*/;
  assign _7141_ = ~q[0] /*27463*/;
  assign _7142_ = sum_32[23] & q[0] /*27462*/;
  assign _7143_ = m_32[23] & _7141_ /*27461*/;
  assign r_32[23] = _7143_ | _7142_ /*27460*/;
  assign _7144_ = ~q[0] /*27459*/;
  assign _7145_ = sum_32[24] & q[0] /*27458*/;
  assign _7146_ = m_32[24] & _7144_ /*27457*/;
  assign r_32[24] = _7146_ | _7145_ /*27456*/;
  assign _7147_ = ~q[0] /*27455*/;
  assign _7148_ = sum_32[25] & q[0] /*27454*/;
  assign _7149_ = m_32[25] & _7147_ /*27453*/;
  assign r_32[25] = _7149_ | _7148_ /*27452*/;
  assign _7150_ = ~q[0] /*27451*/;
  assign _7151_ = sum_32[26] & q[0] /*27450*/;
  assign _7152_ = m_32[26] & _7150_ /*27449*/;
  assign r_32[26] = _7152_ | _7151_ /*27448*/;
  assign _7153_ = ~q[0] /*27447*/;
  assign _7154_ = sum_32[27] & q[0] /*27446*/;
  assign _7155_ = m_32[27] & _7153_ /*27445*/;
  assign r_32[27] = _7155_ | _7154_ /*27444*/;
  assign _7156_ = ~q[0] /*27443*/;
  assign _7157_ = sum_32[28] & q[0] /*27442*/;
  assign _7158_ = m_32[28] & _7156_ /*27441*/;
  assign r_32[28] = _7158_ | _7157_ /*27440*/;
  assign _7159_ = ~q[0] /*27439*/;
  assign _7160_ = sum_32[29] & q[0] /*27438*/;
  assign _7161_ = m_32[29] & _7159_ /*27437*/;
  assign r_32[29] = _7161_ | _7160_ /*27436*/;
  assign _7162_ = ~q[0] /*27435*/;
  assign _7163_ = sum_32[30] & q[0] /*27434*/;
  assign _7164_ = m_32[30] & _7162_ /*27433*/;
  assign r_32[30] = _7164_ | _7163_ /*27432*/;
  assign _7165_ = ~q[0] /*27431*/;
  assign _7166_ = sum_32[31] & q[0] /*27430*/;
  assign _7167_ = m_32[31] & _7165_ /*27429*/;
  assign r_32[31] = _7167_ | _7166_ /*27428*/;
  assign rout[0] = r_32[0] /*0*/;
  assign rout[1] = r_32[1] /*1*/;
  assign rout[2] = r_32[2] /*2*/;
  assign rout[3] = r_32[3] /*3*/;
  assign rout[4] = r_32[4] /*4*/;
  assign rout[5] = r_32[5] /*5*/;
  assign rout[6] = r_32[6] /*6*/;
  assign rout[7] = r_32[7] /*7*/;
  assign rout[8] = r_32[8] /*8*/;
  assign rout[9] = r_32[9] /*9*/;
  assign rout[10] = r_32[10] /*10*/;
  assign rout[11] = r_32[11] /*11*/;
  assign rout[12] = r_32[12] /*12*/;
  assign rout[13] = r_32[13] /*13*/;
  assign rout[14] = r_32[14] /*14*/;
  assign rout[15] = r_32[15] /*15*/;
  assign rout[16] = r_32[16] /*16*/;
  assign rout[17] = r_32[17] /*17*/;
  assign rout[18] = r_32[18] /*18*/;
  assign rout[19] = r_32[19] /*19*/;
  assign rout[20] = r_32[20] /*20*/;
  assign rout[21] = r_32[21] /*21*/;
  assign rout[22] = r_32[22] /*22*/;
  assign rout[23] = r_32[23] /*23*/;
  assign rout[24] = r_32[24] /*24*/;
  assign rout[25] = r_32[25] /*25*/;
  assign rout[26] = r_32[26] /*26*/;
  assign rout[27] = r_32[27] /*27*/;
  assign rout[28] = r_32[28] /*28*/;
  assign rout[29] = r_32[29] /*29*/;
  assign rout[30] = r_32[30] /*30*/;
  assign rout[31] = r_32[31] /*31*/;
endmodule