module nonresdivReduced(R_0, D, Q, R_n1);
input [61:0] R_0;
input [30:0] D;
output [31:0] Q;
output [30:0] R_n1;
wire _0_;
wire _1_;
wire _2_;
wire _3_;
wire _4_;
wire _5_;
wire _6_;
wire _7_;
wire _8_;
wire _9_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire _30_;
wire _31_;
wire _32_;
wire _33_;
wire _34_;
wire _35_;
wire _36_;
wire _37_;
wire _38_;
wire _39_;
wire _40_;
wire _41_;
wire _42_;
wire _43_;
wire _44_;
wire _45_;
wire _46_;
wire _47_;
wire _48_;
wire _49_;
wire _50_;
wire _51_;
wire _52_;
wire _53_;
wire _54_;
wire _55_;
wire _56_;
wire _57_;
wire _58_;
wire _59_;
wire _60_;
wire _61_;
wire _62_;
wire _63_;
wire _64_;
wire _65_;
wire _66_;
wire _67_;
wire _68_;
wire _69_;
wire _70_;
wire _71_;
wire _72_;
wire _73_;
wire _74_;
wire _75_;
wire _76_;
wire _77_;
wire _78_;
wire _79_;
wire _80_;
wire _81_;
wire _82_;
wire _83_;
wire _84_;
wire _85_;
wire _86_;
wire _87_;
wire _88_;
wire _89_;
wire _90_;
wire _91_;
wire _92_;
wire _93_;
wire _94_;
wire _95_;
wire _96_;
wire _97_;
wire _98_;
wire _99_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
wire _255_;
wire _256_;
wire _257_;
wire _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire _267_;
wire _268_;
wire _269_;
wire _270_;
wire _271_;
wire _272_;
wire _273_;
wire _274_;
wire _275_;
wire _276_;
wire _277_;
wire _278_;
wire _279_;
wire _280_;
wire _281_;
wire _282_;
wire _283_;
wire _284_;
wire _285_;
wire _286_;
wire _287_;
wire _288_;
wire _289_;
wire _290_;
wire _291_;
wire _292_;
wire _293_;
wire _294_;
wire _295_;
wire _296_;
wire _297_;
wire _298_;
wire _299_;
wire _300_;
wire _301_;
wire _302_;
wire _303_;
wire _304_;
wire _305_;
wire _306_;
wire _307_;
wire _308_;
wire _309_;
wire _310_;
wire _311_;
wire _312_;
wire _313_;
wire _314_;
wire _315_;
wire _316_;
wire _317_;
wire _318_;
wire _319_;
wire _320_;
wire _321_;
wire _322_;
wire _323_;
wire _324_;
wire _325_;
wire _326_;
wire _327_;
wire _328_;
wire _329_;
wire _330_;
wire _331_;
wire _332_;
wire _333_;
wire _334_;
wire _335_;
wire _336_;
wire _337_;
wire _338_;
wire _339_;
wire _340_;
wire _341_;
wire _342_;
wire _343_;
wire _344_;
wire _345_;
wire _346_;
wire _347_;
wire _348_;
wire _349_;
wire _350_;
wire _351_;
wire _352_;
wire _353_;
wire _354_;
wire _355_;
wire _356_;
wire _357_;
wire _358_;
wire _359_;
wire _360_;
wire _361_;
wire _362_;
wire _363_;
wire _364_;
wire _365_;
wire _366_;
wire _367_;
wire _368_;
wire _369_;
wire _370_;
wire _371_;
wire _372_;
wire _373_;
wire _374_;
wire _375_;
wire _376_;
wire _377_;
wire _378_;
wire _379_;
wire _380_;
wire _381_;
wire _382_;
wire _383_;
wire _384_;
wire _385_;
wire _386_;
wire _387_;
wire _388_;
wire _389_;
wire _390_;
wire _391_;
wire _392_;
wire _393_;
wire _394_;
wire _395_;
wire _396_;
wire _397_;
wire _398_;
wire _399_;
wire _400_;
wire _401_;
wire _402_;
wire _403_;
wire _404_;
wire _405_;
wire _406_;
wire _407_;
wire _408_;
wire _409_;
wire _410_;
wire _411_;
wire _412_;
wire _413_;
wire _414_;
wire _415_;
wire _416_;
wire _417_;
wire _418_;
wire _419_;
wire _420_;
wire _421_;
wire _422_;
wire _423_;
wire _424_;
wire _425_;
wire _426_;
wire _427_;
wire _428_;
wire _429_;
wire _430_;
wire _431_;
wire _432_;
wire _433_;
wire _434_;
wire _435_;
wire _436_;
wire _437_;
wire _438_;
wire _439_;
wire _440_;
wire _441_;
wire _442_;
wire _443_;
wire _444_;
wire _445_;
wire _446_;
wire _447_;
wire _448_;
wire _449_;
wire _450_;
wire _451_;
wire _452_;
wire _453_;
wire _454_;
wire _455_;
wire _456_;
wire _457_;
wire _458_;
wire _459_;
wire _460_;
wire _461_;
wire _462_;
wire _463_;
wire _464_;
wire _465_;
wire _466_;
wire _467_;
wire _468_;
wire _469_;
wire _470_;
wire _471_;
wire _472_;
wire _473_;
wire _474_;
wire _475_;
wire _476_;
wire _477_;
wire _478_;
wire _479_;
wire _480_;
wire _481_;
wire _482_;
wire _483_;
wire _484_;
wire _485_;
wire _486_;
wire _487_;
wire _488_;
wire _489_;
wire _490_;
wire _491_;
wire _492_;
wire _493_;
wire _494_;
wire _495_;
wire _496_;
wire _497_;
wire _498_;
wire _499_;
wire _500_;
wire _501_;
wire _502_;
wire _503_;
wire _504_;
wire _505_;
wire _506_;
wire _507_;
wire _508_;
wire _509_;
wire _510_;
wire _511_;
wire _512_;
wire _513_;
wire _514_;
wire _515_;
wire _516_;
wire _517_;
wire _518_;
wire _519_;
wire _520_;
wire _521_;
wire _522_;
wire _523_;
wire _524_;
wire _525_;
wire _526_;
wire _527_;
wire _528_;
wire _529_;
wire _530_;
wire _531_;
wire _532_;
wire _533_;
wire _534_;
wire _535_;
wire _536_;
wire _537_;
wire _538_;
wire _539_;
wire _540_;
wire _541_;
wire _542_;
wire _543_;
wire _544_;
wire _545_;
wire _546_;
wire _547_;
wire _548_;
wire _549_;
wire _550_;
wire _551_;
wire _552_;
wire _553_;
wire _554_;
wire _555_;
wire _556_;
wire _557_;
wire _558_;
wire _559_;
wire _560_;
wire _561_;
wire _562_;
wire _563_;
wire _564_;
wire _565_;
wire _566_;
wire _567_;
wire _568_;
wire _569_;
wire _570_;
wire _571_;
wire _572_;
wire _573_;
wire _574_;
wire _575_;
wire _576_;
wire _577_;
wire _578_;
wire _579_;
wire _580_;
wire _581_;
wire _582_;
wire _583_;
wire _584_;
wire _585_;
wire _586_;
wire _587_;
wire _588_;
wire _589_;
wire _590_;
wire _591_;
wire _592_;
wire _593_;
wire _594_;
wire _595_;
wire _596_;
wire _597_;
wire _598_;
wire _599_;
wire _600_;
wire _601_;
wire _602_;
wire _603_;
wire _604_;
wire _605_;
wire _606_;
wire _607_;
wire _608_;
wire _609_;
wire _610_;
wire _611_;
wire _612_;
wire _613_;
wire _614_;
wire _615_;
wire _616_;
wire _617_;
wire _618_;
wire _619_;
wire _620_;
wire _621_;
wire _622_;
wire _623_;
wire _624_;
wire _625_;
wire _626_;
wire _627_;
wire _628_;
wire _629_;
wire _630_;
wire _631_;
wire _632_;
wire _633_;
wire _634_;
wire _635_;
wire _636_;
wire _637_;
wire _638_;
wire _639_;
wire _640_;
wire _641_;
wire _642_;
wire _643_;
wire _644_;
wire _645_;
wire _646_;
wire _647_;
wire _648_;
wire _649_;
wire _650_;
wire _651_;
wire _652_;
wire _653_;
wire _654_;
wire _655_;
wire _656_;
wire _657_;
wire _658_;
wire _659_;
wire _660_;
wire _661_;
wire _662_;
wire _663_;
wire _664_;
wire _665_;
wire _666_;
wire _667_;
wire _668_;
wire _669_;
wire _670_;
wire _671_;
wire _672_;
wire _673_;
wire _674_;
wire _675_;
wire _676_;
wire _677_;
wire _678_;
wire _679_;
wire _680_;
wire _681_;
wire _682_;
wire _683_;
wire _684_;
wire _685_;
wire _686_;
wire _687_;
wire _688_;
wire _689_;
wire _690_;
wire _691_;
wire _692_;
wire _693_;
wire _694_;
wire _695_;
wire _696_;
wire _697_;
wire _698_;
wire _699_;
wire _700_;
wire _701_;
wire _702_;
wire _703_;
wire _704_;
wire _705_;
wire _706_;
wire _707_;
wire _708_;
wire _709_;
wire _710_;
wire _711_;
wire _712_;
wire _713_;
wire _714_;
wire _715_;
wire _716_;
wire _717_;
wire _718_;
wire _719_;
wire _720_;
wire _721_;
wire _722_;
wire _723_;
wire _724_;
wire _725_;
wire _726_;
wire _727_;
wire _728_;
wire _729_;
wire _730_;
wire _731_;
wire _732_;
wire _733_;
wire _734_;
wire _735_;
wire _736_;
wire _737_;
wire _738_;
wire _739_;
wire _740_;
wire _741_;
wire _742_;
wire _743_;
wire _744_;
wire _745_;
wire _746_;
wire _747_;
wire _748_;
wire _749_;
wire _750_;
wire _751_;
wire _752_;
wire _753_;
wire _754_;
wire _755_;
wire _756_;
wire _757_;
wire _758_;
wire _759_;
wire _760_;
wire _761_;
wire _762_;
wire _763_;
wire _764_;
wire _765_;
wire _766_;
wire _767_;
wire _768_;
wire _769_;
wire _770_;
wire _771_;
wire _772_;
wire _773_;
wire _774_;
wire _775_;
wire _776_;
wire _777_;
wire _778_;
wire _779_;
wire _780_;
wire _781_;
wire _782_;
wire _783_;
wire _784_;
wire _785_;
wire _786_;
wire _787_;
wire _788_;
wire _789_;
wire _790_;
wire _791_;
wire _792_;
wire _793_;
wire _794_;
wire _795_;
wire _796_;
wire _797_;
wire _798_;
wire _799_;
wire _800_;
wire _801_;
wire _802_;
wire _803_;
wire _804_;
wire _805_;
wire _806_;
wire _807_;
wire _808_;
wire _809_;
wire _810_;
wire _811_;
wire _812_;
wire _813_;
wire _814_;
wire _815_;
wire _816_;
wire _817_;
wire _818_;
wire _819_;
wire _820_;
wire _821_;
wire _822_;
wire _823_;
wire _824_;
wire _825_;
wire _826_;
wire _827_;
wire _828_;
wire _829_;
wire _830_;
wire _831_;
wire _832_;
wire _833_;
wire _834_;
wire _835_;
wire _836_;
wire _837_;
wire _838_;
wire _839_;
wire _840_;
wire _841_;
wire _842_;
wire _843_;
wire _844_;
wire _845_;
wire _846_;
wire _847_;
wire _848_;
wire _849_;
wire _850_;
wire _851_;
wire _852_;
wire _853_;
wire _854_;
wire _855_;
wire _856_;
wire _857_;
wire _858_;
wire _859_;
wire _860_;
wire _861_;
wire _862_;
wire _863_;
wire _864_;
wire _865_;
wire _866_;
wire _867_;
wire _868_;
wire _869_;
wire _870_;
wire _871_;
wire _872_;
wire _873_;
wire _874_;
wire _875_;
wire _876_;
wire _877_;
wire _878_;
wire _879_;
wire _880_;
wire _881_;
wire _882_;
wire _883_;
wire _884_;
wire _885_;
wire _886_;
wire _887_;
wire _888_;
wire _889_;
wire _890_;
wire _891_;
wire _892_;
wire _893_;
wire _894_;
wire _895_;
wire _896_;
wire _897_;
wire _898_;
wire _899_;
wire _900_;
wire _901_;
wire _902_;
wire _903_;
wire _904_;
wire _905_;
wire _906_;
wire _907_;
wire _908_;
wire _909_;
wire _910_;
wire _911_;
wire _912_;
wire _913_;
wire _914_;
wire _915_;
wire _916_;
wire _917_;
wire _918_;
wire _919_;
wire _920_;
wire _921_;
wire _922_;
wire _923_;
wire _924_;
wire _925_;
wire _926_;
wire _927_;
wire _928_;
wire _929_;
wire _930_;
wire _931_;
wire _932_;
wire _933_;
wire _934_;
wire _935_;
wire _936_;
wire _937_;
wire _938_;
wire _939_;
wire _940_;
wire _941_;
wire _942_;
wire _943_;
wire _944_;
wire _945_;
wire _946_;
wire _947_;
wire _948_;
wire _949_;
wire _950_;
wire _951_;
wire _952_;
wire _953_;
wire _954_;
wire _955_;
wire _956_;
wire _957_;
wire _958_;
wire _959_;
wire _960_;
wire _961_;
wire _962_;
wire _963_;
wire _964_;
wire _965_;
wire _966_;
wire _967_;
wire _968_;
wire _969_;
wire _970_;
wire _971_;
wire _972_;
wire _973_;
wire _974_;
wire _975_;
wire _976_;
wire _977_;
wire _978_;
wire _979_;
wire _980_;
wire _981_;
wire _982_;
wire _983_;
wire _984_;
wire _985_;
wire _986_;
wire _987_;
wire _988_;
wire _989_;
wire _990_;
wire _991_;
wire _992_;
wire _993_;
wire _994_;
wire _995_;
wire _996_;
wire _997_;
wire _998_;
wire _999_;
wire _1000_;
wire _1001_;
wire _1002_;
wire _1003_;
wire _1004_;
wire _1005_;
wire _1006_;
wire _1007_;
wire _1008_;
wire _1009_;
wire _1010_;
wire _1011_;
wire _1012_;
wire _1013_;
wire _1014_;
wire _1015_;
wire _1016_;
wire _1017_;
wire _1018_;
wire _1019_;
wire _1020_;
wire _1021_;
wire _1022_;
wire _1023_;
wire _1024_;
wire _1025_;
wire _1026_;
wire _1027_;
wire _1028_;
wire _1029_;
wire _1030_;
wire _1031_;
wire _1032_;
wire _1033_;
wire _1034_;
wire _1035_;
wire _1036_;
wire _1037_;
wire _1038_;
wire _1039_;
wire _1040_;
wire _1041_;
wire _1042_;
wire _1043_;
wire _1044_;
wire _1045_;
wire _1046_;
wire _1047_;
wire _1048_;
wire _1049_;
wire _1050_;
wire _1051_;
wire _1052_;
wire _1053_;
wire _1054_;
wire _1055_;
wire _1056_;
wire _1057_;
wire _1058_;
wire _1059_;
wire _1060_;
wire _1061_;
wire _1062_;
wire _1063_;
wire _1064_;
wire _1065_;
wire _1066_;
wire _1067_;
wire _1068_;
wire _1069_;
wire _1070_;
wire _1071_;
wire _1072_;
wire _1073_;
wire _1074_;
wire _1075_;
wire _1076_;
wire _1077_;
wire _1078_;
wire _1079_;
wire _1080_;
wire _1081_;
wire _1082_;
wire _1083_;
wire _1084_;
wire _1085_;
wire _1086_;
wire _1087_;
wire _1088_;
wire _1089_;
wire _1090_;
wire _1091_;
wire _1092_;
wire _1093_;
wire _1094_;
wire _1095_;
wire _1096_;
wire _1097_;
wire _1098_;
wire _1099_;
wire _1100_;
wire _1101_;
wire _1102_;
wire _1103_;
wire _1104_;
wire _1105_;
wire _1106_;
wire _1107_;
wire _1108_;
wire _1109_;
wire _1110_;
wire _1111_;
wire _1112_;
wire _1113_;
wire _1114_;
wire _1115_;
wire _1116_;
wire _1117_;
wire _1118_;
wire _1119_;
wire _1120_;
wire _1121_;
wire _1122_;
wire _1123_;
wire _1124_;
wire _1125_;
wire _1126_;
wire _1127_;
wire _1128_;
wire _1129_;
wire _1130_;
wire _1131_;
wire _1132_;
wire _1133_;
wire _1134_;
wire _1135_;
wire _1136_;
wire _1137_;
wire _1138_;
wire _1139_;
wire _1140_;
wire _1141_;
wire _1142_;
wire _1143_;
wire _1144_;
wire _1145_;
wire _1146_;
wire _1147_;
wire _1148_;
wire _1149_;
wire _1150_;
wire _1151_;
wire _1152_;
wire _1153_;
wire _1154_;
wire _1155_;
wire _1156_;
wire _1157_;
wire _1158_;
wire _1159_;
wire _1160_;
wire _1161_;
wire _1162_;
wire _1163_;
wire _1164_;
wire _1165_;
wire _1166_;
wire _1167_;
wire _1168_;
wire _1169_;
wire _1170_;
wire _1171_;
wire _1172_;
wire _1173_;
wire _1174_;
wire _1175_;
wire _1176_;
wire _1177_;
wire _1178_;
wire _1179_;
wire _1180_;
wire _1181_;
wire _1182_;
wire _1183_;
wire _1184_;
wire _1185_;
wire _1186_;
wire _1187_;
wire _1188_;
wire _1189_;
wire _1190_;
wire _1191_;
wire _1192_;
wire _1193_;
wire _1194_;
wire _1195_;
wire _1196_;
wire _1197_;
wire _1198_;
wire _1199_;
wire _1200_;
wire _1201_;
wire _1202_;
wire _1203_;
wire _1204_;
wire _1205_;
wire _1206_;
wire _1207_;
wire _1208_;
wire _1209_;
wire _1210_;
wire _1211_;
wire _1212_;
wire _1213_;
wire _1214_;
wire _1215_;
wire _1216_;
wire _1217_;
wire _1218_;
wire _1219_;
wire _1220_;
wire _1221_;
wire _1222_;
wire _1223_;
wire _1224_;
wire _1225_;
wire _1226_;
wire _1227_;
wire _1228_;
wire _1229_;
wire _1230_;
wire _1231_;
wire _1232_;
wire _1233_;
wire _1234_;
wire _1235_;
wire _1236_;
wire _1237_;
wire _1238_;
wire _1239_;
wire _1240_;
wire _1241_;
wire _1242_;
wire _1243_;
wire _1244_;
wire _1245_;
wire _1246_;
wire _1247_;
wire _1248_;
wire _1249_;
wire _1250_;
wire _1251_;
wire _1252_;
wire _1253_;
wire _1254_;
wire _1255_;
wire _1256_;
wire _1257_;
wire _1258_;
wire _1259_;
wire _1260_;
wire _1261_;
wire _1262_;
wire _1263_;
wire _1264_;
wire _1265_;
wire _1266_;
wire _1267_;
wire _1268_;
wire _1269_;
wire _1270_;
wire _1271_;
wire _1272_;
wire _1273_;
wire _1274_;
wire _1275_;
wire _1276_;
wire _1277_;
wire _1278_;
wire _1279_;
wire _1280_;
wire _1281_;
wire _1282_;
wire _1283_;
wire _1284_;
wire _1285_;
wire _1286_;
wire _1287_;
wire _1288_;
wire _1289_;
wire _1290_;
wire _1291_;
wire _1292_;
wire _1293_;
wire _1294_;
wire _1295_;
wire _1296_;
wire _1297_;
wire _1298_;
wire _1299_;
wire _1300_;
wire _1301_;
wire _1302_;
wire _1303_;
wire _1304_;
wire _1305_;
wire _1306_;
wire _1307_;
wire _1308_;
wire _1309_;
wire _1310_;
wire _1311_;
wire _1312_;
wire _1313_;
wire _1314_;
wire _1315_;
wire _1316_;
wire _1317_;
wire _1318_;
wire _1319_;
wire _1320_;
wire _1321_;
wire _1322_;
wire _1323_;
wire _1324_;
wire _1325_;
wire _1326_;
wire _1327_;
wire _1328_;
wire _1329_;
wire _1330_;
wire _1331_;
wire _1332_;
wire _1333_;
wire _1334_;
wire _1335_;
wire _1336_;
wire _1337_;
wire _1338_;
wire _1339_;
wire _1340_;
wire _1341_;
wire _1342_;
wire _1343_;
wire _1344_;
wire _1345_;
wire _1346_;
wire _1347_;
wire _1348_;
wire _1349_;
wire _1350_;
wire _1351_;
wire _1352_;
wire _1353_;
wire _1354_;
wire _1355_;
wire _1356_;
wire _1357_;
wire _1358_;
wire _1359_;
wire _1360_;
wire _1361_;
wire _1362_;
wire _1363_;
wire _1364_;
wire _1365_;
wire _1366_;
wire _1367_;
wire _1368_;
wire _1369_;
wire _1370_;
wire _1371_;
wire _1372_;
wire _1373_;
wire _1374_;
wire _1375_;
wire _1376_;
wire _1377_;
wire _1378_;
wire _1379_;
wire _1380_;
wire _1381_;
wire _1382_;
wire _1383_;
wire _1384_;
wire _1385_;
wire _1386_;
wire _1387_;
wire _1388_;
wire _1389_;
wire _1390_;
wire _1391_;
wire _1392_;
wire _1393_;
wire _1394_;
wire _1395_;
wire _1396_;
wire _1397_;
wire _1398_;
wire _1399_;
wire _1400_;
wire _1401_;
wire _1402_;
wire _1403_;
wire _1404_;
wire _1405_;
wire _1406_;
wire _1407_;
wire _1408_;
wire _1409_;
wire _1410_;
wire _1411_;
wire _1412_;
wire _1413_;
wire _1414_;
wire _1415_;
wire _1416_;
wire _1417_;
wire _1418_;
wire _1419_;
wire _1420_;
wire _1421_;
wire _1422_;
wire _1423_;
wire _1424_;
wire _1425_;
wire _1426_;
wire _1427_;
wire _1428_;
wire _1429_;
wire _1430_;
wire _1431_;
wire _1432_;
wire _1433_;
wire _1434_;
wire _1435_;
wire _1436_;
wire _1437_;
wire _1438_;
wire _1439_;
wire _1440_;
wire _1441_;
wire _1442_;
wire _1443_;
wire _1444_;
wire _1445_;
wire _1446_;
wire _1447_;
wire _1448_;
wire _1449_;
wire _1450_;
wire _1451_;
wire _1452_;
wire _1453_;
wire _1454_;
wire _1455_;
wire _1456_;
wire _1457_;
wire _1458_;
wire _1459_;
wire _1460_;
wire _1461_;
wire _1462_;
wire _1463_;
wire _1464_;
wire _1465_;
wire _1466_;
wire _1467_;
wire _1468_;
wire _1469_;
wire _1470_;
wire _1471_;
wire _1472_;
wire _1473_;
wire _1474_;
wire _1475_;
wire _1476_;
wire _1477_;
wire _1478_;
wire _1479_;
wire _1480_;
wire _1481_;
wire _1482_;
wire _1483_;
wire _1484_;
wire _1485_;
wire _1486_;
wire _1487_;
wire _1488_;
wire _1489_;
wire _1490_;
wire _1491_;
wire _1492_;
wire _1493_;
wire _1494_;
wire _1495_;
wire _1496_;
wire _1497_;
wire _1498_;
wire _1499_;
wire _1500_;
wire _1501_;
wire _1502_;
wire _1503_;
wire _1504_;
wire _1505_;
wire _1506_;
wire _1507_;
wire _1508_;
wire _1509_;
wire _1510_;
wire _1511_;
wire _1512_;
wire _1513_;
wire _1514_;
wire _1515_;
wire _1516_;
wire _1517_;
wire _1518_;
wire _1519_;
wire _1520_;
wire _1521_;
wire _1522_;
wire _1523_;
wire _1524_;
wire _1525_;
wire _1526_;
wire _1527_;
wire _1528_;
wire _1529_;
wire _1530_;
wire _1531_;
wire _1532_;
wire _1533_;
wire _1534_;
wire _1535_;
wire _1536_;
wire _1537_;
wire _1538_;
wire _1539_;
wire _1540_;
wire _1541_;
wire _1542_;
wire _1543_;
wire _1544_;
wire _1545_;
wire _1546_;
wire _1547_;
wire _1548_;
wire _1549_;
wire _1550_;
wire _1551_;
wire _1552_;
wire _1553_;
wire _1554_;
wire _1555_;
wire _1556_;
wire _1557_;
wire _1558_;
wire _1559_;
wire _1560_;
wire _1561_;
wire _1562_;
wire _1563_;
wire _1564_;
wire _1565_;
wire _1566_;
wire _1567_;
wire _1568_;
wire _1569_;
wire _1570_;
wire _1571_;
wire _1572_;
wire _1573_;
wire _1574_;
wire _1575_;
wire _1576_;
wire _1577_;
wire _1578_;
wire _1579_;
wire _1580_;
wire _1581_;
wire _1582_;
wire _1583_;
wire _1584_;
wire _1585_;
wire _1586_;
wire _1587_;
wire _1588_;
wire _1589_;
wire _1590_;
wire _1591_;
wire _1592_;
wire _1593_;
wire _1594_;
wire _1595_;
wire _1596_;
wire _1597_;
wire _1598_;
wire _1599_;
wire _1600_;
wire _1601_;
wire _1602_;
wire _1603_;
wire _1604_;
wire _1605_;
wire _1606_;
wire _1607_;
wire _1608_;
wire _1609_;
wire _1610_;
wire _1611_;
wire _1612_;
wire _1613_;
wire _1614_;
wire _1615_;
wire _1616_;
wire _1617_;
wire _1618_;
wire _1619_;
wire _1620_;
wire _1621_;
wire _1622_;
wire _1623_;
wire _1624_;
wire _1625_;
wire _1626_;
wire _1627_;
wire _1628_;
wire _1629_;
wire _1630_;
wire _1631_;
wire _1632_;
wire _1633_;
wire _1634_;
wire _1635_;
wire _1636_;
wire _1637_;
wire _1638_;
wire _1639_;
wire _1640_;
wire _1641_;
wire _1642_;
wire _1643_;
wire _1644_;
wire _1645_;
wire _1646_;
wire _1647_;
wire _1648_;
wire _1649_;
wire _1650_;
wire _1651_;
wire _1652_;
wire _1653_;
wire _1654_;
wire _1655_;
wire _1656_;
wire _1657_;
wire _1658_;
wire _1659_;
wire _1660_;
wire _1661_;
wire _1662_;
wire _1663_;
wire _1664_;
wire _1665_;
wire _1666_;
wire _1667_;
wire _1668_;
wire _1669_;
wire _1670_;
wire _1671_;
wire _1672_;
wire _1673_;
wire _1674_;
wire _1675_;
wire _1676_;
wire _1677_;
wire _1678_;
wire _1679_;
wire _1680_;
wire _1681_;
wire _1682_;
wire _1683_;
wire _1684_;
wire _1685_;
wire _1686_;
wire _1687_;
wire _1688_;
wire _1689_;
wire _1690_;
wire _1691_;
wire _1692_;
wire _1693_;
wire _1694_;
wire _1695_;
wire _1696_;
wire _1697_;
wire _1698_;
wire _1699_;
wire _1700_;
wire _1701_;
wire _1702_;
wire _1703_;
wire _1704_;
wire _1705_;
wire _1706_;
wire _1707_;
wire _1708_;
wire _1709_;
wire _1710_;
wire _1711_;
wire _1712_;
wire _1713_;
wire _1714_;
wire _1715_;
wire _1716_;
wire _1717_;
wire _1718_;
wire _1719_;
wire _1720_;
wire _1721_;
wire _1722_;
wire _1723_;
wire _1724_;
wire _1725_;
wire _1726_;
wire _1727_;
wire _1728_;
wire _1729_;
wire _1730_;
wire _1731_;
wire _1732_;
wire _1733_;
wire _1734_;
wire _1735_;
wire _1736_;
wire _1737_;
wire _1738_;
wire _1739_;
wire _1740_;
wire _1741_;
wire _1742_;
wire _1743_;
wire _1744_;
wire _1745_;
wire _1746_;
wire _1747_;
wire _1748_;
wire _1749_;
wire _1750_;
wire _1751_;
wire _1752_;
wire _1753_;
wire _1754_;
wire _1755_;
wire _1756_;
wire _1757_;
wire _1758_;
wire _1759_;
wire _1760_;
wire _1761_;
wire _1762_;
wire _1763_;
wire _1764_;
wire _1765_;
wire _1766_;
wire _1767_;
wire _1768_;
wire _1769_;
wire _1770_;
wire _1771_;
wire _1772_;
wire _1773_;
wire _1774_;
wire _1775_;
wire _1776_;
wire _1777_;
wire _1778_;
wire _1779_;
wire _1780_;
wire _1781_;
wire _1782_;
wire _1783_;
wire _1784_;
wire _1785_;
wire _1786_;
wire _1787_;
wire _1788_;
wire _1789_;
wire _1790_;
wire _1791_;
wire _1792_;
wire _1793_;
wire _1794_;
wire _1795_;
wire _1796_;
wire _1797_;
wire _1798_;
wire _1799_;
wire _1800_;
wire _1801_;
wire _1802_;
wire _1803_;
wire _1804_;
wire _1805_;
wire _1806_;
wire _1807_;
wire _1808_;
wire _1809_;
wire _1810_;
wire _1811_;
wire _1812_;
wire _1813_;
wire _1814_;
wire _1815_;
wire _1816_;
wire _1817_;
wire _1818_;
wire _1819_;
wire _1820_;
wire _1821_;
wire _1822_;
wire _1823_;
wire _1824_;
wire _1825_;
wire _1826_;
wire _1827_;
wire _1828_;
wire _1829_;
wire _1830_;
wire _1831_;
wire _1832_;
wire _1833_;
wire _1834_;
wire _1835_;
wire _1836_;
wire _1837_;
wire _1838_;
wire _1839_;
wire _1840_;
wire _1841_;
wire _1842_;
wire _1843_;
wire _1844_;
wire _1845_;
wire _1846_;
wire _1847_;
wire _1848_;
wire _1849_;
wire _1850_;
wire _1851_;
wire _1852_;
wire _1853_;
wire _1854_;
wire _1855_;
wire _1856_;
wire _1857_;
wire _1858_;
wire _1859_;
wire _1860_;
wire _1861_;
wire _1862_;
wire _1863_;
wire _1864_;
wire _1865_;
wire _1866_;
wire _1867_;
wire _1868_;
wire _1869_;
wire _1870_;
wire _1871_;
wire _1872_;
wire _1873_;
wire _1874_;
wire _1875_;
wire _1876_;
wire _1877_;
wire _1878_;
wire _1879_;
wire _1880_;
wire _1881_;
wire _1882_;
wire _1883_;
wire _1884_;
wire _1885_;
wire _1886_;
wire _1887_;
wire _1888_;
wire _1889_;
wire _1890_;
wire _1891_;
wire _1892_;
wire _1893_;
wire _1894_;
wire _1895_;
wire _1896_;
wire _1897_;
wire _1898_;
wire _1899_;
wire _1900_;
wire _1901_;
wire _1902_;
wire _1903_;
wire _1904_;
wire _1905_;
wire _1906_;
wire _1907_;
wire _1908_;
wire _1909_;
wire _1910_;
wire _1911_;
wire _1912_;
wire _1913_;
wire _1914_;
wire _1915_;
wire _1916_;
wire _1917_;
wire _1918_;
wire _1919_;
wire _1920_;
wire _1921_;
wire _1922_;
wire _1923_;
wire _1924_;
wire _1925_;
wire _1926_;
wire _1927_;
wire _1928_;
wire _1929_;
wire _1930_;
wire _1931_;
wire _1932_;
wire _1933_;
wire _1934_;
wire _1935_;
wire _1936_;
wire _1937_;
wire _1938_;
wire _1939_;
wire _1940_;
wire _1941_;
wire _1942_;
wire _1943_;
wire _1944_;
wire _1945_;
wire _1946_;
wire _1947_;
wire _1948_;
wire _1949_;
wire _1950_;
wire _1951_;
wire _1952_;
wire _1953_;
wire _1954_;
wire _1955_;
wire _1956_;
wire _1957_;
wire _1958_;
wire _1959_;
wire _1960_;
wire _1961_;
wire _1962_;
wire _1963_;
wire _1964_;
wire _1965_;
wire _1966_;
wire _1967_;
wire _1968_;
wire _1969_;
wire _1970_;
wire _1971_;
wire _1972_;
wire _1973_;
wire _1974_;
wire _1975_;
wire _1976_;
wire _1977_;
wire _1978_;
wire _1979_;
wire _1980_;
wire _1981_;
wire _1982_;
wire _1983_;
wire _1984_;
wire _1985_;
wire _1986_;
wire _1987_;
wire _1988_;
wire _1989_;
wire _1990_;
wire _1991_;
wire _1992_;
wire _1993_;
wire _1994_;
wire _1995_;
wire _1996_;
wire _1997_;
wire _1998_;
wire _1999_;
wire _2000_;
wire _2001_;
wire _2002_;
wire _2003_;
wire _2004_;
wire _2005_;
wire _2006_;
wire _2007_;
wire _2008_;
wire _2009_;
wire _2010_;
wire _2011_;
wire _2012_;
wire _2013_;
wire _2014_;
wire _2015_;
wire _2016_;
wire _2017_;
wire _2018_;
wire _2019_;
wire _2020_;
wire _2021_;
wire _2022_;
wire _2023_;
wire _2024_;
wire _2025_;
wire _2026_;
wire _2027_;
wire _2028_;
wire _2029_;
wire _2030_;
wire _2031_;
wire _2032_;
wire _2033_;
wire _2034_;
wire _2035_;
wire _2036_;
wire _2037_;
wire _2038_;
wire _2039_;
wire _2040_;
wire _2041_;
wire _2042_;
wire _2043_;
wire _2044_;
wire _2045_;
wire _2046_;
wire _2047_;
wire _2048_;
wire _2049_;
wire _2050_;
wire _2051_;
wire _2052_;
wire _2053_;
wire _2054_;
wire _2055_;
wire _2056_;
wire _2057_;
wire _2058_;
wire _2059_;
wire _2060_;
wire _2061_;
wire _2062_;
wire _2063_;
wire _2064_;
wire _2065_;
wire _2066_;
wire _2067_;
wire _2068_;
wire _2069_;
wire _2070_;
wire _2071_;
wire _2072_;
wire _2073_;
wire _2074_;
wire _2075_;
wire _2076_;
wire _2077_;
wire _2078_;
wire _2079_;
wire _2080_;
wire _2081_;
wire _2082_;
wire _2083_;
wire _2084_;
wire _2085_;
wire _2086_;
wire _2087_;
wire _2088_;
wire _2089_;
wire _2090_;
wire _2091_;
wire _2092_;
wire _2093_;
wire _2094_;
wire _2095_;
wire _2096_;
wire _2097_;
wire _2098_;
wire _2099_;
wire _2100_;
wire _2101_;
wire _2102_;
wire _2103_;
wire _2104_;
wire _2105_;
wire _2106_;
wire _2107_;
wire _2108_;
wire _2109_;
wire _2110_;
wire _2111_;
wire _2112_;
wire _2113_;
wire _2114_;
wire _2115_;
wire _2116_;
wire _2117_;
wire _2118_;
wire _2119_;
wire _2120_;
wire _2121_;
wire _2122_;
wire _2123_;
wire _2124_;
wire _2125_;
wire _2126_;
wire _2127_;
wire _2128_;
wire _2129_;
wire _2130_;
wire _2131_;
wire _2132_;
wire _2133_;
wire _2134_;
wire _2135_;
wire _2136_;
wire _2137_;
wire _2138_;
wire _2139_;
wire _2140_;
wire _2141_;
wire _2142_;
wire _2143_;
wire _2144_;
wire _2145_;
wire _2146_;
wire _2147_;
wire _2148_;
wire _2149_;
wire _2150_;
wire _2151_;
wire _2152_;
wire _2153_;
wire _2154_;
wire _2155_;
wire _2156_;
wire _2157_;
wire _2158_;
wire _2159_;
wire _2160_;
wire _2161_;
wire _2162_;
wire _2163_;
wire _2164_;
wire _2165_;
wire _2166_;
wire _2167_;
wire _2168_;
wire _2169_;
wire _2170_;
wire _2171_;
wire _2172_;
wire _2173_;
wire _2174_;
wire _2175_;
wire _2176_;
wire _2177_;
wire _2178_;
wire _2179_;
wire _2180_;
wire _2181_;
wire _2182_;
wire _2183_;
wire _2184_;
wire _2185_;
wire _2186_;
wire _2187_;
wire _2188_;
wire _2189_;
wire _2190_;
wire _2191_;
wire _2192_;
wire _2193_;
wire _2194_;
wire _2195_;
wire _2196_;
wire _2197_;
wire _2198_;
wire _2199_;
wire _2200_;
wire _2201_;
wire _2202_;
wire _2203_;
wire _2204_;
wire _2205_;
wire _2206_;
wire _2207_;
wire _2208_;
wire _2209_;
wire _2210_;
wire _2211_;
wire _2212_;
wire _2213_;
wire _2214_;
wire _2215_;
wire _2216_;
wire _2217_;
wire _2218_;
wire _2219_;
wire _2220_;
wire _2221_;
wire _2222_;
wire _2223_;
wire _2224_;
wire _2225_;
wire _2226_;
wire _2227_;
wire _2228_;
wire _2229_;
wire _2230_;
wire _2231_;
wire _2232_;
wire _2233_;
wire _2234_;
wire _2235_;
wire _2236_;
wire _2237_;
wire _2238_;
wire _2239_;
wire _2240_;
wire _2241_;
wire _2242_;
wire _2243_;
wire _2244_;
wire _2245_;
wire _2246_;
wire _2247_;
wire _2248_;
wire _2249_;
wire _2250_;
wire _2251_;
wire _2252_;
wire _2253_;
wire _2254_;
wire _2255_;
wire _2256_;
wire _2257_;
wire _2258_;
wire _2259_;
wire _2260_;
wire _2261_;
wire _2262_;
wire _2263_;
wire _2264_;
wire _2265_;
wire _2266_;
wire _2267_;
wire _2268_;
wire _2269_;
wire _2270_;
wire _2271_;
wire _2272_;
wire _2273_;
wire _2274_;
wire _2275_;
wire _2276_;
wire _2277_;
wire _2278_;
wire _2279_;
wire _2280_;
wire _2281_;
wire _2282_;
wire _2283_;
wire _2284_;
wire _2285_;
wire _2286_;
wire _2287_;
wire _2288_;
wire _2289_;
wire _2290_;
wire _2291_;
wire _2292_;
wire _2293_;
wire _2294_;
wire _2295_;
wire _2296_;
wire _2297_;
wire _2298_;
wire _2299_;
wire _2300_;
wire _2301_;
wire _2302_;
wire _2303_;
wire _2304_;
wire _2305_;
wire _2306_;
wire _2307_;
wire _2308_;
wire _2309_;
wire _2310_;
wire _2311_;
wire _2312_;
wire _2313_;
wire _2314_;
wire _2315_;
wire _2316_;
wire _2317_;
wire _2318_;
wire _2319_;
wire _2320_;
wire _2321_;
wire _2322_;
wire _2323_;
wire _2324_;
wire _2325_;
wire _2326_;
wire _2327_;
wire _2328_;
wire _2329_;
wire _2330_;
wire _2331_;
wire _2332_;
wire _2333_;
wire _2334_;
wire _2335_;
wire _2336_;
wire _2337_;
wire _2338_;
wire _2339_;
wire _2340_;
wire _2341_;
wire _2342_;
wire _2343_;
wire _2344_;
wire _2345_;
wire _2346_;
wire _2347_;
wire _2348_;
wire _2349_;
wire _2350_;
wire _2351_;
wire _2352_;
wire _2353_;
wire _2354_;
wire _2355_;
wire _2356_;
wire _2357_;
wire _2358_;
wire _2359_;
wire _2360_;
wire _2361_;
wire _2362_;
wire _2363_;
wire _2364_;
wire _2365_;
wire _2366_;
wire _2367_;
wire _2368_;
wire _2369_;
wire _2370_;
wire _2371_;
wire _2372_;
wire _2373_;
wire _2374_;
wire _2375_;
wire _2376_;
wire _2377_;
wire _2378_;
wire _2379_;
wire _2380_;
wire _2381_;
wire _2382_;
wire _2383_;
wire _2384_;
wire _2385_;
wire _2386_;
wire _2387_;
wire _2388_;
wire _2389_;
wire _2390_;
wire _2391_;
wire _2392_;
wire _2393_;
wire _2394_;
wire _2395_;
wire _2396_;
wire _2397_;
wire _2398_;
wire _2399_;
wire _2400_;
wire _2401_;
wire _2402_;
wire _2403_;
wire _2404_;
wire _2405_;
wire _2406_;
wire _2407_;
wire _2408_;
wire _2409_;
wire _2410_;
wire _2411_;
wire _2412_;
wire _2413_;
wire _2414_;
wire _2415_;
wire _2416_;
wire _2417_;
wire _2418_;
wire _2419_;
wire _2420_;
wire _2421_;
wire _2422_;
wire _2423_;
wire _2424_;
wire _2425_;
wire _2426_;
wire _2427_;
wire _2428_;
wire _2429_;
wire _2430_;
wire _2431_;
wire _2432_;
wire _2433_;
wire _2434_;
wire _2435_;
wire _2436_;
wire _2437_;
wire _2438_;
wire _2439_;
wire _2440_;
wire _2441_;
wire _2442_;
wire _2443_;
wire _2444_;
wire _2445_;
wire _2446_;
wire _2447_;
wire _2448_;
wire _2449_;
wire _2450_;
wire _2451_;
wire _2452_;
wire _2453_;
wire _2454_;
wire _2455_;
wire _2456_;
wire _2457_;
wire _2458_;
wire _2459_;
wire _2460_;
wire _2461_;
wire _2462_;
wire _2463_;
wire _2464_;
wire _2465_;
wire _2466_;
wire _2467_;
wire _2468_;
wire _2469_;
wire _2470_;
wire _2471_;
wire _2472_;
wire _2473_;
wire _2474_;
wire _2475_;
wire _2476_;
wire _2477_;
wire _2478_;
wire _2479_;
wire _2480_;
wire _2481_;
wire _2482_;
wire _2483_;
wire _2484_;
wire _2485_;
wire _2486_;
wire _2487_;
wire _2488_;
wire _2489_;
wire _2490_;
wire _2491_;
wire _2492_;
wire _2493_;
wire _2494_;
wire _2495_;
wire _2496_;
wire _2497_;
wire _2498_;
wire _2499_;
wire _2500_;
wire _2501_;
wire _2502_;
wire _2503_;
wire _2504_;
wire _2505_;
wire _2506_;
wire _2507_;
wire _2508_;
wire _2509_;
wire _2510_;
wire _2511_;
wire _2512_;
wire _2513_;
wire _2514_;
wire _2515_;
wire _2516_;
wire _2517_;
wire _2518_;
wire _2519_;
wire _2520_;
wire _2521_;
wire _2522_;
wire _2523_;
wire _2524_;
wire _2525_;
wire _2526_;
wire _2527_;
wire _2528_;
wire _2529_;
wire _2530_;
wire _2531_;
wire _2532_;
wire _2533_;
wire _2534_;
wire _2535_;
wire _2536_;
wire _2537_;
wire _2538_;
wire _2539_;
wire _2540_;
wire _2541_;
wire _2542_;
wire _2543_;
wire _2544_;
wire _2545_;
wire _2546_;
wire _2547_;
wire _2548_;
wire _2549_;
wire _2550_;
wire _2551_;
wire _2552_;
wire _2553_;
wire _2554_;
wire _2555_;
wire _2556_;
wire _2557_;
wire _2558_;
wire _2559_;
wire _2560_;
wire _2561_;
wire _2562_;
wire _2563_;
wire _2564_;
wire _2565_;
wire _2566_;
wire _2567_;
wire _2568_;
wire _2569_;
wire _2570_;
wire _2571_;
wire _2572_;
wire _2573_;
wire _2574_;
wire _2575_;
wire _2576_;
wire _2577_;
wire _2578_;
wire _2579_;
wire _2580_;
wire _2581_;
wire _2582_;
wire _2583_;
wire _2584_;
wire _2585_;
wire _2586_;
wire _2587_;
wire _2588_;
wire _2589_;
wire _2590_;
wire _2591_;
wire _2592_;
wire _2593_;
wire _2594_;
wire _2595_;
wire _2596_;
wire _2597_;
wire _2598_;
wire _2599_;
wire _2600_;
wire _2601_;
wire _2602_;
wire _2603_;
wire _2604_;
wire _2605_;
wire _2606_;
wire _2607_;
wire _2608_;
wire _2609_;
wire _2610_;
wire _2611_;
wire _2612_;
wire _2613_;
wire _2614_;
wire _2615_;
wire _2616_;
wire _2617_;
wire _2618_;
wire _2619_;
wire _2620_;
wire _2621_;
wire _2622_;
wire _2623_;
wire _2624_;
wire _2625_;
wire _2626_;
wire _2627_;
wire _2628_;
wire _2629_;
wire _2630_;
wire _2631_;
wire _2632_;
wire _2633_;
wire _2634_;
wire _2635_;
wire _2636_;
wire _2637_;
wire _2638_;
wire _2639_;
wire _2640_;
wire _2641_;
wire _2642_;
wire _2643_;
wire _2644_;
wire _2645_;
wire _2646_;
wire _2647_;
wire _2648_;
wire _2649_;
wire _2650_;
wire _2651_;
wire _2652_;
wire _2653_;
wire _2654_;
wire _2655_;
wire _2656_;
wire _2657_;
wire _2658_;
wire _2659_;
wire _2660_;
wire _2661_;
wire _2662_;
wire _2663_;
wire _2664_;
wire _2665_;
wire _2666_;
wire _2667_;
wire _2668_;
wire _2669_;
wire _2670_;
wire _2671_;
wire _2672_;
wire _2673_;
wire _2674_;
wire _2675_;
wire _2676_;
wire _2677_;
wire _2678_;
wire _2679_;
wire _2680_;
wire _2681_;
wire _2682_;
wire _2683_;
wire _2684_;
wire _2685_;
wire _2686_;
wire _2687_;
wire _2688_;
wire _2689_;
wire _2690_;
wire _2691_;
wire _2692_;
wire _2693_;
wire _2694_;
wire _2695_;
wire _2696_;
wire _2697_;
wire _2698_;
wire _2699_;
wire _2700_;
wire _2701_;
wire _2702_;
wire _2703_;
wire _2704_;
wire _2705_;
wire _2706_;
wire _2707_;
wire _2708_;
wire _2709_;
wire _2710_;
wire _2711_;
wire _2712_;
wire _2713_;
wire _2714_;
wire _2715_;
wire _2716_;
wire _2717_;
wire _2718_;
wire _2719_;
wire _2720_;
wire _2721_;
wire _2722_;
wire _2723_;
wire _2724_;
wire _2725_;
wire _2726_;
wire _2727_;
wire _2728_;
wire _2729_;
wire _2730_;
wire _2731_;
wire _2732_;
wire _2733_;
wire _2734_;
wire _2735_;
wire _2736_;
wire _2737_;
wire _2738_;
wire _2739_;
wire _2740_;
wire _2741_;
wire _2742_;
wire _2743_;
wire _2744_;
wire _2745_;
wire _2746_;
wire _2747_;
wire _2748_;
wire _2749_;
wire _2750_;
wire _2751_;
wire _2752_;
wire _2753_;
wire _2754_;
wire _2755_;
wire _2756_;
wire _2757_;
wire _2758_;
wire _2759_;
wire _2760_;
wire _2761_;
wire _2762_;
wire _2763_;
wire _2764_;
wire _2765_;
wire _2766_;
wire _2767_;
wire _2768_;
wire _2769_;
wire _2770_;
wire _2771_;
wire _2772_;
wire _2773_;
wire _2774_;
wire _2775_;
wire _2776_;
wire _2777_;
wire _2778_;
wire _2779_;
wire _2780_;
wire _2781_;
wire _2782_;
wire _2783_;
wire _2784_;
wire _2785_;
wire _2786_;
wire _2787_;
wire _2788_;
wire _2789_;
wire _2790_;
wire _2791_;
wire _2792_;
wire _2793_;
wire _2794_;
wire _2795_;
wire _2796_;
wire _2797_;
wire _2798_;
wire _2799_;
wire _2800_;
wire _2801_;
wire _2802_;
wire _2803_;
wire _2804_;
wire _2805_;
wire _2806_;
wire _2807_;
wire _2808_;
wire _2809_;
wire _2810_;
wire _2811_;
wire _2812_;
wire _2813_;
wire _2814_;
wire _2815_;
wire _2816_;
wire _2817_;
wire _2818_;
wire _2819_;
wire _2820_;
wire _2821_;
wire _2822_;
wire _2823_;
wire _2824_;
wire _2825_;
wire _2826_;
wire _2827_;
wire _2828_;
wire _2829_;
wire _2830_;
wire _2831_;
wire _2832_;
wire _2833_;
wire _2834_;
wire _2835_;
wire _2836_;
wire _2837_;
wire _2838_;
wire _2839_;
wire _2840_;
wire _2841_;
wire _2842_;
wire _2843_;
wire _2844_;
wire _2845_;
wire _2846_;
wire _2847_;
wire _2848_;
wire _2849_;
wire _2850_;
wire _2851_;
wire _2852_;
wire _2853_;
wire _2854_;
wire _2855_;
wire _2856_;
wire _2857_;
wire _2858_;
wire _2859_;
wire _2860_;
wire _2861_;
wire _2862_;
wire _2863_;
wire _2864_;
wire _2865_;
wire _2866_;
wire _2867_;
wire _2868_;
wire _2869_;
wire _2870_;
wire _2871_;
wire _2872_;
wire _2873_;
wire _2874_;
wire _2875_;
wire _2876_;
wire _2877_;
wire _2878_;
wire _2879_;
wire _2880_;
wire _2881_;
wire _2882_;
wire _2883_;
wire _2884_;
wire _2885_;
wire _2886_;
wire _2887_;
wire _2888_;
wire _2889_;
wire _2890_;
wire _2891_;
wire _2892_;
wire _2893_;
wire _2894_;
wire _2895_;
wire _2896_;
wire _2897_;
wire _2898_;
wire _2899_;
wire _2900_;
wire _2901_;
wire _2902_;
wire _2903_;
wire _2904_;
wire _2905_;
wire _2906_;
wire _2907_;
wire _2908_;
wire _2909_;
wire _2910_;
wire _2911_;
wire _2912_;
wire _2913_;
wire _2914_;
wire _2915_;
wire _2916_;
wire _2917_;
wire _2918_;
wire _2919_;
wire _2920_;
wire _2921_;
wire _2922_;
wire _2923_;
wire _2924_;
wire _2925_;
wire _2926_;
wire _2927_;
wire _2928_;
wire _2929_;
wire _2930_;
wire _2931_;
wire _2932_;
wire _2933_;
wire _2934_;
wire _2935_;
wire _2936_;
wire _2937_;
wire _2938_;
wire _2939_;
wire _2940_;
wire _2941_;
wire _2942_;
wire _2943_;
wire _2944_;
wire _2945_;
wire _2946_;
wire _2947_;
wire _2948_;
wire _2949_;
wire _2950_;
wire _2951_;
wire _2952_;
wire _2953_;
wire _2954_;
wire _2955_;
wire _2956_;
wire _2957_;
wire _2958_;
wire _2959_;
wire _2960_;
wire _2961_;
wire _2962_;
wire _2963_;
wire _2964_;
wire _2965_;
wire _2966_;
wire _2967_;
wire _2968_;
wire _2969_;
wire _2970_;
wire _2971_;
wire _2972_;
wire _2973_;
wire _2974_;
wire _2975_;
wire _2976_;
wire _2977_;
wire _2978_;
wire _2979_;
wire _2980_;
wire _2981_;
wire _2982_;
wire _2983_;
wire _2984_;
wire _2985_;
wire _2986_;
wire _2987_;
wire _2988_;
wire _2989_;
wire _2990_;
wire _2991_;
wire _2992_;
wire _2993_;
wire _2994_;
wire _2995_;
wire _2996_;
wire _2997_;
wire _2998_;
wire _2999_;
wire _3000_;
wire _3001_;
wire _3002_;
wire _3003_;
wire _3004_;
wire _3005_;
wire _3006_;
wire _3007_;
wire _3008_;
wire _3009_;
wire _3010_;
wire _3011_;
wire _3012_;
wire _3013_;
wire _3014_;
wire _3015_;
wire _3016_;
wire _3017_;
wire _3018_;
wire _3019_;
wire _3020_;
wire _3021_;
wire _3022_;
wire _3023_;
wire _3024_;
wire _3025_;
wire _3026_;
wire _3027_;
wire _3028_;
wire _3029_;
wire _3030_;
wire _3031_;
wire _3032_;
wire _3033_;
wire _3034_;
wire _3035_;
wire _3036_;
wire _3037_;
wire _3038_;
wire _3039_;
wire _3040_;
wire _3041_;
wire _3042_;
wire _3043_;
wire _3044_;
wire _3045_;
wire _3046_;
wire _3047_;
wire _3048_;
wire _3049_;
wire _3050_;
wire _3051_;
wire _3052_;
wire _3053_;
wire _3054_;
wire _3055_;
wire _3056_;
wire _3057_;
wire _3058_;
wire _3059_;
wire _3060_;
wire _3061_;
wire _3062_;
wire _3063_;
wire _3064_;
wire _3065_;
wire _3066_;
wire _3067_;
wire _3068_;
wire _3069_;
wire _3070_;
wire _3071_;
wire _3072_;
wire _3073_;
wire _3074_;
wire _3075_;
wire _3076_;
wire _3077_;
wire _3078_;
wire _3079_;
wire _3080_;
wire _3081_;
wire _3082_;
wire _3083_;
wire _3084_;
wire _3085_;
wire _3086_;
wire _3087_;
wire _3088_;
wire _3089_;
wire _3090_;
wire _3091_;
wire _3092_;
wire _3093_;
wire _3094_;
wire _3095_;
wire _3096_;
wire _3097_;
wire _3098_;
wire _3099_;
wire _3100_;
wire _3101_;
wire _3102_;
wire _3103_;
wire _3104_;
wire _3105_;
wire _3106_;
wire _3107_;
wire _3108_;
wire _3109_;
wire _3110_;
wire _3111_;
wire _3112_;
wire _3113_;
wire _3114_;
wire _3115_;
wire _3116_;
wire _3117_;
wire _3118_;
wire _3119_;
wire _3120_;
wire _3121_;
wire _3122_;
wire _3123_;
wire _3124_;
wire _3125_;
wire _3126_;
wire _3127_;
wire _3128_;
wire _3129_;
wire _3130_;
wire _3131_;
wire _3132_;
wire _3133_;
wire _3134_;
wire _3135_;
wire _3136_;
wire _3137_;
wire _3138_;
wire _3139_;
wire _3140_;
wire _3141_;
wire _3142_;
wire _3143_;
wire _3144_;
wire _3145_;
wire _3146_;
wire _3147_;
wire _3148_;
wire _3149_;
wire _3150_;
wire _3151_;
wire _3152_;
wire _3153_;
wire _3154_;
wire _3155_;
wire _3156_;
wire _3157_;
wire _3158_;
wire _3159_;
wire _3160_;
wire _3161_;
wire _3162_;
wire _3163_;
wire _3164_;
wire _3165_;
wire _3166_;
wire _3167_;
wire _3168_;
wire _3169_;
wire _3170_;
wire _3171_;
wire _3172_;
wire _3173_;
wire _3174_;
wire _3175_;
wire _3176_;
wire _3177_;
wire _3178_;
wire _3179_;
wire _3180_;
wire _3181_;
wire _3182_;
wire _3183_;
wire _3184_;
wire _3185_;
wire _3186_;
wire _3187_;
wire _3188_;
wire _3189_;
wire _3190_;
wire _3191_;
wire _3192_;
wire _3193_;
wire _3194_;
wire _3195_;
wire _3196_;
wire _3197_;
wire _3198_;
wire _3199_;
wire _3200_;
wire _3201_;
wire _3202_;
wire _3203_;
wire _3204_;
wire _3205_;
wire _3206_;
wire _3207_;
wire _3208_;
wire _3209_;
wire _3210_;
wire _3211_;
wire _3212_;
wire _3213_;
wire _3214_;
wire _3215_;
wire _3216_;
wire _3217_;
wire _3218_;
wire _3219_;
wire _3220_;
wire _3221_;
wire _3222_;
wire _3223_;
wire _3224_;
wire _3225_;
wire _3226_;
wire _3227_;
wire _3228_;
wire _3229_;
wire _3230_;
wire _3231_;
wire _3232_;
wire _3233_;
wire _3234_;
wire _3235_;
wire _3236_;
wire _3237_;
wire _3238_;
wire _3239_;
wire _3240_;
wire _3241_;
wire _3242_;
wire _3243_;
wire _3244_;
wire _3245_;
wire _3246_;
wire _3247_;
wire _3248_;
wire _3249_;
wire _3250_;
wire _3251_;
wire _3252_;
wire _3253_;
wire _3254_;
wire _3255_;
wire _3256_;
wire _3257_;
wire _3258_;
wire _3259_;
wire _3260_;
wire _3261_;
wire _3262_;
wire _3263_;
wire _3264_;
wire _3265_;
wire _3266_;
wire _3267_;
wire _3268_;
wire _3269_;
wire _3270_;
wire _3271_;
wire _3272_;
wire _3273_;
wire _3274_;
wire _3275_;
wire _3276_;
wire _3277_;
wire _3278_;
wire _3279_;
wire _3280_;
wire _3281_;
wire _3282_;
wire _3283_;
wire _3284_;
wire _3285_;
wire _3286_;
wire _3287_;
wire _3288_;
wire _3289_;
wire _3290_;
wire _3291_;
wire _3292_;
wire _3293_;
wire _3294_;
wire _3295_;
wire _3296_;
wire _3297_;
wire _3298_;
wire _3299_;
wire _3300_;
wire _3301_;
wire _3302_;
wire _3303_;
wire _3304_;
wire _3305_;
wire _3306_;
wire _3307_;
wire _3308_;
wire _3309_;
wire _3310_;
wire _3311_;
wire _3312_;
wire _3313_;
wire _3314_;
wire _3315_;
wire _3316_;
wire _3317_;
wire _3318_;
wire _3319_;
wire _3320_;
wire _3321_;
wire _3322_;
wire _3323_;
wire _3324_;
wire _3325_;
wire _3326_;
wire _3327_;
wire _3328_;
wire _3329_;
wire _3330_;
wire _3331_;
wire _3332_;
wire _3333_;
wire _3334_;
wire _3335_;
wire _3336_;
wire _3337_;
wire _3338_;
wire _3339_;
wire _3340_;
wire _3341_;
wire _3342_;
wire _3343_;
wire _3344_;
wire _3345_;
wire _3346_;
wire _3347_;
wire _3348_;
wire _3349_;
wire _3350_;
wire _3351_;
wire _3352_;
wire _3353_;
wire _3354_;
wire _3355_;
wire _3356_;
wire _3357_;
wire _3358_;
wire _3359_;
wire _3360_;
wire _3361_;
wire _3362_;
wire _3363_;
wire _3364_;
wire _3365_;
wire _3366_;
wire _3367_;
wire _3368_;
wire _3369_;
wire _3370_;
wire _3371_;
wire _3372_;
wire _3373_;
wire _3374_;
wire _3375_;
wire _3376_;
wire _3377_;
wire _3378_;
wire _3379_;
wire _3380_;
wire _3381_;
wire _3382_;
wire _3383_;
wire _3384_;
wire _3385_;
wire _3386_;
wire _3387_;
wire _3388_;
wire _3389_;
wire _3390_;
wire _3391_;
wire _3392_;
wire _3393_;
wire _3394_;
wire _3395_;
wire _3396_;
wire _3397_;
wire _3398_;
wire _3399_;
wire _3400_;
wire _3401_;
wire _3402_;
wire _3403_;
wire _3404_;
wire _3405_;
wire _3406_;
wire _3407_;
wire _3408_;
wire _3409_;
wire _3410_;
wire _3411_;
wire _3412_;
wire _3413_;
wire _3414_;
wire _3415_;
wire _3416_;
wire _3417_;
wire _3418_;
wire _3419_;
wire _3420_;
wire _3421_;
wire _3422_;
wire _3423_;
wire _3424_;
wire _3425_;
wire _3426_;
wire _3427_;
wire _3428_;
wire _3429_;
wire _3430_;
wire _3431_;
wire _3432_;
wire _3433_;
wire _3434_;
wire _3435_;
wire _3436_;
wire _3437_;
wire _3438_;
wire _3439_;
wire _3440_;
wire _3441_;
wire _3442_;
wire _3443_;
wire _3444_;
wire _3445_;
wire _3446_;
wire _3447_;
wire _3448_;
wire _3449_;
wire _3450_;
wire _3451_;
wire _3452_;
wire _3453_;
wire _3454_;
wire _3455_;
wire _3456_;
wire _3457_;
wire _3458_;
wire _3459_;
wire _3460_;
wire _3461_;
wire _3462_;
wire _3463_;
wire _3464_;
wire _3465_;
wire _3466_;
wire _3467_;
wire _3468_;
wire _3469_;
wire _3470_;
wire _3471_;
wire _3472_;
wire _3473_;
wire _3474_;
wire _3475_;
wire _3476_;
wire _3477_;
wire _3478_;
wire _3479_;
wire _3480_;
wire _3481_;
wire _3482_;
wire _3483_;
wire _3484_;
wire _3485_;
wire _3486_;
wire _3487_;
wire _3488_;
wire _3489_;
wire _3490_;
wire _3491_;
wire _3492_;
wire _3493_;
wire _3494_;
wire _3495_;
wire _3496_;
wire _3497_;
wire _3498_;
wire _3499_;
wire _3500_;
wire _3501_;
wire _3502_;
wire _3503_;
wire _3504_;
wire _3505_;
wire _3506_;
wire _3507_;
wire _3508_;
wire _3509_;
wire _3510_;
wire _3511_;
wire _3512_;
wire _3513_;
wire _3514_;
wire _3515_;
wire _3516_;
wire _3517_;
wire _3518_;
wire _3519_;
wire _3520_;
wire _3521_;
wire _3522_;
wire _3523_;
wire _3524_;
wire _3525_;
wire _3526_;
wire _3527_;
wire _3528_;
wire _3529_;
wire _3530_;
wire _3531_;
wire _3532_;
wire _3533_;
wire _3534_;
wire _3535_;
wire _3536_;
wire _3537_;
wire _3538_;
wire _3539_;
wire _3540_;
wire _3541_;
wire _3542_;
wire _3543_;
wire _3544_;
wire _3545_;
wire _3546_;
wire _3547_;
wire _3548_;
wire _3549_;
wire _3550_;
wire _3551_;
wire _3552_;
wire _3553_;
wire _3554_;
wire _3555_;
wire _3556_;
wire _3557_;
wire _3558_;
wire _3559_;
wire _3560_;
wire _3561_;
wire _3562_;
wire _3563_;
wire _3564_;
wire _3565_;
wire _3566_;
wire _3567_;
wire _3568_;
wire _3569_;
wire _3570_;
wire _3571_;
wire _3572_;
wire _3573_;
wire _3574_;
wire _3575_;
wire _3576_;
wire _3577_;
wire _3578_;
wire _3579_;
wire _3580_;
wire _3581_;
wire _3582_;
wire _3583_;
wire _3584_;
wire _3585_;
wire _3586_;
wire _3587_;
wire _3588_;
wire _3589_;
wire _3590_;
wire _3591_;
wire _3592_;
wire _3593_;
wire _3594_;
wire _3595_;
wire _3596_;
wire _3597_;
wire _3598_;
wire _3599_;
wire _3600_;
wire _3601_;
wire _3602_;
wire _3603_;
wire _3604_;
wire _3605_;
wire _3606_;
wire _3607_;
wire _3608_;
wire _3609_;
wire _3610_;
wire _3611_;
wire _3612_;
wire _3613_;
wire _3614_;
wire _3615_;
wire _3616_;
wire _3617_;
wire _3618_;
wire _3619_;
wire _3620_;
wire _3621_;
wire _3622_;
wire _3623_;
wire _3624_;
wire _3625_;
wire _3626_;
wire _3627_;
wire _3628_;
wire _3629_;
wire _3630_;
wire _3631_;
wire _3632_;
wire _3633_;
wire _3634_;
wire _3635_;
wire _3636_;
wire _3637_;
wire _3638_;
wire _3639_;
wire _3640_;
wire _3641_;
wire _3642_;
wire _3643_;
wire _3644_;
wire _3645_;
wire _3646_;
wire _3647_;
wire _3648_;
wire _3649_;
wire _3650_;
wire _3651_;
wire _3652_;
wire _3653_;
wire _3654_;
wire _3655_;
wire _3656_;
wire _3657_;
wire _3658_;
wire _3659_;
wire _3660_;
wire _3661_;
wire _3662_;
wire _3663_;
wire _3664_;
wire _3665_;
wire _3666_;
wire _3667_;
wire _3668_;
wire _3669_;
wire _3670_;
wire _3671_;
wire _3672_;
wire _3673_;
wire _3674_;
wire _3675_;
wire _3676_;
wire _3677_;
wire _3678_;
wire _3679_;
wire _3680_;
wire _3681_;
wire _3682_;
wire _3683_;
wire _3684_;
wire _3685_;
wire _3686_;
wire _3687_;
wire _3688_;
wire _3689_;
wire _3690_;
wire _3691_;
wire _3692_;
wire _3693_;
wire _3694_;
wire _3695_;
wire _3696_;
wire _3697_;
wire _3698_;
wire _3699_;
wire _3700_;
wire _3701_;
wire _3702_;
wire _3703_;
wire _3704_;
wire _3705_;
wire _3706_;
wire _3707_;
wire _3708_;
wire _3709_;
wire _3710_;
wire _3711_;
wire _3712_;
wire _3713_;
wire _3714_;
wire _3715_;
wire _3716_;
wire _3717_;
wire _3718_;
wire _3719_;
wire _3720_;
wire _3721_;
wire _3722_;
wire _3723_;
wire _3724_;
wire _3725_;
wire _3726_;
wire _3727_;
wire _3728_;
wire _3729_;
wire _3730_;
wire _3731_;
wire _3732_;
wire _3733_;
wire _3734_;
wire _3735_;
wire _3736_;
wire _3737_;
wire _3738_;
wire _3739_;
wire _3740_;
wire _3741_;
wire _3742_;
wire _3743_;
wire _3744_;
wire _3745_;
wire _3746_;
wire _3747_;
wire _3748_;
wire _3749_;
wire _3750_;
wire _3751_;
wire _3752_;
wire _3753_;
wire _3754_;
wire _3755_;
wire _3756_;
wire _3757_;
wire _3758_;
wire _3759_;
wire _3760_;
wire _3761_;
wire _3762_;
wire _3763_;
wire _3764_;
wire _3765_;
wire _3766_;
wire _3767_;
wire _3768_;
wire _3769_;
wire _3770_;
wire _3771_;
wire _3772_;
wire _3773_;
wire _3774_;
wire _3775_;
wire _3776_;
wire _3777_;
wire _3778_;
wire _3779_;
wire _3780_;
wire _3781_;
wire _3782_;
wire _3783_;
wire _3784_;
wire _3785_;
wire _3786_;
wire _3787_;
wire _3788_;
wire _3789_;
wire _3790_;
wire _3791_;
wire _3792_;
wire _3793_;
wire _3794_;
wire _3795_;
wire _3796_;
wire _3797_;
wire _3798_;
wire _3799_;
wire _3800_;
wire _3801_;
wire _3802_;
wire _3803_;
wire _3804_;
wire _3805_;
wire _3806_;
wire _3807_;
wire _3808_;
wire _3809_;
wire _3810_;
wire _3811_;
wire _3812_;
wire _3813_;
wire _3814_;
wire _3815_;
wire _3816_;
wire _3817_;
wire _3818_;
wire _3819_;
wire _3820_;
wire _3821_;
wire _3822_;
wire _3823_;
wire _3824_;
wire _3825_;
wire _3826_;
wire _3827_;
wire _3828_;
wire _3829_;
wire _3830_;
wire _3831_;
wire _3832_;
wire _3833_;
wire _3834_;
wire _3835_;
wire _3836_;
wire _3837_;
wire _3838_;
wire _3839_;
wire _3840_;
wire _3841_;
wire _3842_;
wire _3843_;
wire _3844_;
wire _3845_;
wire _3846_;
wire _3847_;
wire _3848_;
wire _3849_;
wire _3850_;
wire _3851_;
wire _3852_;
wire _3853_;
wire _3854_;
wire _3855_;
wire _3856_;
wire _3857_;
wire _3858_;
wire _3859_;
wire _3860_;
wire _3861_;
wire _3862_;
wire _3863_;
wire _3864_;
wire _3865_;
wire _3866_;
wire _3867_;
wire _3868_;
wire _3869_;
wire _3870_;
wire _3871_;
wire _3872_;
wire _3873_;
wire _3874_;
wire _3875_;
wire _3876_;
wire _3877_;
wire _3878_;
wire _3879_;
wire _3880_;
wire _3881_;
wire _3882_;
wire _3883_;
wire _3884_;
wire _3885_;
wire _3886_;
wire _3887_;
wire _3888_;
wire _3889_;
wire _3890_;
wire _3891_;
wire _3892_;
wire _3893_;
wire _3894_;
wire _3895_;
wire _3896_;
wire _3897_;
wire _3898_;
wire _3899_;
wire _3900_;
wire _3901_;
wire _3902_;
wire _3903_;
wire _3904_;
wire _3905_;
wire _3906_;
wire _3907_;
wire _3908_;
wire _3909_;
wire _3910_;
wire _3911_;
wire _3912_;
wire _3913_;
wire _3914_;
wire _3915_;
wire _3916_;
wire _3917_;
wire _3918_;
wire _3919_;
wire _3920_;
wire _3921_;
wire _3922_;
wire _3923_;
wire _3924_;
wire _3925_;
wire _3926_;
wire _3927_;
wire _3928_;
wire _3929_;
wire _3930_;
wire _3931_;
wire _3932_;
wire _3933_;
wire _3934_;
wire _3935_;
wire _3936_;
wire _3937_;
wire _3938_;
wire _3939_;
wire _3940_;
wire _3941_;
wire _3942_;
wire _3943_;
wire _3944_;
wire _3945_;
wire _3946_;
wire _3947_;
wire _3948_;
wire _3949_;
wire _3950_;
wire _3951_;
wire _3952_;
wire _3953_;
wire _3954_;
wire _3955_;
wire _3956_;
wire _3957_;
wire _3958_;
wire _3959_;
wire _3960_;
wire _3961_;
wire _3962_;
wire _3963_;
wire _3964_;
wire _3965_;
wire _3966_;
wire _3967_;
wire _3968_;
wire _3969_;
wire _3970_;
wire _3971_;
wire _3972_;
wire _3973_;
wire _3974_;
wire _3975_;
wire _3976_;
wire _3977_;
wire _3978_;
wire _3979_;
wire _3980_;
wire _3981_;
wire _3982_;
wire _3983_;
wire _3984_;
wire _3985_;
wire _3986_;
wire _3987_;
wire _3988_;
wire _3989_;
wire _3990_;
wire _3991_;
wire _3992_;
wire _3993_;
wire _3994_;
wire _3995_;
wire _3996_;
wire _3997_;
wire _3998_;
wire _3999_;
wire _4000_;
wire _4001_;
wire _4002_;
wire _4003_;
wire _4004_;
wire _4005_;
wire _4006_;
wire _4007_;
wire _4008_;
wire _4009_;
wire _4010_;
wire _4011_;
wire _4012_;
wire _4013_;
wire _4014_;
wire _4015_;
wire _4016_;
wire _4017_;
wire _4018_;
wire _4019_;
wire _4020_;
wire _4021_;
wire _4022_;
wire _4023_;
wire _4024_;
wire _4025_;
wire _4026_;
wire _4027_;
wire _4028_;
wire _4029_;
wire _4030_;
wire _4031_;
wire _4032_;
wire _4033_;
wire _4034_;
wire _4035_;
wire _4036_;
wire _4037_;
wire _4038_;
wire _4039_;
wire _4040_;
wire _4041_;
wire _4042_;
wire _4043_;
wire _4044_;
wire _4045_;
wire _4046_;
wire _4047_;
wire _4048_;
wire _4049_;
wire _4050_;
wire _4051_;
wire _4052_;
wire _4053_;
wire _4054_;
wire _4055_;
wire _4056_;
wire _4057_;
wire _4058_;
wire _4059_;
wire _4060_;
wire _4061_;
wire _4062_;
wire _4063_;
wire _4064_;
wire _4065_;
wire _4066_;
wire _4067_;
wire _4068_;
wire _4069_;
wire _4070_;
wire _4071_;
wire _4072_;
wire _4073_;
wire _4074_;
wire _4075_;
wire _4076_;
wire _4077_;
wire _4078_;
wire _4079_;
wire _4080_;
wire _4081_;
wire _4082_;
wire _4083_;
wire _4084_;
wire _4085_;
wire _4086_;
wire _4087_;
wire _4088_;
wire _4089_;
wire _4090_;
wire _4091_;
wire _4092_;
wire _4093_;
wire _4094_;
wire _4095_;
wire _4096_;
wire _4097_;
wire _4098_;
wire _4099_;
wire _4100_;
wire _4101_;
wire _4102_;
wire _4103_;
wire _4104_;
wire _4105_;
wire _4106_;
wire _4107_;
wire _4108_;
wire _4109_;
wire _4110_;
wire _4111_;
wire _4112_;
wire _4113_;
wire _4114_;
wire _4115_;
wire _4116_;
wire _4117_;
wire _4118_;
wire _4119_;
wire _4120_;
wire _4121_;
wire _4122_;
wire _4123_;
wire _4124_;
wire _4125_;
wire _4126_;
wire _4127_;
wire _4128_;
wire _4129_;
wire _4130_;
wire _4131_;
wire _4132_;
wire _4133_;
wire _4134_;
wire _4135_;
wire _4136_;
wire _4137_;
wire _4138_;
wire _4139_;
wire _4140_;
wire _4141_;
wire _4142_;
wire _4143_;
wire _4144_;
wire _4145_;
wire _4146_;
wire _4147_;
wire _4148_;
wire _4149_;
wire _4150_;
wire _4151_;
wire _4152_;
wire _4153_;
wire _4154_;
wire _4155_;
wire _4156_;
wire _4157_;
wire _4158_;
wire _4159_;
wire _4160_;
wire _4161_;
wire _4162_;
wire _4163_;
wire _4164_;
wire _4165_;
wire _4166_;
wire _4167_;
wire _4168_;
wire _4169_;
wire _4170_;
wire _4171_;
wire _4172_;
wire _4173_;
wire _4174_;
wire _4175_;
wire _4176_;
wire _4177_;
wire _4178_;
wire _4179_;
wire _4180_;
wire _4181_;
wire _4182_;
wire _4183_;
wire _4184_;
wire _4185_;
wire _4186_;
wire _4187_;
wire _4188_;
wire _4189_;
wire _4190_;
wire _4191_;
wire _4192_;
wire _4193_;
wire _4194_;
wire _4195_;
wire _4196_;
wire _4197_;
wire _4198_;
wire _4199_;
wire _4200_;
wire _4201_;
wire _4202_;
wire _4203_;
wire _4204_;
wire _4205_;
wire _4206_;
wire _4207_;
wire _4208_;
wire _4209_;
wire _4210_;
wire _4211_;
wire _4212_;
wire _4213_;
wire _4214_;
wire _4215_;
wire _4216_;
wire _4217_;
wire _4218_;
wire _4219_;
wire _4220_;
wire _4221_;
wire _4222_;
wire _4223_;
wire _4224_;
wire _4225_;
wire _4226_;
wire _4227_;
wire _4228_;
wire _4229_;
wire _4230_;
wire _4231_;
wire _4232_;
wire _4233_;
wire _4234_;
wire _4235_;
wire _4236_;
wire _4237_;
wire _4238_;
wire _4239_;
wire _4240_;
wire _4241_;
wire _4242_;
wire _4243_;
wire _4244_;
wire _4245_;
wire _4246_;
wire _4247_;
wire _4248_;
wire _4249_;
wire _4250_;
wire _4251_;
wire _4252_;
wire _4253_;
wire _4254_;
wire _4255_;
wire _4256_;
wire _4257_;
wire _4258_;
wire _4259_;
wire _4260_;
wire _4261_;
wire _4262_;
wire _4263_;
wire _4264_;
wire _4265_;
wire _4266_;
wire _4267_;
wire _4268_;
wire _4269_;
wire _4270_;
wire _4271_;
wire _4272_;
wire _4273_;
wire _4274_;
wire _4275_;
wire _4276_;
wire _4277_;
wire _4278_;
wire _4279_;
wire _4280_;
wire _4281_;
wire _4282_;
wire _4283_;
wire _4284_;
wire _4285_;
wire _4286_;
wire _4287_;
wire _4288_;
wire _4289_;
wire _4290_;
wire _4291_;
wire _4292_;
wire _4293_;
wire _4294_;
wire _4295_;
wire _4296_;
wire _4297_;
wire _4298_;
wire _4299_;
wire _4300_;
wire _4301_;
wire _4302_;
wire _4303_;
wire _4304_;
wire _4305_;
wire _4306_;
wire _4307_;
wire _4308_;
wire _4309_;
wire _4310_;
wire _4311_;
wire _4312_;
wire _4313_;
wire _4314_;
wire _4315_;
wire _4316_;
wire _4317_;
wire _4318_;
wire _4319_;
wire _4320_;
wire _4321_;
wire _4322_;
wire _4323_;
wire _4324_;
wire _4325_;
wire _4326_;
wire _4327_;
wire _4328_;
wire _4329_;
wire _4330_;
wire _4331_;
wire _4332_;
wire _4333_;
wire _4334_;
wire _4335_;
wire _4336_;
wire _4337_;
wire _4338_;
wire _4339_;
wire _4340_;
wire _4341_;
wire _4342_;
wire _4343_;
wire _4344_;
wire _4345_;
wire _4346_;
wire _4347_;
wire _4348_;
wire _4349_;
wire _4350_;
wire _4351_;
wire _4352_;
wire _4353_;
wire _4354_;
wire _4355_;
wire _4356_;
wire _4357_;
wire _4358_;
wire _4359_;
wire _4360_;
wire _4361_;
wire _4362_;
wire _4363_;
wire _4364_;
wire _4365_;
wire _4366_;
wire _4367_;
wire _4368_;
wire _4369_;
wire _4370_;
wire _4371_;
wire _4372_;
wire _4373_;
wire _4374_;
wire _4375_;
wire _4376_;
wire _4377_;
wire _4378_;
wire _4379_;
wire _4380_;
wire _4381_;
wire _4382_;
wire _4383_;
wire _4384_;
wire _4385_;
wire _4386_;
wire _4387_;
wire _4388_;
wire _4389_;
wire _4390_;
wire _4391_;
wire _4392_;
wire _4393_;
wire _4394_;
wire _4395_;
wire _4396_;
wire _4397_;
wire _4398_;
wire _4399_;
wire _4400_;
wire _4401_;
wire _4402_;
wire _4403_;
wire _4404_;
wire _4405_;
wire _4406_;
wire _4407_;
wire _4408_;
wire _4409_;
wire _4410_;
wire _4411_;
wire _4412_;
wire _4413_;
wire _4414_;
wire _4415_;
wire _4416_;
wire _4417_;
wire _4418_;
wire _4419_;
wire _4420_;
wire _4421_;
wire _4422_;
wire _4423_;
wire _4424_;
wire _4425_;
wire _4426_;
wire _4427_;
wire _4428_;
wire _4429_;
wire _4430_;
wire _4431_;
wire _4432_;
wire _4433_;
wire _4434_;
wire _4435_;
wire _4436_;
wire _4437_;
wire _4438_;
wire _4439_;
wire _4440_;
wire _4441_;
wire _4442_;
wire _4443_;
wire _4444_;
wire _4445_;
wire _4446_;
wire _4447_;
wire _4448_;
wire _4449_;
wire _4450_;
wire _4451_;
wire _4452_;
wire _4453_;
wire _4454_;
wire _4455_;
wire _4456_;
wire _4457_;
wire _4458_;
wire _4459_;
wire _4460_;
wire _4461_;
wire _4462_;
wire _4463_;
wire _4464_;
wire _4465_;
wire _4466_;
wire _4467_;
wire _4468_;
wire _4469_;
wire _4470_;
wire _4471_;
wire _4472_;
wire _4473_;
wire _4474_;
wire _4475_;
wire _4476_;
wire _4477_;
wire _4478_;
wire _4479_;
wire _4480_;
wire _4481_;
wire _4482_;
wire _4483_;
wire _4484_;
wire _4485_;
wire _4486_;
wire _4487_;
wire _4488_;
wire _4489_;
wire _4490_;
wire _4491_;
wire _4492_;
wire _4493_;
wire _4494_;
wire _4495_;
wire _4496_;
wire _4497_;
wire _4498_;
wire _4499_;
wire _4500_;
wire _4501_;
wire _4502_;
wire _4503_;
wire _4504_;
wire _4505_;
wire _4506_;
wire _4507_;
wire _4508_;
wire _4509_;
wire _4510_;
wire _4511_;
wire _4512_;
wire _4513_;
wire _4514_;
wire _4515_;
wire _4516_;
wire _4517_;
wire _4518_;
wire _4519_;
wire _4520_;
wire _4521_;
wire _4522_;
wire _4523_;
wire _4524_;
wire _4525_;
wire _4526_;
wire _4527_;
wire _4528_;
wire _4529_;
wire _4530_;
wire _4531_;
wire _4532_;
wire _4533_;
wire _4534_;
wire _4535_;
wire _4536_;
wire _4537_;
wire _4538_;
wire _4539_;
wire _4540_;
wire _4541_;
wire _4542_;
wire _4543_;
wire _4544_;
wire _4545_;
wire _4546_;
wire _4547_;
wire _4548_;
wire _4549_;
wire _4550_;
wire _4551_;
wire _4552_;
wire _4553_;
wire _4554_;
wire _4555_;
wire _4556_;
wire _4557_;
wire _4558_;
wire _4559_;
wire _4560_;
wire _4561_;
wire _4562_;
wire _4563_;
wire _4564_;
wire _4565_;
wire _4566_;
wire _4567_;
wire _4568_;
wire _4569_;
wire _4570_;
wire _4571_;
wire _4572_;
wire _4573_;
wire _4574_;
wire _4575_;
wire _4576_;
wire _4577_;
wire _4578_;
wire _4579_;
wire _4580_;
wire _4581_;
wire _4582_;
wire _4583_;
wire _4584_;
wire _4585_;
wire _4586_;
wire _4587_;
wire _4588_;
wire _4589_;
wire _4590_;
wire _4591_;
wire _4592_;
wire _4593_;
wire _4594_;
wire _4595_;
wire _4596_;
wire _4597_;
wire _4598_;
wire _4599_;
wire _4600_;
wire _4601_;
wire _4602_;
wire _4603_;
wire _4604_;
wire _4605_;
wire _4606_;
wire _4607_;
wire _4608_;
wire _4609_;
wire _4610_;
wire _4611_;
wire _4612_;
wire _4613_;
wire _4614_;
wire _4615_;
wire _4616_;
wire _4617_;
wire _4618_;
wire _4619_;
wire _4620_;
wire _4621_;
wire _4622_;
wire _4623_;
wire _4624_;
wire _4625_;
wire _4626_;
wire _4627_;
wire _4628_;
wire _4629_;
wire _4630_;
wire _4631_;
wire _4632_;
wire _4633_;
wire _4634_;
wire _4635_;
wire _4636_;
wire _4637_;
wire _4638_;
wire _4639_;
wire _4640_;
wire _4641_;
wire _4642_;
wire _4643_;
wire _4644_;
wire _4645_;
wire _4646_;
wire _4647_;
wire _4648_;
wire _4649_;
wire _4650_;
wire _4651_;
wire _4652_;
wire _4653_;
wire _4654_;
wire _4655_;
wire _4656_;
wire _4657_;
wire _4658_;
wire _4659_;
wire _4660_;
wire _4661_;
wire _4662_;
wire _4663_;
wire _4664_;
wire _4665_;
wire _4666_;
wire _4667_;
wire _4668_;
wire _4669_;
wire _4670_;
wire _4671_;
wire _4672_;
wire _4673_;
wire _4674_;
wire _4675_;
wire _4676_;
wire _4677_;
wire _4678_;
wire _4679_;
wire _4680_;
wire _4681_;
wire _4682_;
wire _4683_;
wire _4684_;
wire _4685_;
wire _4686_;
wire _4687_;
wire _4688_;
wire _4689_;
wire _4690_;
wire _4691_;
wire _4692_;
wire _4693_;
wire _4694_;
wire _4695_;
wire _4696_;
wire _4697_;
wire _4698_;
wire _4699_;
wire _4700_;
wire _4701_;
wire _4702_;
wire _4703_;
wire _4704_;
wire _4705_;
wire _4706_;
wire _4707_;
wire _4708_;
wire _4709_;
wire _4710_;
wire _4711_;
wire _4712_;
wire _4713_;
wire _4714_;
wire _4715_;
wire _4716_;
wire _4717_;
wire _4718_;
wire _4719_;
wire _4720_;
wire _4721_;
wire _4722_;
wire _4723_;
wire _4724_;
wire _4725_;
wire _4726_;
wire _4727_;
wire _4728_;
wire _4729_;
wire _4730_;
wire _4731_;
wire _4732_;
wire _4733_;
wire _4734_;
wire _4735_;
wire _4736_;
wire _4737_;
wire _4738_;
wire _4739_;
wire _4740_;
wire _4741_;
wire _4742_;
wire _4743_;
wire _4744_;
wire _4745_;
wire _4746_;
wire _4747_;
wire _4748_;
wire _4749_;
wire _4750_;
wire _4751_;
wire _4752_;
wire _4753_;
wire _4754_;
wire _4755_;
wire _4756_;
wire _4757_;
wire _4758_;
wire _4759_;
wire _4760_;
wire _4761_;
wire _4762_;
wire _4763_;
wire _4764_;
wire _4765_;
wire _4766_;
wire _4767_;
wire _4768_;
wire _4769_;
wire _4770_;
wire _4771_;
wire _4772_;
wire _4773_;
wire _4774_;
wire _4775_;
wire _4776_;
wire _4777_;
wire _4778_;
wire _4779_;
wire _4780_;
wire _4781_;
wire _4782_;
wire _4783_;
wire _4784_;
wire _4785_;
wire _4786_;
wire _4787_;
wire _4788_;
wire _4789_;
wire _4790_;
wire _4791_;
wire _4792_;
wire _4793_;
wire _4794_;
wire _4795_;
wire _4796_;
wire _4797_;
wire _4798_;
wire _4799_;
wire _4800_;
wire _4801_;
wire _4802_;
wire _4803_;
wire _4804_;
wire _4805_;
wire _4806_;
wire _4807_;
wire _4808_;
wire _4809_;
wire _4810_;
wire _4811_;
wire _4812_;
wire _4813_;
wire _4814_;
wire _4815_;
wire _4816_;
wire _4817_;
wire _4818_;
wire _4819_;
wire _4820_;
wire _4821_;
wire _4822_;
wire _4823_;
wire _4824_;
wire _4825_;
wire _4826_;
wire _4827_;
wire _4828_;
wire _4829_;
wire _4830_;
wire _4831_;
wire _4832_;
wire _4833_;
wire _4834_;
wire _4835_;
wire _4836_;
wire _4837_;
wire _4838_;
wire _4839_;
wire _4840_;
wire _4841_;
wire _4842_;
wire _4843_;
wire _4844_;
wire _4845_;
wire _4846_;
wire _4847_;
wire _4848_;
wire _4849_;
wire _4850_;
wire _4851_;
wire _4852_;
wire _4853_;
wire _4854_;
wire _4855_;
wire _4856_;
wire _4857_;
wire _4858_;
wire _4859_;
wire _4860_;
wire _4861_;
wire _4862_;
wire _4863_;
wire _4864_;
wire _4865_;
wire _4866_;
wire _4867_;
wire _4868_;
wire _4869_;
wire _4870_;
wire _4871_;
wire _4872_;
wire _4873_;
wire _4874_;
wire _4875_;
wire _4876_;
wire _4877_;
wire _4878_;
wire _4879_;
wire _4880_;
wire _4881_;
wire _4882_;
wire _4883_;
wire _4884_;
wire _4885_;
wire _4886_;
wire _4887_;
wire _4888_;
wire _4889_;
wire _4890_;
wire _4891_;
wire _4892_;
wire _4893_;
wire _4894_;
wire _4895_;
wire _4896_;
wire _4897_;
wire _4898_;
wire _4899_;
wire _4900_;
wire _4901_;
wire _4902_;
wire _4903_;
wire _4904_;
wire _4905_;
wire _4906_;
wire _4907_;
wire _4908_;
wire _4909_;
wire _4910_;
wire _4911_;
wire _4912_;
wire _4913_;
wire _4914_;
wire _4915_;
wire _4916_;
wire _4917_;
wire _4918_;
wire _4919_;
wire _4920_;
wire _4921_;
wire _4922_;
wire _4923_;
wire _4924_;
wire _4925_;
wire _4926_;
wire _4927_;
wire _4928_;
wire _4929_;
wire _4930_;
wire _4931_;
wire _4932_;
wire _4933_;
wire _4934_;
wire _4935_;
wire _4936_;
wire _4937_;
wire _4938_;
wire _4939_;
wire _4940_;
wire _4941_;
wire _4942_;
wire _4943_;
wire _4944_;
wire _4945_;
wire _4946_;
wire _4947_;
wire _4948_;
wire _4949_;
wire _4950_;
wire _4951_;
wire _4952_;
wire _4953_;
wire _4954_;
wire _4955_;
wire _4956_;
wire _4957_;
wire _4958_;
wire _4959_;
wire _4960_;
wire _4961_;
wire _4962_;
wire _4963_;
wire _4964_;
wire _4965_;
wire _4966_;
wire _4967_;
wire _4968_;
wire _4969_;
wire _4970_;
wire _4971_;
wire _4972_;
wire _4973_;
wire _4974_;
wire _4975_;
wire _4976_;
wire _4977_;
wire _4978_;
wire _4979_;
wire _4980_;
wire _4981_;
wire _4982_;
wire _4983_;
wire _4984_;
wire _4985_;
wire _4986_;
wire _4987_;
wire _4988_;
wire _4989_;
wire _4990_;
wire _4991_;
wire _4992_;
wire _4993_;
wire _4994_;
wire _4995_;
wire _4996_;
wire _4997_;
wire _4998_;
wire _4999_;
wire _5000_;
wire _5001_;
wire _5002_;
wire _5003_;
wire _5004_;
wire _5005_;
wire _5006_;
wire _5007_;
wire _5008_;
wire _5009_;
wire _5010_;
wire _5011_;
wire _5012_;
wire _5013_;
wire _5014_;
wire _5015_;
wire _5016_;
wire _5017_;
wire _5018_;
wire _5019_;
wire _5020_;
wire _5021_;
wire _5022_;
wire _5023_;
wire _5024_;
wire _5025_;
wire _5026_;
wire _5027_;
wire _5028_;
wire _5029_;
wire _5030_;
wire _5031_;
wire _5032_;
wire _5033_;
wire _5034_;
wire _5035_;
wire _5036_;
wire _5037_;
wire _5038_;
wire _5039_;
wire _5040_;
wire _5041_;
wire _5042_;
wire _5043_;
wire _5044_;
wire _5045_;
wire _5046_;
wire _5047_;
wire _5048_;
wire _5049_;
wire _5050_;
wire _5051_;
wire _5052_;
wire _5053_;
wire _5054_;
wire _5055_;
wire _5056_;
wire _5057_;
wire _5058_;
wire _5059_;
wire _5060_;
wire _5061_;
wire _5062_;
wire _5063_;
wire _5064_;
wire _5065_;
wire _5066_;
wire _5067_;
wire _5068_;
wire _5069_;
wire _5070_;
wire _5071_;
wire _5072_;
wire _5073_;
wire _5074_;
wire _5075_;
wire _5076_;
wire _5077_;
wire _5078_;
wire _5079_;
wire _5080_;
wire _5081_;
wire _5082_;
wire _5083_;
wire _5084_;
wire _5085_;
wire _5086_;
wire _5087_;
wire _5088_;
wire _5089_;
wire _5090_;
wire _5091_;
wire _5092_;
wire _5093_;
wire _5094_;
wire _5095_;
wire _5096_;
wire _5097_;
wire _5098_;
wire _5099_;
wire _5100_;
wire _5101_;
wire _5102_;
wire _5103_;
wire _5104_;
wire _5105_;
wire _5106_;
wire _5107_;
wire _5108_;
wire _5109_;
wire _5110_;
wire _5111_;
wire _5112_;
wire _5113_;
wire _5114_;
wire _5115_;
wire _5116_;
wire _5117_;
wire _5118_;
wire _5119_;
wire _5120_;
wire _5121_;
wire _5122_;
wire _5123_;
wire _5124_;
wire _5125_;
wire _5126_;
wire _5127_;
wire _5128_;
wire _5129_;
wire _5130_;
wire _5131_;
wire _5132_;
wire _5133_;
wire _5134_;
wire _5135_;
wire _5136_;
wire _5137_;
wire _5138_;
wire _5139_;
wire _5140_;
wire _5141_;
wire _5142_;
wire _5143_;
wire _5144_;
wire _5145_;
wire _5146_;
wire _5147_;
wire _5148_;
wire _5149_;
wire _5150_;
wire _5151_;
wire _5152_;
wire _5153_;
wire _5154_;
wire _5155_;
wire _5156_;
wire _5157_;
wire _5158_;
wire _5159_;
wire _5160_;
wire _5161_;
wire _5162_;
wire _5163_;
wire _5164_;
wire _5165_;
wire _5166_;
wire _5167_;
wire _5168_;
wire _5169_;
wire _5170_;
wire _5171_;
wire _5172_;
wire _5173_;
wire _5174_;
wire _5175_;
wire _5176_;
wire _5177_;
wire _5178_;
wire _5179_;
wire _5180_;
wire _5181_;
wire _5182_;
wire _5183_;
wire _5184_;
wire _5185_;
wire _5186_;
wire _5187_;
wire _5188_;
wire _5189_;
wire _5190_;
wire _5191_;
wire _5192_;
wire _5193_;
wire _5194_;
wire _5195_;
wire _5196_;
wire _5197_;
wire _5198_;
wire _5199_;
wire _5200_;
wire _5201_;
wire _5202_;
wire _5203_;
wire _5204_;
wire _5205_;
wire _5206_;
wire _5207_;
wire _5208_;
wire _5209_;
wire _5210_;
wire _5211_;
wire _5212_;
wire _5213_;
wire _5214_;
wire _5215_;
wire _5216_;
wire _5217_;
wire _5218_;
wire _5219_;
wire _5220_;
wire _5221_;
wire _5222_;
wire _5223_;
wire _5224_;
wire _5225_;
wire _5226_;
wire _5227_;
wire _5228_;
wire _5229_;
wire _5230_;
wire _5231_;
wire _5232_;
wire _5233_;
wire _5234_;
wire _5235_;
wire _5236_;
wire _5237_;
wire _5238_;
wire _5239_;
wire _5240_;
wire _5241_;
wire _5242_;
wire _5243_;
wire _5244_;
wire _5245_;
wire _5246_;
wire _5247_;
wire _5248_;
wire _5249_;
wire _5250_;
wire _5251_;
wire _5252_;
wire _5253_;
wire _5254_;
wire _5255_;
wire _5256_;
wire _5257_;
wire _5258_;
wire _5259_;
wire _5260_;
wire _5261_;
wire _5262_;
wire _5263_;
wire _5264_;
wire _5265_;
wire _5266_;
wire _5267_;
wire _5268_;
wire _5269_;
wire _5270_;
wire _5271_;
wire _5272_;
wire _5273_;
wire _5274_;
wire _5275_;
wire _5276_;
wire _5277_;
wire _5278_;
wire _5279_;
wire _5280_;
wire _5281_;
wire _5282_;
wire _5283_;
wire _5284_;
wire _5285_;
wire _5286_;
wire _5287_;
wire _5288_;
wire _5289_;
wire _5290_;
wire _5291_;
wire _5292_;
wire _5293_;
wire _5294_;
wire _5295_;
wire _5296_;
wire _5297_;
wire _5298_;
wire _5299_;
wire _5300_;
wire _5301_;
wire _5302_;
wire _5303_;
wire _5304_;
wire _5305_;
wire _5306_;
wire _5307_;
wire _5308_;
wire _5309_;
wire _5310_;
wire _5311_;
wire _5312_;
wire _5313_;
wire _5314_;
wire _5315_;
wire _5316_;
wire _5317_;
wire _5318_;
wire _5319_;
wire _5320_;
wire _5321_;
wire _5322_;
wire _5323_;
wire _5324_;
wire _5325_;
wire _5326_;
wire _5327_;
wire _5328_;
wire _5329_;
wire _5330_;
wire _5331_;
wire _5332_;
wire _5333_;
wire _5334_;
wire _5335_;
wire _5336_;
wire _5337_;
wire _5338_;
wire _5339_;
wire _5340_;
wire _5341_;
wire _5342_;
wire _5343_;
wire _5344_;
wire _5345_;
wire _5346_;
wire _5347_;
wire _5348_;
wire _5349_;
wire _5350_;
wire _5351_;
wire _5352_;
wire _5353_;
wire _5354_;
wire _5355_;
wire _5356_;
wire _5357_;
wire _5358_;
wire _5359_;
wire _5360_;
wire _5361_;
wire _5362_;
wire _5363_;
wire _5364_;
wire _5365_;
wire _5366_;
wire _5367_;
wire _5368_;
wire _5369_;
wire _5370_;
wire _5371_;
wire _5372_;
wire _5373_;
wire _5374_;
wire _5375_;
wire _5376_;
wire _5377_;
wire _5378_;
wire _5379_;
wire _5380_;
wire _5381_;
wire _5382_;
wire _5383_;
wire _5384_;
wire _5385_;
wire _5386_;
wire _5387_;
wire _5388_;
wire _5389_;
wire _5390_;
wire _5391_;
wire _5392_;
wire _5393_;
wire _5394_;
wire _5395_;
wire _5396_;
wire _5397_;
wire _5398_;
wire _5399_;
wire _5400_;
wire _5401_;
wire _5402_;
wire _5403_;
wire _5404_;
wire _5405_;
wire _5406_;
wire _5407_;
wire _5408_;
wire _5409_;
wire _5410_;
wire _5411_;
wire _5412_;
wire _5413_;
wire _5414_;
wire _5415_;
wire _5416_;
wire _5417_;
wire _5418_;
wire _5419_;
wire _5420_;
wire _5421_;
wire _5422_;
wire _5423_;
wire _5424_;
wire _5425_;
wire _5426_;
wire _5427_;
wire _5428_;
wire _5429_;
wire _5430_;
wire _5431_;
wire _5432_;
wire _5433_;
wire _5434_;
wire _5435_;
wire _5436_;
wire _5437_;
wire _5438_;
wire _5439_;
wire _5440_;
wire _5441_;
wire _5442_;
wire _5443_;
wire _5444_;
wire _5445_;
wire _5446_;
wire _5447_;
wire _5448_;
wire _5449_;
wire _5450_;
wire _5451_;
wire _5452_;
wire _5453_;
wire _5454_;
wire _5455_;
wire _5456_;
wire _5457_;
wire _5458_;
wire _5459_;
wire _5460_;
wire _5461_;
wire _5462_;
wire _5463_;
wire _5464_;
wire _5465_;
wire _5466_;
wire _5467_;
wire _5468_;
wire _5469_;
wire _5470_;
wire _5471_;
wire _5472_;
wire _5473_;
wire _5474_;
wire _5475_;
wire _5476_;
wire _5477_;
wire _5478_;
wire _5479_;
wire _5480_;
wire _5481_;
wire _5482_;
wire _5483_;
wire _5484_;
wire _5485_;
wire _5486_;
wire _5487_;
wire _5488_;
wire _5489_;
wire _5490_;
wire _5491_;
wire _5492_;
wire _5493_;
wire _5494_;
wire _5495_;
wire _5496_;
wire _5497_;
wire _5498_;
wire _5499_;
wire _5500_;
wire _5501_;
wire _5502_;
wire _5503_;
wire _5504_;
wire _5505_;
wire _5506_;
wire _5507_;
wire _5508_;
wire _5509_;
wire _5510_;
wire _5511_;
wire _5512_;
wire _5513_;
wire _5514_;
wire _5515_;
wire _5516_;
wire _5517_;
wire _5518_;
wire _5519_;
wire _5520_;
wire _5521_;
wire _5522_;
wire _5523_;
wire _5524_;
wire _5525_;
wire _5526_;
wire _5527_;
wire _5528_;
wire _5529_;
wire _5530_;
wire _5531_;
wire _5532_;
wire _5533_;
wire _5534_;
wire _5535_;
wire _5536_;
wire _5537_;
wire _5538_;
wire _5539_;
wire _5540_;
wire _5541_;
wire _5542_;
wire _5543_;
wire _5544_;
wire _5545_;
wire _5546_;
wire _5547_;
wire _5548_;
wire _5549_;
wire _5550_;
wire _5551_;
wire _5552_;
wire _5553_;
wire _5554_;
wire _5555_;
wire _5556_;
wire _5557_;
wire _5558_;
wire _5559_;
wire _5560_;
wire _5561_;
wire _5562_;
wire _5563_;
wire _5564_;
wire _5565_;
wire _5566_;
wire _5567_;
wire _5568_;
wire _5569_;
wire _5570_;
wire _5571_;
wire _5572_;
wire _5573_;
wire _5574_;
wire _5575_;
wire _5576_;
wire _5577_;
wire _5578_;
wire _5579_;
wire _5580_;
wire _5581_;
wire _5582_;
wire _5583_;
wire _5584_;
wire _5585_;
wire _5586_;
wire _5587_;
wire _5588_;
wire _5589_;
wire _5590_;
wire _5591_;
wire _5592_;
wire _5593_;
wire _5594_;
wire _5595_;
wire _5596_;
wire _5597_;
wire _5598_;
wire _5599_;
wire _5600_;
wire _5601_;
wire _5602_;
wire _5603_;
wire _5604_;
wire _5605_;
wire _5606_;
wire _5607_;
wire _5608_;
wire _5609_;
wire _5610_;
wire _5611_;
wire _5612_;
wire _5613_;
wire _5614_;
wire _5615_;
wire _5616_;
wire _5617_;
wire _5618_;
wire _5619_;
wire _5620_;
wire _5621_;
wire _5622_;
wire _5623_;
wire _5624_;
wire _5625_;
wire _5626_;
wire _5627_;
wire _5628_;
wire _5629_;
wire _5630_;
wire _5631_;
wire _5632_;
wire _5633_;
wire _5634_;
wire _5635_;
wire _5636_;
wire _5637_;
wire _5638_;
wire _5639_;
wire _5640_;
wire _5641_;
wire _5642_;
wire _5643_;
wire _5644_;
wire _5645_;
wire _5646_;
wire _5647_;
wire _5648_;
wire _5649_;
wire _5650_;
wire _5651_;
wire _5652_;
wire _5653_;
wire _5654_;
wire _5655_;
wire _5656_;
wire _5657_;
wire _5658_;
wire _5659_;
wire _5660_;
wire _5661_;
wire _5662_;
wire _5663_;
wire _5664_;
wire _5665_;
wire _5666_;
wire _5667_;
wire _5668_;
wire _5669_;
wire _5670_;
wire _5671_;
wire _5672_;
wire _5673_;
wire _5674_;
wire _5675_;
wire _5676_;
wire _5677_;
wire _5678_;
wire _5679_;
wire _5680_;
wire _5681_;
wire _5682_;
wire _5683_;
wire _5684_;
wire _5685_;
wire _5686_;
wire _5687_;
wire _5688_;
wire _5689_;
wire _5690_;
wire _5691_;
wire _5692_;
wire _5693_;
wire _5694_;
wire _5695_;
wire _5696_;
wire _5697_;
wire _5698_;
wire _5699_;
wire _5700_;
wire _5701_;
wire _5702_;
wire _5703_;
wire _5704_;
wire _5705_;
wire _5706_;
wire _5707_;
wire _5708_;
wire _5709_;
wire _5710_;
wire _5711_;
wire _5712_;
wire _5713_;
wire _5714_;
wire _5715_;
wire _5716_;
wire _5717_;
wire _5718_;
wire _5719_;
wire _5720_;
wire _5721_;
wire _5722_;
wire _5723_;
wire _5724_;
wire _5725_;
wire _5726_;
wire _5727_;
wire _5728_;
wire _5729_;
wire _5730_;
wire _5731_;
wire _5732_;
wire _5733_;
wire _5734_;
wire _5735_;
wire _5736_;
wire _5737_;
wire _5738_;
wire _5739_;
wire _5740_;
wire _5741_;
wire _5742_;
wire _5743_;
wire _5744_;
wire _5745_;
wire _5746_;
wire _5747_;
wire _5748_;
wire _5749_;
wire _5750_;
wire _5751_;
wire _5752_;
wire _5753_;
wire _5754_;
wire _5755_;
wire _5756_;
wire _5757_;
wire _5758_;
wire _5759_;
wire _5760_;
wire _5761_;
wire _5762_;
wire _5763_;
wire _5764_;
wire _5765_;
wire _5766_;
wire _5767_;
wire _5768_;
wire _5769_;
wire _5770_;
wire _5771_;
wire _5772_;
wire _5773_;
wire _5774_;
wire _5775_;
wire _5776_;
wire _5777_;
wire _5778_;
wire _5779_;
wire _5780_;
wire _5781_;
wire _5782_;
wire _5783_;
wire _5784_;
wire _5785_;
wire _5786_;
wire _5787_;
wire _5788_;
wire _5789_;
wire _5790_;
wire _5791_;
wire _5792_;
wire _5793_;
wire _5794_;
wire _5795_;
wire _5796_;
wire _5797_;
wire _5798_;
wire _5799_;
wire _5800_;
wire _5801_;
wire _5802_;
wire _5803_;
wire _5804_;
wire _5805_;
wire _5806_;
wire _5807_;
wire _5808_;
wire _5809_;
wire _5810_;
wire _5811_;
wire _5812_;
wire _5813_;
wire _5814_;
wire _5815_;
wire _5816_;
wire _5817_;
wire _5818_;
wire _5819_;
wire _5820_;
wire _5821_;
wire _5822_;
wire _5823_;
wire _5824_;
wire _5825_;
wire _5826_;
wire _5827_;
wire _5828_;
wire _5829_;
wire _5830_;
wire _5831_;
wire _5832_;
wire _5833_;
wire _5834_;
wire _5835_;
wire _5836_;
wire _5837_;
wire _5838_;
wire _5839_;
wire _5840_;
wire _5841_;
wire _5842_;
wire _5843_;
wire _5844_;
wire _5845_;
wire _5846_;
wire _5847_;
wire _5848_;
wire _5849_;
wire _5850_;
wire _5851_;
wire _5852_;
wire _5853_;
wire _5854_;
wire _5855_;
wire _5856_;
wire _5857_;
wire _5858_;
wire _5859_;
wire _5860_;
wire _5861_;
wire _5862_;
wire _5863_;
wire _5864_;
wire _5865_;
wire _5866_;
wire _5867_;
wire _5868_;
wire _5869_;
wire _5870_;
wire _5871_;
wire _5872_;
wire _5873_;
wire _5874_;
wire _5875_;
wire _5876_;
wire _5877_;
wire _5878_;
wire _5879_;
wire _5880_;
wire _5881_;
wire _5882_;
wire _5883_;
wire _5884_;
wire _5885_;
wire _5886_;
wire _5887_;
wire _5888_;
wire _5889_;
wire _5890_;
wire _5891_;
wire _5892_;
wire _5893_;
wire _5894_;
wire _5895_;
wire _5896_;
wire _5897_;
wire _5898_;
wire _5899_;
wire _5900_;
wire _5901_;
wire _5902_;
wire _5903_;
wire _5904_;
wire _5905_;
wire _5906_;
wire _5907_;
wire _5908_;
wire _5909_;
wire _5910_;
wire _5911_;
wire _5912_;
wire _5913_;
wire _5914_;
wire _5915_;
wire _5916_;
wire _5917_;
wire _5918_;
wire _5919_;
wire _5920_;
wire _5921_;
wire _5922_;
wire _5923_;
wire _5924_;
wire _5925_;
wire _5926_;
wire _5927_;
wire _5928_;
wire _5929_;
wire _5930_;
wire _5931_;
wire _5932_;
wire _5933_;
wire _5934_;
wire _5935_;
wire _5936_;
wire _5937_;
wire _5938_;
wire _5939_;
wire _5940_;
wire _5941_;
wire _5942_;
wire _5943_;
wire _5944_;
wire _5945_;
wire _5946_;
wire _5947_;
wire _5948_;
wire _5949_;
wire _5950_;
wire _5951_;
wire _5952_;
wire _5953_;
wire _5954_;
wire _5955_;
wire _5956_;
wire _5957_;
wire _5958_;
wire _5959_;
wire _5960_;
wire _5961_;
wire _5962_;
wire _5963_;
wire _5964_;
wire _5965_;
wire _5966_;
wire _5967_;
wire _5968_;
wire _5969_;
wire _5970_;
wire _5971_;
wire _5972_;
wire _5973_;
wire _5974_;
wire _5975_;
wire _5976_;
wire _5977_;
wire _5978_;
wire _5979_;
wire _5980_;
wire _5981_;
wire _5982_;
wire _5983_;
wire _5984_;
wire _5985_;
wire _5986_;
wire _5987_;
wire _5988_;
wire _5989_;
wire _5990_;
wire _5991_;
wire _5992_;
wire _5993_;
wire _5994_;
wire _5995_;
wire _5996_;
wire _5997_;
wire _5998_;
wire _5999_;
wire _6000_;
wire _6001_;
wire _6002_;
wire _6003_;
wire _6004_;
wire _6005_;
wire _6006_;
wire _6007_;
wire _6008_;
wire _6009_;
wire _6010_;
wire _6011_;
wire _6012_;
wire _6013_;
wire _6014_;
wire _6015_;
wire _6016_;
wire _6017_;
wire _6018_;
wire _6019_;
wire _6020_;
wire _6021_;
wire _6022_;
wire _6023_;
wire _6024_;
wire _6025_;
wire _6026_;
wire _6027_;
wire _6028_;
wire _6029_;
wire _6030_;
wire _6031_;
wire _6032_;
wire _6033_;
wire _6034_;
wire _6035_;
wire _6036_;
wire _6037_;
wire _6038_;
wire _6039_;
wire _6040_;
wire _6041_;
wire _6042_;
wire _6043_;
wire _6044_;
wire _6045_;
wire _6046_;
wire _6047_;
wire _6048_;
wire _6049_;
wire _6050_;
wire _6051_;
wire _6052_;
wire _6053_;
wire _6054_;
wire _6055_;
wire _6056_;
wire _6057_;
wire _6058_;
wire _6059_;
wire _6060_;
wire _6061_;
wire _6062_;
wire _6063_;
wire _6064_;
wire _6065_;
wire _6066_;
wire _6067_;
wire _6068_;
wire _6069_;
wire _6070_;
wire _6071_;
wire _6072_;
wire _6073_;
wire _6074_;
wire _6075_;
wire _6076_;
wire _6077_;
wire _6078_;
wire _6079_;
wire _6080_;
wire _6081_;
wire _6082_;
wire _6083_;
wire _6084_;
wire _6085_;
wire _6086_;
wire _6087_;
wire _6088_;
wire _6089_;
wire _6090_;
wire _6091_;
wire _6092_;
wire _6093_;
wire _6094_;
wire _6095_;
wire _6096_;
wire _6097_;
wire _6098_;
wire _6099_;
wire _6100_;
wire _6101_;
wire _6102_;
wire _6103_;
wire _6104_;
wire _6105_;
wire _6106_;
wire _6107_;
wire _6108_;
wire _6109_;
wire _6110_;
wire _6111_;
wire _6112_;
wire _6113_;
wire _6114_;
wire _6115_;
wire _6116_;
wire _6117_;
wire _6118_;
wire _6119_;
wire _6120_;
wire _6121_;
wire _6122_;
wire _6123_;
wire _6124_;
wire _6125_;
wire _6126_;
wire _6127_;
wire _6128_;
wire _6129_;
wire _6130_;
wire _6131_;
wire _6132_;
wire _6133_;
wire _6134_;
wire _6135_;
wire _6136_;
wire _6137_;
wire _6138_;
wire _6139_;
wire _6140_;
wire _6141_;
wire _6142_;
wire _6143_;
wire _6144_;
wire _6145_;
wire _6146_;
wire _6147_;
wire _6148_;
wire _6149_;
wire _6150_;
wire _6151_;
wire _6152_;
wire _6153_;
wire _6154_;
wire _6155_;
wire _6156_;
wire _6157_;
wire _6158_;
wire _6159_;
wire _6160_;
wire _6161_;
wire _6162_;
wire _6163_;
wire _6164_;
wire _6165_;
wire _6166_;
wire _6167_;
wire _6168_;
wire _6169_;
wire _6170_;
wire _6171_;
wire _6172_;
wire _6173_;
wire _6174_;
wire _6175_;
wire _6176_;
wire _6177_;
wire _6178_;
wire _6179_;
wire _6180_;
wire _6181_;
wire _6182_;
wire _6183_;
wire _6184_;
wire _6185_;
wire _6186_;
wire _6187_;
wire _6188_;
wire _6189_;
wire _6190_;
wire _6191_;
wire _6192_;
wire _6193_;
wire _6194_;
wire _6195_;
wire _6196_;
wire _6197_;
wire _6198_;
wire _6199_;
wire _6200_;
wire _6201_;
wire _6202_;
wire _6203_;
wire _6204_;
wire _6205_;
wire _6206_;
wire _6207_;
wire _6208_;
wire _6209_;
wire _6210_;
wire _6211_;
wire _6212_;
wire _6213_;
wire _6214_;
wire _6215_;
wire _6216_;
wire _6217_;
wire _6218_;
wire _6219_;
wire _6220_;
wire _6221_;
wire _6222_;
wire _6223_;
wire _6224_;
wire _6225_;
wire _6226_;
wire _6227_;
wire _6228_;
wire _6229_;
wire _6230_;
wire _6231_;
wire _6232_;
wire _6233_;
wire _6234_;
wire _6235_;
wire _6236_;
wire _6237_;
wire _6238_;
wire _6239_;
wire _6240_;
wire _6241_;
wire _6242_;
wire _6243_;
wire _6244_;
wire _6245_;
wire _6246_;
wire _6247_;
wire _6248_;
wire _6249_;
wire _6250_;
wire _6251_;
wire _6252_;
wire _6253_;
wire _6254_;
wire _6255_;
wire _6256_;
wire _6257_;
wire _6258_;
wire _6259_;
wire _6260_;
wire _6261_;
wire _6262_;
wire _6263_;
wire _6264_;
wire _6265_;
wire _6266_;
wire _6267_;
wire _6268_;
wire _6269_;
wire _6270_;
wire _6271_;
wire _6272_;
wire _6273_;
wire _6274_;
wire _6275_;
wire _6276_;
wire _6277_;
wire _6278_;
wire _6279_;
wire _6280_;
wire _6281_;
wire _6282_;
wire _6283_;
wire _6284_;
wire _6285_;
wire _6286_;
wire _6287_;
wire _6288_;
wire _6289_;
wire _6290_;
wire _6291_;
wire _6292_;
wire _6293_;
wire _6294_;
wire _6295_;
wire _6296_;
wire _6297_;
wire _6298_;
wire _6299_;
wire _6300_;
wire _6301_;
wire _6302_;
wire _6303_;
wire _6304_;
wire _6305_;
wire _6306_;
wire _6307_;
wire _6308_;
wire _6309_;
wire _6310_;
wire _6311_;
wire _6312_;
wire _6313_;
wire _6314_;
wire _6315_;
wire _6316_;
wire _6317_;
wire _6318_;
wire _6319_;
wire _6320_;
wire _6321_;
wire _6322_;
wire _6323_;
wire _6324_;
wire _6325_;
wire _6326_;
wire _6327_;
wire _6328_;
wire _6329_;
wire _6330_;
wire _6331_;
wire _6332_;
wire _6333_;
wire _6334_;
wire _6335_;
wire _6336_;
wire _6337_;
wire _6338_;
wire _6339_;
wire _6340_;
wire _6341_;
wire _6342_;
wire _6343_;
wire _6344_;
wire _6345_;
wire _6346_;
wire _6347_;
wire _6348_;
wire _6349_;
wire _6350_;
wire _6351_;
wire _6352_;
wire _6353_;
wire _6354_;
wire _6355_;
wire _6356_;
wire _6357_;
wire _6358_;
wire _6359_;
wire _6360_;
wire _6361_;
wire _6362_;
wire _6363_;
wire _6364_;
wire _6365_;
wire _6366_;
wire _6367_;
wire _6368_;
wire _6369_;
wire _6370_;
wire _6371_;
wire _6372_;
wire _6373_;
wire _6374_;
wire _6375_;
wire _6376_;
wire _6377_;
wire _6378_;
wire _6379_;
wire _6380_;
wire _6381_;
wire _6382_;
wire _6383_;
wire _6384_;
wire _6385_;
wire _6386_;
wire _6387_;
wire _6388_;
wire _6389_;
wire _6390_;
wire _6391_;
wire _6392_;
wire _6393_;
wire _6394_;
wire _6395_;
wire _6396_;
wire _6397_;
wire _6398_;
wire _6399_;
wire _6400_;
wire _6401_;
wire _6402_;
wire _6403_;
wire _6404_;
wire _6405_;
wire _6406_;
wire _6407_;
wire _6408_;
wire _6409_;
wire _6410_;
wire _6411_;
wire _6412_;
wire _6413_;
wire _6414_;
wire _6415_;
wire _6416_;
wire _6417_;
wire _6418_;
wire _6419_;
wire _6420_;
wire _6421_;
wire _6422_;
wire _6423_;
wire _6424_;
wire _6425_;
wire _6426_;
wire _6427_;
wire _6428_;
wire _6429_;
wire _6430_;
wire _6431_;
wire _6432_;
wire _6433_;
wire _6434_;
wire _6435_;
wire _6436_;
wire _6437_;
wire _6438_;
wire _6439_;
wire _6440_;
wire _6441_;
wire _6442_;
wire _6443_;
wire _6444_;
wire _6445_;
wire _6446_;
wire _6447_;
wire _6448_;
wire _6449_;
wire _6450_;
wire _6451_;
wire _6452_;
wire _6453_;
wire _6454_;
wire _6455_;
wire _6456_;
wire _6457_;
wire _6458_;
wire _6459_;
wire _6460_;
wire _6461_;
wire _6462_;
wire _6463_;
wire _6464_;
wire _6465_;
wire _6466_;
wire _6467_;
wire _6468_;
wire _6469_;
wire _6470_;
wire _6471_;
wire _6472_;
wire _6473_;
wire _6474_;
wire _6475_;
wire _6476_;
wire _6477_;
wire _6478_;
wire _6479_;
wire _6480_;
wire _6481_;
wire _6482_;
wire _6483_;
wire _6484_;
wire _6485_;
wire _6486_;
wire _6487_;
wire _6488_;
wire _6489_;
wire _6490_;
wire _6491_;
wire _6492_;
wire _6493_;
wire _6494_;
wire _6495_;
wire _6496_;
wire _6497_;
wire _6498_;
wire _6499_;
wire _6500_;
wire _6501_;
wire _6502_;
wire _6503_;
wire _6504_;
wire _6505_;
wire _6506_;
wire _6507_;
wire _6508_;
wire _6509_;
wire _6510_;
wire _6511_;
wire _6512_;
wire _6513_;
wire _6514_;
wire _6515_;
wire _6516_;
wire _6517_;
wire _6518_;
wire _6519_;
wire _6520_;
wire _6521_;
wire _6522_;
wire _6523_;
wire _6524_;
wire _6525_;
wire _6526_;
wire _6527_;
wire _6528_;
wire _6529_;
wire _6530_;
wire _6531_;
wire _6532_;
wire _6533_;
wire _6534_;
wire _6535_;
wire _6536_;
wire _6537_;
wire _6538_;
wire _6539_;
wire _6540_;
wire _6541_;
wire _6542_;
wire _6543_;
wire _6544_;
wire _6545_;
wire _6546_;
wire _6547_;
wire _6548_;
wire _6549_;
wire _6550_;
wire _6551_;
wire _6552_;
wire _6553_;
wire _6554_;
wire _6555_;
wire _6556_;
wire _6557_;
wire _6558_;
wire _6559_;
wire _6560_;
wire _6561_;
wire _6562_;
wire _6563_;
wire _6564_;
wire _6565_;
wire _6566_;
wire _6567_;
wire _6568_;
wire _6569_;
wire _6570_;
wire _6571_;
wire _6572_;
wire _6573_;
wire _6574_;
wire _6575_;
wire _6576_;
wire _6577_;
wire _6578_;
wire _6579_;
wire _6580_;
wire _6581_;
wire _6582_;
wire _6583_;
wire _6584_;
wire _6585_;
wire _6586_;
wire _6587_;
wire _6588_;
wire _6589_;
wire _6590_;
wire _6591_;
wire _6592_;
wire _6593_;
wire _6594_;
wire _6595_;
wire _6596_;
wire _6597_;
wire _6598_;
wire _6599_;
wire _6600_;
wire _6601_;
wire _6602_;
wire _6603_;
wire _6604_;
wire _6605_;
wire _6606_;
wire _6607_;
wire _6608_;
wire _6609_;
wire _6610_;
wire _6611_;
wire _6612_;
wire _6613_;
wire _6614_;
wire _6615_;
wire _6616_;
wire _6617_;
wire _6618_;
wire _6619_;
wire _6620_;
wire _6621_;
wire _6622_;
wire _6623_;
wire _6624_;
wire _6625_;
wire _6626_;
wire _6627_;
wire _6628_;
wire _6629_;
wire _6630_;
wire _6631_;
wire _6632_;
wire _6633_;
wire _6634_;
wire _6635_;
wire _6636_;
wire _6637_;
wire _6638_;
wire _6639_;
wire _6640_;
wire _6641_;
wire _6642_;
wire _6643_;
wire _6644_;
wire _6645_;
wire _6646_;
wire _6647_;
wire _6648_;
wire _6649_;
wire _6650_;
wire _6651_;
wire _6652_;
wire _6653_;
wire _6654_;
wire _6655_;
wire _6656_;
wire _6657_;
wire _6658_;
wire _6659_;
wire _6660_;
wire _6661_;
wire _6662_;
wire _6663_;
wire _6664_;
wire _6665_;
wire _6666_;
wire _6667_;
wire _6668_;
wire _6669_;
wire _6670_;
wire _6671_;
wire _6672_;
wire _6673_;
wire _6674_;
wire _6675_;
wire _6676_;
wire _6677_;
wire _6678_;
wire _6679_;
wire _6680_;
wire _6681_;
wire _6682_;
wire _6683_;
wire _6684_;
wire _6685_;
wire _6686_;
wire _6687_;
wire _6688_;
wire _6689_;
wire _6690_;
wire _6691_;
wire _6692_;
wire _6693_;
wire _6694_;
wire _6695_;
wire _6696_;
wire _6697_;
wire _6698_;
wire _6699_;
wire _6700_;
wire _6701_;
wire _6702_;
wire _6703_;
wire _6704_;
wire _6705_;
wire _6706_;
wire _6707_;
wire _6708_;
wire _6709_;
wire _6710_;
wire _6711_;
wire _6712_;
wire _6713_;
wire _6714_;
wire _6715_;
wire _6716_;
wire _6717_;
wire _6718_;
wire _6719_;
wire _6720_;
wire _6721_;
wire _6722_;
wire _6723_;
wire _6724_;
wire _6725_;
wire _6726_;
wire _6727_;
wire _6728_;
wire _6729_;
wire _6730_;
wire _6731_;
wire _6732_;
wire _6733_;
wire _6734_;
wire _6735_;
wire _6736_;
wire _6737_;
wire _6738_;
wire _6739_;
wire _6740_;
wire _6741_;
wire _6742_;
wire _6743_;
wire _6744_;
wire _6745_;
wire _6746_;
wire _6747_;
wire _6748_;
wire _6749_;
wire _6750_;
wire _6751_;
wire _6752_;
wire _6753_;
wire _6754_;
wire _6755_;
wire _6756_;
wire _6757_;
wire _6758_;
wire _6759_;
wire _6760_;
wire _6761_;
wire _6762_;
wire _6763_;
wire _6764_;
wire _6765_;
wire _6766_;
wire _6767_;
wire _6768_;
wire _6769_;
wire _6770_;
wire _6771_;
wire _6772_;
wire _6773_;
wire _6774_;
wire _6775_;
wire _6776_;
wire _6777_;
wire _6778_;
wire _6779_;
wire _6780_;
wire _6781_;
wire _6782_;
wire _6783_;
wire _6784_;
wire _6785_;
wire _6786_;
wire _6787_;
wire _6788_;
wire _6789_;
wire _6790_;
wire _6791_;
wire _6792_;
wire _6793_;
wire _6794_;
wire _6795_;
wire _6796_;
wire _6797_;
wire _6798_;
wire _6799_;
wire _6800_;
wire _6801_;
wire _6802_;
wire _6803_;
wire _6804_;
wire _6805_;
wire _6806_;
wire _6807_;
wire _6808_;
wire _6809_;
wire _6810_;
wire _6811_;
wire _6812_;
wire _6813_;
wire _6814_;
wire _6815_;
wire _6816_;
wire _6817_;
wire _6818_;
wire _6819_;
wire _6820_;
wire _6821_;
wire _6822_;
wire _6823_;
wire _6824_;
wire _6825_;
wire _6826_;
wire _6827_;
wire _6828_;
wire _6829_;
wire _6830_;
wire _6831_;
wire _6832_;
wire _6833_;
wire _6834_;
wire _6835_;
wire _6836_;
wire _6837_;
wire _6838_;
wire _6839_;
wire _6840_;
wire _6841_;
wire _6842_;
wire _6843_;
wire _6844_;
wire _6845_;
wire _6846_;
wire _6847_;
wire _6848_;
wire _6849_;
wire _6850_;
wire _6851_;
wire _6852_;
wire _6853_;
wire _6854_;
wire _6855_;
wire _6856_;
wire _6857_;
wire _6858_;
wire _6859_;
wire _6860_;
wire _6861_;
wire _6862_;
wire _6863_;
wire _6864_;
wire _6865_;
wire _6866_;
wire _6867_;
wire _6868_;
wire _6869_;
wire _6870_;
wire _6871_;
wire _6872_;
wire _6873_;
wire _6874_;
wire _6875_;
wire _6876_;
wire _6877_;
wire _6878_;
wire _6879_;
wire _6880_;
wire _6881_;
wire _6882_;
wire _6883_;
wire _6884_;
wire _6885_;
wire _6886_;
wire _6887_;
wire _6888_;
wire _6889_;
wire _6890_;
wire _6891_;
wire _6892_;
wire _6893_;
wire _6894_;
wire _6895_;
wire _6896_;
wire _6897_;
wire _6898_;
wire _6899_;
wire _6900_;
wire _6901_;
wire _6902_;
wire _6903_;
wire _6904_;
wire _6905_;
wire _6906_;
wire _6907_;
wire _6908_;
wire _6909_;
wire _6910_;
wire _6911_;
wire _6912_;
wire _6913_;
wire _6914_;
wire _6915_;
wire _6916_;
wire _6917_;
wire _6918_;
wire _6919_;
wire _6920_;
wire _6921_;
wire _6922_;
wire _6923_;
wire _6924_;
wire _6925_;
wire _6926_;
wire _6927_;
wire _6928_;
wire _6929_;
wire _6930_;
wire _6931_;
wire _6932_;
wire _6933_;
wire _6934_;
wire _6935_;
wire _6936_;
wire _6937_;
wire _6938_;
wire _6939_;
wire _6940_;
wire _6941_;
wire _6942_;
wire _6943_;
wire _6944_;
wire _6945_;
wire _6946_;
wire _6947_;
wire _6948_;
wire _6949_;
wire _6950_;
wire _6951_;
wire _6952_;
wire _6953_;
wire _6954_;
wire _6955_;
wire _6956_;
wire _6957_;
wire _6958_;
wire _6959_;
wire _6960_;
wire _6961_;
wire _6962_;
wire _6963_;
wire _6964_;
wire _6965_;
wire _6966_;
wire _6967_;
wire _6968_;
wire _6969_;
wire _6970_;
wire _6971_;
wire _6972_;
wire _6973_;
wire _6974_;
wire _6975_;
wire _6976_;
wire _6977_;
wire _6978_;
wire _6979_;
wire _6980_;
wire _6981_;
wire _6982_;
wire _6983_;
wire _6984_;
wire _6985_;
wire _6986_;
wire _6987_;
wire _6988_;
wire _6989_;
wire _6990_;
wire _6991_;
wire _6992_;
wire _6993_;
wire _6994_;
wire _6995_;
wire _6996_;
wire _6997_;
wire _6998_;
wire _6999_;
wire _7000_;
wire _7001_;
wire _7002_;
wire _7003_;
wire _7004_;
wire _7005_;
wire _7006_;
wire _7007_;
wire _7008_;
wire _7009_;
wire _7010_;
wire _7011_;
wire _7012_;
wire _7013_;
wire _7014_;
wire _7015_;
wire _7016_;
wire _7017_;
wire _7018_;
wire _7019_;
wire _7020_;
wire _7021_;
wire _7022_;
wire _7023_;
wire _7024_;
wire _7025_;
wire _7026_;
wire _7027_;
wire _7028_;
wire _7029_;
wire _7030_;
wire _7031_;
wire _7032_;
wire _7033_;
wire _7034_;
wire _7035_;
wire _7036_;
wire _7037_;
wire _7038_;
wire _7039_;
wire _7040_;
wire _7041_;
wire _7042_;
wire _7043_;
wire _7044_;
wire _7045_;
wire _7046_;
wire _7047_;
wire _7048_;
wire _7049_;
wire _7050_;
wire _7051_;
wire _7052_;
wire _7053_;
wire _7054_;
wire _7055_;
wire _7056_;
wire _7057_;
wire _7058_;
wire _7059_;
wire _7060_;
wire _7061_;
wire _7062_;
wire _7063_;
wire _7064_;
wire _7065_;
wire _7066_;
wire _7067_;
wire _7068_;
wire _7069_;
wire _7070_;
wire _7071_;
wire _7072_;
wire _7073_;
wire _7074_;
wire _7075_;
wire _7076_;
wire _7077_;
wire _7078_;
wire _7079_;
wire _7080_;
wire _7081_;
wire _7082_;
wire _7083_;
wire _7084_;
wire _7085_;
wire _7086_;
wire _7087_;
wire _7088_;
wire _7089_;
wire _7090_;
wire _7091_;
wire _7092_;
wire _7093_;
wire _7094_;
wire _7095_;
wire _7096_;
wire _7097_;
wire _7098_;
wire _7099_;
wire _7100_;
wire _7101_;
wire _7102_;
wire _7103_;
wire _7104_;
wire _7105_;
wire _7106_;
wire _7107_;
wire _7108_;
wire _7109_;
wire _7110_;
wire _7111_;
wire _7112_;
wire _7113_;
wire _7114_;
wire _7115_;
wire _7116_;
wire _7117_;
wire _7118_;
wire _7119_;
wire _7120_;
wire _7121_;
wire _7122_;
wire _7123_;
wire _7124_;
wire _7125_;
wire _7126_;
wire _7127_;
wire _7128_;
wire _7129_;
wire _7130_;
wire _7131_;
wire _7132_;
wire _7133_;
wire _7134_;
wire _7135_;
wire _7136_;
wire _7137_;
wire _7138_;
wire _7139_;
wire _7140_;
wire _7141_;
wire _7142_;
wire _7143_;
wire _7144_;
wire _7145_;
wire _7146_;
wire _7147_;
wire _7148_;
wire _7149_;
wire _7150_;
wire _7151_;
wire _7152_;
wire _7153_;
wire _7154_;
wire _7155_;
wire _7156_;
wire _7157_;
wire _7158_;
wire _7159_;
wire _7160_;
wire _7161_;
wire _7162_;
wire _7163_;
wire _7164_;
wire _7165_;
wire _7166_;
wire _7167_;
wire _7168_;
wire _7169_;
wire _7170_;
wire _7171_;
wire _7172_;
wire _7173_;
wire _7174_;
wire _7175_;
wire _7176_;
wire _7177_;
wire _7178_;
wire _7179_;
wire _7180_;
wire _7181_;
wire _7182_;
wire _7183_;
wire _7184_;
wire _7185_;
wire _7186_;
wire _7187_;
wire _7188_;
wire _7189_;
wire _7190_;
wire _7191_;
wire _7192_;
wire _7193_;
wire _7194_;
wire _7195_;
wire _7196_;
wire _7197_;
wire _7198_;
wire _7199_;
wire _7200_;
wire _7201_;
wire _7202_;
wire _7203_;
wire _7204_;
wire _7205_;
wire _7206_;
wire _7207_;
wire _7208_;
wire _7209_;
wire _7210_;
wire _7211_;
wire _7212_;
wire _7213_;
wire _7214_;
wire _7215_;
wire _7216_;
wire _7217_;
wire _7218_;
wire _7219_;
wire _7220_;
wire _7221_;
wire _7222_;
wire _7223_;
wire _7224_;
wire _7225_;
wire _7226_;
wire _7227_;
wire _7228_;
wire _7229_;
wire _7230_;
wire _7231_;
wire _7232_;
wire _7233_;
wire _7234_;
wire _7235_;
wire _7236_;
wire _7237_;
wire _7238_;
wire _7239_;
wire _7240_;
wire _7241_;
wire _7242_;
wire _7243_;
wire _7244_;
wire _7245_;
wire _7246_;
wire _7247_;
wire _7248_;
wire _7249_;
wire _7250_;
wire _7251_;
wire _7252_;
wire _7253_;
wire _7254_;
wire _7255_;
wire _7256_;
wire _7257_;
wire _7258_;
wire _7259_;
wire _7260_;
wire _7261_;
wire _7262_;
wire _7263_;
wire _7264_;
wire _7265_;
wire _7266_;
wire _7267_;
wire _7268_;
wire _7269_;
wire _7270_;
wire _7271_;
wire _7272_;
wire _7273_;
wire _7274_;
wire _7275_;
wire _7276_;
wire _7277_;
wire _7278_;
wire _7279_;
wire _7280_;
wire _7281_;
wire _7282_;
wire _7283_;
wire _7284_;
wire _7285_;
wire _7286_;
wire _7287_;
wire _7288_;
wire _7289_;
wire _7290_;
wire _7291_;
wire _7292_;
wire _7293_;
wire _7294_;
wire _7295_;
wire _7296_;
wire _7297_;
wire _7298_;
wire _7299_;
wire _7300_;
wire _7301_;
wire _7302_;
wire _7303_;
wire _7304_;
wire _7305_;
wire _7306_;
wire _7307_;
wire _7308_;
wire _7309_;
wire _7310_;
wire _7311_;
wire _7312_;
wire _7313_;
wire _7314_;
wire _7315_;
wire _7316_;
wire _7317_;
wire _7318_;
wire _7319_;
wire _7320_;
wire _7321_;
wire _7322_;
wire _7323_;
wire _7324_;
wire _7325_;
wire _7326_;
wire zeroWire;
wire oneWire;
assign zeroWire = 1'b0 /*12827*/;
assign oneWire = 1'b1 /*12827*/;
assign _37_ = ~D[0] /*12633*/;
assign _34_ = R_0[31] & _37_ /*12629*/;
assign _35_ = R_0[31] ^ _37_ /*12632*/;
assign _36_ = oneWire & _35_ /*12630*/;
assign _0_ = oneWire ^ _35_ /*12631*/;
assign _33_ = _34_ | _36_ /*12628*/;
assign _42_ = ~D[1] /*12627*/;
assign _39_ = R_0[32] & _42_ /*12623*/;
assign _40_ = R_0[32] ^ _42_ /*12626*/;
assign _41_ = _33_ & _40_ /*12624*/;
assign _1_ = _33_ ^ _40_ /*12625*/;
assign _38_ = _39_ | _41_ /*12622*/;
assign _47_ = ~D[2] /*12621*/;
assign _44_ = R_0[33] & _47_ /*12617*/;
assign _45_ = R_0[33] ^ _47_ /*12620*/;
assign _46_ = _38_ & _45_ /*12618*/;
assign _2_ = _38_ ^ _45_ /*12619*/;
assign _43_ = _44_ | _46_ /*12616*/;
assign _52_ = ~D[3] /*12615*/;
assign _49_ = R_0[34] & _52_ /*12611*/;
assign _50_ = R_0[34] ^ _52_ /*12614*/;
assign _51_ = _43_ & _50_ /*12612*/;
assign _3_ = _43_ ^ _50_ /*12613*/;
assign _48_ = _49_ | _51_ /*12610*/;
assign _57_ = ~D[4] /*12609*/;
assign _54_ = R_0[35] & _57_ /*12605*/;
assign _55_ = R_0[35] ^ _57_ /*12608*/;
assign _56_ = _48_ & _55_ /*12606*/;
assign _4_ = _48_ ^ _55_ /*12607*/;
assign _53_ = _54_ | _56_ /*12604*/;
assign _62_ = ~D[5] /*12603*/;
assign _59_ = R_0[36] & _62_ /*12599*/;
assign _60_ = R_0[36] ^ _62_ /*12602*/;
assign _61_ = _53_ & _60_ /*12600*/;
assign _5_ = _53_ ^ _60_ /*12601*/;
assign _58_ = _59_ | _61_ /*12598*/;
assign _67_ = ~D[6] /*12597*/;
assign _64_ = R_0[37] & _67_ /*12593*/;
assign _65_ = R_0[37] ^ _67_ /*12596*/;
assign _66_ = _58_ & _65_ /*12594*/;
assign _6_ = _58_ ^ _65_ /*12595*/;
assign _63_ = _64_ | _66_ /*12592*/;
assign _72_ = ~D[7] /*12591*/;
assign _69_ = R_0[38] & _72_ /*12587*/;
assign _70_ = R_0[38] ^ _72_ /*12590*/;
assign _71_ = _63_ & _70_ /*12588*/;
assign _7_ = _63_ ^ _70_ /*12589*/;
assign _68_ = _69_ | _71_ /*12586*/;
assign _77_ = ~D[8] /*12585*/;
assign _74_ = R_0[39] & _77_ /*12581*/;
assign _75_ = R_0[39] ^ _77_ /*12584*/;
assign _76_ = _68_ & _75_ /*12582*/;
assign _8_ = _68_ ^ _75_ /*12583*/;
assign _73_ = _74_ | _76_ /*12580*/;
assign _82_ = ~D[9] /*12579*/;
assign _79_ = R_0[40] & _82_ /*12575*/;
assign _80_ = R_0[40] ^ _82_ /*12578*/;
assign _81_ = _73_ & _80_ /*12576*/;
assign _9_ = _73_ ^ _80_ /*12577*/;
assign _78_ = _79_ | _81_ /*12574*/;
assign _87_ = ~D[10] /*12573*/;
assign _84_ = R_0[41] & _87_ /*12569*/;
assign _85_ = R_0[41] ^ _87_ /*12572*/;
assign _86_ = _78_ & _85_ /*12570*/;
assign _10_ = _78_ ^ _85_ /*12571*/;
assign _83_ = _84_ | _86_ /*12568*/;
assign _92_ = ~D[11] /*12567*/;
assign _89_ = R_0[42] & _92_ /*12563*/;
assign _90_ = R_0[42] ^ _92_ /*12566*/;
assign _91_ = _83_ & _90_ /*12564*/;
assign _11_ = _83_ ^ _90_ /*12565*/;
assign _88_ = _89_ | _91_ /*12562*/;
assign _97_ = ~D[12] /*12561*/;
assign _94_ = R_0[43] & _97_ /*12557*/;
assign _95_ = R_0[43] ^ _97_ /*12560*/;
assign _96_ = _88_ & _95_ /*12558*/;
assign _12_ = _88_ ^ _95_ /*12559*/;
assign _93_ = _94_ | _96_ /*12556*/;
assign _102_ = ~D[13] /*12555*/;
assign _99_ = R_0[44] & _102_ /*12551*/;
assign _100_ = R_0[44] ^ _102_ /*12554*/;
assign _101_ = _93_ & _100_ /*12552*/;
assign _13_ = _93_ ^ _100_ /*12553*/;
assign _98_ = _99_ | _101_ /*12550*/;
assign _107_ = ~D[14] /*12549*/;
assign _104_ = R_0[45] & _107_ /*12545*/;
assign _105_ = R_0[45] ^ _107_ /*12548*/;
assign _106_ = _98_ & _105_ /*12546*/;
assign _14_ = _98_ ^ _105_ /*12547*/;
assign _103_ = _104_ | _106_ /*12544*/;
assign _112_ = ~D[15] /*12543*/;
assign _109_ = R_0[46] & _112_ /*12539*/;
assign _110_ = R_0[46] ^ _112_ /*12542*/;
assign _111_ = _103_ & _110_ /*12540*/;
assign _15_ = _103_ ^ _110_ /*12541*/;
assign _108_ = _109_ | _111_ /*12538*/;
assign _117_ = ~D[16] /*12537*/;
assign _114_ = R_0[47] & _117_ /*12533*/;
assign _115_ = R_0[47] ^ _117_ /*12536*/;
assign _116_ = _108_ & _115_ /*12534*/;
assign _16_ = _108_ ^ _115_ /*12535*/;
assign _113_ = _114_ | _116_ /*12532*/;
assign _122_ = ~D[17] /*12531*/;
assign _119_ = R_0[48] & _122_ /*12527*/;
assign _120_ = R_0[48] ^ _122_ /*12530*/;
assign _121_ = _113_ & _120_ /*12528*/;
assign _17_ = _113_ ^ _120_ /*12529*/;
assign _118_ = _119_ | _121_ /*12526*/;
assign _127_ = ~D[18] /*12525*/;
assign _124_ = R_0[49] & _127_ /*12521*/;
assign _125_ = R_0[49] ^ _127_ /*12524*/;
assign _126_ = _118_ & _125_ /*12522*/;
assign _18_ = _118_ ^ _125_ /*12523*/;
assign _123_ = _124_ | _126_ /*12520*/;
assign _132_ = ~D[19] /*12519*/;
assign _129_ = R_0[50] & _132_ /*12515*/;
assign _130_ = R_0[50] ^ _132_ /*12518*/;
assign _131_ = _123_ & _130_ /*12516*/;
assign _19_ = _123_ ^ _130_ /*12517*/;
assign _128_ = _129_ | _131_ /*12514*/;
assign _137_ = ~D[20] /*12513*/;
assign _134_ = R_0[51] & _137_ /*12509*/;
assign _135_ = R_0[51] ^ _137_ /*12512*/;
assign _136_ = _128_ & _135_ /*12510*/;
assign _20_ = _128_ ^ _135_ /*12511*/;
assign _133_ = _134_ | _136_ /*12508*/;
assign _142_ = ~D[21] /*12507*/;
assign _139_ = R_0[52] & _142_ /*12503*/;
assign _140_ = R_0[52] ^ _142_ /*12506*/;
assign _141_ = _133_ & _140_ /*12504*/;
assign _21_ = _133_ ^ _140_ /*12505*/;
assign _138_ = _139_ | _141_ /*12502*/;
assign _147_ = ~D[22] /*12501*/;
assign _144_ = R_0[53] & _147_ /*12497*/;
assign _145_ = R_0[53] ^ _147_ /*12500*/;
assign _146_ = _138_ & _145_ /*12498*/;
assign _22_ = _138_ ^ _145_ /*12499*/;
assign _143_ = _144_ | _146_ /*12496*/;
assign _152_ = ~D[23] /*12495*/;
assign _149_ = R_0[54] & _152_ /*12491*/;
assign _150_ = R_0[54] ^ _152_ /*12494*/;
assign _151_ = _143_ & _150_ /*12492*/;
assign _23_ = _143_ ^ _150_ /*12493*/;
assign _148_ = _149_ | _151_ /*12490*/;
assign _157_ = ~D[24] /*12489*/;
assign _154_ = R_0[55] & _157_ /*12485*/;
assign _155_ = R_0[55] ^ _157_ /*12488*/;
assign _156_ = _148_ & _155_ /*12486*/;
assign _24_ = _148_ ^ _155_ /*12487*/;
assign _153_ = _154_ | _156_ /*12484*/;
assign _162_ = ~D[25] /*12483*/;
assign _159_ = R_0[56] & _162_ /*12479*/;
assign _160_ = R_0[56] ^ _162_ /*12482*/;
assign _161_ = _153_ & _160_ /*12480*/;
assign _25_ = _153_ ^ _160_ /*12481*/;
assign _158_ = _159_ | _161_ /*12478*/;
assign _167_ = ~D[26] /*12477*/;
assign _164_ = R_0[57] & _167_ /*12473*/;
assign _165_ = R_0[57] ^ _167_ /*12476*/;
assign _166_ = _158_ & _165_ /*12474*/;
assign _26_ = _158_ ^ _165_ /*12475*/;
assign _163_ = _164_ | _166_ /*12472*/;
assign _172_ = ~D[27] /*12471*/;
assign _169_ = R_0[58] & _172_ /*12467*/;
assign _170_ = R_0[58] ^ _172_ /*12470*/;
assign _171_ = _163_ & _170_ /*12468*/;
assign _27_ = _163_ ^ _170_ /*12469*/;
assign _168_ = _169_ | _171_ /*12466*/;
assign _177_ = ~D[28] /*12465*/;
assign _174_ = R_0[59] & _177_ /*12461*/;
assign _175_ = R_0[59] ^ _177_ /*12464*/;
assign _176_ = _168_ & _175_ /*12462*/;
assign _28_ = _168_ ^ _175_ /*12463*/;
assign _173_ = _174_ | _176_ /*12460*/;
assign _182_ = ~D[29] /*12459*/;
assign _179_ = R_0[60] & _182_ /*12455*/;
assign _180_ = R_0[60] ^ _182_ /*12458*/;
assign _181_ = _173_ & _180_ /*12456*/;
assign _29_ = _173_ ^ _180_ /*12457*/;
assign _178_ = _179_ | _181_ /*12454*/;
assign _187_ = ~D[30] /*12453*/;
assign _184_ = R_0[61] & _187_ /*12449*/;
assign _185_ = R_0[61] ^ _187_ /*12452*/;
assign _186_ = _178_ & _185_ /*12450*/;
assign _30_ = _178_ ^ _185_ /*12451*/;
assign _183_ = _184_ | _186_ /*12448*/;
assign _188_ = zeroWire & oneWire /*12443*/;
assign _189_ = zeroWire ^ oneWire /*12446*/;
assign _190_ = _183_ & _189_ /*12444*/;
assign _31_ = _183_ ^ _189_ /*12445*/;
assign Q[31] = _188_ | _190_ /*12442*/;
assign _230_ = D[0] ^ Q[31] /*12250*/;
assign _227_ = R_0[30] & _230_ /*12246*/;
assign _228_ = R_0[30] ^ _230_ /*12249*/;
assign _229_ = Q[31] & _228_ /*12247*/;
assign _193_ = Q[31] ^ _228_ /*12248*/;
assign _226_ = _227_ | _229_ /*12245*/;
assign _235_ = D[1] ^ Q[31] /*12244*/;
assign _232_ = _0_ & _235_ /*12240*/;
assign _233_ = _0_ ^ _235_ /*12243*/;
assign _234_ = _226_ & _233_ /*12241*/;
assign _194_ = _226_ ^ _233_ /*12242*/;
assign _231_ = _232_ | _234_ /*12239*/;
assign _240_ = D[2] ^ Q[31] /*12238*/;
assign _237_ = _1_ & _240_ /*12234*/;
assign _238_ = _1_ ^ _240_ /*12237*/;
assign _239_ = _231_ & _238_ /*12235*/;
assign _195_ = _231_ ^ _238_ /*12236*/;
assign _236_ = _237_ | _239_ /*12233*/;
assign _245_ = D[3] ^ Q[31] /*12232*/;
assign _242_ = _2_ & _245_ /*12228*/;
assign _243_ = _2_ ^ _245_ /*12231*/;
assign _244_ = _236_ & _243_ /*12229*/;
assign _196_ = _236_ ^ _243_ /*12230*/;
assign _241_ = _242_ | _244_ /*12227*/;
assign _250_ = D[4] ^ Q[31] /*12226*/;
assign _247_ = _3_ & _250_ /*12222*/;
assign _248_ = _3_ ^ _250_ /*12225*/;
assign _249_ = _241_ & _248_ /*12223*/;
assign _197_ = _241_ ^ _248_ /*12224*/;
assign _246_ = _247_ | _249_ /*12221*/;
assign _255_ = D[5] ^ Q[31] /*12220*/;
assign _252_ = _4_ & _255_ /*12216*/;
assign _253_ = _4_ ^ _255_ /*12219*/;
assign _254_ = _246_ & _253_ /*12217*/;
assign _198_ = _246_ ^ _253_ /*12218*/;
assign _251_ = _252_ | _254_ /*12215*/;
assign _260_ = D[6] ^ Q[31] /*12214*/;
assign _257_ = _5_ & _260_ /*12210*/;
assign _258_ = _5_ ^ _260_ /*12213*/;
assign _259_ = _251_ & _258_ /*12211*/;
assign _199_ = _251_ ^ _258_ /*12212*/;
assign _256_ = _257_ | _259_ /*12209*/;
assign _265_ = D[7] ^ Q[31] /*12208*/;
assign _262_ = _6_ & _265_ /*12204*/;
assign _263_ = _6_ ^ _265_ /*12207*/;
assign _264_ = _256_ & _263_ /*12205*/;
assign _200_ = _256_ ^ _263_ /*12206*/;
assign _261_ = _262_ | _264_ /*12203*/;
assign _270_ = D[8] ^ Q[31] /*12202*/;
assign _267_ = _7_ & _270_ /*12198*/;
assign _268_ = _7_ ^ _270_ /*12201*/;
assign _269_ = _261_ & _268_ /*12199*/;
assign _201_ = _261_ ^ _268_ /*12200*/;
assign _266_ = _267_ | _269_ /*12197*/;
assign _275_ = D[9] ^ Q[31] /*12196*/;
assign _272_ = _8_ & _275_ /*12192*/;
assign _273_ = _8_ ^ _275_ /*12195*/;
assign _274_ = _266_ & _273_ /*12193*/;
assign _202_ = _266_ ^ _273_ /*12194*/;
assign _271_ = _272_ | _274_ /*12191*/;
assign _280_ = D[10] ^ Q[31] /*12190*/;
assign _277_ = _9_ & _280_ /*12186*/;
assign _278_ = _9_ ^ _280_ /*12189*/;
assign _279_ = _271_ & _278_ /*12187*/;
assign _203_ = _271_ ^ _278_ /*12188*/;
assign _276_ = _277_ | _279_ /*12185*/;
assign _285_ = D[11] ^ Q[31] /*12184*/;
assign _282_ = _10_ & _285_ /*12180*/;
assign _283_ = _10_ ^ _285_ /*12183*/;
assign _284_ = _276_ & _283_ /*12181*/;
assign _204_ = _276_ ^ _283_ /*12182*/;
assign _281_ = _282_ | _284_ /*12179*/;
assign _290_ = D[12] ^ Q[31] /*12178*/;
assign _287_ = _11_ & _290_ /*12174*/;
assign _288_ = _11_ ^ _290_ /*12177*/;
assign _289_ = _281_ & _288_ /*12175*/;
assign _205_ = _281_ ^ _288_ /*12176*/;
assign _286_ = _287_ | _289_ /*12173*/;
assign _295_ = D[13] ^ Q[31] /*12172*/;
assign _292_ = _12_ & _295_ /*12168*/;
assign _293_ = _12_ ^ _295_ /*12171*/;
assign _294_ = _286_ & _293_ /*12169*/;
assign _206_ = _286_ ^ _293_ /*12170*/;
assign _291_ = _292_ | _294_ /*12167*/;
assign _300_ = D[14] ^ Q[31] /*12166*/;
assign _297_ = _13_ & _300_ /*12162*/;
assign _298_ = _13_ ^ _300_ /*12165*/;
assign _299_ = _291_ & _298_ /*12163*/;
assign _207_ = _291_ ^ _298_ /*12164*/;
assign _296_ = _297_ | _299_ /*12161*/;
assign _305_ = D[15] ^ Q[31] /*12160*/;
assign _302_ = _14_ & _305_ /*12156*/;
assign _303_ = _14_ ^ _305_ /*12159*/;
assign _304_ = _296_ & _303_ /*12157*/;
assign _208_ = _296_ ^ _303_ /*12158*/;
assign _301_ = _302_ | _304_ /*12155*/;
assign _310_ = D[16] ^ Q[31] /*12154*/;
assign _307_ = _15_ & _310_ /*12150*/;
assign _308_ = _15_ ^ _310_ /*12153*/;
assign _309_ = _301_ & _308_ /*12151*/;
assign _209_ = _301_ ^ _308_ /*12152*/;
assign _306_ = _307_ | _309_ /*12149*/;
assign _315_ = D[17] ^ Q[31] /*12148*/;
assign _312_ = _16_ & _315_ /*12144*/;
assign _313_ = _16_ ^ _315_ /*12147*/;
assign _314_ = _306_ & _313_ /*12145*/;
assign _210_ = _306_ ^ _313_ /*12146*/;
assign _311_ = _312_ | _314_ /*12143*/;
assign _320_ = D[18] ^ Q[31] /*12142*/;
assign _317_ = _17_ & _320_ /*12138*/;
assign _318_ = _17_ ^ _320_ /*12141*/;
assign _319_ = _311_ & _318_ /*12139*/;
assign _211_ = _311_ ^ _318_ /*12140*/;
assign _316_ = _317_ | _319_ /*12137*/;
assign _325_ = D[19] ^ Q[31] /*12136*/;
assign _322_ = _18_ & _325_ /*12132*/;
assign _323_ = _18_ ^ _325_ /*12135*/;
assign _324_ = _316_ & _323_ /*12133*/;
assign _212_ = _316_ ^ _323_ /*12134*/;
assign _321_ = _322_ | _324_ /*12131*/;
assign _330_ = D[20] ^ Q[31] /*12130*/;
assign _327_ = _19_ & _330_ /*12126*/;
assign _328_ = _19_ ^ _330_ /*12129*/;
assign _329_ = _321_ & _328_ /*12127*/;
assign _213_ = _321_ ^ _328_ /*12128*/;
assign _326_ = _327_ | _329_ /*12125*/;
assign _335_ = D[21] ^ Q[31] /*12124*/;
assign _332_ = _20_ & _335_ /*12120*/;
assign _333_ = _20_ ^ _335_ /*12123*/;
assign _334_ = _326_ & _333_ /*12121*/;
assign _214_ = _326_ ^ _333_ /*12122*/;
assign _331_ = _332_ | _334_ /*12119*/;
assign _340_ = D[22] ^ Q[31] /*12118*/;
assign _337_ = _21_ & _340_ /*12114*/;
assign _338_ = _21_ ^ _340_ /*12117*/;
assign _339_ = _331_ & _338_ /*12115*/;
assign _215_ = _331_ ^ _338_ /*12116*/;
assign _336_ = _337_ | _339_ /*12113*/;
assign _345_ = D[23] ^ Q[31] /*12112*/;
assign _342_ = _22_ & _345_ /*12108*/;
assign _343_ = _22_ ^ _345_ /*12111*/;
assign _344_ = _336_ & _343_ /*12109*/;
assign _216_ = _336_ ^ _343_ /*12110*/;
assign _341_ = _342_ | _344_ /*12107*/;
assign _350_ = D[24] ^ Q[31] /*12106*/;
assign _347_ = _23_ & _350_ /*12102*/;
assign _348_ = _23_ ^ _350_ /*12105*/;
assign _349_ = _341_ & _348_ /*12103*/;
assign _217_ = _341_ ^ _348_ /*12104*/;
assign _346_ = _347_ | _349_ /*12101*/;
assign _355_ = D[25] ^ Q[31] /*12100*/;
assign _352_ = _24_ & _355_ /*12096*/;
assign _353_ = _24_ ^ _355_ /*12099*/;
assign _354_ = _346_ & _353_ /*12097*/;
assign _218_ = _346_ ^ _353_ /*12098*/;
assign _351_ = _352_ | _354_ /*12095*/;
assign _360_ = D[26] ^ Q[31] /*12094*/;
assign _357_ = _25_ & _360_ /*12090*/;
assign _358_ = _25_ ^ _360_ /*12093*/;
assign _359_ = _351_ & _358_ /*12091*/;
assign _219_ = _351_ ^ _358_ /*12092*/;
assign _356_ = _357_ | _359_ /*12089*/;
assign _365_ = D[27] ^ Q[31] /*12088*/;
assign _362_ = _26_ & _365_ /*12084*/;
assign _363_ = _26_ ^ _365_ /*12087*/;
assign _364_ = _356_ & _363_ /*12085*/;
assign _220_ = _356_ ^ _363_ /*12086*/;
assign _361_ = _362_ | _364_ /*12083*/;
assign _370_ = D[28] ^ Q[31] /*12082*/;
assign _367_ = _27_ & _370_ /*12078*/;
assign _368_ = _27_ ^ _370_ /*12081*/;
assign _369_ = _361_ & _368_ /*12079*/;
assign _221_ = _361_ ^ _368_ /*12080*/;
assign _366_ = _367_ | _369_ /*12077*/;
assign _375_ = D[29] ^ Q[31] /*12076*/;
assign _372_ = _28_ & _375_ /*12072*/;
assign _373_ = _28_ ^ _375_ /*12075*/;
assign _374_ = _366_ & _373_ /*12073*/;
assign _222_ = _366_ ^ _373_ /*12074*/;
assign _371_ = _372_ | _374_ /*12071*/;
assign _380_ = D[30] ^ Q[31] /*12070*/;
assign _377_ = _29_ & _380_ /*12066*/;
assign _378_ = _29_ ^ _380_ /*12069*/;
assign _379_ = _371_ & _378_ /*12067*/;
assign _223_ = _371_ ^ _378_ /*12068*/;
assign _376_ = _377_ | _379_ /*12065*/;
assign _384_ = zeroWire ^ Q[31] /*12064*/;
assign _381_ = _30_ & _384_ /*12060*/;
assign _382_ = _30_ ^ _384_ /*12063*/;
assign _383_ = _376_ & _382_ /*12061*/;
assign _224_ = _376_ ^ _382_ /*12062*/;
assign Q[30] = _381_ | _383_ /*12059*/;
assign _423_ = D[0] ^ Q[30] /*11865*/;
assign _420_ = R_0[29] & _423_ /*11861*/;
assign _421_ = R_0[29] ^ _423_ /*11864*/;
assign _422_ = Q[30] & _421_ /*11862*/;
assign _386_ = Q[30] ^ _421_ /*11863*/;
assign _419_ = _420_ | _422_ /*11860*/;
assign _428_ = D[1] ^ Q[30] /*11859*/;
assign _425_ = _193_ & _428_ /*11855*/;
assign _426_ = _193_ ^ _428_ /*11858*/;
assign _427_ = _419_ & _426_ /*11856*/;
assign _387_ = _419_ ^ _426_ /*11857*/;
assign _424_ = _425_ | _427_ /*11854*/;
assign _433_ = D[2] ^ Q[30] /*11853*/;
assign _430_ = _194_ & _433_ /*11849*/;
assign _431_ = _194_ ^ _433_ /*11852*/;
assign _432_ = _424_ & _431_ /*11850*/;
assign _388_ = _424_ ^ _431_ /*11851*/;
assign _429_ = _430_ | _432_ /*11848*/;
assign _438_ = D[3] ^ Q[30] /*11847*/;
assign _435_ = _195_ & _438_ /*11843*/;
assign _436_ = _195_ ^ _438_ /*11846*/;
assign _437_ = _429_ & _436_ /*11844*/;
assign _389_ = _429_ ^ _436_ /*11845*/;
assign _434_ = _435_ | _437_ /*11842*/;
assign _443_ = D[4] ^ Q[30] /*11841*/;
assign _440_ = _196_ & _443_ /*11837*/;
assign _441_ = _196_ ^ _443_ /*11840*/;
assign _442_ = _434_ & _441_ /*11838*/;
assign _390_ = _434_ ^ _441_ /*11839*/;
assign _439_ = _440_ | _442_ /*11836*/;
assign _448_ = D[5] ^ Q[30] /*11835*/;
assign _445_ = _197_ & _448_ /*11831*/;
assign _446_ = _197_ ^ _448_ /*11834*/;
assign _447_ = _439_ & _446_ /*11832*/;
assign _391_ = _439_ ^ _446_ /*11833*/;
assign _444_ = _445_ | _447_ /*11830*/;
assign _453_ = D[6] ^ Q[30] /*11829*/;
assign _450_ = _198_ & _453_ /*11825*/;
assign _451_ = _198_ ^ _453_ /*11828*/;
assign _452_ = _444_ & _451_ /*11826*/;
assign _392_ = _444_ ^ _451_ /*11827*/;
assign _449_ = _450_ | _452_ /*11824*/;
assign _458_ = D[7] ^ Q[30] /*11823*/;
assign _455_ = _199_ & _458_ /*11819*/;
assign _456_ = _199_ ^ _458_ /*11822*/;
assign _457_ = _449_ & _456_ /*11820*/;
assign _393_ = _449_ ^ _456_ /*11821*/;
assign _454_ = _455_ | _457_ /*11818*/;
assign _463_ = D[8] ^ Q[30] /*11817*/;
assign _460_ = _200_ & _463_ /*11813*/;
assign _461_ = _200_ ^ _463_ /*11816*/;
assign _462_ = _454_ & _461_ /*11814*/;
assign _394_ = _454_ ^ _461_ /*11815*/;
assign _459_ = _460_ | _462_ /*11812*/;
assign _468_ = D[9] ^ Q[30] /*11811*/;
assign _465_ = _201_ & _468_ /*11807*/;
assign _466_ = _201_ ^ _468_ /*11810*/;
assign _467_ = _459_ & _466_ /*11808*/;
assign _395_ = _459_ ^ _466_ /*11809*/;
assign _464_ = _465_ | _467_ /*11806*/;
assign _473_ = D[10] ^ Q[30] /*11805*/;
assign _470_ = _202_ & _473_ /*11801*/;
assign _471_ = _202_ ^ _473_ /*11804*/;
assign _472_ = _464_ & _471_ /*11802*/;
assign _396_ = _464_ ^ _471_ /*11803*/;
assign _469_ = _470_ | _472_ /*11800*/;
assign _478_ = D[11] ^ Q[30] /*11799*/;
assign _475_ = _203_ & _478_ /*11795*/;
assign _476_ = _203_ ^ _478_ /*11798*/;
assign _477_ = _469_ & _476_ /*11796*/;
assign _397_ = _469_ ^ _476_ /*11797*/;
assign _474_ = _475_ | _477_ /*11794*/;
assign _483_ = D[12] ^ Q[30] /*11793*/;
assign _480_ = _204_ & _483_ /*11789*/;
assign _481_ = _204_ ^ _483_ /*11792*/;
assign _482_ = _474_ & _481_ /*11790*/;
assign _398_ = _474_ ^ _481_ /*11791*/;
assign _479_ = _480_ | _482_ /*11788*/;
assign _488_ = D[13] ^ Q[30] /*11787*/;
assign _485_ = _205_ & _488_ /*11783*/;
assign _486_ = _205_ ^ _488_ /*11786*/;
assign _487_ = _479_ & _486_ /*11784*/;
assign _399_ = _479_ ^ _486_ /*11785*/;
assign _484_ = _485_ | _487_ /*11782*/;
assign _493_ = D[14] ^ Q[30] /*11781*/;
assign _490_ = _206_ & _493_ /*11777*/;
assign _491_ = _206_ ^ _493_ /*11780*/;
assign _492_ = _484_ & _491_ /*11778*/;
assign _400_ = _484_ ^ _491_ /*11779*/;
assign _489_ = _490_ | _492_ /*11776*/;
assign _498_ = D[15] ^ Q[30] /*11775*/;
assign _495_ = _207_ & _498_ /*11771*/;
assign _496_ = _207_ ^ _498_ /*11774*/;
assign _497_ = _489_ & _496_ /*11772*/;
assign _401_ = _489_ ^ _496_ /*11773*/;
assign _494_ = _495_ | _497_ /*11770*/;
assign _503_ = D[16] ^ Q[30] /*11769*/;
assign _500_ = _208_ & _503_ /*11765*/;
assign _501_ = _208_ ^ _503_ /*11768*/;
assign _502_ = _494_ & _501_ /*11766*/;
assign _402_ = _494_ ^ _501_ /*11767*/;
assign _499_ = _500_ | _502_ /*11764*/;
assign _508_ = D[17] ^ Q[30] /*11763*/;
assign _505_ = _209_ & _508_ /*11759*/;
assign _506_ = _209_ ^ _508_ /*11762*/;
assign _507_ = _499_ & _506_ /*11760*/;
assign _403_ = _499_ ^ _506_ /*11761*/;
assign _504_ = _505_ | _507_ /*11758*/;
assign _513_ = D[18] ^ Q[30] /*11757*/;
assign _510_ = _210_ & _513_ /*11753*/;
assign _511_ = _210_ ^ _513_ /*11756*/;
assign _512_ = _504_ & _511_ /*11754*/;
assign _404_ = _504_ ^ _511_ /*11755*/;
assign _509_ = _510_ | _512_ /*11752*/;
assign _518_ = D[19] ^ Q[30] /*11751*/;
assign _515_ = _211_ & _518_ /*11747*/;
assign _516_ = _211_ ^ _518_ /*11750*/;
assign _517_ = _509_ & _516_ /*11748*/;
assign _405_ = _509_ ^ _516_ /*11749*/;
assign _514_ = _515_ | _517_ /*11746*/;
assign _523_ = D[20] ^ Q[30] /*11745*/;
assign _520_ = _212_ & _523_ /*11741*/;
assign _521_ = _212_ ^ _523_ /*11744*/;
assign _522_ = _514_ & _521_ /*11742*/;
assign _406_ = _514_ ^ _521_ /*11743*/;
assign _519_ = _520_ | _522_ /*11740*/;
assign _528_ = D[21] ^ Q[30] /*11739*/;
assign _525_ = _213_ & _528_ /*11735*/;
assign _526_ = _213_ ^ _528_ /*11738*/;
assign _527_ = _519_ & _526_ /*11736*/;
assign _407_ = _519_ ^ _526_ /*11737*/;
assign _524_ = _525_ | _527_ /*11734*/;
assign _533_ = D[22] ^ Q[30] /*11733*/;
assign _530_ = _214_ & _533_ /*11729*/;
assign _531_ = _214_ ^ _533_ /*11732*/;
assign _532_ = _524_ & _531_ /*11730*/;
assign _408_ = _524_ ^ _531_ /*11731*/;
assign _529_ = _530_ | _532_ /*11728*/;
assign _538_ = D[23] ^ Q[30] /*11727*/;
assign _535_ = _215_ & _538_ /*11723*/;
assign _536_ = _215_ ^ _538_ /*11726*/;
assign _537_ = _529_ & _536_ /*11724*/;
assign _409_ = _529_ ^ _536_ /*11725*/;
assign _534_ = _535_ | _537_ /*11722*/;
assign _543_ = D[24] ^ Q[30] /*11721*/;
assign _540_ = _216_ & _543_ /*11717*/;
assign _541_ = _216_ ^ _543_ /*11720*/;
assign _542_ = _534_ & _541_ /*11718*/;
assign _410_ = _534_ ^ _541_ /*11719*/;
assign _539_ = _540_ | _542_ /*11716*/;
assign _548_ = D[25] ^ Q[30] /*11715*/;
assign _545_ = _217_ & _548_ /*11711*/;
assign _546_ = _217_ ^ _548_ /*11714*/;
assign _547_ = _539_ & _546_ /*11712*/;
assign _411_ = _539_ ^ _546_ /*11713*/;
assign _544_ = _545_ | _547_ /*11710*/;
assign _553_ = D[26] ^ Q[30] /*11709*/;
assign _550_ = _218_ & _553_ /*11705*/;
assign _551_ = _218_ ^ _553_ /*11708*/;
assign _552_ = _544_ & _551_ /*11706*/;
assign _412_ = _544_ ^ _551_ /*11707*/;
assign _549_ = _550_ | _552_ /*11704*/;
assign _558_ = D[27] ^ Q[30] /*11703*/;
assign _555_ = _219_ & _558_ /*11699*/;
assign _556_ = _219_ ^ _558_ /*11702*/;
assign _557_ = _549_ & _556_ /*11700*/;
assign _413_ = _549_ ^ _556_ /*11701*/;
assign _554_ = _555_ | _557_ /*11698*/;
assign _563_ = D[28] ^ Q[30] /*11697*/;
assign _560_ = _220_ & _563_ /*11693*/;
assign _561_ = _220_ ^ _563_ /*11696*/;
assign _562_ = _554_ & _561_ /*11694*/;
assign _414_ = _554_ ^ _561_ /*11695*/;
assign _559_ = _560_ | _562_ /*11692*/;
assign _568_ = D[29] ^ Q[30] /*11691*/;
assign _565_ = _221_ & _568_ /*11687*/;
assign _566_ = _221_ ^ _568_ /*11690*/;
assign _567_ = _559_ & _566_ /*11688*/;
assign _415_ = _559_ ^ _566_ /*11689*/;
assign _564_ = _565_ | _567_ /*11686*/;
assign _573_ = D[30] ^ Q[30] /*11685*/;
assign _570_ = _222_ & _573_ /*11681*/;
assign _571_ = _222_ ^ _573_ /*11684*/;
assign _572_ = _564_ & _571_ /*11682*/;
assign _416_ = _564_ ^ _571_ /*11683*/;
assign _569_ = _570_ | _572_ /*11680*/;
assign _577_ = zeroWire ^ Q[30] /*11679*/;
assign _574_ = _223_ & _577_ /*11675*/;
assign _575_ = _223_ ^ _577_ /*11678*/;
assign _576_ = _569_ & _575_ /*11676*/;
assign _417_ = _569_ ^ _575_ /*11677*/;
assign Q[29] = _574_ | _576_ /*11674*/;
assign _616_ = D[0] ^ Q[29] /*11480*/;
assign _613_ = R_0[28] & _616_ /*11476*/;
assign _614_ = R_0[28] ^ _616_ /*11479*/;
assign _615_ = Q[29] & _614_ /*11477*/;
assign _579_ = Q[29] ^ _614_ /*11478*/;
assign _612_ = _613_ | _615_ /*11475*/;
assign _621_ = D[1] ^ Q[29] /*11474*/;
assign _618_ = _386_ & _621_ /*11470*/;
assign _619_ = _386_ ^ _621_ /*11473*/;
assign _620_ = _612_ & _619_ /*11471*/;
assign _580_ = _612_ ^ _619_ /*11472*/;
assign _617_ = _618_ | _620_ /*11469*/;
assign _626_ = D[2] ^ Q[29] /*11468*/;
assign _623_ = _387_ & _626_ /*11464*/;
assign _624_ = _387_ ^ _626_ /*11467*/;
assign _625_ = _617_ & _624_ /*11465*/;
assign _581_ = _617_ ^ _624_ /*11466*/;
assign _622_ = _623_ | _625_ /*11463*/;
assign _631_ = D[3] ^ Q[29] /*11462*/;
assign _628_ = _388_ & _631_ /*11458*/;
assign _629_ = _388_ ^ _631_ /*11461*/;
assign _630_ = _622_ & _629_ /*11459*/;
assign _582_ = _622_ ^ _629_ /*11460*/;
assign _627_ = _628_ | _630_ /*11457*/;
assign _636_ = D[4] ^ Q[29] /*11456*/;
assign _633_ = _389_ & _636_ /*11452*/;
assign _634_ = _389_ ^ _636_ /*11455*/;
assign _635_ = _627_ & _634_ /*11453*/;
assign _583_ = _627_ ^ _634_ /*11454*/;
assign _632_ = _633_ | _635_ /*11451*/;
assign _641_ = D[5] ^ Q[29] /*11450*/;
assign _638_ = _390_ & _641_ /*11446*/;
assign _639_ = _390_ ^ _641_ /*11449*/;
assign _640_ = _632_ & _639_ /*11447*/;
assign _584_ = _632_ ^ _639_ /*11448*/;
assign _637_ = _638_ | _640_ /*11445*/;
assign _646_ = D[6] ^ Q[29] /*11444*/;
assign _643_ = _391_ & _646_ /*11440*/;
assign _644_ = _391_ ^ _646_ /*11443*/;
assign _645_ = _637_ & _644_ /*11441*/;
assign _585_ = _637_ ^ _644_ /*11442*/;
assign _642_ = _643_ | _645_ /*11439*/;
assign _651_ = D[7] ^ Q[29] /*11438*/;
assign _648_ = _392_ & _651_ /*11434*/;
assign _649_ = _392_ ^ _651_ /*11437*/;
assign _650_ = _642_ & _649_ /*11435*/;
assign _586_ = _642_ ^ _649_ /*11436*/;
assign _647_ = _648_ | _650_ /*11433*/;
assign _656_ = D[8] ^ Q[29] /*11432*/;
assign _653_ = _393_ & _656_ /*11428*/;
assign _654_ = _393_ ^ _656_ /*11431*/;
assign _655_ = _647_ & _654_ /*11429*/;
assign _587_ = _647_ ^ _654_ /*11430*/;
assign _652_ = _653_ | _655_ /*11427*/;
assign _661_ = D[9] ^ Q[29] /*11426*/;
assign _658_ = _394_ & _661_ /*11422*/;
assign _659_ = _394_ ^ _661_ /*11425*/;
assign _660_ = _652_ & _659_ /*11423*/;
assign _588_ = _652_ ^ _659_ /*11424*/;
assign _657_ = _658_ | _660_ /*11421*/;
assign _666_ = D[10] ^ Q[29] /*11420*/;
assign _663_ = _395_ & _666_ /*11416*/;
assign _664_ = _395_ ^ _666_ /*11419*/;
assign _665_ = _657_ & _664_ /*11417*/;
assign _589_ = _657_ ^ _664_ /*11418*/;
assign _662_ = _663_ | _665_ /*11415*/;
assign _671_ = D[11] ^ Q[29] /*11414*/;
assign _668_ = _396_ & _671_ /*11410*/;
assign _669_ = _396_ ^ _671_ /*11413*/;
assign _670_ = _662_ & _669_ /*11411*/;
assign _590_ = _662_ ^ _669_ /*11412*/;
assign _667_ = _668_ | _670_ /*11409*/;
assign _676_ = D[12] ^ Q[29] /*11408*/;
assign _673_ = _397_ & _676_ /*11404*/;
assign _674_ = _397_ ^ _676_ /*11407*/;
assign _675_ = _667_ & _674_ /*11405*/;
assign _591_ = _667_ ^ _674_ /*11406*/;
assign _672_ = _673_ | _675_ /*11403*/;
assign _681_ = D[13] ^ Q[29] /*11402*/;
assign _678_ = _398_ & _681_ /*11398*/;
assign _679_ = _398_ ^ _681_ /*11401*/;
assign _680_ = _672_ & _679_ /*11399*/;
assign _592_ = _672_ ^ _679_ /*11400*/;
assign _677_ = _678_ | _680_ /*11397*/;
assign _686_ = D[14] ^ Q[29] /*11396*/;
assign _683_ = _399_ & _686_ /*11392*/;
assign _684_ = _399_ ^ _686_ /*11395*/;
assign _685_ = _677_ & _684_ /*11393*/;
assign _593_ = _677_ ^ _684_ /*11394*/;
assign _682_ = _683_ | _685_ /*11391*/;
assign _691_ = D[15] ^ Q[29] /*11390*/;
assign _688_ = _400_ & _691_ /*11386*/;
assign _689_ = _400_ ^ _691_ /*11389*/;
assign _690_ = _682_ & _689_ /*11387*/;
assign _594_ = _682_ ^ _689_ /*11388*/;
assign _687_ = _688_ | _690_ /*11385*/;
assign _696_ = D[16] ^ Q[29] /*11384*/;
assign _693_ = _401_ & _696_ /*11380*/;
assign _694_ = _401_ ^ _696_ /*11383*/;
assign _695_ = _687_ & _694_ /*11381*/;
assign _595_ = _687_ ^ _694_ /*11382*/;
assign _692_ = _693_ | _695_ /*11379*/;
assign _701_ = D[17] ^ Q[29] /*11378*/;
assign _698_ = _402_ & _701_ /*11374*/;
assign _699_ = _402_ ^ _701_ /*11377*/;
assign _700_ = _692_ & _699_ /*11375*/;
assign _596_ = _692_ ^ _699_ /*11376*/;
assign _697_ = _698_ | _700_ /*11373*/;
assign _706_ = D[18] ^ Q[29] /*11372*/;
assign _703_ = _403_ & _706_ /*11368*/;
assign _704_ = _403_ ^ _706_ /*11371*/;
assign _705_ = _697_ & _704_ /*11369*/;
assign _597_ = _697_ ^ _704_ /*11370*/;
assign _702_ = _703_ | _705_ /*11367*/;
assign _711_ = D[19] ^ Q[29] /*11366*/;
assign _708_ = _404_ & _711_ /*11362*/;
assign _709_ = _404_ ^ _711_ /*11365*/;
assign _710_ = _702_ & _709_ /*11363*/;
assign _598_ = _702_ ^ _709_ /*11364*/;
assign _707_ = _708_ | _710_ /*11361*/;
assign _716_ = D[20] ^ Q[29] /*11360*/;
assign _713_ = _405_ & _716_ /*11356*/;
assign _714_ = _405_ ^ _716_ /*11359*/;
assign _715_ = _707_ & _714_ /*11357*/;
assign _599_ = _707_ ^ _714_ /*11358*/;
assign _712_ = _713_ | _715_ /*11355*/;
assign _721_ = D[21] ^ Q[29] /*11354*/;
assign _718_ = _406_ & _721_ /*11350*/;
assign _719_ = _406_ ^ _721_ /*11353*/;
assign _720_ = _712_ & _719_ /*11351*/;
assign _600_ = _712_ ^ _719_ /*11352*/;
assign _717_ = _718_ | _720_ /*11349*/;
assign _726_ = D[22] ^ Q[29] /*11348*/;
assign _723_ = _407_ & _726_ /*11344*/;
assign _724_ = _407_ ^ _726_ /*11347*/;
assign _725_ = _717_ & _724_ /*11345*/;
assign _601_ = _717_ ^ _724_ /*11346*/;
assign _722_ = _723_ | _725_ /*11343*/;
assign _731_ = D[23] ^ Q[29] /*11342*/;
assign _728_ = _408_ & _731_ /*11338*/;
assign _729_ = _408_ ^ _731_ /*11341*/;
assign _730_ = _722_ & _729_ /*11339*/;
assign _602_ = _722_ ^ _729_ /*11340*/;
assign _727_ = _728_ | _730_ /*11337*/;
assign _736_ = D[24] ^ Q[29] /*11336*/;
assign _733_ = _409_ & _736_ /*11332*/;
assign _734_ = _409_ ^ _736_ /*11335*/;
assign _735_ = _727_ & _734_ /*11333*/;
assign _603_ = _727_ ^ _734_ /*11334*/;
assign _732_ = _733_ | _735_ /*11331*/;
assign _741_ = D[25] ^ Q[29] /*11330*/;
assign _738_ = _410_ & _741_ /*11326*/;
assign _739_ = _410_ ^ _741_ /*11329*/;
assign _740_ = _732_ & _739_ /*11327*/;
assign _604_ = _732_ ^ _739_ /*11328*/;
assign _737_ = _738_ | _740_ /*11325*/;
assign _746_ = D[26] ^ Q[29] /*11324*/;
assign _743_ = _411_ & _746_ /*11320*/;
assign _744_ = _411_ ^ _746_ /*11323*/;
assign _745_ = _737_ & _744_ /*11321*/;
assign _605_ = _737_ ^ _744_ /*11322*/;
assign _742_ = _743_ | _745_ /*11319*/;
assign _751_ = D[27] ^ Q[29] /*11318*/;
assign _748_ = _412_ & _751_ /*11314*/;
assign _749_ = _412_ ^ _751_ /*11317*/;
assign _750_ = _742_ & _749_ /*11315*/;
assign _606_ = _742_ ^ _749_ /*11316*/;
assign _747_ = _748_ | _750_ /*11313*/;
assign _756_ = D[28] ^ Q[29] /*11312*/;
assign _753_ = _413_ & _756_ /*11308*/;
assign _754_ = _413_ ^ _756_ /*11311*/;
assign _755_ = _747_ & _754_ /*11309*/;
assign _607_ = _747_ ^ _754_ /*11310*/;
assign _752_ = _753_ | _755_ /*11307*/;
assign _761_ = D[29] ^ Q[29] /*11306*/;
assign _758_ = _414_ & _761_ /*11302*/;
assign _759_ = _414_ ^ _761_ /*11305*/;
assign _760_ = _752_ & _759_ /*11303*/;
assign _608_ = _752_ ^ _759_ /*11304*/;
assign _757_ = _758_ | _760_ /*11301*/;
assign _766_ = D[30] ^ Q[29] /*11300*/;
assign _763_ = _415_ & _766_ /*11296*/;
assign _764_ = _415_ ^ _766_ /*11299*/;
assign _765_ = _757_ & _764_ /*11297*/;
assign _609_ = _757_ ^ _764_ /*11298*/;
assign _762_ = _763_ | _765_ /*11295*/;
assign _770_ = zeroWire ^ Q[29] /*11294*/;
assign _767_ = _416_ & _770_ /*11290*/;
assign _768_ = _416_ ^ _770_ /*11293*/;
assign _769_ = _762_ & _768_ /*11291*/;
assign _610_ = _762_ ^ _768_ /*11292*/;
assign Q[28] = _767_ | _769_ /*11289*/;
assign _809_ = D[0] ^ Q[28] /*11095*/;
assign _806_ = R_0[27] & _809_ /*11091*/;
assign _807_ = R_0[27] ^ _809_ /*11094*/;
assign _808_ = Q[28] & _807_ /*11092*/;
assign _772_ = Q[28] ^ _807_ /*11093*/;
assign _805_ = _806_ | _808_ /*11090*/;
assign _814_ = D[1] ^ Q[28] /*11089*/;
assign _811_ = _579_ & _814_ /*11085*/;
assign _812_ = _579_ ^ _814_ /*11088*/;
assign _813_ = _805_ & _812_ /*11086*/;
assign _773_ = _805_ ^ _812_ /*11087*/;
assign _810_ = _811_ | _813_ /*11084*/;
assign _819_ = D[2] ^ Q[28] /*11083*/;
assign _816_ = _580_ & _819_ /*11079*/;
assign _817_ = _580_ ^ _819_ /*11082*/;
assign _818_ = _810_ & _817_ /*11080*/;
assign _774_ = _810_ ^ _817_ /*11081*/;
assign _815_ = _816_ | _818_ /*11078*/;
assign _824_ = D[3] ^ Q[28] /*11077*/;
assign _821_ = _581_ & _824_ /*11073*/;
assign _822_ = _581_ ^ _824_ /*11076*/;
assign _823_ = _815_ & _822_ /*11074*/;
assign _775_ = _815_ ^ _822_ /*11075*/;
assign _820_ = _821_ | _823_ /*11072*/;
assign _829_ = D[4] ^ Q[28] /*11071*/;
assign _826_ = _582_ & _829_ /*11067*/;
assign _827_ = _582_ ^ _829_ /*11070*/;
assign _828_ = _820_ & _827_ /*11068*/;
assign _776_ = _820_ ^ _827_ /*11069*/;
assign _825_ = _826_ | _828_ /*11066*/;
assign _834_ = D[5] ^ Q[28] /*11065*/;
assign _831_ = _583_ & _834_ /*11061*/;
assign _832_ = _583_ ^ _834_ /*11064*/;
assign _833_ = _825_ & _832_ /*11062*/;
assign _777_ = _825_ ^ _832_ /*11063*/;
assign _830_ = _831_ | _833_ /*11060*/;
assign _839_ = D[6] ^ Q[28] /*11059*/;
assign _836_ = _584_ & _839_ /*11055*/;
assign _837_ = _584_ ^ _839_ /*11058*/;
assign _838_ = _830_ & _837_ /*11056*/;
assign _778_ = _830_ ^ _837_ /*11057*/;
assign _835_ = _836_ | _838_ /*11054*/;
assign _844_ = D[7] ^ Q[28] /*11053*/;
assign _841_ = _585_ & _844_ /*11049*/;
assign _842_ = _585_ ^ _844_ /*11052*/;
assign _843_ = _835_ & _842_ /*11050*/;
assign _779_ = _835_ ^ _842_ /*11051*/;
assign _840_ = _841_ | _843_ /*11048*/;
assign _849_ = D[8] ^ Q[28] /*11047*/;
assign _846_ = _586_ & _849_ /*11043*/;
assign _847_ = _586_ ^ _849_ /*11046*/;
assign _848_ = _840_ & _847_ /*11044*/;
assign _780_ = _840_ ^ _847_ /*11045*/;
assign _845_ = _846_ | _848_ /*11042*/;
assign _854_ = D[9] ^ Q[28] /*11041*/;
assign _851_ = _587_ & _854_ /*11037*/;
assign _852_ = _587_ ^ _854_ /*11040*/;
assign _853_ = _845_ & _852_ /*11038*/;
assign _781_ = _845_ ^ _852_ /*11039*/;
assign _850_ = _851_ | _853_ /*11036*/;
assign _859_ = D[10] ^ Q[28] /*11035*/;
assign _856_ = _588_ & _859_ /*11031*/;
assign _857_ = _588_ ^ _859_ /*11034*/;
assign _858_ = _850_ & _857_ /*11032*/;
assign _782_ = _850_ ^ _857_ /*11033*/;
assign _855_ = _856_ | _858_ /*11030*/;
assign _864_ = D[11] ^ Q[28] /*11029*/;
assign _861_ = _589_ & _864_ /*11025*/;
assign _862_ = _589_ ^ _864_ /*11028*/;
assign _863_ = _855_ & _862_ /*11026*/;
assign _783_ = _855_ ^ _862_ /*11027*/;
assign _860_ = _861_ | _863_ /*11024*/;
assign _869_ = D[12] ^ Q[28] /*11023*/;
assign _866_ = _590_ & _869_ /*11019*/;
assign _867_ = _590_ ^ _869_ /*11022*/;
assign _868_ = _860_ & _867_ /*11020*/;
assign _784_ = _860_ ^ _867_ /*11021*/;
assign _865_ = _866_ | _868_ /*11018*/;
assign _874_ = D[13] ^ Q[28] /*11017*/;
assign _871_ = _591_ & _874_ /*11013*/;
assign _872_ = _591_ ^ _874_ /*11016*/;
assign _873_ = _865_ & _872_ /*11014*/;
assign _785_ = _865_ ^ _872_ /*11015*/;
assign _870_ = _871_ | _873_ /*11012*/;
assign _879_ = D[14] ^ Q[28] /*11011*/;
assign _876_ = _592_ & _879_ /*11007*/;
assign _877_ = _592_ ^ _879_ /*11010*/;
assign _878_ = _870_ & _877_ /*11008*/;
assign _786_ = _870_ ^ _877_ /*11009*/;
assign _875_ = _876_ | _878_ /*11006*/;
assign _884_ = D[15] ^ Q[28] /*11005*/;
assign _881_ = _593_ & _884_ /*11001*/;
assign _882_ = _593_ ^ _884_ /*11004*/;
assign _883_ = _875_ & _882_ /*11002*/;
assign _787_ = _875_ ^ _882_ /*11003*/;
assign _880_ = _881_ | _883_ /*11000*/;
assign _889_ = D[16] ^ Q[28] /*10999*/;
assign _886_ = _594_ & _889_ /*10995*/;
assign _887_ = _594_ ^ _889_ /*10998*/;
assign _888_ = _880_ & _887_ /*10996*/;
assign _788_ = _880_ ^ _887_ /*10997*/;
assign _885_ = _886_ | _888_ /*10994*/;
assign _894_ = D[17] ^ Q[28] /*10993*/;
assign _891_ = _595_ & _894_ /*10989*/;
assign _892_ = _595_ ^ _894_ /*10992*/;
assign _893_ = _885_ & _892_ /*10990*/;
assign _789_ = _885_ ^ _892_ /*10991*/;
assign _890_ = _891_ | _893_ /*10988*/;
assign _899_ = D[18] ^ Q[28] /*10987*/;
assign _896_ = _596_ & _899_ /*10983*/;
assign _897_ = _596_ ^ _899_ /*10986*/;
assign _898_ = _890_ & _897_ /*10984*/;
assign _790_ = _890_ ^ _897_ /*10985*/;
assign _895_ = _896_ | _898_ /*10982*/;
assign _904_ = D[19] ^ Q[28] /*10981*/;
assign _901_ = _597_ & _904_ /*10977*/;
assign _902_ = _597_ ^ _904_ /*10980*/;
assign _903_ = _895_ & _902_ /*10978*/;
assign _791_ = _895_ ^ _902_ /*10979*/;
assign _900_ = _901_ | _903_ /*10976*/;
assign _909_ = D[20] ^ Q[28] /*10975*/;
assign _906_ = _598_ & _909_ /*10971*/;
assign _907_ = _598_ ^ _909_ /*10974*/;
assign _908_ = _900_ & _907_ /*10972*/;
assign _792_ = _900_ ^ _907_ /*10973*/;
assign _905_ = _906_ | _908_ /*10970*/;
assign _914_ = D[21] ^ Q[28] /*10969*/;
assign _911_ = _599_ & _914_ /*10965*/;
assign _912_ = _599_ ^ _914_ /*10968*/;
assign _913_ = _905_ & _912_ /*10966*/;
assign _793_ = _905_ ^ _912_ /*10967*/;
assign _910_ = _911_ | _913_ /*10964*/;
assign _919_ = D[22] ^ Q[28] /*10963*/;
assign _916_ = _600_ & _919_ /*10959*/;
assign _917_ = _600_ ^ _919_ /*10962*/;
assign _918_ = _910_ & _917_ /*10960*/;
assign _794_ = _910_ ^ _917_ /*10961*/;
assign _915_ = _916_ | _918_ /*10958*/;
assign _924_ = D[23] ^ Q[28] /*10957*/;
assign _921_ = _601_ & _924_ /*10953*/;
assign _922_ = _601_ ^ _924_ /*10956*/;
assign _923_ = _915_ & _922_ /*10954*/;
assign _795_ = _915_ ^ _922_ /*10955*/;
assign _920_ = _921_ | _923_ /*10952*/;
assign _929_ = D[24] ^ Q[28] /*10951*/;
assign _926_ = _602_ & _929_ /*10947*/;
assign _927_ = _602_ ^ _929_ /*10950*/;
assign _928_ = _920_ & _927_ /*10948*/;
assign _796_ = _920_ ^ _927_ /*10949*/;
assign _925_ = _926_ | _928_ /*10946*/;
assign _934_ = D[25] ^ Q[28] /*10945*/;
assign _931_ = _603_ & _934_ /*10941*/;
assign _932_ = _603_ ^ _934_ /*10944*/;
assign _933_ = _925_ & _932_ /*10942*/;
assign _797_ = _925_ ^ _932_ /*10943*/;
assign _930_ = _931_ | _933_ /*10940*/;
assign _939_ = D[26] ^ Q[28] /*10939*/;
assign _936_ = _604_ & _939_ /*10935*/;
assign _937_ = _604_ ^ _939_ /*10938*/;
assign _938_ = _930_ & _937_ /*10936*/;
assign _798_ = _930_ ^ _937_ /*10937*/;
assign _935_ = _936_ | _938_ /*10934*/;
assign _944_ = D[27] ^ Q[28] /*10933*/;
assign _941_ = _605_ & _944_ /*10929*/;
assign _942_ = _605_ ^ _944_ /*10932*/;
assign _943_ = _935_ & _942_ /*10930*/;
assign _799_ = _935_ ^ _942_ /*10931*/;
assign _940_ = _941_ | _943_ /*10928*/;
assign _949_ = D[28] ^ Q[28] /*10927*/;
assign _946_ = _606_ & _949_ /*10923*/;
assign _947_ = _606_ ^ _949_ /*10926*/;
assign _948_ = _940_ & _947_ /*10924*/;
assign _800_ = _940_ ^ _947_ /*10925*/;
assign _945_ = _946_ | _948_ /*10922*/;
assign _954_ = D[29] ^ Q[28] /*10921*/;
assign _951_ = _607_ & _954_ /*10917*/;
assign _952_ = _607_ ^ _954_ /*10920*/;
assign _953_ = _945_ & _952_ /*10918*/;
assign _801_ = _945_ ^ _952_ /*10919*/;
assign _950_ = _951_ | _953_ /*10916*/;
assign _959_ = D[30] ^ Q[28] /*10915*/;
assign _956_ = _608_ & _959_ /*10911*/;
assign _957_ = _608_ ^ _959_ /*10914*/;
assign _958_ = _950_ & _957_ /*10912*/;
assign _802_ = _950_ ^ _957_ /*10913*/;
assign _955_ = _956_ | _958_ /*10910*/;
assign _963_ = zeroWire ^ Q[28] /*10909*/;
assign _960_ = _609_ & _963_ /*10905*/;
assign _961_ = _609_ ^ _963_ /*10908*/;
assign _962_ = _955_ & _961_ /*10906*/;
assign _803_ = _955_ ^ _961_ /*10907*/;
assign Q[27] = _960_ | _962_ /*10904*/;
assign _1002_ = D[0] ^ Q[27] /*10710*/;
assign _999_ = R_0[26] & _1002_ /*10706*/;
assign _1000_ = R_0[26] ^ _1002_ /*10709*/;
assign _1001_ = Q[27] & _1000_ /*10707*/;
assign _965_ = Q[27] ^ _1000_ /*10708*/;
assign _998_ = _999_ | _1001_ /*10705*/;
assign _1007_ = D[1] ^ Q[27] /*10704*/;
assign _1004_ = _772_ & _1007_ /*10700*/;
assign _1005_ = _772_ ^ _1007_ /*10703*/;
assign _1006_ = _998_ & _1005_ /*10701*/;
assign _966_ = _998_ ^ _1005_ /*10702*/;
assign _1003_ = _1004_ | _1006_ /*10699*/;
assign _1012_ = D[2] ^ Q[27] /*10698*/;
assign _1009_ = _773_ & _1012_ /*10694*/;
assign _1010_ = _773_ ^ _1012_ /*10697*/;
assign _1011_ = _1003_ & _1010_ /*10695*/;
assign _967_ = _1003_ ^ _1010_ /*10696*/;
assign _1008_ = _1009_ | _1011_ /*10693*/;
assign _1017_ = D[3] ^ Q[27] /*10692*/;
assign _1014_ = _774_ & _1017_ /*10688*/;
assign _1015_ = _774_ ^ _1017_ /*10691*/;
assign _1016_ = _1008_ & _1015_ /*10689*/;
assign _968_ = _1008_ ^ _1015_ /*10690*/;
assign _1013_ = _1014_ | _1016_ /*10687*/;
assign _1022_ = D[4] ^ Q[27] /*10686*/;
assign _1019_ = _775_ & _1022_ /*10682*/;
assign _1020_ = _775_ ^ _1022_ /*10685*/;
assign _1021_ = _1013_ & _1020_ /*10683*/;
assign _969_ = _1013_ ^ _1020_ /*10684*/;
assign _1018_ = _1019_ | _1021_ /*10681*/;
assign _1027_ = D[5] ^ Q[27] /*10680*/;
assign _1024_ = _776_ & _1027_ /*10676*/;
assign _1025_ = _776_ ^ _1027_ /*10679*/;
assign _1026_ = _1018_ & _1025_ /*10677*/;
assign _970_ = _1018_ ^ _1025_ /*10678*/;
assign _1023_ = _1024_ | _1026_ /*10675*/;
assign _1032_ = D[6] ^ Q[27] /*10674*/;
assign _1029_ = _777_ & _1032_ /*10670*/;
assign _1030_ = _777_ ^ _1032_ /*10673*/;
assign _1031_ = _1023_ & _1030_ /*10671*/;
assign _971_ = _1023_ ^ _1030_ /*10672*/;
assign _1028_ = _1029_ | _1031_ /*10669*/;
assign _1037_ = D[7] ^ Q[27] /*10668*/;
assign _1034_ = _778_ & _1037_ /*10664*/;
assign _1035_ = _778_ ^ _1037_ /*10667*/;
assign _1036_ = _1028_ & _1035_ /*10665*/;
assign _972_ = _1028_ ^ _1035_ /*10666*/;
assign _1033_ = _1034_ | _1036_ /*10663*/;
assign _1042_ = D[8] ^ Q[27] /*10662*/;
assign _1039_ = _779_ & _1042_ /*10658*/;
assign _1040_ = _779_ ^ _1042_ /*10661*/;
assign _1041_ = _1033_ & _1040_ /*10659*/;
assign _973_ = _1033_ ^ _1040_ /*10660*/;
assign _1038_ = _1039_ | _1041_ /*10657*/;
assign _1047_ = D[9] ^ Q[27] /*10656*/;
assign _1044_ = _780_ & _1047_ /*10652*/;
assign _1045_ = _780_ ^ _1047_ /*10655*/;
assign _1046_ = _1038_ & _1045_ /*10653*/;
assign _974_ = _1038_ ^ _1045_ /*10654*/;
assign _1043_ = _1044_ | _1046_ /*10651*/;
assign _1052_ = D[10] ^ Q[27] /*10650*/;
assign _1049_ = _781_ & _1052_ /*10646*/;
assign _1050_ = _781_ ^ _1052_ /*10649*/;
assign _1051_ = _1043_ & _1050_ /*10647*/;
assign _975_ = _1043_ ^ _1050_ /*10648*/;
assign _1048_ = _1049_ | _1051_ /*10645*/;
assign _1057_ = D[11] ^ Q[27] /*10644*/;
assign _1054_ = _782_ & _1057_ /*10640*/;
assign _1055_ = _782_ ^ _1057_ /*10643*/;
assign _1056_ = _1048_ & _1055_ /*10641*/;
assign _976_ = _1048_ ^ _1055_ /*10642*/;
assign _1053_ = _1054_ | _1056_ /*10639*/;
assign _1062_ = D[12] ^ Q[27] /*10638*/;
assign _1059_ = _783_ & _1062_ /*10634*/;
assign _1060_ = _783_ ^ _1062_ /*10637*/;
assign _1061_ = _1053_ & _1060_ /*10635*/;
assign _977_ = _1053_ ^ _1060_ /*10636*/;
assign _1058_ = _1059_ | _1061_ /*10633*/;
assign _1067_ = D[13] ^ Q[27] /*10632*/;
assign _1064_ = _784_ & _1067_ /*10628*/;
assign _1065_ = _784_ ^ _1067_ /*10631*/;
assign _1066_ = _1058_ & _1065_ /*10629*/;
assign _978_ = _1058_ ^ _1065_ /*10630*/;
assign _1063_ = _1064_ | _1066_ /*10627*/;
assign _1072_ = D[14] ^ Q[27] /*10626*/;
assign _1069_ = _785_ & _1072_ /*10622*/;
assign _1070_ = _785_ ^ _1072_ /*10625*/;
assign _1071_ = _1063_ & _1070_ /*10623*/;
assign _979_ = _1063_ ^ _1070_ /*10624*/;
assign _1068_ = _1069_ | _1071_ /*10621*/;
assign _1077_ = D[15] ^ Q[27] /*10620*/;
assign _1074_ = _786_ & _1077_ /*10616*/;
assign _1075_ = _786_ ^ _1077_ /*10619*/;
assign _1076_ = _1068_ & _1075_ /*10617*/;
assign _980_ = _1068_ ^ _1075_ /*10618*/;
assign _1073_ = _1074_ | _1076_ /*10615*/;
assign _1082_ = D[16] ^ Q[27] /*10614*/;
assign _1079_ = _787_ & _1082_ /*10610*/;
assign _1080_ = _787_ ^ _1082_ /*10613*/;
assign _1081_ = _1073_ & _1080_ /*10611*/;
assign _981_ = _1073_ ^ _1080_ /*10612*/;
assign _1078_ = _1079_ | _1081_ /*10609*/;
assign _1087_ = D[17] ^ Q[27] /*10608*/;
assign _1084_ = _788_ & _1087_ /*10604*/;
assign _1085_ = _788_ ^ _1087_ /*10607*/;
assign _1086_ = _1078_ & _1085_ /*10605*/;
assign _982_ = _1078_ ^ _1085_ /*10606*/;
assign _1083_ = _1084_ | _1086_ /*10603*/;
assign _1092_ = D[18] ^ Q[27] /*10602*/;
assign _1089_ = _789_ & _1092_ /*10598*/;
assign _1090_ = _789_ ^ _1092_ /*10601*/;
assign _1091_ = _1083_ & _1090_ /*10599*/;
assign _983_ = _1083_ ^ _1090_ /*10600*/;
assign _1088_ = _1089_ | _1091_ /*10597*/;
assign _1097_ = D[19] ^ Q[27] /*10596*/;
assign _1094_ = _790_ & _1097_ /*10592*/;
assign _1095_ = _790_ ^ _1097_ /*10595*/;
assign _1096_ = _1088_ & _1095_ /*10593*/;
assign _984_ = _1088_ ^ _1095_ /*10594*/;
assign _1093_ = _1094_ | _1096_ /*10591*/;
assign _1102_ = D[20] ^ Q[27] /*10590*/;
assign _1099_ = _791_ & _1102_ /*10586*/;
assign _1100_ = _791_ ^ _1102_ /*10589*/;
assign _1101_ = _1093_ & _1100_ /*10587*/;
assign _985_ = _1093_ ^ _1100_ /*10588*/;
assign _1098_ = _1099_ | _1101_ /*10585*/;
assign _1107_ = D[21] ^ Q[27] /*10584*/;
assign _1104_ = _792_ & _1107_ /*10580*/;
assign _1105_ = _792_ ^ _1107_ /*10583*/;
assign _1106_ = _1098_ & _1105_ /*10581*/;
assign _986_ = _1098_ ^ _1105_ /*10582*/;
assign _1103_ = _1104_ | _1106_ /*10579*/;
assign _1112_ = D[22] ^ Q[27] /*10578*/;
assign _1109_ = _793_ & _1112_ /*10574*/;
assign _1110_ = _793_ ^ _1112_ /*10577*/;
assign _1111_ = _1103_ & _1110_ /*10575*/;
assign _987_ = _1103_ ^ _1110_ /*10576*/;
assign _1108_ = _1109_ | _1111_ /*10573*/;
assign _1117_ = D[23] ^ Q[27] /*10572*/;
assign _1114_ = _794_ & _1117_ /*10568*/;
assign _1115_ = _794_ ^ _1117_ /*10571*/;
assign _1116_ = _1108_ & _1115_ /*10569*/;
assign _988_ = _1108_ ^ _1115_ /*10570*/;
assign _1113_ = _1114_ | _1116_ /*10567*/;
assign _1122_ = D[24] ^ Q[27] /*10566*/;
assign _1119_ = _795_ & _1122_ /*10562*/;
assign _1120_ = _795_ ^ _1122_ /*10565*/;
assign _1121_ = _1113_ & _1120_ /*10563*/;
assign _989_ = _1113_ ^ _1120_ /*10564*/;
assign _1118_ = _1119_ | _1121_ /*10561*/;
assign _1127_ = D[25] ^ Q[27] /*10560*/;
assign _1124_ = _796_ & _1127_ /*10556*/;
assign _1125_ = _796_ ^ _1127_ /*10559*/;
assign _1126_ = _1118_ & _1125_ /*10557*/;
assign _990_ = _1118_ ^ _1125_ /*10558*/;
assign _1123_ = _1124_ | _1126_ /*10555*/;
assign _1132_ = D[26] ^ Q[27] /*10554*/;
assign _1129_ = _797_ & _1132_ /*10550*/;
assign _1130_ = _797_ ^ _1132_ /*10553*/;
assign _1131_ = _1123_ & _1130_ /*10551*/;
assign _991_ = _1123_ ^ _1130_ /*10552*/;
assign _1128_ = _1129_ | _1131_ /*10549*/;
assign _1137_ = D[27] ^ Q[27] /*10548*/;
assign _1134_ = _798_ & _1137_ /*10544*/;
assign _1135_ = _798_ ^ _1137_ /*10547*/;
assign _1136_ = _1128_ & _1135_ /*10545*/;
assign _992_ = _1128_ ^ _1135_ /*10546*/;
assign _1133_ = _1134_ | _1136_ /*10543*/;
assign _1142_ = D[28] ^ Q[27] /*10542*/;
assign _1139_ = _799_ & _1142_ /*10538*/;
assign _1140_ = _799_ ^ _1142_ /*10541*/;
assign _1141_ = _1133_ & _1140_ /*10539*/;
assign _993_ = _1133_ ^ _1140_ /*10540*/;
assign _1138_ = _1139_ | _1141_ /*10537*/;
assign _1147_ = D[29] ^ Q[27] /*10536*/;
assign _1144_ = _800_ & _1147_ /*10532*/;
assign _1145_ = _800_ ^ _1147_ /*10535*/;
assign _1146_ = _1138_ & _1145_ /*10533*/;
assign _994_ = _1138_ ^ _1145_ /*10534*/;
assign _1143_ = _1144_ | _1146_ /*10531*/;
assign _1152_ = D[30] ^ Q[27] /*10530*/;
assign _1149_ = _801_ & _1152_ /*10526*/;
assign _1150_ = _801_ ^ _1152_ /*10529*/;
assign _1151_ = _1143_ & _1150_ /*10527*/;
assign _995_ = _1143_ ^ _1150_ /*10528*/;
assign _1148_ = _1149_ | _1151_ /*10525*/;
assign _1156_ = zeroWire ^ Q[27] /*10524*/;
assign _1153_ = _802_ & _1156_ /*10520*/;
assign _1154_ = _802_ ^ _1156_ /*10523*/;
assign _1155_ = _1148_ & _1154_ /*10521*/;
assign _996_ = _1148_ ^ _1154_ /*10522*/;
assign Q[26] = _1153_ | _1155_ /*10519*/;
assign _1195_ = D[0] ^ Q[26] /*10325*/;
assign _1192_ = R_0[25] & _1195_ /*10321*/;
assign _1193_ = R_0[25] ^ _1195_ /*10324*/;
assign _1194_ = Q[26] & _1193_ /*10322*/;
assign _1158_ = Q[26] ^ _1193_ /*10323*/;
assign _1191_ = _1192_ | _1194_ /*10320*/;
assign _1200_ = D[1] ^ Q[26] /*10319*/;
assign _1197_ = _965_ & _1200_ /*10315*/;
assign _1198_ = _965_ ^ _1200_ /*10318*/;
assign _1199_ = _1191_ & _1198_ /*10316*/;
assign _1159_ = _1191_ ^ _1198_ /*10317*/;
assign _1196_ = _1197_ | _1199_ /*10314*/;
assign _1205_ = D[2] ^ Q[26] /*10313*/;
assign _1202_ = _966_ & _1205_ /*10309*/;
assign _1203_ = _966_ ^ _1205_ /*10312*/;
assign _1204_ = _1196_ & _1203_ /*10310*/;
assign _1160_ = _1196_ ^ _1203_ /*10311*/;
assign _1201_ = _1202_ | _1204_ /*10308*/;
assign _1210_ = D[3] ^ Q[26] /*10307*/;
assign _1207_ = _967_ & _1210_ /*10303*/;
assign _1208_ = _967_ ^ _1210_ /*10306*/;
assign _1209_ = _1201_ & _1208_ /*10304*/;
assign _1161_ = _1201_ ^ _1208_ /*10305*/;
assign _1206_ = _1207_ | _1209_ /*10302*/;
assign _1215_ = D[4] ^ Q[26] /*10301*/;
assign _1212_ = _968_ & _1215_ /*10297*/;
assign _1213_ = _968_ ^ _1215_ /*10300*/;
assign _1214_ = _1206_ & _1213_ /*10298*/;
assign _1162_ = _1206_ ^ _1213_ /*10299*/;
assign _1211_ = _1212_ | _1214_ /*10296*/;
assign _1220_ = D[5] ^ Q[26] /*10295*/;
assign _1217_ = _969_ & _1220_ /*10291*/;
assign _1218_ = _969_ ^ _1220_ /*10294*/;
assign _1219_ = _1211_ & _1218_ /*10292*/;
assign _1163_ = _1211_ ^ _1218_ /*10293*/;
assign _1216_ = _1217_ | _1219_ /*10290*/;
assign _1225_ = D[6] ^ Q[26] /*10289*/;
assign _1222_ = _970_ & _1225_ /*10285*/;
assign _1223_ = _970_ ^ _1225_ /*10288*/;
assign _1224_ = _1216_ & _1223_ /*10286*/;
assign _1164_ = _1216_ ^ _1223_ /*10287*/;
assign _1221_ = _1222_ | _1224_ /*10284*/;
assign _1230_ = D[7] ^ Q[26] /*10283*/;
assign _1227_ = _971_ & _1230_ /*10279*/;
assign _1228_ = _971_ ^ _1230_ /*10282*/;
assign _1229_ = _1221_ & _1228_ /*10280*/;
assign _1165_ = _1221_ ^ _1228_ /*10281*/;
assign _1226_ = _1227_ | _1229_ /*10278*/;
assign _1235_ = D[8] ^ Q[26] /*10277*/;
assign _1232_ = _972_ & _1235_ /*10273*/;
assign _1233_ = _972_ ^ _1235_ /*10276*/;
assign _1234_ = _1226_ & _1233_ /*10274*/;
assign _1166_ = _1226_ ^ _1233_ /*10275*/;
assign _1231_ = _1232_ | _1234_ /*10272*/;
assign _1240_ = D[9] ^ Q[26] /*10271*/;
assign _1237_ = _973_ & _1240_ /*10267*/;
assign _1238_ = _973_ ^ _1240_ /*10270*/;
assign _1239_ = _1231_ & _1238_ /*10268*/;
assign _1167_ = _1231_ ^ _1238_ /*10269*/;
assign _1236_ = _1237_ | _1239_ /*10266*/;
assign _1245_ = D[10] ^ Q[26] /*10265*/;
assign _1242_ = _974_ & _1245_ /*10261*/;
assign _1243_ = _974_ ^ _1245_ /*10264*/;
assign _1244_ = _1236_ & _1243_ /*10262*/;
assign _1168_ = _1236_ ^ _1243_ /*10263*/;
assign _1241_ = _1242_ | _1244_ /*10260*/;
assign _1250_ = D[11] ^ Q[26] /*10259*/;
assign _1247_ = _975_ & _1250_ /*10255*/;
assign _1248_ = _975_ ^ _1250_ /*10258*/;
assign _1249_ = _1241_ & _1248_ /*10256*/;
assign _1169_ = _1241_ ^ _1248_ /*10257*/;
assign _1246_ = _1247_ | _1249_ /*10254*/;
assign _1255_ = D[12] ^ Q[26] /*10253*/;
assign _1252_ = _976_ & _1255_ /*10249*/;
assign _1253_ = _976_ ^ _1255_ /*10252*/;
assign _1254_ = _1246_ & _1253_ /*10250*/;
assign _1170_ = _1246_ ^ _1253_ /*10251*/;
assign _1251_ = _1252_ | _1254_ /*10248*/;
assign _1260_ = D[13] ^ Q[26] /*10247*/;
assign _1257_ = _977_ & _1260_ /*10243*/;
assign _1258_ = _977_ ^ _1260_ /*10246*/;
assign _1259_ = _1251_ & _1258_ /*10244*/;
assign _1171_ = _1251_ ^ _1258_ /*10245*/;
assign _1256_ = _1257_ | _1259_ /*10242*/;
assign _1265_ = D[14] ^ Q[26] /*10241*/;
assign _1262_ = _978_ & _1265_ /*10237*/;
assign _1263_ = _978_ ^ _1265_ /*10240*/;
assign _1264_ = _1256_ & _1263_ /*10238*/;
assign _1172_ = _1256_ ^ _1263_ /*10239*/;
assign _1261_ = _1262_ | _1264_ /*10236*/;
assign _1270_ = D[15] ^ Q[26] /*10235*/;
assign _1267_ = _979_ & _1270_ /*10231*/;
assign _1268_ = _979_ ^ _1270_ /*10234*/;
assign _1269_ = _1261_ & _1268_ /*10232*/;
assign _1173_ = _1261_ ^ _1268_ /*10233*/;
assign _1266_ = _1267_ | _1269_ /*10230*/;
assign _1275_ = D[16] ^ Q[26] /*10229*/;
assign _1272_ = _980_ & _1275_ /*10225*/;
assign _1273_ = _980_ ^ _1275_ /*10228*/;
assign _1274_ = _1266_ & _1273_ /*10226*/;
assign _1174_ = _1266_ ^ _1273_ /*10227*/;
assign _1271_ = _1272_ | _1274_ /*10224*/;
assign _1280_ = D[17] ^ Q[26] /*10223*/;
assign _1277_ = _981_ & _1280_ /*10219*/;
assign _1278_ = _981_ ^ _1280_ /*10222*/;
assign _1279_ = _1271_ & _1278_ /*10220*/;
assign _1175_ = _1271_ ^ _1278_ /*10221*/;
assign _1276_ = _1277_ | _1279_ /*10218*/;
assign _1285_ = D[18] ^ Q[26] /*10217*/;
assign _1282_ = _982_ & _1285_ /*10213*/;
assign _1283_ = _982_ ^ _1285_ /*10216*/;
assign _1284_ = _1276_ & _1283_ /*10214*/;
assign _1176_ = _1276_ ^ _1283_ /*10215*/;
assign _1281_ = _1282_ | _1284_ /*10212*/;
assign _1290_ = D[19] ^ Q[26] /*10211*/;
assign _1287_ = _983_ & _1290_ /*10207*/;
assign _1288_ = _983_ ^ _1290_ /*10210*/;
assign _1289_ = _1281_ & _1288_ /*10208*/;
assign _1177_ = _1281_ ^ _1288_ /*10209*/;
assign _1286_ = _1287_ | _1289_ /*10206*/;
assign _1295_ = D[20] ^ Q[26] /*10205*/;
assign _1292_ = _984_ & _1295_ /*10201*/;
assign _1293_ = _984_ ^ _1295_ /*10204*/;
assign _1294_ = _1286_ & _1293_ /*10202*/;
assign _1178_ = _1286_ ^ _1293_ /*10203*/;
assign _1291_ = _1292_ | _1294_ /*10200*/;
assign _1300_ = D[21] ^ Q[26] /*10199*/;
assign _1297_ = _985_ & _1300_ /*10195*/;
assign _1298_ = _985_ ^ _1300_ /*10198*/;
assign _1299_ = _1291_ & _1298_ /*10196*/;
assign _1179_ = _1291_ ^ _1298_ /*10197*/;
assign _1296_ = _1297_ | _1299_ /*10194*/;
assign _1305_ = D[22] ^ Q[26] /*10193*/;
assign _1302_ = _986_ & _1305_ /*10189*/;
assign _1303_ = _986_ ^ _1305_ /*10192*/;
assign _1304_ = _1296_ & _1303_ /*10190*/;
assign _1180_ = _1296_ ^ _1303_ /*10191*/;
assign _1301_ = _1302_ | _1304_ /*10188*/;
assign _1310_ = D[23] ^ Q[26] /*10187*/;
assign _1307_ = _987_ & _1310_ /*10183*/;
assign _1308_ = _987_ ^ _1310_ /*10186*/;
assign _1309_ = _1301_ & _1308_ /*10184*/;
assign _1181_ = _1301_ ^ _1308_ /*10185*/;
assign _1306_ = _1307_ | _1309_ /*10182*/;
assign _1315_ = D[24] ^ Q[26] /*10181*/;
assign _1312_ = _988_ & _1315_ /*10177*/;
assign _1313_ = _988_ ^ _1315_ /*10180*/;
assign _1314_ = _1306_ & _1313_ /*10178*/;
assign _1182_ = _1306_ ^ _1313_ /*10179*/;
assign _1311_ = _1312_ | _1314_ /*10176*/;
assign _1320_ = D[25] ^ Q[26] /*10175*/;
assign _1317_ = _989_ & _1320_ /*10171*/;
assign _1318_ = _989_ ^ _1320_ /*10174*/;
assign _1319_ = _1311_ & _1318_ /*10172*/;
assign _1183_ = _1311_ ^ _1318_ /*10173*/;
assign _1316_ = _1317_ | _1319_ /*10170*/;
assign _1325_ = D[26] ^ Q[26] /*10169*/;
assign _1322_ = _990_ & _1325_ /*10165*/;
assign _1323_ = _990_ ^ _1325_ /*10168*/;
assign _1324_ = _1316_ & _1323_ /*10166*/;
assign _1184_ = _1316_ ^ _1323_ /*10167*/;
assign _1321_ = _1322_ | _1324_ /*10164*/;
assign _1330_ = D[27] ^ Q[26] /*10163*/;
assign _1327_ = _991_ & _1330_ /*10159*/;
assign _1328_ = _991_ ^ _1330_ /*10162*/;
assign _1329_ = _1321_ & _1328_ /*10160*/;
assign _1185_ = _1321_ ^ _1328_ /*10161*/;
assign _1326_ = _1327_ | _1329_ /*10158*/;
assign _1335_ = D[28] ^ Q[26] /*10157*/;
assign _1332_ = _992_ & _1335_ /*10153*/;
assign _1333_ = _992_ ^ _1335_ /*10156*/;
assign _1334_ = _1326_ & _1333_ /*10154*/;
assign _1186_ = _1326_ ^ _1333_ /*10155*/;
assign _1331_ = _1332_ | _1334_ /*10152*/;
assign _1340_ = D[29] ^ Q[26] /*10151*/;
assign _1337_ = _993_ & _1340_ /*10147*/;
assign _1338_ = _993_ ^ _1340_ /*10150*/;
assign _1339_ = _1331_ & _1338_ /*10148*/;
assign _1187_ = _1331_ ^ _1338_ /*10149*/;
assign _1336_ = _1337_ | _1339_ /*10146*/;
assign _1345_ = D[30] ^ Q[26] /*10145*/;
assign _1342_ = _994_ & _1345_ /*10141*/;
assign _1343_ = _994_ ^ _1345_ /*10144*/;
assign _1344_ = _1336_ & _1343_ /*10142*/;
assign _1188_ = _1336_ ^ _1343_ /*10143*/;
assign _1341_ = _1342_ | _1344_ /*10140*/;
assign _1349_ = zeroWire ^ Q[26] /*10139*/;
assign _1346_ = _995_ & _1349_ /*10135*/;
assign _1347_ = _995_ ^ _1349_ /*10138*/;
assign _1348_ = _1341_ & _1347_ /*10136*/;
assign _1189_ = _1341_ ^ _1347_ /*10137*/;
assign Q[25] = _1346_ | _1348_ /*10134*/;
assign _1388_ = D[0] ^ Q[25] /*9940*/;
assign _1385_ = R_0[24] & _1388_ /*9936*/;
assign _1386_ = R_0[24] ^ _1388_ /*9939*/;
assign _1387_ = Q[25] & _1386_ /*9937*/;
assign _1351_ = Q[25] ^ _1386_ /*9938*/;
assign _1384_ = _1385_ | _1387_ /*9935*/;
assign _1393_ = D[1] ^ Q[25] /*9934*/;
assign _1390_ = _1158_ & _1393_ /*9930*/;
assign _1391_ = _1158_ ^ _1393_ /*9933*/;
assign _1392_ = _1384_ & _1391_ /*9931*/;
assign _1352_ = _1384_ ^ _1391_ /*9932*/;
assign _1389_ = _1390_ | _1392_ /*9929*/;
assign _1398_ = D[2] ^ Q[25] /*9928*/;
assign _1395_ = _1159_ & _1398_ /*9924*/;
assign _1396_ = _1159_ ^ _1398_ /*9927*/;
assign _1397_ = _1389_ & _1396_ /*9925*/;
assign _1353_ = _1389_ ^ _1396_ /*9926*/;
assign _1394_ = _1395_ | _1397_ /*9923*/;
assign _1403_ = D[3] ^ Q[25] /*9922*/;
assign _1400_ = _1160_ & _1403_ /*9918*/;
assign _1401_ = _1160_ ^ _1403_ /*9921*/;
assign _1402_ = _1394_ & _1401_ /*9919*/;
assign _1354_ = _1394_ ^ _1401_ /*9920*/;
assign _1399_ = _1400_ | _1402_ /*9917*/;
assign _1408_ = D[4] ^ Q[25] /*9916*/;
assign _1405_ = _1161_ & _1408_ /*9912*/;
assign _1406_ = _1161_ ^ _1408_ /*9915*/;
assign _1407_ = _1399_ & _1406_ /*9913*/;
assign _1355_ = _1399_ ^ _1406_ /*9914*/;
assign _1404_ = _1405_ | _1407_ /*9911*/;
assign _1413_ = D[5] ^ Q[25] /*9910*/;
assign _1410_ = _1162_ & _1413_ /*9906*/;
assign _1411_ = _1162_ ^ _1413_ /*9909*/;
assign _1412_ = _1404_ & _1411_ /*9907*/;
assign _1356_ = _1404_ ^ _1411_ /*9908*/;
assign _1409_ = _1410_ | _1412_ /*9905*/;
assign _1418_ = D[6] ^ Q[25] /*9904*/;
assign _1415_ = _1163_ & _1418_ /*9900*/;
assign _1416_ = _1163_ ^ _1418_ /*9903*/;
assign _1417_ = _1409_ & _1416_ /*9901*/;
assign _1357_ = _1409_ ^ _1416_ /*9902*/;
assign _1414_ = _1415_ | _1417_ /*9899*/;
assign _1423_ = D[7] ^ Q[25] /*9898*/;
assign _1420_ = _1164_ & _1423_ /*9894*/;
assign _1421_ = _1164_ ^ _1423_ /*9897*/;
assign _1422_ = _1414_ & _1421_ /*9895*/;
assign _1358_ = _1414_ ^ _1421_ /*9896*/;
assign _1419_ = _1420_ | _1422_ /*9893*/;
assign _1428_ = D[8] ^ Q[25] /*9892*/;
assign _1425_ = _1165_ & _1428_ /*9888*/;
assign _1426_ = _1165_ ^ _1428_ /*9891*/;
assign _1427_ = _1419_ & _1426_ /*9889*/;
assign _1359_ = _1419_ ^ _1426_ /*9890*/;
assign _1424_ = _1425_ | _1427_ /*9887*/;
assign _1433_ = D[9] ^ Q[25] /*9886*/;
assign _1430_ = _1166_ & _1433_ /*9882*/;
assign _1431_ = _1166_ ^ _1433_ /*9885*/;
assign _1432_ = _1424_ & _1431_ /*9883*/;
assign _1360_ = _1424_ ^ _1431_ /*9884*/;
assign _1429_ = _1430_ | _1432_ /*9881*/;
assign _1438_ = D[10] ^ Q[25] /*9880*/;
assign _1435_ = _1167_ & _1438_ /*9876*/;
assign _1436_ = _1167_ ^ _1438_ /*9879*/;
assign _1437_ = _1429_ & _1436_ /*9877*/;
assign _1361_ = _1429_ ^ _1436_ /*9878*/;
assign _1434_ = _1435_ | _1437_ /*9875*/;
assign _1443_ = D[11] ^ Q[25] /*9874*/;
assign _1440_ = _1168_ & _1443_ /*9870*/;
assign _1441_ = _1168_ ^ _1443_ /*9873*/;
assign _1442_ = _1434_ & _1441_ /*9871*/;
assign _1362_ = _1434_ ^ _1441_ /*9872*/;
assign _1439_ = _1440_ | _1442_ /*9869*/;
assign _1448_ = D[12] ^ Q[25] /*9868*/;
assign _1445_ = _1169_ & _1448_ /*9864*/;
assign _1446_ = _1169_ ^ _1448_ /*9867*/;
assign _1447_ = _1439_ & _1446_ /*9865*/;
assign _1363_ = _1439_ ^ _1446_ /*9866*/;
assign _1444_ = _1445_ | _1447_ /*9863*/;
assign _1453_ = D[13] ^ Q[25] /*9862*/;
assign _1450_ = _1170_ & _1453_ /*9858*/;
assign _1451_ = _1170_ ^ _1453_ /*9861*/;
assign _1452_ = _1444_ & _1451_ /*9859*/;
assign _1364_ = _1444_ ^ _1451_ /*9860*/;
assign _1449_ = _1450_ | _1452_ /*9857*/;
assign _1458_ = D[14] ^ Q[25] /*9856*/;
assign _1455_ = _1171_ & _1458_ /*9852*/;
assign _1456_ = _1171_ ^ _1458_ /*9855*/;
assign _1457_ = _1449_ & _1456_ /*9853*/;
assign _1365_ = _1449_ ^ _1456_ /*9854*/;
assign _1454_ = _1455_ | _1457_ /*9851*/;
assign _1463_ = D[15] ^ Q[25] /*9850*/;
assign _1460_ = _1172_ & _1463_ /*9846*/;
assign _1461_ = _1172_ ^ _1463_ /*9849*/;
assign _1462_ = _1454_ & _1461_ /*9847*/;
assign _1366_ = _1454_ ^ _1461_ /*9848*/;
assign _1459_ = _1460_ | _1462_ /*9845*/;
assign _1468_ = D[16] ^ Q[25] /*9844*/;
assign _1465_ = _1173_ & _1468_ /*9840*/;
assign _1466_ = _1173_ ^ _1468_ /*9843*/;
assign _1467_ = _1459_ & _1466_ /*9841*/;
assign _1367_ = _1459_ ^ _1466_ /*9842*/;
assign _1464_ = _1465_ | _1467_ /*9839*/;
assign _1473_ = D[17] ^ Q[25] /*9838*/;
assign _1470_ = _1174_ & _1473_ /*9834*/;
assign _1471_ = _1174_ ^ _1473_ /*9837*/;
assign _1472_ = _1464_ & _1471_ /*9835*/;
assign _1368_ = _1464_ ^ _1471_ /*9836*/;
assign _1469_ = _1470_ | _1472_ /*9833*/;
assign _1478_ = D[18] ^ Q[25] /*9832*/;
assign _1475_ = _1175_ & _1478_ /*9828*/;
assign _1476_ = _1175_ ^ _1478_ /*9831*/;
assign _1477_ = _1469_ & _1476_ /*9829*/;
assign _1369_ = _1469_ ^ _1476_ /*9830*/;
assign _1474_ = _1475_ | _1477_ /*9827*/;
assign _1483_ = D[19] ^ Q[25] /*9826*/;
assign _1480_ = _1176_ & _1483_ /*9822*/;
assign _1481_ = _1176_ ^ _1483_ /*9825*/;
assign _1482_ = _1474_ & _1481_ /*9823*/;
assign _1370_ = _1474_ ^ _1481_ /*9824*/;
assign _1479_ = _1480_ | _1482_ /*9821*/;
assign _1488_ = D[20] ^ Q[25] /*9820*/;
assign _1485_ = _1177_ & _1488_ /*9816*/;
assign _1486_ = _1177_ ^ _1488_ /*9819*/;
assign _1487_ = _1479_ & _1486_ /*9817*/;
assign _1371_ = _1479_ ^ _1486_ /*9818*/;
assign _1484_ = _1485_ | _1487_ /*9815*/;
assign _1493_ = D[21] ^ Q[25] /*9814*/;
assign _1490_ = _1178_ & _1493_ /*9810*/;
assign _1491_ = _1178_ ^ _1493_ /*9813*/;
assign _1492_ = _1484_ & _1491_ /*9811*/;
assign _1372_ = _1484_ ^ _1491_ /*9812*/;
assign _1489_ = _1490_ | _1492_ /*9809*/;
assign _1498_ = D[22] ^ Q[25] /*9808*/;
assign _1495_ = _1179_ & _1498_ /*9804*/;
assign _1496_ = _1179_ ^ _1498_ /*9807*/;
assign _1497_ = _1489_ & _1496_ /*9805*/;
assign _1373_ = _1489_ ^ _1496_ /*9806*/;
assign _1494_ = _1495_ | _1497_ /*9803*/;
assign _1503_ = D[23] ^ Q[25] /*9802*/;
assign _1500_ = _1180_ & _1503_ /*9798*/;
assign _1501_ = _1180_ ^ _1503_ /*9801*/;
assign _1502_ = _1494_ & _1501_ /*9799*/;
assign _1374_ = _1494_ ^ _1501_ /*9800*/;
assign _1499_ = _1500_ | _1502_ /*9797*/;
assign _1508_ = D[24] ^ Q[25] /*9796*/;
assign _1505_ = _1181_ & _1508_ /*9792*/;
assign _1506_ = _1181_ ^ _1508_ /*9795*/;
assign _1507_ = _1499_ & _1506_ /*9793*/;
assign _1375_ = _1499_ ^ _1506_ /*9794*/;
assign _1504_ = _1505_ | _1507_ /*9791*/;
assign _1513_ = D[25] ^ Q[25] /*9790*/;
assign _1510_ = _1182_ & _1513_ /*9786*/;
assign _1511_ = _1182_ ^ _1513_ /*9789*/;
assign _1512_ = _1504_ & _1511_ /*9787*/;
assign _1376_ = _1504_ ^ _1511_ /*9788*/;
assign _1509_ = _1510_ | _1512_ /*9785*/;
assign _1518_ = D[26] ^ Q[25] /*9784*/;
assign _1515_ = _1183_ & _1518_ /*9780*/;
assign _1516_ = _1183_ ^ _1518_ /*9783*/;
assign _1517_ = _1509_ & _1516_ /*9781*/;
assign _1377_ = _1509_ ^ _1516_ /*9782*/;
assign _1514_ = _1515_ | _1517_ /*9779*/;
assign _1523_ = D[27] ^ Q[25] /*9778*/;
assign _1520_ = _1184_ & _1523_ /*9774*/;
assign _1521_ = _1184_ ^ _1523_ /*9777*/;
assign _1522_ = _1514_ & _1521_ /*9775*/;
assign _1378_ = _1514_ ^ _1521_ /*9776*/;
assign _1519_ = _1520_ | _1522_ /*9773*/;
assign _1528_ = D[28] ^ Q[25] /*9772*/;
assign _1525_ = _1185_ & _1528_ /*9768*/;
assign _1526_ = _1185_ ^ _1528_ /*9771*/;
assign _1527_ = _1519_ & _1526_ /*9769*/;
assign _1379_ = _1519_ ^ _1526_ /*9770*/;
assign _1524_ = _1525_ | _1527_ /*9767*/;
assign _1533_ = D[29] ^ Q[25] /*9766*/;
assign _1530_ = _1186_ & _1533_ /*9762*/;
assign _1531_ = _1186_ ^ _1533_ /*9765*/;
assign _1532_ = _1524_ & _1531_ /*9763*/;
assign _1380_ = _1524_ ^ _1531_ /*9764*/;
assign _1529_ = _1530_ | _1532_ /*9761*/;
assign _1538_ = D[30] ^ Q[25] /*9760*/;
assign _1535_ = _1187_ & _1538_ /*9756*/;
assign _1536_ = _1187_ ^ _1538_ /*9759*/;
assign _1537_ = _1529_ & _1536_ /*9757*/;
assign _1381_ = _1529_ ^ _1536_ /*9758*/;
assign _1534_ = _1535_ | _1537_ /*9755*/;
assign _1542_ = zeroWire ^ Q[25] /*9754*/;
assign _1539_ = _1188_ & _1542_ /*9750*/;
assign _1540_ = _1188_ ^ _1542_ /*9753*/;
assign _1541_ = _1534_ & _1540_ /*9751*/;
assign _1382_ = _1534_ ^ _1540_ /*9752*/;
assign Q[24] = _1539_ | _1541_ /*9749*/;
assign _1581_ = D[0] ^ Q[24] /*9555*/;
assign _1578_ = R_0[23] & _1581_ /*9551*/;
assign _1579_ = R_0[23] ^ _1581_ /*9554*/;
assign _1580_ = Q[24] & _1579_ /*9552*/;
assign _1544_ = Q[24] ^ _1579_ /*9553*/;
assign _1577_ = _1578_ | _1580_ /*9550*/;
assign _1586_ = D[1] ^ Q[24] /*9549*/;
assign _1583_ = _1351_ & _1586_ /*9545*/;
assign _1584_ = _1351_ ^ _1586_ /*9548*/;
assign _1585_ = _1577_ & _1584_ /*9546*/;
assign _1545_ = _1577_ ^ _1584_ /*9547*/;
assign _1582_ = _1583_ | _1585_ /*9544*/;
assign _1591_ = D[2] ^ Q[24] /*9543*/;
assign _1588_ = _1352_ & _1591_ /*9539*/;
assign _1589_ = _1352_ ^ _1591_ /*9542*/;
assign _1590_ = _1582_ & _1589_ /*9540*/;
assign _1546_ = _1582_ ^ _1589_ /*9541*/;
assign _1587_ = _1588_ | _1590_ /*9538*/;
assign _1596_ = D[3] ^ Q[24] /*9537*/;
assign _1593_ = _1353_ & _1596_ /*9533*/;
assign _1594_ = _1353_ ^ _1596_ /*9536*/;
assign _1595_ = _1587_ & _1594_ /*9534*/;
assign _1547_ = _1587_ ^ _1594_ /*9535*/;
assign _1592_ = _1593_ | _1595_ /*9532*/;
assign _1601_ = D[4] ^ Q[24] /*9531*/;
assign _1598_ = _1354_ & _1601_ /*9527*/;
assign _1599_ = _1354_ ^ _1601_ /*9530*/;
assign _1600_ = _1592_ & _1599_ /*9528*/;
assign _1548_ = _1592_ ^ _1599_ /*9529*/;
assign _1597_ = _1598_ | _1600_ /*9526*/;
assign _1606_ = D[5] ^ Q[24] /*9525*/;
assign _1603_ = _1355_ & _1606_ /*9521*/;
assign _1604_ = _1355_ ^ _1606_ /*9524*/;
assign _1605_ = _1597_ & _1604_ /*9522*/;
assign _1549_ = _1597_ ^ _1604_ /*9523*/;
assign _1602_ = _1603_ | _1605_ /*9520*/;
assign _1611_ = D[6] ^ Q[24] /*9519*/;
assign _1608_ = _1356_ & _1611_ /*9515*/;
assign _1609_ = _1356_ ^ _1611_ /*9518*/;
assign _1610_ = _1602_ & _1609_ /*9516*/;
assign _1550_ = _1602_ ^ _1609_ /*9517*/;
assign _1607_ = _1608_ | _1610_ /*9514*/;
assign _1616_ = D[7] ^ Q[24] /*9513*/;
assign _1613_ = _1357_ & _1616_ /*9509*/;
assign _1614_ = _1357_ ^ _1616_ /*9512*/;
assign _1615_ = _1607_ & _1614_ /*9510*/;
assign _1551_ = _1607_ ^ _1614_ /*9511*/;
assign _1612_ = _1613_ | _1615_ /*9508*/;
assign _1621_ = D[8] ^ Q[24] /*9507*/;
assign _1618_ = _1358_ & _1621_ /*9503*/;
assign _1619_ = _1358_ ^ _1621_ /*9506*/;
assign _1620_ = _1612_ & _1619_ /*9504*/;
assign _1552_ = _1612_ ^ _1619_ /*9505*/;
assign _1617_ = _1618_ | _1620_ /*9502*/;
assign _1626_ = D[9] ^ Q[24] /*9501*/;
assign _1623_ = _1359_ & _1626_ /*9497*/;
assign _1624_ = _1359_ ^ _1626_ /*9500*/;
assign _1625_ = _1617_ & _1624_ /*9498*/;
assign _1553_ = _1617_ ^ _1624_ /*9499*/;
assign _1622_ = _1623_ | _1625_ /*9496*/;
assign _1631_ = D[10] ^ Q[24] /*9495*/;
assign _1628_ = _1360_ & _1631_ /*9491*/;
assign _1629_ = _1360_ ^ _1631_ /*9494*/;
assign _1630_ = _1622_ & _1629_ /*9492*/;
assign _1554_ = _1622_ ^ _1629_ /*9493*/;
assign _1627_ = _1628_ | _1630_ /*9490*/;
assign _1636_ = D[11] ^ Q[24] /*9489*/;
assign _1633_ = _1361_ & _1636_ /*9485*/;
assign _1634_ = _1361_ ^ _1636_ /*9488*/;
assign _1635_ = _1627_ & _1634_ /*9486*/;
assign _1555_ = _1627_ ^ _1634_ /*9487*/;
assign _1632_ = _1633_ | _1635_ /*9484*/;
assign _1641_ = D[12] ^ Q[24] /*9483*/;
assign _1638_ = _1362_ & _1641_ /*9479*/;
assign _1639_ = _1362_ ^ _1641_ /*9482*/;
assign _1640_ = _1632_ & _1639_ /*9480*/;
assign _1556_ = _1632_ ^ _1639_ /*9481*/;
assign _1637_ = _1638_ | _1640_ /*9478*/;
assign _1646_ = D[13] ^ Q[24] /*9477*/;
assign _1643_ = _1363_ & _1646_ /*9473*/;
assign _1644_ = _1363_ ^ _1646_ /*9476*/;
assign _1645_ = _1637_ & _1644_ /*9474*/;
assign _1557_ = _1637_ ^ _1644_ /*9475*/;
assign _1642_ = _1643_ | _1645_ /*9472*/;
assign _1651_ = D[14] ^ Q[24] /*9471*/;
assign _1648_ = _1364_ & _1651_ /*9467*/;
assign _1649_ = _1364_ ^ _1651_ /*9470*/;
assign _1650_ = _1642_ & _1649_ /*9468*/;
assign _1558_ = _1642_ ^ _1649_ /*9469*/;
assign _1647_ = _1648_ | _1650_ /*9466*/;
assign _1656_ = D[15] ^ Q[24] /*9465*/;
assign _1653_ = _1365_ & _1656_ /*9461*/;
assign _1654_ = _1365_ ^ _1656_ /*9464*/;
assign _1655_ = _1647_ & _1654_ /*9462*/;
assign _1559_ = _1647_ ^ _1654_ /*9463*/;
assign _1652_ = _1653_ | _1655_ /*9460*/;
assign _1661_ = D[16] ^ Q[24] /*9459*/;
assign _1658_ = _1366_ & _1661_ /*9455*/;
assign _1659_ = _1366_ ^ _1661_ /*9458*/;
assign _1660_ = _1652_ & _1659_ /*9456*/;
assign _1560_ = _1652_ ^ _1659_ /*9457*/;
assign _1657_ = _1658_ | _1660_ /*9454*/;
assign _1666_ = D[17] ^ Q[24] /*9453*/;
assign _1663_ = _1367_ & _1666_ /*9449*/;
assign _1664_ = _1367_ ^ _1666_ /*9452*/;
assign _1665_ = _1657_ & _1664_ /*9450*/;
assign _1561_ = _1657_ ^ _1664_ /*9451*/;
assign _1662_ = _1663_ | _1665_ /*9448*/;
assign _1671_ = D[18] ^ Q[24] /*9447*/;
assign _1668_ = _1368_ & _1671_ /*9443*/;
assign _1669_ = _1368_ ^ _1671_ /*9446*/;
assign _1670_ = _1662_ & _1669_ /*9444*/;
assign _1562_ = _1662_ ^ _1669_ /*9445*/;
assign _1667_ = _1668_ | _1670_ /*9442*/;
assign _1676_ = D[19] ^ Q[24] /*9441*/;
assign _1673_ = _1369_ & _1676_ /*9437*/;
assign _1674_ = _1369_ ^ _1676_ /*9440*/;
assign _1675_ = _1667_ & _1674_ /*9438*/;
assign _1563_ = _1667_ ^ _1674_ /*9439*/;
assign _1672_ = _1673_ | _1675_ /*9436*/;
assign _1681_ = D[20] ^ Q[24] /*9435*/;
assign _1678_ = _1370_ & _1681_ /*9431*/;
assign _1679_ = _1370_ ^ _1681_ /*9434*/;
assign _1680_ = _1672_ & _1679_ /*9432*/;
assign _1564_ = _1672_ ^ _1679_ /*9433*/;
assign _1677_ = _1678_ | _1680_ /*9430*/;
assign _1686_ = D[21] ^ Q[24] /*9429*/;
assign _1683_ = _1371_ & _1686_ /*9425*/;
assign _1684_ = _1371_ ^ _1686_ /*9428*/;
assign _1685_ = _1677_ & _1684_ /*9426*/;
assign _1565_ = _1677_ ^ _1684_ /*9427*/;
assign _1682_ = _1683_ | _1685_ /*9424*/;
assign _1691_ = D[22] ^ Q[24] /*9423*/;
assign _1688_ = _1372_ & _1691_ /*9419*/;
assign _1689_ = _1372_ ^ _1691_ /*9422*/;
assign _1690_ = _1682_ & _1689_ /*9420*/;
assign _1566_ = _1682_ ^ _1689_ /*9421*/;
assign _1687_ = _1688_ | _1690_ /*9418*/;
assign _1696_ = D[23] ^ Q[24] /*9417*/;
assign _1693_ = _1373_ & _1696_ /*9413*/;
assign _1694_ = _1373_ ^ _1696_ /*9416*/;
assign _1695_ = _1687_ & _1694_ /*9414*/;
assign _1567_ = _1687_ ^ _1694_ /*9415*/;
assign _1692_ = _1693_ | _1695_ /*9412*/;
assign _1701_ = D[24] ^ Q[24] /*9411*/;
assign _1698_ = _1374_ & _1701_ /*9407*/;
assign _1699_ = _1374_ ^ _1701_ /*9410*/;
assign _1700_ = _1692_ & _1699_ /*9408*/;
assign _1568_ = _1692_ ^ _1699_ /*9409*/;
assign _1697_ = _1698_ | _1700_ /*9406*/;
assign _1706_ = D[25] ^ Q[24] /*9405*/;
assign _1703_ = _1375_ & _1706_ /*9401*/;
assign _1704_ = _1375_ ^ _1706_ /*9404*/;
assign _1705_ = _1697_ & _1704_ /*9402*/;
assign _1569_ = _1697_ ^ _1704_ /*9403*/;
assign _1702_ = _1703_ | _1705_ /*9400*/;
assign _1711_ = D[26] ^ Q[24] /*9399*/;
assign _1708_ = _1376_ & _1711_ /*9395*/;
assign _1709_ = _1376_ ^ _1711_ /*9398*/;
assign _1710_ = _1702_ & _1709_ /*9396*/;
assign _1570_ = _1702_ ^ _1709_ /*9397*/;
assign _1707_ = _1708_ | _1710_ /*9394*/;
assign _1716_ = D[27] ^ Q[24] /*9393*/;
assign _1713_ = _1377_ & _1716_ /*9389*/;
assign _1714_ = _1377_ ^ _1716_ /*9392*/;
assign _1715_ = _1707_ & _1714_ /*9390*/;
assign _1571_ = _1707_ ^ _1714_ /*9391*/;
assign _1712_ = _1713_ | _1715_ /*9388*/;
assign _1721_ = D[28] ^ Q[24] /*9387*/;
assign _1718_ = _1378_ & _1721_ /*9383*/;
assign _1719_ = _1378_ ^ _1721_ /*9386*/;
assign _1720_ = _1712_ & _1719_ /*9384*/;
assign _1572_ = _1712_ ^ _1719_ /*9385*/;
assign _1717_ = _1718_ | _1720_ /*9382*/;
assign _1726_ = D[29] ^ Q[24] /*9381*/;
assign _1723_ = _1379_ & _1726_ /*9377*/;
assign _1724_ = _1379_ ^ _1726_ /*9380*/;
assign _1725_ = _1717_ & _1724_ /*9378*/;
assign _1573_ = _1717_ ^ _1724_ /*9379*/;
assign _1722_ = _1723_ | _1725_ /*9376*/;
assign _1731_ = D[30] ^ Q[24] /*9375*/;
assign _1728_ = _1380_ & _1731_ /*9371*/;
assign _1729_ = _1380_ ^ _1731_ /*9374*/;
assign _1730_ = _1722_ & _1729_ /*9372*/;
assign _1574_ = _1722_ ^ _1729_ /*9373*/;
assign _1727_ = _1728_ | _1730_ /*9370*/;
assign _1735_ = zeroWire ^ Q[24] /*9369*/;
assign _1732_ = _1381_ & _1735_ /*9365*/;
assign _1733_ = _1381_ ^ _1735_ /*9368*/;
assign _1734_ = _1727_ & _1733_ /*9366*/;
assign _1575_ = _1727_ ^ _1733_ /*9367*/;
assign Q[23] = _1732_ | _1734_ /*9364*/;
assign _1774_ = D[0] ^ Q[23] /*9170*/;
assign _1771_ = R_0[22] & _1774_ /*9166*/;
assign _1772_ = R_0[22] ^ _1774_ /*9169*/;
assign _1773_ = Q[23] & _1772_ /*9167*/;
assign _1737_ = Q[23] ^ _1772_ /*9168*/;
assign _1770_ = _1771_ | _1773_ /*9165*/;
assign _1779_ = D[1] ^ Q[23] /*9164*/;
assign _1776_ = _1544_ & _1779_ /*9160*/;
assign _1777_ = _1544_ ^ _1779_ /*9163*/;
assign _1778_ = _1770_ & _1777_ /*9161*/;
assign _1738_ = _1770_ ^ _1777_ /*9162*/;
assign _1775_ = _1776_ | _1778_ /*9159*/;
assign _1784_ = D[2] ^ Q[23] /*9158*/;
assign _1781_ = _1545_ & _1784_ /*9154*/;
assign _1782_ = _1545_ ^ _1784_ /*9157*/;
assign _1783_ = _1775_ & _1782_ /*9155*/;
assign _1739_ = _1775_ ^ _1782_ /*9156*/;
assign _1780_ = _1781_ | _1783_ /*9153*/;
assign _1789_ = D[3] ^ Q[23] /*9152*/;
assign _1786_ = _1546_ & _1789_ /*9148*/;
assign _1787_ = _1546_ ^ _1789_ /*9151*/;
assign _1788_ = _1780_ & _1787_ /*9149*/;
assign _1740_ = _1780_ ^ _1787_ /*9150*/;
assign _1785_ = _1786_ | _1788_ /*9147*/;
assign _1794_ = D[4] ^ Q[23] /*9146*/;
assign _1791_ = _1547_ & _1794_ /*9142*/;
assign _1792_ = _1547_ ^ _1794_ /*9145*/;
assign _1793_ = _1785_ & _1792_ /*9143*/;
assign _1741_ = _1785_ ^ _1792_ /*9144*/;
assign _1790_ = _1791_ | _1793_ /*9141*/;
assign _1799_ = D[5] ^ Q[23] /*9140*/;
assign _1796_ = _1548_ & _1799_ /*9136*/;
assign _1797_ = _1548_ ^ _1799_ /*9139*/;
assign _1798_ = _1790_ & _1797_ /*9137*/;
assign _1742_ = _1790_ ^ _1797_ /*9138*/;
assign _1795_ = _1796_ | _1798_ /*9135*/;
assign _1804_ = D[6] ^ Q[23] /*9134*/;
assign _1801_ = _1549_ & _1804_ /*9130*/;
assign _1802_ = _1549_ ^ _1804_ /*9133*/;
assign _1803_ = _1795_ & _1802_ /*9131*/;
assign _1743_ = _1795_ ^ _1802_ /*9132*/;
assign _1800_ = _1801_ | _1803_ /*9129*/;
assign _1809_ = D[7] ^ Q[23] /*9128*/;
assign _1806_ = _1550_ & _1809_ /*9124*/;
assign _1807_ = _1550_ ^ _1809_ /*9127*/;
assign _1808_ = _1800_ & _1807_ /*9125*/;
assign _1744_ = _1800_ ^ _1807_ /*9126*/;
assign _1805_ = _1806_ | _1808_ /*9123*/;
assign _1814_ = D[8] ^ Q[23] /*9122*/;
assign _1811_ = _1551_ & _1814_ /*9118*/;
assign _1812_ = _1551_ ^ _1814_ /*9121*/;
assign _1813_ = _1805_ & _1812_ /*9119*/;
assign _1745_ = _1805_ ^ _1812_ /*9120*/;
assign _1810_ = _1811_ | _1813_ /*9117*/;
assign _1819_ = D[9] ^ Q[23] /*9116*/;
assign _1816_ = _1552_ & _1819_ /*9112*/;
assign _1817_ = _1552_ ^ _1819_ /*9115*/;
assign _1818_ = _1810_ & _1817_ /*9113*/;
assign _1746_ = _1810_ ^ _1817_ /*9114*/;
assign _1815_ = _1816_ | _1818_ /*9111*/;
assign _1824_ = D[10] ^ Q[23] /*9110*/;
assign _1821_ = _1553_ & _1824_ /*9106*/;
assign _1822_ = _1553_ ^ _1824_ /*9109*/;
assign _1823_ = _1815_ & _1822_ /*9107*/;
assign _1747_ = _1815_ ^ _1822_ /*9108*/;
assign _1820_ = _1821_ | _1823_ /*9105*/;
assign _1829_ = D[11] ^ Q[23] /*9104*/;
assign _1826_ = _1554_ & _1829_ /*9100*/;
assign _1827_ = _1554_ ^ _1829_ /*9103*/;
assign _1828_ = _1820_ & _1827_ /*9101*/;
assign _1748_ = _1820_ ^ _1827_ /*9102*/;
assign _1825_ = _1826_ | _1828_ /*9099*/;
assign _1834_ = D[12] ^ Q[23] /*9098*/;
assign _1831_ = _1555_ & _1834_ /*9094*/;
assign _1832_ = _1555_ ^ _1834_ /*9097*/;
assign _1833_ = _1825_ & _1832_ /*9095*/;
assign _1749_ = _1825_ ^ _1832_ /*9096*/;
assign _1830_ = _1831_ | _1833_ /*9093*/;
assign _1839_ = D[13] ^ Q[23] /*9092*/;
assign _1836_ = _1556_ & _1839_ /*9088*/;
assign _1837_ = _1556_ ^ _1839_ /*9091*/;
assign _1838_ = _1830_ & _1837_ /*9089*/;
assign _1750_ = _1830_ ^ _1837_ /*9090*/;
assign _1835_ = _1836_ | _1838_ /*9087*/;
assign _1844_ = D[14] ^ Q[23] /*9086*/;
assign _1841_ = _1557_ & _1844_ /*9082*/;
assign _1842_ = _1557_ ^ _1844_ /*9085*/;
assign _1843_ = _1835_ & _1842_ /*9083*/;
assign _1751_ = _1835_ ^ _1842_ /*9084*/;
assign _1840_ = _1841_ | _1843_ /*9081*/;
assign _1849_ = D[15] ^ Q[23] /*9080*/;
assign _1846_ = _1558_ & _1849_ /*9076*/;
assign _1847_ = _1558_ ^ _1849_ /*9079*/;
assign _1848_ = _1840_ & _1847_ /*9077*/;
assign _1752_ = _1840_ ^ _1847_ /*9078*/;
assign _1845_ = _1846_ | _1848_ /*9075*/;
assign _1854_ = D[16] ^ Q[23] /*9074*/;
assign _1851_ = _1559_ & _1854_ /*9070*/;
assign _1852_ = _1559_ ^ _1854_ /*9073*/;
assign _1853_ = _1845_ & _1852_ /*9071*/;
assign _1753_ = _1845_ ^ _1852_ /*9072*/;
assign _1850_ = _1851_ | _1853_ /*9069*/;
assign _1859_ = D[17] ^ Q[23] /*9068*/;
assign _1856_ = _1560_ & _1859_ /*9064*/;
assign _1857_ = _1560_ ^ _1859_ /*9067*/;
assign _1858_ = _1850_ & _1857_ /*9065*/;
assign _1754_ = _1850_ ^ _1857_ /*9066*/;
assign _1855_ = _1856_ | _1858_ /*9063*/;
assign _1864_ = D[18] ^ Q[23] /*9062*/;
assign _1861_ = _1561_ & _1864_ /*9058*/;
assign _1862_ = _1561_ ^ _1864_ /*9061*/;
assign _1863_ = _1855_ & _1862_ /*9059*/;
assign _1755_ = _1855_ ^ _1862_ /*9060*/;
assign _1860_ = _1861_ | _1863_ /*9057*/;
assign _1869_ = D[19] ^ Q[23] /*9056*/;
assign _1866_ = _1562_ & _1869_ /*9052*/;
assign _1867_ = _1562_ ^ _1869_ /*9055*/;
assign _1868_ = _1860_ & _1867_ /*9053*/;
assign _1756_ = _1860_ ^ _1867_ /*9054*/;
assign _1865_ = _1866_ | _1868_ /*9051*/;
assign _1874_ = D[20] ^ Q[23] /*9050*/;
assign _1871_ = _1563_ & _1874_ /*9046*/;
assign _1872_ = _1563_ ^ _1874_ /*9049*/;
assign _1873_ = _1865_ & _1872_ /*9047*/;
assign _1757_ = _1865_ ^ _1872_ /*9048*/;
assign _1870_ = _1871_ | _1873_ /*9045*/;
assign _1879_ = D[21] ^ Q[23] /*9044*/;
assign _1876_ = _1564_ & _1879_ /*9040*/;
assign _1877_ = _1564_ ^ _1879_ /*9043*/;
assign _1878_ = _1870_ & _1877_ /*9041*/;
assign _1758_ = _1870_ ^ _1877_ /*9042*/;
assign _1875_ = _1876_ | _1878_ /*9039*/;
assign _1884_ = D[22] ^ Q[23] /*9038*/;
assign _1881_ = _1565_ & _1884_ /*9034*/;
assign _1882_ = _1565_ ^ _1884_ /*9037*/;
assign _1883_ = _1875_ & _1882_ /*9035*/;
assign _1759_ = _1875_ ^ _1882_ /*9036*/;
assign _1880_ = _1881_ | _1883_ /*9033*/;
assign _1889_ = D[23] ^ Q[23] /*9032*/;
assign _1886_ = _1566_ & _1889_ /*9028*/;
assign _1887_ = _1566_ ^ _1889_ /*9031*/;
assign _1888_ = _1880_ & _1887_ /*9029*/;
assign _1760_ = _1880_ ^ _1887_ /*9030*/;
assign _1885_ = _1886_ | _1888_ /*9027*/;
assign _1894_ = D[24] ^ Q[23] /*9026*/;
assign _1891_ = _1567_ & _1894_ /*9022*/;
assign _1892_ = _1567_ ^ _1894_ /*9025*/;
assign _1893_ = _1885_ & _1892_ /*9023*/;
assign _1761_ = _1885_ ^ _1892_ /*9024*/;
assign _1890_ = _1891_ | _1893_ /*9021*/;
assign _1899_ = D[25] ^ Q[23] /*9020*/;
assign _1896_ = _1568_ & _1899_ /*9016*/;
assign _1897_ = _1568_ ^ _1899_ /*9019*/;
assign _1898_ = _1890_ & _1897_ /*9017*/;
assign _1762_ = _1890_ ^ _1897_ /*9018*/;
assign _1895_ = _1896_ | _1898_ /*9015*/;
assign _1904_ = D[26] ^ Q[23] /*9014*/;
assign _1901_ = _1569_ & _1904_ /*9010*/;
assign _1902_ = _1569_ ^ _1904_ /*9013*/;
assign _1903_ = _1895_ & _1902_ /*9011*/;
assign _1763_ = _1895_ ^ _1902_ /*9012*/;
assign _1900_ = _1901_ | _1903_ /*9009*/;
assign _1909_ = D[27] ^ Q[23] /*9008*/;
assign _1906_ = _1570_ & _1909_ /*9004*/;
assign _1907_ = _1570_ ^ _1909_ /*9007*/;
assign _1908_ = _1900_ & _1907_ /*9005*/;
assign _1764_ = _1900_ ^ _1907_ /*9006*/;
assign _1905_ = _1906_ | _1908_ /*9003*/;
assign _1914_ = D[28] ^ Q[23] /*9002*/;
assign _1911_ = _1571_ & _1914_ /*8998*/;
assign _1912_ = _1571_ ^ _1914_ /*9001*/;
assign _1913_ = _1905_ & _1912_ /*8999*/;
assign _1765_ = _1905_ ^ _1912_ /*9000*/;
assign _1910_ = _1911_ | _1913_ /*8997*/;
assign _1919_ = D[29] ^ Q[23] /*8996*/;
assign _1916_ = _1572_ & _1919_ /*8992*/;
assign _1917_ = _1572_ ^ _1919_ /*8995*/;
assign _1918_ = _1910_ & _1917_ /*8993*/;
assign _1766_ = _1910_ ^ _1917_ /*8994*/;
assign _1915_ = _1916_ | _1918_ /*8991*/;
assign _1924_ = D[30] ^ Q[23] /*8990*/;
assign _1921_ = _1573_ & _1924_ /*8986*/;
assign _1922_ = _1573_ ^ _1924_ /*8989*/;
assign _1923_ = _1915_ & _1922_ /*8987*/;
assign _1767_ = _1915_ ^ _1922_ /*8988*/;
assign _1920_ = _1921_ | _1923_ /*8985*/;
assign _1928_ = zeroWire ^ Q[23] /*8984*/;
assign _1925_ = _1574_ & _1928_ /*8980*/;
assign _1926_ = _1574_ ^ _1928_ /*8983*/;
assign _1927_ = _1920_ & _1926_ /*8981*/;
assign _1768_ = _1920_ ^ _1926_ /*8982*/;
assign Q[22] = _1925_ | _1927_ /*8979*/;
assign _1967_ = D[0] ^ Q[22] /*8785*/;
assign _1964_ = R_0[21] & _1967_ /*8781*/;
assign _1965_ = R_0[21] ^ _1967_ /*8784*/;
assign _1966_ = Q[22] & _1965_ /*8782*/;
assign _1930_ = Q[22] ^ _1965_ /*8783*/;
assign _1963_ = _1964_ | _1966_ /*8780*/;
assign _1972_ = D[1] ^ Q[22] /*8779*/;
assign _1969_ = _1737_ & _1972_ /*8775*/;
assign _1970_ = _1737_ ^ _1972_ /*8778*/;
assign _1971_ = _1963_ & _1970_ /*8776*/;
assign _1931_ = _1963_ ^ _1970_ /*8777*/;
assign _1968_ = _1969_ | _1971_ /*8774*/;
assign _1977_ = D[2] ^ Q[22] /*8773*/;
assign _1974_ = _1738_ & _1977_ /*8769*/;
assign _1975_ = _1738_ ^ _1977_ /*8772*/;
assign _1976_ = _1968_ & _1975_ /*8770*/;
assign _1932_ = _1968_ ^ _1975_ /*8771*/;
assign _1973_ = _1974_ | _1976_ /*8768*/;
assign _1982_ = D[3] ^ Q[22] /*8767*/;
assign _1979_ = _1739_ & _1982_ /*8763*/;
assign _1980_ = _1739_ ^ _1982_ /*8766*/;
assign _1981_ = _1973_ & _1980_ /*8764*/;
assign _1933_ = _1973_ ^ _1980_ /*8765*/;
assign _1978_ = _1979_ | _1981_ /*8762*/;
assign _1987_ = D[4] ^ Q[22] /*8761*/;
assign _1984_ = _1740_ & _1987_ /*8757*/;
assign _1985_ = _1740_ ^ _1987_ /*8760*/;
assign _1986_ = _1978_ & _1985_ /*8758*/;
assign _1934_ = _1978_ ^ _1985_ /*8759*/;
assign _1983_ = _1984_ | _1986_ /*8756*/;
assign _1992_ = D[5] ^ Q[22] /*8755*/;
assign _1989_ = _1741_ & _1992_ /*8751*/;
assign _1990_ = _1741_ ^ _1992_ /*8754*/;
assign _1991_ = _1983_ & _1990_ /*8752*/;
assign _1935_ = _1983_ ^ _1990_ /*8753*/;
assign _1988_ = _1989_ | _1991_ /*8750*/;
assign _1997_ = D[6] ^ Q[22] /*8749*/;
assign _1994_ = _1742_ & _1997_ /*8745*/;
assign _1995_ = _1742_ ^ _1997_ /*8748*/;
assign _1996_ = _1988_ & _1995_ /*8746*/;
assign _1936_ = _1988_ ^ _1995_ /*8747*/;
assign _1993_ = _1994_ | _1996_ /*8744*/;
assign _2002_ = D[7] ^ Q[22] /*8743*/;
assign _1999_ = _1743_ & _2002_ /*8739*/;
assign _2000_ = _1743_ ^ _2002_ /*8742*/;
assign _2001_ = _1993_ & _2000_ /*8740*/;
assign _1937_ = _1993_ ^ _2000_ /*8741*/;
assign _1998_ = _1999_ | _2001_ /*8738*/;
assign _2007_ = D[8] ^ Q[22] /*8737*/;
assign _2004_ = _1744_ & _2007_ /*8733*/;
assign _2005_ = _1744_ ^ _2007_ /*8736*/;
assign _2006_ = _1998_ & _2005_ /*8734*/;
assign _1938_ = _1998_ ^ _2005_ /*8735*/;
assign _2003_ = _2004_ | _2006_ /*8732*/;
assign _2012_ = D[9] ^ Q[22] /*8731*/;
assign _2009_ = _1745_ & _2012_ /*8727*/;
assign _2010_ = _1745_ ^ _2012_ /*8730*/;
assign _2011_ = _2003_ & _2010_ /*8728*/;
assign _1939_ = _2003_ ^ _2010_ /*8729*/;
assign _2008_ = _2009_ | _2011_ /*8726*/;
assign _2017_ = D[10] ^ Q[22] /*8725*/;
assign _2014_ = _1746_ & _2017_ /*8721*/;
assign _2015_ = _1746_ ^ _2017_ /*8724*/;
assign _2016_ = _2008_ & _2015_ /*8722*/;
assign _1940_ = _2008_ ^ _2015_ /*8723*/;
assign _2013_ = _2014_ | _2016_ /*8720*/;
assign _2022_ = D[11] ^ Q[22] /*8719*/;
assign _2019_ = _1747_ & _2022_ /*8715*/;
assign _2020_ = _1747_ ^ _2022_ /*8718*/;
assign _2021_ = _2013_ & _2020_ /*8716*/;
assign _1941_ = _2013_ ^ _2020_ /*8717*/;
assign _2018_ = _2019_ | _2021_ /*8714*/;
assign _2027_ = D[12] ^ Q[22] /*8713*/;
assign _2024_ = _1748_ & _2027_ /*8709*/;
assign _2025_ = _1748_ ^ _2027_ /*8712*/;
assign _2026_ = _2018_ & _2025_ /*8710*/;
assign _1942_ = _2018_ ^ _2025_ /*8711*/;
assign _2023_ = _2024_ | _2026_ /*8708*/;
assign _2032_ = D[13] ^ Q[22] /*8707*/;
assign _2029_ = _1749_ & _2032_ /*8703*/;
assign _2030_ = _1749_ ^ _2032_ /*8706*/;
assign _2031_ = _2023_ & _2030_ /*8704*/;
assign _1943_ = _2023_ ^ _2030_ /*8705*/;
assign _2028_ = _2029_ | _2031_ /*8702*/;
assign _2037_ = D[14] ^ Q[22] /*8701*/;
assign _2034_ = _1750_ & _2037_ /*8697*/;
assign _2035_ = _1750_ ^ _2037_ /*8700*/;
assign _2036_ = _2028_ & _2035_ /*8698*/;
assign _1944_ = _2028_ ^ _2035_ /*8699*/;
assign _2033_ = _2034_ | _2036_ /*8696*/;
assign _2042_ = D[15] ^ Q[22] /*8695*/;
assign _2039_ = _1751_ & _2042_ /*8691*/;
assign _2040_ = _1751_ ^ _2042_ /*8694*/;
assign _2041_ = _2033_ & _2040_ /*8692*/;
assign _1945_ = _2033_ ^ _2040_ /*8693*/;
assign _2038_ = _2039_ | _2041_ /*8690*/;
assign _2047_ = D[16] ^ Q[22] /*8689*/;
assign _2044_ = _1752_ & _2047_ /*8685*/;
assign _2045_ = _1752_ ^ _2047_ /*8688*/;
assign _2046_ = _2038_ & _2045_ /*8686*/;
assign _1946_ = _2038_ ^ _2045_ /*8687*/;
assign _2043_ = _2044_ | _2046_ /*8684*/;
assign _2052_ = D[17] ^ Q[22] /*8683*/;
assign _2049_ = _1753_ & _2052_ /*8679*/;
assign _2050_ = _1753_ ^ _2052_ /*8682*/;
assign _2051_ = _2043_ & _2050_ /*8680*/;
assign _1947_ = _2043_ ^ _2050_ /*8681*/;
assign _2048_ = _2049_ | _2051_ /*8678*/;
assign _2057_ = D[18] ^ Q[22] /*8677*/;
assign _2054_ = _1754_ & _2057_ /*8673*/;
assign _2055_ = _1754_ ^ _2057_ /*8676*/;
assign _2056_ = _2048_ & _2055_ /*8674*/;
assign _1948_ = _2048_ ^ _2055_ /*8675*/;
assign _2053_ = _2054_ | _2056_ /*8672*/;
assign _2062_ = D[19] ^ Q[22] /*8671*/;
assign _2059_ = _1755_ & _2062_ /*8667*/;
assign _2060_ = _1755_ ^ _2062_ /*8670*/;
assign _2061_ = _2053_ & _2060_ /*8668*/;
assign _1949_ = _2053_ ^ _2060_ /*8669*/;
assign _2058_ = _2059_ | _2061_ /*8666*/;
assign _2067_ = D[20] ^ Q[22] /*8665*/;
assign _2064_ = _1756_ & _2067_ /*8661*/;
assign _2065_ = _1756_ ^ _2067_ /*8664*/;
assign _2066_ = _2058_ & _2065_ /*8662*/;
assign _1950_ = _2058_ ^ _2065_ /*8663*/;
assign _2063_ = _2064_ | _2066_ /*8660*/;
assign _2072_ = D[21] ^ Q[22] /*8659*/;
assign _2069_ = _1757_ & _2072_ /*8655*/;
assign _2070_ = _1757_ ^ _2072_ /*8658*/;
assign _2071_ = _2063_ & _2070_ /*8656*/;
assign _1951_ = _2063_ ^ _2070_ /*8657*/;
assign _2068_ = _2069_ | _2071_ /*8654*/;
assign _2077_ = D[22] ^ Q[22] /*8653*/;
assign _2074_ = _1758_ & _2077_ /*8649*/;
assign _2075_ = _1758_ ^ _2077_ /*8652*/;
assign _2076_ = _2068_ & _2075_ /*8650*/;
assign _1952_ = _2068_ ^ _2075_ /*8651*/;
assign _2073_ = _2074_ | _2076_ /*8648*/;
assign _2082_ = D[23] ^ Q[22] /*8647*/;
assign _2079_ = _1759_ & _2082_ /*8643*/;
assign _2080_ = _1759_ ^ _2082_ /*8646*/;
assign _2081_ = _2073_ & _2080_ /*8644*/;
assign _1953_ = _2073_ ^ _2080_ /*8645*/;
assign _2078_ = _2079_ | _2081_ /*8642*/;
assign _2087_ = D[24] ^ Q[22] /*8641*/;
assign _2084_ = _1760_ & _2087_ /*8637*/;
assign _2085_ = _1760_ ^ _2087_ /*8640*/;
assign _2086_ = _2078_ & _2085_ /*8638*/;
assign _1954_ = _2078_ ^ _2085_ /*8639*/;
assign _2083_ = _2084_ | _2086_ /*8636*/;
assign _2092_ = D[25] ^ Q[22] /*8635*/;
assign _2089_ = _1761_ & _2092_ /*8631*/;
assign _2090_ = _1761_ ^ _2092_ /*8634*/;
assign _2091_ = _2083_ & _2090_ /*8632*/;
assign _1955_ = _2083_ ^ _2090_ /*8633*/;
assign _2088_ = _2089_ | _2091_ /*8630*/;
assign _2097_ = D[26] ^ Q[22] /*8629*/;
assign _2094_ = _1762_ & _2097_ /*8625*/;
assign _2095_ = _1762_ ^ _2097_ /*8628*/;
assign _2096_ = _2088_ & _2095_ /*8626*/;
assign _1956_ = _2088_ ^ _2095_ /*8627*/;
assign _2093_ = _2094_ | _2096_ /*8624*/;
assign _2102_ = D[27] ^ Q[22] /*8623*/;
assign _2099_ = _1763_ & _2102_ /*8619*/;
assign _2100_ = _1763_ ^ _2102_ /*8622*/;
assign _2101_ = _2093_ & _2100_ /*8620*/;
assign _1957_ = _2093_ ^ _2100_ /*8621*/;
assign _2098_ = _2099_ | _2101_ /*8618*/;
assign _2107_ = D[28] ^ Q[22] /*8617*/;
assign _2104_ = _1764_ & _2107_ /*8613*/;
assign _2105_ = _1764_ ^ _2107_ /*8616*/;
assign _2106_ = _2098_ & _2105_ /*8614*/;
assign _1958_ = _2098_ ^ _2105_ /*8615*/;
assign _2103_ = _2104_ | _2106_ /*8612*/;
assign _2112_ = D[29] ^ Q[22] /*8611*/;
assign _2109_ = _1765_ & _2112_ /*8607*/;
assign _2110_ = _1765_ ^ _2112_ /*8610*/;
assign _2111_ = _2103_ & _2110_ /*8608*/;
assign _1959_ = _2103_ ^ _2110_ /*8609*/;
assign _2108_ = _2109_ | _2111_ /*8606*/;
assign _2117_ = D[30] ^ Q[22] /*8605*/;
assign _2114_ = _1766_ & _2117_ /*8601*/;
assign _2115_ = _1766_ ^ _2117_ /*8604*/;
assign _2116_ = _2108_ & _2115_ /*8602*/;
assign _1960_ = _2108_ ^ _2115_ /*8603*/;
assign _2113_ = _2114_ | _2116_ /*8600*/;
assign _2121_ = zeroWire ^ Q[22] /*8599*/;
assign _2118_ = _1767_ & _2121_ /*8595*/;
assign _2119_ = _1767_ ^ _2121_ /*8598*/;
assign _2120_ = _2113_ & _2119_ /*8596*/;
assign _1961_ = _2113_ ^ _2119_ /*8597*/;
assign Q[21] = _2118_ | _2120_ /*8594*/;
assign _2160_ = D[0] ^ Q[21] /*8400*/;
assign _2157_ = R_0[20] & _2160_ /*8396*/;
assign _2158_ = R_0[20] ^ _2160_ /*8399*/;
assign _2159_ = Q[21] & _2158_ /*8397*/;
assign _2123_ = Q[21] ^ _2158_ /*8398*/;
assign _2156_ = _2157_ | _2159_ /*8395*/;
assign _2165_ = D[1] ^ Q[21] /*8394*/;
assign _2162_ = _1930_ & _2165_ /*8390*/;
assign _2163_ = _1930_ ^ _2165_ /*8393*/;
assign _2164_ = _2156_ & _2163_ /*8391*/;
assign _2124_ = _2156_ ^ _2163_ /*8392*/;
assign _2161_ = _2162_ | _2164_ /*8389*/;
assign _2170_ = D[2] ^ Q[21] /*8388*/;
assign _2167_ = _1931_ & _2170_ /*8384*/;
assign _2168_ = _1931_ ^ _2170_ /*8387*/;
assign _2169_ = _2161_ & _2168_ /*8385*/;
assign _2125_ = _2161_ ^ _2168_ /*8386*/;
assign _2166_ = _2167_ | _2169_ /*8383*/;
assign _2175_ = D[3] ^ Q[21] /*8382*/;
assign _2172_ = _1932_ & _2175_ /*8378*/;
assign _2173_ = _1932_ ^ _2175_ /*8381*/;
assign _2174_ = _2166_ & _2173_ /*8379*/;
assign _2126_ = _2166_ ^ _2173_ /*8380*/;
assign _2171_ = _2172_ | _2174_ /*8377*/;
assign _2180_ = D[4] ^ Q[21] /*8376*/;
assign _2177_ = _1933_ & _2180_ /*8372*/;
assign _2178_ = _1933_ ^ _2180_ /*8375*/;
assign _2179_ = _2171_ & _2178_ /*8373*/;
assign _2127_ = _2171_ ^ _2178_ /*8374*/;
assign _2176_ = _2177_ | _2179_ /*8371*/;
assign _2185_ = D[5] ^ Q[21] /*8370*/;
assign _2182_ = _1934_ & _2185_ /*8366*/;
assign _2183_ = _1934_ ^ _2185_ /*8369*/;
assign _2184_ = _2176_ & _2183_ /*8367*/;
assign _2128_ = _2176_ ^ _2183_ /*8368*/;
assign _2181_ = _2182_ | _2184_ /*8365*/;
assign _2190_ = D[6] ^ Q[21] /*8364*/;
assign _2187_ = _1935_ & _2190_ /*8360*/;
assign _2188_ = _1935_ ^ _2190_ /*8363*/;
assign _2189_ = _2181_ & _2188_ /*8361*/;
assign _2129_ = _2181_ ^ _2188_ /*8362*/;
assign _2186_ = _2187_ | _2189_ /*8359*/;
assign _2195_ = D[7] ^ Q[21] /*8358*/;
assign _2192_ = _1936_ & _2195_ /*8354*/;
assign _2193_ = _1936_ ^ _2195_ /*8357*/;
assign _2194_ = _2186_ & _2193_ /*8355*/;
assign _2130_ = _2186_ ^ _2193_ /*8356*/;
assign _2191_ = _2192_ | _2194_ /*8353*/;
assign _2200_ = D[8] ^ Q[21] /*8352*/;
assign _2197_ = _1937_ & _2200_ /*8348*/;
assign _2198_ = _1937_ ^ _2200_ /*8351*/;
assign _2199_ = _2191_ & _2198_ /*8349*/;
assign _2131_ = _2191_ ^ _2198_ /*8350*/;
assign _2196_ = _2197_ | _2199_ /*8347*/;
assign _2205_ = D[9] ^ Q[21] /*8346*/;
assign _2202_ = _1938_ & _2205_ /*8342*/;
assign _2203_ = _1938_ ^ _2205_ /*8345*/;
assign _2204_ = _2196_ & _2203_ /*8343*/;
assign _2132_ = _2196_ ^ _2203_ /*8344*/;
assign _2201_ = _2202_ | _2204_ /*8341*/;
assign _2210_ = D[10] ^ Q[21] /*8340*/;
assign _2207_ = _1939_ & _2210_ /*8336*/;
assign _2208_ = _1939_ ^ _2210_ /*8339*/;
assign _2209_ = _2201_ & _2208_ /*8337*/;
assign _2133_ = _2201_ ^ _2208_ /*8338*/;
assign _2206_ = _2207_ | _2209_ /*8335*/;
assign _2215_ = D[11] ^ Q[21] /*8334*/;
assign _2212_ = _1940_ & _2215_ /*8330*/;
assign _2213_ = _1940_ ^ _2215_ /*8333*/;
assign _2214_ = _2206_ & _2213_ /*8331*/;
assign _2134_ = _2206_ ^ _2213_ /*8332*/;
assign _2211_ = _2212_ | _2214_ /*8329*/;
assign _2220_ = D[12] ^ Q[21] /*8328*/;
assign _2217_ = _1941_ & _2220_ /*8324*/;
assign _2218_ = _1941_ ^ _2220_ /*8327*/;
assign _2219_ = _2211_ & _2218_ /*8325*/;
assign _2135_ = _2211_ ^ _2218_ /*8326*/;
assign _2216_ = _2217_ | _2219_ /*8323*/;
assign _2225_ = D[13] ^ Q[21] /*8322*/;
assign _2222_ = _1942_ & _2225_ /*8318*/;
assign _2223_ = _1942_ ^ _2225_ /*8321*/;
assign _2224_ = _2216_ & _2223_ /*8319*/;
assign _2136_ = _2216_ ^ _2223_ /*8320*/;
assign _2221_ = _2222_ | _2224_ /*8317*/;
assign _2230_ = D[14] ^ Q[21] /*8316*/;
assign _2227_ = _1943_ & _2230_ /*8312*/;
assign _2228_ = _1943_ ^ _2230_ /*8315*/;
assign _2229_ = _2221_ & _2228_ /*8313*/;
assign _2137_ = _2221_ ^ _2228_ /*8314*/;
assign _2226_ = _2227_ | _2229_ /*8311*/;
assign _2235_ = D[15] ^ Q[21] /*8310*/;
assign _2232_ = _1944_ & _2235_ /*8306*/;
assign _2233_ = _1944_ ^ _2235_ /*8309*/;
assign _2234_ = _2226_ & _2233_ /*8307*/;
assign _2138_ = _2226_ ^ _2233_ /*8308*/;
assign _2231_ = _2232_ | _2234_ /*8305*/;
assign _2240_ = D[16] ^ Q[21] /*8304*/;
assign _2237_ = _1945_ & _2240_ /*8300*/;
assign _2238_ = _1945_ ^ _2240_ /*8303*/;
assign _2239_ = _2231_ & _2238_ /*8301*/;
assign _2139_ = _2231_ ^ _2238_ /*8302*/;
assign _2236_ = _2237_ | _2239_ /*8299*/;
assign _2245_ = D[17] ^ Q[21] /*8298*/;
assign _2242_ = _1946_ & _2245_ /*8294*/;
assign _2243_ = _1946_ ^ _2245_ /*8297*/;
assign _2244_ = _2236_ & _2243_ /*8295*/;
assign _2140_ = _2236_ ^ _2243_ /*8296*/;
assign _2241_ = _2242_ | _2244_ /*8293*/;
assign _2250_ = D[18] ^ Q[21] /*8292*/;
assign _2247_ = _1947_ & _2250_ /*8288*/;
assign _2248_ = _1947_ ^ _2250_ /*8291*/;
assign _2249_ = _2241_ & _2248_ /*8289*/;
assign _2141_ = _2241_ ^ _2248_ /*8290*/;
assign _2246_ = _2247_ | _2249_ /*8287*/;
assign _2255_ = D[19] ^ Q[21] /*8286*/;
assign _2252_ = _1948_ & _2255_ /*8282*/;
assign _2253_ = _1948_ ^ _2255_ /*8285*/;
assign _2254_ = _2246_ & _2253_ /*8283*/;
assign _2142_ = _2246_ ^ _2253_ /*8284*/;
assign _2251_ = _2252_ | _2254_ /*8281*/;
assign _2260_ = D[20] ^ Q[21] /*8280*/;
assign _2257_ = _1949_ & _2260_ /*8276*/;
assign _2258_ = _1949_ ^ _2260_ /*8279*/;
assign _2259_ = _2251_ & _2258_ /*8277*/;
assign _2143_ = _2251_ ^ _2258_ /*8278*/;
assign _2256_ = _2257_ | _2259_ /*8275*/;
assign _2265_ = D[21] ^ Q[21] /*8274*/;
assign _2262_ = _1950_ & _2265_ /*8270*/;
assign _2263_ = _1950_ ^ _2265_ /*8273*/;
assign _2264_ = _2256_ & _2263_ /*8271*/;
assign _2144_ = _2256_ ^ _2263_ /*8272*/;
assign _2261_ = _2262_ | _2264_ /*8269*/;
assign _2270_ = D[22] ^ Q[21] /*8268*/;
assign _2267_ = _1951_ & _2270_ /*8264*/;
assign _2268_ = _1951_ ^ _2270_ /*8267*/;
assign _2269_ = _2261_ & _2268_ /*8265*/;
assign _2145_ = _2261_ ^ _2268_ /*8266*/;
assign _2266_ = _2267_ | _2269_ /*8263*/;
assign _2275_ = D[23] ^ Q[21] /*8262*/;
assign _2272_ = _1952_ & _2275_ /*8258*/;
assign _2273_ = _1952_ ^ _2275_ /*8261*/;
assign _2274_ = _2266_ & _2273_ /*8259*/;
assign _2146_ = _2266_ ^ _2273_ /*8260*/;
assign _2271_ = _2272_ | _2274_ /*8257*/;
assign _2280_ = D[24] ^ Q[21] /*8256*/;
assign _2277_ = _1953_ & _2280_ /*8252*/;
assign _2278_ = _1953_ ^ _2280_ /*8255*/;
assign _2279_ = _2271_ & _2278_ /*8253*/;
assign _2147_ = _2271_ ^ _2278_ /*8254*/;
assign _2276_ = _2277_ | _2279_ /*8251*/;
assign _2285_ = D[25] ^ Q[21] /*8250*/;
assign _2282_ = _1954_ & _2285_ /*8246*/;
assign _2283_ = _1954_ ^ _2285_ /*8249*/;
assign _2284_ = _2276_ & _2283_ /*8247*/;
assign _2148_ = _2276_ ^ _2283_ /*8248*/;
assign _2281_ = _2282_ | _2284_ /*8245*/;
assign _2290_ = D[26] ^ Q[21] /*8244*/;
assign _2287_ = _1955_ & _2290_ /*8240*/;
assign _2288_ = _1955_ ^ _2290_ /*8243*/;
assign _2289_ = _2281_ & _2288_ /*8241*/;
assign _2149_ = _2281_ ^ _2288_ /*8242*/;
assign _2286_ = _2287_ | _2289_ /*8239*/;
assign _2295_ = D[27] ^ Q[21] /*8238*/;
assign _2292_ = _1956_ & _2295_ /*8234*/;
assign _2293_ = _1956_ ^ _2295_ /*8237*/;
assign _2294_ = _2286_ & _2293_ /*8235*/;
assign _2150_ = _2286_ ^ _2293_ /*8236*/;
assign _2291_ = _2292_ | _2294_ /*8233*/;
assign _2300_ = D[28] ^ Q[21] /*8232*/;
assign _2297_ = _1957_ & _2300_ /*8228*/;
assign _2298_ = _1957_ ^ _2300_ /*8231*/;
assign _2299_ = _2291_ & _2298_ /*8229*/;
assign _2151_ = _2291_ ^ _2298_ /*8230*/;
assign _2296_ = _2297_ | _2299_ /*8227*/;
assign _2305_ = D[29] ^ Q[21] /*8226*/;
assign _2302_ = _1958_ & _2305_ /*8222*/;
assign _2303_ = _1958_ ^ _2305_ /*8225*/;
assign _2304_ = _2296_ & _2303_ /*8223*/;
assign _2152_ = _2296_ ^ _2303_ /*8224*/;
assign _2301_ = _2302_ | _2304_ /*8221*/;
assign _2310_ = D[30] ^ Q[21] /*8220*/;
assign _2307_ = _1959_ & _2310_ /*8216*/;
assign _2308_ = _1959_ ^ _2310_ /*8219*/;
assign _2309_ = _2301_ & _2308_ /*8217*/;
assign _2153_ = _2301_ ^ _2308_ /*8218*/;
assign _2306_ = _2307_ | _2309_ /*8215*/;
assign _2314_ = zeroWire ^ Q[21] /*8214*/;
assign _2311_ = _1960_ & _2314_ /*8210*/;
assign _2312_ = _1960_ ^ _2314_ /*8213*/;
assign _2313_ = _2306_ & _2312_ /*8211*/;
assign _2154_ = _2306_ ^ _2312_ /*8212*/;
assign Q[20] = _2311_ | _2313_ /*8209*/;
assign _2353_ = D[0] ^ Q[20] /*8015*/;
assign _2350_ = R_0[19] & _2353_ /*8011*/;
assign _2351_ = R_0[19] ^ _2353_ /*8014*/;
assign _2352_ = Q[20] & _2351_ /*8012*/;
assign _2316_ = Q[20] ^ _2351_ /*8013*/;
assign _2349_ = _2350_ | _2352_ /*8010*/;
assign _2358_ = D[1] ^ Q[20] /*8009*/;
assign _2355_ = _2123_ & _2358_ /*8005*/;
assign _2356_ = _2123_ ^ _2358_ /*8008*/;
assign _2357_ = _2349_ & _2356_ /*8006*/;
assign _2317_ = _2349_ ^ _2356_ /*8007*/;
assign _2354_ = _2355_ | _2357_ /*8004*/;
assign _2363_ = D[2] ^ Q[20] /*8003*/;
assign _2360_ = _2124_ & _2363_ /*7999*/;
assign _2361_ = _2124_ ^ _2363_ /*8002*/;
assign _2362_ = _2354_ & _2361_ /*8000*/;
assign _2318_ = _2354_ ^ _2361_ /*8001*/;
assign _2359_ = _2360_ | _2362_ /*7998*/;
assign _2368_ = D[3] ^ Q[20] /*7997*/;
assign _2365_ = _2125_ & _2368_ /*7993*/;
assign _2366_ = _2125_ ^ _2368_ /*7996*/;
assign _2367_ = _2359_ & _2366_ /*7994*/;
assign _2319_ = _2359_ ^ _2366_ /*7995*/;
assign _2364_ = _2365_ | _2367_ /*7992*/;
assign _2373_ = D[4] ^ Q[20] /*7991*/;
assign _2370_ = _2126_ & _2373_ /*7987*/;
assign _2371_ = _2126_ ^ _2373_ /*7990*/;
assign _2372_ = _2364_ & _2371_ /*7988*/;
assign _2320_ = _2364_ ^ _2371_ /*7989*/;
assign _2369_ = _2370_ | _2372_ /*7986*/;
assign _2378_ = D[5] ^ Q[20] /*7985*/;
assign _2375_ = _2127_ & _2378_ /*7981*/;
assign _2376_ = _2127_ ^ _2378_ /*7984*/;
assign _2377_ = _2369_ & _2376_ /*7982*/;
assign _2321_ = _2369_ ^ _2376_ /*7983*/;
assign _2374_ = _2375_ | _2377_ /*7980*/;
assign _2383_ = D[6] ^ Q[20] /*7979*/;
assign _2380_ = _2128_ & _2383_ /*7975*/;
assign _2381_ = _2128_ ^ _2383_ /*7978*/;
assign _2382_ = _2374_ & _2381_ /*7976*/;
assign _2322_ = _2374_ ^ _2381_ /*7977*/;
assign _2379_ = _2380_ | _2382_ /*7974*/;
assign _2388_ = D[7] ^ Q[20] /*7973*/;
assign _2385_ = _2129_ & _2388_ /*7969*/;
assign _2386_ = _2129_ ^ _2388_ /*7972*/;
assign _2387_ = _2379_ & _2386_ /*7970*/;
assign _2323_ = _2379_ ^ _2386_ /*7971*/;
assign _2384_ = _2385_ | _2387_ /*7968*/;
assign _2393_ = D[8] ^ Q[20] /*7967*/;
assign _2390_ = _2130_ & _2393_ /*7963*/;
assign _2391_ = _2130_ ^ _2393_ /*7966*/;
assign _2392_ = _2384_ & _2391_ /*7964*/;
assign _2324_ = _2384_ ^ _2391_ /*7965*/;
assign _2389_ = _2390_ | _2392_ /*7962*/;
assign _2398_ = D[9] ^ Q[20] /*7961*/;
assign _2395_ = _2131_ & _2398_ /*7957*/;
assign _2396_ = _2131_ ^ _2398_ /*7960*/;
assign _2397_ = _2389_ & _2396_ /*7958*/;
assign _2325_ = _2389_ ^ _2396_ /*7959*/;
assign _2394_ = _2395_ | _2397_ /*7956*/;
assign _2403_ = D[10] ^ Q[20] /*7955*/;
assign _2400_ = _2132_ & _2403_ /*7951*/;
assign _2401_ = _2132_ ^ _2403_ /*7954*/;
assign _2402_ = _2394_ & _2401_ /*7952*/;
assign _2326_ = _2394_ ^ _2401_ /*7953*/;
assign _2399_ = _2400_ | _2402_ /*7950*/;
assign _2408_ = D[11] ^ Q[20] /*7949*/;
assign _2405_ = _2133_ & _2408_ /*7945*/;
assign _2406_ = _2133_ ^ _2408_ /*7948*/;
assign _2407_ = _2399_ & _2406_ /*7946*/;
assign _2327_ = _2399_ ^ _2406_ /*7947*/;
assign _2404_ = _2405_ | _2407_ /*7944*/;
assign _2413_ = D[12] ^ Q[20] /*7943*/;
assign _2410_ = _2134_ & _2413_ /*7939*/;
assign _2411_ = _2134_ ^ _2413_ /*7942*/;
assign _2412_ = _2404_ & _2411_ /*7940*/;
assign _2328_ = _2404_ ^ _2411_ /*7941*/;
assign _2409_ = _2410_ | _2412_ /*7938*/;
assign _2418_ = D[13] ^ Q[20] /*7937*/;
assign _2415_ = _2135_ & _2418_ /*7933*/;
assign _2416_ = _2135_ ^ _2418_ /*7936*/;
assign _2417_ = _2409_ & _2416_ /*7934*/;
assign _2329_ = _2409_ ^ _2416_ /*7935*/;
assign _2414_ = _2415_ | _2417_ /*7932*/;
assign _2423_ = D[14] ^ Q[20] /*7931*/;
assign _2420_ = _2136_ & _2423_ /*7927*/;
assign _2421_ = _2136_ ^ _2423_ /*7930*/;
assign _2422_ = _2414_ & _2421_ /*7928*/;
assign _2330_ = _2414_ ^ _2421_ /*7929*/;
assign _2419_ = _2420_ | _2422_ /*7926*/;
assign _2428_ = D[15] ^ Q[20] /*7925*/;
assign _2425_ = _2137_ & _2428_ /*7921*/;
assign _2426_ = _2137_ ^ _2428_ /*7924*/;
assign _2427_ = _2419_ & _2426_ /*7922*/;
assign _2331_ = _2419_ ^ _2426_ /*7923*/;
assign _2424_ = _2425_ | _2427_ /*7920*/;
assign _2433_ = D[16] ^ Q[20] /*7919*/;
assign _2430_ = _2138_ & _2433_ /*7915*/;
assign _2431_ = _2138_ ^ _2433_ /*7918*/;
assign _2432_ = _2424_ & _2431_ /*7916*/;
assign _2332_ = _2424_ ^ _2431_ /*7917*/;
assign _2429_ = _2430_ | _2432_ /*7914*/;
assign _2438_ = D[17] ^ Q[20] /*7913*/;
assign _2435_ = _2139_ & _2438_ /*7909*/;
assign _2436_ = _2139_ ^ _2438_ /*7912*/;
assign _2437_ = _2429_ & _2436_ /*7910*/;
assign _2333_ = _2429_ ^ _2436_ /*7911*/;
assign _2434_ = _2435_ | _2437_ /*7908*/;
assign _2443_ = D[18] ^ Q[20] /*7907*/;
assign _2440_ = _2140_ & _2443_ /*7903*/;
assign _2441_ = _2140_ ^ _2443_ /*7906*/;
assign _2442_ = _2434_ & _2441_ /*7904*/;
assign _2334_ = _2434_ ^ _2441_ /*7905*/;
assign _2439_ = _2440_ | _2442_ /*7902*/;
assign _2448_ = D[19] ^ Q[20] /*7901*/;
assign _2445_ = _2141_ & _2448_ /*7897*/;
assign _2446_ = _2141_ ^ _2448_ /*7900*/;
assign _2447_ = _2439_ & _2446_ /*7898*/;
assign _2335_ = _2439_ ^ _2446_ /*7899*/;
assign _2444_ = _2445_ | _2447_ /*7896*/;
assign _2453_ = D[20] ^ Q[20] /*7895*/;
assign _2450_ = _2142_ & _2453_ /*7891*/;
assign _2451_ = _2142_ ^ _2453_ /*7894*/;
assign _2452_ = _2444_ & _2451_ /*7892*/;
assign _2336_ = _2444_ ^ _2451_ /*7893*/;
assign _2449_ = _2450_ | _2452_ /*7890*/;
assign _2458_ = D[21] ^ Q[20] /*7889*/;
assign _2455_ = _2143_ & _2458_ /*7885*/;
assign _2456_ = _2143_ ^ _2458_ /*7888*/;
assign _2457_ = _2449_ & _2456_ /*7886*/;
assign _2337_ = _2449_ ^ _2456_ /*7887*/;
assign _2454_ = _2455_ | _2457_ /*7884*/;
assign _2463_ = D[22] ^ Q[20] /*7883*/;
assign _2460_ = _2144_ & _2463_ /*7879*/;
assign _2461_ = _2144_ ^ _2463_ /*7882*/;
assign _2462_ = _2454_ & _2461_ /*7880*/;
assign _2338_ = _2454_ ^ _2461_ /*7881*/;
assign _2459_ = _2460_ | _2462_ /*7878*/;
assign _2468_ = D[23] ^ Q[20] /*7877*/;
assign _2465_ = _2145_ & _2468_ /*7873*/;
assign _2466_ = _2145_ ^ _2468_ /*7876*/;
assign _2467_ = _2459_ & _2466_ /*7874*/;
assign _2339_ = _2459_ ^ _2466_ /*7875*/;
assign _2464_ = _2465_ | _2467_ /*7872*/;
assign _2473_ = D[24] ^ Q[20] /*7871*/;
assign _2470_ = _2146_ & _2473_ /*7867*/;
assign _2471_ = _2146_ ^ _2473_ /*7870*/;
assign _2472_ = _2464_ & _2471_ /*7868*/;
assign _2340_ = _2464_ ^ _2471_ /*7869*/;
assign _2469_ = _2470_ | _2472_ /*7866*/;
assign _2478_ = D[25] ^ Q[20] /*7865*/;
assign _2475_ = _2147_ & _2478_ /*7861*/;
assign _2476_ = _2147_ ^ _2478_ /*7864*/;
assign _2477_ = _2469_ & _2476_ /*7862*/;
assign _2341_ = _2469_ ^ _2476_ /*7863*/;
assign _2474_ = _2475_ | _2477_ /*7860*/;
assign _2483_ = D[26] ^ Q[20] /*7859*/;
assign _2480_ = _2148_ & _2483_ /*7855*/;
assign _2481_ = _2148_ ^ _2483_ /*7858*/;
assign _2482_ = _2474_ & _2481_ /*7856*/;
assign _2342_ = _2474_ ^ _2481_ /*7857*/;
assign _2479_ = _2480_ | _2482_ /*7854*/;
assign _2488_ = D[27] ^ Q[20] /*7853*/;
assign _2485_ = _2149_ & _2488_ /*7849*/;
assign _2486_ = _2149_ ^ _2488_ /*7852*/;
assign _2487_ = _2479_ & _2486_ /*7850*/;
assign _2343_ = _2479_ ^ _2486_ /*7851*/;
assign _2484_ = _2485_ | _2487_ /*7848*/;
assign _2493_ = D[28] ^ Q[20] /*7847*/;
assign _2490_ = _2150_ & _2493_ /*7843*/;
assign _2491_ = _2150_ ^ _2493_ /*7846*/;
assign _2492_ = _2484_ & _2491_ /*7844*/;
assign _2344_ = _2484_ ^ _2491_ /*7845*/;
assign _2489_ = _2490_ | _2492_ /*7842*/;
assign _2498_ = D[29] ^ Q[20] /*7841*/;
assign _2495_ = _2151_ & _2498_ /*7837*/;
assign _2496_ = _2151_ ^ _2498_ /*7840*/;
assign _2497_ = _2489_ & _2496_ /*7838*/;
assign _2345_ = _2489_ ^ _2496_ /*7839*/;
assign _2494_ = _2495_ | _2497_ /*7836*/;
assign _2503_ = D[30] ^ Q[20] /*7835*/;
assign _2500_ = _2152_ & _2503_ /*7831*/;
assign _2501_ = _2152_ ^ _2503_ /*7834*/;
assign _2502_ = _2494_ & _2501_ /*7832*/;
assign _2346_ = _2494_ ^ _2501_ /*7833*/;
assign _2499_ = _2500_ | _2502_ /*7830*/;
assign _2507_ = zeroWire ^ Q[20] /*7829*/;
assign _2504_ = _2153_ & _2507_ /*7825*/;
assign _2505_ = _2153_ ^ _2507_ /*7828*/;
assign _2506_ = _2499_ & _2505_ /*7826*/;
assign _2347_ = _2499_ ^ _2505_ /*7827*/;
assign Q[19] = _2504_ | _2506_ /*7824*/;
assign _2546_ = D[0] ^ Q[19] /*7630*/;
assign _2543_ = R_0[18] & _2546_ /*7626*/;
assign _2544_ = R_0[18] ^ _2546_ /*7629*/;
assign _2545_ = Q[19] & _2544_ /*7627*/;
assign _2509_ = Q[19] ^ _2544_ /*7628*/;
assign _2542_ = _2543_ | _2545_ /*7625*/;
assign _2551_ = D[1] ^ Q[19] /*7624*/;
assign _2548_ = _2316_ & _2551_ /*7620*/;
assign _2549_ = _2316_ ^ _2551_ /*7623*/;
assign _2550_ = _2542_ & _2549_ /*7621*/;
assign _2510_ = _2542_ ^ _2549_ /*7622*/;
assign _2547_ = _2548_ | _2550_ /*7619*/;
assign _2556_ = D[2] ^ Q[19] /*7618*/;
assign _2553_ = _2317_ & _2556_ /*7614*/;
assign _2554_ = _2317_ ^ _2556_ /*7617*/;
assign _2555_ = _2547_ & _2554_ /*7615*/;
assign _2511_ = _2547_ ^ _2554_ /*7616*/;
assign _2552_ = _2553_ | _2555_ /*7613*/;
assign _2561_ = D[3] ^ Q[19] /*7612*/;
assign _2558_ = _2318_ & _2561_ /*7608*/;
assign _2559_ = _2318_ ^ _2561_ /*7611*/;
assign _2560_ = _2552_ & _2559_ /*7609*/;
assign _2512_ = _2552_ ^ _2559_ /*7610*/;
assign _2557_ = _2558_ | _2560_ /*7607*/;
assign _2566_ = D[4] ^ Q[19] /*7606*/;
assign _2563_ = _2319_ & _2566_ /*7602*/;
assign _2564_ = _2319_ ^ _2566_ /*7605*/;
assign _2565_ = _2557_ & _2564_ /*7603*/;
assign _2513_ = _2557_ ^ _2564_ /*7604*/;
assign _2562_ = _2563_ | _2565_ /*7601*/;
assign _2571_ = D[5] ^ Q[19] /*7600*/;
assign _2568_ = _2320_ & _2571_ /*7596*/;
assign _2569_ = _2320_ ^ _2571_ /*7599*/;
assign _2570_ = _2562_ & _2569_ /*7597*/;
assign _2514_ = _2562_ ^ _2569_ /*7598*/;
assign _2567_ = _2568_ | _2570_ /*7595*/;
assign _2576_ = D[6] ^ Q[19] /*7594*/;
assign _2573_ = _2321_ & _2576_ /*7590*/;
assign _2574_ = _2321_ ^ _2576_ /*7593*/;
assign _2575_ = _2567_ & _2574_ /*7591*/;
assign _2515_ = _2567_ ^ _2574_ /*7592*/;
assign _2572_ = _2573_ | _2575_ /*7589*/;
assign _2581_ = D[7] ^ Q[19] /*7588*/;
assign _2578_ = _2322_ & _2581_ /*7584*/;
assign _2579_ = _2322_ ^ _2581_ /*7587*/;
assign _2580_ = _2572_ & _2579_ /*7585*/;
assign _2516_ = _2572_ ^ _2579_ /*7586*/;
assign _2577_ = _2578_ | _2580_ /*7583*/;
assign _2586_ = D[8] ^ Q[19] /*7582*/;
assign _2583_ = _2323_ & _2586_ /*7578*/;
assign _2584_ = _2323_ ^ _2586_ /*7581*/;
assign _2585_ = _2577_ & _2584_ /*7579*/;
assign _2517_ = _2577_ ^ _2584_ /*7580*/;
assign _2582_ = _2583_ | _2585_ /*7577*/;
assign _2591_ = D[9] ^ Q[19] /*7576*/;
assign _2588_ = _2324_ & _2591_ /*7572*/;
assign _2589_ = _2324_ ^ _2591_ /*7575*/;
assign _2590_ = _2582_ & _2589_ /*7573*/;
assign _2518_ = _2582_ ^ _2589_ /*7574*/;
assign _2587_ = _2588_ | _2590_ /*7571*/;
assign _2596_ = D[10] ^ Q[19] /*7570*/;
assign _2593_ = _2325_ & _2596_ /*7566*/;
assign _2594_ = _2325_ ^ _2596_ /*7569*/;
assign _2595_ = _2587_ & _2594_ /*7567*/;
assign _2519_ = _2587_ ^ _2594_ /*7568*/;
assign _2592_ = _2593_ | _2595_ /*7565*/;
assign _2601_ = D[11] ^ Q[19] /*7564*/;
assign _2598_ = _2326_ & _2601_ /*7560*/;
assign _2599_ = _2326_ ^ _2601_ /*7563*/;
assign _2600_ = _2592_ & _2599_ /*7561*/;
assign _2520_ = _2592_ ^ _2599_ /*7562*/;
assign _2597_ = _2598_ | _2600_ /*7559*/;
assign _2606_ = D[12] ^ Q[19] /*7558*/;
assign _2603_ = _2327_ & _2606_ /*7554*/;
assign _2604_ = _2327_ ^ _2606_ /*7557*/;
assign _2605_ = _2597_ & _2604_ /*7555*/;
assign _2521_ = _2597_ ^ _2604_ /*7556*/;
assign _2602_ = _2603_ | _2605_ /*7553*/;
assign _2611_ = D[13] ^ Q[19] /*7552*/;
assign _2608_ = _2328_ & _2611_ /*7548*/;
assign _2609_ = _2328_ ^ _2611_ /*7551*/;
assign _2610_ = _2602_ & _2609_ /*7549*/;
assign _2522_ = _2602_ ^ _2609_ /*7550*/;
assign _2607_ = _2608_ | _2610_ /*7547*/;
assign _2616_ = D[14] ^ Q[19] /*7546*/;
assign _2613_ = _2329_ & _2616_ /*7542*/;
assign _2614_ = _2329_ ^ _2616_ /*7545*/;
assign _2615_ = _2607_ & _2614_ /*7543*/;
assign _2523_ = _2607_ ^ _2614_ /*7544*/;
assign _2612_ = _2613_ | _2615_ /*7541*/;
assign _2621_ = D[15] ^ Q[19] /*7540*/;
assign _2618_ = _2330_ & _2621_ /*7536*/;
assign _2619_ = _2330_ ^ _2621_ /*7539*/;
assign _2620_ = _2612_ & _2619_ /*7537*/;
assign _2524_ = _2612_ ^ _2619_ /*7538*/;
assign _2617_ = _2618_ | _2620_ /*7535*/;
assign _2626_ = D[16] ^ Q[19] /*7534*/;
assign _2623_ = _2331_ & _2626_ /*7530*/;
assign _2624_ = _2331_ ^ _2626_ /*7533*/;
assign _2625_ = _2617_ & _2624_ /*7531*/;
assign _2525_ = _2617_ ^ _2624_ /*7532*/;
assign _2622_ = _2623_ | _2625_ /*7529*/;
assign _2631_ = D[17] ^ Q[19] /*7528*/;
assign _2628_ = _2332_ & _2631_ /*7524*/;
assign _2629_ = _2332_ ^ _2631_ /*7527*/;
assign _2630_ = _2622_ & _2629_ /*7525*/;
assign _2526_ = _2622_ ^ _2629_ /*7526*/;
assign _2627_ = _2628_ | _2630_ /*7523*/;
assign _2636_ = D[18] ^ Q[19] /*7522*/;
assign _2633_ = _2333_ & _2636_ /*7518*/;
assign _2634_ = _2333_ ^ _2636_ /*7521*/;
assign _2635_ = _2627_ & _2634_ /*7519*/;
assign _2527_ = _2627_ ^ _2634_ /*7520*/;
assign _2632_ = _2633_ | _2635_ /*7517*/;
assign _2641_ = D[19] ^ Q[19] /*7516*/;
assign _2638_ = _2334_ & _2641_ /*7512*/;
assign _2639_ = _2334_ ^ _2641_ /*7515*/;
assign _2640_ = _2632_ & _2639_ /*7513*/;
assign _2528_ = _2632_ ^ _2639_ /*7514*/;
assign _2637_ = _2638_ | _2640_ /*7511*/;
assign _2646_ = D[20] ^ Q[19] /*7510*/;
assign _2643_ = _2335_ & _2646_ /*7506*/;
assign _2644_ = _2335_ ^ _2646_ /*7509*/;
assign _2645_ = _2637_ & _2644_ /*7507*/;
assign _2529_ = _2637_ ^ _2644_ /*7508*/;
assign _2642_ = _2643_ | _2645_ /*7505*/;
assign _2651_ = D[21] ^ Q[19] /*7504*/;
assign _2648_ = _2336_ & _2651_ /*7500*/;
assign _2649_ = _2336_ ^ _2651_ /*7503*/;
assign _2650_ = _2642_ & _2649_ /*7501*/;
assign _2530_ = _2642_ ^ _2649_ /*7502*/;
assign _2647_ = _2648_ | _2650_ /*7499*/;
assign _2656_ = D[22] ^ Q[19] /*7498*/;
assign _2653_ = _2337_ & _2656_ /*7494*/;
assign _2654_ = _2337_ ^ _2656_ /*7497*/;
assign _2655_ = _2647_ & _2654_ /*7495*/;
assign _2531_ = _2647_ ^ _2654_ /*7496*/;
assign _2652_ = _2653_ | _2655_ /*7493*/;
assign _2661_ = D[23] ^ Q[19] /*7492*/;
assign _2658_ = _2338_ & _2661_ /*7488*/;
assign _2659_ = _2338_ ^ _2661_ /*7491*/;
assign _2660_ = _2652_ & _2659_ /*7489*/;
assign _2532_ = _2652_ ^ _2659_ /*7490*/;
assign _2657_ = _2658_ | _2660_ /*7487*/;
assign _2666_ = D[24] ^ Q[19] /*7486*/;
assign _2663_ = _2339_ & _2666_ /*7482*/;
assign _2664_ = _2339_ ^ _2666_ /*7485*/;
assign _2665_ = _2657_ & _2664_ /*7483*/;
assign _2533_ = _2657_ ^ _2664_ /*7484*/;
assign _2662_ = _2663_ | _2665_ /*7481*/;
assign _2671_ = D[25] ^ Q[19] /*7480*/;
assign _2668_ = _2340_ & _2671_ /*7476*/;
assign _2669_ = _2340_ ^ _2671_ /*7479*/;
assign _2670_ = _2662_ & _2669_ /*7477*/;
assign _2534_ = _2662_ ^ _2669_ /*7478*/;
assign _2667_ = _2668_ | _2670_ /*7475*/;
assign _2676_ = D[26] ^ Q[19] /*7474*/;
assign _2673_ = _2341_ & _2676_ /*7470*/;
assign _2674_ = _2341_ ^ _2676_ /*7473*/;
assign _2675_ = _2667_ & _2674_ /*7471*/;
assign _2535_ = _2667_ ^ _2674_ /*7472*/;
assign _2672_ = _2673_ | _2675_ /*7469*/;
assign _2681_ = D[27] ^ Q[19] /*7468*/;
assign _2678_ = _2342_ & _2681_ /*7464*/;
assign _2679_ = _2342_ ^ _2681_ /*7467*/;
assign _2680_ = _2672_ & _2679_ /*7465*/;
assign _2536_ = _2672_ ^ _2679_ /*7466*/;
assign _2677_ = _2678_ | _2680_ /*7463*/;
assign _2686_ = D[28] ^ Q[19] /*7462*/;
assign _2683_ = _2343_ & _2686_ /*7458*/;
assign _2684_ = _2343_ ^ _2686_ /*7461*/;
assign _2685_ = _2677_ & _2684_ /*7459*/;
assign _2537_ = _2677_ ^ _2684_ /*7460*/;
assign _2682_ = _2683_ | _2685_ /*7457*/;
assign _2691_ = D[29] ^ Q[19] /*7456*/;
assign _2688_ = _2344_ & _2691_ /*7452*/;
assign _2689_ = _2344_ ^ _2691_ /*7455*/;
assign _2690_ = _2682_ & _2689_ /*7453*/;
assign _2538_ = _2682_ ^ _2689_ /*7454*/;
assign _2687_ = _2688_ | _2690_ /*7451*/;
assign _2696_ = D[30] ^ Q[19] /*7450*/;
assign _2693_ = _2345_ & _2696_ /*7446*/;
assign _2694_ = _2345_ ^ _2696_ /*7449*/;
assign _2695_ = _2687_ & _2694_ /*7447*/;
assign _2539_ = _2687_ ^ _2694_ /*7448*/;
assign _2692_ = _2693_ | _2695_ /*7445*/;
assign _2700_ = zeroWire ^ Q[19] /*7444*/;
assign _2697_ = _2346_ & _2700_ /*7440*/;
assign _2698_ = _2346_ ^ _2700_ /*7443*/;
assign _2699_ = _2692_ & _2698_ /*7441*/;
assign _2540_ = _2692_ ^ _2698_ /*7442*/;
assign Q[18] = _2697_ | _2699_ /*7439*/;
assign _2739_ = D[0] ^ Q[18] /*7245*/;
assign _2736_ = R_0[17] & _2739_ /*7241*/;
assign _2737_ = R_0[17] ^ _2739_ /*7244*/;
assign _2738_ = Q[18] & _2737_ /*7242*/;
assign _2702_ = Q[18] ^ _2737_ /*7243*/;
assign _2735_ = _2736_ | _2738_ /*7240*/;
assign _2744_ = D[1] ^ Q[18] /*7239*/;
assign _2741_ = _2509_ & _2744_ /*7235*/;
assign _2742_ = _2509_ ^ _2744_ /*7238*/;
assign _2743_ = _2735_ & _2742_ /*7236*/;
assign _2703_ = _2735_ ^ _2742_ /*7237*/;
assign _2740_ = _2741_ | _2743_ /*7234*/;
assign _2749_ = D[2] ^ Q[18] /*7233*/;
assign _2746_ = _2510_ & _2749_ /*7229*/;
assign _2747_ = _2510_ ^ _2749_ /*7232*/;
assign _2748_ = _2740_ & _2747_ /*7230*/;
assign _2704_ = _2740_ ^ _2747_ /*7231*/;
assign _2745_ = _2746_ | _2748_ /*7228*/;
assign _2754_ = D[3] ^ Q[18] /*7227*/;
assign _2751_ = _2511_ & _2754_ /*7223*/;
assign _2752_ = _2511_ ^ _2754_ /*7226*/;
assign _2753_ = _2745_ & _2752_ /*7224*/;
assign _2705_ = _2745_ ^ _2752_ /*7225*/;
assign _2750_ = _2751_ | _2753_ /*7222*/;
assign _2759_ = D[4] ^ Q[18] /*7221*/;
assign _2756_ = _2512_ & _2759_ /*7217*/;
assign _2757_ = _2512_ ^ _2759_ /*7220*/;
assign _2758_ = _2750_ & _2757_ /*7218*/;
assign _2706_ = _2750_ ^ _2757_ /*7219*/;
assign _2755_ = _2756_ | _2758_ /*7216*/;
assign _2764_ = D[5] ^ Q[18] /*7215*/;
assign _2761_ = _2513_ & _2764_ /*7211*/;
assign _2762_ = _2513_ ^ _2764_ /*7214*/;
assign _2763_ = _2755_ & _2762_ /*7212*/;
assign _2707_ = _2755_ ^ _2762_ /*7213*/;
assign _2760_ = _2761_ | _2763_ /*7210*/;
assign _2769_ = D[6] ^ Q[18] /*7209*/;
assign _2766_ = _2514_ & _2769_ /*7205*/;
assign _2767_ = _2514_ ^ _2769_ /*7208*/;
assign _2768_ = _2760_ & _2767_ /*7206*/;
assign _2708_ = _2760_ ^ _2767_ /*7207*/;
assign _2765_ = _2766_ | _2768_ /*7204*/;
assign _2774_ = D[7] ^ Q[18] /*7203*/;
assign _2771_ = _2515_ & _2774_ /*7199*/;
assign _2772_ = _2515_ ^ _2774_ /*7202*/;
assign _2773_ = _2765_ & _2772_ /*7200*/;
assign _2709_ = _2765_ ^ _2772_ /*7201*/;
assign _2770_ = _2771_ | _2773_ /*7198*/;
assign _2779_ = D[8] ^ Q[18] /*7197*/;
assign _2776_ = _2516_ & _2779_ /*7193*/;
assign _2777_ = _2516_ ^ _2779_ /*7196*/;
assign _2778_ = _2770_ & _2777_ /*7194*/;
assign _2710_ = _2770_ ^ _2777_ /*7195*/;
assign _2775_ = _2776_ | _2778_ /*7192*/;
assign _2784_ = D[9] ^ Q[18] /*7191*/;
assign _2781_ = _2517_ & _2784_ /*7187*/;
assign _2782_ = _2517_ ^ _2784_ /*7190*/;
assign _2783_ = _2775_ & _2782_ /*7188*/;
assign _2711_ = _2775_ ^ _2782_ /*7189*/;
assign _2780_ = _2781_ | _2783_ /*7186*/;
assign _2789_ = D[10] ^ Q[18] /*7185*/;
assign _2786_ = _2518_ & _2789_ /*7181*/;
assign _2787_ = _2518_ ^ _2789_ /*7184*/;
assign _2788_ = _2780_ & _2787_ /*7182*/;
assign _2712_ = _2780_ ^ _2787_ /*7183*/;
assign _2785_ = _2786_ | _2788_ /*7180*/;
assign _2794_ = D[11] ^ Q[18] /*7179*/;
assign _2791_ = _2519_ & _2794_ /*7175*/;
assign _2792_ = _2519_ ^ _2794_ /*7178*/;
assign _2793_ = _2785_ & _2792_ /*7176*/;
assign _2713_ = _2785_ ^ _2792_ /*7177*/;
assign _2790_ = _2791_ | _2793_ /*7174*/;
assign _2799_ = D[12] ^ Q[18] /*7173*/;
assign _2796_ = _2520_ & _2799_ /*7169*/;
assign _2797_ = _2520_ ^ _2799_ /*7172*/;
assign _2798_ = _2790_ & _2797_ /*7170*/;
assign _2714_ = _2790_ ^ _2797_ /*7171*/;
assign _2795_ = _2796_ | _2798_ /*7168*/;
assign _2804_ = D[13] ^ Q[18] /*7167*/;
assign _2801_ = _2521_ & _2804_ /*7163*/;
assign _2802_ = _2521_ ^ _2804_ /*7166*/;
assign _2803_ = _2795_ & _2802_ /*7164*/;
assign _2715_ = _2795_ ^ _2802_ /*7165*/;
assign _2800_ = _2801_ | _2803_ /*7162*/;
assign _2809_ = D[14] ^ Q[18] /*7161*/;
assign _2806_ = _2522_ & _2809_ /*7157*/;
assign _2807_ = _2522_ ^ _2809_ /*7160*/;
assign _2808_ = _2800_ & _2807_ /*7158*/;
assign _2716_ = _2800_ ^ _2807_ /*7159*/;
assign _2805_ = _2806_ | _2808_ /*7156*/;
assign _2814_ = D[15] ^ Q[18] /*7155*/;
assign _2811_ = _2523_ & _2814_ /*7151*/;
assign _2812_ = _2523_ ^ _2814_ /*7154*/;
assign _2813_ = _2805_ & _2812_ /*7152*/;
assign _2717_ = _2805_ ^ _2812_ /*7153*/;
assign _2810_ = _2811_ | _2813_ /*7150*/;
assign _2819_ = D[16] ^ Q[18] /*7149*/;
assign _2816_ = _2524_ & _2819_ /*7145*/;
assign _2817_ = _2524_ ^ _2819_ /*7148*/;
assign _2818_ = _2810_ & _2817_ /*7146*/;
assign _2718_ = _2810_ ^ _2817_ /*7147*/;
assign _2815_ = _2816_ | _2818_ /*7144*/;
assign _2824_ = D[17] ^ Q[18] /*7143*/;
assign _2821_ = _2525_ & _2824_ /*7139*/;
assign _2822_ = _2525_ ^ _2824_ /*7142*/;
assign _2823_ = _2815_ & _2822_ /*7140*/;
assign _2719_ = _2815_ ^ _2822_ /*7141*/;
assign _2820_ = _2821_ | _2823_ /*7138*/;
assign _2829_ = D[18] ^ Q[18] /*7137*/;
assign _2826_ = _2526_ & _2829_ /*7133*/;
assign _2827_ = _2526_ ^ _2829_ /*7136*/;
assign _2828_ = _2820_ & _2827_ /*7134*/;
assign _2720_ = _2820_ ^ _2827_ /*7135*/;
assign _2825_ = _2826_ | _2828_ /*7132*/;
assign _2834_ = D[19] ^ Q[18] /*7131*/;
assign _2831_ = _2527_ & _2834_ /*7127*/;
assign _2832_ = _2527_ ^ _2834_ /*7130*/;
assign _2833_ = _2825_ & _2832_ /*7128*/;
assign _2721_ = _2825_ ^ _2832_ /*7129*/;
assign _2830_ = _2831_ | _2833_ /*7126*/;
assign _2839_ = D[20] ^ Q[18] /*7125*/;
assign _2836_ = _2528_ & _2839_ /*7121*/;
assign _2837_ = _2528_ ^ _2839_ /*7124*/;
assign _2838_ = _2830_ & _2837_ /*7122*/;
assign _2722_ = _2830_ ^ _2837_ /*7123*/;
assign _2835_ = _2836_ | _2838_ /*7120*/;
assign _2844_ = D[21] ^ Q[18] /*7119*/;
assign _2841_ = _2529_ & _2844_ /*7115*/;
assign _2842_ = _2529_ ^ _2844_ /*7118*/;
assign _2843_ = _2835_ & _2842_ /*7116*/;
assign _2723_ = _2835_ ^ _2842_ /*7117*/;
assign _2840_ = _2841_ | _2843_ /*7114*/;
assign _2849_ = D[22] ^ Q[18] /*7113*/;
assign _2846_ = _2530_ & _2849_ /*7109*/;
assign _2847_ = _2530_ ^ _2849_ /*7112*/;
assign _2848_ = _2840_ & _2847_ /*7110*/;
assign _2724_ = _2840_ ^ _2847_ /*7111*/;
assign _2845_ = _2846_ | _2848_ /*7108*/;
assign _2854_ = D[23] ^ Q[18] /*7107*/;
assign _2851_ = _2531_ & _2854_ /*7103*/;
assign _2852_ = _2531_ ^ _2854_ /*7106*/;
assign _2853_ = _2845_ & _2852_ /*7104*/;
assign _2725_ = _2845_ ^ _2852_ /*7105*/;
assign _2850_ = _2851_ | _2853_ /*7102*/;
assign _2859_ = D[24] ^ Q[18] /*7101*/;
assign _2856_ = _2532_ & _2859_ /*7097*/;
assign _2857_ = _2532_ ^ _2859_ /*7100*/;
assign _2858_ = _2850_ & _2857_ /*7098*/;
assign _2726_ = _2850_ ^ _2857_ /*7099*/;
assign _2855_ = _2856_ | _2858_ /*7096*/;
assign _2864_ = D[25] ^ Q[18] /*7095*/;
assign _2861_ = _2533_ & _2864_ /*7091*/;
assign _2862_ = _2533_ ^ _2864_ /*7094*/;
assign _2863_ = _2855_ & _2862_ /*7092*/;
assign _2727_ = _2855_ ^ _2862_ /*7093*/;
assign _2860_ = _2861_ | _2863_ /*7090*/;
assign _2869_ = D[26] ^ Q[18] /*7089*/;
assign _2866_ = _2534_ & _2869_ /*7085*/;
assign _2867_ = _2534_ ^ _2869_ /*7088*/;
assign _2868_ = _2860_ & _2867_ /*7086*/;
assign _2728_ = _2860_ ^ _2867_ /*7087*/;
assign _2865_ = _2866_ | _2868_ /*7084*/;
assign _2874_ = D[27] ^ Q[18] /*7083*/;
assign _2871_ = _2535_ & _2874_ /*7079*/;
assign _2872_ = _2535_ ^ _2874_ /*7082*/;
assign _2873_ = _2865_ & _2872_ /*7080*/;
assign _2729_ = _2865_ ^ _2872_ /*7081*/;
assign _2870_ = _2871_ | _2873_ /*7078*/;
assign _2879_ = D[28] ^ Q[18] /*7077*/;
assign _2876_ = _2536_ & _2879_ /*7073*/;
assign _2877_ = _2536_ ^ _2879_ /*7076*/;
assign _2878_ = _2870_ & _2877_ /*7074*/;
assign _2730_ = _2870_ ^ _2877_ /*7075*/;
assign _2875_ = _2876_ | _2878_ /*7072*/;
assign _2884_ = D[29] ^ Q[18] /*7071*/;
assign _2881_ = _2537_ & _2884_ /*7067*/;
assign _2882_ = _2537_ ^ _2884_ /*7070*/;
assign _2883_ = _2875_ & _2882_ /*7068*/;
assign _2731_ = _2875_ ^ _2882_ /*7069*/;
assign _2880_ = _2881_ | _2883_ /*7066*/;
assign _2889_ = D[30] ^ Q[18] /*7065*/;
assign _2886_ = _2538_ & _2889_ /*7061*/;
assign _2887_ = _2538_ ^ _2889_ /*7064*/;
assign _2888_ = _2880_ & _2887_ /*7062*/;
assign _2732_ = _2880_ ^ _2887_ /*7063*/;
assign _2885_ = _2886_ | _2888_ /*7060*/;
assign _2893_ = zeroWire ^ Q[18] /*7059*/;
assign _2890_ = _2539_ & _2893_ /*7055*/;
assign _2891_ = _2539_ ^ _2893_ /*7058*/;
assign _2892_ = _2885_ & _2891_ /*7056*/;
assign _2733_ = _2885_ ^ _2891_ /*7057*/;
assign Q[17] = _2890_ | _2892_ /*7054*/;
assign _2932_ = D[0] ^ Q[17] /*6860*/;
assign _2929_ = R_0[16] & _2932_ /*6856*/;
assign _2930_ = R_0[16] ^ _2932_ /*6859*/;
assign _2931_ = Q[17] & _2930_ /*6857*/;
assign _2895_ = Q[17] ^ _2930_ /*6858*/;
assign _2928_ = _2929_ | _2931_ /*6855*/;
assign _2937_ = D[1] ^ Q[17] /*6854*/;
assign _2934_ = _2702_ & _2937_ /*6850*/;
assign _2935_ = _2702_ ^ _2937_ /*6853*/;
assign _2936_ = _2928_ & _2935_ /*6851*/;
assign _2896_ = _2928_ ^ _2935_ /*6852*/;
assign _2933_ = _2934_ | _2936_ /*6849*/;
assign _2942_ = D[2] ^ Q[17] /*6848*/;
assign _2939_ = _2703_ & _2942_ /*6844*/;
assign _2940_ = _2703_ ^ _2942_ /*6847*/;
assign _2941_ = _2933_ & _2940_ /*6845*/;
assign _2897_ = _2933_ ^ _2940_ /*6846*/;
assign _2938_ = _2939_ | _2941_ /*6843*/;
assign _2947_ = D[3] ^ Q[17] /*6842*/;
assign _2944_ = _2704_ & _2947_ /*6838*/;
assign _2945_ = _2704_ ^ _2947_ /*6841*/;
assign _2946_ = _2938_ & _2945_ /*6839*/;
assign _2898_ = _2938_ ^ _2945_ /*6840*/;
assign _2943_ = _2944_ | _2946_ /*6837*/;
assign _2952_ = D[4] ^ Q[17] /*6836*/;
assign _2949_ = _2705_ & _2952_ /*6832*/;
assign _2950_ = _2705_ ^ _2952_ /*6835*/;
assign _2951_ = _2943_ & _2950_ /*6833*/;
assign _2899_ = _2943_ ^ _2950_ /*6834*/;
assign _2948_ = _2949_ | _2951_ /*6831*/;
assign _2957_ = D[5] ^ Q[17] /*6830*/;
assign _2954_ = _2706_ & _2957_ /*6826*/;
assign _2955_ = _2706_ ^ _2957_ /*6829*/;
assign _2956_ = _2948_ & _2955_ /*6827*/;
assign _2900_ = _2948_ ^ _2955_ /*6828*/;
assign _2953_ = _2954_ | _2956_ /*6825*/;
assign _2962_ = D[6] ^ Q[17] /*6824*/;
assign _2959_ = _2707_ & _2962_ /*6820*/;
assign _2960_ = _2707_ ^ _2962_ /*6823*/;
assign _2961_ = _2953_ & _2960_ /*6821*/;
assign _2901_ = _2953_ ^ _2960_ /*6822*/;
assign _2958_ = _2959_ | _2961_ /*6819*/;
assign _2967_ = D[7] ^ Q[17] /*6818*/;
assign _2964_ = _2708_ & _2967_ /*6814*/;
assign _2965_ = _2708_ ^ _2967_ /*6817*/;
assign _2966_ = _2958_ & _2965_ /*6815*/;
assign _2902_ = _2958_ ^ _2965_ /*6816*/;
assign _2963_ = _2964_ | _2966_ /*6813*/;
assign _2972_ = D[8] ^ Q[17] /*6812*/;
assign _2969_ = _2709_ & _2972_ /*6808*/;
assign _2970_ = _2709_ ^ _2972_ /*6811*/;
assign _2971_ = _2963_ & _2970_ /*6809*/;
assign _2903_ = _2963_ ^ _2970_ /*6810*/;
assign _2968_ = _2969_ | _2971_ /*6807*/;
assign _2977_ = D[9] ^ Q[17] /*6806*/;
assign _2974_ = _2710_ & _2977_ /*6802*/;
assign _2975_ = _2710_ ^ _2977_ /*6805*/;
assign _2976_ = _2968_ & _2975_ /*6803*/;
assign _2904_ = _2968_ ^ _2975_ /*6804*/;
assign _2973_ = _2974_ | _2976_ /*6801*/;
assign _2982_ = D[10] ^ Q[17] /*6800*/;
assign _2979_ = _2711_ & _2982_ /*6796*/;
assign _2980_ = _2711_ ^ _2982_ /*6799*/;
assign _2981_ = _2973_ & _2980_ /*6797*/;
assign _2905_ = _2973_ ^ _2980_ /*6798*/;
assign _2978_ = _2979_ | _2981_ /*6795*/;
assign _2987_ = D[11] ^ Q[17] /*6794*/;
assign _2984_ = _2712_ & _2987_ /*6790*/;
assign _2985_ = _2712_ ^ _2987_ /*6793*/;
assign _2986_ = _2978_ & _2985_ /*6791*/;
assign _2906_ = _2978_ ^ _2985_ /*6792*/;
assign _2983_ = _2984_ | _2986_ /*6789*/;
assign _2992_ = D[12] ^ Q[17] /*6788*/;
assign _2989_ = _2713_ & _2992_ /*6784*/;
assign _2990_ = _2713_ ^ _2992_ /*6787*/;
assign _2991_ = _2983_ & _2990_ /*6785*/;
assign _2907_ = _2983_ ^ _2990_ /*6786*/;
assign _2988_ = _2989_ | _2991_ /*6783*/;
assign _2997_ = D[13] ^ Q[17] /*6782*/;
assign _2994_ = _2714_ & _2997_ /*6778*/;
assign _2995_ = _2714_ ^ _2997_ /*6781*/;
assign _2996_ = _2988_ & _2995_ /*6779*/;
assign _2908_ = _2988_ ^ _2995_ /*6780*/;
assign _2993_ = _2994_ | _2996_ /*6777*/;
assign _3002_ = D[14] ^ Q[17] /*6776*/;
assign _2999_ = _2715_ & _3002_ /*6772*/;
assign _3000_ = _2715_ ^ _3002_ /*6775*/;
assign _3001_ = _2993_ & _3000_ /*6773*/;
assign _2909_ = _2993_ ^ _3000_ /*6774*/;
assign _2998_ = _2999_ | _3001_ /*6771*/;
assign _3007_ = D[15] ^ Q[17] /*6770*/;
assign _3004_ = _2716_ & _3007_ /*6766*/;
assign _3005_ = _2716_ ^ _3007_ /*6769*/;
assign _3006_ = _2998_ & _3005_ /*6767*/;
assign _2910_ = _2998_ ^ _3005_ /*6768*/;
assign _3003_ = _3004_ | _3006_ /*6765*/;
assign _3012_ = D[16] ^ Q[17] /*6764*/;
assign _3009_ = _2717_ & _3012_ /*6760*/;
assign _3010_ = _2717_ ^ _3012_ /*6763*/;
assign _3011_ = _3003_ & _3010_ /*6761*/;
assign _2911_ = _3003_ ^ _3010_ /*6762*/;
assign _3008_ = _3009_ | _3011_ /*6759*/;
assign _3017_ = D[17] ^ Q[17] /*6758*/;
assign _3014_ = _2718_ & _3017_ /*6754*/;
assign _3015_ = _2718_ ^ _3017_ /*6757*/;
assign _3016_ = _3008_ & _3015_ /*6755*/;
assign _2912_ = _3008_ ^ _3015_ /*6756*/;
assign _3013_ = _3014_ | _3016_ /*6753*/;
assign _3022_ = D[18] ^ Q[17] /*6752*/;
assign _3019_ = _2719_ & _3022_ /*6748*/;
assign _3020_ = _2719_ ^ _3022_ /*6751*/;
assign _3021_ = _3013_ & _3020_ /*6749*/;
assign _2913_ = _3013_ ^ _3020_ /*6750*/;
assign _3018_ = _3019_ | _3021_ /*6747*/;
assign _3027_ = D[19] ^ Q[17] /*6746*/;
assign _3024_ = _2720_ & _3027_ /*6742*/;
assign _3025_ = _2720_ ^ _3027_ /*6745*/;
assign _3026_ = _3018_ & _3025_ /*6743*/;
assign _2914_ = _3018_ ^ _3025_ /*6744*/;
assign _3023_ = _3024_ | _3026_ /*6741*/;
assign _3032_ = D[20] ^ Q[17] /*6740*/;
assign _3029_ = _2721_ & _3032_ /*6736*/;
assign _3030_ = _2721_ ^ _3032_ /*6739*/;
assign _3031_ = _3023_ & _3030_ /*6737*/;
assign _2915_ = _3023_ ^ _3030_ /*6738*/;
assign _3028_ = _3029_ | _3031_ /*6735*/;
assign _3037_ = D[21] ^ Q[17] /*6734*/;
assign _3034_ = _2722_ & _3037_ /*6730*/;
assign _3035_ = _2722_ ^ _3037_ /*6733*/;
assign _3036_ = _3028_ & _3035_ /*6731*/;
assign _2916_ = _3028_ ^ _3035_ /*6732*/;
assign _3033_ = _3034_ | _3036_ /*6729*/;
assign _3042_ = D[22] ^ Q[17] /*6728*/;
assign _3039_ = _2723_ & _3042_ /*6724*/;
assign _3040_ = _2723_ ^ _3042_ /*6727*/;
assign _3041_ = _3033_ & _3040_ /*6725*/;
assign _2917_ = _3033_ ^ _3040_ /*6726*/;
assign _3038_ = _3039_ | _3041_ /*6723*/;
assign _3047_ = D[23] ^ Q[17] /*6722*/;
assign _3044_ = _2724_ & _3047_ /*6718*/;
assign _3045_ = _2724_ ^ _3047_ /*6721*/;
assign _3046_ = _3038_ & _3045_ /*6719*/;
assign _2918_ = _3038_ ^ _3045_ /*6720*/;
assign _3043_ = _3044_ | _3046_ /*6717*/;
assign _3052_ = D[24] ^ Q[17] /*6716*/;
assign _3049_ = _2725_ & _3052_ /*6712*/;
assign _3050_ = _2725_ ^ _3052_ /*6715*/;
assign _3051_ = _3043_ & _3050_ /*6713*/;
assign _2919_ = _3043_ ^ _3050_ /*6714*/;
assign _3048_ = _3049_ | _3051_ /*6711*/;
assign _3057_ = D[25] ^ Q[17] /*6710*/;
assign _3054_ = _2726_ & _3057_ /*6706*/;
assign _3055_ = _2726_ ^ _3057_ /*6709*/;
assign _3056_ = _3048_ & _3055_ /*6707*/;
assign _2920_ = _3048_ ^ _3055_ /*6708*/;
assign _3053_ = _3054_ | _3056_ /*6705*/;
assign _3062_ = D[26] ^ Q[17] /*6704*/;
assign _3059_ = _2727_ & _3062_ /*6700*/;
assign _3060_ = _2727_ ^ _3062_ /*6703*/;
assign _3061_ = _3053_ & _3060_ /*6701*/;
assign _2921_ = _3053_ ^ _3060_ /*6702*/;
assign _3058_ = _3059_ | _3061_ /*6699*/;
assign _3067_ = D[27] ^ Q[17] /*6698*/;
assign _3064_ = _2728_ & _3067_ /*6694*/;
assign _3065_ = _2728_ ^ _3067_ /*6697*/;
assign _3066_ = _3058_ & _3065_ /*6695*/;
assign _2922_ = _3058_ ^ _3065_ /*6696*/;
assign _3063_ = _3064_ | _3066_ /*6693*/;
assign _3072_ = D[28] ^ Q[17] /*6692*/;
assign _3069_ = _2729_ & _3072_ /*6688*/;
assign _3070_ = _2729_ ^ _3072_ /*6691*/;
assign _3071_ = _3063_ & _3070_ /*6689*/;
assign _2923_ = _3063_ ^ _3070_ /*6690*/;
assign _3068_ = _3069_ | _3071_ /*6687*/;
assign _3077_ = D[29] ^ Q[17] /*6686*/;
assign _3074_ = _2730_ & _3077_ /*6682*/;
assign _3075_ = _2730_ ^ _3077_ /*6685*/;
assign _3076_ = _3068_ & _3075_ /*6683*/;
assign _2924_ = _3068_ ^ _3075_ /*6684*/;
assign _3073_ = _3074_ | _3076_ /*6681*/;
assign _3082_ = D[30] ^ Q[17] /*6680*/;
assign _3079_ = _2731_ & _3082_ /*6676*/;
assign _3080_ = _2731_ ^ _3082_ /*6679*/;
assign _3081_ = _3073_ & _3080_ /*6677*/;
assign _2925_ = _3073_ ^ _3080_ /*6678*/;
assign _3078_ = _3079_ | _3081_ /*6675*/;
assign _3086_ = zeroWire ^ Q[17] /*6674*/;
assign _3083_ = _2732_ & _3086_ /*6670*/;
assign _3084_ = _2732_ ^ _3086_ /*6673*/;
assign _3085_ = _3078_ & _3084_ /*6671*/;
assign _2926_ = _3078_ ^ _3084_ /*6672*/;
assign Q[16] = _3083_ | _3085_ /*6669*/;
assign _3125_ = D[0] ^ Q[16] /*6475*/;
assign _3122_ = R_0[15] & _3125_ /*6471*/;
assign _3123_ = R_0[15] ^ _3125_ /*6474*/;
assign _3124_ = Q[16] & _3123_ /*6472*/;
assign _3088_ = Q[16] ^ _3123_ /*6473*/;
assign _3121_ = _3122_ | _3124_ /*6470*/;
assign _3130_ = D[1] ^ Q[16] /*6469*/;
assign _3127_ = _2895_ & _3130_ /*6465*/;
assign _3128_ = _2895_ ^ _3130_ /*6468*/;
assign _3129_ = _3121_ & _3128_ /*6466*/;
assign _3089_ = _3121_ ^ _3128_ /*6467*/;
assign _3126_ = _3127_ | _3129_ /*6464*/;
assign _3135_ = D[2] ^ Q[16] /*6463*/;
assign _3132_ = _2896_ & _3135_ /*6459*/;
assign _3133_ = _2896_ ^ _3135_ /*6462*/;
assign _3134_ = _3126_ & _3133_ /*6460*/;
assign _3090_ = _3126_ ^ _3133_ /*6461*/;
assign _3131_ = _3132_ | _3134_ /*6458*/;
assign _3140_ = D[3] ^ Q[16] /*6457*/;
assign _3137_ = _2897_ & _3140_ /*6453*/;
assign _3138_ = _2897_ ^ _3140_ /*6456*/;
assign _3139_ = _3131_ & _3138_ /*6454*/;
assign _3091_ = _3131_ ^ _3138_ /*6455*/;
assign _3136_ = _3137_ | _3139_ /*6452*/;
assign _3145_ = D[4] ^ Q[16] /*6451*/;
assign _3142_ = _2898_ & _3145_ /*6447*/;
assign _3143_ = _2898_ ^ _3145_ /*6450*/;
assign _3144_ = _3136_ & _3143_ /*6448*/;
assign _3092_ = _3136_ ^ _3143_ /*6449*/;
assign _3141_ = _3142_ | _3144_ /*6446*/;
assign _3150_ = D[5] ^ Q[16] /*6445*/;
assign _3147_ = _2899_ & _3150_ /*6441*/;
assign _3148_ = _2899_ ^ _3150_ /*6444*/;
assign _3149_ = _3141_ & _3148_ /*6442*/;
assign _3093_ = _3141_ ^ _3148_ /*6443*/;
assign _3146_ = _3147_ | _3149_ /*6440*/;
assign _3155_ = D[6] ^ Q[16] /*6439*/;
assign _3152_ = _2900_ & _3155_ /*6435*/;
assign _3153_ = _2900_ ^ _3155_ /*6438*/;
assign _3154_ = _3146_ & _3153_ /*6436*/;
assign _3094_ = _3146_ ^ _3153_ /*6437*/;
assign _3151_ = _3152_ | _3154_ /*6434*/;
assign _3160_ = D[7] ^ Q[16] /*6433*/;
assign _3157_ = _2901_ & _3160_ /*6429*/;
assign _3158_ = _2901_ ^ _3160_ /*6432*/;
assign _3159_ = _3151_ & _3158_ /*6430*/;
assign _3095_ = _3151_ ^ _3158_ /*6431*/;
assign _3156_ = _3157_ | _3159_ /*6428*/;
assign _3165_ = D[8] ^ Q[16] /*6427*/;
assign _3162_ = _2902_ & _3165_ /*6423*/;
assign _3163_ = _2902_ ^ _3165_ /*6426*/;
assign _3164_ = _3156_ & _3163_ /*6424*/;
assign _3096_ = _3156_ ^ _3163_ /*6425*/;
assign _3161_ = _3162_ | _3164_ /*6422*/;
assign _3170_ = D[9] ^ Q[16] /*6421*/;
assign _3167_ = _2903_ & _3170_ /*6417*/;
assign _3168_ = _2903_ ^ _3170_ /*6420*/;
assign _3169_ = _3161_ & _3168_ /*6418*/;
assign _3097_ = _3161_ ^ _3168_ /*6419*/;
assign _3166_ = _3167_ | _3169_ /*6416*/;
assign _3175_ = D[10] ^ Q[16] /*6415*/;
assign _3172_ = _2904_ & _3175_ /*6411*/;
assign _3173_ = _2904_ ^ _3175_ /*6414*/;
assign _3174_ = _3166_ & _3173_ /*6412*/;
assign _3098_ = _3166_ ^ _3173_ /*6413*/;
assign _3171_ = _3172_ | _3174_ /*6410*/;
assign _3180_ = D[11] ^ Q[16] /*6409*/;
assign _3177_ = _2905_ & _3180_ /*6405*/;
assign _3178_ = _2905_ ^ _3180_ /*6408*/;
assign _3179_ = _3171_ & _3178_ /*6406*/;
assign _3099_ = _3171_ ^ _3178_ /*6407*/;
assign _3176_ = _3177_ | _3179_ /*6404*/;
assign _3185_ = D[12] ^ Q[16] /*6403*/;
assign _3182_ = _2906_ & _3185_ /*6399*/;
assign _3183_ = _2906_ ^ _3185_ /*6402*/;
assign _3184_ = _3176_ & _3183_ /*6400*/;
assign _3100_ = _3176_ ^ _3183_ /*6401*/;
assign _3181_ = _3182_ | _3184_ /*6398*/;
assign _3190_ = D[13] ^ Q[16] /*6397*/;
assign _3187_ = _2907_ & _3190_ /*6393*/;
assign _3188_ = _2907_ ^ _3190_ /*6396*/;
assign _3189_ = _3181_ & _3188_ /*6394*/;
assign _3101_ = _3181_ ^ _3188_ /*6395*/;
assign _3186_ = _3187_ | _3189_ /*6392*/;
assign _3195_ = D[14] ^ Q[16] /*6391*/;
assign _3192_ = _2908_ & _3195_ /*6387*/;
assign _3193_ = _2908_ ^ _3195_ /*6390*/;
assign _3194_ = _3186_ & _3193_ /*6388*/;
assign _3102_ = _3186_ ^ _3193_ /*6389*/;
assign _3191_ = _3192_ | _3194_ /*6386*/;
assign _3200_ = D[15] ^ Q[16] /*6385*/;
assign _3197_ = _2909_ & _3200_ /*6381*/;
assign _3198_ = _2909_ ^ _3200_ /*6384*/;
assign _3199_ = _3191_ & _3198_ /*6382*/;
assign _3103_ = _3191_ ^ _3198_ /*6383*/;
assign _3196_ = _3197_ | _3199_ /*6380*/;
assign _3205_ = D[16] ^ Q[16] /*6379*/;
assign _3202_ = _2910_ & _3205_ /*6375*/;
assign _3203_ = _2910_ ^ _3205_ /*6378*/;
assign _3204_ = _3196_ & _3203_ /*6376*/;
assign _3104_ = _3196_ ^ _3203_ /*6377*/;
assign _3201_ = _3202_ | _3204_ /*6374*/;
assign _3210_ = D[17] ^ Q[16] /*6373*/;
assign _3207_ = _2911_ & _3210_ /*6369*/;
assign _3208_ = _2911_ ^ _3210_ /*6372*/;
assign _3209_ = _3201_ & _3208_ /*6370*/;
assign _3105_ = _3201_ ^ _3208_ /*6371*/;
assign _3206_ = _3207_ | _3209_ /*6368*/;
assign _3215_ = D[18] ^ Q[16] /*6367*/;
assign _3212_ = _2912_ & _3215_ /*6363*/;
assign _3213_ = _2912_ ^ _3215_ /*6366*/;
assign _3214_ = _3206_ & _3213_ /*6364*/;
assign _3106_ = _3206_ ^ _3213_ /*6365*/;
assign _3211_ = _3212_ | _3214_ /*6362*/;
assign _3220_ = D[19] ^ Q[16] /*6361*/;
assign _3217_ = _2913_ & _3220_ /*6357*/;
assign _3218_ = _2913_ ^ _3220_ /*6360*/;
assign _3219_ = _3211_ & _3218_ /*6358*/;
assign _3107_ = _3211_ ^ _3218_ /*6359*/;
assign _3216_ = _3217_ | _3219_ /*6356*/;
assign _3225_ = D[20] ^ Q[16] /*6355*/;
assign _3222_ = _2914_ & _3225_ /*6351*/;
assign _3223_ = _2914_ ^ _3225_ /*6354*/;
assign _3224_ = _3216_ & _3223_ /*6352*/;
assign _3108_ = _3216_ ^ _3223_ /*6353*/;
assign _3221_ = _3222_ | _3224_ /*6350*/;
assign _3230_ = D[21] ^ Q[16] /*6349*/;
assign _3227_ = _2915_ & _3230_ /*6345*/;
assign _3228_ = _2915_ ^ _3230_ /*6348*/;
assign _3229_ = _3221_ & _3228_ /*6346*/;
assign _3109_ = _3221_ ^ _3228_ /*6347*/;
assign _3226_ = _3227_ | _3229_ /*6344*/;
assign _3235_ = D[22] ^ Q[16] /*6343*/;
assign _3232_ = _2916_ & _3235_ /*6339*/;
assign _3233_ = _2916_ ^ _3235_ /*6342*/;
assign _3234_ = _3226_ & _3233_ /*6340*/;
assign _3110_ = _3226_ ^ _3233_ /*6341*/;
assign _3231_ = _3232_ | _3234_ /*6338*/;
assign _3240_ = D[23] ^ Q[16] /*6337*/;
assign _3237_ = _2917_ & _3240_ /*6333*/;
assign _3238_ = _2917_ ^ _3240_ /*6336*/;
assign _3239_ = _3231_ & _3238_ /*6334*/;
assign _3111_ = _3231_ ^ _3238_ /*6335*/;
assign _3236_ = _3237_ | _3239_ /*6332*/;
assign _3245_ = D[24] ^ Q[16] /*6331*/;
assign _3242_ = _2918_ & _3245_ /*6327*/;
assign _3243_ = _2918_ ^ _3245_ /*6330*/;
assign _3244_ = _3236_ & _3243_ /*6328*/;
assign _3112_ = _3236_ ^ _3243_ /*6329*/;
assign _3241_ = _3242_ | _3244_ /*6326*/;
assign _3250_ = D[25] ^ Q[16] /*6325*/;
assign _3247_ = _2919_ & _3250_ /*6321*/;
assign _3248_ = _2919_ ^ _3250_ /*6324*/;
assign _3249_ = _3241_ & _3248_ /*6322*/;
assign _3113_ = _3241_ ^ _3248_ /*6323*/;
assign _3246_ = _3247_ | _3249_ /*6320*/;
assign _3255_ = D[26] ^ Q[16] /*6319*/;
assign _3252_ = _2920_ & _3255_ /*6315*/;
assign _3253_ = _2920_ ^ _3255_ /*6318*/;
assign _3254_ = _3246_ & _3253_ /*6316*/;
assign _3114_ = _3246_ ^ _3253_ /*6317*/;
assign _3251_ = _3252_ | _3254_ /*6314*/;
assign _3260_ = D[27] ^ Q[16] /*6313*/;
assign _3257_ = _2921_ & _3260_ /*6309*/;
assign _3258_ = _2921_ ^ _3260_ /*6312*/;
assign _3259_ = _3251_ & _3258_ /*6310*/;
assign _3115_ = _3251_ ^ _3258_ /*6311*/;
assign _3256_ = _3257_ | _3259_ /*6308*/;
assign _3265_ = D[28] ^ Q[16] /*6307*/;
assign _3262_ = _2922_ & _3265_ /*6303*/;
assign _3263_ = _2922_ ^ _3265_ /*6306*/;
assign _3264_ = _3256_ & _3263_ /*6304*/;
assign _3116_ = _3256_ ^ _3263_ /*6305*/;
assign _3261_ = _3262_ | _3264_ /*6302*/;
assign _3270_ = D[29] ^ Q[16] /*6301*/;
assign _3267_ = _2923_ & _3270_ /*6297*/;
assign _3268_ = _2923_ ^ _3270_ /*6300*/;
assign _3269_ = _3261_ & _3268_ /*6298*/;
assign _3117_ = _3261_ ^ _3268_ /*6299*/;
assign _3266_ = _3267_ | _3269_ /*6296*/;
assign _3275_ = D[30] ^ Q[16] /*6295*/;
assign _3272_ = _2924_ & _3275_ /*6291*/;
assign _3273_ = _2924_ ^ _3275_ /*6294*/;
assign _3274_ = _3266_ & _3273_ /*6292*/;
assign _3118_ = _3266_ ^ _3273_ /*6293*/;
assign _3271_ = _3272_ | _3274_ /*6290*/;
assign _3279_ = zeroWire ^ Q[16] /*6289*/;
assign _3276_ = _2925_ & _3279_ /*6285*/;
assign _3277_ = _2925_ ^ _3279_ /*6288*/;
assign _3278_ = _3271_ & _3277_ /*6286*/;
assign _3119_ = _3271_ ^ _3277_ /*6287*/;
assign Q[15] = _3276_ | _3278_ /*6284*/;
assign _3318_ = D[0] ^ Q[15] /*6090*/;
assign _3315_ = R_0[14] & _3318_ /*6086*/;
assign _3316_ = R_0[14] ^ _3318_ /*6089*/;
assign _3317_ = Q[15] & _3316_ /*6087*/;
assign _3281_ = Q[15] ^ _3316_ /*6088*/;
assign _3314_ = _3315_ | _3317_ /*6085*/;
assign _3323_ = D[1] ^ Q[15] /*6084*/;
assign _3320_ = _3088_ & _3323_ /*6080*/;
assign _3321_ = _3088_ ^ _3323_ /*6083*/;
assign _3322_ = _3314_ & _3321_ /*6081*/;
assign _3282_ = _3314_ ^ _3321_ /*6082*/;
assign _3319_ = _3320_ | _3322_ /*6079*/;
assign _3328_ = D[2] ^ Q[15] /*6078*/;
assign _3325_ = _3089_ & _3328_ /*6074*/;
assign _3326_ = _3089_ ^ _3328_ /*6077*/;
assign _3327_ = _3319_ & _3326_ /*6075*/;
assign _3283_ = _3319_ ^ _3326_ /*6076*/;
assign _3324_ = _3325_ | _3327_ /*6073*/;
assign _3333_ = D[3] ^ Q[15] /*6072*/;
assign _3330_ = _3090_ & _3333_ /*6068*/;
assign _3331_ = _3090_ ^ _3333_ /*6071*/;
assign _3332_ = _3324_ & _3331_ /*6069*/;
assign _3284_ = _3324_ ^ _3331_ /*6070*/;
assign _3329_ = _3330_ | _3332_ /*6067*/;
assign _3338_ = D[4] ^ Q[15] /*6066*/;
assign _3335_ = _3091_ & _3338_ /*6062*/;
assign _3336_ = _3091_ ^ _3338_ /*6065*/;
assign _3337_ = _3329_ & _3336_ /*6063*/;
assign _3285_ = _3329_ ^ _3336_ /*6064*/;
assign _3334_ = _3335_ | _3337_ /*6061*/;
assign _3343_ = D[5] ^ Q[15] /*6060*/;
assign _3340_ = _3092_ & _3343_ /*6056*/;
assign _3341_ = _3092_ ^ _3343_ /*6059*/;
assign _3342_ = _3334_ & _3341_ /*6057*/;
assign _3286_ = _3334_ ^ _3341_ /*6058*/;
assign _3339_ = _3340_ | _3342_ /*6055*/;
assign _3348_ = D[6] ^ Q[15] /*6054*/;
assign _3345_ = _3093_ & _3348_ /*6050*/;
assign _3346_ = _3093_ ^ _3348_ /*6053*/;
assign _3347_ = _3339_ & _3346_ /*6051*/;
assign _3287_ = _3339_ ^ _3346_ /*6052*/;
assign _3344_ = _3345_ | _3347_ /*6049*/;
assign _3353_ = D[7] ^ Q[15] /*6048*/;
assign _3350_ = _3094_ & _3353_ /*6044*/;
assign _3351_ = _3094_ ^ _3353_ /*6047*/;
assign _3352_ = _3344_ & _3351_ /*6045*/;
assign _3288_ = _3344_ ^ _3351_ /*6046*/;
assign _3349_ = _3350_ | _3352_ /*6043*/;
assign _3358_ = D[8] ^ Q[15] /*6042*/;
assign _3355_ = _3095_ & _3358_ /*6038*/;
assign _3356_ = _3095_ ^ _3358_ /*6041*/;
assign _3357_ = _3349_ & _3356_ /*6039*/;
assign _3289_ = _3349_ ^ _3356_ /*6040*/;
assign _3354_ = _3355_ | _3357_ /*6037*/;
assign _3363_ = D[9] ^ Q[15] /*6036*/;
assign _3360_ = _3096_ & _3363_ /*6032*/;
assign _3361_ = _3096_ ^ _3363_ /*6035*/;
assign _3362_ = _3354_ & _3361_ /*6033*/;
assign _3290_ = _3354_ ^ _3361_ /*6034*/;
assign _3359_ = _3360_ | _3362_ /*6031*/;
assign _3368_ = D[10] ^ Q[15] /*6030*/;
assign _3365_ = _3097_ & _3368_ /*6026*/;
assign _3366_ = _3097_ ^ _3368_ /*6029*/;
assign _3367_ = _3359_ & _3366_ /*6027*/;
assign _3291_ = _3359_ ^ _3366_ /*6028*/;
assign _3364_ = _3365_ | _3367_ /*6025*/;
assign _3373_ = D[11] ^ Q[15] /*6024*/;
assign _3370_ = _3098_ & _3373_ /*6020*/;
assign _3371_ = _3098_ ^ _3373_ /*6023*/;
assign _3372_ = _3364_ & _3371_ /*6021*/;
assign _3292_ = _3364_ ^ _3371_ /*6022*/;
assign _3369_ = _3370_ | _3372_ /*6019*/;
assign _3378_ = D[12] ^ Q[15] /*6018*/;
assign _3375_ = _3099_ & _3378_ /*6014*/;
assign _3376_ = _3099_ ^ _3378_ /*6017*/;
assign _3377_ = _3369_ & _3376_ /*6015*/;
assign _3293_ = _3369_ ^ _3376_ /*6016*/;
assign _3374_ = _3375_ | _3377_ /*6013*/;
assign _3383_ = D[13] ^ Q[15] /*6012*/;
assign _3380_ = _3100_ & _3383_ /*6008*/;
assign _3381_ = _3100_ ^ _3383_ /*6011*/;
assign _3382_ = _3374_ & _3381_ /*6009*/;
assign _3294_ = _3374_ ^ _3381_ /*6010*/;
assign _3379_ = _3380_ | _3382_ /*6007*/;
assign _3388_ = D[14] ^ Q[15] /*6006*/;
assign _3385_ = _3101_ & _3388_ /*6002*/;
assign _3386_ = _3101_ ^ _3388_ /*6005*/;
assign _3387_ = _3379_ & _3386_ /*6003*/;
assign _3295_ = _3379_ ^ _3386_ /*6004*/;
assign _3384_ = _3385_ | _3387_ /*6001*/;
assign _3393_ = D[15] ^ Q[15] /*6000*/;
assign _3390_ = _3102_ & _3393_ /*5996*/;
assign _3391_ = _3102_ ^ _3393_ /*5999*/;
assign _3392_ = _3384_ & _3391_ /*5997*/;
assign _3296_ = _3384_ ^ _3391_ /*5998*/;
assign _3389_ = _3390_ | _3392_ /*5995*/;
assign _3398_ = D[16] ^ Q[15] /*5994*/;
assign _3395_ = _3103_ & _3398_ /*5990*/;
assign _3396_ = _3103_ ^ _3398_ /*5993*/;
assign _3397_ = _3389_ & _3396_ /*5991*/;
assign _3297_ = _3389_ ^ _3396_ /*5992*/;
assign _3394_ = _3395_ | _3397_ /*5989*/;
assign _3403_ = D[17] ^ Q[15] /*5988*/;
assign _3400_ = _3104_ & _3403_ /*5984*/;
assign _3401_ = _3104_ ^ _3403_ /*5987*/;
assign _3402_ = _3394_ & _3401_ /*5985*/;
assign _3298_ = _3394_ ^ _3401_ /*5986*/;
assign _3399_ = _3400_ | _3402_ /*5983*/;
assign _3408_ = D[18] ^ Q[15] /*5982*/;
assign _3405_ = _3105_ & _3408_ /*5978*/;
assign _3406_ = _3105_ ^ _3408_ /*5981*/;
assign _3407_ = _3399_ & _3406_ /*5979*/;
assign _3299_ = _3399_ ^ _3406_ /*5980*/;
assign _3404_ = _3405_ | _3407_ /*5977*/;
assign _3413_ = D[19] ^ Q[15] /*5976*/;
assign _3410_ = _3106_ & _3413_ /*5972*/;
assign _3411_ = _3106_ ^ _3413_ /*5975*/;
assign _3412_ = _3404_ & _3411_ /*5973*/;
assign _3300_ = _3404_ ^ _3411_ /*5974*/;
assign _3409_ = _3410_ | _3412_ /*5971*/;
assign _3418_ = D[20] ^ Q[15] /*5970*/;
assign _3415_ = _3107_ & _3418_ /*5966*/;
assign _3416_ = _3107_ ^ _3418_ /*5969*/;
assign _3417_ = _3409_ & _3416_ /*5967*/;
assign _3301_ = _3409_ ^ _3416_ /*5968*/;
assign _3414_ = _3415_ | _3417_ /*5965*/;
assign _3423_ = D[21] ^ Q[15] /*5964*/;
assign _3420_ = _3108_ & _3423_ /*5960*/;
assign _3421_ = _3108_ ^ _3423_ /*5963*/;
assign _3422_ = _3414_ & _3421_ /*5961*/;
assign _3302_ = _3414_ ^ _3421_ /*5962*/;
assign _3419_ = _3420_ | _3422_ /*5959*/;
assign _3428_ = D[22] ^ Q[15] /*5958*/;
assign _3425_ = _3109_ & _3428_ /*5954*/;
assign _3426_ = _3109_ ^ _3428_ /*5957*/;
assign _3427_ = _3419_ & _3426_ /*5955*/;
assign _3303_ = _3419_ ^ _3426_ /*5956*/;
assign _3424_ = _3425_ | _3427_ /*5953*/;
assign _3433_ = D[23] ^ Q[15] /*5952*/;
assign _3430_ = _3110_ & _3433_ /*5948*/;
assign _3431_ = _3110_ ^ _3433_ /*5951*/;
assign _3432_ = _3424_ & _3431_ /*5949*/;
assign _3304_ = _3424_ ^ _3431_ /*5950*/;
assign _3429_ = _3430_ | _3432_ /*5947*/;
assign _3438_ = D[24] ^ Q[15] /*5946*/;
assign _3435_ = _3111_ & _3438_ /*5942*/;
assign _3436_ = _3111_ ^ _3438_ /*5945*/;
assign _3437_ = _3429_ & _3436_ /*5943*/;
assign _3305_ = _3429_ ^ _3436_ /*5944*/;
assign _3434_ = _3435_ | _3437_ /*5941*/;
assign _3443_ = D[25] ^ Q[15] /*5940*/;
assign _3440_ = _3112_ & _3443_ /*5936*/;
assign _3441_ = _3112_ ^ _3443_ /*5939*/;
assign _3442_ = _3434_ & _3441_ /*5937*/;
assign _3306_ = _3434_ ^ _3441_ /*5938*/;
assign _3439_ = _3440_ | _3442_ /*5935*/;
assign _3448_ = D[26] ^ Q[15] /*5934*/;
assign _3445_ = _3113_ & _3448_ /*5930*/;
assign _3446_ = _3113_ ^ _3448_ /*5933*/;
assign _3447_ = _3439_ & _3446_ /*5931*/;
assign _3307_ = _3439_ ^ _3446_ /*5932*/;
assign _3444_ = _3445_ | _3447_ /*5929*/;
assign _3453_ = D[27] ^ Q[15] /*5928*/;
assign _3450_ = _3114_ & _3453_ /*5924*/;
assign _3451_ = _3114_ ^ _3453_ /*5927*/;
assign _3452_ = _3444_ & _3451_ /*5925*/;
assign _3308_ = _3444_ ^ _3451_ /*5926*/;
assign _3449_ = _3450_ | _3452_ /*5923*/;
assign _3458_ = D[28] ^ Q[15] /*5922*/;
assign _3455_ = _3115_ & _3458_ /*5918*/;
assign _3456_ = _3115_ ^ _3458_ /*5921*/;
assign _3457_ = _3449_ & _3456_ /*5919*/;
assign _3309_ = _3449_ ^ _3456_ /*5920*/;
assign _3454_ = _3455_ | _3457_ /*5917*/;
assign _3463_ = D[29] ^ Q[15] /*5916*/;
assign _3460_ = _3116_ & _3463_ /*5912*/;
assign _3461_ = _3116_ ^ _3463_ /*5915*/;
assign _3462_ = _3454_ & _3461_ /*5913*/;
assign _3310_ = _3454_ ^ _3461_ /*5914*/;
assign _3459_ = _3460_ | _3462_ /*5911*/;
assign _3468_ = D[30] ^ Q[15] /*5910*/;
assign _3465_ = _3117_ & _3468_ /*5906*/;
assign _3466_ = _3117_ ^ _3468_ /*5909*/;
assign _3467_ = _3459_ & _3466_ /*5907*/;
assign _3311_ = _3459_ ^ _3466_ /*5908*/;
assign _3464_ = _3465_ | _3467_ /*5905*/;
assign _3472_ = zeroWire ^ Q[15] /*5904*/;
assign _3469_ = _3118_ & _3472_ /*5900*/;
assign _3470_ = _3118_ ^ _3472_ /*5903*/;
assign _3471_ = _3464_ & _3470_ /*5901*/;
assign _3312_ = _3464_ ^ _3470_ /*5902*/;
assign Q[14] = _3469_ | _3471_ /*5899*/;
assign _3511_ = D[0] ^ Q[14] /*5705*/;
assign _3508_ = R_0[13] & _3511_ /*5701*/;
assign _3509_ = R_0[13] ^ _3511_ /*5704*/;
assign _3510_ = Q[14] & _3509_ /*5702*/;
assign _3474_ = Q[14] ^ _3509_ /*5703*/;
assign _3507_ = _3508_ | _3510_ /*5700*/;
assign _3516_ = D[1] ^ Q[14] /*5699*/;
assign _3513_ = _3281_ & _3516_ /*5695*/;
assign _3514_ = _3281_ ^ _3516_ /*5698*/;
assign _3515_ = _3507_ & _3514_ /*5696*/;
assign _3475_ = _3507_ ^ _3514_ /*5697*/;
assign _3512_ = _3513_ | _3515_ /*5694*/;
assign _3521_ = D[2] ^ Q[14] /*5693*/;
assign _3518_ = _3282_ & _3521_ /*5689*/;
assign _3519_ = _3282_ ^ _3521_ /*5692*/;
assign _3520_ = _3512_ & _3519_ /*5690*/;
assign _3476_ = _3512_ ^ _3519_ /*5691*/;
assign _3517_ = _3518_ | _3520_ /*5688*/;
assign _3526_ = D[3] ^ Q[14] /*5687*/;
assign _3523_ = _3283_ & _3526_ /*5683*/;
assign _3524_ = _3283_ ^ _3526_ /*5686*/;
assign _3525_ = _3517_ & _3524_ /*5684*/;
assign _3477_ = _3517_ ^ _3524_ /*5685*/;
assign _3522_ = _3523_ | _3525_ /*5682*/;
assign _3531_ = D[4] ^ Q[14] /*5681*/;
assign _3528_ = _3284_ & _3531_ /*5677*/;
assign _3529_ = _3284_ ^ _3531_ /*5680*/;
assign _3530_ = _3522_ & _3529_ /*5678*/;
assign _3478_ = _3522_ ^ _3529_ /*5679*/;
assign _3527_ = _3528_ | _3530_ /*5676*/;
assign _3536_ = D[5] ^ Q[14] /*5675*/;
assign _3533_ = _3285_ & _3536_ /*5671*/;
assign _3534_ = _3285_ ^ _3536_ /*5674*/;
assign _3535_ = _3527_ & _3534_ /*5672*/;
assign _3479_ = _3527_ ^ _3534_ /*5673*/;
assign _3532_ = _3533_ | _3535_ /*5670*/;
assign _3541_ = D[6] ^ Q[14] /*5669*/;
assign _3538_ = _3286_ & _3541_ /*5665*/;
assign _3539_ = _3286_ ^ _3541_ /*5668*/;
assign _3540_ = _3532_ & _3539_ /*5666*/;
assign _3480_ = _3532_ ^ _3539_ /*5667*/;
assign _3537_ = _3538_ | _3540_ /*5664*/;
assign _3546_ = D[7] ^ Q[14] /*5663*/;
assign _3543_ = _3287_ & _3546_ /*5659*/;
assign _3544_ = _3287_ ^ _3546_ /*5662*/;
assign _3545_ = _3537_ & _3544_ /*5660*/;
assign _3481_ = _3537_ ^ _3544_ /*5661*/;
assign _3542_ = _3543_ | _3545_ /*5658*/;
assign _3551_ = D[8] ^ Q[14] /*5657*/;
assign _3548_ = _3288_ & _3551_ /*5653*/;
assign _3549_ = _3288_ ^ _3551_ /*5656*/;
assign _3550_ = _3542_ & _3549_ /*5654*/;
assign _3482_ = _3542_ ^ _3549_ /*5655*/;
assign _3547_ = _3548_ | _3550_ /*5652*/;
assign _3556_ = D[9] ^ Q[14] /*5651*/;
assign _3553_ = _3289_ & _3556_ /*5647*/;
assign _3554_ = _3289_ ^ _3556_ /*5650*/;
assign _3555_ = _3547_ & _3554_ /*5648*/;
assign _3483_ = _3547_ ^ _3554_ /*5649*/;
assign _3552_ = _3553_ | _3555_ /*5646*/;
assign _3561_ = D[10] ^ Q[14] /*5645*/;
assign _3558_ = _3290_ & _3561_ /*5641*/;
assign _3559_ = _3290_ ^ _3561_ /*5644*/;
assign _3560_ = _3552_ & _3559_ /*5642*/;
assign _3484_ = _3552_ ^ _3559_ /*5643*/;
assign _3557_ = _3558_ | _3560_ /*5640*/;
assign _3566_ = D[11] ^ Q[14] /*5639*/;
assign _3563_ = _3291_ & _3566_ /*5635*/;
assign _3564_ = _3291_ ^ _3566_ /*5638*/;
assign _3565_ = _3557_ & _3564_ /*5636*/;
assign _3485_ = _3557_ ^ _3564_ /*5637*/;
assign _3562_ = _3563_ | _3565_ /*5634*/;
assign _3571_ = D[12] ^ Q[14] /*5633*/;
assign _3568_ = _3292_ & _3571_ /*5629*/;
assign _3569_ = _3292_ ^ _3571_ /*5632*/;
assign _3570_ = _3562_ & _3569_ /*5630*/;
assign _3486_ = _3562_ ^ _3569_ /*5631*/;
assign _3567_ = _3568_ | _3570_ /*5628*/;
assign _3576_ = D[13] ^ Q[14] /*5627*/;
assign _3573_ = _3293_ & _3576_ /*5623*/;
assign _3574_ = _3293_ ^ _3576_ /*5626*/;
assign _3575_ = _3567_ & _3574_ /*5624*/;
assign _3487_ = _3567_ ^ _3574_ /*5625*/;
assign _3572_ = _3573_ | _3575_ /*5622*/;
assign _3581_ = D[14] ^ Q[14] /*5621*/;
assign _3578_ = _3294_ & _3581_ /*5617*/;
assign _3579_ = _3294_ ^ _3581_ /*5620*/;
assign _3580_ = _3572_ & _3579_ /*5618*/;
assign _3488_ = _3572_ ^ _3579_ /*5619*/;
assign _3577_ = _3578_ | _3580_ /*5616*/;
assign _3586_ = D[15] ^ Q[14] /*5615*/;
assign _3583_ = _3295_ & _3586_ /*5611*/;
assign _3584_ = _3295_ ^ _3586_ /*5614*/;
assign _3585_ = _3577_ & _3584_ /*5612*/;
assign _3489_ = _3577_ ^ _3584_ /*5613*/;
assign _3582_ = _3583_ | _3585_ /*5610*/;
assign _3591_ = D[16] ^ Q[14] /*5609*/;
assign _3588_ = _3296_ & _3591_ /*5605*/;
assign _3589_ = _3296_ ^ _3591_ /*5608*/;
assign _3590_ = _3582_ & _3589_ /*5606*/;
assign _3490_ = _3582_ ^ _3589_ /*5607*/;
assign _3587_ = _3588_ | _3590_ /*5604*/;
assign _3596_ = D[17] ^ Q[14] /*5603*/;
assign _3593_ = _3297_ & _3596_ /*5599*/;
assign _3594_ = _3297_ ^ _3596_ /*5602*/;
assign _3595_ = _3587_ & _3594_ /*5600*/;
assign _3491_ = _3587_ ^ _3594_ /*5601*/;
assign _3592_ = _3593_ | _3595_ /*5598*/;
assign _3601_ = D[18] ^ Q[14] /*5597*/;
assign _3598_ = _3298_ & _3601_ /*5593*/;
assign _3599_ = _3298_ ^ _3601_ /*5596*/;
assign _3600_ = _3592_ & _3599_ /*5594*/;
assign _3492_ = _3592_ ^ _3599_ /*5595*/;
assign _3597_ = _3598_ | _3600_ /*5592*/;
assign _3606_ = D[19] ^ Q[14] /*5591*/;
assign _3603_ = _3299_ & _3606_ /*5587*/;
assign _3604_ = _3299_ ^ _3606_ /*5590*/;
assign _3605_ = _3597_ & _3604_ /*5588*/;
assign _3493_ = _3597_ ^ _3604_ /*5589*/;
assign _3602_ = _3603_ | _3605_ /*5586*/;
assign _3611_ = D[20] ^ Q[14] /*5585*/;
assign _3608_ = _3300_ & _3611_ /*5581*/;
assign _3609_ = _3300_ ^ _3611_ /*5584*/;
assign _3610_ = _3602_ & _3609_ /*5582*/;
assign _3494_ = _3602_ ^ _3609_ /*5583*/;
assign _3607_ = _3608_ | _3610_ /*5580*/;
assign _3616_ = D[21] ^ Q[14] /*5579*/;
assign _3613_ = _3301_ & _3616_ /*5575*/;
assign _3614_ = _3301_ ^ _3616_ /*5578*/;
assign _3615_ = _3607_ & _3614_ /*5576*/;
assign _3495_ = _3607_ ^ _3614_ /*5577*/;
assign _3612_ = _3613_ | _3615_ /*5574*/;
assign _3621_ = D[22] ^ Q[14] /*5573*/;
assign _3618_ = _3302_ & _3621_ /*5569*/;
assign _3619_ = _3302_ ^ _3621_ /*5572*/;
assign _3620_ = _3612_ & _3619_ /*5570*/;
assign _3496_ = _3612_ ^ _3619_ /*5571*/;
assign _3617_ = _3618_ | _3620_ /*5568*/;
assign _3626_ = D[23] ^ Q[14] /*5567*/;
assign _3623_ = _3303_ & _3626_ /*5563*/;
assign _3624_ = _3303_ ^ _3626_ /*5566*/;
assign _3625_ = _3617_ & _3624_ /*5564*/;
assign _3497_ = _3617_ ^ _3624_ /*5565*/;
assign _3622_ = _3623_ | _3625_ /*5562*/;
assign _3631_ = D[24] ^ Q[14] /*5561*/;
assign _3628_ = _3304_ & _3631_ /*5557*/;
assign _3629_ = _3304_ ^ _3631_ /*5560*/;
assign _3630_ = _3622_ & _3629_ /*5558*/;
assign _3498_ = _3622_ ^ _3629_ /*5559*/;
assign _3627_ = _3628_ | _3630_ /*5556*/;
assign _3636_ = D[25] ^ Q[14] /*5555*/;
assign _3633_ = _3305_ & _3636_ /*5551*/;
assign _3634_ = _3305_ ^ _3636_ /*5554*/;
assign _3635_ = _3627_ & _3634_ /*5552*/;
assign _3499_ = _3627_ ^ _3634_ /*5553*/;
assign _3632_ = _3633_ | _3635_ /*5550*/;
assign _3641_ = D[26] ^ Q[14] /*5549*/;
assign _3638_ = _3306_ & _3641_ /*5545*/;
assign _3639_ = _3306_ ^ _3641_ /*5548*/;
assign _3640_ = _3632_ & _3639_ /*5546*/;
assign _3500_ = _3632_ ^ _3639_ /*5547*/;
assign _3637_ = _3638_ | _3640_ /*5544*/;
assign _3646_ = D[27] ^ Q[14] /*5543*/;
assign _3643_ = _3307_ & _3646_ /*5539*/;
assign _3644_ = _3307_ ^ _3646_ /*5542*/;
assign _3645_ = _3637_ & _3644_ /*5540*/;
assign _3501_ = _3637_ ^ _3644_ /*5541*/;
assign _3642_ = _3643_ | _3645_ /*5538*/;
assign _3651_ = D[28] ^ Q[14] /*5537*/;
assign _3648_ = _3308_ & _3651_ /*5533*/;
assign _3649_ = _3308_ ^ _3651_ /*5536*/;
assign _3650_ = _3642_ & _3649_ /*5534*/;
assign _3502_ = _3642_ ^ _3649_ /*5535*/;
assign _3647_ = _3648_ | _3650_ /*5532*/;
assign _3656_ = D[29] ^ Q[14] /*5531*/;
assign _3653_ = _3309_ & _3656_ /*5527*/;
assign _3654_ = _3309_ ^ _3656_ /*5530*/;
assign _3655_ = _3647_ & _3654_ /*5528*/;
assign _3503_ = _3647_ ^ _3654_ /*5529*/;
assign _3652_ = _3653_ | _3655_ /*5526*/;
assign _3661_ = D[30] ^ Q[14] /*5525*/;
assign _3658_ = _3310_ & _3661_ /*5521*/;
assign _3659_ = _3310_ ^ _3661_ /*5524*/;
assign _3660_ = _3652_ & _3659_ /*5522*/;
assign _3504_ = _3652_ ^ _3659_ /*5523*/;
assign _3657_ = _3658_ | _3660_ /*5520*/;
assign _3665_ = zeroWire ^ Q[14] /*5519*/;
assign _3662_ = _3311_ & _3665_ /*5515*/;
assign _3663_ = _3311_ ^ _3665_ /*5518*/;
assign _3664_ = _3657_ & _3663_ /*5516*/;
assign _3505_ = _3657_ ^ _3663_ /*5517*/;
assign Q[13] = _3662_ | _3664_ /*5514*/;
assign _3704_ = D[0] ^ Q[13] /*5320*/;
assign _3701_ = R_0[12] & _3704_ /*5316*/;
assign _3702_ = R_0[12] ^ _3704_ /*5319*/;
assign _3703_ = Q[13] & _3702_ /*5317*/;
assign _3667_ = Q[13] ^ _3702_ /*5318*/;
assign _3700_ = _3701_ | _3703_ /*5315*/;
assign _3709_ = D[1] ^ Q[13] /*5314*/;
assign _3706_ = _3474_ & _3709_ /*5310*/;
assign _3707_ = _3474_ ^ _3709_ /*5313*/;
assign _3708_ = _3700_ & _3707_ /*5311*/;
assign _3668_ = _3700_ ^ _3707_ /*5312*/;
assign _3705_ = _3706_ | _3708_ /*5309*/;
assign _3714_ = D[2] ^ Q[13] /*5308*/;
assign _3711_ = _3475_ & _3714_ /*5304*/;
assign _3712_ = _3475_ ^ _3714_ /*5307*/;
assign _3713_ = _3705_ & _3712_ /*5305*/;
assign _3669_ = _3705_ ^ _3712_ /*5306*/;
assign _3710_ = _3711_ | _3713_ /*5303*/;
assign _3719_ = D[3] ^ Q[13] /*5302*/;
assign _3716_ = _3476_ & _3719_ /*5298*/;
assign _3717_ = _3476_ ^ _3719_ /*5301*/;
assign _3718_ = _3710_ & _3717_ /*5299*/;
assign _3670_ = _3710_ ^ _3717_ /*5300*/;
assign _3715_ = _3716_ | _3718_ /*5297*/;
assign _3724_ = D[4] ^ Q[13] /*5296*/;
assign _3721_ = _3477_ & _3724_ /*5292*/;
assign _3722_ = _3477_ ^ _3724_ /*5295*/;
assign _3723_ = _3715_ & _3722_ /*5293*/;
assign _3671_ = _3715_ ^ _3722_ /*5294*/;
assign _3720_ = _3721_ | _3723_ /*5291*/;
assign _3729_ = D[5] ^ Q[13] /*5290*/;
assign _3726_ = _3478_ & _3729_ /*5286*/;
assign _3727_ = _3478_ ^ _3729_ /*5289*/;
assign _3728_ = _3720_ & _3727_ /*5287*/;
assign _3672_ = _3720_ ^ _3727_ /*5288*/;
assign _3725_ = _3726_ | _3728_ /*5285*/;
assign _3734_ = D[6] ^ Q[13] /*5284*/;
assign _3731_ = _3479_ & _3734_ /*5280*/;
assign _3732_ = _3479_ ^ _3734_ /*5283*/;
assign _3733_ = _3725_ & _3732_ /*5281*/;
assign _3673_ = _3725_ ^ _3732_ /*5282*/;
assign _3730_ = _3731_ | _3733_ /*5279*/;
assign _3739_ = D[7] ^ Q[13] /*5278*/;
assign _3736_ = _3480_ & _3739_ /*5274*/;
assign _3737_ = _3480_ ^ _3739_ /*5277*/;
assign _3738_ = _3730_ & _3737_ /*5275*/;
assign _3674_ = _3730_ ^ _3737_ /*5276*/;
assign _3735_ = _3736_ | _3738_ /*5273*/;
assign _3744_ = D[8] ^ Q[13] /*5272*/;
assign _3741_ = _3481_ & _3744_ /*5268*/;
assign _3742_ = _3481_ ^ _3744_ /*5271*/;
assign _3743_ = _3735_ & _3742_ /*5269*/;
assign _3675_ = _3735_ ^ _3742_ /*5270*/;
assign _3740_ = _3741_ | _3743_ /*5267*/;
assign _3749_ = D[9] ^ Q[13] /*5266*/;
assign _3746_ = _3482_ & _3749_ /*5262*/;
assign _3747_ = _3482_ ^ _3749_ /*5265*/;
assign _3748_ = _3740_ & _3747_ /*5263*/;
assign _3676_ = _3740_ ^ _3747_ /*5264*/;
assign _3745_ = _3746_ | _3748_ /*5261*/;
assign _3754_ = D[10] ^ Q[13] /*5260*/;
assign _3751_ = _3483_ & _3754_ /*5256*/;
assign _3752_ = _3483_ ^ _3754_ /*5259*/;
assign _3753_ = _3745_ & _3752_ /*5257*/;
assign _3677_ = _3745_ ^ _3752_ /*5258*/;
assign _3750_ = _3751_ | _3753_ /*5255*/;
assign _3759_ = D[11] ^ Q[13] /*5254*/;
assign _3756_ = _3484_ & _3759_ /*5250*/;
assign _3757_ = _3484_ ^ _3759_ /*5253*/;
assign _3758_ = _3750_ & _3757_ /*5251*/;
assign _3678_ = _3750_ ^ _3757_ /*5252*/;
assign _3755_ = _3756_ | _3758_ /*5249*/;
assign _3764_ = D[12] ^ Q[13] /*5248*/;
assign _3761_ = _3485_ & _3764_ /*5244*/;
assign _3762_ = _3485_ ^ _3764_ /*5247*/;
assign _3763_ = _3755_ & _3762_ /*5245*/;
assign _3679_ = _3755_ ^ _3762_ /*5246*/;
assign _3760_ = _3761_ | _3763_ /*5243*/;
assign _3769_ = D[13] ^ Q[13] /*5242*/;
assign _3766_ = _3486_ & _3769_ /*5238*/;
assign _3767_ = _3486_ ^ _3769_ /*5241*/;
assign _3768_ = _3760_ & _3767_ /*5239*/;
assign _3680_ = _3760_ ^ _3767_ /*5240*/;
assign _3765_ = _3766_ | _3768_ /*5237*/;
assign _3774_ = D[14] ^ Q[13] /*5236*/;
assign _3771_ = _3487_ & _3774_ /*5232*/;
assign _3772_ = _3487_ ^ _3774_ /*5235*/;
assign _3773_ = _3765_ & _3772_ /*5233*/;
assign _3681_ = _3765_ ^ _3772_ /*5234*/;
assign _3770_ = _3771_ | _3773_ /*5231*/;
assign _3779_ = D[15] ^ Q[13] /*5230*/;
assign _3776_ = _3488_ & _3779_ /*5226*/;
assign _3777_ = _3488_ ^ _3779_ /*5229*/;
assign _3778_ = _3770_ & _3777_ /*5227*/;
assign _3682_ = _3770_ ^ _3777_ /*5228*/;
assign _3775_ = _3776_ | _3778_ /*5225*/;
assign _3784_ = D[16] ^ Q[13] /*5224*/;
assign _3781_ = _3489_ & _3784_ /*5220*/;
assign _3782_ = _3489_ ^ _3784_ /*5223*/;
assign _3783_ = _3775_ & _3782_ /*5221*/;
assign _3683_ = _3775_ ^ _3782_ /*5222*/;
assign _3780_ = _3781_ | _3783_ /*5219*/;
assign _3789_ = D[17] ^ Q[13] /*5218*/;
assign _3786_ = _3490_ & _3789_ /*5214*/;
assign _3787_ = _3490_ ^ _3789_ /*5217*/;
assign _3788_ = _3780_ & _3787_ /*5215*/;
assign _3684_ = _3780_ ^ _3787_ /*5216*/;
assign _3785_ = _3786_ | _3788_ /*5213*/;
assign _3794_ = D[18] ^ Q[13] /*5212*/;
assign _3791_ = _3491_ & _3794_ /*5208*/;
assign _3792_ = _3491_ ^ _3794_ /*5211*/;
assign _3793_ = _3785_ & _3792_ /*5209*/;
assign _3685_ = _3785_ ^ _3792_ /*5210*/;
assign _3790_ = _3791_ | _3793_ /*5207*/;
assign _3799_ = D[19] ^ Q[13] /*5206*/;
assign _3796_ = _3492_ & _3799_ /*5202*/;
assign _3797_ = _3492_ ^ _3799_ /*5205*/;
assign _3798_ = _3790_ & _3797_ /*5203*/;
assign _3686_ = _3790_ ^ _3797_ /*5204*/;
assign _3795_ = _3796_ | _3798_ /*5201*/;
assign _3804_ = D[20] ^ Q[13] /*5200*/;
assign _3801_ = _3493_ & _3804_ /*5196*/;
assign _3802_ = _3493_ ^ _3804_ /*5199*/;
assign _3803_ = _3795_ & _3802_ /*5197*/;
assign _3687_ = _3795_ ^ _3802_ /*5198*/;
assign _3800_ = _3801_ | _3803_ /*5195*/;
assign _3809_ = D[21] ^ Q[13] /*5194*/;
assign _3806_ = _3494_ & _3809_ /*5190*/;
assign _3807_ = _3494_ ^ _3809_ /*5193*/;
assign _3808_ = _3800_ & _3807_ /*5191*/;
assign _3688_ = _3800_ ^ _3807_ /*5192*/;
assign _3805_ = _3806_ | _3808_ /*5189*/;
assign _3814_ = D[22] ^ Q[13] /*5188*/;
assign _3811_ = _3495_ & _3814_ /*5184*/;
assign _3812_ = _3495_ ^ _3814_ /*5187*/;
assign _3813_ = _3805_ & _3812_ /*5185*/;
assign _3689_ = _3805_ ^ _3812_ /*5186*/;
assign _3810_ = _3811_ | _3813_ /*5183*/;
assign _3819_ = D[23] ^ Q[13] /*5182*/;
assign _3816_ = _3496_ & _3819_ /*5178*/;
assign _3817_ = _3496_ ^ _3819_ /*5181*/;
assign _3818_ = _3810_ & _3817_ /*5179*/;
assign _3690_ = _3810_ ^ _3817_ /*5180*/;
assign _3815_ = _3816_ | _3818_ /*5177*/;
assign _3824_ = D[24] ^ Q[13] /*5176*/;
assign _3821_ = _3497_ & _3824_ /*5172*/;
assign _3822_ = _3497_ ^ _3824_ /*5175*/;
assign _3823_ = _3815_ & _3822_ /*5173*/;
assign _3691_ = _3815_ ^ _3822_ /*5174*/;
assign _3820_ = _3821_ | _3823_ /*5171*/;
assign _3829_ = D[25] ^ Q[13] /*5170*/;
assign _3826_ = _3498_ & _3829_ /*5166*/;
assign _3827_ = _3498_ ^ _3829_ /*5169*/;
assign _3828_ = _3820_ & _3827_ /*5167*/;
assign _3692_ = _3820_ ^ _3827_ /*5168*/;
assign _3825_ = _3826_ | _3828_ /*5165*/;
assign _3834_ = D[26] ^ Q[13] /*5164*/;
assign _3831_ = _3499_ & _3834_ /*5160*/;
assign _3832_ = _3499_ ^ _3834_ /*5163*/;
assign _3833_ = _3825_ & _3832_ /*5161*/;
assign _3693_ = _3825_ ^ _3832_ /*5162*/;
assign _3830_ = _3831_ | _3833_ /*5159*/;
assign _3839_ = D[27] ^ Q[13] /*5158*/;
assign _3836_ = _3500_ & _3839_ /*5154*/;
assign _3837_ = _3500_ ^ _3839_ /*5157*/;
assign _3838_ = _3830_ & _3837_ /*5155*/;
assign _3694_ = _3830_ ^ _3837_ /*5156*/;
assign _3835_ = _3836_ | _3838_ /*5153*/;
assign _3844_ = D[28] ^ Q[13] /*5152*/;
assign _3841_ = _3501_ & _3844_ /*5148*/;
assign _3842_ = _3501_ ^ _3844_ /*5151*/;
assign _3843_ = _3835_ & _3842_ /*5149*/;
assign _3695_ = _3835_ ^ _3842_ /*5150*/;
assign _3840_ = _3841_ | _3843_ /*5147*/;
assign _3849_ = D[29] ^ Q[13] /*5146*/;
assign _3846_ = _3502_ & _3849_ /*5142*/;
assign _3847_ = _3502_ ^ _3849_ /*5145*/;
assign _3848_ = _3840_ & _3847_ /*5143*/;
assign _3696_ = _3840_ ^ _3847_ /*5144*/;
assign _3845_ = _3846_ | _3848_ /*5141*/;
assign _3854_ = D[30] ^ Q[13] /*5140*/;
assign _3851_ = _3503_ & _3854_ /*5136*/;
assign _3852_ = _3503_ ^ _3854_ /*5139*/;
assign _3853_ = _3845_ & _3852_ /*5137*/;
assign _3697_ = _3845_ ^ _3852_ /*5138*/;
assign _3850_ = _3851_ | _3853_ /*5135*/;
assign _3858_ = zeroWire ^ Q[13] /*5134*/;
assign _3855_ = _3504_ & _3858_ /*5130*/;
assign _3856_ = _3504_ ^ _3858_ /*5133*/;
assign _3857_ = _3850_ & _3856_ /*5131*/;
assign _3698_ = _3850_ ^ _3856_ /*5132*/;
assign Q[12] = _3855_ | _3857_ /*5129*/;
assign _3897_ = D[0] ^ Q[12] /*4935*/;
assign _3894_ = R_0[11] & _3897_ /*4931*/;
assign _3895_ = R_0[11] ^ _3897_ /*4934*/;
assign _3896_ = Q[12] & _3895_ /*4932*/;
assign _3860_ = Q[12] ^ _3895_ /*4933*/;
assign _3893_ = _3894_ | _3896_ /*4930*/;
assign _3902_ = D[1] ^ Q[12] /*4929*/;
assign _3899_ = _3667_ & _3902_ /*4925*/;
assign _3900_ = _3667_ ^ _3902_ /*4928*/;
assign _3901_ = _3893_ & _3900_ /*4926*/;
assign _3861_ = _3893_ ^ _3900_ /*4927*/;
assign _3898_ = _3899_ | _3901_ /*4924*/;
assign _3907_ = D[2] ^ Q[12] /*4923*/;
assign _3904_ = _3668_ & _3907_ /*4919*/;
assign _3905_ = _3668_ ^ _3907_ /*4922*/;
assign _3906_ = _3898_ & _3905_ /*4920*/;
assign _3862_ = _3898_ ^ _3905_ /*4921*/;
assign _3903_ = _3904_ | _3906_ /*4918*/;
assign _3912_ = D[3] ^ Q[12] /*4917*/;
assign _3909_ = _3669_ & _3912_ /*4913*/;
assign _3910_ = _3669_ ^ _3912_ /*4916*/;
assign _3911_ = _3903_ & _3910_ /*4914*/;
assign _3863_ = _3903_ ^ _3910_ /*4915*/;
assign _3908_ = _3909_ | _3911_ /*4912*/;
assign _3917_ = D[4] ^ Q[12] /*4911*/;
assign _3914_ = _3670_ & _3917_ /*4907*/;
assign _3915_ = _3670_ ^ _3917_ /*4910*/;
assign _3916_ = _3908_ & _3915_ /*4908*/;
assign _3864_ = _3908_ ^ _3915_ /*4909*/;
assign _3913_ = _3914_ | _3916_ /*4906*/;
assign _3922_ = D[5] ^ Q[12] /*4905*/;
assign _3919_ = _3671_ & _3922_ /*4901*/;
assign _3920_ = _3671_ ^ _3922_ /*4904*/;
assign _3921_ = _3913_ & _3920_ /*4902*/;
assign _3865_ = _3913_ ^ _3920_ /*4903*/;
assign _3918_ = _3919_ | _3921_ /*4900*/;
assign _3927_ = D[6] ^ Q[12] /*4899*/;
assign _3924_ = _3672_ & _3927_ /*4895*/;
assign _3925_ = _3672_ ^ _3927_ /*4898*/;
assign _3926_ = _3918_ & _3925_ /*4896*/;
assign _3866_ = _3918_ ^ _3925_ /*4897*/;
assign _3923_ = _3924_ | _3926_ /*4894*/;
assign _3932_ = D[7] ^ Q[12] /*4893*/;
assign _3929_ = _3673_ & _3932_ /*4889*/;
assign _3930_ = _3673_ ^ _3932_ /*4892*/;
assign _3931_ = _3923_ & _3930_ /*4890*/;
assign _3867_ = _3923_ ^ _3930_ /*4891*/;
assign _3928_ = _3929_ | _3931_ /*4888*/;
assign _3937_ = D[8] ^ Q[12] /*4887*/;
assign _3934_ = _3674_ & _3937_ /*4883*/;
assign _3935_ = _3674_ ^ _3937_ /*4886*/;
assign _3936_ = _3928_ & _3935_ /*4884*/;
assign _3868_ = _3928_ ^ _3935_ /*4885*/;
assign _3933_ = _3934_ | _3936_ /*4882*/;
assign _3942_ = D[9] ^ Q[12] /*4881*/;
assign _3939_ = _3675_ & _3942_ /*4877*/;
assign _3940_ = _3675_ ^ _3942_ /*4880*/;
assign _3941_ = _3933_ & _3940_ /*4878*/;
assign _3869_ = _3933_ ^ _3940_ /*4879*/;
assign _3938_ = _3939_ | _3941_ /*4876*/;
assign _3947_ = D[10] ^ Q[12] /*4875*/;
assign _3944_ = _3676_ & _3947_ /*4871*/;
assign _3945_ = _3676_ ^ _3947_ /*4874*/;
assign _3946_ = _3938_ & _3945_ /*4872*/;
assign _3870_ = _3938_ ^ _3945_ /*4873*/;
assign _3943_ = _3944_ | _3946_ /*4870*/;
assign _3952_ = D[11] ^ Q[12] /*4869*/;
assign _3949_ = _3677_ & _3952_ /*4865*/;
assign _3950_ = _3677_ ^ _3952_ /*4868*/;
assign _3951_ = _3943_ & _3950_ /*4866*/;
assign _3871_ = _3943_ ^ _3950_ /*4867*/;
assign _3948_ = _3949_ | _3951_ /*4864*/;
assign _3957_ = D[12] ^ Q[12] /*4863*/;
assign _3954_ = _3678_ & _3957_ /*4859*/;
assign _3955_ = _3678_ ^ _3957_ /*4862*/;
assign _3956_ = _3948_ & _3955_ /*4860*/;
assign _3872_ = _3948_ ^ _3955_ /*4861*/;
assign _3953_ = _3954_ | _3956_ /*4858*/;
assign _3962_ = D[13] ^ Q[12] /*4857*/;
assign _3959_ = _3679_ & _3962_ /*4853*/;
assign _3960_ = _3679_ ^ _3962_ /*4856*/;
assign _3961_ = _3953_ & _3960_ /*4854*/;
assign _3873_ = _3953_ ^ _3960_ /*4855*/;
assign _3958_ = _3959_ | _3961_ /*4852*/;
assign _3967_ = D[14] ^ Q[12] /*4851*/;
assign _3964_ = _3680_ & _3967_ /*4847*/;
assign _3965_ = _3680_ ^ _3967_ /*4850*/;
assign _3966_ = _3958_ & _3965_ /*4848*/;
assign _3874_ = _3958_ ^ _3965_ /*4849*/;
assign _3963_ = _3964_ | _3966_ /*4846*/;
assign _3972_ = D[15] ^ Q[12] /*4845*/;
assign _3969_ = _3681_ & _3972_ /*4841*/;
assign _3970_ = _3681_ ^ _3972_ /*4844*/;
assign _3971_ = _3963_ & _3970_ /*4842*/;
assign _3875_ = _3963_ ^ _3970_ /*4843*/;
assign _3968_ = _3969_ | _3971_ /*4840*/;
assign _3977_ = D[16] ^ Q[12] /*4839*/;
assign _3974_ = _3682_ & _3977_ /*4835*/;
assign _3975_ = _3682_ ^ _3977_ /*4838*/;
assign _3976_ = _3968_ & _3975_ /*4836*/;
assign _3876_ = _3968_ ^ _3975_ /*4837*/;
assign _3973_ = _3974_ | _3976_ /*4834*/;
assign _3982_ = D[17] ^ Q[12] /*4833*/;
assign _3979_ = _3683_ & _3982_ /*4829*/;
assign _3980_ = _3683_ ^ _3982_ /*4832*/;
assign _3981_ = _3973_ & _3980_ /*4830*/;
assign _3877_ = _3973_ ^ _3980_ /*4831*/;
assign _3978_ = _3979_ | _3981_ /*4828*/;
assign _3987_ = D[18] ^ Q[12] /*4827*/;
assign _3984_ = _3684_ & _3987_ /*4823*/;
assign _3985_ = _3684_ ^ _3987_ /*4826*/;
assign _3986_ = _3978_ & _3985_ /*4824*/;
assign _3878_ = _3978_ ^ _3985_ /*4825*/;
assign _3983_ = _3984_ | _3986_ /*4822*/;
assign _3992_ = D[19] ^ Q[12] /*4821*/;
assign _3989_ = _3685_ & _3992_ /*4817*/;
assign _3990_ = _3685_ ^ _3992_ /*4820*/;
assign _3991_ = _3983_ & _3990_ /*4818*/;
assign _3879_ = _3983_ ^ _3990_ /*4819*/;
assign _3988_ = _3989_ | _3991_ /*4816*/;
assign _3997_ = D[20] ^ Q[12] /*4815*/;
assign _3994_ = _3686_ & _3997_ /*4811*/;
assign _3995_ = _3686_ ^ _3997_ /*4814*/;
assign _3996_ = _3988_ & _3995_ /*4812*/;
assign _3880_ = _3988_ ^ _3995_ /*4813*/;
assign _3993_ = _3994_ | _3996_ /*4810*/;
assign _4002_ = D[21] ^ Q[12] /*4809*/;
assign _3999_ = _3687_ & _4002_ /*4805*/;
assign _4000_ = _3687_ ^ _4002_ /*4808*/;
assign _4001_ = _3993_ & _4000_ /*4806*/;
assign _3881_ = _3993_ ^ _4000_ /*4807*/;
assign _3998_ = _3999_ | _4001_ /*4804*/;
assign _4007_ = D[22] ^ Q[12] /*4803*/;
assign _4004_ = _3688_ & _4007_ /*4799*/;
assign _4005_ = _3688_ ^ _4007_ /*4802*/;
assign _4006_ = _3998_ & _4005_ /*4800*/;
assign _3882_ = _3998_ ^ _4005_ /*4801*/;
assign _4003_ = _4004_ | _4006_ /*4798*/;
assign _4012_ = D[23] ^ Q[12] /*4797*/;
assign _4009_ = _3689_ & _4012_ /*4793*/;
assign _4010_ = _3689_ ^ _4012_ /*4796*/;
assign _4011_ = _4003_ & _4010_ /*4794*/;
assign _3883_ = _4003_ ^ _4010_ /*4795*/;
assign _4008_ = _4009_ | _4011_ /*4792*/;
assign _4017_ = D[24] ^ Q[12] /*4791*/;
assign _4014_ = _3690_ & _4017_ /*4787*/;
assign _4015_ = _3690_ ^ _4017_ /*4790*/;
assign _4016_ = _4008_ & _4015_ /*4788*/;
assign _3884_ = _4008_ ^ _4015_ /*4789*/;
assign _4013_ = _4014_ | _4016_ /*4786*/;
assign _4022_ = D[25] ^ Q[12] /*4785*/;
assign _4019_ = _3691_ & _4022_ /*4781*/;
assign _4020_ = _3691_ ^ _4022_ /*4784*/;
assign _4021_ = _4013_ & _4020_ /*4782*/;
assign _3885_ = _4013_ ^ _4020_ /*4783*/;
assign _4018_ = _4019_ | _4021_ /*4780*/;
assign _4027_ = D[26] ^ Q[12] /*4779*/;
assign _4024_ = _3692_ & _4027_ /*4775*/;
assign _4025_ = _3692_ ^ _4027_ /*4778*/;
assign _4026_ = _4018_ & _4025_ /*4776*/;
assign _3886_ = _4018_ ^ _4025_ /*4777*/;
assign _4023_ = _4024_ | _4026_ /*4774*/;
assign _4032_ = D[27] ^ Q[12] /*4773*/;
assign _4029_ = _3693_ & _4032_ /*4769*/;
assign _4030_ = _3693_ ^ _4032_ /*4772*/;
assign _4031_ = _4023_ & _4030_ /*4770*/;
assign _3887_ = _4023_ ^ _4030_ /*4771*/;
assign _4028_ = _4029_ | _4031_ /*4768*/;
assign _4037_ = D[28] ^ Q[12] /*4767*/;
assign _4034_ = _3694_ & _4037_ /*4763*/;
assign _4035_ = _3694_ ^ _4037_ /*4766*/;
assign _4036_ = _4028_ & _4035_ /*4764*/;
assign _3888_ = _4028_ ^ _4035_ /*4765*/;
assign _4033_ = _4034_ | _4036_ /*4762*/;
assign _4042_ = D[29] ^ Q[12] /*4761*/;
assign _4039_ = _3695_ & _4042_ /*4757*/;
assign _4040_ = _3695_ ^ _4042_ /*4760*/;
assign _4041_ = _4033_ & _4040_ /*4758*/;
assign _3889_ = _4033_ ^ _4040_ /*4759*/;
assign _4038_ = _4039_ | _4041_ /*4756*/;
assign _4047_ = D[30] ^ Q[12] /*4755*/;
assign _4044_ = _3696_ & _4047_ /*4751*/;
assign _4045_ = _3696_ ^ _4047_ /*4754*/;
assign _4046_ = _4038_ & _4045_ /*4752*/;
assign _3890_ = _4038_ ^ _4045_ /*4753*/;
assign _4043_ = _4044_ | _4046_ /*4750*/;
assign _4051_ = zeroWire ^ Q[12] /*4749*/;
assign _4048_ = _3697_ & _4051_ /*4745*/;
assign _4049_ = _3697_ ^ _4051_ /*4748*/;
assign _4050_ = _4043_ & _4049_ /*4746*/;
assign _3891_ = _4043_ ^ _4049_ /*4747*/;
assign Q[11] = _4048_ | _4050_ /*4744*/;
assign _4090_ = D[0] ^ Q[11] /*4550*/;
assign _4087_ = R_0[10] & _4090_ /*4546*/;
assign _4088_ = R_0[10] ^ _4090_ /*4549*/;
assign _4089_ = Q[11] & _4088_ /*4547*/;
assign _4053_ = Q[11] ^ _4088_ /*4548*/;
assign _4086_ = _4087_ | _4089_ /*4545*/;
assign _4095_ = D[1] ^ Q[11] /*4544*/;
assign _4092_ = _3860_ & _4095_ /*4540*/;
assign _4093_ = _3860_ ^ _4095_ /*4543*/;
assign _4094_ = _4086_ & _4093_ /*4541*/;
assign _4054_ = _4086_ ^ _4093_ /*4542*/;
assign _4091_ = _4092_ | _4094_ /*4539*/;
assign _4100_ = D[2] ^ Q[11] /*4538*/;
assign _4097_ = _3861_ & _4100_ /*4534*/;
assign _4098_ = _3861_ ^ _4100_ /*4537*/;
assign _4099_ = _4091_ & _4098_ /*4535*/;
assign _4055_ = _4091_ ^ _4098_ /*4536*/;
assign _4096_ = _4097_ | _4099_ /*4533*/;
assign _4105_ = D[3] ^ Q[11] /*4532*/;
assign _4102_ = _3862_ & _4105_ /*4528*/;
assign _4103_ = _3862_ ^ _4105_ /*4531*/;
assign _4104_ = _4096_ & _4103_ /*4529*/;
assign _4056_ = _4096_ ^ _4103_ /*4530*/;
assign _4101_ = _4102_ | _4104_ /*4527*/;
assign _4110_ = D[4] ^ Q[11] /*4526*/;
assign _4107_ = _3863_ & _4110_ /*4522*/;
assign _4108_ = _3863_ ^ _4110_ /*4525*/;
assign _4109_ = _4101_ & _4108_ /*4523*/;
assign _4057_ = _4101_ ^ _4108_ /*4524*/;
assign _4106_ = _4107_ | _4109_ /*4521*/;
assign _4115_ = D[5] ^ Q[11] /*4520*/;
assign _4112_ = _3864_ & _4115_ /*4516*/;
assign _4113_ = _3864_ ^ _4115_ /*4519*/;
assign _4114_ = _4106_ & _4113_ /*4517*/;
assign _4058_ = _4106_ ^ _4113_ /*4518*/;
assign _4111_ = _4112_ | _4114_ /*4515*/;
assign _4120_ = D[6] ^ Q[11] /*4514*/;
assign _4117_ = _3865_ & _4120_ /*4510*/;
assign _4118_ = _3865_ ^ _4120_ /*4513*/;
assign _4119_ = _4111_ & _4118_ /*4511*/;
assign _4059_ = _4111_ ^ _4118_ /*4512*/;
assign _4116_ = _4117_ | _4119_ /*4509*/;
assign _4125_ = D[7] ^ Q[11] /*4508*/;
assign _4122_ = _3866_ & _4125_ /*4504*/;
assign _4123_ = _3866_ ^ _4125_ /*4507*/;
assign _4124_ = _4116_ & _4123_ /*4505*/;
assign _4060_ = _4116_ ^ _4123_ /*4506*/;
assign _4121_ = _4122_ | _4124_ /*4503*/;
assign _4130_ = D[8] ^ Q[11] /*4502*/;
assign _4127_ = _3867_ & _4130_ /*4498*/;
assign _4128_ = _3867_ ^ _4130_ /*4501*/;
assign _4129_ = _4121_ & _4128_ /*4499*/;
assign _4061_ = _4121_ ^ _4128_ /*4500*/;
assign _4126_ = _4127_ | _4129_ /*4497*/;
assign _4135_ = D[9] ^ Q[11] /*4496*/;
assign _4132_ = _3868_ & _4135_ /*4492*/;
assign _4133_ = _3868_ ^ _4135_ /*4495*/;
assign _4134_ = _4126_ & _4133_ /*4493*/;
assign _4062_ = _4126_ ^ _4133_ /*4494*/;
assign _4131_ = _4132_ | _4134_ /*4491*/;
assign _4140_ = D[10] ^ Q[11] /*4490*/;
assign _4137_ = _3869_ & _4140_ /*4486*/;
assign _4138_ = _3869_ ^ _4140_ /*4489*/;
assign _4139_ = _4131_ & _4138_ /*4487*/;
assign _4063_ = _4131_ ^ _4138_ /*4488*/;
assign _4136_ = _4137_ | _4139_ /*4485*/;
assign _4145_ = D[11] ^ Q[11] /*4484*/;
assign _4142_ = _3870_ & _4145_ /*4480*/;
assign _4143_ = _3870_ ^ _4145_ /*4483*/;
assign _4144_ = _4136_ & _4143_ /*4481*/;
assign _4064_ = _4136_ ^ _4143_ /*4482*/;
assign _4141_ = _4142_ | _4144_ /*4479*/;
assign _4150_ = D[12] ^ Q[11] /*4478*/;
assign _4147_ = _3871_ & _4150_ /*4474*/;
assign _4148_ = _3871_ ^ _4150_ /*4477*/;
assign _4149_ = _4141_ & _4148_ /*4475*/;
assign _4065_ = _4141_ ^ _4148_ /*4476*/;
assign _4146_ = _4147_ | _4149_ /*4473*/;
assign _4155_ = D[13] ^ Q[11] /*4472*/;
assign _4152_ = _3872_ & _4155_ /*4468*/;
assign _4153_ = _3872_ ^ _4155_ /*4471*/;
assign _4154_ = _4146_ & _4153_ /*4469*/;
assign _4066_ = _4146_ ^ _4153_ /*4470*/;
assign _4151_ = _4152_ | _4154_ /*4467*/;
assign _4160_ = D[14] ^ Q[11] /*4466*/;
assign _4157_ = _3873_ & _4160_ /*4462*/;
assign _4158_ = _3873_ ^ _4160_ /*4465*/;
assign _4159_ = _4151_ & _4158_ /*4463*/;
assign _4067_ = _4151_ ^ _4158_ /*4464*/;
assign _4156_ = _4157_ | _4159_ /*4461*/;
assign _4165_ = D[15] ^ Q[11] /*4460*/;
assign _4162_ = _3874_ & _4165_ /*4456*/;
assign _4163_ = _3874_ ^ _4165_ /*4459*/;
assign _4164_ = _4156_ & _4163_ /*4457*/;
assign _4068_ = _4156_ ^ _4163_ /*4458*/;
assign _4161_ = _4162_ | _4164_ /*4455*/;
assign _4170_ = D[16] ^ Q[11] /*4454*/;
assign _4167_ = _3875_ & _4170_ /*4450*/;
assign _4168_ = _3875_ ^ _4170_ /*4453*/;
assign _4169_ = _4161_ & _4168_ /*4451*/;
assign _4069_ = _4161_ ^ _4168_ /*4452*/;
assign _4166_ = _4167_ | _4169_ /*4449*/;
assign _4175_ = D[17] ^ Q[11] /*4448*/;
assign _4172_ = _3876_ & _4175_ /*4444*/;
assign _4173_ = _3876_ ^ _4175_ /*4447*/;
assign _4174_ = _4166_ & _4173_ /*4445*/;
assign _4070_ = _4166_ ^ _4173_ /*4446*/;
assign _4171_ = _4172_ | _4174_ /*4443*/;
assign _4180_ = D[18] ^ Q[11] /*4442*/;
assign _4177_ = _3877_ & _4180_ /*4438*/;
assign _4178_ = _3877_ ^ _4180_ /*4441*/;
assign _4179_ = _4171_ & _4178_ /*4439*/;
assign _4071_ = _4171_ ^ _4178_ /*4440*/;
assign _4176_ = _4177_ | _4179_ /*4437*/;
assign _4185_ = D[19] ^ Q[11] /*4436*/;
assign _4182_ = _3878_ & _4185_ /*4432*/;
assign _4183_ = _3878_ ^ _4185_ /*4435*/;
assign _4184_ = _4176_ & _4183_ /*4433*/;
assign _4072_ = _4176_ ^ _4183_ /*4434*/;
assign _4181_ = _4182_ | _4184_ /*4431*/;
assign _4190_ = D[20] ^ Q[11] /*4430*/;
assign _4187_ = _3879_ & _4190_ /*4426*/;
assign _4188_ = _3879_ ^ _4190_ /*4429*/;
assign _4189_ = _4181_ & _4188_ /*4427*/;
assign _4073_ = _4181_ ^ _4188_ /*4428*/;
assign _4186_ = _4187_ | _4189_ /*4425*/;
assign _4195_ = D[21] ^ Q[11] /*4424*/;
assign _4192_ = _3880_ & _4195_ /*4420*/;
assign _4193_ = _3880_ ^ _4195_ /*4423*/;
assign _4194_ = _4186_ & _4193_ /*4421*/;
assign _4074_ = _4186_ ^ _4193_ /*4422*/;
assign _4191_ = _4192_ | _4194_ /*4419*/;
assign _4200_ = D[22] ^ Q[11] /*4418*/;
assign _4197_ = _3881_ & _4200_ /*4414*/;
assign _4198_ = _3881_ ^ _4200_ /*4417*/;
assign _4199_ = _4191_ & _4198_ /*4415*/;
assign _4075_ = _4191_ ^ _4198_ /*4416*/;
assign _4196_ = _4197_ | _4199_ /*4413*/;
assign _4205_ = D[23] ^ Q[11] /*4412*/;
assign _4202_ = _3882_ & _4205_ /*4408*/;
assign _4203_ = _3882_ ^ _4205_ /*4411*/;
assign _4204_ = _4196_ & _4203_ /*4409*/;
assign _4076_ = _4196_ ^ _4203_ /*4410*/;
assign _4201_ = _4202_ | _4204_ /*4407*/;
assign _4210_ = D[24] ^ Q[11] /*4406*/;
assign _4207_ = _3883_ & _4210_ /*4402*/;
assign _4208_ = _3883_ ^ _4210_ /*4405*/;
assign _4209_ = _4201_ & _4208_ /*4403*/;
assign _4077_ = _4201_ ^ _4208_ /*4404*/;
assign _4206_ = _4207_ | _4209_ /*4401*/;
assign _4215_ = D[25] ^ Q[11] /*4400*/;
assign _4212_ = _3884_ & _4215_ /*4396*/;
assign _4213_ = _3884_ ^ _4215_ /*4399*/;
assign _4214_ = _4206_ & _4213_ /*4397*/;
assign _4078_ = _4206_ ^ _4213_ /*4398*/;
assign _4211_ = _4212_ | _4214_ /*4395*/;
assign _4220_ = D[26] ^ Q[11] /*4394*/;
assign _4217_ = _3885_ & _4220_ /*4390*/;
assign _4218_ = _3885_ ^ _4220_ /*4393*/;
assign _4219_ = _4211_ & _4218_ /*4391*/;
assign _4079_ = _4211_ ^ _4218_ /*4392*/;
assign _4216_ = _4217_ | _4219_ /*4389*/;
assign _4225_ = D[27] ^ Q[11] /*4388*/;
assign _4222_ = _3886_ & _4225_ /*4384*/;
assign _4223_ = _3886_ ^ _4225_ /*4387*/;
assign _4224_ = _4216_ & _4223_ /*4385*/;
assign _4080_ = _4216_ ^ _4223_ /*4386*/;
assign _4221_ = _4222_ | _4224_ /*4383*/;
assign _4230_ = D[28] ^ Q[11] /*4382*/;
assign _4227_ = _3887_ & _4230_ /*4378*/;
assign _4228_ = _3887_ ^ _4230_ /*4381*/;
assign _4229_ = _4221_ & _4228_ /*4379*/;
assign _4081_ = _4221_ ^ _4228_ /*4380*/;
assign _4226_ = _4227_ | _4229_ /*4377*/;
assign _4235_ = D[29] ^ Q[11] /*4376*/;
assign _4232_ = _3888_ & _4235_ /*4372*/;
assign _4233_ = _3888_ ^ _4235_ /*4375*/;
assign _4234_ = _4226_ & _4233_ /*4373*/;
assign _4082_ = _4226_ ^ _4233_ /*4374*/;
assign _4231_ = _4232_ | _4234_ /*4371*/;
assign _4240_ = D[30] ^ Q[11] /*4370*/;
assign _4237_ = _3889_ & _4240_ /*4366*/;
assign _4238_ = _3889_ ^ _4240_ /*4369*/;
assign _4239_ = _4231_ & _4238_ /*4367*/;
assign _4083_ = _4231_ ^ _4238_ /*4368*/;
assign _4236_ = _4237_ | _4239_ /*4365*/;
assign _4244_ = zeroWire ^ Q[11] /*4364*/;
assign _4241_ = _3890_ & _4244_ /*4360*/;
assign _4242_ = _3890_ ^ _4244_ /*4363*/;
assign _4243_ = _4236_ & _4242_ /*4361*/;
assign _4084_ = _4236_ ^ _4242_ /*4362*/;
assign Q[10] = _4241_ | _4243_ /*4359*/;
assign _4283_ = D[0] ^ Q[10] /*4165*/;
assign _4280_ = R_0[9] & _4283_ /*4161*/;
assign _4281_ = R_0[9] ^ _4283_ /*4164*/;
assign _4282_ = Q[10] & _4281_ /*4162*/;
assign _4246_ = Q[10] ^ _4281_ /*4163*/;
assign _4279_ = _4280_ | _4282_ /*4160*/;
assign _4288_ = D[1] ^ Q[10] /*4159*/;
assign _4285_ = _4053_ & _4288_ /*4155*/;
assign _4286_ = _4053_ ^ _4288_ /*4158*/;
assign _4287_ = _4279_ & _4286_ /*4156*/;
assign _4247_ = _4279_ ^ _4286_ /*4157*/;
assign _4284_ = _4285_ | _4287_ /*4154*/;
assign _4293_ = D[2] ^ Q[10] /*4153*/;
assign _4290_ = _4054_ & _4293_ /*4149*/;
assign _4291_ = _4054_ ^ _4293_ /*4152*/;
assign _4292_ = _4284_ & _4291_ /*4150*/;
assign _4248_ = _4284_ ^ _4291_ /*4151*/;
assign _4289_ = _4290_ | _4292_ /*4148*/;
assign _4298_ = D[3] ^ Q[10] /*4147*/;
assign _4295_ = _4055_ & _4298_ /*4143*/;
assign _4296_ = _4055_ ^ _4298_ /*4146*/;
assign _4297_ = _4289_ & _4296_ /*4144*/;
assign _4249_ = _4289_ ^ _4296_ /*4145*/;
assign _4294_ = _4295_ | _4297_ /*4142*/;
assign _4303_ = D[4] ^ Q[10] /*4141*/;
assign _4300_ = _4056_ & _4303_ /*4137*/;
assign _4301_ = _4056_ ^ _4303_ /*4140*/;
assign _4302_ = _4294_ & _4301_ /*4138*/;
assign _4250_ = _4294_ ^ _4301_ /*4139*/;
assign _4299_ = _4300_ | _4302_ /*4136*/;
assign _4308_ = D[5] ^ Q[10] /*4135*/;
assign _4305_ = _4057_ & _4308_ /*4131*/;
assign _4306_ = _4057_ ^ _4308_ /*4134*/;
assign _4307_ = _4299_ & _4306_ /*4132*/;
assign _4251_ = _4299_ ^ _4306_ /*4133*/;
assign _4304_ = _4305_ | _4307_ /*4130*/;
assign _4313_ = D[6] ^ Q[10] /*4129*/;
assign _4310_ = _4058_ & _4313_ /*4125*/;
assign _4311_ = _4058_ ^ _4313_ /*4128*/;
assign _4312_ = _4304_ & _4311_ /*4126*/;
assign _4252_ = _4304_ ^ _4311_ /*4127*/;
assign _4309_ = _4310_ | _4312_ /*4124*/;
assign _4318_ = D[7] ^ Q[10] /*4123*/;
assign _4315_ = _4059_ & _4318_ /*4119*/;
assign _4316_ = _4059_ ^ _4318_ /*4122*/;
assign _4317_ = _4309_ & _4316_ /*4120*/;
assign _4253_ = _4309_ ^ _4316_ /*4121*/;
assign _4314_ = _4315_ | _4317_ /*4118*/;
assign _4323_ = D[8] ^ Q[10] /*4117*/;
assign _4320_ = _4060_ & _4323_ /*4113*/;
assign _4321_ = _4060_ ^ _4323_ /*4116*/;
assign _4322_ = _4314_ & _4321_ /*4114*/;
assign _4254_ = _4314_ ^ _4321_ /*4115*/;
assign _4319_ = _4320_ | _4322_ /*4112*/;
assign _4328_ = D[9] ^ Q[10] /*4111*/;
assign _4325_ = _4061_ & _4328_ /*4107*/;
assign _4326_ = _4061_ ^ _4328_ /*4110*/;
assign _4327_ = _4319_ & _4326_ /*4108*/;
assign _4255_ = _4319_ ^ _4326_ /*4109*/;
assign _4324_ = _4325_ | _4327_ /*4106*/;
assign _4333_ = D[10] ^ Q[10] /*4105*/;
assign _4330_ = _4062_ & _4333_ /*4101*/;
assign _4331_ = _4062_ ^ _4333_ /*4104*/;
assign _4332_ = _4324_ & _4331_ /*4102*/;
assign _4256_ = _4324_ ^ _4331_ /*4103*/;
assign _4329_ = _4330_ | _4332_ /*4100*/;
assign _4338_ = D[11] ^ Q[10] /*4099*/;
assign _4335_ = _4063_ & _4338_ /*4095*/;
assign _4336_ = _4063_ ^ _4338_ /*4098*/;
assign _4337_ = _4329_ & _4336_ /*4096*/;
assign _4257_ = _4329_ ^ _4336_ /*4097*/;
assign _4334_ = _4335_ | _4337_ /*4094*/;
assign _4343_ = D[12] ^ Q[10] /*4093*/;
assign _4340_ = _4064_ & _4343_ /*4089*/;
assign _4341_ = _4064_ ^ _4343_ /*4092*/;
assign _4342_ = _4334_ & _4341_ /*4090*/;
assign _4258_ = _4334_ ^ _4341_ /*4091*/;
assign _4339_ = _4340_ | _4342_ /*4088*/;
assign _4348_ = D[13] ^ Q[10] /*4087*/;
assign _4345_ = _4065_ & _4348_ /*4083*/;
assign _4346_ = _4065_ ^ _4348_ /*4086*/;
assign _4347_ = _4339_ & _4346_ /*4084*/;
assign _4259_ = _4339_ ^ _4346_ /*4085*/;
assign _4344_ = _4345_ | _4347_ /*4082*/;
assign _4353_ = D[14] ^ Q[10] /*4081*/;
assign _4350_ = _4066_ & _4353_ /*4077*/;
assign _4351_ = _4066_ ^ _4353_ /*4080*/;
assign _4352_ = _4344_ & _4351_ /*4078*/;
assign _4260_ = _4344_ ^ _4351_ /*4079*/;
assign _4349_ = _4350_ | _4352_ /*4076*/;
assign _4358_ = D[15] ^ Q[10] /*4075*/;
assign _4355_ = _4067_ & _4358_ /*4071*/;
assign _4356_ = _4067_ ^ _4358_ /*4074*/;
assign _4357_ = _4349_ & _4356_ /*4072*/;
assign _4261_ = _4349_ ^ _4356_ /*4073*/;
assign _4354_ = _4355_ | _4357_ /*4070*/;
assign _4363_ = D[16] ^ Q[10] /*4069*/;
assign _4360_ = _4068_ & _4363_ /*4065*/;
assign _4361_ = _4068_ ^ _4363_ /*4068*/;
assign _4362_ = _4354_ & _4361_ /*4066*/;
assign _4262_ = _4354_ ^ _4361_ /*4067*/;
assign _4359_ = _4360_ | _4362_ /*4064*/;
assign _4368_ = D[17] ^ Q[10] /*4063*/;
assign _4365_ = _4069_ & _4368_ /*4059*/;
assign _4366_ = _4069_ ^ _4368_ /*4062*/;
assign _4367_ = _4359_ & _4366_ /*4060*/;
assign _4263_ = _4359_ ^ _4366_ /*4061*/;
assign _4364_ = _4365_ | _4367_ /*4058*/;
assign _4373_ = D[18] ^ Q[10] /*4057*/;
assign _4370_ = _4070_ & _4373_ /*4053*/;
assign _4371_ = _4070_ ^ _4373_ /*4056*/;
assign _4372_ = _4364_ & _4371_ /*4054*/;
assign _4264_ = _4364_ ^ _4371_ /*4055*/;
assign _4369_ = _4370_ | _4372_ /*4052*/;
assign _4378_ = D[19] ^ Q[10] /*4051*/;
assign _4375_ = _4071_ & _4378_ /*4047*/;
assign _4376_ = _4071_ ^ _4378_ /*4050*/;
assign _4377_ = _4369_ & _4376_ /*4048*/;
assign _4265_ = _4369_ ^ _4376_ /*4049*/;
assign _4374_ = _4375_ | _4377_ /*4046*/;
assign _4383_ = D[20] ^ Q[10] /*4045*/;
assign _4380_ = _4072_ & _4383_ /*4041*/;
assign _4381_ = _4072_ ^ _4383_ /*4044*/;
assign _4382_ = _4374_ & _4381_ /*4042*/;
assign _4266_ = _4374_ ^ _4381_ /*4043*/;
assign _4379_ = _4380_ | _4382_ /*4040*/;
assign _4388_ = D[21] ^ Q[10] /*4039*/;
assign _4385_ = _4073_ & _4388_ /*4035*/;
assign _4386_ = _4073_ ^ _4388_ /*4038*/;
assign _4387_ = _4379_ & _4386_ /*4036*/;
assign _4267_ = _4379_ ^ _4386_ /*4037*/;
assign _4384_ = _4385_ | _4387_ /*4034*/;
assign _4393_ = D[22] ^ Q[10] /*4033*/;
assign _4390_ = _4074_ & _4393_ /*4029*/;
assign _4391_ = _4074_ ^ _4393_ /*4032*/;
assign _4392_ = _4384_ & _4391_ /*4030*/;
assign _4268_ = _4384_ ^ _4391_ /*4031*/;
assign _4389_ = _4390_ | _4392_ /*4028*/;
assign _4398_ = D[23] ^ Q[10] /*4027*/;
assign _4395_ = _4075_ & _4398_ /*4023*/;
assign _4396_ = _4075_ ^ _4398_ /*4026*/;
assign _4397_ = _4389_ & _4396_ /*4024*/;
assign _4269_ = _4389_ ^ _4396_ /*4025*/;
assign _4394_ = _4395_ | _4397_ /*4022*/;
assign _4403_ = D[24] ^ Q[10] /*4021*/;
assign _4400_ = _4076_ & _4403_ /*4017*/;
assign _4401_ = _4076_ ^ _4403_ /*4020*/;
assign _4402_ = _4394_ & _4401_ /*4018*/;
assign _4270_ = _4394_ ^ _4401_ /*4019*/;
assign _4399_ = _4400_ | _4402_ /*4016*/;
assign _4408_ = D[25] ^ Q[10] /*4015*/;
assign _4405_ = _4077_ & _4408_ /*4011*/;
assign _4406_ = _4077_ ^ _4408_ /*4014*/;
assign _4407_ = _4399_ & _4406_ /*4012*/;
assign _4271_ = _4399_ ^ _4406_ /*4013*/;
assign _4404_ = _4405_ | _4407_ /*4010*/;
assign _4413_ = D[26] ^ Q[10] /*4009*/;
assign _4410_ = _4078_ & _4413_ /*4005*/;
assign _4411_ = _4078_ ^ _4413_ /*4008*/;
assign _4412_ = _4404_ & _4411_ /*4006*/;
assign _4272_ = _4404_ ^ _4411_ /*4007*/;
assign _4409_ = _4410_ | _4412_ /*4004*/;
assign _4418_ = D[27] ^ Q[10] /*4003*/;
assign _4415_ = _4079_ & _4418_ /*3999*/;
assign _4416_ = _4079_ ^ _4418_ /*4002*/;
assign _4417_ = _4409_ & _4416_ /*4000*/;
assign _4273_ = _4409_ ^ _4416_ /*4001*/;
assign _4414_ = _4415_ | _4417_ /*3998*/;
assign _4423_ = D[28] ^ Q[10] /*3997*/;
assign _4420_ = _4080_ & _4423_ /*3993*/;
assign _4421_ = _4080_ ^ _4423_ /*3996*/;
assign _4422_ = _4414_ & _4421_ /*3994*/;
assign _4274_ = _4414_ ^ _4421_ /*3995*/;
assign _4419_ = _4420_ | _4422_ /*3992*/;
assign _4428_ = D[29] ^ Q[10] /*3991*/;
assign _4425_ = _4081_ & _4428_ /*3987*/;
assign _4426_ = _4081_ ^ _4428_ /*3990*/;
assign _4427_ = _4419_ & _4426_ /*3988*/;
assign _4275_ = _4419_ ^ _4426_ /*3989*/;
assign _4424_ = _4425_ | _4427_ /*3986*/;
assign _4433_ = D[30] ^ Q[10] /*3985*/;
assign _4430_ = _4082_ & _4433_ /*3981*/;
assign _4431_ = _4082_ ^ _4433_ /*3984*/;
assign _4432_ = _4424_ & _4431_ /*3982*/;
assign _4276_ = _4424_ ^ _4431_ /*3983*/;
assign _4429_ = _4430_ | _4432_ /*3980*/;
assign _4437_ = zeroWire ^ Q[10] /*3979*/;
assign _4434_ = _4083_ & _4437_ /*3975*/;
assign _4435_ = _4083_ ^ _4437_ /*3978*/;
assign _4436_ = _4429_ & _4435_ /*3976*/;
assign _4277_ = _4429_ ^ _4435_ /*3977*/;
assign Q[9] = _4434_ | _4436_ /*3974*/;
assign _4476_ = D[0] ^ Q[9] /*3780*/;
assign _4473_ = R_0[8] & _4476_ /*3776*/;
assign _4474_ = R_0[8] ^ _4476_ /*3779*/;
assign _4475_ = Q[9] & _4474_ /*3777*/;
assign _4439_ = Q[9] ^ _4474_ /*3778*/;
assign _4472_ = _4473_ | _4475_ /*3775*/;
assign _4481_ = D[1] ^ Q[9] /*3774*/;
assign _4478_ = _4246_ & _4481_ /*3770*/;
assign _4479_ = _4246_ ^ _4481_ /*3773*/;
assign _4480_ = _4472_ & _4479_ /*3771*/;
assign _4440_ = _4472_ ^ _4479_ /*3772*/;
assign _4477_ = _4478_ | _4480_ /*3769*/;
assign _4486_ = D[2] ^ Q[9] /*3768*/;
assign _4483_ = _4247_ & _4486_ /*3764*/;
assign _4484_ = _4247_ ^ _4486_ /*3767*/;
assign _4485_ = _4477_ & _4484_ /*3765*/;
assign _4441_ = _4477_ ^ _4484_ /*3766*/;
assign _4482_ = _4483_ | _4485_ /*3763*/;
assign _4491_ = D[3] ^ Q[9] /*3762*/;
assign _4488_ = _4248_ & _4491_ /*3758*/;
assign _4489_ = _4248_ ^ _4491_ /*3761*/;
assign _4490_ = _4482_ & _4489_ /*3759*/;
assign _4442_ = _4482_ ^ _4489_ /*3760*/;
assign _4487_ = _4488_ | _4490_ /*3757*/;
assign _4496_ = D[4] ^ Q[9] /*3756*/;
assign _4493_ = _4249_ & _4496_ /*3752*/;
assign _4494_ = _4249_ ^ _4496_ /*3755*/;
assign _4495_ = _4487_ & _4494_ /*3753*/;
assign _4443_ = _4487_ ^ _4494_ /*3754*/;
assign _4492_ = _4493_ | _4495_ /*3751*/;
assign _4501_ = D[5] ^ Q[9] /*3750*/;
assign _4498_ = _4250_ & _4501_ /*3746*/;
assign _4499_ = _4250_ ^ _4501_ /*3749*/;
assign _4500_ = _4492_ & _4499_ /*3747*/;
assign _4444_ = _4492_ ^ _4499_ /*3748*/;
assign _4497_ = _4498_ | _4500_ /*3745*/;
assign _4506_ = D[6] ^ Q[9] /*3744*/;
assign _4503_ = _4251_ & _4506_ /*3740*/;
assign _4504_ = _4251_ ^ _4506_ /*3743*/;
assign _4505_ = _4497_ & _4504_ /*3741*/;
assign _4445_ = _4497_ ^ _4504_ /*3742*/;
assign _4502_ = _4503_ | _4505_ /*3739*/;
assign _4511_ = D[7] ^ Q[9] /*3738*/;
assign _4508_ = _4252_ & _4511_ /*3734*/;
assign _4509_ = _4252_ ^ _4511_ /*3737*/;
assign _4510_ = _4502_ & _4509_ /*3735*/;
assign _4446_ = _4502_ ^ _4509_ /*3736*/;
assign _4507_ = _4508_ | _4510_ /*3733*/;
assign _4516_ = D[8] ^ Q[9] /*3732*/;
assign _4513_ = _4253_ & _4516_ /*3728*/;
assign _4514_ = _4253_ ^ _4516_ /*3731*/;
assign _4515_ = _4507_ & _4514_ /*3729*/;
assign _4447_ = _4507_ ^ _4514_ /*3730*/;
assign _4512_ = _4513_ | _4515_ /*3727*/;
assign _4521_ = D[9] ^ Q[9] /*3726*/;
assign _4518_ = _4254_ & _4521_ /*3722*/;
assign _4519_ = _4254_ ^ _4521_ /*3725*/;
assign _4520_ = _4512_ & _4519_ /*3723*/;
assign _4448_ = _4512_ ^ _4519_ /*3724*/;
assign _4517_ = _4518_ | _4520_ /*3721*/;
assign _4526_ = D[10] ^ Q[9] /*3720*/;
assign _4523_ = _4255_ & _4526_ /*3716*/;
assign _4524_ = _4255_ ^ _4526_ /*3719*/;
assign _4525_ = _4517_ & _4524_ /*3717*/;
assign _4449_ = _4517_ ^ _4524_ /*3718*/;
assign _4522_ = _4523_ | _4525_ /*3715*/;
assign _4531_ = D[11] ^ Q[9] /*3714*/;
assign _4528_ = _4256_ & _4531_ /*3710*/;
assign _4529_ = _4256_ ^ _4531_ /*3713*/;
assign _4530_ = _4522_ & _4529_ /*3711*/;
assign _4450_ = _4522_ ^ _4529_ /*3712*/;
assign _4527_ = _4528_ | _4530_ /*3709*/;
assign _4536_ = D[12] ^ Q[9] /*3708*/;
assign _4533_ = _4257_ & _4536_ /*3704*/;
assign _4534_ = _4257_ ^ _4536_ /*3707*/;
assign _4535_ = _4527_ & _4534_ /*3705*/;
assign _4451_ = _4527_ ^ _4534_ /*3706*/;
assign _4532_ = _4533_ | _4535_ /*3703*/;
assign _4541_ = D[13] ^ Q[9] /*3702*/;
assign _4538_ = _4258_ & _4541_ /*3698*/;
assign _4539_ = _4258_ ^ _4541_ /*3701*/;
assign _4540_ = _4532_ & _4539_ /*3699*/;
assign _4452_ = _4532_ ^ _4539_ /*3700*/;
assign _4537_ = _4538_ | _4540_ /*3697*/;
assign _4546_ = D[14] ^ Q[9] /*3696*/;
assign _4543_ = _4259_ & _4546_ /*3692*/;
assign _4544_ = _4259_ ^ _4546_ /*3695*/;
assign _4545_ = _4537_ & _4544_ /*3693*/;
assign _4453_ = _4537_ ^ _4544_ /*3694*/;
assign _4542_ = _4543_ | _4545_ /*3691*/;
assign _4551_ = D[15] ^ Q[9] /*3690*/;
assign _4548_ = _4260_ & _4551_ /*3686*/;
assign _4549_ = _4260_ ^ _4551_ /*3689*/;
assign _4550_ = _4542_ & _4549_ /*3687*/;
assign _4454_ = _4542_ ^ _4549_ /*3688*/;
assign _4547_ = _4548_ | _4550_ /*3685*/;
assign _4556_ = D[16] ^ Q[9] /*3684*/;
assign _4553_ = _4261_ & _4556_ /*3680*/;
assign _4554_ = _4261_ ^ _4556_ /*3683*/;
assign _4555_ = _4547_ & _4554_ /*3681*/;
assign _4455_ = _4547_ ^ _4554_ /*3682*/;
assign _4552_ = _4553_ | _4555_ /*3679*/;
assign _4561_ = D[17] ^ Q[9] /*3678*/;
assign _4558_ = _4262_ & _4561_ /*3674*/;
assign _4559_ = _4262_ ^ _4561_ /*3677*/;
assign _4560_ = _4552_ & _4559_ /*3675*/;
assign _4456_ = _4552_ ^ _4559_ /*3676*/;
assign _4557_ = _4558_ | _4560_ /*3673*/;
assign _4566_ = D[18] ^ Q[9] /*3672*/;
assign _4563_ = _4263_ & _4566_ /*3668*/;
assign _4564_ = _4263_ ^ _4566_ /*3671*/;
assign _4565_ = _4557_ & _4564_ /*3669*/;
assign _4457_ = _4557_ ^ _4564_ /*3670*/;
assign _4562_ = _4563_ | _4565_ /*3667*/;
assign _4571_ = D[19] ^ Q[9] /*3666*/;
assign _4568_ = _4264_ & _4571_ /*3662*/;
assign _4569_ = _4264_ ^ _4571_ /*3665*/;
assign _4570_ = _4562_ & _4569_ /*3663*/;
assign _4458_ = _4562_ ^ _4569_ /*3664*/;
assign _4567_ = _4568_ | _4570_ /*3661*/;
assign _4576_ = D[20] ^ Q[9] /*3660*/;
assign _4573_ = _4265_ & _4576_ /*3656*/;
assign _4574_ = _4265_ ^ _4576_ /*3659*/;
assign _4575_ = _4567_ & _4574_ /*3657*/;
assign _4459_ = _4567_ ^ _4574_ /*3658*/;
assign _4572_ = _4573_ | _4575_ /*3655*/;
assign _4581_ = D[21] ^ Q[9] /*3654*/;
assign _4578_ = _4266_ & _4581_ /*3650*/;
assign _4579_ = _4266_ ^ _4581_ /*3653*/;
assign _4580_ = _4572_ & _4579_ /*3651*/;
assign _4460_ = _4572_ ^ _4579_ /*3652*/;
assign _4577_ = _4578_ | _4580_ /*3649*/;
assign _4586_ = D[22] ^ Q[9] /*3648*/;
assign _4583_ = _4267_ & _4586_ /*3644*/;
assign _4584_ = _4267_ ^ _4586_ /*3647*/;
assign _4585_ = _4577_ & _4584_ /*3645*/;
assign _4461_ = _4577_ ^ _4584_ /*3646*/;
assign _4582_ = _4583_ | _4585_ /*3643*/;
assign _4591_ = D[23] ^ Q[9] /*3642*/;
assign _4588_ = _4268_ & _4591_ /*3638*/;
assign _4589_ = _4268_ ^ _4591_ /*3641*/;
assign _4590_ = _4582_ & _4589_ /*3639*/;
assign _4462_ = _4582_ ^ _4589_ /*3640*/;
assign _4587_ = _4588_ | _4590_ /*3637*/;
assign _4596_ = D[24] ^ Q[9] /*3636*/;
assign _4593_ = _4269_ & _4596_ /*3632*/;
assign _4594_ = _4269_ ^ _4596_ /*3635*/;
assign _4595_ = _4587_ & _4594_ /*3633*/;
assign _4463_ = _4587_ ^ _4594_ /*3634*/;
assign _4592_ = _4593_ | _4595_ /*3631*/;
assign _4601_ = D[25] ^ Q[9] /*3630*/;
assign _4598_ = _4270_ & _4601_ /*3626*/;
assign _4599_ = _4270_ ^ _4601_ /*3629*/;
assign _4600_ = _4592_ & _4599_ /*3627*/;
assign _4464_ = _4592_ ^ _4599_ /*3628*/;
assign _4597_ = _4598_ | _4600_ /*3625*/;
assign _4606_ = D[26] ^ Q[9] /*3624*/;
assign _4603_ = _4271_ & _4606_ /*3620*/;
assign _4604_ = _4271_ ^ _4606_ /*3623*/;
assign _4605_ = _4597_ & _4604_ /*3621*/;
assign _4465_ = _4597_ ^ _4604_ /*3622*/;
assign _4602_ = _4603_ | _4605_ /*3619*/;
assign _4611_ = D[27] ^ Q[9] /*3618*/;
assign _4608_ = _4272_ & _4611_ /*3614*/;
assign _4609_ = _4272_ ^ _4611_ /*3617*/;
assign _4610_ = _4602_ & _4609_ /*3615*/;
assign _4466_ = _4602_ ^ _4609_ /*3616*/;
assign _4607_ = _4608_ | _4610_ /*3613*/;
assign _4616_ = D[28] ^ Q[9] /*3612*/;
assign _4613_ = _4273_ & _4616_ /*3608*/;
assign _4614_ = _4273_ ^ _4616_ /*3611*/;
assign _4615_ = _4607_ & _4614_ /*3609*/;
assign _4467_ = _4607_ ^ _4614_ /*3610*/;
assign _4612_ = _4613_ | _4615_ /*3607*/;
assign _4621_ = D[29] ^ Q[9] /*3606*/;
assign _4618_ = _4274_ & _4621_ /*3602*/;
assign _4619_ = _4274_ ^ _4621_ /*3605*/;
assign _4620_ = _4612_ & _4619_ /*3603*/;
assign _4468_ = _4612_ ^ _4619_ /*3604*/;
assign _4617_ = _4618_ | _4620_ /*3601*/;
assign _4626_ = D[30] ^ Q[9] /*3600*/;
assign _4623_ = _4275_ & _4626_ /*3596*/;
assign _4624_ = _4275_ ^ _4626_ /*3599*/;
assign _4625_ = _4617_ & _4624_ /*3597*/;
assign _4469_ = _4617_ ^ _4624_ /*3598*/;
assign _4622_ = _4623_ | _4625_ /*3595*/;
assign _4630_ = zeroWire ^ Q[9] /*3594*/;
assign _4627_ = _4276_ & _4630_ /*3590*/;
assign _4628_ = _4276_ ^ _4630_ /*3593*/;
assign _4629_ = _4622_ & _4628_ /*3591*/;
assign _4470_ = _4622_ ^ _4628_ /*3592*/;
assign Q[8] = _4627_ | _4629_ /*3589*/;
assign _4669_ = D[0] ^ Q[8] /*3395*/;
assign _4666_ = R_0[7] & _4669_ /*3391*/;
assign _4667_ = R_0[7] ^ _4669_ /*3394*/;
assign _4668_ = Q[8] & _4667_ /*3392*/;
assign _4632_ = Q[8] ^ _4667_ /*3393*/;
assign _4665_ = _4666_ | _4668_ /*3390*/;
assign _4674_ = D[1] ^ Q[8] /*3389*/;
assign _4671_ = _4439_ & _4674_ /*3385*/;
assign _4672_ = _4439_ ^ _4674_ /*3388*/;
assign _4673_ = _4665_ & _4672_ /*3386*/;
assign _4633_ = _4665_ ^ _4672_ /*3387*/;
assign _4670_ = _4671_ | _4673_ /*3384*/;
assign _4679_ = D[2] ^ Q[8] /*3383*/;
assign _4676_ = _4440_ & _4679_ /*3379*/;
assign _4677_ = _4440_ ^ _4679_ /*3382*/;
assign _4678_ = _4670_ & _4677_ /*3380*/;
assign _4634_ = _4670_ ^ _4677_ /*3381*/;
assign _4675_ = _4676_ | _4678_ /*3378*/;
assign _4684_ = D[3] ^ Q[8] /*3377*/;
assign _4681_ = _4441_ & _4684_ /*3373*/;
assign _4682_ = _4441_ ^ _4684_ /*3376*/;
assign _4683_ = _4675_ & _4682_ /*3374*/;
assign _4635_ = _4675_ ^ _4682_ /*3375*/;
assign _4680_ = _4681_ | _4683_ /*3372*/;
assign _4689_ = D[4] ^ Q[8] /*3371*/;
assign _4686_ = _4442_ & _4689_ /*3367*/;
assign _4687_ = _4442_ ^ _4689_ /*3370*/;
assign _4688_ = _4680_ & _4687_ /*3368*/;
assign _4636_ = _4680_ ^ _4687_ /*3369*/;
assign _4685_ = _4686_ | _4688_ /*3366*/;
assign _4694_ = D[5] ^ Q[8] /*3365*/;
assign _4691_ = _4443_ & _4694_ /*3361*/;
assign _4692_ = _4443_ ^ _4694_ /*3364*/;
assign _4693_ = _4685_ & _4692_ /*3362*/;
assign _4637_ = _4685_ ^ _4692_ /*3363*/;
assign _4690_ = _4691_ | _4693_ /*3360*/;
assign _4699_ = D[6] ^ Q[8] /*3359*/;
assign _4696_ = _4444_ & _4699_ /*3355*/;
assign _4697_ = _4444_ ^ _4699_ /*3358*/;
assign _4698_ = _4690_ & _4697_ /*3356*/;
assign _4638_ = _4690_ ^ _4697_ /*3357*/;
assign _4695_ = _4696_ | _4698_ /*3354*/;
assign _4704_ = D[7] ^ Q[8] /*3353*/;
assign _4701_ = _4445_ & _4704_ /*3349*/;
assign _4702_ = _4445_ ^ _4704_ /*3352*/;
assign _4703_ = _4695_ & _4702_ /*3350*/;
assign _4639_ = _4695_ ^ _4702_ /*3351*/;
assign _4700_ = _4701_ | _4703_ /*3348*/;
assign _4709_ = D[8] ^ Q[8] /*3347*/;
assign _4706_ = _4446_ & _4709_ /*3343*/;
assign _4707_ = _4446_ ^ _4709_ /*3346*/;
assign _4708_ = _4700_ & _4707_ /*3344*/;
assign _4640_ = _4700_ ^ _4707_ /*3345*/;
assign _4705_ = _4706_ | _4708_ /*3342*/;
assign _4714_ = D[9] ^ Q[8] /*3341*/;
assign _4711_ = _4447_ & _4714_ /*3337*/;
assign _4712_ = _4447_ ^ _4714_ /*3340*/;
assign _4713_ = _4705_ & _4712_ /*3338*/;
assign _4641_ = _4705_ ^ _4712_ /*3339*/;
assign _4710_ = _4711_ | _4713_ /*3336*/;
assign _4719_ = D[10] ^ Q[8] /*3335*/;
assign _4716_ = _4448_ & _4719_ /*3331*/;
assign _4717_ = _4448_ ^ _4719_ /*3334*/;
assign _4718_ = _4710_ & _4717_ /*3332*/;
assign _4642_ = _4710_ ^ _4717_ /*3333*/;
assign _4715_ = _4716_ | _4718_ /*3330*/;
assign _4724_ = D[11] ^ Q[8] /*3329*/;
assign _4721_ = _4449_ & _4724_ /*3325*/;
assign _4722_ = _4449_ ^ _4724_ /*3328*/;
assign _4723_ = _4715_ & _4722_ /*3326*/;
assign _4643_ = _4715_ ^ _4722_ /*3327*/;
assign _4720_ = _4721_ | _4723_ /*3324*/;
assign _4729_ = D[12] ^ Q[8] /*3323*/;
assign _4726_ = _4450_ & _4729_ /*3319*/;
assign _4727_ = _4450_ ^ _4729_ /*3322*/;
assign _4728_ = _4720_ & _4727_ /*3320*/;
assign _4644_ = _4720_ ^ _4727_ /*3321*/;
assign _4725_ = _4726_ | _4728_ /*3318*/;
assign _4734_ = D[13] ^ Q[8] /*3317*/;
assign _4731_ = _4451_ & _4734_ /*3313*/;
assign _4732_ = _4451_ ^ _4734_ /*3316*/;
assign _4733_ = _4725_ & _4732_ /*3314*/;
assign _4645_ = _4725_ ^ _4732_ /*3315*/;
assign _4730_ = _4731_ | _4733_ /*3312*/;
assign _4739_ = D[14] ^ Q[8] /*3311*/;
assign _4736_ = _4452_ & _4739_ /*3307*/;
assign _4737_ = _4452_ ^ _4739_ /*3310*/;
assign _4738_ = _4730_ & _4737_ /*3308*/;
assign _4646_ = _4730_ ^ _4737_ /*3309*/;
assign _4735_ = _4736_ | _4738_ /*3306*/;
assign _4744_ = D[15] ^ Q[8] /*3305*/;
assign _4741_ = _4453_ & _4744_ /*3301*/;
assign _4742_ = _4453_ ^ _4744_ /*3304*/;
assign _4743_ = _4735_ & _4742_ /*3302*/;
assign _4647_ = _4735_ ^ _4742_ /*3303*/;
assign _4740_ = _4741_ | _4743_ /*3300*/;
assign _4749_ = D[16] ^ Q[8] /*3299*/;
assign _4746_ = _4454_ & _4749_ /*3295*/;
assign _4747_ = _4454_ ^ _4749_ /*3298*/;
assign _4748_ = _4740_ & _4747_ /*3296*/;
assign _4648_ = _4740_ ^ _4747_ /*3297*/;
assign _4745_ = _4746_ | _4748_ /*3294*/;
assign _4754_ = D[17] ^ Q[8] /*3293*/;
assign _4751_ = _4455_ & _4754_ /*3289*/;
assign _4752_ = _4455_ ^ _4754_ /*3292*/;
assign _4753_ = _4745_ & _4752_ /*3290*/;
assign _4649_ = _4745_ ^ _4752_ /*3291*/;
assign _4750_ = _4751_ | _4753_ /*3288*/;
assign _4759_ = D[18] ^ Q[8] /*3287*/;
assign _4756_ = _4456_ & _4759_ /*3283*/;
assign _4757_ = _4456_ ^ _4759_ /*3286*/;
assign _4758_ = _4750_ & _4757_ /*3284*/;
assign _4650_ = _4750_ ^ _4757_ /*3285*/;
assign _4755_ = _4756_ | _4758_ /*3282*/;
assign _4764_ = D[19] ^ Q[8] /*3281*/;
assign _4761_ = _4457_ & _4764_ /*3277*/;
assign _4762_ = _4457_ ^ _4764_ /*3280*/;
assign _4763_ = _4755_ & _4762_ /*3278*/;
assign _4651_ = _4755_ ^ _4762_ /*3279*/;
assign _4760_ = _4761_ | _4763_ /*3276*/;
assign _4769_ = D[20] ^ Q[8] /*3275*/;
assign _4766_ = _4458_ & _4769_ /*3271*/;
assign _4767_ = _4458_ ^ _4769_ /*3274*/;
assign _4768_ = _4760_ & _4767_ /*3272*/;
assign _4652_ = _4760_ ^ _4767_ /*3273*/;
assign _4765_ = _4766_ | _4768_ /*3270*/;
assign _4774_ = D[21] ^ Q[8] /*3269*/;
assign _4771_ = _4459_ & _4774_ /*3265*/;
assign _4772_ = _4459_ ^ _4774_ /*3268*/;
assign _4773_ = _4765_ & _4772_ /*3266*/;
assign _4653_ = _4765_ ^ _4772_ /*3267*/;
assign _4770_ = _4771_ | _4773_ /*3264*/;
assign _4779_ = D[22] ^ Q[8] /*3263*/;
assign _4776_ = _4460_ & _4779_ /*3259*/;
assign _4777_ = _4460_ ^ _4779_ /*3262*/;
assign _4778_ = _4770_ & _4777_ /*3260*/;
assign _4654_ = _4770_ ^ _4777_ /*3261*/;
assign _4775_ = _4776_ | _4778_ /*3258*/;
assign _4784_ = D[23] ^ Q[8] /*3257*/;
assign _4781_ = _4461_ & _4784_ /*3253*/;
assign _4782_ = _4461_ ^ _4784_ /*3256*/;
assign _4783_ = _4775_ & _4782_ /*3254*/;
assign _4655_ = _4775_ ^ _4782_ /*3255*/;
assign _4780_ = _4781_ | _4783_ /*3252*/;
assign _4789_ = D[24] ^ Q[8] /*3251*/;
assign _4786_ = _4462_ & _4789_ /*3247*/;
assign _4787_ = _4462_ ^ _4789_ /*3250*/;
assign _4788_ = _4780_ & _4787_ /*3248*/;
assign _4656_ = _4780_ ^ _4787_ /*3249*/;
assign _4785_ = _4786_ | _4788_ /*3246*/;
assign _4794_ = D[25] ^ Q[8] /*3245*/;
assign _4791_ = _4463_ & _4794_ /*3241*/;
assign _4792_ = _4463_ ^ _4794_ /*3244*/;
assign _4793_ = _4785_ & _4792_ /*3242*/;
assign _4657_ = _4785_ ^ _4792_ /*3243*/;
assign _4790_ = _4791_ | _4793_ /*3240*/;
assign _4799_ = D[26] ^ Q[8] /*3239*/;
assign _4796_ = _4464_ & _4799_ /*3235*/;
assign _4797_ = _4464_ ^ _4799_ /*3238*/;
assign _4798_ = _4790_ & _4797_ /*3236*/;
assign _4658_ = _4790_ ^ _4797_ /*3237*/;
assign _4795_ = _4796_ | _4798_ /*3234*/;
assign _4804_ = D[27] ^ Q[8] /*3233*/;
assign _4801_ = _4465_ & _4804_ /*3229*/;
assign _4802_ = _4465_ ^ _4804_ /*3232*/;
assign _4803_ = _4795_ & _4802_ /*3230*/;
assign _4659_ = _4795_ ^ _4802_ /*3231*/;
assign _4800_ = _4801_ | _4803_ /*3228*/;
assign _4809_ = D[28] ^ Q[8] /*3227*/;
assign _4806_ = _4466_ & _4809_ /*3223*/;
assign _4807_ = _4466_ ^ _4809_ /*3226*/;
assign _4808_ = _4800_ & _4807_ /*3224*/;
assign _4660_ = _4800_ ^ _4807_ /*3225*/;
assign _4805_ = _4806_ | _4808_ /*3222*/;
assign _4814_ = D[29] ^ Q[8] /*3221*/;
assign _4811_ = _4467_ & _4814_ /*3217*/;
assign _4812_ = _4467_ ^ _4814_ /*3220*/;
assign _4813_ = _4805_ & _4812_ /*3218*/;
assign _4661_ = _4805_ ^ _4812_ /*3219*/;
assign _4810_ = _4811_ | _4813_ /*3216*/;
assign _4819_ = D[30] ^ Q[8] /*3215*/;
assign _4816_ = _4468_ & _4819_ /*3211*/;
assign _4817_ = _4468_ ^ _4819_ /*3214*/;
assign _4818_ = _4810_ & _4817_ /*3212*/;
assign _4662_ = _4810_ ^ _4817_ /*3213*/;
assign _4815_ = _4816_ | _4818_ /*3210*/;
assign _4823_ = zeroWire ^ Q[8] /*3209*/;
assign _4820_ = _4469_ & _4823_ /*3205*/;
assign _4821_ = _4469_ ^ _4823_ /*3208*/;
assign _4822_ = _4815_ & _4821_ /*3206*/;
assign _4663_ = _4815_ ^ _4821_ /*3207*/;
assign Q[7] = _4820_ | _4822_ /*3204*/;
assign _4862_ = D[0] ^ Q[7] /*3010*/;
assign _4859_ = R_0[6] & _4862_ /*3006*/;
assign _4860_ = R_0[6] ^ _4862_ /*3009*/;
assign _4861_ = Q[7] & _4860_ /*3007*/;
assign _4825_ = Q[7] ^ _4860_ /*3008*/;
assign _4858_ = _4859_ | _4861_ /*3005*/;
assign _4867_ = D[1] ^ Q[7] /*3004*/;
assign _4864_ = _4632_ & _4867_ /*3000*/;
assign _4865_ = _4632_ ^ _4867_ /*3003*/;
assign _4866_ = _4858_ & _4865_ /*3001*/;
assign _4826_ = _4858_ ^ _4865_ /*3002*/;
assign _4863_ = _4864_ | _4866_ /*2999*/;
assign _4872_ = D[2] ^ Q[7] /*2998*/;
assign _4869_ = _4633_ & _4872_ /*2994*/;
assign _4870_ = _4633_ ^ _4872_ /*2997*/;
assign _4871_ = _4863_ & _4870_ /*2995*/;
assign _4827_ = _4863_ ^ _4870_ /*2996*/;
assign _4868_ = _4869_ | _4871_ /*2993*/;
assign _4877_ = D[3] ^ Q[7] /*2992*/;
assign _4874_ = _4634_ & _4877_ /*2988*/;
assign _4875_ = _4634_ ^ _4877_ /*2991*/;
assign _4876_ = _4868_ & _4875_ /*2989*/;
assign _4828_ = _4868_ ^ _4875_ /*2990*/;
assign _4873_ = _4874_ | _4876_ /*2987*/;
assign _4882_ = D[4] ^ Q[7] /*2986*/;
assign _4879_ = _4635_ & _4882_ /*2982*/;
assign _4880_ = _4635_ ^ _4882_ /*2985*/;
assign _4881_ = _4873_ & _4880_ /*2983*/;
assign _4829_ = _4873_ ^ _4880_ /*2984*/;
assign _4878_ = _4879_ | _4881_ /*2981*/;
assign _4887_ = D[5] ^ Q[7] /*2980*/;
assign _4884_ = _4636_ & _4887_ /*2976*/;
assign _4885_ = _4636_ ^ _4887_ /*2979*/;
assign _4886_ = _4878_ & _4885_ /*2977*/;
assign _4830_ = _4878_ ^ _4885_ /*2978*/;
assign _4883_ = _4884_ | _4886_ /*2975*/;
assign _4892_ = D[6] ^ Q[7] /*2974*/;
assign _4889_ = _4637_ & _4892_ /*2970*/;
assign _4890_ = _4637_ ^ _4892_ /*2973*/;
assign _4891_ = _4883_ & _4890_ /*2971*/;
assign _4831_ = _4883_ ^ _4890_ /*2972*/;
assign _4888_ = _4889_ | _4891_ /*2969*/;
assign _4897_ = D[7] ^ Q[7] /*2968*/;
assign _4894_ = _4638_ & _4897_ /*2964*/;
assign _4895_ = _4638_ ^ _4897_ /*2967*/;
assign _4896_ = _4888_ & _4895_ /*2965*/;
assign _4832_ = _4888_ ^ _4895_ /*2966*/;
assign _4893_ = _4894_ | _4896_ /*2963*/;
assign _4902_ = D[8] ^ Q[7] /*2962*/;
assign _4899_ = _4639_ & _4902_ /*2958*/;
assign _4900_ = _4639_ ^ _4902_ /*2961*/;
assign _4901_ = _4893_ & _4900_ /*2959*/;
assign _4833_ = _4893_ ^ _4900_ /*2960*/;
assign _4898_ = _4899_ | _4901_ /*2957*/;
assign _4907_ = D[9] ^ Q[7] /*2956*/;
assign _4904_ = _4640_ & _4907_ /*2952*/;
assign _4905_ = _4640_ ^ _4907_ /*2955*/;
assign _4906_ = _4898_ & _4905_ /*2953*/;
assign _4834_ = _4898_ ^ _4905_ /*2954*/;
assign _4903_ = _4904_ | _4906_ /*2951*/;
assign _4912_ = D[10] ^ Q[7] /*2950*/;
assign _4909_ = _4641_ & _4912_ /*2946*/;
assign _4910_ = _4641_ ^ _4912_ /*2949*/;
assign _4911_ = _4903_ & _4910_ /*2947*/;
assign _4835_ = _4903_ ^ _4910_ /*2948*/;
assign _4908_ = _4909_ | _4911_ /*2945*/;
assign _4917_ = D[11] ^ Q[7] /*2944*/;
assign _4914_ = _4642_ & _4917_ /*2940*/;
assign _4915_ = _4642_ ^ _4917_ /*2943*/;
assign _4916_ = _4908_ & _4915_ /*2941*/;
assign _4836_ = _4908_ ^ _4915_ /*2942*/;
assign _4913_ = _4914_ | _4916_ /*2939*/;
assign _4922_ = D[12] ^ Q[7] /*2938*/;
assign _4919_ = _4643_ & _4922_ /*2934*/;
assign _4920_ = _4643_ ^ _4922_ /*2937*/;
assign _4921_ = _4913_ & _4920_ /*2935*/;
assign _4837_ = _4913_ ^ _4920_ /*2936*/;
assign _4918_ = _4919_ | _4921_ /*2933*/;
assign _4927_ = D[13] ^ Q[7] /*2932*/;
assign _4924_ = _4644_ & _4927_ /*2928*/;
assign _4925_ = _4644_ ^ _4927_ /*2931*/;
assign _4926_ = _4918_ & _4925_ /*2929*/;
assign _4838_ = _4918_ ^ _4925_ /*2930*/;
assign _4923_ = _4924_ | _4926_ /*2927*/;
assign _4932_ = D[14] ^ Q[7] /*2926*/;
assign _4929_ = _4645_ & _4932_ /*2922*/;
assign _4930_ = _4645_ ^ _4932_ /*2925*/;
assign _4931_ = _4923_ & _4930_ /*2923*/;
assign _4839_ = _4923_ ^ _4930_ /*2924*/;
assign _4928_ = _4929_ | _4931_ /*2921*/;
assign _4937_ = D[15] ^ Q[7] /*2920*/;
assign _4934_ = _4646_ & _4937_ /*2916*/;
assign _4935_ = _4646_ ^ _4937_ /*2919*/;
assign _4936_ = _4928_ & _4935_ /*2917*/;
assign _4840_ = _4928_ ^ _4935_ /*2918*/;
assign _4933_ = _4934_ | _4936_ /*2915*/;
assign _4942_ = D[16] ^ Q[7] /*2914*/;
assign _4939_ = _4647_ & _4942_ /*2910*/;
assign _4940_ = _4647_ ^ _4942_ /*2913*/;
assign _4941_ = _4933_ & _4940_ /*2911*/;
assign _4841_ = _4933_ ^ _4940_ /*2912*/;
assign _4938_ = _4939_ | _4941_ /*2909*/;
assign _4947_ = D[17] ^ Q[7] /*2908*/;
assign _4944_ = _4648_ & _4947_ /*2904*/;
assign _4945_ = _4648_ ^ _4947_ /*2907*/;
assign _4946_ = _4938_ & _4945_ /*2905*/;
assign _4842_ = _4938_ ^ _4945_ /*2906*/;
assign _4943_ = _4944_ | _4946_ /*2903*/;
assign _4952_ = D[18] ^ Q[7] /*2902*/;
assign _4949_ = _4649_ & _4952_ /*2898*/;
assign _4950_ = _4649_ ^ _4952_ /*2901*/;
assign _4951_ = _4943_ & _4950_ /*2899*/;
assign _4843_ = _4943_ ^ _4950_ /*2900*/;
assign _4948_ = _4949_ | _4951_ /*2897*/;
assign _4957_ = D[19] ^ Q[7] /*2896*/;
assign _4954_ = _4650_ & _4957_ /*2892*/;
assign _4955_ = _4650_ ^ _4957_ /*2895*/;
assign _4956_ = _4948_ & _4955_ /*2893*/;
assign _4844_ = _4948_ ^ _4955_ /*2894*/;
assign _4953_ = _4954_ | _4956_ /*2891*/;
assign _4962_ = D[20] ^ Q[7] /*2890*/;
assign _4959_ = _4651_ & _4962_ /*2886*/;
assign _4960_ = _4651_ ^ _4962_ /*2889*/;
assign _4961_ = _4953_ & _4960_ /*2887*/;
assign _4845_ = _4953_ ^ _4960_ /*2888*/;
assign _4958_ = _4959_ | _4961_ /*2885*/;
assign _4967_ = D[21] ^ Q[7] /*2884*/;
assign _4964_ = _4652_ & _4967_ /*2880*/;
assign _4965_ = _4652_ ^ _4967_ /*2883*/;
assign _4966_ = _4958_ & _4965_ /*2881*/;
assign _4846_ = _4958_ ^ _4965_ /*2882*/;
assign _4963_ = _4964_ | _4966_ /*2879*/;
assign _4972_ = D[22] ^ Q[7] /*2878*/;
assign _4969_ = _4653_ & _4972_ /*2874*/;
assign _4970_ = _4653_ ^ _4972_ /*2877*/;
assign _4971_ = _4963_ & _4970_ /*2875*/;
assign _4847_ = _4963_ ^ _4970_ /*2876*/;
assign _4968_ = _4969_ | _4971_ /*2873*/;
assign _4977_ = D[23] ^ Q[7] /*2872*/;
assign _4974_ = _4654_ & _4977_ /*2868*/;
assign _4975_ = _4654_ ^ _4977_ /*2871*/;
assign _4976_ = _4968_ & _4975_ /*2869*/;
assign _4848_ = _4968_ ^ _4975_ /*2870*/;
assign _4973_ = _4974_ | _4976_ /*2867*/;
assign _4982_ = D[24] ^ Q[7] /*2866*/;
assign _4979_ = _4655_ & _4982_ /*2862*/;
assign _4980_ = _4655_ ^ _4982_ /*2865*/;
assign _4981_ = _4973_ & _4980_ /*2863*/;
assign _4849_ = _4973_ ^ _4980_ /*2864*/;
assign _4978_ = _4979_ | _4981_ /*2861*/;
assign _4987_ = D[25] ^ Q[7] /*2860*/;
assign _4984_ = _4656_ & _4987_ /*2856*/;
assign _4985_ = _4656_ ^ _4987_ /*2859*/;
assign _4986_ = _4978_ & _4985_ /*2857*/;
assign _4850_ = _4978_ ^ _4985_ /*2858*/;
assign _4983_ = _4984_ | _4986_ /*2855*/;
assign _4992_ = D[26] ^ Q[7] /*2854*/;
assign _4989_ = _4657_ & _4992_ /*2850*/;
assign _4990_ = _4657_ ^ _4992_ /*2853*/;
assign _4991_ = _4983_ & _4990_ /*2851*/;
assign _4851_ = _4983_ ^ _4990_ /*2852*/;
assign _4988_ = _4989_ | _4991_ /*2849*/;
assign _4997_ = D[27] ^ Q[7] /*2848*/;
assign _4994_ = _4658_ & _4997_ /*2844*/;
assign _4995_ = _4658_ ^ _4997_ /*2847*/;
assign _4996_ = _4988_ & _4995_ /*2845*/;
assign _4852_ = _4988_ ^ _4995_ /*2846*/;
assign _4993_ = _4994_ | _4996_ /*2843*/;
assign _5002_ = D[28] ^ Q[7] /*2842*/;
assign _4999_ = _4659_ & _5002_ /*2838*/;
assign _5000_ = _4659_ ^ _5002_ /*2841*/;
assign _5001_ = _4993_ & _5000_ /*2839*/;
assign _4853_ = _4993_ ^ _5000_ /*2840*/;
assign _4998_ = _4999_ | _5001_ /*2837*/;
assign _5007_ = D[29] ^ Q[7] /*2836*/;
assign _5004_ = _4660_ & _5007_ /*2832*/;
assign _5005_ = _4660_ ^ _5007_ /*2835*/;
assign _5006_ = _4998_ & _5005_ /*2833*/;
assign _4854_ = _4998_ ^ _5005_ /*2834*/;
assign _5003_ = _5004_ | _5006_ /*2831*/;
assign _5012_ = D[30] ^ Q[7] /*2830*/;
assign _5009_ = _4661_ & _5012_ /*2826*/;
assign _5010_ = _4661_ ^ _5012_ /*2829*/;
assign _5011_ = _5003_ & _5010_ /*2827*/;
assign _4855_ = _5003_ ^ _5010_ /*2828*/;
assign _5008_ = _5009_ | _5011_ /*2825*/;
assign _5016_ = zeroWire ^ Q[7] /*2824*/;
assign _5013_ = _4662_ & _5016_ /*2820*/;
assign _5014_ = _4662_ ^ _5016_ /*2823*/;
assign _5015_ = _5008_ & _5014_ /*2821*/;
assign _4856_ = _5008_ ^ _5014_ /*2822*/;
assign Q[6] = _5013_ | _5015_ /*2819*/;
assign _5055_ = D[0] ^ Q[6] /*2625*/;
assign _5052_ = R_0[5] & _5055_ /*2621*/;
assign _5053_ = R_0[5] ^ _5055_ /*2624*/;
assign _5054_ = Q[6] & _5053_ /*2622*/;
assign _5018_ = Q[6] ^ _5053_ /*2623*/;
assign _5051_ = _5052_ | _5054_ /*2620*/;
assign _5060_ = D[1] ^ Q[6] /*2619*/;
assign _5057_ = _4825_ & _5060_ /*2615*/;
assign _5058_ = _4825_ ^ _5060_ /*2618*/;
assign _5059_ = _5051_ & _5058_ /*2616*/;
assign _5019_ = _5051_ ^ _5058_ /*2617*/;
assign _5056_ = _5057_ | _5059_ /*2614*/;
assign _5065_ = D[2] ^ Q[6] /*2613*/;
assign _5062_ = _4826_ & _5065_ /*2609*/;
assign _5063_ = _4826_ ^ _5065_ /*2612*/;
assign _5064_ = _5056_ & _5063_ /*2610*/;
assign _5020_ = _5056_ ^ _5063_ /*2611*/;
assign _5061_ = _5062_ | _5064_ /*2608*/;
assign _5070_ = D[3] ^ Q[6] /*2607*/;
assign _5067_ = _4827_ & _5070_ /*2603*/;
assign _5068_ = _4827_ ^ _5070_ /*2606*/;
assign _5069_ = _5061_ & _5068_ /*2604*/;
assign _5021_ = _5061_ ^ _5068_ /*2605*/;
assign _5066_ = _5067_ | _5069_ /*2602*/;
assign _5075_ = D[4] ^ Q[6] /*2601*/;
assign _5072_ = _4828_ & _5075_ /*2597*/;
assign _5073_ = _4828_ ^ _5075_ /*2600*/;
assign _5074_ = _5066_ & _5073_ /*2598*/;
assign _5022_ = _5066_ ^ _5073_ /*2599*/;
assign _5071_ = _5072_ | _5074_ /*2596*/;
assign _5080_ = D[5] ^ Q[6] /*2595*/;
assign _5077_ = _4829_ & _5080_ /*2591*/;
assign _5078_ = _4829_ ^ _5080_ /*2594*/;
assign _5079_ = _5071_ & _5078_ /*2592*/;
assign _5023_ = _5071_ ^ _5078_ /*2593*/;
assign _5076_ = _5077_ | _5079_ /*2590*/;
assign _5085_ = D[6] ^ Q[6] /*2589*/;
assign _5082_ = _4830_ & _5085_ /*2585*/;
assign _5083_ = _4830_ ^ _5085_ /*2588*/;
assign _5084_ = _5076_ & _5083_ /*2586*/;
assign _5024_ = _5076_ ^ _5083_ /*2587*/;
assign _5081_ = _5082_ | _5084_ /*2584*/;
assign _5090_ = D[7] ^ Q[6] /*2583*/;
assign _5087_ = _4831_ & _5090_ /*2579*/;
assign _5088_ = _4831_ ^ _5090_ /*2582*/;
assign _5089_ = _5081_ & _5088_ /*2580*/;
assign _5025_ = _5081_ ^ _5088_ /*2581*/;
assign _5086_ = _5087_ | _5089_ /*2578*/;
assign _5095_ = D[8] ^ Q[6] /*2577*/;
assign _5092_ = _4832_ & _5095_ /*2573*/;
assign _5093_ = _4832_ ^ _5095_ /*2576*/;
assign _5094_ = _5086_ & _5093_ /*2574*/;
assign _5026_ = _5086_ ^ _5093_ /*2575*/;
assign _5091_ = _5092_ | _5094_ /*2572*/;
assign _5100_ = D[9] ^ Q[6] /*2571*/;
assign _5097_ = _4833_ & _5100_ /*2567*/;
assign _5098_ = _4833_ ^ _5100_ /*2570*/;
assign _5099_ = _5091_ & _5098_ /*2568*/;
assign _5027_ = _5091_ ^ _5098_ /*2569*/;
assign _5096_ = _5097_ | _5099_ /*2566*/;
assign _5105_ = D[10] ^ Q[6] /*2565*/;
assign _5102_ = _4834_ & _5105_ /*2561*/;
assign _5103_ = _4834_ ^ _5105_ /*2564*/;
assign _5104_ = _5096_ & _5103_ /*2562*/;
assign _5028_ = _5096_ ^ _5103_ /*2563*/;
assign _5101_ = _5102_ | _5104_ /*2560*/;
assign _5110_ = D[11] ^ Q[6] /*2559*/;
assign _5107_ = _4835_ & _5110_ /*2555*/;
assign _5108_ = _4835_ ^ _5110_ /*2558*/;
assign _5109_ = _5101_ & _5108_ /*2556*/;
assign _5029_ = _5101_ ^ _5108_ /*2557*/;
assign _5106_ = _5107_ | _5109_ /*2554*/;
assign _5115_ = D[12] ^ Q[6] /*2553*/;
assign _5112_ = _4836_ & _5115_ /*2549*/;
assign _5113_ = _4836_ ^ _5115_ /*2552*/;
assign _5114_ = _5106_ & _5113_ /*2550*/;
assign _5030_ = _5106_ ^ _5113_ /*2551*/;
assign _5111_ = _5112_ | _5114_ /*2548*/;
assign _5120_ = D[13] ^ Q[6] /*2547*/;
assign _5117_ = _4837_ & _5120_ /*2543*/;
assign _5118_ = _4837_ ^ _5120_ /*2546*/;
assign _5119_ = _5111_ & _5118_ /*2544*/;
assign _5031_ = _5111_ ^ _5118_ /*2545*/;
assign _5116_ = _5117_ | _5119_ /*2542*/;
assign _5125_ = D[14] ^ Q[6] /*2541*/;
assign _5122_ = _4838_ & _5125_ /*2537*/;
assign _5123_ = _4838_ ^ _5125_ /*2540*/;
assign _5124_ = _5116_ & _5123_ /*2538*/;
assign _5032_ = _5116_ ^ _5123_ /*2539*/;
assign _5121_ = _5122_ | _5124_ /*2536*/;
assign _5130_ = D[15] ^ Q[6] /*2535*/;
assign _5127_ = _4839_ & _5130_ /*2531*/;
assign _5128_ = _4839_ ^ _5130_ /*2534*/;
assign _5129_ = _5121_ & _5128_ /*2532*/;
assign _5033_ = _5121_ ^ _5128_ /*2533*/;
assign _5126_ = _5127_ | _5129_ /*2530*/;
assign _5135_ = D[16] ^ Q[6] /*2529*/;
assign _5132_ = _4840_ & _5135_ /*2525*/;
assign _5133_ = _4840_ ^ _5135_ /*2528*/;
assign _5134_ = _5126_ & _5133_ /*2526*/;
assign _5034_ = _5126_ ^ _5133_ /*2527*/;
assign _5131_ = _5132_ | _5134_ /*2524*/;
assign _5140_ = D[17] ^ Q[6] /*2523*/;
assign _5137_ = _4841_ & _5140_ /*2519*/;
assign _5138_ = _4841_ ^ _5140_ /*2522*/;
assign _5139_ = _5131_ & _5138_ /*2520*/;
assign _5035_ = _5131_ ^ _5138_ /*2521*/;
assign _5136_ = _5137_ | _5139_ /*2518*/;
assign _5145_ = D[18] ^ Q[6] /*2517*/;
assign _5142_ = _4842_ & _5145_ /*2513*/;
assign _5143_ = _4842_ ^ _5145_ /*2516*/;
assign _5144_ = _5136_ & _5143_ /*2514*/;
assign _5036_ = _5136_ ^ _5143_ /*2515*/;
assign _5141_ = _5142_ | _5144_ /*2512*/;
assign _5150_ = D[19] ^ Q[6] /*2511*/;
assign _5147_ = _4843_ & _5150_ /*2507*/;
assign _5148_ = _4843_ ^ _5150_ /*2510*/;
assign _5149_ = _5141_ & _5148_ /*2508*/;
assign _5037_ = _5141_ ^ _5148_ /*2509*/;
assign _5146_ = _5147_ | _5149_ /*2506*/;
assign _5155_ = D[20] ^ Q[6] /*2505*/;
assign _5152_ = _4844_ & _5155_ /*2501*/;
assign _5153_ = _4844_ ^ _5155_ /*2504*/;
assign _5154_ = _5146_ & _5153_ /*2502*/;
assign _5038_ = _5146_ ^ _5153_ /*2503*/;
assign _5151_ = _5152_ | _5154_ /*2500*/;
assign _5160_ = D[21] ^ Q[6] /*2499*/;
assign _5157_ = _4845_ & _5160_ /*2495*/;
assign _5158_ = _4845_ ^ _5160_ /*2498*/;
assign _5159_ = _5151_ & _5158_ /*2496*/;
assign _5039_ = _5151_ ^ _5158_ /*2497*/;
assign _5156_ = _5157_ | _5159_ /*2494*/;
assign _5165_ = D[22] ^ Q[6] /*2493*/;
assign _5162_ = _4846_ & _5165_ /*2489*/;
assign _5163_ = _4846_ ^ _5165_ /*2492*/;
assign _5164_ = _5156_ & _5163_ /*2490*/;
assign _5040_ = _5156_ ^ _5163_ /*2491*/;
assign _5161_ = _5162_ | _5164_ /*2488*/;
assign _5170_ = D[23] ^ Q[6] /*2487*/;
assign _5167_ = _4847_ & _5170_ /*2483*/;
assign _5168_ = _4847_ ^ _5170_ /*2486*/;
assign _5169_ = _5161_ & _5168_ /*2484*/;
assign _5041_ = _5161_ ^ _5168_ /*2485*/;
assign _5166_ = _5167_ | _5169_ /*2482*/;
assign _5175_ = D[24] ^ Q[6] /*2481*/;
assign _5172_ = _4848_ & _5175_ /*2477*/;
assign _5173_ = _4848_ ^ _5175_ /*2480*/;
assign _5174_ = _5166_ & _5173_ /*2478*/;
assign _5042_ = _5166_ ^ _5173_ /*2479*/;
assign _5171_ = _5172_ | _5174_ /*2476*/;
assign _5180_ = D[25] ^ Q[6] /*2475*/;
assign _5177_ = _4849_ & _5180_ /*2471*/;
assign _5178_ = _4849_ ^ _5180_ /*2474*/;
assign _5179_ = _5171_ & _5178_ /*2472*/;
assign _5043_ = _5171_ ^ _5178_ /*2473*/;
assign _5176_ = _5177_ | _5179_ /*2470*/;
assign _5185_ = D[26] ^ Q[6] /*2469*/;
assign _5182_ = _4850_ & _5185_ /*2465*/;
assign _5183_ = _4850_ ^ _5185_ /*2468*/;
assign _5184_ = _5176_ & _5183_ /*2466*/;
assign _5044_ = _5176_ ^ _5183_ /*2467*/;
assign _5181_ = _5182_ | _5184_ /*2464*/;
assign _5190_ = D[27] ^ Q[6] /*2463*/;
assign _5187_ = _4851_ & _5190_ /*2459*/;
assign _5188_ = _4851_ ^ _5190_ /*2462*/;
assign _5189_ = _5181_ & _5188_ /*2460*/;
assign _5045_ = _5181_ ^ _5188_ /*2461*/;
assign _5186_ = _5187_ | _5189_ /*2458*/;
assign _5195_ = D[28] ^ Q[6] /*2457*/;
assign _5192_ = _4852_ & _5195_ /*2453*/;
assign _5193_ = _4852_ ^ _5195_ /*2456*/;
assign _5194_ = _5186_ & _5193_ /*2454*/;
assign _5046_ = _5186_ ^ _5193_ /*2455*/;
assign _5191_ = _5192_ | _5194_ /*2452*/;
assign _5200_ = D[29] ^ Q[6] /*2451*/;
assign _5197_ = _4853_ & _5200_ /*2447*/;
assign _5198_ = _4853_ ^ _5200_ /*2450*/;
assign _5199_ = _5191_ & _5198_ /*2448*/;
assign _5047_ = _5191_ ^ _5198_ /*2449*/;
assign _5196_ = _5197_ | _5199_ /*2446*/;
assign _5205_ = D[30] ^ Q[6] /*2445*/;
assign _5202_ = _4854_ & _5205_ /*2441*/;
assign _5203_ = _4854_ ^ _5205_ /*2444*/;
assign _5204_ = _5196_ & _5203_ /*2442*/;
assign _5048_ = _5196_ ^ _5203_ /*2443*/;
assign _5201_ = _5202_ | _5204_ /*2440*/;
assign _5209_ = zeroWire ^ Q[6] /*2439*/;
assign _5206_ = _4855_ & _5209_ /*2435*/;
assign _5207_ = _4855_ ^ _5209_ /*2438*/;
assign _5208_ = _5201_ & _5207_ /*2436*/;
assign _5049_ = _5201_ ^ _5207_ /*2437*/;
assign Q[5] = _5206_ | _5208_ /*2434*/;
assign _5248_ = D[0] ^ Q[5] /*2240*/;
assign _5245_ = R_0[4] & _5248_ /*2236*/;
assign _5246_ = R_0[4] ^ _5248_ /*2239*/;
assign _5247_ = Q[5] & _5246_ /*2237*/;
assign _5211_ = Q[5] ^ _5246_ /*2238*/;
assign _5244_ = _5245_ | _5247_ /*2235*/;
assign _5253_ = D[1] ^ Q[5] /*2234*/;
assign _5250_ = _5018_ & _5253_ /*2230*/;
assign _5251_ = _5018_ ^ _5253_ /*2233*/;
assign _5252_ = _5244_ & _5251_ /*2231*/;
assign _5212_ = _5244_ ^ _5251_ /*2232*/;
assign _5249_ = _5250_ | _5252_ /*2229*/;
assign _5258_ = D[2] ^ Q[5] /*2228*/;
assign _5255_ = _5019_ & _5258_ /*2224*/;
assign _5256_ = _5019_ ^ _5258_ /*2227*/;
assign _5257_ = _5249_ & _5256_ /*2225*/;
assign _5213_ = _5249_ ^ _5256_ /*2226*/;
assign _5254_ = _5255_ | _5257_ /*2223*/;
assign _5263_ = D[3] ^ Q[5] /*2222*/;
assign _5260_ = _5020_ & _5263_ /*2218*/;
assign _5261_ = _5020_ ^ _5263_ /*2221*/;
assign _5262_ = _5254_ & _5261_ /*2219*/;
assign _5214_ = _5254_ ^ _5261_ /*2220*/;
assign _5259_ = _5260_ | _5262_ /*2217*/;
assign _5268_ = D[4] ^ Q[5] /*2216*/;
assign _5265_ = _5021_ & _5268_ /*2212*/;
assign _5266_ = _5021_ ^ _5268_ /*2215*/;
assign _5267_ = _5259_ & _5266_ /*2213*/;
assign _5215_ = _5259_ ^ _5266_ /*2214*/;
assign _5264_ = _5265_ | _5267_ /*2211*/;
assign _5273_ = D[5] ^ Q[5] /*2210*/;
assign _5270_ = _5022_ & _5273_ /*2206*/;
assign _5271_ = _5022_ ^ _5273_ /*2209*/;
assign _5272_ = _5264_ & _5271_ /*2207*/;
assign _5216_ = _5264_ ^ _5271_ /*2208*/;
assign _5269_ = _5270_ | _5272_ /*2205*/;
assign _5278_ = D[6] ^ Q[5] /*2204*/;
assign _5275_ = _5023_ & _5278_ /*2200*/;
assign _5276_ = _5023_ ^ _5278_ /*2203*/;
assign _5277_ = _5269_ & _5276_ /*2201*/;
assign _5217_ = _5269_ ^ _5276_ /*2202*/;
assign _5274_ = _5275_ | _5277_ /*2199*/;
assign _5283_ = D[7] ^ Q[5] /*2198*/;
assign _5280_ = _5024_ & _5283_ /*2194*/;
assign _5281_ = _5024_ ^ _5283_ /*2197*/;
assign _5282_ = _5274_ & _5281_ /*2195*/;
assign _5218_ = _5274_ ^ _5281_ /*2196*/;
assign _5279_ = _5280_ | _5282_ /*2193*/;
assign _5288_ = D[8] ^ Q[5] /*2192*/;
assign _5285_ = _5025_ & _5288_ /*2188*/;
assign _5286_ = _5025_ ^ _5288_ /*2191*/;
assign _5287_ = _5279_ & _5286_ /*2189*/;
assign _5219_ = _5279_ ^ _5286_ /*2190*/;
assign _5284_ = _5285_ | _5287_ /*2187*/;
assign _5293_ = D[9] ^ Q[5] /*2186*/;
assign _5290_ = _5026_ & _5293_ /*2182*/;
assign _5291_ = _5026_ ^ _5293_ /*2185*/;
assign _5292_ = _5284_ & _5291_ /*2183*/;
assign _5220_ = _5284_ ^ _5291_ /*2184*/;
assign _5289_ = _5290_ | _5292_ /*2181*/;
assign _5298_ = D[10] ^ Q[5] /*2180*/;
assign _5295_ = _5027_ & _5298_ /*2176*/;
assign _5296_ = _5027_ ^ _5298_ /*2179*/;
assign _5297_ = _5289_ & _5296_ /*2177*/;
assign _5221_ = _5289_ ^ _5296_ /*2178*/;
assign _5294_ = _5295_ | _5297_ /*2175*/;
assign _5303_ = D[11] ^ Q[5] /*2174*/;
assign _5300_ = _5028_ & _5303_ /*2170*/;
assign _5301_ = _5028_ ^ _5303_ /*2173*/;
assign _5302_ = _5294_ & _5301_ /*2171*/;
assign _5222_ = _5294_ ^ _5301_ /*2172*/;
assign _5299_ = _5300_ | _5302_ /*2169*/;
assign _5308_ = D[12] ^ Q[5] /*2168*/;
assign _5305_ = _5029_ & _5308_ /*2164*/;
assign _5306_ = _5029_ ^ _5308_ /*2167*/;
assign _5307_ = _5299_ & _5306_ /*2165*/;
assign _5223_ = _5299_ ^ _5306_ /*2166*/;
assign _5304_ = _5305_ | _5307_ /*2163*/;
assign _5313_ = D[13] ^ Q[5] /*2162*/;
assign _5310_ = _5030_ & _5313_ /*2158*/;
assign _5311_ = _5030_ ^ _5313_ /*2161*/;
assign _5312_ = _5304_ & _5311_ /*2159*/;
assign _5224_ = _5304_ ^ _5311_ /*2160*/;
assign _5309_ = _5310_ | _5312_ /*2157*/;
assign _5318_ = D[14] ^ Q[5] /*2156*/;
assign _5315_ = _5031_ & _5318_ /*2152*/;
assign _5316_ = _5031_ ^ _5318_ /*2155*/;
assign _5317_ = _5309_ & _5316_ /*2153*/;
assign _5225_ = _5309_ ^ _5316_ /*2154*/;
assign _5314_ = _5315_ | _5317_ /*2151*/;
assign _5323_ = D[15] ^ Q[5] /*2150*/;
assign _5320_ = _5032_ & _5323_ /*2146*/;
assign _5321_ = _5032_ ^ _5323_ /*2149*/;
assign _5322_ = _5314_ & _5321_ /*2147*/;
assign _5226_ = _5314_ ^ _5321_ /*2148*/;
assign _5319_ = _5320_ | _5322_ /*2145*/;
assign _5328_ = D[16] ^ Q[5] /*2144*/;
assign _5325_ = _5033_ & _5328_ /*2140*/;
assign _5326_ = _5033_ ^ _5328_ /*2143*/;
assign _5327_ = _5319_ & _5326_ /*2141*/;
assign _5227_ = _5319_ ^ _5326_ /*2142*/;
assign _5324_ = _5325_ | _5327_ /*2139*/;
assign _5333_ = D[17] ^ Q[5] /*2138*/;
assign _5330_ = _5034_ & _5333_ /*2134*/;
assign _5331_ = _5034_ ^ _5333_ /*2137*/;
assign _5332_ = _5324_ & _5331_ /*2135*/;
assign _5228_ = _5324_ ^ _5331_ /*2136*/;
assign _5329_ = _5330_ | _5332_ /*2133*/;
assign _5338_ = D[18] ^ Q[5] /*2132*/;
assign _5335_ = _5035_ & _5338_ /*2128*/;
assign _5336_ = _5035_ ^ _5338_ /*2131*/;
assign _5337_ = _5329_ & _5336_ /*2129*/;
assign _5229_ = _5329_ ^ _5336_ /*2130*/;
assign _5334_ = _5335_ | _5337_ /*2127*/;
assign _5343_ = D[19] ^ Q[5] /*2126*/;
assign _5340_ = _5036_ & _5343_ /*2122*/;
assign _5341_ = _5036_ ^ _5343_ /*2125*/;
assign _5342_ = _5334_ & _5341_ /*2123*/;
assign _5230_ = _5334_ ^ _5341_ /*2124*/;
assign _5339_ = _5340_ | _5342_ /*2121*/;
assign _5348_ = D[20] ^ Q[5] /*2120*/;
assign _5345_ = _5037_ & _5348_ /*2116*/;
assign _5346_ = _5037_ ^ _5348_ /*2119*/;
assign _5347_ = _5339_ & _5346_ /*2117*/;
assign _5231_ = _5339_ ^ _5346_ /*2118*/;
assign _5344_ = _5345_ | _5347_ /*2115*/;
assign _5353_ = D[21] ^ Q[5] /*2114*/;
assign _5350_ = _5038_ & _5353_ /*2110*/;
assign _5351_ = _5038_ ^ _5353_ /*2113*/;
assign _5352_ = _5344_ & _5351_ /*2111*/;
assign _5232_ = _5344_ ^ _5351_ /*2112*/;
assign _5349_ = _5350_ | _5352_ /*2109*/;
assign _5358_ = D[22] ^ Q[5] /*2108*/;
assign _5355_ = _5039_ & _5358_ /*2104*/;
assign _5356_ = _5039_ ^ _5358_ /*2107*/;
assign _5357_ = _5349_ & _5356_ /*2105*/;
assign _5233_ = _5349_ ^ _5356_ /*2106*/;
assign _5354_ = _5355_ | _5357_ /*2103*/;
assign _5363_ = D[23] ^ Q[5] /*2102*/;
assign _5360_ = _5040_ & _5363_ /*2098*/;
assign _5361_ = _5040_ ^ _5363_ /*2101*/;
assign _5362_ = _5354_ & _5361_ /*2099*/;
assign _5234_ = _5354_ ^ _5361_ /*2100*/;
assign _5359_ = _5360_ | _5362_ /*2097*/;
assign _5368_ = D[24] ^ Q[5] /*2096*/;
assign _5365_ = _5041_ & _5368_ /*2092*/;
assign _5366_ = _5041_ ^ _5368_ /*2095*/;
assign _5367_ = _5359_ & _5366_ /*2093*/;
assign _5235_ = _5359_ ^ _5366_ /*2094*/;
assign _5364_ = _5365_ | _5367_ /*2091*/;
assign _5373_ = D[25] ^ Q[5] /*2090*/;
assign _5370_ = _5042_ & _5373_ /*2086*/;
assign _5371_ = _5042_ ^ _5373_ /*2089*/;
assign _5372_ = _5364_ & _5371_ /*2087*/;
assign _5236_ = _5364_ ^ _5371_ /*2088*/;
assign _5369_ = _5370_ | _5372_ /*2085*/;
assign _5378_ = D[26] ^ Q[5] /*2084*/;
assign _5375_ = _5043_ & _5378_ /*2080*/;
assign _5376_ = _5043_ ^ _5378_ /*2083*/;
assign _5377_ = _5369_ & _5376_ /*2081*/;
assign _5237_ = _5369_ ^ _5376_ /*2082*/;
assign _5374_ = _5375_ | _5377_ /*2079*/;
assign _5383_ = D[27] ^ Q[5] /*2078*/;
assign _5380_ = _5044_ & _5383_ /*2074*/;
assign _5381_ = _5044_ ^ _5383_ /*2077*/;
assign _5382_ = _5374_ & _5381_ /*2075*/;
assign _5238_ = _5374_ ^ _5381_ /*2076*/;
assign _5379_ = _5380_ | _5382_ /*2073*/;
assign _5388_ = D[28] ^ Q[5] /*2072*/;
assign _5385_ = _5045_ & _5388_ /*2068*/;
assign _5386_ = _5045_ ^ _5388_ /*2071*/;
assign _5387_ = _5379_ & _5386_ /*2069*/;
assign _5239_ = _5379_ ^ _5386_ /*2070*/;
assign _5384_ = _5385_ | _5387_ /*2067*/;
assign _5393_ = D[29] ^ Q[5] /*2066*/;
assign _5390_ = _5046_ & _5393_ /*2062*/;
assign _5391_ = _5046_ ^ _5393_ /*2065*/;
assign _5392_ = _5384_ & _5391_ /*2063*/;
assign _5240_ = _5384_ ^ _5391_ /*2064*/;
assign _5389_ = _5390_ | _5392_ /*2061*/;
assign _5398_ = D[30] ^ Q[5] /*2060*/;
assign _5395_ = _5047_ & _5398_ /*2056*/;
assign _5396_ = _5047_ ^ _5398_ /*2059*/;
assign _5397_ = _5389_ & _5396_ /*2057*/;
assign _5241_ = _5389_ ^ _5396_ /*2058*/;
assign _5394_ = _5395_ | _5397_ /*2055*/;
assign _5402_ = zeroWire ^ Q[5] /*2054*/;
assign _5399_ = _5048_ & _5402_ /*2050*/;
assign _5400_ = _5048_ ^ _5402_ /*2053*/;
assign _5401_ = _5394_ & _5400_ /*2051*/;
assign _5242_ = _5394_ ^ _5400_ /*2052*/;
assign Q[4] = _5399_ | _5401_ /*2049*/;
assign _5441_ = D[0] ^ Q[4] /*1855*/;
assign _5438_ = R_0[3] & _5441_ /*1851*/;
assign _5439_ = R_0[3] ^ _5441_ /*1854*/;
assign _5440_ = Q[4] & _5439_ /*1852*/;
assign _5404_ = Q[4] ^ _5439_ /*1853*/;
assign _5437_ = _5438_ | _5440_ /*1850*/;
assign _5446_ = D[1] ^ Q[4] /*1849*/;
assign _5443_ = _5211_ & _5446_ /*1845*/;
assign _5444_ = _5211_ ^ _5446_ /*1848*/;
assign _5445_ = _5437_ & _5444_ /*1846*/;
assign _5405_ = _5437_ ^ _5444_ /*1847*/;
assign _5442_ = _5443_ | _5445_ /*1844*/;
assign _5451_ = D[2] ^ Q[4] /*1843*/;
assign _5448_ = _5212_ & _5451_ /*1839*/;
assign _5449_ = _5212_ ^ _5451_ /*1842*/;
assign _5450_ = _5442_ & _5449_ /*1840*/;
assign _5406_ = _5442_ ^ _5449_ /*1841*/;
assign _5447_ = _5448_ | _5450_ /*1838*/;
assign _5456_ = D[3] ^ Q[4] /*1837*/;
assign _5453_ = _5213_ & _5456_ /*1833*/;
assign _5454_ = _5213_ ^ _5456_ /*1836*/;
assign _5455_ = _5447_ & _5454_ /*1834*/;
assign _5407_ = _5447_ ^ _5454_ /*1835*/;
assign _5452_ = _5453_ | _5455_ /*1832*/;
assign _5461_ = D[4] ^ Q[4] /*1831*/;
assign _5458_ = _5214_ & _5461_ /*1827*/;
assign _5459_ = _5214_ ^ _5461_ /*1830*/;
assign _5460_ = _5452_ & _5459_ /*1828*/;
assign _5408_ = _5452_ ^ _5459_ /*1829*/;
assign _5457_ = _5458_ | _5460_ /*1826*/;
assign _5466_ = D[5] ^ Q[4] /*1825*/;
assign _5463_ = _5215_ & _5466_ /*1821*/;
assign _5464_ = _5215_ ^ _5466_ /*1824*/;
assign _5465_ = _5457_ & _5464_ /*1822*/;
assign _5409_ = _5457_ ^ _5464_ /*1823*/;
assign _5462_ = _5463_ | _5465_ /*1820*/;
assign _5471_ = D[6] ^ Q[4] /*1819*/;
assign _5468_ = _5216_ & _5471_ /*1815*/;
assign _5469_ = _5216_ ^ _5471_ /*1818*/;
assign _5470_ = _5462_ & _5469_ /*1816*/;
assign _5410_ = _5462_ ^ _5469_ /*1817*/;
assign _5467_ = _5468_ | _5470_ /*1814*/;
assign _5476_ = D[7] ^ Q[4] /*1813*/;
assign _5473_ = _5217_ & _5476_ /*1809*/;
assign _5474_ = _5217_ ^ _5476_ /*1812*/;
assign _5475_ = _5467_ & _5474_ /*1810*/;
assign _5411_ = _5467_ ^ _5474_ /*1811*/;
assign _5472_ = _5473_ | _5475_ /*1808*/;
assign _5481_ = D[8] ^ Q[4] /*1807*/;
assign _5478_ = _5218_ & _5481_ /*1803*/;
assign _5479_ = _5218_ ^ _5481_ /*1806*/;
assign _5480_ = _5472_ & _5479_ /*1804*/;
assign _5412_ = _5472_ ^ _5479_ /*1805*/;
assign _5477_ = _5478_ | _5480_ /*1802*/;
assign _5486_ = D[9] ^ Q[4] /*1801*/;
assign _5483_ = _5219_ & _5486_ /*1797*/;
assign _5484_ = _5219_ ^ _5486_ /*1800*/;
assign _5485_ = _5477_ & _5484_ /*1798*/;
assign _5413_ = _5477_ ^ _5484_ /*1799*/;
assign _5482_ = _5483_ | _5485_ /*1796*/;
assign _5491_ = D[10] ^ Q[4] /*1795*/;
assign _5488_ = _5220_ & _5491_ /*1791*/;
assign _5489_ = _5220_ ^ _5491_ /*1794*/;
assign _5490_ = _5482_ & _5489_ /*1792*/;
assign _5414_ = _5482_ ^ _5489_ /*1793*/;
assign _5487_ = _5488_ | _5490_ /*1790*/;
assign _5496_ = D[11] ^ Q[4] /*1789*/;
assign _5493_ = _5221_ & _5496_ /*1785*/;
assign _5494_ = _5221_ ^ _5496_ /*1788*/;
assign _5495_ = _5487_ & _5494_ /*1786*/;
assign _5415_ = _5487_ ^ _5494_ /*1787*/;
assign _5492_ = _5493_ | _5495_ /*1784*/;
assign _5501_ = D[12] ^ Q[4] /*1783*/;
assign _5498_ = _5222_ & _5501_ /*1779*/;
assign _5499_ = _5222_ ^ _5501_ /*1782*/;
assign _5500_ = _5492_ & _5499_ /*1780*/;
assign _5416_ = _5492_ ^ _5499_ /*1781*/;
assign _5497_ = _5498_ | _5500_ /*1778*/;
assign _5506_ = D[13] ^ Q[4] /*1777*/;
assign _5503_ = _5223_ & _5506_ /*1773*/;
assign _5504_ = _5223_ ^ _5506_ /*1776*/;
assign _5505_ = _5497_ & _5504_ /*1774*/;
assign _5417_ = _5497_ ^ _5504_ /*1775*/;
assign _5502_ = _5503_ | _5505_ /*1772*/;
assign _5511_ = D[14] ^ Q[4] /*1771*/;
assign _5508_ = _5224_ & _5511_ /*1767*/;
assign _5509_ = _5224_ ^ _5511_ /*1770*/;
assign _5510_ = _5502_ & _5509_ /*1768*/;
assign _5418_ = _5502_ ^ _5509_ /*1769*/;
assign _5507_ = _5508_ | _5510_ /*1766*/;
assign _5516_ = D[15] ^ Q[4] /*1765*/;
assign _5513_ = _5225_ & _5516_ /*1761*/;
assign _5514_ = _5225_ ^ _5516_ /*1764*/;
assign _5515_ = _5507_ & _5514_ /*1762*/;
assign _5419_ = _5507_ ^ _5514_ /*1763*/;
assign _5512_ = _5513_ | _5515_ /*1760*/;
assign _5521_ = D[16] ^ Q[4] /*1759*/;
assign _5518_ = _5226_ & _5521_ /*1755*/;
assign _5519_ = _5226_ ^ _5521_ /*1758*/;
assign _5520_ = _5512_ & _5519_ /*1756*/;
assign _5420_ = _5512_ ^ _5519_ /*1757*/;
assign _5517_ = _5518_ | _5520_ /*1754*/;
assign _5526_ = D[17] ^ Q[4] /*1753*/;
assign _5523_ = _5227_ & _5526_ /*1749*/;
assign _5524_ = _5227_ ^ _5526_ /*1752*/;
assign _5525_ = _5517_ & _5524_ /*1750*/;
assign _5421_ = _5517_ ^ _5524_ /*1751*/;
assign _5522_ = _5523_ | _5525_ /*1748*/;
assign _5531_ = D[18] ^ Q[4] /*1747*/;
assign _5528_ = _5228_ & _5531_ /*1743*/;
assign _5529_ = _5228_ ^ _5531_ /*1746*/;
assign _5530_ = _5522_ & _5529_ /*1744*/;
assign _5422_ = _5522_ ^ _5529_ /*1745*/;
assign _5527_ = _5528_ | _5530_ /*1742*/;
assign _5536_ = D[19] ^ Q[4] /*1741*/;
assign _5533_ = _5229_ & _5536_ /*1737*/;
assign _5534_ = _5229_ ^ _5536_ /*1740*/;
assign _5535_ = _5527_ & _5534_ /*1738*/;
assign _5423_ = _5527_ ^ _5534_ /*1739*/;
assign _5532_ = _5533_ | _5535_ /*1736*/;
assign _5541_ = D[20] ^ Q[4] /*1735*/;
assign _5538_ = _5230_ & _5541_ /*1731*/;
assign _5539_ = _5230_ ^ _5541_ /*1734*/;
assign _5540_ = _5532_ & _5539_ /*1732*/;
assign _5424_ = _5532_ ^ _5539_ /*1733*/;
assign _5537_ = _5538_ | _5540_ /*1730*/;
assign _5546_ = D[21] ^ Q[4] /*1729*/;
assign _5543_ = _5231_ & _5546_ /*1725*/;
assign _5544_ = _5231_ ^ _5546_ /*1728*/;
assign _5545_ = _5537_ & _5544_ /*1726*/;
assign _5425_ = _5537_ ^ _5544_ /*1727*/;
assign _5542_ = _5543_ | _5545_ /*1724*/;
assign _5551_ = D[22] ^ Q[4] /*1723*/;
assign _5548_ = _5232_ & _5551_ /*1719*/;
assign _5549_ = _5232_ ^ _5551_ /*1722*/;
assign _5550_ = _5542_ & _5549_ /*1720*/;
assign _5426_ = _5542_ ^ _5549_ /*1721*/;
assign _5547_ = _5548_ | _5550_ /*1718*/;
assign _5556_ = D[23] ^ Q[4] /*1717*/;
assign _5553_ = _5233_ & _5556_ /*1713*/;
assign _5554_ = _5233_ ^ _5556_ /*1716*/;
assign _5555_ = _5547_ & _5554_ /*1714*/;
assign _5427_ = _5547_ ^ _5554_ /*1715*/;
assign _5552_ = _5553_ | _5555_ /*1712*/;
assign _5561_ = D[24] ^ Q[4] /*1711*/;
assign _5558_ = _5234_ & _5561_ /*1707*/;
assign _5559_ = _5234_ ^ _5561_ /*1710*/;
assign _5560_ = _5552_ & _5559_ /*1708*/;
assign _5428_ = _5552_ ^ _5559_ /*1709*/;
assign _5557_ = _5558_ | _5560_ /*1706*/;
assign _5566_ = D[25] ^ Q[4] /*1705*/;
assign _5563_ = _5235_ & _5566_ /*1701*/;
assign _5564_ = _5235_ ^ _5566_ /*1704*/;
assign _5565_ = _5557_ & _5564_ /*1702*/;
assign _5429_ = _5557_ ^ _5564_ /*1703*/;
assign _5562_ = _5563_ | _5565_ /*1700*/;
assign _5571_ = D[26] ^ Q[4] /*1699*/;
assign _5568_ = _5236_ & _5571_ /*1695*/;
assign _5569_ = _5236_ ^ _5571_ /*1698*/;
assign _5570_ = _5562_ & _5569_ /*1696*/;
assign _5430_ = _5562_ ^ _5569_ /*1697*/;
assign _5567_ = _5568_ | _5570_ /*1694*/;
assign _5576_ = D[27] ^ Q[4] /*1693*/;
assign _5573_ = _5237_ & _5576_ /*1689*/;
assign _5574_ = _5237_ ^ _5576_ /*1692*/;
assign _5575_ = _5567_ & _5574_ /*1690*/;
assign _5431_ = _5567_ ^ _5574_ /*1691*/;
assign _5572_ = _5573_ | _5575_ /*1688*/;
assign _5581_ = D[28] ^ Q[4] /*1687*/;
assign _5578_ = _5238_ & _5581_ /*1683*/;
assign _5579_ = _5238_ ^ _5581_ /*1686*/;
assign _5580_ = _5572_ & _5579_ /*1684*/;
assign _5432_ = _5572_ ^ _5579_ /*1685*/;
assign _5577_ = _5578_ | _5580_ /*1682*/;
assign _5586_ = D[29] ^ Q[4] /*1681*/;
assign _5583_ = _5239_ & _5586_ /*1677*/;
assign _5584_ = _5239_ ^ _5586_ /*1680*/;
assign _5585_ = _5577_ & _5584_ /*1678*/;
assign _5433_ = _5577_ ^ _5584_ /*1679*/;
assign _5582_ = _5583_ | _5585_ /*1676*/;
assign _5591_ = D[30] ^ Q[4] /*1675*/;
assign _5588_ = _5240_ & _5591_ /*1671*/;
assign _5589_ = _5240_ ^ _5591_ /*1674*/;
assign _5590_ = _5582_ & _5589_ /*1672*/;
assign _5434_ = _5582_ ^ _5589_ /*1673*/;
assign _5587_ = _5588_ | _5590_ /*1670*/;
assign _5595_ = zeroWire ^ Q[4] /*1669*/;
assign _5592_ = _5241_ & _5595_ /*1665*/;
assign _5593_ = _5241_ ^ _5595_ /*1668*/;
assign _5594_ = _5587_ & _5593_ /*1666*/;
assign _5435_ = _5587_ ^ _5593_ /*1667*/;
assign Q[3] = _5592_ | _5594_ /*1664*/;
assign _5634_ = D[0] ^ Q[3] /*1470*/;
assign _5631_ = R_0[2] & _5634_ /*1466*/;
assign _5632_ = R_0[2] ^ _5634_ /*1469*/;
assign _5633_ = Q[3] & _5632_ /*1467*/;
assign _5597_ = Q[3] ^ _5632_ /*1468*/;
assign _5630_ = _5631_ | _5633_ /*1465*/;
assign _5639_ = D[1] ^ Q[3] /*1464*/;
assign _5636_ = _5404_ & _5639_ /*1460*/;
assign _5637_ = _5404_ ^ _5639_ /*1463*/;
assign _5638_ = _5630_ & _5637_ /*1461*/;
assign _5598_ = _5630_ ^ _5637_ /*1462*/;
assign _5635_ = _5636_ | _5638_ /*1459*/;
assign _5644_ = D[2] ^ Q[3] /*1458*/;
assign _5641_ = _5405_ & _5644_ /*1454*/;
assign _5642_ = _5405_ ^ _5644_ /*1457*/;
assign _5643_ = _5635_ & _5642_ /*1455*/;
assign _5599_ = _5635_ ^ _5642_ /*1456*/;
assign _5640_ = _5641_ | _5643_ /*1453*/;
assign _5649_ = D[3] ^ Q[3] /*1452*/;
assign _5646_ = _5406_ & _5649_ /*1448*/;
assign _5647_ = _5406_ ^ _5649_ /*1451*/;
assign _5648_ = _5640_ & _5647_ /*1449*/;
assign _5600_ = _5640_ ^ _5647_ /*1450*/;
assign _5645_ = _5646_ | _5648_ /*1447*/;
assign _5654_ = D[4] ^ Q[3] /*1446*/;
assign _5651_ = _5407_ & _5654_ /*1442*/;
assign _5652_ = _5407_ ^ _5654_ /*1445*/;
assign _5653_ = _5645_ & _5652_ /*1443*/;
assign _5601_ = _5645_ ^ _5652_ /*1444*/;
assign _5650_ = _5651_ | _5653_ /*1441*/;
assign _5659_ = D[5] ^ Q[3] /*1440*/;
assign _5656_ = _5408_ & _5659_ /*1436*/;
assign _5657_ = _5408_ ^ _5659_ /*1439*/;
assign _5658_ = _5650_ & _5657_ /*1437*/;
assign _5602_ = _5650_ ^ _5657_ /*1438*/;
assign _5655_ = _5656_ | _5658_ /*1435*/;
assign _5664_ = D[6] ^ Q[3] /*1434*/;
assign _5661_ = _5409_ & _5664_ /*1430*/;
assign _5662_ = _5409_ ^ _5664_ /*1433*/;
assign _5663_ = _5655_ & _5662_ /*1431*/;
assign _5603_ = _5655_ ^ _5662_ /*1432*/;
assign _5660_ = _5661_ | _5663_ /*1429*/;
assign _5669_ = D[7] ^ Q[3] /*1428*/;
assign _5666_ = _5410_ & _5669_ /*1424*/;
assign _5667_ = _5410_ ^ _5669_ /*1427*/;
assign _5668_ = _5660_ & _5667_ /*1425*/;
assign _5604_ = _5660_ ^ _5667_ /*1426*/;
assign _5665_ = _5666_ | _5668_ /*1423*/;
assign _5674_ = D[8] ^ Q[3] /*1422*/;
assign _5671_ = _5411_ & _5674_ /*1418*/;
assign _5672_ = _5411_ ^ _5674_ /*1421*/;
assign _5673_ = _5665_ & _5672_ /*1419*/;
assign _5605_ = _5665_ ^ _5672_ /*1420*/;
assign _5670_ = _5671_ | _5673_ /*1417*/;
assign _5679_ = D[9] ^ Q[3] /*1416*/;
assign _5676_ = _5412_ & _5679_ /*1412*/;
assign _5677_ = _5412_ ^ _5679_ /*1415*/;
assign _5678_ = _5670_ & _5677_ /*1413*/;
assign _5606_ = _5670_ ^ _5677_ /*1414*/;
assign _5675_ = _5676_ | _5678_ /*1411*/;
assign _5684_ = D[10] ^ Q[3] /*1410*/;
assign _5681_ = _5413_ & _5684_ /*1406*/;
assign _5682_ = _5413_ ^ _5684_ /*1409*/;
assign _5683_ = _5675_ & _5682_ /*1407*/;
assign _5607_ = _5675_ ^ _5682_ /*1408*/;
assign _5680_ = _5681_ | _5683_ /*1405*/;
assign _5689_ = D[11] ^ Q[3] /*1404*/;
assign _5686_ = _5414_ & _5689_ /*1400*/;
assign _5687_ = _5414_ ^ _5689_ /*1403*/;
assign _5688_ = _5680_ & _5687_ /*1401*/;
assign _5608_ = _5680_ ^ _5687_ /*1402*/;
assign _5685_ = _5686_ | _5688_ /*1399*/;
assign _5694_ = D[12] ^ Q[3] /*1398*/;
assign _5691_ = _5415_ & _5694_ /*1394*/;
assign _5692_ = _5415_ ^ _5694_ /*1397*/;
assign _5693_ = _5685_ & _5692_ /*1395*/;
assign _5609_ = _5685_ ^ _5692_ /*1396*/;
assign _5690_ = _5691_ | _5693_ /*1393*/;
assign _5699_ = D[13] ^ Q[3] /*1392*/;
assign _5696_ = _5416_ & _5699_ /*1388*/;
assign _5697_ = _5416_ ^ _5699_ /*1391*/;
assign _5698_ = _5690_ & _5697_ /*1389*/;
assign _5610_ = _5690_ ^ _5697_ /*1390*/;
assign _5695_ = _5696_ | _5698_ /*1387*/;
assign _5704_ = D[14] ^ Q[3] /*1386*/;
assign _5701_ = _5417_ & _5704_ /*1382*/;
assign _5702_ = _5417_ ^ _5704_ /*1385*/;
assign _5703_ = _5695_ & _5702_ /*1383*/;
assign _5611_ = _5695_ ^ _5702_ /*1384*/;
assign _5700_ = _5701_ | _5703_ /*1381*/;
assign _5709_ = D[15] ^ Q[3] /*1380*/;
assign _5706_ = _5418_ & _5709_ /*1376*/;
assign _5707_ = _5418_ ^ _5709_ /*1379*/;
assign _5708_ = _5700_ & _5707_ /*1377*/;
assign _5612_ = _5700_ ^ _5707_ /*1378*/;
assign _5705_ = _5706_ | _5708_ /*1375*/;
assign _5714_ = D[16] ^ Q[3] /*1374*/;
assign _5711_ = _5419_ & _5714_ /*1370*/;
assign _5712_ = _5419_ ^ _5714_ /*1373*/;
assign _5713_ = _5705_ & _5712_ /*1371*/;
assign _5613_ = _5705_ ^ _5712_ /*1372*/;
assign _5710_ = _5711_ | _5713_ /*1369*/;
assign _5719_ = D[17] ^ Q[3] /*1368*/;
assign _5716_ = _5420_ & _5719_ /*1364*/;
assign _5717_ = _5420_ ^ _5719_ /*1367*/;
assign _5718_ = _5710_ & _5717_ /*1365*/;
assign _5614_ = _5710_ ^ _5717_ /*1366*/;
assign _5715_ = _5716_ | _5718_ /*1363*/;
assign _5724_ = D[18] ^ Q[3] /*1362*/;
assign _5721_ = _5421_ & _5724_ /*1358*/;
assign _5722_ = _5421_ ^ _5724_ /*1361*/;
assign _5723_ = _5715_ & _5722_ /*1359*/;
assign _5615_ = _5715_ ^ _5722_ /*1360*/;
assign _5720_ = _5721_ | _5723_ /*1357*/;
assign _5729_ = D[19] ^ Q[3] /*1356*/;
assign _5726_ = _5422_ & _5729_ /*1352*/;
assign _5727_ = _5422_ ^ _5729_ /*1355*/;
assign _5728_ = _5720_ & _5727_ /*1353*/;
assign _5616_ = _5720_ ^ _5727_ /*1354*/;
assign _5725_ = _5726_ | _5728_ /*1351*/;
assign _5734_ = D[20] ^ Q[3] /*1350*/;
assign _5731_ = _5423_ & _5734_ /*1346*/;
assign _5732_ = _5423_ ^ _5734_ /*1349*/;
assign _5733_ = _5725_ & _5732_ /*1347*/;
assign _5617_ = _5725_ ^ _5732_ /*1348*/;
assign _5730_ = _5731_ | _5733_ /*1345*/;
assign _5739_ = D[21] ^ Q[3] /*1344*/;
assign _5736_ = _5424_ & _5739_ /*1340*/;
assign _5737_ = _5424_ ^ _5739_ /*1343*/;
assign _5738_ = _5730_ & _5737_ /*1341*/;
assign _5618_ = _5730_ ^ _5737_ /*1342*/;
assign _5735_ = _5736_ | _5738_ /*1339*/;
assign _5744_ = D[22] ^ Q[3] /*1338*/;
assign _5741_ = _5425_ & _5744_ /*1334*/;
assign _5742_ = _5425_ ^ _5744_ /*1337*/;
assign _5743_ = _5735_ & _5742_ /*1335*/;
assign _5619_ = _5735_ ^ _5742_ /*1336*/;
assign _5740_ = _5741_ | _5743_ /*1333*/;
assign _5749_ = D[23] ^ Q[3] /*1332*/;
assign _5746_ = _5426_ & _5749_ /*1328*/;
assign _5747_ = _5426_ ^ _5749_ /*1331*/;
assign _5748_ = _5740_ & _5747_ /*1329*/;
assign _5620_ = _5740_ ^ _5747_ /*1330*/;
assign _5745_ = _5746_ | _5748_ /*1327*/;
assign _5754_ = D[24] ^ Q[3] /*1326*/;
assign _5751_ = _5427_ & _5754_ /*1322*/;
assign _5752_ = _5427_ ^ _5754_ /*1325*/;
assign _5753_ = _5745_ & _5752_ /*1323*/;
assign _5621_ = _5745_ ^ _5752_ /*1324*/;
assign _5750_ = _5751_ | _5753_ /*1321*/;
assign _5759_ = D[25] ^ Q[3] /*1320*/;
assign _5756_ = _5428_ & _5759_ /*1316*/;
assign _5757_ = _5428_ ^ _5759_ /*1319*/;
assign _5758_ = _5750_ & _5757_ /*1317*/;
assign _5622_ = _5750_ ^ _5757_ /*1318*/;
assign _5755_ = _5756_ | _5758_ /*1315*/;
assign _5764_ = D[26] ^ Q[3] /*1314*/;
assign _5761_ = _5429_ & _5764_ /*1310*/;
assign _5762_ = _5429_ ^ _5764_ /*1313*/;
assign _5763_ = _5755_ & _5762_ /*1311*/;
assign _5623_ = _5755_ ^ _5762_ /*1312*/;
assign _5760_ = _5761_ | _5763_ /*1309*/;
assign _5769_ = D[27] ^ Q[3] /*1308*/;
assign _5766_ = _5430_ & _5769_ /*1304*/;
assign _5767_ = _5430_ ^ _5769_ /*1307*/;
assign _5768_ = _5760_ & _5767_ /*1305*/;
assign _5624_ = _5760_ ^ _5767_ /*1306*/;
assign _5765_ = _5766_ | _5768_ /*1303*/;
assign _5774_ = D[28] ^ Q[3] /*1302*/;
assign _5771_ = _5431_ & _5774_ /*1298*/;
assign _5772_ = _5431_ ^ _5774_ /*1301*/;
assign _5773_ = _5765_ & _5772_ /*1299*/;
assign _5625_ = _5765_ ^ _5772_ /*1300*/;
assign _5770_ = _5771_ | _5773_ /*1297*/;
assign _5779_ = D[29] ^ Q[3] /*1296*/;
assign _5776_ = _5432_ & _5779_ /*1292*/;
assign _5777_ = _5432_ ^ _5779_ /*1295*/;
assign _5778_ = _5770_ & _5777_ /*1293*/;
assign _5626_ = _5770_ ^ _5777_ /*1294*/;
assign _5775_ = _5776_ | _5778_ /*1291*/;
assign _5784_ = D[30] ^ Q[3] /*1290*/;
assign _5781_ = _5433_ & _5784_ /*1286*/;
assign _5782_ = _5433_ ^ _5784_ /*1289*/;
assign _5783_ = _5775_ & _5782_ /*1287*/;
assign _5627_ = _5775_ ^ _5782_ /*1288*/;
assign _5780_ = _5781_ | _5783_ /*1285*/;
assign _5788_ = zeroWire ^ Q[3] /*1284*/;
assign _5785_ = _5434_ & _5788_ /*1280*/;
assign _5786_ = _5434_ ^ _5788_ /*1283*/;
assign _5787_ = _5780_ & _5786_ /*1281*/;
assign _5628_ = _5780_ ^ _5786_ /*1282*/;
assign Q[2] = _5785_ | _5787_ /*1279*/;
assign _5827_ = D[0] ^ Q[2] /*1085*/;
assign _5824_ = R_0[1] & _5827_ /*1081*/;
assign _5825_ = R_0[1] ^ _5827_ /*1084*/;
assign _5826_ = Q[2] & _5825_ /*1082*/;
assign _5790_ = Q[2] ^ _5825_ /*1083*/;
assign _5823_ = _5824_ | _5826_ /*1080*/;
assign _5832_ = D[1] ^ Q[2] /*1079*/;
assign _5829_ = _5597_ & _5832_ /*1075*/;
assign _5830_ = _5597_ ^ _5832_ /*1078*/;
assign _5831_ = _5823_ & _5830_ /*1076*/;
assign _5791_ = _5823_ ^ _5830_ /*1077*/;
assign _5828_ = _5829_ | _5831_ /*1074*/;
assign _5837_ = D[2] ^ Q[2] /*1073*/;
assign _5834_ = _5598_ & _5837_ /*1069*/;
assign _5835_ = _5598_ ^ _5837_ /*1072*/;
assign _5836_ = _5828_ & _5835_ /*1070*/;
assign _5792_ = _5828_ ^ _5835_ /*1071*/;
assign _5833_ = _5834_ | _5836_ /*1068*/;
assign _5842_ = D[3] ^ Q[2] /*1067*/;
assign _5839_ = _5599_ & _5842_ /*1063*/;
assign _5840_ = _5599_ ^ _5842_ /*1066*/;
assign _5841_ = _5833_ & _5840_ /*1064*/;
assign _5793_ = _5833_ ^ _5840_ /*1065*/;
assign _5838_ = _5839_ | _5841_ /*1062*/;
assign _5847_ = D[4] ^ Q[2] /*1061*/;
assign _5844_ = _5600_ & _5847_ /*1057*/;
assign _5845_ = _5600_ ^ _5847_ /*1060*/;
assign _5846_ = _5838_ & _5845_ /*1058*/;
assign _5794_ = _5838_ ^ _5845_ /*1059*/;
assign _5843_ = _5844_ | _5846_ /*1056*/;
assign _5852_ = D[5] ^ Q[2] /*1055*/;
assign _5849_ = _5601_ & _5852_ /*1051*/;
assign _5850_ = _5601_ ^ _5852_ /*1054*/;
assign _5851_ = _5843_ & _5850_ /*1052*/;
assign _5795_ = _5843_ ^ _5850_ /*1053*/;
assign _5848_ = _5849_ | _5851_ /*1050*/;
assign _5857_ = D[6] ^ Q[2] /*1049*/;
assign _5854_ = _5602_ & _5857_ /*1045*/;
assign _5855_ = _5602_ ^ _5857_ /*1048*/;
assign _5856_ = _5848_ & _5855_ /*1046*/;
assign _5796_ = _5848_ ^ _5855_ /*1047*/;
assign _5853_ = _5854_ | _5856_ /*1044*/;
assign _5862_ = D[7] ^ Q[2] /*1043*/;
assign _5859_ = _5603_ & _5862_ /*1039*/;
assign _5860_ = _5603_ ^ _5862_ /*1042*/;
assign _5861_ = _5853_ & _5860_ /*1040*/;
assign _5797_ = _5853_ ^ _5860_ /*1041*/;
assign _5858_ = _5859_ | _5861_ /*1038*/;
assign _5867_ = D[8] ^ Q[2] /*1037*/;
assign _5864_ = _5604_ & _5867_ /*1033*/;
assign _5865_ = _5604_ ^ _5867_ /*1036*/;
assign _5866_ = _5858_ & _5865_ /*1034*/;
assign _5798_ = _5858_ ^ _5865_ /*1035*/;
assign _5863_ = _5864_ | _5866_ /*1032*/;
assign _5872_ = D[9] ^ Q[2] /*1031*/;
assign _5869_ = _5605_ & _5872_ /*1027*/;
assign _5870_ = _5605_ ^ _5872_ /*1030*/;
assign _5871_ = _5863_ & _5870_ /*1028*/;
assign _5799_ = _5863_ ^ _5870_ /*1029*/;
assign _5868_ = _5869_ | _5871_ /*1026*/;
assign _5877_ = D[10] ^ Q[2] /*1025*/;
assign _5874_ = _5606_ & _5877_ /*1021*/;
assign _5875_ = _5606_ ^ _5877_ /*1024*/;
assign _5876_ = _5868_ & _5875_ /*1022*/;
assign _5800_ = _5868_ ^ _5875_ /*1023*/;
assign _5873_ = _5874_ | _5876_ /*1020*/;
assign _5882_ = D[11] ^ Q[2] /*1019*/;
assign _5879_ = _5607_ & _5882_ /*1015*/;
assign _5880_ = _5607_ ^ _5882_ /*1018*/;
assign _5881_ = _5873_ & _5880_ /*1016*/;
assign _5801_ = _5873_ ^ _5880_ /*1017*/;
assign _5878_ = _5879_ | _5881_ /*1014*/;
assign _5887_ = D[12] ^ Q[2] /*1013*/;
assign _5884_ = _5608_ & _5887_ /*1009*/;
assign _5885_ = _5608_ ^ _5887_ /*1012*/;
assign _5886_ = _5878_ & _5885_ /*1010*/;
assign _5802_ = _5878_ ^ _5885_ /*1011*/;
assign _5883_ = _5884_ | _5886_ /*1008*/;
assign _5892_ = D[13] ^ Q[2] /*1007*/;
assign _5889_ = _5609_ & _5892_ /*1003*/;
assign _5890_ = _5609_ ^ _5892_ /*1006*/;
assign _5891_ = _5883_ & _5890_ /*1004*/;
assign _5803_ = _5883_ ^ _5890_ /*1005*/;
assign _5888_ = _5889_ | _5891_ /*1002*/;
assign _5897_ = D[14] ^ Q[2] /*1001*/;
assign _5894_ = _5610_ & _5897_ /*997*/;
assign _5895_ = _5610_ ^ _5897_ /*1000*/;
assign _5896_ = _5888_ & _5895_ /*998*/;
assign _5804_ = _5888_ ^ _5895_ /*999*/;
assign _5893_ = _5894_ | _5896_ /*996*/;
assign _5902_ = D[15] ^ Q[2] /*995*/;
assign _5899_ = _5611_ & _5902_ /*991*/;
assign _5900_ = _5611_ ^ _5902_ /*994*/;
assign _5901_ = _5893_ & _5900_ /*992*/;
assign _5805_ = _5893_ ^ _5900_ /*993*/;
assign _5898_ = _5899_ | _5901_ /*990*/;
assign _5907_ = D[16] ^ Q[2] /*989*/;
assign _5904_ = _5612_ & _5907_ /*985*/;
assign _5905_ = _5612_ ^ _5907_ /*988*/;
assign _5906_ = _5898_ & _5905_ /*986*/;
assign _5806_ = _5898_ ^ _5905_ /*987*/;
assign _5903_ = _5904_ | _5906_ /*984*/;
assign _5912_ = D[17] ^ Q[2] /*983*/;
assign _5909_ = _5613_ & _5912_ /*979*/;
assign _5910_ = _5613_ ^ _5912_ /*982*/;
assign _5911_ = _5903_ & _5910_ /*980*/;
assign _5807_ = _5903_ ^ _5910_ /*981*/;
assign _5908_ = _5909_ | _5911_ /*978*/;
assign _5917_ = D[18] ^ Q[2] /*977*/;
assign _5914_ = _5614_ & _5917_ /*973*/;
assign _5915_ = _5614_ ^ _5917_ /*976*/;
assign _5916_ = _5908_ & _5915_ /*974*/;
assign _5808_ = _5908_ ^ _5915_ /*975*/;
assign _5913_ = _5914_ | _5916_ /*972*/;
assign _5922_ = D[19] ^ Q[2] /*971*/;
assign _5919_ = _5615_ & _5922_ /*967*/;
assign _5920_ = _5615_ ^ _5922_ /*970*/;
assign _5921_ = _5913_ & _5920_ /*968*/;
assign _5809_ = _5913_ ^ _5920_ /*969*/;
assign _5918_ = _5919_ | _5921_ /*966*/;
assign _5927_ = D[20] ^ Q[2] /*965*/;
assign _5924_ = _5616_ & _5927_ /*961*/;
assign _5925_ = _5616_ ^ _5927_ /*964*/;
assign _5926_ = _5918_ & _5925_ /*962*/;
assign _5810_ = _5918_ ^ _5925_ /*963*/;
assign _5923_ = _5924_ | _5926_ /*960*/;
assign _5932_ = D[21] ^ Q[2] /*959*/;
assign _5929_ = _5617_ & _5932_ /*955*/;
assign _5930_ = _5617_ ^ _5932_ /*958*/;
assign _5931_ = _5923_ & _5930_ /*956*/;
assign _5811_ = _5923_ ^ _5930_ /*957*/;
assign _5928_ = _5929_ | _5931_ /*954*/;
assign _5937_ = D[22] ^ Q[2] /*953*/;
assign _5934_ = _5618_ & _5937_ /*949*/;
assign _5935_ = _5618_ ^ _5937_ /*952*/;
assign _5936_ = _5928_ & _5935_ /*950*/;
assign _5812_ = _5928_ ^ _5935_ /*951*/;
assign _5933_ = _5934_ | _5936_ /*948*/;
assign _5942_ = D[23] ^ Q[2] /*947*/;
assign _5939_ = _5619_ & _5942_ /*943*/;
assign _5940_ = _5619_ ^ _5942_ /*946*/;
assign _5941_ = _5933_ & _5940_ /*944*/;
assign _5813_ = _5933_ ^ _5940_ /*945*/;
assign _5938_ = _5939_ | _5941_ /*942*/;
assign _5947_ = D[24] ^ Q[2] /*941*/;
assign _5944_ = _5620_ & _5947_ /*937*/;
assign _5945_ = _5620_ ^ _5947_ /*940*/;
assign _5946_ = _5938_ & _5945_ /*938*/;
assign _5814_ = _5938_ ^ _5945_ /*939*/;
assign _5943_ = _5944_ | _5946_ /*936*/;
assign _5952_ = D[25] ^ Q[2] /*935*/;
assign _5949_ = _5621_ & _5952_ /*931*/;
assign _5950_ = _5621_ ^ _5952_ /*934*/;
assign _5951_ = _5943_ & _5950_ /*932*/;
assign _5815_ = _5943_ ^ _5950_ /*933*/;
assign _5948_ = _5949_ | _5951_ /*930*/;
assign _5957_ = D[26] ^ Q[2] /*929*/;
assign _5954_ = _5622_ & _5957_ /*925*/;
assign _5955_ = _5622_ ^ _5957_ /*928*/;
assign _5956_ = _5948_ & _5955_ /*926*/;
assign _5816_ = _5948_ ^ _5955_ /*927*/;
assign _5953_ = _5954_ | _5956_ /*924*/;
assign _5962_ = D[27] ^ Q[2] /*923*/;
assign _5959_ = _5623_ & _5962_ /*919*/;
assign _5960_ = _5623_ ^ _5962_ /*922*/;
assign _5961_ = _5953_ & _5960_ /*920*/;
assign _5817_ = _5953_ ^ _5960_ /*921*/;
assign _5958_ = _5959_ | _5961_ /*918*/;
assign _5967_ = D[28] ^ Q[2] /*917*/;
assign _5964_ = _5624_ & _5967_ /*913*/;
assign _5965_ = _5624_ ^ _5967_ /*916*/;
assign _5966_ = _5958_ & _5965_ /*914*/;
assign _5818_ = _5958_ ^ _5965_ /*915*/;
assign _5963_ = _5964_ | _5966_ /*912*/;
assign _5972_ = D[29] ^ Q[2] /*911*/;
assign _5969_ = _5625_ & _5972_ /*907*/;
assign _5970_ = _5625_ ^ _5972_ /*910*/;
assign _5971_ = _5963_ & _5970_ /*908*/;
assign _5819_ = _5963_ ^ _5970_ /*909*/;
assign _5968_ = _5969_ | _5971_ /*906*/;
assign _5977_ = D[30] ^ Q[2] /*905*/;
assign _5974_ = _5626_ & _5977_ /*901*/;
assign _5975_ = _5626_ ^ _5977_ /*904*/;
assign _5976_ = _5968_ & _5975_ /*902*/;
assign _5820_ = _5968_ ^ _5975_ /*903*/;
assign _5973_ = _5974_ | _5976_ /*900*/;
assign _5981_ = zeroWire ^ Q[2] /*899*/;
assign _5978_ = _5627_ & _5981_ /*895*/;
assign _5979_ = _5627_ ^ _5981_ /*898*/;
assign _5980_ = _5973_ & _5979_ /*896*/;
assign _5821_ = _5973_ ^ _5979_ /*897*/;
assign Q[1] = _5978_ | _5980_ /*894*/;
assign _6020_ = D[0] ^ Q[1] /*700*/;
assign _6017_ = R_0[0] & _6020_ /*696*/;
assign _6018_ = R_0[0] ^ _6020_ /*699*/;
assign _6019_ = Q[1] & _6018_ /*697*/;
assign _5983_ = Q[1] ^ _6018_ /*698*/;
assign _6016_ = _6017_ | _6019_ /*695*/;
assign _6025_ = D[1] ^ Q[1] /*694*/;
assign _6022_ = _5790_ & _6025_ /*690*/;
assign _6023_ = _5790_ ^ _6025_ /*693*/;
assign _6024_ = _6016_ & _6023_ /*691*/;
assign _5984_ = _6016_ ^ _6023_ /*692*/;
assign _6021_ = _6022_ | _6024_ /*689*/;
assign _6030_ = D[2] ^ Q[1] /*688*/;
assign _6027_ = _5791_ & _6030_ /*684*/;
assign _6028_ = _5791_ ^ _6030_ /*687*/;
assign _6029_ = _6021_ & _6028_ /*685*/;
assign _5985_ = _6021_ ^ _6028_ /*686*/;
assign _6026_ = _6027_ | _6029_ /*683*/;
assign _6035_ = D[3] ^ Q[1] /*682*/;
assign _6032_ = _5792_ & _6035_ /*678*/;
assign _6033_ = _5792_ ^ _6035_ /*681*/;
assign _6034_ = _6026_ & _6033_ /*679*/;
assign _5986_ = _6026_ ^ _6033_ /*680*/;
assign _6031_ = _6032_ | _6034_ /*677*/;
assign _6040_ = D[4] ^ Q[1] /*676*/;
assign _6037_ = _5793_ & _6040_ /*672*/;
assign _6038_ = _5793_ ^ _6040_ /*675*/;
assign _6039_ = _6031_ & _6038_ /*673*/;
assign _5987_ = _6031_ ^ _6038_ /*674*/;
assign _6036_ = _6037_ | _6039_ /*671*/;
assign _6045_ = D[5] ^ Q[1] /*670*/;
assign _6042_ = _5794_ & _6045_ /*666*/;
assign _6043_ = _5794_ ^ _6045_ /*669*/;
assign _6044_ = _6036_ & _6043_ /*667*/;
assign _5988_ = _6036_ ^ _6043_ /*668*/;
assign _6041_ = _6042_ | _6044_ /*665*/;
assign _6050_ = D[6] ^ Q[1] /*664*/;
assign _6047_ = _5795_ & _6050_ /*660*/;
assign _6048_ = _5795_ ^ _6050_ /*663*/;
assign _6049_ = _6041_ & _6048_ /*661*/;
assign _5989_ = _6041_ ^ _6048_ /*662*/;
assign _6046_ = _6047_ | _6049_ /*659*/;
assign _6055_ = D[7] ^ Q[1] /*658*/;
assign _6052_ = _5796_ & _6055_ /*654*/;
assign _6053_ = _5796_ ^ _6055_ /*657*/;
assign _6054_ = _6046_ & _6053_ /*655*/;
assign _5990_ = _6046_ ^ _6053_ /*656*/;
assign _6051_ = _6052_ | _6054_ /*653*/;
assign _6060_ = D[8] ^ Q[1] /*652*/;
assign _6057_ = _5797_ & _6060_ /*648*/;
assign _6058_ = _5797_ ^ _6060_ /*651*/;
assign _6059_ = _6051_ & _6058_ /*649*/;
assign _5991_ = _6051_ ^ _6058_ /*650*/;
assign _6056_ = _6057_ | _6059_ /*647*/;
assign _6065_ = D[9] ^ Q[1] /*646*/;
assign _6062_ = _5798_ & _6065_ /*642*/;
assign _6063_ = _5798_ ^ _6065_ /*645*/;
assign _6064_ = _6056_ & _6063_ /*643*/;
assign _5992_ = _6056_ ^ _6063_ /*644*/;
assign _6061_ = _6062_ | _6064_ /*641*/;
assign _6070_ = D[10] ^ Q[1] /*640*/;
assign _6067_ = _5799_ & _6070_ /*636*/;
assign _6068_ = _5799_ ^ _6070_ /*639*/;
assign _6069_ = _6061_ & _6068_ /*637*/;
assign _5993_ = _6061_ ^ _6068_ /*638*/;
assign _6066_ = _6067_ | _6069_ /*635*/;
assign _6075_ = D[11] ^ Q[1] /*634*/;
assign _6072_ = _5800_ & _6075_ /*630*/;
assign _6073_ = _5800_ ^ _6075_ /*633*/;
assign _6074_ = _6066_ & _6073_ /*631*/;
assign _5994_ = _6066_ ^ _6073_ /*632*/;
assign _6071_ = _6072_ | _6074_ /*629*/;
assign _6080_ = D[12] ^ Q[1] /*628*/;
assign _6077_ = _5801_ & _6080_ /*624*/;
assign _6078_ = _5801_ ^ _6080_ /*627*/;
assign _6079_ = _6071_ & _6078_ /*625*/;
assign _5995_ = _6071_ ^ _6078_ /*626*/;
assign _6076_ = _6077_ | _6079_ /*623*/;
assign _6085_ = D[13] ^ Q[1] /*622*/;
assign _6082_ = _5802_ & _6085_ /*618*/;
assign _6083_ = _5802_ ^ _6085_ /*621*/;
assign _6084_ = _6076_ & _6083_ /*619*/;
assign _5996_ = _6076_ ^ _6083_ /*620*/;
assign _6081_ = _6082_ | _6084_ /*617*/;
assign _6090_ = D[14] ^ Q[1] /*616*/;
assign _6087_ = _5803_ & _6090_ /*612*/;
assign _6088_ = _5803_ ^ _6090_ /*615*/;
assign _6089_ = _6081_ & _6088_ /*613*/;
assign _5997_ = _6081_ ^ _6088_ /*614*/;
assign _6086_ = _6087_ | _6089_ /*611*/;
assign _6095_ = D[15] ^ Q[1] /*610*/;
assign _6092_ = _5804_ & _6095_ /*606*/;
assign _6093_ = _5804_ ^ _6095_ /*609*/;
assign _6094_ = _6086_ & _6093_ /*607*/;
assign _5998_ = _6086_ ^ _6093_ /*608*/;
assign _6091_ = _6092_ | _6094_ /*605*/;
assign _6100_ = D[16] ^ Q[1] /*604*/;
assign _6097_ = _5805_ & _6100_ /*600*/;
assign _6098_ = _5805_ ^ _6100_ /*603*/;
assign _6099_ = _6091_ & _6098_ /*601*/;
assign _5999_ = _6091_ ^ _6098_ /*602*/;
assign _6096_ = _6097_ | _6099_ /*599*/;
assign _6105_ = D[17] ^ Q[1] /*598*/;
assign _6102_ = _5806_ & _6105_ /*594*/;
assign _6103_ = _5806_ ^ _6105_ /*597*/;
assign _6104_ = _6096_ & _6103_ /*595*/;
assign _6000_ = _6096_ ^ _6103_ /*596*/;
assign _6101_ = _6102_ | _6104_ /*593*/;
assign _6110_ = D[18] ^ Q[1] /*592*/;
assign _6107_ = _5807_ & _6110_ /*588*/;
assign _6108_ = _5807_ ^ _6110_ /*591*/;
assign _6109_ = _6101_ & _6108_ /*589*/;
assign _6001_ = _6101_ ^ _6108_ /*590*/;
assign _6106_ = _6107_ | _6109_ /*587*/;
assign _6115_ = D[19] ^ Q[1] /*586*/;
assign _6112_ = _5808_ & _6115_ /*582*/;
assign _6113_ = _5808_ ^ _6115_ /*585*/;
assign _6114_ = _6106_ & _6113_ /*583*/;
assign _6002_ = _6106_ ^ _6113_ /*584*/;
assign _6111_ = _6112_ | _6114_ /*581*/;
assign _6120_ = D[20] ^ Q[1] /*580*/;
assign _6117_ = _5809_ & _6120_ /*576*/;
assign _6118_ = _5809_ ^ _6120_ /*579*/;
assign _6119_ = _6111_ & _6118_ /*577*/;
assign _6003_ = _6111_ ^ _6118_ /*578*/;
assign _6116_ = _6117_ | _6119_ /*575*/;
assign _6125_ = D[21] ^ Q[1] /*574*/;
assign _6122_ = _5810_ & _6125_ /*570*/;
assign _6123_ = _5810_ ^ _6125_ /*573*/;
assign _6124_ = _6116_ & _6123_ /*571*/;
assign _6004_ = _6116_ ^ _6123_ /*572*/;
assign _6121_ = _6122_ | _6124_ /*569*/;
assign _6130_ = D[22] ^ Q[1] /*568*/;
assign _6127_ = _5811_ & _6130_ /*564*/;
assign _6128_ = _5811_ ^ _6130_ /*567*/;
assign _6129_ = _6121_ & _6128_ /*565*/;
assign _6005_ = _6121_ ^ _6128_ /*566*/;
assign _6126_ = _6127_ | _6129_ /*563*/;
assign _6135_ = D[23] ^ Q[1] /*562*/;
assign _6132_ = _5812_ & _6135_ /*558*/;
assign _6133_ = _5812_ ^ _6135_ /*561*/;
assign _6134_ = _6126_ & _6133_ /*559*/;
assign _6006_ = _6126_ ^ _6133_ /*560*/;
assign _6131_ = _6132_ | _6134_ /*557*/;
assign _6140_ = D[24] ^ Q[1] /*556*/;
assign _6137_ = _5813_ & _6140_ /*552*/;
assign _6138_ = _5813_ ^ _6140_ /*555*/;
assign _6139_ = _6131_ & _6138_ /*553*/;
assign _6007_ = _6131_ ^ _6138_ /*554*/;
assign _6136_ = _6137_ | _6139_ /*551*/;
assign _6145_ = D[25] ^ Q[1] /*550*/;
assign _6142_ = _5814_ & _6145_ /*546*/;
assign _6143_ = _5814_ ^ _6145_ /*549*/;
assign _6144_ = _6136_ & _6143_ /*547*/;
assign _6008_ = _6136_ ^ _6143_ /*548*/;
assign _6141_ = _6142_ | _6144_ /*545*/;
assign _6150_ = D[26] ^ Q[1] /*544*/;
assign _6147_ = _5815_ & _6150_ /*540*/;
assign _6148_ = _5815_ ^ _6150_ /*543*/;
assign _6149_ = _6141_ & _6148_ /*541*/;
assign _6009_ = _6141_ ^ _6148_ /*542*/;
assign _6146_ = _6147_ | _6149_ /*539*/;
assign _6155_ = D[27] ^ Q[1] /*538*/;
assign _6152_ = _5816_ & _6155_ /*534*/;
assign _6153_ = _5816_ ^ _6155_ /*537*/;
assign _6154_ = _6146_ & _6153_ /*535*/;
assign _6010_ = _6146_ ^ _6153_ /*536*/;
assign _6151_ = _6152_ | _6154_ /*533*/;
assign _6160_ = D[28] ^ Q[1] /*532*/;
assign _6157_ = _5817_ & _6160_ /*528*/;
assign _6158_ = _5817_ ^ _6160_ /*531*/;
assign _6159_ = _6151_ & _6158_ /*529*/;
assign _6011_ = _6151_ ^ _6158_ /*530*/;
assign _6156_ = _6157_ | _6159_ /*527*/;
assign _6165_ = D[29] ^ Q[1] /*526*/;
assign _6162_ = _5818_ & _6165_ /*522*/;
assign _6163_ = _5818_ ^ _6165_ /*525*/;
assign _6164_ = _6156_ & _6163_ /*523*/;
assign _6012_ = _6156_ ^ _6163_ /*524*/;
assign _6161_ = _6162_ | _6164_ /*521*/;
assign _6170_ = D[30] ^ Q[1] /*520*/;
assign _6167_ = _5819_ & _6170_ /*516*/;
assign _6168_ = _5819_ ^ _6170_ /*519*/;
assign _6169_ = _6161_ & _6168_ /*517*/;
assign _6013_ = _6161_ ^ _6168_ /*518*/;
assign _6166_ = _6167_ | _6169_ /*515*/;
assign _6174_ = zeroWire ^ Q[1] /*514*/;
assign _6171_ = _5820_ & _6174_ /*510*/;
assign _6172_ = _5820_ ^ _6174_ /*513*/;
assign _6173_ = _6166_ & _6172_ /*511*/;
assign _6014_ = _6166_ ^ _6172_ /*512*/;
assign Q[0] = _6171_ | _6173_ /*509*/;
assign _6178_ = ~Q[0] /*314*/;
assign _6177_ = _6178_ & D[0] /*313*/;
assign _6180_ = _5983_ & _6177_ /*308*/;
assign _6181_ = _5983_ ^ _6177_ /*311*/;
assign _6182_ = zeroWire & _6181_ /*309*/;
assign R_n1[0] = zeroWire ^ _6181_ /*310*/;
assign _6179_ = _6180_ | _6182_ /*307*/;
assign _6184_ = ~Q[0] /*306*/;
assign _6183_ = _6184_ & D[1] /*305*/;
assign _6186_ = _5984_ & _6183_ /*300*/;
assign _6187_ = _5984_ ^ _6183_ /*303*/;
assign _6188_ = _6179_ & _6187_ /*301*/;
assign R_n1[1] = _6179_ ^ _6187_ /*302*/;
assign _6185_ = _6186_ | _6188_ /*299*/;
assign _6190_ = ~Q[0] /*298*/;
assign _6189_ = _6190_ & D[2] /*297*/;
assign _6192_ = _5985_ & _6189_ /*292*/;
assign _6193_ = _5985_ ^ _6189_ /*295*/;
assign _6194_ = _6185_ & _6193_ /*293*/;
assign R_n1[2] = _6185_ ^ _6193_ /*294*/;
assign _6191_ = _6192_ | _6194_ /*291*/;
assign _6196_ = ~Q[0] /*290*/;
assign _6195_ = _6196_ & D[3] /*289*/;
assign _6198_ = _5986_ & _6195_ /*284*/;
assign _6199_ = _5986_ ^ _6195_ /*287*/;
assign _6200_ = _6191_ & _6199_ /*285*/;
assign R_n1[3] = _6191_ ^ _6199_ /*286*/;
assign _6197_ = _6198_ | _6200_ /*283*/;
assign _6202_ = ~Q[0] /*282*/;
assign _6201_ = _6202_ & D[4] /*281*/;
assign _6204_ = _5987_ & _6201_ /*276*/;
assign _6205_ = _5987_ ^ _6201_ /*279*/;
assign _6206_ = _6197_ & _6205_ /*277*/;
assign R_n1[4] = _6197_ ^ _6205_ /*278*/;
assign _6203_ = _6204_ | _6206_ /*275*/;
assign _6208_ = ~Q[0] /*274*/;
assign _6207_ = _6208_ & D[5] /*273*/;
assign _6210_ = _5988_ & _6207_ /*268*/;
assign _6211_ = _5988_ ^ _6207_ /*271*/;
assign _6212_ = _6203_ & _6211_ /*269*/;
assign R_n1[5] = _6203_ ^ _6211_ /*270*/;
assign _6209_ = _6210_ | _6212_ /*267*/;
assign _6214_ = ~Q[0] /*266*/;
assign _6213_ = _6214_ & D[6] /*265*/;
assign _6216_ = _5989_ & _6213_ /*260*/;
assign _6217_ = _5989_ ^ _6213_ /*263*/;
assign _6218_ = _6209_ & _6217_ /*261*/;
assign R_n1[6] = _6209_ ^ _6217_ /*262*/;
assign _6215_ = _6216_ | _6218_ /*259*/;
assign _6220_ = ~Q[0] /*258*/;
assign _6219_ = _6220_ & D[7] /*257*/;
assign _6222_ = _5990_ & _6219_ /*252*/;
assign _6223_ = _5990_ ^ _6219_ /*255*/;
assign _6224_ = _6215_ & _6223_ /*253*/;
assign R_n1[7] = _6215_ ^ _6223_ /*254*/;
assign _6221_ = _6222_ | _6224_ /*251*/;
assign _6226_ = ~Q[0] /*250*/;
assign _6225_ = _6226_ & D[8] /*249*/;
assign _6228_ = _5991_ & _6225_ /*244*/;
assign _6229_ = _5991_ ^ _6225_ /*247*/;
assign _6230_ = _6221_ & _6229_ /*245*/;
assign R_n1[8] = _6221_ ^ _6229_ /*246*/;
assign _6227_ = _6228_ | _6230_ /*243*/;
assign _6232_ = ~Q[0] /*242*/;
assign _6231_ = _6232_ & D[9] /*241*/;
assign _6234_ = _5992_ & _6231_ /*236*/;
assign _6235_ = _5992_ ^ _6231_ /*239*/;
assign _6236_ = _6227_ & _6235_ /*237*/;
assign R_n1[9] = _6227_ ^ _6235_ /*238*/;
assign _6233_ = _6234_ | _6236_ /*235*/;
assign _6238_ = ~Q[0] /*234*/;
assign _6237_ = _6238_ & D[10] /*233*/;
assign _6240_ = _5993_ & _6237_ /*228*/;
assign _6241_ = _5993_ ^ _6237_ /*231*/;
assign _6242_ = _6233_ & _6241_ /*229*/;
assign R_n1[10] = _6233_ ^ _6241_ /*230*/;
assign _6239_ = _6240_ | _6242_ /*227*/;
assign _6244_ = ~Q[0] /*226*/;
assign _6243_ = _6244_ & D[11] /*225*/;
assign _6246_ = _5994_ & _6243_ /*220*/;
assign _6247_ = _5994_ ^ _6243_ /*223*/;
assign _6248_ = _6239_ & _6247_ /*221*/;
assign R_n1[11] = _6239_ ^ _6247_ /*222*/;
assign _6245_ = _6246_ | _6248_ /*219*/;
assign _6250_ = ~Q[0] /*218*/;
assign _6249_ = _6250_ & D[12] /*217*/;
assign _6252_ = _5995_ & _6249_ /*212*/;
assign _6253_ = _5995_ ^ _6249_ /*215*/;
assign _6254_ = _6245_ & _6253_ /*213*/;
assign R_n1[12] = _6245_ ^ _6253_ /*214*/;
assign _6251_ = _6252_ | _6254_ /*211*/;
assign _6256_ = ~Q[0] /*210*/;
assign _6255_ = _6256_ & D[13] /*209*/;
assign _6258_ = _5996_ & _6255_ /*204*/;
assign _6259_ = _5996_ ^ _6255_ /*207*/;
assign _6260_ = _6251_ & _6259_ /*205*/;
assign R_n1[13] = _6251_ ^ _6259_ /*206*/;
assign _6257_ = _6258_ | _6260_ /*203*/;
assign _6262_ = ~Q[0] /*202*/;
assign _6261_ = _6262_ & D[14] /*201*/;
assign _6264_ = _5997_ & _6261_ /*196*/;
assign _6265_ = _5997_ ^ _6261_ /*199*/;
assign _6266_ = _6257_ & _6265_ /*197*/;
assign R_n1[14] = _6257_ ^ _6265_ /*198*/;
assign _6263_ = _6264_ | _6266_ /*195*/;
assign _6268_ = ~Q[0] /*194*/;
assign _6267_ = _6268_ & D[15] /*193*/;
assign _6270_ = _5998_ & _6267_ /*188*/;
assign _6271_ = _5998_ ^ _6267_ /*191*/;
assign _6272_ = _6263_ & _6271_ /*189*/;
assign R_n1[15] = _6263_ ^ _6271_ /*190*/;
assign _6269_ = _6270_ | _6272_ /*187*/;
assign _6274_ = ~Q[0] /*186*/;
assign _6273_ = _6274_ & D[16] /*185*/;
assign _6276_ = _5999_ & _6273_ /*180*/;
assign _6277_ = _5999_ ^ _6273_ /*183*/;
assign _6278_ = _6269_ & _6277_ /*181*/;
assign R_n1[16] = _6269_ ^ _6277_ /*182*/;
assign _6275_ = _6276_ | _6278_ /*179*/;
assign _6280_ = ~Q[0] /*178*/;
assign _6279_ = _6280_ & D[17] /*177*/;
assign _6282_ = _6000_ & _6279_ /*172*/;
assign _6283_ = _6000_ ^ _6279_ /*175*/;
assign _6284_ = _6275_ & _6283_ /*173*/;
assign R_n1[17] = _6275_ ^ _6283_ /*174*/;
assign _6281_ = _6282_ | _6284_ /*171*/;
assign _6286_ = ~Q[0] /*170*/;
assign _6285_ = _6286_ & D[18] /*169*/;
assign _6288_ = _6001_ & _6285_ /*164*/;
assign _6289_ = _6001_ ^ _6285_ /*167*/;
assign _6290_ = _6281_ & _6289_ /*165*/;
assign R_n1[18] = _6281_ ^ _6289_ /*166*/;
assign _6287_ = _6288_ | _6290_ /*163*/;
assign _6292_ = ~Q[0] /*162*/;
assign _6291_ = _6292_ & D[19] /*161*/;
assign _6294_ = _6002_ & _6291_ /*156*/;
assign _6295_ = _6002_ ^ _6291_ /*159*/;
assign _6296_ = _6287_ & _6295_ /*157*/;
assign R_n1[19] = _6287_ ^ _6295_ /*158*/;
assign _6293_ = _6294_ | _6296_ /*155*/;
assign _6298_ = ~Q[0] /*154*/;
assign _6297_ = _6298_ & D[20] /*153*/;
assign _6300_ = _6003_ & _6297_ /*148*/;
assign _6301_ = _6003_ ^ _6297_ /*151*/;
assign _6302_ = _6293_ & _6301_ /*149*/;
assign R_n1[20] = _6293_ ^ _6301_ /*150*/;
assign _6299_ = _6300_ | _6302_ /*147*/;
assign _6304_ = ~Q[0] /*146*/;
assign _6303_ = _6304_ & D[21] /*145*/;
assign _6306_ = _6004_ & _6303_ /*140*/;
assign _6307_ = _6004_ ^ _6303_ /*143*/;
assign _6308_ = _6299_ & _6307_ /*141*/;
assign R_n1[21] = _6299_ ^ _6307_ /*142*/;
assign _6305_ = _6306_ | _6308_ /*139*/;
assign _6310_ = ~Q[0] /*138*/;
assign _6309_ = _6310_ & D[22] /*137*/;
assign _6312_ = _6005_ & _6309_ /*132*/;
assign _6313_ = _6005_ ^ _6309_ /*135*/;
assign _6314_ = _6305_ & _6313_ /*133*/;
assign R_n1[22] = _6305_ ^ _6313_ /*134*/;
assign _6311_ = _6312_ | _6314_ /*131*/;
assign _6316_ = ~Q[0] /*130*/;
assign _6315_ = _6316_ & D[23] /*129*/;
assign _6318_ = _6006_ & _6315_ /*124*/;
assign _6319_ = _6006_ ^ _6315_ /*127*/;
assign _6320_ = _6311_ & _6319_ /*125*/;
assign R_n1[23] = _6311_ ^ _6319_ /*126*/;
assign _6317_ = _6318_ | _6320_ /*123*/;
assign _6322_ = ~Q[0] /*122*/;
assign _6321_ = _6322_ & D[24] /*121*/;
assign _6324_ = _6007_ & _6321_ /*116*/;
assign _6325_ = _6007_ ^ _6321_ /*119*/;
assign _6326_ = _6317_ & _6325_ /*117*/;
assign R_n1[24] = _6317_ ^ _6325_ /*118*/;
assign _6323_ = _6324_ | _6326_ /*115*/;
assign _6328_ = ~Q[0] /*114*/;
assign _6327_ = _6328_ & D[25] /*113*/;
assign _6330_ = _6008_ & _6327_ /*108*/;
assign _6331_ = _6008_ ^ _6327_ /*111*/;
assign _6332_ = _6323_ & _6331_ /*109*/;
assign R_n1[25] = _6323_ ^ _6331_ /*110*/;
assign _6329_ = _6330_ | _6332_ /*107*/;
assign _6334_ = ~Q[0] /*106*/;
assign _6333_ = _6334_ & D[26] /*105*/;
assign _6336_ = _6009_ & _6333_ /*100*/;
assign _6337_ = _6009_ ^ _6333_ /*103*/;
assign _6338_ = _6329_ & _6337_ /*101*/;
assign R_n1[26] = _6329_ ^ _6337_ /*102*/;
assign _6335_ = _6336_ | _6338_ /*99*/;
assign _6340_ = ~Q[0] /*98*/;
assign _6339_ = _6340_ & D[27] /*97*/;
assign _6342_ = _6010_ & _6339_ /*92*/;
assign _6343_ = _6010_ ^ _6339_ /*95*/;
assign _6344_ = _6335_ & _6343_ /*93*/;
assign R_n1[27] = _6335_ ^ _6343_ /*94*/;
assign _6341_ = _6342_ | _6344_ /*91*/;
assign _6346_ = ~Q[0] /*90*/;
assign _6345_ = _6346_ & D[28] /*89*/;
assign _6348_ = _6011_ & _6345_ /*84*/;
assign _6349_ = _6011_ ^ _6345_ /*87*/;
assign _6350_ = _6341_ & _6349_ /*85*/;
assign R_n1[28] = _6341_ ^ _6349_ /*86*/;
assign _6347_ = _6348_ | _6350_ /*83*/;
assign _6352_ = ~Q[0] /*82*/;
assign _6351_ = _6352_ & D[29] /*81*/;
assign _6354_ = _6012_ & _6351_ /*76*/;
assign _6355_ = _6012_ ^ _6351_ /*79*/;
assign _6356_ = _6347_ & _6355_ /*77*/;
assign R_n1[29] = _6347_ ^ _6355_ /*78*/;
assign _6353_ = _6354_ | _6356_ /*75*/;
assign _6358_ = ~Q[0] /*74*/;
assign _6357_ = _6358_ & D[30] /*73*/;
assign _6360_ = _6013_ & _6357_ /*68*/;
assign _6361_ = _6013_ ^ _6357_ /*71*/;
assign _6362_ = _6353_ & _6361_ /*69*/;
assign R_n1[30] = _6353_ ^ _6361_ /*70*/;
assign _6359_ = _6360_ | _6362_ /*67*/;
endmodule
