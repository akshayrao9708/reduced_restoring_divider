module divider(q, rout, rin, div);
  wire _0_;
  wire _1_;
  wire _2_;
  wire _3_;
  wire _4_;
  wire _5_;
  wire _6_;
  wire _7_;
  wire _8_;
  wire _9_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  wire _38_;
  wire _39_;
  wire _40_;
  wire _41_;
  wire _42_;
  wire _43_;
  wire _44_;
  wire _45_;
  wire _46_;
  wire _47_;
  wire _48_;
  wire _49_;
  wire _50_;
  wire _51_;
  wire _52_;
  wire _53_;
  wire _54_;
  wire _55_;
  wire _56_;
  wire _57_;
  wire _58_;
  wire _59_;
  wire _60_;
  wire _61_;
  wire _62_;
  wire _63_;
  wire _64_;
  wire _65_;
  wire _66_;
  wire _67_;
  wire _68_;
  wire _69_;
  wire _70_;
  wire _71_;
  wire _72_;
  wire _73_;
  wire _74_;
  wire _75_;
  wire _76_;
  wire _77_;
  wire _78_;
  wire _79_;
  wire _80_;
  wire _81_;
  wire _82_;
  wire _83_;
  wire _84_;
  wire _85_;
  wire _86_;
  wire _87_;
  wire _88_;
  wire _89_;
  wire _90_;
  wire _91_;
  wire _92_;
  wire _93_;
  wire _94_;
  wire _95_;
  wire _96_;
  wire _97_;
  wire _98_;
  wire _99_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire _304_;
  wire _305_;
  wire _306_;
  wire _307_;
  wire _308_;
  wire _309_;
  wire _310_;
  wire _311_;
  wire _312_;
  wire _313_;
  wire _314_;
  wire _315_;
  wire _316_;
  wire _317_;
  wire _318_;
  wire _319_;
  wire _320_;
  wire _321_;
  wire _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire _326_;
  wire _327_;
  wire _328_;
  wire _329_;
  wire _330_;
  wire _331_;
  wire _332_;
  wire _333_;
  wire _334_;
  wire _335_;
  wire _336_;
  wire _337_;
  wire _338_;
  wire _339_;
  wire _340_;
  wire _341_;
  wire _342_;
  wire _343_;
  wire _344_;
  wire _345_;
  wire _346_;
  wire _347_;
  wire _348_;
  wire _349_;
  wire _350_;
  wire _351_;
  wire _352_;
  wire _353_;
  wire _354_;
  wire _355_;
  wire _356_;
  wire _357_;
  wire _358_;
  wire _359_;
  wire _360_;
  wire _361_;
  wire _362_;
  wire _363_;
  wire _364_;
  wire _365_;
  wire _366_;
  wire _367_;
  wire _368_;
  wire _369_;
  wire _370_;
  wire _371_;
  wire _372_;
  wire _373_;
  wire _374_;
  wire _375_;
  wire _376_;
  wire _377_;
  wire _378_;
  wire _379_;
  wire _380_;
  wire _381_;
  wire _382_;
  wire _383_;
  wire _384_;
  wire _385_;
  wire _386_;
  wire _387_;
  wire _388_;
  wire _389_;
  wire _390_;
  wire _391_;
  wire _392_;
  wire _393_;
  wire _394_;
  wire _395_;
  wire _396_;
  wire _397_;
  wire _398_;
  wire _399_;
  wire _400_;
  wire _401_;
  wire _402_;
  wire _403_;
  wire _404_;
  wire _405_;
  wire _406_;
  wire _407_;
  wire _408_;
  wire _409_;
  wire _410_;
  wire _411_;
  wire _412_;
  wire _413_;
  wire _414_;
  wire _415_;
  wire _416_;
  wire _417_;
  wire _418_;
  wire _419_;
  wire _420_;
  wire _421_;
  wire _422_;
  wire _423_;
  wire _424_;
  wire _425_;
  wire _426_;
  wire _427_;
  wire _428_;
  wire _429_;
  wire _430_;
  wire _431_;
  wire _432_;
  wire _433_;
  wire _434_;
  wire _435_;
  wire _436_;
  wire _437_;
  wire _438_;
  wire _439_;
  wire _440_;
  wire _441_;
  wire _442_;
  wire _443_;
  wire _444_;
  wire _445_;
  wire _446_;
  wire _447_;
  wire _448_;
  wire _449_;
  wire _450_;
  wire _451_;
  wire _452_;
  wire _453_;
  wire _454_;
  wire _455_;
  wire _456_;
  wire _457_;
  wire _458_;
  wire _459_;
  wire _460_;
  wire _461_;
  wire _462_;
  wire _463_;
  wire _464_;
  wire _465_;
  wire _466_;
  wire _467_;
  wire _468_;
  wire _469_;
  wire _470_;
  wire _471_;
  wire _472_;
  wire _473_;
  wire _474_;
  wire _475_;
  wire _476_;
  wire _477_;
  wire _478_;
  wire _479_;
  wire _480_;
  wire _481_;
  wire _482_;
  wire _483_;
  wire _484_;
  wire _485_;
  wire _486_;
  wire _487_;
  wire _488_;
  wire _489_;
  wire _490_;
  wire _491_;
  wire _492_;
  wire _493_;
  wire _494_;
  wire _495_;
  wire _496_;
  wire _497_;
  wire _498_;
  wire _499_;
  wire _500_;
  wire _501_;
  wire _502_;
  wire _503_;
  wire _504_;
  wire _505_;
  wire _506_;
  wire _507_;
  wire _508_;
  wire _509_;
  wire _510_;
  wire _511_;
  wire _512_;
  wire _513_;
  wire _514_;
  wire _515_;
  wire _516_;
  wire _517_;
  wire _518_;
  wire _519_;
  wire _520_;
  wire _521_;
  wire _522_;
  wire _523_;
  wire _524_;
  wire _525_;
  wire _526_;
  wire _527_;
  wire _528_;
  wire _529_;
  wire _530_;
  wire _531_;
  wire _532_;
  wire _533_;
  wire _534_;
  wire _535_;
  wire _536_;
  wire _537_;
  wire _538_;
  wire _539_;
  wire _540_;
  wire _541_;
  wire _542_;
  wire _543_;
  wire _544_;
  wire _545_;
  wire _546_;
  wire _547_;
  wire _548_;
  wire _549_;
  wire _550_;
  wire _551_;
  wire _552_;
  wire _553_;
  wire _554_;
  wire _555_;
  wire _556_;
  wire _557_;
  wire _558_;
  wire _559_;
  wire _560_;
  wire _561_;
  wire _562_;
  wire _563_;
  wire _564_;
  wire _565_;
  wire _566_;
  wire _567_;
  wire _568_;
  wire _569_;
  wire _570_;
  wire _571_;
  wire _572_;
  wire _573_;
  wire _574_;
  wire _575_;
  wire _576_;
  wire _577_;
  wire _578_;
  wire _579_;
  wire _580_;
  wire _581_;
  wire _582_;
  wire _583_;
  wire _584_;
  wire _585_;
  wire _586_;
  wire _587_;
  wire _588_;
  wire _589_;
  wire _590_;
  wire _591_;
  wire _592_;
  wire _593_;
  wire _594_;
  wire _595_;
  wire _596_;
  wire _597_;
  wire _598_;
  wire _599_;
  wire _600_;
  wire _601_;
  wire _602_;
  wire _603_;
  wire _604_;
  wire _605_;
  wire _606_;
  wire _607_;
  wire _608_;
  wire _609_;
  wire _610_;
  wire _611_;
  wire _612_;
  wire _613_;
  wire _614_;
  wire _615_;
  wire _616_;
  wire _617_;
  wire _618_;
  wire _619_;
  wire _620_;
  wire _621_;
  wire _622_;
  wire _623_;
  wire _624_;
  wire _625_;
  wire _626_;
  wire _627_;
  wire _628_;
  wire _629_;
  wire _630_;
  wire _631_;
  wire _632_;
  wire _633_;
  wire _634_;
  wire _635_;
  wire _636_;
  wire _637_;
  wire _638_;
  wire _639_;
  wire _640_;
  wire _641_;
  wire _642_;
  wire _643_;
  wire _644_;
  wire _645_;
  wire _646_;
  wire _647_;
  wire _648_;
  wire _649_;
  wire _650_;
  wire _651_;
  wire _652_;
  wire _653_;
  wire _654_;
  wire _655_;
  wire _656_;
  wire _657_;
  wire _658_;
  wire _659_;
  wire _660_;
  wire _661_;
  wire _662_;
  wire _663_;
  wire _664_;
  wire _665_;
  wire _666_;
  wire _667_;
  wire _668_;
  wire _669_;
  wire _670_;
  wire _671_;
  wire _672_;
  wire _673_;
  wire _674_;
  wire _675_;
  wire _676_;
  wire _677_;
  wire _678_;
  wire _679_;
  wire _680_;
  wire _681_;
  wire _682_;
  wire _683_;
  wire _684_;
  wire _685_;
  wire _686_;
  wire _687_;
  wire _688_;
  wire _689_;
  wire _690_;
  wire _691_;
  wire _692_;
  wire _693_;
  wire _694_;
  wire _695_;
  wire _696_;
  wire _697_;
  wire _698_;
  wire _699_;
  wire _700_;
  wire _701_;
  wire _702_;
  wire _703_;
  wire _704_;
  wire _705_;
  wire _706_;
  wire _707_;
  wire _708_;
  wire _709_;
  wire _710_;
  wire _711_;
  wire _712_;
  wire _713_;
  wire _714_;
  wire _715_;
  wire _716_;
  wire _717_;
  wire _718_;
  wire _719_;
  wire _720_;
  wire _721_;
  wire _722_;
  wire _723_;
  wire _724_;
  wire _725_;
  wire _726_;
  wire _727_;
  wire _728_;
  wire _729_;
  wire _730_;
  wire _731_;
  wire _732_;
  wire _733_;
  wire _734_;
  wire _735_;
  wire _736_;
  wire _737_;
  wire _738_;
  wire _739_;
  wire _740_;
  wire _741_;
  wire _742_;
  wire _743_;
  wire _744_;
  wire _745_;
  wire _746_;
  wire _747_;
  wire _748_;
  wire _749_;
  wire _750_;
  wire _751_;
  wire _752_;
  wire _753_;
  wire _754_;
  wire _755_;
  wire _756_;
  wire _757_;
  wire _758_;
  wire _759_;
  wire _760_;
  wire _761_;
  wire _762_;
  wire _763_;
  wire _764_;
  wire _765_;
  wire _766_;
  wire _767_;
  wire _768_;
  wire _769_;
  wire _770_;
  wire _771_;
  wire _772_;
  wire _773_;
  wire _774_;
  wire _775_;
  wire _776_;
  wire _777_;
  wire _778_;
  wire _779_;
  wire _780_;
  wire _781_;
  wire _782_;
  wire _783_;
  wire _784_;
  wire _785_;
  wire _786_;
  wire _787_;
  wire _788_;
  wire _789_;
  wire _790_;
  wire _791_;
  wire _792_;
  wire _793_;
  wire _794_;
  wire _795_;
  wire _796_;
  wire _797_;
  wire _798_;
  wire _799_;
  wire _800_;
  wire _801_;
  wire _802_;
  wire _803_;
  wire _804_;
  wire _805_;
  wire _806_;
  wire _807_;
  wire _808_;
  wire _809_;
  wire _810_;
  wire _811_;
  wire _812_;
  wire _813_;
  wire _814_;
  wire _815_;
  wire _816_;
  wire _817_;
  wire _818_;
  wire _819_;
  wire _820_;
  wire _821_;
  wire _822_;
  wire _823_;
  wire _824_;
  wire _825_;
  wire _826_;
  wire _827_;
  wire _828_;
  wire _829_;
  wire _830_;
  wire _831_;
  wire _832_;
  wire _833_;
  wire _834_;
  wire _835_;
  wire _836_;
  wire _837_;
  wire _838_;
  wire _839_;
  wire _840_;
  wire _841_;
  wire _842_;
  wire _843_;
  wire _844_;
  wire _845_;
  wire _846_;
  wire _847_;
  wire _848_;
  wire _849_;
  wire _850_;
  wire _851_;
  wire _852_;
  wire _853_;
  wire _854_;
  wire _855_;
  wire _856_;
  wire _857_;
  wire _858_;
  wire _859_;
  wire _860_;
  wire _861_;
  wire _862_;
  wire _863_;
  wire _864_;
  wire _865_;
  wire _866_;
  wire _867_;
  wire _868_;
  wire _869_;
  wire _870_;
  wire _871_;
  wire _872_;
  wire _873_;
  wire _874_;
  wire _875_;
  wire _876_;
  wire _877_;
  wire _878_;
  wire _879_;
  wire _880_;
  wire _881_;
  wire _882_;
  wire _883_;
  wire _884_;
  wire _885_;
  wire _886_;
  wire _887_;
  wire _888_;
  wire _889_;
  wire _890_;
  wire _891_;
  wire _892_;
  wire _893_;
  wire _894_;
  wire _895_;
  wire _896_;
  wire _897_;
  wire _898_;
  wire _899_;
  wire _900_;
  wire _901_;
  wire _902_;
  wire _903_;
  wire _904_;
  wire _905_;
  wire _906_;
  wire _907_;
  wire _908_;
  wire _909_;
  wire _910_;
  wire _911_;
  wire _912_;
  wire _913_;
  wire _914_;
  wire _915_;
  wire _916_;
  wire _917_;
  wire _918_;
  wire _919_;
  wire _920_;
  wire _921_;
  wire _922_;
  wire _923_;
  wire _924_;
  wire _925_;
  wire _926_;
  wire _927_;
  wire _928_;
  wire _929_;
  wire _930_;
  wire _931_;
  wire _932_;
  wire _933_;
  wire _934_;
  wire _935_;
  wire _936_;
  wire _937_;
  wire _938_;
  wire _939_;
  wire _940_;
  wire _941_;
  wire _942_;
  wire _943_;
  wire _944_;
  wire _945_;
  wire _946_;
  wire _947_;
  wire _948_;
  wire _949_;
  wire _950_;
  wire _951_;
  wire _952_;
  wire _953_;
  wire _954_;
  wire _955_;
  wire _956_;
  wire _957_;
  wire _958_;
  wire _959_;
  wire _960_;
  wire _961_;
  wire _962_;
  wire _963_;
  wire _964_;
  wire _965_;
  wire _966_;
  wire _967_;
  wire _968_;
  wire _969_;
  wire _970_;
  wire _971_;
  wire _972_;
  wire _973_;
  wire _974_;
  wire _975_;
  wire _976_;
  wire _977_;
  wire _978_;
  wire _979_;
  wire _980_;
  wire _981_;
  wire _982_;
  wire _983_;
  wire _984_;
  wire _985_;
  wire _986_;
  wire _987_;
  wire _988_;
  wire _989_;
  wire _990_;
  wire _991_;
  wire _992_;
  wire _993_;
  wire _994_;
  wire _995_;
  wire _996_;
  wire _997_;
  wire _998_;
  wire _999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire _1601_;
  wire _1602_;
  wire _1603_;
  wire _1604_;
  wire _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire _1611_;
  wire _1612_;
  wire _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire _1629_;
  wire _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire _1720_;
  wire _1721_;
  wire _1722_;
  wire _1723_;
  wire _1724_;
  wire _1725_;
  wire _1726_;
  wire _1727_;
  wire _1728_;
  wire _1729_;
  wire _1730_;
  wire _1731_;
  wire _1732_;
  wire _1733_;
  wire _1734_;
  wire _1735_;
  wire _1736_;
  wire _1737_;
  wire _1738_;
  wire _1739_;
  wire _1740_;
  wire _1741_;
  wire _1742_;
  wire _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire _1751_;
  wire _1752_;
  wire _1753_;
  wire _1754_;
  wire _1755_;
  wire _1756_;
  wire _1757_;
  wire _1758_;
  wire _1759_;
  wire _1760_;
  wire _1761_;
  wire _1762_;
  wire _1763_;
  wire _1764_;
  wire _1765_;
  wire _1766_;
  wire _1767_;
  wire _1768_;
  wire _1769_;
  wire _1770_;
  wire _1771_;
  wire _1772_;
  wire _1773_;
  wire _1774_;
  wire _1775_;
  wire _1776_;
  wire _1777_;
  wire _1778_;
  wire _1779_;
  wire _1780_;
  wire _1781_;
  wire _1782_;
  wire _1783_;
  wire _1784_;
  wire _1785_;
  wire _1786_;
  wire _1787_;
  wire _1788_;
  wire _1789_;
  wire _1790_;
  wire _1791_;
  wire _1792_;
  wire _1793_;
  wire _1794_;
  wire _1795_;
  wire _1796_;
  wire _1797_;
  wire _1798_;
  wire _1799_;
  wire _1800_;
  wire _1801_;
  wire _1802_;
  wire _1803_;
  wire _1804_;
  wire _1805_;
  wire _1806_;
  wire _1807_;
  wire _1808_;
  wire _1809_;
  wire _1810_;
  wire _1811_;
  wire _1812_;
  wire _1813_;
  wire _1814_;
  wire _1815_;
  wire _1816_;
  wire _1817_;
  wire _1818_;
  wire _1819_;
  wire _1820_;
  wire _1821_;
  wire _1822_;
  wire _1823_;
  wire _1824_;
  wire _1825_;
  wire _1826_;
  wire _1827_;
  wire _1828_;
  wire _1829_;
  wire _1830_;
  wire _1831_;
  wire _1832_;
  wire _1833_;
  wire _1834_;
  wire _1835_;
  wire _1836_;
  wire _1837_;
  wire _1838_;
  wire _1839_;
  wire _1840_;
  wire _1841_;
  wire _1842_;
  wire _1843_;
  wire _1844_;
  wire _1845_;
  wire _1846_;
  wire _1847_;
  wire _1848_;
  wire _1849_;
  wire _1850_;
  wire _1851_;
  wire _1852_;
  wire _1853_;
  wire _1854_;
  wire _1855_;
  wire _1856_;
  wire _1857_;
  wire _1858_;
  wire _1859_;
  wire _1860_;
  wire _1861_;
  wire _1862_;
  wire _1863_;
  wire _1864_;
  wire _1865_;
  wire _1866_;
  wire _1867_;
  wire _1868_;
  wire _1869_;
  wire _1870_;
  wire _1871_;
  wire _1872_;
  wire _1873_;
  wire _1874_;
  wire _1875_;
  wire _1876_;
  wire _1877_;
  wire _1878_;
  wire _1879_;
  wire _1880_;
  wire _1881_;
  wire _1882_;
  wire _1883_;
  wire _1884_;
  wire _1885_;
  wire _1886_;
  wire _1887_;
  wire _1888_;
  wire _1889_;
  wire _1890_;
  wire _1891_;
  wire _1892_;
  wire _1893_;
  wire _1894_;
  wire _1895_;
  wire _1896_;
  wire _1897_;
  wire _1898_;
  wire _1899_;
  wire _1900_;
  wire _1901_;
  wire _1902_;
  wire _1903_;
  wire _1904_;
  wire _1905_;
  wire _1906_;
  wire _1907_;
  wire _1908_;
  wire _1909_;
  wire _1910_;
  wire _1911_;
  wire _1912_;
  wire _1913_;
  wire _1914_;
  wire _1915_;
  wire _1916_;
  wire _1917_;
  wire _1918_;
  wire _1919_;
  wire _1920_;
  wire _1921_;
  wire _1922_;
  wire _1923_;
  wire _1924_;
  wire _1925_;
  wire _1926_;
  wire _1927_;
  wire _1928_;
  wire _1929_;
  wire _1930_;
  wire _1931_;
  wire _1932_;
  wire _1933_;
  wire _1934_;
  wire _1935_;
  wire _1936_;
  wire _1937_;
  wire _1938_;
  wire _1939_;
  wire _1940_;
  wire _1941_;
  wire _1942_;
  wire _1943_;
  wire _1944_;
  wire _1945_;
  wire _1946_;
  wire _1947_;
  wire _1948_;
  wire _1949_;
  wire _1950_;
  wire _1951_;
  wire _1952_;
  wire _1953_;
  wire _1954_;
  wire _1955_;
  wire _1956_;
  wire _1957_;
  wire _1958_;
  wire _1959_;
  wire _1960_;
  wire _1961_;
  wire _1962_;
  wire _1963_;
  wire _1964_;
  wire _1965_;
  wire _1966_;
  wire _1967_;
  wire _1968_;
  wire _1969_;
  wire _1970_;
  wire _1971_;
  wire _1972_;
  wire _1973_;
  wire _1974_;
  wire _1975_;
  wire _1976_;
  wire _1977_;
  wire _1978_;
  wire _1979_;
  wire _1980_;
  wire _1981_;
  wire _1982_;
  wire _1983_;
  wire _1984_;
  wire _1985_;
  wire _1986_;
  wire _1987_;
  wire _1988_;
  wire _1989_;
  wire _1990_;
  wire _1991_;
  wire _1992_;
  wire _1993_;
  wire _1994_;
  wire _1995_;
  wire _1996_;
  wire _1997_;
  wire _1998_;
  wire _1999_;
  wire _2000_;
  wire _2001_;
  wire _2002_;
  wire _2003_;
  wire _2004_;
  wire _2005_;
  wire _2006_;
  wire _2007_;
  wire _2008_;
  wire _2009_;
  wire _2010_;
  wire _2011_;
  wire _2012_;
  wire _2013_;
  wire _2014_;
  wire _2015_;
  wire _2016_;
  wire _2017_;
  wire _2018_;
  wire _2019_;
  wire _2020_;
  wire _2021_;
  wire _2022_;
  wire _2023_;
  wire _2024_;
  wire _2025_;
  wire _2026_;
  wire _2027_;
  wire _2028_;
  wire _2029_;
  wire _2030_;
  wire _2031_;
  wire _2032_;
  wire _2033_;
  wire _2034_;
  wire _2035_;
  wire _2036_;
  wire _2037_;
  wire _2038_;
  wire _2039_;
  wire _2040_;
  wire _2041_;
  wire _2042_;
  wire _2043_;
  wire _2044_;
  wire _2045_;
  wire _2046_;
  wire _2047_;
  wire _2048_;
  wire _2049_;
  wire _2050_;
  wire _2051_;
  wire _2052_;
  wire _2053_;
  wire _2054_;
  wire _2055_;
  wire _2056_;
  wire _2057_;
  wire _2058_;
  wire _2059_;
  wire _2060_;
  wire _2061_;
  wire _2062_;
  wire _2063_;
  wire _2064_;
  wire _2065_;
  wire _2066_;
  wire _2067_;
  wire _2068_;
  wire _2069_;
  wire _2070_;
  wire _2071_;
  wire _2072_;
  wire _2073_;
  wire _2074_;
  wire _2075_;
  wire _2076_;
  wire _2077_;
  wire _2078_;
  wire _2079_;
  wire _2080_;
  wire _2081_;
  wire _2082_;
  wire _2083_;
  wire _2084_;
  wire _2085_;
  wire _2086_;
  wire _2087_;
  wire _2088_;
  wire _2089_;
  wire _2090_;
  wire _2091_;
  wire _2092_;
  wire _2093_;
  wire _2094_;
  wire _2095_;
  wire _2096_;
  wire _2097_;
  wire _2098_;
  wire _2099_;
  wire _2100_;
  wire _2101_;
  wire _2102_;
  wire _2103_;
  wire _2104_;
  wire _2105_;
  wire _2106_;
  wire _2107_;
  wire _2108_;
  wire _2109_;
  wire _2110_;
  wire _2111_;
  wire _2112_;
  wire _2113_;
  wire _2114_;
  wire _2115_;
  wire _2116_;
  wire _2117_;
  wire _2118_;
  wire _2119_;
  wire _2120_;
  wire _2121_;
  wire _2122_;
  wire _2123_;
  wire _2124_;
  wire _2125_;
  wire _2126_;
  wire _2127_;
  wire _2128_;
  wire _2129_;
  wire _2130_;
  wire _2131_;
  wire _2132_;
  wire _2133_;
  wire _2134_;
  wire _2135_;
  wire _2136_;
  wire _2137_;
  wire _2138_;
  wire _2139_;
  wire _2140_;
  wire _2141_;
  wire _2142_;
  wire _2143_;
  wire _2144_;
  wire _2145_;
  wire _2146_;
  wire _2147_;
  wire _2148_;
  wire _2149_;
  wire _2150_;
  wire _2151_;
  wire _2152_;
  wire _2153_;
  wire _2154_;
  wire _2155_;
  wire _2156_;
  wire _2157_;
  wire _2158_;
  wire _2159_;
  wire _2160_;
  wire _2161_;
  wire _2162_;
  wire _2163_;
  wire _2164_;
  wire _2165_;
  wire _2166_;
  wire _2167_;
  wire _2168_;
  wire _2169_;
  wire _2170_;
  wire _2171_;
  wire _2172_;
  wire _2173_;
  wire _2174_;
  wire _2175_;
  wire _2176_;
  wire _2177_;
  wire _2178_;
  wire _2179_;
  wire _2180_;
  wire _2181_;
  wire _2182_;
  wire _2183_;
  wire _2184_;
  wire _2185_;
  wire _2186_;
  wire _2187_;
  wire _2188_;
  wire _2189_;
  wire _2190_;
  wire _2191_;
  wire _2192_;
  wire _2193_;
  wire _2194_;
  wire _2195_;
  wire _2196_;
  wire _2197_;
  wire _2198_;
  wire _2199_;
  wire _2200_;
  wire _2201_;
  wire _2202_;
  wire _2203_;
  wire _2204_;
  wire _2205_;
  wire _2206_;
  wire _2207_;
  wire _2208_;
  wire _2209_;
  wire _2210_;
  wire _2211_;
  wire _2212_;
  wire _2213_;
  wire _2214_;
  wire _2215_;
  wire _2216_;
  wire _2217_;
  wire _2218_;
  wire _2219_;
  wire _2220_;
  wire _2221_;
  wire _2222_;
  wire _2223_;
  wire _2224_;
  wire _2225_;
  wire _2226_;
  wire _2227_;
  wire _2228_;
  wire _2229_;
  wire _2230_;
  wire _2231_;
  wire _2232_;
  wire _2233_;
  wire _2234_;
  wire _2235_;
  wire _2236_;
  wire _2237_;
  wire _2238_;
  wire _2239_;
  wire _2240_;
  wire _2241_;
  wire _2242_;
  wire _2243_;
  wire _2244_;
  wire _2245_;
  wire _2246_;
  wire _2247_;
  wire _2248_;
  wire _2249_;
  wire _2250_;
  wire _2251_;
  wire _2252_;
  wire _2253_;
  wire _2254_;
  wire _2255_;
  wire _2256_;
  wire _2257_;
  wire _2258_;
  wire _2259_;
  wire _2260_;
  wire _2261_;
  wire _2262_;
  wire _2263_;
  wire _2264_;
  wire _2265_;
  wire _2266_;
  wire _2267_;
  wire _2268_;
  wire _2269_;
  wire _2270_;
  wire _2271_;
  wire _2272_;
  wire _2273_;
  wire _2274_;
  wire _2275_;
  wire _2276_;
  wire _2277_;
  wire _2278_;
  wire _2279_;
  wire _2280_;
  wire _2281_;
  wire _2282_;
  wire _2283_;
  wire _2284_;
  wire _2285_;
  wire _2286_;
  wire _2287_;
  wire _2288_;
  wire _2289_;
  wire _2290_;
  wire _2291_;
  wire _2292_;
  wire _2293_;
  wire _2294_;
  wire _2295_;
  wire _2296_;
  wire _2297_;
  wire _2298_;
  wire _2299_;
  wire _2300_;
  wire _2301_;
  wire _2302_;
  wire _2303_;
  wire _2304_;
  wire _2305_;
  wire _2306_;
  wire _2307_;
  wire _2308_;
  wire _2309_;
  wire _2310_;
  wire _2311_;
  wire _2312_;
  wire _2313_;
  wire _2314_;
  wire _2315_;
  wire _2316_;
  wire _2317_;
  wire _2318_;
  wire _2319_;
  wire _2320_;
  wire _2321_;
  wire _2322_;
  wire _2323_;
  wire _2324_;
  wire _2325_;
  wire _2326_;
  wire _2327_;
  wire _2328_;
  wire _2329_;
  wire _2330_;
  wire _2331_;
  wire _2332_;
  wire _2333_;
  wire _2334_;
  wire _2335_;
  wire _2336_;
  wire _2337_;
  wire _2338_;
  wire _2339_;
  wire _2340_;
  wire _2341_;
  wire _2342_;
  wire _2343_;
  wire _2344_;
  wire _2345_;
  wire _2346_;
  wire _2347_;
  wire _2348_;
  wire _2349_;
  wire _2350_;
  wire _2351_;
  wire _2352_;
  wire _2353_;
  wire _2354_;
  wire _2355_;
  wire _2356_;
  wire _2357_;
  wire _2358_;
  wire _2359_;
  wire _2360_;
  wire _2361_;
  wire _2362_;
  wire _2363_;
  wire _2364_;
  wire _2365_;
  wire _2366_;
  wire _2367_;
  wire _2368_;
  wire _2369_;
  wire _2370_;
  wire _2371_;
  wire _2372_;
  wire _2373_;
  wire _2374_;
  wire _2375_;
  wire _2376_;
  wire _2377_;
  wire _2378_;
  wire _2379_;
  wire _2380_;
  wire _2381_;
  wire _2382_;
  wire _2383_;
  wire _2384_;
  wire _2385_;
  wire _2386_;
  wire _2387_;
  wire _2388_;
  wire _2389_;
  wire _2390_;
  wire _2391_;
  wire _2392_;
  wire _2393_;
  wire _2394_;
  wire _2395_;
  wire _2396_;
  wire _2397_;
  wire _2398_;
  wire _2399_;
  wire _2400_;
  wire _2401_;
  wire _2402_;
  wire _2403_;
  wire _2404_;
  wire _2405_;
  wire _2406_;
  wire _2407_;
  wire _2408_;
  wire _2409_;
  wire _2410_;
  wire _2411_;
  wire _2412_;
  wire _2413_;
  wire _2414_;
  wire _2415_;
  wire _2416_;
  wire _2417_;
  wire _2418_;
  wire _2419_;
  wire _2420_;
  wire _2421_;
  wire _2422_;
  wire _2423_;
  wire _2424_;
  wire _2425_;
  wire _2426_;
  wire _2427_;
  wire _2428_;
  wire _2429_;
  wire _2430_;
  wire _2431_;
  wire _2432_;
  wire _2433_;
  wire _2434_;
  wire _2435_;
  wire _2436_;
  wire _2437_;
  wire _2438_;
  wire _2439_;
  wire _2440_;
  wire _2441_;
  wire _2442_;
  wire _2443_;
  wire _2444_;
  wire _2445_;
  wire _2446_;
  wire _2447_;
  wire _2448_;
  wire _2449_;
  wire _2450_;
  wire _2451_;
  wire _2452_;
  wire _2453_;
  wire _2454_;
  wire _2455_;
  wire _2456_;
  wire _2457_;
  wire _2458_;
  wire _2459_;
  wire _2460_;
  wire _2461_;
  wire _2462_;
  wire _2463_;
  wire _2464_;
  wire _2465_;
  wire _2466_;
  wire _2467_;
  wire _2468_;
  wire _2469_;
  wire _2470_;
  wire _2471_;
  wire _2472_;
  wire _2473_;
  wire _2474_;
  wire _2475_;
  wire _2476_;
  wire _2477_;
  wire _2478_;
  wire _2479_;
  wire _2480_;
  wire _2481_;
  wire _2482_;
  wire _2483_;
  wire _2484_;
  wire _2485_;
  wire _2486_;
  wire _2487_;
  wire _2488_;
  wire _2489_;
  wire _2490_;
  wire _2491_;
  wire _2492_;
  wire _2493_;
  wire _2494_;
  wire _2495_;
  wire _2496_;
  wire _2497_;
  wire _2498_;
  wire _2499_;
  wire _2500_;
  wire _2501_;
  wire _2502_;
  wire _2503_;
  wire _2504_;
  wire _2505_;
  wire _2506_;
  wire _2507_;
  wire _2508_;
  wire _2509_;
  wire _2510_;
  wire _2511_;
  wire _2512_;
  wire _2513_;
  wire _2514_;
  wire _2515_;
  wire _2516_;
  wire _2517_;
  wire _2518_;
  wire _2519_;
  wire _2520_;
  wire _2521_;
  wire _2522_;
  wire _2523_;
  wire _2524_;
  wire _2525_;
  wire _2526_;
  wire _2527_;
  wire _2528_;
  wire _2529_;
  wire _2530_;
  wire _2531_;
  wire _2532_;
  wire _2533_;
  wire _2534_;
  wire _2535_;
  wire _2536_;
  wire _2537_;
  wire _2538_;
  wire _2539_;
  wire _2540_;
  wire _2541_;
  wire _2542_;
  wire _2543_;
  wire _2544_;
  wire _2545_;
  wire _2546_;
  wire _2547_;
  wire _2548_;
  wire _2549_;
  wire _2550_;
  wire _2551_;
  wire _2552_;
  wire _2553_;
  wire _2554_;
  wire _2555_;
  wire _2556_;
  wire _2557_;
  wire _2558_;
  wire _2559_;
  wire _2560_;
  wire _2561_;
  wire _2562_;
  wire _2563_;
  wire _2564_;
  wire _2565_;
  wire _2566_;
  wire _2567_;
  wire _2568_;
  wire _2569_;
  wire _2570_;
  wire _2571_;
  wire _2572_;
  wire _2573_;
  wire _2574_;
  wire _2575_;
  wire _2576_;
  wire _2577_;
  wire _2578_;
  wire _2579_;
  wire _2580_;
  wire _2581_;
  wire _2582_;
  wire _2583_;
  wire _2584_;
  wire _2585_;
  wire _2586_;
  wire _2587_;
  wire _2588_;
  wire _2589_;
  wire _2590_;
  wire _2591_;
  wire _2592_;
  wire _2593_;
  wire _2594_;
  wire _2595_;
  wire _2596_;
  wire _2597_;
  wire _2598_;
  wire _2599_;
  wire _2600_;
  wire _2601_;
  wire _2602_;
  wire _2603_;
  wire _2604_;
  wire _2605_;
  wire _2606_;
  wire _2607_;
  wire _2608_;
  wire _2609_;
  wire _2610_;
  wire _2611_;
  wire _2612_;
  wire _2613_;
  wire _2614_;
  wire _2615_;
  wire _2616_;
  wire _2617_;
  wire _2618_;
  wire _2619_;
  wire _2620_;
  wire _2621_;
  wire _2622_;
  wire _2623_;
  wire _2624_;
  wire _2625_;
  wire _2626_;
  wire _2627_;
  wire _2628_;
  wire _2629_;
  wire _2630_;
  wire _2631_;
  wire _2632_;
  wire _2633_;
  wire _2634_;
  wire _2635_;
  wire _2636_;
  wire _2637_;
  wire _2638_;
  wire _2639_;
  wire _2640_;
  wire _2641_;
  wire _2642_;
  wire _2643_;
  wire _2644_;
  wire _2645_;
  wire _2646_;
  wire _2647_;
  wire _2648_;
  wire _2649_;
  wire _2650_;
  wire _2651_;
  wire _2652_;
  wire _2653_;
  wire _2654_;
  wire _2655_;
  wire _2656_;
  wire _2657_;
  wire _2658_;
  wire _2659_;
  wire _2660_;
  wire _2661_;
  wire _2662_;
  wire _2663_;
  wire _2664_;
  wire _2665_;
  wire _2666_;
  wire _2667_;
  wire _2668_;
  wire _2669_;
  wire _2670_;
  wire _2671_;
  wire _2672_;
  wire _2673_;
  wire _2674_;
  wire _2675_;
  wire _2676_;
  wire _2677_;
  wire _2678_;
  wire _2679_;
  wire _2680_;
  wire _2681_;
  wire _2682_;
  wire _2683_;
  wire _2684_;
  wire _2685_;
  wire _2686_;
  wire _2687_;
  wire _2688_;
  wire _2689_;
  wire _2690_;
  wire _2691_;
  wire _2692_;
  wire _2693_;
  wire _2694_;
  wire _2695_;
  wire _2696_;
  wire _2697_;
  wire _2698_;
  wire _2699_;
  wire _2700_;
  wire _2701_;
  wire _2702_;
  wire _2703_;
  wire _2704_;
  wire _2705_;
  wire _2706_;
  wire _2707_;
  wire _2708_;
  wire _2709_;
  wire _2710_;
  wire _2711_;
  wire _2712_;
  wire _2713_;
  wire _2714_;
  wire _2715_;
  wire _2716_;
  wire _2717_;
  wire _2718_;
  wire _2719_;
  wire _2720_;
  wire _2721_;
  wire _2722_;
  wire _2723_;
  wire _2724_;
  wire _2725_;
  wire _2726_;
  wire _2727_;
  wire _2728_;
  wire _2729_;
  wire _2730_;
  wire _2731_;
  wire _2732_;
  wire _2733_;
  wire _2734_;
  wire _2735_;
  wire _2736_;
  wire _2737_;
  wire _2738_;
  wire _2739_;
  wire _2740_;
  wire _2741_;
  wire _2742_;
  wire _2743_;
  wire _2744_;
  wire _2745_;
  wire _2746_;
  wire _2747_;
  wire _2748_;
  wire _2749_;
  wire _2750_;
  wire _2751_;
  wire _2752_;
  wire _2753_;
  wire _2754_;
  wire _2755_;
  wire _2756_;
  wire _2757_;
  wire _2758_;
  wire _2759_;
  wire _2760_;
  wire _2761_;
  wire _2762_;
  wire _2763_;
  wire _2764_;
  wire _2765_;
  wire _2766_;
  wire _2767_;
  wire _2768_;
  wire _2769_;
  wire _2770_;
  wire _2771_;
  wire _2772_;
  wire _2773_;
  wire _2774_;
  wire _2775_;
  wire _2776_;
  wire _2777_;
  wire _2778_;
  wire _2779_;
  wire _2780_;
  wire _2781_;
  wire _2782_;
  wire _2783_;
  wire _2784_;
  wire _2785_;
  wire _2786_;
  wire _2787_;
  wire _2788_;
  wire _2789_;
  wire _2790_;
  wire _2791_;
  wire _2792_;
  wire _2793_;
  wire _2794_;
  wire _2795_;
  wire _2796_;
  wire _2797_;
  wire _2798_;
  wire _2799_;
  wire _2800_;
  wire _2801_;
  wire _2802_;
  wire _2803_;
  wire _2804_;
  wire _2805_;
  wire _2806_;
  wire _2807_;
  wire _2808_;
  wire _2809_;
  wire _2810_;
  wire _2811_;
  wire _2812_;
  wire _2813_;
  wire _2814_;
  wire _2815_;
  wire _2816_;
  wire _2817_;
  wire _2818_;
  wire _2819_;
  wire _2820_;
  wire _2821_;
  wire _2822_;
  wire _2823_;
  wire _2824_;
  wire _2825_;
  wire _2826_;
  wire _2827_;
  wire _2828_;
  wire _2829_;
  wire _2830_;
  wire _2831_;
  wire _2832_;
  wire _2833_;
  wire _2834_;
  wire _2835_;
  wire _2836_;
  wire _2837_;
  wire _2838_;
  wire _2839_;
  wire _2840_;
  wire _2841_;
  wire _2842_;
  wire _2843_;
  wire _2844_;
  wire _2845_;
  wire _2846_;
  wire _2847_;
  wire _2848_;
  wire _2849_;
  wire _2850_;
  wire _2851_;
  wire _2852_;
  wire _2853_;
  wire _2854_;
  wire _2855_;
  wire _2856_;
  wire _2857_;
  wire _2858_;
  wire _2859_;
  wire _2860_;
  wire _2861_;
  wire _2862_;
  wire _2863_;
  wire _2864_;
  wire _2865_;
  wire _2866_;
  wire _2867_;
  wire _2868_;
  wire _2869_;
  wire _2870_;
  wire _2871_;
  wire _2872_;
  wire _2873_;
  wire _2874_;
  wire _2875_;
  wire _2876_;
  wire _2877_;
  wire _2878_;
  wire _2879_;
  wire _2880_;
  wire _2881_;
  wire _2882_;
  wire _2883_;
  wire _2884_;
  wire _2885_;
  wire _2886_;
  wire _2887_;
  wire _2888_;
  wire _2889_;
  wire _2890_;
  wire _2891_;
  wire _2892_;
  wire _2893_;
  wire _2894_;
  wire _2895_;
  wire _2896_;
  wire _2897_;
  wire _2898_;
  wire _2899_;
  wire _2900_;
  wire _2901_;
  wire _2902_;
  wire _2903_;
  wire _2904_;
  wire _2905_;
  wire _2906_;
  wire _2907_;
  wire _2908_;
  wire _2909_;
  wire _2910_;
  wire _2911_;
  wire _2912_;
  wire _2913_;
  wire _2914_;
  wire _2915_;
  wire _2916_;
  wire _2917_;
  wire _2918_;
  wire _2919_;
  wire _2920_;
  wire _2921_;
  wire _2922_;
  wire _2923_;
  wire _2924_;
  wire _2925_;
  wire _2926_;
  wire _2927_;
  wire _2928_;
  wire _2929_;
  wire _2930_;
  wire _2931_;
  wire _2932_;
  wire _2933_;
  wire _2934_;
  wire _2935_;
  wire _2936_;
  wire _2937_;
  wire _2938_;
  wire _2939_;
  wire _2940_;
  wire _2941_;
  wire _2942_;
  wire _2943_;
  wire _2944_;
  wire _2945_;
  wire _2946_;
  wire _2947_;
  wire _2948_;
  wire _2949_;
  wire _2950_;
  wire _2951_;
  wire _2952_;
  wire _2953_;
  wire _2954_;
  wire _2955_;
  wire _2956_;
  wire _2957_;
  wire _2958_;
  wire _2959_;
  wire _2960_;
  wire _2961_;
  wire _2962_;
  wire _2963_;
  wire _2964_;
  wire _2965_;
  wire _2966_;
  wire _2967_;
  wire _2968_;
  wire _2969_;
  wire _2970_;
  wire _2971_;
  wire _2972_;
  wire _2973_;
  wire _2974_;
  wire _2975_;
  wire _2976_;
  wire _2977_;
  wire _2978_;
  wire _2979_;
  wire _2980_;
  wire _2981_;
  wire _2982_;
  wire _2983_;
  wire _2984_;
  wire _2985_;
  wire _2986_;
  wire _2987_;
  wire _2988_;
  wire _2989_;
  wire _2990_;
  wire _2991_;
  wire _2992_;
  wire _2993_;
  wire _2994_;
  wire _2995_;
  wire _2996_;
  wire _2997_;
  wire _2998_;
  wire _2999_;
  wire _3000_;
  wire _3001_;
  wire _3002_;
  wire _3003_;
  wire _3004_;
  wire _3005_;
  wire _3006_;
  wire _3007_;
  wire _3008_;
  wire _3009_;
  wire _3010_;
  wire _3011_;
  wire _3012_;
  wire _3013_;
  wire _3014_;
  wire _3015_;
  wire _3016_;
  wire _3017_;
  wire _3018_;
  wire _3019_;
  wire _3020_;
  wire _3021_;
  wire _3022_;
  wire _3023_;
  wire _3024_;
  wire _3025_;
  wire _3026_;
  wire _3027_;
  wire _3028_;
  wire _3029_;
  wire _3030_;
  wire _3031_;
  wire _3032_;
  wire _3033_;
  wire _3034_;
  wire _3035_;
  wire _3036_;
  wire _3037_;
  wire _3038_;
  wire _3039_;
  wire _3040_;
  wire _3041_;
  wire _3042_;
  wire _3043_;
  wire _3044_;
  wire _3045_;
  wire _3046_;
  wire _3047_;
  wire _3048_;
  wire _3049_;
  wire _3050_;
  wire _3051_;
  wire _3052_;
  wire _3053_;
  wire _3054_;
  wire _3055_;
  wire _3056_;
  wire _3057_;
  wire _3058_;
  wire _3059_;
  wire _3060_;
  wire _3061_;
  wire _3062_;
  wire _3063_;
  wire _3064_;
  wire _3065_;
  wire _3066_;
  wire _3067_;
  wire _3068_;
  wire _3069_;
  wire _3070_;
  wire _3071_;
  wire _3072_;
  wire _3073_;
  wire _3074_;
  wire _3075_;
  wire _3076_;
  wire _3077_;
  wire _3078_;
  wire _3079_;
  wire _3080_;
  wire _3081_;
  wire _3082_;
  wire _3083_;
  wire _3084_;
  wire _3085_;
  wire _3086_;
  wire _3087_;
  wire _3088_;
  wire _3089_;
  wire _3090_;
  wire _3091_;
  wire _3092_;
  wire _3093_;
  wire _3094_;
  wire _3095_;
  wire _3096_;
  wire _3097_;
  wire _3098_;
  wire _3099_;
  wire _3100_;
  wire _3101_;
  wire _3102_;
  wire _3103_;
  wire _3104_;
  wire _3105_;
  wire _3106_;
  wire _3107_;
  wire _3108_;
  wire _3109_;
  wire _3110_;
  wire _3111_;
  wire _3112_;
  wire _3113_;
  wire _3114_;
  wire _3115_;
  wire _3116_;
  wire _3117_;
  wire _3118_;
  wire _3119_;
  wire _3120_;
  wire _3121_;
  wire _3122_;
  wire _3123_;
  wire _3124_;
  wire _3125_;
  wire _3126_;
  wire _3127_;
  wire _3128_;
  wire _3129_;
  wire _3130_;
  wire _3131_;
  wire _3132_;
  wire _3133_;
  wire _3134_;
  wire _3135_;
  wire _3136_;
  wire _3137_;
  wire _3138_;
  wire _3139_;
  wire _3140_;
  wire _3141_;
  wire _3142_;
  wire _3143_;
  wire _3144_;
  wire _3145_;
  wire _3146_;
  wire _3147_;
  wire _3148_;
  wire _3149_;
  wire _3150_;
  wire _3151_;
  wire _3152_;
  wire _3153_;
  wire _3154_;
  wire _3155_;
  wire _3156_;
  wire _3157_;
  wire _3158_;
  wire _3159_;
  wire _3160_;
  wire _3161_;
  wire _3162_;
  wire _3163_;
  wire _3164_;
  wire _3165_;
  wire _3166_;
  wire _3167_;
  wire _3168_;
  wire _3169_;
  wire _3170_;
  wire _3171_;
  wire _3172_;
  wire _3173_;
  wire _3174_;
  wire _3175_;
  wire _3176_;
  wire _3177_;
  wire _3178_;
  wire _3179_;
  wire _3180_;
  wire _3181_;
  wire _3182_;
  wire _3183_;
  wire _3184_;
  wire _3185_;
  wire _3186_;
  wire _3187_;
  wire _3188_;
  wire _3189_;
  wire _3190_;
  wire _3191_;
  wire _3192_;
  wire _3193_;
  wire _3194_;
  wire _3195_;
  wire _3196_;
  wire _3197_;
  wire _3198_;
  wire _3199_;
  wire _3200_;
  wire _3201_;
  wire _3202_;
  wire _3203_;
  wire _3204_;
  wire _3205_;
  wire _3206_;
  wire _3207_;
  wire _3208_;
  wire _3209_;
  wire _3210_;
  wire _3211_;
  wire _3212_;
  wire _3213_;
  wire _3214_;
  wire _3215_;
  wire _3216_;
  wire _3217_;
  wire _3218_;
  wire _3219_;
  wire _3220_;
  wire _3221_;
  wire _3222_;
  wire _3223_;
  wire _3224_;
  wire _3225_;
  wire _3226_;
  wire _3227_;
  wire _3228_;
  wire _3229_;
  wire _3230_;
  wire _3231_;
  wire _3232_;
  wire _3233_;
  wire _3234_;
  wire _3235_;
  wire _3236_;
  wire _3237_;
  wire _3238_;
  wire _3239_;
  wire _3240_;
  wire _3241_;
  wire _3242_;
  wire _3243_;
  wire _3244_;
  wire _3245_;
  wire _3246_;
  wire _3247_;
  wire _3248_;
  wire _3249_;
  wire _3250_;
  wire _3251_;
  wire _3252_;
  wire _3253_;
  wire _3254_;
  wire _3255_;
  wire _3256_;
  wire _3257_;
  wire _3258_;
  wire _3259_;
  wire _3260_;
  wire _3261_;
  wire _3262_;
  wire _3263_;
  wire _3264_;
  wire _3265_;
  wire _3266_;
  wire _3267_;
  wire _3268_;
  wire _3269_;
  wire _3270_;
  wire _3271_;
  wire _3272_;
  wire _3273_;
  wire _3274_;
  wire _3275_;
  wire _3276_;
  wire _3277_;
  wire _3278_;
  wire _3279_;
  wire _3280_;
  wire _3281_;
  wire _3282_;
  wire _3283_;
  wire _3284_;
  wire _3285_;
  wire _3286_;
  wire _3287_;
  wire _3288_;
  wire _3289_;
  wire _3290_;
  wire _3291_;
  wire _3292_;
  wire _3293_;
  wire _3294_;
  wire _3295_;
  wire _3296_;
  wire _3297_;
  wire _3298_;
  wire _3299_;
  wire _3300_;
  wire _3301_;
  wire _3302_;
  wire _3303_;
  wire _3304_;
  wire _3305_;
  wire _3306_;
  wire _3307_;
  wire _3308_;
  wire _3309_;
  wire _3310_;
  wire _3311_;
  wire _3312_;
  wire _3313_;
  wire _3314_;
  wire _3315_;
  wire _3316_;
  wire _3317_;
  wire _3318_;
  wire _3319_;
  wire _3320_;
  wire _3321_;
  wire _3322_;
  wire _3323_;
  wire _3324_;
  wire _3325_;
  wire _3326_;
  wire _3327_;
  wire _3328_;
  wire _3329_;
  wire _3330_;
  wire _3331_;
  wire _3332_;
  wire _3333_;
  wire _3334_;
  wire _3335_;
  wire _3336_;
  wire _3337_;
  wire _3338_;
  wire _3339_;
  wire _3340_;
  wire _3341_;
  wire _3342_;
  wire _3343_;
  wire _3344_;
  wire _3345_;
  wire _3346_;
  wire _3347_;
  wire _3348_;
  wire _3349_;
  wire _3350_;
  wire _3351_;
  wire _3352_;
  wire _3353_;
  wire _3354_;
  wire _3355_;
  wire _3356_;
  wire _3357_;
  wire _3358_;
  wire _3359_;
  wire _3360_;
  wire _3361_;
  wire _3362_;
  wire _3363_;
  wire _3364_;
  wire _3365_;
  wire _3366_;
  wire _3367_;
  wire _3368_;
  wire _3369_;
  wire _3370_;
  wire _3371_;
  wire _3372_;
  wire _3373_;
  wire _3374_;
  wire _3375_;
  wire _3376_;
  wire _3377_;
  wire _3378_;
  wire _3379_;
  wire _3380_;
  wire _3381_;
  wire _3382_;
  wire _3383_;
  wire _3384_;
  wire _3385_;
  wire _3386_;
  wire _3387_;
  wire _3388_;
  wire _3389_;
  wire _3390_;
  wire _3391_;
  wire _3392_;
  wire _3393_;
  wire _3394_;
  wire _3395_;
  wire _3396_;
  wire _3397_;
  wire _3398_;
  wire _3399_;
  wire _3400_;
  wire _3401_;
  wire _3402_;
  wire _3403_;
  wire _3404_;
  wire _3405_;
  wire _3406_;
  wire _3407_;
  wire _3408_;
  wire _3409_;
  wire _3410_;
  wire _3411_;
  wire _3412_;
  wire _3413_;
  wire _3414_;
  wire _3415_;
  wire _3416_;
  wire _3417_;
  wire _3418_;
  wire _3419_;
  wire _3420_;
  wire _3421_;
  wire _3422_;
  wire _3423_;
  wire _3424_;
  wire _3425_;
  wire _3426_;
  wire _3427_;
  wire _3428_;
  wire _3429_;
  wire _3430_;
  wire _3431_;
  wire _3432_;
  wire _3433_;
  wire _3434_;
  wire _3435_;
  wire _3436_;
  wire _3437_;
  wire _3438_;
  wire _3439_;
  wire _3440_;
  wire _3441_;
  wire _3442_;
  wire _3443_;
  wire _3444_;
  wire _3445_;
  wire _3446_;
  wire _3447_;
  wire _3448_;
  wire _3449_;
  wire _3450_;
  wire _3451_;
  wire _3452_;
  wire _3453_;
  wire _3454_;
  wire _3455_;
  wire _3456_;
  wire _3457_;
  wire _3458_;
  wire _3459_;
  wire _3460_;
  wire _3461_;
  wire _3462_;
  wire _3463_;
  wire _3464_;
  wire _3465_;
  wire _3466_;
  wire _3467_;
  wire _3468_;
  wire _3469_;
  wire _3470_;
  wire _3471_;
  wire _3472_;
  wire _3473_;
  wire _3474_;
  wire _3475_;
  wire _3476_;
  wire _3477_;
  wire _3478_;
  wire _3479_;
  wire _3480_;
  wire _3481_;
  wire _3482_;
  wire _3483_;
  wire _3484_;
  wire _3485_;
  wire _3486_;
  wire _3487_;
  wire _3488_;
  wire _3489_;
  wire _3490_;
  wire _3491_;
  wire _3492_;
  wire _3493_;
  wire _3494_;
  wire _3495_;
  wire _3496_;
  wire _3497_;
  wire _3498_;
  wire _3499_;
  wire _3500_;
  wire _3501_;
  wire _3502_;
  wire _3503_;
  wire _3504_;
  wire _3505_;
  wire _3506_;
  wire _3507_;
  wire _3508_;
  wire _3509_;
  wire _3510_;
  wire _3511_;
  wire _3512_;
  wire _3513_;
  wire _3514_;
  wire _3515_;
  wire _3516_;
  wire _3517_;
  wire _3518_;
  wire _3519_;
  wire _3520_;
  wire _3521_;
  wire _3522_;
  wire _3523_;
  wire _3524_;
  wire _3525_;
  wire _3526_;
  wire _3527_;
  wire _3528_;
  wire _3529_;
  wire _3530_;
  wire _3531_;
  wire _3532_;
  wire _3533_;
  wire _3534_;
  wire _3535_;
  wire _3536_;
  wire _3537_;
  wire _3538_;
  wire _3539_;
  wire _3540_;
  wire _3541_;
  wire _3542_;
  wire _3543_;
  wire _3544_;
  wire _3545_;
  wire _3546_;
  wire _3547_;
  wire _3548_;
  wire _3549_;
  wire _3550_;
  wire _3551_;
  wire _3552_;
  wire _3553_;
  wire _3554_;
  wire _3555_;
  wire _3556_;
  wire _3557_;
  wire _3558_;
  wire _3559_;
  wire _3560_;
  wire _3561_;
  wire _3562_;
  wire _3563_;
  wire _3564_;
  wire _3565_;
  wire _3566_;
  wire _3567_;
  wire _3568_;
  wire _3569_;
  wire _3570_;
  wire _3571_;
  wire _3572_;
  wire _3573_;
  wire _3574_;
  wire _3575_;
  wire _3576_;
  wire _3577_;
  wire _3578_;
  wire _3579_;
  wire _3580_;
  wire _3581_;
  wire _3582_;
  wire _3583_;
  wire _3584_;
  wire _3585_;
  wire _3586_;
  wire _3587_;
  wire _3588_;
  wire _3589_;
  wire _3590_;
  wire _3591_;
  wire _3592_;
  wire _3593_;
  wire _3594_;
  wire _3595_;
  wire _3596_;
  wire _3597_;
  wire _3598_;
  wire _3599_;
  wire _3600_;
  wire _3601_;
  wire _3602_;
  wire _3603_;
  wire _3604_;
  wire _3605_;
  wire _3606_;
  wire _3607_;
  wire _3608_;
  wire _3609_;
  wire _3610_;
  wire _3611_;
  wire _3612_;
  wire _3613_;
  wire _3614_;
  wire _3615_;
  wire _3616_;
  wire _3617_;
  wire _3618_;
  wire _3619_;
  wire _3620_;
  wire _3621_;
  wire _3622_;
  wire _3623_;
  wire _3624_;
  wire _3625_;
  wire _3626_;
  wire _3627_;
  wire _3628_;
  wire _3629_;
  wire _3630_;
  wire _3631_;
  wire _3632_;
  wire _3633_;
  wire _3634_;
  wire _3635_;
  wire _3636_;
  wire _3637_;
  wire _3638_;
  wire _3639_;
  wire _3640_;
  wire _3641_;
  wire _3642_;
  wire _3643_;
  wire _3644_;
  wire _3645_;
  wire _3646_;
  wire _3647_;
  wire _3648_;
  wire _3649_;
  wire _3650_;
  wire _3651_;
  wire _3652_;
  wire _3653_;
  wire _3654_;
  wire _3655_;
  wire _3656_;
  wire _3657_;
  wire _3658_;
  wire _3659_;
  wire _3660_;
  wire _3661_;
  wire _3662_;
  wire _3663_;
  wire _3664_;
  wire _3665_;
  wire _3666_;
  wire _3667_;
  wire _3668_;
  wire _3669_;
  wire _3670_;
  wire _3671_;
  wire _3672_;
  wire _3673_;
  wire _3674_;
  wire _3675_;
  wire _3676_;
  wire _3677_;
  wire _3678_;
  wire _3679_;
  wire _3680_;
  wire _3681_;
  wire _3682_;
  wire _3683_;
  wire _3684_;
  wire _3685_;
  wire _3686_;
  wire _3687_;
  wire _3688_;
  wire _3689_;
  wire _3690_;
  wire _3691_;
  wire _3692_;
  wire _3693_;
  wire _3694_;
  wire _3695_;
  wire _3696_;
  wire _3697_;
  wire _3698_;
  wire _3699_;
  wire _3700_;
  wire _3701_;
  wire _3702_;
  wire _3703_;
  wire _3704_;
  wire _3705_;
  wire _3706_;
  wire _3707_;
  wire _3708_;
  wire _3709_;
  wire _3710_;
  wire _3711_;
  wire _3712_;
  wire _3713_;
  wire _3714_;
  wire _3715_;
  wire _3716_;
  wire _3717_;
  wire _3718_;
  wire _3719_;
  wire _3720_;
  wire _3721_;
  wire _3722_;
  wire _3723_;
  wire _3724_;
  wire _3725_;
  wire _3726_;
  wire _3727_;
  wire _3728_;
  wire _3729_;
  wire _3730_;
  wire _3731_;
  wire _3732_;
  wire _3733_;
  wire _3734_;
  wire _3735_;
  wire _3736_;
  wire _3737_;
  wire _3738_;
  wire _3739_;
  wire _3740_;
  wire _3741_;
  wire _3742_;
  wire _3743_;
  wire _3744_;
  wire _3745_;
  wire _3746_;
  wire _3747_;
  wire _3748_;
  wire _3749_;
  wire _3750_;
  wire _3751_;
  wire _3752_;
  wire _3753_;
  wire _3754_;
  wire _3755_;
  wire _3756_;
  wire _3757_;
  wire _3758_;
  wire _3759_;
  wire _3760_;
  wire _3761_;
  wire _3762_;
  wire _3763_;
  wire _3764_;
  wire _3765_;
  wire _3766_;
  wire _3767_;
  wire _3768_;
  wire _3769_;
  wire _3770_;
  wire _3771_;
  wire _3772_;
  wire _3773_;
  wire _3774_;
  wire _3775_;
  wire _3776_;
  wire _3777_;
  wire _3778_;
  wire _3779_;
  wire _3780_;
  wire _3781_;
  wire _3782_;
  wire _3783_;
  wire _3784_;
  wire _3785_;
  wire _3786_;
  wire _3787_;
  wire _3788_;
  wire _3789_;
  wire _3790_;
  wire _3791_;
  wire _3792_;
  wire _3793_;
  wire _3794_;
  wire _3795_;
  wire _3796_;
  wire _3797_;
  wire _3798_;
  wire _3799_;
  wire _3800_;
  wire _3801_;
  wire _3802_;
  wire _3803_;
  wire _3804_;
  wire _3805_;
  wire _3806_;
  wire _3807_;
  wire _3808_;
  wire _3809_;
  wire _3810_;
  wire _3811_;
  wire _3812_;
  wire _3813_;
  wire _3814_;
  wire _3815_;
  wire _3816_;
  wire _3817_;
  wire _3818_;
  wire _3819_;
  wire _3820_;
  wire _3821_;
  wire _3822_;
  wire _3823_;
  wire _3824_;
  wire _3825_;
  wire _3826_;
  wire _3827_;
  wire _3828_;
  wire _3829_;
  wire _3830_;
  wire _3831_;
  wire _3832_;
  wire _3833_;
  wire _3834_;
  wire _3835_;
  wire _3836_;
  wire _3837_;
  wire _3838_;
  wire _3839_;
  wire _3840_;
  wire _3841_;
  wire _3842_;
  wire _3843_;
  wire _3844_;
  wire _3845_;
  wire _3846_;
  wire _3847_;
  wire _3848_;
  wire _3849_;
  wire _3850_;
  wire _3851_;
  wire _3852_;
  wire _3853_;
  wire _3854_;
  wire _3855_;
  wire _3856_;
  wire _3857_;
  wire _3858_;
  wire _3859_;
  wire _3860_;
  wire _3861_;
  wire _3862_;
  wire _3863_;
  wire _3864_;
  wire _3865_;
  wire _3866_;
  wire _3867_;
  wire _3868_;
  wire _3869_;
  wire _3870_;
  wire _3871_;
  wire _3872_;
  wire _3873_;
  wire _3874_;
  wire _3875_;
  wire _3876_;
  wire _3877_;
  wire _3878_;
  wire _3879_;
  wire _3880_;
  wire _3881_;
  wire _3882_;
  wire _3883_;
  wire _3884_;
  wire _3885_;
  wire _3886_;
  wire _3887_;
  wire _3888_;
  wire _3889_;
  wire _3890_;
  wire _3891_;
  wire _3892_;
  wire _3893_;
  wire _3894_;
  wire _3895_;
  wire _3896_;
  wire _3897_;
  wire _3898_;
  wire _3899_;
  wire _3900_;
  wire _3901_;
  wire _3902_;
  wire _3903_;
  wire _3904_;
  wire _3905_;
  wire _3906_;
  wire _3907_;
  wire _3908_;
  wire _3909_;
  wire _3910_;
  wire _3911_;
  wire _3912_;
  wire _3913_;
  wire _3914_;
  wire _3915_;
  wire _3916_;
  wire _3917_;
  wire _3918_;
  wire _3919_;
  wire _3920_;
  wire _3921_;
  wire _3922_;
  wire _3923_;
  wire _3924_;
  wire _3925_;
  wire _3926_;
  wire _3927_;
  wire _3928_;
  wire _3929_;
  wire _3930_;
  wire _3931_;
  wire _3932_;
  wire _3933_;
  wire _3934_;
  wire _3935_;
  wire _3936_;
  wire _3937_;
  wire _3938_;
  wire _3939_;
  wire _3940_;
  wire _3941_;
  wire _3942_;
  wire _3943_;
  wire _3944_;
  wire _3945_;
  wire _3946_;
  wire _3947_;
  wire _3948_;
  wire _3949_;
  wire _3950_;
  wire _3951_;
  wire _3952_;
  wire _3953_;
  wire _3954_;
  wire _3955_;
  wire _3956_;
  wire _3957_;
  wire _3958_;
  wire _3959_;
  wire _3960_;
  wire _3961_;
  wire _3962_;
  wire _3963_;
  wire _3964_;
  wire _3965_;
  wire _3966_;
  wire _3967_;
  wire _3968_;
  wire _3969_;
  wire _3970_;
  wire _3971_;
  wire _3972_;
  wire _3973_;
  wire _3974_;
  wire _3975_;
  wire _3976_;
  wire _3977_;
  wire _3978_;
  wire _3979_;
  wire _3980_;
  wire _3981_;
  wire _3982_;
  wire _3983_;
  wire _3984_;
  wire _3985_;
  wire _3986_;
  wire _3987_;
  wire _3988_;
  wire _3989_;
  wire _3990_;
  wire _3991_;
  wire _3992_;
  wire _3993_;
  wire _3994_;
  wire _3995_;
  wire _3996_;
  wire _3997_;
  wire _3998_;
  wire _3999_;
  wire _4000_;
  wire _4001_;
  wire _4002_;
  wire _4003_;
  wire _4004_;
  wire _4005_;
  wire _4006_;
  wire _4007_;
  wire _4008_;
  wire _4009_;
  wire _4010_;
  wire _4011_;
  wire _4012_;
  wire _4013_;
  wire _4014_;
  wire _4015_;
  wire _4016_;
  wire _4017_;
  wire _4018_;
  wire _4019_;
  wire _4020_;
  wire _4021_;
  wire _4022_;
  wire _4023_;
  wire _4024_;
  wire _4025_;
  wire _4026_;
  wire _4027_;
  wire _4028_;
  wire _4029_;
  wire _4030_;
  wire _4031_;
  wire _4032_;
  wire _4033_;
  wire _4034_;
  wire _4035_;
  wire _4036_;
  wire _4037_;
  wire _4038_;
  wire _4039_;
  wire _4040_;
  wire _4041_;
  wire _4042_;
  wire _4043_;
  wire _4044_;
  wire _4045_;
  wire _4046_;
  wire _4047_;
  wire _4048_;
  wire _4049_;
  wire _4050_;
  wire _4051_;
  wire _4052_;
  wire _4053_;
  wire _4054_;
  wire _4055_;
  wire _4056_;
  wire _4057_;
  wire _4058_;
  wire _4059_;
  wire _4060_;
  wire _4061_;
  wire _4062_;
  wire _4063_;
  wire _4064_;
  wire _4065_;
  wire _4066_;
  wire _4067_;
  wire _4068_;
  wire _4069_;
  wire _4070_;
  wire _4071_;
  wire _4072_;
  wire _4073_;
  wire _4074_;
  wire _4075_;
  wire _4076_;
  wire _4077_;
  wire _4078_;
  wire _4079_;
  wire _4080_;
  wire _4081_;
  wire _4082_;
  wire _4083_;
  wire _4084_;
  wire _4085_;
  wire _4086_;
  wire _4087_;
  wire _4088_;
  wire _4089_;
  wire _4090_;
  wire _4091_;
  wire _4092_;
  wire _4093_;
  wire _4094_;
  wire _4095_;
  wire _4096_;
  wire _4097_;
  wire _4098_;
  wire _4099_;
  wire _4100_;
  wire _4101_;
  wire _4102_;
  wire _4103_;
  wire _4104_;
  wire _4105_;
  wire _4106_;
  wire _4107_;
  wire _4108_;
  wire _4109_;
  wire _4110_;
  wire _4111_;
  wire _4112_;
  wire _4113_;
  wire _4114_;
  wire _4115_;
  wire _4116_;
  wire _4117_;
  wire _4118_;
  wire _4119_;
  wire _4120_;
  wire _4121_;
  wire _4122_;
  wire _4123_;
  wire _4124_;
  wire _4125_;
  wire _4126_;
  wire _4127_;
  wire _4128_;
  wire _4129_;
  wire _4130_;
  wire _4131_;
  wire _4132_;
  wire _4133_;
  wire _4134_;
  wire _4135_;
  wire _4136_;
  wire _4137_;
  wire _4138_;
  wire _4139_;
  wire _4140_;
  wire _4141_;
  wire _4142_;
  wire _4143_;
  wire _4144_;
  wire _4145_;
  wire _4146_;
  wire _4147_;
  wire _4148_;
  wire _4149_;
  wire _4150_;
  wire _4151_;
  wire _4152_;
  wire _4153_;
  wire _4154_;
  wire _4155_;
  wire _4156_;
  wire _4157_;
  wire _4158_;
  wire _4159_;
  wire _4160_;
  wire _4161_;
  wire _4162_;
  wire _4163_;
  wire _4164_;
  wire _4165_;
  wire _4166_;
  wire _4167_;
  wire _4168_;
  wire _4169_;
  wire _4170_;
  wire _4171_;
  wire _4172_;
  wire _4173_;
  wire _4174_;
  wire _4175_;
  wire _4176_;
  wire _4177_;
  wire _4178_;
  wire _4179_;
  wire _4180_;
  wire _4181_;
  wire _4182_;
  wire _4183_;
  wire _4184_;
  wire _4185_;
  wire _4186_;
  wire _4187_;
  wire _4188_;
  wire _4189_;
  wire _4190_;
  wire _4191_;
  wire _4192_;
  wire _4193_;
  wire _4194_;
  wire _4195_;
  wire _4196_;
  wire _4197_;
  wire _4198_;
  wire _4199_;
  wire _4200_;
  wire _4201_;
  wire _4202_;
  wire _4203_;
  wire _4204_;
  wire _4205_;
  wire _4206_;
  wire _4207_;
  wire _4208_;
  wire _4209_;
  wire _4210_;
  wire _4211_;
  wire _4212_;
  wire _4213_;
  wire _4214_;
  wire _4215_;
  wire _4216_;
  wire _4217_;
  wire _4218_;
  wire _4219_;
  wire _4220_;
  wire _4221_;
  wire _4222_;
  wire _4223_;
  wire _4224_;
  wire _4225_;
  wire _4226_;
  wire _4227_;
  wire _4228_;
  wire _4229_;
  wire _4230_;
  wire _4231_;
  wire _4232_;
  wire _4233_;
  wire _4234_;
  wire _4235_;
  wire _4236_;
  wire _4237_;
  wire _4238_;
  wire _4239_;
  wire _4240_;
  wire _4241_;
  wire _4242_;
  wire _4243_;
  wire _4244_;
  wire _4245_;
  wire _4246_;
  wire _4247_;
  wire _4248_;
  wire _4249_;
  wire _4250_;
  wire _4251_;
  wire _4252_;
  wire _4253_;
  wire _4254_;
  wire _4255_;
  wire _4256_;
  wire _4257_;
  wire _4258_;
  wire _4259_;
  wire _4260_;
  wire _4261_;
  wire _4262_;
  wire _4263_;
  wire _4264_;
  wire _4265_;
  wire _4266_;
  wire _4267_;
  wire _4268_;
  wire _4269_;
  wire _4270_;
  wire _4271_;
  wire _4272_;
  wire _4273_;
  wire _4274_;
  wire _4275_;
  wire _4276_;
  wire _4277_;
  wire _4278_;
  wire _4279_;
  wire _4280_;
  wire _4281_;
  wire _4282_;
  wire _4283_;
  wire _4284_;
  wire _4285_;
  wire _4286_;
  wire _4287_;
  wire _4288_;
  wire _4289_;
  wire _4290_;
  wire _4291_;
  wire _4292_;
  wire _4293_;
  wire _4294_;
  wire _4295_;
  wire _4296_;
  wire _4297_;
  wire _4298_;
  wire _4299_;
  wire _4300_;
  wire _4301_;
  wire _4302_;
  wire _4303_;
  wire _4304_;
  wire _4305_;
  wire _4306_;
  wire _4307_;
  wire _4308_;
  wire _4309_;
  wire _4310_;
  wire _4311_;
  wire _4312_;
  wire _4313_;
  wire _4314_;
  wire _4315_;
  wire _4316_;
  wire _4317_;
  wire _4318_;
  wire _4319_;
  wire _4320_;
  wire _4321_;
  wire _4322_;
  wire _4323_;
  wire _4324_;
  wire _4325_;
  wire _4326_;
  wire _4327_;
  wire _4328_;
  wire _4329_;
  wire _4330_;
  wire _4331_;
  wire _4332_;
  wire _4333_;
  wire _4334_;
  wire _4335_;
  wire _4336_;
  wire _4337_;
  wire _4338_;
  wire _4339_;
  wire _4340_;
  wire _4341_;
  wire _4342_;
  wire _4343_;
  wire _4344_;
  wire _4345_;
  wire _4346_;
  wire _4347_;
  wire _4348_;
  wire _4349_;
  wire _4350_;
  wire _4351_;
  wire _4352_;
  wire _4353_;
  wire _4354_;
  wire _4355_;
  wire _4356_;
  wire _4357_;
  wire _4358_;
  wire _4359_;
  wire _4360_;
  wire _4361_;
  wire _4362_;
  wire _4363_;
  wire _4364_;
  wire _4365_;
  wire _4366_;
  wire _4367_;
  wire _4368_;
  wire _4369_;
  wire _4370_;
  wire _4371_;
  wire _4372_;
  wire _4373_;
  wire _4374_;
  wire _4375_;
  wire _4376_;
  wire _4377_;
  wire _4378_;
  wire _4379_;
  wire _4380_;
  wire _4381_;
  wire _4382_;
  wire _4383_;
  wire _4384_;
  wire _4385_;
  wire _4386_;
  wire _4387_;
  wire _4388_;
  wire _4389_;
  wire _4390_;
  wire _4391_;
  wire _4392_;
  wire _4393_;
  wire _4394_;
  wire _4395_;
  wire _4396_;
  wire _4397_;
  wire _4398_;
  wire _4399_;
  wire _4400_;
  wire _4401_;
  wire _4402_;
  wire _4403_;
  wire _4404_;
  wire _4405_;
  wire _4406_;
  wire _4407_;
  wire _4408_;
  wire _4409_;
  wire _4410_;
  wire _4411_;
  wire _4412_;
  wire _4413_;
  wire _4414_;
  wire _4415_;
  wire _4416_;
  wire _4417_;
  wire _4418_;
  wire _4419_;
  wire _4420_;
  wire _4421_;
  wire _4422_;
  wire _4423_;
  wire _4424_;
  wire _4425_;
  wire _4426_;
  wire _4427_;
  wire _4428_;
  wire _4429_;
  wire _4430_;
  wire _4431_;
  wire _4432_;
  wire _4433_;
  wire _4434_;
  wire _4435_;
  wire _4436_;
  wire _4437_;
  wire _4438_;
  wire _4439_;
  wire _4440_;
  wire _4441_;
  wire _4442_;
  wire _4443_;
  wire _4444_;
  wire _4445_;
  wire _4446_;
  wire _4447_;
  wire _4448_;
  wire _4449_;
  wire _4450_;
  wire _4451_;
  wire _4452_;
  wire _4453_;
  wire _4454_;
  wire _4455_;
  wire _4456_;
  wire _4457_;
  wire _4458_;
  wire _4459_;
  wire _4460_;
  wire _4461_;
  wire _4462_;
  wire _4463_;
  wire _4464_;
  wire _4465_;
  wire _4466_;
  wire _4467_;
  wire _4468_;
  wire _4469_;
  wire _4470_;
  wire _4471_;
  wire _4472_;
  wire _4473_;
  wire _4474_;
  wire _4475_;
  wire _4476_;
  wire _4477_;
  wire _4478_;
  wire _4479_;
  wire _4480_;
  wire _4481_;
  wire _4482_;
  wire _4483_;
  wire _4484_;
  wire _4485_;
  wire _4486_;
  wire _4487_;
  wire _4488_;
  wire _4489_;
  wire _4490_;
  wire _4491_;
  wire _4492_;
  wire _4493_;
  wire _4494_;
  wire _4495_;
  wire _4496_;
  wire _4497_;
  wire _4498_;
  wire _4499_;
  wire _4500_;
  wire _4501_;
  wire _4502_;
  wire _4503_;
  wire _4504_;
  wire _4505_;
  wire _4506_;
  wire _4507_;
  wire _4508_;
  wire _4509_;
  wire _4510_;
  wire _4511_;
  wire _4512_;
  wire _4513_;
  wire _4514_;
  wire _4515_;
  wire _4516_;
  wire _4517_;
  wire _4518_;
  wire _4519_;
  wire _4520_;
  wire _4521_;
  wire _4522_;
  wire _4523_;
  wire _4524_;
  wire _4525_;
  wire _4526_;
  wire _4527_;
  wire _4528_;
  wire _4529_;
  wire _4530_;
  wire _4531_;
  wire _4532_;
  wire _4533_;
  wire _4534_;
  wire _4535_;
  wire _4536_;
  wire _4537_;
  wire _4538_;
  wire _4539_;
  wire _4540_;
  wire _4541_;
  wire _4542_;
  wire _4543_;
  wire _4544_;
  wire _4545_;
  wire _4546_;
  wire _4547_;
  wire _4548_;
  wire _4549_;
  wire _4550_;
  wire _4551_;
  wire _4552_;
  wire _4553_;
  wire _4554_;
  wire _4555_;
  wire _4556_;
  wire _4557_;
  wire _4558_;
  wire _4559_;
  wire _4560_;
  wire _4561_;
  wire _4562_;
  wire _4563_;
  wire _4564_;
  wire _4565_;
  wire _4566_;
  wire _4567_;
  wire _4568_;
  wire _4569_;
  wire _4570_;
  wire _4571_;
  wire _4572_;
  wire _4573_;
  wire _4574_;
  wire _4575_;
  wire _4576_;
  wire _4577_;
  wire _4578_;
  wire _4579_;
  wire _4580_;
  wire _4581_;
  wire _4582_;
  wire _4583_;
  wire _4584_;
  wire _4585_;
  wire _4586_;
  wire _4587_;
  wire _4588_;
  wire _4589_;
  wire _4590_;
  wire _4591_;
  wire _4592_;
  wire _4593_;
  wire _4594_;
  wire _4595_;
  wire _4596_;
  wire _4597_;
  wire _4598_;
  wire _4599_;
  wire _4600_;
  wire _4601_;
  wire _4602_;
  wire _4603_;
  wire _4604_;
  wire _4605_;
  wire _4606_;
  wire _4607_;
  wire _4608_;
  wire _4609_;
  wire _4610_;
  wire _4611_;
  wire _4612_;
  wire _4613_;
  wire _4614_;
  wire _4615_;
  wire _4616_;
  wire _4617_;
  wire _4618_;
  wire _4619_;
  wire _4620_;
  wire _4621_;
  wire _4622_;
  wire _4623_;
  wire _4624_;
  wire _4625_;
  wire _4626_;
  wire _4627_;
  wire _4628_;
  wire _4629_;
  wire _4630_;
  wire _4631_;
  wire _4632_;
  wire _4633_;
  wire _4634_;
  wire _4635_;
  wire _4636_;
  wire _4637_;
  wire _4638_;
  wire _4639_;
  wire _4640_;
  wire _4641_;
  wire _4642_;
  wire _4643_;
  wire _4644_;
  wire _4645_;
  wire _4646_;
  wire _4647_;
  wire _4648_;
  wire _4649_;
  wire _4650_;
  wire _4651_;
  wire _4652_;
  wire _4653_;
  wire _4654_;
  wire _4655_;
  wire _4656_;
  wire _4657_;
  wire _4658_;
  wire _4659_;
  wire _4660_;
  wire _4661_;
  wire _4662_;
  wire _4663_;
  wire _4664_;
  wire _4665_;
  wire _4666_;
  wire _4667_;
  wire _4668_;
  wire _4669_;
  wire _4670_;
  wire _4671_;
  wire _4672_;
  wire _4673_;
  wire _4674_;
  wire _4675_;
  wire _4676_;
  wire _4677_;
  wire _4678_;
  wire _4679_;
  wire _4680_;
  wire _4681_;
  wire _4682_;
  wire _4683_;
  wire _4684_;
  wire _4685_;
  wire _4686_;
  wire _4687_;
  wire _4688_;
  wire _4689_;
  wire _4690_;
  wire _4691_;
  wire _4692_;
  wire _4693_;
  wire _4694_;
  wire _4695_;
  wire _4696_;
  wire _4697_;
  wire _4698_;
  wire _4699_;
  wire _4700_;
  wire _4701_;
  wire _4702_;
  wire _4703_;
  wire _4704_;
  wire _4705_;
  wire _4706_;
  wire _4707_;
  wire _4708_;
  wire _4709_;
  wire _4710_;
  wire _4711_;
  wire _4712_;
  wire _4713_;
  wire _4714_;
  wire _4715_;
  wire _4716_;
  wire _4717_;
  wire _4718_;
  wire _4719_;
  wire _4720_;
  wire _4721_;
  wire _4722_;
  wire _4723_;
  wire _4724_;
  wire _4725_;
  wire _4726_;
  wire _4727_;
  wire _4728_;
  wire _4729_;
  wire _4730_;
  wire _4731_;
  wire _4732_;
  wire _4733_;
  wire _4734_;
  wire _4735_;
  wire _4736_;
  wire _4737_;
  wire _4738_;
  wire _4739_;
  wire _4740_;
  wire _4741_;
  wire _4742_;
  wire _4743_;
  wire _4744_;
  wire _4745_;
  wire _4746_;
  wire _4747_;
  wire _4748_;
  wire _4749_;
  wire _4750_;
  wire _4751_;
  wire _4752_;
  wire _4753_;
  wire _4754_;
  wire _4755_;
  wire _4756_;
  wire _4757_;
  wire _4758_;
  wire _4759_;
  wire _4760_;
  wire _4761_;
  wire _4762_;
  wire _4763_;
  wire _4764_;
  wire _4765_;
  wire _4766_;
  wire _4767_;
  wire _4768_;
  wire _4769_;
  wire _4770_;
  wire _4771_;
  wire _4772_;
  wire _4773_;
  wire _4774_;
  wire _4775_;
  wire _4776_;
  wire _4777_;
  wire _4778_;
  wire _4779_;
  wire _4780_;
  wire _4781_;
  wire _4782_;
  wire _4783_;
  wire _4784_;
  wire _4785_;
  wire _4786_;
  wire _4787_;
  wire _4788_;
  wire _4789_;
  wire _4790_;
  wire _4791_;
  wire _4792_;
  wire _4793_;
  wire _4794_;
  wire _4795_;
  wire _4796_;
  wire _4797_;
  wire _4798_;
  wire _4799_;
  wire _4800_;
  wire _4801_;
  wire _4802_;
  wire _4803_;
  wire _4804_;
  wire _4805_;
  wire _4806_;
  wire _4807_;
  wire _4808_;
  wire _4809_;
  wire _4810_;
  wire _4811_;
  wire _4812_;
  wire _4813_;
  wire _4814_;
  wire _4815_;
  wire _4816_;
  wire _4817_;
  wire _4818_;
  wire _4819_;
  wire _4820_;
  wire _4821_;
  wire _4822_;
  wire _4823_;
  wire _4824_;
  wire _4825_;
  wire _4826_;
  wire _4827_;
  wire _4828_;
  wire _4829_;
  wire _4830_;
  wire _4831_;
  wire _4832_;
  wire _4833_;
  wire _4834_;
  wire _4835_;
  wire _4836_;
  wire _4837_;
  wire _4838_;
  wire _4839_;
  wire _4840_;
  wire _4841_;
  wire _4842_;
  wire _4843_;
  wire _4844_;
  wire _4845_;
  wire _4846_;
  wire _4847_;
  wire _4848_;
  wire _4849_;
  wire _4850_;
  wire _4851_;
  wire _4852_;
  wire _4853_;
  wire _4854_;
  wire _4855_;
  wire _4856_;
  wire _4857_;
  wire _4858_;
  wire _4859_;
  wire _4860_;
  wire _4861_;
  wire _4862_;
  wire _4863_;
  wire _4864_;
  wire _4865_;
  wire _4866_;
  wire _4867_;
  wire _4868_;
  wire _4869_;
  wire _4870_;
  wire _4871_;
  wire _4872_;
  wire _4873_;
  wire _4874_;
  wire _4875_;
  wire _4876_;
  wire _4877_;
  wire _4878_;
  wire _4879_;
  wire _4880_;
  wire _4881_;
  wire _4882_;
  wire _4883_;
  wire _4884_;
  wire _4885_;
  wire _4886_;
  wire _4887_;
  wire _4888_;
  wire _4889_;
  wire _4890_;
  wire _4891_;
  wire _4892_;
  wire _4893_;
  wire _4894_;
  wire _4895_;
  wire _4896_;
  wire _4897_;
  wire _4898_;
  wire _4899_;
  wire _4900_;
  wire _4901_;
  wire _4902_;
  wire _4903_;
  wire _4904_;
  wire _4905_;
  wire _4906_;
  wire _4907_;
  wire _4908_;
  wire _4909_;
  wire _4910_;
  wire _4911_;
  wire _4912_;
  wire _4913_;
  wire _4914_;
  wire _4915_;
  wire _4916_;
  wire _4917_;
  wire _4918_;
  wire _4919_;
  wire _4920_;
  wire _4921_;
  wire _4922_;
  wire _4923_;
  wire _4924_;
  wire _4925_;
  wire _4926_;
  wire _4927_;
  wire _4928_;
  wire _4929_;
  wire _4930_;
  wire _4931_;
  wire _4932_;
  wire _4933_;
  wire _4934_;
  wire _4935_;
  wire _4936_;
  wire _4937_;
  wire _4938_;
  wire _4939_;
  wire _4940_;
  wire _4941_;
  wire _4942_;
  wire _4943_;
  wire _4944_;
  wire _4945_;
  wire _4946_;
  wire _4947_;
  wire _4948_;
  wire _4949_;
  wire _4950_;
  wire _4951_;
  wire _4952_;
  wire _4953_;
  wire _4954_;
  wire _4955_;
  wire _4956_;
  wire _4957_;
  wire _4958_;
  wire _4959_;
  wire _4960_;
  wire _4961_;
  wire _4962_;
  wire _4963_;
  wire _4964_;
  wire _4965_;
  wire _4966_;
  wire _4967_;
  wire _4968_;
  wire _4969_;
  wire _4970_;
  wire _4971_;
  wire _4972_;
  wire _4973_;
  wire _4974_;
  wire _4975_;
  wire _4976_;
  wire _4977_;
  wire _4978_;
  wire _4979_;
  wire _4980_;
  wire _4981_;
  wire _4982_;
  wire _4983_;
  wire _4984_;
  wire _4985_;
  wire _4986_;
  wire _4987_;
  wire _4988_;
  wire _4989_;
  wire _4990_;
  wire _4991_;
  wire _4992_;
  wire _4993_;
  wire _4994_;
  wire _4995_;
  wire _4996_;
  wire _4997_;
  wire _4998_;
  wire _4999_;
  wire _5000_;
  wire _5001_;
  wire _5002_;
  wire _5003_;
  wire _5004_;
  wire _5005_;
  wire _5006_;
  wire _5007_;
  wire _5008_;
  wire _5009_;
  wire _5010_;
  wire _5011_;
  wire _5012_;
  wire _5013_;
  wire _5014_;
  wire _5015_;
  wire _5016_;
  wire _5017_;
  wire _5018_;
  wire _5019_;
  wire _5020_;
  wire _5021_;
  wire _5022_;
  wire _5023_;
  wire _5024_;
  wire _5025_;
  wire _5026_;
  wire _5027_;
  wire _5028_;
  wire _5029_;
  wire _5030_;
  wire _5031_;
  wire _5032_;
  wire _5033_;
  wire _5034_;
  wire _5035_;
  wire _5036_;
  wire _5037_;
  wire _5038_;
  wire _5039_;
  wire _5040_;
  wire _5041_;
  wire _5042_;
  wire _5043_;
  wire _5044_;
  wire _5045_;
  wire _5046_;
  wire _5047_;
  wire _5048_;
  wire _5049_;
  wire _5050_;
  wire _5051_;
  wire _5052_;
  wire _5053_;
  wire _5054_;
  wire _5055_;
  wire [30:0] r_0;
  wire [31:0] r_1;
  wire [31:0] m_1;
  wire [31:0] sum_1;
  wire [30:0] inv_1;
  wire [32:0] r_2;
  wire [32:0] m_2;
  wire [32:0] sum_2;
  wire [31:0] inv_2;
  wire [33:0] r_3;
  wire [33:0] m_3;
  wire [33:0] sum_3;
  wire [32:0] inv_3;
  wire [34:0] r_4;
  wire [34:0] m_4;
  wire [34:0] sum_4;
  wire [33:0] inv_4;
  wire [35:0] r_5;
  wire [35:0] m_5;
  wire [35:0] sum_5;
  wire [34:0] inv_5;
  wire [36:0] r_6;
  wire [36:0] m_6;
  wire [36:0] sum_6;
  wire [35:0] inv_6;
  wire [37:0] r_7;
  wire [37:0] m_7;
  wire [37:0] sum_7;
  wire [36:0] inv_7;
  wire [38:0] r_8;
  wire [38:0] m_8;
  wire [38:0] sum_8;
  wire [37:0] inv_8;
  wire [39:0] r_9;
  wire [39:0] m_9;
  wire [39:0] sum_9;
  wire [38:0] inv_9;
  wire [40:0] r_10;
  wire [40:0] m_10;
  wire [40:0] sum_10;
  wire [39:0] inv_10;
  wire [41:0] r_11;
  wire [41:0] m_11;
  wire [41:0] sum_11;
  wire [40:0] inv_11;
  wire [42:0] r_12;
  wire [42:0] m_12;
  wire [42:0] sum_12;
  wire [41:0] inv_12;
  wire [43:0] r_13;
  wire [43:0] m_13;
  wire [43:0] sum_13;
  wire [42:0] inv_13;
  wire [44:0] r_14;
  wire [44:0] m_14;
  wire [44:0] sum_14;
  wire [43:0] inv_14;
  wire [45:0] r_15;
  wire [45:0] m_15;
  wire [45:0] sum_15;
  wire [44:0] inv_15;
  wire [46:0] r_16;
  wire [46:0] m_16;
  wire [46:0] sum_16;
  wire [45:0] inv_16;
  wire zeroWire;
  wire oneWire;
  input [29:0] rin;
  input [14:0] div;
  output [15:0] q;
  output [46:0] rout;
  assign zeroWire = 1'b0 /*0*/;
  assign oneWire = 1'b1 /*0*/;
  assign r_0[0] = rin[0] /*9168*/;
  assign r_0[1] = rin[1] /*9167*/;
  assign r_0[2] = rin[2] /*9166*/;
  assign r_0[3] = rin[3] /*9165*/;
  assign r_0[4] = rin[4] /*9164*/;
  assign r_0[5] = rin[5] /*9163*/;
  assign r_0[6] = rin[6] /*9162*/;
  assign r_0[7] = rin[7] /*9161*/;
  assign r_0[8] = rin[8] /*9160*/;
  assign r_0[9] = rin[9] /*9159*/;
  assign r_0[10] = rin[10] /*9158*/;
  assign r_0[11] = rin[11] /*9157*/;
  assign r_0[12] = rin[12] /*9156*/;
  assign r_0[13] = rin[13] /*9155*/;
  assign r_0[14] = rin[14] /*9154*/;
  assign r_0[15] = rin[15] /*9153*/;
  assign r_0[16] = rin[16] /*9152*/;
  assign r_0[17] = rin[17] /*9151*/;
  assign r_0[18] = rin[18] /*9150*/;
  assign r_0[19] = rin[19] /*9149*/;
  assign r_0[20] = rin[20] /*9148*/;
  assign r_0[21] = rin[21] /*9147*/;
  assign r_0[22] = rin[22] /*9146*/;
  assign r_0[23] = rin[23] /*9145*/;
  assign r_0[24] = rin[24] /*9144*/;
  assign r_0[25] = rin[25] /*9143*/;
  assign r_0[26] = rin[26] /*9142*/;
  assign r_0[27] = rin[27] /*9141*/;
  assign r_0[28] = rin[28] /*9140*/;
  assign r_0[29] = rin[29] /*9139*/;
  assign r_0[30] = zeroWire /*9138*/;
  assign inv_1[0] = oneWire /*8544*/;
  assign inv_1[1] = oneWire /*8538*/;
  assign inv_1[2] = oneWire /*8532*/;
  assign inv_1[3] = oneWire /*8526*/;
  assign inv_1[4] = oneWire /*8520*/;
  assign inv_1[5] = oneWire /*8514*/;
  assign inv_1[6] = oneWire /*8508*/;
  assign inv_1[7] = oneWire /*8502*/;
  assign inv_1[8] = oneWire /*8496*/;
  assign inv_1[9] = oneWire /*8490*/;
  assign inv_1[10] = oneWire /*8484*/;
  assign inv_1[11] = oneWire /*8478*/;
  assign inv_1[12] = oneWire /*8472*/;
  assign inv_1[13] = oneWire /*8466*/;
  assign inv_1[14] = oneWire /*8460*/;
  assign inv_1[15] = ~div[0] /*8454*/;
  assign inv_1[16] = ~div[1] /*8448*/;
  assign inv_1[17] = ~div[2] /*8442*/;
  assign inv_1[18] = ~div[3] /*8436*/;
  assign inv_1[19] = ~div[4] /*8430*/;
  assign inv_1[20] = ~div[5] /*8424*/;
  assign inv_1[21] = ~div[6] /*8418*/;
  assign inv_1[22] = ~div[7] /*8412*/;
  assign inv_1[23] = ~div[8] /*8406*/;
  assign inv_1[24] = ~div[9] /*8400*/;
  assign inv_1[25] = ~div[10] /*8394*/;
  assign inv_1[26] = ~div[11] /*8388*/;
  assign inv_1[27] = ~div[12] /*8382*/;
  assign inv_1[28] = ~div[13] /*8376*/;
  assign inv_1[29] = ~div[14] /*8370*/;
  assign inv_1[30] = oneWire /*8364*/;
  assign _0_ = inv_1[0] ^ r_0[0] /*8543*/;
  assign sum_1[0] = _0_ ^ oneWire /*8542*/;
  assign _1_ = _0_ & oneWire /*8541*/;
  assign _2_ = inv_1[0] & r_0[0] /*8540*/;
  assign _3_ = _1_ | _2_ /*8539*/;
  assign _4_ = inv_1[1] ^ r_0[1] /*8537*/;
  assign sum_1[1] = _4_ ^ _3_ /*8536*/;
  assign _5_ = _4_ & _3_ /*8535*/;
  assign _6_ = inv_1[1] & r_0[1] /*8534*/;
  assign _7_ = _5_ | _6_ /*8533*/;
  assign _8_ = inv_1[2] ^ r_0[2] /*8531*/;
  assign sum_1[2] = _8_ ^ _7_ /*8530*/;
  assign _9_ = _8_ & _7_ /*8529*/;
  assign _10_ = inv_1[2] & r_0[2] /*8528*/;
  assign _11_ = _9_ | _10_ /*8527*/;
  assign _12_ = inv_1[3] ^ r_0[3] /*8525*/;
  assign sum_1[3] = _12_ ^ _11_ /*8524*/;
  assign _13_ = _12_ & _11_ /*8523*/;
  assign _14_ = inv_1[3] & r_0[3] /*8522*/;
  assign _15_ = _13_ | _14_ /*8521*/;
  assign _16_ = inv_1[4] ^ r_0[4] /*8519*/;
  assign sum_1[4] = _16_ ^ _15_ /*8518*/;
  assign _17_ = _16_ & _15_ /*8517*/;
  assign _18_ = inv_1[4] & r_0[4] /*8516*/;
  assign _19_ = _17_ | _18_ /*8515*/;
  assign _20_ = inv_1[5] ^ r_0[5] /*8513*/;
  assign sum_1[5] = _20_ ^ _19_ /*8512*/;
  assign _21_ = _20_ & _19_ /*8511*/;
  assign _22_ = inv_1[5] & r_0[5] /*8510*/;
  assign _23_ = _21_ | _22_ /*8509*/;
  assign _24_ = inv_1[6] ^ r_0[6] /*8507*/;
  assign sum_1[6] = _24_ ^ _23_ /*8506*/;
  assign _25_ = _24_ & _23_ /*8505*/;
  assign _26_ = inv_1[6] & r_0[6] /*8504*/;
  assign _27_ = _25_ | _26_ /*8503*/;
  assign _28_ = inv_1[7] ^ r_0[7] /*8501*/;
  assign sum_1[7] = _28_ ^ _27_ /*8500*/;
  assign _29_ = _28_ & _27_ /*8499*/;
  assign _30_ = inv_1[7] & r_0[7] /*8498*/;
  assign _31_ = _29_ | _30_ /*8497*/;
  assign _32_ = inv_1[8] ^ r_0[8] /*8495*/;
  assign sum_1[8] = _32_ ^ _31_ /*8494*/;
  assign _33_ = _32_ & _31_ /*8493*/;
  assign _34_ = inv_1[8] & r_0[8] /*8492*/;
  assign _35_ = _33_ | _34_ /*8491*/;
  assign _36_ = inv_1[9] ^ r_0[9] /*8489*/;
  assign sum_1[9] = _36_ ^ _35_ /*8488*/;
  assign _37_ = _36_ & _35_ /*8487*/;
  assign _38_ = inv_1[9] & r_0[9] /*8486*/;
  assign _39_ = _37_ | _38_ /*8485*/;
  assign _40_ = inv_1[10] ^ r_0[10] /*8483*/;
  assign sum_1[10] = _40_ ^ _39_ /*8482*/;
  assign _41_ = _40_ & _39_ /*8481*/;
  assign _42_ = inv_1[10] & r_0[10] /*8480*/;
  assign _43_ = _41_ | _42_ /*8479*/;
  assign _44_ = inv_1[11] ^ r_0[11] /*8477*/;
  assign sum_1[11] = _44_ ^ _43_ /*8476*/;
  assign _45_ = _44_ & _43_ /*8475*/;
  assign _46_ = inv_1[11] & r_0[11] /*8474*/;
  assign _47_ = _45_ | _46_ /*8473*/;
  assign _48_ = inv_1[12] ^ r_0[12] /*8471*/;
  assign sum_1[12] = _48_ ^ _47_ /*8470*/;
  assign _49_ = _48_ & _47_ /*8469*/;
  assign _50_ = inv_1[12] & r_0[12] /*8468*/;
  assign _51_ = _49_ | _50_ /*8467*/;
  assign _52_ = inv_1[13] ^ r_0[13] /*8465*/;
  assign sum_1[13] = _52_ ^ _51_ /*8464*/;
  assign _53_ = _52_ & _51_ /*8463*/;
  assign _54_ = inv_1[13] & r_0[13] /*8462*/;
  assign _55_ = _53_ | _54_ /*8461*/;
  assign _56_ = inv_1[14] ^ r_0[14] /*8459*/;
  assign sum_1[14] = _56_ ^ _55_ /*8458*/;
  assign _57_ = _56_ & _55_ /*8457*/;
  assign _58_ = inv_1[14] & r_0[14] /*8456*/;
  assign _59_ = _57_ | _58_ /*8455*/;
  assign _60_ = inv_1[15] ^ r_0[15] /*8453*/;
  assign sum_1[15] = _60_ ^ _59_ /*8452*/;
  assign _61_ = _60_ & _59_ /*8451*/;
  assign _62_ = inv_1[15] & r_0[15] /*8450*/;
  assign _63_ = _61_ | _62_ /*8449*/;
  assign _64_ = inv_1[16] ^ r_0[16] /*8447*/;
  assign sum_1[16] = _64_ ^ _63_ /*8446*/;
  assign _65_ = _64_ & _63_ /*8445*/;
  assign _66_ = inv_1[16] & r_0[16] /*8444*/;
  assign _67_ = _65_ | _66_ /*8443*/;
  assign _68_ = inv_1[17] ^ r_0[17] /*8441*/;
  assign sum_1[17] = _68_ ^ _67_ /*8440*/;
  assign _69_ = _68_ & _67_ /*8439*/;
  assign _70_ = inv_1[17] & r_0[17] /*8438*/;
  assign _71_ = _69_ | _70_ /*8437*/;
  assign _72_ = inv_1[18] ^ r_0[18] /*8435*/;
  assign sum_1[18] = _72_ ^ _71_ /*8434*/;
  assign _73_ = _72_ & _71_ /*8433*/;
  assign _74_ = inv_1[18] & r_0[18] /*8432*/;
  assign _75_ = _73_ | _74_ /*8431*/;
  assign _76_ = inv_1[19] ^ r_0[19] /*8429*/;
  assign sum_1[19] = _76_ ^ _75_ /*8428*/;
  assign _77_ = _76_ & _75_ /*8427*/;
  assign _78_ = inv_1[19] & r_0[19] /*8426*/;
  assign _79_ = _77_ | _78_ /*8425*/;
  assign _80_ = inv_1[20] ^ r_0[20] /*8423*/;
  assign sum_1[20] = _80_ ^ _79_ /*8422*/;
  assign _81_ = _80_ & _79_ /*8421*/;
  assign _82_ = inv_1[20] & r_0[20] /*8420*/;
  assign _83_ = _81_ | _82_ /*8419*/;
  assign _84_ = inv_1[21] ^ r_0[21] /*8417*/;
  assign sum_1[21] = _84_ ^ _83_ /*8416*/;
  assign _85_ = _84_ & _83_ /*8415*/;
  assign _86_ = inv_1[21] & r_0[21] /*8414*/;
  assign _87_ = _85_ | _86_ /*8413*/;
  assign _88_ = inv_1[22] ^ r_0[22] /*8411*/;
  assign sum_1[22] = _88_ ^ _87_ /*8410*/;
  assign _89_ = _88_ & _87_ /*8409*/;
  assign _90_ = inv_1[22] & r_0[22] /*8408*/;
  assign _91_ = _89_ | _90_ /*8407*/;
  assign _92_ = inv_1[23] ^ r_0[23] /*8405*/;
  assign sum_1[23] = _92_ ^ _91_ /*8404*/;
  assign _93_ = _92_ & _91_ /*8403*/;
  assign _94_ = inv_1[23] & r_0[23] /*8402*/;
  assign _95_ = _93_ | _94_ /*8401*/;
  assign _96_ = inv_1[24] ^ r_0[24] /*8399*/;
  assign sum_1[24] = _96_ ^ _95_ /*8398*/;
  assign _97_ = _96_ & _95_ /*8397*/;
  assign _98_ = inv_1[24] & r_0[24] /*8396*/;
  assign _99_ = _97_ | _98_ /*8395*/;
  assign _100_ = inv_1[25] ^ r_0[25] /*8393*/;
  assign sum_1[25] = _100_ ^ _99_ /*8392*/;
  assign _101_ = _100_ & _99_ /*8391*/;
  assign _102_ = inv_1[25] & r_0[25] /*8390*/;
  assign _103_ = _101_ | _102_ /*8389*/;
  assign _104_ = inv_1[26] ^ r_0[26] /*8387*/;
  assign sum_1[26] = _104_ ^ _103_ /*8386*/;
  assign _105_ = _104_ & _103_ /*8385*/;
  assign _106_ = inv_1[26] & r_0[26] /*8384*/;
  assign _107_ = _105_ | _106_ /*8383*/;
  assign _108_ = inv_1[27] ^ r_0[27] /*8381*/;
  assign sum_1[27] = _108_ ^ _107_ /*8380*/;
  assign _109_ = _108_ & _107_ /*8379*/;
  assign _110_ = inv_1[27] & r_0[27] /*8378*/;
  assign _111_ = _109_ | _110_ /*8377*/;
  assign _112_ = inv_1[28] ^ r_0[28] /*8375*/;
  assign sum_1[28] = _112_ ^ _111_ /*8374*/;
  assign _113_ = _112_ & _111_ /*8373*/;
  assign _114_ = inv_1[28] & r_0[28] /*8372*/;
  assign _115_ = _113_ | _114_ /*8371*/;
  assign _116_ = inv_1[29] ^ r_0[29] /*8369*/;
  assign sum_1[29] = _116_ ^ _115_ /*8368*/;
  assign _117_ = _116_ & _115_ /*8367*/;
  assign _118_ = inv_1[29] & r_0[29] /*8366*/;
  assign _119_ = _117_ | _118_ /*8365*/;
  assign _120_ = inv_1[30] ^ r_0[30] /*8363*/;
  assign sum_1[30] = _120_ ^ _119_ /*8362*/;
  assign _121_ = _120_ & _119_ /*8361*/;
  assign _122_ = inv_1[30] & r_0[30] /*8360*/;
  assign _123_ = _121_ | _122_ /*8359*/;
  assign _124_ = _123_ ^ _119_ /*8358*/;
  assign _125_ = ~_124_ /*8357*/;
  assign _126_ = sum_1[30] & _125_ /*8356*/;
  assign _127_ = _124_ & _123_ /*8355*/;
  assign sum_1[31] = _127_ | _126_ /*8354*/;
  assign q[15] = ~sum_1[31] /*8353*/;
  assign m_1[0] = r_0[0] /*8352*/;
  assign m_1[1] = r_0[1] /*8351*/;
  assign m_1[2] = r_0[2] /*8350*/;
  assign m_1[3] = r_0[3] /*8349*/;
  assign m_1[4] = r_0[4] /*8348*/;
  assign m_1[5] = r_0[5] /*8347*/;
  assign m_1[6] = r_0[6] /*8346*/;
  assign m_1[7] = r_0[7] /*8345*/;
  assign m_1[8] = r_0[8] /*8344*/;
  assign m_1[9] = r_0[9] /*8343*/;
  assign m_1[10] = r_0[10] /*8342*/;
  assign m_1[11] = r_0[11] /*8341*/;
  assign m_1[12] = r_0[12] /*8340*/;
  assign m_1[13] = r_0[13] /*8339*/;
  assign m_1[14] = r_0[14] /*8338*/;
  assign m_1[15] = r_0[15] /*8337*/;
  assign m_1[16] = r_0[16] /*8336*/;
  assign m_1[17] = r_0[17] /*8335*/;
  assign m_1[18] = r_0[18] /*8334*/;
  assign m_1[19] = r_0[19] /*8333*/;
  assign m_1[20] = r_0[20] /*8332*/;
  assign m_1[21] = r_0[21] /*8331*/;
  assign m_1[22] = r_0[22] /*8330*/;
  assign m_1[23] = r_0[23] /*8329*/;
  assign m_1[24] = r_0[24] /*8328*/;
  assign m_1[25] = r_0[25] /*8327*/;
  assign m_1[26] = r_0[26] /*8326*/;
  assign m_1[27] = r_0[27] /*8325*/;
  assign m_1[28] = r_0[28] /*8324*/;
  assign m_1[29] = r_0[29] /*8323*/;
  assign m_1[30] = r_0[30] /*8322*/;
  assign m_1[31] = r_0[30] /*8321*/;
  assign _129_ = ~q[15] /*8320*/;
  assign _130_ = sum_1[0] & q[15] /*8319*/;
  assign _131_ = m_1[0] & _129_ /*8318*/;
  assign r_1[0] = _131_ | _130_ /*8317*/;
  assign _132_ = ~q[15] /*8316*/;
  assign _133_ = sum_1[1] & q[15] /*8315*/;
  assign _134_ = m_1[1] & _132_ /*8314*/;
  assign r_1[1] = _134_ | _133_ /*8313*/;
  assign _135_ = ~q[15] /*8312*/;
  assign _136_ = sum_1[2] & q[15] /*8311*/;
  assign _137_ = m_1[2] & _135_ /*8310*/;
  assign r_1[2] = _137_ | _136_ /*8309*/;
  assign _138_ = ~q[15] /*8308*/;
  assign _139_ = sum_1[3] & q[15] /*8307*/;
  assign _140_ = m_1[3] & _138_ /*8306*/;
  assign r_1[3] = _140_ | _139_ /*8305*/;
  assign _141_ = ~q[15] /*8304*/;
  assign _142_ = sum_1[4] & q[15] /*8303*/;
  assign _143_ = m_1[4] & _141_ /*8302*/;
  assign r_1[4] = _143_ | _142_ /*8301*/;
  assign _144_ = ~q[15] /*8300*/;
  assign _145_ = sum_1[5] & q[15] /*8299*/;
  assign _146_ = m_1[5] & _144_ /*8298*/;
  assign r_1[5] = _146_ | _145_ /*8297*/;
  assign _147_ = ~q[15] /*8296*/;
  assign _148_ = sum_1[6] & q[15] /*8295*/;
  assign _149_ = m_1[6] & _147_ /*8294*/;
  assign r_1[6] = _149_ | _148_ /*8293*/;
  assign _150_ = ~q[15] /*8292*/;
  assign _151_ = sum_1[7] & q[15] /*8291*/;
  assign _152_ = m_1[7] & _150_ /*8290*/;
  assign r_1[7] = _152_ | _151_ /*8289*/;
  assign _153_ = ~q[15] /*8288*/;
  assign _154_ = sum_1[8] & q[15] /*8287*/;
  assign _155_ = m_1[8] & _153_ /*8286*/;
  assign r_1[8] = _155_ | _154_ /*8285*/;
  assign _156_ = ~q[15] /*8284*/;
  assign _157_ = sum_1[9] & q[15] /*8283*/;
  assign _158_ = m_1[9] & _156_ /*8282*/;
  assign r_1[9] = _158_ | _157_ /*8281*/;
  assign _159_ = ~q[15] /*8280*/;
  assign _160_ = sum_1[10] & q[15] /*8279*/;
  assign _161_ = m_1[10] & _159_ /*8278*/;
  assign r_1[10] = _161_ | _160_ /*8277*/;
  assign _162_ = ~q[15] /*8276*/;
  assign _163_ = sum_1[11] & q[15] /*8275*/;
  assign _164_ = m_1[11] & _162_ /*8274*/;
  assign r_1[11] = _164_ | _163_ /*8273*/;
  assign _165_ = ~q[15] /*8272*/;
  assign _166_ = sum_1[12] & q[15] /*8271*/;
  assign _167_ = m_1[12] & _165_ /*8270*/;
  assign r_1[12] = _167_ | _166_ /*8269*/;
  assign _168_ = ~q[15] /*8268*/;
  assign _169_ = sum_1[13] & q[15] /*8267*/;
  assign _170_ = m_1[13] & _168_ /*8266*/;
  assign r_1[13] = _170_ | _169_ /*8265*/;
  assign _171_ = ~q[15] /*8264*/;
  assign _172_ = sum_1[14] & q[15] /*8263*/;
  assign _173_ = m_1[14] & _171_ /*8262*/;
  assign r_1[14] = _173_ | _172_ /*8261*/;
  assign _174_ = ~q[15] /*8260*/;
  assign _175_ = sum_1[15] & q[15] /*8259*/;
  assign _176_ = m_1[15] & _174_ /*8258*/;
  assign r_1[15] = _176_ | _175_ /*8257*/;
  assign _177_ = ~q[15] /*8256*/;
  assign _178_ = sum_1[16] & q[15] /*8255*/;
  assign _179_ = m_1[16] & _177_ /*8254*/;
  assign r_1[16] = _179_ | _178_ /*8253*/;
  assign _180_ = ~q[15] /*8252*/;
  assign _181_ = sum_1[17] & q[15] /*8251*/;
  assign _182_ = m_1[17] & _180_ /*8250*/;
  assign r_1[17] = _182_ | _181_ /*8249*/;
  assign _183_ = ~q[15] /*8248*/;
  assign _184_ = sum_1[18] & q[15] /*8247*/;
  assign _185_ = m_1[18] & _183_ /*8246*/;
  assign r_1[18] = _185_ | _184_ /*8245*/;
  assign _186_ = ~q[15] /*8244*/;
  assign _187_ = sum_1[19] & q[15] /*8243*/;
  assign _188_ = m_1[19] & _186_ /*8242*/;
  assign r_1[19] = _188_ | _187_ /*8241*/;
  assign _189_ = ~q[15] /*8240*/;
  assign _190_ = sum_1[20] & q[15] /*8239*/;
  assign _191_ = m_1[20] & _189_ /*8238*/;
  assign r_1[20] = _191_ | _190_ /*8237*/;
  assign _192_ = ~q[15] /*8236*/;
  assign _193_ = sum_1[21] & q[15] /*8235*/;
  assign _194_ = m_1[21] & _192_ /*8234*/;
  assign r_1[21] = _194_ | _193_ /*8233*/;
  assign _195_ = ~q[15] /*8232*/;
  assign _196_ = sum_1[22] & q[15] /*8231*/;
  assign _197_ = m_1[22] & _195_ /*8230*/;
  assign r_1[22] = _197_ | _196_ /*8229*/;
  assign _198_ = ~q[15] /*8228*/;
  assign _199_ = sum_1[23] & q[15] /*8227*/;
  assign _200_ = m_1[23] & _198_ /*8226*/;
  assign r_1[23] = _200_ | _199_ /*8225*/;
  assign _201_ = ~q[15] /*8224*/;
  assign _202_ = sum_1[24] & q[15] /*8223*/;
  assign _203_ = m_1[24] & _201_ /*8222*/;
  assign r_1[24] = _203_ | _202_ /*8221*/;
  assign _204_ = ~q[15] /*8220*/;
  assign _205_ = sum_1[25] & q[15] /*8219*/;
  assign _206_ = m_1[25] & _204_ /*8218*/;
  assign r_1[25] = _206_ | _205_ /*8217*/;
  assign _207_ = ~q[15] /*8216*/;
  assign _208_ = sum_1[26] & q[15] /*8215*/;
  assign _209_ = m_1[26] & _207_ /*8214*/;
  assign r_1[26] = _209_ | _208_ /*8213*/;
  assign _210_ = ~q[15] /*8212*/;
  assign _211_ = sum_1[27] & q[15] /*8211*/;
  assign _212_ = m_1[27] & _210_ /*8210*/;
  assign r_1[27] = _212_ | _211_ /*8209*/;
  assign _213_ = ~q[15] /*8208*/;
  assign _214_ = sum_1[28] & q[15] /*8207*/;
  assign _215_ = m_1[28] & _213_ /*8206*/;
  assign r_1[28] = _215_ | _214_ /*8205*/;
  assign _216_ = ~q[15] /*8204*/;
  assign _217_ = sum_1[29] & q[15] /*8203*/;
  assign _218_ = m_1[29] & _216_ /*8202*/;
  assign r_1[29] = _218_ | _217_ /*8201*/;
  assign _219_ = ~q[15] /*8200*/;
  assign _220_ = sum_1[30] & q[15] /*8199*/;
  assign _221_ = m_1[30] & _219_ /*8198*/;
  assign r_1[30] = _221_ | _220_ /*8197*/;
  assign _222_ = ~q[15] /*8196*/;
  assign _223_ = sum_1[31] & q[15] /*8195*/;
  assign _224_ = m_1[31] & _222_ /*8194*/;
  assign r_1[31] = _224_ | _223_ /*8193*/;
  assign inv_2[0] = oneWire /*8012*/;
  assign inv_2[1] = oneWire /*8006*/;
  assign inv_2[2] = oneWire /*8000*/;
  assign inv_2[3] = oneWire /*7994*/;
  assign inv_2[4] = oneWire /*7988*/;
  assign inv_2[5] = oneWire /*7982*/;
  assign inv_2[6] = oneWire /*7976*/;
  assign inv_2[7] = oneWire /*7970*/;
  assign inv_2[8] = oneWire /*7964*/;
  assign inv_2[9] = oneWire /*7958*/;
  assign inv_2[10] = oneWire /*7952*/;
  assign inv_2[11] = oneWire /*7946*/;
  assign inv_2[12] = oneWire /*7940*/;
  assign inv_2[13] = oneWire /*7934*/;
  assign inv_2[14] = ~div[0] /*7928*/;
  assign inv_2[15] = ~div[1] /*7922*/;
  assign inv_2[16] = ~div[2] /*7916*/;
  assign inv_2[17] = ~div[3] /*7910*/;
  assign inv_2[18] = ~div[4] /*7904*/;
  assign inv_2[19] = ~div[5] /*7898*/;
  assign inv_2[20] = ~div[6] /*7892*/;
  assign inv_2[21] = ~div[7] /*7886*/;
  assign inv_2[22] = ~div[8] /*7880*/;
  assign inv_2[23] = ~div[9] /*7874*/;
  assign inv_2[24] = ~div[10] /*7868*/;
  assign inv_2[25] = ~div[11] /*7862*/;
  assign inv_2[26] = ~div[12] /*7856*/;
  assign inv_2[27] = ~div[13] /*7850*/;
  assign inv_2[28] = ~div[14] /*7844*/;
  assign inv_2[29] = oneWire /*7838*/;
  assign inv_2[30] = oneWire /*7832*/;
  assign inv_2[31] = oneWire /*7826*/;
  assign _225_ = inv_2[0] ^ r_1[0] /*8011*/;
  assign sum_2[0] = _225_ ^ oneWire /*8010*/;
  assign _226_ = _225_ & oneWire /*8009*/;
  assign _227_ = inv_2[0] & r_1[0] /*8008*/;
  assign _228_ = _226_ | _227_ /*8007*/;
  assign _229_ = inv_2[1] ^ r_1[1] /*8005*/;
  assign sum_2[1] = _229_ ^ _228_ /*8004*/;
  assign _230_ = _229_ & _228_ /*8003*/;
  assign _231_ = inv_2[1] & r_1[1] /*8002*/;
  assign _232_ = _230_ | _231_ /*8001*/;
  assign _233_ = inv_2[2] ^ r_1[2] /*7999*/;
  assign sum_2[2] = _233_ ^ _232_ /*7998*/;
  assign _234_ = _233_ & _232_ /*7997*/;
  assign _235_ = inv_2[2] & r_1[2] /*7996*/;
  assign _236_ = _234_ | _235_ /*7995*/;
  assign _237_ = inv_2[3] ^ r_1[3] /*7993*/;
  assign sum_2[3] = _237_ ^ _236_ /*7992*/;
  assign _238_ = _237_ & _236_ /*7991*/;
  assign _239_ = inv_2[3] & r_1[3] /*7990*/;
  assign _240_ = _238_ | _239_ /*7989*/;
  assign _241_ = inv_2[4] ^ r_1[4] /*7987*/;
  assign sum_2[4] = _241_ ^ _240_ /*7986*/;
  assign _242_ = _241_ & _240_ /*7985*/;
  assign _243_ = inv_2[4] & r_1[4] /*7984*/;
  assign _244_ = _242_ | _243_ /*7983*/;
  assign _245_ = inv_2[5] ^ r_1[5] /*7981*/;
  assign sum_2[5] = _245_ ^ _244_ /*7980*/;
  assign _246_ = _245_ & _244_ /*7979*/;
  assign _247_ = inv_2[5] & r_1[5] /*7978*/;
  assign _248_ = _246_ | _247_ /*7977*/;
  assign _249_ = inv_2[6] ^ r_1[6] /*7975*/;
  assign sum_2[6] = _249_ ^ _248_ /*7974*/;
  assign _250_ = _249_ & _248_ /*7973*/;
  assign _251_ = inv_2[6] & r_1[6] /*7972*/;
  assign _252_ = _250_ | _251_ /*7971*/;
  assign _253_ = inv_2[7] ^ r_1[7] /*7969*/;
  assign sum_2[7] = _253_ ^ _252_ /*7968*/;
  assign _254_ = _253_ & _252_ /*7967*/;
  assign _255_ = inv_2[7] & r_1[7] /*7966*/;
  assign _256_ = _254_ | _255_ /*7965*/;
  assign _257_ = inv_2[8] ^ r_1[8] /*7963*/;
  assign sum_2[8] = _257_ ^ _256_ /*7962*/;
  assign _258_ = _257_ & _256_ /*7961*/;
  assign _259_ = inv_2[8] & r_1[8] /*7960*/;
  assign _260_ = _258_ | _259_ /*7959*/;
  assign _261_ = inv_2[9] ^ r_1[9] /*7957*/;
  assign sum_2[9] = _261_ ^ _260_ /*7956*/;
  assign _262_ = _261_ & _260_ /*7955*/;
  assign _263_ = inv_2[9] & r_1[9] /*7954*/;
  assign _264_ = _262_ | _263_ /*7953*/;
  assign _265_ = inv_2[10] ^ r_1[10] /*7951*/;
  assign sum_2[10] = _265_ ^ _264_ /*7950*/;
  assign _266_ = _265_ & _264_ /*7949*/;
  assign _267_ = inv_2[10] & r_1[10] /*7948*/;
  assign _268_ = _266_ | _267_ /*7947*/;
  assign _269_ = inv_2[11] ^ r_1[11] /*7945*/;
  assign sum_2[11] = _269_ ^ _268_ /*7944*/;
  assign _270_ = _269_ & _268_ /*7943*/;
  assign _271_ = inv_2[11] & r_1[11] /*7942*/;
  assign _272_ = _270_ | _271_ /*7941*/;
  assign _273_ = inv_2[12] ^ r_1[12] /*7939*/;
  assign sum_2[12] = _273_ ^ _272_ /*7938*/;
  assign _274_ = _273_ & _272_ /*7937*/;
  assign _275_ = inv_2[12] & r_1[12] /*7936*/;
  assign _276_ = _274_ | _275_ /*7935*/;
  assign _277_ = inv_2[13] ^ r_1[13] /*7933*/;
  assign sum_2[13] = _277_ ^ _276_ /*7932*/;
  assign _278_ = _277_ & _276_ /*7931*/;
  assign _279_ = inv_2[13] & r_1[13] /*7930*/;
  assign _280_ = _278_ | _279_ /*7929*/;
  assign _281_ = inv_2[14] ^ r_1[14] /*7927*/;
  assign sum_2[14] = _281_ ^ _280_ /*7926*/;
  assign _282_ = _281_ & _280_ /*7925*/;
  assign _283_ = inv_2[14] & r_1[14] /*7924*/;
  assign _284_ = _282_ | _283_ /*7923*/;
  assign _285_ = inv_2[15] ^ r_1[15] /*7921*/;
  assign sum_2[15] = _285_ ^ _284_ /*7920*/;
  assign _286_ = _285_ & _284_ /*7919*/;
  assign _287_ = inv_2[15] & r_1[15] /*7918*/;
  assign _288_ = _286_ | _287_ /*7917*/;
  assign _289_ = inv_2[16] ^ r_1[16] /*7915*/;
  assign sum_2[16] = _289_ ^ _288_ /*7914*/;
  assign _290_ = _289_ & _288_ /*7913*/;
  assign _291_ = inv_2[16] & r_1[16] /*7912*/;
  assign _292_ = _290_ | _291_ /*7911*/;
  assign _293_ = inv_2[17] ^ r_1[17] /*7909*/;
  assign sum_2[17] = _293_ ^ _292_ /*7908*/;
  assign _294_ = _293_ & _292_ /*7907*/;
  assign _295_ = inv_2[17] & r_1[17] /*7906*/;
  assign _296_ = _294_ | _295_ /*7905*/;
  assign _297_ = inv_2[18] ^ r_1[18] /*7903*/;
  assign sum_2[18] = _297_ ^ _296_ /*7902*/;
  assign _298_ = _297_ & _296_ /*7901*/;
  assign _299_ = inv_2[18] & r_1[18] /*7900*/;
  assign _300_ = _298_ | _299_ /*7899*/;
  assign _301_ = inv_2[19] ^ r_1[19] /*7897*/;
  assign sum_2[19] = _301_ ^ _300_ /*7896*/;
  assign _302_ = _301_ & _300_ /*7895*/;
  assign _303_ = inv_2[19] & r_1[19] /*7894*/;
  assign _304_ = _302_ | _303_ /*7893*/;
  assign _305_ = inv_2[20] ^ r_1[20] /*7891*/;
  assign sum_2[20] = _305_ ^ _304_ /*7890*/;
  assign _306_ = _305_ & _304_ /*7889*/;
  assign _307_ = inv_2[20] & r_1[20] /*7888*/;
  assign _308_ = _306_ | _307_ /*7887*/;
  assign _309_ = inv_2[21] ^ r_1[21] /*7885*/;
  assign sum_2[21] = _309_ ^ _308_ /*7884*/;
  assign _310_ = _309_ & _308_ /*7883*/;
  assign _311_ = inv_2[21] & r_1[21] /*7882*/;
  assign _312_ = _310_ | _311_ /*7881*/;
  assign _313_ = inv_2[22] ^ r_1[22] /*7879*/;
  assign sum_2[22] = _313_ ^ _312_ /*7878*/;
  assign _314_ = _313_ & _312_ /*7877*/;
  assign _315_ = inv_2[22] & r_1[22] /*7876*/;
  assign _316_ = _314_ | _315_ /*7875*/;
  assign _317_ = inv_2[23] ^ r_1[23] /*7873*/;
  assign sum_2[23] = _317_ ^ _316_ /*7872*/;
  assign _318_ = _317_ & _316_ /*7871*/;
  assign _319_ = inv_2[23] & r_1[23] /*7870*/;
  assign _320_ = _318_ | _319_ /*7869*/;
  assign _321_ = inv_2[24] ^ r_1[24] /*7867*/;
  assign sum_2[24] = _321_ ^ _320_ /*7866*/;
  assign _322_ = _321_ & _320_ /*7865*/;
  assign _323_ = inv_2[24] & r_1[24] /*7864*/;
  assign _324_ = _322_ | _323_ /*7863*/;
  assign _325_ = inv_2[25] ^ r_1[25] /*7861*/;
  assign sum_2[25] = _325_ ^ _324_ /*7860*/;
  assign _326_ = _325_ & _324_ /*7859*/;
  assign _327_ = inv_2[25] & r_1[25] /*7858*/;
  assign _328_ = _326_ | _327_ /*7857*/;
  assign _329_ = inv_2[26] ^ r_1[26] /*7855*/;
  assign sum_2[26] = _329_ ^ _328_ /*7854*/;
  assign _330_ = _329_ & _328_ /*7853*/;
  assign _331_ = inv_2[26] & r_1[26] /*7852*/;
  assign _332_ = _330_ | _331_ /*7851*/;
  assign _333_ = inv_2[27] ^ r_1[27] /*7849*/;
  assign sum_2[27] = _333_ ^ _332_ /*7848*/;
  assign _334_ = _333_ & _332_ /*7847*/;
  assign _335_ = inv_2[27] & r_1[27] /*7846*/;
  assign _336_ = _334_ | _335_ /*7845*/;
  assign _337_ = inv_2[28] ^ r_1[28] /*7843*/;
  assign sum_2[28] = _337_ ^ _336_ /*7842*/;
  assign _338_ = _337_ & _336_ /*7841*/;
  assign _339_ = inv_2[28] & r_1[28] /*7840*/;
  assign _340_ = _338_ | _339_ /*7839*/;
  assign _341_ = inv_2[29] ^ r_1[29] /*7837*/;
  assign sum_2[29] = _341_ ^ _340_ /*7836*/;
  assign _342_ = _341_ & _340_ /*7835*/;
  assign _343_ = inv_2[29] & r_1[29] /*7834*/;
  assign _344_ = _342_ | _343_ /*7833*/;
  assign _345_ = inv_2[30] ^ r_1[30] /*7831*/;
  assign sum_2[30] = _345_ ^ _344_ /*7830*/;
  assign _346_ = _345_ & _344_ /*7829*/;
  assign _347_ = inv_2[30] & r_1[30] /*7828*/;
  assign _348_ = _346_ | _347_ /*7827*/;
  assign _349_ = inv_2[31] ^ r_1[31] /*7825*/;
  assign sum_2[31] = _349_ ^ _348_ /*7824*/;
  assign _350_ = _349_ & _348_ /*7823*/;
  assign _351_ = inv_2[31] & r_1[31] /*7822*/;
  assign _352_ = _350_ | _351_ /*7821*/;
  assign _353_ = _352_ ^ _348_ /*7820*/;
  assign _354_ = ~_353_ /*7819*/;
  assign _355_ = sum_2[31] & _354_ /*7818*/;
  assign _356_ = _353_ & _352_ /*7817*/;
  assign sum_2[32] = _356_ | _355_ /*7816*/;
  assign q[14] = ~sum_2[32] /*7815*/;
  assign m_2[0] = r_1[0] /*7814*/;
  assign m_2[1] = r_1[1] /*7813*/;
  assign m_2[2] = r_1[2] /*7812*/;
  assign m_2[3] = r_1[3] /*7811*/;
  assign m_2[4] = r_1[4] /*7810*/;
  assign m_2[5] = r_1[5] /*7809*/;
  assign m_2[6] = r_1[6] /*7808*/;
  assign m_2[7] = r_1[7] /*7807*/;
  assign m_2[8] = r_1[8] /*7806*/;
  assign m_2[9] = r_1[9] /*7805*/;
  assign m_2[10] = r_1[10] /*7804*/;
  assign m_2[11] = r_1[11] /*7803*/;
  assign m_2[12] = r_1[12] /*7802*/;
  assign m_2[13] = r_1[13] /*7801*/;
  assign m_2[14] = r_1[14] /*7800*/;
  assign m_2[15] = r_1[15] /*7799*/;
  assign m_2[16] = r_1[16] /*7798*/;
  assign m_2[17] = r_1[17] /*7797*/;
  assign m_2[18] = r_1[18] /*7796*/;
  assign m_2[19] = r_1[19] /*7795*/;
  assign m_2[20] = r_1[20] /*7794*/;
  assign m_2[21] = r_1[21] /*7793*/;
  assign m_2[22] = r_1[22] /*7792*/;
  assign m_2[23] = r_1[23] /*7791*/;
  assign m_2[24] = r_1[24] /*7790*/;
  assign m_2[25] = r_1[25] /*7789*/;
  assign m_2[26] = r_1[26] /*7788*/;
  assign m_2[27] = r_1[27] /*7787*/;
  assign m_2[28] = r_1[28] /*7786*/;
  assign m_2[29] = r_1[29] /*7785*/;
  assign m_2[30] = r_1[30] /*7784*/;
  assign m_2[31] = r_1[31] /*7783*/;
  assign m_2[32] = r_1[31] /*7782*/;
  assign _358_ = ~q[14] /*7781*/;
  assign _359_ = sum_2[0] & q[14] /*7780*/;
  assign _360_ = m_2[0] & _358_ /*7779*/;
  assign r_2[0] = _360_ | _359_ /*7778*/;
  assign _361_ = ~q[14] /*7777*/;
  assign _362_ = sum_2[1] & q[14] /*7776*/;
  assign _363_ = m_2[1] & _361_ /*7775*/;
  assign r_2[1] = _363_ | _362_ /*7774*/;
  assign _364_ = ~q[14] /*7773*/;
  assign _365_ = sum_2[2] & q[14] /*7772*/;
  assign _366_ = m_2[2] & _364_ /*7771*/;
  assign r_2[2] = _366_ | _365_ /*7770*/;
  assign _367_ = ~q[14] /*7769*/;
  assign _368_ = sum_2[3] & q[14] /*7768*/;
  assign _369_ = m_2[3] & _367_ /*7767*/;
  assign r_2[3] = _369_ | _368_ /*7766*/;
  assign _370_ = ~q[14] /*7765*/;
  assign _371_ = sum_2[4] & q[14] /*7764*/;
  assign _372_ = m_2[4] & _370_ /*7763*/;
  assign r_2[4] = _372_ | _371_ /*7762*/;
  assign _373_ = ~q[14] /*7761*/;
  assign _374_ = sum_2[5] & q[14] /*7760*/;
  assign _375_ = m_2[5] & _373_ /*7759*/;
  assign r_2[5] = _375_ | _374_ /*7758*/;
  assign _376_ = ~q[14] /*7757*/;
  assign _377_ = sum_2[6] & q[14] /*7756*/;
  assign _378_ = m_2[6] & _376_ /*7755*/;
  assign r_2[6] = _378_ | _377_ /*7754*/;
  assign _379_ = ~q[14] /*7753*/;
  assign _380_ = sum_2[7] & q[14] /*7752*/;
  assign _381_ = m_2[7] & _379_ /*7751*/;
  assign r_2[7] = _381_ | _380_ /*7750*/;
  assign _382_ = ~q[14] /*7749*/;
  assign _383_ = sum_2[8] & q[14] /*7748*/;
  assign _384_ = m_2[8] & _382_ /*7747*/;
  assign r_2[8] = _384_ | _383_ /*7746*/;
  assign _385_ = ~q[14] /*7745*/;
  assign _386_ = sum_2[9] & q[14] /*7744*/;
  assign _387_ = m_2[9] & _385_ /*7743*/;
  assign r_2[9] = _387_ | _386_ /*7742*/;
  assign _388_ = ~q[14] /*7741*/;
  assign _389_ = sum_2[10] & q[14] /*7740*/;
  assign _390_ = m_2[10] & _388_ /*7739*/;
  assign r_2[10] = _390_ | _389_ /*7738*/;
  assign _391_ = ~q[14] /*7737*/;
  assign _392_ = sum_2[11] & q[14] /*7736*/;
  assign _393_ = m_2[11] & _391_ /*7735*/;
  assign r_2[11] = _393_ | _392_ /*7734*/;
  assign _394_ = ~q[14] /*7733*/;
  assign _395_ = sum_2[12] & q[14] /*7732*/;
  assign _396_ = m_2[12] & _394_ /*7731*/;
  assign r_2[12] = _396_ | _395_ /*7730*/;
  assign _397_ = ~q[14] /*7729*/;
  assign _398_ = sum_2[13] & q[14] /*7728*/;
  assign _399_ = m_2[13] & _397_ /*7727*/;
  assign r_2[13] = _399_ | _398_ /*7726*/;
  assign _400_ = ~q[14] /*7725*/;
  assign _401_ = sum_2[14] & q[14] /*7724*/;
  assign _402_ = m_2[14] & _400_ /*7723*/;
  assign r_2[14] = _402_ | _401_ /*7722*/;
  assign _403_ = ~q[14] /*7721*/;
  assign _404_ = sum_2[15] & q[14] /*7720*/;
  assign _405_ = m_2[15] & _403_ /*7719*/;
  assign r_2[15] = _405_ | _404_ /*7718*/;
  assign _406_ = ~q[14] /*7717*/;
  assign _407_ = sum_2[16] & q[14] /*7716*/;
  assign _408_ = m_2[16] & _406_ /*7715*/;
  assign r_2[16] = _408_ | _407_ /*7714*/;
  assign _409_ = ~q[14] /*7713*/;
  assign _410_ = sum_2[17] & q[14] /*7712*/;
  assign _411_ = m_2[17] & _409_ /*7711*/;
  assign r_2[17] = _411_ | _410_ /*7710*/;
  assign _412_ = ~q[14] /*7709*/;
  assign _413_ = sum_2[18] & q[14] /*7708*/;
  assign _414_ = m_2[18] & _412_ /*7707*/;
  assign r_2[18] = _414_ | _413_ /*7706*/;
  assign _415_ = ~q[14] /*7705*/;
  assign _416_ = sum_2[19] & q[14] /*7704*/;
  assign _417_ = m_2[19] & _415_ /*7703*/;
  assign r_2[19] = _417_ | _416_ /*7702*/;
  assign _418_ = ~q[14] /*7701*/;
  assign _419_ = sum_2[20] & q[14] /*7700*/;
  assign _420_ = m_2[20] & _418_ /*7699*/;
  assign r_2[20] = _420_ | _419_ /*7698*/;
  assign _421_ = ~q[14] /*7697*/;
  assign _422_ = sum_2[21] & q[14] /*7696*/;
  assign _423_ = m_2[21] & _421_ /*7695*/;
  assign r_2[21] = _423_ | _422_ /*7694*/;
  assign _424_ = ~q[14] /*7693*/;
  assign _425_ = sum_2[22] & q[14] /*7692*/;
  assign _426_ = m_2[22] & _424_ /*7691*/;
  assign r_2[22] = _426_ | _425_ /*7690*/;
  assign _427_ = ~q[14] /*7689*/;
  assign _428_ = sum_2[23] & q[14] /*7688*/;
  assign _429_ = m_2[23] & _427_ /*7687*/;
  assign r_2[23] = _429_ | _428_ /*7686*/;
  assign _430_ = ~q[14] /*7685*/;
  assign _431_ = sum_2[24] & q[14] /*7684*/;
  assign _432_ = m_2[24] & _430_ /*7683*/;
  assign r_2[24] = _432_ | _431_ /*7682*/;
  assign _433_ = ~q[14] /*7681*/;
  assign _434_ = sum_2[25] & q[14] /*7680*/;
  assign _435_ = m_2[25] & _433_ /*7679*/;
  assign r_2[25] = _435_ | _434_ /*7678*/;
  assign _436_ = ~q[14] /*7677*/;
  assign _437_ = sum_2[26] & q[14] /*7676*/;
  assign _438_ = m_2[26] & _436_ /*7675*/;
  assign r_2[26] = _438_ | _437_ /*7674*/;
  assign _439_ = ~q[14] /*7673*/;
  assign _440_ = sum_2[27] & q[14] /*7672*/;
  assign _441_ = m_2[27] & _439_ /*7671*/;
  assign r_2[27] = _441_ | _440_ /*7670*/;
  assign _442_ = ~q[14] /*7669*/;
  assign _443_ = sum_2[28] & q[14] /*7668*/;
  assign _444_ = m_2[28] & _442_ /*7667*/;
  assign r_2[28] = _444_ | _443_ /*7666*/;
  assign _445_ = ~q[14] /*7665*/;
  assign _446_ = sum_2[29] & q[14] /*7664*/;
  assign _447_ = m_2[29] & _445_ /*7663*/;
  assign r_2[29] = _447_ | _446_ /*7662*/;
  assign _448_ = ~q[14] /*7661*/;
  assign _449_ = sum_2[30] & q[14] /*7660*/;
  assign _450_ = m_2[30] & _448_ /*7659*/;
  assign r_2[30] = _450_ | _449_ /*7658*/;
  assign _451_ = ~q[14] /*7657*/;
  assign _452_ = sum_2[31] & q[14] /*7656*/;
  assign _453_ = m_2[31] & _451_ /*7655*/;
  assign r_2[31] = _453_ | _452_ /*7654*/;
  assign _454_ = ~q[14] /*7653*/;
  assign _455_ = sum_2[32] & q[14] /*7652*/;
  assign _456_ = m_2[32] & _454_ /*7651*/;
  assign r_2[32] = _456_ | _455_ /*7650*/;
  assign inv_3[0] = oneWire /*7480*/;
  assign inv_3[1] = oneWire /*7474*/;
  assign inv_3[2] = oneWire /*7468*/;
  assign inv_3[3] = oneWire /*7462*/;
  assign inv_3[4] = oneWire /*7456*/;
  assign inv_3[5] = oneWire /*7450*/;
  assign inv_3[6] = oneWire /*7444*/;
  assign inv_3[7] = oneWire /*7438*/;
  assign inv_3[8] = oneWire /*7432*/;
  assign inv_3[9] = oneWire /*7426*/;
  assign inv_3[10] = oneWire /*7420*/;
  assign inv_3[11] = oneWire /*7414*/;
  assign inv_3[12] = oneWire /*7408*/;
  assign inv_3[13] = ~div[0] /*7402*/;
  assign inv_3[14] = ~div[1] /*7396*/;
  assign inv_3[15] = ~div[2] /*7390*/;
  assign inv_3[16] = ~div[3] /*7384*/;
  assign inv_3[17] = ~div[4] /*7378*/;
  assign inv_3[18] = ~div[5] /*7372*/;
  assign inv_3[19] = ~div[6] /*7366*/;
  assign inv_3[20] = ~div[7] /*7360*/;
  assign inv_3[21] = ~div[8] /*7354*/;
  assign inv_3[22] = ~div[9] /*7348*/;
  assign inv_3[23] = ~div[10] /*7342*/;
  assign inv_3[24] = ~div[11] /*7336*/;
  assign inv_3[25] = ~div[12] /*7330*/;
  assign inv_3[26] = ~div[13] /*7324*/;
  assign inv_3[27] = ~div[14] /*7318*/;
  assign inv_3[28] = oneWire /*7312*/;
  assign inv_3[29] = oneWire /*7306*/;
  assign inv_3[30] = oneWire /*7300*/;
  assign inv_3[31] = oneWire /*7294*/;
  assign inv_3[32] = oneWire /*7288*/;
  assign _457_ = inv_3[0] ^ r_2[0] /*7479*/;
  assign sum_3[0] = _457_ ^ oneWire /*7478*/;
  assign _458_ = _457_ & oneWire /*7477*/;
  assign _459_ = inv_3[0] & r_2[0] /*7476*/;
  assign _460_ = _458_ | _459_ /*7475*/;
  assign _461_ = inv_3[1] ^ r_2[1] /*7473*/;
  assign sum_3[1] = _461_ ^ _460_ /*7472*/;
  assign _462_ = _461_ & _460_ /*7471*/;
  assign _463_ = inv_3[1] & r_2[1] /*7470*/;
  assign _464_ = _462_ | _463_ /*7469*/;
  assign _465_ = inv_3[2] ^ r_2[2] /*7467*/;
  assign sum_3[2] = _465_ ^ _464_ /*7466*/;
  assign _466_ = _465_ & _464_ /*7465*/;
  assign _467_ = inv_3[2] & r_2[2] /*7464*/;
  assign _468_ = _466_ | _467_ /*7463*/;
  assign _469_ = inv_3[3] ^ r_2[3] /*7461*/;
  assign sum_3[3] = _469_ ^ _468_ /*7460*/;
  assign _470_ = _469_ & _468_ /*7459*/;
  assign _471_ = inv_3[3] & r_2[3] /*7458*/;
  assign _472_ = _470_ | _471_ /*7457*/;
  assign _473_ = inv_3[4] ^ r_2[4] /*7455*/;
  assign sum_3[4] = _473_ ^ _472_ /*7454*/;
  assign _474_ = _473_ & _472_ /*7453*/;
  assign _475_ = inv_3[4] & r_2[4] /*7452*/;
  assign _476_ = _474_ | _475_ /*7451*/;
  assign _477_ = inv_3[5] ^ r_2[5] /*7449*/;
  assign sum_3[5] = _477_ ^ _476_ /*7448*/;
  assign _478_ = _477_ & _476_ /*7447*/;
  assign _479_ = inv_3[5] & r_2[5] /*7446*/;
  assign _480_ = _478_ | _479_ /*7445*/;
  assign _481_ = inv_3[6] ^ r_2[6] /*7443*/;
  assign sum_3[6] = _481_ ^ _480_ /*7442*/;
  assign _482_ = _481_ & _480_ /*7441*/;
  assign _483_ = inv_3[6] & r_2[6] /*7440*/;
  assign _484_ = _482_ | _483_ /*7439*/;
  assign _485_ = inv_3[7] ^ r_2[7] /*7437*/;
  assign sum_3[7] = _485_ ^ _484_ /*7436*/;
  assign _486_ = _485_ & _484_ /*7435*/;
  assign _487_ = inv_3[7] & r_2[7] /*7434*/;
  assign _488_ = _486_ | _487_ /*7433*/;
  assign _489_ = inv_3[8] ^ r_2[8] /*7431*/;
  assign sum_3[8] = _489_ ^ _488_ /*7430*/;
  assign _490_ = _489_ & _488_ /*7429*/;
  assign _491_ = inv_3[8] & r_2[8] /*7428*/;
  assign _492_ = _490_ | _491_ /*7427*/;
  assign _493_ = inv_3[9] ^ r_2[9] /*7425*/;
  assign sum_3[9] = _493_ ^ _492_ /*7424*/;
  assign _494_ = _493_ & _492_ /*7423*/;
  assign _495_ = inv_3[9] & r_2[9] /*7422*/;
  assign _496_ = _494_ | _495_ /*7421*/;
  assign _497_ = inv_3[10] ^ r_2[10] /*7419*/;
  assign sum_3[10] = _497_ ^ _496_ /*7418*/;
  assign _498_ = _497_ & _496_ /*7417*/;
  assign _499_ = inv_3[10] & r_2[10] /*7416*/;
  assign _500_ = _498_ | _499_ /*7415*/;
  assign _501_ = inv_3[11] ^ r_2[11] /*7413*/;
  assign sum_3[11] = _501_ ^ _500_ /*7412*/;
  assign _502_ = _501_ & _500_ /*7411*/;
  assign _503_ = inv_3[11] & r_2[11] /*7410*/;
  assign _504_ = _502_ | _503_ /*7409*/;
  assign _505_ = inv_3[12] ^ r_2[12] /*7407*/;
  assign sum_3[12] = _505_ ^ _504_ /*7406*/;
  assign _506_ = _505_ & _504_ /*7405*/;
  assign _507_ = inv_3[12] & r_2[12] /*7404*/;
  assign _508_ = _506_ | _507_ /*7403*/;
  assign _509_ = inv_3[13] ^ r_2[13] /*7401*/;
  assign sum_3[13] = _509_ ^ _508_ /*7400*/;
  assign _510_ = _509_ & _508_ /*7399*/;
  assign _511_ = inv_3[13] & r_2[13] /*7398*/;
  assign _512_ = _510_ | _511_ /*7397*/;
  assign _513_ = inv_3[14] ^ r_2[14] /*7395*/;
  assign sum_3[14] = _513_ ^ _512_ /*7394*/;
  assign _514_ = _513_ & _512_ /*7393*/;
  assign _515_ = inv_3[14] & r_2[14] /*7392*/;
  assign _516_ = _514_ | _515_ /*7391*/;
  assign _517_ = inv_3[15] ^ r_2[15] /*7389*/;
  assign sum_3[15] = _517_ ^ _516_ /*7388*/;
  assign _518_ = _517_ & _516_ /*7387*/;
  assign _519_ = inv_3[15] & r_2[15] /*7386*/;
  assign _520_ = _518_ | _519_ /*7385*/;
  assign _521_ = inv_3[16] ^ r_2[16] /*7383*/;
  assign sum_3[16] = _521_ ^ _520_ /*7382*/;
  assign _522_ = _521_ & _520_ /*7381*/;
  assign _523_ = inv_3[16] & r_2[16] /*7380*/;
  assign _524_ = _522_ | _523_ /*7379*/;
  assign _525_ = inv_3[17] ^ r_2[17] /*7377*/;
  assign sum_3[17] = _525_ ^ _524_ /*7376*/;
  assign _526_ = _525_ & _524_ /*7375*/;
  assign _527_ = inv_3[17] & r_2[17] /*7374*/;
  assign _528_ = _526_ | _527_ /*7373*/;
  assign _529_ = inv_3[18] ^ r_2[18] /*7371*/;
  assign sum_3[18] = _529_ ^ _528_ /*7370*/;
  assign _530_ = _529_ & _528_ /*7369*/;
  assign _531_ = inv_3[18] & r_2[18] /*7368*/;
  assign _532_ = _530_ | _531_ /*7367*/;
  assign _533_ = inv_3[19] ^ r_2[19] /*7365*/;
  assign sum_3[19] = _533_ ^ _532_ /*7364*/;
  assign _534_ = _533_ & _532_ /*7363*/;
  assign _535_ = inv_3[19] & r_2[19] /*7362*/;
  assign _536_ = _534_ | _535_ /*7361*/;
  assign _537_ = inv_3[20] ^ r_2[20] /*7359*/;
  assign sum_3[20] = _537_ ^ _536_ /*7358*/;
  assign _538_ = _537_ & _536_ /*7357*/;
  assign _539_ = inv_3[20] & r_2[20] /*7356*/;
  assign _540_ = _538_ | _539_ /*7355*/;
  assign _541_ = inv_3[21] ^ r_2[21] /*7353*/;
  assign sum_3[21] = _541_ ^ _540_ /*7352*/;
  assign _542_ = _541_ & _540_ /*7351*/;
  assign _543_ = inv_3[21] & r_2[21] /*7350*/;
  assign _544_ = _542_ | _543_ /*7349*/;
  assign _545_ = inv_3[22] ^ r_2[22] /*7347*/;
  assign sum_3[22] = _545_ ^ _544_ /*7346*/;
  assign _546_ = _545_ & _544_ /*7345*/;
  assign _547_ = inv_3[22] & r_2[22] /*7344*/;
  assign _548_ = _546_ | _547_ /*7343*/;
  assign _549_ = inv_3[23] ^ r_2[23] /*7341*/;
  assign sum_3[23] = _549_ ^ _548_ /*7340*/;
  assign _550_ = _549_ & _548_ /*7339*/;
  assign _551_ = inv_3[23] & r_2[23] /*7338*/;
  assign _552_ = _550_ | _551_ /*7337*/;
  assign _553_ = inv_3[24] ^ r_2[24] /*7335*/;
  assign sum_3[24] = _553_ ^ _552_ /*7334*/;
  assign _554_ = _553_ & _552_ /*7333*/;
  assign _555_ = inv_3[24] & r_2[24] /*7332*/;
  assign _556_ = _554_ | _555_ /*7331*/;
  assign _557_ = inv_3[25] ^ r_2[25] /*7329*/;
  assign sum_3[25] = _557_ ^ _556_ /*7328*/;
  assign _558_ = _557_ & _556_ /*7327*/;
  assign _559_ = inv_3[25] & r_2[25] /*7326*/;
  assign _560_ = _558_ | _559_ /*7325*/;
  assign _561_ = inv_3[26] ^ r_2[26] /*7323*/;
  assign sum_3[26] = _561_ ^ _560_ /*7322*/;
  assign _562_ = _561_ & _560_ /*7321*/;
  assign _563_ = inv_3[26] & r_2[26] /*7320*/;
  assign _564_ = _562_ | _563_ /*7319*/;
  assign _565_ = inv_3[27] ^ r_2[27] /*7317*/;
  assign sum_3[27] = _565_ ^ _564_ /*7316*/;
  assign _566_ = _565_ & _564_ /*7315*/;
  assign _567_ = inv_3[27] & r_2[27] /*7314*/;
  assign _568_ = _566_ | _567_ /*7313*/;
  assign _569_ = inv_3[28] ^ r_2[28] /*7311*/;
  assign sum_3[28] = _569_ ^ _568_ /*7310*/;
  assign _570_ = _569_ & _568_ /*7309*/;
  assign _571_ = inv_3[28] & r_2[28] /*7308*/;
  assign _572_ = _570_ | _571_ /*7307*/;
  assign _573_ = inv_3[29] ^ r_2[29] /*7305*/;
  assign sum_3[29] = _573_ ^ _572_ /*7304*/;
  assign _574_ = _573_ & _572_ /*7303*/;
  assign _575_ = inv_3[29] & r_2[29] /*7302*/;
  assign _576_ = _574_ | _575_ /*7301*/;
  assign _577_ = inv_3[30] ^ r_2[30] /*7299*/;
  assign sum_3[30] = _577_ ^ _576_ /*7298*/;
  assign _578_ = _577_ & _576_ /*7297*/;
  assign _579_ = inv_3[30] & r_2[30] /*7296*/;
  assign _580_ = _578_ | _579_ /*7295*/;
  assign _581_ = inv_3[31] ^ r_2[31] /*7293*/;
  assign sum_3[31] = _581_ ^ _580_ /*7292*/;
  assign _582_ = _581_ & _580_ /*7291*/;
  assign _583_ = inv_3[31] & r_2[31] /*7290*/;
  assign _584_ = _582_ | _583_ /*7289*/;
  assign _585_ = inv_3[32] ^ r_2[32] /*7287*/;
  assign sum_3[32] = _585_ ^ _584_ /*7286*/;
  assign _586_ = _585_ & _584_ /*7285*/;
  assign _587_ = inv_3[32] & r_2[32] /*7284*/;
  assign _588_ = _586_ | _587_ /*7283*/;
  assign _589_ = _588_ ^ _584_ /*7282*/;
  assign _590_ = ~_589_ /*7281*/;
  assign _591_ = sum_3[32] & _590_ /*7280*/;
  assign _592_ = _589_ & _588_ /*7279*/;
  assign sum_3[33] = _592_ | _591_ /*7278*/;
  assign q[13] = ~sum_3[33] /*7277*/;
  assign m_3[0] = r_2[0] /*7276*/;
  assign m_3[1] = r_2[1] /*7275*/;
  assign m_3[2] = r_2[2] /*7274*/;
  assign m_3[3] = r_2[3] /*7273*/;
  assign m_3[4] = r_2[4] /*7272*/;
  assign m_3[5] = r_2[5] /*7271*/;
  assign m_3[6] = r_2[6] /*7270*/;
  assign m_3[7] = r_2[7] /*7269*/;
  assign m_3[8] = r_2[8] /*7268*/;
  assign m_3[9] = r_2[9] /*7267*/;
  assign m_3[10] = r_2[10] /*7266*/;
  assign m_3[11] = r_2[11] /*7265*/;
  assign m_3[12] = r_2[12] /*7264*/;
  assign m_3[13] = r_2[13] /*7263*/;
  assign m_3[14] = r_2[14] /*7262*/;
  assign m_3[15] = r_2[15] /*7261*/;
  assign m_3[16] = r_2[16] /*7260*/;
  assign m_3[17] = r_2[17] /*7259*/;
  assign m_3[18] = r_2[18] /*7258*/;
  assign m_3[19] = r_2[19] /*7257*/;
  assign m_3[20] = r_2[20] /*7256*/;
  assign m_3[21] = r_2[21] /*7255*/;
  assign m_3[22] = r_2[22] /*7254*/;
  assign m_3[23] = r_2[23] /*7253*/;
  assign m_3[24] = r_2[24] /*7252*/;
  assign m_3[25] = r_2[25] /*7251*/;
  assign m_3[26] = r_2[26] /*7250*/;
  assign m_3[27] = r_2[27] /*7249*/;
  assign m_3[28] = r_2[28] /*7248*/;
  assign m_3[29] = r_2[29] /*7247*/;
  assign m_3[30] = r_2[30] /*7246*/;
  assign m_3[31] = r_2[31] /*7245*/;
  assign m_3[32] = r_2[32] /*7244*/;
  assign m_3[33] = r_2[32] /*7243*/;
  assign _594_ = ~q[13] /*7242*/;
  assign _595_ = sum_3[0] & q[13] /*7241*/;
  assign _596_ = m_3[0] & _594_ /*7240*/;
  assign r_3[0] = _596_ | _595_ /*7239*/;
  assign _597_ = ~q[13] /*7238*/;
  assign _598_ = sum_3[1] & q[13] /*7237*/;
  assign _599_ = m_3[1] & _597_ /*7236*/;
  assign r_3[1] = _599_ | _598_ /*7235*/;
  assign _600_ = ~q[13] /*7234*/;
  assign _601_ = sum_3[2] & q[13] /*7233*/;
  assign _602_ = m_3[2] & _600_ /*7232*/;
  assign r_3[2] = _602_ | _601_ /*7231*/;
  assign _603_ = ~q[13] /*7230*/;
  assign _604_ = sum_3[3] & q[13] /*7229*/;
  assign _605_ = m_3[3] & _603_ /*7228*/;
  assign r_3[3] = _605_ | _604_ /*7227*/;
  assign _606_ = ~q[13] /*7226*/;
  assign _607_ = sum_3[4] & q[13] /*7225*/;
  assign _608_ = m_3[4] & _606_ /*7224*/;
  assign r_3[4] = _608_ | _607_ /*7223*/;
  assign _609_ = ~q[13] /*7222*/;
  assign _610_ = sum_3[5] & q[13] /*7221*/;
  assign _611_ = m_3[5] & _609_ /*7220*/;
  assign r_3[5] = _611_ | _610_ /*7219*/;
  assign _612_ = ~q[13] /*7218*/;
  assign _613_ = sum_3[6] & q[13] /*7217*/;
  assign _614_ = m_3[6] & _612_ /*7216*/;
  assign r_3[6] = _614_ | _613_ /*7215*/;
  assign _615_ = ~q[13] /*7214*/;
  assign _616_ = sum_3[7] & q[13] /*7213*/;
  assign _617_ = m_3[7] & _615_ /*7212*/;
  assign r_3[7] = _617_ | _616_ /*7211*/;
  assign _618_ = ~q[13] /*7210*/;
  assign _619_ = sum_3[8] & q[13] /*7209*/;
  assign _620_ = m_3[8] & _618_ /*7208*/;
  assign r_3[8] = _620_ | _619_ /*7207*/;
  assign _621_ = ~q[13] /*7206*/;
  assign _622_ = sum_3[9] & q[13] /*7205*/;
  assign _623_ = m_3[9] & _621_ /*7204*/;
  assign r_3[9] = _623_ | _622_ /*7203*/;
  assign _624_ = ~q[13] /*7202*/;
  assign _625_ = sum_3[10] & q[13] /*7201*/;
  assign _626_ = m_3[10] & _624_ /*7200*/;
  assign r_3[10] = _626_ | _625_ /*7199*/;
  assign _627_ = ~q[13] /*7198*/;
  assign _628_ = sum_3[11] & q[13] /*7197*/;
  assign _629_ = m_3[11] & _627_ /*7196*/;
  assign r_3[11] = _629_ | _628_ /*7195*/;
  assign _630_ = ~q[13] /*7194*/;
  assign _631_ = sum_3[12] & q[13] /*7193*/;
  assign _632_ = m_3[12] & _630_ /*7192*/;
  assign r_3[12] = _632_ | _631_ /*7191*/;
  assign _633_ = ~q[13] /*7190*/;
  assign _634_ = sum_3[13] & q[13] /*7189*/;
  assign _635_ = m_3[13] & _633_ /*7188*/;
  assign r_3[13] = _635_ | _634_ /*7187*/;
  assign _636_ = ~q[13] /*7186*/;
  assign _637_ = sum_3[14] & q[13] /*7185*/;
  assign _638_ = m_3[14] & _636_ /*7184*/;
  assign r_3[14] = _638_ | _637_ /*7183*/;
  assign _639_ = ~q[13] /*7182*/;
  assign _640_ = sum_3[15] & q[13] /*7181*/;
  assign _641_ = m_3[15] & _639_ /*7180*/;
  assign r_3[15] = _641_ | _640_ /*7179*/;
  assign _642_ = ~q[13] /*7178*/;
  assign _643_ = sum_3[16] & q[13] /*7177*/;
  assign _644_ = m_3[16] & _642_ /*7176*/;
  assign r_3[16] = _644_ | _643_ /*7175*/;
  assign _645_ = ~q[13] /*7174*/;
  assign _646_ = sum_3[17] & q[13] /*7173*/;
  assign _647_ = m_3[17] & _645_ /*7172*/;
  assign r_3[17] = _647_ | _646_ /*7171*/;
  assign _648_ = ~q[13] /*7170*/;
  assign _649_ = sum_3[18] & q[13] /*7169*/;
  assign _650_ = m_3[18] & _648_ /*7168*/;
  assign r_3[18] = _650_ | _649_ /*7167*/;
  assign _651_ = ~q[13] /*7166*/;
  assign _652_ = sum_3[19] & q[13] /*7165*/;
  assign _653_ = m_3[19] & _651_ /*7164*/;
  assign r_3[19] = _653_ | _652_ /*7163*/;
  assign _654_ = ~q[13] /*7162*/;
  assign _655_ = sum_3[20] & q[13] /*7161*/;
  assign _656_ = m_3[20] & _654_ /*7160*/;
  assign r_3[20] = _656_ | _655_ /*7159*/;
  assign _657_ = ~q[13] /*7158*/;
  assign _658_ = sum_3[21] & q[13] /*7157*/;
  assign _659_ = m_3[21] & _657_ /*7156*/;
  assign r_3[21] = _659_ | _658_ /*7155*/;
  assign _660_ = ~q[13] /*7154*/;
  assign _661_ = sum_3[22] & q[13] /*7153*/;
  assign _662_ = m_3[22] & _660_ /*7152*/;
  assign r_3[22] = _662_ | _661_ /*7151*/;
  assign _663_ = ~q[13] /*7150*/;
  assign _664_ = sum_3[23] & q[13] /*7149*/;
  assign _665_ = m_3[23] & _663_ /*7148*/;
  assign r_3[23] = _665_ | _664_ /*7147*/;
  assign _666_ = ~q[13] /*7146*/;
  assign _667_ = sum_3[24] & q[13] /*7145*/;
  assign _668_ = m_3[24] & _666_ /*7144*/;
  assign r_3[24] = _668_ | _667_ /*7143*/;
  assign _669_ = ~q[13] /*7142*/;
  assign _670_ = sum_3[25] & q[13] /*7141*/;
  assign _671_ = m_3[25] & _669_ /*7140*/;
  assign r_3[25] = _671_ | _670_ /*7139*/;
  assign _672_ = ~q[13] /*7138*/;
  assign _673_ = sum_3[26] & q[13] /*7137*/;
  assign _674_ = m_3[26] & _672_ /*7136*/;
  assign r_3[26] = _674_ | _673_ /*7135*/;
  assign _675_ = ~q[13] /*7134*/;
  assign _676_ = sum_3[27] & q[13] /*7133*/;
  assign _677_ = m_3[27] & _675_ /*7132*/;
  assign r_3[27] = _677_ | _676_ /*7131*/;
  assign _678_ = ~q[13] /*7130*/;
  assign _679_ = sum_3[28] & q[13] /*7129*/;
  assign _680_ = m_3[28] & _678_ /*7128*/;
  assign r_3[28] = _680_ | _679_ /*7127*/;
  assign _681_ = ~q[13] /*7126*/;
  assign _682_ = sum_3[29] & q[13] /*7125*/;
  assign _683_ = m_3[29] & _681_ /*7124*/;
  assign r_3[29] = _683_ | _682_ /*7123*/;
  assign _684_ = ~q[13] /*7122*/;
  assign _685_ = sum_3[30] & q[13] /*7121*/;
  assign _686_ = m_3[30] & _684_ /*7120*/;
  assign r_3[30] = _686_ | _685_ /*7119*/;
  assign _687_ = ~q[13] /*7118*/;
  assign _688_ = sum_3[31] & q[13] /*7117*/;
  assign _689_ = m_3[31] & _687_ /*7116*/;
  assign r_3[31] = _689_ | _688_ /*7115*/;
  assign _690_ = ~q[13] /*7114*/;
  assign _691_ = sum_3[32] & q[13] /*7113*/;
  assign _692_ = m_3[32] & _690_ /*7112*/;
  assign r_3[32] = _692_ | _691_ /*7111*/;
  assign _693_ = ~q[13] /*7110*/;
  assign _694_ = sum_3[33] & q[13] /*7109*/;
  assign _695_ = m_3[33] & _693_ /*7108*/;
  assign r_3[33] = _695_ | _694_ /*7107*/;
  assign inv_4[0] = oneWire /*6948*/;
  assign inv_4[1] = oneWire /*6942*/;
  assign inv_4[2] = oneWire /*6936*/;
  assign inv_4[3] = oneWire /*6930*/;
  assign inv_4[4] = oneWire /*6924*/;
  assign inv_4[5] = oneWire /*6918*/;
  assign inv_4[6] = oneWire /*6912*/;
  assign inv_4[7] = oneWire /*6906*/;
  assign inv_4[8] = oneWire /*6900*/;
  assign inv_4[9] = oneWire /*6894*/;
  assign inv_4[10] = oneWire /*6888*/;
  assign inv_4[11] = oneWire /*6882*/;
  assign inv_4[12] = ~div[0] /*6876*/;
  assign inv_4[13] = ~div[1] /*6870*/;
  assign inv_4[14] = ~div[2] /*6864*/;
  assign inv_4[15] = ~div[3] /*6858*/;
  assign inv_4[16] = ~div[4] /*6852*/;
  assign inv_4[17] = ~div[5] /*6846*/;
  assign inv_4[18] = ~div[6] /*6840*/;
  assign inv_4[19] = ~div[7] /*6834*/;
  assign inv_4[20] = ~div[8] /*6828*/;
  assign inv_4[21] = ~div[9] /*6822*/;
  assign inv_4[22] = ~div[10] /*6816*/;
  assign inv_4[23] = ~div[11] /*6810*/;
  assign inv_4[24] = ~div[12] /*6804*/;
  assign inv_4[25] = ~div[13] /*6798*/;
  assign inv_4[26] = ~div[14] /*6792*/;
  assign inv_4[27] = oneWire /*6786*/;
  assign inv_4[28] = oneWire /*6780*/;
  assign inv_4[29] = oneWire /*6774*/;
  assign inv_4[30] = oneWire /*6768*/;
  assign inv_4[31] = oneWire /*6762*/;
  assign inv_4[32] = oneWire /*6756*/;
  assign inv_4[33] = oneWire /*6750*/;
  assign _696_ = inv_4[0] ^ r_3[0] /*6947*/;
  assign sum_4[0] = _696_ ^ oneWire /*6946*/;
  assign _697_ = _696_ & oneWire /*6945*/;
  assign _698_ = inv_4[0] & r_3[0] /*6944*/;
  assign _699_ = _697_ | _698_ /*6943*/;
  assign _700_ = inv_4[1] ^ r_3[1] /*6941*/;
  assign sum_4[1] = _700_ ^ _699_ /*6940*/;
  assign _701_ = _700_ & _699_ /*6939*/;
  assign _702_ = inv_4[1] & r_3[1] /*6938*/;
  assign _703_ = _701_ | _702_ /*6937*/;
  assign _704_ = inv_4[2] ^ r_3[2] /*6935*/;
  assign sum_4[2] = _704_ ^ _703_ /*6934*/;
  assign _705_ = _704_ & _703_ /*6933*/;
  assign _706_ = inv_4[2] & r_3[2] /*6932*/;
  assign _707_ = _705_ | _706_ /*6931*/;
  assign _708_ = inv_4[3] ^ r_3[3] /*6929*/;
  assign sum_4[3] = _708_ ^ _707_ /*6928*/;
  assign _709_ = _708_ & _707_ /*6927*/;
  assign _710_ = inv_4[3] & r_3[3] /*6926*/;
  assign _711_ = _709_ | _710_ /*6925*/;
  assign _712_ = inv_4[4] ^ r_3[4] /*6923*/;
  assign sum_4[4] = _712_ ^ _711_ /*6922*/;
  assign _713_ = _712_ & _711_ /*6921*/;
  assign _714_ = inv_4[4] & r_3[4] /*6920*/;
  assign _715_ = _713_ | _714_ /*6919*/;
  assign _716_ = inv_4[5] ^ r_3[5] /*6917*/;
  assign sum_4[5] = _716_ ^ _715_ /*6916*/;
  assign _717_ = _716_ & _715_ /*6915*/;
  assign _718_ = inv_4[5] & r_3[5] /*6914*/;
  assign _719_ = _717_ | _718_ /*6913*/;
  assign _720_ = inv_4[6] ^ r_3[6] /*6911*/;
  assign sum_4[6] = _720_ ^ _719_ /*6910*/;
  assign _721_ = _720_ & _719_ /*6909*/;
  assign _722_ = inv_4[6] & r_3[6] /*6908*/;
  assign _723_ = _721_ | _722_ /*6907*/;
  assign _724_ = inv_4[7] ^ r_3[7] /*6905*/;
  assign sum_4[7] = _724_ ^ _723_ /*6904*/;
  assign _725_ = _724_ & _723_ /*6903*/;
  assign _726_ = inv_4[7] & r_3[7] /*6902*/;
  assign _727_ = _725_ | _726_ /*6901*/;
  assign _728_ = inv_4[8] ^ r_3[8] /*6899*/;
  assign sum_4[8] = _728_ ^ _727_ /*6898*/;
  assign _729_ = _728_ & _727_ /*6897*/;
  assign _730_ = inv_4[8] & r_3[8] /*6896*/;
  assign _731_ = _729_ | _730_ /*6895*/;
  assign _732_ = inv_4[9] ^ r_3[9] /*6893*/;
  assign sum_4[9] = _732_ ^ _731_ /*6892*/;
  assign _733_ = _732_ & _731_ /*6891*/;
  assign _734_ = inv_4[9] & r_3[9] /*6890*/;
  assign _735_ = _733_ | _734_ /*6889*/;
  assign _736_ = inv_4[10] ^ r_3[10] /*6887*/;
  assign sum_4[10] = _736_ ^ _735_ /*6886*/;
  assign _737_ = _736_ & _735_ /*6885*/;
  assign _738_ = inv_4[10] & r_3[10] /*6884*/;
  assign _739_ = _737_ | _738_ /*6883*/;
  assign _740_ = inv_4[11] ^ r_3[11] /*6881*/;
  assign sum_4[11] = _740_ ^ _739_ /*6880*/;
  assign _741_ = _740_ & _739_ /*6879*/;
  assign _742_ = inv_4[11] & r_3[11] /*6878*/;
  assign _743_ = _741_ | _742_ /*6877*/;
  assign _744_ = inv_4[12] ^ r_3[12] /*6875*/;
  assign sum_4[12] = _744_ ^ _743_ /*6874*/;
  assign _745_ = _744_ & _743_ /*6873*/;
  assign _746_ = inv_4[12] & r_3[12] /*6872*/;
  assign _747_ = _745_ | _746_ /*6871*/;
  assign _748_ = inv_4[13] ^ r_3[13] /*6869*/;
  assign sum_4[13] = _748_ ^ _747_ /*6868*/;
  assign _749_ = _748_ & _747_ /*6867*/;
  assign _750_ = inv_4[13] & r_3[13] /*6866*/;
  assign _751_ = _749_ | _750_ /*6865*/;
  assign _752_ = inv_4[14] ^ r_3[14] /*6863*/;
  assign sum_4[14] = _752_ ^ _751_ /*6862*/;
  assign _753_ = _752_ & _751_ /*6861*/;
  assign _754_ = inv_4[14] & r_3[14] /*6860*/;
  assign _755_ = _753_ | _754_ /*6859*/;
  assign _756_ = inv_4[15] ^ r_3[15] /*6857*/;
  assign sum_4[15] = _756_ ^ _755_ /*6856*/;
  assign _757_ = _756_ & _755_ /*6855*/;
  assign _758_ = inv_4[15] & r_3[15] /*6854*/;
  assign _759_ = _757_ | _758_ /*6853*/;
  assign _760_ = inv_4[16] ^ r_3[16] /*6851*/;
  assign sum_4[16] = _760_ ^ _759_ /*6850*/;
  assign _761_ = _760_ & _759_ /*6849*/;
  assign _762_ = inv_4[16] & r_3[16] /*6848*/;
  assign _763_ = _761_ | _762_ /*6847*/;
  assign _764_ = inv_4[17] ^ r_3[17] /*6845*/;
  assign sum_4[17] = _764_ ^ _763_ /*6844*/;
  assign _765_ = _764_ & _763_ /*6843*/;
  assign _766_ = inv_4[17] & r_3[17] /*6842*/;
  assign _767_ = _765_ | _766_ /*6841*/;
  assign _768_ = inv_4[18] ^ r_3[18] /*6839*/;
  assign sum_4[18] = _768_ ^ _767_ /*6838*/;
  assign _769_ = _768_ & _767_ /*6837*/;
  assign _770_ = inv_4[18] & r_3[18] /*6836*/;
  assign _771_ = _769_ | _770_ /*6835*/;
  assign _772_ = inv_4[19] ^ r_3[19] /*6833*/;
  assign sum_4[19] = _772_ ^ _771_ /*6832*/;
  assign _773_ = _772_ & _771_ /*6831*/;
  assign _774_ = inv_4[19] & r_3[19] /*6830*/;
  assign _775_ = _773_ | _774_ /*6829*/;
  assign _776_ = inv_4[20] ^ r_3[20] /*6827*/;
  assign sum_4[20] = _776_ ^ _775_ /*6826*/;
  assign _777_ = _776_ & _775_ /*6825*/;
  assign _778_ = inv_4[20] & r_3[20] /*6824*/;
  assign _779_ = _777_ | _778_ /*6823*/;
  assign _780_ = inv_4[21] ^ r_3[21] /*6821*/;
  assign sum_4[21] = _780_ ^ _779_ /*6820*/;
  assign _781_ = _780_ & _779_ /*6819*/;
  assign _782_ = inv_4[21] & r_3[21] /*6818*/;
  assign _783_ = _781_ | _782_ /*6817*/;
  assign _784_ = inv_4[22] ^ r_3[22] /*6815*/;
  assign sum_4[22] = _784_ ^ _783_ /*6814*/;
  assign _785_ = _784_ & _783_ /*6813*/;
  assign _786_ = inv_4[22] & r_3[22] /*6812*/;
  assign _787_ = _785_ | _786_ /*6811*/;
  assign _788_ = inv_4[23] ^ r_3[23] /*6809*/;
  assign sum_4[23] = _788_ ^ _787_ /*6808*/;
  assign _789_ = _788_ & _787_ /*6807*/;
  assign _790_ = inv_4[23] & r_3[23] /*6806*/;
  assign _791_ = _789_ | _790_ /*6805*/;
  assign _792_ = inv_4[24] ^ r_3[24] /*6803*/;
  assign sum_4[24] = _792_ ^ _791_ /*6802*/;
  assign _793_ = _792_ & _791_ /*6801*/;
  assign _794_ = inv_4[24] & r_3[24] /*6800*/;
  assign _795_ = _793_ | _794_ /*6799*/;
  assign _796_ = inv_4[25] ^ r_3[25] /*6797*/;
  assign sum_4[25] = _796_ ^ _795_ /*6796*/;
  assign _797_ = _796_ & _795_ /*6795*/;
  assign _798_ = inv_4[25] & r_3[25] /*6794*/;
  assign _799_ = _797_ | _798_ /*6793*/;
  assign _800_ = inv_4[26] ^ r_3[26] /*6791*/;
  assign sum_4[26] = _800_ ^ _799_ /*6790*/;
  assign _801_ = _800_ & _799_ /*6789*/;
  assign _802_ = inv_4[26] & r_3[26] /*6788*/;
  assign _803_ = _801_ | _802_ /*6787*/;
  assign _804_ = inv_4[27] ^ r_3[27] /*6785*/;
  assign sum_4[27] = _804_ ^ _803_ /*6784*/;
  assign _805_ = _804_ & _803_ /*6783*/;
  assign _806_ = inv_4[27] & r_3[27] /*6782*/;
  assign _807_ = _805_ | _806_ /*6781*/;
  assign _808_ = inv_4[28] ^ r_3[28] /*6779*/;
  assign sum_4[28] = _808_ ^ _807_ /*6778*/;
  assign _809_ = _808_ & _807_ /*6777*/;
  assign _810_ = inv_4[28] & r_3[28] /*6776*/;
  assign _811_ = _809_ | _810_ /*6775*/;
  assign _812_ = inv_4[29] ^ r_3[29] /*6773*/;
  assign sum_4[29] = _812_ ^ _811_ /*6772*/;
  assign _813_ = _812_ & _811_ /*6771*/;
  assign _814_ = inv_4[29] & r_3[29] /*6770*/;
  assign _815_ = _813_ | _814_ /*6769*/;
  assign _816_ = inv_4[30] ^ r_3[30] /*6767*/;
  assign sum_4[30] = _816_ ^ _815_ /*6766*/;
  assign _817_ = _816_ & _815_ /*6765*/;
  assign _818_ = inv_4[30] & r_3[30] /*6764*/;
  assign _819_ = _817_ | _818_ /*6763*/;
  assign _820_ = inv_4[31] ^ r_3[31] /*6761*/;
  assign sum_4[31] = _820_ ^ _819_ /*6760*/;
  assign _821_ = _820_ & _819_ /*6759*/;
  assign _822_ = inv_4[31] & r_3[31] /*6758*/;
  assign _823_ = _821_ | _822_ /*6757*/;
  assign _824_ = inv_4[32] ^ r_3[32] /*6755*/;
  assign sum_4[32] = _824_ ^ _823_ /*6754*/;
  assign _825_ = _824_ & _823_ /*6753*/;
  assign _826_ = inv_4[32] & r_3[32] /*6752*/;
  assign _827_ = _825_ | _826_ /*6751*/;
  assign _828_ = inv_4[33] ^ r_3[33] /*6749*/;
  assign sum_4[33] = _828_ ^ _827_ /*6748*/;
  assign _829_ = _828_ & _827_ /*6747*/;
  assign _830_ = inv_4[33] & r_3[33] /*6746*/;
  assign _831_ = _829_ | _830_ /*6745*/;
  assign _832_ = _831_ ^ _827_ /*6744*/;
  assign _833_ = ~_832_ /*6743*/;
  assign _834_ = sum_4[33] & _833_ /*6742*/;
  assign _835_ = _832_ & _831_ /*6741*/;
  assign sum_4[34] = _835_ | _834_ /*6740*/;
  assign q[12] = ~sum_4[34] /*6739*/;
  assign m_4[0] = r_3[0] /*6738*/;
  assign m_4[1] = r_3[1] /*6737*/;
  assign m_4[2] = r_3[2] /*6736*/;
  assign m_4[3] = r_3[3] /*6735*/;
  assign m_4[4] = r_3[4] /*6734*/;
  assign m_4[5] = r_3[5] /*6733*/;
  assign m_4[6] = r_3[6] /*6732*/;
  assign m_4[7] = r_3[7] /*6731*/;
  assign m_4[8] = r_3[8] /*6730*/;
  assign m_4[9] = r_3[9] /*6729*/;
  assign m_4[10] = r_3[10] /*6728*/;
  assign m_4[11] = r_3[11] /*6727*/;
  assign m_4[12] = r_3[12] /*6726*/;
  assign m_4[13] = r_3[13] /*6725*/;
  assign m_4[14] = r_3[14] /*6724*/;
  assign m_4[15] = r_3[15] /*6723*/;
  assign m_4[16] = r_3[16] /*6722*/;
  assign m_4[17] = r_3[17] /*6721*/;
  assign m_4[18] = r_3[18] /*6720*/;
  assign m_4[19] = r_3[19] /*6719*/;
  assign m_4[20] = r_3[20] /*6718*/;
  assign m_4[21] = r_3[21] /*6717*/;
  assign m_4[22] = r_3[22] /*6716*/;
  assign m_4[23] = r_3[23] /*6715*/;
  assign m_4[24] = r_3[24] /*6714*/;
  assign m_4[25] = r_3[25] /*6713*/;
  assign m_4[26] = r_3[26] /*6712*/;
  assign m_4[27] = r_3[27] /*6711*/;
  assign m_4[28] = r_3[28] /*6710*/;
  assign m_4[29] = r_3[29] /*6709*/;
  assign m_4[30] = r_3[30] /*6708*/;
  assign m_4[31] = r_3[31] /*6707*/;
  assign m_4[32] = r_3[32] /*6706*/;
  assign m_4[33] = r_3[33] /*6705*/;
  assign m_4[34] = r_3[33] /*6704*/;
  assign _837_ = ~q[12] /*6703*/;
  assign _838_ = sum_4[0] & q[12] /*6702*/;
  assign _839_ = m_4[0] & _837_ /*6701*/;
  assign r_4[0] = _839_ | _838_ /*6700*/;
  assign _840_ = ~q[12] /*6699*/;
  assign _841_ = sum_4[1] & q[12] /*6698*/;
  assign _842_ = m_4[1] & _840_ /*6697*/;
  assign r_4[1] = _842_ | _841_ /*6696*/;
  assign _843_ = ~q[12] /*6695*/;
  assign _844_ = sum_4[2] & q[12] /*6694*/;
  assign _845_ = m_4[2] & _843_ /*6693*/;
  assign r_4[2] = _845_ | _844_ /*6692*/;
  assign _846_ = ~q[12] /*6691*/;
  assign _847_ = sum_4[3] & q[12] /*6690*/;
  assign _848_ = m_4[3] & _846_ /*6689*/;
  assign r_4[3] = _848_ | _847_ /*6688*/;
  assign _849_ = ~q[12] /*6687*/;
  assign _850_ = sum_4[4] & q[12] /*6686*/;
  assign _851_ = m_4[4] & _849_ /*6685*/;
  assign r_4[4] = _851_ | _850_ /*6684*/;
  assign _852_ = ~q[12] /*6683*/;
  assign _853_ = sum_4[5] & q[12] /*6682*/;
  assign _854_ = m_4[5] & _852_ /*6681*/;
  assign r_4[5] = _854_ | _853_ /*6680*/;
  assign _855_ = ~q[12] /*6679*/;
  assign _856_ = sum_4[6] & q[12] /*6678*/;
  assign _857_ = m_4[6] & _855_ /*6677*/;
  assign r_4[6] = _857_ | _856_ /*6676*/;
  assign _858_ = ~q[12] /*6675*/;
  assign _859_ = sum_4[7] & q[12] /*6674*/;
  assign _860_ = m_4[7] & _858_ /*6673*/;
  assign r_4[7] = _860_ | _859_ /*6672*/;
  assign _861_ = ~q[12] /*6671*/;
  assign _862_ = sum_4[8] & q[12] /*6670*/;
  assign _863_ = m_4[8] & _861_ /*6669*/;
  assign r_4[8] = _863_ | _862_ /*6668*/;
  assign _864_ = ~q[12] /*6667*/;
  assign _865_ = sum_4[9] & q[12] /*6666*/;
  assign _866_ = m_4[9] & _864_ /*6665*/;
  assign r_4[9] = _866_ | _865_ /*6664*/;
  assign _867_ = ~q[12] /*6663*/;
  assign _868_ = sum_4[10] & q[12] /*6662*/;
  assign _869_ = m_4[10] & _867_ /*6661*/;
  assign r_4[10] = _869_ | _868_ /*6660*/;
  assign _870_ = ~q[12] /*6659*/;
  assign _871_ = sum_4[11] & q[12] /*6658*/;
  assign _872_ = m_4[11] & _870_ /*6657*/;
  assign r_4[11] = _872_ | _871_ /*6656*/;
  assign _873_ = ~q[12] /*6655*/;
  assign _874_ = sum_4[12] & q[12] /*6654*/;
  assign _875_ = m_4[12] & _873_ /*6653*/;
  assign r_4[12] = _875_ | _874_ /*6652*/;
  assign _876_ = ~q[12] /*6651*/;
  assign _877_ = sum_4[13] & q[12] /*6650*/;
  assign _878_ = m_4[13] & _876_ /*6649*/;
  assign r_4[13] = _878_ | _877_ /*6648*/;
  assign _879_ = ~q[12] /*6647*/;
  assign _880_ = sum_4[14] & q[12] /*6646*/;
  assign _881_ = m_4[14] & _879_ /*6645*/;
  assign r_4[14] = _881_ | _880_ /*6644*/;
  assign _882_ = ~q[12] /*6643*/;
  assign _883_ = sum_4[15] & q[12] /*6642*/;
  assign _884_ = m_4[15] & _882_ /*6641*/;
  assign r_4[15] = _884_ | _883_ /*6640*/;
  assign _885_ = ~q[12] /*6639*/;
  assign _886_ = sum_4[16] & q[12] /*6638*/;
  assign _887_ = m_4[16] & _885_ /*6637*/;
  assign r_4[16] = _887_ | _886_ /*6636*/;
  assign _888_ = ~q[12] /*6635*/;
  assign _889_ = sum_4[17] & q[12] /*6634*/;
  assign _890_ = m_4[17] & _888_ /*6633*/;
  assign r_4[17] = _890_ | _889_ /*6632*/;
  assign _891_ = ~q[12] /*6631*/;
  assign _892_ = sum_4[18] & q[12] /*6630*/;
  assign _893_ = m_4[18] & _891_ /*6629*/;
  assign r_4[18] = _893_ | _892_ /*6628*/;
  assign _894_ = ~q[12] /*6627*/;
  assign _895_ = sum_4[19] & q[12] /*6626*/;
  assign _896_ = m_4[19] & _894_ /*6625*/;
  assign r_4[19] = _896_ | _895_ /*6624*/;
  assign _897_ = ~q[12] /*6623*/;
  assign _898_ = sum_4[20] & q[12] /*6622*/;
  assign _899_ = m_4[20] & _897_ /*6621*/;
  assign r_4[20] = _899_ | _898_ /*6620*/;
  assign _900_ = ~q[12] /*6619*/;
  assign _901_ = sum_4[21] & q[12] /*6618*/;
  assign _902_ = m_4[21] & _900_ /*6617*/;
  assign r_4[21] = _902_ | _901_ /*6616*/;
  assign _903_ = ~q[12] /*6615*/;
  assign _904_ = sum_4[22] & q[12] /*6614*/;
  assign _905_ = m_4[22] & _903_ /*6613*/;
  assign r_4[22] = _905_ | _904_ /*6612*/;
  assign _906_ = ~q[12] /*6611*/;
  assign _907_ = sum_4[23] & q[12] /*6610*/;
  assign _908_ = m_4[23] & _906_ /*6609*/;
  assign r_4[23] = _908_ | _907_ /*6608*/;
  assign _909_ = ~q[12] /*6607*/;
  assign _910_ = sum_4[24] & q[12] /*6606*/;
  assign _911_ = m_4[24] & _909_ /*6605*/;
  assign r_4[24] = _911_ | _910_ /*6604*/;
  assign _912_ = ~q[12] /*6603*/;
  assign _913_ = sum_4[25] & q[12] /*6602*/;
  assign _914_ = m_4[25] & _912_ /*6601*/;
  assign r_4[25] = _914_ | _913_ /*6600*/;
  assign _915_ = ~q[12] /*6599*/;
  assign _916_ = sum_4[26] & q[12] /*6598*/;
  assign _917_ = m_4[26] & _915_ /*6597*/;
  assign r_4[26] = _917_ | _916_ /*6596*/;
  assign _918_ = ~q[12] /*6595*/;
  assign _919_ = sum_4[27] & q[12] /*6594*/;
  assign _920_ = m_4[27] & _918_ /*6593*/;
  assign r_4[27] = _920_ | _919_ /*6592*/;
  assign _921_ = ~q[12] /*6591*/;
  assign _922_ = sum_4[28] & q[12] /*6590*/;
  assign _923_ = m_4[28] & _921_ /*6589*/;
  assign r_4[28] = _923_ | _922_ /*6588*/;
  assign _924_ = ~q[12] /*6587*/;
  assign _925_ = sum_4[29] & q[12] /*6586*/;
  assign _926_ = m_4[29] & _924_ /*6585*/;
  assign r_4[29] = _926_ | _925_ /*6584*/;
  assign _927_ = ~q[12] /*6583*/;
  assign _928_ = sum_4[30] & q[12] /*6582*/;
  assign _929_ = m_4[30] & _927_ /*6581*/;
  assign r_4[30] = _929_ | _928_ /*6580*/;
  assign _930_ = ~q[12] /*6579*/;
  assign _931_ = sum_4[31] & q[12] /*6578*/;
  assign _932_ = m_4[31] & _930_ /*6577*/;
  assign r_4[31] = _932_ | _931_ /*6576*/;
  assign _933_ = ~q[12] /*6575*/;
  assign _934_ = sum_4[32] & q[12] /*6574*/;
  assign _935_ = m_4[32] & _933_ /*6573*/;
  assign r_4[32] = _935_ | _934_ /*6572*/;
  assign _936_ = ~q[12] /*6571*/;
  assign _937_ = sum_4[33] & q[12] /*6570*/;
  assign _938_ = m_4[33] & _936_ /*6569*/;
  assign r_4[33] = _938_ | _937_ /*6568*/;
  assign _939_ = ~q[12] /*6567*/;
  assign _940_ = sum_4[34] & q[12] /*6566*/;
  assign _941_ = m_4[34] & _939_ /*6565*/;
  assign r_4[34] = _941_ | _940_ /*6564*/;
  assign inv_5[0] = oneWire /*6416*/;
  assign inv_5[1] = oneWire /*6410*/;
  assign inv_5[2] = oneWire /*6404*/;
  assign inv_5[3] = oneWire /*6398*/;
  assign inv_5[4] = oneWire /*6392*/;
  assign inv_5[5] = oneWire /*6386*/;
  assign inv_5[6] = oneWire /*6380*/;
  assign inv_5[7] = oneWire /*6374*/;
  assign inv_5[8] = oneWire /*6368*/;
  assign inv_5[9] = oneWire /*6362*/;
  assign inv_5[10] = oneWire /*6356*/;
  assign inv_5[11] = ~div[0] /*6350*/;
  assign inv_5[12] = ~div[1] /*6344*/;
  assign inv_5[13] = ~div[2] /*6338*/;
  assign inv_5[14] = ~div[3] /*6332*/;
  assign inv_5[15] = ~div[4] /*6326*/;
  assign inv_5[16] = ~div[5] /*6320*/;
  assign inv_5[17] = ~div[6] /*6314*/;
  assign inv_5[18] = ~div[7] /*6308*/;
  assign inv_5[19] = ~div[8] /*6302*/;
  assign inv_5[20] = ~div[9] /*6296*/;
  assign inv_5[21] = ~div[10] /*6290*/;
  assign inv_5[22] = ~div[11] /*6284*/;
  assign inv_5[23] = ~div[12] /*6278*/;
  assign inv_5[24] = ~div[13] /*6272*/;
  assign inv_5[25] = ~div[14] /*6266*/;
  assign inv_5[26] = oneWire /*6260*/;
  assign inv_5[27] = oneWire /*6254*/;
  assign inv_5[28] = oneWire /*6248*/;
  assign inv_5[29] = oneWire /*6242*/;
  assign inv_5[30] = oneWire /*6236*/;
  assign inv_5[31] = oneWire /*6230*/;
  assign inv_5[32] = oneWire /*6224*/;
  assign inv_5[33] = oneWire /*6218*/;
  assign inv_5[34] = oneWire /*6212*/;
  assign _942_ = inv_5[0] ^ r_4[0] /*6415*/;
  assign sum_5[0] = _942_ ^ oneWire /*6414*/;
  assign _943_ = _942_ & oneWire /*6413*/;
  assign _944_ = inv_5[0] & r_4[0] /*6412*/;
  assign _945_ = _943_ | _944_ /*6411*/;
  assign _946_ = inv_5[1] ^ r_4[1] /*6409*/;
  assign sum_5[1] = _946_ ^ _945_ /*6408*/;
  assign _947_ = _946_ & _945_ /*6407*/;
  assign _948_ = inv_5[1] & r_4[1] /*6406*/;
  assign _949_ = _947_ | _948_ /*6405*/;
  assign _950_ = inv_5[2] ^ r_4[2] /*6403*/;
  assign sum_5[2] = _950_ ^ _949_ /*6402*/;
  assign _951_ = _950_ & _949_ /*6401*/;
  assign _952_ = inv_5[2] & r_4[2] /*6400*/;
  assign _953_ = _951_ | _952_ /*6399*/;
  assign _954_ = inv_5[3] ^ r_4[3] /*6397*/;
  assign sum_5[3] = _954_ ^ _953_ /*6396*/;
  assign _955_ = _954_ & _953_ /*6395*/;
  assign _956_ = inv_5[3] & r_4[3] /*6394*/;
  assign _957_ = _955_ | _956_ /*6393*/;
  assign _958_ = inv_5[4] ^ r_4[4] /*6391*/;
  assign sum_5[4] = _958_ ^ _957_ /*6390*/;
  assign _959_ = _958_ & _957_ /*6389*/;
  assign _960_ = inv_5[4] & r_4[4] /*6388*/;
  assign _961_ = _959_ | _960_ /*6387*/;
  assign _962_ = inv_5[5] ^ r_4[5] /*6385*/;
  assign sum_5[5] = _962_ ^ _961_ /*6384*/;
  assign _963_ = _962_ & _961_ /*6383*/;
  assign _964_ = inv_5[5] & r_4[5] /*6382*/;
  assign _965_ = _963_ | _964_ /*6381*/;
  assign _966_ = inv_5[6] ^ r_4[6] /*6379*/;
  assign sum_5[6] = _966_ ^ _965_ /*6378*/;
  assign _967_ = _966_ & _965_ /*6377*/;
  assign _968_ = inv_5[6] & r_4[6] /*6376*/;
  assign _969_ = _967_ | _968_ /*6375*/;
  assign _970_ = inv_5[7] ^ r_4[7] /*6373*/;
  assign sum_5[7] = _970_ ^ _969_ /*6372*/;
  assign _971_ = _970_ & _969_ /*6371*/;
  assign _972_ = inv_5[7] & r_4[7] /*6370*/;
  assign _973_ = _971_ | _972_ /*6369*/;
  assign _974_ = inv_5[8] ^ r_4[8] /*6367*/;
  assign sum_5[8] = _974_ ^ _973_ /*6366*/;
  assign _975_ = _974_ & _973_ /*6365*/;
  assign _976_ = inv_5[8] & r_4[8] /*6364*/;
  assign _977_ = _975_ | _976_ /*6363*/;
  assign _978_ = inv_5[9] ^ r_4[9] /*6361*/;
  assign sum_5[9] = _978_ ^ _977_ /*6360*/;
  assign _979_ = _978_ & _977_ /*6359*/;
  assign _980_ = inv_5[9] & r_4[9] /*6358*/;
  assign _981_ = _979_ | _980_ /*6357*/;
  assign _982_ = inv_5[10] ^ r_4[10] /*6355*/;
  assign sum_5[10] = _982_ ^ _981_ /*6354*/;
  assign _983_ = _982_ & _981_ /*6353*/;
  assign _984_ = inv_5[10] & r_4[10] /*6352*/;
  assign _985_ = _983_ | _984_ /*6351*/;
  assign _986_ = inv_5[11] ^ r_4[11] /*6349*/;
  assign sum_5[11] = _986_ ^ _985_ /*6348*/;
  assign _987_ = _986_ & _985_ /*6347*/;
  assign _988_ = inv_5[11] & r_4[11] /*6346*/;
  assign _989_ = _987_ | _988_ /*6345*/;
  assign _990_ = inv_5[12] ^ r_4[12] /*6343*/;
  assign sum_5[12] = _990_ ^ _989_ /*6342*/;
  assign _991_ = _990_ & _989_ /*6341*/;
  assign _992_ = inv_5[12] & r_4[12] /*6340*/;
  assign _993_ = _991_ | _992_ /*6339*/;
  assign _994_ = inv_5[13] ^ r_4[13] /*6337*/;
  assign sum_5[13] = _994_ ^ _993_ /*6336*/;
  assign _995_ = _994_ & _993_ /*6335*/;
  assign _996_ = inv_5[13] & r_4[13] /*6334*/;
  assign _997_ = _995_ | _996_ /*6333*/;
  assign _998_ = inv_5[14] ^ r_4[14] /*6331*/;
  assign sum_5[14] = _998_ ^ _997_ /*6330*/;
  assign _999_ = _998_ & _997_ /*6329*/;
  assign _1000_ = inv_5[14] & r_4[14] /*6328*/;
  assign _1001_ = _999_ | _1000_ /*6327*/;
  assign _1002_ = inv_5[15] ^ r_4[15] /*6325*/;
  assign sum_5[15] = _1002_ ^ _1001_ /*6324*/;
  assign _1003_ = _1002_ & _1001_ /*6323*/;
  assign _1004_ = inv_5[15] & r_4[15] /*6322*/;
  assign _1005_ = _1003_ | _1004_ /*6321*/;
  assign _1006_ = inv_5[16] ^ r_4[16] /*6319*/;
  assign sum_5[16] = _1006_ ^ _1005_ /*6318*/;
  assign _1007_ = _1006_ & _1005_ /*6317*/;
  assign _1008_ = inv_5[16] & r_4[16] /*6316*/;
  assign _1009_ = _1007_ | _1008_ /*6315*/;
  assign _1010_ = inv_5[17] ^ r_4[17] /*6313*/;
  assign sum_5[17] = _1010_ ^ _1009_ /*6312*/;
  assign _1011_ = _1010_ & _1009_ /*6311*/;
  assign _1012_ = inv_5[17] & r_4[17] /*6310*/;
  assign _1013_ = _1011_ | _1012_ /*6309*/;
  assign _1014_ = inv_5[18] ^ r_4[18] /*6307*/;
  assign sum_5[18] = _1014_ ^ _1013_ /*6306*/;
  assign _1015_ = _1014_ & _1013_ /*6305*/;
  assign _1016_ = inv_5[18] & r_4[18] /*6304*/;
  assign _1017_ = _1015_ | _1016_ /*6303*/;
  assign _1018_ = inv_5[19] ^ r_4[19] /*6301*/;
  assign sum_5[19] = _1018_ ^ _1017_ /*6300*/;
  assign _1019_ = _1018_ & _1017_ /*6299*/;
  assign _1020_ = inv_5[19] & r_4[19] /*6298*/;
  assign _1021_ = _1019_ | _1020_ /*6297*/;
  assign _1022_ = inv_5[20] ^ r_4[20] /*6295*/;
  assign sum_5[20] = _1022_ ^ _1021_ /*6294*/;
  assign _1023_ = _1022_ & _1021_ /*6293*/;
  assign _1024_ = inv_5[20] & r_4[20] /*6292*/;
  assign _1025_ = _1023_ | _1024_ /*6291*/;
  assign _1026_ = inv_5[21] ^ r_4[21] /*6289*/;
  assign sum_5[21] = _1026_ ^ _1025_ /*6288*/;
  assign _1027_ = _1026_ & _1025_ /*6287*/;
  assign _1028_ = inv_5[21] & r_4[21] /*6286*/;
  assign _1029_ = _1027_ | _1028_ /*6285*/;
  assign _1030_ = inv_5[22] ^ r_4[22] /*6283*/;
  assign sum_5[22] = _1030_ ^ _1029_ /*6282*/;
  assign _1031_ = _1030_ & _1029_ /*6281*/;
  assign _1032_ = inv_5[22] & r_4[22] /*6280*/;
  assign _1033_ = _1031_ | _1032_ /*6279*/;
  assign _1034_ = inv_5[23] ^ r_4[23] /*6277*/;
  assign sum_5[23] = _1034_ ^ _1033_ /*6276*/;
  assign _1035_ = _1034_ & _1033_ /*6275*/;
  assign _1036_ = inv_5[23] & r_4[23] /*6274*/;
  assign _1037_ = _1035_ | _1036_ /*6273*/;
  assign _1038_ = inv_5[24] ^ r_4[24] /*6271*/;
  assign sum_5[24] = _1038_ ^ _1037_ /*6270*/;
  assign _1039_ = _1038_ & _1037_ /*6269*/;
  assign _1040_ = inv_5[24] & r_4[24] /*6268*/;
  assign _1041_ = _1039_ | _1040_ /*6267*/;
  assign _1042_ = inv_5[25] ^ r_4[25] /*6265*/;
  assign sum_5[25] = _1042_ ^ _1041_ /*6264*/;
  assign _1043_ = _1042_ & _1041_ /*6263*/;
  assign _1044_ = inv_5[25] & r_4[25] /*6262*/;
  assign _1045_ = _1043_ | _1044_ /*6261*/;
  assign _1046_ = inv_5[26] ^ r_4[26] /*6259*/;
  assign sum_5[26] = _1046_ ^ _1045_ /*6258*/;
  assign _1047_ = _1046_ & _1045_ /*6257*/;
  assign _1048_ = inv_5[26] & r_4[26] /*6256*/;
  assign _1049_ = _1047_ | _1048_ /*6255*/;
  assign _1050_ = inv_5[27] ^ r_4[27] /*6253*/;
  assign sum_5[27] = _1050_ ^ _1049_ /*6252*/;
  assign _1051_ = _1050_ & _1049_ /*6251*/;
  assign _1052_ = inv_5[27] & r_4[27] /*6250*/;
  assign _1053_ = _1051_ | _1052_ /*6249*/;
  assign _1054_ = inv_5[28] ^ r_4[28] /*6247*/;
  assign sum_5[28] = _1054_ ^ _1053_ /*6246*/;
  assign _1055_ = _1054_ & _1053_ /*6245*/;
  assign _1056_ = inv_5[28] & r_4[28] /*6244*/;
  assign _1057_ = _1055_ | _1056_ /*6243*/;
  assign _1058_ = inv_5[29] ^ r_4[29] /*6241*/;
  assign sum_5[29] = _1058_ ^ _1057_ /*6240*/;
  assign _1059_ = _1058_ & _1057_ /*6239*/;
  assign _1060_ = inv_5[29] & r_4[29] /*6238*/;
  assign _1061_ = _1059_ | _1060_ /*6237*/;
  assign _1062_ = inv_5[30] ^ r_4[30] /*6235*/;
  assign sum_5[30] = _1062_ ^ _1061_ /*6234*/;
  assign _1063_ = _1062_ & _1061_ /*6233*/;
  assign _1064_ = inv_5[30] & r_4[30] /*6232*/;
  assign _1065_ = _1063_ | _1064_ /*6231*/;
  assign _1066_ = inv_5[31] ^ r_4[31] /*6229*/;
  assign sum_5[31] = _1066_ ^ _1065_ /*6228*/;
  assign _1067_ = _1066_ & _1065_ /*6227*/;
  assign _1068_ = inv_5[31] & r_4[31] /*6226*/;
  assign _1069_ = _1067_ | _1068_ /*6225*/;
  assign _1070_ = inv_5[32] ^ r_4[32] /*6223*/;
  assign sum_5[32] = _1070_ ^ _1069_ /*6222*/;
  assign _1071_ = _1070_ & _1069_ /*6221*/;
  assign _1072_ = inv_5[32] & r_4[32] /*6220*/;
  assign _1073_ = _1071_ | _1072_ /*6219*/;
  assign _1074_ = inv_5[33] ^ r_4[33] /*6217*/;
  assign sum_5[33] = _1074_ ^ _1073_ /*6216*/;
  assign _1075_ = _1074_ & _1073_ /*6215*/;
  assign _1076_ = inv_5[33] & r_4[33] /*6214*/;
  assign _1077_ = _1075_ | _1076_ /*6213*/;
  assign _1078_ = inv_5[34] ^ r_4[34] /*6211*/;
  assign sum_5[34] = _1078_ ^ _1077_ /*6210*/;
  assign _1079_ = _1078_ & _1077_ /*6209*/;
  assign _1080_ = inv_5[34] & r_4[34] /*6208*/;
  assign _1081_ = _1079_ | _1080_ /*6207*/;
  assign _1082_ = _1081_ ^ _1077_ /*6206*/;
  assign _1083_ = ~_1082_ /*6205*/;
  assign _1084_ = sum_5[34] & _1083_ /*6204*/;
  assign _1085_ = _1082_ & _1081_ /*6203*/;
  assign sum_5[35] = _1085_ | _1084_ /*6202*/;
  assign q[11] = ~sum_5[35] /*6201*/;
  assign m_5[0] = r_4[0] /*6200*/;
  assign m_5[1] = r_4[1] /*6199*/;
  assign m_5[2] = r_4[2] /*6198*/;
  assign m_5[3] = r_4[3] /*6197*/;
  assign m_5[4] = r_4[4] /*6196*/;
  assign m_5[5] = r_4[5] /*6195*/;
  assign m_5[6] = r_4[6] /*6194*/;
  assign m_5[7] = r_4[7] /*6193*/;
  assign m_5[8] = r_4[8] /*6192*/;
  assign m_5[9] = r_4[9] /*6191*/;
  assign m_5[10] = r_4[10] /*6190*/;
  assign m_5[11] = r_4[11] /*6189*/;
  assign m_5[12] = r_4[12] /*6188*/;
  assign m_5[13] = r_4[13] /*6187*/;
  assign m_5[14] = r_4[14] /*6186*/;
  assign m_5[15] = r_4[15] /*6185*/;
  assign m_5[16] = r_4[16] /*6184*/;
  assign m_5[17] = r_4[17] /*6183*/;
  assign m_5[18] = r_4[18] /*6182*/;
  assign m_5[19] = r_4[19] /*6181*/;
  assign m_5[20] = r_4[20] /*6180*/;
  assign m_5[21] = r_4[21] /*6179*/;
  assign m_5[22] = r_4[22] /*6178*/;
  assign m_5[23] = r_4[23] /*6177*/;
  assign m_5[24] = r_4[24] /*6176*/;
  assign m_5[25] = r_4[25] /*6175*/;
  assign m_5[26] = r_4[26] /*6174*/;
  assign m_5[27] = r_4[27] /*6173*/;
  assign m_5[28] = r_4[28] /*6172*/;
  assign m_5[29] = r_4[29] /*6171*/;
  assign m_5[30] = r_4[30] /*6170*/;
  assign m_5[31] = r_4[31] /*6169*/;
  assign m_5[32] = r_4[32] /*6168*/;
  assign m_5[33] = r_4[33] /*6167*/;
  assign m_5[34] = r_4[34] /*6166*/;
  assign m_5[35] = r_4[34] /*6165*/;
  assign _1087_ = ~q[11] /*6164*/;
  assign _1088_ = sum_5[0] & q[11] /*6163*/;
  assign _1089_ = m_5[0] & _1087_ /*6162*/;
  assign r_5[0] = _1089_ | _1088_ /*6161*/;
  assign _1090_ = ~q[11] /*6160*/;
  assign _1091_ = sum_5[1] & q[11] /*6159*/;
  assign _1092_ = m_5[1] & _1090_ /*6158*/;
  assign r_5[1] = _1092_ | _1091_ /*6157*/;
  assign _1093_ = ~q[11] /*6156*/;
  assign _1094_ = sum_5[2] & q[11] /*6155*/;
  assign _1095_ = m_5[2] & _1093_ /*6154*/;
  assign r_5[2] = _1095_ | _1094_ /*6153*/;
  assign _1096_ = ~q[11] /*6152*/;
  assign _1097_ = sum_5[3] & q[11] /*6151*/;
  assign _1098_ = m_5[3] & _1096_ /*6150*/;
  assign r_5[3] = _1098_ | _1097_ /*6149*/;
  assign _1099_ = ~q[11] /*6148*/;
  assign _1100_ = sum_5[4] & q[11] /*6147*/;
  assign _1101_ = m_5[4] & _1099_ /*6146*/;
  assign r_5[4] = _1101_ | _1100_ /*6145*/;
  assign _1102_ = ~q[11] /*6144*/;
  assign _1103_ = sum_5[5] & q[11] /*6143*/;
  assign _1104_ = m_5[5] & _1102_ /*6142*/;
  assign r_5[5] = _1104_ | _1103_ /*6141*/;
  assign _1105_ = ~q[11] /*6140*/;
  assign _1106_ = sum_5[6] & q[11] /*6139*/;
  assign _1107_ = m_5[6] & _1105_ /*6138*/;
  assign r_5[6] = _1107_ | _1106_ /*6137*/;
  assign _1108_ = ~q[11] /*6136*/;
  assign _1109_ = sum_5[7] & q[11] /*6135*/;
  assign _1110_ = m_5[7] & _1108_ /*6134*/;
  assign r_5[7] = _1110_ | _1109_ /*6133*/;
  assign _1111_ = ~q[11] /*6132*/;
  assign _1112_ = sum_5[8] & q[11] /*6131*/;
  assign _1113_ = m_5[8] & _1111_ /*6130*/;
  assign r_5[8] = _1113_ | _1112_ /*6129*/;
  assign _1114_ = ~q[11] /*6128*/;
  assign _1115_ = sum_5[9] & q[11] /*6127*/;
  assign _1116_ = m_5[9] & _1114_ /*6126*/;
  assign r_5[9] = _1116_ | _1115_ /*6125*/;
  assign _1117_ = ~q[11] /*6124*/;
  assign _1118_ = sum_5[10] & q[11] /*6123*/;
  assign _1119_ = m_5[10] & _1117_ /*6122*/;
  assign r_5[10] = _1119_ | _1118_ /*6121*/;
  assign _1120_ = ~q[11] /*6120*/;
  assign _1121_ = sum_5[11] & q[11] /*6119*/;
  assign _1122_ = m_5[11] & _1120_ /*6118*/;
  assign r_5[11] = _1122_ | _1121_ /*6117*/;
  assign _1123_ = ~q[11] /*6116*/;
  assign _1124_ = sum_5[12] & q[11] /*6115*/;
  assign _1125_ = m_5[12] & _1123_ /*6114*/;
  assign r_5[12] = _1125_ | _1124_ /*6113*/;
  assign _1126_ = ~q[11] /*6112*/;
  assign _1127_ = sum_5[13] & q[11] /*6111*/;
  assign _1128_ = m_5[13] & _1126_ /*6110*/;
  assign r_5[13] = _1128_ | _1127_ /*6109*/;
  assign _1129_ = ~q[11] /*6108*/;
  assign _1130_ = sum_5[14] & q[11] /*6107*/;
  assign _1131_ = m_5[14] & _1129_ /*6106*/;
  assign r_5[14] = _1131_ | _1130_ /*6105*/;
  assign _1132_ = ~q[11] /*6104*/;
  assign _1133_ = sum_5[15] & q[11] /*6103*/;
  assign _1134_ = m_5[15] & _1132_ /*6102*/;
  assign r_5[15] = _1134_ | _1133_ /*6101*/;
  assign _1135_ = ~q[11] /*6100*/;
  assign _1136_ = sum_5[16] & q[11] /*6099*/;
  assign _1137_ = m_5[16] & _1135_ /*6098*/;
  assign r_5[16] = _1137_ | _1136_ /*6097*/;
  assign _1138_ = ~q[11] /*6096*/;
  assign _1139_ = sum_5[17] & q[11] /*6095*/;
  assign _1140_ = m_5[17] & _1138_ /*6094*/;
  assign r_5[17] = _1140_ | _1139_ /*6093*/;
  assign _1141_ = ~q[11] /*6092*/;
  assign _1142_ = sum_5[18] & q[11] /*6091*/;
  assign _1143_ = m_5[18] & _1141_ /*6090*/;
  assign r_5[18] = _1143_ | _1142_ /*6089*/;
  assign _1144_ = ~q[11] /*6088*/;
  assign _1145_ = sum_5[19] & q[11] /*6087*/;
  assign _1146_ = m_5[19] & _1144_ /*6086*/;
  assign r_5[19] = _1146_ | _1145_ /*6085*/;
  assign _1147_ = ~q[11] /*6084*/;
  assign _1148_ = sum_5[20] & q[11] /*6083*/;
  assign _1149_ = m_5[20] & _1147_ /*6082*/;
  assign r_5[20] = _1149_ | _1148_ /*6081*/;
  assign _1150_ = ~q[11] /*6080*/;
  assign _1151_ = sum_5[21] & q[11] /*6079*/;
  assign _1152_ = m_5[21] & _1150_ /*6078*/;
  assign r_5[21] = _1152_ | _1151_ /*6077*/;
  assign _1153_ = ~q[11] /*6076*/;
  assign _1154_ = sum_5[22] & q[11] /*6075*/;
  assign _1155_ = m_5[22] & _1153_ /*6074*/;
  assign r_5[22] = _1155_ | _1154_ /*6073*/;
  assign _1156_ = ~q[11] /*6072*/;
  assign _1157_ = sum_5[23] & q[11] /*6071*/;
  assign _1158_ = m_5[23] & _1156_ /*6070*/;
  assign r_5[23] = _1158_ | _1157_ /*6069*/;
  assign _1159_ = ~q[11] /*6068*/;
  assign _1160_ = sum_5[24] & q[11] /*6067*/;
  assign _1161_ = m_5[24] & _1159_ /*6066*/;
  assign r_5[24] = _1161_ | _1160_ /*6065*/;
  assign _1162_ = ~q[11] /*6064*/;
  assign _1163_ = sum_5[25] & q[11] /*6063*/;
  assign _1164_ = m_5[25] & _1162_ /*6062*/;
  assign r_5[25] = _1164_ | _1163_ /*6061*/;
  assign _1165_ = ~q[11] /*6060*/;
  assign _1166_ = sum_5[26] & q[11] /*6059*/;
  assign _1167_ = m_5[26] & _1165_ /*6058*/;
  assign r_5[26] = _1167_ | _1166_ /*6057*/;
  assign _1168_ = ~q[11] /*6056*/;
  assign _1169_ = sum_5[27] & q[11] /*6055*/;
  assign _1170_ = m_5[27] & _1168_ /*6054*/;
  assign r_5[27] = _1170_ | _1169_ /*6053*/;
  assign _1171_ = ~q[11] /*6052*/;
  assign _1172_ = sum_5[28] & q[11] /*6051*/;
  assign _1173_ = m_5[28] & _1171_ /*6050*/;
  assign r_5[28] = _1173_ | _1172_ /*6049*/;
  assign _1174_ = ~q[11] /*6048*/;
  assign _1175_ = sum_5[29] & q[11] /*6047*/;
  assign _1176_ = m_5[29] & _1174_ /*6046*/;
  assign r_5[29] = _1176_ | _1175_ /*6045*/;
  assign _1177_ = ~q[11] /*6044*/;
  assign _1178_ = sum_5[30] & q[11] /*6043*/;
  assign _1179_ = m_5[30] & _1177_ /*6042*/;
  assign r_5[30] = _1179_ | _1178_ /*6041*/;
  assign _1180_ = ~q[11] /*6040*/;
  assign _1181_ = sum_5[31] & q[11] /*6039*/;
  assign _1182_ = m_5[31] & _1180_ /*6038*/;
  assign r_5[31] = _1182_ | _1181_ /*6037*/;
  assign _1183_ = ~q[11] /*6036*/;
  assign _1184_ = sum_5[32] & q[11] /*6035*/;
  assign _1185_ = m_5[32] & _1183_ /*6034*/;
  assign r_5[32] = _1185_ | _1184_ /*6033*/;
  assign _1186_ = ~q[11] /*6032*/;
  assign _1187_ = sum_5[33] & q[11] /*6031*/;
  assign _1188_ = m_5[33] & _1186_ /*6030*/;
  assign r_5[33] = _1188_ | _1187_ /*6029*/;
  assign _1189_ = ~q[11] /*6028*/;
  assign _1190_ = sum_5[34] & q[11] /*6027*/;
  assign _1191_ = m_5[34] & _1189_ /*6026*/;
  assign r_5[34] = _1191_ | _1190_ /*6025*/;
  assign _1192_ = ~q[11] /*6024*/;
  assign _1193_ = sum_5[35] & q[11] /*6023*/;
  assign _1194_ = m_5[35] & _1192_ /*6022*/;
  assign r_5[35] = _1194_ | _1193_ /*6021*/;
  assign inv_6[0] = oneWire /*5884*/;
  assign inv_6[1] = oneWire /*5878*/;
  assign inv_6[2] = oneWire /*5872*/;
  assign inv_6[3] = oneWire /*5866*/;
  assign inv_6[4] = oneWire /*5860*/;
  assign inv_6[5] = oneWire /*5854*/;
  assign inv_6[6] = oneWire /*5848*/;
  assign inv_6[7] = oneWire /*5842*/;
  assign inv_6[8] = oneWire /*5836*/;
  assign inv_6[9] = oneWire /*5830*/;
  assign inv_6[10] = ~div[0] /*5824*/;
  assign inv_6[11] = ~div[1] /*5818*/;
  assign inv_6[12] = ~div[2] /*5812*/;
  assign inv_6[13] = ~div[3] /*5806*/;
  assign inv_6[14] = ~div[4] /*5800*/;
  assign inv_6[15] = ~div[5] /*5794*/;
  assign inv_6[16] = ~div[6] /*5788*/;
  assign inv_6[17] = ~div[7] /*5782*/;
  assign inv_6[18] = ~div[8] /*5776*/;
  assign inv_6[19] = ~div[9] /*5770*/;
  assign inv_6[20] = ~div[10] /*5764*/;
  assign inv_6[21] = ~div[11] /*5758*/;
  assign inv_6[22] = ~div[12] /*5752*/;
  assign inv_6[23] = ~div[13] /*5746*/;
  assign inv_6[24] = ~div[14] /*5740*/;
  assign inv_6[25] = oneWire /*5734*/;
  assign inv_6[26] = oneWire /*5728*/;
  assign inv_6[27] = oneWire /*5722*/;
  assign inv_6[28] = oneWire /*5716*/;
  assign inv_6[29] = oneWire /*5710*/;
  assign inv_6[30] = oneWire /*5704*/;
  assign inv_6[31] = oneWire /*5698*/;
  assign inv_6[32] = oneWire /*5692*/;
  assign inv_6[33] = oneWire /*5686*/;
  assign inv_6[34] = oneWire /*5680*/;
  assign inv_6[35] = oneWire /*5674*/;
  assign _1195_ = inv_6[0] ^ r_5[0] /*5883*/;
  assign sum_6[0] = _1195_ ^ oneWire /*5882*/;
  assign _1196_ = _1195_ & oneWire /*5881*/;
  assign _1197_ = inv_6[0] & r_5[0] /*5880*/;
  assign _1198_ = _1196_ | _1197_ /*5879*/;
  assign _1199_ = inv_6[1] ^ r_5[1] /*5877*/;
  assign sum_6[1] = _1199_ ^ _1198_ /*5876*/;
  assign _1200_ = _1199_ & _1198_ /*5875*/;
  assign _1201_ = inv_6[1] & r_5[1] /*5874*/;
  assign _1202_ = _1200_ | _1201_ /*5873*/;
  assign _1203_ = inv_6[2] ^ r_5[2] /*5871*/;
  assign sum_6[2] = _1203_ ^ _1202_ /*5870*/;
  assign _1204_ = _1203_ & _1202_ /*5869*/;
  assign _1205_ = inv_6[2] & r_5[2] /*5868*/;
  assign _1206_ = _1204_ | _1205_ /*5867*/;
  assign _1207_ = inv_6[3] ^ r_5[3] /*5865*/;
  assign sum_6[3] = _1207_ ^ _1206_ /*5864*/;
  assign _1208_ = _1207_ & _1206_ /*5863*/;
  assign _1209_ = inv_6[3] & r_5[3] /*5862*/;
  assign _1210_ = _1208_ | _1209_ /*5861*/;
  assign _1211_ = inv_6[4] ^ r_5[4] /*5859*/;
  assign sum_6[4] = _1211_ ^ _1210_ /*5858*/;
  assign _1212_ = _1211_ & _1210_ /*5857*/;
  assign _1213_ = inv_6[4] & r_5[4] /*5856*/;
  assign _1214_ = _1212_ | _1213_ /*5855*/;
  assign _1215_ = inv_6[5] ^ r_5[5] /*5853*/;
  assign sum_6[5] = _1215_ ^ _1214_ /*5852*/;
  assign _1216_ = _1215_ & _1214_ /*5851*/;
  assign _1217_ = inv_6[5] & r_5[5] /*5850*/;
  assign _1218_ = _1216_ | _1217_ /*5849*/;
  assign _1219_ = inv_6[6] ^ r_5[6] /*5847*/;
  assign sum_6[6] = _1219_ ^ _1218_ /*5846*/;
  assign _1220_ = _1219_ & _1218_ /*5845*/;
  assign _1221_ = inv_6[6] & r_5[6] /*5844*/;
  assign _1222_ = _1220_ | _1221_ /*5843*/;
  assign _1223_ = inv_6[7] ^ r_5[7] /*5841*/;
  assign sum_6[7] = _1223_ ^ _1222_ /*5840*/;
  assign _1224_ = _1223_ & _1222_ /*5839*/;
  assign _1225_ = inv_6[7] & r_5[7] /*5838*/;
  assign _1226_ = _1224_ | _1225_ /*5837*/;
  assign _1227_ = inv_6[8] ^ r_5[8] /*5835*/;
  assign sum_6[8] = _1227_ ^ _1226_ /*5834*/;
  assign _1228_ = _1227_ & _1226_ /*5833*/;
  assign _1229_ = inv_6[8] & r_5[8] /*5832*/;
  assign _1230_ = _1228_ | _1229_ /*5831*/;
  assign _1231_ = inv_6[9] ^ r_5[9] /*5829*/;
  assign sum_6[9] = _1231_ ^ _1230_ /*5828*/;
  assign _1232_ = _1231_ & _1230_ /*5827*/;
  assign _1233_ = inv_6[9] & r_5[9] /*5826*/;
  assign _1234_ = _1232_ | _1233_ /*5825*/;
  assign _1235_ = inv_6[10] ^ r_5[10] /*5823*/;
  assign sum_6[10] = _1235_ ^ _1234_ /*5822*/;
  assign _1236_ = _1235_ & _1234_ /*5821*/;
  assign _1237_ = inv_6[10] & r_5[10] /*5820*/;
  assign _1238_ = _1236_ | _1237_ /*5819*/;
  assign _1239_ = inv_6[11] ^ r_5[11] /*5817*/;
  assign sum_6[11] = _1239_ ^ _1238_ /*5816*/;
  assign _1240_ = _1239_ & _1238_ /*5815*/;
  assign _1241_ = inv_6[11] & r_5[11] /*5814*/;
  assign _1242_ = _1240_ | _1241_ /*5813*/;
  assign _1243_ = inv_6[12] ^ r_5[12] /*5811*/;
  assign sum_6[12] = _1243_ ^ _1242_ /*5810*/;
  assign _1244_ = _1243_ & _1242_ /*5809*/;
  assign _1245_ = inv_6[12] & r_5[12] /*5808*/;
  assign _1246_ = _1244_ | _1245_ /*5807*/;
  assign _1247_ = inv_6[13] ^ r_5[13] /*5805*/;
  assign sum_6[13] = _1247_ ^ _1246_ /*5804*/;
  assign _1248_ = _1247_ & _1246_ /*5803*/;
  assign _1249_ = inv_6[13] & r_5[13] /*5802*/;
  assign _1250_ = _1248_ | _1249_ /*5801*/;
  assign _1251_ = inv_6[14] ^ r_5[14] /*5799*/;
  assign sum_6[14] = _1251_ ^ _1250_ /*5798*/;
  assign _1252_ = _1251_ & _1250_ /*5797*/;
  assign _1253_ = inv_6[14] & r_5[14] /*5796*/;
  assign _1254_ = _1252_ | _1253_ /*5795*/;
  assign _1255_ = inv_6[15] ^ r_5[15] /*5793*/;
  assign sum_6[15] = _1255_ ^ _1254_ /*5792*/;
  assign _1256_ = _1255_ & _1254_ /*5791*/;
  assign _1257_ = inv_6[15] & r_5[15] /*5790*/;
  assign _1258_ = _1256_ | _1257_ /*5789*/;
  assign _1259_ = inv_6[16] ^ r_5[16] /*5787*/;
  assign sum_6[16] = _1259_ ^ _1258_ /*5786*/;
  assign _1260_ = _1259_ & _1258_ /*5785*/;
  assign _1261_ = inv_6[16] & r_5[16] /*5784*/;
  assign _1262_ = _1260_ | _1261_ /*5783*/;
  assign _1263_ = inv_6[17] ^ r_5[17] /*5781*/;
  assign sum_6[17] = _1263_ ^ _1262_ /*5780*/;
  assign _1264_ = _1263_ & _1262_ /*5779*/;
  assign _1265_ = inv_6[17] & r_5[17] /*5778*/;
  assign _1266_ = _1264_ | _1265_ /*5777*/;
  assign _1267_ = inv_6[18] ^ r_5[18] /*5775*/;
  assign sum_6[18] = _1267_ ^ _1266_ /*5774*/;
  assign _1268_ = _1267_ & _1266_ /*5773*/;
  assign _1269_ = inv_6[18] & r_5[18] /*5772*/;
  assign _1270_ = _1268_ | _1269_ /*5771*/;
  assign _1271_ = inv_6[19] ^ r_5[19] /*5769*/;
  assign sum_6[19] = _1271_ ^ _1270_ /*5768*/;
  assign _1272_ = _1271_ & _1270_ /*5767*/;
  assign _1273_ = inv_6[19] & r_5[19] /*5766*/;
  assign _1274_ = _1272_ | _1273_ /*5765*/;
  assign _1275_ = inv_6[20] ^ r_5[20] /*5763*/;
  assign sum_6[20] = _1275_ ^ _1274_ /*5762*/;
  assign _1276_ = _1275_ & _1274_ /*5761*/;
  assign _1277_ = inv_6[20] & r_5[20] /*5760*/;
  assign _1278_ = _1276_ | _1277_ /*5759*/;
  assign _1279_ = inv_6[21] ^ r_5[21] /*5757*/;
  assign sum_6[21] = _1279_ ^ _1278_ /*5756*/;
  assign _1280_ = _1279_ & _1278_ /*5755*/;
  assign _1281_ = inv_6[21] & r_5[21] /*5754*/;
  assign _1282_ = _1280_ | _1281_ /*5753*/;
  assign _1283_ = inv_6[22] ^ r_5[22] /*5751*/;
  assign sum_6[22] = _1283_ ^ _1282_ /*5750*/;
  assign _1284_ = _1283_ & _1282_ /*5749*/;
  assign _1285_ = inv_6[22] & r_5[22] /*5748*/;
  assign _1286_ = _1284_ | _1285_ /*5747*/;
  assign _1287_ = inv_6[23] ^ r_5[23] /*5745*/;
  assign sum_6[23] = _1287_ ^ _1286_ /*5744*/;
  assign _1288_ = _1287_ & _1286_ /*5743*/;
  assign _1289_ = inv_6[23] & r_5[23] /*5742*/;
  assign _1290_ = _1288_ | _1289_ /*5741*/;
  assign _1291_ = inv_6[24] ^ r_5[24] /*5739*/;
  assign sum_6[24] = _1291_ ^ _1290_ /*5738*/;
  assign _1292_ = _1291_ & _1290_ /*5737*/;
  assign _1293_ = inv_6[24] & r_5[24] /*5736*/;
  assign _1294_ = _1292_ | _1293_ /*5735*/;
  assign _1295_ = inv_6[25] ^ r_5[25] /*5733*/;
  assign sum_6[25] = _1295_ ^ _1294_ /*5732*/;
  assign _1296_ = _1295_ & _1294_ /*5731*/;
  assign _1297_ = inv_6[25] & r_5[25] /*5730*/;
  assign _1298_ = _1296_ | _1297_ /*5729*/;
  assign _1299_ = inv_6[26] ^ r_5[26] /*5727*/;
  assign sum_6[26] = _1299_ ^ _1298_ /*5726*/;
  assign _1300_ = _1299_ & _1298_ /*5725*/;
  assign _1301_ = inv_6[26] & r_5[26] /*5724*/;
  assign _1302_ = _1300_ | _1301_ /*5723*/;
  assign _1303_ = inv_6[27] ^ r_5[27] /*5721*/;
  assign sum_6[27] = _1303_ ^ _1302_ /*5720*/;
  assign _1304_ = _1303_ & _1302_ /*5719*/;
  assign _1305_ = inv_6[27] & r_5[27] /*5718*/;
  assign _1306_ = _1304_ | _1305_ /*5717*/;
  assign _1307_ = inv_6[28] ^ r_5[28] /*5715*/;
  assign sum_6[28] = _1307_ ^ _1306_ /*5714*/;
  assign _1308_ = _1307_ & _1306_ /*5713*/;
  assign _1309_ = inv_6[28] & r_5[28] /*5712*/;
  assign _1310_ = _1308_ | _1309_ /*5711*/;
  assign _1311_ = inv_6[29] ^ r_5[29] /*5709*/;
  assign sum_6[29] = _1311_ ^ _1310_ /*5708*/;
  assign _1312_ = _1311_ & _1310_ /*5707*/;
  assign _1313_ = inv_6[29] & r_5[29] /*5706*/;
  assign _1314_ = _1312_ | _1313_ /*5705*/;
  assign _1315_ = inv_6[30] ^ r_5[30] /*5703*/;
  assign sum_6[30] = _1315_ ^ _1314_ /*5702*/;
  assign _1316_ = _1315_ & _1314_ /*5701*/;
  assign _1317_ = inv_6[30] & r_5[30] /*5700*/;
  assign _1318_ = _1316_ | _1317_ /*5699*/;
  assign _1319_ = inv_6[31] ^ r_5[31] /*5697*/;
  assign sum_6[31] = _1319_ ^ _1318_ /*5696*/;
  assign _1320_ = _1319_ & _1318_ /*5695*/;
  assign _1321_ = inv_6[31] & r_5[31] /*5694*/;
  assign _1322_ = _1320_ | _1321_ /*5693*/;
  assign _1323_ = inv_6[32] ^ r_5[32] /*5691*/;
  assign sum_6[32] = _1323_ ^ _1322_ /*5690*/;
  assign _1324_ = _1323_ & _1322_ /*5689*/;
  assign _1325_ = inv_6[32] & r_5[32] /*5688*/;
  assign _1326_ = _1324_ | _1325_ /*5687*/;
  assign _1327_ = inv_6[33] ^ r_5[33] /*5685*/;
  assign sum_6[33] = _1327_ ^ _1326_ /*5684*/;
  assign _1328_ = _1327_ & _1326_ /*5683*/;
  assign _1329_ = inv_6[33] & r_5[33] /*5682*/;
  assign _1330_ = _1328_ | _1329_ /*5681*/;
  assign _1331_ = inv_6[34] ^ r_5[34] /*5679*/;
  assign sum_6[34] = _1331_ ^ _1330_ /*5678*/;
  assign _1332_ = _1331_ & _1330_ /*5677*/;
  assign _1333_ = inv_6[34] & r_5[34] /*5676*/;
  assign _1334_ = _1332_ | _1333_ /*5675*/;
  assign _1335_ = inv_6[35] ^ r_5[35] /*5673*/;
  assign sum_6[35] = _1335_ ^ _1334_ /*5672*/;
  assign _1336_ = _1335_ & _1334_ /*5671*/;
  assign _1337_ = inv_6[35] & r_5[35] /*5670*/;
  assign _1338_ = _1336_ | _1337_ /*5669*/;
  assign _1339_ = _1338_ ^ _1334_ /*5668*/;
  assign _1340_ = ~_1339_ /*5667*/;
  assign _1341_ = sum_6[35] & _1340_ /*5666*/;
  assign _1342_ = _1339_ & _1338_ /*5665*/;
  assign sum_6[36] = _1342_ | _1341_ /*5664*/;
  assign q[10] = ~sum_6[36] /*5663*/;
  assign m_6[0] = r_5[0] /*5662*/;
  assign m_6[1] = r_5[1] /*5661*/;
  assign m_6[2] = r_5[2] /*5660*/;
  assign m_6[3] = r_5[3] /*5659*/;
  assign m_6[4] = r_5[4] /*5658*/;
  assign m_6[5] = r_5[5] /*5657*/;
  assign m_6[6] = r_5[6] /*5656*/;
  assign m_6[7] = r_5[7] /*5655*/;
  assign m_6[8] = r_5[8] /*5654*/;
  assign m_6[9] = r_5[9] /*5653*/;
  assign m_6[10] = r_5[10] /*5652*/;
  assign m_6[11] = r_5[11] /*5651*/;
  assign m_6[12] = r_5[12] /*5650*/;
  assign m_6[13] = r_5[13] /*5649*/;
  assign m_6[14] = r_5[14] /*5648*/;
  assign m_6[15] = r_5[15] /*5647*/;
  assign m_6[16] = r_5[16] /*5646*/;
  assign m_6[17] = r_5[17] /*5645*/;
  assign m_6[18] = r_5[18] /*5644*/;
  assign m_6[19] = r_5[19] /*5643*/;
  assign m_6[20] = r_5[20] /*5642*/;
  assign m_6[21] = r_5[21] /*5641*/;
  assign m_6[22] = r_5[22] /*5640*/;
  assign m_6[23] = r_5[23] /*5639*/;
  assign m_6[24] = r_5[24] /*5638*/;
  assign m_6[25] = r_5[25] /*5637*/;
  assign m_6[26] = r_5[26] /*5636*/;
  assign m_6[27] = r_5[27] /*5635*/;
  assign m_6[28] = r_5[28] /*5634*/;
  assign m_6[29] = r_5[29] /*5633*/;
  assign m_6[30] = r_5[30] /*5632*/;
  assign m_6[31] = r_5[31] /*5631*/;
  assign m_6[32] = r_5[32] /*5630*/;
  assign m_6[33] = r_5[33] /*5629*/;
  assign m_6[34] = r_5[34] /*5628*/;
  assign m_6[35] = r_5[35] /*5627*/;
  assign m_6[36] = r_5[35] /*5626*/;
  assign _1344_ = ~q[10] /*5625*/;
  assign _1345_ = sum_6[0] & q[10] /*5624*/;
  assign _1346_ = m_6[0] & _1344_ /*5623*/;
  assign r_6[0] = _1346_ | _1345_ /*5622*/;
  assign _1347_ = ~q[10] /*5621*/;
  assign _1348_ = sum_6[1] & q[10] /*5620*/;
  assign _1349_ = m_6[1] & _1347_ /*5619*/;
  assign r_6[1] = _1349_ | _1348_ /*5618*/;
  assign _1350_ = ~q[10] /*5617*/;
  assign _1351_ = sum_6[2] & q[10] /*5616*/;
  assign _1352_ = m_6[2] & _1350_ /*5615*/;
  assign r_6[2] = _1352_ | _1351_ /*5614*/;
  assign _1353_ = ~q[10] /*5613*/;
  assign _1354_ = sum_6[3] & q[10] /*5612*/;
  assign _1355_ = m_6[3] & _1353_ /*5611*/;
  assign r_6[3] = _1355_ | _1354_ /*5610*/;
  assign _1356_ = ~q[10] /*5609*/;
  assign _1357_ = sum_6[4] & q[10] /*5608*/;
  assign _1358_ = m_6[4] & _1356_ /*5607*/;
  assign r_6[4] = _1358_ | _1357_ /*5606*/;
  assign _1359_ = ~q[10] /*5605*/;
  assign _1360_ = sum_6[5] & q[10] /*5604*/;
  assign _1361_ = m_6[5] & _1359_ /*5603*/;
  assign r_6[5] = _1361_ | _1360_ /*5602*/;
  assign _1362_ = ~q[10] /*5601*/;
  assign _1363_ = sum_6[6] & q[10] /*5600*/;
  assign _1364_ = m_6[6] & _1362_ /*5599*/;
  assign r_6[6] = _1364_ | _1363_ /*5598*/;
  assign _1365_ = ~q[10] /*5597*/;
  assign _1366_ = sum_6[7] & q[10] /*5596*/;
  assign _1367_ = m_6[7] & _1365_ /*5595*/;
  assign r_6[7] = _1367_ | _1366_ /*5594*/;
  assign _1368_ = ~q[10] /*5593*/;
  assign _1369_ = sum_6[8] & q[10] /*5592*/;
  assign _1370_ = m_6[8] & _1368_ /*5591*/;
  assign r_6[8] = _1370_ | _1369_ /*5590*/;
  assign _1371_ = ~q[10] /*5589*/;
  assign _1372_ = sum_6[9] & q[10] /*5588*/;
  assign _1373_ = m_6[9] & _1371_ /*5587*/;
  assign r_6[9] = _1373_ | _1372_ /*5586*/;
  assign _1374_ = ~q[10] /*5585*/;
  assign _1375_ = sum_6[10] & q[10] /*5584*/;
  assign _1376_ = m_6[10] & _1374_ /*5583*/;
  assign r_6[10] = _1376_ | _1375_ /*5582*/;
  assign _1377_ = ~q[10] /*5581*/;
  assign _1378_ = sum_6[11] & q[10] /*5580*/;
  assign _1379_ = m_6[11] & _1377_ /*5579*/;
  assign r_6[11] = _1379_ | _1378_ /*5578*/;
  assign _1380_ = ~q[10] /*5577*/;
  assign _1381_ = sum_6[12] & q[10] /*5576*/;
  assign _1382_ = m_6[12] & _1380_ /*5575*/;
  assign r_6[12] = _1382_ | _1381_ /*5574*/;
  assign _1383_ = ~q[10] /*5573*/;
  assign _1384_ = sum_6[13] & q[10] /*5572*/;
  assign _1385_ = m_6[13] & _1383_ /*5571*/;
  assign r_6[13] = _1385_ | _1384_ /*5570*/;
  assign _1386_ = ~q[10] /*5569*/;
  assign _1387_ = sum_6[14] & q[10] /*5568*/;
  assign _1388_ = m_6[14] & _1386_ /*5567*/;
  assign r_6[14] = _1388_ | _1387_ /*5566*/;
  assign _1389_ = ~q[10] /*5565*/;
  assign _1390_ = sum_6[15] & q[10] /*5564*/;
  assign _1391_ = m_6[15] & _1389_ /*5563*/;
  assign r_6[15] = _1391_ | _1390_ /*5562*/;
  assign _1392_ = ~q[10] /*5561*/;
  assign _1393_ = sum_6[16] & q[10] /*5560*/;
  assign _1394_ = m_6[16] & _1392_ /*5559*/;
  assign r_6[16] = _1394_ | _1393_ /*5558*/;
  assign _1395_ = ~q[10] /*5557*/;
  assign _1396_ = sum_6[17] & q[10] /*5556*/;
  assign _1397_ = m_6[17] & _1395_ /*5555*/;
  assign r_6[17] = _1397_ | _1396_ /*5554*/;
  assign _1398_ = ~q[10] /*5553*/;
  assign _1399_ = sum_6[18] & q[10] /*5552*/;
  assign _1400_ = m_6[18] & _1398_ /*5551*/;
  assign r_6[18] = _1400_ | _1399_ /*5550*/;
  assign _1401_ = ~q[10] /*5549*/;
  assign _1402_ = sum_6[19] & q[10] /*5548*/;
  assign _1403_ = m_6[19] & _1401_ /*5547*/;
  assign r_6[19] = _1403_ | _1402_ /*5546*/;
  assign _1404_ = ~q[10] /*5545*/;
  assign _1405_ = sum_6[20] & q[10] /*5544*/;
  assign _1406_ = m_6[20] & _1404_ /*5543*/;
  assign r_6[20] = _1406_ | _1405_ /*5542*/;
  assign _1407_ = ~q[10] /*5541*/;
  assign _1408_ = sum_6[21] & q[10] /*5540*/;
  assign _1409_ = m_6[21] & _1407_ /*5539*/;
  assign r_6[21] = _1409_ | _1408_ /*5538*/;
  assign _1410_ = ~q[10] /*5537*/;
  assign _1411_ = sum_6[22] & q[10] /*5536*/;
  assign _1412_ = m_6[22] & _1410_ /*5535*/;
  assign r_6[22] = _1412_ | _1411_ /*5534*/;
  assign _1413_ = ~q[10] /*5533*/;
  assign _1414_ = sum_6[23] & q[10] /*5532*/;
  assign _1415_ = m_6[23] & _1413_ /*5531*/;
  assign r_6[23] = _1415_ | _1414_ /*5530*/;
  assign _1416_ = ~q[10] /*5529*/;
  assign _1417_ = sum_6[24] & q[10] /*5528*/;
  assign _1418_ = m_6[24] & _1416_ /*5527*/;
  assign r_6[24] = _1418_ | _1417_ /*5526*/;
  assign _1419_ = ~q[10] /*5525*/;
  assign _1420_ = sum_6[25] & q[10] /*5524*/;
  assign _1421_ = m_6[25] & _1419_ /*5523*/;
  assign r_6[25] = _1421_ | _1420_ /*5522*/;
  assign _1422_ = ~q[10] /*5521*/;
  assign _1423_ = sum_6[26] & q[10] /*5520*/;
  assign _1424_ = m_6[26] & _1422_ /*5519*/;
  assign r_6[26] = _1424_ | _1423_ /*5518*/;
  assign _1425_ = ~q[10] /*5517*/;
  assign _1426_ = sum_6[27] & q[10] /*5516*/;
  assign _1427_ = m_6[27] & _1425_ /*5515*/;
  assign r_6[27] = _1427_ | _1426_ /*5514*/;
  assign _1428_ = ~q[10] /*5513*/;
  assign _1429_ = sum_6[28] & q[10] /*5512*/;
  assign _1430_ = m_6[28] & _1428_ /*5511*/;
  assign r_6[28] = _1430_ | _1429_ /*5510*/;
  assign _1431_ = ~q[10] /*5509*/;
  assign _1432_ = sum_6[29] & q[10] /*5508*/;
  assign _1433_ = m_6[29] & _1431_ /*5507*/;
  assign r_6[29] = _1433_ | _1432_ /*5506*/;
  assign _1434_ = ~q[10] /*5505*/;
  assign _1435_ = sum_6[30] & q[10] /*5504*/;
  assign _1436_ = m_6[30] & _1434_ /*5503*/;
  assign r_6[30] = _1436_ | _1435_ /*5502*/;
  assign _1437_ = ~q[10] /*5501*/;
  assign _1438_ = sum_6[31] & q[10] /*5500*/;
  assign _1439_ = m_6[31] & _1437_ /*5499*/;
  assign r_6[31] = _1439_ | _1438_ /*5498*/;
  assign _1440_ = ~q[10] /*5497*/;
  assign _1441_ = sum_6[32] & q[10] /*5496*/;
  assign _1442_ = m_6[32] & _1440_ /*5495*/;
  assign r_6[32] = _1442_ | _1441_ /*5494*/;
  assign _1443_ = ~q[10] /*5493*/;
  assign _1444_ = sum_6[33] & q[10] /*5492*/;
  assign _1445_ = m_6[33] & _1443_ /*5491*/;
  assign r_6[33] = _1445_ | _1444_ /*5490*/;
  assign _1446_ = ~q[10] /*5489*/;
  assign _1447_ = sum_6[34] & q[10] /*5488*/;
  assign _1448_ = m_6[34] & _1446_ /*5487*/;
  assign r_6[34] = _1448_ | _1447_ /*5486*/;
  assign _1449_ = ~q[10] /*5485*/;
  assign _1450_ = sum_6[35] & q[10] /*5484*/;
  assign _1451_ = m_6[35] & _1449_ /*5483*/;
  assign r_6[35] = _1451_ | _1450_ /*5482*/;
  assign _1452_ = ~q[10] /*5481*/;
  assign _1453_ = sum_6[36] & q[10] /*5480*/;
  assign _1454_ = m_6[36] & _1452_ /*5479*/;
  assign r_6[36] = _1454_ | _1453_ /*5478*/;
  assign inv_7[0] = oneWire /*5352*/;
  assign inv_7[1] = oneWire /*5346*/;
  assign inv_7[2] = oneWire /*5340*/;
  assign inv_7[3] = oneWire /*5334*/;
  assign inv_7[4] = oneWire /*5328*/;
  assign inv_7[5] = oneWire /*5322*/;
  assign inv_7[6] = oneWire /*5316*/;
  assign inv_7[7] = oneWire /*5310*/;
  assign inv_7[8] = oneWire /*5304*/;
  assign inv_7[9] = ~div[0] /*5298*/;
  assign inv_7[10] = ~div[1] /*5292*/;
  assign inv_7[11] = ~div[2] /*5286*/;
  assign inv_7[12] = ~div[3] /*5280*/;
  assign inv_7[13] = ~div[4] /*5274*/;
  assign inv_7[14] = ~div[5] /*5268*/;
  assign inv_7[15] = ~div[6] /*5262*/;
  assign inv_7[16] = ~div[7] /*5256*/;
  assign inv_7[17] = ~div[8] /*5250*/;
  assign inv_7[18] = ~div[9] /*5244*/;
  assign inv_7[19] = ~div[10] /*5238*/;
  assign inv_7[20] = ~div[11] /*5232*/;
  assign inv_7[21] = ~div[12] /*5226*/;
  assign inv_7[22] = ~div[13] /*5220*/;
  assign inv_7[23] = ~div[14] /*5214*/;
  assign inv_7[24] = oneWire /*5208*/;
  assign inv_7[25] = oneWire /*5202*/;
  assign inv_7[26] = oneWire /*5196*/;
  assign inv_7[27] = oneWire /*5190*/;
  assign inv_7[28] = oneWire /*5184*/;
  assign inv_7[29] = oneWire /*5178*/;
  assign inv_7[30] = oneWire /*5172*/;
  assign inv_7[31] = oneWire /*5166*/;
  assign inv_7[32] = oneWire /*5160*/;
  assign inv_7[33] = oneWire /*5154*/;
  assign inv_7[34] = oneWire /*5148*/;
  assign inv_7[35] = oneWire /*5142*/;
  assign inv_7[36] = oneWire /*5136*/;
  assign _1455_ = inv_7[0] ^ r_6[0] /*5351*/;
  assign sum_7[0] = _1455_ ^ oneWire /*5350*/;
  assign _1456_ = _1455_ & oneWire /*5349*/;
  assign _1457_ = inv_7[0] & r_6[0] /*5348*/;
  assign _1458_ = _1456_ | _1457_ /*5347*/;
  assign _1459_ = inv_7[1] ^ r_6[1] /*5345*/;
  assign sum_7[1] = _1459_ ^ _1458_ /*5344*/;
  assign _1460_ = _1459_ & _1458_ /*5343*/;
  assign _1461_ = inv_7[1] & r_6[1] /*5342*/;
  assign _1462_ = _1460_ | _1461_ /*5341*/;
  assign _1463_ = inv_7[2] ^ r_6[2] /*5339*/;
  assign sum_7[2] = _1463_ ^ _1462_ /*5338*/;
  assign _1464_ = _1463_ & _1462_ /*5337*/;
  assign _1465_ = inv_7[2] & r_6[2] /*5336*/;
  assign _1466_ = _1464_ | _1465_ /*5335*/;
  assign _1467_ = inv_7[3] ^ r_6[3] /*5333*/;
  assign sum_7[3] = _1467_ ^ _1466_ /*5332*/;
  assign _1468_ = _1467_ & _1466_ /*5331*/;
  assign _1469_ = inv_7[3] & r_6[3] /*5330*/;
  assign _1470_ = _1468_ | _1469_ /*5329*/;
  assign _1471_ = inv_7[4] ^ r_6[4] /*5327*/;
  assign sum_7[4] = _1471_ ^ _1470_ /*5326*/;
  assign _1472_ = _1471_ & _1470_ /*5325*/;
  assign _1473_ = inv_7[4] & r_6[4] /*5324*/;
  assign _1474_ = _1472_ | _1473_ /*5323*/;
  assign _1475_ = inv_7[5] ^ r_6[5] /*5321*/;
  assign sum_7[5] = _1475_ ^ _1474_ /*5320*/;
  assign _1476_ = _1475_ & _1474_ /*5319*/;
  assign _1477_ = inv_7[5] & r_6[5] /*5318*/;
  assign _1478_ = _1476_ | _1477_ /*5317*/;
  assign _1479_ = inv_7[6] ^ r_6[6] /*5315*/;
  assign sum_7[6] = _1479_ ^ _1478_ /*5314*/;
  assign _1480_ = _1479_ & _1478_ /*5313*/;
  assign _1481_ = inv_7[6] & r_6[6] /*5312*/;
  assign _1482_ = _1480_ | _1481_ /*5311*/;
  assign _1483_ = inv_7[7] ^ r_6[7] /*5309*/;
  assign sum_7[7] = _1483_ ^ _1482_ /*5308*/;
  assign _1484_ = _1483_ & _1482_ /*5307*/;
  assign _1485_ = inv_7[7] & r_6[7] /*5306*/;
  assign _1486_ = _1484_ | _1485_ /*5305*/;
  assign _1487_ = inv_7[8] ^ r_6[8] /*5303*/;
  assign sum_7[8] = _1487_ ^ _1486_ /*5302*/;
  assign _1488_ = _1487_ & _1486_ /*5301*/;
  assign _1489_ = inv_7[8] & r_6[8] /*5300*/;
  assign _1490_ = _1488_ | _1489_ /*5299*/;
  assign _1491_ = inv_7[9] ^ r_6[9] /*5297*/;
  assign sum_7[9] = _1491_ ^ _1490_ /*5296*/;
  assign _1492_ = _1491_ & _1490_ /*5295*/;
  assign _1493_ = inv_7[9] & r_6[9] /*5294*/;
  assign _1494_ = _1492_ | _1493_ /*5293*/;
  assign _1495_ = inv_7[10] ^ r_6[10] /*5291*/;
  assign sum_7[10] = _1495_ ^ _1494_ /*5290*/;
  assign _1496_ = _1495_ & _1494_ /*5289*/;
  assign _1497_ = inv_7[10] & r_6[10] /*5288*/;
  assign _1498_ = _1496_ | _1497_ /*5287*/;
  assign _1499_ = inv_7[11] ^ r_6[11] /*5285*/;
  assign sum_7[11] = _1499_ ^ _1498_ /*5284*/;
  assign _1500_ = _1499_ & _1498_ /*5283*/;
  assign _1501_ = inv_7[11] & r_6[11] /*5282*/;
  assign _1502_ = _1500_ | _1501_ /*5281*/;
  assign _1503_ = inv_7[12] ^ r_6[12] /*5279*/;
  assign sum_7[12] = _1503_ ^ _1502_ /*5278*/;
  assign _1504_ = _1503_ & _1502_ /*5277*/;
  assign _1505_ = inv_7[12] & r_6[12] /*5276*/;
  assign _1506_ = _1504_ | _1505_ /*5275*/;
  assign _1507_ = inv_7[13] ^ r_6[13] /*5273*/;
  assign sum_7[13] = _1507_ ^ _1506_ /*5272*/;
  assign _1508_ = _1507_ & _1506_ /*5271*/;
  assign _1509_ = inv_7[13] & r_6[13] /*5270*/;
  assign _1510_ = _1508_ | _1509_ /*5269*/;
  assign _1511_ = inv_7[14] ^ r_6[14] /*5267*/;
  assign sum_7[14] = _1511_ ^ _1510_ /*5266*/;
  assign _1512_ = _1511_ & _1510_ /*5265*/;
  assign _1513_ = inv_7[14] & r_6[14] /*5264*/;
  assign _1514_ = _1512_ | _1513_ /*5263*/;
  assign _1515_ = inv_7[15] ^ r_6[15] /*5261*/;
  assign sum_7[15] = _1515_ ^ _1514_ /*5260*/;
  assign _1516_ = _1515_ & _1514_ /*5259*/;
  assign _1517_ = inv_7[15] & r_6[15] /*5258*/;
  assign _1518_ = _1516_ | _1517_ /*5257*/;
  assign _1519_ = inv_7[16] ^ r_6[16] /*5255*/;
  assign sum_7[16] = _1519_ ^ _1518_ /*5254*/;
  assign _1520_ = _1519_ & _1518_ /*5253*/;
  assign _1521_ = inv_7[16] & r_6[16] /*5252*/;
  assign _1522_ = _1520_ | _1521_ /*5251*/;
  assign _1523_ = inv_7[17] ^ r_6[17] /*5249*/;
  assign sum_7[17] = _1523_ ^ _1522_ /*5248*/;
  assign _1524_ = _1523_ & _1522_ /*5247*/;
  assign _1525_ = inv_7[17] & r_6[17] /*5246*/;
  assign _1526_ = _1524_ | _1525_ /*5245*/;
  assign _1527_ = inv_7[18] ^ r_6[18] /*5243*/;
  assign sum_7[18] = _1527_ ^ _1526_ /*5242*/;
  assign _1528_ = _1527_ & _1526_ /*5241*/;
  assign _1529_ = inv_7[18] & r_6[18] /*5240*/;
  assign _1530_ = _1528_ | _1529_ /*5239*/;
  assign _1531_ = inv_7[19] ^ r_6[19] /*5237*/;
  assign sum_7[19] = _1531_ ^ _1530_ /*5236*/;
  assign _1532_ = _1531_ & _1530_ /*5235*/;
  assign _1533_ = inv_7[19] & r_6[19] /*5234*/;
  assign _1534_ = _1532_ | _1533_ /*5233*/;
  assign _1535_ = inv_7[20] ^ r_6[20] /*5231*/;
  assign sum_7[20] = _1535_ ^ _1534_ /*5230*/;
  assign _1536_ = _1535_ & _1534_ /*5229*/;
  assign _1537_ = inv_7[20] & r_6[20] /*5228*/;
  assign _1538_ = _1536_ | _1537_ /*5227*/;
  assign _1539_ = inv_7[21] ^ r_6[21] /*5225*/;
  assign sum_7[21] = _1539_ ^ _1538_ /*5224*/;
  assign _1540_ = _1539_ & _1538_ /*5223*/;
  assign _1541_ = inv_7[21] & r_6[21] /*5222*/;
  assign _1542_ = _1540_ | _1541_ /*5221*/;
  assign _1543_ = inv_7[22] ^ r_6[22] /*5219*/;
  assign sum_7[22] = _1543_ ^ _1542_ /*5218*/;
  assign _1544_ = _1543_ & _1542_ /*5217*/;
  assign _1545_ = inv_7[22] & r_6[22] /*5216*/;
  assign _1546_ = _1544_ | _1545_ /*5215*/;
  assign _1547_ = inv_7[23] ^ r_6[23] /*5213*/;
  assign sum_7[23] = _1547_ ^ _1546_ /*5212*/;
  assign _1548_ = _1547_ & _1546_ /*5211*/;
  assign _1549_ = inv_7[23] & r_6[23] /*5210*/;
  assign _1550_ = _1548_ | _1549_ /*5209*/;
  assign _1551_ = inv_7[24] ^ r_6[24] /*5207*/;
  assign sum_7[24] = _1551_ ^ _1550_ /*5206*/;
  assign _1552_ = _1551_ & _1550_ /*5205*/;
  assign _1553_ = inv_7[24] & r_6[24] /*5204*/;
  assign _1554_ = _1552_ | _1553_ /*5203*/;
  assign _1555_ = inv_7[25] ^ r_6[25] /*5201*/;
  assign sum_7[25] = _1555_ ^ _1554_ /*5200*/;
  assign _1556_ = _1555_ & _1554_ /*5199*/;
  assign _1557_ = inv_7[25] & r_6[25] /*5198*/;
  assign _1558_ = _1556_ | _1557_ /*5197*/;
  assign _1559_ = inv_7[26] ^ r_6[26] /*5195*/;
  assign sum_7[26] = _1559_ ^ _1558_ /*5194*/;
  assign _1560_ = _1559_ & _1558_ /*5193*/;
  assign _1561_ = inv_7[26] & r_6[26] /*5192*/;
  assign _1562_ = _1560_ | _1561_ /*5191*/;
  assign _1563_ = inv_7[27] ^ r_6[27] /*5189*/;
  assign sum_7[27] = _1563_ ^ _1562_ /*5188*/;
  assign _1564_ = _1563_ & _1562_ /*5187*/;
  assign _1565_ = inv_7[27] & r_6[27] /*5186*/;
  assign _1566_ = _1564_ | _1565_ /*5185*/;
  assign _1567_ = inv_7[28] ^ r_6[28] /*5183*/;
  assign sum_7[28] = _1567_ ^ _1566_ /*5182*/;
  assign _1568_ = _1567_ & _1566_ /*5181*/;
  assign _1569_ = inv_7[28] & r_6[28] /*5180*/;
  assign _1570_ = _1568_ | _1569_ /*5179*/;
  assign _1571_ = inv_7[29] ^ r_6[29] /*5177*/;
  assign sum_7[29] = _1571_ ^ _1570_ /*5176*/;
  assign _1572_ = _1571_ & _1570_ /*5175*/;
  assign _1573_ = inv_7[29] & r_6[29] /*5174*/;
  assign _1574_ = _1572_ | _1573_ /*5173*/;
  assign _1575_ = inv_7[30] ^ r_6[30] /*5171*/;
  assign sum_7[30] = _1575_ ^ _1574_ /*5170*/;
  assign _1576_ = _1575_ & _1574_ /*5169*/;
  assign _1577_ = inv_7[30] & r_6[30] /*5168*/;
  assign _1578_ = _1576_ | _1577_ /*5167*/;
  assign _1579_ = inv_7[31] ^ r_6[31] /*5165*/;
  assign sum_7[31] = _1579_ ^ _1578_ /*5164*/;
  assign _1580_ = _1579_ & _1578_ /*5163*/;
  assign _1581_ = inv_7[31] & r_6[31] /*5162*/;
  assign _1582_ = _1580_ | _1581_ /*5161*/;
  assign _1583_ = inv_7[32] ^ r_6[32] /*5159*/;
  assign sum_7[32] = _1583_ ^ _1582_ /*5158*/;
  assign _1584_ = _1583_ & _1582_ /*5157*/;
  assign _1585_ = inv_7[32] & r_6[32] /*5156*/;
  assign _1586_ = _1584_ | _1585_ /*5155*/;
  assign _1587_ = inv_7[33] ^ r_6[33] /*5153*/;
  assign sum_7[33] = _1587_ ^ _1586_ /*5152*/;
  assign _1588_ = _1587_ & _1586_ /*5151*/;
  assign _1589_ = inv_7[33] & r_6[33] /*5150*/;
  assign _1590_ = _1588_ | _1589_ /*5149*/;
  assign _1591_ = inv_7[34] ^ r_6[34] /*5147*/;
  assign sum_7[34] = _1591_ ^ _1590_ /*5146*/;
  assign _1592_ = _1591_ & _1590_ /*5145*/;
  assign _1593_ = inv_7[34] & r_6[34] /*5144*/;
  assign _1594_ = _1592_ | _1593_ /*5143*/;
  assign _1595_ = inv_7[35] ^ r_6[35] /*5141*/;
  assign sum_7[35] = _1595_ ^ _1594_ /*5140*/;
  assign _1596_ = _1595_ & _1594_ /*5139*/;
  assign _1597_ = inv_7[35] & r_6[35] /*5138*/;
  assign _1598_ = _1596_ | _1597_ /*5137*/;
  assign _1599_ = inv_7[36] ^ r_6[36] /*5135*/;
  assign sum_7[36] = _1599_ ^ _1598_ /*5134*/;
  assign _1600_ = _1599_ & _1598_ /*5133*/;
  assign _1601_ = inv_7[36] & r_6[36] /*5132*/;
  assign _1602_ = _1600_ | _1601_ /*5131*/;
  assign _1603_ = _1602_ ^ _1598_ /*5130*/;
  assign _1604_ = ~_1603_ /*5129*/;
  assign _1605_ = sum_7[36] & _1604_ /*5128*/;
  assign _1606_ = _1603_ & _1602_ /*5127*/;
  assign sum_7[37] = _1606_ | _1605_ /*5126*/;
  assign q[9] = ~sum_7[37] /*5125*/;
  assign m_7[0] = r_6[0] /*5124*/;
  assign m_7[1] = r_6[1] /*5123*/;
  assign m_7[2] = r_6[2] /*5122*/;
  assign m_7[3] = r_6[3] /*5121*/;
  assign m_7[4] = r_6[4] /*5120*/;
  assign m_7[5] = r_6[5] /*5119*/;
  assign m_7[6] = r_6[6] /*5118*/;
  assign m_7[7] = r_6[7] /*5117*/;
  assign m_7[8] = r_6[8] /*5116*/;
  assign m_7[9] = r_6[9] /*5115*/;
  assign m_7[10] = r_6[10] /*5114*/;
  assign m_7[11] = r_6[11] /*5113*/;
  assign m_7[12] = r_6[12] /*5112*/;
  assign m_7[13] = r_6[13] /*5111*/;
  assign m_7[14] = r_6[14] /*5110*/;
  assign m_7[15] = r_6[15] /*5109*/;
  assign m_7[16] = r_6[16] /*5108*/;
  assign m_7[17] = r_6[17] /*5107*/;
  assign m_7[18] = r_6[18] /*5106*/;
  assign m_7[19] = r_6[19] /*5105*/;
  assign m_7[20] = r_6[20] /*5104*/;
  assign m_7[21] = r_6[21] /*5103*/;
  assign m_7[22] = r_6[22] /*5102*/;
  assign m_7[23] = r_6[23] /*5101*/;
  assign m_7[24] = r_6[24] /*5100*/;
  assign m_7[25] = r_6[25] /*5099*/;
  assign m_7[26] = r_6[26] /*5098*/;
  assign m_7[27] = r_6[27] /*5097*/;
  assign m_7[28] = r_6[28] /*5096*/;
  assign m_7[29] = r_6[29] /*5095*/;
  assign m_7[30] = r_6[30] /*5094*/;
  assign m_7[31] = r_6[31] /*5093*/;
  assign m_7[32] = r_6[32] /*5092*/;
  assign m_7[33] = r_6[33] /*5091*/;
  assign m_7[34] = r_6[34] /*5090*/;
  assign m_7[35] = r_6[35] /*5089*/;
  assign m_7[36] = r_6[36] /*5088*/;
  assign m_7[37] = r_6[36] /*5087*/;
  assign _1608_ = ~q[9] /*5086*/;
  assign _1609_ = sum_7[0] & q[9] /*5085*/;
  assign _1610_ = m_7[0] & _1608_ /*5084*/;
  assign r_7[0] = _1610_ | _1609_ /*5083*/;
  assign _1611_ = ~q[9] /*5082*/;
  assign _1612_ = sum_7[1] & q[9] /*5081*/;
  assign _1613_ = m_7[1] & _1611_ /*5080*/;
  assign r_7[1] = _1613_ | _1612_ /*5079*/;
  assign _1614_ = ~q[9] /*5078*/;
  assign _1615_ = sum_7[2] & q[9] /*5077*/;
  assign _1616_ = m_7[2] & _1614_ /*5076*/;
  assign r_7[2] = _1616_ | _1615_ /*5075*/;
  assign _1617_ = ~q[9] /*5074*/;
  assign _1618_ = sum_7[3] & q[9] /*5073*/;
  assign _1619_ = m_7[3] & _1617_ /*5072*/;
  assign r_7[3] = _1619_ | _1618_ /*5071*/;
  assign _1620_ = ~q[9] /*5070*/;
  assign _1621_ = sum_7[4] & q[9] /*5069*/;
  assign _1622_ = m_7[4] & _1620_ /*5068*/;
  assign r_7[4] = _1622_ | _1621_ /*5067*/;
  assign _1623_ = ~q[9] /*5066*/;
  assign _1624_ = sum_7[5] & q[9] /*5065*/;
  assign _1625_ = m_7[5] & _1623_ /*5064*/;
  assign r_7[5] = _1625_ | _1624_ /*5063*/;
  assign _1626_ = ~q[9] /*5062*/;
  assign _1627_ = sum_7[6] & q[9] /*5061*/;
  assign _1628_ = m_7[6] & _1626_ /*5060*/;
  assign r_7[6] = _1628_ | _1627_ /*5059*/;
  assign _1629_ = ~q[9] /*5058*/;
  assign _1630_ = sum_7[7] & q[9] /*5057*/;
  assign _1631_ = m_7[7] & _1629_ /*5056*/;
  assign r_7[7] = _1631_ | _1630_ /*5055*/;
  assign _1632_ = ~q[9] /*5054*/;
  assign _1633_ = sum_7[8] & q[9] /*5053*/;
  assign _1634_ = m_7[8] & _1632_ /*5052*/;
  assign r_7[8] = _1634_ | _1633_ /*5051*/;
  assign _1635_ = ~q[9] /*5050*/;
  assign _1636_ = sum_7[9] & q[9] /*5049*/;
  assign _1637_ = m_7[9] & _1635_ /*5048*/;
  assign r_7[9] = _1637_ | _1636_ /*5047*/;
  assign _1638_ = ~q[9] /*5046*/;
  assign _1639_ = sum_7[10] & q[9] /*5045*/;
  assign _1640_ = m_7[10] & _1638_ /*5044*/;
  assign r_7[10] = _1640_ | _1639_ /*5043*/;
  assign _1641_ = ~q[9] /*5042*/;
  assign _1642_ = sum_7[11] & q[9] /*5041*/;
  assign _1643_ = m_7[11] & _1641_ /*5040*/;
  assign r_7[11] = _1643_ | _1642_ /*5039*/;
  assign _1644_ = ~q[9] /*5038*/;
  assign _1645_ = sum_7[12] & q[9] /*5037*/;
  assign _1646_ = m_7[12] & _1644_ /*5036*/;
  assign r_7[12] = _1646_ | _1645_ /*5035*/;
  assign _1647_ = ~q[9] /*5034*/;
  assign _1648_ = sum_7[13] & q[9] /*5033*/;
  assign _1649_ = m_7[13] & _1647_ /*5032*/;
  assign r_7[13] = _1649_ | _1648_ /*5031*/;
  assign _1650_ = ~q[9] /*5030*/;
  assign _1651_ = sum_7[14] & q[9] /*5029*/;
  assign _1652_ = m_7[14] & _1650_ /*5028*/;
  assign r_7[14] = _1652_ | _1651_ /*5027*/;
  assign _1653_ = ~q[9] /*5026*/;
  assign _1654_ = sum_7[15] & q[9] /*5025*/;
  assign _1655_ = m_7[15] & _1653_ /*5024*/;
  assign r_7[15] = _1655_ | _1654_ /*5023*/;
  assign _1656_ = ~q[9] /*5022*/;
  assign _1657_ = sum_7[16] & q[9] /*5021*/;
  assign _1658_ = m_7[16] & _1656_ /*5020*/;
  assign r_7[16] = _1658_ | _1657_ /*5019*/;
  assign _1659_ = ~q[9] /*5018*/;
  assign _1660_ = sum_7[17] & q[9] /*5017*/;
  assign _1661_ = m_7[17] & _1659_ /*5016*/;
  assign r_7[17] = _1661_ | _1660_ /*5015*/;
  assign _1662_ = ~q[9] /*5014*/;
  assign _1663_ = sum_7[18] & q[9] /*5013*/;
  assign _1664_ = m_7[18] & _1662_ /*5012*/;
  assign r_7[18] = _1664_ | _1663_ /*5011*/;
  assign _1665_ = ~q[9] /*5010*/;
  assign _1666_ = sum_7[19] & q[9] /*5009*/;
  assign _1667_ = m_7[19] & _1665_ /*5008*/;
  assign r_7[19] = _1667_ | _1666_ /*5007*/;
  assign _1668_ = ~q[9] /*5006*/;
  assign _1669_ = sum_7[20] & q[9] /*5005*/;
  assign _1670_ = m_7[20] & _1668_ /*5004*/;
  assign r_7[20] = _1670_ | _1669_ /*5003*/;
  assign _1671_ = ~q[9] /*5002*/;
  assign _1672_ = sum_7[21] & q[9] /*5001*/;
  assign _1673_ = m_7[21] & _1671_ /*5000*/;
  assign r_7[21] = _1673_ | _1672_ /*4999*/;
  assign _1674_ = ~q[9] /*4998*/;
  assign _1675_ = sum_7[22] & q[9] /*4997*/;
  assign _1676_ = m_7[22] & _1674_ /*4996*/;
  assign r_7[22] = _1676_ | _1675_ /*4995*/;
  assign _1677_ = ~q[9] /*4994*/;
  assign _1678_ = sum_7[23] & q[9] /*4993*/;
  assign _1679_ = m_7[23] & _1677_ /*4992*/;
  assign r_7[23] = _1679_ | _1678_ /*4991*/;
  assign _1680_ = ~q[9] /*4990*/;
  assign _1681_ = sum_7[24] & q[9] /*4989*/;
  assign _1682_ = m_7[24] & _1680_ /*4988*/;
  assign r_7[24] = _1682_ | _1681_ /*4987*/;
  assign _1683_ = ~q[9] /*4986*/;
  assign _1684_ = sum_7[25] & q[9] /*4985*/;
  assign _1685_ = m_7[25] & _1683_ /*4984*/;
  assign r_7[25] = _1685_ | _1684_ /*4983*/;
  assign _1686_ = ~q[9] /*4982*/;
  assign _1687_ = sum_7[26] & q[9] /*4981*/;
  assign _1688_ = m_7[26] & _1686_ /*4980*/;
  assign r_7[26] = _1688_ | _1687_ /*4979*/;
  assign _1689_ = ~q[9] /*4978*/;
  assign _1690_ = sum_7[27] & q[9] /*4977*/;
  assign _1691_ = m_7[27] & _1689_ /*4976*/;
  assign r_7[27] = _1691_ | _1690_ /*4975*/;
  assign _1692_ = ~q[9] /*4974*/;
  assign _1693_ = sum_7[28] & q[9] /*4973*/;
  assign _1694_ = m_7[28] & _1692_ /*4972*/;
  assign r_7[28] = _1694_ | _1693_ /*4971*/;
  assign _1695_ = ~q[9] /*4970*/;
  assign _1696_ = sum_7[29] & q[9] /*4969*/;
  assign _1697_ = m_7[29] & _1695_ /*4968*/;
  assign r_7[29] = _1697_ | _1696_ /*4967*/;
  assign _1698_ = ~q[9] /*4966*/;
  assign _1699_ = sum_7[30] & q[9] /*4965*/;
  assign _1700_ = m_7[30] & _1698_ /*4964*/;
  assign r_7[30] = _1700_ | _1699_ /*4963*/;
  assign _1701_ = ~q[9] /*4962*/;
  assign _1702_ = sum_7[31] & q[9] /*4961*/;
  assign _1703_ = m_7[31] & _1701_ /*4960*/;
  assign r_7[31] = _1703_ | _1702_ /*4959*/;
  assign _1704_ = ~q[9] /*4958*/;
  assign _1705_ = sum_7[32] & q[9] /*4957*/;
  assign _1706_ = m_7[32] & _1704_ /*4956*/;
  assign r_7[32] = _1706_ | _1705_ /*4955*/;
  assign _1707_ = ~q[9] /*4954*/;
  assign _1708_ = sum_7[33] & q[9] /*4953*/;
  assign _1709_ = m_7[33] & _1707_ /*4952*/;
  assign r_7[33] = _1709_ | _1708_ /*4951*/;
  assign _1710_ = ~q[9] /*4950*/;
  assign _1711_ = sum_7[34] & q[9] /*4949*/;
  assign _1712_ = m_7[34] & _1710_ /*4948*/;
  assign r_7[34] = _1712_ | _1711_ /*4947*/;
  assign _1713_ = ~q[9] /*4946*/;
  assign _1714_ = sum_7[35] & q[9] /*4945*/;
  assign _1715_ = m_7[35] & _1713_ /*4944*/;
  assign r_7[35] = _1715_ | _1714_ /*4943*/;
  assign _1716_ = ~q[9] /*4942*/;
  assign _1717_ = sum_7[36] & q[9] /*4941*/;
  assign _1718_ = m_7[36] & _1716_ /*4940*/;
  assign r_7[36] = _1718_ | _1717_ /*4939*/;
  assign _1719_ = ~q[9] /*4938*/;
  assign _1720_ = sum_7[37] & q[9] /*4937*/;
  assign _1721_ = m_7[37] & _1719_ /*4936*/;
  assign r_7[37] = _1721_ | _1720_ /*4935*/;
  assign inv_8[0] = oneWire /*4820*/;
  assign inv_8[1] = oneWire /*4814*/;
  assign inv_8[2] = oneWire /*4808*/;
  assign inv_8[3] = oneWire /*4802*/;
  assign inv_8[4] = oneWire /*4796*/;
  assign inv_8[5] = oneWire /*4790*/;
  assign inv_8[6] = oneWire /*4784*/;
  assign inv_8[7] = oneWire /*4778*/;
  assign inv_8[8] = ~div[0] /*4772*/;
  assign inv_8[9] = ~div[1] /*4766*/;
  assign inv_8[10] = ~div[2] /*4760*/;
  assign inv_8[11] = ~div[3] /*4754*/;
  assign inv_8[12] = ~div[4] /*4748*/;
  assign inv_8[13] = ~div[5] /*4742*/;
  assign inv_8[14] = ~div[6] /*4736*/;
  assign inv_8[15] = ~div[7] /*4730*/;
  assign inv_8[16] = ~div[8] /*4724*/;
  assign inv_8[17] = ~div[9] /*4718*/;
  assign inv_8[18] = ~div[10] /*4712*/;
  assign inv_8[19] = ~div[11] /*4706*/;
  assign inv_8[20] = ~div[12] /*4700*/;
  assign inv_8[21] = ~div[13] /*4694*/;
  assign inv_8[22] = ~div[14] /*4688*/;
  assign inv_8[23] = oneWire /*4682*/;
  assign inv_8[24] = oneWire /*4676*/;
  assign inv_8[25] = oneWire /*4670*/;
  assign inv_8[26] = oneWire /*4664*/;
  assign inv_8[27] = oneWire /*4658*/;
  assign inv_8[28] = oneWire /*4652*/;
  assign inv_8[29] = oneWire /*4646*/;
  assign inv_8[30] = oneWire /*4640*/;
  assign inv_8[31] = oneWire /*4634*/;
  assign inv_8[32] = oneWire /*4628*/;
  assign inv_8[33] = oneWire /*4622*/;
  assign inv_8[34] = oneWire /*4616*/;
  assign inv_8[35] = oneWire /*4610*/;
  assign inv_8[36] = oneWire /*4604*/;
  assign inv_8[37] = oneWire /*4598*/;
  assign _1722_ = inv_8[0] ^ r_7[0] /*4819*/;
  assign sum_8[0] = _1722_ ^ oneWire /*4818*/;
  assign _1723_ = _1722_ & oneWire /*4817*/;
  assign _1724_ = inv_8[0] & r_7[0] /*4816*/;
  assign _1725_ = _1723_ | _1724_ /*4815*/;
  assign _1726_ = inv_8[1] ^ r_7[1] /*4813*/;
  assign sum_8[1] = _1726_ ^ _1725_ /*4812*/;
  assign _1727_ = _1726_ & _1725_ /*4811*/;
  assign _1728_ = inv_8[1] & r_7[1] /*4810*/;
  assign _1729_ = _1727_ | _1728_ /*4809*/;
  assign _1730_ = inv_8[2] ^ r_7[2] /*4807*/;
  assign sum_8[2] = _1730_ ^ _1729_ /*4806*/;
  assign _1731_ = _1730_ & _1729_ /*4805*/;
  assign _1732_ = inv_8[2] & r_7[2] /*4804*/;
  assign _1733_ = _1731_ | _1732_ /*4803*/;
  assign _1734_ = inv_8[3] ^ r_7[3] /*4801*/;
  assign sum_8[3] = _1734_ ^ _1733_ /*4800*/;
  assign _1735_ = _1734_ & _1733_ /*4799*/;
  assign _1736_ = inv_8[3] & r_7[3] /*4798*/;
  assign _1737_ = _1735_ | _1736_ /*4797*/;
  assign _1738_ = inv_8[4] ^ r_7[4] /*4795*/;
  assign sum_8[4] = _1738_ ^ _1737_ /*4794*/;
  assign _1739_ = _1738_ & _1737_ /*4793*/;
  assign _1740_ = inv_8[4] & r_7[4] /*4792*/;
  assign _1741_ = _1739_ | _1740_ /*4791*/;
  assign _1742_ = inv_8[5] ^ r_7[5] /*4789*/;
  assign sum_8[5] = _1742_ ^ _1741_ /*4788*/;
  assign _1743_ = _1742_ & _1741_ /*4787*/;
  assign _1744_ = inv_8[5] & r_7[5] /*4786*/;
  assign _1745_ = _1743_ | _1744_ /*4785*/;
  assign _1746_ = inv_8[6] ^ r_7[6] /*4783*/;
  assign sum_8[6] = _1746_ ^ _1745_ /*4782*/;
  assign _1747_ = _1746_ & _1745_ /*4781*/;
  assign _1748_ = inv_8[6] & r_7[6] /*4780*/;
  assign _1749_ = _1747_ | _1748_ /*4779*/;
  assign _1750_ = inv_8[7] ^ r_7[7] /*4777*/;
  assign sum_8[7] = _1750_ ^ _1749_ /*4776*/;
  assign _1751_ = _1750_ & _1749_ /*4775*/;
  assign _1752_ = inv_8[7] & r_7[7] /*4774*/;
  assign _1753_ = _1751_ | _1752_ /*4773*/;
  assign _1754_ = inv_8[8] ^ r_7[8] /*4771*/;
  assign sum_8[8] = _1754_ ^ _1753_ /*4770*/;
  assign _1755_ = _1754_ & _1753_ /*4769*/;
  assign _1756_ = inv_8[8] & r_7[8] /*4768*/;
  assign _1757_ = _1755_ | _1756_ /*4767*/;
  assign _1758_ = inv_8[9] ^ r_7[9] /*4765*/;
  assign sum_8[9] = _1758_ ^ _1757_ /*4764*/;
  assign _1759_ = _1758_ & _1757_ /*4763*/;
  assign _1760_ = inv_8[9] & r_7[9] /*4762*/;
  assign _1761_ = _1759_ | _1760_ /*4761*/;
  assign _1762_ = inv_8[10] ^ r_7[10] /*4759*/;
  assign sum_8[10] = _1762_ ^ _1761_ /*4758*/;
  assign _1763_ = _1762_ & _1761_ /*4757*/;
  assign _1764_ = inv_8[10] & r_7[10] /*4756*/;
  assign _1765_ = _1763_ | _1764_ /*4755*/;
  assign _1766_ = inv_8[11] ^ r_7[11] /*4753*/;
  assign sum_8[11] = _1766_ ^ _1765_ /*4752*/;
  assign _1767_ = _1766_ & _1765_ /*4751*/;
  assign _1768_ = inv_8[11] & r_7[11] /*4750*/;
  assign _1769_ = _1767_ | _1768_ /*4749*/;
  assign _1770_ = inv_8[12] ^ r_7[12] /*4747*/;
  assign sum_8[12] = _1770_ ^ _1769_ /*4746*/;
  assign _1771_ = _1770_ & _1769_ /*4745*/;
  assign _1772_ = inv_8[12] & r_7[12] /*4744*/;
  assign _1773_ = _1771_ | _1772_ /*4743*/;
  assign _1774_ = inv_8[13] ^ r_7[13] /*4741*/;
  assign sum_8[13] = _1774_ ^ _1773_ /*4740*/;
  assign _1775_ = _1774_ & _1773_ /*4739*/;
  assign _1776_ = inv_8[13] & r_7[13] /*4738*/;
  assign _1777_ = _1775_ | _1776_ /*4737*/;
  assign _1778_ = inv_8[14] ^ r_7[14] /*4735*/;
  assign sum_8[14] = _1778_ ^ _1777_ /*4734*/;
  assign _1779_ = _1778_ & _1777_ /*4733*/;
  assign _1780_ = inv_8[14] & r_7[14] /*4732*/;
  assign _1781_ = _1779_ | _1780_ /*4731*/;
  assign _1782_ = inv_8[15] ^ r_7[15] /*4729*/;
  assign sum_8[15] = _1782_ ^ _1781_ /*4728*/;
  assign _1783_ = _1782_ & _1781_ /*4727*/;
  assign _1784_ = inv_8[15] & r_7[15] /*4726*/;
  assign _1785_ = _1783_ | _1784_ /*4725*/;
  assign _1786_ = inv_8[16] ^ r_7[16] /*4723*/;
  assign sum_8[16] = _1786_ ^ _1785_ /*4722*/;
  assign _1787_ = _1786_ & _1785_ /*4721*/;
  assign _1788_ = inv_8[16] & r_7[16] /*4720*/;
  assign _1789_ = _1787_ | _1788_ /*4719*/;
  assign _1790_ = inv_8[17] ^ r_7[17] /*4717*/;
  assign sum_8[17] = _1790_ ^ _1789_ /*4716*/;
  assign _1791_ = _1790_ & _1789_ /*4715*/;
  assign _1792_ = inv_8[17] & r_7[17] /*4714*/;
  assign _1793_ = _1791_ | _1792_ /*4713*/;
  assign _1794_ = inv_8[18] ^ r_7[18] /*4711*/;
  assign sum_8[18] = _1794_ ^ _1793_ /*4710*/;
  assign _1795_ = _1794_ & _1793_ /*4709*/;
  assign _1796_ = inv_8[18] & r_7[18] /*4708*/;
  assign _1797_ = _1795_ | _1796_ /*4707*/;
  assign _1798_ = inv_8[19] ^ r_7[19] /*4705*/;
  assign sum_8[19] = _1798_ ^ _1797_ /*4704*/;
  assign _1799_ = _1798_ & _1797_ /*4703*/;
  assign _1800_ = inv_8[19] & r_7[19] /*4702*/;
  assign _1801_ = _1799_ | _1800_ /*4701*/;
  assign _1802_ = inv_8[20] ^ r_7[20] /*4699*/;
  assign sum_8[20] = _1802_ ^ _1801_ /*4698*/;
  assign _1803_ = _1802_ & _1801_ /*4697*/;
  assign _1804_ = inv_8[20] & r_7[20] /*4696*/;
  assign _1805_ = _1803_ | _1804_ /*4695*/;
  assign _1806_ = inv_8[21] ^ r_7[21] /*4693*/;
  assign sum_8[21] = _1806_ ^ _1805_ /*4692*/;
  assign _1807_ = _1806_ & _1805_ /*4691*/;
  assign _1808_ = inv_8[21] & r_7[21] /*4690*/;
  assign _1809_ = _1807_ | _1808_ /*4689*/;
  assign _1810_ = inv_8[22] ^ r_7[22] /*4687*/;
  assign sum_8[22] = _1810_ ^ _1809_ /*4686*/;
  assign _1811_ = _1810_ & _1809_ /*4685*/;
  assign _1812_ = inv_8[22] & r_7[22] /*4684*/;
  assign _1813_ = _1811_ | _1812_ /*4683*/;
  assign _1814_ = inv_8[23] ^ r_7[23] /*4681*/;
  assign sum_8[23] = _1814_ ^ _1813_ /*4680*/;
  assign _1815_ = _1814_ & _1813_ /*4679*/;
  assign _1816_ = inv_8[23] & r_7[23] /*4678*/;
  assign _1817_ = _1815_ | _1816_ /*4677*/;
  assign _1818_ = inv_8[24] ^ r_7[24] /*4675*/;
  assign sum_8[24] = _1818_ ^ _1817_ /*4674*/;
  assign _1819_ = _1818_ & _1817_ /*4673*/;
  assign _1820_ = inv_8[24] & r_7[24] /*4672*/;
  assign _1821_ = _1819_ | _1820_ /*4671*/;
  assign _1822_ = inv_8[25] ^ r_7[25] /*4669*/;
  assign sum_8[25] = _1822_ ^ _1821_ /*4668*/;
  assign _1823_ = _1822_ & _1821_ /*4667*/;
  assign _1824_ = inv_8[25] & r_7[25] /*4666*/;
  assign _1825_ = _1823_ | _1824_ /*4665*/;
  assign _1826_ = inv_8[26] ^ r_7[26] /*4663*/;
  assign sum_8[26] = _1826_ ^ _1825_ /*4662*/;
  assign _1827_ = _1826_ & _1825_ /*4661*/;
  assign _1828_ = inv_8[26] & r_7[26] /*4660*/;
  assign _1829_ = _1827_ | _1828_ /*4659*/;
  assign _1830_ = inv_8[27] ^ r_7[27] /*4657*/;
  assign sum_8[27] = _1830_ ^ _1829_ /*4656*/;
  assign _1831_ = _1830_ & _1829_ /*4655*/;
  assign _1832_ = inv_8[27] & r_7[27] /*4654*/;
  assign _1833_ = _1831_ | _1832_ /*4653*/;
  assign _1834_ = inv_8[28] ^ r_7[28] /*4651*/;
  assign sum_8[28] = _1834_ ^ _1833_ /*4650*/;
  assign _1835_ = _1834_ & _1833_ /*4649*/;
  assign _1836_ = inv_8[28] & r_7[28] /*4648*/;
  assign _1837_ = _1835_ | _1836_ /*4647*/;
  assign _1838_ = inv_8[29] ^ r_7[29] /*4645*/;
  assign sum_8[29] = _1838_ ^ _1837_ /*4644*/;
  assign _1839_ = _1838_ & _1837_ /*4643*/;
  assign _1840_ = inv_8[29] & r_7[29] /*4642*/;
  assign _1841_ = _1839_ | _1840_ /*4641*/;
  assign _1842_ = inv_8[30] ^ r_7[30] /*4639*/;
  assign sum_8[30] = _1842_ ^ _1841_ /*4638*/;
  assign _1843_ = _1842_ & _1841_ /*4637*/;
  assign _1844_ = inv_8[30] & r_7[30] /*4636*/;
  assign _1845_ = _1843_ | _1844_ /*4635*/;
  assign _1846_ = inv_8[31] ^ r_7[31] /*4633*/;
  assign sum_8[31] = _1846_ ^ _1845_ /*4632*/;
  assign _1847_ = _1846_ & _1845_ /*4631*/;
  assign _1848_ = inv_8[31] & r_7[31] /*4630*/;
  assign _1849_ = _1847_ | _1848_ /*4629*/;
  assign _1850_ = inv_8[32] ^ r_7[32] /*4627*/;
  assign sum_8[32] = _1850_ ^ _1849_ /*4626*/;
  assign _1851_ = _1850_ & _1849_ /*4625*/;
  assign _1852_ = inv_8[32] & r_7[32] /*4624*/;
  assign _1853_ = _1851_ | _1852_ /*4623*/;
  assign _1854_ = inv_8[33] ^ r_7[33] /*4621*/;
  assign sum_8[33] = _1854_ ^ _1853_ /*4620*/;
  assign _1855_ = _1854_ & _1853_ /*4619*/;
  assign _1856_ = inv_8[33] & r_7[33] /*4618*/;
  assign _1857_ = _1855_ | _1856_ /*4617*/;
  assign _1858_ = inv_8[34] ^ r_7[34] /*4615*/;
  assign sum_8[34] = _1858_ ^ _1857_ /*4614*/;
  assign _1859_ = _1858_ & _1857_ /*4613*/;
  assign _1860_ = inv_8[34] & r_7[34] /*4612*/;
  assign _1861_ = _1859_ | _1860_ /*4611*/;
  assign _1862_ = inv_8[35] ^ r_7[35] /*4609*/;
  assign sum_8[35] = _1862_ ^ _1861_ /*4608*/;
  assign _1863_ = _1862_ & _1861_ /*4607*/;
  assign _1864_ = inv_8[35] & r_7[35] /*4606*/;
  assign _1865_ = _1863_ | _1864_ /*4605*/;
  assign _1866_ = inv_8[36] ^ r_7[36] /*4603*/;
  assign sum_8[36] = _1866_ ^ _1865_ /*4602*/;
  assign _1867_ = _1866_ & _1865_ /*4601*/;
  assign _1868_ = inv_8[36] & r_7[36] /*4600*/;
  assign _1869_ = _1867_ | _1868_ /*4599*/;
  assign _1870_ = inv_8[37] ^ r_7[37] /*4597*/;
  assign sum_8[37] = _1870_ ^ _1869_ /*4596*/;
  assign _1871_ = _1870_ & _1869_ /*4595*/;
  assign _1872_ = inv_8[37] & r_7[37] /*4594*/;
  assign _1873_ = _1871_ | _1872_ /*4593*/;
  assign _1874_ = _1873_ ^ _1869_ /*4592*/;
  assign _1875_ = ~_1874_ /*4591*/;
  assign _1876_ = sum_8[37] & _1875_ /*4590*/;
  assign _1877_ = _1874_ & _1873_ /*4589*/;
  assign sum_8[38] = _1877_ | _1876_ /*4588*/;
  assign q[8] = ~sum_8[38] /*4587*/;
  assign m_8[0] = r_7[0] /*4586*/;
  assign m_8[1] = r_7[1] /*4585*/;
  assign m_8[2] = r_7[2] /*4584*/;
  assign m_8[3] = r_7[3] /*4583*/;
  assign m_8[4] = r_7[4] /*4582*/;
  assign m_8[5] = r_7[5] /*4581*/;
  assign m_8[6] = r_7[6] /*4580*/;
  assign m_8[7] = r_7[7] /*4579*/;
  assign m_8[8] = r_7[8] /*4578*/;
  assign m_8[9] = r_7[9] /*4577*/;
  assign m_8[10] = r_7[10] /*4576*/;
  assign m_8[11] = r_7[11] /*4575*/;
  assign m_8[12] = r_7[12] /*4574*/;
  assign m_8[13] = r_7[13] /*4573*/;
  assign m_8[14] = r_7[14] /*4572*/;
  assign m_8[15] = r_7[15] /*4571*/;
  assign m_8[16] = r_7[16] /*4570*/;
  assign m_8[17] = r_7[17] /*4569*/;
  assign m_8[18] = r_7[18] /*4568*/;
  assign m_8[19] = r_7[19] /*4567*/;
  assign m_8[20] = r_7[20] /*4566*/;
  assign m_8[21] = r_7[21] /*4565*/;
  assign m_8[22] = r_7[22] /*4564*/;
  assign m_8[23] = r_7[23] /*4563*/;
  assign m_8[24] = r_7[24] /*4562*/;
  assign m_8[25] = r_7[25] /*4561*/;
  assign m_8[26] = r_7[26] /*4560*/;
  assign m_8[27] = r_7[27] /*4559*/;
  assign m_8[28] = r_7[28] /*4558*/;
  assign m_8[29] = r_7[29] /*4557*/;
  assign m_8[30] = r_7[30] /*4556*/;
  assign m_8[31] = r_7[31] /*4555*/;
  assign m_8[32] = r_7[32] /*4554*/;
  assign m_8[33] = r_7[33] /*4553*/;
  assign m_8[34] = r_7[34] /*4552*/;
  assign m_8[35] = r_7[35] /*4551*/;
  assign m_8[36] = r_7[36] /*4550*/;
  assign m_8[37] = r_7[37] /*4549*/;
  assign m_8[38] = r_7[37] /*4548*/;
  assign _1879_ = ~q[8] /*4547*/;
  assign _1880_ = sum_8[0] & q[8] /*4546*/;
  assign _1881_ = m_8[0] & _1879_ /*4545*/;
  assign r_8[0] = _1881_ | _1880_ /*4544*/;
  assign _1882_ = ~q[8] /*4543*/;
  assign _1883_ = sum_8[1] & q[8] /*4542*/;
  assign _1884_ = m_8[1] & _1882_ /*4541*/;
  assign r_8[1] = _1884_ | _1883_ /*4540*/;
  assign _1885_ = ~q[8] /*4539*/;
  assign _1886_ = sum_8[2] & q[8] /*4538*/;
  assign _1887_ = m_8[2] & _1885_ /*4537*/;
  assign r_8[2] = _1887_ | _1886_ /*4536*/;
  assign _1888_ = ~q[8] /*4535*/;
  assign _1889_ = sum_8[3] & q[8] /*4534*/;
  assign _1890_ = m_8[3] & _1888_ /*4533*/;
  assign r_8[3] = _1890_ | _1889_ /*4532*/;
  assign _1891_ = ~q[8] /*4531*/;
  assign _1892_ = sum_8[4] & q[8] /*4530*/;
  assign _1893_ = m_8[4] & _1891_ /*4529*/;
  assign r_8[4] = _1893_ | _1892_ /*4528*/;
  assign _1894_ = ~q[8] /*4527*/;
  assign _1895_ = sum_8[5] & q[8] /*4526*/;
  assign _1896_ = m_8[5] & _1894_ /*4525*/;
  assign r_8[5] = _1896_ | _1895_ /*4524*/;
  assign _1897_ = ~q[8] /*4523*/;
  assign _1898_ = sum_8[6] & q[8] /*4522*/;
  assign _1899_ = m_8[6] & _1897_ /*4521*/;
  assign r_8[6] = _1899_ | _1898_ /*4520*/;
  assign _1900_ = ~q[8] /*4519*/;
  assign _1901_ = sum_8[7] & q[8] /*4518*/;
  assign _1902_ = m_8[7] & _1900_ /*4517*/;
  assign r_8[7] = _1902_ | _1901_ /*4516*/;
  assign _1903_ = ~q[8] /*4515*/;
  assign _1904_ = sum_8[8] & q[8] /*4514*/;
  assign _1905_ = m_8[8] & _1903_ /*4513*/;
  assign r_8[8] = _1905_ | _1904_ /*4512*/;
  assign _1906_ = ~q[8] /*4511*/;
  assign _1907_ = sum_8[9] & q[8] /*4510*/;
  assign _1908_ = m_8[9] & _1906_ /*4509*/;
  assign r_8[9] = _1908_ | _1907_ /*4508*/;
  assign _1909_ = ~q[8] /*4507*/;
  assign _1910_ = sum_8[10] & q[8] /*4506*/;
  assign _1911_ = m_8[10] & _1909_ /*4505*/;
  assign r_8[10] = _1911_ | _1910_ /*4504*/;
  assign _1912_ = ~q[8] /*4503*/;
  assign _1913_ = sum_8[11] & q[8] /*4502*/;
  assign _1914_ = m_8[11] & _1912_ /*4501*/;
  assign r_8[11] = _1914_ | _1913_ /*4500*/;
  assign _1915_ = ~q[8] /*4499*/;
  assign _1916_ = sum_8[12] & q[8] /*4498*/;
  assign _1917_ = m_8[12] & _1915_ /*4497*/;
  assign r_8[12] = _1917_ | _1916_ /*4496*/;
  assign _1918_ = ~q[8] /*4495*/;
  assign _1919_ = sum_8[13] & q[8] /*4494*/;
  assign _1920_ = m_8[13] & _1918_ /*4493*/;
  assign r_8[13] = _1920_ | _1919_ /*4492*/;
  assign _1921_ = ~q[8] /*4491*/;
  assign _1922_ = sum_8[14] & q[8] /*4490*/;
  assign _1923_ = m_8[14] & _1921_ /*4489*/;
  assign r_8[14] = _1923_ | _1922_ /*4488*/;
  assign _1924_ = ~q[8] /*4487*/;
  assign _1925_ = sum_8[15] & q[8] /*4486*/;
  assign _1926_ = m_8[15] & _1924_ /*4485*/;
  assign r_8[15] = _1926_ | _1925_ /*4484*/;
  assign _1927_ = ~q[8] /*4483*/;
  assign _1928_ = sum_8[16] & q[8] /*4482*/;
  assign _1929_ = m_8[16] & _1927_ /*4481*/;
  assign r_8[16] = _1929_ | _1928_ /*4480*/;
  assign _1930_ = ~q[8] /*4479*/;
  assign _1931_ = sum_8[17] & q[8] /*4478*/;
  assign _1932_ = m_8[17] & _1930_ /*4477*/;
  assign r_8[17] = _1932_ | _1931_ /*4476*/;
  assign _1933_ = ~q[8] /*4475*/;
  assign _1934_ = sum_8[18] & q[8] /*4474*/;
  assign _1935_ = m_8[18] & _1933_ /*4473*/;
  assign r_8[18] = _1935_ | _1934_ /*4472*/;
  assign _1936_ = ~q[8] /*4471*/;
  assign _1937_ = sum_8[19] & q[8] /*4470*/;
  assign _1938_ = m_8[19] & _1936_ /*4469*/;
  assign r_8[19] = _1938_ | _1937_ /*4468*/;
  assign _1939_ = ~q[8] /*4467*/;
  assign _1940_ = sum_8[20] & q[8] /*4466*/;
  assign _1941_ = m_8[20] & _1939_ /*4465*/;
  assign r_8[20] = _1941_ | _1940_ /*4464*/;
  assign _1942_ = ~q[8] /*4463*/;
  assign _1943_ = sum_8[21] & q[8] /*4462*/;
  assign _1944_ = m_8[21] & _1942_ /*4461*/;
  assign r_8[21] = _1944_ | _1943_ /*4460*/;
  assign _1945_ = ~q[8] /*4459*/;
  assign _1946_ = sum_8[22] & q[8] /*4458*/;
  assign _1947_ = m_8[22] & _1945_ /*4457*/;
  assign r_8[22] = _1947_ | _1946_ /*4456*/;
  assign _1948_ = ~q[8] /*4455*/;
  assign _1949_ = sum_8[23] & q[8] /*4454*/;
  assign _1950_ = m_8[23] & _1948_ /*4453*/;
  assign r_8[23] = _1950_ | _1949_ /*4452*/;
  assign _1951_ = ~q[8] /*4451*/;
  assign _1952_ = sum_8[24] & q[8] /*4450*/;
  assign _1953_ = m_8[24] & _1951_ /*4449*/;
  assign r_8[24] = _1953_ | _1952_ /*4448*/;
  assign _1954_ = ~q[8] /*4447*/;
  assign _1955_ = sum_8[25] & q[8] /*4446*/;
  assign _1956_ = m_8[25] & _1954_ /*4445*/;
  assign r_8[25] = _1956_ | _1955_ /*4444*/;
  assign _1957_ = ~q[8] /*4443*/;
  assign _1958_ = sum_8[26] & q[8] /*4442*/;
  assign _1959_ = m_8[26] & _1957_ /*4441*/;
  assign r_8[26] = _1959_ | _1958_ /*4440*/;
  assign _1960_ = ~q[8] /*4439*/;
  assign _1961_ = sum_8[27] & q[8] /*4438*/;
  assign _1962_ = m_8[27] & _1960_ /*4437*/;
  assign r_8[27] = _1962_ | _1961_ /*4436*/;
  assign _1963_ = ~q[8] /*4435*/;
  assign _1964_ = sum_8[28] & q[8] /*4434*/;
  assign _1965_ = m_8[28] & _1963_ /*4433*/;
  assign r_8[28] = _1965_ | _1964_ /*4432*/;
  assign _1966_ = ~q[8] /*4431*/;
  assign _1967_ = sum_8[29] & q[8] /*4430*/;
  assign _1968_ = m_8[29] & _1966_ /*4429*/;
  assign r_8[29] = _1968_ | _1967_ /*4428*/;
  assign _1969_ = ~q[8] /*4427*/;
  assign _1970_ = sum_8[30] & q[8] /*4426*/;
  assign _1971_ = m_8[30] & _1969_ /*4425*/;
  assign r_8[30] = _1971_ | _1970_ /*4424*/;
  assign _1972_ = ~q[8] /*4423*/;
  assign _1973_ = sum_8[31] & q[8] /*4422*/;
  assign _1974_ = m_8[31] & _1972_ /*4421*/;
  assign r_8[31] = _1974_ | _1973_ /*4420*/;
  assign _1975_ = ~q[8] /*4419*/;
  assign _1976_ = sum_8[32] & q[8] /*4418*/;
  assign _1977_ = m_8[32] & _1975_ /*4417*/;
  assign r_8[32] = _1977_ | _1976_ /*4416*/;
  assign _1978_ = ~q[8] /*4415*/;
  assign _1979_ = sum_8[33] & q[8] /*4414*/;
  assign _1980_ = m_8[33] & _1978_ /*4413*/;
  assign r_8[33] = _1980_ | _1979_ /*4412*/;
  assign _1981_ = ~q[8] /*4411*/;
  assign _1982_ = sum_8[34] & q[8] /*4410*/;
  assign _1983_ = m_8[34] & _1981_ /*4409*/;
  assign r_8[34] = _1983_ | _1982_ /*4408*/;
  assign _1984_ = ~q[8] /*4407*/;
  assign _1985_ = sum_8[35] & q[8] /*4406*/;
  assign _1986_ = m_8[35] & _1984_ /*4405*/;
  assign r_8[35] = _1986_ | _1985_ /*4404*/;
  assign _1987_ = ~q[8] /*4403*/;
  assign _1988_ = sum_8[36] & q[8] /*4402*/;
  assign _1989_ = m_8[36] & _1987_ /*4401*/;
  assign r_8[36] = _1989_ | _1988_ /*4400*/;
  assign _1990_ = ~q[8] /*4399*/;
  assign _1991_ = sum_8[37] & q[8] /*4398*/;
  assign _1992_ = m_8[37] & _1990_ /*4397*/;
  assign r_8[37] = _1992_ | _1991_ /*4396*/;
  assign _1993_ = ~q[8] /*4395*/;
  assign _1994_ = sum_8[38] & q[8] /*4394*/;
  assign _1995_ = m_8[38] & _1993_ /*4393*/;
  assign r_8[38] = _1995_ | _1994_ /*4392*/;
  assign inv_9[0] = oneWire /*4288*/;
  assign inv_9[1] = oneWire /*4282*/;
  assign inv_9[2] = oneWire /*4276*/;
  assign inv_9[3] = oneWire /*4270*/;
  assign inv_9[4] = oneWire /*4264*/;
  assign inv_9[5] = oneWire /*4258*/;
  assign inv_9[6] = oneWire /*4252*/;
  assign inv_9[7] = ~div[0] /*4246*/;
  assign inv_9[8] = ~div[1] /*4240*/;
  assign inv_9[9] = ~div[2] /*4234*/;
  assign inv_9[10] = ~div[3] /*4228*/;
  assign inv_9[11] = ~div[4] /*4222*/;
  assign inv_9[12] = ~div[5] /*4216*/;
  assign inv_9[13] = ~div[6] /*4210*/;
  assign inv_9[14] = ~div[7] /*4204*/;
  assign inv_9[15] = ~div[8] /*4198*/;
  assign inv_9[16] = ~div[9] /*4192*/;
  assign inv_9[17] = ~div[10] /*4186*/;
  assign inv_9[18] = ~div[11] /*4180*/;
  assign inv_9[19] = ~div[12] /*4174*/;
  assign inv_9[20] = ~div[13] /*4168*/;
  assign inv_9[21] = ~div[14] /*4162*/;
  assign inv_9[22] = oneWire /*4156*/;
  assign inv_9[23] = oneWire /*4150*/;
  assign inv_9[24] = oneWire /*4144*/;
  assign inv_9[25] = oneWire /*4138*/;
  assign inv_9[26] = oneWire /*4132*/;
  assign inv_9[27] = oneWire /*4126*/;
  assign inv_9[28] = oneWire /*4120*/;
  assign inv_9[29] = oneWire /*4114*/;
  assign inv_9[30] = oneWire /*4108*/;
  assign inv_9[31] = oneWire /*4102*/;
  assign inv_9[32] = oneWire /*4096*/;
  assign inv_9[33] = oneWire /*4090*/;
  assign inv_9[34] = oneWire /*4084*/;
  assign inv_9[35] = oneWire /*4078*/;
  assign inv_9[36] = oneWire /*4072*/;
  assign inv_9[37] = oneWire /*4066*/;
  assign inv_9[38] = oneWire /*4060*/;
  assign _1996_ = inv_9[0] ^ r_8[0] /*4287*/;
  assign sum_9[0] = _1996_ ^ oneWire /*4286*/;
  assign _1997_ = _1996_ & oneWire /*4285*/;
  assign _1998_ = inv_9[0] & r_8[0] /*4284*/;
  assign _1999_ = _1997_ | _1998_ /*4283*/;
  assign _2000_ = inv_9[1] ^ r_8[1] /*4281*/;
  assign sum_9[1] = _2000_ ^ _1999_ /*4280*/;
  assign _2001_ = _2000_ & _1999_ /*4279*/;
  assign _2002_ = inv_9[1] & r_8[1] /*4278*/;
  assign _2003_ = _2001_ | _2002_ /*4277*/;
  assign _2004_ = inv_9[2] ^ r_8[2] /*4275*/;
  assign sum_9[2] = _2004_ ^ _2003_ /*4274*/;
  assign _2005_ = _2004_ & _2003_ /*4273*/;
  assign _2006_ = inv_9[2] & r_8[2] /*4272*/;
  assign _2007_ = _2005_ | _2006_ /*4271*/;
  assign _2008_ = inv_9[3] ^ r_8[3] /*4269*/;
  assign sum_9[3] = _2008_ ^ _2007_ /*4268*/;
  assign _2009_ = _2008_ & _2007_ /*4267*/;
  assign _2010_ = inv_9[3] & r_8[3] /*4266*/;
  assign _2011_ = _2009_ | _2010_ /*4265*/;
  assign _2012_ = inv_9[4] ^ r_8[4] /*4263*/;
  assign sum_9[4] = _2012_ ^ _2011_ /*4262*/;
  assign _2013_ = _2012_ & _2011_ /*4261*/;
  assign _2014_ = inv_9[4] & r_8[4] /*4260*/;
  assign _2015_ = _2013_ | _2014_ /*4259*/;
  assign _2016_ = inv_9[5] ^ r_8[5] /*4257*/;
  assign sum_9[5] = _2016_ ^ _2015_ /*4256*/;
  assign _2017_ = _2016_ & _2015_ /*4255*/;
  assign _2018_ = inv_9[5] & r_8[5] /*4254*/;
  assign _2019_ = _2017_ | _2018_ /*4253*/;
  assign _2020_ = inv_9[6] ^ r_8[6] /*4251*/;
  assign sum_9[6] = _2020_ ^ _2019_ /*4250*/;
  assign _2021_ = _2020_ & _2019_ /*4249*/;
  assign _2022_ = inv_9[6] & r_8[6] /*4248*/;
  assign _2023_ = _2021_ | _2022_ /*4247*/;
  assign _2024_ = inv_9[7] ^ r_8[7] /*4245*/;
  assign sum_9[7] = _2024_ ^ _2023_ /*4244*/;
  assign _2025_ = _2024_ & _2023_ /*4243*/;
  assign _2026_ = inv_9[7] & r_8[7] /*4242*/;
  assign _2027_ = _2025_ | _2026_ /*4241*/;
  assign _2028_ = inv_9[8] ^ r_8[8] /*4239*/;
  assign sum_9[8] = _2028_ ^ _2027_ /*4238*/;
  assign _2029_ = _2028_ & _2027_ /*4237*/;
  assign _2030_ = inv_9[8] & r_8[8] /*4236*/;
  assign _2031_ = _2029_ | _2030_ /*4235*/;
  assign _2032_ = inv_9[9] ^ r_8[9] /*4233*/;
  assign sum_9[9] = _2032_ ^ _2031_ /*4232*/;
  assign _2033_ = _2032_ & _2031_ /*4231*/;
  assign _2034_ = inv_9[9] & r_8[9] /*4230*/;
  assign _2035_ = _2033_ | _2034_ /*4229*/;
  assign _2036_ = inv_9[10] ^ r_8[10] /*4227*/;
  assign sum_9[10] = _2036_ ^ _2035_ /*4226*/;
  assign _2037_ = _2036_ & _2035_ /*4225*/;
  assign _2038_ = inv_9[10] & r_8[10] /*4224*/;
  assign _2039_ = _2037_ | _2038_ /*4223*/;
  assign _2040_ = inv_9[11] ^ r_8[11] /*4221*/;
  assign sum_9[11] = _2040_ ^ _2039_ /*4220*/;
  assign _2041_ = _2040_ & _2039_ /*4219*/;
  assign _2042_ = inv_9[11] & r_8[11] /*4218*/;
  assign _2043_ = _2041_ | _2042_ /*4217*/;
  assign _2044_ = inv_9[12] ^ r_8[12] /*4215*/;
  assign sum_9[12] = _2044_ ^ _2043_ /*4214*/;
  assign _2045_ = _2044_ & _2043_ /*4213*/;
  assign _2046_ = inv_9[12] & r_8[12] /*4212*/;
  assign _2047_ = _2045_ | _2046_ /*4211*/;
  assign _2048_ = inv_9[13] ^ r_8[13] /*4209*/;
  assign sum_9[13] = _2048_ ^ _2047_ /*4208*/;
  assign _2049_ = _2048_ & _2047_ /*4207*/;
  assign _2050_ = inv_9[13] & r_8[13] /*4206*/;
  assign _2051_ = _2049_ | _2050_ /*4205*/;
  assign _2052_ = inv_9[14] ^ r_8[14] /*4203*/;
  assign sum_9[14] = _2052_ ^ _2051_ /*4202*/;
  assign _2053_ = _2052_ & _2051_ /*4201*/;
  assign _2054_ = inv_9[14] & r_8[14] /*4200*/;
  assign _2055_ = _2053_ | _2054_ /*4199*/;
  assign _2056_ = inv_9[15] ^ r_8[15] /*4197*/;
  assign sum_9[15] = _2056_ ^ _2055_ /*4196*/;
  assign _2057_ = _2056_ & _2055_ /*4195*/;
  assign _2058_ = inv_9[15] & r_8[15] /*4194*/;
  assign _2059_ = _2057_ | _2058_ /*4193*/;
  assign _2060_ = inv_9[16] ^ r_8[16] /*4191*/;
  assign sum_9[16] = _2060_ ^ _2059_ /*4190*/;
  assign _2061_ = _2060_ & _2059_ /*4189*/;
  assign _2062_ = inv_9[16] & r_8[16] /*4188*/;
  assign _2063_ = _2061_ | _2062_ /*4187*/;
  assign _2064_ = inv_9[17] ^ r_8[17] /*4185*/;
  assign sum_9[17] = _2064_ ^ _2063_ /*4184*/;
  assign _2065_ = _2064_ & _2063_ /*4183*/;
  assign _2066_ = inv_9[17] & r_8[17] /*4182*/;
  assign _2067_ = _2065_ | _2066_ /*4181*/;
  assign _2068_ = inv_9[18] ^ r_8[18] /*4179*/;
  assign sum_9[18] = _2068_ ^ _2067_ /*4178*/;
  assign _2069_ = _2068_ & _2067_ /*4177*/;
  assign _2070_ = inv_9[18] & r_8[18] /*4176*/;
  assign _2071_ = _2069_ | _2070_ /*4175*/;
  assign _2072_ = inv_9[19] ^ r_8[19] /*4173*/;
  assign sum_9[19] = _2072_ ^ _2071_ /*4172*/;
  assign _2073_ = _2072_ & _2071_ /*4171*/;
  assign _2074_ = inv_9[19] & r_8[19] /*4170*/;
  assign _2075_ = _2073_ | _2074_ /*4169*/;
  assign _2076_ = inv_9[20] ^ r_8[20] /*4167*/;
  assign sum_9[20] = _2076_ ^ _2075_ /*4166*/;
  assign _2077_ = _2076_ & _2075_ /*4165*/;
  assign _2078_ = inv_9[20] & r_8[20] /*4164*/;
  assign _2079_ = _2077_ | _2078_ /*4163*/;
  assign _2080_ = inv_9[21] ^ r_8[21] /*4161*/;
  assign sum_9[21] = _2080_ ^ _2079_ /*4160*/;
  assign _2081_ = _2080_ & _2079_ /*4159*/;
  assign _2082_ = inv_9[21] & r_8[21] /*4158*/;
  assign _2083_ = _2081_ | _2082_ /*4157*/;
  assign _2084_ = inv_9[22] ^ r_8[22] /*4155*/;
  assign sum_9[22] = _2084_ ^ _2083_ /*4154*/;
  assign _2085_ = _2084_ & _2083_ /*4153*/;
  assign _2086_ = inv_9[22] & r_8[22] /*4152*/;
  assign _2087_ = _2085_ | _2086_ /*4151*/;
  assign _2088_ = inv_9[23] ^ r_8[23] /*4149*/;
  assign sum_9[23] = _2088_ ^ _2087_ /*4148*/;
  assign _2089_ = _2088_ & _2087_ /*4147*/;
  assign _2090_ = inv_9[23] & r_8[23] /*4146*/;
  assign _2091_ = _2089_ | _2090_ /*4145*/;
  assign _2092_ = inv_9[24] ^ r_8[24] /*4143*/;
  assign sum_9[24] = _2092_ ^ _2091_ /*4142*/;
  assign _2093_ = _2092_ & _2091_ /*4141*/;
  assign _2094_ = inv_9[24] & r_8[24] /*4140*/;
  assign _2095_ = _2093_ | _2094_ /*4139*/;
  assign _2096_ = inv_9[25] ^ r_8[25] /*4137*/;
  assign sum_9[25] = _2096_ ^ _2095_ /*4136*/;
  assign _2097_ = _2096_ & _2095_ /*4135*/;
  assign _2098_ = inv_9[25] & r_8[25] /*4134*/;
  assign _2099_ = _2097_ | _2098_ /*4133*/;
  assign _2100_ = inv_9[26] ^ r_8[26] /*4131*/;
  assign sum_9[26] = _2100_ ^ _2099_ /*4130*/;
  assign _2101_ = _2100_ & _2099_ /*4129*/;
  assign _2102_ = inv_9[26] & r_8[26] /*4128*/;
  assign _2103_ = _2101_ | _2102_ /*4127*/;
  assign _2104_ = inv_9[27] ^ r_8[27] /*4125*/;
  assign sum_9[27] = _2104_ ^ _2103_ /*4124*/;
  assign _2105_ = _2104_ & _2103_ /*4123*/;
  assign _2106_ = inv_9[27] & r_8[27] /*4122*/;
  assign _2107_ = _2105_ | _2106_ /*4121*/;
  assign _2108_ = inv_9[28] ^ r_8[28] /*4119*/;
  assign sum_9[28] = _2108_ ^ _2107_ /*4118*/;
  assign _2109_ = _2108_ & _2107_ /*4117*/;
  assign _2110_ = inv_9[28] & r_8[28] /*4116*/;
  assign _2111_ = _2109_ | _2110_ /*4115*/;
  assign _2112_ = inv_9[29] ^ r_8[29] /*4113*/;
  assign sum_9[29] = _2112_ ^ _2111_ /*4112*/;
  assign _2113_ = _2112_ & _2111_ /*4111*/;
  assign _2114_ = inv_9[29] & r_8[29] /*4110*/;
  assign _2115_ = _2113_ | _2114_ /*4109*/;
  assign _2116_ = inv_9[30] ^ r_8[30] /*4107*/;
  assign sum_9[30] = _2116_ ^ _2115_ /*4106*/;
  assign _2117_ = _2116_ & _2115_ /*4105*/;
  assign _2118_ = inv_9[30] & r_8[30] /*4104*/;
  assign _2119_ = _2117_ | _2118_ /*4103*/;
  assign _2120_ = inv_9[31] ^ r_8[31] /*4101*/;
  assign sum_9[31] = _2120_ ^ _2119_ /*4100*/;
  assign _2121_ = _2120_ & _2119_ /*4099*/;
  assign _2122_ = inv_9[31] & r_8[31] /*4098*/;
  assign _2123_ = _2121_ | _2122_ /*4097*/;
  assign _2124_ = inv_9[32] ^ r_8[32] /*4095*/;
  assign sum_9[32] = _2124_ ^ _2123_ /*4094*/;
  assign _2125_ = _2124_ & _2123_ /*4093*/;
  assign _2126_ = inv_9[32] & r_8[32] /*4092*/;
  assign _2127_ = _2125_ | _2126_ /*4091*/;
  assign _2128_ = inv_9[33] ^ r_8[33] /*4089*/;
  assign sum_9[33] = _2128_ ^ _2127_ /*4088*/;
  assign _2129_ = _2128_ & _2127_ /*4087*/;
  assign _2130_ = inv_9[33] & r_8[33] /*4086*/;
  assign _2131_ = _2129_ | _2130_ /*4085*/;
  assign _2132_ = inv_9[34] ^ r_8[34] /*4083*/;
  assign sum_9[34] = _2132_ ^ _2131_ /*4082*/;
  assign _2133_ = _2132_ & _2131_ /*4081*/;
  assign _2134_ = inv_9[34] & r_8[34] /*4080*/;
  assign _2135_ = _2133_ | _2134_ /*4079*/;
  assign _2136_ = inv_9[35] ^ r_8[35] /*4077*/;
  assign sum_9[35] = _2136_ ^ _2135_ /*4076*/;
  assign _2137_ = _2136_ & _2135_ /*4075*/;
  assign _2138_ = inv_9[35] & r_8[35] /*4074*/;
  assign _2139_ = _2137_ | _2138_ /*4073*/;
  assign _2140_ = inv_9[36] ^ r_8[36] /*4071*/;
  assign sum_9[36] = _2140_ ^ _2139_ /*4070*/;
  assign _2141_ = _2140_ & _2139_ /*4069*/;
  assign _2142_ = inv_9[36] & r_8[36] /*4068*/;
  assign _2143_ = _2141_ | _2142_ /*4067*/;
  assign _2144_ = inv_9[37] ^ r_8[37] /*4065*/;
  assign sum_9[37] = _2144_ ^ _2143_ /*4064*/;
  assign _2145_ = _2144_ & _2143_ /*4063*/;
  assign _2146_ = inv_9[37] & r_8[37] /*4062*/;
  assign _2147_ = _2145_ | _2146_ /*4061*/;
  assign _2148_ = inv_9[38] ^ r_8[38] /*4059*/;
  assign sum_9[38] = _2148_ ^ _2147_ /*4058*/;
  assign _2149_ = _2148_ & _2147_ /*4057*/;
  assign _2150_ = inv_9[38] & r_8[38] /*4056*/;
  assign _2151_ = _2149_ | _2150_ /*4055*/;
  assign _2152_ = _2151_ ^ _2147_ /*4054*/;
  assign _2153_ = ~_2152_ /*4053*/;
  assign _2154_ = sum_9[38] & _2153_ /*4052*/;
  assign _2155_ = _2152_ & _2151_ /*4051*/;
  assign sum_9[39] = _2155_ | _2154_ /*4050*/;
  assign q[7] = ~sum_9[39] /*4049*/;
  assign m_9[0] = r_8[0] /*4048*/;
  assign m_9[1] = r_8[1] /*4047*/;
  assign m_9[2] = r_8[2] /*4046*/;
  assign m_9[3] = r_8[3] /*4045*/;
  assign m_9[4] = r_8[4] /*4044*/;
  assign m_9[5] = r_8[5] /*4043*/;
  assign m_9[6] = r_8[6] /*4042*/;
  assign m_9[7] = r_8[7] /*4041*/;
  assign m_9[8] = r_8[8] /*4040*/;
  assign m_9[9] = r_8[9] /*4039*/;
  assign m_9[10] = r_8[10] /*4038*/;
  assign m_9[11] = r_8[11] /*4037*/;
  assign m_9[12] = r_8[12] /*4036*/;
  assign m_9[13] = r_8[13] /*4035*/;
  assign m_9[14] = r_8[14] /*4034*/;
  assign m_9[15] = r_8[15] /*4033*/;
  assign m_9[16] = r_8[16] /*4032*/;
  assign m_9[17] = r_8[17] /*4031*/;
  assign m_9[18] = r_8[18] /*4030*/;
  assign m_9[19] = r_8[19] /*4029*/;
  assign m_9[20] = r_8[20] /*4028*/;
  assign m_9[21] = r_8[21] /*4027*/;
  assign m_9[22] = r_8[22] /*4026*/;
  assign m_9[23] = r_8[23] /*4025*/;
  assign m_9[24] = r_8[24] /*4024*/;
  assign m_9[25] = r_8[25] /*4023*/;
  assign m_9[26] = r_8[26] /*4022*/;
  assign m_9[27] = r_8[27] /*4021*/;
  assign m_9[28] = r_8[28] /*4020*/;
  assign m_9[29] = r_8[29] /*4019*/;
  assign m_9[30] = r_8[30] /*4018*/;
  assign m_9[31] = r_8[31] /*4017*/;
  assign m_9[32] = r_8[32] /*4016*/;
  assign m_9[33] = r_8[33] /*4015*/;
  assign m_9[34] = r_8[34] /*4014*/;
  assign m_9[35] = r_8[35] /*4013*/;
  assign m_9[36] = r_8[36] /*4012*/;
  assign m_9[37] = r_8[37] /*4011*/;
  assign m_9[38] = r_8[38] /*4010*/;
  assign m_9[39] = r_8[38] /*4009*/;
  assign _2157_ = ~q[7] /*4008*/;
  assign _2158_ = sum_9[0] & q[7] /*4007*/;
  assign _2159_ = m_9[0] & _2157_ /*4006*/;
  assign r_9[0] = _2159_ | _2158_ /*4005*/;
  assign _2160_ = ~q[7] /*4004*/;
  assign _2161_ = sum_9[1] & q[7] /*4003*/;
  assign _2162_ = m_9[1] & _2160_ /*4002*/;
  assign r_9[1] = _2162_ | _2161_ /*4001*/;
  assign _2163_ = ~q[7] /*4000*/;
  assign _2164_ = sum_9[2] & q[7] /*3999*/;
  assign _2165_ = m_9[2] & _2163_ /*3998*/;
  assign r_9[2] = _2165_ | _2164_ /*3997*/;
  assign _2166_ = ~q[7] /*3996*/;
  assign _2167_ = sum_9[3] & q[7] /*3995*/;
  assign _2168_ = m_9[3] & _2166_ /*3994*/;
  assign r_9[3] = _2168_ | _2167_ /*3993*/;
  assign _2169_ = ~q[7] /*3992*/;
  assign _2170_ = sum_9[4] & q[7] /*3991*/;
  assign _2171_ = m_9[4] & _2169_ /*3990*/;
  assign r_9[4] = _2171_ | _2170_ /*3989*/;
  assign _2172_ = ~q[7] /*3988*/;
  assign _2173_ = sum_9[5] & q[7] /*3987*/;
  assign _2174_ = m_9[5] & _2172_ /*3986*/;
  assign r_9[5] = _2174_ | _2173_ /*3985*/;
  assign _2175_ = ~q[7] /*3984*/;
  assign _2176_ = sum_9[6] & q[7] /*3983*/;
  assign _2177_ = m_9[6] & _2175_ /*3982*/;
  assign r_9[6] = _2177_ | _2176_ /*3981*/;
  assign _2178_ = ~q[7] /*3980*/;
  assign _2179_ = sum_9[7] & q[7] /*3979*/;
  assign _2180_ = m_9[7] & _2178_ /*3978*/;
  assign r_9[7] = _2180_ | _2179_ /*3977*/;
  assign _2181_ = ~q[7] /*3976*/;
  assign _2182_ = sum_9[8] & q[7] /*3975*/;
  assign _2183_ = m_9[8] & _2181_ /*3974*/;
  assign r_9[8] = _2183_ | _2182_ /*3973*/;
  assign _2184_ = ~q[7] /*3972*/;
  assign _2185_ = sum_9[9] & q[7] /*3971*/;
  assign _2186_ = m_9[9] & _2184_ /*3970*/;
  assign r_9[9] = _2186_ | _2185_ /*3969*/;
  assign _2187_ = ~q[7] /*3968*/;
  assign _2188_ = sum_9[10] & q[7] /*3967*/;
  assign _2189_ = m_9[10] & _2187_ /*3966*/;
  assign r_9[10] = _2189_ | _2188_ /*3965*/;
  assign _2190_ = ~q[7] /*3964*/;
  assign _2191_ = sum_9[11] & q[7] /*3963*/;
  assign _2192_ = m_9[11] & _2190_ /*3962*/;
  assign r_9[11] = _2192_ | _2191_ /*3961*/;
  assign _2193_ = ~q[7] /*3960*/;
  assign _2194_ = sum_9[12] & q[7] /*3959*/;
  assign _2195_ = m_9[12] & _2193_ /*3958*/;
  assign r_9[12] = _2195_ | _2194_ /*3957*/;
  assign _2196_ = ~q[7] /*3956*/;
  assign _2197_ = sum_9[13] & q[7] /*3955*/;
  assign _2198_ = m_9[13] & _2196_ /*3954*/;
  assign r_9[13] = _2198_ | _2197_ /*3953*/;
  assign _2199_ = ~q[7] /*3952*/;
  assign _2200_ = sum_9[14] & q[7] /*3951*/;
  assign _2201_ = m_9[14] & _2199_ /*3950*/;
  assign r_9[14] = _2201_ | _2200_ /*3949*/;
  assign _2202_ = ~q[7] /*3948*/;
  assign _2203_ = sum_9[15] & q[7] /*3947*/;
  assign _2204_ = m_9[15] & _2202_ /*3946*/;
  assign r_9[15] = _2204_ | _2203_ /*3945*/;
  assign _2205_ = ~q[7] /*3944*/;
  assign _2206_ = sum_9[16] & q[7] /*3943*/;
  assign _2207_ = m_9[16] & _2205_ /*3942*/;
  assign r_9[16] = _2207_ | _2206_ /*3941*/;
  assign _2208_ = ~q[7] /*3940*/;
  assign _2209_ = sum_9[17] & q[7] /*3939*/;
  assign _2210_ = m_9[17] & _2208_ /*3938*/;
  assign r_9[17] = _2210_ | _2209_ /*3937*/;
  assign _2211_ = ~q[7] /*3936*/;
  assign _2212_ = sum_9[18] & q[7] /*3935*/;
  assign _2213_ = m_9[18] & _2211_ /*3934*/;
  assign r_9[18] = _2213_ | _2212_ /*3933*/;
  assign _2214_ = ~q[7] /*3932*/;
  assign _2215_ = sum_9[19] & q[7] /*3931*/;
  assign _2216_ = m_9[19] & _2214_ /*3930*/;
  assign r_9[19] = _2216_ | _2215_ /*3929*/;
  assign _2217_ = ~q[7] /*3928*/;
  assign _2218_ = sum_9[20] & q[7] /*3927*/;
  assign _2219_ = m_9[20] & _2217_ /*3926*/;
  assign r_9[20] = _2219_ | _2218_ /*3925*/;
  assign _2220_ = ~q[7] /*3924*/;
  assign _2221_ = sum_9[21] & q[7] /*3923*/;
  assign _2222_ = m_9[21] & _2220_ /*3922*/;
  assign r_9[21] = _2222_ | _2221_ /*3921*/;
  assign _2223_ = ~q[7] /*3920*/;
  assign _2224_ = sum_9[22] & q[7] /*3919*/;
  assign _2225_ = m_9[22] & _2223_ /*3918*/;
  assign r_9[22] = _2225_ | _2224_ /*3917*/;
  assign _2226_ = ~q[7] /*3916*/;
  assign _2227_ = sum_9[23] & q[7] /*3915*/;
  assign _2228_ = m_9[23] & _2226_ /*3914*/;
  assign r_9[23] = _2228_ | _2227_ /*3913*/;
  assign _2229_ = ~q[7] /*3912*/;
  assign _2230_ = sum_9[24] & q[7] /*3911*/;
  assign _2231_ = m_9[24] & _2229_ /*3910*/;
  assign r_9[24] = _2231_ | _2230_ /*3909*/;
  assign _2232_ = ~q[7] /*3908*/;
  assign _2233_ = sum_9[25] & q[7] /*3907*/;
  assign _2234_ = m_9[25] & _2232_ /*3906*/;
  assign r_9[25] = _2234_ | _2233_ /*3905*/;
  assign _2235_ = ~q[7] /*3904*/;
  assign _2236_ = sum_9[26] & q[7] /*3903*/;
  assign _2237_ = m_9[26] & _2235_ /*3902*/;
  assign r_9[26] = _2237_ | _2236_ /*3901*/;
  assign _2238_ = ~q[7] /*3900*/;
  assign _2239_ = sum_9[27] & q[7] /*3899*/;
  assign _2240_ = m_9[27] & _2238_ /*3898*/;
  assign r_9[27] = _2240_ | _2239_ /*3897*/;
  assign _2241_ = ~q[7] /*3896*/;
  assign _2242_ = sum_9[28] & q[7] /*3895*/;
  assign _2243_ = m_9[28] & _2241_ /*3894*/;
  assign r_9[28] = _2243_ | _2242_ /*3893*/;
  assign _2244_ = ~q[7] /*3892*/;
  assign _2245_ = sum_9[29] & q[7] /*3891*/;
  assign _2246_ = m_9[29] & _2244_ /*3890*/;
  assign r_9[29] = _2246_ | _2245_ /*3889*/;
  assign _2247_ = ~q[7] /*3888*/;
  assign _2248_ = sum_9[30] & q[7] /*3887*/;
  assign _2249_ = m_9[30] & _2247_ /*3886*/;
  assign r_9[30] = _2249_ | _2248_ /*3885*/;
  assign _2250_ = ~q[7] /*3884*/;
  assign _2251_ = sum_9[31] & q[7] /*3883*/;
  assign _2252_ = m_9[31] & _2250_ /*3882*/;
  assign r_9[31] = _2252_ | _2251_ /*3881*/;
  assign _2253_ = ~q[7] /*3880*/;
  assign _2254_ = sum_9[32] & q[7] /*3879*/;
  assign _2255_ = m_9[32] & _2253_ /*3878*/;
  assign r_9[32] = _2255_ | _2254_ /*3877*/;
  assign _2256_ = ~q[7] /*3876*/;
  assign _2257_ = sum_9[33] & q[7] /*3875*/;
  assign _2258_ = m_9[33] & _2256_ /*3874*/;
  assign r_9[33] = _2258_ | _2257_ /*3873*/;
  assign _2259_ = ~q[7] /*3872*/;
  assign _2260_ = sum_9[34] & q[7] /*3871*/;
  assign _2261_ = m_9[34] & _2259_ /*3870*/;
  assign r_9[34] = _2261_ | _2260_ /*3869*/;
  assign _2262_ = ~q[7] /*3868*/;
  assign _2263_ = sum_9[35] & q[7] /*3867*/;
  assign _2264_ = m_9[35] & _2262_ /*3866*/;
  assign r_9[35] = _2264_ | _2263_ /*3865*/;
  assign _2265_ = ~q[7] /*3864*/;
  assign _2266_ = sum_9[36] & q[7] /*3863*/;
  assign _2267_ = m_9[36] & _2265_ /*3862*/;
  assign r_9[36] = _2267_ | _2266_ /*3861*/;
  assign _2268_ = ~q[7] /*3860*/;
  assign _2269_ = sum_9[37] & q[7] /*3859*/;
  assign _2270_ = m_9[37] & _2268_ /*3858*/;
  assign r_9[37] = _2270_ | _2269_ /*3857*/;
  assign _2271_ = ~q[7] /*3856*/;
  assign _2272_ = sum_9[38] & q[7] /*3855*/;
  assign _2273_ = m_9[38] & _2271_ /*3854*/;
  assign r_9[38] = _2273_ | _2272_ /*3853*/;
  assign _2274_ = ~q[7] /*3852*/;
  assign _2275_ = sum_9[39] & q[7] /*3851*/;
  assign _2276_ = m_9[39] & _2274_ /*3850*/;
  assign r_9[39] = _2276_ | _2275_ /*3849*/;
  assign inv_10[0] = oneWire /*3756*/;
  assign inv_10[1] = oneWire /*3750*/;
  assign inv_10[2] = oneWire /*3744*/;
  assign inv_10[3] = oneWire /*3738*/;
  assign inv_10[4] = oneWire /*3732*/;
  assign inv_10[5] = oneWire /*3726*/;
  assign inv_10[6] = ~div[0] /*3720*/;
  assign inv_10[7] = ~div[1] /*3714*/;
  assign inv_10[8] = ~div[2] /*3708*/;
  assign inv_10[9] = ~div[3] /*3702*/;
  assign inv_10[10] = ~div[4] /*3696*/;
  assign inv_10[11] = ~div[5] /*3690*/;
  assign inv_10[12] = ~div[6] /*3684*/;
  assign inv_10[13] = ~div[7] /*3678*/;
  assign inv_10[14] = ~div[8] /*3672*/;
  assign inv_10[15] = ~div[9] /*3666*/;
  assign inv_10[16] = ~div[10] /*3660*/;
  assign inv_10[17] = ~div[11] /*3654*/;
  assign inv_10[18] = ~div[12] /*3648*/;
  assign inv_10[19] = ~div[13] /*3642*/;
  assign inv_10[20] = ~div[14] /*3636*/;
  assign inv_10[21] = oneWire /*3630*/;
  assign inv_10[22] = oneWire /*3624*/;
  assign inv_10[23] = oneWire /*3618*/;
  assign inv_10[24] = oneWire /*3612*/;
  assign inv_10[25] = oneWire /*3606*/;
  assign inv_10[26] = oneWire /*3600*/;
  assign inv_10[27] = oneWire /*3594*/;
  assign inv_10[28] = oneWire /*3588*/;
  assign inv_10[29] = oneWire /*3582*/;
  assign inv_10[30] = oneWire /*3576*/;
  assign inv_10[31] = oneWire /*3570*/;
  assign inv_10[32] = oneWire /*3564*/;
  assign inv_10[33] = oneWire /*3558*/;
  assign inv_10[34] = oneWire /*3552*/;
  assign inv_10[35] = oneWire /*3546*/;
  assign inv_10[36] = oneWire /*3540*/;
  assign inv_10[37] = oneWire /*3534*/;
  assign inv_10[38] = oneWire /*3528*/;
  assign inv_10[39] = oneWire /*3522*/;
  assign _2277_ = inv_10[0] ^ r_9[0] /*3755*/;
  assign sum_10[0] = _2277_ ^ oneWire /*3754*/;
  assign _2278_ = _2277_ & oneWire /*3753*/;
  assign _2279_ = inv_10[0] & r_9[0] /*3752*/;
  assign _2280_ = _2278_ | _2279_ /*3751*/;
  assign _2281_ = inv_10[1] ^ r_9[1] /*3749*/;
  assign sum_10[1] = _2281_ ^ _2280_ /*3748*/;
  assign _2282_ = _2281_ & _2280_ /*3747*/;
  assign _2283_ = inv_10[1] & r_9[1] /*3746*/;
  assign _2284_ = _2282_ | _2283_ /*3745*/;
  assign _2285_ = inv_10[2] ^ r_9[2] /*3743*/;
  assign sum_10[2] = _2285_ ^ _2284_ /*3742*/;
  assign _2286_ = _2285_ & _2284_ /*3741*/;
  assign _2287_ = inv_10[2] & r_9[2] /*3740*/;
  assign _2288_ = _2286_ | _2287_ /*3739*/;
  assign _2289_ = inv_10[3] ^ r_9[3] /*3737*/;
  assign sum_10[3] = _2289_ ^ _2288_ /*3736*/;
  assign _2290_ = _2289_ & _2288_ /*3735*/;
  assign _2291_ = inv_10[3] & r_9[3] /*3734*/;
  assign _2292_ = _2290_ | _2291_ /*3733*/;
  assign _2293_ = inv_10[4] ^ r_9[4] /*3731*/;
  assign sum_10[4] = _2293_ ^ _2292_ /*3730*/;
  assign _2294_ = _2293_ & _2292_ /*3729*/;
  assign _2295_ = inv_10[4] & r_9[4] /*3728*/;
  assign _2296_ = _2294_ | _2295_ /*3727*/;
  assign _2297_ = inv_10[5] ^ r_9[5] /*3725*/;
  assign sum_10[5] = _2297_ ^ _2296_ /*3724*/;
  assign _2298_ = _2297_ & _2296_ /*3723*/;
  assign _2299_ = inv_10[5] & r_9[5] /*3722*/;
  assign _2300_ = _2298_ | _2299_ /*3721*/;
  assign _2301_ = inv_10[6] ^ r_9[6] /*3719*/;
  assign sum_10[6] = _2301_ ^ _2300_ /*3718*/;
  assign _2302_ = _2301_ & _2300_ /*3717*/;
  assign _2303_ = inv_10[6] & r_9[6] /*3716*/;
  assign _2304_ = _2302_ | _2303_ /*3715*/;
  assign _2305_ = inv_10[7] ^ r_9[7] /*3713*/;
  assign sum_10[7] = _2305_ ^ _2304_ /*3712*/;
  assign _2306_ = _2305_ & _2304_ /*3711*/;
  assign _2307_ = inv_10[7] & r_9[7] /*3710*/;
  assign _2308_ = _2306_ | _2307_ /*3709*/;
  assign _2309_ = inv_10[8] ^ r_9[8] /*3707*/;
  assign sum_10[8] = _2309_ ^ _2308_ /*3706*/;
  assign _2310_ = _2309_ & _2308_ /*3705*/;
  assign _2311_ = inv_10[8] & r_9[8] /*3704*/;
  assign _2312_ = _2310_ | _2311_ /*3703*/;
  assign _2313_ = inv_10[9] ^ r_9[9] /*3701*/;
  assign sum_10[9] = _2313_ ^ _2312_ /*3700*/;
  assign _2314_ = _2313_ & _2312_ /*3699*/;
  assign _2315_ = inv_10[9] & r_9[9] /*3698*/;
  assign _2316_ = _2314_ | _2315_ /*3697*/;
  assign _2317_ = inv_10[10] ^ r_9[10] /*3695*/;
  assign sum_10[10] = _2317_ ^ _2316_ /*3694*/;
  assign _2318_ = _2317_ & _2316_ /*3693*/;
  assign _2319_ = inv_10[10] & r_9[10] /*3692*/;
  assign _2320_ = _2318_ | _2319_ /*3691*/;
  assign _2321_ = inv_10[11] ^ r_9[11] /*3689*/;
  assign sum_10[11] = _2321_ ^ _2320_ /*3688*/;
  assign _2322_ = _2321_ & _2320_ /*3687*/;
  assign _2323_ = inv_10[11] & r_9[11] /*3686*/;
  assign _2324_ = _2322_ | _2323_ /*3685*/;
  assign _2325_ = inv_10[12] ^ r_9[12] /*3683*/;
  assign sum_10[12] = _2325_ ^ _2324_ /*3682*/;
  assign _2326_ = _2325_ & _2324_ /*3681*/;
  assign _2327_ = inv_10[12] & r_9[12] /*3680*/;
  assign _2328_ = _2326_ | _2327_ /*3679*/;
  assign _2329_ = inv_10[13] ^ r_9[13] /*3677*/;
  assign sum_10[13] = _2329_ ^ _2328_ /*3676*/;
  assign _2330_ = _2329_ & _2328_ /*3675*/;
  assign _2331_ = inv_10[13] & r_9[13] /*3674*/;
  assign _2332_ = _2330_ | _2331_ /*3673*/;
  assign _2333_ = inv_10[14] ^ r_9[14] /*3671*/;
  assign sum_10[14] = _2333_ ^ _2332_ /*3670*/;
  assign _2334_ = _2333_ & _2332_ /*3669*/;
  assign _2335_ = inv_10[14] & r_9[14] /*3668*/;
  assign _2336_ = _2334_ | _2335_ /*3667*/;
  assign _2337_ = inv_10[15] ^ r_9[15] /*3665*/;
  assign sum_10[15] = _2337_ ^ _2336_ /*3664*/;
  assign _2338_ = _2337_ & _2336_ /*3663*/;
  assign _2339_ = inv_10[15] & r_9[15] /*3662*/;
  assign _2340_ = _2338_ | _2339_ /*3661*/;
  assign _2341_ = inv_10[16] ^ r_9[16] /*3659*/;
  assign sum_10[16] = _2341_ ^ _2340_ /*3658*/;
  assign _2342_ = _2341_ & _2340_ /*3657*/;
  assign _2343_ = inv_10[16] & r_9[16] /*3656*/;
  assign _2344_ = _2342_ | _2343_ /*3655*/;
  assign _2345_ = inv_10[17] ^ r_9[17] /*3653*/;
  assign sum_10[17] = _2345_ ^ _2344_ /*3652*/;
  assign _2346_ = _2345_ & _2344_ /*3651*/;
  assign _2347_ = inv_10[17] & r_9[17] /*3650*/;
  assign _2348_ = _2346_ | _2347_ /*3649*/;
  assign _2349_ = inv_10[18] ^ r_9[18] /*3647*/;
  assign sum_10[18] = _2349_ ^ _2348_ /*3646*/;
  assign _2350_ = _2349_ & _2348_ /*3645*/;
  assign _2351_ = inv_10[18] & r_9[18] /*3644*/;
  assign _2352_ = _2350_ | _2351_ /*3643*/;
  assign _2353_ = inv_10[19] ^ r_9[19] /*3641*/;
  assign sum_10[19] = _2353_ ^ _2352_ /*3640*/;
  assign _2354_ = _2353_ & _2352_ /*3639*/;
  assign _2355_ = inv_10[19] & r_9[19] /*3638*/;
  assign _2356_ = _2354_ | _2355_ /*3637*/;
  assign _2357_ = inv_10[20] ^ r_9[20] /*3635*/;
  assign sum_10[20] = _2357_ ^ _2356_ /*3634*/;
  assign _2358_ = _2357_ & _2356_ /*3633*/;
  assign _2359_ = inv_10[20] & r_9[20] /*3632*/;
  assign _2360_ = _2358_ | _2359_ /*3631*/;
  assign _2361_ = inv_10[21] ^ r_9[21] /*3629*/;
  assign sum_10[21] = _2361_ ^ _2360_ /*3628*/;
  assign _2362_ = _2361_ & _2360_ /*3627*/;
  assign _2363_ = inv_10[21] & r_9[21] /*3626*/;
  assign _2364_ = _2362_ | _2363_ /*3625*/;
  assign _2365_ = inv_10[22] ^ r_9[22] /*3623*/;
  assign sum_10[22] = _2365_ ^ _2364_ /*3622*/;
  assign _2366_ = _2365_ & _2364_ /*3621*/;
  assign _2367_ = inv_10[22] & r_9[22] /*3620*/;
  assign _2368_ = _2366_ | _2367_ /*3619*/;
  assign _2369_ = inv_10[23] ^ r_9[23] /*3617*/;
  assign sum_10[23] = _2369_ ^ _2368_ /*3616*/;
  assign _2370_ = _2369_ & _2368_ /*3615*/;
  assign _2371_ = inv_10[23] & r_9[23] /*3614*/;
  assign _2372_ = _2370_ | _2371_ /*3613*/;
  assign _2373_ = inv_10[24] ^ r_9[24] /*3611*/;
  assign sum_10[24] = _2373_ ^ _2372_ /*3610*/;
  assign _2374_ = _2373_ & _2372_ /*3609*/;
  assign _2375_ = inv_10[24] & r_9[24] /*3608*/;
  assign _2376_ = _2374_ | _2375_ /*3607*/;
  assign _2377_ = inv_10[25] ^ r_9[25] /*3605*/;
  assign sum_10[25] = _2377_ ^ _2376_ /*3604*/;
  assign _2378_ = _2377_ & _2376_ /*3603*/;
  assign _2379_ = inv_10[25] & r_9[25] /*3602*/;
  assign _2380_ = _2378_ | _2379_ /*3601*/;
  assign _2381_ = inv_10[26] ^ r_9[26] /*3599*/;
  assign sum_10[26] = _2381_ ^ _2380_ /*3598*/;
  assign _2382_ = _2381_ & _2380_ /*3597*/;
  assign _2383_ = inv_10[26] & r_9[26] /*3596*/;
  assign _2384_ = _2382_ | _2383_ /*3595*/;
  assign _2385_ = inv_10[27] ^ r_9[27] /*3593*/;
  assign sum_10[27] = _2385_ ^ _2384_ /*3592*/;
  assign _2386_ = _2385_ & _2384_ /*3591*/;
  assign _2387_ = inv_10[27] & r_9[27] /*3590*/;
  assign _2388_ = _2386_ | _2387_ /*3589*/;
  assign _2389_ = inv_10[28] ^ r_9[28] /*3587*/;
  assign sum_10[28] = _2389_ ^ _2388_ /*3586*/;
  assign _2390_ = _2389_ & _2388_ /*3585*/;
  assign _2391_ = inv_10[28] & r_9[28] /*3584*/;
  assign _2392_ = _2390_ | _2391_ /*3583*/;
  assign _2393_ = inv_10[29] ^ r_9[29] /*3581*/;
  assign sum_10[29] = _2393_ ^ _2392_ /*3580*/;
  assign _2394_ = _2393_ & _2392_ /*3579*/;
  assign _2395_ = inv_10[29] & r_9[29] /*3578*/;
  assign _2396_ = _2394_ | _2395_ /*3577*/;
  assign _2397_ = inv_10[30] ^ r_9[30] /*3575*/;
  assign sum_10[30] = _2397_ ^ _2396_ /*3574*/;
  assign _2398_ = _2397_ & _2396_ /*3573*/;
  assign _2399_ = inv_10[30] & r_9[30] /*3572*/;
  assign _2400_ = _2398_ | _2399_ /*3571*/;
  assign _2401_ = inv_10[31] ^ r_9[31] /*3569*/;
  assign sum_10[31] = _2401_ ^ _2400_ /*3568*/;
  assign _2402_ = _2401_ & _2400_ /*3567*/;
  assign _2403_ = inv_10[31] & r_9[31] /*3566*/;
  assign _2404_ = _2402_ | _2403_ /*3565*/;
  assign _2405_ = inv_10[32] ^ r_9[32] /*3563*/;
  assign sum_10[32] = _2405_ ^ _2404_ /*3562*/;
  assign _2406_ = _2405_ & _2404_ /*3561*/;
  assign _2407_ = inv_10[32] & r_9[32] /*3560*/;
  assign _2408_ = _2406_ | _2407_ /*3559*/;
  assign _2409_ = inv_10[33] ^ r_9[33] /*3557*/;
  assign sum_10[33] = _2409_ ^ _2408_ /*3556*/;
  assign _2410_ = _2409_ & _2408_ /*3555*/;
  assign _2411_ = inv_10[33] & r_9[33] /*3554*/;
  assign _2412_ = _2410_ | _2411_ /*3553*/;
  assign _2413_ = inv_10[34] ^ r_9[34] /*3551*/;
  assign sum_10[34] = _2413_ ^ _2412_ /*3550*/;
  assign _2414_ = _2413_ & _2412_ /*3549*/;
  assign _2415_ = inv_10[34] & r_9[34] /*3548*/;
  assign _2416_ = _2414_ | _2415_ /*3547*/;
  assign _2417_ = inv_10[35] ^ r_9[35] /*3545*/;
  assign sum_10[35] = _2417_ ^ _2416_ /*3544*/;
  assign _2418_ = _2417_ & _2416_ /*3543*/;
  assign _2419_ = inv_10[35] & r_9[35] /*3542*/;
  assign _2420_ = _2418_ | _2419_ /*3541*/;
  assign _2421_ = inv_10[36] ^ r_9[36] /*3539*/;
  assign sum_10[36] = _2421_ ^ _2420_ /*3538*/;
  assign _2422_ = _2421_ & _2420_ /*3537*/;
  assign _2423_ = inv_10[36] & r_9[36] /*3536*/;
  assign _2424_ = _2422_ | _2423_ /*3535*/;
  assign _2425_ = inv_10[37] ^ r_9[37] /*3533*/;
  assign sum_10[37] = _2425_ ^ _2424_ /*3532*/;
  assign _2426_ = _2425_ & _2424_ /*3531*/;
  assign _2427_ = inv_10[37] & r_9[37] /*3530*/;
  assign _2428_ = _2426_ | _2427_ /*3529*/;
  assign _2429_ = inv_10[38] ^ r_9[38] /*3527*/;
  assign sum_10[38] = _2429_ ^ _2428_ /*3526*/;
  assign _2430_ = _2429_ & _2428_ /*3525*/;
  assign _2431_ = inv_10[38] & r_9[38] /*3524*/;
  assign _2432_ = _2430_ | _2431_ /*3523*/;
  assign _2433_ = inv_10[39] ^ r_9[39] /*3521*/;
  assign sum_10[39] = _2433_ ^ _2432_ /*3520*/;
  assign _2434_ = _2433_ & _2432_ /*3519*/;
  assign _2435_ = inv_10[39] & r_9[39] /*3518*/;
  assign _2436_ = _2434_ | _2435_ /*3517*/;
  assign _2437_ = _2436_ ^ _2432_ /*3516*/;
  assign _2438_ = ~_2437_ /*3515*/;
  assign _2439_ = sum_10[39] & _2438_ /*3514*/;
  assign _2440_ = _2437_ & _2436_ /*3513*/;
  assign sum_10[40] = _2440_ | _2439_ /*3512*/;
  assign q[6] = ~sum_10[40] /*3511*/;
  assign m_10[0] = r_9[0] /*3510*/;
  assign m_10[1] = r_9[1] /*3509*/;
  assign m_10[2] = r_9[2] /*3508*/;
  assign m_10[3] = r_9[3] /*3507*/;
  assign m_10[4] = r_9[4] /*3506*/;
  assign m_10[5] = r_9[5] /*3505*/;
  assign m_10[6] = r_9[6] /*3504*/;
  assign m_10[7] = r_9[7] /*3503*/;
  assign m_10[8] = r_9[8] /*3502*/;
  assign m_10[9] = r_9[9] /*3501*/;
  assign m_10[10] = r_9[10] /*3500*/;
  assign m_10[11] = r_9[11] /*3499*/;
  assign m_10[12] = r_9[12] /*3498*/;
  assign m_10[13] = r_9[13] /*3497*/;
  assign m_10[14] = r_9[14] /*3496*/;
  assign m_10[15] = r_9[15] /*3495*/;
  assign m_10[16] = r_9[16] /*3494*/;
  assign m_10[17] = r_9[17] /*3493*/;
  assign m_10[18] = r_9[18] /*3492*/;
  assign m_10[19] = r_9[19] /*3491*/;
  assign m_10[20] = r_9[20] /*3490*/;
  assign m_10[21] = r_9[21] /*3489*/;
  assign m_10[22] = r_9[22] /*3488*/;
  assign m_10[23] = r_9[23] /*3487*/;
  assign m_10[24] = r_9[24] /*3486*/;
  assign m_10[25] = r_9[25] /*3485*/;
  assign m_10[26] = r_9[26] /*3484*/;
  assign m_10[27] = r_9[27] /*3483*/;
  assign m_10[28] = r_9[28] /*3482*/;
  assign m_10[29] = r_9[29] /*3481*/;
  assign m_10[30] = r_9[30] /*3480*/;
  assign m_10[31] = r_9[31] /*3479*/;
  assign m_10[32] = r_9[32] /*3478*/;
  assign m_10[33] = r_9[33] /*3477*/;
  assign m_10[34] = r_9[34] /*3476*/;
  assign m_10[35] = r_9[35] /*3475*/;
  assign m_10[36] = r_9[36] /*3474*/;
  assign m_10[37] = r_9[37] /*3473*/;
  assign m_10[38] = r_9[38] /*3472*/;
  assign m_10[39] = r_9[39] /*3471*/;
  assign m_10[40] = r_9[39] /*3470*/;
  assign _2442_ = ~q[6] /*3469*/;
  assign _2443_ = sum_10[0] & q[6] /*3468*/;
  assign _2444_ = m_10[0] & _2442_ /*3467*/;
  assign r_10[0] = _2444_ | _2443_ /*3466*/;
  assign _2445_ = ~q[6] /*3465*/;
  assign _2446_ = sum_10[1] & q[6] /*3464*/;
  assign _2447_ = m_10[1] & _2445_ /*3463*/;
  assign r_10[1] = _2447_ | _2446_ /*3462*/;
  assign _2448_ = ~q[6] /*3461*/;
  assign _2449_ = sum_10[2] & q[6] /*3460*/;
  assign _2450_ = m_10[2] & _2448_ /*3459*/;
  assign r_10[2] = _2450_ | _2449_ /*3458*/;
  assign _2451_ = ~q[6] /*3457*/;
  assign _2452_ = sum_10[3] & q[6] /*3456*/;
  assign _2453_ = m_10[3] & _2451_ /*3455*/;
  assign r_10[3] = _2453_ | _2452_ /*3454*/;
  assign _2454_ = ~q[6] /*3453*/;
  assign _2455_ = sum_10[4] & q[6] /*3452*/;
  assign _2456_ = m_10[4] & _2454_ /*3451*/;
  assign r_10[4] = _2456_ | _2455_ /*3450*/;
  assign _2457_ = ~q[6] /*3449*/;
  assign _2458_ = sum_10[5] & q[6] /*3448*/;
  assign _2459_ = m_10[5] & _2457_ /*3447*/;
  assign r_10[5] = _2459_ | _2458_ /*3446*/;
  assign _2460_ = ~q[6] /*3445*/;
  assign _2461_ = sum_10[6] & q[6] /*3444*/;
  assign _2462_ = m_10[6] & _2460_ /*3443*/;
  assign r_10[6] = _2462_ | _2461_ /*3442*/;
  assign _2463_ = ~q[6] /*3441*/;
  assign _2464_ = sum_10[7] & q[6] /*3440*/;
  assign _2465_ = m_10[7] & _2463_ /*3439*/;
  assign r_10[7] = _2465_ | _2464_ /*3438*/;
  assign _2466_ = ~q[6] /*3437*/;
  assign _2467_ = sum_10[8] & q[6] /*3436*/;
  assign _2468_ = m_10[8] & _2466_ /*3435*/;
  assign r_10[8] = _2468_ | _2467_ /*3434*/;
  assign _2469_ = ~q[6] /*3433*/;
  assign _2470_ = sum_10[9] & q[6] /*3432*/;
  assign _2471_ = m_10[9] & _2469_ /*3431*/;
  assign r_10[9] = _2471_ | _2470_ /*3430*/;
  assign _2472_ = ~q[6] /*3429*/;
  assign _2473_ = sum_10[10] & q[6] /*3428*/;
  assign _2474_ = m_10[10] & _2472_ /*3427*/;
  assign r_10[10] = _2474_ | _2473_ /*3426*/;
  assign _2475_ = ~q[6] /*3425*/;
  assign _2476_ = sum_10[11] & q[6] /*3424*/;
  assign _2477_ = m_10[11] & _2475_ /*3423*/;
  assign r_10[11] = _2477_ | _2476_ /*3422*/;
  assign _2478_ = ~q[6] /*3421*/;
  assign _2479_ = sum_10[12] & q[6] /*3420*/;
  assign _2480_ = m_10[12] & _2478_ /*3419*/;
  assign r_10[12] = _2480_ | _2479_ /*3418*/;
  assign _2481_ = ~q[6] /*3417*/;
  assign _2482_ = sum_10[13] & q[6] /*3416*/;
  assign _2483_ = m_10[13] & _2481_ /*3415*/;
  assign r_10[13] = _2483_ | _2482_ /*3414*/;
  assign _2484_ = ~q[6] /*3413*/;
  assign _2485_ = sum_10[14] & q[6] /*3412*/;
  assign _2486_ = m_10[14] & _2484_ /*3411*/;
  assign r_10[14] = _2486_ | _2485_ /*3410*/;
  assign _2487_ = ~q[6] /*3409*/;
  assign _2488_ = sum_10[15] & q[6] /*3408*/;
  assign _2489_ = m_10[15] & _2487_ /*3407*/;
  assign r_10[15] = _2489_ | _2488_ /*3406*/;
  assign _2490_ = ~q[6] /*3405*/;
  assign _2491_ = sum_10[16] & q[6] /*3404*/;
  assign _2492_ = m_10[16] & _2490_ /*3403*/;
  assign r_10[16] = _2492_ | _2491_ /*3402*/;
  assign _2493_ = ~q[6] /*3401*/;
  assign _2494_ = sum_10[17] & q[6] /*3400*/;
  assign _2495_ = m_10[17] & _2493_ /*3399*/;
  assign r_10[17] = _2495_ | _2494_ /*3398*/;
  assign _2496_ = ~q[6] /*3397*/;
  assign _2497_ = sum_10[18] & q[6] /*3396*/;
  assign _2498_ = m_10[18] & _2496_ /*3395*/;
  assign r_10[18] = _2498_ | _2497_ /*3394*/;
  assign _2499_ = ~q[6] /*3393*/;
  assign _2500_ = sum_10[19] & q[6] /*3392*/;
  assign _2501_ = m_10[19] & _2499_ /*3391*/;
  assign r_10[19] = _2501_ | _2500_ /*3390*/;
  assign _2502_ = ~q[6] /*3389*/;
  assign _2503_ = sum_10[20] & q[6] /*3388*/;
  assign _2504_ = m_10[20] & _2502_ /*3387*/;
  assign r_10[20] = _2504_ | _2503_ /*3386*/;
  assign _2505_ = ~q[6] /*3385*/;
  assign _2506_ = sum_10[21] & q[6] /*3384*/;
  assign _2507_ = m_10[21] & _2505_ /*3383*/;
  assign r_10[21] = _2507_ | _2506_ /*3382*/;
  assign _2508_ = ~q[6] /*3381*/;
  assign _2509_ = sum_10[22] & q[6] /*3380*/;
  assign _2510_ = m_10[22] & _2508_ /*3379*/;
  assign r_10[22] = _2510_ | _2509_ /*3378*/;
  assign _2511_ = ~q[6] /*3377*/;
  assign _2512_ = sum_10[23] & q[6] /*3376*/;
  assign _2513_ = m_10[23] & _2511_ /*3375*/;
  assign r_10[23] = _2513_ | _2512_ /*3374*/;
  assign _2514_ = ~q[6] /*3373*/;
  assign _2515_ = sum_10[24] & q[6] /*3372*/;
  assign _2516_ = m_10[24] & _2514_ /*3371*/;
  assign r_10[24] = _2516_ | _2515_ /*3370*/;
  assign _2517_ = ~q[6] /*3369*/;
  assign _2518_ = sum_10[25] & q[6] /*3368*/;
  assign _2519_ = m_10[25] & _2517_ /*3367*/;
  assign r_10[25] = _2519_ | _2518_ /*3366*/;
  assign _2520_ = ~q[6] /*3365*/;
  assign _2521_ = sum_10[26] & q[6] /*3364*/;
  assign _2522_ = m_10[26] & _2520_ /*3363*/;
  assign r_10[26] = _2522_ | _2521_ /*3362*/;
  assign _2523_ = ~q[6] /*3361*/;
  assign _2524_ = sum_10[27] & q[6] /*3360*/;
  assign _2525_ = m_10[27] & _2523_ /*3359*/;
  assign r_10[27] = _2525_ | _2524_ /*3358*/;
  assign _2526_ = ~q[6] /*3357*/;
  assign _2527_ = sum_10[28] & q[6] /*3356*/;
  assign _2528_ = m_10[28] & _2526_ /*3355*/;
  assign r_10[28] = _2528_ | _2527_ /*3354*/;
  assign _2529_ = ~q[6] /*3353*/;
  assign _2530_ = sum_10[29] & q[6] /*3352*/;
  assign _2531_ = m_10[29] & _2529_ /*3351*/;
  assign r_10[29] = _2531_ | _2530_ /*3350*/;
  assign _2532_ = ~q[6] /*3349*/;
  assign _2533_ = sum_10[30] & q[6] /*3348*/;
  assign _2534_ = m_10[30] & _2532_ /*3347*/;
  assign r_10[30] = _2534_ | _2533_ /*3346*/;
  assign _2535_ = ~q[6] /*3345*/;
  assign _2536_ = sum_10[31] & q[6] /*3344*/;
  assign _2537_ = m_10[31] & _2535_ /*3343*/;
  assign r_10[31] = _2537_ | _2536_ /*3342*/;
  assign _2538_ = ~q[6] /*3341*/;
  assign _2539_ = sum_10[32] & q[6] /*3340*/;
  assign _2540_ = m_10[32] & _2538_ /*3339*/;
  assign r_10[32] = _2540_ | _2539_ /*3338*/;
  assign _2541_ = ~q[6] /*3337*/;
  assign _2542_ = sum_10[33] & q[6] /*3336*/;
  assign _2543_ = m_10[33] & _2541_ /*3335*/;
  assign r_10[33] = _2543_ | _2542_ /*3334*/;
  assign _2544_ = ~q[6] /*3333*/;
  assign _2545_ = sum_10[34] & q[6] /*3332*/;
  assign _2546_ = m_10[34] & _2544_ /*3331*/;
  assign r_10[34] = _2546_ | _2545_ /*3330*/;
  assign _2547_ = ~q[6] /*3329*/;
  assign _2548_ = sum_10[35] & q[6] /*3328*/;
  assign _2549_ = m_10[35] & _2547_ /*3327*/;
  assign r_10[35] = _2549_ | _2548_ /*3326*/;
  assign _2550_ = ~q[6] /*3325*/;
  assign _2551_ = sum_10[36] & q[6] /*3324*/;
  assign _2552_ = m_10[36] & _2550_ /*3323*/;
  assign r_10[36] = _2552_ | _2551_ /*3322*/;
  assign _2553_ = ~q[6] /*3321*/;
  assign _2554_ = sum_10[37] & q[6] /*3320*/;
  assign _2555_ = m_10[37] & _2553_ /*3319*/;
  assign r_10[37] = _2555_ | _2554_ /*3318*/;
  assign _2556_ = ~q[6] /*3317*/;
  assign _2557_ = sum_10[38] & q[6] /*3316*/;
  assign _2558_ = m_10[38] & _2556_ /*3315*/;
  assign r_10[38] = _2558_ | _2557_ /*3314*/;
  assign _2559_ = ~q[6] /*3313*/;
  assign _2560_ = sum_10[39] & q[6] /*3312*/;
  assign _2561_ = m_10[39] & _2559_ /*3311*/;
  assign r_10[39] = _2561_ | _2560_ /*3310*/;
  assign _2562_ = ~q[6] /*3309*/;
  assign _2563_ = sum_10[40] & q[6] /*3308*/;
  assign _2564_ = m_10[40] & _2562_ /*3307*/;
  assign r_10[40] = _2564_ | _2563_ /*3306*/;
  assign inv_11[0] = oneWire /*3224*/;
  assign inv_11[1] = oneWire /*3218*/;
  assign inv_11[2] = oneWire /*3212*/;
  assign inv_11[3] = oneWire /*3206*/;
  assign inv_11[4] = oneWire /*3200*/;
  assign inv_11[5] = ~div[0] /*3194*/;
  assign inv_11[6] = ~div[1] /*3188*/;
  assign inv_11[7] = ~div[2] /*3182*/;
  assign inv_11[8] = ~div[3] /*3176*/;
  assign inv_11[9] = ~div[4] /*3170*/;
  assign inv_11[10] = ~div[5] /*3164*/;
  assign inv_11[11] = ~div[6] /*3158*/;
  assign inv_11[12] = ~div[7] /*3152*/;
  assign inv_11[13] = ~div[8] /*3146*/;
  assign inv_11[14] = ~div[9] /*3140*/;
  assign inv_11[15] = ~div[10] /*3134*/;
  assign inv_11[16] = ~div[11] /*3128*/;
  assign inv_11[17] = ~div[12] /*3122*/;
  assign inv_11[18] = ~div[13] /*3116*/;
  assign inv_11[19] = ~div[14] /*3110*/;
  assign inv_11[20] = oneWire /*3104*/;
  assign inv_11[21] = oneWire /*3098*/;
  assign inv_11[22] = oneWire /*3092*/;
  assign inv_11[23] = oneWire /*3086*/;
  assign inv_11[24] = oneWire /*3080*/;
  assign inv_11[25] = oneWire /*3074*/;
  assign inv_11[26] = oneWire /*3068*/;
  assign inv_11[27] = oneWire /*3062*/;
  assign inv_11[28] = oneWire /*3056*/;
  assign inv_11[29] = oneWire /*3050*/;
  assign inv_11[30] = oneWire /*3044*/;
  assign inv_11[31] = oneWire /*3038*/;
  assign inv_11[32] = oneWire /*3032*/;
  assign inv_11[33] = oneWire /*3026*/;
  assign inv_11[34] = oneWire /*3020*/;
  assign inv_11[35] = oneWire /*3014*/;
  assign inv_11[36] = oneWire /*3008*/;
  assign inv_11[37] = oneWire /*3002*/;
  assign inv_11[38] = oneWire /*2996*/;
  assign inv_11[39] = oneWire /*2990*/;
  assign inv_11[40] = oneWire /*2984*/;
  assign _2565_ = inv_11[0] ^ r_10[0] /*3223*/;
  assign sum_11[0] = _2565_ ^ oneWire /*3222*/;
  assign _2566_ = _2565_ & oneWire /*3221*/;
  assign _2567_ = inv_11[0] & r_10[0] /*3220*/;
  assign _2568_ = _2566_ | _2567_ /*3219*/;
  assign _2569_ = inv_11[1] ^ r_10[1] /*3217*/;
  assign sum_11[1] = _2569_ ^ _2568_ /*3216*/;
  assign _2570_ = _2569_ & _2568_ /*3215*/;
  assign _2571_ = inv_11[1] & r_10[1] /*3214*/;
  assign _2572_ = _2570_ | _2571_ /*3213*/;
  assign _2573_ = inv_11[2] ^ r_10[2] /*3211*/;
  assign sum_11[2] = _2573_ ^ _2572_ /*3210*/;
  assign _2574_ = _2573_ & _2572_ /*3209*/;
  assign _2575_ = inv_11[2] & r_10[2] /*3208*/;
  assign _2576_ = _2574_ | _2575_ /*3207*/;
  assign _2577_ = inv_11[3] ^ r_10[3] /*3205*/;
  assign sum_11[3] = _2577_ ^ _2576_ /*3204*/;
  assign _2578_ = _2577_ & _2576_ /*3203*/;
  assign _2579_ = inv_11[3] & r_10[3] /*3202*/;
  assign _2580_ = _2578_ | _2579_ /*3201*/;
  assign _2581_ = inv_11[4] ^ r_10[4] /*3199*/;
  assign sum_11[4] = _2581_ ^ _2580_ /*3198*/;
  assign _2582_ = _2581_ & _2580_ /*3197*/;
  assign _2583_ = inv_11[4] & r_10[4] /*3196*/;
  assign _2584_ = _2582_ | _2583_ /*3195*/;
  assign _2585_ = inv_11[5] ^ r_10[5] /*3193*/;
  assign sum_11[5] = _2585_ ^ _2584_ /*3192*/;
  assign _2586_ = _2585_ & _2584_ /*3191*/;
  assign _2587_ = inv_11[5] & r_10[5] /*3190*/;
  assign _2588_ = _2586_ | _2587_ /*3189*/;
  assign _2589_ = inv_11[6] ^ r_10[6] /*3187*/;
  assign sum_11[6] = _2589_ ^ _2588_ /*3186*/;
  assign _2590_ = _2589_ & _2588_ /*3185*/;
  assign _2591_ = inv_11[6] & r_10[6] /*3184*/;
  assign _2592_ = _2590_ | _2591_ /*3183*/;
  assign _2593_ = inv_11[7] ^ r_10[7] /*3181*/;
  assign sum_11[7] = _2593_ ^ _2592_ /*3180*/;
  assign _2594_ = _2593_ & _2592_ /*3179*/;
  assign _2595_ = inv_11[7] & r_10[7] /*3178*/;
  assign _2596_ = _2594_ | _2595_ /*3177*/;
  assign _2597_ = inv_11[8] ^ r_10[8] /*3175*/;
  assign sum_11[8] = _2597_ ^ _2596_ /*3174*/;
  assign _2598_ = _2597_ & _2596_ /*3173*/;
  assign _2599_ = inv_11[8] & r_10[8] /*3172*/;
  assign _2600_ = _2598_ | _2599_ /*3171*/;
  assign _2601_ = inv_11[9] ^ r_10[9] /*3169*/;
  assign sum_11[9] = _2601_ ^ _2600_ /*3168*/;
  assign _2602_ = _2601_ & _2600_ /*3167*/;
  assign _2603_ = inv_11[9] & r_10[9] /*3166*/;
  assign _2604_ = _2602_ | _2603_ /*3165*/;
  assign _2605_ = inv_11[10] ^ r_10[10] /*3163*/;
  assign sum_11[10] = _2605_ ^ _2604_ /*3162*/;
  assign _2606_ = _2605_ & _2604_ /*3161*/;
  assign _2607_ = inv_11[10] & r_10[10] /*3160*/;
  assign _2608_ = _2606_ | _2607_ /*3159*/;
  assign _2609_ = inv_11[11] ^ r_10[11] /*3157*/;
  assign sum_11[11] = _2609_ ^ _2608_ /*3156*/;
  assign _2610_ = _2609_ & _2608_ /*3155*/;
  assign _2611_ = inv_11[11] & r_10[11] /*3154*/;
  assign _2612_ = _2610_ | _2611_ /*3153*/;
  assign _2613_ = inv_11[12] ^ r_10[12] /*3151*/;
  assign sum_11[12] = _2613_ ^ _2612_ /*3150*/;
  assign _2614_ = _2613_ & _2612_ /*3149*/;
  assign _2615_ = inv_11[12] & r_10[12] /*3148*/;
  assign _2616_ = _2614_ | _2615_ /*3147*/;
  assign _2617_ = inv_11[13] ^ r_10[13] /*3145*/;
  assign sum_11[13] = _2617_ ^ _2616_ /*3144*/;
  assign _2618_ = _2617_ & _2616_ /*3143*/;
  assign _2619_ = inv_11[13] & r_10[13] /*3142*/;
  assign _2620_ = _2618_ | _2619_ /*3141*/;
  assign _2621_ = inv_11[14] ^ r_10[14] /*3139*/;
  assign sum_11[14] = _2621_ ^ _2620_ /*3138*/;
  assign _2622_ = _2621_ & _2620_ /*3137*/;
  assign _2623_ = inv_11[14] & r_10[14] /*3136*/;
  assign _2624_ = _2622_ | _2623_ /*3135*/;
  assign _2625_ = inv_11[15] ^ r_10[15] /*3133*/;
  assign sum_11[15] = _2625_ ^ _2624_ /*3132*/;
  assign _2626_ = _2625_ & _2624_ /*3131*/;
  assign _2627_ = inv_11[15] & r_10[15] /*3130*/;
  assign _2628_ = _2626_ | _2627_ /*3129*/;
  assign _2629_ = inv_11[16] ^ r_10[16] /*3127*/;
  assign sum_11[16] = _2629_ ^ _2628_ /*3126*/;
  assign _2630_ = _2629_ & _2628_ /*3125*/;
  assign _2631_ = inv_11[16] & r_10[16] /*3124*/;
  assign _2632_ = _2630_ | _2631_ /*3123*/;
  assign _2633_ = inv_11[17] ^ r_10[17] /*3121*/;
  assign sum_11[17] = _2633_ ^ _2632_ /*3120*/;
  assign _2634_ = _2633_ & _2632_ /*3119*/;
  assign _2635_ = inv_11[17] & r_10[17] /*3118*/;
  assign _2636_ = _2634_ | _2635_ /*3117*/;
  assign _2637_ = inv_11[18] ^ r_10[18] /*3115*/;
  assign sum_11[18] = _2637_ ^ _2636_ /*3114*/;
  assign _2638_ = _2637_ & _2636_ /*3113*/;
  assign _2639_ = inv_11[18] & r_10[18] /*3112*/;
  assign _2640_ = _2638_ | _2639_ /*3111*/;
  assign _2641_ = inv_11[19] ^ r_10[19] /*3109*/;
  assign sum_11[19] = _2641_ ^ _2640_ /*3108*/;
  assign _2642_ = _2641_ & _2640_ /*3107*/;
  assign _2643_ = inv_11[19] & r_10[19] /*3106*/;
  assign _2644_ = _2642_ | _2643_ /*3105*/;
  assign _2645_ = inv_11[20] ^ r_10[20] /*3103*/;
  assign sum_11[20] = _2645_ ^ _2644_ /*3102*/;
  assign _2646_ = _2645_ & _2644_ /*3101*/;
  assign _2647_ = inv_11[20] & r_10[20] /*3100*/;
  assign _2648_ = _2646_ | _2647_ /*3099*/;
  assign _2649_ = inv_11[21] ^ r_10[21] /*3097*/;
  assign sum_11[21] = _2649_ ^ _2648_ /*3096*/;
  assign _2650_ = _2649_ & _2648_ /*3095*/;
  assign _2651_ = inv_11[21] & r_10[21] /*3094*/;
  assign _2652_ = _2650_ | _2651_ /*3093*/;
  assign _2653_ = inv_11[22] ^ r_10[22] /*3091*/;
  assign sum_11[22] = _2653_ ^ _2652_ /*3090*/;
  assign _2654_ = _2653_ & _2652_ /*3089*/;
  assign _2655_ = inv_11[22] & r_10[22] /*3088*/;
  assign _2656_ = _2654_ | _2655_ /*3087*/;
  assign _2657_ = inv_11[23] ^ r_10[23] /*3085*/;
  assign sum_11[23] = _2657_ ^ _2656_ /*3084*/;
  assign _2658_ = _2657_ & _2656_ /*3083*/;
  assign _2659_ = inv_11[23] & r_10[23] /*3082*/;
  assign _2660_ = _2658_ | _2659_ /*3081*/;
  assign _2661_ = inv_11[24] ^ r_10[24] /*3079*/;
  assign sum_11[24] = _2661_ ^ _2660_ /*3078*/;
  assign _2662_ = _2661_ & _2660_ /*3077*/;
  assign _2663_ = inv_11[24] & r_10[24] /*3076*/;
  assign _2664_ = _2662_ | _2663_ /*3075*/;
  assign _2665_ = inv_11[25] ^ r_10[25] /*3073*/;
  assign sum_11[25] = _2665_ ^ _2664_ /*3072*/;
  assign _2666_ = _2665_ & _2664_ /*3071*/;
  assign _2667_ = inv_11[25] & r_10[25] /*3070*/;
  assign _2668_ = _2666_ | _2667_ /*3069*/;
  assign _2669_ = inv_11[26] ^ r_10[26] /*3067*/;
  assign sum_11[26] = _2669_ ^ _2668_ /*3066*/;
  assign _2670_ = _2669_ & _2668_ /*3065*/;
  assign _2671_ = inv_11[26] & r_10[26] /*3064*/;
  assign _2672_ = _2670_ | _2671_ /*3063*/;
  assign _2673_ = inv_11[27] ^ r_10[27] /*3061*/;
  assign sum_11[27] = _2673_ ^ _2672_ /*3060*/;
  assign _2674_ = _2673_ & _2672_ /*3059*/;
  assign _2675_ = inv_11[27] & r_10[27] /*3058*/;
  assign _2676_ = _2674_ | _2675_ /*3057*/;
  assign _2677_ = inv_11[28] ^ r_10[28] /*3055*/;
  assign sum_11[28] = _2677_ ^ _2676_ /*3054*/;
  assign _2678_ = _2677_ & _2676_ /*3053*/;
  assign _2679_ = inv_11[28] & r_10[28] /*3052*/;
  assign _2680_ = _2678_ | _2679_ /*3051*/;
  assign _2681_ = inv_11[29] ^ r_10[29] /*3049*/;
  assign sum_11[29] = _2681_ ^ _2680_ /*3048*/;
  assign _2682_ = _2681_ & _2680_ /*3047*/;
  assign _2683_ = inv_11[29] & r_10[29] /*3046*/;
  assign _2684_ = _2682_ | _2683_ /*3045*/;
  assign _2685_ = inv_11[30] ^ r_10[30] /*3043*/;
  assign sum_11[30] = _2685_ ^ _2684_ /*3042*/;
  assign _2686_ = _2685_ & _2684_ /*3041*/;
  assign _2687_ = inv_11[30] & r_10[30] /*3040*/;
  assign _2688_ = _2686_ | _2687_ /*3039*/;
  assign _2689_ = inv_11[31] ^ r_10[31] /*3037*/;
  assign sum_11[31] = _2689_ ^ _2688_ /*3036*/;
  assign _2690_ = _2689_ & _2688_ /*3035*/;
  assign _2691_ = inv_11[31] & r_10[31] /*3034*/;
  assign _2692_ = _2690_ | _2691_ /*3033*/;
  assign _2693_ = inv_11[32] ^ r_10[32] /*3031*/;
  assign sum_11[32] = _2693_ ^ _2692_ /*3030*/;
  assign _2694_ = _2693_ & _2692_ /*3029*/;
  assign _2695_ = inv_11[32] & r_10[32] /*3028*/;
  assign _2696_ = _2694_ | _2695_ /*3027*/;
  assign _2697_ = inv_11[33] ^ r_10[33] /*3025*/;
  assign sum_11[33] = _2697_ ^ _2696_ /*3024*/;
  assign _2698_ = _2697_ & _2696_ /*3023*/;
  assign _2699_ = inv_11[33] & r_10[33] /*3022*/;
  assign _2700_ = _2698_ | _2699_ /*3021*/;
  assign _2701_ = inv_11[34] ^ r_10[34] /*3019*/;
  assign sum_11[34] = _2701_ ^ _2700_ /*3018*/;
  assign _2702_ = _2701_ & _2700_ /*3017*/;
  assign _2703_ = inv_11[34] & r_10[34] /*3016*/;
  assign _2704_ = _2702_ | _2703_ /*3015*/;
  assign _2705_ = inv_11[35] ^ r_10[35] /*3013*/;
  assign sum_11[35] = _2705_ ^ _2704_ /*3012*/;
  assign _2706_ = _2705_ & _2704_ /*3011*/;
  assign _2707_ = inv_11[35] & r_10[35] /*3010*/;
  assign _2708_ = _2706_ | _2707_ /*3009*/;
  assign _2709_ = inv_11[36] ^ r_10[36] /*3007*/;
  assign sum_11[36] = _2709_ ^ _2708_ /*3006*/;
  assign _2710_ = _2709_ & _2708_ /*3005*/;
  assign _2711_ = inv_11[36] & r_10[36] /*3004*/;
  assign _2712_ = _2710_ | _2711_ /*3003*/;
  assign _2713_ = inv_11[37] ^ r_10[37] /*3001*/;
  assign sum_11[37] = _2713_ ^ _2712_ /*3000*/;
  assign _2714_ = _2713_ & _2712_ /*2999*/;
  assign _2715_ = inv_11[37] & r_10[37] /*2998*/;
  assign _2716_ = _2714_ | _2715_ /*2997*/;
  assign _2717_ = inv_11[38] ^ r_10[38] /*2995*/;
  assign sum_11[38] = _2717_ ^ _2716_ /*2994*/;
  assign _2718_ = _2717_ & _2716_ /*2993*/;
  assign _2719_ = inv_11[38] & r_10[38] /*2992*/;
  assign _2720_ = _2718_ | _2719_ /*2991*/;
  assign _2721_ = inv_11[39] ^ r_10[39] /*2989*/;
  assign sum_11[39] = _2721_ ^ _2720_ /*2988*/;
  assign _2722_ = _2721_ & _2720_ /*2987*/;
  assign _2723_ = inv_11[39] & r_10[39] /*2986*/;
  assign _2724_ = _2722_ | _2723_ /*2985*/;
  assign _2725_ = inv_11[40] ^ r_10[40] /*2983*/;
  assign sum_11[40] = _2725_ ^ _2724_ /*2982*/;
  assign _2726_ = _2725_ & _2724_ /*2981*/;
  assign _2727_ = inv_11[40] & r_10[40] /*2980*/;
  assign _2728_ = _2726_ | _2727_ /*2979*/;
  assign _2729_ = _2728_ ^ _2724_ /*2978*/;
  assign _2730_ = ~_2729_ /*2977*/;
  assign _2731_ = sum_11[40] & _2730_ /*2976*/;
  assign _2732_ = _2729_ & _2728_ /*2975*/;
  assign sum_11[41] = _2732_ | _2731_ /*2974*/;
  assign q[5] = ~sum_11[41] /*2973*/;
  assign m_11[0] = r_10[0] /*2972*/;
  assign m_11[1] = r_10[1] /*2971*/;
  assign m_11[2] = r_10[2] /*2970*/;
  assign m_11[3] = r_10[3] /*2969*/;
  assign m_11[4] = r_10[4] /*2968*/;
  assign m_11[5] = r_10[5] /*2967*/;
  assign m_11[6] = r_10[6] /*2966*/;
  assign m_11[7] = r_10[7] /*2965*/;
  assign m_11[8] = r_10[8] /*2964*/;
  assign m_11[9] = r_10[9] /*2963*/;
  assign m_11[10] = r_10[10] /*2962*/;
  assign m_11[11] = r_10[11] /*2961*/;
  assign m_11[12] = r_10[12] /*2960*/;
  assign m_11[13] = r_10[13] /*2959*/;
  assign m_11[14] = r_10[14] /*2958*/;
  assign m_11[15] = r_10[15] /*2957*/;
  assign m_11[16] = r_10[16] /*2956*/;
  assign m_11[17] = r_10[17] /*2955*/;
  assign m_11[18] = r_10[18] /*2954*/;
  assign m_11[19] = r_10[19] /*2953*/;
  assign m_11[20] = r_10[20] /*2952*/;
  assign m_11[21] = r_10[21] /*2951*/;
  assign m_11[22] = r_10[22] /*2950*/;
  assign m_11[23] = r_10[23] /*2949*/;
  assign m_11[24] = r_10[24] /*2948*/;
  assign m_11[25] = r_10[25] /*2947*/;
  assign m_11[26] = r_10[26] /*2946*/;
  assign m_11[27] = r_10[27] /*2945*/;
  assign m_11[28] = r_10[28] /*2944*/;
  assign m_11[29] = r_10[29] /*2943*/;
  assign m_11[30] = r_10[30] /*2942*/;
  assign m_11[31] = r_10[31] /*2941*/;
  assign m_11[32] = r_10[32] /*2940*/;
  assign m_11[33] = r_10[33] /*2939*/;
  assign m_11[34] = r_10[34] /*2938*/;
  assign m_11[35] = r_10[35] /*2937*/;
  assign m_11[36] = r_10[36] /*2936*/;
  assign m_11[37] = r_10[37] /*2935*/;
  assign m_11[38] = r_10[38] /*2934*/;
  assign m_11[39] = r_10[39] /*2933*/;
  assign m_11[40] = r_10[40] /*2932*/;
  assign m_11[41] = r_10[40] /*2931*/;
  assign _2734_ = ~q[5] /*2930*/;
  assign _2735_ = sum_11[0] & q[5] /*2929*/;
  assign _2736_ = m_11[0] & _2734_ /*2928*/;
  assign r_11[0] = _2736_ | _2735_ /*2927*/;
  assign _2737_ = ~q[5] /*2926*/;
  assign _2738_ = sum_11[1] & q[5] /*2925*/;
  assign _2739_ = m_11[1] & _2737_ /*2924*/;
  assign r_11[1] = _2739_ | _2738_ /*2923*/;
  assign _2740_ = ~q[5] /*2922*/;
  assign _2741_ = sum_11[2] & q[5] /*2921*/;
  assign _2742_ = m_11[2] & _2740_ /*2920*/;
  assign r_11[2] = _2742_ | _2741_ /*2919*/;
  assign _2743_ = ~q[5] /*2918*/;
  assign _2744_ = sum_11[3] & q[5] /*2917*/;
  assign _2745_ = m_11[3] & _2743_ /*2916*/;
  assign r_11[3] = _2745_ | _2744_ /*2915*/;
  assign _2746_ = ~q[5] /*2914*/;
  assign _2747_ = sum_11[4] & q[5] /*2913*/;
  assign _2748_ = m_11[4] & _2746_ /*2912*/;
  assign r_11[4] = _2748_ | _2747_ /*2911*/;
  assign _2749_ = ~q[5] /*2910*/;
  assign _2750_ = sum_11[5] & q[5] /*2909*/;
  assign _2751_ = m_11[5] & _2749_ /*2908*/;
  assign r_11[5] = _2751_ | _2750_ /*2907*/;
  assign _2752_ = ~q[5] /*2906*/;
  assign _2753_ = sum_11[6] & q[5] /*2905*/;
  assign _2754_ = m_11[6] & _2752_ /*2904*/;
  assign r_11[6] = _2754_ | _2753_ /*2903*/;
  assign _2755_ = ~q[5] /*2902*/;
  assign _2756_ = sum_11[7] & q[5] /*2901*/;
  assign _2757_ = m_11[7] & _2755_ /*2900*/;
  assign r_11[7] = _2757_ | _2756_ /*2899*/;
  assign _2758_ = ~q[5] /*2898*/;
  assign _2759_ = sum_11[8] & q[5] /*2897*/;
  assign _2760_ = m_11[8] & _2758_ /*2896*/;
  assign r_11[8] = _2760_ | _2759_ /*2895*/;
  assign _2761_ = ~q[5] /*2894*/;
  assign _2762_ = sum_11[9] & q[5] /*2893*/;
  assign _2763_ = m_11[9] & _2761_ /*2892*/;
  assign r_11[9] = _2763_ | _2762_ /*2891*/;
  assign _2764_ = ~q[5] /*2890*/;
  assign _2765_ = sum_11[10] & q[5] /*2889*/;
  assign _2766_ = m_11[10] & _2764_ /*2888*/;
  assign r_11[10] = _2766_ | _2765_ /*2887*/;
  assign _2767_ = ~q[5] /*2886*/;
  assign _2768_ = sum_11[11] & q[5] /*2885*/;
  assign _2769_ = m_11[11] & _2767_ /*2884*/;
  assign r_11[11] = _2769_ | _2768_ /*2883*/;
  assign _2770_ = ~q[5] /*2882*/;
  assign _2771_ = sum_11[12] & q[5] /*2881*/;
  assign _2772_ = m_11[12] & _2770_ /*2880*/;
  assign r_11[12] = _2772_ | _2771_ /*2879*/;
  assign _2773_ = ~q[5] /*2878*/;
  assign _2774_ = sum_11[13] & q[5] /*2877*/;
  assign _2775_ = m_11[13] & _2773_ /*2876*/;
  assign r_11[13] = _2775_ | _2774_ /*2875*/;
  assign _2776_ = ~q[5] /*2874*/;
  assign _2777_ = sum_11[14] & q[5] /*2873*/;
  assign _2778_ = m_11[14] & _2776_ /*2872*/;
  assign r_11[14] = _2778_ | _2777_ /*2871*/;
  assign _2779_ = ~q[5] /*2870*/;
  assign _2780_ = sum_11[15] & q[5] /*2869*/;
  assign _2781_ = m_11[15] & _2779_ /*2868*/;
  assign r_11[15] = _2781_ | _2780_ /*2867*/;
  assign _2782_ = ~q[5] /*2866*/;
  assign _2783_ = sum_11[16] & q[5] /*2865*/;
  assign _2784_ = m_11[16] & _2782_ /*2864*/;
  assign r_11[16] = _2784_ | _2783_ /*2863*/;
  assign _2785_ = ~q[5] /*2862*/;
  assign _2786_ = sum_11[17] & q[5] /*2861*/;
  assign _2787_ = m_11[17] & _2785_ /*2860*/;
  assign r_11[17] = _2787_ | _2786_ /*2859*/;
  assign _2788_ = ~q[5] /*2858*/;
  assign _2789_ = sum_11[18] & q[5] /*2857*/;
  assign _2790_ = m_11[18] & _2788_ /*2856*/;
  assign r_11[18] = _2790_ | _2789_ /*2855*/;
  assign _2791_ = ~q[5] /*2854*/;
  assign _2792_ = sum_11[19] & q[5] /*2853*/;
  assign _2793_ = m_11[19] & _2791_ /*2852*/;
  assign r_11[19] = _2793_ | _2792_ /*2851*/;
  assign _2794_ = ~q[5] /*2850*/;
  assign _2795_ = sum_11[20] & q[5] /*2849*/;
  assign _2796_ = m_11[20] & _2794_ /*2848*/;
  assign r_11[20] = _2796_ | _2795_ /*2847*/;
  assign _2797_ = ~q[5] /*2846*/;
  assign _2798_ = sum_11[21] & q[5] /*2845*/;
  assign _2799_ = m_11[21] & _2797_ /*2844*/;
  assign r_11[21] = _2799_ | _2798_ /*2843*/;
  assign _2800_ = ~q[5] /*2842*/;
  assign _2801_ = sum_11[22] & q[5] /*2841*/;
  assign _2802_ = m_11[22] & _2800_ /*2840*/;
  assign r_11[22] = _2802_ | _2801_ /*2839*/;
  assign _2803_ = ~q[5] /*2838*/;
  assign _2804_ = sum_11[23] & q[5] /*2837*/;
  assign _2805_ = m_11[23] & _2803_ /*2836*/;
  assign r_11[23] = _2805_ | _2804_ /*2835*/;
  assign _2806_ = ~q[5] /*2834*/;
  assign _2807_ = sum_11[24] & q[5] /*2833*/;
  assign _2808_ = m_11[24] & _2806_ /*2832*/;
  assign r_11[24] = _2808_ | _2807_ /*2831*/;
  assign _2809_ = ~q[5] /*2830*/;
  assign _2810_ = sum_11[25] & q[5] /*2829*/;
  assign _2811_ = m_11[25] & _2809_ /*2828*/;
  assign r_11[25] = _2811_ | _2810_ /*2827*/;
  assign _2812_ = ~q[5] /*2826*/;
  assign _2813_ = sum_11[26] & q[5] /*2825*/;
  assign _2814_ = m_11[26] & _2812_ /*2824*/;
  assign r_11[26] = _2814_ | _2813_ /*2823*/;
  assign _2815_ = ~q[5] /*2822*/;
  assign _2816_ = sum_11[27] & q[5] /*2821*/;
  assign _2817_ = m_11[27] & _2815_ /*2820*/;
  assign r_11[27] = _2817_ | _2816_ /*2819*/;
  assign _2818_ = ~q[5] /*2818*/;
  assign _2819_ = sum_11[28] & q[5] /*2817*/;
  assign _2820_ = m_11[28] & _2818_ /*2816*/;
  assign r_11[28] = _2820_ | _2819_ /*2815*/;
  assign _2821_ = ~q[5] /*2814*/;
  assign _2822_ = sum_11[29] & q[5] /*2813*/;
  assign _2823_ = m_11[29] & _2821_ /*2812*/;
  assign r_11[29] = _2823_ | _2822_ /*2811*/;
  assign _2824_ = ~q[5] /*2810*/;
  assign _2825_ = sum_11[30] & q[5] /*2809*/;
  assign _2826_ = m_11[30] & _2824_ /*2808*/;
  assign r_11[30] = _2826_ | _2825_ /*2807*/;
  assign _2827_ = ~q[5] /*2806*/;
  assign _2828_ = sum_11[31] & q[5] /*2805*/;
  assign _2829_ = m_11[31] & _2827_ /*2804*/;
  assign r_11[31] = _2829_ | _2828_ /*2803*/;
  assign _2830_ = ~q[5] /*2802*/;
  assign _2831_ = sum_11[32] & q[5] /*2801*/;
  assign _2832_ = m_11[32] & _2830_ /*2800*/;
  assign r_11[32] = _2832_ | _2831_ /*2799*/;
  assign _2833_ = ~q[5] /*2798*/;
  assign _2834_ = sum_11[33] & q[5] /*2797*/;
  assign _2835_ = m_11[33] & _2833_ /*2796*/;
  assign r_11[33] = _2835_ | _2834_ /*2795*/;
  assign _2836_ = ~q[5] /*2794*/;
  assign _2837_ = sum_11[34] & q[5] /*2793*/;
  assign _2838_ = m_11[34] & _2836_ /*2792*/;
  assign r_11[34] = _2838_ | _2837_ /*2791*/;
  assign _2839_ = ~q[5] /*2790*/;
  assign _2840_ = sum_11[35] & q[5] /*2789*/;
  assign _2841_ = m_11[35] & _2839_ /*2788*/;
  assign r_11[35] = _2841_ | _2840_ /*2787*/;
  assign _2842_ = ~q[5] /*2786*/;
  assign _2843_ = sum_11[36] & q[5] /*2785*/;
  assign _2844_ = m_11[36] & _2842_ /*2784*/;
  assign r_11[36] = _2844_ | _2843_ /*2783*/;
  assign _2845_ = ~q[5] /*2782*/;
  assign _2846_ = sum_11[37] & q[5] /*2781*/;
  assign _2847_ = m_11[37] & _2845_ /*2780*/;
  assign r_11[37] = _2847_ | _2846_ /*2779*/;
  assign _2848_ = ~q[5] /*2778*/;
  assign _2849_ = sum_11[38] & q[5] /*2777*/;
  assign _2850_ = m_11[38] & _2848_ /*2776*/;
  assign r_11[38] = _2850_ | _2849_ /*2775*/;
  assign _2851_ = ~q[5] /*2774*/;
  assign _2852_ = sum_11[39] & q[5] /*2773*/;
  assign _2853_ = m_11[39] & _2851_ /*2772*/;
  assign r_11[39] = _2853_ | _2852_ /*2771*/;
  assign _2854_ = ~q[5] /*2770*/;
  assign _2855_ = sum_11[40] & q[5] /*2769*/;
  assign _2856_ = m_11[40] & _2854_ /*2768*/;
  assign r_11[40] = _2856_ | _2855_ /*2767*/;
  assign _2857_ = ~q[5] /*2766*/;
  assign _2858_ = sum_11[41] & q[5] /*2765*/;
  assign _2859_ = m_11[41] & _2857_ /*2764*/;
  assign r_11[41] = _2859_ | _2858_ /*2763*/;
  assign inv_12[0] = oneWire /*2692*/;
  assign inv_12[1] = oneWire /*2686*/;
  assign inv_12[2] = oneWire /*2680*/;
  assign inv_12[3] = oneWire /*2674*/;
  assign inv_12[4] = ~div[0] /*2668*/;
  assign inv_12[5] = ~div[1] /*2662*/;
  assign inv_12[6] = ~div[2] /*2656*/;
  assign inv_12[7] = ~div[3] /*2650*/;
  assign inv_12[8] = ~div[4] /*2644*/;
  assign inv_12[9] = ~div[5] /*2638*/;
  assign inv_12[10] = ~div[6] /*2632*/;
  assign inv_12[11] = ~div[7] /*2626*/;
  assign inv_12[12] = ~div[8] /*2620*/;
  assign inv_12[13] = ~div[9] /*2614*/;
  assign inv_12[14] = ~div[10] /*2608*/;
  assign inv_12[15] = ~div[11] /*2602*/;
  assign inv_12[16] = ~div[12] /*2596*/;
  assign inv_12[17] = ~div[13] /*2590*/;
  assign inv_12[18] = ~div[14] /*2584*/;
  assign inv_12[19] = oneWire /*2578*/;
  assign inv_12[20] = oneWire /*2572*/;
  assign inv_12[21] = oneWire /*2566*/;
  assign inv_12[22] = oneWire /*2560*/;
  assign inv_12[23] = oneWire /*2554*/;
  assign inv_12[24] = oneWire /*2548*/;
  assign inv_12[25] = oneWire /*2542*/;
  assign inv_12[26] = oneWire /*2536*/;
  assign inv_12[27] = oneWire /*2530*/;
  assign inv_12[28] = oneWire /*2524*/;
  assign inv_12[29] = oneWire /*2518*/;
  assign inv_12[30] = oneWire /*2512*/;
  assign inv_12[31] = oneWire /*2506*/;
  assign inv_12[32] = oneWire /*2500*/;
  assign inv_12[33] = oneWire /*2494*/;
  assign inv_12[34] = oneWire /*2488*/;
  assign inv_12[35] = oneWire /*2482*/;
  assign inv_12[36] = oneWire /*2476*/;
  assign inv_12[37] = oneWire /*2470*/;
  assign inv_12[38] = oneWire /*2464*/;
  assign inv_12[39] = oneWire /*2458*/;
  assign inv_12[40] = oneWire /*2452*/;
  assign inv_12[41] = oneWire /*2446*/;
  assign _2860_ = inv_12[0] ^ r_11[0] /*2691*/;
  assign sum_12[0] = _2860_ ^ oneWire /*2690*/;
  assign _2861_ = _2860_ & oneWire /*2689*/;
  assign _2862_ = inv_12[0] & r_11[0] /*2688*/;
  assign _2863_ = _2861_ | _2862_ /*2687*/;
  assign _2864_ = inv_12[1] ^ r_11[1] /*2685*/;
  assign sum_12[1] = _2864_ ^ _2863_ /*2684*/;
  assign _2865_ = _2864_ & _2863_ /*2683*/;
  assign _2866_ = inv_12[1] & r_11[1] /*2682*/;
  assign _2867_ = _2865_ | _2866_ /*2681*/;
  assign _2868_ = inv_12[2] ^ r_11[2] /*2679*/;
  assign sum_12[2] = _2868_ ^ _2867_ /*2678*/;
  assign _2869_ = _2868_ & _2867_ /*2677*/;
  assign _2870_ = inv_12[2] & r_11[2] /*2676*/;
  assign _2871_ = _2869_ | _2870_ /*2675*/;
  assign _2872_ = inv_12[3] ^ r_11[3] /*2673*/;
  assign sum_12[3] = _2872_ ^ _2871_ /*2672*/;
  assign _2873_ = _2872_ & _2871_ /*2671*/;
  assign _2874_ = inv_12[3] & r_11[3] /*2670*/;
  assign _2875_ = _2873_ | _2874_ /*2669*/;
  assign _2876_ = inv_12[4] ^ r_11[4] /*2667*/;
  assign sum_12[4] = _2876_ ^ _2875_ /*2666*/;
  assign _2877_ = _2876_ & _2875_ /*2665*/;
  assign _2878_ = inv_12[4] & r_11[4] /*2664*/;
  assign _2879_ = _2877_ | _2878_ /*2663*/;
  assign _2880_ = inv_12[5] ^ r_11[5] /*2661*/;
  assign sum_12[5] = _2880_ ^ _2879_ /*2660*/;
  assign _2881_ = _2880_ & _2879_ /*2659*/;
  assign _2882_ = inv_12[5] & r_11[5] /*2658*/;
  assign _2883_ = _2881_ | _2882_ /*2657*/;
  assign _2884_ = inv_12[6] ^ r_11[6] /*2655*/;
  assign sum_12[6] = _2884_ ^ _2883_ /*2654*/;
  assign _2885_ = _2884_ & _2883_ /*2653*/;
  assign _2886_ = inv_12[6] & r_11[6] /*2652*/;
  assign _2887_ = _2885_ | _2886_ /*2651*/;
  assign _2888_ = inv_12[7] ^ r_11[7] /*2649*/;
  assign sum_12[7] = _2888_ ^ _2887_ /*2648*/;
  assign _2889_ = _2888_ & _2887_ /*2647*/;
  assign _2890_ = inv_12[7] & r_11[7] /*2646*/;
  assign _2891_ = _2889_ | _2890_ /*2645*/;
  assign _2892_ = inv_12[8] ^ r_11[8] /*2643*/;
  assign sum_12[8] = _2892_ ^ _2891_ /*2642*/;
  assign _2893_ = _2892_ & _2891_ /*2641*/;
  assign _2894_ = inv_12[8] & r_11[8] /*2640*/;
  assign _2895_ = _2893_ | _2894_ /*2639*/;
  assign _2896_ = inv_12[9] ^ r_11[9] /*2637*/;
  assign sum_12[9] = _2896_ ^ _2895_ /*2636*/;
  assign _2897_ = _2896_ & _2895_ /*2635*/;
  assign _2898_ = inv_12[9] & r_11[9] /*2634*/;
  assign _2899_ = _2897_ | _2898_ /*2633*/;
  assign _2900_ = inv_12[10] ^ r_11[10] /*2631*/;
  assign sum_12[10] = _2900_ ^ _2899_ /*2630*/;
  assign _2901_ = _2900_ & _2899_ /*2629*/;
  assign _2902_ = inv_12[10] & r_11[10] /*2628*/;
  assign _2903_ = _2901_ | _2902_ /*2627*/;
  assign _2904_ = inv_12[11] ^ r_11[11] /*2625*/;
  assign sum_12[11] = _2904_ ^ _2903_ /*2624*/;
  assign _2905_ = _2904_ & _2903_ /*2623*/;
  assign _2906_ = inv_12[11] & r_11[11] /*2622*/;
  assign _2907_ = _2905_ | _2906_ /*2621*/;
  assign _2908_ = inv_12[12] ^ r_11[12] /*2619*/;
  assign sum_12[12] = _2908_ ^ _2907_ /*2618*/;
  assign _2909_ = _2908_ & _2907_ /*2617*/;
  assign _2910_ = inv_12[12] & r_11[12] /*2616*/;
  assign _2911_ = _2909_ | _2910_ /*2615*/;
  assign _2912_ = inv_12[13] ^ r_11[13] /*2613*/;
  assign sum_12[13] = _2912_ ^ _2911_ /*2612*/;
  assign _2913_ = _2912_ & _2911_ /*2611*/;
  assign _2914_ = inv_12[13] & r_11[13] /*2610*/;
  assign _2915_ = _2913_ | _2914_ /*2609*/;
  assign _2916_ = inv_12[14] ^ r_11[14] /*2607*/;
  assign sum_12[14] = _2916_ ^ _2915_ /*2606*/;
  assign _2917_ = _2916_ & _2915_ /*2605*/;
  assign _2918_ = inv_12[14] & r_11[14] /*2604*/;
  assign _2919_ = _2917_ | _2918_ /*2603*/;
  assign _2920_ = inv_12[15] ^ r_11[15] /*2601*/;
  assign sum_12[15] = _2920_ ^ _2919_ /*2600*/;
  assign _2921_ = _2920_ & _2919_ /*2599*/;
  assign _2922_ = inv_12[15] & r_11[15] /*2598*/;
  assign _2923_ = _2921_ | _2922_ /*2597*/;
  assign _2924_ = inv_12[16] ^ r_11[16] /*2595*/;
  assign sum_12[16] = _2924_ ^ _2923_ /*2594*/;
  assign _2925_ = _2924_ & _2923_ /*2593*/;
  assign _2926_ = inv_12[16] & r_11[16] /*2592*/;
  assign _2927_ = _2925_ | _2926_ /*2591*/;
  assign _2928_ = inv_12[17] ^ r_11[17] /*2589*/;
  assign sum_12[17] = _2928_ ^ _2927_ /*2588*/;
  assign _2929_ = _2928_ & _2927_ /*2587*/;
  assign _2930_ = inv_12[17] & r_11[17] /*2586*/;
  assign _2931_ = _2929_ | _2930_ /*2585*/;
  assign _2932_ = inv_12[18] ^ r_11[18] /*2583*/;
  assign sum_12[18] = _2932_ ^ _2931_ /*2582*/;
  assign _2933_ = _2932_ & _2931_ /*2581*/;
  assign _2934_ = inv_12[18] & r_11[18] /*2580*/;
  assign _2935_ = _2933_ | _2934_ /*2579*/;
  assign _2936_ = inv_12[19] ^ r_11[19] /*2577*/;
  assign sum_12[19] = _2936_ ^ _2935_ /*2576*/;
  assign _2937_ = _2936_ & _2935_ /*2575*/;
  assign _2938_ = inv_12[19] & r_11[19] /*2574*/;
  assign _2939_ = _2937_ | _2938_ /*2573*/;
  assign _2940_ = inv_12[20] ^ r_11[20] /*2571*/;
  assign sum_12[20] = _2940_ ^ _2939_ /*2570*/;
  assign _2941_ = _2940_ & _2939_ /*2569*/;
  assign _2942_ = inv_12[20] & r_11[20] /*2568*/;
  assign _2943_ = _2941_ | _2942_ /*2567*/;
  assign _2944_ = inv_12[21] ^ r_11[21] /*2565*/;
  assign sum_12[21] = _2944_ ^ _2943_ /*2564*/;
  assign _2945_ = _2944_ & _2943_ /*2563*/;
  assign _2946_ = inv_12[21] & r_11[21] /*2562*/;
  assign _2947_ = _2945_ | _2946_ /*2561*/;
  assign _2948_ = inv_12[22] ^ r_11[22] /*2559*/;
  assign sum_12[22] = _2948_ ^ _2947_ /*2558*/;
  assign _2949_ = _2948_ & _2947_ /*2557*/;
  assign _2950_ = inv_12[22] & r_11[22] /*2556*/;
  assign _2951_ = _2949_ | _2950_ /*2555*/;
  assign _2952_ = inv_12[23] ^ r_11[23] /*2553*/;
  assign sum_12[23] = _2952_ ^ _2951_ /*2552*/;
  assign _2953_ = _2952_ & _2951_ /*2551*/;
  assign _2954_ = inv_12[23] & r_11[23] /*2550*/;
  assign _2955_ = _2953_ | _2954_ /*2549*/;
  assign _2956_ = inv_12[24] ^ r_11[24] /*2547*/;
  assign sum_12[24] = _2956_ ^ _2955_ /*2546*/;
  assign _2957_ = _2956_ & _2955_ /*2545*/;
  assign _2958_ = inv_12[24] & r_11[24] /*2544*/;
  assign _2959_ = _2957_ | _2958_ /*2543*/;
  assign _2960_ = inv_12[25] ^ r_11[25] /*2541*/;
  assign sum_12[25] = _2960_ ^ _2959_ /*2540*/;
  assign _2961_ = _2960_ & _2959_ /*2539*/;
  assign _2962_ = inv_12[25] & r_11[25] /*2538*/;
  assign _2963_ = _2961_ | _2962_ /*2537*/;
  assign _2964_ = inv_12[26] ^ r_11[26] /*2535*/;
  assign sum_12[26] = _2964_ ^ _2963_ /*2534*/;
  assign _2965_ = _2964_ & _2963_ /*2533*/;
  assign _2966_ = inv_12[26] & r_11[26] /*2532*/;
  assign _2967_ = _2965_ | _2966_ /*2531*/;
  assign _2968_ = inv_12[27] ^ r_11[27] /*2529*/;
  assign sum_12[27] = _2968_ ^ _2967_ /*2528*/;
  assign _2969_ = _2968_ & _2967_ /*2527*/;
  assign _2970_ = inv_12[27] & r_11[27] /*2526*/;
  assign _2971_ = _2969_ | _2970_ /*2525*/;
  assign _2972_ = inv_12[28] ^ r_11[28] /*2523*/;
  assign sum_12[28] = _2972_ ^ _2971_ /*2522*/;
  assign _2973_ = _2972_ & _2971_ /*2521*/;
  assign _2974_ = inv_12[28] & r_11[28] /*2520*/;
  assign _2975_ = _2973_ | _2974_ /*2519*/;
  assign _2976_ = inv_12[29] ^ r_11[29] /*2517*/;
  assign sum_12[29] = _2976_ ^ _2975_ /*2516*/;
  assign _2977_ = _2976_ & _2975_ /*2515*/;
  assign _2978_ = inv_12[29] & r_11[29] /*2514*/;
  assign _2979_ = _2977_ | _2978_ /*2513*/;
  assign _2980_ = inv_12[30] ^ r_11[30] /*2511*/;
  assign sum_12[30] = _2980_ ^ _2979_ /*2510*/;
  assign _2981_ = _2980_ & _2979_ /*2509*/;
  assign _2982_ = inv_12[30] & r_11[30] /*2508*/;
  assign _2983_ = _2981_ | _2982_ /*2507*/;
  assign _2984_ = inv_12[31] ^ r_11[31] /*2505*/;
  assign sum_12[31] = _2984_ ^ _2983_ /*2504*/;
  assign _2985_ = _2984_ & _2983_ /*2503*/;
  assign _2986_ = inv_12[31] & r_11[31] /*2502*/;
  assign _2987_ = _2985_ | _2986_ /*2501*/;
  assign _2988_ = inv_12[32] ^ r_11[32] /*2499*/;
  assign sum_12[32] = _2988_ ^ _2987_ /*2498*/;
  assign _2989_ = _2988_ & _2987_ /*2497*/;
  assign _2990_ = inv_12[32] & r_11[32] /*2496*/;
  assign _2991_ = _2989_ | _2990_ /*2495*/;
  assign _2992_ = inv_12[33] ^ r_11[33] /*2493*/;
  assign sum_12[33] = _2992_ ^ _2991_ /*2492*/;
  assign _2993_ = _2992_ & _2991_ /*2491*/;
  assign _2994_ = inv_12[33] & r_11[33] /*2490*/;
  assign _2995_ = _2993_ | _2994_ /*2489*/;
  assign _2996_ = inv_12[34] ^ r_11[34] /*2487*/;
  assign sum_12[34] = _2996_ ^ _2995_ /*2486*/;
  assign _2997_ = _2996_ & _2995_ /*2485*/;
  assign _2998_ = inv_12[34] & r_11[34] /*2484*/;
  assign _2999_ = _2997_ | _2998_ /*2483*/;
  assign _3000_ = inv_12[35] ^ r_11[35] /*2481*/;
  assign sum_12[35] = _3000_ ^ _2999_ /*2480*/;
  assign _3001_ = _3000_ & _2999_ /*2479*/;
  assign _3002_ = inv_12[35] & r_11[35] /*2478*/;
  assign _3003_ = _3001_ | _3002_ /*2477*/;
  assign _3004_ = inv_12[36] ^ r_11[36] /*2475*/;
  assign sum_12[36] = _3004_ ^ _3003_ /*2474*/;
  assign _3005_ = _3004_ & _3003_ /*2473*/;
  assign _3006_ = inv_12[36] & r_11[36] /*2472*/;
  assign _3007_ = _3005_ | _3006_ /*2471*/;
  assign _3008_ = inv_12[37] ^ r_11[37] /*2469*/;
  assign sum_12[37] = _3008_ ^ _3007_ /*2468*/;
  assign _3009_ = _3008_ & _3007_ /*2467*/;
  assign _3010_ = inv_12[37] & r_11[37] /*2466*/;
  assign _3011_ = _3009_ | _3010_ /*2465*/;
  assign _3012_ = inv_12[38] ^ r_11[38] /*2463*/;
  assign sum_12[38] = _3012_ ^ _3011_ /*2462*/;
  assign _3013_ = _3012_ & _3011_ /*2461*/;
  assign _3014_ = inv_12[38] & r_11[38] /*2460*/;
  assign _3015_ = _3013_ | _3014_ /*2459*/;
  assign _3016_ = inv_12[39] ^ r_11[39] /*2457*/;
  assign sum_12[39] = _3016_ ^ _3015_ /*2456*/;
  assign _3017_ = _3016_ & _3015_ /*2455*/;
  assign _3018_ = inv_12[39] & r_11[39] /*2454*/;
  assign _3019_ = _3017_ | _3018_ /*2453*/;
  assign _3020_ = inv_12[40] ^ r_11[40] /*2451*/;
  assign sum_12[40] = _3020_ ^ _3019_ /*2450*/;
  assign _3021_ = _3020_ & _3019_ /*2449*/;
  assign _3022_ = inv_12[40] & r_11[40] /*2448*/;
  assign _3023_ = _3021_ | _3022_ /*2447*/;
  assign _3024_ = inv_12[41] ^ r_11[41] /*2445*/;
  assign sum_12[41] = _3024_ ^ _3023_ /*2444*/;
  assign _3025_ = _3024_ & _3023_ /*2443*/;
  assign _3026_ = inv_12[41] & r_11[41] /*2442*/;
  assign _3027_ = _3025_ | _3026_ /*2441*/;
  assign _3028_ = _3027_ ^ _3023_ /*2440*/;
  assign _3029_ = ~_3028_ /*2439*/;
  assign _3030_ = sum_12[41] & _3029_ /*2438*/;
  assign _3031_ = _3028_ & _3027_ /*2437*/;
  assign sum_12[42] = _3031_ | _3030_ /*2436*/;
  assign q[4] = ~sum_12[42] /*2435*/;
  assign m_12[0] = r_11[0] /*2434*/;
  assign m_12[1] = r_11[1] /*2433*/;
  assign m_12[2] = r_11[2] /*2432*/;
  assign m_12[3] = r_11[3] /*2431*/;
  assign m_12[4] = r_11[4] /*2430*/;
  assign m_12[5] = r_11[5] /*2429*/;
  assign m_12[6] = r_11[6] /*2428*/;
  assign m_12[7] = r_11[7] /*2427*/;
  assign m_12[8] = r_11[8] /*2426*/;
  assign m_12[9] = r_11[9] /*2425*/;
  assign m_12[10] = r_11[10] /*2424*/;
  assign m_12[11] = r_11[11] /*2423*/;
  assign m_12[12] = r_11[12] /*2422*/;
  assign m_12[13] = r_11[13] /*2421*/;
  assign m_12[14] = r_11[14] /*2420*/;
  assign m_12[15] = r_11[15] /*2419*/;
  assign m_12[16] = r_11[16] /*2418*/;
  assign m_12[17] = r_11[17] /*2417*/;
  assign m_12[18] = r_11[18] /*2416*/;
  assign m_12[19] = r_11[19] /*2415*/;
  assign m_12[20] = r_11[20] /*2414*/;
  assign m_12[21] = r_11[21] /*2413*/;
  assign m_12[22] = r_11[22] /*2412*/;
  assign m_12[23] = r_11[23] /*2411*/;
  assign m_12[24] = r_11[24] /*2410*/;
  assign m_12[25] = r_11[25] /*2409*/;
  assign m_12[26] = r_11[26] /*2408*/;
  assign m_12[27] = r_11[27] /*2407*/;
  assign m_12[28] = r_11[28] /*2406*/;
  assign m_12[29] = r_11[29] /*2405*/;
  assign m_12[30] = r_11[30] /*2404*/;
  assign m_12[31] = r_11[31] /*2403*/;
  assign m_12[32] = r_11[32] /*2402*/;
  assign m_12[33] = r_11[33] /*2401*/;
  assign m_12[34] = r_11[34] /*2400*/;
  assign m_12[35] = r_11[35] /*2399*/;
  assign m_12[36] = r_11[36] /*2398*/;
  assign m_12[37] = r_11[37] /*2397*/;
  assign m_12[38] = r_11[38] /*2396*/;
  assign m_12[39] = r_11[39] /*2395*/;
  assign m_12[40] = r_11[40] /*2394*/;
  assign m_12[41] = r_11[41] /*2393*/;
  assign m_12[42] = r_11[41] /*2392*/;
  assign _3033_ = ~q[4] /*2391*/;
  assign _3034_ = sum_12[0] & q[4] /*2390*/;
  assign _3035_ = m_12[0] & _3033_ /*2389*/;
  assign r_12[0] = _3035_ | _3034_ /*2388*/;
  assign _3036_ = ~q[4] /*2387*/;
  assign _3037_ = sum_12[1] & q[4] /*2386*/;
  assign _3038_ = m_12[1] & _3036_ /*2385*/;
  assign r_12[1] = _3038_ | _3037_ /*2384*/;
  assign _3039_ = ~q[4] /*2383*/;
  assign _3040_ = sum_12[2] & q[4] /*2382*/;
  assign _3041_ = m_12[2] & _3039_ /*2381*/;
  assign r_12[2] = _3041_ | _3040_ /*2380*/;
  assign _3042_ = ~q[4] /*2379*/;
  assign _3043_ = sum_12[3] & q[4] /*2378*/;
  assign _3044_ = m_12[3] & _3042_ /*2377*/;
  assign r_12[3] = _3044_ | _3043_ /*2376*/;
  assign _3045_ = ~q[4] /*2375*/;
  assign _3046_ = sum_12[4] & q[4] /*2374*/;
  assign _3047_ = m_12[4] & _3045_ /*2373*/;
  assign r_12[4] = _3047_ | _3046_ /*2372*/;
  assign _3048_ = ~q[4] /*2371*/;
  assign _3049_ = sum_12[5] & q[4] /*2370*/;
  assign _3050_ = m_12[5] & _3048_ /*2369*/;
  assign r_12[5] = _3050_ | _3049_ /*2368*/;
  assign _3051_ = ~q[4] /*2367*/;
  assign _3052_ = sum_12[6] & q[4] /*2366*/;
  assign _3053_ = m_12[6] & _3051_ /*2365*/;
  assign r_12[6] = _3053_ | _3052_ /*2364*/;
  assign _3054_ = ~q[4] /*2363*/;
  assign _3055_ = sum_12[7] & q[4] /*2362*/;
  assign _3056_ = m_12[7] & _3054_ /*2361*/;
  assign r_12[7] = _3056_ | _3055_ /*2360*/;
  assign _3057_ = ~q[4] /*2359*/;
  assign _3058_ = sum_12[8] & q[4] /*2358*/;
  assign _3059_ = m_12[8] & _3057_ /*2357*/;
  assign r_12[8] = _3059_ | _3058_ /*2356*/;
  assign _3060_ = ~q[4] /*2355*/;
  assign _3061_ = sum_12[9] & q[4] /*2354*/;
  assign _3062_ = m_12[9] & _3060_ /*2353*/;
  assign r_12[9] = _3062_ | _3061_ /*2352*/;
  assign _3063_ = ~q[4] /*2351*/;
  assign _3064_ = sum_12[10] & q[4] /*2350*/;
  assign _3065_ = m_12[10] & _3063_ /*2349*/;
  assign r_12[10] = _3065_ | _3064_ /*2348*/;
  assign _3066_ = ~q[4] /*2347*/;
  assign _3067_ = sum_12[11] & q[4] /*2346*/;
  assign _3068_ = m_12[11] & _3066_ /*2345*/;
  assign r_12[11] = _3068_ | _3067_ /*2344*/;
  assign _3069_ = ~q[4] /*2343*/;
  assign _3070_ = sum_12[12] & q[4] /*2342*/;
  assign _3071_ = m_12[12] & _3069_ /*2341*/;
  assign r_12[12] = _3071_ | _3070_ /*2340*/;
  assign _3072_ = ~q[4] /*2339*/;
  assign _3073_ = sum_12[13] & q[4] /*2338*/;
  assign _3074_ = m_12[13] & _3072_ /*2337*/;
  assign r_12[13] = _3074_ | _3073_ /*2336*/;
  assign _3075_ = ~q[4] /*2335*/;
  assign _3076_ = sum_12[14] & q[4] /*2334*/;
  assign _3077_ = m_12[14] & _3075_ /*2333*/;
  assign r_12[14] = _3077_ | _3076_ /*2332*/;
  assign _3078_ = ~q[4] /*2331*/;
  assign _3079_ = sum_12[15] & q[4] /*2330*/;
  assign _3080_ = m_12[15] & _3078_ /*2329*/;
  assign r_12[15] = _3080_ | _3079_ /*2328*/;
  assign _3081_ = ~q[4] /*2327*/;
  assign _3082_ = sum_12[16] & q[4] /*2326*/;
  assign _3083_ = m_12[16] & _3081_ /*2325*/;
  assign r_12[16] = _3083_ | _3082_ /*2324*/;
  assign _3084_ = ~q[4] /*2323*/;
  assign _3085_ = sum_12[17] & q[4] /*2322*/;
  assign _3086_ = m_12[17] & _3084_ /*2321*/;
  assign r_12[17] = _3086_ | _3085_ /*2320*/;
  assign _3087_ = ~q[4] /*2319*/;
  assign _3088_ = sum_12[18] & q[4] /*2318*/;
  assign _3089_ = m_12[18] & _3087_ /*2317*/;
  assign r_12[18] = _3089_ | _3088_ /*2316*/;
  assign _3090_ = ~q[4] /*2315*/;
  assign _3091_ = sum_12[19] & q[4] /*2314*/;
  assign _3092_ = m_12[19] & _3090_ /*2313*/;
  assign r_12[19] = _3092_ | _3091_ /*2312*/;
  assign _3093_ = ~q[4] /*2311*/;
  assign _3094_ = sum_12[20] & q[4] /*2310*/;
  assign _3095_ = m_12[20] & _3093_ /*2309*/;
  assign r_12[20] = _3095_ | _3094_ /*2308*/;
  assign _3096_ = ~q[4] /*2307*/;
  assign _3097_ = sum_12[21] & q[4] /*2306*/;
  assign _3098_ = m_12[21] & _3096_ /*2305*/;
  assign r_12[21] = _3098_ | _3097_ /*2304*/;
  assign _3099_ = ~q[4] /*2303*/;
  assign _3100_ = sum_12[22] & q[4] /*2302*/;
  assign _3101_ = m_12[22] & _3099_ /*2301*/;
  assign r_12[22] = _3101_ | _3100_ /*2300*/;
  assign _3102_ = ~q[4] /*2299*/;
  assign _3103_ = sum_12[23] & q[4] /*2298*/;
  assign _3104_ = m_12[23] & _3102_ /*2297*/;
  assign r_12[23] = _3104_ | _3103_ /*2296*/;
  assign _3105_ = ~q[4] /*2295*/;
  assign _3106_ = sum_12[24] & q[4] /*2294*/;
  assign _3107_ = m_12[24] & _3105_ /*2293*/;
  assign r_12[24] = _3107_ | _3106_ /*2292*/;
  assign _3108_ = ~q[4] /*2291*/;
  assign _3109_ = sum_12[25] & q[4] /*2290*/;
  assign _3110_ = m_12[25] & _3108_ /*2289*/;
  assign r_12[25] = _3110_ | _3109_ /*2288*/;
  assign _3111_ = ~q[4] /*2287*/;
  assign _3112_ = sum_12[26] & q[4] /*2286*/;
  assign _3113_ = m_12[26] & _3111_ /*2285*/;
  assign r_12[26] = _3113_ | _3112_ /*2284*/;
  assign _3114_ = ~q[4] /*2283*/;
  assign _3115_ = sum_12[27] & q[4] /*2282*/;
  assign _3116_ = m_12[27] & _3114_ /*2281*/;
  assign r_12[27] = _3116_ | _3115_ /*2280*/;
  assign _3117_ = ~q[4] /*2279*/;
  assign _3118_ = sum_12[28] & q[4] /*2278*/;
  assign _3119_ = m_12[28] & _3117_ /*2277*/;
  assign r_12[28] = _3119_ | _3118_ /*2276*/;
  assign _3120_ = ~q[4] /*2275*/;
  assign _3121_ = sum_12[29] & q[4] /*2274*/;
  assign _3122_ = m_12[29] & _3120_ /*2273*/;
  assign r_12[29] = _3122_ | _3121_ /*2272*/;
  assign _3123_ = ~q[4] /*2271*/;
  assign _3124_ = sum_12[30] & q[4] /*2270*/;
  assign _3125_ = m_12[30] & _3123_ /*2269*/;
  assign r_12[30] = _3125_ | _3124_ /*2268*/;
  assign _3126_ = ~q[4] /*2267*/;
  assign _3127_ = sum_12[31] & q[4] /*2266*/;
  assign _3128_ = m_12[31] & _3126_ /*2265*/;
  assign r_12[31] = _3128_ | _3127_ /*2264*/;
  assign _3129_ = ~q[4] /*2263*/;
  assign _3130_ = sum_12[32] & q[4] /*2262*/;
  assign _3131_ = m_12[32] & _3129_ /*2261*/;
  assign r_12[32] = _3131_ | _3130_ /*2260*/;
  assign _3132_ = ~q[4] /*2259*/;
  assign _3133_ = sum_12[33] & q[4] /*2258*/;
  assign _3134_ = m_12[33] & _3132_ /*2257*/;
  assign r_12[33] = _3134_ | _3133_ /*2256*/;
  assign _3135_ = ~q[4] /*2255*/;
  assign _3136_ = sum_12[34] & q[4] /*2254*/;
  assign _3137_ = m_12[34] & _3135_ /*2253*/;
  assign r_12[34] = _3137_ | _3136_ /*2252*/;
  assign _3138_ = ~q[4] /*2251*/;
  assign _3139_ = sum_12[35] & q[4] /*2250*/;
  assign _3140_ = m_12[35] & _3138_ /*2249*/;
  assign r_12[35] = _3140_ | _3139_ /*2248*/;
  assign _3141_ = ~q[4] /*2247*/;
  assign _3142_ = sum_12[36] & q[4] /*2246*/;
  assign _3143_ = m_12[36] & _3141_ /*2245*/;
  assign r_12[36] = _3143_ | _3142_ /*2244*/;
  assign _3144_ = ~q[4] /*2243*/;
  assign _3145_ = sum_12[37] & q[4] /*2242*/;
  assign _3146_ = m_12[37] & _3144_ /*2241*/;
  assign r_12[37] = _3146_ | _3145_ /*2240*/;
  assign _3147_ = ~q[4] /*2239*/;
  assign _3148_ = sum_12[38] & q[4] /*2238*/;
  assign _3149_ = m_12[38] & _3147_ /*2237*/;
  assign r_12[38] = _3149_ | _3148_ /*2236*/;
  assign _3150_ = ~q[4] /*2235*/;
  assign _3151_ = sum_12[39] & q[4] /*2234*/;
  assign _3152_ = m_12[39] & _3150_ /*2233*/;
  assign r_12[39] = _3152_ | _3151_ /*2232*/;
  assign _3153_ = ~q[4] /*2231*/;
  assign _3154_ = sum_12[40] & q[4] /*2230*/;
  assign _3155_ = m_12[40] & _3153_ /*2229*/;
  assign r_12[40] = _3155_ | _3154_ /*2228*/;
  assign _3156_ = ~q[4] /*2227*/;
  assign _3157_ = sum_12[41] & q[4] /*2226*/;
  assign _3158_ = m_12[41] & _3156_ /*2225*/;
  assign r_12[41] = _3158_ | _3157_ /*2224*/;
  assign _3159_ = ~q[4] /*2223*/;
  assign _3160_ = sum_12[42] & q[4] /*2222*/;
  assign _3161_ = m_12[42] & _3159_ /*2221*/;
  assign r_12[42] = _3161_ | _3160_ /*2220*/;
  assign inv_13[0] = oneWire /*2160*/;
  assign inv_13[1] = oneWire /*2154*/;
  assign inv_13[2] = oneWire /*2148*/;
  assign inv_13[3] = ~div[0] /*2142*/;
  assign inv_13[4] = ~div[1] /*2136*/;
  assign inv_13[5] = ~div[2] /*2130*/;
  assign inv_13[6] = ~div[3] /*2124*/;
  assign inv_13[7] = ~div[4] /*2118*/;
  assign inv_13[8] = ~div[5] /*2112*/;
  assign inv_13[9] = ~div[6] /*2106*/;
  assign inv_13[10] = ~div[7] /*2100*/;
  assign inv_13[11] = ~div[8] /*2094*/;
  assign inv_13[12] = ~div[9] /*2088*/;
  assign inv_13[13] = ~div[10] /*2082*/;
  assign inv_13[14] = ~div[11] /*2076*/;
  assign inv_13[15] = ~div[12] /*2070*/;
  assign inv_13[16] = ~div[13] /*2064*/;
  assign inv_13[17] = ~div[14] /*2058*/;
  assign inv_13[18] = oneWire /*2052*/;
  assign inv_13[19] = oneWire /*2046*/;
  assign inv_13[20] = oneWire /*2040*/;
  assign inv_13[21] = oneWire /*2034*/;
  assign inv_13[22] = oneWire /*2028*/;
  assign inv_13[23] = oneWire /*2022*/;
  assign inv_13[24] = oneWire /*2016*/;
  assign inv_13[25] = oneWire /*2010*/;
  assign inv_13[26] = oneWire /*2004*/;
  assign inv_13[27] = oneWire /*1998*/;
  assign inv_13[28] = oneWire /*1992*/;
  assign inv_13[29] = oneWire /*1986*/;
  assign inv_13[30] = oneWire /*1980*/;
  assign inv_13[31] = oneWire /*1974*/;
  assign inv_13[32] = oneWire /*1968*/;
  assign inv_13[33] = oneWire /*1962*/;
  assign inv_13[34] = oneWire /*1956*/;
  assign inv_13[35] = oneWire /*1950*/;
  assign inv_13[36] = oneWire /*1944*/;
  assign inv_13[37] = oneWire /*1938*/;
  assign inv_13[38] = oneWire /*1932*/;
  assign inv_13[39] = oneWire /*1926*/;
  assign inv_13[40] = oneWire /*1920*/;
  assign inv_13[41] = oneWire /*1914*/;
  assign inv_13[42] = oneWire /*1908*/;
  assign _3162_ = inv_13[0] ^ r_12[0] /*2159*/;
  assign sum_13[0] = _3162_ ^ oneWire /*2158*/;
  assign _3163_ = _3162_ & oneWire /*2157*/;
  assign _3164_ = inv_13[0] & r_12[0] /*2156*/;
  assign _3165_ = _3163_ | _3164_ /*2155*/;
  assign _3166_ = inv_13[1] ^ r_12[1] /*2153*/;
  assign sum_13[1] = _3166_ ^ _3165_ /*2152*/;
  assign _3167_ = _3166_ & _3165_ /*2151*/;
  assign _3168_ = inv_13[1] & r_12[1] /*2150*/;
  assign _3169_ = _3167_ | _3168_ /*2149*/;
  assign _3170_ = inv_13[2] ^ r_12[2] /*2147*/;
  assign sum_13[2] = _3170_ ^ _3169_ /*2146*/;
  assign _3171_ = _3170_ & _3169_ /*2145*/;
  assign _3172_ = inv_13[2] & r_12[2] /*2144*/;
  assign _3173_ = _3171_ | _3172_ /*2143*/;
  assign _3174_ = inv_13[3] ^ r_12[3] /*2141*/;
  assign sum_13[3] = _3174_ ^ _3173_ /*2140*/;
  assign _3175_ = _3174_ & _3173_ /*2139*/;
  assign _3176_ = inv_13[3] & r_12[3] /*2138*/;
  assign _3177_ = _3175_ | _3176_ /*2137*/;
  assign _3178_ = inv_13[4] ^ r_12[4] /*2135*/;
  assign sum_13[4] = _3178_ ^ _3177_ /*2134*/;
  assign _3179_ = _3178_ & _3177_ /*2133*/;
  assign _3180_ = inv_13[4] & r_12[4] /*2132*/;
  assign _3181_ = _3179_ | _3180_ /*2131*/;
  assign _3182_ = inv_13[5] ^ r_12[5] /*2129*/;
  assign sum_13[5] = _3182_ ^ _3181_ /*2128*/;
  assign _3183_ = _3182_ & _3181_ /*2127*/;
  assign _3184_ = inv_13[5] & r_12[5] /*2126*/;
  assign _3185_ = _3183_ | _3184_ /*2125*/;
  assign _3186_ = inv_13[6] ^ r_12[6] /*2123*/;
  assign sum_13[6] = _3186_ ^ _3185_ /*2122*/;
  assign _3187_ = _3186_ & _3185_ /*2121*/;
  assign _3188_ = inv_13[6] & r_12[6] /*2120*/;
  assign _3189_ = _3187_ | _3188_ /*2119*/;
  assign _3190_ = inv_13[7] ^ r_12[7] /*2117*/;
  assign sum_13[7] = _3190_ ^ _3189_ /*2116*/;
  assign _3191_ = _3190_ & _3189_ /*2115*/;
  assign _3192_ = inv_13[7] & r_12[7] /*2114*/;
  assign _3193_ = _3191_ | _3192_ /*2113*/;
  assign _3194_ = inv_13[8] ^ r_12[8] /*2111*/;
  assign sum_13[8] = _3194_ ^ _3193_ /*2110*/;
  assign _3195_ = _3194_ & _3193_ /*2109*/;
  assign _3196_ = inv_13[8] & r_12[8] /*2108*/;
  assign _3197_ = _3195_ | _3196_ /*2107*/;
  assign _3198_ = inv_13[9] ^ r_12[9] /*2105*/;
  assign sum_13[9] = _3198_ ^ _3197_ /*2104*/;
  assign _3199_ = _3198_ & _3197_ /*2103*/;
  assign _3200_ = inv_13[9] & r_12[9] /*2102*/;
  assign _3201_ = _3199_ | _3200_ /*2101*/;
  assign _3202_ = inv_13[10] ^ r_12[10] /*2099*/;
  assign sum_13[10] = _3202_ ^ _3201_ /*2098*/;
  assign _3203_ = _3202_ & _3201_ /*2097*/;
  assign _3204_ = inv_13[10] & r_12[10] /*2096*/;
  assign _3205_ = _3203_ | _3204_ /*2095*/;
  assign _3206_ = inv_13[11] ^ r_12[11] /*2093*/;
  assign sum_13[11] = _3206_ ^ _3205_ /*2092*/;
  assign _3207_ = _3206_ & _3205_ /*2091*/;
  assign _3208_ = inv_13[11] & r_12[11] /*2090*/;
  assign _3209_ = _3207_ | _3208_ /*2089*/;
  assign _3210_ = inv_13[12] ^ r_12[12] /*2087*/;
  assign sum_13[12] = _3210_ ^ _3209_ /*2086*/;
  assign _3211_ = _3210_ & _3209_ /*2085*/;
  assign _3212_ = inv_13[12] & r_12[12] /*2084*/;
  assign _3213_ = _3211_ | _3212_ /*2083*/;
  assign _3214_ = inv_13[13] ^ r_12[13] /*2081*/;
  assign sum_13[13] = _3214_ ^ _3213_ /*2080*/;
  assign _3215_ = _3214_ & _3213_ /*2079*/;
  assign _3216_ = inv_13[13] & r_12[13] /*2078*/;
  assign _3217_ = _3215_ | _3216_ /*2077*/;
  assign _3218_ = inv_13[14] ^ r_12[14] /*2075*/;
  assign sum_13[14] = _3218_ ^ _3217_ /*2074*/;
  assign _3219_ = _3218_ & _3217_ /*2073*/;
  assign _3220_ = inv_13[14] & r_12[14] /*2072*/;
  assign _3221_ = _3219_ | _3220_ /*2071*/;
  assign _3222_ = inv_13[15] ^ r_12[15] /*2069*/;
  assign sum_13[15] = _3222_ ^ _3221_ /*2068*/;
  assign _3223_ = _3222_ & _3221_ /*2067*/;
  assign _3224_ = inv_13[15] & r_12[15] /*2066*/;
  assign _3225_ = _3223_ | _3224_ /*2065*/;
  assign _3226_ = inv_13[16] ^ r_12[16] /*2063*/;
  assign sum_13[16] = _3226_ ^ _3225_ /*2062*/;
  assign _3227_ = _3226_ & _3225_ /*2061*/;
  assign _3228_ = inv_13[16] & r_12[16] /*2060*/;
  assign _3229_ = _3227_ | _3228_ /*2059*/;
  assign _3230_ = inv_13[17] ^ r_12[17] /*2057*/;
  assign sum_13[17] = _3230_ ^ _3229_ /*2056*/;
  assign _3231_ = _3230_ & _3229_ /*2055*/;
  assign _3232_ = inv_13[17] & r_12[17] /*2054*/;
  assign _3233_ = _3231_ | _3232_ /*2053*/;
  assign _3234_ = inv_13[18] ^ r_12[18] /*2051*/;
  assign sum_13[18] = _3234_ ^ _3233_ /*2050*/;
  assign _3235_ = _3234_ & _3233_ /*2049*/;
  assign _3236_ = inv_13[18] & r_12[18] /*2048*/;
  assign _3237_ = _3235_ | _3236_ /*2047*/;
  assign _3238_ = inv_13[19] ^ r_12[19] /*2045*/;
  assign sum_13[19] = _3238_ ^ _3237_ /*2044*/;
  assign _3239_ = _3238_ & _3237_ /*2043*/;
  assign _3240_ = inv_13[19] & r_12[19] /*2042*/;
  assign _3241_ = _3239_ | _3240_ /*2041*/;
  assign _3242_ = inv_13[20] ^ r_12[20] /*2039*/;
  assign sum_13[20] = _3242_ ^ _3241_ /*2038*/;
  assign _3243_ = _3242_ & _3241_ /*2037*/;
  assign _3244_ = inv_13[20] & r_12[20] /*2036*/;
  assign _3245_ = _3243_ | _3244_ /*2035*/;
  assign _3246_ = inv_13[21] ^ r_12[21] /*2033*/;
  assign sum_13[21] = _3246_ ^ _3245_ /*2032*/;
  assign _3247_ = _3246_ & _3245_ /*2031*/;
  assign _3248_ = inv_13[21] & r_12[21] /*2030*/;
  assign _3249_ = _3247_ | _3248_ /*2029*/;
  assign _3250_ = inv_13[22] ^ r_12[22] /*2027*/;
  assign sum_13[22] = _3250_ ^ _3249_ /*2026*/;
  assign _3251_ = _3250_ & _3249_ /*2025*/;
  assign _3252_ = inv_13[22] & r_12[22] /*2024*/;
  assign _3253_ = _3251_ | _3252_ /*2023*/;
  assign _3254_ = inv_13[23] ^ r_12[23] /*2021*/;
  assign sum_13[23] = _3254_ ^ _3253_ /*2020*/;
  assign _3255_ = _3254_ & _3253_ /*2019*/;
  assign _3256_ = inv_13[23] & r_12[23] /*2018*/;
  assign _3257_ = _3255_ | _3256_ /*2017*/;
  assign _3258_ = inv_13[24] ^ r_12[24] /*2015*/;
  assign sum_13[24] = _3258_ ^ _3257_ /*2014*/;
  assign _3259_ = _3258_ & _3257_ /*2013*/;
  assign _3260_ = inv_13[24] & r_12[24] /*2012*/;
  assign _3261_ = _3259_ | _3260_ /*2011*/;
  assign _3262_ = inv_13[25] ^ r_12[25] /*2009*/;
  assign sum_13[25] = _3262_ ^ _3261_ /*2008*/;
  assign _3263_ = _3262_ & _3261_ /*2007*/;
  assign _3264_ = inv_13[25] & r_12[25] /*2006*/;
  assign _3265_ = _3263_ | _3264_ /*2005*/;
  assign _3266_ = inv_13[26] ^ r_12[26] /*2003*/;
  assign sum_13[26] = _3266_ ^ _3265_ /*2002*/;
  assign _3267_ = _3266_ & _3265_ /*2001*/;
  assign _3268_ = inv_13[26] & r_12[26] /*2000*/;
  assign _3269_ = _3267_ | _3268_ /*1999*/;
  assign _3270_ = inv_13[27] ^ r_12[27] /*1997*/;
  assign sum_13[27] = _3270_ ^ _3269_ /*1996*/;
  assign _3271_ = _3270_ & _3269_ /*1995*/;
  assign _3272_ = inv_13[27] & r_12[27] /*1994*/;
  assign _3273_ = _3271_ | _3272_ /*1993*/;
  assign _3274_ = inv_13[28] ^ r_12[28] /*1991*/;
  assign sum_13[28] = _3274_ ^ _3273_ /*1990*/;
  assign _3275_ = _3274_ & _3273_ /*1989*/;
  assign _3276_ = inv_13[28] & r_12[28] /*1988*/;
  assign _3277_ = _3275_ | _3276_ /*1987*/;
  assign _3278_ = inv_13[29] ^ r_12[29] /*1985*/;
  assign sum_13[29] = _3278_ ^ _3277_ /*1984*/;
  assign _3279_ = _3278_ & _3277_ /*1983*/;
  assign _3280_ = inv_13[29] & r_12[29] /*1982*/;
  assign _3281_ = _3279_ | _3280_ /*1981*/;
  assign _3282_ = inv_13[30] ^ r_12[30] /*1979*/;
  assign sum_13[30] = _3282_ ^ _3281_ /*1978*/;
  assign _3283_ = _3282_ & _3281_ /*1977*/;
  assign _3284_ = inv_13[30] & r_12[30] /*1976*/;
  assign _3285_ = _3283_ | _3284_ /*1975*/;
  assign _3286_ = inv_13[31] ^ r_12[31] /*1973*/;
  assign sum_13[31] = _3286_ ^ _3285_ /*1972*/;
  assign _3287_ = _3286_ & _3285_ /*1971*/;
  assign _3288_ = inv_13[31] & r_12[31] /*1970*/;
  assign _3289_ = _3287_ | _3288_ /*1969*/;
  assign _3290_ = inv_13[32] ^ r_12[32] /*1967*/;
  assign sum_13[32] = _3290_ ^ _3289_ /*1966*/;
  assign _3291_ = _3290_ & _3289_ /*1965*/;
  assign _3292_ = inv_13[32] & r_12[32] /*1964*/;
  assign _3293_ = _3291_ | _3292_ /*1963*/;
  assign _3294_ = inv_13[33] ^ r_12[33] /*1961*/;
  assign sum_13[33] = _3294_ ^ _3293_ /*1960*/;
  assign _3295_ = _3294_ & _3293_ /*1959*/;
  assign _3296_ = inv_13[33] & r_12[33] /*1958*/;
  assign _3297_ = _3295_ | _3296_ /*1957*/;
  assign _3298_ = inv_13[34] ^ r_12[34] /*1955*/;
  assign sum_13[34] = _3298_ ^ _3297_ /*1954*/;
  assign _3299_ = _3298_ & _3297_ /*1953*/;
  assign _3300_ = inv_13[34] & r_12[34] /*1952*/;
  assign _3301_ = _3299_ | _3300_ /*1951*/;
  assign _3302_ = inv_13[35] ^ r_12[35] /*1949*/;
  assign sum_13[35] = _3302_ ^ _3301_ /*1948*/;
  assign _3303_ = _3302_ & _3301_ /*1947*/;
  assign _3304_ = inv_13[35] & r_12[35] /*1946*/;
  assign _3305_ = _3303_ | _3304_ /*1945*/;
  assign _3306_ = inv_13[36] ^ r_12[36] /*1943*/;
  assign sum_13[36] = _3306_ ^ _3305_ /*1942*/;
  assign _3307_ = _3306_ & _3305_ /*1941*/;
  assign _3308_ = inv_13[36] & r_12[36] /*1940*/;
  assign _3309_ = _3307_ | _3308_ /*1939*/;
  assign _3310_ = inv_13[37] ^ r_12[37] /*1937*/;
  assign sum_13[37] = _3310_ ^ _3309_ /*1936*/;
  assign _3311_ = _3310_ & _3309_ /*1935*/;
  assign _3312_ = inv_13[37] & r_12[37] /*1934*/;
  assign _3313_ = _3311_ | _3312_ /*1933*/;
  assign _3314_ = inv_13[38] ^ r_12[38] /*1931*/;
  assign sum_13[38] = _3314_ ^ _3313_ /*1930*/;
  assign _3315_ = _3314_ & _3313_ /*1929*/;
  assign _3316_ = inv_13[38] & r_12[38] /*1928*/;
  assign _3317_ = _3315_ | _3316_ /*1927*/;
  assign _3318_ = inv_13[39] ^ r_12[39] /*1925*/;
  assign sum_13[39] = _3318_ ^ _3317_ /*1924*/;
  assign _3319_ = _3318_ & _3317_ /*1923*/;
  assign _3320_ = inv_13[39] & r_12[39] /*1922*/;
  assign _3321_ = _3319_ | _3320_ /*1921*/;
  assign _3322_ = inv_13[40] ^ r_12[40] /*1919*/;
  assign sum_13[40] = _3322_ ^ _3321_ /*1918*/;
  assign _3323_ = _3322_ & _3321_ /*1917*/;
  assign _3324_ = inv_13[40] & r_12[40] /*1916*/;
  assign _3325_ = _3323_ | _3324_ /*1915*/;
  assign _3326_ = inv_13[41] ^ r_12[41] /*1913*/;
  assign sum_13[41] = _3326_ ^ _3325_ /*1912*/;
  assign _3327_ = _3326_ & _3325_ /*1911*/;
  assign _3328_ = inv_13[41] & r_12[41] /*1910*/;
  assign _3329_ = _3327_ | _3328_ /*1909*/;
  assign _3330_ = inv_13[42] ^ r_12[42] /*1907*/;
  assign sum_13[42] = _3330_ ^ _3329_ /*1906*/;
  assign _3331_ = _3330_ & _3329_ /*1905*/;
  assign _3332_ = inv_13[42] & r_12[42] /*1904*/;
  assign _3333_ = _3331_ | _3332_ /*1903*/;
  assign _3334_ = _3333_ ^ _3329_ /*1902*/;
  assign _3335_ = ~_3334_ /*1901*/;
  assign _3336_ = sum_13[42] & _3335_ /*1900*/;
  assign _3337_ = _3334_ & _3333_ /*1899*/;
  assign sum_13[43] = _3337_ | _3336_ /*1898*/;
  assign q[3] = ~sum_13[43] /*1897*/;
  assign m_13[0] = r_12[0] /*1896*/;
  assign m_13[1] = r_12[1] /*1895*/;
  assign m_13[2] = r_12[2] /*1894*/;
  assign m_13[3] = r_12[3] /*1893*/;
  assign m_13[4] = r_12[4] /*1892*/;
  assign m_13[5] = r_12[5] /*1891*/;
  assign m_13[6] = r_12[6] /*1890*/;
  assign m_13[7] = r_12[7] /*1889*/;
  assign m_13[8] = r_12[8] /*1888*/;
  assign m_13[9] = r_12[9] /*1887*/;
  assign m_13[10] = r_12[10] /*1886*/;
  assign m_13[11] = r_12[11] /*1885*/;
  assign m_13[12] = r_12[12] /*1884*/;
  assign m_13[13] = r_12[13] /*1883*/;
  assign m_13[14] = r_12[14] /*1882*/;
  assign m_13[15] = r_12[15] /*1881*/;
  assign m_13[16] = r_12[16] /*1880*/;
  assign m_13[17] = r_12[17] /*1879*/;
  assign m_13[18] = r_12[18] /*1878*/;
  assign m_13[19] = r_12[19] /*1877*/;
  assign m_13[20] = r_12[20] /*1876*/;
  assign m_13[21] = r_12[21] /*1875*/;
  assign m_13[22] = r_12[22] /*1874*/;
  assign m_13[23] = r_12[23] /*1873*/;
  assign m_13[24] = r_12[24] /*1872*/;
  assign m_13[25] = r_12[25] /*1871*/;
  assign m_13[26] = r_12[26] /*1870*/;
  assign m_13[27] = r_12[27] /*1869*/;
  assign m_13[28] = r_12[28] /*1868*/;
  assign m_13[29] = r_12[29] /*1867*/;
  assign m_13[30] = r_12[30] /*1866*/;
  assign m_13[31] = r_12[31] /*1865*/;
  assign m_13[32] = r_12[32] /*1864*/;
  assign m_13[33] = r_12[33] /*1863*/;
  assign m_13[34] = r_12[34] /*1862*/;
  assign m_13[35] = r_12[35] /*1861*/;
  assign m_13[36] = r_12[36] /*1860*/;
  assign m_13[37] = r_12[37] /*1859*/;
  assign m_13[38] = r_12[38] /*1858*/;
  assign m_13[39] = r_12[39] /*1857*/;
  assign m_13[40] = r_12[40] /*1856*/;
  assign m_13[41] = r_12[41] /*1855*/;
  assign m_13[42] = r_12[42] /*1854*/;
  assign m_13[43] = r_12[42] /*1853*/;
  assign _3339_ = ~q[3] /*1852*/;
  assign _3340_ = sum_13[0] & q[3] /*1851*/;
  assign _3341_ = m_13[0] & _3339_ /*1850*/;
  assign r_13[0] = _3341_ | _3340_ /*1849*/;
  assign _3342_ = ~q[3] /*1848*/;
  assign _3343_ = sum_13[1] & q[3] /*1847*/;
  assign _3344_ = m_13[1] & _3342_ /*1846*/;
  assign r_13[1] = _3344_ | _3343_ /*1845*/;
  assign _3345_ = ~q[3] /*1844*/;
  assign _3346_ = sum_13[2] & q[3] /*1843*/;
  assign _3347_ = m_13[2] & _3345_ /*1842*/;
  assign r_13[2] = _3347_ | _3346_ /*1841*/;
  assign _3348_ = ~q[3] /*1840*/;
  assign _3349_ = sum_13[3] & q[3] /*1839*/;
  assign _3350_ = m_13[3] & _3348_ /*1838*/;
  assign r_13[3] = _3350_ | _3349_ /*1837*/;
  assign _3351_ = ~q[3] /*1836*/;
  assign _3352_ = sum_13[4] & q[3] /*1835*/;
  assign _3353_ = m_13[4] & _3351_ /*1834*/;
  assign r_13[4] = _3353_ | _3352_ /*1833*/;
  assign _3354_ = ~q[3] /*1832*/;
  assign _3355_ = sum_13[5] & q[3] /*1831*/;
  assign _3356_ = m_13[5] & _3354_ /*1830*/;
  assign r_13[5] = _3356_ | _3355_ /*1829*/;
  assign _3357_ = ~q[3] /*1828*/;
  assign _3358_ = sum_13[6] & q[3] /*1827*/;
  assign _3359_ = m_13[6] & _3357_ /*1826*/;
  assign r_13[6] = _3359_ | _3358_ /*1825*/;
  assign _3360_ = ~q[3] /*1824*/;
  assign _3361_ = sum_13[7] & q[3] /*1823*/;
  assign _3362_ = m_13[7] & _3360_ /*1822*/;
  assign r_13[7] = _3362_ | _3361_ /*1821*/;
  assign _3363_ = ~q[3] /*1820*/;
  assign _3364_ = sum_13[8] & q[3] /*1819*/;
  assign _3365_ = m_13[8] & _3363_ /*1818*/;
  assign r_13[8] = _3365_ | _3364_ /*1817*/;
  assign _3366_ = ~q[3] /*1816*/;
  assign _3367_ = sum_13[9] & q[3] /*1815*/;
  assign _3368_ = m_13[9] & _3366_ /*1814*/;
  assign r_13[9] = _3368_ | _3367_ /*1813*/;
  assign _3369_ = ~q[3] /*1812*/;
  assign _3370_ = sum_13[10] & q[3] /*1811*/;
  assign _3371_ = m_13[10] & _3369_ /*1810*/;
  assign r_13[10] = _3371_ | _3370_ /*1809*/;
  assign _3372_ = ~q[3] /*1808*/;
  assign _3373_ = sum_13[11] & q[3] /*1807*/;
  assign _3374_ = m_13[11] & _3372_ /*1806*/;
  assign r_13[11] = _3374_ | _3373_ /*1805*/;
  assign _3375_ = ~q[3] /*1804*/;
  assign _3376_ = sum_13[12] & q[3] /*1803*/;
  assign _3377_ = m_13[12] & _3375_ /*1802*/;
  assign r_13[12] = _3377_ | _3376_ /*1801*/;
  assign _3378_ = ~q[3] /*1800*/;
  assign _3379_ = sum_13[13] & q[3] /*1799*/;
  assign _3380_ = m_13[13] & _3378_ /*1798*/;
  assign r_13[13] = _3380_ | _3379_ /*1797*/;
  assign _3381_ = ~q[3] /*1796*/;
  assign _3382_ = sum_13[14] & q[3] /*1795*/;
  assign _3383_ = m_13[14] & _3381_ /*1794*/;
  assign r_13[14] = _3383_ | _3382_ /*1793*/;
  assign _3384_ = ~q[3] /*1792*/;
  assign _3385_ = sum_13[15] & q[3] /*1791*/;
  assign _3386_ = m_13[15] & _3384_ /*1790*/;
  assign r_13[15] = _3386_ | _3385_ /*1789*/;
  assign _3387_ = ~q[3] /*1788*/;
  assign _3388_ = sum_13[16] & q[3] /*1787*/;
  assign _3389_ = m_13[16] & _3387_ /*1786*/;
  assign r_13[16] = _3389_ | _3388_ /*1785*/;
  assign _3390_ = ~q[3] /*1784*/;
  assign _3391_ = sum_13[17] & q[3] /*1783*/;
  assign _3392_ = m_13[17] & _3390_ /*1782*/;
  assign r_13[17] = _3392_ | _3391_ /*1781*/;
  assign _3393_ = ~q[3] /*1780*/;
  assign _3394_ = sum_13[18] & q[3] /*1779*/;
  assign _3395_ = m_13[18] & _3393_ /*1778*/;
  assign r_13[18] = _3395_ | _3394_ /*1777*/;
  assign _3396_ = ~q[3] /*1776*/;
  assign _3397_ = sum_13[19] & q[3] /*1775*/;
  assign _3398_ = m_13[19] & _3396_ /*1774*/;
  assign r_13[19] = _3398_ | _3397_ /*1773*/;
  assign _3399_ = ~q[3] /*1772*/;
  assign _3400_ = sum_13[20] & q[3] /*1771*/;
  assign _3401_ = m_13[20] & _3399_ /*1770*/;
  assign r_13[20] = _3401_ | _3400_ /*1769*/;
  assign _3402_ = ~q[3] /*1768*/;
  assign _3403_ = sum_13[21] & q[3] /*1767*/;
  assign _3404_ = m_13[21] & _3402_ /*1766*/;
  assign r_13[21] = _3404_ | _3403_ /*1765*/;
  assign _3405_ = ~q[3] /*1764*/;
  assign _3406_ = sum_13[22] & q[3] /*1763*/;
  assign _3407_ = m_13[22] & _3405_ /*1762*/;
  assign r_13[22] = _3407_ | _3406_ /*1761*/;
  assign _3408_ = ~q[3] /*1760*/;
  assign _3409_ = sum_13[23] & q[3] /*1759*/;
  assign _3410_ = m_13[23] & _3408_ /*1758*/;
  assign r_13[23] = _3410_ | _3409_ /*1757*/;
  assign _3411_ = ~q[3] /*1756*/;
  assign _3412_ = sum_13[24] & q[3] /*1755*/;
  assign _3413_ = m_13[24] & _3411_ /*1754*/;
  assign r_13[24] = _3413_ | _3412_ /*1753*/;
  assign _3414_ = ~q[3] /*1752*/;
  assign _3415_ = sum_13[25] & q[3] /*1751*/;
  assign _3416_ = m_13[25] & _3414_ /*1750*/;
  assign r_13[25] = _3416_ | _3415_ /*1749*/;
  assign _3417_ = ~q[3] /*1748*/;
  assign _3418_ = sum_13[26] & q[3] /*1747*/;
  assign _3419_ = m_13[26] & _3417_ /*1746*/;
  assign r_13[26] = _3419_ | _3418_ /*1745*/;
  assign _3420_ = ~q[3] /*1744*/;
  assign _3421_ = sum_13[27] & q[3] /*1743*/;
  assign _3422_ = m_13[27] & _3420_ /*1742*/;
  assign r_13[27] = _3422_ | _3421_ /*1741*/;
  assign _3423_ = ~q[3] /*1740*/;
  assign _3424_ = sum_13[28] & q[3] /*1739*/;
  assign _3425_ = m_13[28] & _3423_ /*1738*/;
  assign r_13[28] = _3425_ | _3424_ /*1737*/;
  assign _3426_ = ~q[3] /*1736*/;
  assign _3427_ = sum_13[29] & q[3] /*1735*/;
  assign _3428_ = m_13[29] & _3426_ /*1734*/;
  assign r_13[29] = _3428_ | _3427_ /*1733*/;
  assign _3429_ = ~q[3] /*1732*/;
  assign _3430_ = sum_13[30] & q[3] /*1731*/;
  assign _3431_ = m_13[30] & _3429_ /*1730*/;
  assign r_13[30] = _3431_ | _3430_ /*1729*/;
  assign _3432_ = ~q[3] /*1728*/;
  assign _3433_ = sum_13[31] & q[3] /*1727*/;
  assign _3434_ = m_13[31] & _3432_ /*1726*/;
  assign r_13[31] = _3434_ | _3433_ /*1725*/;
  assign _3435_ = ~q[3] /*1724*/;
  assign _3436_ = sum_13[32] & q[3] /*1723*/;
  assign _3437_ = m_13[32] & _3435_ /*1722*/;
  assign r_13[32] = _3437_ | _3436_ /*1721*/;
  assign _3438_ = ~q[3] /*1720*/;
  assign _3439_ = sum_13[33] & q[3] /*1719*/;
  assign _3440_ = m_13[33] & _3438_ /*1718*/;
  assign r_13[33] = _3440_ | _3439_ /*1717*/;
  assign _3441_ = ~q[3] /*1716*/;
  assign _3442_ = sum_13[34] & q[3] /*1715*/;
  assign _3443_ = m_13[34] & _3441_ /*1714*/;
  assign r_13[34] = _3443_ | _3442_ /*1713*/;
  assign _3444_ = ~q[3] /*1712*/;
  assign _3445_ = sum_13[35] & q[3] /*1711*/;
  assign _3446_ = m_13[35] & _3444_ /*1710*/;
  assign r_13[35] = _3446_ | _3445_ /*1709*/;
  assign _3447_ = ~q[3] /*1708*/;
  assign _3448_ = sum_13[36] & q[3] /*1707*/;
  assign _3449_ = m_13[36] & _3447_ /*1706*/;
  assign r_13[36] = _3449_ | _3448_ /*1705*/;
  assign _3450_ = ~q[3] /*1704*/;
  assign _3451_ = sum_13[37] & q[3] /*1703*/;
  assign _3452_ = m_13[37] & _3450_ /*1702*/;
  assign r_13[37] = _3452_ | _3451_ /*1701*/;
  assign _3453_ = ~q[3] /*1700*/;
  assign _3454_ = sum_13[38] & q[3] /*1699*/;
  assign _3455_ = m_13[38] & _3453_ /*1698*/;
  assign r_13[38] = _3455_ | _3454_ /*1697*/;
  assign _3456_ = ~q[3] /*1696*/;
  assign _3457_ = sum_13[39] & q[3] /*1695*/;
  assign _3458_ = m_13[39] & _3456_ /*1694*/;
  assign r_13[39] = _3458_ | _3457_ /*1693*/;
  assign _3459_ = ~q[3] /*1692*/;
  assign _3460_ = sum_13[40] & q[3] /*1691*/;
  assign _3461_ = m_13[40] & _3459_ /*1690*/;
  assign r_13[40] = _3461_ | _3460_ /*1689*/;
  assign _3462_ = ~q[3] /*1688*/;
  assign _3463_ = sum_13[41] & q[3] /*1687*/;
  assign _3464_ = m_13[41] & _3462_ /*1686*/;
  assign r_13[41] = _3464_ | _3463_ /*1685*/;
  assign _3465_ = ~q[3] /*1684*/;
  assign _3466_ = sum_13[42] & q[3] /*1683*/;
  assign _3467_ = m_13[42] & _3465_ /*1682*/;
  assign r_13[42] = _3467_ | _3466_ /*1681*/;
  assign _3468_ = ~q[3] /*1680*/;
  assign _3469_ = sum_13[43] & q[3] /*1679*/;
  assign _3470_ = m_13[43] & _3468_ /*1678*/;
  assign r_13[43] = _3470_ | _3469_ /*1677*/;
  assign inv_14[0] = oneWire /*1628*/;
  assign inv_14[1] = oneWire /*1622*/;
  assign inv_14[2] = ~div[0] /*1616*/;
  assign inv_14[3] = ~div[1] /*1610*/;
  assign inv_14[4] = ~div[2] /*1604*/;
  assign inv_14[5] = ~div[3] /*1598*/;
  assign inv_14[6] = ~div[4] /*1592*/;
  assign inv_14[7] = ~div[5] /*1586*/;
  assign inv_14[8] = ~div[6] /*1580*/;
  assign inv_14[9] = ~div[7] /*1574*/;
  assign inv_14[10] = ~div[8] /*1568*/;
  assign inv_14[11] = ~div[9] /*1562*/;
  assign inv_14[12] = ~div[10] /*1556*/;
  assign inv_14[13] = ~div[11] /*1550*/;
  assign inv_14[14] = ~div[12] /*1544*/;
  assign inv_14[15] = ~div[13] /*1538*/;
  assign inv_14[16] = ~div[14] /*1532*/;
  assign inv_14[17] = oneWire /*1526*/;
  assign inv_14[18] = oneWire /*1520*/;
  assign inv_14[19] = oneWire /*1514*/;
  assign inv_14[20] = oneWire /*1508*/;
  assign inv_14[21] = oneWire /*1502*/;
  assign inv_14[22] = oneWire /*1496*/;
  assign inv_14[23] = oneWire /*1490*/;
  assign inv_14[24] = oneWire /*1484*/;
  assign inv_14[25] = oneWire /*1478*/;
  assign inv_14[26] = oneWire /*1472*/;
  assign inv_14[27] = oneWire /*1466*/;
  assign inv_14[28] = oneWire /*1460*/;
  assign inv_14[29] = oneWire /*1454*/;
  assign inv_14[30] = oneWire /*1448*/;
  assign inv_14[31] = oneWire /*1442*/;
  assign inv_14[32] = oneWire /*1436*/;
  assign inv_14[33] = oneWire /*1430*/;
  assign inv_14[34] = oneWire /*1424*/;
  assign inv_14[35] = oneWire /*1418*/;
  assign inv_14[36] = oneWire /*1412*/;
  assign inv_14[37] = oneWire /*1406*/;
  assign inv_14[38] = oneWire /*1400*/;
  assign inv_14[39] = oneWire /*1394*/;
  assign inv_14[40] = oneWire /*1388*/;
  assign inv_14[41] = oneWire /*1382*/;
  assign inv_14[42] = oneWire /*1376*/;
  assign inv_14[43] = oneWire /*1370*/;
  assign _3471_ = inv_14[0] ^ r_13[0] /*1627*/;
  assign sum_14[0] = _3471_ ^ oneWire /*1626*/;
  assign _3472_ = _3471_ & oneWire /*1625*/;
  assign _3473_ = inv_14[0] & r_13[0] /*1624*/;
  assign _3474_ = _3472_ | _3473_ /*1623*/;
  assign _3475_ = inv_14[1] ^ r_13[1] /*1621*/;
  assign sum_14[1] = _3475_ ^ _3474_ /*1620*/;
  assign _3476_ = _3475_ & _3474_ /*1619*/;
  assign _3477_ = inv_14[1] & r_13[1] /*1618*/;
  assign _3478_ = _3476_ | _3477_ /*1617*/;
  assign _3479_ = inv_14[2] ^ r_13[2] /*1615*/;
  assign sum_14[2] = _3479_ ^ _3478_ /*1614*/;
  assign _3480_ = _3479_ & _3478_ /*1613*/;
  assign _3481_ = inv_14[2] & r_13[2] /*1612*/;
  assign _3482_ = _3480_ | _3481_ /*1611*/;
  assign _3483_ = inv_14[3] ^ r_13[3] /*1609*/;
  assign sum_14[3] = _3483_ ^ _3482_ /*1608*/;
  assign _3484_ = _3483_ & _3482_ /*1607*/;
  assign _3485_ = inv_14[3] & r_13[3] /*1606*/;
  assign _3486_ = _3484_ | _3485_ /*1605*/;
  assign _3487_ = inv_14[4] ^ r_13[4] /*1603*/;
  assign sum_14[4] = _3487_ ^ _3486_ /*1602*/;
  assign _3488_ = _3487_ & _3486_ /*1601*/;
  assign _3489_ = inv_14[4] & r_13[4] /*1600*/;
  assign _3490_ = _3488_ | _3489_ /*1599*/;
  assign _3491_ = inv_14[5] ^ r_13[5] /*1597*/;
  assign sum_14[5] = _3491_ ^ _3490_ /*1596*/;
  assign _3492_ = _3491_ & _3490_ /*1595*/;
  assign _3493_ = inv_14[5] & r_13[5] /*1594*/;
  assign _3494_ = _3492_ | _3493_ /*1593*/;
  assign _3495_ = inv_14[6] ^ r_13[6] /*1591*/;
  assign sum_14[6] = _3495_ ^ _3494_ /*1590*/;
  assign _3496_ = _3495_ & _3494_ /*1589*/;
  assign _3497_ = inv_14[6] & r_13[6] /*1588*/;
  assign _3498_ = _3496_ | _3497_ /*1587*/;
  assign _3499_ = inv_14[7] ^ r_13[7] /*1585*/;
  assign sum_14[7] = _3499_ ^ _3498_ /*1584*/;
  assign _3500_ = _3499_ & _3498_ /*1583*/;
  assign _3501_ = inv_14[7] & r_13[7] /*1582*/;
  assign _3502_ = _3500_ | _3501_ /*1581*/;
  assign _3503_ = inv_14[8] ^ r_13[8] /*1579*/;
  assign sum_14[8] = _3503_ ^ _3502_ /*1578*/;
  assign _3504_ = _3503_ & _3502_ /*1577*/;
  assign _3505_ = inv_14[8] & r_13[8] /*1576*/;
  assign _3506_ = _3504_ | _3505_ /*1575*/;
  assign _3507_ = inv_14[9] ^ r_13[9] /*1573*/;
  assign sum_14[9] = _3507_ ^ _3506_ /*1572*/;
  assign _3508_ = _3507_ & _3506_ /*1571*/;
  assign _3509_ = inv_14[9] & r_13[9] /*1570*/;
  assign _3510_ = _3508_ | _3509_ /*1569*/;
  assign _3511_ = inv_14[10] ^ r_13[10] /*1567*/;
  assign sum_14[10] = _3511_ ^ _3510_ /*1566*/;
  assign _3512_ = _3511_ & _3510_ /*1565*/;
  assign _3513_ = inv_14[10] & r_13[10] /*1564*/;
  assign _3514_ = _3512_ | _3513_ /*1563*/;
  assign _3515_ = inv_14[11] ^ r_13[11] /*1561*/;
  assign sum_14[11] = _3515_ ^ _3514_ /*1560*/;
  assign _3516_ = _3515_ & _3514_ /*1559*/;
  assign _3517_ = inv_14[11] & r_13[11] /*1558*/;
  assign _3518_ = _3516_ | _3517_ /*1557*/;
  assign _3519_ = inv_14[12] ^ r_13[12] /*1555*/;
  assign sum_14[12] = _3519_ ^ _3518_ /*1554*/;
  assign _3520_ = _3519_ & _3518_ /*1553*/;
  assign _3521_ = inv_14[12] & r_13[12] /*1552*/;
  assign _3522_ = _3520_ | _3521_ /*1551*/;
  assign _3523_ = inv_14[13] ^ r_13[13] /*1549*/;
  assign sum_14[13] = _3523_ ^ _3522_ /*1548*/;
  assign _3524_ = _3523_ & _3522_ /*1547*/;
  assign _3525_ = inv_14[13] & r_13[13] /*1546*/;
  assign _3526_ = _3524_ | _3525_ /*1545*/;
  assign _3527_ = inv_14[14] ^ r_13[14] /*1543*/;
  assign sum_14[14] = _3527_ ^ _3526_ /*1542*/;
  assign _3528_ = _3527_ & _3526_ /*1541*/;
  assign _3529_ = inv_14[14] & r_13[14] /*1540*/;
  assign _3530_ = _3528_ | _3529_ /*1539*/;
  assign _3531_ = inv_14[15] ^ r_13[15] /*1537*/;
  assign sum_14[15] = _3531_ ^ _3530_ /*1536*/;
  assign _3532_ = _3531_ & _3530_ /*1535*/;
  assign _3533_ = inv_14[15] & r_13[15] /*1534*/;
  assign _3534_ = _3532_ | _3533_ /*1533*/;
  assign _3535_ = inv_14[16] ^ r_13[16] /*1531*/;
  assign sum_14[16] = _3535_ ^ _3534_ /*1530*/;
  assign _3536_ = _3535_ & _3534_ /*1529*/;
  assign _3537_ = inv_14[16] & r_13[16] /*1528*/;
  assign _3538_ = _3536_ | _3537_ /*1527*/;
  assign _3539_ = inv_14[17] ^ r_13[17] /*1525*/;
  assign sum_14[17] = _3539_ ^ _3538_ /*1524*/;
  assign _3540_ = _3539_ & _3538_ /*1523*/;
  assign _3541_ = inv_14[17] & r_13[17] /*1522*/;
  assign _3542_ = _3540_ | _3541_ /*1521*/;
  assign _3543_ = inv_14[18] ^ r_13[18] /*1519*/;
  assign sum_14[18] = _3543_ ^ _3542_ /*1518*/;
  assign _3544_ = _3543_ & _3542_ /*1517*/;
  assign _3545_ = inv_14[18] & r_13[18] /*1516*/;
  assign _3546_ = _3544_ | _3545_ /*1515*/;
  assign _3547_ = inv_14[19] ^ r_13[19] /*1513*/;
  assign sum_14[19] = _3547_ ^ _3546_ /*1512*/;
  assign _3548_ = _3547_ & _3546_ /*1511*/;
  assign _3549_ = inv_14[19] & r_13[19] /*1510*/;
  assign _3550_ = _3548_ | _3549_ /*1509*/;
  assign _3551_ = inv_14[20] ^ r_13[20] /*1507*/;
  assign sum_14[20] = _3551_ ^ _3550_ /*1506*/;
  assign _3552_ = _3551_ & _3550_ /*1505*/;
  assign _3553_ = inv_14[20] & r_13[20] /*1504*/;
  assign _3554_ = _3552_ | _3553_ /*1503*/;
  assign _3555_ = inv_14[21] ^ r_13[21] /*1501*/;
  assign sum_14[21] = _3555_ ^ _3554_ /*1500*/;
  assign _3556_ = _3555_ & _3554_ /*1499*/;
  assign _3557_ = inv_14[21] & r_13[21] /*1498*/;
  assign _3558_ = _3556_ | _3557_ /*1497*/;
  assign _3559_ = inv_14[22] ^ r_13[22] /*1495*/;
  assign sum_14[22] = _3559_ ^ _3558_ /*1494*/;
  assign _3560_ = _3559_ & _3558_ /*1493*/;
  assign _3561_ = inv_14[22] & r_13[22] /*1492*/;
  assign _3562_ = _3560_ | _3561_ /*1491*/;
  assign _3563_ = inv_14[23] ^ r_13[23] /*1489*/;
  assign sum_14[23] = _3563_ ^ _3562_ /*1488*/;
  assign _3564_ = _3563_ & _3562_ /*1487*/;
  assign _3565_ = inv_14[23] & r_13[23] /*1486*/;
  assign _3566_ = _3564_ | _3565_ /*1485*/;
  assign _3567_ = inv_14[24] ^ r_13[24] /*1483*/;
  assign sum_14[24] = _3567_ ^ _3566_ /*1482*/;
  assign _3568_ = _3567_ & _3566_ /*1481*/;
  assign _3569_ = inv_14[24] & r_13[24] /*1480*/;
  assign _3570_ = _3568_ | _3569_ /*1479*/;
  assign _3571_ = inv_14[25] ^ r_13[25] /*1477*/;
  assign sum_14[25] = _3571_ ^ _3570_ /*1476*/;
  assign _3572_ = _3571_ & _3570_ /*1475*/;
  assign _3573_ = inv_14[25] & r_13[25] /*1474*/;
  assign _3574_ = _3572_ | _3573_ /*1473*/;
  assign _3575_ = inv_14[26] ^ r_13[26] /*1471*/;
  assign sum_14[26] = _3575_ ^ _3574_ /*1470*/;
  assign _3576_ = _3575_ & _3574_ /*1469*/;
  assign _3577_ = inv_14[26] & r_13[26] /*1468*/;
  assign _3578_ = _3576_ | _3577_ /*1467*/;
  assign _3579_ = inv_14[27] ^ r_13[27] /*1465*/;
  assign sum_14[27] = _3579_ ^ _3578_ /*1464*/;
  assign _3580_ = _3579_ & _3578_ /*1463*/;
  assign _3581_ = inv_14[27] & r_13[27] /*1462*/;
  assign _3582_ = _3580_ | _3581_ /*1461*/;
  assign _3583_ = inv_14[28] ^ r_13[28] /*1459*/;
  assign sum_14[28] = _3583_ ^ _3582_ /*1458*/;
  assign _3584_ = _3583_ & _3582_ /*1457*/;
  assign _3585_ = inv_14[28] & r_13[28] /*1456*/;
  assign _3586_ = _3584_ | _3585_ /*1455*/;
  assign _3587_ = inv_14[29] ^ r_13[29] /*1453*/;
  assign sum_14[29] = _3587_ ^ _3586_ /*1452*/;
  assign _3588_ = _3587_ & _3586_ /*1451*/;
  assign _3589_ = inv_14[29] & r_13[29] /*1450*/;
  assign _3590_ = _3588_ | _3589_ /*1449*/;
  assign _3591_ = inv_14[30] ^ r_13[30] /*1447*/;
  assign sum_14[30] = _3591_ ^ _3590_ /*1446*/;
  assign _3592_ = _3591_ & _3590_ /*1445*/;
  assign _3593_ = inv_14[30] & r_13[30] /*1444*/;
  assign _3594_ = _3592_ | _3593_ /*1443*/;
  assign _3595_ = inv_14[31] ^ r_13[31] /*1441*/;
  assign sum_14[31] = _3595_ ^ _3594_ /*1440*/;
  assign _3596_ = _3595_ & _3594_ /*1439*/;
  assign _3597_ = inv_14[31] & r_13[31] /*1438*/;
  assign _3598_ = _3596_ | _3597_ /*1437*/;
  assign _3599_ = inv_14[32] ^ r_13[32] /*1435*/;
  assign sum_14[32] = _3599_ ^ _3598_ /*1434*/;
  assign _3600_ = _3599_ & _3598_ /*1433*/;
  assign _3601_ = inv_14[32] & r_13[32] /*1432*/;
  assign _3602_ = _3600_ | _3601_ /*1431*/;
  assign _3603_ = inv_14[33] ^ r_13[33] /*1429*/;
  assign sum_14[33] = _3603_ ^ _3602_ /*1428*/;
  assign _3604_ = _3603_ & _3602_ /*1427*/;
  assign _3605_ = inv_14[33] & r_13[33] /*1426*/;
  assign _3606_ = _3604_ | _3605_ /*1425*/;
  assign _3607_ = inv_14[34] ^ r_13[34] /*1423*/;
  assign sum_14[34] = _3607_ ^ _3606_ /*1422*/;
  assign _3608_ = _3607_ & _3606_ /*1421*/;
  assign _3609_ = inv_14[34] & r_13[34] /*1420*/;
  assign _3610_ = _3608_ | _3609_ /*1419*/;
  assign _3611_ = inv_14[35] ^ r_13[35] /*1417*/;
  assign sum_14[35] = _3611_ ^ _3610_ /*1416*/;
  assign _3612_ = _3611_ & _3610_ /*1415*/;
  assign _3613_ = inv_14[35] & r_13[35] /*1414*/;
  assign _3614_ = _3612_ | _3613_ /*1413*/;
  assign _3615_ = inv_14[36] ^ r_13[36] /*1411*/;
  assign sum_14[36] = _3615_ ^ _3614_ /*1410*/;
  assign _3616_ = _3615_ & _3614_ /*1409*/;
  assign _3617_ = inv_14[36] & r_13[36] /*1408*/;
  assign _3618_ = _3616_ | _3617_ /*1407*/;
  assign _3619_ = inv_14[37] ^ r_13[37] /*1405*/;
  assign sum_14[37] = _3619_ ^ _3618_ /*1404*/;
  assign _3620_ = _3619_ & _3618_ /*1403*/;
  assign _3621_ = inv_14[37] & r_13[37] /*1402*/;
  assign _3622_ = _3620_ | _3621_ /*1401*/;
  assign _3623_ = inv_14[38] ^ r_13[38] /*1399*/;
  assign sum_14[38] = _3623_ ^ _3622_ /*1398*/;
  assign _3624_ = _3623_ & _3622_ /*1397*/;
  assign _3625_ = inv_14[38] & r_13[38] /*1396*/;
  assign _3626_ = _3624_ | _3625_ /*1395*/;
  assign _3627_ = inv_14[39] ^ r_13[39] /*1393*/;
  assign sum_14[39] = _3627_ ^ _3626_ /*1392*/;
  assign _3628_ = _3627_ & _3626_ /*1391*/;
  assign _3629_ = inv_14[39] & r_13[39] /*1390*/;
  assign _3630_ = _3628_ | _3629_ /*1389*/;
  assign _3631_ = inv_14[40] ^ r_13[40] /*1387*/;
  assign sum_14[40] = _3631_ ^ _3630_ /*1386*/;
  assign _3632_ = _3631_ & _3630_ /*1385*/;
  assign _3633_ = inv_14[40] & r_13[40] /*1384*/;
  assign _3634_ = _3632_ | _3633_ /*1383*/;
  assign _3635_ = inv_14[41] ^ r_13[41] /*1381*/;
  assign sum_14[41] = _3635_ ^ _3634_ /*1380*/;
  assign _3636_ = _3635_ & _3634_ /*1379*/;
  assign _3637_ = inv_14[41] & r_13[41] /*1378*/;
  assign _3638_ = _3636_ | _3637_ /*1377*/;
  assign _3639_ = inv_14[42] ^ r_13[42] /*1375*/;
  assign sum_14[42] = _3639_ ^ _3638_ /*1374*/;
  assign _3640_ = _3639_ & _3638_ /*1373*/;
  assign _3641_ = inv_14[42] & r_13[42] /*1372*/;
  assign _3642_ = _3640_ | _3641_ /*1371*/;
  assign _3643_ = inv_14[43] ^ r_13[43] /*1369*/;
  assign sum_14[43] = _3643_ ^ _3642_ /*1368*/;
  assign _3644_ = _3643_ & _3642_ /*1367*/;
  assign _3645_ = inv_14[43] & r_13[43] /*1366*/;
  assign _3646_ = _3644_ | _3645_ /*1365*/;
  assign _3647_ = _3646_ ^ _3642_ /*1364*/;
  assign _3648_ = ~_3647_ /*1363*/;
  assign _3649_ = sum_14[43] & _3648_ /*1362*/;
  assign _3650_ = _3647_ & _3646_ /*1361*/;
  assign sum_14[44] = _3650_ | _3649_ /*1360*/;
  assign q[2] = ~sum_14[44] /*1359*/;
  assign m_14[0] = r_13[0] /*1358*/;
  assign m_14[1] = r_13[1] /*1357*/;
  assign m_14[2] = r_13[2] /*1356*/;
  assign m_14[3] = r_13[3] /*1355*/;
  assign m_14[4] = r_13[4] /*1354*/;
  assign m_14[5] = r_13[5] /*1353*/;
  assign m_14[6] = r_13[6] /*1352*/;
  assign m_14[7] = r_13[7] /*1351*/;
  assign m_14[8] = r_13[8] /*1350*/;
  assign m_14[9] = r_13[9] /*1349*/;
  assign m_14[10] = r_13[10] /*1348*/;
  assign m_14[11] = r_13[11] /*1347*/;
  assign m_14[12] = r_13[12] /*1346*/;
  assign m_14[13] = r_13[13] /*1345*/;
  assign m_14[14] = r_13[14] /*1344*/;
  assign m_14[15] = r_13[15] /*1343*/;
  assign m_14[16] = r_13[16] /*1342*/;
  assign m_14[17] = r_13[17] /*1341*/;
  assign m_14[18] = r_13[18] /*1340*/;
  assign m_14[19] = r_13[19] /*1339*/;
  assign m_14[20] = r_13[20] /*1338*/;
  assign m_14[21] = r_13[21] /*1337*/;
  assign m_14[22] = r_13[22] /*1336*/;
  assign m_14[23] = r_13[23] /*1335*/;
  assign m_14[24] = r_13[24] /*1334*/;
  assign m_14[25] = r_13[25] /*1333*/;
  assign m_14[26] = r_13[26] /*1332*/;
  assign m_14[27] = r_13[27] /*1331*/;
  assign m_14[28] = r_13[28] /*1330*/;
  assign m_14[29] = r_13[29] /*1329*/;
  assign m_14[30] = r_13[30] /*1328*/;
  assign m_14[31] = r_13[31] /*1327*/;
  assign m_14[32] = r_13[32] /*1326*/;
  assign m_14[33] = r_13[33] /*1325*/;
  assign m_14[34] = r_13[34] /*1324*/;
  assign m_14[35] = r_13[35] /*1323*/;
  assign m_14[36] = r_13[36] /*1322*/;
  assign m_14[37] = r_13[37] /*1321*/;
  assign m_14[38] = r_13[38] /*1320*/;
  assign m_14[39] = r_13[39] /*1319*/;
  assign m_14[40] = r_13[40] /*1318*/;
  assign m_14[41] = r_13[41] /*1317*/;
  assign m_14[42] = r_13[42] /*1316*/;
  assign m_14[43] = r_13[43] /*1315*/;
  assign m_14[44] = r_13[43] /*1314*/;
  assign _3652_ = ~q[2] /*1313*/;
  assign _3653_ = sum_14[0] & q[2] /*1312*/;
  assign _3654_ = m_14[0] & _3652_ /*1311*/;
  assign r_14[0] = _3654_ | _3653_ /*1310*/;
  assign _3655_ = ~q[2] /*1309*/;
  assign _3656_ = sum_14[1] & q[2] /*1308*/;
  assign _3657_ = m_14[1] & _3655_ /*1307*/;
  assign r_14[1] = _3657_ | _3656_ /*1306*/;
  assign _3658_ = ~q[2] /*1305*/;
  assign _3659_ = sum_14[2] & q[2] /*1304*/;
  assign _3660_ = m_14[2] & _3658_ /*1303*/;
  assign r_14[2] = _3660_ | _3659_ /*1302*/;
  assign _3661_ = ~q[2] /*1301*/;
  assign _3662_ = sum_14[3] & q[2] /*1300*/;
  assign _3663_ = m_14[3] & _3661_ /*1299*/;
  assign r_14[3] = _3663_ | _3662_ /*1298*/;
  assign _3664_ = ~q[2] /*1297*/;
  assign _3665_ = sum_14[4] & q[2] /*1296*/;
  assign _3666_ = m_14[4] & _3664_ /*1295*/;
  assign r_14[4] = _3666_ | _3665_ /*1294*/;
  assign _3667_ = ~q[2] /*1293*/;
  assign _3668_ = sum_14[5] & q[2] /*1292*/;
  assign _3669_ = m_14[5] & _3667_ /*1291*/;
  assign r_14[5] = _3669_ | _3668_ /*1290*/;
  assign _3670_ = ~q[2] /*1289*/;
  assign _3671_ = sum_14[6] & q[2] /*1288*/;
  assign _3672_ = m_14[6] & _3670_ /*1287*/;
  assign r_14[6] = _3672_ | _3671_ /*1286*/;
  assign _3673_ = ~q[2] /*1285*/;
  assign _3674_ = sum_14[7] & q[2] /*1284*/;
  assign _3675_ = m_14[7] & _3673_ /*1283*/;
  assign r_14[7] = _3675_ | _3674_ /*1282*/;
  assign _3676_ = ~q[2] /*1281*/;
  assign _3677_ = sum_14[8] & q[2] /*1280*/;
  assign _3678_ = m_14[8] & _3676_ /*1279*/;
  assign r_14[8] = _3678_ | _3677_ /*1278*/;
  assign _3679_ = ~q[2] /*1277*/;
  assign _3680_ = sum_14[9] & q[2] /*1276*/;
  assign _3681_ = m_14[9] & _3679_ /*1275*/;
  assign r_14[9] = _3681_ | _3680_ /*1274*/;
  assign _3682_ = ~q[2] /*1273*/;
  assign _3683_ = sum_14[10] & q[2] /*1272*/;
  assign _3684_ = m_14[10] & _3682_ /*1271*/;
  assign r_14[10] = _3684_ | _3683_ /*1270*/;
  assign _3685_ = ~q[2] /*1269*/;
  assign _3686_ = sum_14[11] & q[2] /*1268*/;
  assign _3687_ = m_14[11] & _3685_ /*1267*/;
  assign r_14[11] = _3687_ | _3686_ /*1266*/;
  assign _3688_ = ~q[2] /*1265*/;
  assign _3689_ = sum_14[12] & q[2] /*1264*/;
  assign _3690_ = m_14[12] & _3688_ /*1263*/;
  assign r_14[12] = _3690_ | _3689_ /*1262*/;
  assign _3691_ = ~q[2] /*1261*/;
  assign _3692_ = sum_14[13] & q[2] /*1260*/;
  assign _3693_ = m_14[13] & _3691_ /*1259*/;
  assign r_14[13] = _3693_ | _3692_ /*1258*/;
  assign _3694_ = ~q[2] /*1257*/;
  assign _3695_ = sum_14[14] & q[2] /*1256*/;
  assign _3696_ = m_14[14] & _3694_ /*1255*/;
  assign r_14[14] = _3696_ | _3695_ /*1254*/;
  assign _3697_ = ~q[2] /*1253*/;
  assign _3698_ = sum_14[15] & q[2] /*1252*/;
  assign _3699_ = m_14[15] & _3697_ /*1251*/;
  assign r_14[15] = _3699_ | _3698_ /*1250*/;
  assign _3700_ = ~q[2] /*1249*/;
  assign _3701_ = sum_14[16] & q[2] /*1248*/;
  assign _3702_ = m_14[16] & _3700_ /*1247*/;
  assign r_14[16] = _3702_ | _3701_ /*1246*/;
  assign _3703_ = ~q[2] /*1245*/;
  assign _3704_ = sum_14[17] & q[2] /*1244*/;
  assign _3705_ = m_14[17] & _3703_ /*1243*/;
  assign r_14[17] = _3705_ | _3704_ /*1242*/;
  assign _3706_ = ~q[2] /*1241*/;
  assign _3707_ = sum_14[18] & q[2] /*1240*/;
  assign _3708_ = m_14[18] & _3706_ /*1239*/;
  assign r_14[18] = _3708_ | _3707_ /*1238*/;
  assign _3709_ = ~q[2] /*1237*/;
  assign _3710_ = sum_14[19] & q[2] /*1236*/;
  assign _3711_ = m_14[19] & _3709_ /*1235*/;
  assign r_14[19] = _3711_ | _3710_ /*1234*/;
  assign _3712_ = ~q[2] /*1233*/;
  assign _3713_ = sum_14[20] & q[2] /*1232*/;
  assign _3714_ = m_14[20] & _3712_ /*1231*/;
  assign r_14[20] = _3714_ | _3713_ /*1230*/;
  assign _3715_ = ~q[2] /*1229*/;
  assign _3716_ = sum_14[21] & q[2] /*1228*/;
  assign _3717_ = m_14[21] & _3715_ /*1227*/;
  assign r_14[21] = _3717_ | _3716_ /*1226*/;
  assign _3718_ = ~q[2] /*1225*/;
  assign _3719_ = sum_14[22] & q[2] /*1224*/;
  assign _3720_ = m_14[22] & _3718_ /*1223*/;
  assign r_14[22] = _3720_ | _3719_ /*1222*/;
  assign _3721_ = ~q[2] /*1221*/;
  assign _3722_ = sum_14[23] & q[2] /*1220*/;
  assign _3723_ = m_14[23] & _3721_ /*1219*/;
  assign r_14[23] = _3723_ | _3722_ /*1218*/;
  assign _3724_ = ~q[2] /*1217*/;
  assign _3725_ = sum_14[24] & q[2] /*1216*/;
  assign _3726_ = m_14[24] & _3724_ /*1215*/;
  assign r_14[24] = _3726_ | _3725_ /*1214*/;
  assign _3727_ = ~q[2] /*1213*/;
  assign _3728_ = sum_14[25] & q[2] /*1212*/;
  assign _3729_ = m_14[25] & _3727_ /*1211*/;
  assign r_14[25] = _3729_ | _3728_ /*1210*/;
  assign _3730_ = ~q[2] /*1209*/;
  assign _3731_ = sum_14[26] & q[2] /*1208*/;
  assign _3732_ = m_14[26] & _3730_ /*1207*/;
  assign r_14[26] = _3732_ | _3731_ /*1206*/;
  assign _3733_ = ~q[2] /*1205*/;
  assign _3734_ = sum_14[27] & q[2] /*1204*/;
  assign _3735_ = m_14[27] & _3733_ /*1203*/;
  assign r_14[27] = _3735_ | _3734_ /*1202*/;
  assign _3736_ = ~q[2] /*1201*/;
  assign _3737_ = sum_14[28] & q[2] /*1200*/;
  assign _3738_ = m_14[28] & _3736_ /*1199*/;
  assign r_14[28] = _3738_ | _3737_ /*1198*/;
  assign _3739_ = ~q[2] /*1197*/;
  assign _3740_ = sum_14[29] & q[2] /*1196*/;
  assign _3741_ = m_14[29] & _3739_ /*1195*/;
  assign r_14[29] = _3741_ | _3740_ /*1194*/;
  assign _3742_ = ~q[2] /*1193*/;
  assign _3743_ = sum_14[30] & q[2] /*1192*/;
  assign _3744_ = m_14[30] & _3742_ /*1191*/;
  assign r_14[30] = _3744_ | _3743_ /*1190*/;
  assign _3745_ = ~q[2] /*1189*/;
  assign _3746_ = sum_14[31] & q[2] /*1188*/;
  assign _3747_ = m_14[31] & _3745_ /*1187*/;
  assign r_14[31] = _3747_ | _3746_ /*1186*/;
  assign _3748_ = ~q[2] /*1185*/;
  assign _3749_ = sum_14[32] & q[2] /*1184*/;
  assign _3750_ = m_14[32] & _3748_ /*1183*/;
  assign r_14[32] = _3750_ | _3749_ /*1182*/;
  assign _3751_ = ~q[2] /*1181*/;
  assign _3752_ = sum_14[33] & q[2] /*1180*/;
  assign _3753_ = m_14[33] & _3751_ /*1179*/;
  assign r_14[33] = _3753_ | _3752_ /*1178*/;
  assign _3754_ = ~q[2] /*1177*/;
  assign _3755_ = sum_14[34] & q[2] /*1176*/;
  assign _3756_ = m_14[34] & _3754_ /*1175*/;
  assign r_14[34] = _3756_ | _3755_ /*1174*/;
  assign _3757_ = ~q[2] /*1173*/;
  assign _3758_ = sum_14[35] & q[2] /*1172*/;
  assign _3759_ = m_14[35] & _3757_ /*1171*/;
  assign r_14[35] = _3759_ | _3758_ /*1170*/;
  assign _3760_ = ~q[2] /*1169*/;
  assign _3761_ = sum_14[36] & q[2] /*1168*/;
  assign _3762_ = m_14[36] & _3760_ /*1167*/;
  assign r_14[36] = _3762_ | _3761_ /*1166*/;
  assign _3763_ = ~q[2] /*1165*/;
  assign _3764_ = sum_14[37] & q[2] /*1164*/;
  assign _3765_ = m_14[37] & _3763_ /*1163*/;
  assign r_14[37] = _3765_ | _3764_ /*1162*/;
  assign _3766_ = ~q[2] /*1161*/;
  assign _3767_ = sum_14[38] & q[2] /*1160*/;
  assign _3768_ = m_14[38] & _3766_ /*1159*/;
  assign r_14[38] = _3768_ | _3767_ /*1158*/;
  assign _3769_ = ~q[2] /*1157*/;
  assign _3770_ = sum_14[39] & q[2] /*1156*/;
  assign _3771_ = m_14[39] & _3769_ /*1155*/;
  assign r_14[39] = _3771_ | _3770_ /*1154*/;
  assign _3772_ = ~q[2] /*1153*/;
  assign _3773_ = sum_14[40] & q[2] /*1152*/;
  assign _3774_ = m_14[40] & _3772_ /*1151*/;
  assign r_14[40] = _3774_ | _3773_ /*1150*/;
  assign _3775_ = ~q[2] /*1149*/;
  assign _3776_ = sum_14[41] & q[2] /*1148*/;
  assign _3777_ = m_14[41] & _3775_ /*1147*/;
  assign r_14[41] = _3777_ | _3776_ /*1146*/;
  assign _3778_ = ~q[2] /*1145*/;
  assign _3779_ = sum_14[42] & q[2] /*1144*/;
  assign _3780_ = m_14[42] & _3778_ /*1143*/;
  assign r_14[42] = _3780_ | _3779_ /*1142*/;
  assign _3781_ = ~q[2] /*1141*/;
  assign _3782_ = sum_14[43] & q[2] /*1140*/;
  assign _3783_ = m_14[43] & _3781_ /*1139*/;
  assign r_14[43] = _3783_ | _3782_ /*1138*/;
  assign _3784_ = ~q[2] /*1137*/;
  assign _3785_ = sum_14[44] & q[2] /*1136*/;
  assign _3786_ = m_14[44] & _3784_ /*1135*/;
  assign r_14[44] = _3786_ | _3785_ /*1134*/;
  assign inv_15[0] = oneWire /*1096*/;
  assign inv_15[1] = ~div[0] /*1090*/;
  assign inv_15[2] = ~div[1] /*1084*/;
  assign inv_15[3] = ~div[2] /*1078*/;
  assign inv_15[4] = ~div[3] /*1072*/;
  assign inv_15[5] = ~div[4] /*1066*/;
  assign inv_15[6] = ~div[5] /*1060*/;
  assign inv_15[7] = ~div[6] /*1054*/;
  assign inv_15[8] = ~div[7] /*1048*/;
  assign inv_15[9] = ~div[8] /*1042*/;
  assign inv_15[10] = ~div[9] /*1036*/;
  assign inv_15[11] = ~div[10] /*1030*/;
  assign inv_15[12] = ~div[11] /*1024*/;
  assign inv_15[13] = ~div[12] /*1018*/;
  assign inv_15[14] = ~div[13] /*1012*/;
  assign inv_15[15] = ~div[14] /*1006*/;
  assign inv_15[16] = oneWire /*1000*/;
  assign inv_15[17] = oneWire /*994*/;
  assign inv_15[18] = oneWire /*988*/;
  assign inv_15[19] = oneWire /*982*/;
  assign inv_15[20] = oneWire /*976*/;
  assign inv_15[21] = oneWire /*970*/;
  assign inv_15[22] = oneWire /*964*/;
  assign inv_15[23] = oneWire /*958*/;
  assign inv_15[24] = oneWire /*952*/;
  assign inv_15[25] = oneWire /*946*/;
  assign inv_15[26] = oneWire /*940*/;
  assign inv_15[27] = oneWire /*934*/;
  assign inv_15[28] = oneWire /*928*/;
  assign inv_15[29] = oneWire /*922*/;
  assign inv_15[30] = oneWire /*916*/;
  assign inv_15[31] = oneWire /*910*/;
  assign inv_15[32] = oneWire /*904*/;
  assign inv_15[33] = oneWire /*898*/;
  assign inv_15[34] = oneWire /*892*/;
  assign inv_15[35] = oneWire /*886*/;
  assign inv_15[36] = oneWire /*880*/;
  assign inv_15[37] = oneWire /*874*/;
  assign inv_15[38] = oneWire /*868*/;
  assign inv_15[39] = oneWire /*862*/;
  assign inv_15[40] = oneWire /*856*/;
  assign inv_15[41] = oneWire /*850*/;
  assign inv_15[42] = oneWire /*844*/;
  assign inv_15[43] = oneWire /*838*/;
  assign inv_15[44] = oneWire /*832*/;
  assign _3787_ = inv_15[0] ^ r_14[0] /*1095*/;
  assign sum_15[0] = _3787_ ^ oneWire /*1094*/;
  assign _3788_ = _3787_ & oneWire /*1093*/;
  assign _3789_ = inv_15[0] & r_14[0] /*1092*/;
  assign _3790_ = _3788_ | _3789_ /*1091*/;
  assign _3791_ = inv_15[1] ^ r_14[1] /*1089*/;
  assign sum_15[1] = _3791_ ^ _3790_ /*1088*/;
  assign _3792_ = _3791_ & _3790_ /*1087*/;
  assign _3793_ = inv_15[1] & r_14[1] /*1086*/;
  assign _3794_ = _3792_ | _3793_ /*1085*/;
  assign _3795_ = inv_15[2] ^ r_14[2] /*1083*/;
  assign sum_15[2] = _3795_ ^ _3794_ /*1082*/;
  assign _3796_ = _3795_ & _3794_ /*1081*/;
  assign _3797_ = inv_15[2] & r_14[2] /*1080*/;
  assign _3798_ = _3796_ | _3797_ /*1079*/;
  assign _3799_ = inv_15[3] ^ r_14[3] /*1077*/;
  assign sum_15[3] = _3799_ ^ _3798_ /*1076*/;
  assign _3800_ = _3799_ & _3798_ /*1075*/;
  assign _3801_ = inv_15[3] & r_14[3] /*1074*/;
  assign _3802_ = _3800_ | _3801_ /*1073*/;
  assign _3803_ = inv_15[4] ^ r_14[4] /*1071*/;
  assign sum_15[4] = _3803_ ^ _3802_ /*1070*/;
  assign _3804_ = _3803_ & _3802_ /*1069*/;
  assign _3805_ = inv_15[4] & r_14[4] /*1068*/;
  assign _3806_ = _3804_ | _3805_ /*1067*/;
  assign _3807_ = inv_15[5] ^ r_14[5] /*1065*/;
  assign sum_15[5] = _3807_ ^ _3806_ /*1064*/;
  assign _3808_ = _3807_ & _3806_ /*1063*/;
  assign _3809_ = inv_15[5] & r_14[5] /*1062*/;
  assign _3810_ = _3808_ | _3809_ /*1061*/;
  assign _3811_ = inv_15[6] ^ r_14[6] /*1059*/;
  assign sum_15[6] = _3811_ ^ _3810_ /*1058*/;
  assign _3812_ = _3811_ & _3810_ /*1057*/;
  assign _3813_ = inv_15[6] & r_14[6] /*1056*/;
  assign _3814_ = _3812_ | _3813_ /*1055*/;
  assign _3815_ = inv_15[7] ^ r_14[7] /*1053*/;
  assign sum_15[7] = _3815_ ^ _3814_ /*1052*/;
  assign _3816_ = _3815_ & _3814_ /*1051*/;
  assign _3817_ = inv_15[7] & r_14[7] /*1050*/;
  assign _3818_ = _3816_ | _3817_ /*1049*/;
  assign _3819_ = inv_15[8] ^ r_14[8] /*1047*/;
  assign sum_15[8] = _3819_ ^ _3818_ /*1046*/;
  assign _3820_ = _3819_ & _3818_ /*1045*/;
  assign _3821_ = inv_15[8] & r_14[8] /*1044*/;
  assign _3822_ = _3820_ | _3821_ /*1043*/;
  assign _3823_ = inv_15[9] ^ r_14[9] /*1041*/;
  assign sum_15[9] = _3823_ ^ _3822_ /*1040*/;
  assign _3824_ = _3823_ & _3822_ /*1039*/;
  assign _3825_ = inv_15[9] & r_14[9] /*1038*/;
  assign _3826_ = _3824_ | _3825_ /*1037*/;
  assign _3827_ = inv_15[10] ^ r_14[10] /*1035*/;
  assign sum_15[10] = _3827_ ^ _3826_ /*1034*/;
  assign _3828_ = _3827_ & _3826_ /*1033*/;
  assign _3829_ = inv_15[10] & r_14[10] /*1032*/;
  assign _3830_ = _3828_ | _3829_ /*1031*/;
  assign _3831_ = inv_15[11] ^ r_14[11] /*1029*/;
  assign sum_15[11] = _3831_ ^ _3830_ /*1028*/;
  assign _3832_ = _3831_ & _3830_ /*1027*/;
  assign _3833_ = inv_15[11] & r_14[11] /*1026*/;
  assign _3834_ = _3832_ | _3833_ /*1025*/;
  assign _3835_ = inv_15[12] ^ r_14[12] /*1023*/;
  assign sum_15[12] = _3835_ ^ _3834_ /*1022*/;
  assign _3836_ = _3835_ & _3834_ /*1021*/;
  assign _3837_ = inv_15[12] & r_14[12] /*1020*/;
  assign _3838_ = _3836_ | _3837_ /*1019*/;
  assign _3839_ = inv_15[13] ^ r_14[13] /*1017*/;
  assign sum_15[13] = _3839_ ^ _3838_ /*1016*/;
  assign _3840_ = _3839_ & _3838_ /*1015*/;
  assign _3841_ = inv_15[13] & r_14[13] /*1014*/;
  assign _3842_ = _3840_ | _3841_ /*1013*/;
  assign _3843_ = inv_15[14] ^ r_14[14] /*1011*/;
  assign sum_15[14] = _3843_ ^ _3842_ /*1010*/;
  assign _3844_ = _3843_ & _3842_ /*1009*/;
  assign _3845_ = inv_15[14] & r_14[14] /*1008*/;
  assign _3846_ = _3844_ | _3845_ /*1007*/;
  assign _3847_ = inv_15[15] ^ r_14[15] /*1005*/;
  assign sum_15[15] = _3847_ ^ _3846_ /*1004*/;
  assign _3848_ = _3847_ & _3846_ /*1003*/;
  assign _3849_ = inv_15[15] & r_14[15] /*1002*/;
  assign _3850_ = _3848_ | _3849_ /*1001*/;
  assign _3851_ = inv_15[16] ^ r_14[16] /*999*/;
  assign sum_15[16] = _3851_ ^ _3850_ /*998*/;
  assign _3852_ = _3851_ & _3850_ /*997*/;
  assign _3853_ = inv_15[16] & r_14[16] /*996*/;
  assign _3854_ = _3852_ | _3853_ /*995*/;
  assign _3855_ = inv_15[17] ^ r_14[17] /*993*/;
  assign sum_15[17] = _3855_ ^ _3854_ /*992*/;
  assign _3856_ = _3855_ & _3854_ /*991*/;
  assign _3857_ = inv_15[17] & r_14[17] /*990*/;
  assign _3858_ = _3856_ | _3857_ /*989*/;
  assign _3859_ = inv_15[18] ^ r_14[18] /*987*/;
  assign sum_15[18] = _3859_ ^ _3858_ /*986*/;
  assign _3860_ = _3859_ & _3858_ /*985*/;
  assign _3861_ = inv_15[18] & r_14[18] /*984*/;
  assign _3862_ = _3860_ | _3861_ /*983*/;
  assign _3863_ = inv_15[19] ^ r_14[19] /*981*/;
  assign sum_15[19] = _3863_ ^ _3862_ /*980*/;
  assign _3864_ = _3863_ & _3862_ /*979*/;
  assign _3865_ = inv_15[19] & r_14[19] /*978*/;
  assign _3866_ = _3864_ | _3865_ /*977*/;
  assign _3867_ = inv_15[20] ^ r_14[20] /*975*/;
  assign sum_15[20] = _3867_ ^ _3866_ /*974*/;
  assign _3868_ = _3867_ & _3866_ /*973*/;
  assign _3869_ = inv_15[20] & r_14[20] /*972*/;
  assign _3870_ = _3868_ | _3869_ /*971*/;
  assign _3871_ = inv_15[21] ^ r_14[21] /*969*/;
  assign sum_15[21] = _3871_ ^ _3870_ /*968*/;
  assign _3872_ = _3871_ & _3870_ /*967*/;
  assign _3873_ = inv_15[21] & r_14[21] /*966*/;
  assign _3874_ = _3872_ | _3873_ /*965*/;
  assign _3875_ = inv_15[22] ^ r_14[22] /*963*/;
  assign sum_15[22] = _3875_ ^ _3874_ /*962*/;
  assign _3876_ = _3875_ & _3874_ /*961*/;
  assign _3877_ = inv_15[22] & r_14[22] /*960*/;
  assign _3878_ = _3876_ | _3877_ /*959*/;
  assign _3879_ = inv_15[23] ^ r_14[23] /*957*/;
  assign sum_15[23] = _3879_ ^ _3878_ /*956*/;
  assign _3880_ = _3879_ & _3878_ /*955*/;
  assign _3881_ = inv_15[23] & r_14[23] /*954*/;
  assign _3882_ = _3880_ | _3881_ /*953*/;
  assign _3883_ = inv_15[24] ^ r_14[24] /*951*/;
  assign sum_15[24] = _3883_ ^ _3882_ /*950*/;
  assign _3884_ = _3883_ & _3882_ /*949*/;
  assign _3885_ = inv_15[24] & r_14[24] /*948*/;
  assign _3886_ = _3884_ | _3885_ /*947*/;
  assign _3887_ = inv_15[25] ^ r_14[25] /*945*/;
  assign sum_15[25] = _3887_ ^ _3886_ /*944*/;
  assign _3888_ = _3887_ & _3886_ /*943*/;
  assign _3889_ = inv_15[25] & r_14[25] /*942*/;
  assign _3890_ = _3888_ | _3889_ /*941*/;
  assign _3891_ = inv_15[26] ^ r_14[26] /*939*/;
  assign sum_15[26] = _3891_ ^ _3890_ /*938*/;
  assign _3892_ = _3891_ & _3890_ /*937*/;
  assign _3893_ = inv_15[26] & r_14[26] /*936*/;
  assign _3894_ = _3892_ | _3893_ /*935*/;
  assign _3895_ = inv_15[27] ^ r_14[27] /*933*/;
  assign sum_15[27] = _3895_ ^ _3894_ /*932*/;
  assign _3896_ = _3895_ & _3894_ /*931*/;
  assign _3897_ = inv_15[27] & r_14[27] /*930*/;
  assign _3898_ = _3896_ | _3897_ /*929*/;
  assign _3899_ = inv_15[28] ^ r_14[28] /*927*/;
  assign sum_15[28] = _3899_ ^ _3898_ /*926*/;
  assign _3900_ = _3899_ & _3898_ /*925*/;
  assign _3901_ = inv_15[28] & r_14[28] /*924*/;
  assign _3902_ = _3900_ | _3901_ /*923*/;
  assign _3903_ = inv_15[29] ^ r_14[29] /*921*/;
  assign sum_15[29] = _3903_ ^ _3902_ /*920*/;
  assign _3904_ = _3903_ & _3902_ /*919*/;
  assign _3905_ = inv_15[29] & r_14[29] /*918*/;
  assign _3906_ = _3904_ | _3905_ /*917*/;
  assign _3907_ = inv_15[30] ^ r_14[30] /*915*/;
  assign sum_15[30] = _3907_ ^ _3906_ /*914*/;
  assign _3908_ = _3907_ & _3906_ /*913*/;
  assign _3909_ = inv_15[30] & r_14[30] /*912*/;
  assign _3910_ = _3908_ | _3909_ /*911*/;
  assign _3911_ = inv_15[31] ^ r_14[31] /*909*/;
  assign sum_15[31] = _3911_ ^ _3910_ /*908*/;
  assign _3912_ = _3911_ & _3910_ /*907*/;
  assign _3913_ = inv_15[31] & r_14[31] /*906*/;
  assign _3914_ = _3912_ | _3913_ /*905*/;
  assign _3915_ = inv_15[32] ^ r_14[32] /*903*/;
  assign sum_15[32] = _3915_ ^ _3914_ /*902*/;
  assign _3916_ = _3915_ & _3914_ /*901*/;
  assign _3917_ = inv_15[32] & r_14[32] /*900*/;
  assign _3918_ = _3916_ | _3917_ /*899*/;
  assign _3919_ = inv_15[33] ^ r_14[33] /*897*/;
  assign sum_15[33] = _3919_ ^ _3918_ /*896*/;
  assign _3920_ = _3919_ & _3918_ /*895*/;
  assign _3921_ = inv_15[33] & r_14[33] /*894*/;
  assign _3922_ = _3920_ | _3921_ /*893*/;
  assign _3923_ = inv_15[34] ^ r_14[34] /*891*/;
  assign sum_15[34] = _3923_ ^ _3922_ /*890*/;
  assign _3924_ = _3923_ & _3922_ /*889*/;
  assign _3925_ = inv_15[34] & r_14[34] /*888*/;
  assign _3926_ = _3924_ | _3925_ /*887*/;
  assign _3927_ = inv_15[35] ^ r_14[35] /*885*/;
  assign sum_15[35] = _3927_ ^ _3926_ /*884*/;
  assign _3928_ = _3927_ & _3926_ /*883*/;
  assign _3929_ = inv_15[35] & r_14[35] /*882*/;
  assign _3930_ = _3928_ | _3929_ /*881*/;
  assign _3931_ = inv_15[36] ^ r_14[36] /*879*/;
  assign sum_15[36] = _3931_ ^ _3930_ /*878*/;
  assign _3932_ = _3931_ & _3930_ /*877*/;
  assign _3933_ = inv_15[36] & r_14[36] /*876*/;
  assign _3934_ = _3932_ | _3933_ /*875*/;
  assign _3935_ = inv_15[37] ^ r_14[37] /*873*/;
  assign sum_15[37] = _3935_ ^ _3934_ /*872*/;
  assign _3936_ = _3935_ & _3934_ /*871*/;
  assign _3937_ = inv_15[37] & r_14[37] /*870*/;
  assign _3938_ = _3936_ | _3937_ /*869*/;
  assign _3939_ = inv_15[38] ^ r_14[38] /*867*/;
  assign sum_15[38] = _3939_ ^ _3938_ /*866*/;
  assign _3940_ = _3939_ & _3938_ /*865*/;
  assign _3941_ = inv_15[38] & r_14[38] /*864*/;
  assign _3942_ = _3940_ | _3941_ /*863*/;
  assign _3943_ = inv_15[39] ^ r_14[39] /*861*/;
  assign sum_15[39] = _3943_ ^ _3942_ /*860*/;
  assign _3944_ = _3943_ & _3942_ /*859*/;
  assign _3945_ = inv_15[39] & r_14[39] /*858*/;
  assign _3946_ = _3944_ | _3945_ /*857*/;
  assign _3947_ = inv_15[40] ^ r_14[40] /*855*/;
  assign sum_15[40] = _3947_ ^ _3946_ /*854*/;
  assign _3948_ = _3947_ & _3946_ /*853*/;
  assign _3949_ = inv_15[40] & r_14[40] /*852*/;
  assign _3950_ = _3948_ | _3949_ /*851*/;
  assign _3951_ = inv_15[41] ^ r_14[41] /*849*/;
  assign sum_15[41] = _3951_ ^ _3950_ /*848*/;
  assign _3952_ = _3951_ & _3950_ /*847*/;
  assign _3953_ = inv_15[41] & r_14[41] /*846*/;
  assign _3954_ = _3952_ | _3953_ /*845*/;
  assign _3955_ = inv_15[42] ^ r_14[42] /*843*/;
  assign sum_15[42] = _3955_ ^ _3954_ /*842*/;
  assign _3956_ = _3955_ & _3954_ /*841*/;
  assign _3957_ = inv_15[42] & r_14[42] /*840*/;
  assign _3958_ = _3956_ | _3957_ /*839*/;
  assign _3959_ = inv_15[43] ^ r_14[43] /*837*/;
  assign sum_15[43] = _3959_ ^ _3958_ /*836*/;
  assign _3960_ = _3959_ & _3958_ /*835*/;
  assign _3961_ = inv_15[43] & r_14[43] /*834*/;
  assign _3962_ = _3960_ | _3961_ /*833*/;
  assign _3963_ = inv_15[44] ^ r_14[44] /*831*/;
  assign sum_15[44] = _3963_ ^ _3962_ /*830*/;
  assign _3964_ = _3963_ & _3962_ /*829*/;
  assign _3965_ = inv_15[44] & r_14[44] /*828*/;
  assign _3966_ = _3964_ | _3965_ /*827*/;
  assign _3967_ = _3966_ ^ _3962_ /*826*/;
  assign _3968_ = ~_3967_ /*825*/;
  assign _3969_ = sum_15[44] & _3968_ /*824*/;
  assign _3970_ = _3967_ & _3966_ /*823*/;
  assign sum_15[45] = _3970_ | _3969_ /*822*/;
  assign q[1] = ~sum_15[45] /*821*/;
  assign m_15[0] = r_14[0] /*820*/;
  assign m_15[1] = r_14[1] /*819*/;
  assign m_15[2] = r_14[2] /*818*/;
  assign m_15[3] = r_14[3] /*817*/;
  assign m_15[4] = r_14[4] /*816*/;
  assign m_15[5] = r_14[5] /*815*/;
  assign m_15[6] = r_14[6] /*814*/;
  assign m_15[7] = r_14[7] /*813*/;
  assign m_15[8] = r_14[8] /*812*/;
  assign m_15[9] = r_14[9] /*811*/;
  assign m_15[10] = r_14[10] /*810*/;
  assign m_15[11] = r_14[11] /*809*/;
  assign m_15[12] = r_14[12] /*808*/;
  assign m_15[13] = r_14[13] /*807*/;
  assign m_15[14] = r_14[14] /*806*/;
  assign m_15[15] = r_14[15] /*805*/;
  assign m_15[16] = r_14[16] /*804*/;
  assign m_15[17] = r_14[17] /*803*/;
  assign m_15[18] = r_14[18] /*802*/;
  assign m_15[19] = r_14[19] /*801*/;
  assign m_15[20] = r_14[20] /*800*/;
  assign m_15[21] = r_14[21] /*799*/;
  assign m_15[22] = r_14[22] /*798*/;
  assign m_15[23] = r_14[23] /*797*/;
  assign m_15[24] = r_14[24] /*796*/;
  assign m_15[25] = r_14[25] /*795*/;
  assign m_15[26] = r_14[26] /*794*/;
  assign m_15[27] = r_14[27] /*793*/;
  assign m_15[28] = r_14[28] /*792*/;
  assign m_15[29] = r_14[29] /*791*/;
  assign m_15[30] = r_14[30] /*790*/;
  assign m_15[31] = r_14[31] /*789*/;
  assign m_15[32] = r_14[32] /*788*/;
  assign m_15[33] = r_14[33] /*787*/;
  assign m_15[34] = r_14[34] /*786*/;
  assign m_15[35] = r_14[35] /*785*/;
  assign m_15[36] = r_14[36] /*784*/;
  assign m_15[37] = r_14[37] /*783*/;
  assign m_15[38] = r_14[38] /*782*/;
  assign m_15[39] = r_14[39] /*781*/;
  assign m_15[40] = r_14[40] /*780*/;
  assign m_15[41] = r_14[41] /*779*/;
  assign m_15[42] = r_14[42] /*778*/;
  assign m_15[43] = r_14[43] /*777*/;
  assign m_15[44] = r_14[44] /*776*/;
  assign m_15[45] = r_14[44] /*775*/;
  assign _3972_ = ~q[1] /*774*/;
  assign _3973_ = sum_15[0] & q[1] /*773*/;
  assign _3974_ = m_15[0] & _3972_ /*772*/;
  assign r_15[0] = _3974_ | _3973_ /*771*/;
  assign _3975_ = ~q[1] /*770*/;
  assign _3976_ = sum_15[1] & q[1] /*769*/;
  assign _3977_ = m_15[1] & _3975_ /*768*/;
  assign r_15[1] = _3977_ | _3976_ /*767*/;
  assign _3978_ = ~q[1] /*766*/;
  assign _3979_ = sum_15[2] & q[1] /*765*/;
  assign _3980_ = m_15[2] & _3978_ /*764*/;
  assign r_15[2] = _3980_ | _3979_ /*763*/;
  assign _3981_ = ~q[1] /*762*/;
  assign _3982_ = sum_15[3] & q[1] /*761*/;
  assign _3983_ = m_15[3] & _3981_ /*760*/;
  assign r_15[3] = _3983_ | _3982_ /*759*/;
  assign _3984_ = ~q[1] /*758*/;
  assign _3985_ = sum_15[4] & q[1] /*757*/;
  assign _3986_ = m_15[4] & _3984_ /*756*/;
  assign r_15[4] = _3986_ | _3985_ /*755*/;
  assign _3987_ = ~q[1] /*754*/;
  assign _3988_ = sum_15[5] & q[1] /*753*/;
  assign _3989_ = m_15[5] & _3987_ /*752*/;
  assign r_15[5] = _3989_ | _3988_ /*751*/;
  assign _3990_ = ~q[1] /*750*/;
  assign _3991_ = sum_15[6] & q[1] /*749*/;
  assign _3992_ = m_15[6] & _3990_ /*748*/;
  assign r_15[6] = _3992_ | _3991_ /*747*/;
  assign _3993_ = ~q[1] /*746*/;
  assign _3994_ = sum_15[7] & q[1] /*745*/;
  assign _3995_ = m_15[7] & _3993_ /*744*/;
  assign r_15[7] = _3995_ | _3994_ /*743*/;
  assign _3996_ = ~q[1] /*742*/;
  assign _3997_ = sum_15[8] & q[1] /*741*/;
  assign _3998_ = m_15[8] & _3996_ /*740*/;
  assign r_15[8] = _3998_ | _3997_ /*739*/;
  assign _3999_ = ~q[1] /*738*/;
  assign _4000_ = sum_15[9] & q[1] /*737*/;
  assign _4001_ = m_15[9] & _3999_ /*736*/;
  assign r_15[9] = _4001_ | _4000_ /*735*/;
  assign _4002_ = ~q[1] /*734*/;
  assign _4003_ = sum_15[10] & q[1] /*733*/;
  assign _4004_ = m_15[10] & _4002_ /*732*/;
  assign r_15[10] = _4004_ | _4003_ /*731*/;
  assign _4005_ = ~q[1] /*730*/;
  assign _4006_ = sum_15[11] & q[1] /*729*/;
  assign _4007_ = m_15[11] & _4005_ /*728*/;
  assign r_15[11] = _4007_ | _4006_ /*727*/;
  assign _4008_ = ~q[1] /*726*/;
  assign _4009_ = sum_15[12] & q[1] /*725*/;
  assign _4010_ = m_15[12] & _4008_ /*724*/;
  assign r_15[12] = _4010_ | _4009_ /*723*/;
  assign _4011_ = ~q[1] /*722*/;
  assign _4012_ = sum_15[13] & q[1] /*721*/;
  assign _4013_ = m_15[13] & _4011_ /*720*/;
  assign r_15[13] = _4013_ | _4012_ /*719*/;
  assign _4014_ = ~q[1] /*718*/;
  assign _4015_ = sum_15[14] & q[1] /*717*/;
  assign _4016_ = m_15[14] & _4014_ /*716*/;
  assign r_15[14] = _4016_ | _4015_ /*715*/;
  assign _4017_ = ~q[1] /*714*/;
  assign _4018_ = sum_15[15] & q[1] /*713*/;
  assign _4019_ = m_15[15] & _4017_ /*712*/;
  assign r_15[15] = _4019_ | _4018_ /*711*/;
  assign _4020_ = ~q[1] /*710*/;
  assign _4021_ = sum_15[16] & q[1] /*709*/;
  assign _4022_ = m_15[16] & _4020_ /*708*/;
  assign r_15[16] = _4022_ | _4021_ /*707*/;
  assign _4023_ = ~q[1] /*706*/;
  assign _4024_ = sum_15[17] & q[1] /*705*/;
  assign _4025_ = m_15[17] & _4023_ /*704*/;
  assign r_15[17] = _4025_ | _4024_ /*703*/;
  assign _4026_ = ~q[1] /*702*/;
  assign _4027_ = sum_15[18] & q[1] /*701*/;
  assign _4028_ = m_15[18] & _4026_ /*700*/;
  assign r_15[18] = _4028_ | _4027_ /*699*/;
  assign _4029_ = ~q[1] /*698*/;
  assign _4030_ = sum_15[19] & q[1] /*697*/;
  assign _4031_ = m_15[19] & _4029_ /*696*/;
  assign r_15[19] = _4031_ | _4030_ /*695*/;
  assign _4032_ = ~q[1] /*694*/;
  assign _4033_ = sum_15[20] & q[1] /*693*/;
  assign _4034_ = m_15[20] & _4032_ /*692*/;
  assign r_15[20] = _4034_ | _4033_ /*691*/;
  assign _4035_ = ~q[1] /*690*/;
  assign _4036_ = sum_15[21] & q[1] /*689*/;
  assign _4037_ = m_15[21] & _4035_ /*688*/;
  assign r_15[21] = _4037_ | _4036_ /*687*/;
  assign _4038_ = ~q[1] /*686*/;
  assign _4039_ = sum_15[22] & q[1] /*685*/;
  assign _4040_ = m_15[22] & _4038_ /*684*/;
  assign r_15[22] = _4040_ | _4039_ /*683*/;
  assign _4041_ = ~q[1] /*682*/;
  assign _4042_ = sum_15[23] & q[1] /*681*/;
  assign _4043_ = m_15[23] & _4041_ /*680*/;
  assign r_15[23] = _4043_ | _4042_ /*679*/;
  assign _4044_ = ~q[1] /*678*/;
  assign _4045_ = sum_15[24] & q[1] /*677*/;
  assign _4046_ = m_15[24] & _4044_ /*676*/;
  assign r_15[24] = _4046_ | _4045_ /*675*/;
  assign _4047_ = ~q[1] /*674*/;
  assign _4048_ = sum_15[25] & q[1] /*673*/;
  assign _4049_ = m_15[25] & _4047_ /*672*/;
  assign r_15[25] = _4049_ | _4048_ /*671*/;
  assign _4050_ = ~q[1] /*670*/;
  assign _4051_ = sum_15[26] & q[1] /*669*/;
  assign _4052_ = m_15[26] & _4050_ /*668*/;
  assign r_15[26] = _4052_ | _4051_ /*667*/;
  assign _4053_ = ~q[1] /*666*/;
  assign _4054_ = sum_15[27] & q[1] /*665*/;
  assign _4055_ = m_15[27] & _4053_ /*664*/;
  assign r_15[27] = _4055_ | _4054_ /*663*/;
  assign _4056_ = ~q[1] /*662*/;
  assign _4057_ = sum_15[28] & q[1] /*661*/;
  assign _4058_ = m_15[28] & _4056_ /*660*/;
  assign r_15[28] = _4058_ | _4057_ /*659*/;
  assign _4059_ = ~q[1] /*658*/;
  assign _4060_ = sum_15[29] & q[1] /*657*/;
  assign _4061_ = m_15[29] & _4059_ /*656*/;
  assign r_15[29] = _4061_ | _4060_ /*655*/;
  assign _4062_ = ~q[1] /*654*/;
  assign _4063_ = sum_15[30] & q[1] /*653*/;
  assign _4064_ = m_15[30] & _4062_ /*652*/;
  assign r_15[30] = _4064_ | _4063_ /*651*/;
  assign _4065_ = ~q[1] /*650*/;
  assign _4066_ = sum_15[31] & q[1] /*649*/;
  assign _4067_ = m_15[31] & _4065_ /*648*/;
  assign r_15[31] = _4067_ | _4066_ /*647*/;
  assign _4068_ = ~q[1] /*646*/;
  assign _4069_ = sum_15[32] & q[1] /*645*/;
  assign _4070_ = m_15[32] & _4068_ /*644*/;
  assign r_15[32] = _4070_ | _4069_ /*643*/;
  assign _4071_ = ~q[1] /*642*/;
  assign _4072_ = sum_15[33] & q[1] /*641*/;
  assign _4073_ = m_15[33] & _4071_ /*640*/;
  assign r_15[33] = _4073_ | _4072_ /*639*/;
  assign _4074_ = ~q[1] /*638*/;
  assign _4075_ = sum_15[34] & q[1] /*637*/;
  assign _4076_ = m_15[34] & _4074_ /*636*/;
  assign r_15[34] = _4076_ | _4075_ /*635*/;
  assign _4077_ = ~q[1] /*634*/;
  assign _4078_ = sum_15[35] & q[1] /*633*/;
  assign _4079_ = m_15[35] & _4077_ /*632*/;
  assign r_15[35] = _4079_ | _4078_ /*631*/;
  assign _4080_ = ~q[1] /*630*/;
  assign _4081_ = sum_15[36] & q[1] /*629*/;
  assign _4082_ = m_15[36] & _4080_ /*628*/;
  assign r_15[36] = _4082_ | _4081_ /*627*/;
  assign _4083_ = ~q[1] /*626*/;
  assign _4084_ = sum_15[37] & q[1] /*625*/;
  assign _4085_ = m_15[37] & _4083_ /*624*/;
  assign r_15[37] = _4085_ | _4084_ /*623*/;
  assign _4086_ = ~q[1] /*622*/;
  assign _4087_ = sum_15[38] & q[1] /*621*/;
  assign _4088_ = m_15[38] & _4086_ /*620*/;
  assign r_15[38] = _4088_ | _4087_ /*619*/;
  assign _4089_ = ~q[1] /*618*/;
  assign _4090_ = sum_15[39] & q[1] /*617*/;
  assign _4091_ = m_15[39] & _4089_ /*616*/;
  assign r_15[39] = _4091_ | _4090_ /*615*/;
  assign _4092_ = ~q[1] /*614*/;
  assign _4093_ = sum_15[40] & q[1] /*613*/;
  assign _4094_ = m_15[40] & _4092_ /*612*/;
  assign r_15[40] = _4094_ | _4093_ /*611*/;
  assign _4095_ = ~q[1] /*610*/;
  assign _4096_ = sum_15[41] & q[1] /*609*/;
  assign _4097_ = m_15[41] & _4095_ /*608*/;
  assign r_15[41] = _4097_ | _4096_ /*607*/;
  assign _4098_ = ~q[1] /*606*/;
  assign _4099_ = sum_15[42] & q[1] /*605*/;
  assign _4100_ = m_15[42] & _4098_ /*604*/;
  assign r_15[42] = _4100_ | _4099_ /*603*/;
  assign _4101_ = ~q[1] /*602*/;
  assign _4102_ = sum_15[43] & q[1] /*601*/;
  assign _4103_ = m_15[43] & _4101_ /*600*/;
  assign r_15[43] = _4103_ | _4102_ /*599*/;
  assign _4104_ = ~q[1] /*598*/;
  assign _4105_ = sum_15[44] & q[1] /*597*/;
  assign _4106_ = m_15[44] & _4104_ /*596*/;
  assign r_15[44] = _4106_ | _4105_ /*595*/;
  assign _4107_ = ~q[1] /*594*/;
  assign _4108_ = sum_15[45] & q[1] /*593*/;
  assign _4109_ = m_15[45] & _4107_ /*592*/;
  assign r_15[45] = _4109_ | _4108_ /*591*/;
  assign inv_16[0] = ~div[0] /*564*/;
  assign inv_16[1] = ~div[1] /*558*/;
  assign inv_16[2] = ~div[2] /*552*/;
  assign inv_16[3] = ~div[3] /*546*/;
  assign inv_16[4] = ~div[4] /*540*/;
  assign inv_16[5] = ~div[5] /*534*/;
  assign inv_16[6] = ~div[6] /*528*/;
  assign inv_16[7] = ~div[7] /*522*/;
  assign inv_16[8] = ~div[8] /*516*/;
  assign inv_16[9] = ~div[9] /*510*/;
  assign inv_16[10] = ~div[10] /*504*/;
  assign inv_16[11] = ~div[11] /*498*/;
  assign inv_16[12] = ~div[12] /*492*/;
  assign inv_16[13] = ~div[13] /*486*/;
  assign inv_16[14] = ~div[14] /*480*/;
  assign inv_16[15] = oneWire /*474*/;
  assign inv_16[16] = oneWire /*468*/;
  assign inv_16[17] = oneWire /*462*/;
  assign inv_16[18] = oneWire /*456*/;
  assign inv_16[19] = oneWire /*450*/;
  assign inv_16[20] = oneWire /*444*/;
  assign inv_16[21] = oneWire /*438*/;
  assign inv_16[22] = oneWire /*432*/;
  assign inv_16[23] = oneWire /*426*/;
  assign inv_16[24] = oneWire /*420*/;
  assign inv_16[25] = oneWire /*414*/;
  assign inv_16[26] = oneWire /*408*/;
  assign inv_16[27] = oneWire /*402*/;
  assign inv_16[28] = oneWire /*396*/;
  assign inv_16[29] = oneWire /*390*/;
  assign inv_16[30] = oneWire /*384*/;
  assign inv_16[31] = oneWire /*378*/;
  assign inv_16[32] = oneWire /*372*/;
  assign inv_16[33] = oneWire /*366*/;
  assign inv_16[34] = oneWire /*360*/;
  assign inv_16[35] = oneWire /*354*/;
  assign inv_16[36] = oneWire /*348*/;
  assign inv_16[37] = oneWire /*342*/;
  assign inv_16[38] = oneWire /*336*/;
  assign inv_16[39] = oneWire /*330*/;
  assign inv_16[40] = oneWire /*324*/;
  assign inv_16[41] = oneWire /*318*/;
  assign inv_16[42] = oneWire /*312*/;
  assign inv_16[43] = oneWire /*306*/;
  assign inv_16[44] = oneWire /*300*/;
  assign inv_16[45] = oneWire /*294*/;
  assign _4110_ = inv_16[0] ^ r_15[0] /*563*/;
  assign sum_16[0] = _4110_ ^ oneWire /*562*/;
  assign _4111_ = _4110_ & oneWire /*561*/;
  assign _4112_ = inv_16[0] & r_15[0] /*560*/;
  assign _4113_ = _4111_ | _4112_ /*559*/;
  assign _4114_ = inv_16[1] ^ r_15[1] /*557*/;
  assign sum_16[1] = _4114_ ^ _4113_ /*556*/;
  assign _4115_ = _4114_ & _4113_ /*555*/;
  assign _4116_ = inv_16[1] & r_15[1] /*554*/;
  assign _4117_ = _4115_ | _4116_ /*553*/;
  assign _4118_ = inv_16[2] ^ r_15[2] /*551*/;
  assign sum_16[2] = _4118_ ^ _4117_ /*550*/;
  assign _4119_ = _4118_ & _4117_ /*549*/;
  assign _4120_ = inv_16[2] & r_15[2] /*548*/;
  assign _4121_ = _4119_ | _4120_ /*547*/;
  assign _4122_ = inv_16[3] ^ r_15[3] /*545*/;
  assign sum_16[3] = _4122_ ^ _4121_ /*544*/;
  assign _4123_ = _4122_ & _4121_ /*543*/;
  assign _4124_ = inv_16[3] & r_15[3] /*542*/;
  assign _4125_ = _4123_ | _4124_ /*541*/;
  assign _4126_ = inv_16[4] ^ r_15[4] /*539*/;
  assign sum_16[4] = _4126_ ^ _4125_ /*538*/;
  assign _4127_ = _4126_ & _4125_ /*537*/;
  assign _4128_ = inv_16[4] & r_15[4] /*536*/;
  assign _4129_ = _4127_ | _4128_ /*535*/;
  assign _4130_ = inv_16[5] ^ r_15[5] /*533*/;
  assign sum_16[5] = _4130_ ^ _4129_ /*532*/;
  assign _4131_ = _4130_ & _4129_ /*531*/;
  assign _4132_ = inv_16[5] & r_15[5] /*530*/;
  assign _4133_ = _4131_ | _4132_ /*529*/;
  assign _4134_ = inv_16[6] ^ r_15[6] /*527*/;
  assign sum_16[6] = _4134_ ^ _4133_ /*526*/;
  assign _4135_ = _4134_ & _4133_ /*525*/;
  assign _4136_ = inv_16[6] & r_15[6] /*524*/;
  assign _4137_ = _4135_ | _4136_ /*523*/;
  assign _4138_ = inv_16[7] ^ r_15[7] /*521*/;
  assign sum_16[7] = _4138_ ^ _4137_ /*520*/;
  assign _4139_ = _4138_ & _4137_ /*519*/;
  assign _4140_ = inv_16[7] & r_15[7] /*518*/;
  assign _4141_ = _4139_ | _4140_ /*517*/;
  assign _4142_ = inv_16[8] ^ r_15[8] /*515*/;
  assign sum_16[8] = _4142_ ^ _4141_ /*514*/;
  assign _4143_ = _4142_ & _4141_ /*513*/;
  assign _4144_ = inv_16[8] & r_15[8] /*512*/;
  assign _4145_ = _4143_ | _4144_ /*511*/;
  assign _4146_ = inv_16[9] ^ r_15[9] /*509*/;
  assign sum_16[9] = _4146_ ^ _4145_ /*508*/;
  assign _4147_ = _4146_ & _4145_ /*507*/;
  assign _4148_ = inv_16[9] & r_15[9] /*506*/;
  assign _4149_ = _4147_ | _4148_ /*505*/;
  assign _4150_ = inv_16[10] ^ r_15[10] /*503*/;
  assign sum_16[10] = _4150_ ^ _4149_ /*502*/;
  assign _4151_ = _4150_ & _4149_ /*501*/;
  assign _4152_ = inv_16[10] & r_15[10] /*500*/;
  assign _4153_ = _4151_ | _4152_ /*499*/;
  assign _4154_ = inv_16[11] ^ r_15[11] /*497*/;
  assign sum_16[11] = _4154_ ^ _4153_ /*496*/;
  assign _4155_ = _4154_ & _4153_ /*495*/;
  assign _4156_ = inv_16[11] & r_15[11] /*494*/;
  assign _4157_ = _4155_ | _4156_ /*493*/;
  assign _4158_ = inv_16[12] ^ r_15[12] /*491*/;
  assign sum_16[12] = _4158_ ^ _4157_ /*490*/;
  assign _4159_ = _4158_ & _4157_ /*489*/;
  assign _4160_ = inv_16[12] & r_15[12] /*488*/;
  assign _4161_ = _4159_ | _4160_ /*487*/;
  assign _4162_ = inv_16[13] ^ r_15[13] /*485*/;
  assign sum_16[13] = _4162_ ^ _4161_ /*484*/;
  assign _4163_ = _4162_ & _4161_ /*483*/;
  assign _4164_ = inv_16[13] & r_15[13] /*482*/;
  assign _4165_ = _4163_ | _4164_ /*481*/;
  assign _4166_ = inv_16[14] ^ r_15[14] /*479*/;
  assign sum_16[14] = _4166_ ^ _4165_ /*478*/;
  assign _4167_ = _4166_ & _4165_ /*477*/;
  assign _4168_ = inv_16[14] & r_15[14] /*476*/;
  assign _4169_ = _4167_ | _4168_ /*475*/;
  assign _4170_ = inv_16[15] ^ r_15[15] /*473*/;
  assign sum_16[15] = _4170_ ^ _4169_ /*472*/;
  assign _4171_ = _4170_ & _4169_ /*471*/;
  assign _4172_ = inv_16[15] & r_15[15] /*470*/;
  assign _4173_ = _4171_ | _4172_ /*469*/;
  assign _4174_ = inv_16[16] ^ r_15[16] /*467*/;
  assign sum_16[16] = _4174_ ^ _4173_ /*466*/;
  assign _4175_ = _4174_ & _4173_ /*465*/;
  assign _4176_ = inv_16[16] & r_15[16] /*464*/;
  assign _4177_ = _4175_ | _4176_ /*463*/;
  assign _4178_ = inv_16[17] ^ r_15[17] /*461*/;
  assign sum_16[17] = _4178_ ^ _4177_ /*460*/;
  assign _4179_ = _4178_ & _4177_ /*459*/;
  assign _4180_ = inv_16[17] & r_15[17] /*458*/;
  assign _4181_ = _4179_ | _4180_ /*457*/;
  assign _4182_ = inv_16[18] ^ r_15[18] /*455*/;
  assign sum_16[18] = _4182_ ^ _4181_ /*454*/;
  assign _4183_ = _4182_ & _4181_ /*453*/;
  assign _4184_ = inv_16[18] & r_15[18] /*452*/;
  assign _4185_ = _4183_ | _4184_ /*451*/;
  assign _4186_ = inv_16[19] ^ r_15[19] /*449*/;
  assign sum_16[19] = _4186_ ^ _4185_ /*448*/;
  assign _4187_ = _4186_ & _4185_ /*447*/;
  assign _4188_ = inv_16[19] & r_15[19] /*446*/;
  assign _4189_ = _4187_ | _4188_ /*445*/;
  assign _4190_ = inv_16[20] ^ r_15[20] /*443*/;
  assign sum_16[20] = _4190_ ^ _4189_ /*442*/;
  assign _4191_ = _4190_ & _4189_ /*441*/;
  assign _4192_ = inv_16[20] & r_15[20] /*440*/;
  assign _4193_ = _4191_ | _4192_ /*439*/;
  assign _4194_ = inv_16[21] ^ r_15[21] /*437*/;
  assign sum_16[21] = _4194_ ^ _4193_ /*436*/;
  assign _4195_ = _4194_ & _4193_ /*435*/;
  assign _4196_ = inv_16[21] & r_15[21] /*434*/;
  assign _4197_ = _4195_ | _4196_ /*433*/;
  assign _4198_ = inv_16[22] ^ r_15[22] /*431*/;
  assign sum_16[22] = _4198_ ^ _4197_ /*430*/;
  assign _4199_ = _4198_ & _4197_ /*429*/;
  assign _4200_ = inv_16[22] & r_15[22] /*428*/;
  assign _4201_ = _4199_ | _4200_ /*427*/;
  assign _4202_ = inv_16[23] ^ r_15[23] /*425*/;
  assign sum_16[23] = _4202_ ^ _4201_ /*424*/;
  assign _4203_ = _4202_ & _4201_ /*423*/;
  assign _4204_ = inv_16[23] & r_15[23] /*422*/;
  assign _4205_ = _4203_ | _4204_ /*421*/;
  assign _4206_ = inv_16[24] ^ r_15[24] /*419*/;
  assign sum_16[24] = _4206_ ^ _4205_ /*418*/;
  assign _4207_ = _4206_ & _4205_ /*417*/;
  assign _4208_ = inv_16[24] & r_15[24] /*416*/;
  assign _4209_ = _4207_ | _4208_ /*415*/;
  assign _4210_ = inv_16[25] ^ r_15[25] /*413*/;
  assign sum_16[25] = _4210_ ^ _4209_ /*412*/;
  assign _4211_ = _4210_ & _4209_ /*411*/;
  assign _4212_ = inv_16[25] & r_15[25] /*410*/;
  assign _4213_ = _4211_ | _4212_ /*409*/;
  assign _4214_ = inv_16[26] ^ r_15[26] /*407*/;
  assign sum_16[26] = _4214_ ^ _4213_ /*406*/;
  assign _4215_ = _4214_ & _4213_ /*405*/;
  assign _4216_ = inv_16[26] & r_15[26] /*404*/;
  assign _4217_ = _4215_ | _4216_ /*403*/;
  assign _4218_ = inv_16[27] ^ r_15[27] /*401*/;
  assign sum_16[27] = _4218_ ^ _4217_ /*400*/;
  assign _4219_ = _4218_ & _4217_ /*399*/;
  assign _4220_ = inv_16[27] & r_15[27] /*398*/;
  assign _4221_ = _4219_ | _4220_ /*397*/;
  assign _4222_ = inv_16[28] ^ r_15[28] /*395*/;
  assign sum_16[28] = _4222_ ^ _4221_ /*394*/;
  assign _4223_ = _4222_ & _4221_ /*393*/;
  assign _4224_ = inv_16[28] & r_15[28] /*392*/;
  assign _4225_ = _4223_ | _4224_ /*391*/;
  assign _4226_ = inv_16[29] ^ r_15[29] /*389*/;
  assign sum_16[29] = _4226_ ^ _4225_ /*388*/;
  assign _4227_ = _4226_ & _4225_ /*387*/;
  assign _4228_ = inv_16[29] & r_15[29] /*386*/;
  assign _4229_ = _4227_ | _4228_ /*385*/;
  assign _4230_ = inv_16[30] ^ r_15[30] /*383*/;
  assign sum_16[30] = _4230_ ^ _4229_ /*382*/;
  assign _4231_ = _4230_ & _4229_ /*381*/;
  assign _4232_ = inv_16[30] & r_15[30] /*380*/;
  assign _4233_ = _4231_ | _4232_ /*379*/;
  assign _4234_ = inv_16[31] ^ r_15[31] /*377*/;
  assign sum_16[31] = _4234_ ^ _4233_ /*376*/;
  assign _4235_ = _4234_ & _4233_ /*375*/;
  assign _4236_ = inv_16[31] & r_15[31] /*374*/;
  assign _4237_ = _4235_ | _4236_ /*373*/;
  assign _4238_ = inv_16[32] ^ r_15[32] /*371*/;
  assign sum_16[32] = _4238_ ^ _4237_ /*370*/;
  assign _4239_ = _4238_ & _4237_ /*369*/;
  assign _4240_ = inv_16[32] & r_15[32] /*368*/;
  assign _4241_ = _4239_ | _4240_ /*367*/;
  assign _4242_ = inv_16[33] ^ r_15[33] /*365*/;
  assign sum_16[33] = _4242_ ^ _4241_ /*364*/;
  assign _4243_ = _4242_ & _4241_ /*363*/;
  assign _4244_ = inv_16[33] & r_15[33] /*362*/;
  assign _4245_ = _4243_ | _4244_ /*361*/;
  assign _4246_ = inv_16[34] ^ r_15[34] /*359*/;
  assign sum_16[34] = _4246_ ^ _4245_ /*358*/;
  assign _4247_ = _4246_ & _4245_ /*357*/;
  assign _4248_ = inv_16[34] & r_15[34] /*356*/;
  assign _4249_ = _4247_ | _4248_ /*355*/;
  assign _4250_ = inv_16[35] ^ r_15[35] /*353*/;
  assign sum_16[35] = _4250_ ^ _4249_ /*352*/;
  assign _4251_ = _4250_ & _4249_ /*351*/;
  assign _4252_ = inv_16[35] & r_15[35] /*350*/;
  assign _4253_ = _4251_ | _4252_ /*349*/;
  assign _4254_ = inv_16[36] ^ r_15[36] /*347*/;
  assign sum_16[36] = _4254_ ^ _4253_ /*346*/;
  assign _4255_ = _4254_ & _4253_ /*345*/;
  assign _4256_ = inv_16[36] & r_15[36] /*344*/;
  assign _4257_ = _4255_ | _4256_ /*343*/;
  assign _4258_ = inv_16[37] ^ r_15[37] /*341*/;
  assign sum_16[37] = _4258_ ^ _4257_ /*340*/;
  assign _4259_ = _4258_ & _4257_ /*339*/;
  assign _4260_ = inv_16[37] & r_15[37] /*338*/;
  assign _4261_ = _4259_ | _4260_ /*337*/;
  assign _4262_ = inv_16[38] ^ r_15[38] /*335*/;
  assign sum_16[38] = _4262_ ^ _4261_ /*334*/;
  assign _4263_ = _4262_ & _4261_ /*333*/;
  assign _4264_ = inv_16[38] & r_15[38] /*332*/;
  assign _4265_ = _4263_ | _4264_ /*331*/;
  assign _4266_ = inv_16[39] ^ r_15[39] /*329*/;
  assign sum_16[39] = _4266_ ^ _4265_ /*328*/;
  assign _4267_ = _4266_ & _4265_ /*327*/;
  assign _4268_ = inv_16[39] & r_15[39] /*326*/;
  assign _4269_ = _4267_ | _4268_ /*325*/;
  assign _4270_ = inv_16[40] ^ r_15[40] /*323*/;
  assign sum_16[40] = _4270_ ^ _4269_ /*322*/;
  assign _4271_ = _4270_ & _4269_ /*321*/;
  assign _4272_ = inv_16[40] & r_15[40] /*320*/;
  assign _4273_ = _4271_ | _4272_ /*319*/;
  assign _4274_ = inv_16[41] ^ r_15[41] /*317*/;
  assign sum_16[41] = _4274_ ^ _4273_ /*316*/;
  assign _4275_ = _4274_ & _4273_ /*315*/;
  assign _4276_ = inv_16[41] & r_15[41] /*314*/;
  assign _4277_ = _4275_ | _4276_ /*313*/;
  assign _4278_ = inv_16[42] ^ r_15[42] /*311*/;
  assign sum_16[42] = _4278_ ^ _4277_ /*310*/;
  assign _4279_ = _4278_ & _4277_ /*309*/;
  assign _4280_ = inv_16[42] & r_15[42] /*308*/;
  assign _4281_ = _4279_ | _4280_ /*307*/;
  assign _4282_ = inv_16[43] ^ r_15[43] /*305*/;
  assign sum_16[43] = _4282_ ^ _4281_ /*304*/;
  assign _4283_ = _4282_ & _4281_ /*303*/;
  assign _4284_ = inv_16[43] & r_15[43] /*302*/;
  assign _4285_ = _4283_ | _4284_ /*301*/;
  assign _4286_ = inv_16[44] ^ r_15[44] /*299*/;
  assign sum_16[44] = _4286_ ^ _4285_ /*298*/;
  assign _4287_ = _4286_ & _4285_ /*297*/;
  assign _4288_ = inv_16[44] & r_15[44] /*296*/;
  assign _4289_ = _4287_ | _4288_ /*295*/;
  assign _4290_ = inv_16[45] ^ r_15[45] /*293*/;
  assign sum_16[45] = _4290_ ^ _4289_ /*292*/;
  assign _4291_ = _4290_ & _4289_ /*291*/;
  assign _4292_ = inv_16[45] & r_15[45] /*290*/;
  assign _4293_ = _4291_ | _4292_ /*289*/;
  assign _4294_ = _4293_ ^ _4289_ /*288*/;
  assign _4295_ = ~_4294_ /*287*/;
  assign _4296_ = sum_16[45] & _4295_ /*286*/;
  assign _4297_ = _4294_ & _4293_ /*285*/;
  assign sum_16[46] = _4297_ | _4296_ /*284*/;
  assign q[0] = ~sum_16[46] /*283*/;
  assign m_16[0] = r_15[0] /*282*/;
  assign m_16[1] = r_15[1] /*281*/;
  assign m_16[2] = r_15[2] /*280*/;
  assign m_16[3] = r_15[3] /*279*/;
  assign m_16[4] = r_15[4] /*278*/;
  assign m_16[5] = r_15[5] /*277*/;
  assign m_16[6] = r_15[6] /*276*/;
  assign m_16[7] = r_15[7] /*275*/;
  assign m_16[8] = r_15[8] /*274*/;
  assign m_16[9] = r_15[9] /*273*/;
  assign m_16[10] = r_15[10] /*272*/;
  assign m_16[11] = r_15[11] /*271*/;
  assign m_16[12] = r_15[12] /*270*/;
  assign m_16[13] = r_15[13] /*269*/;
  assign m_16[14] = r_15[14] /*268*/;
  assign m_16[15] = r_15[15] /*267*/;
  assign m_16[16] = r_15[16] /*266*/;
  assign m_16[17] = r_15[17] /*265*/;
  assign m_16[18] = r_15[18] /*264*/;
  assign m_16[19] = r_15[19] /*263*/;
  assign m_16[20] = r_15[20] /*262*/;
  assign m_16[21] = r_15[21] /*261*/;
  assign m_16[22] = r_15[22] /*260*/;
  assign m_16[23] = r_15[23] /*259*/;
  assign m_16[24] = r_15[24] /*258*/;
  assign m_16[25] = r_15[25] /*257*/;
  assign m_16[26] = r_15[26] /*256*/;
  assign m_16[27] = r_15[27] /*255*/;
  assign m_16[28] = r_15[28] /*254*/;
  assign m_16[29] = r_15[29] /*253*/;
  assign m_16[30] = r_15[30] /*252*/;
  assign m_16[31] = r_15[31] /*251*/;
  assign m_16[32] = r_15[32] /*250*/;
  assign m_16[33] = r_15[33] /*249*/;
  assign m_16[34] = r_15[34] /*248*/;
  assign m_16[35] = r_15[35] /*247*/;
  assign m_16[36] = r_15[36] /*246*/;
  assign m_16[37] = r_15[37] /*245*/;
  assign m_16[38] = r_15[38] /*244*/;
  assign m_16[39] = r_15[39] /*243*/;
  assign m_16[40] = r_15[40] /*242*/;
  assign m_16[41] = r_15[41] /*241*/;
  assign m_16[42] = r_15[42] /*240*/;
  assign m_16[43] = r_15[43] /*239*/;
  assign m_16[44] = r_15[44] /*238*/;
  assign m_16[45] = r_15[45] /*237*/;
  assign m_16[46] = r_15[45] /*236*/;
  assign _4299_ = ~q[0] /*235*/;
  assign _4300_ = sum_16[0] & q[0] /*234*/;
  assign _4301_ = m_16[0] & _4299_ /*233*/;
  assign r_16[0] = _4301_ | _4300_ /*232*/;
  assign _4302_ = ~q[0] /*231*/;
  assign _4303_ = sum_16[1] & q[0] /*230*/;
  assign _4304_ = m_16[1] & _4302_ /*229*/;
  assign r_16[1] = _4304_ | _4303_ /*228*/;
  assign _4305_ = ~q[0] /*227*/;
  assign _4306_ = sum_16[2] & q[0] /*226*/;
  assign _4307_ = m_16[2] & _4305_ /*225*/;
  assign r_16[2] = _4307_ | _4306_ /*224*/;
  assign _4308_ = ~q[0] /*223*/;
  assign _4309_ = sum_16[3] & q[0] /*222*/;
  assign _4310_ = m_16[3] & _4308_ /*221*/;
  assign r_16[3] = _4310_ | _4309_ /*220*/;
  assign _4311_ = ~q[0] /*219*/;
  assign _4312_ = sum_16[4] & q[0] /*218*/;
  assign _4313_ = m_16[4] & _4311_ /*217*/;
  assign r_16[4] = _4313_ | _4312_ /*216*/;
  assign _4314_ = ~q[0] /*215*/;
  assign _4315_ = sum_16[5] & q[0] /*214*/;
  assign _4316_ = m_16[5] & _4314_ /*213*/;
  assign r_16[5] = _4316_ | _4315_ /*212*/;
  assign _4317_ = ~q[0] /*211*/;
  assign _4318_ = sum_16[6] & q[0] /*210*/;
  assign _4319_ = m_16[6] & _4317_ /*209*/;
  assign r_16[6] = _4319_ | _4318_ /*208*/;
  assign _4320_ = ~q[0] /*207*/;
  assign _4321_ = sum_16[7] & q[0] /*206*/;
  assign _4322_ = m_16[7] & _4320_ /*205*/;
  assign r_16[7] = _4322_ | _4321_ /*204*/;
  assign _4323_ = ~q[0] /*203*/;
  assign _4324_ = sum_16[8] & q[0] /*202*/;
  assign _4325_ = m_16[8] & _4323_ /*201*/;
  assign r_16[8] = _4325_ | _4324_ /*200*/;
  assign _4326_ = ~q[0] /*199*/;
  assign _4327_ = sum_16[9] & q[0] /*198*/;
  assign _4328_ = m_16[9] & _4326_ /*197*/;
  assign r_16[9] = _4328_ | _4327_ /*196*/;
  assign _4329_ = ~q[0] /*195*/;
  assign _4330_ = sum_16[10] & q[0] /*194*/;
  assign _4331_ = m_16[10] & _4329_ /*193*/;
  assign r_16[10] = _4331_ | _4330_ /*192*/;
  assign _4332_ = ~q[0] /*191*/;
  assign _4333_ = sum_16[11] & q[0] /*190*/;
  assign _4334_ = m_16[11] & _4332_ /*189*/;
  assign r_16[11] = _4334_ | _4333_ /*188*/;
  assign _4335_ = ~q[0] /*187*/;
  assign _4336_ = sum_16[12] & q[0] /*186*/;
  assign _4337_ = m_16[12] & _4335_ /*185*/;
  assign r_16[12] = _4337_ | _4336_ /*184*/;
  assign _4338_ = ~q[0] /*183*/;
  assign _4339_ = sum_16[13] & q[0] /*182*/;
  assign _4340_ = m_16[13] & _4338_ /*181*/;
  assign r_16[13] = _4340_ | _4339_ /*180*/;
  assign _4341_ = ~q[0] /*179*/;
  assign _4342_ = sum_16[14] & q[0] /*178*/;
  assign _4343_ = m_16[14] & _4341_ /*177*/;
  assign r_16[14] = _4343_ | _4342_ /*176*/;
  assign _4344_ = ~q[0] /*175*/;
  assign _4345_ = sum_16[15] & q[0] /*174*/;
  assign _4346_ = m_16[15] & _4344_ /*173*/;
  assign r_16[15] = _4346_ | _4345_ /*172*/;
  assign _4347_ = ~q[0] /*171*/;
  assign _4348_ = sum_16[16] & q[0] /*170*/;
  assign _4349_ = m_16[16] & _4347_ /*169*/;
  assign r_16[16] = _4349_ | _4348_ /*168*/;
  assign _4350_ = ~q[0] /*167*/;
  assign _4351_ = sum_16[17] & q[0] /*166*/;
  assign _4352_ = m_16[17] & _4350_ /*165*/;
  assign r_16[17] = _4352_ | _4351_ /*164*/;
  assign _4353_ = ~q[0] /*163*/;
  assign _4354_ = sum_16[18] & q[0] /*162*/;
  assign _4355_ = m_16[18] & _4353_ /*161*/;
  assign r_16[18] = _4355_ | _4354_ /*160*/;
  assign _4356_ = ~q[0] /*159*/;
  assign _4357_ = sum_16[19] & q[0] /*158*/;
  assign _4358_ = m_16[19] & _4356_ /*157*/;
  assign r_16[19] = _4358_ | _4357_ /*156*/;
  assign _4359_ = ~q[0] /*155*/;
  assign _4360_ = sum_16[20] & q[0] /*154*/;
  assign _4361_ = m_16[20] & _4359_ /*153*/;
  assign r_16[20] = _4361_ | _4360_ /*152*/;
  assign _4362_ = ~q[0] /*151*/;
  assign _4363_ = sum_16[21] & q[0] /*150*/;
  assign _4364_ = m_16[21] & _4362_ /*149*/;
  assign r_16[21] = _4364_ | _4363_ /*148*/;
  assign _4365_ = ~q[0] /*147*/;
  assign _4366_ = sum_16[22] & q[0] /*146*/;
  assign _4367_ = m_16[22] & _4365_ /*145*/;
  assign r_16[22] = _4367_ | _4366_ /*144*/;
  assign _4368_ = ~q[0] /*143*/;
  assign _4369_ = sum_16[23] & q[0] /*142*/;
  assign _4370_ = m_16[23] & _4368_ /*141*/;
  assign r_16[23] = _4370_ | _4369_ /*140*/;
  assign _4371_ = ~q[0] /*139*/;
  assign _4372_ = sum_16[24] & q[0] /*138*/;
  assign _4373_ = m_16[24] & _4371_ /*137*/;
  assign r_16[24] = _4373_ | _4372_ /*136*/;
  assign _4374_ = ~q[0] /*135*/;
  assign _4375_ = sum_16[25] & q[0] /*134*/;
  assign _4376_ = m_16[25] & _4374_ /*133*/;
  assign r_16[25] = _4376_ | _4375_ /*132*/;
  assign _4377_ = ~q[0] /*131*/;
  assign _4378_ = sum_16[26] & q[0] /*130*/;
  assign _4379_ = m_16[26] & _4377_ /*129*/;
  assign r_16[26] = _4379_ | _4378_ /*128*/;
  assign _4380_ = ~q[0] /*127*/;
  assign _4381_ = sum_16[27] & q[0] /*126*/;
  assign _4382_ = m_16[27] & _4380_ /*125*/;
  assign r_16[27] = _4382_ | _4381_ /*124*/;
  assign _4383_ = ~q[0] /*123*/;
  assign _4384_ = sum_16[28] & q[0] /*122*/;
  assign _4385_ = m_16[28] & _4383_ /*121*/;
  assign r_16[28] = _4385_ | _4384_ /*120*/;
  assign _4386_ = ~q[0] /*119*/;
  assign _4387_ = sum_16[29] & q[0] /*118*/;
  assign _4388_ = m_16[29] & _4386_ /*117*/;
  assign r_16[29] = _4388_ | _4387_ /*116*/;
  assign _4389_ = ~q[0] /*115*/;
  assign _4390_ = sum_16[30] & q[0] /*114*/;
  assign _4391_ = m_16[30] & _4389_ /*113*/;
  assign r_16[30] = _4391_ | _4390_ /*112*/;
  assign _4392_ = ~q[0] /*111*/;
  assign _4393_ = sum_16[31] & q[0] /*110*/;
  assign _4394_ = m_16[31] & _4392_ /*109*/;
  assign r_16[31] = _4394_ | _4393_ /*108*/;
  assign _4395_ = ~q[0] /*107*/;
  assign _4396_ = sum_16[32] & q[0] /*106*/;
  assign _4397_ = m_16[32] & _4395_ /*105*/;
  assign r_16[32] = _4397_ | _4396_ /*104*/;
  assign _4398_ = ~q[0] /*103*/;
  assign _4399_ = sum_16[33] & q[0] /*102*/;
  assign _4400_ = m_16[33] & _4398_ /*101*/;
  assign r_16[33] = _4400_ | _4399_ /*100*/;
  assign _4401_ = ~q[0] /*99*/;
  assign _4402_ = sum_16[34] & q[0] /*98*/;
  assign _4403_ = m_16[34] & _4401_ /*97*/;
  assign r_16[34] = _4403_ | _4402_ /*96*/;
  assign _4404_ = ~q[0] /*95*/;
  assign _4405_ = sum_16[35] & q[0] /*94*/;
  assign _4406_ = m_16[35] & _4404_ /*93*/;
  assign r_16[35] = _4406_ | _4405_ /*92*/;
  assign _4407_ = ~q[0] /*91*/;
  assign _4408_ = sum_16[36] & q[0] /*90*/;
  assign _4409_ = m_16[36] & _4407_ /*89*/;
  assign r_16[36] = _4409_ | _4408_ /*88*/;
  assign _4410_ = ~q[0] /*87*/;
  assign _4411_ = sum_16[37] & q[0] /*86*/;
  assign _4412_ = m_16[37] & _4410_ /*85*/;
  assign r_16[37] = _4412_ | _4411_ /*84*/;
  assign _4413_ = ~q[0] /*83*/;
  assign _4414_ = sum_16[38] & q[0] /*82*/;
  assign _4415_ = m_16[38] & _4413_ /*81*/;
  assign r_16[38] = _4415_ | _4414_ /*80*/;
  assign _4416_ = ~q[0] /*79*/;
  assign _4417_ = sum_16[39] & q[0] /*78*/;
  assign _4418_ = m_16[39] & _4416_ /*77*/;
  assign r_16[39] = _4418_ | _4417_ /*76*/;
  assign _4419_ = ~q[0] /*75*/;
  assign _4420_ = sum_16[40] & q[0] /*74*/;
  assign _4421_ = m_16[40] & _4419_ /*73*/;
  assign r_16[40] = _4421_ | _4420_ /*72*/;
  assign _4422_ = ~q[0] /*71*/;
  assign _4423_ = sum_16[41] & q[0] /*70*/;
  assign _4424_ = m_16[41] & _4422_ /*69*/;
  assign r_16[41] = _4424_ | _4423_ /*68*/;
  assign _4425_ = ~q[0] /*67*/;
  assign _4426_ = sum_16[42] & q[0] /*66*/;
  assign _4427_ = m_16[42] & _4425_ /*65*/;
  assign r_16[42] = _4427_ | _4426_ /*64*/;
  assign _4428_ = ~q[0] /*63*/;
  assign _4429_ = sum_16[43] & q[0] /*62*/;
  assign _4430_ = m_16[43] & _4428_ /*61*/;
  assign r_16[43] = _4430_ | _4429_ /*60*/;
  assign _4431_ = ~q[0] /*59*/;
  assign _4432_ = sum_16[44] & q[0] /*58*/;
  assign _4433_ = m_16[44] & _4431_ /*57*/;
  assign r_16[44] = _4433_ | _4432_ /*56*/;
  assign _4434_ = ~q[0] /*55*/;
  assign _4435_ = sum_16[45] & q[0] /*54*/;
  assign _4436_ = m_16[45] & _4434_ /*53*/;
  assign r_16[45] = _4436_ | _4435_ /*52*/;
  assign _4437_ = ~q[0] /*51*/;
  assign _4438_ = sum_16[46] & q[0] /*50*/;
  assign _4439_ = m_16[46] & _4437_ /*49*/;
  assign r_16[46] = _4439_ | _4438_ /*48*/;
  assign rout[0] = r_16[0] /*0*/;
  assign rout[1] = r_16[1] /*1*/;
  assign rout[2] = r_16[2] /*2*/;
  assign rout[3] = r_16[3] /*3*/;
  assign rout[4] = r_16[4] /*4*/;
  assign rout[5] = r_16[5] /*5*/;
  assign rout[6] = r_16[6] /*6*/;
  assign rout[7] = r_16[7] /*7*/;
  assign rout[8] = r_16[8] /*8*/;
  assign rout[9] = r_16[9] /*9*/;
  assign rout[10] = r_16[10] /*10*/;
  assign rout[11] = r_16[11] /*11*/;
  assign rout[12] = r_16[12] /*12*/;
  assign rout[13] = r_16[13] /*13*/;
  assign rout[14] = r_16[14] /*14*/;
  assign rout[15] = r_16[15] /*15*/;
  assign rout[16] = r_16[16] /*16*/;
  assign rout[17] = r_16[17] /*17*/;
  assign rout[18] = r_16[18] /*18*/;
  assign rout[19] = r_16[19] /*19*/;
  assign rout[20] = r_16[20] /*20*/;
  assign rout[21] = r_16[21] /*21*/;
  assign rout[22] = r_16[22] /*22*/;
  assign rout[23] = r_16[23] /*23*/;
  assign rout[24] = r_16[24] /*24*/;
  assign rout[25] = r_16[25] /*25*/;
  assign rout[26] = r_16[26] /*26*/;
  assign rout[27] = r_16[27] /*27*/;
  assign rout[28] = r_16[28] /*28*/;
  assign rout[29] = r_16[29] /*29*/;
  assign rout[30] = r_16[30] /*30*/;
  assign rout[31] = r_16[31] /*31*/;
  assign rout[32] = r_16[32] /*32*/;
  assign rout[33] = r_16[33] /*33*/;
  assign rout[34] = r_16[34] /*34*/;
  assign rout[35] = r_16[35] /*35*/;
  assign rout[36] = r_16[36] /*36*/;
  assign rout[37] = r_16[37] /*37*/;
  assign rout[38] = r_16[38] /*38*/;
  assign rout[39] = r_16[39] /*39*/;
  assign rout[40] = r_16[40] /*40*/;
  assign rout[41] = r_16[41] /*41*/;
  assign rout[42] = r_16[42] /*42*/;
  assign rout[43] = r_16[43] /*43*/;
  assign rout[44] = r_16[44] /*44*/;
  assign rout[45] = r_16[45] /*45*/;
  assign rout[46] = r_16[46] /*46*/;
endmodule