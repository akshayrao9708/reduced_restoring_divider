module divider(q, rout, rin, div);
  wire _0_;
  wire _1_;
  wire _2_;
  wire _3_;
  wire _4_;
  wire _5_;
  wire _6_;
  wire _7_;
  wire _8_;
  wire _9_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  wire _38_;
  wire _39_;
  wire _40_;
  wire _41_;
  wire _42_;
  wire _43_;
  wire _44_;
  wire _45_;
  wire _46_;
  wire _47_;
  wire _48_;
  wire _49_;
  wire _50_;
  wire _51_;
  wire _52_;
  wire _53_;
  wire _54_;
  wire _55_;
  wire _56_;
  wire _57_;
  wire _58_;
  wire _59_;
  wire _60_;
  wire _61_;
  wire _62_;
  wire _63_;
  wire _64_;
  wire _65_;
  wire _66_;
  wire _67_;
  wire _68_;
  wire _69_;
  wire _70_;
  wire _71_;
  wire [2:0] r_0;
  wire [3:0] r_1;
  wire [3:0] m_1;
  wire [3:0] sum_1;
  wire [2:0] inv_1;
  wire [4:0] r_2;
  wire [4:0] m_2;
  wire [4:0] sum_2;
  wire [3:0] inv_2;
  wire zeroWire;
  wire oneWire;
  input [1:0] rin;
  input [0:0] div;
  output [1:0] q;
  output [4:0] rout;
  assign zeroWire = 1'b0 /*0*/;
  assign oneWire = 1'b1 /*0*/;
  assign r_0[0] = rin[0] /*194*/;
  assign r_0[1] = rin[1] /*193*/;
  assign r_0[2] = zeroWire /*192*/;
  assign inv_1[0] = oneWire /*116*/;
  assign inv_1[1] = ~div[0] /*110*/;
  assign inv_1[2] = oneWire /*104*/;
  assign _0_ = inv_1[0] ^ r_0[0] /*115*/;
  assign sum_1[0] = _0_ ^ oneWire /*114*/;
  assign _1_ = _0_ & oneWire /*113*/;
  assign _2_ = inv_1[0] & r_0[0] /*112*/;
  assign _3_ = _1_ | _2_ /*111*/;
  assign _4_ = inv_1[1] ^ r_0[1] /*109*/;
  assign sum_1[1] = _4_ ^ _3_ /*108*/;
  assign _5_ = _4_ & _3_ /*107*/;
  assign _6_ = inv_1[1] & r_0[1] /*106*/;
  assign _7_ = _5_ | _6_ /*105*/;
  assign _8_ = inv_1[2] ^ r_0[2] /*103*/;
  assign sum_1[2] = _8_ ^ _7_ /*102*/;
  assign _9_ = _8_ & _7_ /*101*/;
  assign _10_ = inv_1[2] & r_0[2] /*100*/;
  assign _11_ = _9_ | _10_ /*99*/;
  assign _12_ = _11_ ^ _7_ /*98*/;
  assign _13_ = ~_12_ /*97*/;
  assign _14_ = sum_1[2] & _13_ /*96*/;
  assign _15_ = _12_ & _11_ /*95*/;
  assign sum_1[3] = _15_ | _14_ /*94*/;
  assign q[1] = ~sum_1[3] /*93*/;
  assign m_1[0] = r_0[0] /*92*/;
  assign m_1[1] = r_0[1] /*91*/;
  assign m_1[2] = r_0[2] /*90*/;
  assign m_1[3] = r_0[2] /*89*/;
  assign _17_ = ~q[1] /*88*/;
  assign _18_ = sum_1[0] & q[1] /*87*/;
  assign _19_ = m_1[0] & _17_ /*86*/;
  assign r_1[0] = _19_ | _18_ /*85*/;
  assign _20_ = ~q[1] /*84*/;
  assign _21_ = sum_1[1] & q[1] /*83*/;
  assign _22_ = m_1[1] & _20_ /*82*/;
  assign r_1[1] = _22_ | _21_ /*81*/;
  assign _23_ = ~q[1] /*80*/;
  assign _24_ = sum_1[2] & q[1] /*79*/;
  assign _25_ = m_1[2] & _23_ /*78*/;
  assign r_1[2] = _25_ | _24_ /*77*/;
  assign _26_ = ~q[1] /*76*/;
  assign _27_ = sum_1[3] & q[1] /*75*/;
  assign _28_ = m_1[3] & _26_ /*74*/;
  assign r_1[3] = _28_ | _27_ /*73*/;
  assign inv_2[0] = ~div[0] /*60*/;
  assign inv_2[1] = oneWire /*54*/;
  assign inv_2[2] = oneWire /*48*/;
  assign inv_2[3] = oneWire /*42*/;
  assign _29_ = inv_2[0] ^ r_1[0] /*59*/;
  assign sum_2[0] = _29_ ^ oneWire /*58*/;
  assign _30_ = _29_ & oneWire /*57*/;
  assign _31_ = inv_2[0] & r_1[0] /*56*/;
  assign _32_ = _30_ | _31_ /*55*/;
  assign _33_ = inv_2[1] ^ r_1[1] /*53*/;
  assign sum_2[1] = _33_ ^ _32_ /*52*/;
  assign _34_ = _33_ & _32_ /*51*/;
  assign _35_ = inv_2[1] & r_1[1] /*50*/;
  assign _36_ = _34_ | _35_ /*49*/;
  assign _37_ = inv_2[2] ^ r_1[2] /*47*/;
  assign sum_2[2] = _37_ ^ _36_ /*46*/;
  assign _38_ = _37_ & _36_ /*45*/;
  assign _39_ = inv_2[2] & r_1[2] /*44*/;
  assign _40_ = _38_ | _39_ /*43*/;
  assign _41_ = inv_2[3] ^ r_1[3] /*41*/;
  assign sum_2[3] = _41_ ^ _40_ /*40*/;
  assign _42_ = _41_ & _40_ /*39*/;
  assign _43_ = inv_2[3] & r_1[3] /*38*/;
  assign _44_ = _42_ | _43_ /*37*/;
  assign _45_ = _44_ ^ _40_ /*36*/;
  assign _46_ = ~_45_ /*35*/;
  assign _47_ = sum_2[3] & _46_ /*34*/;
  assign _48_ = _45_ & _44_ /*33*/;
  assign sum_2[4] = _48_ | _47_ /*32*/;
  assign q[0] = ~sum_2[4] /*31*/;
  assign m_2[0] = r_1[0] /*30*/;
  assign m_2[1] = r_1[1] /*29*/;
  assign m_2[2] = r_1[2] /*28*/;
  assign m_2[3] = r_1[3] /*27*/;
  assign m_2[4] = r_1[3] /*26*/;
  assign _50_ = ~q[0] /*25*/;
  assign _51_ = sum_2[0] & q[0] /*24*/;
  assign _52_ = m_2[0] & _50_ /*23*/;
  assign r_2[0] = _52_ | _51_ /*22*/;
  assign _53_ = ~q[0] /*21*/;
  assign _54_ = sum_2[1] & q[0] /*20*/;
  assign _55_ = m_2[1] & _53_ /*19*/;
  assign r_2[1] = _55_ | _54_ /*18*/;
  assign _56_ = ~q[0] /*17*/;
  assign _57_ = sum_2[2] & q[0] /*16*/;
  assign _58_ = m_2[2] & _56_ /*15*/;
  assign r_2[2] = _58_ | _57_ /*14*/;
  assign _59_ = ~q[0] /*13*/;
  assign _60_ = sum_2[3] & q[0] /*12*/;
  assign _61_ = m_2[3] & _59_ /*11*/;
  assign r_2[3] = _61_ | _60_ /*10*/;
  assign _62_ = ~q[0] /*9*/;
  assign _63_ = sum_2[4] & q[0] /*8*/;
  assign _64_ = m_2[4] & _62_ /*7*/;
  assign r_2[4] = _64_ | _63_ /*6*/;
  assign rout[0] = r_2[0] /*0*/;
  assign rout[1] = r_2[1] /*1*/;
  assign rout[2] = r_2[2] /*2*/;
  assign rout[3] = r_2[3] /*3*/;
  assign rout[4] = r_2[4] /*4*/;
endmodule