module nonresdivReduced(R_0, D, Q, R_n1);
input [29:0] R_0;
input [14:0] D;
output [15:0] Q;
output [14:0] R_n1;
wire _0_;
wire _1_;
wire _2_;
wire _3_;
wire _4_;
wire _5_;
wire _6_;
wire _7_;
wire _8_;
wire _9_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire _30_;
wire _31_;
wire _32_;
wire _33_;
wire _34_;
wire _35_;
wire _36_;
wire _37_;
wire _38_;
wire _39_;
wire _40_;
wire _41_;
wire _42_;
wire _43_;
wire _44_;
wire _45_;
wire _46_;
wire _47_;
wire _48_;
wire _49_;
wire _50_;
wire _51_;
wire _52_;
wire _53_;
wire _54_;
wire _55_;
wire _56_;
wire _57_;
wire _58_;
wire _59_;
wire _60_;
wire _61_;
wire _62_;
wire _63_;
wire _64_;
wire _65_;
wire _66_;
wire _67_;
wire _68_;
wire _69_;
wire _70_;
wire _71_;
wire _72_;
wire _73_;
wire _74_;
wire _75_;
wire _76_;
wire _77_;
wire _78_;
wire _79_;
wire _80_;
wire _81_;
wire _82_;
wire _83_;
wire _84_;
wire _85_;
wire _86_;
wire _87_;
wire _88_;
wire _89_;
wire _90_;
wire _91_;
wire _92_;
wire _93_;
wire _94_;
wire _95_;
wire _96_;
wire _97_;
wire _98_;
wire _99_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
wire _255_;
wire _256_;
wire _257_;
wire _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire _267_;
wire _268_;
wire _269_;
wire _270_;
wire _271_;
wire _272_;
wire _273_;
wire _274_;
wire _275_;
wire _276_;
wire _277_;
wire _278_;
wire _279_;
wire _280_;
wire _281_;
wire _282_;
wire _283_;
wire _284_;
wire _285_;
wire _286_;
wire _287_;
wire _288_;
wire _289_;
wire _290_;
wire _291_;
wire _292_;
wire _293_;
wire _294_;
wire _295_;
wire _296_;
wire _297_;
wire _298_;
wire _299_;
wire _300_;
wire _301_;
wire _302_;
wire _303_;
wire _304_;
wire _305_;
wire _306_;
wire _307_;
wire _308_;
wire _309_;
wire _310_;
wire _311_;
wire _312_;
wire _313_;
wire _314_;
wire _315_;
wire _316_;
wire _317_;
wire _318_;
wire _319_;
wire _320_;
wire _321_;
wire _322_;
wire _323_;
wire _324_;
wire _325_;
wire _326_;
wire _327_;
wire _328_;
wire _329_;
wire _330_;
wire _331_;
wire _332_;
wire _333_;
wire _334_;
wire _335_;
wire _336_;
wire _337_;
wire _338_;
wire _339_;
wire _340_;
wire _341_;
wire _342_;
wire _343_;
wire _344_;
wire _345_;
wire _346_;
wire _347_;
wire _348_;
wire _349_;
wire _350_;
wire _351_;
wire _352_;
wire _353_;
wire _354_;
wire _355_;
wire _356_;
wire _357_;
wire _358_;
wire _359_;
wire _360_;
wire _361_;
wire _362_;
wire _363_;
wire _364_;
wire _365_;
wire _366_;
wire _367_;
wire _368_;
wire _369_;
wire _370_;
wire _371_;
wire _372_;
wire _373_;
wire _374_;
wire _375_;
wire _376_;
wire _377_;
wire _378_;
wire _379_;
wire _380_;
wire _381_;
wire _382_;
wire _383_;
wire _384_;
wire _385_;
wire _386_;
wire _387_;
wire _388_;
wire _389_;
wire _390_;
wire _391_;
wire _392_;
wire _393_;
wire _394_;
wire _395_;
wire _396_;
wire _397_;
wire _398_;
wire _399_;
wire _400_;
wire _401_;
wire _402_;
wire _403_;
wire _404_;
wire _405_;
wire _406_;
wire _407_;
wire _408_;
wire _409_;
wire _410_;
wire _411_;
wire _412_;
wire _413_;
wire _414_;
wire _415_;
wire _416_;
wire _417_;
wire _418_;
wire _419_;
wire _420_;
wire _421_;
wire _422_;
wire _423_;
wire _424_;
wire _425_;
wire _426_;
wire _427_;
wire _428_;
wire _429_;
wire _430_;
wire _431_;
wire _432_;
wire _433_;
wire _434_;
wire _435_;
wire _436_;
wire _437_;
wire _438_;
wire _439_;
wire _440_;
wire _441_;
wire _442_;
wire _443_;
wire _444_;
wire _445_;
wire _446_;
wire _447_;
wire _448_;
wire _449_;
wire _450_;
wire _451_;
wire _452_;
wire _453_;
wire _454_;
wire _455_;
wire _456_;
wire _457_;
wire _458_;
wire _459_;
wire _460_;
wire _461_;
wire _462_;
wire _463_;
wire _464_;
wire _465_;
wire _466_;
wire _467_;
wire _468_;
wire _469_;
wire _470_;
wire _471_;
wire _472_;
wire _473_;
wire _474_;
wire _475_;
wire _476_;
wire _477_;
wire _478_;
wire _479_;
wire _480_;
wire _481_;
wire _482_;
wire _483_;
wire _484_;
wire _485_;
wire _486_;
wire _487_;
wire _488_;
wire _489_;
wire _490_;
wire _491_;
wire _492_;
wire _493_;
wire _494_;
wire _495_;
wire _496_;
wire _497_;
wire _498_;
wire _499_;
wire _500_;
wire _501_;
wire _502_;
wire _503_;
wire _504_;
wire _505_;
wire _506_;
wire _507_;
wire _508_;
wire _509_;
wire _510_;
wire _511_;
wire _512_;
wire _513_;
wire _514_;
wire _515_;
wire _516_;
wire _517_;
wire _518_;
wire _519_;
wire _520_;
wire _521_;
wire _522_;
wire _523_;
wire _524_;
wire _525_;
wire _526_;
wire _527_;
wire _528_;
wire _529_;
wire _530_;
wire _531_;
wire _532_;
wire _533_;
wire _534_;
wire _535_;
wire _536_;
wire _537_;
wire _538_;
wire _539_;
wire _540_;
wire _541_;
wire _542_;
wire _543_;
wire _544_;
wire _545_;
wire _546_;
wire _547_;
wire _548_;
wire _549_;
wire _550_;
wire _551_;
wire _552_;
wire _553_;
wire _554_;
wire _555_;
wire _556_;
wire _557_;
wire _558_;
wire _559_;
wire _560_;
wire _561_;
wire _562_;
wire _563_;
wire _564_;
wire _565_;
wire _566_;
wire _567_;
wire _568_;
wire _569_;
wire _570_;
wire _571_;
wire _572_;
wire _573_;
wire _574_;
wire _575_;
wire _576_;
wire _577_;
wire _578_;
wire _579_;
wire _580_;
wire _581_;
wire _582_;
wire _583_;
wire _584_;
wire _585_;
wire _586_;
wire _587_;
wire _588_;
wire _589_;
wire _590_;
wire _591_;
wire _592_;
wire _593_;
wire _594_;
wire _595_;
wire _596_;
wire _597_;
wire _598_;
wire _599_;
wire _600_;
wire _601_;
wire _602_;
wire _603_;
wire _604_;
wire _605_;
wire _606_;
wire _607_;
wire _608_;
wire _609_;
wire _610_;
wire _611_;
wire _612_;
wire _613_;
wire _614_;
wire _615_;
wire _616_;
wire _617_;
wire _618_;
wire _619_;
wire _620_;
wire _621_;
wire _622_;
wire _623_;
wire _624_;
wire _625_;
wire _626_;
wire _627_;
wire _628_;
wire _629_;
wire _630_;
wire _631_;
wire _632_;
wire _633_;
wire _634_;
wire _635_;
wire _636_;
wire _637_;
wire _638_;
wire _639_;
wire _640_;
wire _641_;
wire _642_;
wire _643_;
wire _644_;
wire _645_;
wire _646_;
wire _647_;
wire _648_;
wire _649_;
wire _650_;
wire _651_;
wire _652_;
wire _653_;
wire _654_;
wire _655_;
wire _656_;
wire _657_;
wire _658_;
wire _659_;
wire _660_;
wire _661_;
wire _662_;
wire _663_;
wire _664_;
wire _665_;
wire _666_;
wire _667_;
wire _668_;
wire _669_;
wire _670_;
wire _671_;
wire _672_;
wire _673_;
wire _674_;
wire _675_;
wire _676_;
wire _677_;
wire _678_;
wire _679_;
wire _680_;
wire _681_;
wire _682_;
wire _683_;
wire _684_;
wire _685_;
wire _686_;
wire _687_;
wire _688_;
wire _689_;
wire _690_;
wire _691_;
wire _692_;
wire _693_;
wire _694_;
wire _695_;
wire _696_;
wire _697_;
wire _698_;
wire _699_;
wire _700_;
wire _701_;
wire _702_;
wire _703_;
wire _704_;
wire _705_;
wire _706_;
wire _707_;
wire _708_;
wire _709_;
wire _710_;
wire _711_;
wire _712_;
wire _713_;
wire _714_;
wire _715_;
wire _716_;
wire _717_;
wire _718_;
wire _719_;
wire _720_;
wire _721_;
wire _722_;
wire _723_;
wire _724_;
wire _725_;
wire _726_;
wire _727_;
wire _728_;
wire _729_;
wire _730_;
wire _731_;
wire _732_;
wire _733_;
wire _734_;
wire _735_;
wire _736_;
wire _737_;
wire _738_;
wire _739_;
wire _740_;
wire _741_;
wire _742_;
wire _743_;
wire _744_;
wire _745_;
wire _746_;
wire _747_;
wire _748_;
wire _749_;
wire _750_;
wire _751_;
wire _752_;
wire _753_;
wire _754_;
wire _755_;
wire _756_;
wire _757_;
wire _758_;
wire _759_;
wire _760_;
wire _761_;
wire _762_;
wire _763_;
wire _764_;
wire _765_;
wire _766_;
wire _767_;
wire _768_;
wire _769_;
wire _770_;
wire _771_;
wire _772_;
wire _773_;
wire _774_;
wire _775_;
wire _776_;
wire _777_;
wire _778_;
wire _779_;
wire _780_;
wire _781_;
wire _782_;
wire _783_;
wire _784_;
wire _785_;
wire _786_;
wire _787_;
wire _788_;
wire _789_;
wire _790_;
wire _791_;
wire _792_;
wire _793_;
wire _794_;
wire _795_;
wire _796_;
wire _797_;
wire _798_;
wire _799_;
wire _800_;
wire _801_;
wire _802_;
wire _803_;
wire _804_;
wire _805_;
wire _806_;
wire _807_;
wire _808_;
wire _809_;
wire _810_;
wire _811_;
wire _812_;
wire _813_;
wire _814_;
wire _815_;
wire _816_;
wire _817_;
wire _818_;
wire _819_;
wire _820_;
wire _821_;
wire _822_;
wire _823_;
wire _824_;
wire _825_;
wire _826_;
wire _827_;
wire _828_;
wire _829_;
wire _830_;
wire _831_;
wire _832_;
wire _833_;
wire _834_;
wire _835_;
wire _836_;
wire _837_;
wire _838_;
wire _839_;
wire _840_;
wire _841_;
wire _842_;
wire _843_;
wire _844_;
wire _845_;
wire _846_;
wire _847_;
wire _848_;
wire _849_;
wire _850_;
wire _851_;
wire _852_;
wire _853_;
wire _854_;
wire _855_;
wire _856_;
wire _857_;
wire _858_;
wire _859_;
wire _860_;
wire _861_;
wire _862_;
wire _863_;
wire _864_;
wire _865_;
wire _866_;
wire _867_;
wire _868_;
wire _869_;
wire _870_;
wire _871_;
wire _872_;
wire _873_;
wire _874_;
wire _875_;
wire _876_;
wire _877_;
wire _878_;
wire _879_;
wire _880_;
wire _881_;
wire _882_;
wire _883_;
wire _884_;
wire _885_;
wire _886_;
wire _887_;
wire _888_;
wire _889_;
wire _890_;
wire _891_;
wire _892_;
wire _893_;
wire _894_;
wire _895_;
wire _896_;
wire _897_;
wire _898_;
wire _899_;
wire _900_;
wire _901_;
wire _902_;
wire _903_;
wire _904_;
wire _905_;
wire _906_;
wire _907_;
wire _908_;
wire _909_;
wire _910_;
wire _911_;
wire _912_;
wire _913_;
wire _914_;
wire _915_;
wire _916_;
wire _917_;
wire _918_;
wire _919_;
wire _920_;
wire _921_;
wire _922_;
wire _923_;
wire _924_;
wire _925_;
wire _926_;
wire _927_;
wire _928_;
wire _929_;
wire _930_;
wire _931_;
wire _932_;
wire _933_;
wire _934_;
wire _935_;
wire _936_;
wire _937_;
wire _938_;
wire _939_;
wire _940_;
wire _941_;
wire _942_;
wire _943_;
wire _944_;
wire _945_;
wire _946_;
wire _947_;
wire _948_;
wire _949_;
wire _950_;
wire _951_;
wire _952_;
wire _953_;
wire _954_;
wire _955_;
wire _956_;
wire _957_;
wire _958_;
wire _959_;
wire _960_;
wire _961_;
wire _962_;
wire _963_;
wire _964_;
wire _965_;
wire _966_;
wire _967_;
wire _968_;
wire _969_;
wire _970_;
wire _971_;
wire _972_;
wire _973_;
wire _974_;
wire _975_;
wire _976_;
wire _977_;
wire _978_;
wire _979_;
wire _980_;
wire _981_;
wire _982_;
wire _983_;
wire _984_;
wire _985_;
wire _986_;
wire _987_;
wire _988_;
wire _989_;
wire _990_;
wire _991_;
wire _992_;
wire _993_;
wire _994_;
wire _995_;
wire _996_;
wire _997_;
wire _998_;
wire _999_;
wire _1000_;
wire _1001_;
wire _1002_;
wire _1003_;
wire _1004_;
wire _1005_;
wire _1006_;
wire _1007_;
wire _1008_;
wire _1009_;
wire _1010_;
wire _1011_;
wire _1012_;
wire _1013_;
wire _1014_;
wire _1015_;
wire _1016_;
wire _1017_;
wire _1018_;
wire _1019_;
wire _1020_;
wire _1021_;
wire _1022_;
wire _1023_;
wire _1024_;
wire _1025_;
wire _1026_;
wire _1027_;
wire _1028_;
wire _1029_;
wire _1030_;
wire _1031_;
wire _1032_;
wire _1033_;
wire _1034_;
wire _1035_;
wire _1036_;
wire _1037_;
wire _1038_;
wire _1039_;
wire _1040_;
wire _1041_;
wire _1042_;
wire _1043_;
wire _1044_;
wire _1045_;
wire _1046_;
wire _1047_;
wire _1048_;
wire _1049_;
wire _1050_;
wire _1051_;
wire _1052_;
wire _1053_;
wire _1054_;
wire _1055_;
wire _1056_;
wire _1057_;
wire _1058_;
wire _1059_;
wire _1060_;
wire _1061_;
wire _1062_;
wire _1063_;
wire _1064_;
wire _1065_;
wire _1066_;
wire _1067_;
wire _1068_;
wire _1069_;
wire _1070_;
wire _1071_;
wire _1072_;
wire _1073_;
wire _1074_;
wire _1075_;
wire _1076_;
wire _1077_;
wire _1078_;
wire _1079_;
wire _1080_;
wire _1081_;
wire _1082_;
wire _1083_;
wire _1084_;
wire _1085_;
wire _1086_;
wire _1087_;
wire _1088_;
wire _1089_;
wire _1090_;
wire _1091_;
wire _1092_;
wire _1093_;
wire _1094_;
wire _1095_;
wire _1096_;
wire _1097_;
wire _1098_;
wire _1099_;
wire _1100_;
wire _1101_;
wire _1102_;
wire _1103_;
wire _1104_;
wire _1105_;
wire _1106_;
wire _1107_;
wire _1108_;
wire _1109_;
wire _1110_;
wire _1111_;
wire _1112_;
wire _1113_;
wire _1114_;
wire _1115_;
wire _1116_;
wire _1117_;
wire _1118_;
wire _1119_;
wire _1120_;
wire _1121_;
wire _1122_;
wire _1123_;
wire _1124_;
wire _1125_;
wire _1126_;
wire _1127_;
wire _1128_;
wire _1129_;
wire _1130_;
wire _1131_;
wire _1132_;
wire _1133_;
wire _1134_;
wire _1135_;
wire _1136_;
wire _1137_;
wire _1138_;
wire _1139_;
wire _1140_;
wire _1141_;
wire _1142_;
wire _1143_;
wire _1144_;
wire _1145_;
wire _1146_;
wire _1147_;
wire _1148_;
wire _1149_;
wire _1150_;
wire _1151_;
wire _1152_;
wire _1153_;
wire _1154_;
wire _1155_;
wire _1156_;
wire _1157_;
wire _1158_;
wire _1159_;
wire _1160_;
wire _1161_;
wire _1162_;
wire _1163_;
wire _1164_;
wire _1165_;
wire _1166_;
wire _1167_;
wire _1168_;
wire _1169_;
wire _1170_;
wire _1171_;
wire _1172_;
wire _1173_;
wire _1174_;
wire _1175_;
wire _1176_;
wire _1177_;
wire _1178_;
wire _1179_;
wire _1180_;
wire _1181_;
wire _1182_;
wire _1183_;
wire _1184_;
wire _1185_;
wire _1186_;
wire _1187_;
wire _1188_;
wire _1189_;
wire _1190_;
wire _1191_;
wire _1192_;
wire _1193_;
wire _1194_;
wire _1195_;
wire _1196_;
wire _1197_;
wire _1198_;
wire _1199_;
wire _1200_;
wire _1201_;
wire _1202_;
wire _1203_;
wire _1204_;
wire _1205_;
wire _1206_;
wire _1207_;
wire _1208_;
wire _1209_;
wire _1210_;
wire _1211_;
wire _1212_;
wire _1213_;
wire _1214_;
wire _1215_;
wire _1216_;
wire _1217_;
wire _1218_;
wire _1219_;
wire _1220_;
wire _1221_;
wire _1222_;
wire _1223_;
wire _1224_;
wire _1225_;
wire _1226_;
wire _1227_;
wire _1228_;
wire _1229_;
wire _1230_;
wire _1231_;
wire _1232_;
wire _1233_;
wire _1234_;
wire _1235_;
wire _1236_;
wire _1237_;
wire _1238_;
wire _1239_;
wire _1240_;
wire _1241_;
wire _1242_;
wire _1243_;
wire _1244_;
wire _1245_;
wire _1246_;
wire _1247_;
wire _1248_;
wire _1249_;
wire _1250_;
wire _1251_;
wire _1252_;
wire _1253_;
wire _1254_;
wire _1255_;
wire _1256_;
wire _1257_;
wire _1258_;
wire _1259_;
wire _1260_;
wire _1261_;
wire _1262_;
wire _1263_;
wire _1264_;
wire _1265_;
wire _1266_;
wire _1267_;
wire _1268_;
wire _1269_;
wire _1270_;
wire _1271_;
wire _1272_;
wire _1273_;
wire _1274_;
wire _1275_;
wire _1276_;
wire _1277_;
wire _1278_;
wire _1279_;
wire _1280_;
wire _1281_;
wire _1282_;
wire _1283_;
wire _1284_;
wire _1285_;
wire _1286_;
wire _1287_;
wire _1288_;
wire _1289_;
wire _1290_;
wire _1291_;
wire _1292_;
wire _1293_;
wire _1294_;
wire _1295_;
wire _1296_;
wire _1297_;
wire _1298_;
wire _1299_;
wire _1300_;
wire _1301_;
wire _1302_;
wire _1303_;
wire _1304_;
wire _1305_;
wire _1306_;
wire _1307_;
wire _1308_;
wire _1309_;
wire _1310_;
wire _1311_;
wire _1312_;
wire _1313_;
wire _1314_;
wire _1315_;
wire _1316_;
wire _1317_;
wire _1318_;
wire _1319_;
wire _1320_;
wire _1321_;
wire _1322_;
wire _1323_;
wire _1324_;
wire _1325_;
wire _1326_;
wire _1327_;
wire _1328_;
wire _1329_;
wire _1330_;
wire _1331_;
wire _1332_;
wire _1333_;
wire _1334_;
wire _1335_;
wire _1336_;
wire _1337_;
wire _1338_;
wire _1339_;
wire _1340_;
wire _1341_;
wire _1342_;
wire _1343_;
wire _1344_;
wire _1345_;
wire _1346_;
wire _1347_;
wire _1348_;
wire _1349_;
wire _1350_;
wire _1351_;
wire _1352_;
wire _1353_;
wire _1354_;
wire _1355_;
wire _1356_;
wire _1357_;
wire _1358_;
wire _1359_;
wire _1360_;
wire _1361_;
wire _1362_;
wire _1363_;
wire _1364_;
wire _1365_;
wire _1366_;
wire _1367_;
wire _1368_;
wire _1369_;
wire _1370_;
wire _1371_;
wire _1372_;
wire _1373_;
wire _1374_;
wire _1375_;
wire _1376_;
wire _1377_;
wire _1378_;
wire _1379_;
wire _1380_;
wire _1381_;
wire _1382_;
wire _1383_;
wire _1384_;
wire _1385_;
wire _1386_;
wire _1387_;
wire _1388_;
wire _1389_;
wire _1390_;
wire _1391_;
wire _1392_;
wire _1393_;
wire _1394_;
wire _1395_;
wire _1396_;
wire _1397_;
wire _1398_;
wire _1399_;
wire _1400_;
wire _1401_;
wire _1402_;
wire _1403_;
wire _1404_;
wire _1405_;
wire _1406_;
wire _1407_;
wire _1408_;
wire _1409_;
wire _1410_;
wire _1411_;
wire _1412_;
wire _1413_;
wire _1414_;
wire _1415_;
wire _1416_;
wire _1417_;
wire _1418_;
wire _1419_;
wire _1420_;
wire _1421_;
wire _1422_;
wire _1423_;
wire _1424_;
wire _1425_;
wire _1426_;
wire _1427_;
wire _1428_;
wire _1429_;
wire _1430_;
wire _1431_;
wire _1432_;
wire _1433_;
wire _1434_;
wire _1435_;
wire _1436_;
wire _1437_;
wire _1438_;
wire _1439_;
wire _1440_;
wire _1441_;
wire _1442_;
wire _1443_;
wire _1444_;
wire _1445_;
wire _1446_;
wire _1447_;
wire _1448_;
wire _1449_;
wire _1450_;
wire _1451_;
wire _1452_;
wire _1453_;
wire _1454_;
wire _1455_;
wire _1456_;
wire _1457_;
wire _1458_;
wire _1459_;
wire _1460_;
wire _1461_;
wire _1462_;
wire _1463_;
wire _1464_;
wire _1465_;
wire _1466_;
wire _1467_;
wire _1468_;
wire _1469_;
wire _1470_;
wire _1471_;
wire _1472_;
wire _1473_;
wire _1474_;
wire _1475_;
wire _1476_;
wire _1477_;
wire _1478_;
wire _1479_;
wire _1480_;
wire _1481_;
wire _1482_;
wire _1483_;
wire _1484_;
wire _1485_;
wire _1486_;
wire _1487_;
wire _1488_;
wire _1489_;
wire _1490_;
wire _1491_;
wire _1492_;
wire _1493_;
wire _1494_;
wire _1495_;
wire _1496_;
wire _1497_;
wire _1498_;
wire _1499_;
wire _1500_;
wire _1501_;
wire _1502_;
wire _1503_;
wire _1504_;
wire _1505_;
wire _1506_;
wire _1507_;
wire _1508_;
wire _1509_;
wire _1510_;
wire _1511_;
wire _1512_;
wire _1513_;
wire _1514_;
wire _1515_;
wire _1516_;
wire _1517_;
wire _1518_;
wire _1519_;
wire _1520_;
wire _1521_;
wire _1522_;
wire _1523_;
wire _1524_;
wire _1525_;
wire _1526_;
wire _1527_;
wire _1528_;
wire _1529_;
wire _1530_;
wire _1531_;
wire _1532_;
wire _1533_;
wire _1534_;
wire _1535_;
wire _1536_;
wire _1537_;
wire _1538_;
wire _1539_;
wire _1540_;
wire _1541_;
wire _1542_;
wire _1543_;
wire _1544_;
wire _1545_;
wire _1546_;
wire _1547_;
wire _1548_;
wire _1549_;
wire _1550_;
wire _1551_;
wire _1552_;
wire _1553_;
wire _1554_;
wire _1555_;
wire _1556_;
wire _1557_;
wire _1558_;
wire _1559_;
wire _1560_;
wire _1561_;
wire _1562_;
wire _1563_;
wire _1564_;
wire _1565_;
wire _1566_;
wire _1567_;
wire _1568_;
wire _1569_;
wire _1570_;
wire _1571_;
wire _1572_;
wire _1573_;
wire _1574_;
wire _1575_;
wire _1576_;
wire _1577_;
wire _1578_;
wire _1579_;
wire _1580_;
wire _1581_;
wire _1582_;
wire _1583_;
wire _1584_;
wire _1585_;
wire _1586_;
wire _1587_;
wire _1588_;
wire _1589_;
wire _1590_;
wire _1591_;
wire _1592_;
wire _1593_;
wire _1594_;
wire _1595_;
wire _1596_;
wire _1597_;
wire _1598_;
wire _1599_;
wire _1600_;
wire _1601_;
wire _1602_;
wire _1603_;
wire _1604_;
wire _1605_;
wire _1606_;
wire _1607_;
wire _1608_;
wire _1609_;
wire _1610_;
wire _1611_;
wire _1612_;
wire _1613_;
wire _1614_;
wire _1615_;
wire _1616_;
wire _1617_;
wire _1618_;
wire _1619_;
wire _1620_;
wire _1621_;
wire _1622_;
wire _1623_;
wire _1624_;
wire _1625_;
wire _1626_;
wire _1627_;
wire _1628_;
wire _1629_;
wire _1630_;
wire _1631_;
wire _1632_;
wire _1633_;
wire _1634_;
wire _1635_;
wire _1636_;
wire _1637_;
wire _1638_;
wire _1639_;
wire _1640_;
wire _1641_;
wire _1642_;
wire _1643_;
wire _1644_;
wire _1645_;
wire _1646_;
wire _1647_;
wire _1648_;
wire _1649_;
wire _1650_;
wire _1651_;
wire _1652_;
wire _1653_;
wire _1654_;
wire _1655_;
wire _1656_;
wire _1657_;
wire _1658_;
wire _1659_;
wire _1660_;
wire _1661_;
wire _1662_;
wire _1663_;
wire _1664_;
wire _1665_;
wire _1666_;
wire _1667_;
wire _1668_;
wire _1669_;
wire _1670_;
wire _1671_;
wire _1672_;
wire _1673_;
wire _1674_;
wire _1675_;
wire _1676_;
wire _1677_;
wire _1678_;
wire _1679_;
wire _1680_;
wire _1681_;
wire _1682_;
wire _1683_;
wire _1684_;
wire _1685_;
wire _1686_;
wire _1687_;
wire _1688_;
wire _1689_;
wire _1690_;
wire _1691_;
wire _1692_;
wire _1693_;
wire _1694_;
wire _1695_;
wire _1696_;
wire _1697_;
wire _1698_;
wire _1699_;
wire _1700_;
wire _1701_;
wire _1702_;
wire _1703_;
wire _1704_;
wire _1705_;
wire _1706_;
wire _1707_;
wire _1708_;
wire _1709_;
wire _1710_;
wire _1711_;
wire _1712_;
wire _1713_;
wire _1714_;
wire _1715_;
wire _1716_;
wire _1717_;
wire _1718_;
wire _1719_;
wire _1720_;
wire _1721_;
wire _1722_;
wire _1723_;
wire _1724_;
wire _1725_;
wire _1726_;
wire _1727_;
wire _1728_;
wire _1729_;
wire _1730_;
wire _1731_;
wire _1732_;
wire _1733_;
wire _1734_;
wire _1735_;
wire _1736_;
wire _1737_;
wire _1738_;
wire _1739_;
wire _1740_;
wire _1741_;
wire _1742_;
wire _1743_;
wire _1744_;
wire _1745_;
wire _1746_;
wire _1747_;
wire _1748_;
wire _1749_;
wire _1750_;
wire _1751_;
wire _1752_;
wire _1753_;
wire _1754_;
wire _1755_;
wire _1756_;
wire _1757_;
wire _1758_;
wire _1759_;
wire _1760_;
wire _1761_;
wire _1762_;
wire _1763_;
wire _1764_;
wire _1765_;
wire _1766_;
wire _1767_;
wire _1768_;
wire _1769_;
wire _1770_;
wire _1771_;
wire _1772_;
wire _1773_;
wire _1774_;
wire _1775_;
wire _1776_;
wire _1777_;
wire _1778_;
wire _1779_;
wire _1780_;
wire _1781_;
wire _1782_;
wire _1783_;
wire _1784_;
wire _1785_;
wire _1786_;
wire _1787_;
wire _1788_;
wire _1789_;
wire _1790_;
wire _1791_;
wire _1792_;
wire _1793_;
wire _1794_;
wire _1795_;
wire _1796_;
wire _1797_;
wire _1798_;
wire _1799_;
wire _1800_;
wire _1801_;
wire _1802_;
wire _1803_;
wire _1804_;
wire _1805_;
wire _1806_;
wire _1807_;
wire _1808_;
wire _1809_;
wire _1810_;
wire _1811_;
wire _1812_;
wire _1813_;
wire _1814_;
wire _1815_;
wire _1816_;
wire _1817_;
wire _1818_;
wire _1819_;
wire _1820_;
wire _1821_;
wire _1822_;
wire _1823_;
wire _1824_;
wire _1825_;
wire _1826_;
wire _1827_;
wire _1828_;
wire _1829_;
wire _1830_;
wire _1831_;
wire _1832_;
wire _1833_;
wire _1834_;
wire _1835_;
wire _1836_;
wire _1837_;
wire _1838_;
wire _1839_;
wire _1840_;
wire _1841_;
wire _1842_;
wire _1843_;
wire _1844_;
wire _1845_;
wire _1846_;
wire _1847_;
wire _1848_;
wire _1849_;
wire _1850_;
wire _1851_;
wire _1852_;
wire _1853_;
wire _1854_;
wire _1855_;
wire _1856_;
wire _1857_;
wire _1858_;
wire _1859_;
wire _1860_;
wire _1861_;
wire _1862_;
wire _1863_;
wire _1864_;
wire _1865_;
wire _1866_;
wire _1867_;
wire _1868_;
wire _1869_;
wire _1870_;
wire zeroWire;
wire oneWire;
assign zeroWire = 1'b0 /*3339*/;
assign oneWire = 1'b1 /*3339*/;
assign _21_ = ~D[0] /*3241*/;
assign _18_ = R_0[15] & _21_ /*3237*/;
assign _19_ = R_0[15] ^ _21_ /*3240*/;
assign _20_ = oneWire & _19_ /*3238*/;
assign _0_ = oneWire ^ _19_ /*3239*/;
assign _17_ = _18_ | _20_ /*3236*/;
assign _26_ = ~D[1] /*3235*/;
assign _23_ = R_0[16] & _26_ /*3231*/;
assign _24_ = R_0[16] ^ _26_ /*3234*/;
assign _25_ = _17_ & _24_ /*3232*/;
assign _1_ = _17_ ^ _24_ /*3233*/;
assign _22_ = _23_ | _25_ /*3230*/;
assign _31_ = ~D[2] /*3229*/;
assign _28_ = R_0[17] & _31_ /*3225*/;
assign _29_ = R_0[17] ^ _31_ /*3228*/;
assign _30_ = _22_ & _29_ /*3226*/;
assign _2_ = _22_ ^ _29_ /*3227*/;
assign _27_ = _28_ | _30_ /*3224*/;
assign _36_ = ~D[3] /*3223*/;
assign _33_ = R_0[18] & _36_ /*3219*/;
assign _34_ = R_0[18] ^ _36_ /*3222*/;
assign _35_ = _27_ & _34_ /*3220*/;
assign _3_ = _27_ ^ _34_ /*3221*/;
assign _32_ = _33_ | _35_ /*3218*/;
assign _41_ = ~D[4] /*3217*/;
assign _38_ = R_0[19] & _41_ /*3213*/;
assign _39_ = R_0[19] ^ _41_ /*3216*/;
assign _40_ = _32_ & _39_ /*3214*/;
assign _4_ = _32_ ^ _39_ /*3215*/;
assign _37_ = _38_ | _40_ /*3212*/;
assign _46_ = ~D[5] /*3211*/;
assign _43_ = R_0[20] & _46_ /*3207*/;
assign _44_ = R_0[20] ^ _46_ /*3210*/;
assign _45_ = _37_ & _44_ /*3208*/;
assign _5_ = _37_ ^ _44_ /*3209*/;
assign _42_ = _43_ | _45_ /*3206*/;
assign _51_ = ~D[6] /*3205*/;
assign _48_ = R_0[21] & _51_ /*3201*/;
assign _49_ = R_0[21] ^ _51_ /*3204*/;
assign _50_ = _42_ & _49_ /*3202*/;
assign _6_ = _42_ ^ _49_ /*3203*/;
assign _47_ = _48_ | _50_ /*3200*/;
assign _56_ = ~D[7] /*3199*/;
assign _53_ = R_0[22] & _56_ /*3195*/;
assign _54_ = R_0[22] ^ _56_ /*3198*/;
assign _55_ = _47_ & _54_ /*3196*/;
assign _7_ = _47_ ^ _54_ /*3197*/;
assign _52_ = _53_ | _55_ /*3194*/;
assign _61_ = ~D[8] /*3193*/;
assign _58_ = R_0[23] & _61_ /*3189*/;
assign _59_ = R_0[23] ^ _61_ /*3192*/;
assign _60_ = _52_ & _59_ /*3190*/;
assign _8_ = _52_ ^ _59_ /*3191*/;
assign _57_ = _58_ | _60_ /*3188*/;
assign _66_ = ~D[9] /*3187*/;
assign _63_ = R_0[24] & _66_ /*3183*/;
assign _64_ = R_0[24] ^ _66_ /*3186*/;
assign _65_ = _57_ & _64_ /*3184*/;
assign _9_ = _57_ ^ _64_ /*3185*/;
assign _62_ = _63_ | _65_ /*3182*/;
assign _71_ = ~D[10] /*3181*/;
assign _68_ = R_0[25] & _71_ /*3177*/;
assign _69_ = R_0[25] ^ _71_ /*3180*/;
assign _70_ = _62_ & _69_ /*3178*/;
assign _10_ = _62_ ^ _69_ /*3179*/;
assign _67_ = _68_ | _70_ /*3176*/;
assign _76_ = ~D[11] /*3175*/;
assign _73_ = R_0[26] & _76_ /*3171*/;
assign _74_ = R_0[26] ^ _76_ /*3174*/;
assign _75_ = _67_ & _74_ /*3172*/;
assign _11_ = _67_ ^ _74_ /*3173*/;
assign _72_ = _73_ | _75_ /*3170*/;
assign _81_ = ~D[12] /*3169*/;
assign _78_ = R_0[27] & _81_ /*3165*/;
assign _79_ = R_0[27] ^ _81_ /*3168*/;
assign _80_ = _72_ & _79_ /*3166*/;
assign _12_ = _72_ ^ _79_ /*3167*/;
assign _77_ = _78_ | _80_ /*3164*/;
assign _86_ = ~D[13] /*3163*/;
assign _83_ = R_0[28] & _86_ /*3159*/;
assign _84_ = R_0[28] ^ _86_ /*3162*/;
assign _85_ = _77_ & _84_ /*3160*/;
assign _13_ = _77_ ^ _84_ /*3161*/;
assign _82_ = _83_ | _85_ /*3158*/;
assign _91_ = ~D[14] /*3157*/;
assign _88_ = R_0[29] & _91_ /*3153*/;
assign _89_ = R_0[29] ^ _91_ /*3156*/;
assign _90_ = _82_ & _89_ /*3154*/;
assign _14_ = _82_ ^ _89_ /*3155*/;
assign _87_ = _88_ | _90_ /*3152*/;
assign _92_ = zeroWire & oneWire /*3147*/;
assign _93_ = zeroWire ^ oneWire /*3150*/;
assign _94_ = _87_ & _93_ /*3148*/;
assign _15_ = _87_ ^ _93_ /*3149*/;
assign Q[15] = _92_ | _94_ /*3146*/;
assign _118_ = D[0] ^ Q[15] /*3050*/;
assign _115_ = R_0[14] & _118_ /*3046*/;
assign _116_ = R_0[14] ^ _118_ /*3049*/;
assign _117_ = Q[15] & _116_ /*3047*/;
assign _97_ = Q[15] ^ _116_ /*3048*/;
assign _114_ = _115_ | _117_ /*3045*/;
assign _123_ = D[1] ^ Q[15] /*3044*/;
assign _120_ = _0_ & _123_ /*3040*/;
assign _121_ = _0_ ^ _123_ /*3043*/;
assign _122_ = _114_ & _121_ /*3041*/;
assign _98_ = _114_ ^ _121_ /*3042*/;
assign _119_ = _120_ | _122_ /*3039*/;
assign _128_ = D[2] ^ Q[15] /*3038*/;
assign _125_ = _1_ & _128_ /*3034*/;
assign _126_ = _1_ ^ _128_ /*3037*/;
assign _127_ = _119_ & _126_ /*3035*/;
assign _99_ = _119_ ^ _126_ /*3036*/;
assign _124_ = _125_ | _127_ /*3033*/;
assign _133_ = D[3] ^ Q[15] /*3032*/;
assign _130_ = _2_ & _133_ /*3028*/;
assign _131_ = _2_ ^ _133_ /*3031*/;
assign _132_ = _124_ & _131_ /*3029*/;
assign _100_ = _124_ ^ _131_ /*3030*/;
assign _129_ = _130_ | _132_ /*3027*/;
assign _138_ = D[4] ^ Q[15] /*3026*/;
assign _135_ = _3_ & _138_ /*3022*/;
assign _136_ = _3_ ^ _138_ /*3025*/;
assign _137_ = _129_ & _136_ /*3023*/;
assign _101_ = _129_ ^ _136_ /*3024*/;
assign _134_ = _135_ | _137_ /*3021*/;
assign _143_ = D[5] ^ Q[15] /*3020*/;
assign _140_ = _4_ & _143_ /*3016*/;
assign _141_ = _4_ ^ _143_ /*3019*/;
assign _142_ = _134_ & _141_ /*3017*/;
assign _102_ = _134_ ^ _141_ /*3018*/;
assign _139_ = _140_ | _142_ /*3015*/;
assign _148_ = D[6] ^ Q[15] /*3014*/;
assign _145_ = _5_ & _148_ /*3010*/;
assign _146_ = _5_ ^ _148_ /*3013*/;
assign _147_ = _139_ & _146_ /*3011*/;
assign _103_ = _139_ ^ _146_ /*3012*/;
assign _144_ = _145_ | _147_ /*3009*/;
assign _153_ = D[7] ^ Q[15] /*3008*/;
assign _150_ = _6_ & _153_ /*3004*/;
assign _151_ = _6_ ^ _153_ /*3007*/;
assign _152_ = _144_ & _151_ /*3005*/;
assign _104_ = _144_ ^ _151_ /*3006*/;
assign _149_ = _150_ | _152_ /*3003*/;
assign _158_ = D[8] ^ Q[15] /*3002*/;
assign _155_ = _7_ & _158_ /*2998*/;
assign _156_ = _7_ ^ _158_ /*3001*/;
assign _157_ = _149_ & _156_ /*2999*/;
assign _105_ = _149_ ^ _156_ /*3000*/;
assign _154_ = _155_ | _157_ /*2997*/;
assign _163_ = D[9] ^ Q[15] /*2996*/;
assign _160_ = _8_ & _163_ /*2992*/;
assign _161_ = _8_ ^ _163_ /*2995*/;
assign _162_ = _154_ & _161_ /*2993*/;
assign _106_ = _154_ ^ _161_ /*2994*/;
assign _159_ = _160_ | _162_ /*2991*/;
assign _168_ = D[10] ^ Q[15] /*2990*/;
assign _165_ = _9_ & _168_ /*2986*/;
assign _166_ = _9_ ^ _168_ /*2989*/;
assign _167_ = _159_ & _166_ /*2987*/;
assign _107_ = _159_ ^ _166_ /*2988*/;
assign _164_ = _165_ | _167_ /*2985*/;
assign _173_ = D[11] ^ Q[15] /*2984*/;
assign _170_ = _10_ & _173_ /*2980*/;
assign _171_ = _10_ ^ _173_ /*2983*/;
assign _172_ = _164_ & _171_ /*2981*/;
assign _108_ = _164_ ^ _171_ /*2982*/;
assign _169_ = _170_ | _172_ /*2979*/;
assign _178_ = D[12] ^ Q[15] /*2978*/;
assign _175_ = _11_ & _178_ /*2974*/;
assign _176_ = _11_ ^ _178_ /*2977*/;
assign _177_ = _169_ & _176_ /*2975*/;
assign _109_ = _169_ ^ _176_ /*2976*/;
assign _174_ = _175_ | _177_ /*2973*/;
assign _183_ = D[13] ^ Q[15] /*2972*/;
assign _180_ = _12_ & _183_ /*2968*/;
assign _181_ = _12_ ^ _183_ /*2971*/;
assign _182_ = _174_ & _181_ /*2969*/;
assign _110_ = _174_ ^ _181_ /*2970*/;
assign _179_ = _180_ | _182_ /*2967*/;
assign _188_ = D[14] ^ Q[15] /*2966*/;
assign _185_ = _13_ & _188_ /*2962*/;
assign _186_ = _13_ ^ _188_ /*2965*/;
assign _187_ = _179_ & _186_ /*2963*/;
assign _111_ = _179_ ^ _186_ /*2964*/;
assign _184_ = _185_ | _187_ /*2961*/;
assign _192_ = zeroWire ^ Q[15] /*2960*/;
assign _189_ = _14_ & _192_ /*2956*/;
assign _190_ = _14_ ^ _192_ /*2959*/;
assign _191_ = _184_ & _190_ /*2957*/;
assign _112_ = _184_ ^ _190_ /*2958*/;
assign Q[14] = _189_ | _191_ /*2955*/;
assign _215_ = D[0] ^ Q[14] /*2857*/;
assign _212_ = R_0[13] & _215_ /*2853*/;
assign _213_ = R_0[13] ^ _215_ /*2856*/;
assign _214_ = Q[14] & _213_ /*2854*/;
assign _194_ = Q[14] ^ _213_ /*2855*/;
assign _211_ = _212_ | _214_ /*2852*/;
assign _220_ = D[1] ^ Q[14] /*2851*/;
assign _217_ = _97_ & _220_ /*2847*/;
assign _218_ = _97_ ^ _220_ /*2850*/;
assign _219_ = _211_ & _218_ /*2848*/;
assign _195_ = _211_ ^ _218_ /*2849*/;
assign _216_ = _217_ | _219_ /*2846*/;
assign _225_ = D[2] ^ Q[14] /*2845*/;
assign _222_ = _98_ & _225_ /*2841*/;
assign _223_ = _98_ ^ _225_ /*2844*/;
assign _224_ = _216_ & _223_ /*2842*/;
assign _196_ = _216_ ^ _223_ /*2843*/;
assign _221_ = _222_ | _224_ /*2840*/;
assign _230_ = D[3] ^ Q[14] /*2839*/;
assign _227_ = _99_ & _230_ /*2835*/;
assign _228_ = _99_ ^ _230_ /*2838*/;
assign _229_ = _221_ & _228_ /*2836*/;
assign _197_ = _221_ ^ _228_ /*2837*/;
assign _226_ = _227_ | _229_ /*2834*/;
assign _235_ = D[4] ^ Q[14] /*2833*/;
assign _232_ = _100_ & _235_ /*2829*/;
assign _233_ = _100_ ^ _235_ /*2832*/;
assign _234_ = _226_ & _233_ /*2830*/;
assign _198_ = _226_ ^ _233_ /*2831*/;
assign _231_ = _232_ | _234_ /*2828*/;
assign _240_ = D[5] ^ Q[14] /*2827*/;
assign _237_ = _101_ & _240_ /*2823*/;
assign _238_ = _101_ ^ _240_ /*2826*/;
assign _239_ = _231_ & _238_ /*2824*/;
assign _199_ = _231_ ^ _238_ /*2825*/;
assign _236_ = _237_ | _239_ /*2822*/;
assign _245_ = D[6] ^ Q[14] /*2821*/;
assign _242_ = _102_ & _245_ /*2817*/;
assign _243_ = _102_ ^ _245_ /*2820*/;
assign _244_ = _236_ & _243_ /*2818*/;
assign _200_ = _236_ ^ _243_ /*2819*/;
assign _241_ = _242_ | _244_ /*2816*/;
assign _250_ = D[7] ^ Q[14] /*2815*/;
assign _247_ = _103_ & _250_ /*2811*/;
assign _248_ = _103_ ^ _250_ /*2814*/;
assign _249_ = _241_ & _248_ /*2812*/;
assign _201_ = _241_ ^ _248_ /*2813*/;
assign _246_ = _247_ | _249_ /*2810*/;
assign _255_ = D[8] ^ Q[14] /*2809*/;
assign _252_ = _104_ & _255_ /*2805*/;
assign _253_ = _104_ ^ _255_ /*2808*/;
assign _254_ = _246_ & _253_ /*2806*/;
assign _202_ = _246_ ^ _253_ /*2807*/;
assign _251_ = _252_ | _254_ /*2804*/;
assign _260_ = D[9] ^ Q[14] /*2803*/;
assign _257_ = _105_ & _260_ /*2799*/;
assign _258_ = _105_ ^ _260_ /*2802*/;
assign _259_ = _251_ & _258_ /*2800*/;
assign _203_ = _251_ ^ _258_ /*2801*/;
assign _256_ = _257_ | _259_ /*2798*/;
assign _265_ = D[10] ^ Q[14] /*2797*/;
assign _262_ = _106_ & _265_ /*2793*/;
assign _263_ = _106_ ^ _265_ /*2796*/;
assign _264_ = _256_ & _263_ /*2794*/;
assign _204_ = _256_ ^ _263_ /*2795*/;
assign _261_ = _262_ | _264_ /*2792*/;
assign _270_ = D[11] ^ Q[14] /*2791*/;
assign _267_ = _107_ & _270_ /*2787*/;
assign _268_ = _107_ ^ _270_ /*2790*/;
assign _269_ = _261_ & _268_ /*2788*/;
assign _205_ = _261_ ^ _268_ /*2789*/;
assign _266_ = _267_ | _269_ /*2786*/;
assign _275_ = D[12] ^ Q[14] /*2785*/;
assign _272_ = _108_ & _275_ /*2781*/;
assign _273_ = _108_ ^ _275_ /*2784*/;
assign _274_ = _266_ & _273_ /*2782*/;
assign _206_ = _266_ ^ _273_ /*2783*/;
assign _271_ = _272_ | _274_ /*2780*/;
assign _280_ = D[13] ^ Q[14] /*2779*/;
assign _277_ = _109_ & _280_ /*2775*/;
assign _278_ = _109_ ^ _280_ /*2778*/;
assign _279_ = _271_ & _278_ /*2776*/;
assign _207_ = _271_ ^ _278_ /*2777*/;
assign _276_ = _277_ | _279_ /*2774*/;
assign _285_ = D[14] ^ Q[14] /*2773*/;
assign _282_ = _110_ & _285_ /*2769*/;
assign _283_ = _110_ ^ _285_ /*2772*/;
assign _284_ = _276_ & _283_ /*2770*/;
assign _208_ = _276_ ^ _283_ /*2771*/;
assign _281_ = _282_ | _284_ /*2768*/;
assign _289_ = zeroWire ^ Q[14] /*2767*/;
assign _286_ = _111_ & _289_ /*2763*/;
assign _287_ = _111_ ^ _289_ /*2766*/;
assign _288_ = _281_ & _287_ /*2764*/;
assign _209_ = _281_ ^ _287_ /*2765*/;
assign Q[13] = _286_ | _288_ /*2762*/;
assign _312_ = D[0] ^ Q[13] /*2664*/;
assign _309_ = R_0[12] & _312_ /*2660*/;
assign _310_ = R_0[12] ^ _312_ /*2663*/;
assign _311_ = Q[13] & _310_ /*2661*/;
assign _291_ = Q[13] ^ _310_ /*2662*/;
assign _308_ = _309_ | _311_ /*2659*/;
assign _317_ = D[1] ^ Q[13] /*2658*/;
assign _314_ = _194_ & _317_ /*2654*/;
assign _315_ = _194_ ^ _317_ /*2657*/;
assign _316_ = _308_ & _315_ /*2655*/;
assign _292_ = _308_ ^ _315_ /*2656*/;
assign _313_ = _314_ | _316_ /*2653*/;
assign _322_ = D[2] ^ Q[13] /*2652*/;
assign _319_ = _195_ & _322_ /*2648*/;
assign _320_ = _195_ ^ _322_ /*2651*/;
assign _321_ = _313_ & _320_ /*2649*/;
assign _293_ = _313_ ^ _320_ /*2650*/;
assign _318_ = _319_ | _321_ /*2647*/;
assign _327_ = D[3] ^ Q[13] /*2646*/;
assign _324_ = _196_ & _327_ /*2642*/;
assign _325_ = _196_ ^ _327_ /*2645*/;
assign _326_ = _318_ & _325_ /*2643*/;
assign _294_ = _318_ ^ _325_ /*2644*/;
assign _323_ = _324_ | _326_ /*2641*/;
assign _332_ = D[4] ^ Q[13] /*2640*/;
assign _329_ = _197_ & _332_ /*2636*/;
assign _330_ = _197_ ^ _332_ /*2639*/;
assign _331_ = _323_ & _330_ /*2637*/;
assign _295_ = _323_ ^ _330_ /*2638*/;
assign _328_ = _329_ | _331_ /*2635*/;
assign _337_ = D[5] ^ Q[13] /*2634*/;
assign _334_ = _198_ & _337_ /*2630*/;
assign _335_ = _198_ ^ _337_ /*2633*/;
assign _336_ = _328_ & _335_ /*2631*/;
assign _296_ = _328_ ^ _335_ /*2632*/;
assign _333_ = _334_ | _336_ /*2629*/;
assign _342_ = D[6] ^ Q[13] /*2628*/;
assign _339_ = _199_ & _342_ /*2624*/;
assign _340_ = _199_ ^ _342_ /*2627*/;
assign _341_ = _333_ & _340_ /*2625*/;
assign _297_ = _333_ ^ _340_ /*2626*/;
assign _338_ = _339_ | _341_ /*2623*/;
assign _347_ = D[7] ^ Q[13] /*2622*/;
assign _344_ = _200_ & _347_ /*2618*/;
assign _345_ = _200_ ^ _347_ /*2621*/;
assign _346_ = _338_ & _345_ /*2619*/;
assign _298_ = _338_ ^ _345_ /*2620*/;
assign _343_ = _344_ | _346_ /*2617*/;
assign _352_ = D[8] ^ Q[13] /*2616*/;
assign _349_ = _201_ & _352_ /*2612*/;
assign _350_ = _201_ ^ _352_ /*2615*/;
assign _351_ = _343_ & _350_ /*2613*/;
assign _299_ = _343_ ^ _350_ /*2614*/;
assign _348_ = _349_ | _351_ /*2611*/;
assign _357_ = D[9] ^ Q[13] /*2610*/;
assign _354_ = _202_ & _357_ /*2606*/;
assign _355_ = _202_ ^ _357_ /*2609*/;
assign _356_ = _348_ & _355_ /*2607*/;
assign _300_ = _348_ ^ _355_ /*2608*/;
assign _353_ = _354_ | _356_ /*2605*/;
assign _362_ = D[10] ^ Q[13] /*2604*/;
assign _359_ = _203_ & _362_ /*2600*/;
assign _360_ = _203_ ^ _362_ /*2603*/;
assign _361_ = _353_ & _360_ /*2601*/;
assign _301_ = _353_ ^ _360_ /*2602*/;
assign _358_ = _359_ | _361_ /*2599*/;
assign _367_ = D[11] ^ Q[13] /*2598*/;
assign _364_ = _204_ & _367_ /*2594*/;
assign _365_ = _204_ ^ _367_ /*2597*/;
assign _366_ = _358_ & _365_ /*2595*/;
assign _302_ = _358_ ^ _365_ /*2596*/;
assign _363_ = _364_ | _366_ /*2593*/;
assign _372_ = D[12] ^ Q[13] /*2592*/;
assign _369_ = _205_ & _372_ /*2588*/;
assign _370_ = _205_ ^ _372_ /*2591*/;
assign _371_ = _363_ & _370_ /*2589*/;
assign _303_ = _363_ ^ _370_ /*2590*/;
assign _368_ = _369_ | _371_ /*2587*/;
assign _377_ = D[13] ^ Q[13] /*2586*/;
assign _374_ = _206_ & _377_ /*2582*/;
assign _375_ = _206_ ^ _377_ /*2585*/;
assign _376_ = _368_ & _375_ /*2583*/;
assign _304_ = _368_ ^ _375_ /*2584*/;
assign _373_ = _374_ | _376_ /*2581*/;
assign _382_ = D[14] ^ Q[13] /*2580*/;
assign _379_ = _207_ & _382_ /*2576*/;
assign _380_ = _207_ ^ _382_ /*2579*/;
assign _381_ = _373_ & _380_ /*2577*/;
assign _305_ = _373_ ^ _380_ /*2578*/;
assign _378_ = _379_ | _381_ /*2575*/;
assign _386_ = zeroWire ^ Q[13] /*2574*/;
assign _383_ = _208_ & _386_ /*2570*/;
assign _384_ = _208_ ^ _386_ /*2573*/;
assign _385_ = _378_ & _384_ /*2571*/;
assign _306_ = _378_ ^ _384_ /*2572*/;
assign Q[12] = _383_ | _385_ /*2569*/;
assign _409_ = D[0] ^ Q[12] /*2471*/;
assign _406_ = R_0[11] & _409_ /*2467*/;
assign _407_ = R_0[11] ^ _409_ /*2470*/;
assign _408_ = Q[12] & _407_ /*2468*/;
assign _388_ = Q[12] ^ _407_ /*2469*/;
assign _405_ = _406_ | _408_ /*2466*/;
assign _414_ = D[1] ^ Q[12] /*2465*/;
assign _411_ = _291_ & _414_ /*2461*/;
assign _412_ = _291_ ^ _414_ /*2464*/;
assign _413_ = _405_ & _412_ /*2462*/;
assign _389_ = _405_ ^ _412_ /*2463*/;
assign _410_ = _411_ | _413_ /*2460*/;
assign _419_ = D[2] ^ Q[12] /*2459*/;
assign _416_ = _292_ & _419_ /*2455*/;
assign _417_ = _292_ ^ _419_ /*2458*/;
assign _418_ = _410_ & _417_ /*2456*/;
assign _390_ = _410_ ^ _417_ /*2457*/;
assign _415_ = _416_ | _418_ /*2454*/;
assign _424_ = D[3] ^ Q[12] /*2453*/;
assign _421_ = _293_ & _424_ /*2449*/;
assign _422_ = _293_ ^ _424_ /*2452*/;
assign _423_ = _415_ & _422_ /*2450*/;
assign _391_ = _415_ ^ _422_ /*2451*/;
assign _420_ = _421_ | _423_ /*2448*/;
assign _429_ = D[4] ^ Q[12] /*2447*/;
assign _426_ = _294_ & _429_ /*2443*/;
assign _427_ = _294_ ^ _429_ /*2446*/;
assign _428_ = _420_ & _427_ /*2444*/;
assign _392_ = _420_ ^ _427_ /*2445*/;
assign _425_ = _426_ | _428_ /*2442*/;
assign _434_ = D[5] ^ Q[12] /*2441*/;
assign _431_ = _295_ & _434_ /*2437*/;
assign _432_ = _295_ ^ _434_ /*2440*/;
assign _433_ = _425_ & _432_ /*2438*/;
assign _393_ = _425_ ^ _432_ /*2439*/;
assign _430_ = _431_ | _433_ /*2436*/;
assign _439_ = D[6] ^ Q[12] /*2435*/;
assign _436_ = _296_ & _439_ /*2431*/;
assign _437_ = _296_ ^ _439_ /*2434*/;
assign _438_ = _430_ & _437_ /*2432*/;
assign _394_ = _430_ ^ _437_ /*2433*/;
assign _435_ = _436_ | _438_ /*2430*/;
assign _444_ = D[7] ^ Q[12] /*2429*/;
assign _441_ = _297_ & _444_ /*2425*/;
assign _442_ = _297_ ^ _444_ /*2428*/;
assign _443_ = _435_ & _442_ /*2426*/;
assign _395_ = _435_ ^ _442_ /*2427*/;
assign _440_ = _441_ | _443_ /*2424*/;
assign _449_ = D[8] ^ Q[12] /*2423*/;
assign _446_ = _298_ & _449_ /*2419*/;
assign _447_ = _298_ ^ _449_ /*2422*/;
assign _448_ = _440_ & _447_ /*2420*/;
assign _396_ = _440_ ^ _447_ /*2421*/;
assign _445_ = _446_ | _448_ /*2418*/;
assign _454_ = D[9] ^ Q[12] /*2417*/;
assign _451_ = _299_ & _454_ /*2413*/;
assign _452_ = _299_ ^ _454_ /*2416*/;
assign _453_ = _445_ & _452_ /*2414*/;
assign _397_ = _445_ ^ _452_ /*2415*/;
assign _450_ = _451_ | _453_ /*2412*/;
assign _459_ = D[10] ^ Q[12] /*2411*/;
assign _456_ = _300_ & _459_ /*2407*/;
assign _457_ = _300_ ^ _459_ /*2410*/;
assign _458_ = _450_ & _457_ /*2408*/;
assign _398_ = _450_ ^ _457_ /*2409*/;
assign _455_ = _456_ | _458_ /*2406*/;
assign _464_ = D[11] ^ Q[12] /*2405*/;
assign _461_ = _301_ & _464_ /*2401*/;
assign _462_ = _301_ ^ _464_ /*2404*/;
assign _463_ = _455_ & _462_ /*2402*/;
assign _399_ = _455_ ^ _462_ /*2403*/;
assign _460_ = _461_ | _463_ /*2400*/;
assign _469_ = D[12] ^ Q[12] /*2399*/;
assign _466_ = _302_ & _469_ /*2395*/;
assign _467_ = _302_ ^ _469_ /*2398*/;
assign _468_ = _460_ & _467_ /*2396*/;
assign _400_ = _460_ ^ _467_ /*2397*/;
assign _465_ = _466_ | _468_ /*2394*/;
assign _474_ = D[13] ^ Q[12] /*2393*/;
assign _471_ = _303_ & _474_ /*2389*/;
assign _472_ = _303_ ^ _474_ /*2392*/;
assign _473_ = _465_ & _472_ /*2390*/;
assign _401_ = _465_ ^ _472_ /*2391*/;
assign _470_ = _471_ | _473_ /*2388*/;
assign _479_ = D[14] ^ Q[12] /*2387*/;
assign _476_ = _304_ & _479_ /*2383*/;
assign _477_ = _304_ ^ _479_ /*2386*/;
assign _478_ = _470_ & _477_ /*2384*/;
assign _402_ = _470_ ^ _477_ /*2385*/;
assign _475_ = _476_ | _478_ /*2382*/;
assign _483_ = zeroWire ^ Q[12] /*2381*/;
assign _480_ = _305_ & _483_ /*2377*/;
assign _481_ = _305_ ^ _483_ /*2380*/;
assign _482_ = _475_ & _481_ /*2378*/;
assign _403_ = _475_ ^ _481_ /*2379*/;
assign Q[11] = _480_ | _482_ /*2376*/;
assign _506_ = D[0] ^ Q[11] /*2278*/;
assign _503_ = R_0[10] & _506_ /*2274*/;
assign _504_ = R_0[10] ^ _506_ /*2277*/;
assign _505_ = Q[11] & _504_ /*2275*/;
assign _485_ = Q[11] ^ _504_ /*2276*/;
assign _502_ = _503_ | _505_ /*2273*/;
assign _511_ = D[1] ^ Q[11] /*2272*/;
assign _508_ = _388_ & _511_ /*2268*/;
assign _509_ = _388_ ^ _511_ /*2271*/;
assign _510_ = _502_ & _509_ /*2269*/;
assign _486_ = _502_ ^ _509_ /*2270*/;
assign _507_ = _508_ | _510_ /*2267*/;
assign _516_ = D[2] ^ Q[11] /*2266*/;
assign _513_ = _389_ & _516_ /*2262*/;
assign _514_ = _389_ ^ _516_ /*2265*/;
assign _515_ = _507_ & _514_ /*2263*/;
assign _487_ = _507_ ^ _514_ /*2264*/;
assign _512_ = _513_ | _515_ /*2261*/;
assign _521_ = D[3] ^ Q[11] /*2260*/;
assign _518_ = _390_ & _521_ /*2256*/;
assign _519_ = _390_ ^ _521_ /*2259*/;
assign _520_ = _512_ & _519_ /*2257*/;
assign _488_ = _512_ ^ _519_ /*2258*/;
assign _517_ = _518_ | _520_ /*2255*/;
assign _526_ = D[4] ^ Q[11] /*2254*/;
assign _523_ = _391_ & _526_ /*2250*/;
assign _524_ = _391_ ^ _526_ /*2253*/;
assign _525_ = _517_ & _524_ /*2251*/;
assign _489_ = _517_ ^ _524_ /*2252*/;
assign _522_ = _523_ | _525_ /*2249*/;
assign _531_ = D[5] ^ Q[11] /*2248*/;
assign _528_ = _392_ & _531_ /*2244*/;
assign _529_ = _392_ ^ _531_ /*2247*/;
assign _530_ = _522_ & _529_ /*2245*/;
assign _490_ = _522_ ^ _529_ /*2246*/;
assign _527_ = _528_ | _530_ /*2243*/;
assign _536_ = D[6] ^ Q[11] /*2242*/;
assign _533_ = _393_ & _536_ /*2238*/;
assign _534_ = _393_ ^ _536_ /*2241*/;
assign _535_ = _527_ & _534_ /*2239*/;
assign _491_ = _527_ ^ _534_ /*2240*/;
assign _532_ = _533_ | _535_ /*2237*/;
assign _541_ = D[7] ^ Q[11] /*2236*/;
assign _538_ = _394_ & _541_ /*2232*/;
assign _539_ = _394_ ^ _541_ /*2235*/;
assign _540_ = _532_ & _539_ /*2233*/;
assign _492_ = _532_ ^ _539_ /*2234*/;
assign _537_ = _538_ | _540_ /*2231*/;
assign _546_ = D[8] ^ Q[11] /*2230*/;
assign _543_ = _395_ & _546_ /*2226*/;
assign _544_ = _395_ ^ _546_ /*2229*/;
assign _545_ = _537_ & _544_ /*2227*/;
assign _493_ = _537_ ^ _544_ /*2228*/;
assign _542_ = _543_ | _545_ /*2225*/;
assign _551_ = D[9] ^ Q[11] /*2224*/;
assign _548_ = _396_ & _551_ /*2220*/;
assign _549_ = _396_ ^ _551_ /*2223*/;
assign _550_ = _542_ & _549_ /*2221*/;
assign _494_ = _542_ ^ _549_ /*2222*/;
assign _547_ = _548_ | _550_ /*2219*/;
assign _556_ = D[10] ^ Q[11] /*2218*/;
assign _553_ = _397_ & _556_ /*2214*/;
assign _554_ = _397_ ^ _556_ /*2217*/;
assign _555_ = _547_ & _554_ /*2215*/;
assign _495_ = _547_ ^ _554_ /*2216*/;
assign _552_ = _553_ | _555_ /*2213*/;
assign _561_ = D[11] ^ Q[11] /*2212*/;
assign _558_ = _398_ & _561_ /*2208*/;
assign _559_ = _398_ ^ _561_ /*2211*/;
assign _560_ = _552_ & _559_ /*2209*/;
assign _496_ = _552_ ^ _559_ /*2210*/;
assign _557_ = _558_ | _560_ /*2207*/;
assign _566_ = D[12] ^ Q[11] /*2206*/;
assign _563_ = _399_ & _566_ /*2202*/;
assign _564_ = _399_ ^ _566_ /*2205*/;
assign _565_ = _557_ & _564_ /*2203*/;
assign _497_ = _557_ ^ _564_ /*2204*/;
assign _562_ = _563_ | _565_ /*2201*/;
assign _571_ = D[13] ^ Q[11] /*2200*/;
assign _568_ = _400_ & _571_ /*2196*/;
assign _569_ = _400_ ^ _571_ /*2199*/;
assign _570_ = _562_ & _569_ /*2197*/;
assign _498_ = _562_ ^ _569_ /*2198*/;
assign _567_ = _568_ | _570_ /*2195*/;
assign _576_ = D[14] ^ Q[11] /*2194*/;
assign _573_ = _401_ & _576_ /*2190*/;
assign _574_ = _401_ ^ _576_ /*2193*/;
assign _575_ = _567_ & _574_ /*2191*/;
assign _499_ = _567_ ^ _574_ /*2192*/;
assign _572_ = _573_ | _575_ /*2189*/;
assign _580_ = zeroWire ^ Q[11] /*2188*/;
assign _577_ = _402_ & _580_ /*2184*/;
assign _578_ = _402_ ^ _580_ /*2187*/;
assign _579_ = _572_ & _578_ /*2185*/;
assign _500_ = _572_ ^ _578_ /*2186*/;
assign Q[10] = _577_ | _579_ /*2183*/;
assign _603_ = D[0] ^ Q[10] /*2085*/;
assign _600_ = R_0[9] & _603_ /*2081*/;
assign _601_ = R_0[9] ^ _603_ /*2084*/;
assign _602_ = Q[10] & _601_ /*2082*/;
assign _582_ = Q[10] ^ _601_ /*2083*/;
assign _599_ = _600_ | _602_ /*2080*/;
assign _608_ = D[1] ^ Q[10] /*2079*/;
assign _605_ = _485_ & _608_ /*2075*/;
assign _606_ = _485_ ^ _608_ /*2078*/;
assign _607_ = _599_ & _606_ /*2076*/;
assign _583_ = _599_ ^ _606_ /*2077*/;
assign _604_ = _605_ | _607_ /*2074*/;
assign _613_ = D[2] ^ Q[10] /*2073*/;
assign _610_ = _486_ & _613_ /*2069*/;
assign _611_ = _486_ ^ _613_ /*2072*/;
assign _612_ = _604_ & _611_ /*2070*/;
assign _584_ = _604_ ^ _611_ /*2071*/;
assign _609_ = _610_ | _612_ /*2068*/;
assign _618_ = D[3] ^ Q[10] /*2067*/;
assign _615_ = _487_ & _618_ /*2063*/;
assign _616_ = _487_ ^ _618_ /*2066*/;
assign _617_ = _609_ & _616_ /*2064*/;
assign _585_ = _609_ ^ _616_ /*2065*/;
assign _614_ = _615_ | _617_ /*2062*/;
assign _623_ = D[4] ^ Q[10] /*2061*/;
assign _620_ = _488_ & _623_ /*2057*/;
assign _621_ = _488_ ^ _623_ /*2060*/;
assign _622_ = _614_ & _621_ /*2058*/;
assign _586_ = _614_ ^ _621_ /*2059*/;
assign _619_ = _620_ | _622_ /*2056*/;
assign _628_ = D[5] ^ Q[10] /*2055*/;
assign _625_ = _489_ & _628_ /*2051*/;
assign _626_ = _489_ ^ _628_ /*2054*/;
assign _627_ = _619_ & _626_ /*2052*/;
assign _587_ = _619_ ^ _626_ /*2053*/;
assign _624_ = _625_ | _627_ /*2050*/;
assign _633_ = D[6] ^ Q[10] /*2049*/;
assign _630_ = _490_ & _633_ /*2045*/;
assign _631_ = _490_ ^ _633_ /*2048*/;
assign _632_ = _624_ & _631_ /*2046*/;
assign _588_ = _624_ ^ _631_ /*2047*/;
assign _629_ = _630_ | _632_ /*2044*/;
assign _638_ = D[7] ^ Q[10] /*2043*/;
assign _635_ = _491_ & _638_ /*2039*/;
assign _636_ = _491_ ^ _638_ /*2042*/;
assign _637_ = _629_ & _636_ /*2040*/;
assign _589_ = _629_ ^ _636_ /*2041*/;
assign _634_ = _635_ | _637_ /*2038*/;
assign _643_ = D[8] ^ Q[10] /*2037*/;
assign _640_ = _492_ & _643_ /*2033*/;
assign _641_ = _492_ ^ _643_ /*2036*/;
assign _642_ = _634_ & _641_ /*2034*/;
assign _590_ = _634_ ^ _641_ /*2035*/;
assign _639_ = _640_ | _642_ /*2032*/;
assign _648_ = D[9] ^ Q[10] /*2031*/;
assign _645_ = _493_ & _648_ /*2027*/;
assign _646_ = _493_ ^ _648_ /*2030*/;
assign _647_ = _639_ & _646_ /*2028*/;
assign _591_ = _639_ ^ _646_ /*2029*/;
assign _644_ = _645_ | _647_ /*2026*/;
assign _653_ = D[10] ^ Q[10] /*2025*/;
assign _650_ = _494_ & _653_ /*2021*/;
assign _651_ = _494_ ^ _653_ /*2024*/;
assign _652_ = _644_ & _651_ /*2022*/;
assign _592_ = _644_ ^ _651_ /*2023*/;
assign _649_ = _650_ | _652_ /*2020*/;
assign _658_ = D[11] ^ Q[10] /*2019*/;
assign _655_ = _495_ & _658_ /*2015*/;
assign _656_ = _495_ ^ _658_ /*2018*/;
assign _657_ = _649_ & _656_ /*2016*/;
assign _593_ = _649_ ^ _656_ /*2017*/;
assign _654_ = _655_ | _657_ /*2014*/;
assign _663_ = D[12] ^ Q[10] /*2013*/;
assign _660_ = _496_ & _663_ /*2009*/;
assign _661_ = _496_ ^ _663_ /*2012*/;
assign _662_ = _654_ & _661_ /*2010*/;
assign _594_ = _654_ ^ _661_ /*2011*/;
assign _659_ = _660_ | _662_ /*2008*/;
assign _668_ = D[13] ^ Q[10] /*2007*/;
assign _665_ = _497_ & _668_ /*2003*/;
assign _666_ = _497_ ^ _668_ /*2006*/;
assign _667_ = _659_ & _666_ /*2004*/;
assign _595_ = _659_ ^ _666_ /*2005*/;
assign _664_ = _665_ | _667_ /*2002*/;
assign _673_ = D[14] ^ Q[10] /*2001*/;
assign _670_ = _498_ & _673_ /*1997*/;
assign _671_ = _498_ ^ _673_ /*2000*/;
assign _672_ = _664_ & _671_ /*1998*/;
assign _596_ = _664_ ^ _671_ /*1999*/;
assign _669_ = _670_ | _672_ /*1996*/;
assign _677_ = zeroWire ^ Q[10] /*1995*/;
assign _674_ = _499_ & _677_ /*1991*/;
assign _675_ = _499_ ^ _677_ /*1994*/;
assign _676_ = _669_ & _675_ /*1992*/;
assign _597_ = _669_ ^ _675_ /*1993*/;
assign Q[9] = _674_ | _676_ /*1990*/;
assign _700_ = D[0] ^ Q[9] /*1892*/;
assign _697_ = R_0[8] & _700_ /*1888*/;
assign _698_ = R_0[8] ^ _700_ /*1891*/;
assign _699_ = Q[9] & _698_ /*1889*/;
assign _679_ = Q[9] ^ _698_ /*1890*/;
assign _696_ = _697_ | _699_ /*1887*/;
assign _705_ = D[1] ^ Q[9] /*1886*/;
assign _702_ = _582_ & _705_ /*1882*/;
assign _703_ = _582_ ^ _705_ /*1885*/;
assign _704_ = _696_ & _703_ /*1883*/;
assign _680_ = _696_ ^ _703_ /*1884*/;
assign _701_ = _702_ | _704_ /*1881*/;
assign _710_ = D[2] ^ Q[9] /*1880*/;
assign _707_ = _583_ & _710_ /*1876*/;
assign _708_ = _583_ ^ _710_ /*1879*/;
assign _709_ = _701_ & _708_ /*1877*/;
assign _681_ = _701_ ^ _708_ /*1878*/;
assign _706_ = _707_ | _709_ /*1875*/;
assign _715_ = D[3] ^ Q[9] /*1874*/;
assign _712_ = _584_ & _715_ /*1870*/;
assign _713_ = _584_ ^ _715_ /*1873*/;
assign _714_ = _706_ & _713_ /*1871*/;
assign _682_ = _706_ ^ _713_ /*1872*/;
assign _711_ = _712_ | _714_ /*1869*/;
assign _720_ = D[4] ^ Q[9] /*1868*/;
assign _717_ = _585_ & _720_ /*1864*/;
assign _718_ = _585_ ^ _720_ /*1867*/;
assign _719_ = _711_ & _718_ /*1865*/;
assign _683_ = _711_ ^ _718_ /*1866*/;
assign _716_ = _717_ | _719_ /*1863*/;
assign _725_ = D[5] ^ Q[9] /*1862*/;
assign _722_ = _586_ & _725_ /*1858*/;
assign _723_ = _586_ ^ _725_ /*1861*/;
assign _724_ = _716_ & _723_ /*1859*/;
assign _684_ = _716_ ^ _723_ /*1860*/;
assign _721_ = _722_ | _724_ /*1857*/;
assign _730_ = D[6] ^ Q[9] /*1856*/;
assign _727_ = _587_ & _730_ /*1852*/;
assign _728_ = _587_ ^ _730_ /*1855*/;
assign _729_ = _721_ & _728_ /*1853*/;
assign _685_ = _721_ ^ _728_ /*1854*/;
assign _726_ = _727_ | _729_ /*1851*/;
assign _735_ = D[7] ^ Q[9] /*1850*/;
assign _732_ = _588_ & _735_ /*1846*/;
assign _733_ = _588_ ^ _735_ /*1849*/;
assign _734_ = _726_ & _733_ /*1847*/;
assign _686_ = _726_ ^ _733_ /*1848*/;
assign _731_ = _732_ | _734_ /*1845*/;
assign _740_ = D[8] ^ Q[9] /*1844*/;
assign _737_ = _589_ & _740_ /*1840*/;
assign _738_ = _589_ ^ _740_ /*1843*/;
assign _739_ = _731_ & _738_ /*1841*/;
assign _687_ = _731_ ^ _738_ /*1842*/;
assign _736_ = _737_ | _739_ /*1839*/;
assign _745_ = D[9] ^ Q[9] /*1838*/;
assign _742_ = _590_ & _745_ /*1834*/;
assign _743_ = _590_ ^ _745_ /*1837*/;
assign _744_ = _736_ & _743_ /*1835*/;
assign _688_ = _736_ ^ _743_ /*1836*/;
assign _741_ = _742_ | _744_ /*1833*/;
assign _750_ = D[10] ^ Q[9] /*1832*/;
assign _747_ = _591_ & _750_ /*1828*/;
assign _748_ = _591_ ^ _750_ /*1831*/;
assign _749_ = _741_ & _748_ /*1829*/;
assign _689_ = _741_ ^ _748_ /*1830*/;
assign _746_ = _747_ | _749_ /*1827*/;
assign _755_ = D[11] ^ Q[9] /*1826*/;
assign _752_ = _592_ & _755_ /*1822*/;
assign _753_ = _592_ ^ _755_ /*1825*/;
assign _754_ = _746_ & _753_ /*1823*/;
assign _690_ = _746_ ^ _753_ /*1824*/;
assign _751_ = _752_ | _754_ /*1821*/;
assign _760_ = D[12] ^ Q[9] /*1820*/;
assign _757_ = _593_ & _760_ /*1816*/;
assign _758_ = _593_ ^ _760_ /*1819*/;
assign _759_ = _751_ & _758_ /*1817*/;
assign _691_ = _751_ ^ _758_ /*1818*/;
assign _756_ = _757_ | _759_ /*1815*/;
assign _765_ = D[13] ^ Q[9] /*1814*/;
assign _762_ = _594_ & _765_ /*1810*/;
assign _763_ = _594_ ^ _765_ /*1813*/;
assign _764_ = _756_ & _763_ /*1811*/;
assign _692_ = _756_ ^ _763_ /*1812*/;
assign _761_ = _762_ | _764_ /*1809*/;
assign _770_ = D[14] ^ Q[9] /*1808*/;
assign _767_ = _595_ & _770_ /*1804*/;
assign _768_ = _595_ ^ _770_ /*1807*/;
assign _769_ = _761_ & _768_ /*1805*/;
assign _693_ = _761_ ^ _768_ /*1806*/;
assign _766_ = _767_ | _769_ /*1803*/;
assign _774_ = zeroWire ^ Q[9] /*1802*/;
assign _771_ = _596_ & _774_ /*1798*/;
assign _772_ = _596_ ^ _774_ /*1801*/;
assign _773_ = _766_ & _772_ /*1799*/;
assign _694_ = _766_ ^ _772_ /*1800*/;
assign Q[8] = _771_ | _773_ /*1797*/;
assign _797_ = D[0] ^ Q[8] /*1699*/;
assign _794_ = R_0[7] & _797_ /*1695*/;
assign _795_ = R_0[7] ^ _797_ /*1698*/;
assign _796_ = Q[8] & _795_ /*1696*/;
assign _776_ = Q[8] ^ _795_ /*1697*/;
assign _793_ = _794_ | _796_ /*1694*/;
assign _802_ = D[1] ^ Q[8] /*1693*/;
assign _799_ = _679_ & _802_ /*1689*/;
assign _800_ = _679_ ^ _802_ /*1692*/;
assign _801_ = _793_ & _800_ /*1690*/;
assign _777_ = _793_ ^ _800_ /*1691*/;
assign _798_ = _799_ | _801_ /*1688*/;
assign _807_ = D[2] ^ Q[8] /*1687*/;
assign _804_ = _680_ & _807_ /*1683*/;
assign _805_ = _680_ ^ _807_ /*1686*/;
assign _806_ = _798_ & _805_ /*1684*/;
assign _778_ = _798_ ^ _805_ /*1685*/;
assign _803_ = _804_ | _806_ /*1682*/;
assign _812_ = D[3] ^ Q[8] /*1681*/;
assign _809_ = _681_ & _812_ /*1677*/;
assign _810_ = _681_ ^ _812_ /*1680*/;
assign _811_ = _803_ & _810_ /*1678*/;
assign _779_ = _803_ ^ _810_ /*1679*/;
assign _808_ = _809_ | _811_ /*1676*/;
assign _817_ = D[4] ^ Q[8] /*1675*/;
assign _814_ = _682_ & _817_ /*1671*/;
assign _815_ = _682_ ^ _817_ /*1674*/;
assign _816_ = _808_ & _815_ /*1672*/;
assign _780_ = _808_ ^ _815_ /*1673*/;
assign _813_ = _814_ | _816_ /*1670*/;
assign _822_ = D[5] ^ Q[8] /*1669*/;
assign _819_ = _683_ & _822_ /*1665*/;
assign _820_ = _683_ ^ _822_ /*1668*/;
assign _821_ = _813_ & _820_ /*1666*/;
assign _781_ = _813_ ^ _820_ /*1667*/;
assign _818_ = _819_ | _821_ /*1664*/;
assign _827_ = D[6] ^ Q[8] /*1663*/;
assign _824_ = _684_ & _827_ /*1659*/;
assign _825_ = _684_ ^ _827_ /*1662*/;
assign _826_ = _818_ & _825_ /*1660*/;
assign _782_ = _818_ ^ _825_ /*1661*/;
assign _823_ = _824_ | _826_ /*1658*/;
assign _832_ = D[7] ^ Q[8] /*1657*/;
assign _829_ = _685_ & _832_ /*1653*/;
assign _830_ = _685_ ^ _832_ /*1656*/;
assign _831_ = _823_ & _830_ /*1654*/;
assign _783_ = _823_ ^ _830_ /*1655*/;
assign _828_ = _829_ | _831_ /*1652*/;
assign _837_ = D[8] ^ Q[8] /*1651*/;
assign _834_ = _686_ & _837_ /*1647*/;
assign _835_ = _686_ ^ _837_ /*1650*/;
assign _836_ = _828_ & _835_ /*1648*/;
assign _784_ = _828_ ^ _835_ /*1649*/;
assign _833_ = _834_ | _836_ /*1646*/;
assign _842_ = D[9] ^ Q[8] /*1645*/;
assign _839_ = _687_ & _842_ /*1641*/;
assign _840_ = _687_ ^ _842_ /*1644*/;
assign _841_ = _833_ & _840_ /*1642*/;
assign _785_ = _833_ ^ _840_ /*1643*/;
assign _838_ = _839_ | _841_ /*1640*/;
assign _847_ = D[10] ^ Q[8] /*1639*/;
assign _844_ = _688_ & _847_ /*1635*/;
assign _845_ = _688_ ^ _847_ /*1638*/;
assign _846_ = _838_ & _845_ /*1636*/;
assign _786_ = _838_ ^ _845_ /*1637*/;
assign _843_ = _844_ | _846_ /*1634*/;
assign _852_ = D[11] ^ Q[8] /*1633*/;
assign _849_ = _689_ & _852_ /*1629*/;
assign _850_ = _689_ ^ _852_ /*1632*/;
assign _851_ = _843_ & _850_ /*1630*/;
assign _787_ = _843_ ^ _850_ /*1631*/;
assign _848_ = _849_ | _851_ /*1628*/;
assign _857_ = D[12] ^ Q[8] /*1627*/;
assign _854_ = _690_ & _857_ /*1623*/;
assign _855_ = _690_ ^ _857_ /*1626*/;
assign _856_ = _848_ & _855_ /*1624*/;
assign _788_ = _848_ ^ _855_ /*1625*/;
assign _853_ = _854_ | _856_ /*1622*/;
assign _862_ = D[13] ^ Q[8] /*1621*/;
assign _859_ = _691_ & _862_ /*1617*/;
assign _860_ = _691_ ^ _862_ /*1620*/;
assign _861_ = _853_ & _860_ /*1618*/;
assign _789_ = _853_ ^ _860_ /*1619*/;
assign _858_ = _859_ | _861_ /*1616*/;
assign _867_ = D[14] ^ Q[8] /*1615*/;
assign _864_ = _692_ & _867_ /*1611*/;
assign _865_ = _692_ ^ _867_ /*1614*/;
assign _866_ = _858_ & _865_ /*1612*/;
assign _790_ = _858_ ^ _865_ /*1613*/;
assign _863_ = _864_ | _866_ /*1610*/;
assign _871_ = zeroWire ^ Q[8] /*1609*/;
assign _868_ = _693_ & _871_ /*1605*/;
assign _869_ = _693_ ^ _871_ /*1608*/;
assign _870_ = _863_ & _869_ /*1606*/;
assign _791_ = _863_ ^ _869_ /*1607*/;
assign Q[7] = _868_ | _870_ /*1604*/;
assign _894_ = D[0] ^ Q[7] /*1506*/;
assign _891_ = R_0[6] & _894_ /*1502*/;
assign _892_ = R_0[6] ^ _894_ /*1505*/;
assign _893_ = Q[7] & _892_ /*1503*/;
assign _873_ = Q[7] ^ _892_ /*1504*/;
assign _890_ = _891_ | _893_ /*1501*/;
assign _899_ = D[1] ^ Q[7] /*1500*/;
assign _896_ = _776_ & _899_ /*1496*/;
assign _897_ = _776_ ^ _899_ /*1499*/;
assign _898_ = _890_ & _897_ /*1497*/;
assign _874_ = _890_ ^ _897_ /*1498*/;
assign _895_ = _896_ | _898_ /*1495*/;
assign _904_ = D[2] ^ Q[7] /*1494*/;
assign _901_ = _777_ & _904_ /*1490*/;
assign _902_ = _777_ ^ _904_ /*1493*/;
assign _903_ = _895_ & _902_ /*1491*/;
assign _875_ = _895_ ^ _902_ /*1492*/;
assign _900_ = _901_ | _903_ /*1489*/;
assign _909_ = D[3] ^ Q[7] /*1488*/;
assign _906_ = _778_ & _909_ /*1484*/;
assign _907_ = _778_ ^ _909_ /*1487*/;
assign _908_ = _900_ & _907_ /*1485*/;
assign _876_ = _900_ ^ _907_ /*1486*/;
assign _905_ = _906_ | _908_ /*1483*/;
assign _914_ = D[4] ^ Q[7] /*1482*/;
assign _911_ = _779_ & _914_ /*1478*/;
assign _912_ = _779_ ^ _914_ /*1481*/;
assign _913_ = _905_ & _912_ /*1479*/;
assign _877_ = _905_ ^ _912_ /*1480*/;
assign _910_ = _911_ | _913_ /*1477*/;
assign _919_ = D[5] ^ Q[7] /*1476*/;
assign _916_ = _780_ & _919_ /*1472*/;
assign _917_ = _780_ ^ _919_ /*1475*/;
assign _918_ = _910_ & _917_ /*1473*/;
assign _878_ = _910_ ^ _917_ /*1474*/;
assign _915_ = _916_ | _918_ /*1471*/;
assign _924_ = D[6] ^ Q[7] /*1470*/;
assign _921_ = _781_ & _924_ /*1466*/;
assign _922_ = _781_ ^ _924_ /*1469*/;
assign _923_ = _915_ & _922_ /*1467*/;
assign _879_ = _915_ ^ _922_ /*1468*/;
assign _920_ = _921_ | _923_ /*1465*/;
assign _929_ = D[7] ^ Q[7] /*1464*/;
assign _926_ = _782_ & _929_ /*1460*/;
assign _927_ = _782_ ^ _929_ /*1463*/;
assign _928_ = _920_ & _927_ /*1461*/;
assign _880_ = _920_ ^ _927_ /*1462*/;
assign _925_ = _926_ | _928_ /*1459*/;
assign _934_ = D[8] ^ Q[7] /*1458*/;
assign _931_ = _783_ & _934_ /*1454*/;
assign _932_ = _783_ ^ _934_ /*1457*/;
assign _933_ = _925_ & _932_ /*1455*/;
assign _881_ = _925_ ^ _932_ /*1456*/;
assign _930_ = _931_ | _933_ /*1453*/;
assign _939_ = D[9] ^ Q[7] /*1452*/;
assign _936_ = _784_ & _939_ /*1448*/;
assign _937_ = _784_ ^ _939_ /*1451*/;
assign _938_ = _930_ & _937_ /*1449*/;
assign _882_ = _930_ ^ _937_ /*1450*/;
assign _935_ = _936_ | _938_ /*1447*/;
assign _944_ = D[10] ^ Q[7] /*1446*/;
assign _941_ = _785_ & _944_ /*1442*/;
assign _942_ = _785_ ^ _944_ /*1445*/;
assign _943_ = _935_ & _942_ /*1443*/;
assign _883_ = _935_ ^ _942_ /*1444*/;
assign _940_ = _941_ | _943_ /*1441*/;
assign _949_ = D[11] ^ Q[7] /*1440*/;
assign _946_ = _786_ & _949_ /*1436*/;
assign _947_ = _786_ ^ _949_ /*1439*/;
assign _948_ = _940_ & _947_ /*1437*/;
assign _884_ = _940_ ^ _947_ /*1438*/;
assign _945_ = _946_ | _948_ /*1435*/;
assign _954_ = D[12] ^ Q[7] /*1434*/;
assign _951_ = _787_ & _954_ /*1430*/;
assign _952_ = _787_ ^ _954_ /*1433*/;
assign _953_ = _945_ & _952_ /*1431*/;
assign _885_ = _945_ ^ _952_ /*1432*/;
assign _950_ = _951_ | _953_ /*1429*/;
assign _959_ = D[13] ^ Q[7] /*1428*/;
assign _956_ = _788_ & _959_ /*1424*/;
assign _957_ = _788_ ^ _959_ /*1427*/;
assign _958_ = _950_ & _957_ /*1425*/;
assign _886_ = _950_ ^ _957_ /*1426*/;
assign _955_ = _956_ | _958_ /*1423*/;
assign _964_ = D[14] ^ Q[7] /*1422*/;
assign _961_ = _789_ & _964_ /*1418*/;
assign _962_ = _789_ ^ _964_ /*1421*/;
assign _963_ = _955_ & _962_ /*1419*/;
assign _887_ = _955_ ^ _962_ /*1420*/;
assign _960_ = _961_ | _963_ /*1417*/;
assign _968_ = zeroWire ^ Q[7] /*1416*/;
assign _965_ = _790_ & _968_ /*1412*/;
assign _966_ = _790_ ^ _968_ /*1415*/;
assign _967_ = _960_ & _966_ /*1413*/;
assign _888_ = _960_ ^ _966_ /*1414*/;
assign Q[6] = _965_ | _967_ /*1411*/;
assign _991_ = D[0] ^ Q[6] /*1313*/;
assign _988_ = R_0[5] & _991_ /*1309*/;
assign _989_ = R_0[5] ^ _991_ /*1312*/;
assign _990_ = Q[6] & _989_ /*1310*/;
assign _970_ = Q[6] ^ _989_ /*1311*/;
assign _987_ = _988_ | _990_ /*1308*/;
assign _996_ = D[1] ^ Q[6] /*1307*/;
assign _993_ = _873_ & _996_ /*1303*/;
assign _994_ = _873_ ^ _996_ /*1306*/;
assign _995_ = _987_ & _994_ /*1304*/;
assign _971_ = _987_ ^ _994_ /*1305*/;
assign _992_ = _993_ | _995_ /*1302*/;
assign _1001_ = D[2] ^ Q[6] /*1301*/;
assign _998_ = _874_ & _1001_ /*1297*/;
assign _999_ = _874_ ^ _1001_ /*1300*/;
assign _1000_ = _992_ & _999_ /*1298*/;
assign _972_ = _992_ ^ _999_ /*1299*/;
assign _997_ = _998_ | _1000_ /*1296*/;
assign _1006_ = D[3] ^ Q[6] /*1295*/;
assign _1003_ = _875_ & _1006_ /*1291*/;
assign _1004_ = _875_ ^ _1006_ /*1294*/;
assign _1005_ = _997_ & _1004_ /*1292*/;
assign _973_ = _997_ ^ _1004_ /*1293*/;
assign _1002_ = _1003_ | _1005_ /*1290*/;
assign _1011_ = D[4] ^ Q[6] /*1289*/;
assign _1008_ = _876_ & _1011_ /*1285*/;
assign _1009_ = _876_ ^ _1011_ /*1288*/;
assign _1010_ = _1002_ & _1009_ /*1286*/;
assign _974_ = _1002_ ^ _1009_ /*1287*/;
assign _1007_ = _1008_ | _1010_ /*1284*/;
assign _1016_ = D[5] ^ Q[6] /*1283*/;
assign _1013_ = _877_ & _1016_ /*1279*/;
assign _1014_ = _877_ ^ _1016_ /*1282*/;
assign _1015_ = _1007_ & _1014_ /*1280*/;
assign _975_ = _1007_ ^ _1014_ /*1281*/;
assign _1012_ = _1013_ | _1015_ /*1278*/;
assign _1021_ = D[6] ^ Q[6] /*1277*/;
assign _1018_ = _878_ & _1021_ /*1273*/;
assign _1019_ = _878_ ^ _1021_ /*1276*/;
assign _1020_ = _1012_ & _1019_ /*1274*/;
assign _976_ = _1012_ ^ _1019_ /*1275*/;
assign _1017_ = _1018_ | _1020_ /*1272*/;
assign _1026_ = D[7] ^ Q[6] /*1271*/;
assign _1023_ = _879_ & _1026_ /*1267*/;
assign _1024_ = _879_ ^ _1026_ /*1270*/;
assign _1025_ = _1017_ & _1024_ /*1268*/;
assign _977_ = _1017_ ^ _1024_ /*1269*/;
assign _1022_ = _1023_ | _1025_ /*1266*/;
assign _1031_ = D[8] ^ Q[6] /*1265*/;
assign _1028_ = _880_ & _1031_ /*1261*/;
assign _1029_ = _880_ ^ _1031_ /*1264*/;
assign _1030_ = _1022_ & _1029_ /*1262*/;
assign _978_ = _1022_ ^ _1029_ /*1263*/;
assign _1027_ = _1028_ | _1030_ /*1260*/;
assign _1036_ = D[9] ^ Q[6] /*1259*/;
assign _1033_ = _881_ & _1036_ /*1255*/;
assign _1034_ = _881_ ^ _1036_ /*1258*/;
assign _1035_ = _1027_ & _1034_ /*1256*/;
assign _979_ = _1027_ ^ _1034_ /*1257*/;
assign _1032_ = _1033_ | _1035_ /*1254*/;
assign _1041_ = D[10] ^ Q[6] /*1253*/;
assign _1038_ = _882_ & _1041_ /*1249*/;
assign _1039_ = _882_ ^ _1041_ /*1252*/;
assign _1040_ = _1032_ & _1039_ /*1250*/;
assign _980_ = _1032_ ^ _1039_ /*1251*/;
assign _1037_ = _1038_ | _1040_ /*1248*/;
assign _1046_ = D[11] ^ Q[6] /*1247*/;
assign _1043_ = _883_ & _1046_ /*1243*/;
assign _1044_ = _883_ ^ _1046_ /*1246*/;
assign _1045_ = _1037_ & _1044_ /*1244*/;
assign _981_ = _1037_ ^ _1044_ /*1245*/;
assign _1042_ = _1043_ | _1045_ /*1242*/;
assign _1051_ = D[12] ^ Q[6] /*1241*/;
assign _1048_ = _884_ & _1051_ /*1237*/;
assign _1049_ = _884_ ^ _1051_ /*1240*/;
assign _1050_ = _1042_ & _1049_ /*1238*/;
assign _982_ = _1042_ ^ _1049_ /*1239*/;
assign _1047_ = _1048_ | _1050_ /*1236*/;
assign _1056_ = D[13] ^ Q[6] /*1235*/;
assign _1053_ = _885_ & _1056_ /*1231*/;
assign _1054_ = _885_ ^ _1056_ /*1234*/;
assign _1055_ = _1047_ & _1054_ /*1232*/;
assign _983_ = _1047_ ^ _1054_ /*1233*/;
assign _1052_ = _1053_ | _1055_ /*1230*/;
assign _1061_ = D[14] ^ Q[6] /*1229*/;
assign _1058_ = _886_ & _1061_ /*1225*/;
assign _1059_ = _886_ ^ _1061_ /*1228*/;
assign _1060_ = _1052_ & _1059_ /*1226*/;
assign _984_ = _1052_ ^ _1059_ /*1227*/;
assign _1057_ = _1058_ | _1060_ /*1224*/;
assign _1065_ = zeroWire ^ Q[6] /*1223*/;
assign _1062_ = _887_ & _1065_ /*1219*/;
assign _1063_ = _887_ ^ _1065_ /*1222*/;
assign _1064_ = _1057_ & _1063_ /*1220*/;
assign _985_ = _1057_ ^ _1063_ /*1221*/;
assign Q[5] = _1062_ | _1064_ /*1218*/;
assign _1088_ = D[0] ^ Q[5] /*1120*/;
assign _1085_ = R_0[4] & _1088_ /*1116*/;
assign _1086_ = R_0[4] ^ _1088_ /*1119*/;
assign _1087_ = Q[5] & _1086_ /*1117*/;
assign _1067_ = Q[5] ^ _1086_ /*1118*/;
assign _1084_ = _1085_ | _1087_ /*1115*/;
assign _1093_ = D[1] ^ Q[5] /*1114*/;
assign _1090_ = _970_ & _1093_ /*1110*/;
assign _1091_ = _970_ ^ _1093_ /*1113*/;
assign _1092_ = _1084_ & _1091_ /*1111*/;
assign _1068_ = _1084_ ^ _1091_ /*1112*/;
assign _1089_ = _1090_ | _1092_ /*1109*/;
assign _1098_ = D[2] ^ Q[5] /*1108*/;
assign _1095_ = _971_ & _1098_ /*1104*/;
assign _1096_ = _971_ ^ _1098_ /*1107*/;
assign _1097_ = _1089_ & _1096_ /*1105*/;
assign _1069_ = _1089_ ^ _1096_ /*1106*/;
assign _1094_ = _1095_ | _1097_ /*1103*/;
assign _1103_ = D[3] ^ Q[5] /*1102*/;
assign _1100_ = _972_ & _1103_ /*1098*/;
assign _1101_ = _972_ ^ _1103_ /*1101*/;
assign _1102_ = _1094_ & _1101_ /*1099*/;
assign _1070_ = _1094_ ^ _1101_ /*1100*/;
assign _1099_ = _1100_ | _1102_ /*1097*/;
assign _1108_ = D[4] ^ Q[5] /*1096*/;
assign _1105_ = _973_ & _1108_ /*1092*/;
assign _1106_ = _973_ ^ _1108_ /*1095*/;
assign _1107_ = _1099_ & _1106_ /*1093*/;
assign _1071_ = _1099_ ^ _1106_ /*1094*/;
assign _1104_ = _1105_ | _1107_ /*1091*/;
assign _1113_ = D[5] ^ Q[5] /*1090*/;
assign _1110_ = _974_ & _1113_ /*1086*/;
assign _1111_ = _974_ ^ _1113_ /*1089*/;
assign _1112_ = _1104_ & _1111_ /*1087*/;
assign _1072_ = _1104_ ^ _1111_ /*1088*/;
assign _1109_ = _1110_ | _1112_ /*1085*/;
assign _1118_ = D[6] ^ Q[5] /*1084*/;
assign _1115_ = _975_ & _1118_ /*1080*/;
assign _1116_ = _975_ ^ _1118_ /*1083*/;
assign _1117_ = _1109_ & _1116_ /*1081*/;
assign _1073_ = _1109_ ^ _1116_ /*1082*/;
assign _1114_ = _1115_ | _1117_ /*1079*/;
assign _1123_ = D[7] ^ Q[5] /*1078*/;
assign _1120_ = _976_ & _1123_ /*1074*/;
assign _1121_ = _976_ ^ _1123_ /*1077*/;
assign _1122_ = _1114_ & _1121_ /*1075*/;
assign _1074_ = _1114_ ^ _1121_ /*1076*/;
assign _1119_ = _1120_ | _1122_ /*1073*/;
assign _1128_ = D[8] ^ Q[5] /*1072*/;
assign _1125_ = _977_ & _1128_ /*1068*/;
assign _1126_ = _977_ ^ _1128_ /*1071*/;
assign _1127_ = _1119_ & _1126_ /*1069*/;
assign _1075_ = _1119_ ^ _1126_ /*1070*/;
assign _1124_ = _1125_ | _1127_ /*1067*/;
assign _1133_ = D[9] ^ Q[5] /*1066*/;
assign _1130_ = _978_ & _1133_ /*1062*/;
assign _1131_ = _978_ ^ _1133_ /*1065*/;
assign _1132_ = _1124_ & _1131_ /*1063*/;
assign _1076_ = _1124_ ^ _1131_ /*1064*/;
assign _1129_ = _1130_ | _1132_ /*1061*/;
assign _1138_ = D[10] ^ Q[5] /*1060*/;
assign _1135_ = _979_ & _1138_ /*1056*/;
assign _1136_ = _979_ ^ _1138_ /*1059*/;
assign _1137_ = _1129_ & _1136_ /*1057*/;
assign _1077_ = _1129_ ^ _1136_ /*1058*/;
assign _1134_ = _1135_ | _1137_ /*1055*/;
assign _1143_ = D[11] ^ Q[5] /*1054*/;
assign _1140_ = _980_ & _1143_ /*1050*/;
assign _1141_ = _980_ ^ _1143_ /*1053*/;
assign _1142_ = _1134_ & _1141_ /*1051*/;
assign _1078_ = _1134_ ^ _1141_ /*1052*/;
assign _1139_ = _1140_ | _1142_ /*1049*/;
assign _1148_ = D[12] ^ Q[5] /*1048*/;
assign _1145_ = _981_ & _1148_ /*1044*/;
assign _1146_ = _981_ ^ _1148_ /*1047*/;
assign _1147_ = _1139_ & _1146_ /*1045*/;
assign _1079_ = _1139_ ^ _1146_ /*1046*/;
assign _1144_ = _1145_ | _1147_ /*1043*/;
assign _1153_ = D[13] ^ Q[5] /*1042*/;
assign _1150_ = _982_ & _1153_ /*1038*/;
assign _1151_ = _982_ ^ _1153_ /*1041*/;
assign _1152_ = _1144_ & _1151_ /*1039*/;
assign _1080_ = _1144_ ^ _1151_ /*1040*/;
assign _1149_ = _1150_ | _1152_ /*1037*/;
assign _1158_ = D[14] ^ Q[5] /*1036*/;
assign _1155_ = _983_ & _1158_ /*1032*/;
assign _1156_ = _983_ ^ _1158_ /*1035*/;
assign _1157_ = _1149_ & _1156_ /*1033*/;
assign _1081_ = _1149_ ^ _1156_ /*1034*/;
assign _1154_ = _1155_ | _1157_ /*1031*/;
assign _1162_ = zeroWire ^ Q[5] /*1030*/;
assign _1159_ = _984_ & _1162_ /*1026*/;
assign _1160_ = _984_ ^ _1162_ /*1029*/;
assign _1161_ = _1154_ & _1160_ /*1027*/;
assign _1082_ = _1154_ ^ _1160_ /*1028*/;
assign Q[4] = _1159_ | _1161_ /*1025*/;
assign _1185_ = D[0] ^ Q[4] /*927*/;
assign _1182_ = R_0[3] & _1185_ /*923*/;
assign _1183_ = R_0[3] ^ _1185_ /*926*/;
assign _1184_ = Q[4] & _1183_ /*924*/;
assign _1164_ = Q[4] ^ _1183_ /*925*/;
assign _1181_ = _1182_ | _1184_ /*922*/;
assign _1190_ = D[1] ^ Q[4] /*921*/;
assign _1187_ = _1067_ & _1190_ /*917*/;
assign _1188_ = _1067_ ^ _1190_ /*920*/;
assign _1189_ = _1181_ & _1188_ /*918*/;
assign _1165_ = _1181_ ^ _1188_ /*919*/;
assign _1186_ = _1187_ | _1189_ /*916*/;
assign _1195_ = D[2] ^ Q[4] /*915*/;
assign _1192_ = _1068_ & _1195_ /*911*/;
assign _1193_ = _1068_ ^ _1195_ /*914*/;
assign _1194_ = _1186_ & _1193_ /*912*/;
assign _1166_ = _1186_ ^ _1193_ /*913*/;
assign _1191_ = _1192_ | _1194_ /*910*/;
assign _1200_ = D[3] ^ Q[4] /*909*/;
assign _1197_ = _1069_ & _1200_ /*905*/;
assign _1198_ = _1069_ ^ _1200_ /*908*/;
assign _1199_ = _1191_ & _1198_ /*906*/;
assign _1167_ = _1191_ ^ _1198_ /*907*/;
assign _1196_ = _1197_ | _1199_ /*904*/;
assign _1205_ = D[4] ^ Q[4] /*903*/;
assign _1202_ = _1070_ & _1205_ /*899*/;
assign _1203_ = _1070_ ^ _1205_ /*902*/;
assign _1204_ = _1196_ & _1203_ /*900*/;
assign _1168_ = _1196_ ^ _1203_ /*901*/;
assign _1201_ = _1202_ | _1204_ /*898*/;
assign _1210_ = D[5] ^ Q[4] /*897*/;
assign _1207_ = _1071_ & _1210_ /*893*/;
assign _1208_ = _1071_ ^ _1210_ /*896*/;
assign _1209_ = _1201_ & _1208_ /*894*/;
assign _1169_ = _1201_ ^ _1208_ /*895*/;
assign _1206_ = _1207_ | _1209_ /*892*/;
assign _1215_ = D[6] ^ Q[4] /*891*/;
assign _1212_ = _1072_ & _1215_ /*887*/;
assign _1213_ = _1072_ ^ _1215_ /*890*/;
assign _1214_ = _1206_ & _1213_ /*888*/;
assign _1170_ = _1206_ ^ _1213_ /*889*/;
assign _1211_ = _1212_ | _1214_ /*886*/;
assign _1220_ = D[7] ^ Q[4] /*885*/;
assign _1217_ = _1073_ & _1220_ /*881*/;
assign _1218_ = _1073_ ^ _1220_ /*884*/;
assign _1219_ = _1211_ & _1218_ /*882*/;
assign _1171_ = _1211_ ^ _1218_ /*883*/;
assign _1216_ = _1217_ | _1219_ /*880*/;
assign _1225_ = D[8] ^ Q[4] /*879*/;
assign _1222_ = _1074_ & _1225_ /*875*/;
assign _1223_ = _1074_ ^ _1225_ /*878*/;
assign _1224_ = _1216_ & _1223_ /*876*/;
assign _1172_ = _1216_ ^ _1223_ /*877*/;
assign _1221_ = _1222_ | _1224_ /*874*/;
assign _1230_ = D[9] ^ Q[4] /*873*/;
assign _1227_ = _1075_ & _1230_ /*869*/;
assign _1228_ = _1075_ ^ _1230_ /*872*/;
assign _1229_ = _1221_ & _1228_ /*870*/;
assign _1173_ = _1221_ ^ _1228_ /*871*/;
assign _1226_ = _1227_ | _1229_ /*868*/;
assign _1235_ = D[10] ^ Q[4] /*867*/;
assign _1232_ = _1076_ & _1235_ /*863*/;
assign _1233_ = _1076_ ^ _1235_ /*866*/;
assign _1234_ = _1226_ & _1233_ /*864*/;
assign _1174_ = _1226_ ^ _1233_ /*865*/;
assign _1231_ = _1232_ | _1234_ /*862*/;
assign _1240_ = D[11] ^ Q[4] /*861*/;
assign _1237_ = _1077_ & _1240_ /*857*/;
assign _1238_ = _1077_ ^ _1240_ /*860*/;
assign _1239_ = _1231_ & _1238_ /*858*/;
assign _1175_ = _1231_ ^ _1238_ /*859*/;
assign _1236_ = _1237_ | _1239_ /*856*/;
assign _1245_ = D[12] ^ Q[4] /*855*/;
assign _1242_ = _1078_ & _1245_ /*851*/;
assign _1243_ = _1078_ ^ _1245_ /*854*/;
assign _1244_ = _1236_ & _1243_ /*852*/;
assign _1176_ = _1236_ ^ _1243_ /*853*/;
assign _1241_ = _1242_ | _1244_ /*850*/;
assign _1250_ = D[13] ^ Q[4] /*849*/;
assign _1247_ = _1079_ & _1250_ /*845*/;
assign _1248_ = _1079_ ^ _1250_ /*848*/;
assign _1249_ = _1241_ & _1248_ /*846*/;
assign _1177_ = _1241_ ^ _1248_ /*847*/;
assign _1246_ = _1247_ | _1249_ /*844*/;
assign _1255_ = D[14] ^ Q[4] /*843*/;
assign _1252_ = _1080_ & _1255_ /*839*/;
assign _1253_ = _1080_ ^ _1255_ /*842*/;
assign _1254_ = _1246_ & _1253_ /*840*/;
assign _1178_ = _1246_ ^ _1253_ /*841*/;
assign _1251_ = _1252_ | _1254_ /*838*/;
assign _1259_ = zeroWire ^ Q[4] /*837*/;
assign _1256_ = _1081_ & _1259_ /*833*/;
assign _1257_ = _1081_ ^ _1259_ /*836*/;
assign _1258_ = _1251_ & _1257_ /*834*/;
assign _1179_ = _1251_ ^ _1257_ /*835*/;
assign Q[3] = _1256_ | _1258_ /*832*/;
assign _1282_ = D[0] ^ Q[3] /*734*/;
assign _1279_ = R_0[2] & _1282_ /*730*/;
assign _1280_ = R_0[2] ^ _1282_ /*733*/;
assign _1281_ = Q[3] & _1280_ /*731*/;
assign _1261_ = Q[3] ^ _1280_ /*732*/;
assign _1278_ = _1279_ | _1281_ /*729*/;
assign _1287_ = D[1] ^ Q[3] /*728*/;
assign _1284_ = _1164_ & _1287_ /*724*/;
assign _1285_ = _1164_ ^ _1287_ /*727*/;
assign _1286_ = _1278_ & _1285_ /*725*/;
assign _1262_ = _1278_ ^ _1285_ /*726*/;
assign _1283_ = _1284_ | _1286_ /*723*/;
assign _1292_ = D[2] ^ Q[3] /*722*/;
assign _1289_ = _1165_ & _1292_ /*718*/;
assign _1290_ = _1165_ ^ _1292_ /*721*/;
assign _1291_ = _1283_ & _1290_ /*719*/;
assign _1263_ = _1283_ ^ _1290_ /*720*/;
assign _1288_ = _1289_ | _1291_ /*717*/;
assign _1297_ = D[3] ^ Q[3] /*716*/;
assign _1294_ = _1166_ & _1297_ /*712*/;
assign _1295_ = _1166_ ^ _1297_ /*715*/;
assign _1296_ = _1288_ & _1295_ /*713*/;
assign _1264_ = _1288_ ^ _1295_ /*714*/;
assign _1293_ = _1294_ | _1296_ /*711*/;
assign _1302_ = D[4] ^ Q[3] /*710*/;
assign _1299_ = _1167_ & _1302_ /*706*/;
assign _1300_ = _1167_ ^ _1302_ /*709*/;
assign _1301_ = _1293_ & _1300_ /*707*/;
assign _1265_ = _1293_ ^ _1300_ /*708*/;
assign _1298_ = _1299_ | _1301_ /*705*/;
assign _1307_ = D[5] ^ Q[3] /*704*/;
assign _1304_ = _1168_ & _1307_ /*700*/;
assign _1305_ = _1168_ ^ _1307_ /*703*/;
assign _1306_ = _1298_ & _1305_ /*701*/;
assign _1266_ = _1298_ ^ _1305_ /*702*/;
assign _1303_ = _1304_ | _1306_ /*699*/;
assign _1312_ = D[6] ^ Q[3] /*698*/;
assign _1309_ = _1169_ & _1312_ /*694*/;
assign _1310_ = _1169_ ^ _1312_ /*697*/;
assign _1311_ = _1303_ & _1310_ /*695*/;
assign _1267_ = _1303_ ^ _1310_ /*696*/;
assign _1308_ = _1309_ | _1311_ /*693*/;
assign _1317_ = D[7] ^ Q[3] /*692*/;
assign _1314_ = _1170_ & _1317_ /*688*/;
assign _1315_ = _1170_ ^ _1317_ /*691*/;
assign _1316_ = _1308_ & _1315_ /*689*/;
assign _1268_ = _1308_ ^ _1315_ /*690*/;
assign _1313_ = _1314_ | _1316_ /*687*/;
assign _1322_ = D[8] ^ Q[3] /*686*/;
assign _1319_ = _1171_ & _1322_ /*682*/;
assign _1320_ = _1171_ ^ _1322_ /*685*/;
assign _1321_ = _1313_ & _1320_ /*683*/;
assign _1269_ = _1313_ ^ _1320_ /*684*/;
assign _1318_ = _1319_ | _1321_ /*681*/;
assign _1327_ = D[9] ^ Q[3] /*680*/;
assign _1324_ = _1172_ & _1327_ /*676*/;
assign _1325_ = _1172_ ^ _1327_ /*679*/;
assign _1326_ = _1318_ & _1325_ /*677*/;
assign _1270_ = _1318_ ^ _1325_ /*678*/;
assign _1323_ = _1324_ | _1326_ /*675*/;
assign _1332_ = D[10] ^ Q[3] /*674*/;
assign _1329_ = _1173_ & _1332_ /*670*/;
assign _1330_ = _1173_ ^ _1332_ /*673*/;
assign _1331_ = _1323_ & _1330_ /*671*/;
assign _1271_ = _1323_ ^ _1330_ /*672*/;
assign _1328_ = _1329_ | _1331_ /*669*/;
assign _1337_ = D[11] ^ Q[3] /*668*/;
assign _1334_ = _1174_ & _1337_ /*664*/;
assign _1335_ = _1174_ ^ _1337_ /*667*/;
assign _1336_ = _1328_ & _1335_ /*665*/;
assign _1272_ = _1328_ ^ _1335_ /*666*/;
assign _1333_ = _1334_ | _1336_ /*663*/;
assign _1342_ = D[12] ^ Q[3] /*662*/;
assign _1339_ = _1175_ & _1342_ /*658*/;
assign _1340_ = _1175_ ^ _1342_ /*661*/;
assign _1341_ = _1333_ & _1340_ /*659*/;
assign _1273_ = _1333_ ^ _1340_ /*660*/;
assign _1338_ = _1339_ | _1341_ /*657*/;
assign _1347_ = D[13] ^ Q[3] /*656*/;
assign _1344_ = _1176_ & _1347_ /*652*/;
assign _1345_ = _1176_ ^ _1347_ /*655*/;
assign _1346_ = _1338_ & _1345_ /*653*/;
assign _1274_ = _1338_ ^ _1345_ /*654*/;
assign _1343_ = _1344_ | _1346_ /*651*/;
assign _1352_ = D[14] ^ Q[3] /*650*/;
assign _1349_ = _1177_ & _1352_ /*646*/;
assign _1350_ = _1177_ ^ _1352_ /*649*/;
assign _1351_ = _1343_ & _1350_ /*647*/;
assign _1275_ = _1343_ ^ _1350_ /*648*/;
assign _1348_ = _1349_ | _1351_ /*645*/;
assign _1356_ = zeroWire ^ Q[3] /*644*/;
assign _1353_ = _1178_ & _1356_ /*640*/;
assign _1354_ = _1178_ ^ _1356_ /*643*/;
assign _1355_ = _1348_ & _1354_ /*641*/;
assign _1276_ = _1348_ ^ _1354_ /*642*/;
assign Q[2] = _1353_ | _1355_ /*639*/;
assign _1379_ = D[0] ^ Q[2] /*541*/;
assign _1376_ = R_0[1] & _1379_ /*537*/;
assign _1377_ = R_0[1] ^ _1379_ /*540*/;
assign _1378_ = Q[2] & _1377_ /*538*/;
assign _1358_ = Q[2] ^ _1377_ /*539*/;
assign _1375_ = _1376_ | _1378_ /*536*/;
assign _1384_ = D[1] ^ Q[2] /*535*/;
assign _1381_ = _1261_ & _1384_ /*531*/;
assign _1382_ = _1261_ ^ _1384_ /*534*/;
assign _1383_ = _1375_ & _1382_ /*532*/;
assign _1359_ = _1375_ ^ _1382_ /*533*/;
assign _1380_ = _1381_ | _1383_ /*530*/;
assign _1389_ = D[2] ^ Q[2] /*529*/;
assign _1386_ = _1262_ & _1389_ /*525*/;
assign _1387_ = _1262_ ^ _1389_ /*528*/;
assign _1388_ = _1380_ & _1387_ /*526*/;
assign _1360_ = _1380_ ^ _1387_ /*527*/;
assign _1385_ = _1386_ | _1388_ /*524*/;
assign _1394_ = D[3] ^ Q[2] /*523*/;
assign _1391_ = _1263_ & _1394_ /*519*/;
assign _1392_ = _1263_ ^ _1394_ /*522*/;
assign _1393_ = _1385_ & _1392_ /*520*/;
assign _1361_ = _1385_ ^ _1392_ /*521*/;
assign _1390_ = _1391_ | _1393_ /*518*/;
assign _1399_ = D[4] ^ Q[2] /*517*/;
assign _1396_ = _1264_ & _1399_ /*513*/;
assign _1397_ = _1264_ ^ _1399_ /*516*/;
assign _1398_ = _1390_ & _1397_ /*514*/;
assign _1362_ = _1390_ ^ _1397_ /*515*/;
assign _1395_ = _1396_ | _1398_ /*512*/;
assign _1404_ = D[5] ^ Q[2] /*511*/;
assign _1401_ = _1265_ & _1404_ /*507*/;
assign _1402_ = _1265_ ^ _1404_ /*510*/;
assign _1403_ = _1395_ & _1402_ /*508*/;
assign _1363_ = _1395_ ^ _1402_ /*509*/;
assign _1400_ = _1401_ | _1403_ /*506*/;
assign _1409_ = D[6] ^ Q[2] /*505*/;
assign _1406_ = _1266_ & _1409_ /*501*/;
assign _1407_ = _1266_ ^ _1409_ /*504*/;
assign _1408_ = _1400_ & _1407_ /*502*/;
assign _1364_ = _1400_ ^ _1407_ /*503*/;
assign _1405_ = _1406_ | _1408_ /*500*/;
assign _1414_ = D[7] ^ Q[2] /*499*/;
assign _1411_ = _1267_ & _1414_ /*495*/;
assign _1412_ = _1267_ ^ _1414_ /*498*/;
assign _1413_ = _1405_ & _1412_ /*496*/;
assign _1365_ = _1405_ ^ _1412_ /*497*/;
assign _1410_ = _1411_ | _1413_ /*494*/;
assign _1419_ = D[8] ^ Q[2] /*493*/;
assign _1416_ = _1268_ & _1419_ /*489*/;
assign _1417_ = _1268_ ^ _1419_ /*492*/;
assign _1418_ = _1410_ & _1417_ /*490*/;
assign _1366_ = _1410_ ^ _1417_ /*491*/;
assign _1415_ = _1416_ | _1418_ /*488*/;
assign _1424_ = D[9] ^ Q[2] /*487*/;
assign _1421_ = _1269_ & _1424_ /*483*/;
assign _1422_ = _1269_ ^ _1424_ /*486*/;
assign _1423_ = _1415_ & _1422_ /*484*/;
assign _1367_ = _1415_ ^ _1422_ /*485*/;
assign _1420_ = _1421_ | _1423_ /*482*/;
assign _1429_ = D[10] ^ Q[2] /*481*/;
assign _1426_ = _1270_ & _1429_ /*477*/;
assign _1427_ = _1270_ ^ _1429_ /*480*/;
assign _1428_ = _1420_ & _1427_ /*478*/;
assign _1368_ = _1420_ ^ _1427_ /*479*/;
assign _1425_ = _1426_ | _1428_ /*476*/;
assign _1434_ = D[11] ^ Q[2] /*475*/;
assign _1431_ = _1271_ & _1434_ /*471*/;
assign _1432_ = _1271_ ^ _1434_ /*474*/;
assign _1433_ = _1425_ & _1432_ /*472*/;
assign _1369_ = _1425_ ^ _1432_ /*473*/;
assign _1430_ = _1431_ | _1433_ /*470*/;
assign _1439_ = D[12] ^ Q[2] /*469*/;
assign _1436_ = _1272_ & _1439_ /*465*/;
assign _1437_ = _1272_ ^ _1439_ /*468*/;
assign _1438_ = _1430_ & _1437_ /*466*/;
assign _1370_ = _1430_ ^ _1437_ /*467*/;
assign _1435_ = _1436_ | _1438_ /*464*/;
assign _1444_ = D[13] ^ Q[2] /*463*/;
assign _1441_ = _1273_ & _1444_ /*459*/;
assign _1442_ = _1273_ ^ _1444_ /*462*/;
assign _1443_ = _1435_ & _1442_ /*460*/;
assign _1371_ = _1435_ ^ _1442_ /*461*/;
assign _1440_ = _1441_ | _1443_ /*458*/;
assign _1449_ = D[14] ^ Q[2] /*457*/;
assign _1446_ = _1274_ & _1449_ /*453*/;
assign _1447_ = _1274_ ^ _1449_ /*456*/;
assign _1448_ = _1440_ & _1447_ /*454*/;
assign _1372_ = _1440_ ^ _1447_ /*455*/;
assign _1445_ = _1446_ | _1448_ /*452*/;
assign _1453_ = zeroWire ^ Q[2] /*451*/;
assign _1450_ = _1275_ & _1453_ /*447*/;
assign _1451_ = _1275_ ^ _1453_ /*450*/;
assign _1452_ = _1445_ & _1451_ /*448*/;
assign _1373_ = _1445_ ^ _1451_ /*449*/;
assign Q[1] = _1450_ | _1452_ /*446*/;
assign _1476_ = D[0] ^ Q[1] /*348*/;
assign _1473_ = R_0[0] & _1476_ /*344*/;
assign _1474_ = R_0[0] ^ _1476_ /*347*/;
assign _1475_ = Q[1] & _1474_ /*345*/;
assign _1455_ = Q[1] ^ _1474_ /*346*/;
assign _1472_ = _1473_ | _1475_ /*343*/;
assign _1481_ = D[1] ^ Q[1] /*342*/;
assign _1478_ = _1358_ & _1481_ /*338*/;
assign _1479_ = _1358_ ^ _1481_ /*341*/;
assign _1480_ = _1472_ & _1479_ /*339*/;
assign _1456_ = _1472_ ^ _1479_ /*340*/;
assign _1477_ = _1478_ | _1480_ /*337*/;
assign _1486_ = D[2] ^ Q[1] /*336*/;
assign _1483_ = _1359_ & _1486_ /*332*/;
assign _1484_ = _1359_ ^ _1486_ /*335*/;
assign _1485_ = _1477_ & _1484_ /*333*/;
assign _1457_ = _1477_ ^ _1484_ /*334*/;
assign _1482_ = _1483_ | _1485_ /*331*/;
assign _1491_ = D[3] ^ Q[1] /*330*/;
assign _1488_ = _1360_ & _1491_ /*326*/;
assign _1489_ = _1360_ ^ _1491_ /*329*/;
assign _1490_ = _1482_ & _1489_ /*327*/;
assign _1458_ = _1482_ ^ _1489_ /*328*/;
assign _1487_ = _1488_ | _1490_ /*325*/;
assign _1496_ = D[4] ^ Q[1] /*324*/;
assign _1493_ = _1361_ & _1496_ /*320*/;
assign _1494_ = _1361_ ^ _1496_ /*323*/;
assign _1495_ = _1487_ & _1494_ /*321*/;
assign _1459_ = _1487_ ^ _1494_ /*322*/;
assign _1492_ = _1493_ | _1495_ /*319*/;
assign _1501_ = D[5] ^ Q[1] /*318*/;
assign _1498_ = _1362_ & _1501_ /*314*/;
assign _1499_ = _1362_ ^ _1501_ /*317*/;
assign _1500_ = _1492_ & _1499_ /*315*/;
assign _1460_ = _1492_ ^ _1499_ /*316*/;
assign _1497_ = _1498_ | _1500_ /*313*/;
assign _1506_ = D[6] ^ Q[1] /*312*/;
assign _1503_ = _1363_ & _1506_ /*308*/;
assign _1504_ = _1363_ ^ _1506_ /*311*/;
assign _1505_ = _1497_ & _1504_ /*309*/;
assign _1461_ = _1497_ ^ _1504_ /*310*/;
assign _1502_ = _1503_ | _1505_ /*307*/;
assign _1511_ = D[7] ^ Q[1] /*306*/;
assign _1508_ = _1364_ & _1511_ /*302*/;
assign _1509_ = _1364_ ^ _1511_ /*305*/;
assign _1510_ = _1502_ & _1509_ /*303*/;
assign _1462_ = _1502_ ^ _1509_ /*304*/;
assign _1507_ = _1508_ | _1510_ /*301*/;
assign _1516_ = D[8] ^ Q[1] /*300*/;
assign _1513_ = _1365_ & _1516_ /*296*/;
assign _1514_ = _1365_ ^ _1516_ /*299*/;
assign _1515_ = _1507_ & _1514_ /*297*/;
assign _1463_ = _1507_ ^ _1514_ /*298*/;
assign _1512_ = _1513_ | _1515_ /*295*/;
assign _1521_ = D[9] ^ Q[1] /*294*/;
assign _1518_ = _1366_ & _1521_ /*290*/;
assign _1519_ = _1366_ ^ _1521_ /*293*/;
assign _1520_ = _1512_ & _1519_ /*291*/;
assign _1464_ = _1512_ ^ _1519_ /*292*/;
assign _1517_ = _1518_ | _1520_ /*289*/;
assign _1526_ = D[10] ^ Q[1] /*288*/;
assign _1523_ = _1367_ & _1526_ /*284*/;
assign _1524_ = _1367_ ^ _1526_ /*287*/;
assign _1525_ = _1517_ & _1524_ /*285*/;
assign _1465_ = _1517_ ^ _1524_ /*286*/;
assign _1522_ = _1523_ | _1525_ /*283*/;
assign _1531_ = D[11] ^ Q[1] /*282*/;
assign _1528_ = _1368_ & _1531_ /*278*/;
assign _1529_ = _1368_ ^ _1531_ /*281*/;
assign _1530_ = _1522_ & _1529_ /*279*/;
assign _1466_ = _1522_ ^ _1529_ /*280*/;
assign _1527_ = _1528_ | _1530_ /*277*/;
assign _1536_ = D[12] ^ Q[1] /*276*/;
assign _1533_ = _1369_ & _1536_ /*272*/;
assign _1534_ = _1369_ ^ _1536_ /*275*/;
assign _1535_ = _1527_ & _1534_ /*273*/;
assign _1467_ = _1527_ ^ _1534_ /*274*/;
assign _1532_ = _1533_ | _1535_ /*271*/;
assign _1541_ = D[13] ^ Q[1] /*270*/;
assign _1538_ = _1370_ & _1541_ /*266*/;
assign _1539_ = _1370_ ^ _1541_ /*269*/;
assign _1540_ = _1532_ & _1539_ /*267*/;
assign _1468_ = _1532_ ^ _1539_ /*268*/;
assign _1537_ = _1538_ | _1540_ /*265*/;
assign _1546_ = D[14] ^ Q[1] /*264*/;
assign _1543_ = _1371_ & _1546_ /*260*/;
assign _1544_ = _1371_ ^ _1546_ /*263*/;
assign _1545_ = _1537_ & _1544_ /*261*/;
assign _1469_ = _1537_ ^ _1544_ /*262*/;
assign _1542_ = _1543_ | _1545_ /*259*/;
assign _1550_ = zeroWire ^ Q[1] /*258*/;
assign _1547_ = _1372_ & _1550_ /*254*/;
assign _1548_ = _1372_ ^ _1550_ /*257*/;
assign _1549_ = _1542_ & _1548_ /*255*/;
assign _1470_ = _1542_ ^ _1548_ /*256*/;
assign Q[0] = _1547_ | _1549_ /*253*/;
assign _1554_ = ~Q[0] /*154*/;
assign _1553_ = _1554_ & D[0] /*153*/;
assign _1556_ = _1455_ & _1553_ /*148*/;
assign _1557_ = _1455_ ^ _1553_ /*151*/;
assign _1558_ = zeroWire & _1557_ /*149*/;
assign R_n1[0] = zeroWire ^ _1557_ /*150*/;
assign _1555_ = _1556_ | _1558_ /*147*/;
assign _1560_ = ~Q[0] /*146*/;
assign _1559_ = _1560_ & D[1] /*145*/;
assign _1562_ = _1456_ & _1559_ /*140*/;
assign _1563_ = _1456_ ^ _1559_ /*143*/;
assign _1564_ = _1555_ & _1563_ /*141*/;
assign R_n1[1] = _1555_ ^ _1563_ /*142*/;
assign _1561_ = _1562_ | _1564_ /*139*/;
assign _1566_ = ~Q[0] /*138*/;
assign _1565_ = _1566_ & D[2] /*137*/;
assign _1568_ = _1457_ & _1565_ /*132*/;
assign _1569_ = _1457_ ^ _1565_ /*135*/;
assign _1570_ = _1561_ & _1569_ /*133*/;
assign R_n1[2] = _1561_ ^ _1569_ /*134*/;
assign _1567_ = _1568_ | _1570_ /*131*/;
assign _1572_ = ~Q[0] /*130*/;
assign _1571_ = _1572_ & D[3] /*129*/;
assign _1574_ = _1458_ & _1571_ /*124*/;
assign _1575_ = _1458_ ^ _1571_ /*127*/;
assign _1576_ = _1567_ & _1575_ /*125*/;
assign R_n1[3] = _1567_ ^ _1575_ /*126*/;
assign _1573_ = _1574_ | _1576_ /*123*/;
assign _1578_ = ~Q[0] /*122*/;
assign _1577_ = _1578_ & D[4] /*121*/;
assign _1580_ = _1459_ & _1577_ /*116*/;
assign _1581_ = _1459_ ^ _1577_ /*119*/;
assign _1582_ = _1573_ & _1581_ /*117*/;
assign R_n1[4] = _1573_ ^ _1581_ /*118*/;
assign _1579_ = _1580_ | _1582_ /*115*/;
assign _1584_ = ~Q[0] /*114*/;
assign _1583_ = _1584_ & D[5] /*113*/;
assign _1586_ = _1460_ & _1583_ /*108*/;
assign _1587_ = _1460_ ^ _1583_ /*111*/;
assign _1588_ = _1579_ & _1587_ /*109*/;
assign R_n1[5] = _1579_ ^ _1587_ /*110*/;
assign _1585_ = _1586_ | _1588_ /*107*/;
assign _1590_ = ~Q[0] /*106*/;
assign _1589_ = _1590_ & D[6] /*105*/;
assign _1592_ = _1461_ & _1589_ /*100*/;
assign _1593_ = _1461_ ^ _1589_ /*103*/;
assign _1594_ = _1585_ & _1593_ /*101*/;
assign R_n1[6] = _1585_ ^ _1593_ /*102*/;
assign _1591_ = _1592_ | _1594_ /*99*/;
assign _1596_ = ~Q[0] /*98*/;
assign _1595_ = _1596_ & D[7] /*97*/;
assign _1598_ = _1462_ & _1595_ /*92*/;
assign _1599_ = _1462_ ^ _1595_ /*95*/;
assign _1600_ = _1591_ & _1599_ /*93*/;
assign R_n1[7] = _1591_ ^ _1599_ /*94*/;
assign _1597_ = _1598_ | _1600_ /*91*/;
assign _1602_ = ~Q[0] /*90*/;
assign _1601_ = _1602_ & D[8] /*89*/;
assign _1604_ = _1463_ & _1601_ /*84*/;
assign _1605_ = _1463_ ^ _1601_ /*87*/;
assign _1606_ = _1597_ & _1605_ /*85*/;
assign R_n1[8] = _1597_ ^ _1605_ /*86*/;
assign _1603_ = _1604_ | _1606_ /*83*/;
assign _1608_ = ~Q[0] /*82*/;
assign _1607_ = _1608_ & D[9] /*81*/;
assign _1610_ = _1464_ & _1607_ /*76*/;
assign _1611_ = _1464_ ^ _1607_ /*79*/;
assign _1612_ = _1603_ & _1611_ /*77*/;
assign R_n1[9] = _1603_ ^ _1611_ /*78*/;
assign _1609_ = _1610_ | _1612_ /*75*/;
assign _1614_ = ~Q[0] /*74*/;
assign _1613_ = _1614_ & D[10] /*73*/;
assign _1616_ = _1465_ & _1613_ /*68*/;
assign _1617_ = _1465_ ^ _1613_ /*71*/;
assign _1618_ = _1609_ & _1617_ /*69*/;
assign R_n1[10] = _1609_ ^ _1617_ /*70*/;
assign _1615_ = _1616_ | _1618_ /*67*/;
assign _1620_ = ~Q[0] /*66*/;
assign _1619_ = _1620_ & D[11] /*65*/;
assign _1622_ = _1466_ & _1619_ /*60*/;
assign _1623_ = _1466_ ^ _1619_ /*63*/;
assign _1624_ = _1615_ & _1623_ /*61*/;
assign R_n1[11] = _1615_ ^ _1623_ /*62*/;
assign _1621_ = _1622_ | _1624_ /*59*/;
assign _1626_ = ~Q[0] /*58*/;
assign _1625_ = _1626_ & D[12] /*57*/;
assign _1628_ = _1467_ & _1625_ /*52*/;
assign _1629_ = _1467_ ^ _1625_ /*55*/;
assign _1630_ = _1621_ & _1629_ /*53*/;
assign R_n1[12] = _1621_ ^ _1629_ /*54*/;
assign _1627_ = _1628_ | _1630_ /*51*/;
assign _1632_ = ~Q[0] /*50*/;
assign _1631_ = _1632_ & D[13] /*49*/;
assign _1634_ = _1468_ & _1631_ /*44*/;
assign _1635_ = _1468_ ^ _1631_ /*47*/;
assign _1636_ = _1627_ & _1635_ /*45*/;
assign R_n1[13] = _1627_ ^ _1635_ /*46*/;
assign _1633_ = _1634_ | _1636_ /*43*/;
assign _1638_ = ~Q[0] /*42*/;
assign _1637_ = _1638_ & D[14] /*41*/;
assign _1640_ = _1469_ & _1637_ /*36*/;
assign _1641_ = _1469_ ^ _1637_ /*39*/;
assign _1642_ = _1633_ & _1641_ /*37*/;
assign R_n1[14] = _1633_ ^ _1641_ /*38*/;
assign _1639_ = _1640_ | _1642_ /*35*/;
endmodule
