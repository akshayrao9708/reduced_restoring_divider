module divider(q, rout, rin, div);
  wire _0_;
  wire _1_;
  wire _2_;
  wire _3_;
  wire _4_;
  wire _5_;
  wire _6_;
  wire _7_;
  wire _8_;
  wire _9_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  wire _38_;
  wire _39_;
  wire _40_;
  wire _41_;
  wire _42_;
  wire _43_;
  wire _44_;
  wire _45_;
  wire _46_;
  wire _47_;
  wire _48_;
  wire _49_;
  wire _50_;
  wire _51_;
  wire _52_;
  wire _53_;
  wire _54_;
  wire _55_;
  wire _56_;
  wire _57_;
  wire _58_;
  wire _59_;
  wire _60_;
  wire _61_;
  wire _62_;
  wire _63_;
  wire _64_;
  wire _65_;
  wire _66_;
  wire _67_;
  wire _68_;
  wire _69_;
  wire _70_;
  wire _71_;
  wire _72_;
  wire _73_;
  wire _74_;
  wire _75_;
  wire _76_;
  wire _77_;
  wire _78_;
  wire _79_;
  wire _80_;
  wire _81_;
  wire _82_;
  wire _83_;
  wire _84_;
  wire _85_;
  wire _86_;
  wire _87_;
  wire _88_;
  wire _89_;
  wire _90_;
  wire _91_;
  wire _92_;
  wire _93_;
  wire _94_;
  wire _95_;
  wire _96_;
  wire _97_;
  wire _98_;
  wire _99_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire _304_;
  wire _305_;
  wire _306_;
  wire _307_;
  wire _308_;
  wire _309_;
  wire _310_;
  wire _311_;
  wire _312_;
  wire _313_;
  wire _314_;
  wire _315_;
  wire _316_;
  wire _317_;
  wire _318_;
  wire _319_;
  wire _320_;
  wire _321_;
  wire _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire _326_;
  wire _327_;
  wire _328_;
  wire _329_;
  wire _330_;
  wire _331_;
  wire _332_;
  wire _333_;
  wire _334_;
  wire _335_;
  wire _336_;
  wire _337_;
  wire _338_;
  wire _339_;
  wire _340_;
  wire _341_;
  wire _342_;
  wire _343_;
  wire _344_;
  wire _345_;
  wire _346_;
  wire _347_;
  wire _348_;
  wire _349_;
  wire _350_;
  wire _351_;
  wire _352_;
  wire _353_;
  wire _354_;
  wire _355_;
  wire _356_;
  wire _357_;
  wire _358_;
  wire _359_;
  wire _360_;
  wire _361_;
  wire _362_;
  wire _363_;
  wire _364_;
  wire _365_;
  wire _366_;
  wire _367_;
  wire _368_;
  wire _369_;
  wire _370_;
  wire _371_;
  wire _372_;
  wire _373_;
  wire _374_;
  wire _375_;
  wire _376_;
  wire _377_;
  wire _378_;
  wire _379_;
  wire _380_;
  wire _381_;
  wire _382_;
  wire _383_;
  wire _384_;
  wire _385_;
  wire _386_;
  wire _387_;
  wire _388_;
  wire _389_;
  wire _390_;
  wire _391_;
  wire _392_;
  wire _393_;
  wire _394_;
  wire _395_;
  wire _396_;
  wire _397_;
  wire _398_;
  wire _399_;
  wire _400_;
  wire _401_;
  wire _402_;
  wire _403_;
  wire _404_;
  wire _405_;
  wire _406_;
  wire _407_;
  wire _408_;
  wire _409_;
  wire _410_;
  wire _411_;
  wire _412_;
  wire _413_;
  wire _414_;
  wire _415_;
  wire _416_;
  wire _417_;
  wire _418_;
  wire _419_;
  wire _420_;
  wire _421_;
  wire _422_;
  wire _423_;
  wire _424_;
  wire _425_;
  wire _426_;
  wire _427_;
  wire _428_;
  wire _429_;
  wire _430_;
  wire _431_;
  wire _432_;
  wire _433_;
  wire _434_;
  wire _435_;
  wire _436_;
  wire _437_;
  wire _438_;
  wire _439_;
  wire _440_;
  wire _441_;
  wire _442_;
  wire _443_;
  wire _444_;
  wire _445_;
  wire _446_;
  wire _447_;
  wire _448_;
  wire _449_;
  wire _450_;
  wire _451_;
  wire _452_;
  wire _453_;
  wire _454_;
  wire _455_;
  wire _456_;
  wire _457_;
  wire _458_;
  wire _459_;
  wire _460_;
  wire _461_;
  wire _462_;
  wire _463_;
  wire _464_;
  wire _465_;
  wire _466_;
  wire _467_;
  wire _468_;
  wire _469_;
  wire _470_;
  wire _471_;
  wire _472_;
  wire _473_;
  wire _474_;
  wire _475_;
  wire _476_;
  wire _477_;
  wire _478_;
  wire _479_;
  wire _480_;
  wire _481_;
  wire _482_;
  wire _483_;
  wire _484_;
  wire _485_;
  wire _486_;
  wire _487_;
  wire _488_;
  wire _489_;
  wire _490_;
  wire _491_;
  wire _492_;
  wire _493_;
  wire _494_;
  wire _495_;
  wire _496_;
  wire _497_;
  wire _498_;
  wire _499_;
  wire _500_;
  wire _501_;
  wire _502_;
  wire _503_;
  wire _504_;
  wire _505_;
  wire _506_;
  wire _507_;
  wire _508_;
  wire _509_;
  wire _510_;
  wire _511_;
  wire _512_;
  wire _513_;
  wire _514_;
  wire _515_;
  wire _516_;
  wire _517_;
  wire _518_;
  wire _519_;
  wire _520_;
  wire _521_;
  wire _522_;
  wire _523_;
  wire _524_;
  wire _525_;
  wire _526_;
  wire _527_;
  wire _528_;
  wire _529_;
  wire _530_;
  wire _531_;
  wire _532_;
  wire _533_;
  wire _534_;
  wire _535_;
  wire _536_;
  wire _537_;
  wire _538_;
  wire _539_;
  wire _540_;
  wire _541_;
  wire _542_;
  wire _543_;
  wire _544_;
  wire _545_;
  wire _546_;
  wire _547_;
  wire _548_;
  wire _549_;
  wire _550_;
  wire _551_;
  wire _552_;
  wire _553_;
  wire _554_;
  wire _555_;
  wire _556_;
  wire _557_;
  wire _558_;
  wire _559_;
  wire _560_;
  wire _561_;
  wire _562_;
  wire _563_;
  wire _564_;
  wire _565_;
  wire _566_;
  wire _567_;
  wire _568_;
  wire _569_;
  wire _570_;
  wire _571_;
  wire _572_;
  wire _573_;
  wire _574_;
  wire _575_;
  wire _576_;
  wire _577_;
  wire _578_;
  wire _579_;
  wire _580_;
  wire _581_;
  wire _582_;
  wire _583_;
  wire _584_;
  wire _585_;
  wire _586_;
  wire _587_;
  wire _588_;
  wire _589_;
  wire _590_;
  wire _591_;
  wire _592_;
  wire _593_;
  wire _594_;
  wire _595_;
  wire _596_;
  wire _597_;
  wire _598_;
  wire _599_;
  wire _600_;
  wire _601_;
  wire _602_;
  wire _603_;
  wire _604_;
  wire _605_;
  wire _606_;
  wire _607_;
  wire _608_;
  wire _609_;
  wire _610_;
  wire _611_;
  wire _612_;
  wire _613_;
  wire _614_;
  wire _615_;
  wire _616_;
  wire _617_;
  wire _618_;
  wire _619_;
  wire _620_;
  wire _621_;
  wire _622_;
  wire _623_;
  wire _624_;
  wire _625_;
  wire _626_;
  wire _627_;
  wire _628_;
  wire _629_;
  wire _630_;
  wire _631_;
  wire _632_;
  wire _633_;
  wire _634_;
  wire _635_;
  wire _636_;
  wire _637_;
  wire _638_;
  wire _639_;
  wire _640_;
  wire _641_;
  wire _642_;
  wire _643_;
  wire _644_;
  wire _645_;
  wire _646_;
  wire _647_;
  wire _648_;
  wire _649_;
  wire _650_;
  wire _651_;
  wire _652_;
  wire _653_;
  wire _654_;
  wire _655_;
  wire _656_;
  wire _657_;
  wire _658_;
  wire _659_;
  wire _660_;
  wire _661_;
  wire _662_;
  wire _663_;
  wire _664_;
  wire _665_;
  wire _666_;
  wire _667_;
  wire _668_;
  wire _669_;
  wire _670_;
  wire _671_;
  wire _672_;
  wire _673_;
  wire _674_;
  wire _675_;
  wire _676_;
  wire _677_;
  wire _678_;
  wire _679_;
  wire _680_;
  wire _681_;
  wire _682_;
  wire _683_;
  wire _684_;
  wire _685_;
  wire _686_;
  wire _687_;
  wire _688_;
  wire _689_;
  wire _690_;
  wire _691_;
  wire _692_;
  wire _693_;
  wire _694_;
  wire _695_;
  wire _696_;
  wire _697_;
  wire _698_;
  wire _699_;
  wire _700_;
  wire _701_;
  wire _702_;
  wire _703_;
  wire _704_;
  wire _705_;
  wire _706_;
  wire _707_;
  wire _708_;
  wire _709_;
  wire _710_;
  wire _711_;
  wire _712_;
  wire _713_;
  wire _714_;
  wire _715_;
  wire _716_;
  wire _717_;
  wire _718_;
  wire _719_;
  wire _720_;
  wire _721_;
  wire _722_;
  wire _723_;
  wire _724_;
  wire _725_;
  wire _726_;
  wire _727_;
  wire _728_;
  wire _729_;
  wire _730_;
  wire _731_;
  wire _732_;
  wire _733_;
  wire _734_;
  wire _735_;
  wire _736_;
  wire _737_;
  wire _738_;
  wire _739_;
  wire _740_;
  wire _741_;
  wire _742_;
  wire _743_;
  wire _744_;
  wire _745_;
  wire _746_;
  wire _747_;
  wire _748_;
  wire _749_;
  wire _750_;
  wire _751_;
  wire _752_;
  wire _753_;
  wire _754_;
  wire _755_;
  wire _756_;
  wire _757_;
  wire _758_;
  wire _759_;
  wire _760_;
  wire _761_;
  wire _762_;
  wire _763_;
  wire _764_;
  wire _765_;
  wire _766_;
  wire _767_;
  wire _768_;
  wire _769_;
  wire _770_;
  wire _771_;
  wire _772_;
  wire _773_;
  wire _774_;
  wire _775_;
  wire _776_;
  wire _777_;
  wire _778_;
  wire _779_;
  wire _780_;
  wire _781_;
  wire _782_;
  wire _783_;
  wire _784_;
  wire _785_;
  wire _786_;
  wire _787_;
  wire _788_;
  wire _789_;
  wire _790_;
  wire _791_;
  wire _792_;
  wire _793_;
  wire _794_;
  wire _795_;
  wire _796_;
  wire _797_;
  wire _798_;
  wire _799_;
  wire _800_;
  wire _801_;
  wire _802_;
  wire _803_;
  wire _804_;
  wire _805_;
  wire _806_;
  wire _807_;
  wire _808_;
  wire _809_;
  wire _810_;
  wire _811_;
  wire _812_;
  wire _813_;
  wire _814_;
  wire _815_;
  wire _816_;
  wire _817_;
  wire _818_;
  wire _819_;
  wire _820_;
  wire _821_;
  wire _822_;
  wire _823_;
  wire _824_;
  wire _825_;
  wire _826_;
  wire _827_;
  wire _828_;
  wire _829_;
  wire _830_;
  wire _831_;
  wire _832_;
  wire _833_;
  wire _834_;
  wire _835_;
  wire _836_;
  wire _837_;
  wire _838_;
  wire _839_;
  wire _840_;
  wire _841_;
  wire _842_;
  wire _843_;
  wire _844_;
  wire _845_;
  wire _846_;
  wire _847_;
  wire _848_;
  wire _849_;
  wire _850_;
  wire _851_;
  wire _852_;
  wire _853_;
  wire _854_;
  wire _855_;
  wire _856_;
  wire _857_;
  wire _858_;
  wire _859_;
  wire _860_;
  wire _861_;
  wire _862_;
  wire _863_;
  wire _864_;
  wire _865_;
  wire _866_;
  wire _867_;
  wire _868_;
  wire _869_;
  wire _870_;
  wire _871_;
  wire _872_;
  wire _873_;
  wire _874_;
  wire _875_;
  wire _876_;
  wire _877_;
  wire _878_;
  wire _879_;
  wire _880_;
  wire _881_;
  wire _882_;
  wire _883_;
  wire _884_;
  wire _885_;
  wire _886_;
  wire _887_;
  wire _888_;
  wire _889_;
  wire _890_;
  wire _891_;
  wire _892_;
  wire _893_;
  wire _894_;
  wire _895_;
  wire _896_;
  wire _897_;
  wire _898_;
  wire _899_;
  wire _900_;
  wire _901_;
  wire _902_;
  wire _903_;
  wire _904_;
  wire _905_;
  wire _906_;
  wire _907_;
  wire _908_;
  wire _909_;
  wire _910_;
  wire _911_;
  wire _912_;
  wire _913_;
  wire _914_;
  wire _915_;
  wire _916_;
  wire _917_;
  wire _918_;
  wire _919_;
  wire _920_;
  wire _921_;
  wire _922_;
  wire _923_;
  wire _924_;
  wire _925_;
  wire _926_;
  wire _927_;
  wire _928_;
  wire _929_;
  wire _930_;
  wire _931_;
  wire _932_;
  wire _933_;
  wire _934_;
  wire _935_;
  wire _936_;
  wire _937_;
  wire _938_;
  wire _939_;
  wire _940_;
  wire _941_;
  wire _942_;
  wire _943_;
  wire _944_;
  wire _945_;
  wire _946_;
  wire _947_;
  wire _948_;
  wire _949_;
  wire _950_;
  wire _951_;
  wire _952_;
  wire _953_;
  wire _954_;
  wire _955_;
  wire _956_;
  wire _957_;
  wire _958_;
  wire _959_;
  wire _960_;
  wire _961_;
  wire _962_;
  wire _963_;
  wire _964_;
  wire _965_;
  wire _966_;
  wire _967_;
  wire _968_;
  wire _969_;
  wire _970_;
  wire _971_;
  wire _972_;
  wire _973_;
  wire _974_;
  wire _975_;
  wire _976_;
  wire _977_;
  wire _978_;
  wire _979_;
  wire _980_;
  wire _981_;
  wire _982_;
  wire _983_;
  wire _984_;
  wire _985_;
  wire _986_;
  wire _987_;
  wire _988_;
  wire _989_;
  wire _990_;
  wire _991_;
  wire _992_;
  wire _993_;
  wire _994_;
  wire _995_;
  wire _996_;
  wire _997_;
  wire _998_;
  wire _999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire _1601_;
  wire _1602_;
  wire _1603_;
  wire _1604_;
  wire _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire _1611_;
  wire _1612_;
  wire _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire _1629_;
  wire _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire _1720_;
  wire _1721_;
  wire _1722_;
  wire _1723_;
  wire _1724_;
  wire _1725_;
  wire _1726_;
  wire _1727_;
  wire _1728_;
  wire _1729_;
  wire _1730_;
  wire _1731_;
  wire _1732_;
  wire _1733_;
  wire _1734_;
  wire _1735_;
  wire _1736_;
  wire _1737_;
  wire _1738_;
  wire _1739_;
  wire _1740_;
  wire _1741_;
  wire _1742_;
  wire _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire _1751_;
  wire _1752_;
  wire _1753_;
  wire _1754_;
  wire _1755_;
  wire _1756_;
  wire _1757_;
  wire _1758_;
  wire _1759_;
  wire _1760_;
  wire _1761_;
  wire _1762_;
  wire _1763_;
  wire _1764_;
  wire _1765_;
  wire _1766_;
  wire _1767_;
  wire _1768_;
  wire _1769_;
  wire _1770_;
  wire _1771_;
  wire _1772_;
  wire _1773_;
  wire _1774_;
  wire _1775_;
  wire _1776_;
  wire _1777_;
  wire _1778_;
  wire _1779_;
  wire _1780_;
  wire _1781_;
  wire _1782_;
  wire _1783_;
  wire _1784_;
  wire _1785_;
  wire _1786_;
  wire _1787_;
  wire _1788_;
  wire _1789_;
  wire _1790_;
  wire _1791_;
  wire _1792_;
  wire _1793_;
  wire _1794_;
  wire _1795_;
  wire _1796_;
  wire _1797_;
  wire _1798_;
  wire _1799_;
  wire _1800_;
  wire _1801_;
  wire _1802_;
  wire _1803_;
  wire _1804_;
  wire _1805_;
  wire _1806_;
  wire _1807_;
  wire _1808_;
  wire _1809_;
  wire _1810_;
  wire _1811_;
  wire _1812_;
  wire _1813_;
  wire _1814_;
  wire _1815_;
  wire _1816_;
  wire _1817_;
  wire _1818_;
  wire _1819_;
  wire _1820_;
  wire _1821_;
  wire _1822_;
  wire _1823_;
  wire _1824_;
  wire _1825_;
  wire _1826_;
  wire _1827_;
  wire _1828_;
  wire _1829_;
  wire _1830_;
  wire _1831_;
  wire _1832_;
  wire _1833_;
  wire _1834_;
  wire _1835_;
  wire _1836_;
  wire _1837_;
  wire _1838_;
  wire _1839_;
  wire _1840_;
  wire _1841_;
  wire _1842_;
  wire _1843_;
  wire _1844_;
  wire _1845_;
  wire _1846_;
  wire _1847_;
  wire _1848_;
  wire _1849_;
  wire _1850_;
  wire _1851_;
  wire _1852_;
  wire _1853_;
  wire _1854_;
  wire _1855_;
  wire _1856_;
  wire _1857_;
  wire _1858_;
  wire _1859_;
  wire _1860_;
  wire _1861_;
  wire _1862_;
  wire _1863_;
  wire _1864_;
  wire _1865_;
  wire _1866_;
  wire _1867_;
  wire _1868_;
  wire _1869_;
  wire _1870_;
  wire _1871_;
  wire _1872_;
  wire _1873_;
  wire _1874_;
  wire _1875_;
  wire _1876_;
  wire _1877_;
  wire _1878_;
  wire _1879_;
  wire _1880_;
  wire _1881_;
  wire _1882_;
  wire _1883_;
  wire _1884_;
  wire _1885_;
  wire _1886_;
  wire _1887_;
  wire _1888_;
  wire _1889_;
  wire _1890_;
  wire _1891_;
  wire _1892_;
  wire _1893_;
  wire _1894_;
  wire _1895_;
  wire _1896_;
  wire _1897_;
  wire _1898_;
  wire _1899_;
  wire _1900_;
  wire _1901_;
  wire _1902_;
  wire _1903_;
  wire _1904_;
  wire _1905_;
  wire _1906_;
  wire _1907_;
  wire _1908_;
  wire _1909_;
  wire _1910_;
  wire _1911_;
  wire _1912_;
  wire _1913_;
  wire _1914_;
  wire _1915_;
  wire _1916_;
  wire _1917_;
  wire _1918_;
  wire _1919_;
  wire _1920_;
  wire _1921_;
  wire _1922_;
  wire _1923_;
  wire _1924_;
  wire _1925_;
  wire _1926_;
  wire _1927_;
  wire _1928_;
  wire _1929_;
  wire _1930_;
  wire _1931_;
  wire _1932_;
  wire _1933_;
  wire _1934_;
  wire _1935_;
  wire _1936_;
  wire _1937_;
  wire _1938_;
  wire _1939_;
  wire _1940_;
  wire _1941_;
  wire _1942_;
  wire _1943_;
  wire _1944_;
  wire _1945_;
  wire _1946_;
  wire _1947_;
  wire _1948_;
  wire _1949_;
  wire _1950_;
  wire _1951_;
  wire _1952_;
  wire _1953_;
  wire _1954_;
  wire _1955_;
  wire _1956_;
  wire _1957_;
  wire _1958_;
  wire _1959_;
  wire _1960_;
  wire _1961_;
  wire _1962_;
  wire _1963_;
  wire _1964_;
  wire _1965_;
  wire _1966_;
  wire _1967_;
  wire _1968_;
  wire _1969_;
  wire _1970_;
  wire _1971_;
  wire _1972_;
  wire _1973_;
  wire _1974_;
  wire _1975_;
  wire _1976_;
  wire _1977_;
  wire _1978_;
  wire _1979_;
  wire _1980_;
  wire _1981_;
  wire _1982_;
  wire _1983_;
  wire _1984_;
  wire _1985_;
  wire _1986_;
  wire _1987_;
  wire _1988_;
  wire _1989_;
  wire _1990_;
  wire _1991_;
  wire _1992_;
  wire _1993_;
  wire _1994_;
  wire _1995_;
  wire _1996_;
  wire _1997_;
  wire _1998_;
  wire _1999_;
  wire _2000_;
  wire _2001_;
  wire _2002_;
  wire _2003_;
  wire _2004_;
  wire _2005_;
  wire _2006_;
  wire _2007_;
  wire _2008_;
  wire _2009_;
  wire _2010_;
  wire _2011_;
  wire _2012_;
  wire _2013_;
  wire _2014_;
  wire _2015_;
  wire _2016_;
  wire _2017_;
  wire _2018_;
  wire _2019_;
  wire _2020_;
  wire _2021_;
  wire _2022_;
  wire _2023_;
  wire _2024_;
  wire _2025_;
  wire _2026_;
  wire _2027_;
  wire _2028_;
  wire _2029_;
  wire _2030_;
  wire _2031_;
  wire _2032_;
  wire _2033_;
  wire _2034_;
  wire _2035_;
  wire _2036_;
  wire _2037_;
  wire _2038_;
  wire _2039_;
  wire _2040_;
  wire _2041_;
  wire _2042_;
  wire _2043_;
  wire _2044_;
  wire _2045_;
  wire _2046_;
  wire _2047_;
  wire _2048_;
  wire _2049_;
  wire _2050_;
  wire _2051_;
  wire _2052_;
  wire _2053_;
  wire _2054_;
  wire _2055_;
  wire _2056_;
  wire _2057_;
  wire _2058_;
  wire _2059_;
  wire _2060_;
  wire _2061_;
  wire _2062_;
  wire _2063_;
  wire _2064_;
  wire _2065_;
  wire _2066_;
  wire _2067_;
  wire _2068_;
  wire _2069_;
  wire _2070_;
  wire _2071_;
  wire _2072_;
  wire _2073_;
  wire _2074_;
  wire _2075_;
  wire _2076_;
  wire _2077_;
  wire _2078_;
  wire _2079_;
  wire _2080_;
  wire _2081_;
  wire _2082_;
  wire _2083_;
  wire _2084_;
  wire _2085_;
  wire _2086_;
  wire _2087_;
  wire _2088_;
  wire _2089_;
  wire _2090_;
  wire _2091_;
  wire _2092_;
  wire _2093_;
  wire _2094_;
  wire _2095_;
  wire _2096_;
  wire _2097_;
  wire _2098_;
  wire _2099_;
  wire _2100_;
  wire _2101_;
  wire _2102_;
  wire _2103_;
  wire _2104_;
  wire _2105_;
  wire _2106_;
  wire _2107_;
  wire _2108_;
  wire _2109_;
  wire _2110_;
  wire _2111_;
  wire _2112_;
  wire _2113_;
  wire _2114_;
  wire _2115_;
  wire _2116_;
  wire _2117_;
  wire _2118_;
  wire _2119_;
  wire _2120_;
  wire _2121_;
  wire _2122_;
  wire _2123_;
  wire _2124_;
  wire _2125_;
  wire _2126_;
  wire _2127_;
  wire _2128_;
  wire _2129_;
  wire _2130_;
  wire _2131_;
  wire _2132_;
  wire _2133_;
  wire _2134_;
  wire _2135_;
  wire _2136_;
  wire _2137_;
  wire _2138_;
  wire _2139_;
  wire _2140_;
  wire _2141_;
  wire _2142_;
  wire _2143_;
  wire _2144_;
  wire _2145_;
  wire _2146_;
  wire _2147_;
  wire _2148_;
  wire _2149_;
  wire _2150_;
  wire _2151_;
  wire _2152_;
  wire _2153_;
  wire _2154_;
  wire _2155_;
  wire _2156_;
  wire _2157_;
  wire _2158_;
  wire _2159_;
  wire _2160_;
  wire _2161_;
  wire _2162_;
  wire _2163_;
  wire _2164_;
  wire _2165_;
  wire _2166_;
  wire _2167_;
  wire _2168_;
  wire _2169_;
  wire _2170_;
  wire _2171_;
  wire _2172_;
  wire _2173_;
  wire _2174_;
  wire _2175_;
  wire _2176_;
  wire _2177_;
  wire _2178_;
  wire _2179_;
  wire _2180_;
  wire _2181_;
  wire _2182_;
  wire _2183_;
  wire _2184_;
  wire _2185_;
  wire _2186_;
  wire _2187_;
  wire _2188_;
  wire _2189_;
  wire _2190_;
  wire _2191_;
  wire _2192_;
  wire _2193_;
  wire _2194_;
  wire _2195_;
  wire _2196_;
  wire _2197_;
  wire _2198_;
  wire _2199_;
  wire _2200_;
  wire _2201_;
  wire _2202_;
  wire _2203_;
  wire _2204_;
  wire _2205_;
  wire _2206_;
  wire _2207_;
  wire _2208_;
  wire _2209_;
  wire _2210_;
  wire _2211_;
  wire _2212_;
  wire _2213_;
  wire _2214_;
  wire _2215_;
  wire _2216_;
  wire _2217_;
  wire _2218_;
  wire _2219_;
  wire _2220_;
  wire _2221_;
  wire _2222_;
  wire _2223_;
  wire _2224_;
  wire _2225_;
  wire _2226_;
  wire _2227_;
  wire _2228_;
  wire _2229_;
  wire _2230_;
  wire _2231_;
  wire _2232_;
  wire _2233_;
  wire _2234_;
  wire _2235_;
  wire _2236_;
  wire _2237_;
  wire _2238_;
  wire _2239_;
  wire _2240_;
  wire _2241_;
  wire _2242_;
  wire _2243_;
  wire _2244_;
  wire _2245_;
  wire _2246_;
  wire _2247_;
  wire _2248_;
  wire _2249_;
  wire _2250_;
  wire _2251_;
  wire _2252_;
  wire _2253_;
  wire _2254_;
  wire _2255_;
  wire _2256_;
  wire _2257_;
  wire _2258_;
  wire _2259_;
  wire _2260_;
  wire _2261_;
  wire _2262_;
  wire _2263_;
  wire _2264_;
  wire _2265_;
  wire _2266_;
  wire _2267_;
  wire _2268_;
  wire _2269_;
  wire _2270_;
  wire _2271_;
  wire _2272_;
  wire _2273_;
  wire _2274_;
  wire _2275_;
  wire _2276_;
  wire _2277_;
  wire _2278_;
  wire _2279_;
  wire _2280_;
  wire _2281_;
  wire _2282_;
  wire _2283_;
  wire _2284_;
  wire _2285_;
  wire _2286_;
  wire _2287_;
  wire _2288_;
  wire _2289_;
  wire _2290_;
  wire _2291_;
  wire _2292_;
  wire _2293_;
  wire _2294_;
  wire _2295_;
  wire _2296_;
  wire _2297_;
  wire _2298_;
  wire _2299_;
  wire _2300_;
  wire _2301_;
  wire _2302_;
  wire _2303_;
  wire _2304_;
  wire _2305_;
  wire _2306_;
  wire _2307_;
  wire _2308_;
  wire _2309_;
  wire _2310_;
  wire _2311_;
  wire _2312_;
  wire _2313_;
  wire _2314_;
  wire _2315_;
  wire _2316_;
  wire _2317_;
  wire _2318_;
  wire _2319_;
  wire _2320_;
  wire _2321_;
  wire _2322_;
  wire _2323_;
  wire _2324_;
  wire _2325_;
  wire _2326_;
  wire _2327_;
  wire _2328_;
  wire _2329_;
  wire _2330_;
  wire _2331_;
  wire _2332_;
  wire _2333_;
  wire _2334_;
  wire _2335_;
  wire _2336_;
  wire _2337_;
  wire _2338_;
  wire _2339_;
  wire _2340_;
  wire _2341_;
  wire _2342_;
  wire _2343_;
  wire _2344_;
  wire _2345_;
  wire _2346_;
  wire _2347_;
  wire _2348_;
  wire _2349_;
  wire _2350_;
  wire _2351_;
  wire _2352_;
  wire _2353_;
  wire _2354_;
  wire _2355_;
  wire _2356_;
  wire _2357_;
  wire _2358_;
  wire _2359_;
  wire _2360_;
  wire _2361_;
  wire _2362_;
  wire _2363_;
  wire _2364_;
  wire _2365_;
  wire _2366_;
  wire _2367_;
  wire _2368_;
  wire _2369_;
  wire _2370_;
  wire _2371_;
  wire _2372_;
  wire _2373_;
  wire _2374_;
  wire _2375_;
  wire _2376_;
  wire _2377_;
  wire _2378_;
  wire _2379_;
  wire _2380_;
  wire _2381_;
  wire _2382_;
  wire _2383_;
  wire _2384_;
  wire _2385_;
  wire _2386_;
  wire _2387_;
  wire _2388_;
  wire _2389_;
  wire _2390_;
  wire _2391_;
  wire _2392_;
  wire _2393_;
  wire _2394_;
  wire _2395_;
  wire _2396_;
  wire _2397_;
  wire _2398_;
  wire _2399_;
  wire _2400_;
  wire _2401_;
  wire _2402_;
  wire _2403_;
  wire _2404_;
  wire _2405_;
  wire _2406_;
  wire _2407_;
  wire _2408_;
  wire _2409_;
  wire _2410_;
  wire _2411_;
  wire _2412_;
  wire _2413_;
  wire _2414_;
  wire _2415_;
  wire _2416_;
  wire _2417_;
  wire _2418_;
  wire _2419_;
  wire _2420_;
  wire _2421_;
  wire _2422_;
  wire _2423_;
  wire _2424_;
  wire _2425_;
  wire _2426_;
  wire _2427_;
  wire _2428_;
  wire _2429_;
  wire _2430_;
  wire _2431_;
  wire _2432_;
  wire _2433_;
  wire _2434_;
  wire _2435_;
  wire _2436_;
  wire _2437_;
  wire _2438_;
  wire _2439_;
  wire _2440_;
  wire _2441_;
  wire _2442_;
  wire _2443_;
  wire _2444_;
  wire _2445_;
  wire _2446_;
  wire _2447_;
  wire _2448_;
  wire _2449_;
  wire _2450_;
  wire _2451_;
  wire _2452_;
  wire _2453_;
  wire _2454_;
  wire _2455_;
  wire _2456_;
  wire _2457_;
  wire _2458_;
  wire _2459_;
  wire _2460_;
  wire _2461_;
  wire _2462_;
  wire _2463_;
  wire _2464_;
  wire _2465_;
  wire _2466_;
  wire _2467_;
  wire _2468_;
  wire _2469_;
  wire _2470_;
  wire _2471_;
  wire _2472_;
  wire _2473_;
  wire _2474_;
  wire _2475_;
  wire _2476_;
  wire _2477_;
  wire _2478_;
  wire _2479_;
  wire _2480_;
  wire _2481_;
  wire _2482_;
  wire _2483_;
  wire _2484_;
  wire _2485_;
  wire _2486_;
  wire _2487_;
  wire _2488_;
  wire _2489_;
  wire _2490_;
  wire _2491_;
  wire _2492_;
  wire _2493_;
  wire _2494_;
  wire _2495_;
  wire _2496_;
  wire _2497_;
  wire _2498_;
  wire _2499_;
  wire _2500_;
  wire _2501_;
  wire _2502_;
  wire _2503_;
  wire _2504_;
  wire _2505_;
  wire _2506_;
  wire _2507_;
  wire _2508_;
  wire _2509_;
  wire _2510_;
  wire _2511_;
  wire _2512_;
  wire _2513_;
  wire _2514_;
  wire _2515_;
  wire _2516_;
  wire _2517_;
  wire _2518_;
  wire _2519_;
  wire _2520_;
  wire _2521_;
  wire _2522_;
  wire _2523_;
  wire _2524_;
  wire _2525_;
  wire _2526_;
  wire _2527_;
  wire _2528_;
  wire _2529_;
  wire _2530_;
  wire _2531_;
  wire _2532_;
  wire _2533_;
  wire _2534_;
  wire _2535_;
  wire _2536_;
  wire _2537_;
  wire _2538_;
  wire _2539_;
  wire _2540_;
  wire _2541_;
  wire _2542_;
  wire _2543_;
  wire _2544_;
  wire _2545_;
  wire _2546_;
  wire _2547_;
  wire _2548_;
  wire _2549_;
  wire _2550_;
  wire _2551_;
  wire _2552_;
  wire _2553_;
  wire _2554_;
  wire _2555_;
  wire _2556_;
  wire _2557_;
  wire _2558_;
  wire _2559_;
  wire _2560_;
  wire _2561_;
  wire _2562_;
  wire _2563_;
  wire _2564_;
  wire _2565_;
  wire _2566_;
  wire _2567_;
  wire _2568_;
  wire _2569_;
  wire _2570_;
  wire _2571_;
  wire _2572_;
  wire _2573_;
  wire _2574_;
  wire _2575_;
  wire _2576_;
  wire _2577_;
  wire _2578_;
  wire _2579_;
  wire _2580_;
  wire _2581_;
  wire _2582_;
  wire _2583_;
  wire _2584_;
  wire _2585_;
  wire _2586_;
  wire _2587_;
  wire _2588_;
  wire _2589_;
  wire _2590_;
  wire _2591_;
  wire _2592_;
  wire _2593_;
  wire _2594_;
  wire _2595_;
  wire _2596_;
  wire _2597_;
  wire _2598_;
  wire _2599_;
  wire _2600_;
  wire _2601_;
  wire _2602_;
  wire _2603_;
  wire _2604_;
  wire _2605_;
  wire _2606_;
  wire _2607_;
  wire _2608_;
  wire _2609_;
  wire _2610_;
  wire _2611_;
  wire _2612_;
  wire _2613_;
  wire _2614_;
  wire _2615_;
  wire _2616_;
  wire _2617_;
  wire _2618_;
  wire _2619_;
  wire _2620_;
  wire _2621_;
  wire _2622_;
  wire _2623_;
  wire _2624_;
  wire _2625_;
  wire _2626_;
  wire _2627_;
  wire _2628_;
  wire _2629_;
  wire _2630_;
  wire _2631_;
  wire _2632_;
  wire _2633_;
  wire _2634_;
  wire _2635_;
  wire _2636_;
  wire _2637_;
  wire _2638_;
  wire _2639_;
  wire _2640_;
  wire _2641_;
  wire _2642_;
  wire _2643_;
  wire _2644_;
  wire _2645_;
  wire _2646_;
  wire _2647_;
  wire _2648_;
  wire _2649_;
  wire _2650_;
  wire _2651_;
  wire _2652_;
  wire _2653_;
  wire _2654_;
  wire _2655_;
  wire _2656_;
  wire _2657_;
  wire _2658_;
  wire _2659_;
  wire _2660_;
  wire _2661_;
  wire _2662_;
  wire _2663_;
  wire _2664_;
  wire _2665_;
  wire _2666_;
  wire _2667_;
  wire _2668_;
  wire _2669_;
  wire _2670_;
  wire _2671_;
  wire _2672_;
  wire _2673_;
  wire _2674_;
  wire _2675_;
  wire _2676_;
  wire _2677_;
  wire _2678_;
  wire _2679_;
  wire _2680_;
  wire _2681_;
  wire _2682_;
  wire _2683_;
  wire _2684_;
  wire _2685_;
  wire _2686_;
  wire _2687_;
  wire _2688_;
  wire _2689_;
  wire _2690_;
  wire _2691_;
  wire _2692_;
  wire _2693_;
  wire _2694_;
  wire _2695_;
  wire _2696_;
  wire _2697_;
  wire _2698_;
  wire _2699_;
  wire _2700_;
  wire _2701_;
  wire _2702_;
  wire _2703_;
  wire _2704_;
  wire _2705_;
  wire _2706_;
  wire _2707_;
  wire _2708_;
  wire _2709_;
  wire _2710_;
  wire _2711_;
  wire _2712_;
  wire _2713_;
  wire _2714_;
  wire _2715_;
  wire _2716_;
  wire _2717_;
  wire _2718_;
  wire _2719_;
  wire _2720_;
  wire _2721_;
  wire _2722_;
  wire _2723_;
  wire _2724_;
  wire _2725_;
  wire _2726_;
  wire _2727_;
  wire _2728_;
  wire _2729_;
  wire _2730_;
  wire _2731_;
  wire _2732_;
  wire _2733_;
  wire _2734_;
  wire _2735_;
  wire _2736_;
  wire _2737_;
  wire _2738_;
  wire _2739_;
  wire _2740_;
  wire _2741_;
  wire _2742_;
  wire _2743_;
  wire _2744_;
  wire _2745_;
  wire _2746_;
  wire _2747_;
  wire _2748_;
  wire _2749_;
  wire _2750_;
  wire _2751_;
  wire _2752_;
  wire _2753_;
  wire _2754_;
  wire _2755_;
  wire _2756_;
  wire _2757_;
  wire _2758_;
  wire _2759_;
  wire _2760_;
  wire _2761_;
  wire _2762_;
  wire _2763_;
  wire _2764_;
  wire _2765_;
  wire _2766_;
  wire _2767_;
  wire _2768_;
  wire _2769_;
  wire _2770_;
  wire _2771_;
  wire _2772_;
  wire _2773_;
  wire _2774_;
  wire _2775_;
  wire _2776_;
  wire _2777_;
  wire _2778_;
  wire _2779_;
  wire _2780_;
  wire _2781_;
  wire _2782_;
  wire _2783_;
  wire _2784_;
  wire _2785_;
  wire _2786_;
  wire _2787_;
  wire _2788_;
  wire _2789_;
  wire _2790_;
  wire _2791_;
  wire _2792_;
  wire _2793_;
  wire _2794_;
  wire _2795_;
  wire _2796_;
  wire _2797_;
  wire _2798_;
  wire _2799_;
  wire _2800_;
  wire _2801_;
  wire _2802_;
  wire _2803_;
  wire _2804_;
  wire _2805_;
  wire _2806_;
  wire _2807_;
  wire _2808_;
  wire _2809_;
  wire _2810_;
  wire _2811_;
  wire _2812_;
  wire _2813_;
  wire _2814_;
  wire _2815_;
  wire _2816_;
  wire _2817_;
  wire _2818_;
  wire _2819_;
  wire _2820_;
  wire _2821_;
  wire _2822_;
  wire _2823_;
  wire _2824_;
  wire _2825_;
  wire _2826_;
  wire _2827_;
  wire _2828_;
  wire _2829_;
  wire _2830_;
  wire _2831_;
  wire _2832_;
  wire _2833_;
  wire _2834_;
  wire _2835_;
  wire _2836_;
  wire _2837_;
  wire _2838_;
  wire _2839_;
  wire _2840_;
  wire _2841_;
  wire _2842_;
  wire _2843_;
  wire _2844_;
  wire _2845_;
  wire _2846_;
  wire _2847_;
  wire _2848_;
  wire _2849_;
  wire _2850_;
  wire _2851_;
  wire _2852_;
  wire _2853_;
  wire _2854_;
  wire _2855_;
  wire _2856_;
  wire _2857_;
  wire _2858_;
  wire _2859_;
  wire _2860_;
  wire _2861_;
  wire _2862_;
  wire _2863_;
  wire _2864_;
  wire _2865_;
  wire _2866_;
  wire _2867_;
  wire _2868_;
  wire _2869_;
  wire _2870_;
  wire _2871_;
  wire _2872_;
  wire _2873_;
  wire _2874_;
  wire _2875_;
  wire _2876_;
  wire _2877_;
  wire _2878_;
  wire _2879_;
  wire _2880_;
  wire _2881_;
  wire _2882_;
  wire _2883_;
  wire _2884_;
  wire _2885_;
  wire _2886_;
  wire _2887_;
  wire _2888_;
  wire _2889_;
  wire _2890_;
  wire _2891_;
  wire _2892_;
  wire _2893_;
  wire _2894_;
  wire _2895_;
  wire _2896_;
  wire _2897_;
  wire _2898_;
  wire _2899_;
  wire _2900_;
  wire _2901_;
  wire _2902_;
  wire _2903_;
  wire _2904_;
  wire _2905_;
  wire _2906_;
  wire _2907_;
  wire _2908_;
  wire _2909_;
  wire _2910_;
  wire _2911_;
  wire _2912_;
  wire _2913_;
  wire _2914_;
  wire _2915_;
  wire _2916_;
  wire _2917_;
  wire _2918_;
  wire _2919_;
  wire _2920_;
  wire _2921_;
  wire _2922_;
  wire _2923_;
  wire _2924_;
  wire _2925_;
  wire _2926_;
  wire _2927_;
  wire _2928_;
  wire _2929_;
  wire _2930_;
  wire _2931_;
  wire _2932_;
  wire _2933_;
  wire _2934_;
  wire _2935_;
  wire _2936_;
  wire _2937_;
  wire _2938_;
  wire _2939_;
  wire _2940_;
  wire _2941_;
  wire _2942_;
  wire _2943_;
  wire _2944_;
  wire _2945_;
  wire _2946_;
  wire _2947_;
  wire _2948_;
  wire _2949_;
  wire _2950_;
  wire _2951_;
  wire _2952_;
  wire _2953_;
  wire _2954_;
  wire _2955_;
  wire _2956_;
  wire _2957_;
  wire _2958_;
  wire _2959_;
  wire _2960_;
  wire _2961_;
  wire _2962_;
  wire _2963_;
  wire _2964_;
  wire _2965_;
  wire _2966_;
  wire _2967_;
  wire _2968_;
  wire _2969_;
  wire _2970_;
  wire _2971_;
  wire _2972_;
  wire _2973_;
  wire _2974_;
  wire _2975_;
  wire _2976_;
  wire _2977_;
  wire _2978_;
  wire _2979_;
  wire _2980_;
  wire _2981_;
  wire _2982_;
  wire _2983_;
  wire _2984_;
  wire _2985_;
  wire _2986_;
  wire _2987_;
  wire _2988_;
  wire _2989_;
  wire _2990_;
  wire _2991_;
  wire _2992_;
  wire _2993_;
  wire _2994_;
  wire _2995_;
  wire _2996_;
  wire _2997_;
  wire _2998_;
  wire _2999_;
  wire _3000_;
  wire _3001_;
  wire _3002_;
  wire _3003_;
  wire _3004_;
  wire _3005_;
  wire _3006_;
  wire _3007_;
  wire _3008_;
  wire _3009_;
  wire _3010_;
  wire _3011_;
  wire _3012_;
  wire _3013_;
  wire _3014_;
  wire _3015_;
  wire _3016_;
  wire _3017_;
  wire _3018_;
  wire _3019_;
  wire _3020_;
  wire _3021_;
  wire _3022_;
  wire _3023_;
  wire _3024_;
  wire _3025_;
  wire _3026_;
  wire _3027_;
  wire _3028_;
  wire _3029_;
  wire _3030_;
  wire _3031_;
  wire _3032_;
  wire _3033_;
  wire _3034_;
  wire _3035_;
  wire _3036_;
  wire _3037_;
  wire _3038_;
  wire _3039_;
  wire _3040_;
  wire _3041_;
  wire _3042_;
  wire _3043_;
  wire _3044_;
  wire _3045_;
  wire _3046_;
  wire _3047_;
  wire _3048_;
  wire _3049_;
  wire _3050_;
  wire _3051_;
  wire _3052_;
  wire _3053_;
  wire _3054_;
  wire _3055_;
  wire _3056_;
  wire _3057_;
  wire _3058_;
  wire _3059_;
  wire _3060_;
  wire _3061_;
  wire _3062_;
  wire _3063_;
  wire _3064_;
  wire _3065_;
  wire _3066_;
  wire _3067_;
  wire _3068_;
  wire _3069_;
  wire _3070_;
  wire _3071_;
  wire _3072_;
  wire _3073_;
  wire _3074_;
  wire _3075_;
  wire _3076_;
  wire _3077_;
  wire _3078_;
  wire _3079_;
  wire _3080_;
  wire _3081_;
  wire _3082_;
  wire _3083_;
  wire _3084_;
  wire _3085_;
  wire _3086_;
  wire _3087_;
  wire _3088_;
  wire _3089_;
  wire _3090_;
  wire _3091_;
  wire _3092_;
  wire _3093_;
  wire _3094_;
  wire _3095_;
  wire _3096_;
  wire _3097_;
  wire _3098_;
  wire _3099_;
  wire _3100_;
  wire _3101_;
  wire _3102_;
  wire _3103_;
  wire _3104_;
  wire _3105_;
  wire _3106_;
  wire _3107_;
  wire _3108_;
  wire _3109_;
  wire _3110_;
  wire _3111_;
  wire _3112_;
  wire _3113_;
  wire _3114_;
  wire _3115_;
  wire _3116_;
  wire _3117_;
  wire _3118_;
  wire _3119_;
  wire _3120_;
  wire _3121_;
  wire _3122_;
  wire _3123_;
  wire _3124_;
  wire _3125_;
  wire _3126_;
  wire _3127_;
  wire _3128_;
  wire _3129_;
  wire _3130_;
  wire _3131_;
  wire _3132_;
  wire _3133_;
  wire _3134_;
  wire _3135_;
  wire _3136_;
  wire _3137_;
  wire _3138_;
  wire _3139_;
  wire _3140_;
  wire _3141_;
  wire _3142_;
  wire _3143_;
  wire _3144_;
  wire _3145_;
  wire _3146_;
  wire _3147_;
  wire _3148_;
  wire _3149_;
  wire _3150_;
  wire _3151_;
  wire _3152_;
  wire _3153_;
  wire _3154_;
  wire _3155_;
  wire _3156_;
  wire _3157_;
  wire _3158_;
  wire _3159_;
  wire _3160_;
  wire _3161_;
  wire _3162_;
  wire _3163_;
  wire _3164_;
  wire _3165_;
  wire _3166_;
  wire _3167_;
  wire _3168_;
  wire _3169_;
  wire _3170_;
  wire _3171_;
  wire _3172_;
  wire _3173_;
  wire _3174_;
  wire _3175_;
  wire _3176_;
  wire _3177_;
  wire _3178_;
  wire _3179_;
  wire _3180_;
  wire _3181_;
  wire _3182_;
  wire _3183_;
  wire _3184_;
  wire _3185_;
  wire _3186_;
  wire _3187_;
  wire _3188_;
  wire _3189_;
  wire _3190_;
  wire _3191_;
  wire _3192_;
  wire _3193_;
  wire _3194_;
  wire _3195_;
  wire _3196_;
  wire _3197_;
  wire _3198_;
  wire _3199_;
  wire _3200_;
  wire _3201_;
  wire _3202_;
  wire _3203_;
  wire _3204_;
  wire _3205_;
  wire _3206_;
  wire _3207_;
  wire _3208_;
  wire _3209_;
  wire _3210_;
  wire _3211_;
  wire _3212_;
  wire _3213_;
  wire _3214_;
  wire _3215_;
  wire _3216_;
  wire _3217_;
  wire _3218_;
  wire _3219_;
  wire _3220_;
  wire _3221_;
  wire _3222_;
  wire _3223_;
  wire _3224_;
  wire _3225_;
  wire _3226_;
  wire _3227_;
  wire _3228_;
  wire _3229_;
  wire _3230_;
  wire _3231_;
  wire _3232_;
  wire _3233_;
  wire _3234_;
  wire _3235_;
  wire _3236_;
  wire _3237_;
  wire _3238_;
  wire _3239_;
  wire _3240_;
  wire _3241_;
  wire _3242_;
  wire _3243_;
  wire _3244_;
  wire _3245_;
  wire _3246_;
  wire _3247_;
  wire _3248_;
  wire _3249_;
  wire _3250_;
  wire _3251_;
  wire _3252_;
  wire _3253_;
  wire _3254_;
  wire _3255_;
  wire _3256_;
  wire _3257_;
  wire _3258_;
  wire _3259_;
  wire _3260_;
  wire _3261_;
  wire _3262_;
  wire _3263_;
  wire _3264_;
  wire _3265_;
  wire _3266_;
  wire _3267_;
  wire _3268_;
  wire _3269_;
  wire _3270_;
  wire _3271_;
  wire _3272_;
  wire _3273_;
  wire _3274_;
  wire _3275_;
  wire _3276_;
  wire _3277_;
  wire _3278_;
  wire _3279_;
  wire _3280_;
  wire _3281_;
  wire _3282_;
  wire _3283_;
  wire _3284_;
  wire _3285_;
  wire _3286_;
  wire _3287_;
  wire _3288_;
  wire _3289_;
  wire _3290_;
  wire _3291_;
  wire _3292_;
  wire _3293_;
  wire _3294_;
  wire _3295_;
  wire _3296_;
  wire _3297_;
  wire _3298_;
  wire _3299_;
  wire _3300_;
  wire _3301_;
  wire _3302_;
  wire _3303_;
  wire _3304_;
  wire _3305_;
  wire _3306_;
  wire _3307_;
  wire _3308_;
  wire _3309_;
  wire _3310_;
  wire _3311_;
  wire _3312_;
  wire _3313_;
  wire _3314_;
  wire _3315_;
  wire _3316_;
  wire _3317_;
  wire _3318_;
  wire _3319_;
  wire _3320_;
  wire _3321_;
  wire _3322_;
  wire _3323_;
  wire _3324_;
  wire _3325_;
  wire _3326_;
  wire _3327_;
  wire _3328_;
  wire _3329_;
  wire _3330_;
  wire _3331_;
  wire _3332_;
  wire _3333_;
  wire _3334_;
  wire _3335_;
  wire _3336_;
  wire _3337_;
  wire _3338_;
  wire _3339_;
  wire _3340_;
  wire _3341_;
  wire _3342_;
  wire _3343_;
  wire _3344_;
  wire _3345_;
  wire _3346_;
  wire _3347_;
  wire _3348_;
  wire _3349_;
  wire _3350_;
  wire _3351_;
  wire _3352_;
  wire _3353_;
  wire _3354_;
  wire _3355_;
  wire _3356_;
  wire _3357_;
  wire _3358_;
  wire _3359_;
  wire _3360_;
  wire _3361_;
  wire _3362_;
  wire _3363_;
  wire _3364_;
  wire _3365_;
  wire _3366_;
  wire _3367_;
  wire _3368_;
  wire _3369_;
  wire _3370_;
  wire _3371_;
  wire _3372_;
  wire _3373_;
  wire _3374_;
  wire _3375_;
  wire _3376_;
  wire _3377_;
  wire _3378_;
  wire _3379_;
  wire _3380_;
  wire _3381_;
  wire _3382_;
  wire _3383_;
  wire _3384_;
  wire _3385_;
  wire _3386_;
  wire _3387_;
  wire _3388_;
  wire _3389_;
  wire _3390_;
  wire _3391_;
  wire _3392_;
  wire _3393_;
  wire _3394_;
  wire _3395_;
  wire _3396_;
  wire _3397_;
  wire _3398_;
  wire _3399_;
  wire _3400_;
  wire _3401_;
  wire _3402_;
  wire _3403_;
  wire _3404_;
  wire _3405_;
  wire _3406_;
  wire _3407_;
  wire _3408_;
  wire _3409_;
  wire _3410_;
  wire _3411_;
  wire _3412_;
  wire _3413_;
  wire _3414_;
  wire _3415_;
  wire _3416_;
  wire _3417_;
  wire _3418_;
  wire _3419_;
  wire _3420_;
  wire _3421_;
  wire _3422_;
  wire _3423_;
  wire _3424_;
  wire _3425_;
  wire _3426_;
  wire _3427_;
  wire _3428_;
  wire _3429_;
  wire _3430_;
  wire _3431_;
  wire _3432_;
  wire _3433_;
  wire _3434_;
  wire _3435_;
  wire _3436_;
  wire _3437_;
  wire _3438_;
  wire _3439_;
  wire _3440_;
  wire _3441_;
  wire _3442_;
  wire _3443_;
  wire _3444_;
  wire _3445_;
  wire _3446_;
  wire _3447_;
  wire _3448_;
  wire _3449_;
  wire _3450_;
  wire _3451_;
  wire _3452_;
  wire _3453_;
  wire _3454_;
  wire _3455_;
  wire _3456_;
  wire _3457_;
  wire _3458_;
  wire _3459_;
  wire _3460_;
  wire _3461_;
  wire _3462_;
  wire _3463_;
  wire _3464_;
  wire _3465_;
  wire _3466_;
  wire _3467_;
  wire _3468_;
  wire _3469_;
  wire _3470_;
  wire _3471_;
  wire _3472_;
  wire _3473_;
  wire _3474_;
  wire _3475_;
  wire _3476_;
  wire _3477_;
  wire _3478_;
  wire _3479_;
  wire _3480_;
  wire _3481_;
  wire _3482_;
  wire _3483_;
  wire _3484_;
  wire _3485_;
  wire _3486_;
  wire _3487_;
  wire _3488_;
  wire _3489_;
  wire _3490_;
  wire _3491_;
  wire _3492_;
  wire _3493_;
  wire _3494_;
  wire _3495_;
  wire _3496_;
  wire _3497_;
  wire _3498_;
  wire _3499_;
  wire _3500_;
  wire _3501_;
  wire _3502_;
  wire _3503_;
  wire _3504_;
  wire _3505_;
  wire _3506_;
  wire _3507_;
  wire _3508_;
  wire _3509_;
  wire _3510_;
  wire _3511_;
  wire _3512_;
  wire _3513_;
  wire _3514_;
  wire _3515_;
  wire _3516_;
  wire _3517_;
  wire _3518_;
  wire _3519_;
  wire _3520_;
  wire _3521_;
  wire _3522_;
  wire _3523_;
  wire _3524_;
  wire _3525_;
  wire _3526_;
  wire _3527_;
  wire _3528_;
  wire _3529_;
  wire _3530_;
  wire _3531_;
  wire _3532_;
  wire _3533_;
  wire _3534_;
  wire _3535_;
  wire _3536_;
  wire _3537_;
  wire _3538_;
  wire _3539_;
  wire _3540_;
  wire _3541_;
  wire _3542_;
  wire _3543_;
  wire _3544_;
  wire _3545_;
  wire _3546_;
  wire _3547_;
  wire _3548_;
  wire _3549_;
  wire _3550_;
  wire _3551_;
  wire _3552_;
  wire _3553_;
  wire _3554_;
  wire _3555_;
  wire _3556_;
  wire _3557_;
  wire _3558_;
  wire _3559_;
  wire _3560_;
  wire _3561_;
  wire _3562_;
  wire _3563_;
  wire _3564_;
  wire _3565_;
  wire _3566_;
  wire _3567_;
  wire _3568_;
  wire _3569_;
  wire _3570_;
  wire _3571_;
  wire _3572_;
  wire _3573_;
  wire _3574_;
  wire _3575_;
  wire _3576_;
  wire _3577_;
  wire _3578_;
  wire _3579_;
  wire _3580_;
  wire _3581_;
  wire _3582_;
  wire _3583_;
  wire _3584_;
  wire _3585_;
  wire _3586_;
  wire _3587_;
  wire _3588_;
  wire _3589_;
  wire _3590_;
  wire _3591_;
  wire _3592_;
  wire _3593_;
  wire _3594_;
  wire _3595_;
  wire _3596_;
  wire _3597_;
  wire _3598_;
  wire _3599_;
  wire _3600_;
  wire _3601_;
  wire _3602_;
  wire _3603_;
  wire _3604_;
  wire _3605_;
  wire _3606_;
  wire _3607_;
  wire _3608_;
  wire _3609_;
  wire _3610_;
  wire _3611_;
  wire _3612_;
  wire _3613_;
  wire _3614_;
  wire _3615_;
  wire _3616_;
  wire _3617_;
  wire _3618_;
  wire _3619_;
  wire _3620_;
  wire _3621_;
  wire _3622_;
  wire _3623_;
  wire _3624_;
  wire _3625_;
  wire _3626_;
  wire _3627_;
  wire _3628_;
  wire _3629_;
  wire _3630_;
  wire _3631_;
  wire _3632_;
  wire _3633_;
  wire _3634_;
  wire _3635_;
  wire _3636_;
  wire _3637_;
  wire _3638_;
  wire _3639_;
  wire _3640_;
  wire _3641_;
  wire _3642_;
  wire _3643_;
  wire _3644_;
  wire _3645_;
  wire _3646_;
  wire _3647_;
  wire _3648_;
  wire _3649_;
  wire _3650_;
  wire _3651_;
  wire _3652_;
  wire _3653_;
  wire _3654_;
  wire _3655_;
  wire _3656_;
  wire _3657_;
  wire _3658_;
  wire _3659_;
  wire _3660_;
  wire _3661_;
  wire _3662_;
  wire _3663_;
  wire _3664_;
  wire _3665_;
  wire _3666_;
  wire _3667_;
  wire _3668_;
  wire _3669_;
  wire _3670_;
  wire _3671_;
  wire _3672_;
  wire _3673_;
  wire _3674_;
  wire _3675_;
  wire _3676_;
  wire _3677_;
  wire _3678_;
  wire _3679_;
  wire _3680_;
  wire _3681_;
  wire _3682_;
  wire _3683_;
  wire _3684_;
  wire _3685_;
  wire _3686_;
  wire _3687_;
  wire _3688_;
  wire _3689_;
  wire _3690_;
  wire _3691_;
  wire _3692_;
  wire _3693_;
  wire _3694_;
  wire _3695_;
  wire _3696_;
  wire _3697_;
  wire _3698_;
  wire _3699_;
  wire _3700_;
  wire _3701_;
  wire _3702_;
  wire _3703_;
  wire _3704_;
  wire _3705_;
  wire _3706_;
  wire _3707_;
  wire _3708_;
  wire _3709_;
  wire _3710_;
  wire _3711_;
  wire _3712_;
  wire _3713_;
  wire _3714_;
  wire _3715_;
  wire _3716_;
  wire _3717_;
  wire _3718_;
  wire _3719_;
  wire _3720_;
  wire _3721_;
  wire _3722_;
  wire _3723_;
  wire _3724_;
  wire _3725_;
  wire _3726_;
  wire _3727_;
  wire _3728_;
  wire _3729_;
  wire _3730_;
  wire _3731_;
  wire _3732_;
  wire _3733_;
  wire _3734_;
  wire _3735_;
  wire _3736_;
  wire _3737_;
  wire _3738_;
  wire _3739_;
  wire _3740_;
  wire _3741_;
  wire _3742_;
  wire _3743_;
  wire _3744_;
  wire _3745_;
  wire _3746_;
  wire _3747_;
  wire _3748_;
  wire _3749_;
  wire _3750_;
  wire _3751_;
  wire _3752_;
  wire _3753_;
  wire _3754_;
  wire _3755_;
  wire _3756_;
  wire _3757_;
  wire _3758_;
  wire _3759_;
  wire _3760_;
  wire _3761_;
  wire _3762_;
  wire _3763_;
  wire _3764_;
  wire _3765_;
  wire _3766_;
  wire _3767_;
  wire _3768_;
  wire _3769_;
  wire _3770_;
  wire _3771_;
  wire _3772_;
  wire _3773_;
  wire _3774_;
  wire _3775_;
  wire _3776_;
  wire _3777_;
  wire _3778_;
  wire _3779_;
  wire _3780_;
  wire _3781_;
  wire _3782_;
  wire _3783_;
  wire _3784_;
  wire _3785_;
  wire _3786_;
  wire _3787_;
  wire _3788_;
  wire _3789_;
  wire _3790_;
  wire _3791_;
  wire _3792_;
  wire _3793_;
  wire _3794_;
  wire _3795_;
  wire _3796_;
  wire _3797_;
  wire _3798_;
  wire _3799_;
  wire _3800_;
  wire _3801_;
  wire _3802_;
  wire _3803_;
  wire _3804_;
  wire _3805_;
  wire _3806_;
  wire _3807_;
  wire _3808_;
  wire _3809_;
  wire _3810_;
  wire _3811_;
  wire _3812_;
  wire _3813_;
  wire _3814_;
  wire _3815_;
  wire _3816_;
  wire _3817_;
  wire _3818_;
  wire _3819_;
  wire _3820_;
  wire _3821_;
  wire _3822_;
  wire _3823_;
  wire _3824_;
  wire _3825_;
  wire _3826_;
  wire _3827_;
  wire _3828_;
  wire _3829_;
  wire _3830_;
  wire _3831_;
  wire _3832_;
  wire _3833_;
  wire _3834_;
  wire _3835_;
  wire _3836_;
  wire _3837_;
  wire _3838_;
  wire _3839_;
  wire _3840_;
  wire _3841_;
  wire _3842_;
  wire _3843_;
  wire _3844_;
  wire _3845_;
  wire _3846_;
  wire _3847_;
  wire _3848_;
  wire _3849_;
  wire _3850_;
  wire _3851_;
  wire _3852_;
  wire _3853_;
  wire _3854_;
  wire _3855_;
  wire _3856_;
  wire _3857_;
  wire _3858_;
  wire _3859_;
  wire _3860_;
  wire _3861_;
  wire _3862_;
  wire _3863_;
  wire _3864_;
  wire _3865_;
  wire _3866_;
  wire _3867_;
  wire _3868_;
  wire _3869_;
  wire _3870_;
  wire _3871_;
  wire _3872_;
  wire _3873_;
  wire _3874_;
  wire _3875_;
  wire _3876_;
  wire _3877_;
  wire _3878_;
  wire _3879_;
  wire _3880_;
  wire _3881_;
  wire _3882_;
  wire _3883_;
  wire _3884_;
  wire _3885_;
  wire _3886_;
  wire _3887_;
  wire _3888_;
  wire _3889_;
  wire _3890_;
  wire _3891_;
  wire _3892_;
  wire _3893_;
  wire _3894_;
  wire _3895_;
  wire _3896_;
  wire _3897_;
  wire _3898_;
  wire _3899_;
  wire _3900_;
  wire _3901_;
  wire _3902_;
  wire _3903_;
  wire _3904_;
  wire _3905_;
  wire _3906_;
  wire _3907_;
  wire _3908_;
  wire _3909_;
  wire _3910_;
  wire _3911_;
  wire _3912_;
  wire _3913_;
  wire _3914_;
  wire _3915_;
  wire _3916_;
  wire _3917_;
  wire _3918_;
  wire _3919_;
  wire _3920_;
  wire _3921_;
  wire _3922_;
  wire _3923_;
  wire _3924_;
  wire _3925_;
  wire _3926_;
  wire _3927_;
  wire _3928_;
  wire _3929_;
  wire _3930_;
  wire _3931_;
  wire _3932_;
  wire _3933_;
  wire _3934_;
  wire _3935_;
  wire _3936_;
  wire _3937_;
  wire _3938_;
  wire _3939_;
  wire _3940_;
  wire _3941_;
  wire _3942_;
  wire _3943_;
  wire _3944_;
  wire _3945_;
  wire _3946_;
  wire _3947_;
  wire _3948_;
  wire _3949_;
  wire _3950_;
  wire _3951_;
  wire _3952_;
  wire _3953_;
  wire _3954_;
  wire _3955_;
  wire _3956_;
  wire _3957_;
  wire _3958_;
  wire _3959_;
  wire _3960_;
  wire _3961_;
  wire _3962_;
  wire _3963_;
  wire _3964_;
  wire _3965_;
  wire _3966_;
  wire _3967_;
  wire _3968_;
  wire _3969_;
  wire _3970_;
  wire _3971_;
  wire _3972_;
  wire _3973_;
  wire _3974_;
  wire _3975_;
  wire _3976_;
  wire _3977_;
  wire _3978_;
  wire _3979_;
  wire _3980_;
  wire _3981_;
  wire _3982_;
  wire _3983_;
  wire _3984_;
  wire _3985_;
  wire _3986_;
  wire _3987_;
  wire _3988_;
  wire _3989_;
  wire _3990_;
  wire _3991_;
  wire _3992_;
  wire _3993_;
  wire _3994_;
  wire _3995_;
  wire _3996_;
  wire _3997_;
  wire _3998_;
  wire _3999_;
  wire _4000_;
  wire _4001_;
  wire _4002_;
  wire _4003_;
  wire _4004_;
  wire _4005_;
  wire _4006_;
  wire _4007_;
  wire _4008_;
  wire _4009_;
  wire _4010_;
  wire _4011_;
  wire _4012_;
  wire _4013_;
  wire _4014_;
  wire _4015_;
  wire _4016_;
  wire _4017_;
  wire _4018_;
  wire _4019_;
  wire _4020_;
  wire _4021_;
  wire _4022_;
  wire _4023_;
  wire _4024_;
  wire _4025_;
  wire _4026_;
  wire _4027_;
  wire _4028_;
  wire _4029_;
  wire _4030_;
  wire _4031_;
  wire [46:0] r_0;
  wire [46:0] r_1;
  wire [23:0] m_1;
  wire [23:0] sum_1;
  wire [23:0] inv_1;
  wire [45:0] r_2;
  wire [23:0] m_2;
  wire [23:0] sum_2;
  wire [23:0] inv_2;
  wire [44:0] r_3;
  wire [23:0] m_3;
  wire [23:0] sum_3;
  wire [23:0] inv_3;
  wire [43:0] r_4;
  wire [23:0] m_4;
  wire [23:0] sum_4;
  wire [23:0] inv_4;
  wire [42:0] r_5;
  wire [23:0] m_5;
  wire [23:0] sum_5;
  wire [23:0] inv_5;
  wire [41:0] r_6;
  wire [23:0] m_6;
  wire [23:0] sum_6;
  wire [23:0] inv_6;
  wire [40:0] r_7;
  wire [23:0] m_7;
  wire [23:0] sum_7;
  wire [23:0] inv_7;
  wire [39:0] r_8;
  wire [23:0] m_8;
  wire [23:0] sum_8;
  wire [23:0] inv_8;
  wire [38:0] r_9;
  wire [23:0] m_9;
  wire [23:0] sum_9;
  wire [23:0] inv_9;
  wire [37:0] r_10;
  wire [23:0] m_10;
  wire [23:0] sum_10;
  wire [23:0] inv_10;
  wire [36:0] r_11;
  wire [23:0] m_11;
  wire [23:0] sum_11;
  wire [23:0] inv_11;
  wire [35:0] r_12;
  wire [23:0] m_12;
  wire [23:0] sum_12;
  wire [23:0] inv_12;
  wire [34:0] r_13;
  wire [23:0] m_13;
  wire [23:0] sum_13;
  wire [23:0] inv_13;
  wire [33:0] r_14;
  wire [23:0] m_14;
  wire [23:0] sum_14;
  wire [23:0] inv_14;
  wire [32:0] r_15;
  wire [23:0] m_15;
  wire [23:0] sum_15;
  wire [23:0] inv_15;
  wire [31:0] r_16;
  wire [23:0] m_16;
  wire [23:0] sum_16;
  wire [23:0] inv_16;
  wire [30:0] r_17;
  wire [23:0] m_17;
  wire [23:0] sum_17;
  wire [23:0] inv_17;
  wire [29:0] r_18;
  wire [23:0] m_18;
  wire [23:0] sum_18;
  wire [23:0] inv_18;
  wire [28:0] r_19;
  wire [23:0] m_19;
  wire [23:0] sum_19;
  wire [23:0] inv_19;
  wire [27:0] r_20;
  wire [23:0] m_20;
  wire [23:0] sum_20;
  wire [23:0] inv_20;
  wire [26:0] r_21;
  wire [23:0] m_21;
  wire [23:0] sum_21;
  wire [23:0] inv_21;
  wire [25:0] r_22;
  wire [23:0] m_22;
  wire [23:0] sum_22;
  wire [23:0] inv_22;
  wire [24:0] r_23;
  wire [23:0] m_23;
  wire [23:0] sum_23;
  wire [23:0] inv_23;
  wire [23:0] r_24;
  wire [23:0] m_24;
  wire [23:0] sum_24;
  wire [23:0] inv_24;
  wire zeroWire;
  wire oneWire;
  input [45:0] rin;
  input [22:0] div;
  output [23:0] q;
  output [23:0] rout;
  assign zeroWire = 1'b0 /*0*/;
  assign oneWire = 1'b1 /*0*/;
  assign r_0[0] = rin[0] /*19007*/;
  assign r_0[1] = rin[1] /*19006*/;
  assign r_0[2] = rin[2] /*19005*/;
  assign r_0[3] = rin[3] /*19004*/;
  assign r_0[4] = rin[4] /*19003*/;
  assign r_0[5] = rin[5] /*19002*/;
  assign r_0[6] = rin[6] /*19001*/;
  assign r_0[7] = rin[7] /*19000*/;
  assign r_0[8] = rin[8] /*18999*/;
  assign r_0[9] = rin[9] /*18998*/;
  assign r_0[10] = rin[10] /*18997*/;
  assign r_0[11] = rin[11] /*18996*/;
  assign r_0[12] = rin[12] /*18995*/;
  assign r_0[13] = rin[13] /*18994*/;
  assign r_0[14] = rin[14] /*18993*/;
  assign r_0[15] = rin[15] /*18992*/;
  assign r_0[16] = rin[16] /*18991*/;
  assign r_0[17] = rin[17] /*18990*/;
  assign r_0[18] = rin[18] /*18989*/;
  assign r_0[19] = rin[19] /*18988*/;
  assign r_0[20] = rin[20] /*18987*/;
  assign r_0[21] = rin[21] /*18986*/;
  assign r_0[22] = rin[22] /*18985*/;
  assign r_0[23] = rin[23] /*18984*/;
  assign r_0[24] = rin[24] /*18983*/;
  assign r_0[25] = rin[25] /*18982*/;
  assign r_0[26] = rin[26] /*18981*/;
  assign r_0[27] = rin[27] /*18980*/;
  assign r_0[28] = rin[28] /*18979*/;
  assign r_0[29] = rin[29] /*18978*/;
  assign r_0[30] = rin[30] /*18977*/;
  assign r_0[31] = rin[31] /*18976*/;
  assign r_0[32] = rin[32] /*18975*/;
  assign r_0[33] = rin[33] /*18974*/;
  assign r_0[34] = rin[34] /*18973*/;
  assign r_0[35] = rin[35] /*18972*/;
  assign r_0[36] = rin[36] /*18971*/;
  assign r_0[37] = rin[37] /*18970*/;
  assign r_0[38] = rin[38] /*18969*/;
  assign r_0[39] = rin[39] /*18968*/;
  assign r_0[40] = rin[40] /*18967*/;
  assign r_0[41] = rin[41] /*18966*/;
  assign r_0[42] = rin[42] /*18965*/;
  assign r_0[43] = rin[43] /*18964*/;
  assign r_0[44] = rin[44] /*18963*/;
  assign r_0[45] = rin[45] /*18962*/;
  assign r_0[46] = zeroWire /*18961*/;
  assign inv_1[0] = ~div[0] /*18960*/;
  assign inv_1[1] = ~div[1] /*18959*/;
  assign inv_1[2] = ~div[2] /*18958*/;
  assign inv_1[3] = ~div[3] /*18957*/;
  assign inv_1[4] = ~div[4] /*18956*/;
  assign inv_1[5] = ~div[5] /*18955*/;
  assign inv_1[6] = ~div[6] /*18954*/;
  assign inv_1[7] = ~div[7] /*18953*/;
  assign inv_1[8] = ~div[8] /*18952*/;
  assign inv_1[9] = ~div[9] /*18951*/;
  assign inv_1[10] = ~div[10] /*18950*/;
  assign inv_1[11] = ~div[11] /*18949*/;
  assign inv_1[12] = ~div[12] /*18948*/;
  assign inv_1[13] = ~div[13] /*18947*/;
  assign inv_1[14] = ~div[14] /*18946*/;
  assign inv_1[15] = ~div[15] /*18945*/;
  assign inv_1[16] = ~div[16] /*18944*/;
  assign inv_1[17] = ~div[17] /*18943*/;
  assign inv_1[18] = ~div[18] /*18942*/;
  assign inv_1[19] = ~div[19] /*18941*/;
  assign inv_1[20] = ~div[20] /*18940*/;
  assign inv_1[21] = ~div[21] /*18939*/;
  assign inv_1[22] = ~div[22] /*18938*/;
assign inv_1[23] = oneWire /*18937*/;
  assign _0_ = inv_1[0] ^ r_0[23] /*18935*/;
  assign sum_1[0] = _0_ ^ oneWire /*18934*/;
  assign _1_ = _0_ & oneWire /*18933*/;
  assign _2_ = inv_1[0] & r_0[23] /*18932*/;
  assign _3_ = _1_ | _2_ /*18931*/;
  assign _4_ = inv_1[1] ^ r_0[24] /*18930*/;
  assign sum_1[1] = _4_ ^ _3_ /*18929*/;
  assign _5_ = _4_ & _3_ /*18928*/;
  assign _6_ = inv_1[1] & r_0[24] /*18927*/;
  assign _7_ = _5_ | _6_ /*18926*/;
  assign _8_ = inv_1[2] ^ r_0[25] /*18924*/;
  assign sum_1[2] = _8_ ^ _7_ /*18923*/;
  assign _9_ = _8_ & _7_ /*18922*/;
  assign _10_ = inv_1[2] & r_0[25] /*18921*/;
  assign _11_ = _9_ | _10_ /*18920*/;
  assign _12_ = inv_1[3] ^ r_0[26] /*18918*/;
  assign sum_1[3] = _12_ ^ _11_ /*18917*/;
  assign _13_ = _12_ & _11_ /*18916*/;
  assign _14_ = inv_1[3] & r_0[26] /*18915*/;
  assign _15_ = _13_ | _14_ /*18914*/;
  assign _16_ = inv_1[4] ^ r_0[27] /*18912*/;
  assign sum_1[4] = _16_ ^ _15_ /*18911*/;
  assign _17_ = _16_ & _15_ /*18910*/;
  assign _18_ = inv_1[4] & r_0[27] /*18909*/;
  assign _19_ = _17_ | _18_ /*18908*/;
  assign _20_ = inv_1[5] ^ r_0[28] /*18906*/;
  assign sum_1[5] = _20_ ^ _19_ /*18905*/;
  assign _21_ = _20_ & _19_ /*18904*/;
  assign _22_ = inv_1[5] & r_0[28] /*18903*/;
  assign _23_ = _21_ | _22_ /*18902*/;
  assign _24_ = inv_1[6] ^ r_0[29] /*18900*/;
  assign sum_1[6] = _24_ ^ _23_ /*18899*/;
  assign _25_ = _24_ & _23_ /*18898*/;
  assign _26_ = inv_1[6] & r_0[29] /*18897*/;
  assign _27_ = _25_ | _26_ /*18896*/;
  assign _28_ = inv_1[7] ^ r_0[30] /*18894*/;
  assign sum_1[7] = _28_ ^ _27_ /*18893*/;
  assign _29_ = _28_ & _27_ /*18892*/;
  assign _30_ = inv_1[7] & r_0[30] /*18891*/;
  assign _31_ = _29_ | _30_ /*18890*/;
  assign _32_ = inv_1[8] ^ r_0[31] /*18888*/;
  assign sum_1[8] = _32_ ^ _31_ /*18887*/;
  assign _33_ = _32_ & _31_ /*18886*/;
  assign _34_ = inv_1[8] & r_0[31] /*18885*/;
  assign _35_ = _33_ | _34_ /*18884*/;
  assign _36_ = inv_1[9] ^ r_0[32] /*18882*/;
  assign sum_1[9] = _36_ ^ _35_ /*18881*/;
  assign _37_ = _36_ & _35_ /*18880*/;
  assign _38_ = inv_1[9] & r_0[32] /*18879*/;
  assign _39_ = _37_ | _38_ /*18878*/;
  assign _40_ = inv_1[10] ^ r_0[33] /*18876*/;
  assign sum_1[10] = _40_ ^ _39_ /*18875*/;
  assign _41_ = _40_ & _39_ /*18874*/;
  assign _42_ = inv_1[10] & r_0[33] /*18873*/;
  assign _43_ = _41_ | _42_ /*18872*/;
  assign _44_ = inv_1[11] ^ r_0[34] /*18870*/;
  assign sum_1[11] = _44_ ^ _43_ /*18869*/;
  assign _45_ = _44_ & _43_ /*18868*/;
  assign _46_ = inv_1[11] & r_0[34] /*18867*/;
  assign _47_ = _45_ | _46_ /*18866*/;
  assign _48_ = inv_1[12] ^ r_0[35] /*18864*/;
  assign sum_1[12] = _48_ ^ _47_ /*18863*/;
  assign _49_ = _48_ & _47_ /*18862*/;
  assign _50_ = inv_1[12] & r_0[35] /*18861*/;
  assign _51_ = _49_ | _50_ /*18860*/;
  assign _52_ = inv_1[13] ^ r_0[36] /*18858*/;
  assign sum_1[13] = _52_ ^ _51_ /*18857*/;
  assign _53_ = _52_ & _51_ /*18856*/;
  assign _54_ = inv_1[13] & r_0[36] /*18855*/;
  assign _55_ = _53_ | _54_ /*18854*/;
  assign _56_ = inv_1[14] ^ r_0[37] /*18852*/;
  assign sum_1[14] = _56_ ^ _55_ /*18851*/;
  assign _57_ = _56_ & _55_ /*18850*/;
  assign _58_ = inv_1[14] & r_0[37] /*18849*/;
  assign _59_ = _57_ | _58_ /*18848*/;
  assign _60_ = inv_1[15] ^ r_0[38] /*18846*/;
  assign sum_1[15] = _60_ ^ _59_ /*18845*/;
  assign _61_ = _60_ & _59_ /*18844*/;
  assign _62_ = inv_1[15] & r_0[38] /*18843*/;
  assign _63_ = _61_ | _62_ /*18842*/;
  assign _64_ = inv_1[16] ^ r_0[39] /*18840*/;
  assign sum_1[16] = _64_ ^ _63_ /*18839*/;
  assign _65_ = _64_ & _63_ /*18838*/;
  assign _66_ = inv_1[16] & r_0[39] /*18837*/;
  assign _67_ = _65_ | _66_ /*18836*/;
  assign _68_ = inv_1[17] ^ r_0[40] /*18834*/;
  assign sum_1[17] = _68_ ^ _67_ /*18833*/;
  assign _69_ = _68_ & _67_ /*18832*/;
  assign _70_ = inv_1[17] & r_0[40] /*18831*/;
  assign _71_ = _69_ | _70_ /*18830*/;
  assign _72_ = inv_1[18] ^ r_0[41] /*18828*/;
  assign sum_1[18] = _72_ ^ _71_ /*18827*/;
  assign _73_ = _72_ & _71_ /*18826*/;
  assign _74_ = inv_1[18] & r_0[41] /*18825*/;
  assign _75_ = _73_ | _74_ /*18824*/;
  assign _76_ = inv_1[19] ^ r_0[42] /*18822*/;
  assign sum_1[19] = _76_ ^ _75_ /*18821*/;
  assign _77_ = _76_ & _75_ /*18820*/;
  assign _78_ = inv_1[19] & r_0[42] /*18819*/;
  assign _79_ = _77_ | _78_ /*18818*/;
  assign _80_ = inv_1[20] ^ r_0[43] /*18816*/;
  assign sum_1[20] = _80_ ^ _79_ /*18815*/;
  assign _81_ = _80_ & _79_ /*18814*/;
  assign _82_ = inv_1[20] & r_0[43] /*18813*/;
  assign _83_ = _81_ | _82_ /*18812*/;
  assign _84_ = inv_1[21] ^ r_0[44] /*18810*/;
  assign sum_1[21] = _84_ ^ _83_ /*18809*/;
  assign _85_ = _84_ & _83_ /*18808*/;
  assign _86_ = inv_1[21] & r_0[44] /*18807*/;
  assign _87_ = _85_ | _86_ /*18806*/;
  assign _88_ = inv_1[22] ^ r_0[45] /*18804*/;
  assign sum_1[22] = _88_ ^ _87_ /*18803*/;
  assign _89_ = _88_ & _87_ /*18802*/;
  assign _90_ = inv_1[22] & r_0[45] /*18801*/;
  assign _91_ = _89_ | _90_ /*18800*/;
  assign _92_ = inv_1[23] ^ r_0[46] /*18798*/;
  assign sum_1[23] = _92_ ^ _91_ /*18797*/;
  assign _93_ = _92_ & _91_ /*18796*/;
  assign _94_ = inv_1[23] & r_0[46] /*18795*/;
  assign _95_ = _93_ | _94_ /*18794*/;
  assign q[23] = ~sum_1[23] /*18813*/;
  assign m_1[0] = r_0[23] /*18812*/;
  assign m_1[1] = r_0[24] /*18811*/;
  assign m_1[2] = r_0[25] /*18810*/;
  assign m_1[3] = r_0[26] /*18809*/;
  assign m_1[4] = r_0[27] /*18808*/;
  assign m_1[5] = r_0[28] /*18807*/;
  assign m_1[6] = r_0[29] /*18806*/;
  assign m_1[7] = r_0[30] /*18805*/;
  assign m_1[8] = r_0[31] /*18804*/;
  assign m_1[9] = r_0[32] /*18803*/;
  assign m_1[10] = r_0[33] /*18802*/;
  assign m_1[11] = r_0[34] /*18801*/;
  assign m_1[12] = r_0[35] /*18800*/;
  assign m_1[13] = r_0[36] /*18799*/;
  assign m_1[14] = r_0[37] /*18798*/;
  assign m_1[15] = r_0[38] /*18797*/;
  assign m_1[16] = r_0[39] /*18796*/;
  assign m_1[17] = r_0[40] /*18795*/;
  assign m_1[18] = r_0[41] /*18794*/;
  assign m_1[19] = r_0[42] /*18793*/;
  assign m_1[20] = r_0[43] /*18792*/;
  assign m_1[21] = r_0[44] /*18791*/;
  assign m_1[22] = r_0[45] /*18790*/;
  assign m_1[23] = r_0[46] /*18789*/;
  assign _96_ = ~q[23] /*18787*/;
  assign _97_ = sum_1[0] & q[23] /*18786*/;
  assign _98_ = m_1[0] & _96_ /*18785*/;
  assign r_1[23] = _98_ | _97_ /*18784*/;
  assign _99_ = ~q[23] /*18783*/;
  assign _100_ = sum_1[1] & q[23] /*18782*/;
  assign _101_ = m_1[1] & _99_ /*18781*/;
  assign r_1[24] = _101_ | _100_ /*18780*/;
  assign _102_ = ~q[23] /*18779*/;
  assign _103_ = sum_1[2] & q[23] /*18778*/;
  assign _104_ = m_1[2] & _102_ /*18777*/;
  assign r_1[25] = _104_ | _103_ /*18776*/;
  assign _105_ = ~q[23] /*18775*/;
  assign _106_ = sum_1[3] & q[23] /*18774*/;
  assign _107_ = m_1[3] & _105_ /*18773*/;
  assign r_1[26] = _107_ | _106_ /*18772*/;
  assign _108_ = ~q[23] /*18771*/;
  assign _109_ = sum_1[4] & q[23] /*18770*/;
  assign _110_ = m_1[4] & _108_ /*18769*/;
  assign r_1[27] = _110_ | _109_ /*18768*/;
  assign _111_ = ~q[23] /*18767*/;
  assign _112_ = sum_1[5] & q[23] /*18766*/;
  assign _113_ = m_1[5] & _111_ /*18765*/;
  assign r_1[28] = _113_ | _112_ /*18764*/;
  assign _114_ = ~q[23] /*18763*/;
  assign _115_ = sum_1[6] & q[23] /*18762*/;
  assign _116_ = m_1[6] & _114_ /*18761*/;
  assign r_1[29] = _116_ | _115_ /*18760*/;
  assign _117_ = ~q[23] /*18759*/;
  assign _118_ = sum_1[7] & q[23] /*18758*/;
  assign _119_ = m_1[7] & _117_ /*18757*/;
  assign r_1[30] = _119_ | _118_ /*18756*/;
  assign _120_ = ~q[23] /*18755*/;
  assign _121_ = sum_1[8] & q[23] /*18754*/;
  assign _122_ = m_1[8] & _120_ /*18753*/;
  assign r_1[31] = _122_ | _121_ /*18752*/;
  assign _123_ = ~q[23] /*18751*/;
  assign _124_ = sum_1[9] & q[23] /*18750*/;
  assign _125_ = m_1[9] & _123_ /*18749*/;
  assign r_1[32] = _125_ | _124_ /*18748*/;
  assign _126_ = ~q[23] /*18747*/;
  assign _127_ = sum_1[10] & q[23] /*18746*/;
  assign _128_ = m_1[10] & _126_ /*18745*/;
  assign r_1[33] = _128_ | _127_ /*18744*/;
  assign _129_ = ~q[23] /*18743*/;
  assign _130_ = sum_1[11] & q[23] /*18742*/;
  assign _131_ = m_1[11] & _129_ /*18741*/;
  assign r_1[34] = _131_ | _130_ /*18740*/;
  assign _132_ = ~q[23] /*18739*/;
  assign _133_ = sum_1[12] & q[23] /*18738*/;
  assign _134_ = m_1[12] & _132_ /*18737*/;
  assign r_1[35] = _134_ | _133_ /*18736*/;
  assign _135_ = ~q[23] /*18735*/;
  assign _136_ = sum_1[13] & q[23] /*18734*/;
  assign _137_ = m_1[13] & _135_ /*18733*/;
  assign r_1[36] = _137_ | _136_ /*18732*/;
  assign _138_ = ~q[23] /*18731*/;
  assign _139_ = sum_1[14] & q[23] /*18730*/;
  assign _140_ = m_1[14] & _138_ /*18729*/;
  assign r_1[37] = _140_ | _139_ /*18728*/;
  assign _141_ = ~q[23] /*18727*/;
  assign _142_ = sum_1[15] & q[23] /*18726*/;
  assign _143_ = m_1[15] & _141_ /*18725*/;
  assign r_1[38] = _143_ | _142_ /*18724*/;
  assign _144_ = ~q[23] /*18723*/;
  assign _145_ = sum_1[16] & q[23] /*18722*/;
  assign _146_ = m_1[16] & _144_ /*18721*/;
  assign r_1[39] = _146_ | _145_ /*18720*/;
  assign _147_ = ~q[23] /*18719*/;
  assign _148_ = sum_1[17] & q[23] /*18718*/;
  assign _149_ = m_1[17] & _147_ /*18717*/;
  assign r_1[40] = _149_ | _148_ /*18716*/;
  assign _150_ = ~q[23] /*18715*/;
  assign _151_ = sum_1[18] & q[23] /*18714*/;
  assign _152_ = m_1[18] & _150_ /*18713*/;
  assign r_1[41] = _152_ | _151_ /*18712*/;
  assign _153_ = ~q[23] /*18711*/;
  assign _154_ = sum_1[19] & q[23] /*18710*/;
  assign _155_ = m_1[19] & _153_ /*18709*/;
  assign r_1[42] = _155_ | _154_ /*18708*/;
  assign _156_ = ~q[23] /*18707*/;
  assign _157_ = sum_1[20] & q[23] /*18706*/;
  assign _158_ = m_1[20] & _156_ /*18705*/;
  assign r_1[43] = _158_ | _157_ /*18704*/;
  assign _159_ = ~q[23] /*18703*/;
  assign _160_ = sum_1[21] & q[23] /*18702*/;
  assign _161_ = m_1[21] & _159_ /*18701*/;
  assign r_1[44] = _161_ | _160_ /*18700*/;
  assign _162_ = ~q[23] /*18699*/;
  assign _163_ = sum_1[22] & q[23] /*18698*/;
  assign _164_ = m_1[22] & _162_ /*18697*/;
  assign r_1[45] = _164_ | _163_ /*18696*/;
  assign _165_ = ~q[23] /*18695*/;
  assign _166_ = sum_1[23] & q[23] /*18694*/;
  assign _167_ = m_1[23] & _165_ /*18693*/;
  assign r_1[46] = _167_ | _166_ /*18692*/;
assign r_1[0]= r_0[0] /*18691*/;
assign r_1[1]= r_0[1] /*18690*/;
assign r_1[2]= r_0[2] /*18689*/;
assign r_1[3]= r_0[3] /*18688*/;
assign r_1[4]= r_0[4] /*18687*/;
assign r_1[5]= r_0[5] /*18686*/;
assign r_1[6]= r_0[6] /*18685*/;
assign r_1[7]= r_0[7] /*18684*/;
assign r_1[8]= r_0[8] /*18683*/;
assign r_1[9]= r_0[9] /*18682*/;
assign r_1[10]= r_0[10] /*18681*/;
assign r_1[11]= r_0[11] /*18680*/;
assign r_1[12]= r_0[12] /*18679*/;
assign r_1[13]= r_0[13] /*18678*/;
assign r_1[14]= r_0[14] /*18677*/;
assign r_1[15]= r_0[15] /*18676*/;
assign r_1[16]= r_0[16] /*18675*/;
assign r_1[17]= r_0[17] /*18674*/;
assign r_1[18]= r_0[18] /*18673*/;
assign r_1[19]= r_0[19] /*18672*/;
assign r_1[20]= r_0[20] /*18671*/;
assign r_1[21]= r_0[21] /*18670*/;
assign r_1[22]= r_0[22] /*18669*/;
  assign inv_2[0] = ~div[0] /*18624*/;
  assign inv_2[1] = ~div[1] /*18623*/;
  assign inv_2[2] = ~div[2] /*18622*/;
  assign inv_2[3] = ~div[3] /*18621*/;
  assign inv_2[4] = ~div[4] /*18620*/;
  assign inv_2[5] = ~div[5] /*18619*/;
  assign inv_2[6] = ~div[6] /*18618*/;
  assign inv_2[7] = ~div[7] /*18617*/;
  assign inv_2[8] = ~div[8] /*18616*/;
  assign inv_2[9] = ~div[9] /*18615*/;
  assign inv_2[10] = ~div[10] /*18614*/;
  assign inv_2[11] = ~div[11] /*18613*/;
  assign inv_2[12] = ~div[12] /*18612*/;
  assign inv_2[13] = ~div[13] /*18611*/;
  assign inv_2[14] = ~div[14] /*18610*/;
  assign inv_2[15] = ~div[15] /*18609*/;
  assign inv_2[16] = ~div[16] /*18608*/;
  assign inv_2[17] = ~div[17] /*18607*/;
  assign inv_2[18] = ~div[18] /*18606*/;
  assign inv_2[19] = ~div[19] /*18605*/;
  assign inv_2[20] = ~div[20] /*18604*/;
  assign inv_2[21] = ~div[21] /*18603*/;
  assign inv_2[22] = ~div[22] /*18602*/;
assign inv_2[23] = oneWire /*18601*/;
  assign _168_ = inv_2[0] ^ r_1[22] /*18599*/;
  assign sum_2[0] = _168_ ^ oneWire /*18598*/;
  assign _169_ = _168_ & oneWire /*18597*/;
  assign _170_ = inv_2[0] & r_1[22] /*18596*/;
  assign _171_ = _169_ | _170_ /*18595*/;
  assign _172_ = inv_2[1] ^ r_1[23] /*18594*/;
  assign sum_2[1] = _172_ ^ _171_ /*18593*/;
  assign _173_ = _172_ & _171_ /*18592*/;
  assign _174_ = inv_2[1] & r_1[23] /*18591*/;
  assign _175_ = _173_ | _174_ /*18590*/;
  assign _176_ = inv_2[2] ^ r_1[24] /*18588*/;
  assign sum_2[2] = _176_ ^ _175_ /*18587*/;
  assign _177_ = _176_ & _175_ /*18586*/;
  assign _178_ = inv_2[2] & r_1[24] /*18585*/;
  assign _179_ = _177_ | _178_ /*18584*/;
  assign _180_ = inv_2[3] ^ r_1[25] /*18582*/;
  assign sum_2[3] = _180_ ^ _179_ /*18581*/;
  assign _181_ = _180_ & _179_ /*18580*/;
  assign _182_ = inv_2[3] & r_1[25] /*18579*/;
  assign _183_ = _181_ | _182_ /*18578*/;
  assign _184_ = inv_2[4] ^ r_1[26] /*18576*/;
  assign sum_2[4] = _184_ ^ _183_ /*18575*/;
  assign _185_ = _184_ & _183_ /*18574*/;
  assign _186_ = inv_2[4] & r_1[26] /*18573*/;
  assign _187_ = _185_ | _186_ /*18572*/;
  assign _188_ = inv_2[5] ^ r_1[27] /*18570*/;
  assign sum_2[5] = _188_ ^ _187_ /*18569*/;
  assign _189_ = _188_ & _187_ /*18568*/;
  assign _190_ = inv_2[5] & r_1[27] /*18567*/;
  assign _191_ = _189_ | _190_ /*18566*/;
  assign _192_ = inv_2[6] ^ r_1[28] /*18564*/;
  assign sum_2[6] = _192_ ^ _191_ /*18563*/;
  assign _193_ = _192_ & _191_ /*18562*/;
  assign _194_ = inv_2[6] & r_1[28] /*18561*/;
  assign _195_ = _193_ | _194_ /*18560*/;
  assign _196_ = inv_2[7] ^ r_1[29] /*18558*/;
  assign sum_2[7] = _196_ ^ _195_ /*18557*/;
  assign _197_ = _196_ & _195_ /*18556*/;
  assign _198_ = inv_2[7] & r_1[29] /*18555*/;
  assign _199_ = _197_ | _198_ /*18554*/;
  assign _200_ = inv_2[8] ^ r_1[30] /*18552*/;
  assign sum_2[8] = _200_ ^ _199_ /*18551*/;
  assign _201_ = _200_ & _199_ /*18550*/;
  assign _202_ = inv_2[8] & r_1[30] /*18549*/;
  assign _203_ = _201_ | _202_ /*18548*/;
  assign _204_ = inv_2[9] ^ r_1[31] /*18546*/;
  assign sum_2[9] = _204_ ^ _203_ /*18545*/;
  assign _205_ = _204_ & _203_ /*18544*/;
  assign _206_ = inv_2[9] & r_1[31] /*18543*/;
  assign _207_ = _205_ | _206_ /*18542*/;
  assign _208_ = inv_2[10] ^ r_1[32] /*18540*/;
  assign sum_2[10] = _208_ ^ _207_ /*18539*/;
  assign _209_ = _208_ & _207_ /*18538*/;
  assign _210_ = inv_2[10] & r_1[32] /*18537*/;
  assign _211_ = _209_ | _210_ /*18536*/;
  assign _212_ = inv_2[11] ^ r_1[33] /*18534*/;
  assign sum_2[11] = _212_ ^ _211_ /*18533*/;
  assign _213_ = _212_ & _211_ /*18532*/;
  assign _214_ = inv_2[11] & r_1[33] /*18531*/;
  assign _215_ = _213_ | _214_ /*18530*/;
  assign _216_ = inv_2[12] ^ r_1[34] /*18528*/;
  assign sum_2[12] = _216_ ^ _215_ /*18527*/;
  assign _217_ = _216_ & _215_ /*18526*/;
  assign _218_ = inv_2[12] & r_1[34] /*18525*/;
  assign _219_ = _217_ | _218_ /*18524*/;
  assign _220_ = inv_2[13] ^ r_1[35] /*18522*/;
  assign sum_2[13] = _220_ ^ _219_ /*18521*/;
  assign _221_ = _220_ & _219_ /*18520*/;
  assign _222_ = inv_2[13] & r_1[35] /*18519*/;
  assign _223_ = _221_ | _222_ /*18518*/;
  assign _224_ = inv_2[14] ^ r_1[36] /*18516*/;
  assign sum_2[14] = _224_ ^ _223_ /*18515*/;
  assign _225_ = _224_ & _223_ /*18514*/;
  assign _226_ = inv_2[14] & r_1[36] /*18513*/;
  assign _227_ = _225_ | _226_ /*18512*/;
  assign _228_ = inv_2[15] ^ r_1[37] /*18510*/;
  assign sum_2[15] = _228_ ^ _227_ /*18509*/;
  assign _229_ = _228_ & _227_ /*18508*/;
  assign _230_ = inv_2[15] & r_1[37] /*18507*/;
  assign _231_ = _229_ | _230_ /*18506*/;
  assign _232_ = inv_2[16] ^ r_1[38] /*18504*/;
  assign sum_2[16] = _232_ ^ _231_ /*18503*/;
  assign _233_ = _232_ & _231_ /*18502*/;
  assign _234_ = inv_2[16] & r_1[38] /*18501*/;
  assign _235_ = _233_ | _234_ /*18500*/;
  assign _236_ = inv_2[17] ^ r_1[39] /*18498*/;
  assign sum_2[17] = _236_ ^ _235_ /*18497*/;
  assign _237_ = _236_ & _235_ /*18496*/;
  assign _238_ = inv_2[17] & r_1[39] /*18495*/;
  assign _239_ = _237_ | _238_ /*18494*/;
  assign _240_ = inv_2[18] ^ r_1[40] /*18492*/;
  assign sum_2[18] = _240_ ^ _239_ /*18491*/;
  assign _241_ = _240_ & _239_ /*18490*/;
  assign _242_ = inv_2[18] & r_1[40] /*18489*/;
  assign _243_ = _241_ | _242_ /*18488*/;
  assign _244_ = inv_2[19] ^ r_1[41] /*18486*/;
  assign sum_2[19] = _244_ ^ _243_ /*18485*/;
  assign _245_ = _244_ & _243_ /*18484*/;
  assign _246_ = inv_2[19] & r_1[41] /*18483*/;
  assign _247_ = _245_ | _246_ /*18482*/;
  assign _248_ = inv_2[20] ^ r_1[42] /*18480*/;
  assign sum_2[20] = _248_ ^ _247_ /*18479*/;
  assign _249_ = _248_ & _247_ /*18478*/;
  assign _250_ = inv_2[20] & r_1[42] /*18477*/;
  assign _251_ = _249_ | _250_ /*18476*/;
  assign _252_ = inv_2[21] ^ r_1[43] /*18474*/;
  assign sum_2[21] = _252_ ^ _251_ /*18473*/;
  assign _253_ = _252_ & _251_ /*18472*/;
  assign _254_ = inv_2[21] & r_1[43] /*18471*/;
  assign _255_ = _253_ | _254_ /*18470*/;
  assign _256_ = inv_2[22] ^ r_1[44] /*18468*/;
  assign sum_2[22] = _256_ ^ _255_ /*18467*/;
  assign _257_ = _256_ & _255_ /*18466*/;
  assign _258_ = inv_2[22] & r_1[44] /*18465*/;
  assign _259_ = _257_ | _258_ /*18464*/;
  assign _260_ = inv_2[23] ^ r_1[45] /*18462*/;
  assign sum_2[23] = _260_ ^ _259_ /*18461*/;
  assign _261_ = _260_ & _259_ /*18460*/;
  assign _262_ = inv_2[23] & r_1[45] /*18459*/;
  assign _263_ = _261_ | _262_ /*18458*/;
  assign q[22] = ~sum_2[23] /*18477*/;
  assign m_2[0] = r_1[22] /*18476*/;
  assign m_2[1] = r_1[23] /*18475*/;
  assign m_2[2] = r_1[24] /*18474*/;
  assign m_2[3] = r_1[25] /*18473*/;
  assign m_2[4] = r_1[26] /*18472*/;
  assign m_2[5] = r_1[27] /*18471*/;
  assign m_2[6] = r_1[28] /*18470*/;
  assign m_2[7] = r_1[29] /*18469*/;
  assign m_2[8] = r_1[30] /*18468*/;
  assign m_2[9] = r_1[31] /*18467*/;
  assign m_2[10] = r_1[32] /*18466*/;
  assign m_2[11] = r_1[33] /*18465*/;
  assign m_2[12] = r_1[34] /*18464*/;
  assign m_2[13] = r_1[35] /*18463*/;
  assign m_2[14] = r_1[36] /*18462*/;
  assign m_2[15] = r_1[37] /*18461*/;
  assign m_2[16] = r_1[38] /*18460*/;
  assign m_2[17] = r_1[39] /*18459*/;
  assign m_2[18] = r_1[40] /*18458*/;
  assign m_2[19] = r_1[41] /*18457*/;
  assign m_2[20] = r_1[42] /*18456*/;
  assign m_2[21] = r_1[43] /*18455*/;
  assign m_2[22] = r_1[44] /*18454*/;
  assign m_2[23] = r_1[45] /*18453*/;
  assign _264_ = ~q[22] /*18451*/;
  assign _265_ = sum_2[0] & q[22] /*18450*/;
  assign _266_ = m_2[0] & _264_ /*18449*/;
  assign r_2[22] = _266_ | _265_ /*18448*/;
  assign _267_ = ~q[22] /*18447*/;
  assign _268_ = sum_2[1] & q[22] /*18446*/;
  assign _269_ = m_2[1] & _267_ /*18445*/;
  assign r_2[23] = _269_ | _268_ /*18444*/;
  assign _270_ = ~q[22] /*18443*/;
  assign _271_ = sum_2[2] & q[22] /*18442*/;
  assign _272_ = m_2[2] & _270_ /*18441*/;
  assign r_2[24] = _272_ | _271_ /*18440*/;
  assign _273_ = ~q[22] /*18439*/;
  assign _274_ = sum_2[3] & q[22] /*18438*/;
  assign _275_ = m_2[3] & _273_ /*18437*/;
  assign r_2[25] = _275_ | _274_ /*18436*/;
  assign _276_ = ~q[22] /*18435*/;
  assign _277_ = sum_2[4] & q[22] /*18434*/;
  assign _278_ = m_2[4] & _276_ /*18433*/;
  assign r_2[26] = _278_ | _277_ /*18432*/;
  assign _279_ = ~q[22] /*18431*/;
  assign _280_ = sum_2[5] & q[22] /*18430*/;
  assign _281_ = m_2[5] & _279_ /*18429*/;
  assign r_2[27] = _281_ | _280_ /*18428*/;
  assign _282_ = ~q[22] /*18427*/;
  assign _283_ = sum_2[6] & q[22] /*18426*/;
  assign _284_ = m_2[6] & _282_ /*18425*/;
  assign r_2[28] = _284_ | _283_ /*18424*/;
  assign _285_ = ~q[22] /*18423*/;
  assign _286_ = sum_2[7] & q[22] /*18422*/;
  assign _287_ = m_2[7] & _285_ /*18421*/;
  assign r_2[29] = _287_ | _286_ /*18420*/;
  assign _288_ = ~q[22] /*18419*/;
  assign _289_ = sum_2[8] & q[22] /*18418*/;
  assign _290_ = m_2[8] & _288_ /*18417*/;
  assign r_2[30] = _290_ | _289_ /*18416*/;
  assign _291_ = ~q[22] /*18415*/;
  assign _292_ = sum_2[9] & q[22] /*18414*/;
  assign _293_ = m_2[9] & _291_ /*18413*/;
  assign r_2[31] = _293_ | _292_ /*18412*/;
  assign _294_ = ~q[22] /*18411*/;
  assign _295_ = sum_2[10] & q[22] /*18410*/;
  assign _296_ = m_2[10] & _294_ /*18409*/;
  assign r_2[32] = _296_ | _295_ /*18408*/;
  assign _297_ = ~q[22] /*18407*/;
  assign _298_ = sum_2[11] & q[22] /*18406*/;
  assign _299_ = m_2[11] & _297_ /*18405*/;
  assign r_2[33] = _299_ | _298_ /*18404*/;
  assign _300_ = ~q[22] /*18403*/;
  assign _301_ = sum_2[12] & q[22] /*18402*/;
  assign _302_ = m_2[12] & _300_ /*18401*/;
  assign r_2[34] = _302_ | _301_ /*18400*/;
  assign _303_ = ~q[22] /*18399*/;
  assign _304_ = sum_2[13] & q[22] /*18398*/;
  assign _305_ = m_2[13] & _303_ /*18397*/;
  assign r_2[35] = _305_ | _304_ /*18396*/;
  assign _306_ = ~q[22] /*18395*/;
  assign _307_ = sum_2[14] & q[22] /*18394*/;
  assign _308_ = m_2[14] & _306_ /*18393*/;
  assign r_2[36] = _308_ | _307_ /*18392*/;
  assign _309_ = ~q[22] /*18391*/;
  assign _310_ = sum_2[15] & q[22] /*18390*/;
  assign _311_ = m_2[15] & _309_ /*18389*/;
  assign r_2[37] = _311_ | _310_ /*18388*/;
  assign _312_ = ~q[22] /*18387*/;
  assign _313_ = sum_2[16] & q[22] /*18386*/;
  assign _314_ = m_2[16] & _312_ /*18385*/;
  assign r_2[38] = _314_ | _313_ /*18384*/;
  assign _315_ = ~q[22] /*18383*/;
  assign _316_ = sum_2[17] & q[22] /*18382*/;
  assign _317_ = m_2[17] & _315_ /*18381*/;
  assign r_2[39] = _317_ | _316_ /*18380*/;
  assign _318_ = ~q[22] /*18379*/;
  assign _319_ = sum_2[18] & q[22] /*18378*/;
  assign _320_ = m_2[18] & _318_ /*18377*/;
  assign r_2[40] = _320_ | _319_ /*18376*/;
  assign _321_ = ~q[22] /*18375*/;
  assign _322_ = sum_2[19] & q[22] /*18374*/;
  assign _323_ = m_2[19] & _321_ /*18373*/;
  assign r_2[41] = _323_ | _322_ /*18372*/;
  assign _324_ = ~q[22] /*18371*/;
  assign _325_ = sum_2[20] & q[22] /*18370*/;
  assign _326_ = m_2[20] & _324_ /*18369*/;
  assign r_2[42] = _326_ | _325_ /*18368*/;
  assign _327_ = ~q[22] /*18367*/;
  assign _328_ = sum_2[21] & q[22] /*18366*/;
  assign _329_ = m_2[21] & _327_ /*18365*/;
  assign r_2[43] = _329_ | _328_ /*18364*/;
  assign _330_ = ~q[22] /*18363*/;
  assign _331_ = sum_2[22] & q[22] /*18362*/;
  assign _332_ = m_2[22] & _330_ /*18361*/;
  assign r_2[44] = _332_ | _331_ /*18360*/;
  assign _333_ = ~q[22] /*18359*/;
  assign _334_ = sum_2[23] & q[22] /*18358*/;
  assign _335_ = m_2[23] & _333_ /*18357*/;
  assign r_2[45] = _335_ | _334_ /*18356*/;
assign r_2[0]= r_1[0] /*18355*/;
assign r_2[1]= r_1[1] /*18354*/;
assign r_2[2]= r_1[2] /*18353*/;
assign r_2[3]= r_1[3] /*18352*/;
assign r_2[4]= r_1[4] /*18351*/;
assign r_2[5]= r_1[5] /*18350*/;
assign r_2[6]= r_1[6] /*18349*/;
assign r_2[7]= r_1[7] /*18348*/;
assign r_2[8]= r_1[8] /*18347*/;
assign r_2[9]= r_1[9] /*18346*/;
assign r_2[10]= r_1[10] /*18345*/;
assign r_2[11]= r_1[11] /*18344*/;
assign r_2[12]= r_1[12] /*18343*/;
assign r_2[13]= r_1[13] /*18342*/;
assign r_2[14]= r_1[14] /*18341*/;
assign r_2[15]= r_1[15] /*18340*/;
assign r_2[16]= r_1[16] /*18339*/;
assign r_2[17]= r_1[17] /*18338*/;
assign r_2[18]= r_1[18] /*18337*/;
assign r_2[19]= r_1[19] /*18336*/;
assign r_2[20]= r_1[20] /*18335*/;
assign r_2[21]= r_1[21] /*18334*/;
  assign inv_3[0] = ~div[0] /*18288*/;
  assign inv_3[1] = ~div[1] /*18287*/;
  assign inv_3[2] = ~div[2] /*18286*/;
  assign inv_3[3] = ~div[3] /*18285*/;
  assign inv_3[4] = ~div[4] /*18284*/;
  assign inv_3[5] = ~div[5] /*18283*/;
  assign inv_3[6] = ~div[6] /*18282*/;
  assign inv_3[7] = ~div[7] /*18281*/;
  assign inv_3[8] = ~div[8] /*18280*/;
  assign inv_3[9] = ~div[9] /*18279*/;
  assign inv_3[10] = ~div[10] /*18278*/;
  assign inv_3[11] = ~div[11] /*18277*/;
  assign inv_3[12] = ~div[12] /*18276*/;
  assign inv_3[13] = ~div[13] /*18275*/;
  assign inv_3[14] = ~div[14] /*18274*/;
  assign inv_3[15] = ~div[15] /*18273*/;
  assign inv_3[16] = ~div[16] /*18272*/;
  assign inv_3[17] = ~div[17] /*18271*/;
  assign inv_3[18] = ~div[18] /*18270*/;
  assign inv_3[19] = ~div[19] /*18269*/;
  assign inv_3[20] = ~div[20] /*18268*/;
  assign inv_3[21] = ~div[21] /*18267*/;
  assign inv_3[22] = ~div[22] /*18266*/;
assign inv_3[23] = oneWire /*18265*/;
  assign _336_ = inv_3[0] ^ r_2[21] /*18263*/;
  assign sum_3[0] = _336_ ^ oneWire /*18262*/;
  assign _337_ = _336_ & oneWire /*18261*/;
  assign _338_ = inv_3[0] & r_2[21] /*18260*/;
  assign _339_ = _337_ | _338_ /*18259*/;
  assign _340_ = inv_3[1] ^ r_2[22] /*18258*/;
  assign sum_3[1] = _340_ ^ _339_ /*18257*/;
  assign _341_ = _340_ & _339_ /*18256*/;
  assign _342_ = inv_3[1] & r_2[22] /*18255*/;
  assign _343_ = _341_ | _342_ /*18254*/;
  assign _344_ = inv_3[2] ^ r_2[23] /*18252*/;
  assign sum_3[2] = _344_ ^ _343_ /*18251*/;
  assign _345_ = _344_ & _343_ /*18250*/;
  assign _346_ = inv_3[2] & r_2[23] /*18249*/;
  assign _347_ = _345_ | _346_ /*18248*/;
  assign _348_ = inv_3[3] ^ r_2[24] /*18246*/;
  assign sum_3[3] = _348_ ^ _347_ /*18245*/;
  assign _349_ = _348_ & _347_ /*18244*/;
  assign _350_ = inv_3[3] & r_2[24] /*18243*/;
  assign _351_ = _349_ | _350_ /*18242*/;
  assign _352_ = inv_3[4] ^ r_2[25] /*18240*/;
  assign sum_3[4] = _352_ ^ _351_ /*18239*/;
  assign _353_ = _352_ & _351_ /*18238*/;
  assign _354_ = inv_3[4] & r_2[25] /*18237*/;
  assign _355_ = _353_ | _354_ /*18236*/;
  assign _356_ = inv_3[5] ^ r_2[26] /*18234*/;
  assign sum_3[5] = _356_ ^ _355_ /*18233*/;
  assign _357_ = _356_ & _355_ /*18232*/;
  assign _358_ = inv_3[5] & r_2[26] /*18231*/;
  assign _359_ = _357_ | _358_ /*18230*/;
  assign _360_ = inv_3[6] ^ r_2[27] /*18228*/;
  assign sum_3[6] = _360_ ^ _359_ /*18227*/;
  assign _361_ = _360_ & _359_ /*18226*/;
  assign _362_ = inv_3[6] & r_2[27] /*18225*/;
  assign _363_ = _361_ | _362_ /*18224*/;
  assign _364_ = inv_3[7] ^ r_2[28] /*18222*/;
  assign sum_3[7] = _364_ ^ _363_ /*18221*/;
  assign _365_ = _364_ & _363_ /*18220*/;
  assign _366_ = inv_3[7] & r_2[28] /*18219*/;
  assign _367_ = _365_ | _366_ /*18218*/;
  assign _368_ = inv_3[8] ^ r_2[29] /*18216*/;
  assign sum_3[8] = _368_ ^ _367_ /*18215*/;
  assign _369_ = _368_ & _367_ /*18214*/;
  assign _370_ = inv_3[8] & r_2[29] /*18213*/;
  assign _371_ = _369_ | _370_ /*18212*/;
  assign _372_ = inv_3[9] ^ r_2[30] /*18210*/;
  assign sum_3[9] = _372_ ^ _371_ /*18209*/;
  assign _373_ = _372_ & _371_ /*18208*/;
  assign _374_ = inv_3[9] & r_2[30] /*18207*/;
  assign _375_ = _373_ | _374_ /*18206*/;
  assign _376_ = inv_3[10] ^ r_2[31] /*18204*/;
  assign sum_3[10] = _376_ ^ _375_ /*18203*/;
  assign _377_ = _376_ & _375_ /*18202*/;
  assign _378_ = inv_3[10] & r_2[31] /*18201*/;
  assign _379_ = _377_ | _378_ /*18200*/;
  assign _380_ = inv_3[11] ^ r_2[32] /*18198*/;
  assign sum_3[11] = _380_ ^ _379_ /*18197*/;
  assign _381_ = _380_ & _379_ /*18196*/;
  assign _382_ = inv_3[11] & r_2[32] /*18195*/;
  assign _383_ = _381_ | _382_ /*18194*/;
  assign _384_ = inv_3[12] ^ r_2[33] /*18192*/;
  assign sum_3[12] = _384_ ^ _383_ /*18191*/;
  assign _385_ = _384_ & _383_ /*18190*/;
  assign _386_ = inv_3[12] & r_2[33] /*18189*/;
  assign _387_ = _385_ | _386_ /*18188*/;
  assign _388_ = inv_3[13] ^ r_2[34] /*18186*/;
  assign sum_3[13] = _388_ ^ _387_ /*18185*/;
  assign _389_ = _388_ & _387_ /*18184*/;
  assign _390_ = inv_3[13] & r_2[34] /*18183*/;
  assign _391_ = _389_ | _390_ /*18182*/;
  assign _392_ = inv_3[14] ^ r_2[35] /*18180*/;
  assign sum_3[14] = _392_ ^ _391_ /*18179*/;
  assign _393_ = _392_ & _391_ /*18178*/;
  assign _394_ = inv_3[14] & r_2[35] /*18177*/;
  assign _395_ = _393_ | _394_ /*18176*/;
  assign _396_ = inv_3[15] ^ r_2[36] /*18174*/;
  assign sum_3[15] = _396_ ^ _395_ /*18173*/;
  assign _397_ = _396_ & _395_ /*18172*/;
  assign _398_ = inv_3[15] & r_2[36] /*18171*/;
  assign _399_ = _397_ | _398_ /*18170*/;
  assign _400_ = inv_3[16] ^ r_2[37] /*18168*/;
  assign sum_3[16] = _400_ ^ _399_ /*18167*/;
  assign _401_ = _400_ & _399_ /*18166*/;
  assign _402_ = inv_3[16] & r_2[37] /*18165*/;
  assign _403_ = _401_ | _402_ /*18164*/;
  assign _404_ = inv_3[17] ^ r_2[38] /*18162*/;
  assign sum_3[17] = _404_ ^ _403_ /*18161*/;
  assign _405_ = _404_ & _403_ /*18160*/;
  assign _406_ = inv_3[17] & r_2[38] /*18159*/;
  assign _407_ = _405_ | _406_ /*18158*/;
  assign _408_ = inv_3[18] ^ r_2[39] /*18156*/;
  assign sum_3[18] = _408_ ^ _407_ /*18155*/;
  assign _409_ = _408_ & _407_ /*18154*/;
  assign _410_ = inv_3[18] & r_2[39] /*18153*/;
  assign _411_ = _409_ | _410_ /*18152*/;
  assign _412_ = inv_3[19] ^ r_2[40] /*18150*/;
  assign sum_3[19] = _412_ ^ _411_ /*18149*/;
  assign _413_ = _412_ & _411_ /*18148*/;
  assign _414_ = inv_3[19] & r_2[40] /*18147*/;
  assign _415_ = _413_ | _414_ /*18146*/;
  assign _416_ = inv_3[20] ^ r_2[41] /*18144*/;
  assign sum_3[20] = _416_ ^ _415_ /*18143*/;
  assign _417_ = _416_ & _415_ /*18142*/;
  assign _418_ = inv_3[20] & r_2[41] /*18141*/;
  assign _419_ = _417_ | _418_ /*18140*/;
  assign _420_ = inv_3[21] ^ r_2[42] /*18138*/;
  assign sum_3[21] = _420_ ^ _419_ /*18137*/;
  assign _421_ = _420_ & _419_ /*18136*/;
  assign _422_ = inv_3[21] & r_2[42] /*18135*/;
  assign _423_ = _421_ | _422_ /*18134*/;
  assign _424_ = inv_3[22] ^ r_2[43] /*18132*/;
  assign sum_3[22] = _424_ ^ _423_ /*18131*/;
  assign _425_ = _424_ & _423_ /*18130*/;
  assign _426_ = inv_3[22] & r_2[43] /*18129*/;
  assign _427_ = _425_ | _426_ /*18128*/;
  assign _428_ = inv_3[23] ^ r_2[44] /*18126*/;
  assign sum_3[23] = _428_ ^ _427_ /*18125*/;
  assign _429_ = _428_ & _427_ /*18124*/;
  assign _430_ = inv_3[23] & r_2[44] /*18123*/;
  assign _431_ = _429_ | _430_ /*18122*/;
  assign q[21] = ~sum_3[23] /*18141*/;
  assign m_3[0] = r_2[21] /*18140*/;
  assign m_3[1] = r_2[22] /*18139*/;
  assign m_3[2] = r_2[23] /*18138*/;
  assign m_3[3] = r_2[24] /*18137*/;
  assign m_3[4] = r_2[25] /*18136*/;
  assign m_3[5] = r_2[26] /*18135*/;
  assign m_3[6] = r_2[27] /*18134*/;
  assign m_3[7] = r_2[28] /*18133*/;
  assign m_3[8] = r_2[29] /*18132*/;
  assign m_3[9] = r_2[30] /*18131*/;
  assign m_3[10] = r_2[31] /*18130*/;
  assign m_3[11] = r_2[32] /*18129*/;
  assign m_3[12] = r_2[33] /*18128*/;
  assign m_3[13] = r_2[34] /*18127*/;
  assign m_3[14] = r_2[35] /*18126*/;
  assign m_3[15] = r_2[36] /*18125*/;
  assign m_3[16] = r_2[37] /*18124*/;
  assign m_3[17] = r_2[38] /*18123*/;
  assign m_3[18] = r_2[39] /*18122*/;
  assign m_3[19] = r_2[40] /*18121*/;
  assign m_3[20] = r_2[41] /*18120*/;
  assign m_3[21] = r_2[42] /*18119*/;
  assign m_3[22] = r_2[43] /*18118*/;
  assign m_3[23] = r_2[44] /*18117*/;
  assign _432_ = ~q[21] /*18115*/;
  assign _433_ = sum_3[0] & q[21] /*18114*/;
  assign _434_ = m_3[0] & _432_ /*18113*/;
  assign r_3[21] = _434_ | _433_ /*18112*/;
  assign _435_ = ~q[21] /*18111*/;
  assign _436_ = sum_3[1] & q[21] /*18110*/;
  assign _437_ = m_3[1] & _435_ /*18109*/;
  assign r_3[22] = _437_ | _436_ /*18108*/;
  assign _438_ = ~q[21] /*18107*/;
  assign _439_ = sum_3[2] & q[21] /*18106*/;
  assign _440_ = m_3[2] & _438_ /*18105*/;
  assign r_3[23] = _440_ | _439_ /*18104*/;
  assign _441_ = ~q[21] /*18103*/;
  assign _442_ = sum_3[3] & q[21] /*18102*/;
  assign _443_ = m_3[3] & _441_ /*18101*/;
  assign r_3[24] = _443_ | _442_ /*18100*/;
  assign _444_ = ~q[21] /*18099*/;
  assign _445_ = sum_3[4] & q[21] /*18098*/;
  assign _446_ = m_3[4] & _444_ /*18097*/;
  assign r_3[25] = _446_ | _445_ /*18096*/;
  assign _447_ = ~q[21] /*18095*/;
  assign _448_ = sum_3[5] & q[21] /*18094*/;
  assign _449_ = m_3[5] & _447_ /*18093*/;
  assign r_3[26] = _449_ | _448_ /*18092*/;
  assign _450_ = ~q[21] /*18091*/;
  assign _451_ = sum_3[6] & q[21] /*18090*/;
  assign _452_ = m_3[6] & _450_ /*18089*/;
  assign r_3[27] = _452_ | _451_ /*18088*/;
  assign _453_ = ~q[21] /*18087*/;
  assign _454_ = sum_3[7] & q[21] /*18086*/;
  assign _455_ = m_3[7] & _453_ /*18085*/;
  assign r_3[28] = _455_ | _454_ /*18084*/;
  assign _456_ = ~q[21] /*18083*/;
  assign _457_ = sum_3[8] & q[21] /*18082*/;
  assign _458_ = m_3[8] & _456_ /*18081*/;
  assign r_3[29] = _458_ | _457_ /*18080*/;
  assign _459_ = ~q[21] /*18079*/;
  assign _460_ = sum_3[9] & q[21] /*18078*/;
  assign _461_ = m_3[9] & _459_ /*18077*/;
  assign r_3[30] = _461_ | _460_ /*18076*/;
  assign _462_ = ~q[21] /*18075*/;
  assign _463_ = sum_3[10] & q[21] /*18074*/;
  assign _464_ = m_3[10] & _462_ /*18073*/;
  assign r_3[31] = _464_ | _463_ /*18072*/;
  assign _465_ = ~q[21] /*18071*/;
  assign _466_ = sum_3[11] & q[21] /*18070*/;
  assign _467_ = m_3[11] & _465_ /*18069*/;
  assign r_3[32] = _467_ | _466_ /*18068*/;
  assign _468_ = ~q[21] /*18067*/;
  assign _469_ = sum_3[12] & q[21] /*18066*/;
  assign _470_ = m_3[12] & _468_ /*18065*/;
  assign r_3[33] = _470_ | _469_ /*18064*/;
  assign _471_ = ~q[21] /*18063*/;
  assign _472_ = sum_3[13] & q[21] /*18062*/;
  assign _473_ = m_3[13] & _471_ /*18061*/;
  assign r_3[34] = _473_ | _472_ /*18060*/;
  assign _474_ = ~q[21] /*18059*/;
  assign _475_ = sum_3[14] & q[21] /*18058*/;
  assign _476_ = m_3[14] & _474_ /*18057*/;
  assign r_3[35] = _476_ | _475_ /*18056*/;
  assign _477_ = ~q[21] /*18055*/;
  assign _478_ = sum_3[15] & q[21] /*18054*/;
  assign _479_ = m_3[15] & _477_ /*18053*/;
  assign r_3[36] = _479_ | _478_ /*18052*/;
  assign _480_ = ~q[21] /*18051*/;
  assign _481_ = sum_3[16] & q[21] /*18050*/;
  assign _482_ = m_3[16] & _480_ /*18049*/;
  assign r_3[37] = _482_ | _481_ /*18048*/;
  assign _483_ = ~q[21] /*18047*/;
  assign _484_ = sum_3[17] & q[21] /*18046*/;
  assign _485_ = m_3[17] & _483_ /*18045*/;
  assign r_3[38] = _485_ | _484_ /*18044*/;
  assign _486_ = ~q[21] /*18043*/;
  assign _487_ = sum_3[18] & q[21] /*18042*/;
  assign _488_ = m_3[18] & _486_ /*18041*/;
  assign r_3[39] = _488_ | _487_ /*18040*/;
  assign _489_ = ~q[21] /*18039*/;
  assign _490_ = sum_3[19] & q[21] /*18038*/;
  assign _491_ = m_3[19] & _489_ /*18037*/;
  assign r_3[40] = _491_ | _490_ /*18036*/;
  assign _492_ = ~q[21] /*18035*/;
  assign _493_ = sum_3[20] & q[21] /*18034*/;
  assign _494_ = m_3[20] & _492_ /*18033*/;
  assign r_3[41] = _494_ | _493_ /*18032*/;
  assign _495_ = ~q[21] /*18031*/;
  assign _496_ = sum_3[21] & q[21] /*18030*/;
  assign _497_ = m_3[21] & _495_ /*18029*/;
  assign r_3[42] = _497_ | _496_ /*18028*/;
  assign _498_ = ~q[21] /*18027*/;
  assign _499_ = sum_3[22] & q[21] /*18026*/;
  assign _500_ = m_3[22] & _498_ /*18025*/;
  assign r_3[43] = _500_ | _499_ /*18024*/;
  assign _501_ = ~q[21] /*18023*/;
  assign _502_ = sum_3[23] & q[21] /*18022*/;
  assign _503_ = m_3[23] & _501_ /*18021*/;
  assign r_3[44] = _503_ | _502_ /*18020*/;
assign r_3[0]= r_2[0] /*18019*/;
assign r_3[1]= r_2[1] /*18018*/;
assign r_3[2]= r_2[2] /*18017*/;
assign r_3[3]= r_2[3] /*18016*/;
assign r_3[4]= r_2[4] /*18015*/;
assign r_3[5]= r_2[5] /*18014*/;
assign r_3[6]= r_2[6] /*18013*/;
assign r_3[7]= r_2[7] /*18012*/;
assign r_3[8]= r_2[8] /*18011*/;
assign r_3[9]= r_2[9] /*18010*/;
assign r_3[10]= r_2[10] /*18009*/;
assign r_3[11]= r_2[11] /*18008*/;
assign r_3[12]= r_2[12] /*18007*/;
assign r_3[13]= r_2[13] /*18006*/;
assign r_3[14]= r_2[14] /*18005*/;
assign r_3[15]= r_2[15] /*18004*/;
assign r_3[16]= r_2[16] /*18003*/;
assign r_3[17]= r_2[17] /*18002*/;
assign r_3[18]= r_2[18] /*18001*/;
assign r_3[19]= r_2[19] /*18000*/;
assign r_3[20]= r_2[20] /*17999*/;
  assign inv_4[0] = ~div[0] /*17952*/;
  assign inv_4[1] = ~div[1] /*17951*/;
  assign inv_4[2] = ~div[2] /*17950*/;
  assign inv_4[3] = ~div[3] /*17949*/;
  assign inv_4[4] = ~div[4] /*17948*/;
  assign inv_4[5] = ~div[5] /*17947*/;
  assign inv_4[6] = ~div[6] /*17946*/;
  assign inv_4[7] = ~div[7] /*17945*/;
  assign inv_4[8] = ~div[8] /*17944*/;
  assign inv_4[9] = ~div[9] /*17943*/;
  assign inv_4[10] = ~div[10] /*17942*/;
  assign inv_4[11] = ~div[11] /*17941*/;
  assign inv_4[12] = ~div[12] /*17940*/;
  assign inv_4[13] = ~div[13] /*17939*/;
  assign inv_4[14] = ~div[14] /*17938*/;
  assign inv_4[15] = ~div[15] /*17937*/;
  assign inv_4[16] = ~div[16] /*17936*/;
  assign inv_4[17] = ~div[17] /*17935*/;
  assign inv_4[18] = ~div[18] /*17934*/;
  assign inv_4[19] = ~div[19] /*17933*/;
  assign inv_4[20] = ~div[20] /*17932*/;
  assign inv_4[21] = ~div[21] /*17931*/;
  assign inv_4[22] = ~div[22] /*17930*/;
assign inv_4[23] = oneWire /*17929*/;
  assign _504_ = inv_4[0] ^ r_3[20] /*17927*/;
  assign sum_4[0] = _504_ ^ oneWire /*17926*/;
  assign _505_ = _504_ & oneWire /*17925*/;
  assign _506_ = inv_4[0] & r_3[20] /*17924*/;
  assign _507_ = _505_ | _506_ /*17923*/;
  assign _508_ = inv_4[1] ^ r_3[21] /*17922*/;
  assign sum_4[1] = _508_ ^ _507_ /*17921*/;
  assign _509_ = _508_ & _507_ /*17920*/;
  assign _510_ = inv_4[1] & r_3[21] /*17919*/;
  assign _511_ = _509_ | _510_ /*17918*/;
  assign _512_ = inv_4[2] ^ r_3[22] /*17916*/;
  assign sum_4[2] = _512_ ^ _511_ /*17915*/;
  assign _513_ = _512_ & _511_ /*17914*/;
  assign _514_ = inv_4[2] & r_3[22] /*17913*/;
  assign _515_ = _513_ | _514_ /*17912*/;
  assign _516_ = inv_4[3] ^ r_3[23] /*17910*/;
  assign sum_4[3] = _516_ ^ _515_ /*17909*/;
  assign _517_ = _516_ & _515_ /*17908*/;
  assign _518_ = inv_4[3] & r_3[23] /*17907*/;
  assign _519_ = _517_ | _518_ /*17906*/;
  assign _520_ = inv_4[4] ^ r_3[24] /*17904*/;
  assign sum_4[4] = _520_ ^ _519_ /*17903*/;
  assign _521_ = _520_ & _519_ /*17902*/;
  assign _522_ = inv_4[4] & r_3[24] /*17901*/;
  assign _523_ = _521_ | _522_ /*17900*/;
  assign _524_ = inv_4[5] ^ r_3[25] /*17898*/;
  assign sum_4[5] = _524_ ^ _523_ /*17897*/;
  assign _525_ = _524_ & _523_ /*17896*/;
  assign _526_ = inv_4[5] & r_3[25] /*17895*/;
  assign _527_ = _525_ | _526_ /*17894*/;
  assign _528_ = inv_4[6] ^ r_3[26] /*17892*/;
  assign sum_4[6] = _528_ ^ _527_ /*17891*/;
  assign _529_ = _528_ & _527_ /*17890*/;
  assign _530_ = inv_4[6] & r_3[26] /*17889*/;
  assign _531_ = _529_ | _530_ /*17888*/;
  assign _532_ = inv_4[7] ^ r_3[27] /*17886*/;
  assign sum_4[7] = _532_ ^ _531_ /*17885*/;
  assign _533_ = _532_ & _531_ /*17884*/;
  assign _534_ = inv_4[7] & r_3[27] /*17883*/;
  assign _535_ = _533_ | _534_ /*17882*/;
  assign _536_ = inv_4[8] ^ r_3[28] /*17880*/;
  assign sum_4[8] = _536_ ^ _535_ /*17879*/;
  assign _537_ = _536_ & _535_ /*17878*/;
  assign _538_ = inv_4[8] & r_3[28] /*17877*/;
  assign _539_ = _537_ | _538_ /*17876*/;
  assign _540_ = inv_4[9] ^ r_3[29] /*17874*/;
  assign sum_4[9] = _540_ ^ _539_ /*17873*/;
  assign _541_ = _540_ & _539_ /*17872*/;
  assign _542_ = inv_4[9] & r_3[29] /*17871*/;
  assign _543_ = _541_ | _542_ /*17870*/;
  assign _544_ = inv_4[10] ^ r_3[30] /*17868*/;
  assign sum_4[10] = _544_ ^ _543_ /*17867*/;
  assign _545_ = _544_ & _543_ /*17866*/;
  assign _546_ = inv_4[10] & r_3[30] /*17865*/;
  assign _547_ = _545_ | _546_ /*17864*/;
  assign _548_ = inv_4[11] ^ r_3[31] /*17862*/;
  assign sum_4[11] = _548_ ^ _547_ /*17861*/;
  assign _549_ = _548_ & _547_ /*17860*/;
  assign _550_ = inv_4[11] & r_3[31] /*17859*/;
  assign _551_ = _549_ | _550_ /*17858*/;
  assign _552_ = inv_4[12] ^ r_3[32] /*17856*/;
  assign sum_4[12] = _552_ ^ _551_ /*17855*/;
  assign _553_ = _552_ & _551_ /*17854*/;
  assign _554_ = inv_4[12] & r_3[32] /*17853*/;
  assign _555_ = _553_ | _554_ /*17852*/;
  assign _556_ = inv_4[13] ^ r_3[33] /*17850*/;
  assign sum_4[13] = _556_ ^ _555_ /*17849*/;
  assign _557_ = _556_ & _555_ /*17848*/;
  assign _558_ = inv_4[13] & r_3[33] /*17847*/;
  assign _559_ = _557_ | _558_ /*17846*/;
  assign _560_ = inv_4[14] ^ r_3[34] /*17844*/;
  assign sum_4[14] = _560_ ^ _559_ /*17843*/;
  assign _561_ = _560_ & _559_ /*17842*/;
  assign _562_ = inv_4[14] & r_3[34] /*17841*/;
  assign _563_ = _561_ | _562_ /*17840*/;
  assign _564_ = inv_4[15] ^ r_3[35] /*17838*/;
  assign sum_4[15] = _564_ ^ _563_ /*17837*/;
  assign _565_ = _564_ & _563_ /*17836*/;
  assign _566_ = inv_4[15] & r_3[35] /*17835*/;
  assign _567_ = _565_ | _566_ /*17834*/;
  assign _568_ = inv_4[16] ^ r_3[36] /*17832*/;
  assign sum_4[16] = _568_ ^ _567_ /*17831*/;
  assign _569_ = _568_ & _567_ /*17830*/;
  assign _570_ = inv_4[16] & r_3[36] /*17829*/;
  assign _571_ = _569_ | _570_ /*17828*/;
  assign _572_ = inv_4[17] ^ r_3[37] /*17826*/;
  assign sum_4[17] = _572_ ^ _571_ /*17825*/;
  assign _573_ = _572_ & _571_ /*17824*/;
  assign _574_ = inv_4[17] & r_3[37] /*17823*/;
  assign _575_ = _573_ | _574_ /*17822*/;
  assign _576_ = inv_4[18] ^ r_3[38] /*17820*/;
  assign sum_4[18] = _576_ ^ _575_ /*17819*/;
  assign _577_ = _576_ & _575_ /*17818*/;
  assign _578_ = inv_4[18] & r_3[38] /*17817*/;
  assign _579_ = _577_ | _578_ /*17816*/;
  assign _580_ = inv_4[19] ^ r_3[39] /*17814*/;
  assign sum_4[19] = _580_ ^ _579_ /*17813*/;
  assign _581_ = _580_ & _579_ /*17812*/;
  assign _582_ = inv_4[19] & r_3[39] /*17811*/;
  assign _583_ = _581_ | _582_ /*17810*/;
  assign _584_ = inv_4[20] ^ r_3[40] /*17808*/;
  assign sum_4[20] = _584_ ^ _583_ /*17807*/;
  assign _585_ = _584_ & _583_ /*17806*/;
  assign _586_ = inv_4[20] & r_3[40] /*17805*/;
  assign _587_ = _585_ | _586_ /*17804*/;
  assign _588_ = inv_4[21] ^ r_3[41] /*17802*/;
  assign sum_4[21] = _588_ ^ _587_ /*17801*/;
  assign _589_ = _588_ & _587_ /*17800*/;
  assign _590_ = inv_4[21] & r_3[41] /*17799*/;
  assign _591_ = _589_ | _590_ /*17798*/;
  assign _592_ = inv_4[22] ^ r_3[42] /*17796*/;
  assign sum_4[22] = _592_ ^ _591_ /*17795*/;
  assign _593_ = _592_ & _591_ /*17794*/;
  assign _594_ = inv_4[22] & r_3[42] /*17793*/;
  assign _595_ = _593_ | _594_ /*17792*/;
  assign _596_ = inv_4[23] ^ r_3[43] /*17790*/;
  assign sum_4[23] = _596_ ^ _595_ /*17789*/;
  assign _597_ = _596_ & _595_ /*17788*/;
  assign _598_ = inv_4[23] & r_3[43] /*17787*/;
  assign _599_ = _597_ | _598_ /*17786*/;
  assign q[20] = ~sum_4[23] /*17805*/;
  assign m_4[0] = r_3[20] /*17804*/;
  assign m_4[1] = r_3[21] /*17803*/;
  assign m_4[2] = r_3[22] /*17802*/;
  assign m_4[3] = r_3[23] /*17801*/;
  assign m_4[4] = r_3[24] /*17800*/;
  assign m_4[5] = r_3[25] /*17799*/;
  assign m_4[6] = r_3[26] /*17798*/;
  assign m_4[7] = r_3[27] /*17797*/;
  assign m_4[8] = r_3[28] /*17796*/;
  assign m_4[9] = r_3[29] /*17795*/;
  assign m_4[10] = r_3[30] /*17794*/;
  assign m_4[11] = r_3[31] /*17793*/;
  assign m_4[12] = r_3[32] /*17792*/;
  assign m_4[13] = r_3[33] /*17791*/;
  assign m_4[14] = r_3[34] /*17790*/;
  assign m_4[15] = r_3[35] /*17789*/;
  assign m_4[16] = r_3[36] /*17788*/;
  assign m_4[17] = r_3[37] /*17787*/;
  assign m_4[18] = r_3[38] /*17786*/;
  assign m_4[19] = r_3[39] /*17785*/;
  assign m_4[20] = r_3[40] /*17784*/;
  assign m_4[21] = r_3[41] /*17783*/;
  assign m_4[22] = r_3[42] /*17782*/;
  assign m_4[23] = r_3[43] /*17781*/;
  assign _600_ = ~q[20] /*17779*/;
  assign _601_ = sum_4[0] & q[20] /*17778*/;
  assign _602_ = m_4[0] & _600_ /*17777*/;
  assign r_4[20] = _602_ | _601_ /*17776*/;
  assign _603_ = ~q[20] /*17775*/;
  assign _604_ = sum_4[1] & q[20] /*17774*/;
  assign _605_ = m_4[1] & _603_ /*17773*/;
  assign r_4[21] = _605_ | _604_ /*17772*/;
  assign _606_ = ~q[20] /*17771*/;
  assign _607_ = sum_4[2] & q[20] /*17770*/;
  assign _608_ = m_4[2] & _606_ /*17769*/;
  assign r_4[22] = _608_ | _607_ /*17768*/;
  assign _609_ = ~q[20] /*17767*/;
  assign _610_ = sum_4[3] & q[20] /*17766*/;
  assign _611_ = m_4[3] & _609_ /*17765*/;
  assign r_4[23] = _611_ | _610_ /*17764*/;
  assign _612_ = ~q[20] /*17763*/;
  assign _613_ = sum_4[4] & q[20] /*17762*/;
  assign _614_ = m_4[4] & _612_ /*17761*/;
  assign r_4[24] = _614_ | _613_ /*17760*/;
  assign _615_ = ~q[20] /*17759*/;
  assign _616_ = sum_4[5] & q[20] /*17758*/;
  assign _617_ = m_4[5] & _615_ /*17757*/;
  assign r_4[25] = _617_ | _616_ /*17756*/;
  assign _618_ = ~q[20] /*17755*/;
  assign _619_ = sum_4[6] & q[20] /*17754*/;
  assign _620_ = m_4[6] & _618_ /*17753*/;
  assign r_4[26] = _620_ | _619_ /*17752*/;
  assign _621_ = ~q[20] /*17751*/;
  assign _622_ = sum_4[7] & q[20] /*17750*/;
  assign _623_ = m_4[7] & _621_ /*17749*/;
  assign r_4[27] = _623_ | _622_ /*17748*/;
  assign _624_ = ~q[20] /*17747*/;
  assign _625_ = sum_4[8] & q[20] /*17746*/;
  assign _626_ = m_4[8] & _624_ /*17745*/;
  assign r_4[28] = _626_ | _625_ /*17744*/;
  assign _627_ = ~q[20] /*17743*/;
  assign _628_ = sum_4[9] & q[20] /*17742*/;
  assign _629_ = m_4[9] & _627_ /*17741*/;
  assign r_4[29] = _629_ | _628_ /*17740*/;
  assign _630_ = ~q[20] /*17739*/;
  assign _631_ = sum_4[10] & q[20] /*17738*/;
  assign _632_ = m_4[10] & _630_ /*17737*/;
  assign r_4[30] = _632_ | _631_ /*17736*/;
  assign _633_ = ~q[20] /*17735*/;
  assign _634_ = sum_4[11] & q[20] /*17734*/;
  assign _635_ = m_4[11] & _633_ /*17733*/;
  assign r_4[31] = _635_ | _634_ /*17732*/;
  assign _636_ = ~q[20] /*17731*/;
  assign _637_ = sum_4[12] & q[20] /*17730*/;
  assign _638_ = m_4[12] & _636_ /*17729*/;
  assign r_4[32] = _638_ | _637_ /*17728*/;
  assign _639_ = ~q[20] /*17727*/;
  assign _640_ = sum_4[13] & q[20] /*17726*/;
  assign _641_ = m_4[13] & _639_ /*17725*/;
  assign r_4[33] = _641_ | _640_ /*17724*/;
  assign _642_ = ~q[20] /*17723*/;
  assign _643_ = sum_4[14] & q[20] /*17722*/;
  assign _644_ = m_4[14] & _642_ /*17721*/;
  assign r_4[34] = _644_ | _643_ /*17720*/;
  assign _645_ = ~q[20] /*17719*/;
  assign _646_ = sum_4[15] & q[20] /*17718*/;
  assign _647_ = m_4[15] & _645_ /*17717*/;
  assign r_4[35] = _647_ | _646_ /*17716*/;
  assign _648_ = ~q[20] /*17715*/;
  assign _649_ = sum_4[16] & q[20] /*17714*/;
  assign _650_ = m_4[16] & _648_ /*17713*/;
  assign r_4[36] = _650_ | _649_ /*17712*/;
  assign _651_ = ~q[20] /*17711*/;
  assign _652_ = sum_4[17] & q[20] /*17710*/;
  assign _653_ = m_4[17] & _651_ /*17709*/;
  assign r_4[37] = _653_ | _652_ /*17708*/;
  assign _654_ = ~q[20] /*17707*/;
  assign _655_ = sum_4[18] & q[20] /*17706*/;
  assign _656_ = m_4[18] & _654_ /*17705*/;
  assign r_4[38] = _656_ | _655_ /*17704*/;
  assign _657_ = ~q[20] /*17703*/;
  assign _658_ = sum_4[19] & q[20] /*17702*/;
  assign _659_ = m_4[19] & _657_ /*17701*/;
  assign r_4[39] = _659_ | _658_ /*17700*/;
  assign _660_ = ~q[20] /*17699*/;
  assign _661_ = sum_4[20] & q[20] /*17698*/;
  assign _662_ = m_4[20] & _660_ /*17697*/;
  assign r_4[40] = _662_ | _661_ /*17696*/;
  assign _663_ = ~q[20] /*17695*/;
  assign _664_ = sum_4[21] & q[20] /*17694*/;
  assign _665_ = m_4[21] & _663_ /*17693*/;
  assign r_4[41] = _665_ | _664_ /*17692*/;
  assign _666_ = ~q[20] /*17691*/;
  assign _667_ = sum_4[22] & q[20] /*17690*/;
  assign _668_ = m_4[22] & _666_ /*17689*/;
  assign r_4[42] = _668_ | _667_ /*17688*/;
  assign _669_ = ~q[20] /*17687*/;
  assign _670_ = sum_4[23] & q[20] /*17686*/;
  assign _671_ = m_4[23] & _669_ /*17685*/;
  assign r_4[43] = _671_ | _670_ /*17684*/;
assign r_4[0]= r_3[0] /*17683*/;
assign r_4[1]= r_3[1] /*17682*/;
assign r_4[2]= r_3[2] /*17681*/;
assign r_4[3]= r_3[3] /*17680*/;
assign r_4[4]= r_3[4] /*17679*/;
assign r_4[5]= r_3[5] /*17678*/;
assign r_4[6]= r_3[6] /*17677*/;
assign r_4[7]= r_3[7] /*17676*/;
assign r_4[8]= r_3[8] /*17675*/;
assign r_4[9]= r_3[9] /*17674*/;
assign r_4[10]= r_3[10] /*17673*/;
assign r_4[11]= r_3[11] /*17672*/;
assign r_4[12]= r_3[12] /*17671*/;
assign r_4[13]= r_3[13] /*17670*/;
assign r_4[14]= r_3[14] /*17669*/;
assign r_4[15]= r_3[15] /*17668*/;
assign r_4[16]= r_3[16] /*17667*/;
assign r_4[17]= r_3[17] /*17666*/;
assign r_4[18]= r_3[18] /*17665*/;
assign r_4[19]= r_3[19] /*17664*/;
  assign inv_5[0] = ~div[0] /*17616*/;
  assign inv_5[1] = ~div[1] /*17615*/;
  assign inv_5[2] = ~div[2] /*17614*/;
  assign inv_5[3] = ~div[3] /*17613*/;
  assign inv_5[4] = ~div[4] /*17612*/;
  assign inv_5[5] = ~div[5] /*17611*/;
  assign inv_5[6] = ~div[6] /*17610*/;
  assign inv_5[7] = ~div[7] /*17609*/;
  assign inv_5[8] = ~div[8] /*17608*/;
  assign inv_5[9] = ~div[9] /*17607*/;
  assign inv_5[10] = ~div[10] /*17606*/;
  assign inv_5[11] = ~div[11] /*17605*/;
  assign inv_5[12] = ~div[12] /*17604*/;
  assign inv_5[13] = ~div[13] /*17603*/;
  assign inv_5[14] = ~div[14] /*17602*/;
  assign inv_5[15] = ~div[15] /*17601*/;
  assign inv_5[16] = ~div[16] /*17600*/;
  assign inv_5[17] = ~div[17] /*17599*/;
  assign inv_5[18] = ~div[18] /*17598*/;
  assign inv_5[19] = ~div[19] /*17597*/;
  assign inv_5[20] = ~div[20] /*17596*/;
  assign inv_5[21] = ~div[21] /*17595*/;
  assign inv_5[22] = ~div[22] /*17594*/;
assign inv_5[23] = oneWire /*17593*/;
  assign _672_ = inv_5[0] ^ r_4[19] /*17591*/;
  assign sum_5[0] = _672_ ^ oneWire /*17590*/;
  assign _673_ = _672_ & oneWire /*17589*/;
  assign _674_ = inv_5[0] & r_4[19] /*17588*/;
  assign _675_ = _673_ | _674_ /*17587*/;
  assign _676_ = inv_5[1] ^ r_4[20] /*17586*/;
  assign sum_5[1] = _676_ ^ _675_ /*17585*/;
  assign _677_ = _676_ & _675_ /*17584*/;
  assign _678_ = inv_5[1] & r_4[20] /*17583*/;
  assign _679_ = _677_ | _678_ /*17582*/;
  assign _680_ = inv_5[2] ^ r_4[21] /*17580*/;
  assign sum_5[2] = _680_ ^ _679_ /*17579*/;
  assign _681_ = _680_ & _679_ /*17578*/;
  assign _682_ = inv_5[2] & r_4[21] /*17577*/;
  assign _683_ = _681_ | _682_ /*17576*/;
  assign _684_ = inv_5[3] ^ r_4[22] /*17574*/;
  assign sum_5[3] = _684_ ^ _683_ /*17573*/;
  assign _685_ = _684_ & _683_ /*17572*/;
  assign _686_ = inv_5[3] & r_4[22] /*17571*/;
  assign _687_ = _685_ | _686_ /*17570*/;
  assign _688_ = inv_5[4] ^ r_4[23] /*17568*/;
  assign sum_5[4] = _688_ ^ _687_ /*17567*/;
  assign _689_ = _688_ & _687_ /*17566*/;
  assign _690_ = inv_5[4] & r_4[23] /*17565*/;
  assign _691_ = _689_ | _690_ /*17564*/;
  assign _692_ = inv_5[5] ^ r_4[24] /*17562*/;
  assign sum_5[5] = _692_ ^ _691_ /*17561*/;
  assign _693_ = _692_ & _691_ /*17560*/;
  assign _694_ = inv_5[5] & r_4[24] /*17559*/;
  assign _695_ = _693_ | _694_ /*17558*/;
  assign _696_ = inv_5[6] ^ r_4[25] /*17556*/;
  assign sum_5[6] = _696_ ^ _695_ /*17555*/;
  assign _697_ = _696_ & _695_ /*17554*/;
  assign _698_ = inv_5[6] & r_4[25] /*17553*/;
  assign _699_ = _697_ | _698_ /*17552*/;
  assign _700_ = inv_5[7] ^ r_4[26] /*17550*/;
  assign sum_5[7] = _700_ ^ _699_ /*17549*/;
  assign _701_ = _700_ & _699_ /*17548*/;
  assign _702_ = inv_5[7] & r_4[26] /*17547*/;
  assign _703_ = _701_ | _702_ /*17546*/;
  assign _704_ = inv_5[8] ^ r_4[27] /*17544*/;
  assign sum_5[8] = _704_ ^ _703_ /*17543*/;
  assign _705_ = _704_ & _703_ /*17542*/;
  assign _706_ = inv_5[8] & r_4[27] /*17541*/;
  assign _707_ = _705_ | _706_ /*17540*/;
  assign _708_ = inv_5[9] ^ r_4[28] /*17538*/;
  assign sum_5[9] = _708_ ^ _707_ /*17537*/;
  assign _709_ = _708_ & _707_ /*17536*/;
  assign _710_ = inv_5[9] & r_4[28] /*17535*/;
  assign _711_ = _709_ | _710_ /*17534*/;
  assign _712_ = inv_5[10] ^ r_4[29] /*17532*/;
  assign sum_5[10] = _712_ ^ _711_ /*17531*/;
  assign _713_ = _712_ & _711_ /*17530*/;
  assign _714_ = inv_5[10] & r_4[29] /*17529*/;
  assign _715_ = _713_ | _714_ /*17528*/;
  assign _716_ = inv_5[11] ^ r_4[30] /*17526*/;
  assign sum_5[11] = _716_ ^ _715_ /*17525*/;
  assign _717_ = _716_ & _715_ /*17524*/;
  assign _718_ = inv_5[11] & r_4[30] /*17523*/;
  assign _719_ = _717_ | _718_ /*17522*/;
  assign _720_ = inv_5[12] ^ r_4[31] /*17520*/;
  assign sum_5[12] = _720_ ^ _719_ /*17519*/;
  assign _721_ = _720_ & _719_ /*17518*/;
  assign _722_ = inv_5[12] & r_4[31] /*17517*/;
  assign _723_ = _721_ | _722_ /*17516*/;
  assign _724_ = inv_5[13] ^ r_4[32] /*17514*/;
  assign sum_5[13] = _724_ ^ _723_ /*17513*/;
  assign _725_ = _724_ & _723_ /*17512*/;
  assign _726_ = inv_5[13] & r_4[32] /*17511*/;
  assign _727_ = _725_ | _726_ /*17510*/;
  assign _728_ = inv_5[14] ^ r_4[33] /*17508*/;
  assign sum_5[14] = _728_ ^ _727_ /*17507*/;
  assign _729_ = _728_ & _727_ /*17506*/;
  assign _730_ = inv_5[14] & r_4[33] /*17505*/;
  assign _731_ = _729_ | _730_ /*17504*/;
  assign _732_ = inv_5[15] ^ r_4[34] /*17502*/;
  assign sum_5[15] = _732_ ^ _731_ /*17501*/;
  assign _733_ = _732_ & _731_ /*17500*/;
  assign _734_ = inv_5[15] & r_4[34] /*17499*/;
  assign _735_ = _733_ | _734_ /*17498*/;
  assign _736_ = inv_5[16] ^ r_4[35] /*17496*/;
  assign sum_5[16] = _736_ ^ _735_ /*17495*/;
  assign _737_ = _736_ & _735_ /*17494*/;
  assign _738_ = inv_5[16] & r_4[35] /*17493*/;
  assign _739_ = _737_ | _738_ /*17492*/;
  assign _740_ = inv_5[17] ^ r_4[36] /*17490*/;
  assign sum_5[17] = _740_ ^ _739_ /*17489*/;
  assign _741_ = _740_ & _739_ /*17488*/;
  assign _742_ = inv_5[17] & r_4[36] /*17487*/;
  assign _743_ = _741_ | _742_ /*17486*/;
  assign _744_ = inv_5[18] ^ r_4[37] /*17484*/;
  assign sum_5[18] = _744_ ^ _743_ /*17483*/;
  assign _745_ = _744_ & _743_ /*17482*/;
  assign _746_ = inv_5[18] & r_4[37] /*17481*/;
  assign _747_ = _745_ | _746_ /*17480*/;
  assign _748_ = inv_5[19] ^ r_4[38] /*17478*/;
  assign sum_5[19] = _748_ ^ _747_ /*17477*/;
  assign _749_ = _748_ & _747_ /*17476*/;
  assign _750_ = inv_5[19] & r_4[38] /*17475*/;
  assign _751_ = _749_ | _750_ /*17474*/;
  assign _752_ = inv_5[20] ^ r_4[39] /*17472*/;
  assign sum_5[20] = _752_ ^ _751_ /*17471*/;
  assign _753_ = _752_ & _751_ /*17470*/;
  assign _754_ = inv_5[20] & r_4[39] /*17469*/;
  assign _755_ = _753_ | _754_ /*17468*/;
  assign _756_ = inv_5[21] ^ r_4[40] /*17466*/;
  assign sum_5[21] = _756_ ^ _755_ /*17465*/;
  assign _757_ = _756_ & _755_ /*17464*/;
  assign _758_ = inv_5[21] & r_4[40] /*17463*/;
  assign _759_ = _757_ | _758_ /*17462*/;
  assign _760_ = inv_5[22] ^ r_4[41] /*17460*/;
  assign sum_5[22] = _760_ ^ _759_ /*17459*/;
  assign _761_ = _760_ & _759_ /*17458*/;
  assign _762_ = inv_5[22] & r_4[41] /*17457*/;
  assign _763_ = _761_ | _762_ /*17456*/;
  assign _764_ = inv_5[23] ^ r_4[42] /*17454*/;
  assign sum_5[23] = _764_ ^ _763_ /*17453*/;
  assign _765_ = _764_ & _763_ /*17452*/;
  assign _766_ = inv_5[23] & r_4[42] /*17451*/;
  assign _767_ = _765_ | _766_ /*17450*/;
  assign q[19] = ~sum_5[23] /*17469*/;
  assign m_5[0] = r_4[19] /*17468*/;
  assign m_5[1] = r_4[20] /*17467*/;
  assign m_5[2] = r_4[21] /*17466*/;
  assign m_5[3] = r_4[22] /*17465*/;
  assign m_5[4] = r_4[23] /*17464*/;
  assign m_5[5] = r_4[24] /*17463*/;
  assign m_5[6] = r_4[25] /*17462*/;
  assign m_5[7] = r_4[26] /*17461*/;
  assign m_5[8] = r_4[27] /*17460*/;
  assign m_5[9] = r_4[28] /*17459*/;
  assign m_5[10] = r_4[29] /*17458*/;
  assign m_5[11] = r_4[30] /*17457*/;
  assign m_5[12] = r_4[31] /*17456*/;
  assign m_5[13] = r_4[32] /*17455*/;
  assign m_5[14] = r_4[33] /*17454*/;
  assign m_5[15] = r_4[34] /*17453*/;
  assign m_5[16] = r_4[35] /*17452*/;
  assign m_5[17] = r_4[36] /*17451*/;
  assign m_5[18] = r_4[37] /*17450*/;
  assign m_5[19] = r_4[38] /*17449*/;
  assign m_5[20] = r_4[39] /*17448*/;
  assign m_5[21] = r_4[40] /*17447*/;
  assign m_5[22] = r_4[41] /*17446*/;
  assign m_5[23] = r_4[42] /*17445*/;
  assign _768_ = ~q[19] /*17443*/;
  assign _769_ = sum_5[0] & q[19] /*17442*/;
  assign _770_ = m_5[0] & _768_ /*17441*/;
  assign r_5[19] = _770_ | _769_ /*17440*/;
  assign _771_ = ~q[19] /*17439*/;
  assign _772_ = sum_5[1] & q[19] /*17438*/;
  assign _773_ = m_5[1] & _771_ /*17437*/;
  assign r_5[20] = _773_ | _772_ /*17436*/;
  assign _774_ = ~q[19] /*17435*/;
  assign _775_ = sum_5[2] & q[19] /*17434*/;
  assign _776_ = m_5[2] & _774_ /*17433*/;
  assign r_5[21] = _776_ | _775_ /*17432*/;
  assign _777_ = ~q[19] /*17431*/;
  assign _778_ = sum_5[3] & q[19] /*17430*/;
  assign _779_ = m_5[3] & _777_ /*17429*/;
  assign r_5[22] = _779_ | _778_ /*17428*/;
  assign _780_ = ~q[19] /*17427*/;
  assign _781_ = sum_5[4] & q[19] /*17426*/;
  assign _782_ = m_5[4] & _780_ /*17425*/;
  assign r_5[23] = _782_ | _781_ /*17424*/;
  assign _783_ = ~q[19] /*17423*/;
  assign _784_ = sum_5[5] & q[19] /*17422*/;
  assign _785_ = m_5[5] & _783_ /*17421*/;
  assign r_5[24] = _785_ | _784_ /*17420*/;
  assign _786_ = ~q[19] /*17419*/;
  assign _787_ = sum_5[6] & q[19] /*17418*/;
  assign _788_ = m_5[6] & _786_ /*17417*/;
  assign r_5[25] = _788_ | _787_ /*17416*/;
  assign _789_ = ~q[19] /*17415*/;
  assign _790_ = sum_5[7] & q[19] /*17414*/;
  assign _791_ = m_5[7] & _789_ /*17413*/;
  assign r_5[26] = _791_ | _790_ /*17412*/;
  assign _792_ = ~q[19] /*17411*/;
  assign _793_ = sum_5[8] & q[19] /*17410*/;
  assign _794_ = m_5[8] & _792_ /*17409*/;
  assign r_5[27] = _794_ | _793_ /*17408*/;
  assign _795_ = ~q[19] /*17407*/;
  assign _796_ = sum_5[9] & q[19] /*17406*/;
  assign _797_ = m_5[9] & _795_ /*17405*/;
  assign r_5[28] = _797_ | _796_ /*17404*/;
  assign _798_ = ~q[19] /*17403*/;
  assign _799_ = sum_5[10] & q[19] /*17402*/;
  assign _800_ = m_5[10] & _798_ /*17401*/;
  assign r_5[29] = _800_ | _799_ /*17400*/;
  assign _801_ = ~q[19] /*17399*/;
  assign _802_ = sum_5[11] & q[19] /*17398*/;
  assign _803_ = m_5[11] & _801_ /*17397*/;
  assign r_5[30] = _803_ | _802_ /*17396*/;
  assign _804_ = ~q[19] /*17395*/;
  assign _805_ = sum_5[12] & q[19] /*17394*/;
  assign _806_ = m_5[12] & _804_ /*17393*/;
  assign r_5[31] = _806_ | _805_ /*17392*/;
  assign _807_ = ~q[19] /*17391*/;
  assign _808_ = sum_5[13] & q[19] /*17390*/;
  assign _809_ = m_5[13] & _807_ /*17389*/;
  assign r_5[32] = _809_ | _808_ /*17388*/;
  assign _810_ = ~q[19] /*17387*/;
  assign _811_ = sum_5[14] & q[19] /*17386*/;
  assign _812_ = m_5[14] & _810_ /*17385*/;
  assign r_5[33] = _812_ | _811_ /*17384*/;
  assign _813_ = ~q[19] /*17383*/;
  assign _814_ = sum_5[15] & q[19] /*17382*/;
  assign _815_ = m_5[15] & _813_ /*17381*/;
  assign r_5[34] = _815_ | _814_ /*17380*/;
  assign _816_ = ~q[19] /*17379*/;
  assign _817_ = sum_5[16] & q[19] /*17378*/;
  assign _818_ = m_5[16] & _816_ /*17377*/;
  assign r_5[35] = _818_ | _817_ /*17376*/;
  assign _819_ = ~q[19] /*17375*/;
  assign _820_ = sum_5[17] & q[19] /*17374*/;
  assign _821_ = m_5[17] & _819_ /*17373*/;
  assign r_5[36] = _821_ | _820_ /*17372*/;
  assign _822_ = ~q[19] /*17371*/;
  assign _823_ = sum_5[18] & q[19] /*17370*/;
  assign _824_ = m_5[18] & _822_ /*17369*/;
  assign r_5[37] = _824_ | _823_ /*17368*/;
  assign _825_ = ~q[19] /*17367*/;
  assign _826_ = sum_5[19] & q[19] /*17366*/;
  assign _827_ = m_5[19] & _825_ /*17365*/;
  assign r_5[38] = _827_ | _826_ /*17364*/;
  assign _828_ = ~q[19] /*17363*/;
  assign _829_ = sum_5[20] & q[19] /*17362*/;
  assign _830_ = m_5[20] & _828_ /*17361*/;
  assign r_5[39] = _830_ | _829_ /*17360*/;
  assign _831_ = ~q[19] /*17359*/;
  assign _832_ = sum_5[21] & q[19] /*17358*/;
  assign _833_ = m_5[21] & _831_ /*17357*/;
  assign r_5[40] = _833_ | _832_ /*17356*/;
  assign _834_ = ~q[19] /*17355*/;
  assign _835_ = sum_5[22] & q[19] /*17354*/;
  assign _836_ = m_5[22] & _834_ /*17353*/;
  assign r_5[41] = _836_ | _835_ /*17352*/;
  assign _837_ = ~q[19] /*17351*/;
  assign _838_ = sum_5[23] & q[19] /*17350*/;
  assign _839_ = m_5[23] & _837_ /*17349*/;
  assign r_5[42] = _839_ | _838_ /*17348*/;
assign r_5[0]= r_4[0] /*17347*/;
assign r_5[1]= r_4[1] /*17346*/;
assign r_5[2]= r_4[2] /*17345*/;
assign r_5[3]= r_4[3] /*17344*/;
assign r_5[4]= r_4[4] /*17343*/;
assign r_5[5]= r_4[5] /*17342*/;
assign r_5[6]= r_4[6] /*17341*/;
assign r_5[7]= r_4[7] /*17340*/;
assign r_5[8]= r_4[8] /*17339*/;
assign r_5[9]= r_4[9] /*17338*/;
assign r_5[10]= r_4[10] /*17337*/;
assign r_5[11]= r_4[11] /*17336*/;
assign r_5[12]= r_4[12] /*17335*/;
assign r_5[13]= r_4[13] /*17334*/;
assign r_5[14]= r_4[14] /*17333*/;
assign r_5[15]= r_4[15] /*17332*/;
assign r_5[16]= r_4[16] /*17331*/;
assign r_5[17]= r_4[17] /*17330*/;
assign r_5[18]= r_4[18] /*17329*/;
  assign inv_6[0] = ~div[0] /*17280*/;
  assign inv_6[1] = ~div[1] /*17279*/;
  assign inv_6[2] = ~div[2] /*17278*/;
  assign inv_6[3] = ~div[3] /*17277*/;
  assign inv_6[4] = ~div[4] /*17276*/;
  assign inv_6[5] = ~div[5] /*17275*/;
  assign inv_6[6] = ~div[6] /*17274*/;
  assign inv_6[7] = ~div[7] /*17273*/;
  assign inv_6[8] = ~div[8] /*17272*/;
  assign inv_6[9] = ~div[9] /*17271*/;
  assign inv_6[10] = ~div[10] /*17270*/;
  assign inv_6[11] = ~div[11] /*17269*/;
  assign inv_6[12] = ~div[12] /*17268*/;
  assign inv_6[13] = ~div[13] /*17267*/;
  assign inv_6[14] = ~div[14] /*17266*/;
  assign inv_6[15] = ~div[15] /*17265*/;
  assign inv_6[16] = ~div[16] /*17264*/;
  assign inv_6[17] = ~div[17] /*17263*/;
  assign inv_6[18] = ~div[18] /*17262*/;
  assign inv_6[19] = ~div[19] /*17261*/;
  assign inv_6[20] = ~div[20] /*17260*/;
  assign inv_6[21] = ~div[21] /*17259*/;
  assign inv_6[22] = ~div[22] /*17258*/;
assign inv_6[23] = oneWire /*17257*/;
  assign _840_ = inv_6[0] ^ r_5[18] /*17255*/;
  assign sum_6[0] = _840_ ^ oneWire /*17254*/;
  assign _841_ = _840_ & oneWire /*17253*/;
  assign _842_ = inv_6[0] & r_5[18] /*17252*/;
  assign _843_ = _841_ | _842_ /*17251*/;
  assign _844_ = inv_6[1] ^ r_5[19] /*17250*/;
  assign sum_6[1] = _844_ ^ _843_ /*17249*/;
  assign _845_ = _844_ & _843_ /*17248*/;
  assign _846_ = inv_6[1] & r_5[19] /*17247*/;
  assign _847_ = _845_ | _846_ /*17246*/;
  assign _848_ = inv_6[2] ^ r_5[20] /*17244*/;
  assign sum_6[2] = _848_ ^ _847_ /*17243*/;
  assign _849_ = _848_ & _847_ /*17242*/;
  assign _850_ = inv_6[2] & r_5[20] /*17241*/;
  assign _851_ = _849_ | _850_ /*17240*/;
  assign _852_ = inv_6[3] ^ r_5[21] /*17238*/;
  assign sum_6[3] = _852_ ^ _851_ /*17237*/;
  assign _853_ = _852_ & _851_ /*17236*/;
  assign _854_ = inv_6[3] & r_5[21] /*17235*/;
  assign _855_ = _853_ | _854_ /*17234*/;
  assign _856_ = inv_6[4] ^ r_5[22] /*17232*/;
  assign sum_6[4] = _856_ ^ _855_ /*17231*/;
  assign _857_ = _856_ & _855_ /*17230*/;
  assign _858_ = inv_6[4] & r_5[22] /*17229*/;
  assign _859_ = _857_ | _858_ /*17228*/;
  assign _860_ = inv_6[5] ^ r_5[23] /*17226*/;
  assign sum_6[5] = _860_ ^ _859_ /*17225*/;
  assign _861_ = _860_ & _859_ /*17224*/;
  assign _862_ = inv_6[5] & r_5[23] /*17223*/;
  assign _863_ = _861_ | _862_ /*17222*/;
  assign _864_ = inv_6[6] ^ r_5[24] /*17220*/;
  assign sum_6[6] = _864_ ^ _863_ /*17219*/;
  assign _865_ = _864_ & _863_ /*17218*/;
  assign _866_ = inv_6[6] & r_5[24] /*17217*/;
  assign _867_ = _865_ | _866_ /*17216*/;
  assign _868_ = inv_6[7] ^ r_5[25] /*17214*/;
  assign sum_6[7] = _868_ ^ _867_ /*17213*/;
  assign _869_ = _868_ & _867_ /*17212*/;
  assign _870_ = inv_6[7] & r_5[25] /*17211*/;
  assign _871_ = _869_ | _870_ /*17210*/;
  assign _872_ = inv_6[8] ^ r_5[26] /*17208*/;
  assign sum_6[8] = _872_ ^ _871_ /*17207*/;
  assign _873_ = _872_ & _871_ /*17206*/;
  assign _874_ = inv_6[8] & r_5[26] /*17205*/;
  assign _875_ = _873_ | _874_ /*17204*/;
  assign _876_ = inv_6[9] ^ r_5[27] /*17202*/;
  assign sum_6[9] = _876_ ^ _875_ /*17201*/;
  assign _877_ = _876_ & _875_ /*17200*/;
  assign _878_ = inv_6[9] & r_5[27] /*17199*/;
  assign _879_ = _877_ | _878_ /*17198*/;
  assign _880_ = inv_6[10] ^ r_5[28] /*17196*/;
  assign sum_6[10] = _880_ ^ _879_ /*17195*/;
  assign _881_ = _880_ & _879_ /*17194*/;
  assign _882_ = inv_6[10] & r_5[28] /*17193*/;
  assign _883_ = _881_ | _882_ /*17192*/;
  assign _884_ = inv_6[11] ^ r_5[29] /*17190*/;
  assign sum_6[11] = _884_ ^ _883_ /*17189*/;
  assign _885_ = _884_ & _883_ /*17188*/;
  assign _886_ = inv_6[11] & r_5[29] /*17187*/;
  assign _887_ = _885_ | _886_ /*17186*/;
  assign _888_ = inv_6[12] ^ r_5[30] /*17184*/;
  assign sum_6[12] = _888_ ^ _887_ /*17183*/;
  assign _889_ = _888_ & _887_ /*17182*/;
  assign _890_ = inv_6[12] & r_5[30] /*17181*/;
  assign _891_ = _889_ | _890_ /*17180*/;
  assign _892_ = inv_6[13] ^ r_5[31] /*17178*/;
  assign sum_6[13] = _892_ ^ _891_ /*17177*/;
  assign _893_ = _892_ & _891_ /*17176*/;
  assign _894_ = inv_6[13] & r_5[31] /*17175*/;
  assign _895_ = _893_ | _894_ /*17174*/;
  assign _896_ = inv_6[14] ^ r_5[32] /*17172*/;
  assign sum_6[14] = _896_ ^ _895_ /*17171*/;
  assign _897_ = _896_ & _895_ /*17170*/;
  assign _898_ = inv_6[14] & r_5[32] /*17169*/;
  assign _899_ = _897_ | _898_ /*17168*/;
  assign _900_ = inv_6[15] ^ r_5[33] /*17166*/;
  assign sum_6[15] = _900_ ^ _899_ /*17165*/;
  assign _901_ = _900_ & _899_ /*17164*/;
  assign _902_ = inv_6[15] & r_5[33] /*17163*/;
  assign _903_ = _901_ | _902_ /*17162*/;
  assign _904_ = inv_6[16] ^ r_5[34] /*17160*/;
  assign sum_6[16] = _904_ ^ _903_ /*17159*/;
  assign _905_ = _904_ & _903_ /*17158*/;
  assign _906_ = inv_6[16] & r_5[34] /*17157*/;
  assign _907_ = _905_ | _906_ /*17156*/;
  assign _908_ = inv_6[17] ^ r_5[35] /*17154*/;
  assign sum_6[17] = _908_ ^ _907_ /*17153*/;
  assign _909_ = _908_ & _907_ /*17152*/;
  assign _910_ = inv_6[17] & r_5[35] /*17151*/;
  assign _911_ = _909_ | _910_ /*17150*/;
  assign _912_ = inv_6[18] ^ r_5[36] /*17148*/;
  assign sum_6[18] = _912_ ^ _911_ /*17147*/;
  assign _913_ = _912_ & _911_ /*17146*/;
  assign _914_ = inv_6[18] & r_5[36] /*17145*/;
  assign _915_ = _913_ | _914_ /*17144*/;
  assign _916_ = inv_6[19] ^ r_5[37] /*17142*/;
  assign sum_6[19] = _916_ ^ _915_ /*17141*/;
  assign _917_ = _916_ & _915_ /*17140*/;
  assign _918_ = inv_6[19] & r_5[37] /*17139*/;
  assign _919_ = _917_ | _918_ /*17138*/;
  assign _920_ = inv_6[20] ^ r_5[38] /*17136*/;
  assign sum_6[20] = _920_ ^ _919_ /*17135*/;
  assign _921_ = _920_ & _919_ /*17134*/;
  assign _922_ = inv_6[20] & r_5[38] /*17133*/;
  assign _923_ = _921_ | _922_ /*17132*/;
  assign _924_ = inv_6[21] ^ r_5[39] /*17130*/;
  assign sum_6[21] = _924_ ^ _923_ /*17129*/;
  assign _925_ = _924_ & _923_ /*17128*/;
  assign _926_ = inv_6[21] & r_5[39] /*17127*/;
  assign _927_ = _925_ | _926_ /*17126*/;
  assign _928_ = inv_6[22] ^ r_5[40] /*17124*/;
  assign sum_6[22] = _928_ ^ _927_ /*17123*/;
  assign _929_ = _928_ & _927_ /*17122*/;
  assign _930_ = inv_6[22] & r_5[40] /*17121*/;
  assign _931_ = _929_ | _930_ /*17120*/;
  assign _932_ = inv_6[23] ^ r_5[41] /*17118*/;
  assign sum_6[23] = _932_ ^ _931_ /*17117*/;
  assign _933_ = _932_ & _931_ /*17116*/;
  assign _934_ = inv_6[23] & r_5[41] /*17115*/;
  assign _935_ = _933_ | _934_ /*17114*/;
  assign q[18] = ~sum_6[23] /*17133*/;
  assign m_6[0] = r_5[18] /*17132*/;
  assign m_6[1] = r_5[19] /*17131*/;
  assign m_6[2] = r_5[20] /*17130*/;
  assign m_6[3] = r_5[21] /*17129*/;
  assign m_6[4] = r_5[22] /*17128*/;
  assign m_6[5] = r_5[23] /*17127*/;
  assign m_6[6] = r_5[24] /*17126*/;
  assign m_6[7] = r_5[25] /*17125*/;
  assign m_6[8] = r_5[26] /*17124*/;
  assign m_6[9] = r_5[27] /*17123*/;
  assign m_6[10] = r_5[28] /*17122*/;
  assign m_6[11] = r_5[29] /*17121*/;
  assign m_6[12] = r_5[30] /*17120*/;
  assign m_6[13] = r_5[31] /*17119*/;
  assign m_6[14] = r_5[32] /*17118*/;
  assign m_6[15] = r_5[33] /*17117*/;
  assign m_6[16] = r_5[34] /*17116*/;
  assign m_6[17] = r_5[35] /*17115*/;
  assign m_6[18] = r_5[36] /*17114*/;
  assign m_6[19] = r_5[37] /*17113*/;
  assign m_6[20] = r_5[38] /*17112*/;
  assign m_6[21] = r_5[39] /*17111*/;
  assign m_6[22] = r_5[40] /*17110*/;
  assign m_6[23] = r_5[41] /*17109*/;
  assign _936_ = ~q[18] /*17107*/;
  assign _937_ = sum_6[0] & q[18] /*17106*/;
  assign _938_ = m_6[0] & _936_ /*17105*/;
  assign r_6[18] = _938_ | _937_ /*17104*/;
  assign _939_ = ~q[18] /*17103*/;
  assign _940_ = sum_6[1] & q[18] /*17102*/;
  assign _941_ = m_6[1] & _939_ /*17101*/;
  assign r_6[19] = _941_ | _940_ /*17100*/;
  assign _942_ = ~q[18] /*17099*/;
  assign _943_ = sum_6[2] & q[18] /*17098*/;
  assign _944_ = m_6[2] & _942_ /*17097*/;
  assign r_6[20] = _944_ | _943_ /*17096*/;
  assign _945_ = ~q[18] /*17095*/;
  assign _946_ = sum_6[3] & q[18] /*17094*/;
  assign _947_ = m_6[3] & _945_ /*17093*/;
  assign r_6[21] = _947_ | _946_ /*17092*/;
  assign _948_ = ~q[18] /*17091*/;
  assign _949_ = sum_6[4] & q[18] /*17090*/;
  assign _950_ = m_6[4] & _948_ /*17089*/;
  assign r_6[22] = _950_ | _949_ /*17088*/;
  assign _951_ = ~q[18] /*17087*/;
  assign _952_ = sum_6[5] & q[18] /*17086*/;
  assign _953_ = m_6[5] & _951_ /*17085*/;
  assign r_6[23] = _953_ | _952_ /*17084*/;
  assign _954_ = ~q[18] /*17083*/;
  assign _955_ = sum_6[6] & q[18] /*17082*/;
  assign _956_ = m_6[6] & _954_ /*17081*/;
  assign r_6[24] = _956_ | _955_ /*17080*/;
  assign _957_ = ~q[18] /*17079*/;
  assign _958_ = sum_6[7] & q[18] /*17078*/;
  assign _959_ = m_6[7] & _957_ /*17077*/;
  assign r_6[25] = _959_ | _958_ /*17076*/;
  assign _960_ = ~q[18] /*17075*/;
  assign _961_ = sum_6[8] & q[18] /*17074*/;
  assign _962_ = m_6[8] & _960_ /*17073*/;
  assign r_6[26] = _962_ | _961_ /*17072*/;
  assign _963_ = ~q[18] /*17071*/;
  assign _964_ = sum_6[9] & q[18] /*17070*/;
  assign _965_ = m_6[9] & _963_ /*17069*/;
  assign r_6[27] = _965_ | _964_ /*17068*/;
  assign _966_ = ~q[18] /*17067*/;
  assign _967_ = sum_6[10] & q[18] /*17066*/;
  assign _968_ = m_6[10] & _966_ /*17065*/;
  assign r_6[28] = _968_ | _967_ /*17064*/;
  assign _969_ = ~q[18] /*17063*/;
  assign _970_ = sum_6[11] & q[18] /*17062*/;
  assign _971_ = m_6[11] & _969_ /*17061*/;
  assign r_6[29] = _971_ | _970_ /*17060*/;
  assign _972_ = ~q[18] /*17059*/;
  assign _973_ = sum_6[12] & q[18] /*17058*/;
  assign _974_ = m_6[12] & _972_ /*17057*/;
  assign r_6[30] = _974_ | _973_ /*17056*/;
  assign _975_ = ~q[18] /*17055*/;
  assign _976_ = sum_6[13] & q[18] /*17054*/;
  assign _977_ = m_6[13] & _975_ /*17053*/;
  assign r_6[31] = _977_ | _976_ /*17052*/;
  assign _978_ = ~q[18] /*17051*/;
  assign _979_ = sum_6[14] & q[18] /*17050*/;
  assign _980_ = m_6[14] & _978_ /*17049*/;
  assign r_6[32] = _980_ | _979_ /*17048*/;
  assign _981_ = ~q[18] /*17047*/;
  assign _982_ = sum_6[15] & q[18] /*17046*/;
  assign _983_ = m_6[15] & _981_ /*17045*/;
  assign r_6[33] = _983_ | _982_ /*17044*/;
  assign _984_ = ~q[18] /*17043*/;
  assign _985_ = sum_6[16] & q[18] /*17042*/;
  assign _986_ = m_6[16] & _984_ /*17041*/;
  assign r_6[34] = _986_ | _985_ /*17040*/;
  assign _987_ = ~q[18] /*17039*/;
  assign _988_ = sum_6[17] & q[18] /*17038*/;
  assign _989_ = m_6[17] & _987_ /*17037*/;
  assign r_6[35] = _989_ | _988_ /*17036*/;
  assign _990_ = ~q[18] /*17035*/;
  assign _991_ = sum_6[18] & q[18] /*17034*/;
  assign _992_ = m_6[18] & _990_ /*17033*/;
  assign r_6[36] = _992_ | _991_ /*17032*/;
  assign _993_ = ~q[18] /*17031*/;
  assign _994_ = sum_6[19] & q[18] /*17030*/;
  assign _995_ = m_6[19] & _993_ /*17029*/;
  assign r_6[37] = _995_ | _994_ /*17028*/;
  assign _996_ = ~q[18] /*17027*/;
  assign _997_ = sum_6[20] & q[18] /*17026*/;
  assign _998_ = m_6[20] & _996_ /*17025*/;
  assign r_6[38] = _998_ | _997_ /*17024*/;
  assign _999_ = ~q[18] /*17023*/;
  assign _1000_ = sum_6[21] & q[18] /*17022*/;
  assign _1001_ = m_6[21] & _999_ /*17021*/;
  assign r_6[39] = _1001_ | _1000_ /*17020*/;
  assign _1002_ = ~q[18] /*17019*/;
  assign _1003_ = sum_6[22] & q[18] /*17018*/;
  assign _1004_ = m_6[22] & _1002_ /*17017*/;
  assign r_6[40] = _1004_ | _1003_ /*17016*/;
  assign _1005_ = ~q[18] /*17015*/;
  assign _1006_ = sum_6[23] & q[18] /*17014*/;
  assign _1007_ = m_6[23] & _1005_ /*17013*/;
  assign r_6[41] = _1007_ | _1006_ /*17012*/;
assign r_6[0]= r_5[0] /*17011*/;
assign r_6[1]= r_5[1] /*17010*/;
assign r_6[2]= r_5[2] /*17009*/;
assign r_6[3]= r_5[3] /*17008*/;
assign r_6[4]= r_5[4] /*17007*/;
assign r_6[5]= r_5[5] /*17006*/;
assign r_6[6]= r_5[6] /*17005*/;
assign r_6[7]= r_5[7] /*17004*/;
assign r_6[8]= r_5[8] /*17003*/;
assign r_6[9]= r_5[9] /*17002*/;
assign r_6[10]= r_5[10] /*17001*/;
assign r_6[11]= r_5[11] /*17000*/;
assign r_6[12]= r_5[12] /*16999*/;
assign r_6[13]= r_5[13] /*16998*/;
assign r_6[14]= r_5[14] /*16997*/;
assign r_6[15]= r_5[15] /*16996*/;
assign r_6[16]= r_5[16] /*16995*/;
assign r_6[17]= r_5[17] /*16994*/;
  assign inv_7[0] = ~div[0] /*16944*/;
  assign inv_7[1] = ~div[1] /*16943*/;
  assign inv_7[2] = ~div[2] /*16942*/;
  assign inv_7[3] = ~div[3] /*16941*/;
  assign inv_7[4] = ~div[4] /*16940*/;
  assign inv_7[5] = ~div[5] /*16939*/;
  assign inv_7[6] = ~div[6] /*16938*/;
  assign inv_7[7] = ~div[7] /*16937*/;
  assign inv_7[8] = ~div[8] /*16936*/;
  assign inv_7[9] = ~div[9] /*16935*/;
  assign inv_7[10] = ~div[10] /*16934*/;
  assign inv_7[11] = ~div[11] /*16933*/;
  assign inv_7[12] = ~div[12] /*16932*/;
  assign inv_7[13] = ~div[13] /*16931*/;
  assign inv_7[14] = ~div[14] /*16930*/;
  assign inv_7[15] = ~div[15] /*16929*/;
  assign inv_7[16] = ~div[16] /*16928*/;
  assign inv_7[17] = ~div[17] /*16927*/;
  assign inv_7[18] = ~div[18] /*16926*/;
  assign inv_7[19] = ~div[19] /*16925*/;
  assign inv_7[20] = ~div[20] /*16924*/;
  assign inv_7[21] = ~div[21] /*16923*/;
  assign inv_7[22] = ~div[22] /*16922*/;
assign inv_7[23] = oneWire /*16921*/;
  assign _1008_ = inv_7[0] ^ r_6[17] /*16919*/;
  assign sum_7[0] = _1008_ ^ oneWire /*16918*/;
  assign _1009_ = _1008_ & oneWire /*16917*/;
  assign _1010_ = inv_7[0] & r_6[17] /*16916*/;
  assign _1011_ = _1009_ | _1010_ /*16915*/;
  assign _1012_ = inv_7[1] ^ r_6[18] /*16914*/;
  assign sum_7[1] = _1012_ ^ _1011_ /*16913*/;
  assign _1013_ = _1012_ & _1011_ /*16912*/;
  assign _1014_ = inv_7[1] & r_6[18] /*16911*/;
  assign _1015_ = _1013_ | _1014_ /*16910*/;
  assign _1016_ = inv_7[2] ^ r_6[19] /*16908*/;
  assign sum_7[2] = _1016_ ^ _1015_ /*16907*/;
  assign _1017_ = _1016_ & _1015_ /*16906*/;
  assign _1018_ = inv_7[2] & r_6[19] /*16905*/;
  assign _1019_ = _1017_ | _1018_ /*16904*/;
  assign _1020_ = inv_7[3] ^ r_6[20] /*16902*/;
  assign sum_7[3] = _1020_ ^ _1019_ /*16901*/;
  assign _1021_ = _1020_ & _1019_ /*16900*/;
  assign _1022_ = inv_7[3] & r_6[20] /*16899*/;
  assign _1023_ = _1021_ | _1022_ /*16898*/;
  assign _1024_ = inv_7[4] ^ r_6[21] /*16896*/;
  assign sum_7[4] = _1024_ ^ _1023_ /*16895*/;
  assign _1025_ = _1024_ & _1023_ /*16894*/;
  assign _1026_ = inv_7[4] & r_6[21] /*16893*/;
  assign _1027_ = _1025_ | _1026_ /*16892*/;
  assign _1028_ = inv_7[5] ^ r_6[22] /*16890*/;
  assign sum_7[5] = _1028_ ^ _1027_ /*16889*/;
  assign _1029_ = _1028_ & _1027_ /*16888*/;
  assign _1030_ = inv_7[5] & r_6[22] /*16887*/;
  assign _1031_ = _1029_ | _1030_ /*16886*/;
  assign _1032_ = inv_7[6] ^ r_6[23] /*16884*/;
  assign sum_7[6] = _1032_ ^ _1031_ /*16883*/;
  assign _1033_ = _1032_ & _1031_ /*16882*/;
  assign _1034_ = inv_7[6] & r_6[23] /*16881*/;
  assign _1035_ = _1033_ | _1034_ /*16880*/;
  assign _1036_ = inv_7[7] ^ r_6[24] /*16878*/;
  assign sum_7[7] = _1036_ ^ _1035_ /*16877*/;
  assign _1037_ = _1036_ & _1035_ /*16876*/;
  assign _1038_ = inv_7[7] & r_6[24] /*16875*/;
  assign _1039_ = _1037_ | _1038_ /*16874*/;
  assign _1040_ = inv_7[8] ^ r_6[25] /*16872*/;
  assign sum_7[8] = _1040_ ^ _1039_ /*16871*/;
  assign _1041_ = _1040_ & _1039_ /*16870*/;
  assign _1042_ = inv_7[8] & r_6[25] /*16869*/;
  assign _1043_ = _1041_ | _1042_ /*16868*/;
  assign _1044_ = inv_7[9] ^ r_6[26] /*16866*/;
  assign sum_7[9] = _1044_ ^ _1043_ /*16865*/;
  assign _1045_ = _1044_ & _1043_ /*16864*/;
  assign _1046_ = inv_7[9] & r_6[26] /*16863*/;
  assign _1047_ = _1045_ | _1046_ /*16862*/;
  assign _1048_ = inv_7[10] ^ r_6[27] /*16860*/;
  assign sum_7[10] = _1048_ ^ _1047_ /*16859*/;
  assign _1049_ = _1048_ & _1047_ /*16858*/;
  assign _1050_ = inv_7[10] & r_6[27] /*16857*/;
  assign _1051_ = _1049_ | _1050_ /*16856*/;
  assign _1052_ = inv_7[11] ^ r_6[28] /*16854*/;
  assign sum_7[11] = _1052_ ^ _1051_ /*16853*/;
  assign _1053_ = _1052_ & _1051_ /*16852*/;
  assign _1054_ = inv_7[11] & r_6[28] /*16851*/;
  assign _1055_ = _1053_ | _1054_ /*16850*/;
  assign _1056_ = inv_7[12] ^ r_6[29] /*16848*/;
  assign sum_7[12] = _1056_ ^ _1055_ /*16847*/;
  assign _1057_ = _1056_ & _1055_ /*16846*/;
  assign _1058_ = inv_7[12] & r_6[29] /*16845*/;
  assign _1059_ = _1057_ | _1058_ /*16844*/;
  assign _1060_ = inv_7[13] ^ r_6[30] /*16842*/;
  assign sum_7[13] = _1060_ ^ _1059_ /*16841*/;
  assign _1061_ = _1060_ & _1059_ /*16840*/;
  assign _1062_ = inv_7[13] & r_6[30] /*16839*/;
  assign _1063_ = _1061_ | _1062_ /*16838*/;
  assign _1064_ = inv_7[14] ^ r_6[31] /*16836*/;
  assign sum_7[14] = _1064_ ^ _1063_ /*16835*/;
  assign _1065_ = _1064_ & _1063_ /*16834*/;
  assign _1066_ = inv_7[14] & r_6[31] /*16833*/;
  assign _1067_ = _1065_ | _1066_ /*16832*/;
  assign _1068_ = inv_7[15] ^ r_6[32] /*16830*/;
  assign sum_7[15] = _1068_ ^ _1067_ /*16829*/;
  assign _1069_ = _1068_ & _1067_ /*16828*/;
  assign _1070_ = inv_7[15] & r_6[32] /*16827*/;
  assign _1071_ = _1069_ | _1070_ /*16826*/;
  assign _1072_ = inv_7[16] ^ r_6[33] /*16824*/;
  assign sum_7[16] = _1072_ ^ _1071_ /*16823*/;
  assign _1073_ = _1072_ & _1071_ /*16822*/;
  assign _1074_ = inv_7[16] & r_6[33] /*16821*/;
  assign _1075_ = _1073_ | _1074_ /*16820*/;
  assign _1076_ = inv_7[17] ^ r_6[34] /*16818*/;
  assign sum_7[17] = _1076_ ^ _1075_ /*16817*/;
  assign _1077_ = _1076_ & _1075_ /*16816*/;
  assign _1078_ = inv_7[17] & r_6[34] /*16815*/;
  assign _1079_ = _1077_ | _1078_ /*16814*/;
  assign _1080_ = inv_7[18] ^ r_6[35] /*16812*/;
  assign sum_7[18] = _1080_ ^ _1079_ /*16811*/;
  assign _1081_ = _1080_ & _1079_ /*16810*/;
  assign _1082_ = inv_7[18] & r_6[35] /*16809*/;
  assign _1083_ = _1081_ | _1082_ /*16808*/;
  assign _1084_ = inv_7[19] ^ r_6[36] /*16806*/;
  assign sum_7[19] = _1084_ ^ _1083_ /*16805*/;
  assign _1085_ = _1084_ & _1083_ /*16804*/;
  assign _1086_ = inv_7[19] & r_6[36] /*16803*/;
  assign _1087_ = _1085_ | _1086_ /*16802*/;
  assign _1088_ = inv_7[20] ^ r_6[37] /*16800*/;
  assign sum_7[20] = _1088_ ^ _1087_ /*16799*/;
  assign _1089_ = _1088_ & _1087_ /*16798*/;
  assign _1090_ = inv_7[20] & r_6[37] /*16797*/;
  assign _1091_ = _1089_ | _1090_ /*16796*/;
  assign _1092_ = inv_7[21] ^ r_6[38] /*16794*/;
  assign sum_7[21] = _1092_ ^ _1091_ /*16793*/;
  assign _1093_ = _1092_ & _1091_ /*16792*/;
  assign _1094_ = inv_7[21] & r_6[38] /*16791*/;
  assign _1095_ = _1093_ | _1094_ /*16790*/;
  assign _1096_ = inv_7[22] ^ r_6[39] /*16788*/;
  assign sum_7[22] = _1096_ ^ _1095_ /*16787*/;
  assign _1097_ = _1096_ & _1095_ /*16786*/;
  assign _1098_ = inv_7[22] & r_6[39] /*16785*/;
  assign _1099_ = _1097_ | _1098_ /*16784*/;
  assign _1100_ = inv_7[23] ^ r_6[40] /*16782*/;
  assign sum_7[23] = _1100_ ^ _1099_ /*16781*/;
  assign _1101_ = _1100_ & _1099_ /*16780*/;
  assign _1102_ = inv_7[23] & r_6[40] /*16779*/;
  assign _1103_ = _1101_ | _1102_ /*16778*/;
  assign q[17] = ~sum_7[23] /*16797*/;
  assign m_7[0] = r_6[17] /*16796*/;
  assign m_7[1] = r_6[18] /*16795*/;
  assign m_7[2] = r_6[19] /*16794*/;
  assign m_7[3] = r_6[20] /*16793*/;
  assign m_7[4] = r_6[21] /*16792*/;
  assign m_7[5] = r_6[22] /*16791*/;
  assign m_7[6] = r_6[23] /*16790*/;
  assign m_7[7] = r_6[24] /*16789*/;
  assign m_7[8] = r_6[25] /*16788*/;
  assign m_7[9] = r_6[26] /*16787*/;
  assign m_7[10] = r_6[27] /*16786*/;
  assign m_7[11] = r_6[28] /*16785*/;
  assign m_7[12] = r_6[29] /*16784*/;
  assign m_7[13] = r_6[30] /*16783*/;
  assign m_7[14] = r_6[31] /*16782*/;
  assign m_7[15] = r_6[32] /*16781*/;
  assign m_7[16] = r_6[33] /*16780*/;
  assign m_7[17] = r_6[34] /*16779*/;
  assign m_7[18] = r_6[35] /*16778*/;
  assign m_7[19] = r_6[36] /*16777*/;
  assign m_7[20] = r_6[37] /*16776*/;
  assign m_7[21] = r_6[38] /*16775*/;
  assign m_7[22] = r_6[39] /*16774*/;
  assign m_7[23] = r_6[40] /*16773*/;
  assign _1104_ = ~q[17] /*16771*/;
  assign _1105_ = sum_7[0] & q[17] /*16770*/;
  assign _1106_ = m_7[0] & _1104_ /*16769*/;
  assign r_7[17] = _1106_ | _1105_ /*16768*/;
  assign _1107_ = ~q[17] /*16767*/;
  assign _1108_ = sum_7[1] & q[17] /*16766*/;
  assign _1109_ = m_7[1] & _1107_ /*16765*/;
  assign r_7[18] = _1109_ | _1108_ /*16764*/;
  assign _1110_ = ~q[17] /*16763*/;
  assign _1111_ = sum_7[2] & q[17] /*16762*/;
  assign _1112_ = m_7[2] & _1110_ /*16761*/;
  assign r_7[19] = _1112_ | _1111_ /*16760*/;
  assign _1113_ = ~q[17] /*16759*/;
  assign _1114_ = sum_7[3] & q[17] /*16758*/;
  assign _1115_ = m_7[3] & _1113_ /*16757*/;
  assign r_7[20] = _1115_ | _1114_ /*16756*/;
  assign _1116_ = ~q[17] /*16755*/;
  assign _1117_ = sum_7[4] & q[17] /*16754*/;
  assign _1118_ = m_7[4] & _1116_ /*16753*/;
  assign r_7[21] = _1118_ | _1117_ /*16752*/;
  assign _1119_ = ~q[17] /*16751*/;
  assign _1120_ = sum_7[5] & q[17] /*16750*/;
  assign _1121_ = m_7[5] & _1119_ /*16749*/;
  assign r_7[22] = _1121_ | _1120_ /*16748*/;
  assign _1122_ = ~q[17] /*16747*/;
  assign _1123_ = sum_7[6] & q[17] /*16746*/;
  assign _1124_ = m_7[6] & _1122_ /*16745*/;
  assign r_7[23] = _1124_ | _1123_ /*16744*/;
  assign _1125_ = ~q[17] /*16743*/;
  assign _1126_ = sum_7[7] & q[17] /*16742*/;
  assign _1127_ = m_7[7] & _1125_ /*16741*/;
  assign r_7[24] = _1127_ | _1126_ /*16740*/;
  assign _1128_ = ~q[17] /*16739*/;
  assign _1129_ = sum_7[8] & q[17] /*16738*/;
  assign _1130_ = m_7[8] & _1128_ /*16737*/;
  assign r_7[25] = _1130_ | _1129_ /*16736*/;
  assign _1131_ = ~q[17] /*16735*/;
  assign _1132_ = sum_7[9] & q[17] /*16734*/;
  assign _1133_ = m_7[9] & _1131_ /*16733*/;
  assign r_7[26] = _1133_ | _1132_ /*16732*/;
  assign _1134_ = ~q[17] /*16731*/;
  assign _1135_ = sum_7[10] & q[17] /*16730*/;
  assign _1136_ = m_7[10] & _1134_ /*16729*/;
  assign r_7[27] = _1136_ | _1135_ /*16728*/;
  assign _1137_ = ~q[17] /*16727*/;
  assign _1138_ = sum_7[11] & q[17] /*16726*/;
  assign _1139_ = m_7[11] & _1137_ /*16725*/;
  assign r_7[28] = _1139_ | _1138_ /*16724*/;
  assign _1140_ = ~q[17] /*16723*/;
  assign _1141_ = sum_7[12] & q[17] /*16722*/;
  assign _1142_ = m_7[12] & _1140_ /*16721*/;
  assign r_7[29] = _1142_ | _1141_ /*16720*/;
  assign _1143_ = ~q[17] /*16719*/;
  assign _1144_ = sum_7[13] & q[17] /*16718*/;
  assign _1145_ = m_7[13] & _1143_ /*16717*/;
  assign r_7[30] = _1145_ | _1144_ /*16716*/;
  assign _1146_ = ~q[17] /*16715*/;
  assign _1147_ = sum_7[14] & q[17] /*16714*/;
  assign _1148_ = m_7[14] & _1146_ /*16713*/;
  assign r_7[31] = _1148_ | _1147_ /*16712*/;
  assign _1149_ = ~q[17] /*16711*/;
  assign _1150_ = sum_7[15] & q[17] /*16710*/;
  assign _1151_ = m_7[15] & _1149_ /*16709*/;
  assign r_7[32] = _1151_ | _1150_ /*16708*/;
  assign _1152_ = ~q[17] /*16707*/;
  assign _1153_ = sum_7[16] & q[17] /*16706*/;
  assign _1154_ = m_7[16] & _1152_ /*16705*/;
  assign r_7[33] = _1154_ | _1153_ /*16704*/;
  assign _1155_ = ~q[17] /*16703*/;
  assign _1156_ = sum_7[17] & q[17] /*16702*/;
  assign _1157_ = m_7[17] & _1155_ /*16701*/;
  assign r_7[34] = _1157_ | _1156_ /*16700*/;
  assign _1158_ = ~q[17] /*16699*/;
  assign _1159_ = sum_7[18] & q[17] /*16698*/;
  assign _1160_ = m_7[18] & _1158_ /*16697*/;
  assign r_7[35] = _1160_ | _1159_ /*16696*/;
  assign _1161_ = ~q[17] /*16695*/;
  assign _1162_ = sum_7[19] & q[17] /*16694*/;
  assign _1163_ = m_7[19] & _1161_ /*16693*/;
  assign r_7[36] = _1163_ | _1162_ /*16692*/;
  assign _1164_ = ~q[17] /*16691*/;
  assign _1165_ = sum_7[20] & q[17] /*16690*/;
  assign _1166_ = m_7[20] & _1164_ /*16689*/;
  assign r_7[37] = _1166_ | _1165_ /*16688*/;
  assign _1167_ = ~q[17] /*16687*/;
  assign _1168_ = sum_7[21] & q[17] /*16686*/;
  assign _1169_ = m_7[21] & _1167_ /*16685*/;
  assign r_7[38] = _1169_ | _1168_ /*16684*/;
  assign _1170_ = ~q[17] /*16683*/;
  assign _1171_ = sum_7[22] & q[17] /*16682*/;
  assign _1172_ = m_7[22] & _1170_ /*16681*/;
  assign r_7[39] = _1172_ | _1171_ /*16680*/;
  assign _1173_ = ~q[17] /*16679*/;
  assign _1174_ = sum_7[23] & q[17] /*16678*/;
  assign _1175_ = m_7[23] & _1173_ /*16677*/;
  assign r_7[40] = _1175_ | _1174_ /*16676*/;
assign r_7[0]= r_6[0] /*16675*/;
assign r_7[1]= r_6[1] /*16674*/;
assign r_7[2]= r_6[2] /*16673*/;
assign r_7[3]= r_6[3] /*16672*/;
assign r_7[4]= r_6[4] /*16671*/;
assign r_7[5]= r_6[5] /*16670*/;
assign r_7[6]= r_6[6] /*16669*/;
assign r_7[7]= r_6[7] /*16668*/;
assign r_7[8]= r_6[8] /*16667*/;
assign r_7[9]= r_6[9] /*16666*/;
assign r_7[10]= r_6[10] /*16665*/;
assign r_7[11]= r_6[11] /*16664*/;
assign r_7[12]= r_6[12] /*16663*/;
assign r_7[13]= r_6[13] /*16662*/;
assign r_7[14]= r_6[14] /*16661*/;
assign r_7[15]= r_6[15] /*16660*/;
assign r_7[16]= r_6[16] /*16659*/;
  assign inv_8[0] = ~div[0] /*16608*/;
  assign inv_8[1] = ~div[1] /*16607*/;
  assign inv_8[2] = ~div[2] /*16606*/;
  assign inv_8[3] = ~div[3] /*16605*/;
  assign inv_8[4] = ~div[4] /*16604*/;
  assign inv_8[5] = ~div[5] /*16603*/;
  assign inv_8[6] = ~div[6] /*16602*/;
  assign inv_8[7] = ~div[7] /*16601*/;
  assign inv_8[8] = ~div[8] /*16600*/;
  assign inv_8[9] = ~div[9] /*16599*/;
  assign inv_8[10] = ~div[10] /*16598*/;
  assign inv_8[11] = ~div[11] /*16597*/;
  assign inv_8[12] = ~div[12] /*16596*/;
  assign inv_8[13] = ~div[13] /*16595*/;
  assign inv_8[14] = ~div[14] /*16594*/;
  assign inv_8[15] = ~div[15] /*16593*/;
  assign inv_8[16] = ~div[16] /*16592*/;
  assign inv_8[17] = ~div[17] /*16591*/;
  assign inv_8[18] = ~div[18] /*16590*/;
  assign inv_8[19] = ~div[19] /*16589*/;
  assign inv_8[20] = ~div[20] /*16588*/;
  assign inv_8[21] = ~div[21] /*16587*/;
  assign inv_8[22] = ~div[22] /*16586*/;
assign inv_8[23] = oneWire /*16585*/;
  assign _1176_ = inv_8[0] ^ r_7[16] /*16583*/;
  assign sum_8[0] = _1176_ ^ oneWire /*16582*/;
  assign _1177_ = _1176_ & oneWire /*16581*/;
  assign _1178_ = inv_8[0] & r_7[16] /*16580*/;
  assign _1179_ = _1177_ | _1178_ /*16579*/;
  assign _1180_ = inv_8[1] ^ r_7[17] /*16578*/;
  assign sum_8[1] = _1180_ ^ _1179_ /*16577*/;
  assign _1181_ = _1180_ & _1179_ /*16576*/;
  assign _1182_ = inv_8[1] & r_7[17] /*16575*/;
  assign _1183_ = _1181_ | _1182_ /*16574*/;
  assign _1184_ = inv_8[2] ^ r_7[18] /*16572*/;
  assign sum_8[2] = _1184_ ^ _1183_ /*16571*/;
  assign _1185_ = _1184_ & _1183_ /*16570*/;
  assign _1186_ = inv_8[2] & r_7[18] /*16569*/;
  assign _1187_ = _1185_ | _1186_ /*16568*/;
  assign _1188_ = inv_8[3] ^ r_7[19] /*16566*/;
  assign sum_8[3] = _1188_ ^ _1187_ /*16565*/;
  assign _1189_ = _1188_ & _1187_ /*16564*/;
  assign _1190_ = inv_8[3] & r_7[19] /*16563*/;
  assign _1191_ = _1189_ | _1190_ /*16562*/;
  assign _1192_ = inv_8[4] ^ r_7[20] /*16560*/;
  assign sum_8[4] = _1192_ ^ _1191_ /*16559*/;
  assign _1193_ = _1192_ & _1191_ /*16558*/;
  assign _1194_ = inv_8[4] & r_7[20] /*16557*/;
  assign _1195_ = _1193_ | _1194_ /*16556*/;
  assign _1196_ = inv_8[5] ^ r_7[21] /*16554*/;
  assign sum_8[5] = _1196_ ^ _1195_ /*16553*/;
  assign _1197_ = _1196_ & _1195_ /*16552*/;
  assign _1198_ = inv_8[5] & r_7[21] /*16551*/;
  assign _1199_ = _1197_ | _1198_ /*16550*/;
  assign _1200_ = inv_8[6] ^ r_7[22] /*16548*/;
  assign sum_8[6] = _1200_ ^ _1199_ /*16547*/;
  assign _1201_ = _1200_ & _1199_ /*16546*/;
  assign _1202_ = inv_8[6] & r_7[22] /*16545*/;
  assign _1203_ = _1201_ | _1202_ /*16544*/;
  assign _1204_ = inv_8[7] ^ r_7[23] /*16542*/;
  assign sum_8[7] = _1204_ ^ _1203_ /*16541*/;
  assign _1205_ = _1204_ & _1203_ /*16540*/;
  assign _1206_ = inv_8[7] & r_7[23] /*16539*/;
  assign _1207_ = _1205_ | _1206_ /*16538*/;
  assign _1208_ = inv_8[8] ^ r_7[24] /*16536*/;
  assign sum_8[8] = _1208_ ^ _1207_ /*16535*/;
  assign _1209_ = _1208_ & _1207_ /*16534*/;
  assign _1210_ = inv_8[8] & r_7[24] /*16533*/;
  assign _1211_ = _1209_ | _1210_ /*16532*/;
  assign _1212_ = inv_8[9] ^ r_7[25] /*16530*/;
  assign sum_8[9] = _1212_ ^ _1211_ /*16529*/;
  assign _1213_ = _1212_ & _1211_ /*16528*/;
  assign _1214_ = inv_8[9] & r_7[25] /*16527*/;
  assign _1215_ = _1213_ | _1214_ /*16526*/;
  assign _1216_ = inv_8[10] ^ r_7[26] /*16524*/;
  assign sum_8[10] = _1216_ ^ _1215_ /*16523*/;
  assign _1217_ = _1216_ & _1215_ /*16522*/;
  assign _1218_ = inv_8[10] & r_7[26] /*16521*/;
  assign _1219_ = _1217_ | _1218_ /*16520*/;
  assign _1220_ = inv_8[11] ^ r_7[27] /*16518*/;
  assign sum_8[11] = _1220_ ^ _1219_ /*16517*/;
  assign _1221_ = _1220_ & _1219_ /*16516*/;
  assign _1222_ = inv_8[11] & r_7[27] /*16515*/;
  assign _1223_ = _1221_ | _1222_ /*16514*/;
  assign _1224_ = inv_8[12] ^ r_7[28] /*16512*/;
  assign sum_8[12] = _1224_ ^ _1223_ /*16511*/;
  assign _1225_ = _1224_ & _1223_ /*16510*/;
  assign _1226_ = inv_8[12] & r_7[28] /*16509*/;
  assign _1227_ = _1225_ | _1226_ /*16508*/;
  assign _1228_ = inv_8[13] ^ r_7[29] /*16506*/;
  assign sum_8[13] = _1228_ ^ _1227_ /*16505*/;
  assign _1229_ = _1228_ & _1227_ /*16504*/;
  assign _1230_ = inv_8[13] & r_7[29] /*16503*/;
  assign _1231_ = _1229_ | _1230_ /*16502*/;
  assign _1232_ = inv_8[14] ^ r_7[30] /*16500*/;
  assign sum_8[14] = _1232_ ^ _1231_ /*16499*/;
  assign _1233_ = _1232_ & _1231_ /*16498*/;
  assign _1234_ = inv_8[14] & r_7[30] /*16497*/;
  assign _1235_ = _1233_ | _1234_ /*16496*/;
  assign _1236_ = inv_8[15] ^ r_7[31] /*16494*/;
  assign sum_8[15] = _1236_ ^ _1235_ /*16493*/;
  assign _1237_ = _1236_ & _1235_ /*16492*/;
  assign _1238_ = inv_8[15] & r_7[31] /*16491*/;
  assign _1239_ = _1237_ | _1238_ /*16490*/;
  assign _1240_ = inv_8[16] ^ r_7[32] /*16488*/;
  assign sum_8[16] = _1240_ ^ _1239_ /*16487*/;
  assign _1241_ = _1240_ & _1239_ /*16486*/;
  assign _1242_ = inv_8[16] & r_7[32] /*16485*/;
  assign _1243_ = _1241_ | _1242_ /*16484*/;
  assign _1244_ = inv_8[17] ^ r_7[33] /*16482*/;
  assign sum_8[17] = _1244_ ^ _1243_ /*16481*/;
  assign _1245_ = _1244_ & _1243_ /*16480*/;
  assign _1246_ = inv_8[17] & r_7[33] /*16479*/;
  assign _1247_ = _1245_ | _1246_ /*16478*/;
  assign _1248_ = inv_8[18] ^ r_7[34] /*16476*/;
  assign sum_8[18] = _1248_ ^ _1247_ /*16475*/;
  assign _1249_ = _1248_ & _1247_ /*16474*/;
  assign _1250_ = inv_8[18] & r_7[34] /*16473*/;
  assign _1251_ = _1249_ | _1250_ /*16472*/;
  assign _1252_ = inv_8[19] ^ r_7[35] /*16470*/;
  assign sum_8[19] = _1252_ ^ _1251_ /*16469*/;
  assign _1253_ = _1252_ & _1251_ /*16468*/;
  assign _1254_ = inv_8[19] & r_7[35] /*16467*/;
  assign _1255_ = _1253_ | _1254_ /*16466*/;
  assign _1256_ = inv_8[20] ^ r_7[36] /*16464*/;
  assign sum_8[20] = _1256_ ^ _1255_ /*16463*/;
  assign _1257_ = _1256_ & _1255_ /*16462*/;
  assign _1258_ = inv_8[20] & r_7[36] /*16461*/;
  assign _1259_ = _1257_ | _1258_ /*16460*/;
  assign _1260_ = inv_8[21] ^ r_7[37] /*16458*/;
  assign sum_8[21] = _1260_ ^ _1259_ /*16457*/;
  assign _1261_ = _1260_ & _1259_ /*16456*/;
  assign _1262_ = inv_8[21] & r_7[37] /*16455*/;
  assign _1263_ = _1261_ | _1262_ /*16454*/;
  assign _1264_ = inv_8[22] ^ r_7[38] /*16452*/;
  assign sum_8[22] = _1264_ ^ _1263_ /*16451*/;
  assign _1265_ = _1264_ & _1263_ /*16450*/;
  assign _1266_ = inv_8[22] & r_7[38] /*16449*/;
  assign _1267_ = _1265_ | _1266_ /*16448*/;
  assign _1268_ = inv_8[23] ^ r_7[39] /*16446*/;
  assign sum_8[23] = _1268_ ^ _1267_ /*16445*/;
  assign _1269_ = _1268_ & _1267_ /*16444*/;
  assign _1270_ = inv_8[23] & r_7[39] /*16443*/;
  assign _1271_ = _1269_ | _1270_ /*16442*/;
  assign q[16] = ~sum_8[23] /*16461*/;
  assign m_8[0] = r_7[16] /*16460*/;
  assign m_8[1] = r_7[17] /*16459*/;
  assign m_8[2] = r_7[18] /*16458*/;
  assign m_8[3] = r_7[19] /*16457*/;
  assign m_8[4] = r_7[20] /*16456*/;
  assign m_8[5] = r_7[21] /*16455*/;
  assign m_8[6] = r_7[22] /*16454*/;
  assign m_8[7] = r_7[23] /*16453*/;
  assign m_8[8] = r_7[24] /*16452*/;
  assign m_8[9] = r_7[25] /*16451*/;
  assign m_8[10] = r_7[26] /*16450*/;
  assign m_8[11] = r_7[27] /*16449*/;
  assign m_8[12] = r_7[28] /*16448*/;
  assign m_8[13] = r_7[29] /*16447*/;
  assign m_8[14] = r_7[30] /*16446*/;
  assign m_8[15] = r_7[31] /*16445*/;
  assign m_8[16] = r_7[32] /*16444*/;
  assign m_8[17] = r_7[33] /*16443*/;
  assign m_8[18] = r_7[34] /*16442*/;
  assign m_8[19] = r_7[35] /*16441*/;
  assign m_8[20] = r_7[36] /*16440*/;
  assign m_8[21] = r_7[37] /*16439*/;
  assign m_8[22] = r_7[38] /*16438*/;
  assign m_8[23] = r_7[39] /*16437*/;
  assign _1272_ = ~q[16] /*16435*/;
  assign _1273_ = sum_8[0] & q[16] /*16434*/;
  assign _1274_ = m_8[0] & _1272_ /*16433*/;
  assign r_8[16] = _1274_ | _1273_ /*16432*/;
  assign _1275_ = ~q[16] /*16431*/;
  assign _1276_ = sum_8[1] & q[16] /*16430*/;
  assign _1277_ = m_8[1] & _1275_ /*16429*/;
  assign r_8[17] = _1277_ | _1276_ /*16428*/;
  assign _1278_ = ~q[16] /*16427*/;
  assign _1279_ = sum_8[2] & q[16] /*16426*/;
  assign _1280_ = m_8[2] & _1278_ /*16425*/;
  assign r_8[18] = _1280_ | _1279_ /*16424*/;
  assign _1281_ = ~q[16] /*16423*/;
  assign _1282_ = sum_8[3] & q[16] /*16422*/;
  assign _1283_ = m_8[3] & _1281_ /*16421*/;
  assign r_8[19] = _1283_ | _1282_ /*16420*/;
  assign _1284_ = ~q[16] /*16419*/;
  assign _1285_ = sum_8[4] & q[16] /*16418*/;
  assign _1286_ = m_8[4] & _1284_ /*16417*/;
  assign r_8[20] = _1286_ | _1285_ /*16416*/;
  assign _1287_ = ~q[16] /*16415*/;
  assign _1288_ = sum_8[5] & q[16] /*16414*/;
  assign _1289_ = m_8[5] & _1287_ /*16413*/;
  assign r_8[21] = _1289_ | _1288_ /*16412*/;
  assign _1290_ = ~q[16] /*16411*/;
  assign _1291_ = sum_8[6] & q[16] /*16410*/;
  assign _1292_ = m_8[6] & _1290_ /*16409*/;
  assign r_8[22] = _1292_ | _1291_ /*16408*/;
  assign _1293_ = ~q[16] /*16407*/;
  assign _1294_ = sum_8[7] & q[16] /*16406*/;
  assign _1295_ = m_8[7] & _1293_ /*16405*/;
  assign r_8[23] = _1295_ | _1294_ /*16404*/;
  assign _1296_ = ~q[16] /*16403*/;
  assign _1297_ = sum_8[8] & q[16] /*16402*/;
  assign _1298_ = m_8[8] & _1296_ /*16401*/;
  assign r_8[24] = _1298_ | _1297_ /*16400*/;
  assign _1299_ = ~q[16] /*16399*/;
  assign _1300_ = sum_8[9] & q[16] /*16398*/;
  assign _1301_ = m_8[9] & _1299_ /*16397*/;
  assign r_8[25] = _1301_ | _1300_ /*16396*/;
  assign _1302_ = ~q[16] /*16395*/;
  assign _1303_ = sum_8[10] & q[16] /*16394*/;
  assign _1304_ = m_8[10] & _1302_ /*16393*/;
  assign r_8[26] = _1304_ | _1303_ /*16392*/;
  assign _1305_ = ~q[16] /*16391*/;
  assign _1306_ = sum_8[11] & q[16] /*16390*/;
  assign _1307_ = m_8[11] & _1305_ /*16389*/;
  assign r_8[27] = _1307_ | _1306_ /*16388*/;
  assign _1308_ = ~q[16] /*16387*/;
  assign _1309_ = sum_8[12] & q[16] /*16386*/;
  assign _1310_ = m_8[12] & _1308_ /*16385*/;
  assign r_8[28] = _1310_ | _1309_ /*16384*/;
  assign _1311_ = ~q[16] /*16383*/;
  assign _1312_ = sum_8[13] & q[16] /*16382*/;
  assign _1313_ = m_8[13] & _1311_ /*16381*/;
  assign r_8[29] = _1313_ | _1312_ /*16380*/;
  assign _1314_ = ~q[16] /*16379*/;
  assign _1315_ = sum_8[14] & q[16] /*16378*/;
  assign _1316_ = m_8[14] & _1314_ /*16377*/;
  assign r_8[30] = _1316_ | _1315_ /*16376*/;
  assign _1317_ = ~q[16] /*16375*/;
  assign _1318_ = sum_8[15] & q[16] /*16374*/;
  assign _1319_ = m_8[15] & _1317_ /*16373*/;
  assign r_8[31] = _1319_ | _1318_ /*16372*/;
  assign _1320_ = ~q[16] /*16371*/;
  assign _1321_ = sum_8[16] & q[16] /*16370*/;
  assign _1322_ = m_8[16] & _1320_ /*16369*/;
  assign r_8[32] = _1322_ | _1321_ /*16368*/;
  assign _1323_ = ~q[16] /*16367*/;
  assign _1324_ = sum_8[17] & q[16] /*16366*/;
  assign _1325_ = m_8[17] & _1323_ /*16365*/;
  assign r_8[33] = _1325_ | _1324_ /*16364*/;
  assign _1326_ = ~q[16] /*16363*/;
  assign _1327_ = sum_8[18] & q[16] /*16362*/;
  assign _1328_ = m_8[18] & _1326_ /*16361*/;
  assign r_8[34] = _1328_ | _1327_ /*16360*/;
  assign _1329_ = ~q[16] /*16359*/;
  assign _1330_ = sum_8[19] & q[16] /*16358*/;
  assign _1331_ = m_8[19] & _1329_ /*16357*/;
  assign r_8[35] = _1331_ | _1330_ /*16356*/;
  assign _1332_ = ~q[16] /*16355*/;
  assign _1333_ = sum_8[20] & q[16] /*16354*/;
  assign _1334_ = m_8[20] & _1332_ /*16353*/;
  assign r_8[36] = _1334_ | _1333_ /*16352*/;
  assign _1335_ = ~q[16] /*16351*/;
  assign _1336_ = sum_8[21] & q[16] /*16350*/;
  assign _1337_ = m_8[21] & _1335_ /*16349*/;
  assign r_8[37] = _1337_ | _1336_ /*16348*/;
  assign _1338_ = ~q[16] /*16347*/;
  assign _1339_ = sum_8[22] & q[16] /*16346*/;
  assign _1340_ = m_8[22] & _1338_ /*16345*/;
  assign r_8[38] = _1340_ | _1339_ /*16344*/;
  assign _1341_ = ~q[16] /*16343*/;
  assign _1342_ = sum_8[23] & q[16] /*16342*/;
  assign _1343_ = m_8[23] & _1341_ /*16341*/;
  assign r_8[39] = _1343_ | _1342_ /*16340*/;
assign r_8[0]= r_7[0] /*16339*/;
assign r_8[1]= r_7[1] /*16338*/;
assign r_8[2]= r_7[2] /*16337*/;
assign r_8[3]= r_7[3] /*16336*/;
assign r_8[4]= r_7[4] /*16335*/;
assign r_8[5]= r_7[5] /*16334*/;
assign r_8[6]= r_7[6] /*16333*/;
assign r_8[7]= r_7[7] /*16332*/;
assign r_8[8]= r_7[8] /*16331*/;
assign r_8[9]= r_7[9] /*16330*/;
assign r_8[10]= r_7[10] /*16329*/;
assign r_8[11]= r_7[11] /*16328*/;
assign r_8[12]= r_7[12] /*16327*/;
assign r_8[13]= r_7[13] /*16326*/;
assign r_8[14]= r_7[14] /*16325*/;
assign r_8[15]= r_7[15] /*16324*/;
  assign inv_9[0] = ~div[0] /*16272*/;
  assign inv_9[1] = ~div[1] /*16271*/;
  assign inv_9[2] = ~div[2] /*16270*/;
  assign inv_9[3] = ~div[3] /*16269*/;
  assign inv_9[4] = ~div[4] /*16268*/;
  assign inv_9[5] = ~div[5] /*16267*/;
  assign inv_9[6] = ~div[6] /*16266*/;
  assign inv_9[7] = ~div[7] /*16265*/;
  assign inv_9[8] = ~div[8] /*16264*/;
  assign inv_9[9] = ~div[9] /*16263*/;
  assign inv_9[10] = ~div[10] /*16262*/;
  assign inv_9[11] = ~div[11] /*16261*/;
  assign inv_9[12] = ~div[12] /*16260*/;
  assign inv_9[13] = ~div[13] /*16259*/;
  assign inv_9[14] = ~div[14] /*16258*/;
  assign inv_9[15] = ~div[15] /*16257*/;
  assign inv_9[16] = ~div[16] /*16256*/;
  assign inv_9[17] = ~div[17] /*16255*/;
  assign inv_9[18] = ~div[18] /*16254*/;
  assign inv_9[19] = ~div[19] /*16253*/;
  assign inv_9[20] = ~div[20] /*16252*/;
  assign inv_9[21] = ~div[21] /*16251*/;
  assign inv_9[22] = ~div[22] /*16250*/;
assign inv_9[23] = oneWire /*16249*/;
  assign _1344_ = inv_9[0] ^ r_8[15] /*16247*/;
  assign sum_9[0] = _1344_ ^ oneWire /*16246*/;
  assign _1345_ = _1344_ & oneWire /*16245*/;
  assign _1346_ = inv_9[0] & r_8[15] /*16244*/;
  assign _1347_ = _1345_ | _1346_ /*16243*/;
  assign _1348_ = inv_9[1] ^ r_8[16] /*16242*/;
  assign sum_9[1] = _1348_ ^ _1347_ /*16241*/;
  assign _1349_ = _1348_ & _1347_ /*16240*/;
  assign _1350_ = inv_9[1] & r_8[16] /*16239*/;
  assign _1351_ = _1349_ | _1350_ /*16238*/;
  assign _1352_ = inv_9[2] ^ r_8[17] /*16236*/;
  assign sum_9[2] = _1352_ ^ _1351_ /*16235*/;
  assign _1353_ = _1352_ & _1351_ /*16234*/;
  assign _1354_ = inv_9[2] & r_8[17] /*16233*/;
  assign _1355_ = _1353_ | _1354_ /*16232*/;
  assign _1356_ = inv_9[3] ^ r_8[18] /*16230*/;
  assign sum_9[3] = _1356_ ^ _1355_ /*16229*/;
  assign _1357_ = _1356_ & _1355_ /*16228*/;
  assign _1358_ = inv_9[3] & r_8[18] /*16227*/;
  assign _1359_ = _1357_ | _1358_ /*16226*/;
  assign _1360_ = inv_9[4] ^ r_8[19] /*16224*/;
  assign sum_9[4] = _1360_ ^ _1359_ /*16223*/;
  assign _1361_ = _1360_ & _1359_ /*16222*/;
  assign _1362_ = inv_9[4] & r_8[19] /*16221*/;
  assign _1363_ = _1361_ | _1362_ /*16220*/;
  assign _1364_ = inv_9[5] ^ r_8[20] /*16218*/;
  assign sum_9[5] = _1364_ ^ _1363_ /*16217*/;
  assign _1365_ = _1364_ & _1363_ /*16216*/;
  assign _1366_ = inv_9[5] & r_8[20] /*16215*/;
  assign _1367_ = _1365_ | _1366_ /*16214*/;
  assign _1368_ = inv_9[6] ^ r_8[21] /*16212*/;
  assign sum_9[6] = _1368_ ^ _1367_ /*16211*/;
  assign _1369_ = _1368_ & _1367_ /*16210*/;
  assign _1370_ = inv_9[6] & r_8[21] /*16209*/;
  assign _1371_ = _1369_ | _1370_ /*16208*/;
  assign _1372_ = inv_9[7] ^ r_8[22] /*16206*/;
  assign sum_9[7] = _1372_ ^ _1371_ /*16205*/;
  assign _1373_ = _1372_ & _1371_ /*16204*/;
  assign _1374_ = inv_9[7] & r_8[22] /*16203*/;
  assign _1375_ = _1373_ | _1374_ /*16202*/;
  assign _1376_ = inv_9[8] ^ r_8[23] /*16200*/;
  assign sum_9[8] = _1376_ ^ _1375_ /*16199*/;
  assign _1377_ = _1376_ & _1375_ /*16198*/;
  assign _1378_ = inv_9[8] & r_8[23] /*16197*/;
  assign _1379_ = _1377_ | _1378_ /*16196*/;
  assign _1380_ = inv_9[9] ^ r_8[24] /*16194*/;
  assign sum_9[9] = _1380_ ^ _1379_ /*16193*/;
  assign _1381_ = _1380_ & _1379_ /*16192*/;
  assign _1382_ = inv_9[9] & r_8[24] /*16191*/;
  assign _1383_ = _1381_ | _1382_ /*16190*/;
  assign _1384_ = inv_9[10] ^ r_8[25] /*16188*/;
  assign sum_9[10] = _1384_ ^ _1383_ /*16187*/;
  assign _1385_ = _1384_ & _1383_ /*16186*/;
  assign _1386_ = inv_9[10] & r_8[25] /*16185*/;
  assign _1387_ = _1385_ | _1386_ /*16184*/;
  assign _1388_ = inv_9[11] ^ r_8[26] /*16182*/;
  assign sum_9[11] = _1388_ ^ _1387_ /*16181*/;
  assign _1389_ = _1388_ & _1387_ /*16180*/;
  assign _1390_ = inv_9[11] & r_8[26] /*16179*/;
  assign _1391_ = _1389_ | _1390_ /*16178*/;
  assign _1392_ = inv_9[12] ^ r_8[27] /*16176*/;
  assign sum_9[12] = _1392_ ^ _1391_ /*16175*/;
  assign _1393_ = _1392_ & _1391_ /*16174*/;
  assign _1394_ = inv_9[12] & r_8[27] /*16173*/;
  assign _1395_ = _1393_ | _1394_ /*16172*/;
  assign _1396_ = inv_9[13] ^ r_8[28] /*16170*/;
  assign sum_9[13] = _1396_ ^ _1395_ /*16169*/;
  assign _1397_ = _1396_ & _1395_ /*16168*/;
  assign _1398_ = inv_9[13] & r_8[28] /*16167*/;
  assign _1399_ = _1397_ | _1398_ /*16166*/;
  assign _1400_ = inv_9[14] ^ r_8[29] /*16164*/;
  assign sum_9[14] = _1400_ ^ _1399_ /*16163*/;
  assign _1401_ = _1400_ & _1399_ /*16162*/;
  assign _1402_ = inv_9[14] & r_8[29] /*16161*/;
  assign _1403_ = _1401_ | _1402_ /*16160*/;
  assign _1404_ = inv_9[15] ^ r_8[30] /*16158*/;
  assign sum_9[15] = _1404_ ^ _1403_ /*16157*/;
  assign _1405_ = _1404_ & _1403_ /*16156*/;
  assign _1406_ = inv_9[15] & r_8[30] /*16155*/;
  assign _1407_ = _1405_ | _1406_ /*16154*/;
  assign _1408_ = inv_9[16] ^ r_8[31] /*16152*/;
  assign sum_9[16] = _1408_ ^ _1407_ /*16151*/;
  assign _1409_ = _1408_ & _1407_ /*16150*/;
  assign _1410_ = inv_9[16] & r_8[31] /*16149*/;
  assign _1411_ = _1409_ | _1410_ /*16148*/;
  assign _1412_ = inv_9[17] ^ r_8[32] /*16146*/;
  assign sum_9[17] = _1412_ ^ _1411_ /*16145*/;
  assign _1413_ = _1412_ & _1411_ /*16144*/;
  assign _1414_ = inv_9[17] & r_8[32] /*16143*/;
  assign _1415_ = _1413_ | _1414_ /*16142*/;
  assign _1416_ = inv_9[18] ^ r_8[33] /*16140*/;
  assign sum_9[18] = _1416_ ^ _1415_ /*16139*/;
  assign _1417_ = _1416_ & _1415_ /*16138*/;
  assign _1418_ = inv_9[18] & r_8[33] /*16137*/;
  assign _1419_ = _1417_ | _1418_ /*16136*/;
  assign _1420_ = inv_9[19] ^ r_8[34] /*16134*/;
  assign sum_9[19] = _1420_ ^ _1419_ /*16133*/;
  assign _1421_ = _1420_ & _1419_ /*16132*/;
  assign _1422_ = inv_9[19] & r_8[34] /*16131*/;
  assign _1423_ = _1421_ | _1422_ /*16130*/;
  assign _1424_ = inv_9[20] ^ r_8[35] /*16128*/;
  assign sum_9[20] = _1424_ ^ _1423_ /*16127*/;
  assign _1425_ = _1424_ & _1423_ /*16126*/;
  assign _1426_ = inv_9[20] & r_8[35] /*16125*/;
  assign _1427_ = _1425_ | _1426_ /*16124*/;
  assign _1428_ = inv_9[21] ^ r_8[36] /*16122*/;
  assign sum_9[21] = _1428_ ^ _1427_ /*16121*/;
  assign _1429_ = _1428_ & _1427_ /*16120*/;
  assign _1430_ = inv_9[21] & r_8[36] /*16119*/;
  assign _1431_ = _1429_ | _1430_ /*16118*/;
  assign _1432_ = inv_9[22] ^ r_8[37] /*16116*/;
  assign sum_9[22] = _1432_ ^ _1431_ /*16115*/;
  assign _1433_ = _1432_ & _1431_ /*16114*/;
  assign _1434_ = inv_9[22] & r_8[37] /*16113*/;
  assign _1435_ = _1433_ | _1434_ /*16112*/;
  assign _1436_ = inv_9[23] ^ r_8[38] /*16110*/;
  assign sum_9[23] = _1436_ ^ _1435_ /*16109*/;
  assign _1437_ = _1436_ & _1435_ /*16108*/;
  assign _1438_ = inv_9[23] & r_8[38] /*16107*/;
  assign _1439_ = _1437_ | _1438_ /*16106*/;
  assign q[15] = ~sum_9[23] /*16125*/;
  assign m_9[0] = r_8[15] /*16124*/;
  assign m_9[1] = r_8[16] /*16123*/;
  assign m_9[2] = r_8[17] /*16122*/;
  assign m_9[3] = r_8[18] /*16121*/;
  assign m_9[4] = r_8[19] /*16120*/;
  assign m_9[5] = r_8[20] /*16119*/;
  assign m_9[6] = r_8[21] /*16118*/;
  assign m_9[7] = r_8[22] /*16117*/;
  assign m_9[8] = r_8[23] /*16116*/;
  assign m_9[9] = r_8[24] /*16115*/;
  assign m_9[10] = r_8[25] /*16114*/;
  assign m_9[11] = r_8[26] /*16113*/;
  assign m_9[12] = r_8[27] /*16112*/;
  assign m_9[13] = r_8[28] /*16111*/;
  assign m_9[14] = r_8[29] /*16110*/;
  assign m_9[15] = r_8[30] /*16109*/;
  assign m_9[16] = r_8[31] /*16108*/;
  assign m_9[17] = r_8[32] /*16107*/;
  assign m_9[18] = r_8[33] /*16106*/;
  assign m_9[19] = r_8[34] /*16105*/;
  assign m_9[20] = r_8[35] /*16104*/;
  assign m_9[21] = r_8[36] /*16103*/;
  assign m_9[22] = r_8[37] /*16102*/;
  assign m_9[23] = r_8[38] /*16101*/;
  assign _1440_ = ~q[15] /*16099*/;
  assign _1441_ = sum_9[0] & q[15] /*16098*/;
  assign _1442_ = m_9[0] & _1440_ /*16097*/;
  assign r_9[15] = _1442_ | _1441_ /*16096*/;
  assign _1443_ = ~q[15] /*16095*/;
  assign _1444_ = sum_9[1] & q[15] /*16094*/;
  assign _1445_ = m_9[1] & _1443_ /*16093*/;
  assign r_9[16] = _1445_ | _1444_ /*16092*/;
  assign _1446_ = ~q[15] /*16091*/;
  assign _1447_ = sum_9[2] & q[15] /*16090*/;
  assign _1448_ = m_9[2] & _1446_ /*16089*/;
  assign r_9[17] = _1448_ | _1447_ /*16088*/;
  assign _1449_ = ~q[15] /*16087*/;
  assign _1450_ = sum_9[3] & q[15] /*16086*/;
  assign _1451_ = m_9[3] & _1449_ /*16085*/;
  assign r_9[18] = _1451_ | _1450_ /*16084*/;
  assign _1452_ = ~q[15] /*16083*/;
  assign _1453_ = sum_9[4] & q[15] /*16082*/;
  assign _1454_ = m_9[4] & _1452_ /*16081*/;
  assign r_9[19] = _1454_ | _1453_ /*16080*/;
  assign _1455_ = ~q[15] /*16079*/;
  assign _1456_ = sum_9[5] & q[15] /*16078*/;
  assign _1457_ = m_9[5] & _1455_ /*16077*/;
  assign r_9[20] = _1457_ | _1456_ /*16076*/;
  assign _1458_ = ~q[15] /*16075*/;
  assign _1459_ = sum_9[6] & q[15] /*16074*/;
  assign _1460_ = m_9[6] & _1458_ /*16073*/;
  assign r_9[21] = _1460_ | _1459_ /*16072*/;
  assign _1461_ = ~q[15] /*16071*/;
  assign _1462_ = sum_9[7] & q[15] /*16070*/;
  assign _1463_ = m_9[7] & _1461_ /*16069*/;
  assign r_9[22] = _1463_ | _1462_ /*16068*/;
  assign _1464_ = ~q[15] /*16067*/;
  assign _1465_ = sum_9[8] & q[15] /*16066*/;
  assign _1466_ = m_9[8] & _1464_ /*16065*/;
  assign r_9[23] = _1466_ | _1465_ /*16064*/;
  assign _1467_ = ~q[15] /*16063*/;
  assign _1468_ = sum_9[9] & q[15] /*16062*/;
  assign _1469_ = m_9[9] & _1467_ /*16061*/;
  assign r_9[24] = _1469_ | _1468_ /*16060*/;
  assign _1470_ = ~q[15] /*16059*/;
  assign _1471_ = sum_9[10] & q[15] /*16058*/;
  assign _1472_ = m_9[10] & _1470_ /*16057*/;
  assign r_9[25] = _1472_ | _1471_ /*16056*/;
  assign _1473_ = ~q[15] /*16055*/;
  assign _1474_ = sum_9[11] & q[15] /*16054*/;
  assign _1475_ = m_9[11] & _1473_ /*16053*/;
  assign r_9[26] = _1475_ | _1474_ /*16052*/;
  assign _1476_ = ~q[15] /*16051*/;
  assign _1477_ = sum_9[12] & q[15] /*16050*/;
  assign _1478_ = m_9[12] & _1476_ /*16049*/;
  assign r_9[27] = _1478_ | _1477_ /*16048*/;
  assign _1479_ = ~q[15] /*16047*/;
  assign _1480_ = sum_9[13] & q[15] /*16046*/;
  assign _1481_ = m_9[13] & _1479_ /*16045*/;
  assign r_9[28] = _1481_ | _1480_ /*16044*/;
  assign _1482_ = ~q[15] /*16043*/;
  assign _1483_ = sum_9[14] & q[15] /*16042*/;
  assign _1484_ = m_9[14] & _1482_ /*16041*/;
  assign r_9[29] = _1484_ | _1483_ /*16040*/;
  assign _1485_ = ~q[15] /*16039*/;
  assign _1486_ = sum_9[15] & q[15] /*16038*/;
  assign _1487_ = m_9[15] & _1485_ /*16037*/;
  assign r_9[30] = _1487_ | _1486_ /*16036*/;
  assign _1488_ = ~q[15] /*16035*/;
  assign _1489_ = sum_9[16] & q[15] /*16034*/;
  assign _1490_ = m_9[16] & _1488_ /*16033*/;
  assign r_9[31] = _1490_ | _1489_ /*16032*/;
  assign _1491_ = ~q[15] /*16031*/;
  assign _1492_ = sum_9[17] & q[15] /*16030*/;
  assign _1493_ = m_9[17] & _1491_ /*16029*/;
  assign r_9[32] = _1493_ | _1492_ /*16028*/;
  assign _1494_ = ~q[15] /*16027*/;
  assign _1495_ = sum_9[18] & q[15] /*16026*/;
  assign _1496_ = m_9[18] & _1494_ /*16025*/;
  assign r_9[33] = _1496_ | _1495_ /*16024*/;
  assign _1497_ = ~q[15] /*16023*/;
  assign _1498_ = sum_9[19] & q[15] /*16022*/;
  assign _1499_ = m_9[19] & _1497_ /*16021*/;
  assign r_9[34] = _1499_ | _1498_ /*16020*/;
  assign _1500_ = ~q[15] /*16019*/;
  assign _1501_ = sum_9[20] & q[15] /*16018*/;
  assign _1502_ = m_9[20] & _1500_ /*16017*/;
  assign r_9[35] = _1502_ | _1501_ /*16016*/;
  assign _1503_ = ~q[15] /*16015*/;
  assign _1504_ = sum_9[21] & q[15] /*16014*/;
  assign _1505_ = m_9[21] & _1503_ /*16013*/;
  assign r_9[36] = _1505_ | _1504_ /*16012*/;
  assign _1506_ = ~q[15] /*16011*/;
  assign _1507_ = sum_9[22] & q[15] /*16010*/;
  assign _1508_ = m_9[22] & _1506_ /*16009*/;
  assign r_9[37] = _1508_ | _1507_ /*16008*/;
  assign _1509_ = ~q[15] /*16007*/;
  assign _1510_ = sum_9[23] & q[15] /*16006*/;
  assign _1511_ = m_9[23] & _1509_ /*16005*/;
  assign r_9[38] = _1511_ | _1510_ /*16004*/;
assign r_9[0]= r_8[0] /*16003*/;
assign r_9[1]= r_8[1] /*16002*/;
assign r_9[2]= r_8[2] /*16001*/;
assign r_9[3]= r_8[3] /*16000*/;
assign r_9[4]= r_8[4] /*15999*/;
assign r_9[5]= r_8[5] /*15998*/;
assign r_9[6]= r_8[6] /*15997*/;
assign r_9[7]= r_8[7] /*15996*/;
assign r_9[8]= r_8[8] /*15995*/;
assign r_9[9]= r_8[9] /*15994*/;
assign r_9[10]= r_8[10] /*15993*/;
assign r_9[11]= r_8[11] /*15992*/;
assign r_9[12]= r_8[12] /*15991*/;
assign r_9[13]= r_8[13] /*15990*/;
assign r_9[14]= r_8[14] /*15989*/;
  assign inv_10[0] = ~div[0] /*15936*/;
  assign inv_10[1] = ~div[1] /*15935*/;
  assign inv_10[2] = ~div[2] /*15934*/;
  assign inv_10[3] = ~div[3] /*15933*/;
  assign inv_10[4] = ~div[4] /*15932*/;
  assign inv_10[5] = ~div[5] /*15931*/;
  assign inv_10[6] = ~div[6] /*15930*/;
  assign inv_10[7] = ~div[7] /*15929*/;
  assign inv_10[8] = ~div[8] /*15928*/;
  assign inv_10[9] = ~div[9] /*15927*/;
  assign inv_10[10] = ~div[10] /*15926*/;
  assign inv_10[11] = ~div[11] /*15925*/;
  assign inv_10[12] = ~div[12] /*15924*/;
  assign inv_10[13] = ~div[13] /*15923*/;
  assign inv_10[14] = ~div[14] /*15922*/;
  assign inv_10[15] = ~div[15] /*15921*/;
  assign inv_10[16] = ~div[16] /*15920*/;
  assign inv_10[17] = ~div[17] /*15919*/;
  assign inv_10[18] = ~div[18] /*15918*/;
  assign inv_10[19] = ~div[19] /*15917*/;
  assign inv_10[20] = ~div[20] /*15916*/;
  assign inv_10[21] = ~div[21] /*15915*/;
  assign inv_10[22] = ~div[22] /*15914*/;
assign inv_10[23] = oneWire /*15913*/;
  assign _1512_ = inv_10[0] ^ r_9[14] /*15911*/;
  assign sum_10[0] = _1512_ ^ oneWire /*15910*/;
  assign _1513_ = _1512_ & oneWire /*15909*/;
  assign _1514_ = inv_10[0] & r_9[14] /*15908*/;
  assign _1515_ = _1513_ | _1514_ /*15907*/;
  assign _1516_ = inv_10[1] ^ r_9[15] /*15906*/;
  assign sum_10[1] = _1516_ ^ _1515_ /*15905*/;
  assign _1517_ = _1516_ & _1515_ /*15904*/;
  assign _1518_ = inv_10[1] & r_9[15] /*15903*/;
  assign _1519_ = _1517_ | _1518_ /*15902*/;
  assign _1520_ = inv_10[2] ^ r_9[16] /*15900*/;
  assign sum_10[2] = _1520_ ^ _1519_ /*15899*/;
  assign _1521_ = _1520_ & _1519_ /*15898*/;
  assign _1522_ = inv_10[2] & r_9[16] /*15897*/;
  assign _1523_ = _1521_ | _1522_ /*15896*/;
  assign _1524_ = inv_10[3] ^ r_9[17] /*15894*/;
  assign sum_10[3] = _1524_ ^ _1523_ /*15893*/;
  assign _1525_ = _1524_ & _1523_ /*15892*/;
  assign _1526_ = inv_10[3] & r_9[17] /*15891*/;
  assign _1527_ = _1525_ | _1526_ /*15890*/;
  assign _1528_ = inv_10[4] ^ r_9[18] /*15888*/;
  assign sum_10[4] = _1528_ ^ _1527_ /*15887*/;
  assign _1529_ = _1528_ & _1527_ /*15886*/;
  assign _1530_ = inv_10[4] & r_9[18] /*15885*/;
  assign _1531_ = _1529_ | _1530_ /*15884*/;
  assign _1532_ = inv_10[5] ^ r_9[19] /*15882*/;
  assign sum_10[5] = _1532_ ^ _1531_ /*15881*/;
  assign _1533_ = _1532_ & _1531_ /*15880*/;
  assign _1534_ = inv_10[5] & r_9[19] /*15879*/;
  assign _1535_ = _1533_ | _1534_ /*15878*/;
  assign _1536_ = inv_10[6] ^ r_9[20] /*15876*/;
  assign sum_10[6] = _1536_ ^ _1535_ /*15875*/;
  assign _1537_ = _1536_ & _1535_ /*15874*/;
  assign _1538_ = inv_10[6] & r_9[20] /*15873*/;
  assign _1539_ = _1537_ | _1538_ /*15872*/;
  assign _1540_ = inv_10[7] ^ r_9[21] /*15870*/;
  assign sum_10[7] = _1540_ ^ _1539_ /*15869*/;
  assign _1541_ = _1540_ & _1539_ /*15868*/;
  assign _1542_ = inv_10[7] & r_9[21] /*15867*/;
  assign _1543_ = _1541_ | _1542_ /*15866*/;
  assign _1544_ = inv_10[8] ^ r_9[22] /*15864*/;
  assign sum_10[8] = _1544_ ^ _1543_ /*15863*/;
  assign _1545_ = _1544_ & _1543_ /*15862*/;
  assign _1546_ = inv_10[8] & r_9[22] /*15861*/;
  assign _1547_ = _1545_ | _1546_ /*15860*/;
  assign _1548_ = inv_10[9] ^ r_9[23] /*15858*/;
  assign sum_10[9] = _1548_ ^ _1547_ /*15857*/;
  assign _1549_ = _1548_ & _1547_ /*15856*/;
  assign _1550_ = inv_10[9] & r_9[23] /*15855*/;
  assign _1551_ = _1549_ | _1550_ /*15854*/;
  assign _1552_ = inv_10[10] ^ r_9[24] /*15852*/;
  assign sum_10[10] = _1552_ ^ _1551_ /*15851*/;
  assign _1553_ = _1552_ & _1551_ /*15850*/;
  assign _1554_ = inv_10[10] & r_9[24] /*15849*/;
  assign _1555_ = _1553_ | _1554_ /*15848*/;
  assign _1556_ = inv_10[11] ^ r_9[25] /*15846*/;
  assign sum_10[11] = _1556_ ^ _1555_ /*15845*/;
  assign _1557_ = _1556_ & _1555_ /*15844*/;
  assign _1558_ = inv_10[11] & r_9[25] /*15843*/;
  assign _1559_ = _1557_ | _1558_ /*15842*/;
  assign _1560_ = inv_10[12] ^ r_9[26] /*15840*/;
  assign sum_10[12] = _1560_ ^ _1559_ /*15839*/;
  assign _1561_ = _1560_ & _1559_ /*15838*/;
  assign _1562_ = inv_10[12] & r_9[26] /*15837*/;
  assign _1563_ = _1561_ | _1562_ /*15836*/;
  assign _1564_ = inv_10[13] ^ r_9[27] /*15834*/;
  assign sum_10[13] = _1564_ ^ _1563_ /*15833*/;
  assign _1565_ = _1564_ & _1563_ /*15832*/;
  assign _1566_ = inv_10[13] & r_9[27] /*15831*/;
  assign _1567_ = _1565_ | _1566_ /*15830*/;
  assign _1568_ = inv_10[14] ^ r_9[28] /*15828*/;
  assign sum_10[14] = _1568_ ^ _1567_ /*15827*/;
  assign _1569_ = _1568_ & _1567_ /*15826*/;
  assign _1570_ = inv_10[14] & r_9[28] /*15825*/;
  assign _1571_ = _1569_ | _1570_ /*15824*/;
  assign _1572_ = inv_10[15] ^ r_9[29] /*15822*/;
  assign sum_10[15] = _1572_ ^ _1571_ /*15821*/;
  assign _1573_ = _1572_ & _1571_ /*15820*/;
  assign _1574_ = inv_10[15] & r_9[29] /*15819*/;
  assign _1575_ = _1573_ | _1574_ /*15818*/;
  assign _1576_ = inv_10[16] ^ r_9[30] /*15816*/;
  assign sum_10[16] = _1576_ ^ _1575_ /*15815*/;
  assign _1577_ = _1576_ & _1575_ /*15814*/;
  assign _1578_ = inv_10[16] & r_9[30] /*15813*/;
  assign _1579_ = _1577_ | _1578_ /*15812*/;
  assign _1580_ = inv_10[17] ^ r_9[31] /*15810*/;
  assign sum_10[17] = _1580_ ^ _1579_ /*15809*/;
  assign _1581_ = _1580_ & _1579_ /*15808*/;
  assign _1582_ = inv_10[17] & r_9[31] /*15807*/;
  assign _1583_ = _1581_ | _1582_ /*15806*/;
  assign _1584_ = inv_10[18] ^ r_9[32] /*15804*/;
  assign sum_10[18] = _1584_ ^ _1583_ /*15803*/;
  assign _1585_ = _1584_ & _1583_ /*15802*/;
  assign _1586_ = inv_10[18] & r_9[32] /*15801*/;
  assign _1587_ = _1585_ | _1586_ /*15800*/;
  assign _1588_ = inv_10[19] ^ r_9[33] /*15798*/;
  assign sum_10[19] = _1588_ ^ _1587_ /*15797*/;
  assign _1589_ = _1588_ & _1587_ /*15796*/;
  assign _1590_ = inv_10[19] & r_9[33] /*15795*/;
  assign _1591_ = _1589_ | _1590_ /*15794*/;
  assign _1592_ = inv_10[20] ^ r_9[34] /*15792*/;
  assign sum_10[20] = _1592_ ^ _1591_ /*15791*/;
  assign _1593_ = _1592_ & _1591_ /*15790*/;
  assign _1594_ = inv_10[20] & r_9[34] /*15789*/;
  assign _1595_ = _1593_ | _1594_ /*15788*/;
  assign _1596_ = inv_10[21] ^ r_9[35] /*15786*/;
  assign sum_10[21] = _1596_ ^ _1595_ /*15785*/;
  assign _1597_ = _1596_ & _1595_ /*15784*/;
  assign _1598_ = inv_10[21] & r_9[35] /*15783*/;
  assign _1599_ = _1597_ | _1598_ /*15782*/;
  assign _1600_ = inv_10[22] ^ r_9[36] /*15780*/;
  assign sum_10[22] = _1600_ ^ _1599_ /*15779*/;
  assign _1601_ = _1600_ & _1599_ /*15778*/;
  assign _1602_ = inv_10[22] & r_9[36] /*15777*/;
  assign _1603_ = _1601_ | _1602_ /*15776*/;
  assign _1604_ = inv_10[23] ^ r_9[37] /*15774*/;
  assign sum_10[23] = _1604_ ^ _1603_ /*15773*/;
  assign _1605_ = _1604_ & _1603_ /*15772*/;
  assign _1606_ = inv_10[23] & r_9[37] /*15771*/;
  assign _1607_ = _1605_ | _1606_ /*15770*/;
  assign q[14] = ~sum_10[23] /*15789*/;
  assign m_10[0] = r_9[14] /*15788*/;
  assign m_10[1] = r_9[15] /*15787*/;
  assign m_10[2] = r_9[16] /*15786*/;
  assign m_10[3] = r_9[17] /*15785*/;
  assign m_10[4] = r_9[18] /*15784*/;
  assign m_10[5] = r_9[19] /*15783*/;
  assign m_10[6] = r_9[20] /*15782*/;
  assign m_10[7] = r_9[21] /*15781*/;
  assign m_10[8] = r_9[22] /*15780*/;
  assign m_10[9] = r_9[23] /*15779*/;
  assign m_10[10] = r_9[24] /*15778*/;
  assign m_10[11] = r_9[25] /*15777*/;
  assign m_10[12] = r_9[26] /*15776*/;
  assign m_10[13] = r_9[27] /*15775*/;
  assign m_10[14] = r_9[28] /*15774*/;
  assign m_10[15] = r_9[29] /*15773*/;
  assign m_10[16] = r_9[30] /*15772*/;
  assign m_10[17] = r_9[31] /*15771*/;
  assign m_10[18] = r_9[32] /*15770*/;
  assign m_10[19] = r_9[33] /*15769*/;
  assign m_10[20] = r_9[34] /*15768*/;
  assign m_10[21] = r_9[35] /*15767*/;
  assign m_10[22] = r_9[36] /*15766*/;
  assign m_10[23] = r_9[37] /*15765*/;
  assign _1608_ = ~q[14] /*15763*/;
  assign _1609_ = sum_10[0] & q[14] /*15762*/;
  assign _1610_ = m_10[0] & _1608_ /*15761*/;
  assign r_10[14] = _1610_ | _1609_ /*15760*/;
  assign _1611_ = ~q[14] /*15759*/;
  assign _1612_ = sum_10[1] & q[14] /*15758*/;
  assign _1613_ = m_10[1] & _1611_ /*15757*/;
  assign r_10[15] = _1613_ | _1612_ /*15756*/;
  assign _1614_ = ~q[14] /*15755*/;
  assign _1615_ = sum_10[2] & q[14] /*15754*/;
  assign _1616_ = m_10[2] & _1614_ /*15753*/;
  assign r_10[16] = _1616_ | _1615_ /*15752*/;
  assign _1617_ = ~q[14] /*15751*/;
  assign _1618_ = sum_10[3] & q[14] /*15750*/;
  assign _1619_ = m_10[3] & _1617_ /*15749*/;
  assign r_10[17] = _1619_ | _1618_ /*15748*/;
  assign _1620_ = ~q[14] /*15747*/;
  assign _1621_ = sum_10[4] & q[14] /*15746*/;
  assign _1622_ = m_10[4] & _1620_ /*15745*/;
  assign r_10[18] = _1622_ | _1621_ /*15744*/;
  assign _1623_ = ~q[14] /*15743*/;
  assign _1624_ = sum_10[5] & q[14] /*15742*/;
  assign _1625_ = m_10[5] & _1623_ /*15741*/;
  assign r_10[19] = _1625_ | _1624_ /*15740*/;
  assign _1626_ = ~q[14] /*15739*/;
  assign _1627_ = sum_10[6] & q[14] /*15738*/;
  assign _1628_ = m_10[6] & _1626_ /*15737*/;
  assign r_10[20] = _1628_ | _1627_ /*15736*/;
  assign _1629_ = ~q[14] /*15735*/;
  assign _1630_ = sum_10[7] & q[14] /*15734*/;
  assign _1631_ = m_10[7] & _1629_ /*15733*/;
  assign r_10[21] = _1631_ | _1630_ /*15732*/;
  assign _1632_ = ~q[14] /*15731*/;
  assign _1633_ = sum_10[8] & q[14] /*15730*/;
  assign _1634_ = m_10[8] & _1632_ /*15729*/;
  assign r_10[22] = _1634_ | _1633_ /*15728*/;
  assign _1635_ = ~q[14] /*15727*/;
  assign _1636_ = sum_10[9] & q[14] /*15726*/;
  assign _1637_ = m_10[9] & _1635_ /*15725*/;
  assign r_10[23] = _1637_ | _1636_ /*15724*/;
  assign _1638_ = ~q[14] /*15723*/;
  assign _1639_ = sum_10[10] & q[14] /*15722*/;
  assign _1640_ = m_10[10] & _1638_ /*15721*/;
  assign r_10[24] = _1640_ | _1639_ /*15720*/;
  assign _1641_ = ~q[14] /*15719*/;
  assign _1642_ = sum_10[11] & q[14] /*15718*/;
  assign _1643_ = m_10[11] & _1641_ /*15717*/;
  assign r_10[25] = _1643_ | _1642_ /*15716*/;
  assign _1644_ = ~q[14] /*15715*/;
  assign _1645_ = sum_10[12] & q[14] /*15714*/;
  assign _1646_ = m_10[12] & _1644_ /*15713*/;
  assign r_10[26] = _1646_ | _1645_ /*15712*/;
  assign _1647_ = ~q[14] /*15711*/;
  assign _1648_ = sum_10[13] & q[14] /*15710*/;
  assign _1649_ = m_10[13] & _1647_ /*15709*/;
  assign r_10[27] = _1649_ | _1648_ /*15708*/;
  assign _1650_ = ~q[14] /*15707*/;
  assign _1651_ = sum_10[14] & q[14] /*15706*/;
  assign _1652_ = m_10[14] & _1650_ /*15705*/;
  assign r_10[28] = _1652_ | _1651_ /*15704*/;
  assign _1653_ = ~q[14] /*15703*/;
  assign _1654_ = sum_10[15] & q[14] /*15702*/;
  assign _1655_ = m_10[15] & _1653_ /*15701*/;
  assign r_10[29] = _1655_ | _1654_ /*15700*/;
  assign _1656_ = ~q[14] /*15699*/;
  assign _1657_ = sum_10[16] & q[14] /*15698*/;
  assign _1658_ = m_10[16] & _1656_ /*15697*/;
  assign r_10[30] = _1658_ | _1657_ /*15696*/;
  assign _1659_ = ~q[14] /*15695*/;
  assign _1660_ = sum_10[17] & q[14] /*15694*/;
  assign _1661_ = m_10[17] & _1659_ /*15693*/;
  assign r_10[31] = _1661_ | _1660_ /*15692*/;
  assign _1662_ = ~q[14] /*15691*/;
  assign _1663_ = sum_10[18] & q[14] /*15690*/;
  assign _1664_ = m_10[18] & _1662_ /*15689*/;
  assign r_10[32] = _1664_ | _1663_ /*15688*/;
  assign _1665_ = ~q[14] /*15687*/;
  assign _1666_ = sum_10[19] & q[14] /*15686*/;
  assign _1667_ = m_10[19] & _1665_ /*15685*/;
  assign r_10[33] = _1667_ | _1666_ /*15684*/;
  assign _1668_ = ~q[14] /*15683*/;
  assign _1669_ = sum_10[20] & q[14] /*15682*/;
  assign _1670_ = m_10[20] & _1668_ /*15681*/;
  assign r_10[34] = _1670_ | _1669_ /*15680*/;
  assign _1671_ = ~q[14] /*15679*/;
  assign _1672_ = sum_10[21] & q[14] /*15678*/;
  assign _1673_ = m_10[21] & _1671_ /*15677*/;
  assign r_10[35] = _1673_ | _1672_ /*15676*/;
  assign _1674_ = ~q[14] /*15675*/;
  assign _1675_ = sum_10[22] & q[14] /*15674*/;
  assign _1676_ = m_10[22] & _1674_ /*15673*/;
  assign r_10[36] = _1676_ | _1675_ /*15672*/;
  assign _1677_ = ~q[14] /*15671*/;
  assign _1678_ = sum_10[23] & q[14] /*15670*/;
  assign _1679_ = m_10[23] & _1677_ /*15669*/;
  assign r_10[37] = _1679_ | _1678_ /*15668*/;
assign r_10[0]= r_9[0] /*15667*/;
assign r_10[1]= r_9[1] /*15666*/;
assign r_10[2]= r_9[2] /*15665*/;
assign r_10[3]= r_9[3] /*15664*/;
assign r_10[4]= r_9[4] /*15663*/;
assign r_10[5]= r_9[5] /*15662*/;
assign r_10[6]= r_9[6] /*15661*/;
assign r_10[7]= r_9[7] /*15660*/;
assign r_10[8]= r_9[8] /*15659*/;
assign r_10[9]= r_9[9] /*15658*/;
assign r_10[10]= r_9[10] /*15657*/;
assign r_10[11]= r_9[11] /*15656*/;
assign r_10[12]= r_9[12] /*15655*/;
assign r_10[13]= r_9[13] /*15654*/;
  assign inv_11[0] = ~div[0] /*15600*/;
  assign inv_11[1] = ~div[1] /*15599*/;
  assign inv_11[2] = ~div[2] /*15598*/;
  assign inv_11[3] = ~div[3] /*15597*/;
  assign inv_11[4] = ~div[4] /*15596*/;
  assign inv_11[5] = ~div[5] /*15595*/;
  assign inv_11[6] = ~div[6] /*15594*/;
  assign inv_11[7] = ~div[7] /*15593*/;
  assign inv_11[8] = ~div[8] /*15592*/;
  assign inv_11[9] = ~div[9] /*15591*/;
  assign inv_11[10] = ~div[10] /*15590*/;
  assign inv_11[11] = ~div[11] /*15589*/;
  assign inv_11[12] = ~div[12] /*15588*/;
  assign inv_11[13] = ~div[13] /*15587*/;
  assign inv_11[14] = ~div[14] /*15586*/;
  assign inv_11[15] = ~div[15] /*15585*/;
  assign inv_11[16] = ~div[16] /*15584*/;
  assign inv_11[17] = ~div[17] /*15583*/;
  assign inv_11[18] = ~div[18] /*15582*/;
  assign inv_11[19] = ~div[19] /*15581*/;
  assign inv_11[20] = ~div[20] /*15580*/;
  assign inv_11[21] = ~div[21] /*15579*/;
  assign inv_11[22] = ~div[22] /*15578*/;
assign inv_11[23] = oneWire /*15577*/;
  assign _1680_ = inv_11[0] ^ r_10[13] /*15575*/;
  assign sum_11[0] = _1680_ ^ oneWire /*15574*/;
  assign _1681_ = _1680_ & oneWire /*15573*/;
  assign _1682_ = inv_11[0] & r_10[13] /*15572*/;
  assign _1683_ = _1681_ | _1682_ /*15571*/;
  assign _1684_ = inv_11[1] ^ r_10[14] /*15570*/;
  assign sum_11[1] = _1684_ ^ _1683_ /*15569*/;
  assign _1685_ = _1684_ & _1683_ /*15568*/;
  assign _1686_ = inv_11[1] & r_10[14] /*15567*/;
  assign _1687_ = _1685_ | _1686_ /*15566*/;
  assign _1688_ = inv_11[2] ^ r_10[15] /*15564*/;
  assign sum_11[2] = _1688_ ^ _1687_ /*15563*/;
  assign _1689_ = _1688_ & _1687_ /*15562*/;
  assign _1690_ = inv_11[2] & r_10[15] /*15561*/;
  assign _1691_ = _1689_ | _1690_ /*15560*/;
  assign _1692_ = inv_11[3] ^ r_10[16] /*15558*/;
  assign sum_11[3] = _1692_ ^ _1691_ /*15557*/;
  assign _1693_ = _1692_ & _1691_ /*15556*/;
  assign _1694_ = inv_11[3] & r_10[16] /*15555*/;
  assign _1695_ = _1693_ | _1694_ /*15554*/;
  assign _1696_ = inv_11[4] ^ r_10[17] /*15552*/;
  assign sum_11[4] = _1696_ ^ _1695_ /*15551*/;
  assign _1697_ = _1696_ & _1695_ /*15550*/;
  assign _1698_ = inv_11[4] & r_10[17] /*15549*/;
  assign _1699_ = _1697_ | _1698_ /*15548*/;
  assign _1700_ = inv_11[5] ^ r_10[18] /*15546*/;
  assign sum_11[5] = _1700_ ^ _1699_ /*15545*/;
  assign _1701_ = _1700_ & _1699_ /*15544*/;
  assign _1702_ = inv_11[5] & r_10[18] /*15543*/;
  assign _1703_ = _1701_ | _1702_ /*15542*/;
  assign _1704_ = inv_11[6] ^ r_10[19] /*15540*/;
  assign sum_11[6] = _1704_ ^ _1703_ /*15539*/;
  assign _1705_ = _1704_ & _1703_ /*15538*/;
  assign _1706_ = inv_11[6] & r_10[19] /*15537*/;
  assign _1707_ = _1705_ | _1706_ /*15536*/;
  assign _1708_ = inv_11[7] ^ r_10[20] /*15534*/;
  assign sum_11[7] = _1708_ ^ _1707_ /*15533*/;
  assign _1709_ = _1708_ & _1707_ /*15532*/;
  assign _1710_ = inv_11[7] & r_10[20] /*15531*/;
  assign _1711_ = _1709_ | _1710_ /*15530*/;
  assign _1712_ = inv_11[8] ^ r_10[21] /*15528*/;
  assign sum_11[8] = _1712_ ^ _1711_ /*15527*/;
  assign _1713_ = _1712_ & _1711_ /*15526*/;
  assign _1714_ = inv_11[8] & r_10[21] /*15525*/;
  assign _1715_ = _1713_ | _1714_ /*15524*/;
  assign _1716_ = inv_11[9] ^ r_10[22] /*15522*/;
  assign sum_11[9] = _1716_ ^ _1715_ /*15521*/;
  assign _1717_ = _1716_ & _1715_ /*15520*/;
  assign _1718_ = inv_11[9] & r_10[22] /*15519*/;
  assign _1719_ = _1717_ | _1718_ /*15518*/;
  assign _1720_ = inv_11[10] ^ r_10[23] /*15516*/;
  assign sum_11[10] = _1720_ ^ _1719_ /*15515*/;
  assign _1721_ = _1720_ & _1719_ /*15514*/;
  assign _1722_ = inv_11[10] & r_10[23] /*15513*/;
  assign _1723_ = _1721_ | _1722_ /*15512*/;
  assign _1724_ = inv_11[11] ^ r_10[24] /*15510*/;
  assign sum_11[11] = _1724_ ^ _1723_ /*15509*/;
  assign _1725_ = _1724_ & _1723_ /*15508*/;
  assign _1726_ = inv_11[11] & r_10[24] /*15507*/;
  assign _1727_ = _1725_ | _1726_ /*15506*/;
  assign _1728_ = inv_11[12] ^ r_10[25] /*15504*/;
  assign sum_11[12] = _1728_ ^ _1727_ /*15503*/;
  assign _1729_ = _1728_ & _1727_ /*15502*/;
  assign _1730_ = inv_11[12] & r_10[25] /*15501*/;
  assign _1731_ = _1729_ | _1730_ /*15500*/;
  assign _1732_ = inv_11[13] ^ r_10[26] /*15498*/;
  assign sum_11[13] = _1732_ ^ _1731_ /*15497*/;
  assign _1733_ = _1732_ & _1731_ /*15496*/;
  assign _1734_ = inv_11[13] & r_10[26] /*15495*/;
  assign _1735_ = _1733_ | _1734_ /*15494*/;
  assign _1736_ = inv_11[14] ^ r_10[27] /*15492*/;
  assign sum_11[14] = _1736_ ^ _1735_ /*15491*/;
  assign _1737_ = _1736_ & _1735_ /*15490*/;
  assign _1738_ = inv_11[14] & r_10[27] /*15489*/;
  assign _1739_ = _1737_ | _1738_ /*15488*/;
  assign _1740_ = inv_11[15] ^ r_10[28] /*15486*/;
  assign sum_11[15] = _1740_ ^ _1739_ /*15485*/;
  assign _1741_ = _1740_ & _1739_ /*15484*/;
  assign _1742_ = inv_11[15] & r_10[28] /*15483*/;
  assign _1743_ = _1741_ | _1742_ /*15482*/;
  assign _1744_ = inv_11[16] ^ r_10[29] /*15480*/;
  assign sum_11[16] = _1744_ ^ _1743_ /*15479*/;
  assign _1745_ = _1744_ & _1743_ /*15478*/;
  assign _1746_ = inv_11[16] & r_10[29] /*15477*/;
  assign _1747_ = _1745_ | _1746_ /*15476*/;
  assign _1748_ = inv_11[17] ^ r_10[30] /*15474*/;
  assign sum_11[17] = _1748_ ^ _1747_ /*15473*/;
  assign _1749_ = _1748_ & _1747_ /*15472*/;
  assign _1750_ = inv_11[17] & r_10[30] /*15471*/;
  assign _1751_ = _1749_ | _1750_ /*15470*/;
  assign _1752_ = inv_11[18] ^ r_10[31] /*15468*/;
  assign sum_11[18] = _1752_ ^ _1751_ /*15467*/;
  assign _1753_ = _1752_ & _1751_ /*15466*/;
  assign _1754_ = inv_11[18] & r_10[31] /*15465*/;
  assign _1755_ = _1753_ | _1754_ /*15464*/;
  assign _1756_ = inv_11[19] ^ r_10[32] /*15462*/;
  assign sum_11[19] = _1756_ ^ _1755_ /*15461*/;
  assign _1757_ = _1756_ & _1755_ /*15460*/;
  assign _1758_ = inv_11[19] & r_10[32] /*15459*/;
  assign _1759_ = _1757_ | _1758_ /*15458*/;
  assign _1760_ = inv_11[20] ^ r_10[33] /*15456*/;
  assign sum_11[20] = _1760_ ^ _1759_ /*15455*/;
  assign _1761_ = _1760_ & _1759_ /*15454*/;
  assign _1762_ = inv_11[20] & r_10[33] /*15453*/;
  assign _1763_ = _1761_ | _1762_ /*15452*/;
  assign _1764_ = inv_11[21] ^ r_10[34] /*15450*/;
  assign sum_11[21] = _1764_ ^ _1763_ /*15449*/;
  assign _1765_ = _1764_ & _1763_ /*15448*/;
  assign _1766_ = inv_11[21] & r_10[34] /*15447*/;
  assign _1767_ = _1765_ | _1766_ /*15446*/;
  assign _1768_ = inv_11[22] ^ r_10[35] /*15444*/;
  assign sum_11[22] = _1768_ ^ _1767_ /*15443*/;
  assign _1769_ = _1768_ & _1767_ /*15442*/;
  assign _1770_ = inv_11[22] & r_10[35] /*15441*/;
  assign _1771_ = _1769_ | _1770_ /*15440*/;
  assign _1772_ = inv_11[23] ^ r_10[36] /*15438*/;
  assign sum_11[23] = _1772_ ^ _1771_ /*15437*/;
  assign _1773_ = _1772_ & _1771_ /*15436*/;
  assign _1774_ = inv_11[23] & r_10[36] /*15435*/;
  assign _1775_ = _1773_ | _1774_ /*15434*/;
  assign q[13] = ~sum_11[23] /*15453*/;
  assign m_11[0] = r_10[13] /*15452*/;
  assign m_11[1] = r_10[14] /*15451*/;
  assign m_11[2] = r_10[15] /*15450*/;
  assign m_11[3] = r_10[16] /*15449*/;
  assign m_11[4] = r_10[17] /*15448*/;
  assign m_11[5] = r_10[18] /*15447*/;
  assign m_11[6] = r_10[19] /*15446*/;
  assign m_11[7] = r_10[20] /*15445*/;
  assign m_11[8] = r_10[21] /*15444*/;
  assign m_11[9] = r_10[22] /*15443*/;
  assign m_11[10] = r_10[23] /*15442*/;
  assign m_11[11] = r_10[24] /*15441*/;
  assign m_11[12] = r_10[25] /*15440*/;
  assign m_11[13] = r_10[26] /*15439*/;
  assign m_11[14] = r_10[27] /*15438*/;
  assign m_11[15] = r_10[28] /*15437*/;
  assign m_11[16] = r_10[29] /*15436*/;
  assign m_11[17] = r_10[30] /*15435*/;
  assign m_11[18] = r_10[31] /*15434*/;
  assign m_11[19] = r_10[32] /*15433*/;
  assign m_11[20] = r_10[33] /*15432*/;
  assign m_11[21] = r_10[34] /*15431*/;
  assign m_11[22] = r_10[35] /*15430*/;
  assign m_11[23] = r_10[36] /*15429*/;
  assign _1776_ = ~q[13] /*15427*/;
  assign _1777_ = sum_11[0] & q[13] /*15426*/;
  assign _1778_ = m_11[0] & _1776_ /*15425*/;
  assign r_11[13] = _1778_ | _1777_ /*15424*/;
  assign _1779_ = ~q[13] /*15423*/;
  assign _1780_ = sum_11[1] & q[13] /*15422*/;
  assign _1781_ = m_11[1] & _1779_ /*15421*/;
  assign r_11[14] = _1781_ | _1780_ /*15420*/;
  assign _1782_ = ~q[13] /*15419*/;
  assign _1783_ = sum_11[2] & q[13] /*15418*/;
  assign _1784_ = m_11[2] & _1782_ /*15417*/;
  assign r_11[15] = _1784_ | _1783_ /*15416*/;
  assign _1785_ = ~q[13] /*15415*/;
  assign _1786_ = sum_11[3] & q[13] /*15414*/;
  assign _1787_ = m_11[3] & _1785_ /*15413*/;
  assign r_11[16] = _1787_ | _1786_ /*15412*/;
  assign _1788_ = ~q[13] /*15411*/;
  assign _1789_ = sum_11[4] & q[13] /*15410*/;
  assign _1790_ = m_11[4] & _1788_ /*15409*/;
  assign r_11[17] = _1790_ | _1789_ /*15408*/;
  assign _1791_ = ~q[13] /*15407*/;
  assign _1792_ = sum_11[5] & q[13] /*15406*/;
  assign _1793_ = m_11[5] & _1791_ /*15405*/;
  assign r_11[18] = _1793_ | _1792_ /*15404*/;
  assign _1794_ = ~q[13] /*15403*/;
  assign _1795_ = sum_11[6] & q[13] /*15402*/;
  assign _1796_ = m_11[6] & _1794_ /*15401*/;
  assign r_11[19] = _1796_ | _1795_ /*15400*/;
  assign _1797_ = ~q[13] /*15399*/;
  assign _1798_ = sum_11[7] & q[13] /*15398*/;
  assign _1799_ = m_11[7] & _1797_ /*15397*/;
  assign r_11[20] = _1799_ | _1798_ /*15396*/;
  assign _1800_ = ~q[13] /*15395*/;
  assign _1801_ = sum_11[8] & q[13] /*15394*/;
  assign _1802_ = m_11[8] & _1800_ /*15393*/;
  assign r_11[21] = _1802_ | _1801_ /*15392*/;
  assign _1803_ = ~q[13] /*15391*/;
  assign _1804_ = sum_11[9] & q[13] /*15390*/;
  assign _1805_ = m_11[9] & _1803_ /*15389*/;
  assign r_11[22] = _1805_ | _1804_ /*15388*/;
  assign _1806_ = ~q[13] /*15387*/;
  assign _1807_ = sum_11[10] & q[13] /*15386*/;
  assign _1808_ = m_11[10] & _1806_ /*15385*/;
  assign r_11[23] = _1808_ | _1807_ /*15384*/;
  assign _1809_ = ~q[13] /*15383*/;
  assign _1810_ = sum_11[11] & q[13] /*15382*/;
  assign _1811_ = m_11[11] & _1809_ /*15381*/;
  assign r_11[24] = _1811_ | _1810_ /*15380*/;
  assign _1812_ = ~q[13] /*15379*/;
  assign _1813_ = sum_11[12] & q[13] /*15378*/;
  assign _1814_ = m_11[12] & _1812_ /*15377*/;
  assign r_11[25] = _1814_ | _1813_ /*15376*/;
  assign _1815_ = ~q[13] /*15375*/;
  assign _1816_ = sum_11[13] & q[13] /*15374*/;
  assign _1817_ = m_11[13] & _1815_ /*15373*/;
  assign r_11[26] = _1817_ | _1816_ /*15372*/;
  assign _1818_ = ~q[13] /*15371*/;
  assign _1819_ = sum_11[14] & q[13] /*15370*/;
  assign _1820_ = m_11[14] & _1818_ /*15369*/;
  assign r_11[27] = _1820_ | _1819_ /*15368*/;
  assign _1821_ = ~q[13] /*15367*/;
  assign _1822_ = sum_11[15] & q[13] /*15366*/;
  assign _1823_ = m_11[15] & _1821_ /*15365*/;
  assign r_11[28] = _1823_ | _1822_ /*15364*/;
  assign _1824_ = ~q[13] /*15363*/;
  assign _1825_ = sum_11[16] & q[13] /*15362*/;
  assign _1826_ = m_11[16] & _1824_ /*15361*/;
  assign r_11[29] = _1826_ | _1825_ /*15360*/;
  assign _1827_ = ~q[13] /*15359*/;
  assign _1828_ = sum_11[17] & q[13] /*15358*/;
  assign _1829_ = m_11[17] & _1827_ /*15357*/;
  assign r_11[30] = _1829_ | _1828_ /*15356*/;
  assign _1830_ = ~q[13] /*15355*/;
  assign _1831_ = sum_11[18] & q[13] /*15354*/;
  assign _1832_ = m_11[18] & _1830_ /*15353*/;
  assign r_11[31] = _1832_ | _1831_ /*15352*/;
  assign _1833_ = ~q[13] /*15351*/;
  assign _1834_ = sum_11[19] & q[13] /*15350*/;
  assign _1835_ = m_11[19] & _1833_ /*15349*/;
  assign r_11[32] = _1835_ | _1834_ /*15348*/;
  assign _1836_ = ~q[13] /*15347*/;
  assign _1837_ = sum_11[20] & q[13] /*15346*/;
  assign _1838_ = m_11[20] & _1836_ /*15345*/;
  assign r_11[33] = _1838_ | _1837_ /*15344*/;
  assign _1839_ = ~q[13] /*15343*/;
  assign _1840_ = sum_11[21] & q[13] /*15342*/;
  assign _1841_ = m_11[21] & _1839_ /*15341*/;
  assign r_11[34] = _1841_ | _1840_ /*15340*/;
  assign _1842_ = ~q[13] /*15339*/;
  assign _1843_ = sum_11[22] & q[13] /*15338*/;
  assign _1844_ = m_11[22] & _1842_ /*15337*/;
  assign r_11[35] = _1844_ | _1843_ /*15336*/;
  assign _1845_ = ~q[13] /*15335*/;
  assign _1846_ = sum_11[23] & q[13] /*15334*/;
  assign _1847_ = m_11[23] & _1845_ /*15333*/;
  assign r_11[36] = _1847_ | _1846_ /*15332*/;
assign r_11[0]= r_10[0] /*15331*/;
assign r_11[1]= r_10[1] /*15330*/;
assign r_11[2]= r_10[2] /*15329*/;
assign r_11[3]= r_10[3] /*15328*/;
assign r_11[4]= r_10[4] /*15327*/;
assign r_11[5]= r_10[5] /*15326*/;
assign r_11[6]= r_10[6] /*15325*/;
assign r_11[7]= r_10[7] /*15324*/;
assign r_11[8]= r_10[8] /*15323*/;
assign r_11[9]= r_10[9] /*15322*/;
assign r_11[10]= r_10[10] /*15321*/;
assign r_11[11]= r_10[11] /*15320*/;
assign r_11[12]= r_10[12] /*15319*/;
  assign inv_12[0] = ~div[0] /*15264*/;
  assign inv_12[1] = ~div[1] /*15263*/;
  assign inv_12[2] = ~div[2] /*15262*/;
  assign inv_12[3] = ~div[3] /*15261*/;
  assign inv_12[4] = ~div[4] /*15260*/;
  assign inv_12[5] = ~div[5] /*15259*/;
  assign inv_12[6] = ~div[6] /*15258*/;
  assign inv_12[7] = ~div[7] /*15257*/;
  assign inv_12[8] = ~div[8] /*15256*/;
  assign inv_12[9] = ~div[9] /*15255*/;
  assign inv_12[10] = ~div[10] /*15254*/;
  assign inv_12[11] = ~div[11] /*15253*/;
  assign inv_12[12] = ~div[12] /*15252*/;
  assign inv_12[13] = ~div[13] /*15251*/;
  assign inv_12[14] = ~div[14] /*15250*/;
  assign inv_12[15] = ~div[15] /*15249*/;
  assign inv_12[16] = ~div[16] /*15248*/;
  assign inv_12[17] = ~div[17] /*15247*/;
  assign inv_12[18] = ~div[18] /*15246*/;
  assign inv_12[19] = ~div[19] /*15245*/;
  assign inv_12[20] = ~div[20] /*15244*/;
  assign inv_12[21] = ~div[21] /*15243*/;
  assign inv_12[22] = ~div[22] /*15242*/;
assign inv_12[23] = oneWire /*15241*/;
  assign _1848_ = inv_12[0] ^ r_11[12] /*15239*/;
  assign sum_12[0] = _1848_ ^ oneWire /*15238*/;
  assign _1849_ = _1848_ & oneWire /*15237*/;
  assign _1850_ = inv_12[0] & r_11[12] /*15236*/;
  assign _1851_ = _1849_ | _1850_ /*15235*/;
  assign _1852_ = inv_12[1] ^ r_11[13] /*15234*/;
  assign sum_12[1] = _1852_ ^ _1851_ /*15233*/;
  assign _1853_ = _1852_ & _1851_ /*15232*/;
  assign _1854_ = inv_12[1] & r_11[13] /*15231*/;
  assign _1855_ = _1853_ | _1854_ /*15230*/;
  assign _1856_ = inv_12[2] ^ r_11[14] /*15228*/;
  assign sum_12[2] = _1856_ ^ _1855_ /*15227*/;
  assign _1857_ = _1856_ & _1855_ /*15226*/;
  assign _1858_ = inv_12[2] & r_11[14] /*15225*/;
  assign _1859_ = _1857_ | _1858_ /*15224*/;
  assign _1860_ = inv_12[3] ^ r_11[15] /*15222*/;
  assign sum_12[3] = _1860_ ^ _1859_ /*15221*/;
  assign _1861_ = _1860_ & _1859_ /*15220*/;
  assign _1862_ = inv_12[3] & r_11[15] /*15219*/;
  assign _1863_ = _1861_ | _1862_ /*15218*/;
  assign _1864_ = inv_12[4] ^ r_11[16] /*15216*/;
  assign sum_12[4] = _1864_ ^ _1863_ /*15215*/;
  assign _1865_ = _1864_ & _1863_ /*15214*/;
  assign _1866_ = inv_12[4] & r_11[16] /*15213*/;
  assign _1867_ = _1865_ | _1866_ /*15212*/;
  assign _1868_ = inv_12[5] ^ r_11[17] /*15210*/;
  assign sum_12[5] = _1868_ ^ _1867_ /*15209*/;
  assign _1869_ = _1868_ & _1867_ /*15208*/;
  assign _1870_ = inv_12[5] & r_11[17] /*15207*/;
  assign _1871_ = _1869_ | _1870_ /*15206*/;
  assign _1872_ = inv_12[6] ^ r_11[18] /*15204*/;
  assign sum_12[6] = _1872_ ^ _1871_ /*15203*/;
  assign _1873_ = _1872_ & _1871_ /*15202*/;
  assign _1874_ = inv_12[6] & r_11[18] /*15201*/;
  assign _1875_ = _1873_ | _1874_ /*15200*/;
  assign _1876_ = inv_12[7] ^ r_11[19] /*15198*/;
  assign sum_12[7] = _1876_ ^ _1875_ /*15197*/;
  assign _1877_ = _1876_ & _1875_ /*15196*/;
  assign _1878_ = inv_12[7] & r_11[19] /*15195*/;
  assign _1879_ = _1877_ | _1878_ /*15194*/;
  assign _1880_ = inv_12[8] ^ r_11[20] /*15192*/;
  assign sum_12[8] = _1880_ ^ _1879_ /*15191*/;
  assign _1881_ = _1880_ & _1879_ /*15190*/;
  assign _1882_ = inv_12[8] & r_11[20] /*15189*/;
  assign _1883_ = _1881_ | _1882_ /*15188*/;
  assign _1884_ = inv_12[9] ^ r_11[21] /*15186*/;
  assign sum_12[9] = _1884_ ^ _1883_ /*15185*/;
  assign _1885_ = _1884_ & _1883_ /*15184*/;
  assign _1886_ = inv_12[9] & r_11[21] /*15183*/;
  assign _1887_ = _1885_ | _1886_ /*15182*/;
  assign _1888_ = inv_12[10] ^ r_11[22] /*15180*/;
  assign sum_12[10] = _1888_ ^ _1887_ /*15179*/;
  assign _1889_ = _1888_ & _1887_ /*15178*/;
  assign _1890_ = inv_12[10] & r_11[22] /*15177*/;
  assign _1891_ = _1889_ | _1890_ /*15176*/;
  assign _1892_ = inv_12[11] ^ r_11[23] /*15174*/;
  assign sum_12[11] = _1892_ ^ _1891_ /*15173*/;
  assign _1893_ = _1892_ & _1891_ /*15172*/;
  assign _1894_ = inv_12[11] & r_11[23] /*15171*/;
  assign _1895_ = _1893_ | _1894_ /*15170*/;
  assign _1896_ = inv_12[12] ^ r_11[24] /*15168*/;
  assign sum_12[12] = _1896_ ^ _1895_ /*15167*/;
  assign _1897_ = _1896_ & _1895_ /*15166*/;
  assign _1898_ = inv_12[12] & r_11[24] /*15165*/;
  assign _1899_ = _1897_ | _1898_ /*15164*/;
  assign _1900_ = inv_12[13] ^ r_11[25] /*15162*/;
  assign sum_12[13] = _1900_ ^ _1899_ /*15161*/;
  assign _1901_ = _1900_ & _1899_ /*15160*/;
  assign _1902_ = inv_12[13] & r_11[25] /*15159*/;
  assign _1903_ = _1901_ | _1902_ /*15158*/;
  assign _1904_ = inv_12[14] ^ r_11[26] /*15156*/;
  assign sum_12[14] = _1904_ ^ _1903_ /*15155*/;
  assign _1905_ = _1904_ & _1903_ /*15154*/;
  assign _1906_ = inv_12[14] & r_11[26] /*15153*/;
  assign _1907_ = _1905_ | _1906_ /*15152*/;
  assign _1908_ = inv_12[15] ^ r_11[27] /*15150*/;
  assign sum_12[15] = _1908_ ^ _1907_ /*15149*/;
  assign _1909_ = _1908_ & _1907_ /*15148*/;
  assign _1910_ = inv_12[15] & r_11[27] /*15147*/;
  assign _1911_ = _1909_ | _1910_ /*15146*/;
  assign _1912_ = inv_12[16] ^ r_11[28] /*15144*/;
  assign sum_12[16] = _1912_ ^ _1911_ /*15143*/;
  assign _1913_ = _1912_ & _1911_ /*15142*/;
  assign _1914_ = inv_12[16] & r_11[28] /*15141*/;
  assign _1915_ = _1913_ | _1914_ /*15140*/;
  assign _1916_ = inv_12[17] ^ r_11[29] /*15138*/;
  assign sum_12[17] = _1916_ ^ _1915_ /*15137*/;
  assign _1917_ = _1916_ & _1915_ /*15136*/;
  assign _1918_ = inv_12[17] & r_11[29] /*15135*/;
  assign _1919_ = _1917_ | _1918_ /*15134*/;
  assign _1920_ = inv_12[18] ^ r_11[30] /*15132*/;
  assign sum_12[18] = _1920_ ^ _1919_ /*15131*/;
  assign _1921_ = _1920_ & _1919_ /*15130*/;
  assign _1922_ = inv_12[18] & r_11[30] /*15129*/;
  assign _1923_ = _1921_ | _1922_ /*15128*/;
  assign _1924_ = inv_12[19] ^ r_11[31] /*15126*/;
  assign sum_12[19] = _1924_ ^ _1923_ /*15125*/;
  assign _1925_ = _1924_ & _1923_ /*15124*/;
  assign _1926_ = inv_12[19] & r_11[31] /*15123*/;
  assign _1927_ = _1925_ | _1926_ /*15122*/;
  assign _1928_ = inv_12[20] ^ r_11[32] /*15120*/;
  assign sum_12[20] = _1928_ ^ _1927_ /*15119*/;
  assign _1929_ = _1928_ & _1927_ /*15118*/;
  assign _1930_ = inv_12[20] & r_11[32] /*15117*/;
  assign _1931_ = _1929_ | _1930_ /*15116*/;
  assign _1932_ = inv_12[21] ^ r_11[33] /*15114*/;
  assign sum_12[21] = _1932_ ^ _1931_ /*15113*/;
  assign _1933_ = _1932_ & _1931_ /*15112*/;
  assign _1934_ = inv_12[21] & r_11[33] /*15111*/;
  assign _1935_ = _1933_ | _1934_ /*15110*/;
  assign _1936_ = inv_12[22] ^ r_11[34] /*15108*/;
  assign sum_12[22] = _1936_ ^ _1935_ /*15107*/;
  assign _1937_ = _1936_ & _1935_ /*15106*/;
  assign _1938_ = inv_12[22] & r_11[34] /*15105*/;
  assign _1939_ = _1937_ | _1938_ /*15104*/;
  assign _1940_ = inv_12[23] ^ r_11[35] /*15102*/;
  assign sum_12[23] = _1940_ ^ _1939_ /*15101*/;
  assign _1941_ = _1940_ & _1939_ /*15100*/;
  assign _1942_ = inv_12[23] & r_11[35] /*15099*/;
  assign _1943_ = _1941_ | _1942_ /*15098*/;
  assign q[12] = ~sum_12[23] /*15117*/;
  assign m_12[0] = r_11[12] /*15116*/;
  assign m_12[1] = r_11[13] /*15115*/;
  assign m_12[2] = r_11[14] /*15114*/;
  assign m_12[3] = r_11[15] /*15113*/;
  assign m_12[4] = r_11[16] /*15112*/;
  assign m_12[5] = r_11[17] /*15111*/;
  assign m_12[6] = r_11[18] /*15110*/;
  assign m_12[7] = r_11[19] /*15109*/;
  assign m_12[8] = r_11[20] /*15108*/;
  assign m_12[9] = r_11[21] /*15107*/;
  assign m_12[10] = r_11[22] /*15106*/;
  assign m_12[11] = r_11[23] /*15105*/;
  assign m_12[12] = r_11[24] /*15104*/;
  assign m_12[13] = r_11[25] /*15103*/;
  assign m_12[14] = r_11[26] /*15102*/;
  assign m_12[15] = r_11[27] /*15101*/;
  assign m_12[16] = r_11[28] /*15100*/;
  assign m_12[17] = r_11[29] /*15099*/;
  assign m_12[18] = r_11[30] /*15098*/;
  assign m_12[19] = r_11[31] /*15097*/;
  assign m_12[20] = r_11[32] /*15096*/;
  assign m_12[21] = r_11[33] /*15095*/;
  assign m_12[22] = r_11[34] /*15094*/;
  assign m_12[23] = r_11[35] /*15093*/;
  assign _1944_ = ~q[12] /*15091*/;
  assign _1945_ = sum_12[0] & q[12] /*15090*/;
  assign _1946_ = m_12[0] & _1944_ /*15089*/;
  assign r_12[12] = _1946_ | _1945_ /*15088*/;
  assign _1947_ = ~q[12] /*15087*/;
  assign _1948_ = sum_12[1] & q[12] /*15086*/;
  assign _1949_ = m_12[1] & _1947_ /*15085*/;
  assign r_12[13] = _1949_ | _1948_ /*15084*/;
  assign _1950_ = ~q[12] /*15083*/;
  assign _1951_ = sum_12[2] & q[12] /*15082*/;
  assign _1952_ = m_12[2] & _1950_ /*15081*/;
  assign r_12[14] = _1952_ | _1951_ /*15080*/;
  assign _1953_ = ~q[12] /*15079*/;
  assign _1954_ = sum_12[3] & q[12] /*15078*/;
  assign _1955_ = m_12[3] & _1953_ /*15077*/;
  assign r_12[15] = _1955_ | _1954_ /*15076*/;
  assign _1956_ = ~q[12] /*15075*/;
  assign _1957_ = sum_12[4] & q[12] /*15074*/;
  assign _1958_ = m_12[4] & _1956_ /*15073*/;
  assign r_12[16] = _1958_ | _1957_ /*15072*/;
  assign _1959_ = ~q[12] /*15071*/;
  assign _1960_ = sum_12[5] & q[12] /*15070*/;
  assign _1961_ = m_12[5] & _1959_ /*15069*/;
  assign r_12[17] = _1961_ | _1960_ /*15068*/;
  assign _1962_ = ~q[12] /*15067*/;
  assign _1963_ = sum_12[6] & q[12] /*15066*/;
  assign _1964_ = m_12[6] & _1962_ /*15065*/;
  assign r_12[18] = _1964_ | _1963_ /*15064*/;
  assign _1965_ = ~q[12] /*15063*/;
  assign _1966_ = sum_12[7] & q[12] /*15062*/;
  assign _1967_ = m_12[7] & _1965_ /*15061*/;
  assign r_12[19] = _1967_ | _1966_ /*15060*/;
  assign _1968_ = ~q[12] /*15059*/;
  assign _1969_ = sum_12[8] & q[12] /*15058*/;
  assign _1970_ = m_12[8] & _1968_ /*15057*/;
  assign r_12[20] = _1970_ | _1969_ /*15056*/;
  assign _1971_ = ~q[12] /*15055*/;
  assign _1972_ = sum_12[9] & q[12] /*15054*/;
  assign _1973_ = m_12[9] & _1971_ /*15053*/;
  assign r_12[21] = _1973_ | _1972_ /*15052*/;
  assign _1974_ = ~q[12] /*15051*/;
  assign _1975_ = sum_12[10] & q[12] /*15050*/;
  assign _1976_ = m_12[10] & _1974_ /*15049*/;
  assign r_12[22] = _1976_ | _1975_ /*15048*/;
  assign _1977_ = ~q[12] /*15047*/;
  assign _1978_ = sum_12[11] & q[12] /*15046*/;
  assign _1979_ = m_12[11] & _1977_ /*15045*/;
  assign r_12[23] = _1979_ | _1978_ /*15044*/;
  assign _1980_ = ~q[12] /*15043*/;
  assign _1981_ = sum_12[12] & q[12] /*15042*/;
  assign _1982_ = m_12[12] & _1980_ /*15041*/;
  assign r_12[24] = _1982_ | _1981_ /*15040*/;
  assign _1983_ = ~q[12] /*15039*/;
  assign _1984_ = sum_12[13] & q[12] /*15038*/;
  assign _1985_ = m_12[13] & _1983_ /*15037*/;
  assign r_12[25] = _1985_ | _1984_ /*15036*/;
  assign _1986_ = ~q[12] /*15035*/;
  assign _1987_ = sum_12[14] & q[12] /*15034*/;
  assign _1988_ = m_12[14] & _1986_ /*15033*/;
  assign r_12[26] = _1988_ | _1987_ /*15032*/;
  assign _1989_ = ~q[12] /*15031*/;
  assign _1990_ = sum_12[15] & q[12] /*15030*/;
  assign _1991_ = m_12[15] & _1989_ /*15029*/;
  assign r_12[27] = _1991_ | _1990_ /*15028*/;
  assign _1992_ = ~q[12] /*15027*/;
  assign _1993_ = sum_12[16] & q[12] /*15026*/;
  assign _1994_ = m_12[16] & _1992_ /*15025*/;
  assign r_12[28] = _1994_ | _1993_ /*15024*/;
  assign _1995_ = ~q[12] /*15023*/;
  assign _1996_ = sum_12[17] & q[12] /*15022*/;
  assign _1997_ = m_12[17] & _1995_ /*15021*/;
  assign r_12[29] = _1997_ | _1996_ /*15020*/;
  assign _1998_ = ~q[12] /*15019*/;
  assign _1999_ = sum_12[18] & q[12] /*15018*/;
  assign _2000_ = m_12[18] & _1998_ /*15017*/;
  assign r_12[30] = _2000_ | _1999_ /*15016*/;
  assign _2001_ = ~q[12] /*15015*/;
  assign _2002_ = sum_12[19] & q[12] /*15014*/;
  assign _2003_ = m_12[19] & _2001_ /*15013*/;
  assign r_12[31] = _2003_ | _2002_ /*15012*/;
  assign _2004_ = ~q[12] /*15011*/;
  assign _2005_ = sum_12[20] & q[12] /*15010*/;
  assign _2006_ = m_12[20] & _2004_ /*15009*/;
  assign r_12[32] = _2006_ | _2005_ /*15008*/;
  assign _2007_ = ~q[12] /*15007*/;
  assign _2008_ = sum_12[21] & q[12] /*15006*/;
  assign _2009_ = m_12[21] & _2007_ /*15005*/;
  assign r_12[33] = _2009_ | _2008_ /*15004*/;
  assign _2010_ = ~q[12] /*15003*/;
  assign _2011_ = sum_12[22] & q[12] /*15002*/;
  assign _2012_ = m_12[22] & _2010_ /*15001*/;
  assign r_12[34] = _2012_ | _2011_ /*15000*/;
  assign _2013_ = ~q[12] /*14999*/;
  assign _2014_ = sum_12[23] & q[12] /*14998*/;
  assign _2015_ = m_12[23] & _2013_ /*14997*/;
  assign r_12[35] = _2015_ | _2014_ /*14996*/;
assign r_12[0]= r_11[0] /*14995*/;
assign r_12[1]= r_11[1] /*14994*/;
assign r_12[2]= r_11[2] /*14993*/;
assign r_12[3]= r_11[3] /*14992*/;
assign r_12[4]= r_11[4] /*14991*/;
assign r_12[5]= r_11[5] /*14990*/;
assign r_12[6]= r_11[6] /*14989*/;
assign r_12[7]= r_11[7] /*14988*/;
assign r_12[8]= r_11[8] /*14987*/;
assign r_12[9]= r_11[9] /*14986*/;
assign r_12[10]= r_11[10] /*14985*/;
assign r_12[11]= r_11[11] /*14984*/;
  assign inv_13[0] = ~div[0] /*14928*/;
  assign inv_13[1] = ~div[1] /*14927*/;
  assign inv_13[2] = ~div[2] /*14926*/;
  assign inv_13[3] = ~div[3] /*14925*/;
  assign inv_13[4] = ~div[4] /*14924*/;
  assign inv_13[5] = ~div[5] /*14923*/;
  assign inv_13[6] = ~div[6] /*14922*/;
  assign inv_13[7] = ~div[7] /*14921*/;
  assign inv_13[8] = ~div[8] /*14920*/;
  assign inv_13[9] = ~div[9] /*14919*/;
  assign inv_13[10] = ~div[10] /*14918*/;
  assign inv_13[11] = ~div[11] /*14917*/;
  assign inv_13[12] = ~div[12] /*14916*/;
  assign inv_13[13] = ~div[13] /*14915*/;
  assign inv_13[14] = ~div[14] /*14914*/;
  assign inv_13[15] = ~div[15] /*14913*/;
  assign inv_13[16] = ~div[16] /*14912*/;
  assign inv_13[17] = ~div[17] /*14911*/;
  assign inv_13[18] = ~div[18] /*14910*/;
  assign inv_13[19] = ~div[19] /*14909*/;
  assign inv_13[20] = ~div[20] /*14908*/;
  assign inv_13[21] = ~div[21] /*14907*/;
  assign inv_13[22] = ~div[22] /*14906*/;
assign inv_13[23] = oneWire /*14905*/;
  assign _2016_ = inv_13[0] ^ r_12[11] /*14903*/;
  assign sum_13[0] = _2016_ ^ oneWire /*14902*/;
  assign _2017_ = _2016_ & oneWire /*14901*/;
  assign _2018_ = inv_13[0] & r_12[11] /*14900*/;
  assign _2019_ = _2017_ | _2018_ /*14899*/;
  assign _2020_ = inv_13[1] ^ r_12[12] /*14898*/;
  assign sum_13[1] = _2020_ ^ _2019_ /*14897*/;
  assign _2021_ = _2020_ & _2019_ /*14896*/;
  assign _2022_ = inv_13[1] & r_12[12] /*14895*/;
  assign _2023_ = _2021_ | _2022_ /*14894*/;
  assign _2024_ = inv_13[2] ^ r_12[13] /*14892*/;
  assign sum_13[2] = _2024_ ^ _2023_ /*14891*/;
  assign _2025_ = _2024_ & _2023_ /*14890*/;
  assign _2026_ = inv_13[2] & r_12[13] /*14889*/;
  assign _2027_ = _2025_ | _2026_ /*14888*/;
  assign _2028_ = inv_13[3] ^ r_12[14] /*14886*/;
  assign sum_13[3] = _2028_ ^ _2027_ /*14885*/;
  assign _2029_ = _2028_ & _2027_ /*14884*/;
  assign _2030_ = inv_13[3] & r_12[14] /*14883*/;
  assign _2031_ = _2029_ | _2030_ /*14882*/;
  assign _2032_ = inv_13[4] ^ r_12[15] /*14880*/;
  assign sum_13[4] = _2032_ ^ _2031_ /*14879*/;
  assign _2033_ = _2032_ & _2031_ /*14878*/;
  assign _2034_ = inv_13[4] & r_12[15] /*14877*/;
  assign _2035_ = _2033_ | _2034_ /*14876*/;
  assign _2036_ = inv_13[5] ^ r_12[16] /*14874*/;
  assign sum_13[5] = _2036_ ^ _2035_ /*14873*/;
  assign _2037_ = _2036_ & _2035_ /*14872*/;
  assign _2038_ = inv_13[5] & r_12[16] /*14871*/;
  assign _2039_ = _2037_ | _2038_ /*14870*/;
  assign _2040_ = inv_13[6] ^ r_12[17] /*14868*/;
  assign sum_13[6] = _2040_ ^ _2039_ /*14867*/;
  assign _2041_ = _2040_ & _2039_ /*14866*/;
  assign _2042_ = inv_13[6] & r_12[17] /*14865*/;
  assign _2043_ = _2041_ | _2042_ /*14864*/;
  assign _2044_ = inv_13[7] ^ r_12[18] /*14862*/;
  assign sum_13[7] = _2044_ ^ _2043_ /*14861*/;
  assign _2045_ = _2044_ & _2043_ /*14860*/;
  assign _2046_ = inv_13[7] & r_12[18] /*14859*/;
  assign _2047_ = _2045_ | _2046_ /*14858*/;
  assign _2048_ = inv_13[8] ^ r_12[19] /*14856*/;
  assign sum_13[8] = _2048_ ^ _2047_ /*14855*/;
  assign _2049_ = _2048_ & _2047_ /*14854*/;
  assign _2050_ = inv_13[8] & r_12[19] /*14853*/;
  assign _2051_ = _2049_ | _2050_ /*14852*/;
  assign _2052_ = inv_13[9] ^ r_12[20] /*14850*/;
  assign sum_13[9] = _2052_ ^ _2051_ /*14849*/;
  assign _2053_ = _2052_ & _2051_ /*14848*/;
  assign _2054_ = inv_13[9] & r_12[20] /*14847*/;
  assign _2055_ = _2053_ | _2054_ /*14846*/;
  assign _2056_ = inv_13[10] ^ r_12[21] /*14844*/;
  assign sum_13[10] = _2056_ ^ _2055_ /*14843*/;
  assign _2057_ = _2056_ & _2055_ /*14842*/;
  assign _2058_ = inv_13[10] & r_12[21] /*14841*/;
  assign _2059_ = _2057_ | _2058_ /*14840*/;
  assign _2060_ = inv_13[11] ^ r_12[22] /*14838*/;
  assign sum_13[11] = _2060_ ^ _2059_ /*14837*/;
  assign _2061_ = _2060_ & _2059_ /*14836*/;
  assign _2062_ = inv_13[11] & r_12[22] /*14835*/;
  assign _2063_ = _2061_ | _2062_ /*14834*/;
  assign _2064_ = inv_13[12] ^ r_12[23] /*14832*/;
  assign sum_13[12] = _2064_ ^ _2063_ /*14831*/;
  assign _2065_ = _2064_ & _2063_ /*14830*/;
  assign _2066_ = inv_13[12] & r_12[23] /*14829*/;
  assign _2067_ = _2065_ | _2066_ /*14828*/;
  assign _2068_ = inv_13[13] ^ r_12[24] /*14826*/;
  assign sum_13[13] = _2068_ ^ _2067_ /*14825*/;
  assign _2069_ = _2068_ & _2067_ /*14824*/;
  assign _2070_ = inv_13[13] & r_12[24] /*14823*/;
  assign _2071_ = _2069_ | _2070_ /*14822*/;
  assign _2072_ = inv_13[14] ^ r_12[25] /*14820*/;
  assign sum_13[14] = _2072_ ^ _2071_ /*14819*/;
  assign _2073_ = _2072_ & _2071_ /*14818*/;
  assign _2074_ = inv_13[14] & r_12[25] /*14817*/;
  assign _2075_ = _2073_ | _2074_ /*14816*/;
  assign _2076_ = inv_13[15] ^ r_12[26] /*14814*/;
  assign sum_13[15] = _2076_ ^ _2075_ /*14813*/;
  assign _2077_ = _2076_ & _2075_ /*14812*/;
  assign _2078_ = inv_13[15] & r_12[26] /*14811*/;
  assign _2079_ = _2077_ | _2078_ /*14810*/;
  assign _2080_ = inv_13[16] ^ r_12[27] /*14808*/;
  assign sum_13[16] = _2080_ ^ _2079_ /*14807*/;
  assign _2081_ = _2080_ & _2079_ /*14806*/;
  assign _2082_ = inv_13[16] & r_12[27] /*14805*/;
  assign _2083_ = _2081_ | _2082_ /*14804*/;
  assign _2084_ = inv_13[17] ^ r_12[28] /*14802*/;
  assign sum_13[17] = _2084_ ^ _2083_ /*14801*/;
  assign _2085_ = _2084_ & _2083_ /*14800*/;
  assign _2086_ = inv_13[17] & r_12[28] /*14799*/;
  assign _2087_ = _2085_ | _2086_ /*14798*/;
  assign _2088_ = inv_13[18] ^ r_12[29] /*14796*/;
  assign sum_13[18] = _2088_ ^ _2087_ /*14795*/;
  assign _2089_ = _2088_ & _2087_ /*14794*/;
  assign _2090_ = inv_13[18] & r_12[29] /*14793*/;
  assign _2091_ = _2089_ | _2090_ /*14792*/;
  assign _2092_ = inv_13[19] ^ r_12[30] /*14790*/;
  assign sum_13[19] = _2092_ ^ _2091_ /*14789*/;
  assign _2093_ = _2092_ & _2091_ /*14788*/;
  assign _2094_ = inv_13[19] & r_12[30] /*14787*/;
  assign _2095_ = _2093_ | _2094_ /*14786*/;
  assign _2096_ = inv_13[20] ^ r_12[31] /*14784*/;
  assign sum_13[20] = _2096_ ^ _2095_ /*14783*/;
  assign _2097_ = _2096_ & _2095_ /*14782*/;
  assign _2098_ = inv_13[20] & r_12[31] /*14781*/;
  assign _2099_ = _2097_ | _2098_ /*14780*/;
  assign _2100_ = inv_13[21] ^ r_12[32] /*14778*/;
  assign sum_13[21] = _2100_ ^ _2099_ /*14777*/;
  assign _2101_ = _2100_ & _2099_ /*14776*/;
  assign _2102_ = inv_13[21] & r_12[32] /*14775*/;
  assign _2103_ = _2101_ | _2102_ /*14774*/;
  assign _2104_ = inv_13[22] ^ r_12[33] /*14772*/;
  assign sum_13[22] = _2104_ ^ _2103_ /*14771*/;
  assign _2105_ = _2104_ & _2103_ /*14770*/;
  assign _2106_ = inv_13[22] & r_12[33] /*14769*/;
  assign _2107_ = _2105_ | _2106_ /*14768*/;
  assign _2108_ = inv_13[23] ^ r_12[34] /*14766*/;
  assign sum_13[23] = _2108_ ^ _2107_ /*14765*/;
  assign _2109_ = _2108_ & _2107_ /*14764*/;
  assign _2110_ = inv_13[23] & r_12[34] /*14763*/;
  assign _2111_ = _2109_ | _2110_ /*14762*/;
  assign q[11] = ~sum_13[23] /*14781*/;
  assign m_13[0] = r_12[11] /*14780*/;
  assign m_13[1] = r_12[12] /*14779*/;
  assign m_13[2] = r_12[13] /*14778*/;
  assign m_13[3] = r_12[14] /*14777*/;
  assign m_13[4] = r_12[15] /*14776*/;
  assign m_13[5] = r_12[16] /*14775*/;
  assign m_13[6] = r_12[17] /*14774*/;
  assign m_13[7] = r_12[18] /*14773*/;
  assign m_13[8] = r_12[19] /*14772*/;
  assign m_13[9] = r_12[20] /*14771*/;
  assign m_13[10] = r_12[21] /*14770*/;
  assign m_13[11] = r_12[22] /*14769*/;
  assign m_13[12] = r_12[23] /*14768*/;
  assign m_13[13] = r_12[24] /*14767*/;
  assign m_13[14] = r_12[25] /*14766*/;
  assign m_13[15] = r_12[26] /*14765*/;
  assign m_13[16] = r_12[27] /*14764*/;
  assign m_13[17] = r_12[28] /*14763*/;
  assign m_13[18] = r_12[29] /*14762*/;
  assign m_13[19] = r_12[30] /*14761*/;
  assign m_13[20] = r_12[31] /*14760*/;
  assign m_13[21] = r_12[32] /*14759*/;
  assign m_13[22] = r_12[33] /*14758*/;
  assign m_13[23] = r_12[34] /*14757*/;
  assign _2112_ = ~q[11] /*14755*/;
  assign _2113_ = sum_13[0] & q[11] /*14754*/;
  assign _2114_ = m_13[0] & _2112_ /*14753*/;
  assign r_13[11] = _2114_ | _2113_ /*14752*/;
  assign _2115_ = ~q[11] /*14751*/;
  assign _2116_ = sum_13[1] & q[11] /*14750*/;
  assign _2117_ = m_13[1] & _2115_ /*14749*/;
  assign r_13[12] = _2117_ | _2116_ /*14748*/;
  assign _2118_ = ~q[11] /*14747*/;
  assign _2119_ = sum_13[2] & q[11] /*14746*/;
  assign _2120_ = m_13[2] & _2118_ /*14745*/;
  assign r_13[13] = _2120_ | _2119_ /*14744*/;
  assign _2121_ = ~q[11] /*14743*/;
  assign _2122_ = sum_13[3] & q[11] /*14742*/;
  assign _2123_ = m_13[3] & _2121_ /*14741*/;
  assign r_13[14] = _2123_ | _2122_ /*14740*/;
  assign _2124_ = ~q[11] /*14739*/;
  assign _2125_ = sum_13[4] & q[11] /*14738*/;
  assign _2126_ = m_13[4] & _2124_ /*14737*/;
  assign r_13[15] = _2126_ | _2125_ /*14736*/;
  assign _2127_ = ~q[11] /*14735*/;
  assign _2128_ = sum_13[5] & q[11] /*14734*/;
  assign _2129_ = m_13[5] & _2127_ /*14733*/;
  assign r_13[16] = _2129_ | _2128_ /*14732*/;
  assign _2130_ = ~q[11] /*14731*/;
  assign _2131_ = sum_13[6] & q[11] /*14730*/;
  assign _2132_ = m_13[6] & _2130_ /*14729*/;
  assign r_13[17] = _2132_ | _2131_ /*14728*/;
  assign _2133_ = ~q[11] /*14727*/;
  assign _2134_ = sum_13[7] & q[11] /*14726*/;
  assign _2135_ = m_13[7] & _2133_ /*14725*/;
  assign r_13[18] = _2135_ | _2134_ /*14724*/;
  assign _2136_ = ~q[11] /*14723*/;
  assign _2137_ = sum_13[8] & q[11] /*14722*/;
  assign _2138_ = m_13[8] & _2136_ /*14721*/;
  assign r_13[19] = _2138_ | _2137_ /*14720*/;
  assign _2139_ = ~q[11] /*14719*/;
  assign _2140_ = sum_13[9] & q[11] /*14718*/;
  assign _2141_ = m_13[9] & _2139_ /*14717*/;
  assign r_13[20] = _2141_ | _2140_ /*14716*/;
  assign _2142_ = ~q[11] /*14715*/;
  assign _2143_ = sum_13[10] & q[11] /*14714*/;
  assign _2144_ = m_13[10] & _2142_ /*14713*/;
  assign r_13[21] = _2144_ | _2143_ /*14712*/;
  assign _2145_ = ~q[11] /*14711*/;
  assign _2146_ = sum_13[11] & q[11] /*14710*/;
  assign _2147_ = m_13[11] & _2145_ /*14709*/;
  assign r_13[22] = _2147_ | _2146_ /*14708*/;
  assign _2148_ = ~q[11] /*14707*/;
  assign _2149_ = sum_13[12] & q[11] /*14706*/;
  assign _2150_ = m_13[12] & _2148_ /*14705*/;
  assign r_13[23] = _2150_ | _2149_ /*14704*/;
  assign _2151_ = ~q[11] /*14703*/;
  assign _2152_ = sum_13[13] & q[11] /*14702*/;
  assign _2153_ = m_13[13] & _2151_ /*14701*/;
  assign r_13[24] = _2153_ | _2152_ /*14700*/;
  assign _2154_ = ~q[11] /*14699*/;
  assign _2155_ = sum_13[14] & q[11] /*14698*/;
  assign _2156_ = m_13[14] & _2154_ /*14697*/;
  assign r_13[25] = _2156_ | _2155_ /*14696*/;
  assign _2157_ = ~q[11] /*14695*/;
  assign _2158_ = sum_13[15] & q[11] /*14694*/;
  assign _2159_ = m_13[15] & _2157_ /*14693*/;
  assign r_13[26] = _2159_ | _2158_ /*14692*/;
  assign _2160_ = ~q[11] /*14691*/;
  assign _2161_ = sum_13[16] & q[11] /*14690*/;
  assign _2162_ = m_13[16] & _2160_ /*14689*/;
  assign r_13[27] = _2162_ | _2161_ /*14688*/;
  assign _2163_ = ~q[11] /*14687*/;
  assign _2164_ = sum_13[17] & q[11] /*14686*/;
  assign _2165_ = m_13[17] & _2163_ /*14685*/;
  assign r_13[28] = _2165_ | _2164_ /*14684*/;
  assign _2166_ = ~q[11] /*14683*/;
  assign _2167_ = sum_13[18] & q[11] /*14682*/;
  assign _2168_ = m_13[18] & _2166_ /*14681*/;
  assign r_13[29] = _2168_ | _2167_ /*14680*/;
  assign _2169_ = ~q[11] /*14679*/;
  assign _2170_ = sum_13[19] & q[11] /*14678*/;
  assign _2171_ = m_13[19] & _2169_ /*14677*/;
  assign r_13[30] = _2171_ | _2170_ /*14676*/;
  assign _2172_ = ~q[11] /*14675*/;
  assign _2173_ = sum_13[20] & q[11] /*14674*/;
  assign _2174_ = m_13[20] & _2172_ /*14673*/;
  assign r_13[31] = _2174_ | _2173_ /*14672*/;
  assign _2175_ = ~q[11] /*14671*/;
  assign _2176_ = sum_13[21] & q[11] /*14670*/;
  assign _2177_ = m_13[21] & _2175_ /*14669*/;
  assign r_13[32] = _2177_ | _2176_ /*14668*/;
  assign _2178_ = ~q[11] /*14667*/;
  assign _2179_ = sum_13[22] & q[11] /*14666*/;
  assign _2180_ = m_13[22] & _2178_ /*14665*/;
  assign r_13[33] = _2180_ | _2179_ /*14664*/;
  assign _2181_ = ~q[11] /*14663*/;
  assign _2182_ = sum_13[23] & q[11] /*14662*/;
  assign _2183_ = m_13[23] & _2181_ /*14661*/;
  assign r_13[34] = _2183_ | _2182_ /*14660*/;
assign r_13[0]= r_12[0] /*14659*/;
assign r_13[1]= r_12[1] /*14658*/;
assign r_13[2]= r_12[2] /*14657*/;
assign r_13[3]= r_12[3] /*14656*/;
assign r_13[4]= r_12[4] /*14655*/;
assign r_13[5]= r_12[5] /*14654*/;
assign r_13[6]= r_12[6] /*14653*/;
assign r_13[7]= r_12[7] /*14652*/;
assign r_13[8]= r_12[8] /*14651*/;
assign r_13[9]= r_12[9] /*14650*/;
assign r_13[10]= r_12[10] /*14649*/;
  assign inv_14[0] = ~div[0] /*14592*/;
  assign inv_14[1] = ~div[1] /*14591*/;
  assign inv_14[2] = ~div[2] /*14590*/;
  assign inv_14[3] = ~div[3] /*14589*/;
  assign inv_14[4] = ~div[4] /*14588*/;
  assign inv_14[5] = ~div[5] /*14587*/;
  assign inv_14[6] = ~div[6] /*14586*/;
  assign inv_14[7] = ~div[7] /*14585*/;
  assign inv_14[8] = ~div[8] /*14584*/;
  assign inv_14[9] = ~div[9] /*14583*/;
  assign inv_14[10] = ~div[10] /*14582*/;
  assign inv_14[11] = ~div[11] /*14581*/;
  assign inv_14[12] = ~div[12] /*14580*/;
  assign inv_14[13] = ~div[13] /*14579*/;
  assign inv_14[14] = ~div[14] /*14578*/;
  assign inv_14[15] = ~div[15] /*14577*/;
  assign inv_14[16] = ~div[16] /*14576*/;
  assign inv_14[17] = ~div[17] /*14575*/;
  assign inv_14[18] = ~div[18] /*14574*/;
  assign inv_14[19] = ~div[19] /*14573*/;
  assign inv_14[20] = ~div[20] /*14572*/;
  assign inv_14[21] = ~div[21] /*14571*/;
  assign inv_14[22] = ~div[22] /*14570*/;
assign inv_14[23] = oneWire /*14569*/;
  assign _2184_ = inv_14[0] ^ r_13[10] /*14567*/;
  assign sum_14[0] = _2184_ ^ oneWire /*14566*/;
  assign _2185_ = _2184_ & oneWire /*14565*/;
  assign _2186_ = inv_14[0] & r_13[10] /*14564*/;
  assign _2187_ = _2185_ | _2186_ /*14563*/;
  assign _2188_ = inv_14[1] ^ r_13[11] /*14562*/;
  assign sum_14[1] = _2188_ ^ _2187_ /*14561*/;
  assign _2189_ = _2188_ & _2187_ /*14560*/;
  assign _2190_ = inv_14[1] & r_13[11] /*14559*/;
  assign _2191_ = _2189_ | _2190_ /*14558*/;
  assign _2192_ = inv_14[2] ^ r_13[12] /*14556*/;
  assign sum_14[2] = _2192_ ^ _2191_ /*14555*/;
  assign _2193_ = _2192_ & _2191_ /*14554*/;
  assign _2194_ = inv_14[2] & r_13[12] /*14553*/;
  assign _2195_ = _2193_ | _2194_ /*14552*/;
  assign _2196_ = inv_14[3] ^ r_13[13] /*14550*/;
  assign sum_14[3] = _2196_ ^ _2195_ /*14549*/;
  assign _2197_ = _2196_ & _2195_ /*14548*/;
  assign _2198_ = inv_14[3] & r_13[13] /*14547*/;
  assign _2199_ = _2197_ | _2198_ /*14546*/;
  assign _2200_ = inv_14[4] ^ r_13[14] /*14544*/;
  assign sum_14[4] = _2200_ ^ _2199_ /*14543*/;
  assign _2201_ = _2200_ & _2199_ /*14542*/;
  assign _2202_ = inv_14[4] & r_13[14] /*14541*/;
  assign _2203_ = _2201_ | _2202_ /*14540*/;
  assign _2204_ = inv_14[5] ^ r_13[15] /*14538*/;
  assign sum_14[5] = _2204_ ^ _2203_ /*14537*/;
  assign _2205_ = _2204_ & _2203_ /*14536*/;
  assign _2206_ = inv_14[5] & r_13[15] /*14535*/;
  assign _2207_ = _2205_ | _2206_ /*14534*/;
  assign _2208_ = inv_14[6] ^ r_13[16] /*14532*/;
  assign sum_14[6] = _2208_ ^ _2207_ /*14531*/;
  assign _2209_ = _2208_ & _2207_ /*14530*/;
  assign _2210_ = inv_14[6] & r_13[16] /*14529*/;
  assign _2211_ = _2209_ | _2210_ /*14528*/;
  assign _2212_ = inv_14[7] ^ r_13[17] /*14526*/;
  assign sum_14[7] = _2212_ ^ _2211_ /*14525*/;
  assign _2213_ = _2212_ & _2211_ /*14524*/;
  assign _2214_ = inv_14[7] & r_13[17] /*14523*/;
  assign _2215_ = _2213_ | _2214_ /*14522*/;
  assign _2216_ = inv_14[8] ^ r_13[18] /*14520*/;
  assign sum_14[8] = _2216_ ^ _2215_ /*14519*/;
  assign _2217_ = _2216_ & _2215_ /*14518*/;
  assign _2218_ = inv_14[8] & r_13[18] /*14517*/;
  assign _2219_ = _2217_ | _2218_ /*14516*/;
  assign _2220_ = inv_14[9] ^ r_13[19] /*14514*/;
  assign sum_14[9] = _2220_ ^ _2219_ /*14513*/;
  assign _2221_ = _2220_ & _2219_ /*14512*/;
  assign _2222_ = inv_14[9] & r_13[19] /*14511*/;
  assign _2223_ = _2221_ | _2222_ /*14510*/;
  assign _2224_ = inv_14[10] ^ r_13[20] /*14508*/;
  assign sum_14[10] = _2224_ ^ _2223_ /*14507*/;
  assign _2225_ = _2224_ & _2223_ /*14506*/;
  assign _2226_ = inv_14[10] & r_13[20] /*14505*/;
  assign _2227_ = _2225_ | _2226_ /*14504*/;
  assign _2228_ = inv_14[11] ^ r_13[21] /*14502*/;
  assign sum_14[11] = _2228_ ^ _2227_ /*14501*/;
  assign _2229_ = _2228_ & _2227_ /*14500*/;
  assign _2230_ = inv_14[11] & r_13[21] /*14499*/;
  assign _2231_ = _2229_ | _2230_ /*14498*/;
  assign _2232_ = inv_14[12] ^ r_13[22] /*14496*/;
  assign sum_14[12] = _2232_ ^ _2231_ /*14495*/;
  assign _2233_ = _2232_ & _2231_ /*14494*/;
  assign _2234_ = inv_14[12] & r_13[22] /*14493*/;
  assign _2235_ = _2233_ | _2234_ /*14492*/;
  assign _2236_ = inv_14[13] ^ r_13[23] /*14490*/;
  assign sum_14[13] = _2236_ ^ _2235_ /*14489*/;
  assign _2237_ = _2236_ & _2235_ /*14488*/;
  assign _2238_ = inv_14[13] & r_13[23] /*14487*/;
  assign _2239_ = _2237_ | _2238_ /*14486*/;
  assign _2240_ = inv_14[14] ^ r_13[24] /*14484*/;
  assign sum_14[14] = _2240_ ^ _2239_ /*14483*/;
  assign _2241_ = _2240_ & _2239_ /*14482*/;
  assign _2242_ = inv_14[14] & r_13[24] /*14481*/;
  assign _2243_ = _2241_ | _2242_ /*14480*/;
  assign _2244_ = inv_14[15] ^ r_13[25] /*14478*/;
  assign sum_14[15] = _2244_ ^ _2243_ /*14477*/;
  assign _2245_ = _2244_ & _2243_ /*14476*/;
  assign _2246_ = inv_14[15] & r_13[25] /*14475*/;
  assign _2247_ = _2245_ | _2246_ /*14474*/;
  assign _2248_ = inv_14[16] ^ r_13[26] /*14472*/;
  assign sum_14[16] = _2248_ ^ _2247_ /*14471*/;
  assign _2249_ = _2248_ & _2247_ /*14470*/;
  assign _2250_ = inv_14[16] & r_13[26] /*14469*/;
  assign _2251_ = _2249_ | _2250_ /*14468*/;
  assign _2252_ = inv_14[17] ^ r_13[27] /*14466*/;
  assign sum_14[17] = _2252_ ^ _2251_ /*14465*/;
  assign _2253_ = _2252_ & _2251_ /*14464*/;
  assign _2254_ = inv_14[17] & r_13[27] /*14463*/;
  assign _2255_ = _2253_ | _2254_ /*14462*/;
  assign _2256_ = inv_14[18] ^ r_13[28] /*14460*/;
  assign sum_14[18] = _2256_ ^ _2255_ /*14459*/;
  assign _2257_ = _2256_ & _2255_ /*14458*/;
  assign _2258_ = inv_14[18] & r_13[28] /*14457*/;
  assign _2259_ = _2257_ | _2258_ /*14456*/;
  assign _2260_ = inv_14[19] ^ r_13[29] /*14454*/;
  assign sum_14[19] = _2260_ ^ _2259_ /*14453*/;
  assign _2261_ = _2260_ & _2259_ /*14452*/;
  assign _2262_ = inv_14[19] & r_13[29] /*14451*/;
  assign _2263_ = _2261_ | _2262_ /*14450*/;
  assign _2264_ = inv_14[20] ^ r_13[30] /*14448*/;
  assign sum_14[20] = _2264_ ^ _2263_ /*14447*/;
  assign _2265_ = _2264_ & _2263_ /*14446*/;
  assign _2266_ = inv_14[20] & r_13[30] /*14445*/;
  assign _2267_ = _2265_ | _2266_ /*14444*/;
  assign _2268_ = inv_14[21] ^ r_13[31] /*14442*/;
  assign sum_14[21] = _2268_ ^ _2267_ /*14441*/;
  assign _2269_ = _2268_ & _2267_ /*14440*/;
  assign _2270_ = inv_14[21] & r_13[31] /*14439*/;
  assign _2271_ = _2269_ | _2270_ /*14438*/;
  assign _2272_ = inv_14[22] ^ r_13[32] /*14436*/;
  assign sum_14[22] = _2272_ ^ _2271_ /*14435*/;
  assign _2273_ = _2272_ & _2271_ /*14434*/;
  assign _2274_ = inv_14[22] & r_13[32] /*14433*/;
  assign _2275_ = _2273_ | _2274_ /*14432*/;
  assign _2276_ = inv_14[23] ^ r_13[33] /*14430*/;
  assign sum_14[23] = _2276_ ^ _2275_ /*14429*/;
  assign _2277_ = _2276_ & _2275_ /*14428*/;
  assign _2278_ = inv_14[23] & r_13[33] /*14427*/;
  assign _2279_ = _2277_ | _2278_ /*14426*/;
  assign q[10] = ~sum_14[23] /*14445*/;
  assign m_14[0] = r_13[10] /*14444*/;
  assign m_14[1] = r_13[11] /*14443*/;
  assign m_14[2] = r_13[12] /*14442*/;
  assign m_14[3] = r_13[13] /*14441*/;
  assign m_14[4] = r_13[14] /*14440*/;
  assign m_14[5] = r_13[15] /*14439*/;
  assign m_14[6] = r_13[16] /*14438*/;
  assign m_14[7] = r_13[17] /*14437*/;
  assign m_14[8] = r_13[18] /*14436*/;
  assign m_14[9] = r_13[19] /*14435*/;
  assign m_14[10] = r_13[20] /*14434*/;
  assign m_14[11] = r_13[21] /*14433*/;
  assign m_14[12] = r_13[22] /*14432*/;
  assign m_14[13] = r_13[23] /*14431*/;
  assign m_14[14] = r_13[24] /*14430*/;
  assign m_14[15] = r_13[25] /*14429*/;
  assign m_14[16] = r_13[26] /*14428*/;
  assign m_14[17] = r_13[27] /*14427*/;
  assign m_14[18] = r_13[28] /*14426*/;
  assign m_14[19] = r_13[29] /*14425*/;
  assign m_14[20] = r_13[30] /*14424*/;
  assign m_14[21] = r_13[31] /*14423*/;
  assign m_14[22] = r_13[32] /*14422*/;
  assign m_14[23] = r_13[33] /*14421*/;
  assign _2280_ = ~q[10] /*14419*/;
  assign _2281_ = sum_14[0] & q[10] /*14418*/;
  assign _2282_ = m_14[0] & _2280_ /*14417*/;
  assign r_14[10] = _2282_ | _2281_ /*14416*/;
  assign _2283_ = ~q[10] /*14415*/;
  assign _2284_ = sum_14[1] & q[10] /*14414*/;
  assign _2285_ = m_14[1] & _2283_ /*14413*/;
  assign r_14[11] = _2285_ | _2284_ /*14412*/;
  assign _2286_ = ~q[10] /*14411*/;
  assign _2287_ = sum_14[2] & q[10] /*14410*/;
  assign _2288_ = m_14[2] & _2286_ /*14409*/;
  assign r_14[12] = _2288_ | _2287_ /*14408*/;
  assign _2289_ = ~q[10] /*14407*/;
  assign _2290_ = sum_14[3] & q[10] /*14406*/;
  assign _2291_ = m_14[3] & _2289_ /*14405*/;
  assign r_14[13] = _2291_ | _2290_ /*14404*/;
  assign _2292_ = ~q[10] /*14403*/;
  assign _2293_ = sum_14[4] & q[10] /*14402*/;
  assign _2294_ = m_14[4] & _2292_ /*14401*/;
  assign r_14[14] = _2294_ | _2293_ /*14400*/;
  assign _2295_ = ~q[10] /*14399*/;
  assign _2296_ = sum_14[5] & q[10] /*14398*/;
  assign _2297_ = m_14[5] & _2295_ /*14397*/;
  assign r_14[15] = _2297_ | _2296_ /*14396*/;
  assign _2298_ = ~q[10] /*14395*/;
  assign _2299_ = sum_14[6] & q[10] /*14394*/;
  assign _2300_ = m_14[6] & _2298_ /*14393*/;
  assign r_14[16] = _2300_ | _2299_ /*14392*/;
  assign _2301_ = ~q[10] /*14391*/;
  assign _2302_ = sum_14[7] & q[10] /*14390*/;
  assign _2303_ = m_14[7] & _2301_ /*14389*/;
  assign r_14[17] = _2303_ | _2302_ /*14388*/;
  assign _2304_ = ~q[10] /*14387*/;
  assign _2305_ = sum_14[8] & q[10] /*14386*/;
  assign _2306_ = m_14[8] & _2304_ /*14385*/;
  assign r_14[18] = _2306_ | _2305_ /*14384*/;
  assign _2307_ = ~q[10] /*14383*/;
  assign _2308_ = sum_14[9] & q[10] /*14382*/;
  assign _2309_ = m_14[9] & _2307_ /*14381*/;
  assign r_14[19] = _2309_ | _2308_ /*14380*/;
  assign _2310_ = ~q[10] /*14379*/;
  assign _2311_ = sum_14[10] & q[10] /*14378*/;
  assign _2312_ = m_14[10] & _2310_ /*14377*/;
  assign r_14[20] = _2312_ | _2311_ /*14376*/;
  assign _2313_ = ~q[10] /*14375*/;
  assign _2314_ = sum_14[11] & q[10] /*14374*/;
  assign _2315_ = m_14[11] & _2313_ /*14373*/;
  assign r_14[21] = _2315_ | _2314_ /*14372*/;
  assign _2316_ = ~q[10] /*14371*/;
  assign _2317_ = sum_14[12] & q[10] /*14370*/;
  assign _2318_ = m_14[12] & _2316_ /*14369*/;
  assign r_14[22] = _2318_ | _2317_ /*14368*/;
  assign _2319_ = ~q[10] /*14367*/;
  assign _2320_ = sum_14[13] & q[10] /*14366*/;
  assign _2321_ = m_14[13] & _2319_ /*14365*/;
  assign r_14[23] = _2321_ | _2320_ /*14364*/;
  assign _2322_ = ~q[10] /*14363*/;
  assign _2323_ = sum_14[14] & q[10] /*14362*/;
  assign _2324_ = m_14[14] & _2322_ /*14361*/;
  assign r_14[24] = _2324_ | _2323_ /*14360*/;
  assign _2325_ = ~q[10] /*14359*/;
  assign _2326_ = sum_14[15] & q[10] /*14358*/;
  assign _2327_ = m_14[15] & _2325_ /*14357*/;
  assign r_14[25] = _2327_ | _2326_ /*14356*/;
  assign _2328_ = ~q[10] /*14355*/;
  assign _2329_ = sum_14[16] & q[10] /*14354*/;
  assign _2330_ = m_14[16] & _2328_ /*14353*/;
  assign r_14[26] = _2330_ | _2329_ /*14352*/;
  assign _2331_ = ~q[10] /*14351*/;
  assign _2332_ = sum_14[17] & q[10] /*14350*/;
  assign _2333_ = m_14[17] & _2331_ /*14349*/;
  assign r_14[27] = _2333_ | _2332_ /*14348*/;
  assign _2334_ = ~q[10] /*14347*/;
  assign _2335_ = sum_14[18] & q[10] /*14346*/;
  assign _2336_ = m_14[18] & _2334_ /*14345*/;
  assign r_14[28] = _2336_ | _2335_ /*14344*/;
  assign _2337_ = ~q[10] /*14343*/;
  assign _2338_ = sum_14[19] & q[10] /*14342*/;
  assign _2339_ = m_14[19] & _2337_ /*14341*/;
  assign r_14[29] = _2339_ | _2338_ /*14340*/;
  assign _2340_ = ~q[10] /*14339*/;
  assign _2341_ = sum_14[20] & q[10] /*14338*/;
  assign _2342_ = m_14[20] & _2340_ /*14337*/;
  assign r_14[30] = _2342_ | _2341_ /*14336*/;
  assign _2343_ = ~q[10] /*14335*/;
  assign _2344_ = sum_14[21] & q[10] /*14334*/;
  assign _2345_ = m_14[21] & _2343_ /*14333*/;
  assign r_14[31] = _2345_ | _2344_ /*14332*/;
  assign _2346_ = ~q[10] /*14331*/;
  assign _2347_ = sum_14[22] & q[10] /*14330*/;
  assign _2348_ = m_14[22] & _2346_ /*14329*/;
  assign r_14[32] = _2348_ | _2347_ /*14328*/;
  assign _2349_ = ~q[10] /*14327*/;
  assign _2350_ = sum_14[23] & q[10] /*14326*/;
  assign _2351_ = m_14[23] & _2349_ /*14325*/;
  assign r_14[33] = _2351_ | _2350_ /*14324*/;
assign r_14[0]= r_13[0] /*14323*/;
assign r_14[1]= r_13[1] /*14322*/;
assign r_14[2]= r_13[2] /*14321*/;
assign r_14[3]= r_13[3] /*14320*/;
assign r_14[4]= r_13[4] /*14319*/;
assign r_14[5]= r_13[5] /*14318*/;
assign r_14[6]= r_13[6] /*14317*/;
assign r_14[7]= r_13[7] /*14316*/;
assign r_14[8]= r_13[8] /*14315*/;
assign r_14[9]= r_13[9] /*14314*/;
  assign inv_15[0] = ~div[0] /*14256*/;
  assign inv_15[1] = ~div[1] /*14255*/;
  assign inv_15[2] = ~div[2] /*14254*/;
  assign inv_15[3] = ~div[3] /*14253*/;
  assign inv_15[4] = ~div[4] /*14252*/;
  assign inv_15[5] = ~div[5] /*14251*/;
  assign inv_15[6] = ~div[6] /*14250*/;
  assign inv_15[7] = ~div[7] /*14249*/;
  assign inv_15[8] = ~div[8] /*14248*/;
  assign inv_15[9] = ~div[9] /*14247*/;
  assign inv_15[10] = ~div[10] /*14246*/;
  assign inv_15[11] = ~div[11] /*14245*/;
  assign inv_15[12] = ~div[12] /*14244*/;
  assign inv_15[13] = ~div[13] /*14243*/;
  assign inv_15[14] = ~div[14] /*14242*/;
  assign inv_15[15] = ~div[15] /*14241*/;
  assign inv_15[16] = ~div[16] /*14240*/;
  assign inv_15[17] = ~div[17] /*14239*/;
  assign inv_15[18] = ~div[18] /*14238*/;
  assign inv_15[19] = ~div[19] /*14237*/;
  assign inv_15[20] = ~div[20] /*14236*/;
  assign inv_15[21] = ~div[21] /*14235*/;
  assign inv_15[22] = ~div[22] /*14234*/;
assign inv_15[23] = oneWire /*14233*/;
  assign _2352_ = inv_15[0] ^ r_14[9] /*14231*/;
  assign sum_15[0] = _2352_ ^ oneWire /*14230*/;
  assign _2353_ = _2352_ & oneWire /*14229*/;
  assign _2354_ = inv_15[0] & r_14[9] /*14228*/;
  assign _2355_ = _2353_ | _2354_ /*14227*/;
  assign _2356_ = inv_15[1] ^ r_14[10] /*14226*/;
  assign sum_15[1] = _2356_ ^ _2355_ /*14225*/;
  assign _2357_ = _2356_ & _2355_ /*14224*/;
  assign _2358_ = inv_15[1] & r_14[10] /*14223*/;
  assign _2359_ = _2357_ | _2358_ /*14222*/;
  assign _2360_ = inv_15[2] ^ r_14[11] /*14220*/;
  assign sum_15[2] = _2360_ ^ _2359_ /*14219*/;
  assign _2361_ = _2360_ & _2359_ /*14218*/;
  assign _2362_ = inv_15[2] & r_14[11] /*14217*/;
  assign _2363_ = _2361_ | _2362_ /*14216*/;
  assign _2364_ = inv_15[3] ^ r_14[12] /*14214*/;
  assign sum_15[3] = _2364_ ^ _2363_ /*14213*/;
  assign _2365_ = _2364_ & _2363_ /*14212*/;
  assign _2366_ = inv_15[3] & r_14[12] /*14211*/;
  assign _2367_ = _2365_ | _2366_ /*14210*/;
  assign _2368_ = inv_15[4] ^ r_14[13] /*14208*/;
  assign sum_15[4] = _2368_ ^ _2367_ /*14207*/;
  assign _2369_ = _2368_ & _2367_ /*14206*/;
  assign _2370_ = inv_15[4] & r_14[13] /*14205*/;
  assign _2371_ = _2369_ | _2370_ /*14204*/;
  assign _2372_ = inv_15[5] ^ r_14[14] /*14202*/;
  assign sum_15[5] = _2372_ ^ _2371_ /*14201*/;
  assign _2373_ = _2372_ & _2371_ /*14200*/;
  assign _2374_ = inv_15[5] & r_14[14] /*14199*/;
  assign _2375_ = _2373_ | _2374_ /*14198*/;
  assign _2376_ = inv_15[6] ^ r_14[15] /*14196*/;
  assign sum_15[6] = _2376_ ^ _2375_ /*14195*/;
  assign _2377_ = _2376_ & _2375_ /*14194*/;
  assign _2378_ = inv_15[6] & r_14[15] /*14193*/;
  assign _2379_ = _2377_ | _2378_ /*14192*/;
  assign _2380_ = inv_15[7] ^ r_14[16] /*14190*/;
  assign sum_15[7] = _2380_ ^ _2379_ /*14189*/;
  assign _2381_ = _2380_ & _2379_ /*14188*/;
  assign _2382_ = inv_15[7] & r_14[16] /*14187*/;
  assign _2383_ = _2381_ | _2382_ /*14186*/;
  assign _2384_ = inv_15[8] ^ r_14[17] /*14184*/;
  assign sum_15[8] = _2384_ ^ _2383_ /*14183*/;
  assign _2385_ = _2384_ & _2383_ /*14182*/;
  assign _2386_ = inv_15[8] & r_14[17] /*14181*/;
  assign _2387_ = _2385_ | _2386_ /*14180*/;
  assign _2388_ = inv_15[9] ^ r_14[18] /*14178*/;
  assign sum_15[9] = _2388_ ^ _2387_ /*14177*/;
  assign _2389_ = _2388_ & _2387_ /*14176*/;
  assign _2390_ = inv_15[9] & r_14[18] /*14175*/;
  assign _2391_ = _2389_ | _2390_ /*14174*/;
  assign _2392_ = inv_15[10] ^ r_14[19] /*14172*/;
  assign sum_15[10] = _2392_ ^ _2391_ /*14171*/;
  assign _2393_ = _2392_ & _2391_ /*14170*/;
  assign _2394_ = inv_15[10] & r_14[19] /*14169*/;
  assign _2395_ = _2393_ | _2394_ /*14168*/;
  assign _2396_ = inv_15[11] ^ r_14[20] /*14166*/;
  assign sum_15[11] = _2396_ ^ _2395_ /*14165*/;
  assign _2397_ = _2396_ & _2395_ /*14164*/;
  assign _2398_ = inv_15[11] & r_14[20] /*14163*/;
  assign _2399_ = _2397_ | _2398_ /*14162*/;
  assign _2400_ = inv_15[12] ^ r_14[21] /*14160*/;
  assign sum_15[12] = _2400_ ^ _2399_ /*14159*/;
  assign _2401_ = _2400_ & _2399_ /*14158*/;
  assign _2402_ = inv_15[12] & r_14[21] /*14157*/;
  assign _2403_ = _2401_ | _2402_ /*14156*/;
  assign _2404_ = inv_15[13] ^ r_14[22] /*14154*/;
  assign sum_15[13] = _2404_ ^ _2403_ /*14153*/;
  assign _2405_ = _2404_ & _2403_ /*14152*/;
  assign _2406_ = inv_15[13] & r_14[22] /*14151*/;
  assign _2407_ = _2405_ | _2406_ /*14150*/;
  assign _2408_ = inv_15[14] ^ r_14[23] /*14148*/;
  assign sum_15[14] = _2408_ ^ _2407_ /*14147*/;
  assign _2409_ = _2408_ & _2407_ /*14146*/;
  assign _2410_ = inv_15[14] & r_14[23] /*14145*/;
  assign _2411_ = _2409_ | _2410_ /*14144*/;
  assign _2412_ = inv_15[15] ^ r_14[24] /*14142*/;
  assign sum_15[15] = _2412_ ^ _2411_ /*14141*/;
  assign _2413_ = _2412_ & _2411_ /*14140*/;
  assign _2414_ = inv_15[15] & r_14[24] /*14139*/;
  assign _2415_ = _2413_ | _2414_ /*14138*/;
  assign _2416_ = inv_15[16] ^ r_14[25] /*14136*/;
  assign sum_15[16] = _2416_ ^ _2415_ /*14135*/;
  assign _2417_ = _2416_ & _2415_ /*14134*/;
  assign _2418_ = inv_15[16] & r_14[25] /*14133*/;
  assign _2419_ = _2417_ | _2418_ /*14132*/;
  assign _2420_ = inv_15[17] ^ r_14[26] /*14130*/;
  assign sum_15[17] = _2420_ ^ _2419_ /*14129*/;
  assign _2421_ = _2420_ & _2419_ /*14128*/;
  assign _2422_ = inv_15[17] & r_14[26] /*14127*/;
  assign _2423_ = _2421_ | _2422_ /*14126*/;
  assign _2424_ = inv_15[18] ^ r_14[27] /*14124*/;
  assign sum_15[18] = _2424_ ^ _2423_ /*14123*/;
  assign _2425_ = _2424_ & _2423_ /*14122*/;
  assign _2426_ = inv_15[18] & r_14[27] /*14121*/;
  assign _2427_ = _2425_ | _2426_ /*14120*/;
  assign _2428_ = inv_15[19] ^ r_14[28] /*14118*/;
  assign sum_15[19] = _2428_ ^ _2427_ /*14117*/;
  assign _2429_ = _2428_ & _2427_ /*14116*/;
  assign _2430_ = inv_15[19] & r_14[28] /*14115*/;
  assign _2431_ = _2429_ | _2430_ /*14114*/;
  assign _2432_ = inv_15[20] ^ r_14[29] /*14112*/;
  assign sum_15[20] = _2432_ ^ _2431_ /*14111*/;
  assign _2433_ = _2432_ & _2431_ /*14110*/;
  assign _2434_ = inv_15[20] & r_14[29] /*14109*/;
  assign _2435_ = _2433_ | _2434_ /*14108*/;
  assign _2436_ = inv_15[21] ^ r_14[30] /*14106*/;
  assign sum_15[21] = _2436_ ^ _2435_ /*14105*/;
  assign _2437_ = _2436_ & _2435_ /*14104*/;
  assign _2438_ = inv_15[21] & r_14[30] /*14103*/;
  assign _2439_ = _2437_ | _2438_ /*14102*/;
  assign _2440_ = inv_15[22] ^ r_14[31] /*14100*/;
  assign sum_15[22] = _2440_ ^ _2439_ /*14099*/;
  assign _2441_ = _2440_ & _2439_ /*14098*/;
  assign _2442_ = inv_15[22] & r_14[31] /*14097*/;
  assign _2443_ = _2441_ | _2442_ /*14096*/;
  assign _2444_ = inv_15[23] ^ r_14[32] /*14094*/;
  assign sum_15[23] = _2444_ ^ _2443_ /*14093*/;
  assign _2445_ = _2444_ & _2443_ /*14092*/;
  assign _2446_ = inv_15[23] & r_14[32] /*14091*/;
  assign _2447_ = _2445_ | _2446_ /*14090*/;
  assign q[9] = ~sum_15[23] /*14109*/;
  assign m_15[0] = r_14[9] /*14108*/;
  assign m_15[1] = r_14[10] /*14107*/;
  assign m_15[2] = r_14[11] /*14106*/;
  assign m_15[3] = r_14[12] /*14105*/;
  assign m_15[4] = r_14[13] /*14104*/;
  assign m_15[5] = r_14[14] /*14103*/;
  assign m_15[6] = r_14[15] /*14102*/;
  assign m_15[7] = r_14[16] /*14101*/;
  assign m_15[8] = r_14[17] /*14100*/;
  assign m_15[9] = r_14[18] /*14099*/;
  assign m_15[10] = r_14[19] /*14098*/;
  assign m_15[11] = r_14[20] /*14097*/;
  assign m_15[12] = r_14[21] /*14096*/;
  assign m_15[13] = r_14[22] /*14095*/;
  assign m_15[14] = r_14[23] /*14094*/;
  assign m_15[15] = r_14[24] /*14093*/;
  assign m_15[16] = r_14[25] /*14092*/;
  assign m_15[17] = r_14[26] /*14091*/;
  assign m_15[18] = r_14[27] /*14090*/;
  assign m_15[19] = r_14[28] /*14089*/;
  assign m_15[20] = r_14[29] /*14088*/;
  assign m_15[21] = r_14[30] /*14087*/;
  assign m_15[22] = r_14[31] /*14086*/;
  assign m_15[23] = r_14[32] /*14085*/;
  assign _2448_ = ~q[9] /*14083*/;
  assign _2449_ = sum_15[0] & q[9] /*14082*/;
  assign _2450_ = m_15[0] & _2448_ /*14081*/;
  assign r_15[9] = _2450_ | _2449_ /*14080*/;
  assign _2451_ = ~q[9] /*14079*/;
  assign _2452_ = sum_15[1] & q[9] /*14078*/;
  assign _2453_ = m_15[1] & _2451_ /*14077*/;
  assign r_15[10] = _2453_ | _2452_ /*14076*/;
  assign _2454_ = ~q[9] /*14075*/;
  assign _2455_ = sum_15[2] & q[9] /*14074*/;
  assign _2456_ = m_15[2] & _2454_ /*14073*/;
  assign r_15[11] = _2456_ | _2455_ /*14072*/;
  assign _2457_ = ~q[9] /*14071*/;
  assign _2458_ = sum_15[3] & q[9] /*14070*/;
  assign _2459_ = m_15[3] & _2457_ /*14069*/;
  assign r_15[12] = _2459_ | _2458_ /*14068*/;
  assign _2460_ = ~q[9] /*14067*/;
  assign _2461_ = sum_15[4] & q[9] /*14066*/;
  assign _2462_ = m_15[4] & _2460_ /*14065*/;
  assign r_15[13] = _2462_ | _2461_ /*14064*/;
  assign _2463_ = ~q[9] /*14063*/;
  assign _2464_ = sum_15[5] & q[9] /*14062*/;
  assign _2465_ = m_15[5] & _2463_ /*14061*/;
  assign r_15[14] = _2465_ | _2464_ /*14060*/;
  assign _2466_ = ~q[9] /*14059*/;
  assign _2467_ = sum_15[6] & q[9] /*14058*/;
  assign _2468_ = m_15[6] & _2466_ /*14057*/;
  assign r_15[15] = _2468_ | _2467_ /*14056*/;
  assign _2469_ = ~q[9] /*14055*/;
  assign _2470_ = sum_15[7] & q[9] /*14054*/;
  assign _2471_ = m_15[7] & _2469_ /*14053*/;
  assign r_15[16] = _2471_ | _2470_ /*14052*/;
  assign _2472_ = ~q[9] /*14051*/;
  assign _2473_ = sum_15[8] & q[9] /*14050*/;
  assign _2474_ = m_15[8] & _2472_ /*14049*/;
  assign r_15[17] = _2474_ | _2473_ /*14048*/;
  assign _2475_ = ~q[9] /*14047*/;
  assign _2476_ = sum_15[9] & q[9] /*14046*/;
  assign _2477_ = m_15[9] & _2475_ /*14045*/;
  assign r_15[18] = _2477_ | _2476_ /*14044*/;
  assign _2478_ = ~q[9] /*14043*/;
  assign _2479_ = sum_15[10] & q[9] /*14042*/;
  assign _2480_ = m_15[10] & _2478_ /*14041*/;
  assign r_15[19] = _2480_ | _2479_ /*14040*/;
  assign _2481_ = ~q[9] /*14039*/;
  assign _2482_ = sum_15[11] & q[9] /*14038*/;
  assign _2483_ = m_15[11] & _2481_ /*14037*/;
  assign r_15[20] = _2483_ | _2482_ /*14036*/;
  assign _2484_ = ~q[9] /*14035*/;
  assign _2485_ = sum_15[12] & q[9] /*14034*/;
  assign _2486_ = m_15[12] & _2484_ /*14033*/;
  assign r_15[21] = _2486_ | _2485_ /*14032*/;
  assign _2487_ = ~q[9] /*14031*/;
  assign _2488_ = sum_15[13] & q[9] /*14030*/;
  assign _2489_ = m_15[13] & _2487_ /*14029*/;
  assign r_15[22] = _2489_ | _2488_ /*14028*/;
  assign _2490_ = ~q[9] /*14027*/;
  assign _2491_ = sum_15[14] & q[9] /*14026*/;
  assign _2492_ = m_15[14] & _2490_ /*14025*/;
  assign r_15[23] = _2492_ | _2491_ /*14024*/;
  assign _2493_ = ~q[9] /*14023*/;
  assign _2494_ = sum_15[15] & q[9] /*14022*/;
  assign _2495_ = m_15[15] & _2493_ /*14021*/;
  assign r_15[24] = _2495_ | _2494_ /*14020*/;
  assign _2496_ = ~q[9] /*14019*/;
  assign _2497_ = sum_15[16] & q[9] /*14018*/;
  assign _2498_ = m_15[16] & _2496_ /*14017*/;
  assign r_15[25] = _2498_ | _2497_ /*14016*/;
  assign _2499_ = ~q[9] /*14015*/;
  assign _2500_ = sum_15[17] & q[9] /*14014*/;
  assign _2501_ = m_15[17] & _2499_ /*14013*/;
  assign r_15[26] = _2501_ | _2500_ /*14012*/;
  assign _2502_ = ~q[9] /*14011*/;
  assign _2503_ = sum_15[18] & q[9] /*14010*/;
  assign _2504_ = m_15[18] & _2502_ /*14009*/;
  assign r_15[27] = _2504_ | _2503_ /*14008*/;
  assign _2505_ = ~q[9] /*14007*/;
  assign _2506_ = sum_15[19] & q[9] /*14006*/;
  assign _2507_ = m_15[19] & _2505_ /*14005*/;
  assign r_15[28] = _2507_ | _2506_ /*14004*/;
  assign _2508_ = ~q[9] /*14003*/;
  assign _2509_ = sum_15[20] & q[9] /*14002*/;
  assign _2510_ = m_15[20] & _2508_ /*14001*/;
  assign r_15[29] = _2510_ | _2509_ /*14000*/;
  assign _2511_ = ~q[9] /*13999*/;
  assign _2512_ = sum_15[21] & q[9] /*13998*/;
  assign _2513_ = m_15[21] & _2511_ /*13997*/;
  assign r_15[30] = _2513_ | _2512_ /*13996*/;
  assign _2514_ = ~q[9] /*13995*/;
  assign _2515_ = sum_15[22] & q[9] /*13994*/;
  assign _2516_ = m_15[22] & _2514_ /*13993*/;
  assign r_15[31] = _2516_ | _2515_ /*13992*/;
  assign _2517_ = ~q[9] /*13991*/;
  assign _2518_ = sum_15[23] & q[9] /*13990*/;
  assign _2519_ = m_15[23] & _2517_ /*13989*/;
  assign r_15[32] = _2519_ | _2518_ /*13988*/;
assign r_15[0]= r_14[0] /*13987*/;
assign r_15[1]= r_14[1] /*13986*/;
assign r_15[2]= r_14[2] /*13985*/;
assign r_15[3]= r_14[3] /*13984*/;
assign r_15[4]= r_14[4] /*13983*/;
assign r_15[5]= r_14[5] /*13982*/;
assign r_15[6]= r_14[6] /*13981*/;
assign r_15[7]= r_14[7] /*13980*/;
assign r_15[8]= r_14[8] /*13979*/;
  assign inv_16[0] = ~div[0] /*13920*/;
  assign inv_16[1] = ~div[1] /*13919*/;
  assign inv_16[2] = ~div[2] /*13918*/;
  assign inv_16[3] = ~div[3] /*13917*/;
  assign inv_16[4] = ~div[4] /*13916*/;
  assign inv_16[5] = ~div[5] /*13915*/;
  assign inv_16[6] = ~div[6] /*13914*/;
  assign inv_16[7] = ~div[7] /*13913*/;
  assign inv_16[8] = ~div[8] /*13912*/;
  assign inv_16[9] = ~div[9] /*13911*/;
  assign inv_16[10] = ~div[10] /*13910*/;
  assign inv_16[11] = ~div[11] /*13909*/;
  assign inv_16[12] = ~div[12] /*13908*/;
  assign inv_16[13] = ~div[13] /*13907*/;
  assign inv_16[14] = ~div[14] /*13906*/;
  assign inv_16[15] = ~div[15] /*13905*/;
  assign inv_16[16] = ~div[16] /*13904*/;
  assign inv_16[17] = ~div[17] /*13903*/;
  assign inv_16[18] = ~div[18] /*13902*/;
  assign inv_16[19] = ~div[19] /*13901*/;
  assign inv_16[20] = ~div[20] /*13900*/;
  assign inv_16[21] = ~div[21] /*13899*/;
  assign inv_16[22] = ~div[22] /*13898*/;
assign inv_16[23] = oneWire /*13897*/;
  assign _2520_ = inv_16[0] ^ r_15[8] /*13895*/;
  assign sum_16[0] = _2520_ ^ oneWire /*13894*/;
  assign _2521_ = _2520_ & oneWire /*13893*/;
  assign _2522_ = inv_16[0] & r_15[8] /*13892*/;
  assign _2523_ = _2521_ | _2522_ /*13891*/;
  assign _2524_ = inv_16[1] ^ r_15[9] /*13890*/;
  assign sum_16[1] = _2524_ ^ _2523_ /*13889*/;
  assign _2525_ = _2524_ & _2523_ /*13888*/;
  assign _2526_ = inv_16[1] & r_15[9] /*13887*/;
  assign _2527_ = _2525_ | _2526_ /*13886*/;
  assign _2528_ = inv_16[2] ^ r_15[10] /*13884*/;
  assign sum_16[2] = _2528_ ^ _2527_ /*13883*/;
  assign _2529_ = _2528_ & _2527_ /*13882*/;
  assign _2530_ = inv_16[2] & r_15[10] /*13881*/;
  assign _2531_ = _2529_ | _2530_ /*13880*/;
  assign _2532_ = inv_16[3] ^ r_15[11] /*13878*/;
  assign sum_16[3] = _2532_ ^ _2531_ /*13877*/;
  assign _2533_ = _2532_ & _2531_ /*13876*/;
  assign _2534_ = inv_16[3] & r_15[11] /*13875*/;
  assign _2535_ = _2533_ | _2534_ /*13874*/;
  assign _2536_ = inv_16[4] ^ r_15[12] /*13872*/;
  assign sum_16[4] = _2536_ ^ _2535_ /*13871*/;
  assign _2537_ = _2536_ & _2535_ /*13870*/;
  assign _2538_ = inv_16[4] & r_15[12] /*13869*/;
  assign _2539_ = _2537_ | _2538_ /*13868*/;
  assign _2540_ = inv_16[5] ^ r_15[13] /*13866*/;
  assign sum_16[5] = _2540_ ^ _2539_ /*13865*/;
  assign _2541_ = _2540_ & _2539_ /*13864*/;
  assign _2542_ = inv_16[5] & r_15[13] /*13863*/;
  assign _2543_ = _2541_ | _2542_ /*13862*/;
  assign _2544_ = inv_16[6] ^ r_15[14] /*13860*/;
  assign sum_16[6] = _2544_ ^ _2543_ /*13859*/;
  assign _2545_ = _2544_ & _2543_ /*13858*/;
  assign _2546_ = inv_16[6] & r_15[14] /*13857*/;
  assign _2547_ = _2545_ | _2546_ /*13856*/;
  assign _2548_ = inv_16[7] ^ r_15[15] /*13854*/;
  assign sum_16[7] = _2548_ ^ _2547_ /*13853*/;
  assign _2549_ = _2548_ & _2547_ /*13852*/;
  assign _2550_ = inv_16[7] & r_15[15] /*13851*/;
  assign _2551_ = _2549_ | _2550_ /*13850*/;
  assign _2552_ = inv_16[8] ^ r_15[16] /*13848*/;
  assign sum_16[8] = _2552_ ^ _2551_ /*13847*/;
  assign _2553_ = _2552_ & _2551_ /*13846*/;
  assign _2554_ = inv_16[8] & r_15[16] /*13845*/;
  assign _2555_ = _2553_ | _2554_ /*13844*/;
  assign _2556_ = inv_16[9] ^ r_15[17] /*13842*/;
  assign sum_16[9] = _2556_ ^ _2555_ /*13841*/;
  assign _2557_ = _2556_ & _2555_ /*13840*/;
  assign _2558_ = inv_16[9] & r_15[17] /*13839*/;
  assign _2559_ = _2557_ | _2558_ /*13838*/;
  assign _2560_ = inv_16[10] ^ r_15[18] /*13836*/;
  assign sum_16[10] = _2560_ ^ _2559_ /*13835*/;
  assign _2561_ = _2560_ & _2559_ /*13834*/;
  assign _2562_ = inv_16[10] & r_15[18] /*13833*/;
  assign _2563_ = _2561_ | _2562_ /*13832*/;
  assign _2564_ = inv_16[11] ^ r_15[19] /*13830*/;
  assign sum_16[11] = _2564_ ^ _2563_ /*13829*/;
  assign _2565_ = _2564_ & _2563_ /*13828*/;
  assign _2566_ = inv_16[11] & r_15[19] /*13827*/;
  assign _2567_ = _2565_ | _2566_ /*13826*/;
  assign _2568_ = inv_16[12] ^ r_15[20] /*13824*/;
  assign sum_16[12] = _2568_ ^ _2567_ /*13823*/;
  assign _2569_ = _2568_ & _2567_ /*13822*/;
  assign _2570_ = inv_16[12] & r_15[20] /*13821*/;
  assign _2571_ = _2569_ | _2570_ /*13820*/;
  assign _2572_ = inv_16[13] ^ r_15[21] /*13818*/;
  assign sum_16[13] = _2572_ ^ _2571_ /*13817*/;
  assign _2573_ = _2572_ & _2571_ /*13816*/;
  assign _2574_ = inv_16[13] & r_15[21] /*13815*/;
  assign _2575_ = _2573_ | _2574_ /*13814*/;
  assign _2576_ = inv_16[14] ^ r_15[22] /*13812*/;
  assign sum_16[14] = _2576_ ^ _2575_ /*13811*/;
  assign _2577_ = _2576_ & _2575_ /*13810*/;
  assign _2578_ = inv_16[14] & r_15[22] /*13809*/;
  assign _2579_ = _2577_ | _2578_ /*13808*/;
  assign _2580_ = inv_16[15] ^ r_15[23] /*13806*/;
  assign sum_16[15] = _2580_ ^ _2579_ /*13805*/;
  assign _2581_ = _2580_ & _2579_ /*13804*/;
  assign _2582_ = inv_16[15] & r_15[23] /*13803*/;
  assign _2583_ = _2581_ | _2582_ /*13802*/;
  assign _2584_ = inv_16[16] ^ r_15[24] /*13800*/;
  assign sum_16[16] = _2584_ ^ _2583_ /*13799*/;
  assign _2585_ = _2584_ & _2583_ /*13798*/;
  assign _2586_ = inv_16[16] & r_15[24] /*13797*/;
  assign _2587_ = _2585_ | _2586_ /*13796*/;
  assign _2588_ = inv_16[17] ^ r_15[25] /*13794*/;
  assign sum_16[17] = _2588_ ^ _2587_ /*13793*/;
  assign _2589_ = _2588_ & _2587_ /*13792*/;
  assign _2590_ = inv_16[17] & r_15[25] /*13791*/;
  assign _2591_ = _2589_ | _2590_ /*13790*/;
  assign _2592_ = inv_16[18] ^ r_15[26] /*13788*/;
  assign sum_16[18] = _2592_ ^ _2591_ /*13787*/;
  assign _2593_ = _2592_ & _2591_ /*13786*/;
  assign _2594_ = inv_16[18] & r_15[26] /*13785*/;
  assign _2595_ = _2593_ | _2594_ /*13784*/;
  assign _2596_ = inv_16[19] ^ r_15[27] /*13782*/;
  assign sum_16[19] = _2596_ ^ _2595_ /*13781*/;
  assign _2597_ = _2596_ & _2595_ /*13780*/;
  assign _2598_ = inv_16[19] & r_15[27] /*13779*/;
  assign _2599_ = _2597_ | _2598_ /*13778*/;
  assign _2600_ = inv_16[20] ^ r_15[28] /*13776*/;
  assign sum_16[20] = _2600_ ^ _2599_ /*13775*/;
  assign _2601_ = _2600_ & _2599_ /*13774*/;
  assign _2602_ = inv_16[20] & r_15[28] /*13773*/;
  assign _2603_ = _2601_ | _2602_ /*13772*/;
  assign _2604_ = inv_16[21] ^ r_15[29] /*13770*/;
  assign sum_16[21] = _2604_ ^ _2603_ /*13769*/;
  assign _2605_ = _2604_ & _2603_ /*13768*/;
  assign _2606_ = inv_16[21] & r_15[29] /*13767*/;
  assign _2607_ = _2605_ | _2606_ /*13766*/;
  assign _2608_ = inv_16[22] ^ r_15[30] /*13764*/;
  assign sum_16[22] = _2608_ ^ _2607_ /*13763*/;
  assign _2609_ = _2608_ & _2607_ /*13762*/;
  assign _2610_ = inv_16[22] & r_15[30] /*13761*/;
  assign _2611_ = _2609_ | _2610_ /*13760*/;
  assign _2612_ = inv_16[23] ^ r_15[31] /*13758*/;
  assign sum_16[23] = _2612_ ^ _2611_ /*13757*/;
  assign _2613_ = _2612_ & _2611_ /*13756*/;
  assign _2614_ = inv_16[23] & r_15[31] /*13755*/;
  assign _2615_ = _2613_ | _2614_ /*13754*/;
  assign q[8] = ~sum_16[23] /*13773*/;
  assign m_16[0] = r_15[8] /*13772*/;
  assign m_16[1] = r_15[9] /*13771*/;
  assign m_16[2] = r_15[10] /*13770*/;
  assign m_16[3] = r_15[11] /*13769*/;
  assign m_16[4] = r_15[12] /*13768*/;
  assign m_16[5] = r_15[13] /*13767*/;
  assign m_16[6] = r_15[14] /*13766*/;
  assign m_16[7] = r_15[15] /*13765*/;
  assign m_16[8] = r_15[16] /*13764*/;
  assign m_16[9] = r_15[17] /*13763*/;
  assign m_16[10] = r_15[18] /*13762*/;
  assign m_16[11] = r_15[19] /*13761*/;
  assign m_16[12] = r_15[20] /*13760*/;
  assign m_16[13] = r_15[21] /*13759*/;
  assign m_16[14] = r_15[22] /*13758*/;
  assign m_16[15] = r_15[23] /*13757*/;
  assign m_16[16] = r_15[24] /*13756*/;
  assign m_16[17] = r_15[25] /*13755*/;
  assign m_16[18] = r_15[26] /*13754*/;
  assign m_16[19] = r_15[27] /*13753*/;
  assign m_16[20] = r_15[28] /*13752*/;
  assign m_16[21] = r_15[29] /*13751*/;
  assign m_16[22] = r_15[30] /*13750*/;
  assign m_16[23] = r_15[31] /*13749*/;
  assign _2616_ = ~q[8] /*13747*/;
  assign _2617_ = sum_16[0] & q[8] /*13746*/;
  assign _2618_ = m_16[0] & _2616_ /*13745*/;
  assign r_16[8] = _2618_ | _2617_ /*13744*/;
  assign _2619_ = ~q[8] /*13743*/;
  assign _2620_ = sum_16[1] & q[8] /*13742*/;
  assign _2621_ = m_16[1] & _2619_ /*13741*/;
  assign r_16[9] = _2621_ | _2620_ /*13740*/;
  assign _2622_ = ~q[8] /*13739*/;
  assign _2623_ = sum_16[2] & q[8] /*13738*/;
  assign _2624_ = m_16[2] & _2622_ /*13737*/;
  assign r_16[10] = _2624_ | _2623_ /*13736*/;
  assign _2625_ = ~q[8] /*13735*/;
  assign _2626_ = sum_16[3] & q[8] /*13734*/;
  assign _2627_ = m_16[3] & _2625_ /*13733*/;
  assign r_16[11] = _2627_ | _2626_ /*13732*/;
  assign _2628_ = ~q[8] /*13731*/;
  assign _2629_ = sum_16[4] & q[8] /*13730*/;
  assign _2630_ = m_16[4] & _2628_ /*13729*/;
  assign r_16[12] = _2630_ | _2629_ /*13728*/;
  assign _2631_ = ~q[8] /*13727*/;
  assign _2632_ = sum_16[5] & q[8] /*13726*/;
  assign _2633_ = m_16[5] & _2631_ /*13725*/;
  assign r_16[13] = _2633_ | _2632_ /*13724*/;
  assign _2634_ = ~q[8] /*13723*/;
  assign _2635_ = sum_16[6] & q[8] /*13722*/;
  assign _2636_ = m_16[6] & _2634_ /*13721*/;
  assign r_16[14] = _2636_ | _2635_ /*13720*/;
  assign _2637_ = ~q[8] /*13719*/;
  assign _2638_ = sum_16[7] & q[8] /*13718*/;
  assign _2639_ = m_16[7] & _2637_ /*13717*/;
  assign r_16[15] = _2639_ | _2638_ /*13716*/;
  assign _2640_ = ~q[8] /*13715*/;
  assign _2641_ = sum_16[8] & q[8] /*13714*/;
  assign _2642_ = m_16[8] & _2640_ /*13713*/;
  assign r_16[16] = _2642_ | _2641_ /*13712*/;
  assign _2643_ = ~q[8] /*13711*/;
  assign _2644_ = sum_16[9] & q[8] /*13710*/;
  assign _2645_ = m_16[9] & _2643_ /*13709*/;
  assign r_16[17] = _2645_ | _2644_ /*13708*/;
  assign _2646_ = ~q[8] /*13707*/;
  assign _2647_ = sum_16[10] & q[8] /*13706*/;
  assign _2648_ = m_16[10] & _2646_ /*13705*/;
  assign r_16[18] = _2648_ | _2647_ /*13704*/;
  assign _2649_ = ~q[8] /*13703*/;
  assign _2650_ = sum_16[11] & q[8] /*13702*/;
  assign _2651_ = m_16[11] & _2649_ /*13701*/;
  assign r_16[19] = _2651_ | _2650_ /*13700*/;
  assign _2652_ = ~q[8] /*13699*/;
  assign _2653_ = sum_16[12] & q[8] /*13698*/;
  assign _2654_ = m_16[12] & _2652_ /*13697*/;
  assign r_16[20] = _2654_ | _2653_ /*13696*/;
  assign _2655_ = ~q[8] /*13695*/;
  assign _2656_ = sum_16[13] & q[8] /*13694*/;
  assign _2657_ = m_16[13] & _2655_ /*13693*/;
  assign r_16[21] = _2657_ | _2656_ /*13692*/;
  assign _2658_ = ~q[8] /*13691*/;
  assign _2659_ = sum_16[14] & q[8] /*13690*/;
  assign _2660_ = m_16[14] & _2658_ /*13689*/;
  assign r_16[22] = _2660_ | _2659_ /*13688*/;
  assign _2661_ = ~q[8] /*13687*/;
  assign _2662_ = sum_16[15] & q[8] /*13686*/;
  assign _2663_ = m_16[15] & _2661_ /*13685*/;
  assign r_16[23] = _2663_ | _2662_ /*13684*/;
  assign _2664_ = ~q[8] /*13683*/;
  assign _2665_ = sum_16[16] & q[8] /*13682*/;
  assign _2666_ = m_16[16] & _2664_ /*13681*/;
  assign r_16[24] = _2666_ | _2665_ /*13680*/;
  assign _2667_ = ~q[8] /*13679*/;
  assign _2668_ = sum_16[17] & q[8] /*13678*/;
  assign _2669_ = m_16[17] & _2667_ /*13677*/;
  assign r_16[25] = _2669_ | _2668_ /*13676*/;
  assign _2670_ = ~q[8] /*13675*/;
  assign _2671_ = sum_16[18] & q[8] /*13674*/;
  assign _2672_ = m_16[18] & _2670_ /*13673*/;
  assign r_16[26] = _2672_ | _2671_ /*13672*/;
  assign _2673_ = ~q[8] /*13671*/;
  assign _2674_ = sum_16[19] & q[8] /*13670*/;
  assign _2675_ = m_16[19] & _2673_ /*13669*/;
  assign r_16[27] = _2675_ | _2674_ /*13668*/;
  assign _2676_ = ~q[8] /*13667*/;
  assign _2677_ = sum_16[20] & q[8] /*13666*/;
  assign _2678_ = m_16[20] & _2676_ /*13665*/;
  assign r_16[28] = _2678_ | _2677_ /*13664*/;
  assign _2679_ = ~q[8] /*13663*/;
  assign _2680_ = sum_16[21] & q[8] /*13662*/;
  assign _2681_ = m_16[21] & _2679_ /*13661*/;
  assign r_16[29] = _2681_ | _2680_ /*13660*/;
  assign _2682_ = ~q[8] /*13659*/;
  assign _2683_ = sum_16[22] & q[8] /*13658*/;
  assign _2684_ = m_16[22] & _2682_ /*13657*/;
  assign r_16[30] = _2684_ | _2683_ /*13656*/;
  assign _2685_ = ~q[8] /*13655*/;
  assign _2686_ = sum_16[23] & q[8] /*13654*/;
  assign _2687_ = m_16[23] & _2685_ /*13653*/;
  assign r_16[31] = _2687_ | _2686_ /*13652*/;
assign r_16[0]= r_15[0] /*13651*/;
assign r_16[1]= r_15[1] /*13650*/;
assign r_16[2]= r_15[2] /*13649*/;
assign r_16[3]= r_15[3] /*13648*/;
assign r_16[4]= r_15[4] /*13647*/;
assign r_16[5]= r_15[5] /*13646*/;
assign r_16[6]= r_15[6] /*13645*/;
assign r_16[7]= r_15[7] /*13644*/;
  assign inv_17[0] = ~div[0] /*13584*/;
  assign inv_17[1] = ~div[1] /*13583*/;
  assign inv_17[2] = ~div[2] /*13582*/;
  assign inv_17[3] = ~div[3] /*13581*/;
  assign inv_17[4] = ~div[4] /*13580*/;
  assign inv_17[5] = ~div[5] /*13579*/;
  assign inv_17[6] = ~div[6] /*13578*/;
  assign inv_17[7] = ~div[7] /*13577*/;
  assign inv_17[8] = ~div[8] /*13576*/;
  assign inv_17[9] = ~div[9] /*13575*/;
  assign inv_17[10] = ~div[10] /*13574*/;
  assign inv_17[11] = ~div[11] /*13573*/;
  assign inv_17[12] = ~div[12] /*13572*/;
  assign inv_17[13] = ~div[13] /*13571*/;
  assign inv_17[14] = ~div[14] /*13570*/;
  assign inv_17[15] = ~div[15] /*13569*/;
  assign inv_17[16] = ~div[16] /*13568*/;
  assign inv_17[17] = ~div[17] /*13567*/;
  assign inv_17[18] = ~div[18] /*13566*/;
  assign inv_17[19] = ~div[19] /*13565*/;
  assign inv_17[20] = ~div[20] /*13564*/;
  assign inv_17[21] = ~div[21] /*13563*/;
  assign inv_17[22] = ~div[22] /*13562*/;
assign inv_17[23] = oneWire /*13561*/;
  assign _2688_ = inv_17[0] ^ r_16[7] /*13559*/;
  assign sum_17[0] = _2688_ ^ oneWire /*13558*/;
  assign _2689_ = _2688_ & oneWire /*13557*/;
  assign _2690_ = inv_17[0] & r_16[7] /*13556*/;
  assign _2691_ = _2689_ | _2690_ /*13555*/;
  assign _2692_ = inv_17[1] ^ r_16[8] /*13554*/;
  assign sum_17[1] = _2692_ ^ _2691_ /*13553*/;
  assign _2693_ = _2692_ & _2691_ /*13552*/;
  assign _2694_ = inv_17[1] & r_16[8] /*13551*/;
  assign _2695_ = _2693_ | _2694_ /*13550*/;
  assign _2696_ = inv_17[2] ^ r_16[9] /*13548*/;
  assign sum_17[2] = _2696_ ^ _2695_ /*13547*/;
  assign _2697_ = _2696_ & _2695_ /*13546*/;
  assign _2698_ = inv_17[2] & r_16[9] /*13545*/;
  assign _2699_ = _2697_ | _2698_ /*13544*/;
  assign _2700_ = inv_17[3] ^ r_16[10] /*13542*/;
  assign sum_17[3] = _2700_ ^ _2699_ /*13541*/;
  assign _2701_ = _2700_ & _2699_ /*13540*/;
  assign _2702_ = inv_17[3] & r_16[10] /*13539*/;
  assign _2703_ = _2701_ | _2702_ /*13538*/;
  assign _2704_ = inv_17[4] ^ r_16[11] /*13536*/;
  assign sum_17[4] = _2704_ ^ _2703_ /*13535*/;
  assign _2705_ = _2704_ & _2703_ /*13534*/;
  assign _2706_ = inv_17[4] & r_16[11] /*13533*/;
  assign _2707_ = _2705_ | _2706_ /*13532*/;
  assign _2708_ = inv_17[5] ^ r_16[12] /*13530*/;
  assign sum_17[5] = _2708_ ^ _2707_ /*13529*/;
  assign _2709_ = _2708_ & _2707_ /*13528*/;
  assign _2710_ = inv_17[5] & r_16[12] /*13527*/;
  assign _2711_ = _2709_ | _2710_ /*13526*/;
  assign _2712_ = inv_17[6] ^ r_16[13] /*13524*/;
  assign sum_17[6] = _2712_ ^ _2711_ /*13523*/;
  assign _2713_ = _2712_ & _2711_ /*13522*/;
  assign _2714_ = inv_17[6] & r_16[13] /*13521*/;
  assign _2715_ = _2713_ | _2714_ /*13520*/;
  assign _2716_ = inv_17[7] ^ r_16[14] /*13518*/;
  assign sum_17[7] = _2716_ ^ _2715_ /*13517*/;
  assign _2717_ = _2716_ & _2715_ /*13516*/;
  assign _2718_ = inv_17[7] & r_16[14] /*13515*/;
  assign _2719_ = _2717_ | _2718_ /*13514*/;
  assign _2720_ = inv_17[8] ^ r_16[15] /*13512*/;
  assign sum_17[8] = _2720_ ^ _2719_ /*13511*/;
  assign _2721_ = _2720_ & _2719_ /*13510*/;
  assign _2722_ = inv_17[8] & r_16[15] /*13509*/;
  assign _2723_ = _2721_ | _2722_ /*13508*/;
  assign _2724_ = inv_17[9] ^ r_16[16] /*13506*/;
  assign sum_17[9] = _2724_ ^ _2723_ /*13505*/;
  assign _2725_ = _2724_ & _2723_ /*13504*/;
  assign _2726_ = inv_17[9] & r_16[16] /*13503*/;
  assign _2727_ = _2725_ | _2726_ /*13502*/;
  assign _2728_ = inv_17[10] ^ r_16[17] /*13500*/;
  assign sum_17[10] = _2728_ ^ _2727_ /*13499*/;
  assign _2729_ = _2728_ & _2727_ /*13498*/;
  assign _2730_ = inv_17[10] & r_16[17] /*13497*/;
  assign _2731_ = _2729_ | _2730_ /*13496*/;
  assign _2732_ = inv_17[11] ^ r_16[18] /*13494*/;
  assign sum_17[11] = _2732_ ^ _2731_ /*13493*/;
  assign _2733_ = _2732_ & _2731_ /*13492*/;
  assign _2734_ = inv_17[11] & r_16[18] /*13491*/;
  assign _2735_ = _2733_ | _2734_ /*13490*/;
  assign _2736_ = inv_17[12] ^ r_16[19] /*13488*/;
  assign sum_17[12] = _2736_ ^ _2735_ /*13487*/;
  assign _2737_ = _2736_ & _2735_ /*13486*/;
  assign _2738_ = inv_17[12] & r_16[19] /*13485*/;
  assign _2739_ = _2737_ | _2738_ /*13484*/;
  assign _2740_ = inv_17[13] ^ r_16[20] /*13482*/;
  assign sum_17[13] = _2740_ ^ _2739_ /*13481*/;
  assign _2741_ = _2740_ & _2739_ /*13480*/;
  assign _2742_ = inv_17[13] & r_16[20] /*13479*/;
  assign _2743_ = _2741_ | _2742_ /*13478*/;
  assign _2744_ = inv_17[14] ^ r_16[21] /*13476*/;
  assign sum_17[14] = _2744_ ^ _2743_ /*13475*/;
  assign _2745_ = _2744_ & _2743_ /*13474*/;
  assign _2746_ = inv_17[14] & r_16[21] /*13473*/;
  assign _2747_ = _2745_ | _2746_ /*13472*/;
  assign _2748_ = inv_17[15] ^ r_16[22] /*13470*/;
  assign sum_17[15] = _2748_ ^ _2747_ /*13469*/;
  assign _2749_ = _2748_ & _2747_ /*13468*/;
  assign _2750_ = inv_17[15] & r_16[22] /*13467*/;
  assign _2751_ = _2749_ | _2750_ /*13466*/;
  assign _2752_ = inv_17[16] ^ r_16[23] /*13464*/;
  assign sum_17[16] = _2752_ ^ _2751_ /*13463*/;
  assign _2753_ = _2752_ & _2751_ /*13462*/;
  assign _2754_ = inv_17[16] & r_16[23] /*13461*/;
  assign _2755_ = _2753_ | _2754_ /*13460*/;
  assign _2756_ = inv_17[17] ^ r_16[24] /*13458*/;
  assign sum_17[17] = _2756_ ^ _2755_ /*13457*/;
  assign _2757_ = _2756_ & _2755_ /*13456*/;
  assign _2758_ = inv_17[17] & r_16[24] /*13455*/;
  assign _2759_ = _2757_ | _2758_ /*13454*/;
  assign _2760_ = inv_17[18] ^ r_16[25] /*13452*/;
  assign sum_17[18] = _2760_ ^ _2759_ /*13451*/;
  assign _2761_ = _2760_ & _2759_ /*13450*/;
  assign _2762_ = inv_17[18] & r_16[25] /*13449*/;
  assign _2763_ = _2761_ | _2762_ /*13448*/;
  assign _2764_ = inv_17[19] ^ r_16[26] /*13446*/;
  assign sum_17[19] = _2764_ ^ _2763_ /*13445*/;
  assign _2765_ = _2764_ & _2763_ /*13444*/;
  assign _2766_ = inv_17[19] & r_16[26] /*13443*/;
  assign _2767_ = _2765_ | _2766_ /*13442*/;
  assign _2768_ = inv_17[20] ^ r_16[27] /*13440*/;
  assign sum_17[20] = _2768_ ^ _2767_ /*13439*/;
  assign _2769_ = _2768_ & _2767_ /*13438*/;
  assign _2770_ = inv_17[20] & r_16[27] /*13437*/;
  assign _2771_ = _2769_ | _2770_ /*13436*/;
  assign _2772_ = inv_17[21] ^ r_16[28] /*13434*/;
  assign sum_17[21] = _2772_ ^ _2771_ /*13433*/;
  assign _2773_ = _2772_ & _2771_ /*13432*/;
  assign _2774_ = inv_17[21] & r_16[28] /*13431*/;
  assign _2775_ = _2773_ | _2774_ /*13430*/;
  assign _2776_ = inv_17[22] ^ r_16[29] /*13428*/;
  assign sum_17[22] = _2776_ ^ _2775_ /*13427*/;
  assign _2777_ = _2776_ & _2775_ /*13426*/;
  assign _2778_ = inv_17[22] & r_16[29] /*13425*/;
  assign _2779_ = _2777_ | _2778_ /*13424*/;
  assign _2780_ = inv_17[23] ^ r_16[30] /*13422*/;
  assign sum_17[23] = _2780_ ^ _2779_ /*13421*/;
  assign _2781_ = _2780_ & _2779_ /*13420*/;
  assign _2782_ = inv_17[23] & r_16[30] /*13419*/;
  assign _2783_ = _2781_ | _2782_ /*13418*/;
  assign q[7] = ~sum_17[23] /*13437*/;
  assign m_17[0] = r_16[7] /*13436*/;
  assign m_17[1] = r_16[8] /*13435*/;
  assign m_17[2] = r_16[9] /*13434*/;
  assign m_17[3] = r_16[10] /*13433*/;
  assign m_17[4] = r_16[11] /*13432*/;
  assign m_17[5] = r_16[12] /*13431*/;
  assign m_17[6] = r_16[13] /*13430*/;
  assign m_17[7] = r_16[14] /*13429*/;
  assign m_17[8] = r_16[15] /*13428*/;
  assign m_17[9] = r_16[16] /*13427*/;
  assign m_17[10] = r_16[17] /*13426*/;
  assign m_17[11] = r_16[18] /*13425*/;
  assign m_17[12] = r_16[19] /*13424*/;
  assign m_17[13] = r_16[20] /*13423*/;
  assign m_17[14] = r_16[21] /*13422*/;
  assign m_17[15] = r_16[22] /*13421*/;
  assign m_17[16] = r_16[23] /*13420*/;
  assign m_17[17] = r_16[24] /*13419*/;
  assign m_17[18] = r_16[25] /*13418*/;
  assign m_17[19] = r_16[26] /*13417*/;
  assign m_17[20] = r_16[27] /*13416*/;
  assign m_17[21] = r_16[28] /*13415*/;
  assign m_17[22] = r_16[29] /*13414*/;
  assign m_17[23] = r_16[30] /*13413*/;
  assign _2784_ = ~q[7] /*13411*/;
  assign _2785_ = sum_17[0] & q[7] /*13410*/;
  assign _2786_ = m_17[0] & _2784_ /*13409*/;
  assign r_17[7] = _2786_ | _2785_ /*13408*/;
  assign _2787_ = ~q[7] /*13407*/;
  assign _2788_ = sum_17[1] & q[7] /*13406*/;
  assign _2789_ = m_17[1] & _2787_ /*13405*/;
  assign r_17[8] = _2789_ | _2788_ /*13404*/;
  assign _2790_ = ~q[7] /*13403*/;
  assign _2791_ = sum_17[2] & q[7] /*13402*/;
  assign _2792_ = m_17[2] & _2790_ /*13401*/;
  assign r_17[9] = _2792_ | _2791_ /*13400*/;
  assign _2793_ = ~q[7] /*13399*/;
  assign _2794_ = sum_17[3] & q[7] /*13398*/;
  assign _2795_ = m_17[3] & _2793_ /*13397*/;
  assign r_17[10] = _2795_ | _2794_ /*13396*/;
  assign _2796_ = ~q[7] /*13395*/;
  assign _2797_ = sum_17[4] & q[7] /*13394*/;
  assign _2798_ = m_17[4] & _2796_ /*13393*/;
  assign r_17[11] = _2798_ | _2797_ /*13392*/;
  assign _2799_ = ~q[7] /*13391*/;
  assign _2800_ = sum_17[5] & q[7] /*13390*/;
  assign _2801_ = m_17[5] & _2799_ /*13389*/;
  assign r_17[12] = _2801_ | _2800_ /*13388*/;
  assign _2802_ = ~q[7] /*13387*/;
  assign _2803_ = sum_17[6] & q[7] /*13386*/;
  assign _2804_ = m_17[6] & _2802_ /*13385*/;
  assign r_17[13] = _2804_ | _2803_ /*13384*/;
  assign _2805_ = ~q[7] /*13383*/;
  assign _2806_ = sum_17[7] & q[7] /*13382*/;
  assign _2807_ = m_17[7] & _2805_ /*13381*/;
  assign r_17[14] = _2807_ | _2806_ /*13380*/;
  assign _2808_ = ~q[7] /*13379*/;
  assign _2809_ = sum_17[8] & q[7] /*13378*/;
  assign _2810_ = m_17[8] & _2808_ /*13377*/;
  assign r_17[15] = _2810_ | _2809_ /*13376*/;
  assign _2811_ = ~q[7] /*13375*/;
  assign _2812_ = sum_17[9] & q[7] /*13374*/;
  assign _2813_ = m_17[9] & _2811_ /*13373*/;
  assign r_17[16] = _2813_ | _2812_ /*13372*/;
  assign _2814_ = ~q[7] /*13371*/;
  assign _2815_ = sum_17[10] & q[7] /*13370*/;
  assign _2816_ = m_17[10] & _2814_ /*13369*/;
  assign r_17[17] = _2816_ | _2815_ /*13368*/;
  assign _2817_ = ~q[7] /*13367*/;
  assign _2818_ = sum_17[11] & q[7] /*13366*/;
  assign _2819_ = m_17[11] & _2817_ /*13365*/;
  assign r_17[18] = _2819_ | _2818_ /*13364*/;
  assign _2820_ = ~q[7] /*13363*/;
  assign _2821_ = sum_17[12] & q[7] /*13362*/;
  assign _2822_ = m_17[12] & _2820_ /*13361*/;
  assign r_17[19] = _2822_ | _2821_ /*13360*/;
  assign _2823_ = ~q[7] /*13359*/;
  assign _2824_ = sum_17[13] & q[7] /*13358*/;
  assign _2825_ = m_17[13] & _2823_ /*13357*/;
  assign r_17[20] = _2825_ | _2824_ /*13356*/;
  assign _2826_ = ~q[7] /*13355*/;
  assign _2827_ = sum_17[14] & q[7] /*13354*/;
  assign _2828_ = m_17[14] & _2826_ /*13353*/;
  assign r_17[21] = _2828_ | _2827_ /*13352*/;
  assign _2829_ = ~q[7] /*13351*/;
  assign _2830_ = sum_17[15] & q[7] /*13350*/;
  assign _2831_ = m_17[15] & _2829_ /*13349*/;
  assign r_17[22] = _2831_ | _2830_ /*13348*/;
  assign _2832_ = ~q[7] /*13347*/;
  assign _2833_ = sum_17[16] & q[7] /*13346*/;
  assign _2834_ = m_17[16] & _2832_ /*13345*/;
  assign r_17[23] = _2834_ | _2833_ /*13344*/;
  assign _2835_ = ~q[7] /*13343*/;
  assign _2836_ = sum_17[17] & q[7] /*13342*/;
  assign _2837_ = m_17[17] & _2835_ /*13341*/;
  assign r_17[24] = _2837_ | _2836_ /*13340*/;
  assign _2838_ = ~q[7] /*13339*/;
  assign _2839_ = sum_17[18] & q[7] /*13338*/;
  assign _2840_ = m_17[18] & _2838_ /*13337*/;
  assign r_17[25] = _2840_ | _2839_ /*13336*/;
  assign _2841_ = ~q[7] /*13335*/;
  assign _2842_ = sum_17[19] & q[7] /*13334*/;
  assign _2843_ = m_17[19] & _2841_ /*13333*/;
  assign r_17[26] = _2843_ | _2842_ /*13332*/;
  assign _2844_ = ~q[7] /*13331*/;
  assign _2845_ = sum_17[20] & q[7] /*13330*/;
  assign _2846_ = m_17[20] & _2844_ /*13329*/;
  assign r_17[27] = _2846_ | _2845_ /*13328*/;
  assign _2847_ = ~q[7] /*13327*/;
  assign _2848_ = sum_17[21] & q[7] /*13326*/;
  assign _2849_ = m_17[21] & _2847_ /*13325*/;
  assign r_17[28] = _2849_ | _2848_ /*13324*/;
  assign _2850_ = ~q[7] /*13323*/;
  assign _2851_ = sum_17[22] & q[7] /*13322*/;
  assign _2852_ = m_17[22] & _2850_ /*13321*/;
  assign r_17[29] = _2852_ | _2851_ /*13320*/;
  assign _2853_ = ~q[7] /*13319*/;
  assign _2854_ = sum_17[23] & q[7] /*13318*/;
  assign _2855_ = m_17[23] & _2853_ /*13317*/;
  assign r_17[30] = _2855_ | _2854_ /*13316*/;
assign r_17[0]= r_16[0] /*13315*/;
assign r_17[1]= r_16[1] /*13314*/;
assign r_17[2]= r_16[2] /*13313*/;
assign r_17[3]= r_16[3] /*13312*/;
assign r_17[4]= r_16[4] /*13311*/;
assign r_17[5]= r_16[5] /*13310*/;
assign r_17[6]= r_16[6] /*13309*/;
  assign inv_18[0] = ~div[0] /*13248*/;
  assign inv_18[1] = ~div[1] /*13247*/;
  assign inv_18[2] = ~div[2] /*13246*/;
  assign inv_18[3] = ~div[3] /*13245*/;
  assign inv_18[4] = ~div[4] /*13244*/;
  assign inv_18[5] = ~div[5] /*13243*/;
  assign inv_18[6] = ~div[6] /*13242*/;
  assign inv_18[7] = ~div[7] /*13241*/;
  assign inv_18[8] = ~div[8] /*13240*/;
  assign inv_18[9] = ~div[9] /*13239*/;
  assign inv_18[10] = ~div[10] /*13238*/;
  assign inv_18[11] = ~div[11] /*13237*/;
  assign inv_18[12] = ~div[12] /*13236*/;
  assign inv_18[13] = ~div[13] /*13235*/;
  assign inv_18[14] = ~div[14] /*13234*/;
  assign inv_18[15] = ~div[15] /*13233*/;
  assign inv_18[16] = ~div[16] /*13232*/;
  assign inv_18[17] = ~div[17] /*13231*/;
  assign inv_18[18] = ~div[18] /*13230*/;
  assign inv_18[19] = ~div[19] /*13229*/;
  assign inv_18[20] = ~div[20] /*13228*/;
  assign inv_18[21] = ~div[21] /*13227*/;
  assign inv_18[22] = ~div[22] /*13226*/;
assign inv_18[23] = oneWire /*13225*/;
  assign _2856_ = inv_18[0] ^ r_17[6] /*13223*/;
  assign sum_18[0] = _2856_ ^ oneWire /*13222*/;
  assign _2857_ = _2856_ & oneWire /*13221*/;
  assign _2858_ = inv_18[0] & r_17[6] /*13220*/;
  assign _2859_ = _2857_ | _2858_ /*13219*/;
  assign _2860_ = inv_18[1] ^ r_17[7] /*13218*/;
  assign sum_18[1] = _2860_ ^ _2859_ /*13217*/;
  assign _2861_ = _2860_ & _2859_ /*13216*/;
  assign _2862_ = inv_18[1] & r_17[7] /*13215*/;
  assign _2863_ = _2861_ | _2862_ /*13214*/;
  assign _2864_ = inv_18[2] ^ r_17[8] /*13212*/;
  assign sum_18[2] = _2864_ ^ _2863_ /*13211*/;
  assign _2865_ = _2864_ & _2863_ /*13210*/;
  assign _2866_ = inv_18[2] & r_17[8] /*13209*/;
  assign _2867_ = _2865_ | _2866_ /*13208*/;
  assign _2868_ = inv_18[3] ^ r_17[9] /*13206*/;
  assign sum_18[3] = _2868_ ^ _2867_ /*13205*/;
  assign _2869_ = _2868_ & _2867_ /*13204*/;
  assign _2870_ = inv_18[3] & r_17[9] /*13203*/;
  assign _2871_ = _2869_ | _2870_ /*13202*/;
  assign _2872_ = inv_18[4] ^ r_17[10] /*13200*/;
  assign sum_18[4] = _2872_ ^ _2871_ /*13199*/;
  assign _2873_ = _2872_ & _2871_ /*13198*/;
  assign _2874_ = inv_18[4] & r_17[10] /*13197*/;
  assign _2875_ = _2873_ | _2874_ /*13196*/;
  assign _2876_ = inv_18[5] ^ r_17[11] /*13194*/;
  assign sum_18[5] = _2876_ ^ _2875_ /*13193*/;
  assign _2877_ = _2876_ & _2875_ /*13192*/;
  assign _2878_ = inv_18[5] & r_17[11] /*13191*/;
  assign _2879_ = _2877_ | _2878_ /*13190*/;
  assign _2880_ = inv_18[6] ^ r_17[12] /*13188*/;
  assign sum_18[6] = _2880_ ^ _2879_ /*13187*/;
  assign _2881_ = _2880_ & _2879_ /*13186*/;
  assign _2882_ = inv_18[6] & r_17[12] /*13185*/;
  assign _2883_ = _2881_ | _2882_ /*13184*/;
  assign _2884_ = inv_18[7] ^ r_17[13] /*13182*/;
  assign sum_18[7] = _2884_ ^ _2883_ /*13181*/;
  assign _2885_ = _2884_ & _2883_ /*13180*/;
  assign _2886_ = inv_18[7] & r_17[13] /*13179*/;
  assign _2887_ = _2885_ | _2886_ /*13178*/;
  assign _2888_ = inv_18[8] ^ r_17[14] /*13176*/;
  assign sum_18[8] = _2888_ ^ _2887_ /*13175*/;
  assign _2889_ = _2888_ & _2887_ /*13174*/;
  assign _2890_ = inv_18[8] & r_17[14] /*13173*/;
  assign _2891_ = _2889_ | _2890_ /*13172*/;
  assign _2892_ = inv_18[9] ^ r_17[15] /*13170*/;
  assign sum_18[9] = _2892_ ^ _2891_ /*13169*/;
  assign _2893_ = _2892_ & _2891_ /*13168*/;
  assign _2894_ = inv_18[9] & r_17[15] /*13167*/;
  assign _2895_ = _2893_ | _2894_ /*13166*/;
  assign _2896_ = inv_18[10] ^ r_17[16] /*13164*/;
  assign sum_18[10] = _2896_ ^ _2895_ /*13163*/;
  assign _2897_ = _2896_ & _2895_ /*13162*/;
  assign _2898_ = inv_18[10] & r_17[16] /*13161*/;
  assign _2899_ = _2897_ | _2898_ /*13160*/;
  assign _2900_ = inv_18[11] ^ r_17[17] /*13158*/;
  assign sum_18[11] = _2900_ ^ _2899_ /*13157*/;
  assign _2901_ = _2900_ & _2899_ /*13156*/;
  assign _2902_ = inv_18[11] & r_17[17] /*13155*/;
  assign _2903_ = _2901_ | _2902_ /*13154*/;
  assign _2904_ = inv_18[12] ^ r_17[18] /*13152*/;
  assign sum_18[12] = _2904_ ^ _2903_ /*13151*/;
  assign _2905_ = _2904_ & _2903_ /*13150*/;
  assign _2906_ = inv_18[12] & r_17[18] /*13149*/;
  assign _2907_ = _2905_ | _2906_ /*13148*/;
  assign _2908_ = inv_18[13] ^ r_17[19] /*13146*/;
  assign sum_18[13] = _2908_ ^ _2907_ /*13145*/;
  assign _2909_ = _2908_ & _2907_ /*13144*/;
  assign _2910_ = inv_18[13] & r_17[19] /*13143*/;
  assign _2911_ = _2909_ | _2910_ /*13142*/;
  assign _2912_ = inv_18[14] ^ r_17[20] /*13140*/;
  assign sum_18[14] = _2912_ ^ _2911_ /*13139*/;
  assign _2913_ = _2912_ & _2911_ /*13138*/;
  assign _2914_ = inv_18[14] & r_17[20] /*13137*/;
  assign _2915_ = _2913_ | _2914_ /*13136*/;
  assign _2916_ = inv_18[15] ^ r_17[21] /*13134*/;
  assign sum_18[15] = _2916_ ^ _2915_ /*13133*/;
  assign _2917_ = _2916_ & _2915_ /*13132*/;
  assign _2918_ = inv_18[15] & r_17[21] /*13131*/;
  assign _2919_ = _2917_ | _2918_ /*13130*/;
  assign _2920_ = inv_18[16] ^ r_17[22] /*13128*/;
  assign sum_18[16] = _2920_ ^ _2919_ /*13127*/;
  assign _2921_ = _2920_ & _2919_ /*13126*/;
  assign _2922_ = inv_18[16] & r_17[22] /*13125*/;
  assign _2923_ = _2921_ | _2922_ /*13124*/;
  assign _2924_ = inv_18[17] ^ r_17[23] /*13122*/;
  assign sum_18[17] = _2924_ ^ _2923_ /*13121*/;
  assign _2925_ = _2924_ & _2923_ /*13120*/;
  assign _2926_ = inv_18[17] & r_17[23] /*13119*/;
  assign _2927_ = _2925_ | _2926_ /*13118*/;
  assign _2928_ = inv_18[18] ^ r_17[24] /*13116*/;
  assign sum_18[18] = _2928_ ^ _2927_ /*13115*/;
  assign _2929_ = _2928_ & _2927_ /*13114*/;
  assign _2930_ = inv_18[18] & r_17[24] /*13113*/;
  assign _2931_ = _2929_ | _2930_ /*13112*/;
  assign _2932_ = inv_18[19] ^ r_17[25] /*13110*/;
  assign sum_18[19] = _2932_ ^ _2931_ /*13109*/;
  assign _2933_ = _2932_ & _2931_ /*13108*/;
  assign _2934_ = inv_18[19] & r_17[25] /*13107*/;
  assign _2935_ = _2933_ | _2934_ /*13106*/;
  assign _2936_ = inv_18[20] ^ r_17[26] /*13104*/;
  assign sum_18[20] = _2936_ ^ _2935_ /*13103*/;
  assign _2937_ = _2936_ & _2935_ /*13102*/;
  assign _2938_ = inv_18[20] & r_17[26] /*13101*/;
  assign _2939_ = _2937_ | _2938_ /*13100*/;
  assign _2940_ = inv_18[21] ^ r_17[27] /*13098*/;
  assign sum_18[21] = _2940_ ^ _2939_ /*13097*/;
  assign _2941_ = _2940_ & _2939_ /*13096*/;
  assign _2942_ = inv_18[21] & r_17[27] /*13095*/;
  assign _2943_ = _2941_ | _2942_ /*13094*/;
  assign _2944_ = inv_18[22] ^ r_17[28] /*13092*/;
  assign sum_18[22] = _2944_ ^ _2943_ /*13091*/;
  assign _2945_ = _2944_ & _2943_ /*13090*/;
  assign _2946_ = inv_18[22] & r_17[28] /*13089*/;
  assign _2947_ = _2945_ | _2946_ /*13088*/;
  assign _2948_ = inv_18[23] ^ r_17[29] /*13086*/;
  assign sum_18[23] = _2948_ ^ _2947_ /*13085*/;
  assign _2949_ = _2948_ & _2947_ /*13084*/;
  assign _2950_ = inv_18[23] & r_17[29] /*13083*/;
  assign _2951_ = _2949_ | _2950_ /*13082*/;
  assign q[6] = ~sum_18[23] /*13101*/;
  assign m_18[0] = r_17[6] /*13100*/;
  assign m_18[1] = r_17[7] /*13099*/;
  assign m_18[2] = r_17[8] /*13098*/;
  assign m_18[3] = r_17[9] /*13097*/;
  assign m_18[4] = r_17[10] /*13096*/;
  assign m_18[5] = r_17[11] /*13095*/;
  assign m_18[6] = r_17[12] /*13094*/;
  assign m_18[7] = r_17[13] /*13093*/;
  assign m_18[8] = r_17[14] /*13092*/;
  assign m_18[9] = r_17[15] /*13091*/;
  assign m_18[10] = r_17[16] /*13090*/;
  assign m_18[11] = r_17[17] /*13089*/;
  assign m_18[12] = r_17[18] /*13088*/;
  assign m_18[13] = r_17[19] /*13087*/;
  assign m_18[14] = r_17[20] /*13086*/;
  assign m_18[15] = r_17[21] /*13085*/;
  assign m_18[16] = r_17[22] /*13084*/;
  assign m_18[17] = r_17[23] /*13083*/;
  assign m_18[18] = r_17[24] /*13082*/;
  assign m_18[19] = r_17[25] /*13081*/;
  assign m_18[20] = r_17[26] /*13080*/;
  assign m_18[21] = r_17[27] /*13079*/;
  assign m_18[22] = r_17[28] /*13078*/;
  assign m_18[23] = r_17[29] /*13077*/;
  assign _2952_ = ~q[6] /*13075*/;
  assign _2953_ = sum_18[0] & q[6] /*13074*/;
  assign _2954_ = m_18[0] & _2952_ /*13073*/;
  assign r_18[6] = _2954_ | _2953_ /*13072*/;
  assign _2955_ = ~q[6] /*13071*/;
  assign _2956_ = sum_18[1] & q[6] /*13070*/;
  assign _2957_ = m_18[1] & _2955_ /*13069*/;
  assign r_18[7] = _2957_ | _2956_ /*13068*/;
  assign _2958_ = ~q[6] /*13067*/;
  assign _2959_ = sum_18[2] & q[6] /*13066*/;
  assign _2960_ = m_18[2] & _2958_ /*13065*/;
  assign r_18[8] = _2960_ | _2959_ /*13064*/;
  assign _2961_ = ~q[6] /*13063*/;
  assign _2962_ = sum_18[3] & q[6] /*13062*/;
  assign _2963_ = m_18[3] & _2961_ /*13061*/;
  assign r_18[9] = _2963_ | _2962_ /*13060*/;
  assign _2964_ = ~q[6] /*13059*/;
  assign _2965_ = sum_18[4] & q[6] /*13058*/;
  assign _2966_ = m_18[4] & _2964_ /*13057*/;
  assign r_18[10] = _2966_ | _2965_ /*13056*/;
  assign _2967_ = ~q[6] /*13055*/;
  assign _2968_ = sum_18[5] & q[6] /*13054*/;
  assign _2969_ = m_18[5] & _2967_ /*13053*/;
  assign r_18[11] = _2969_ | _2968_ /*13052*/;
  assign _2970_ = ~q[6] /*13051*/;
  assign _2971_ = sum_18[6] & q[6] /*13050*/;
  assign _2972_ = m_18[6] & _2970_ /*13049*/;
  assign r_18[12] = _2972_ | _2971_ /*13048*/;
  assign _2973_ = ~q[6] /*13047*/;
  assign _2974_ = sum_18[7] & q[6] /*13046*/;
  assign _2975_ = m_18[7] & _2973_ /*13045*/;
  assign r_18[13] = _2975_ | _2974_ /*13044*/;
  assign _2976_ = ~q[6] /*13043*/;
  assign _2977_ = sum_18[8] & q[6] /*13042*/;
  assign _2978_ = m_18[8] & _2976_ /*13041*/;
  assign r_18[14] = _2978_ | _2977_ /*13040*/;
  assign _2979_ = ~q[6] /*13039*/;
  assign _2980_ = sum_18[9] & q[6] /*13038*/;
  assign _2981_ = m_18[9] & _2979_ /*13037*/;
  assign r_18[15] = _2981_ | _2980_ /*13036*/;
  assign _2982_ = ~q[6] /*13035*/;
  assign _2983_ = sum_18[10] & q[6] /*13034*/;
  assign _2984_ = m_18[10] & _2982_ /*13033*/;
  assign r_18[16] = _2984_ | _2983_ /*13032*/;
  assign _2985_ = ~q[6] /*13031*/;
  assign _2986_ = sum_18[11] & q[6] /*13030*/;
  assign _2987_ = m_18[11] & _2985_ /*13029*/;
  assign r_18[17] = _2987_ | _2986_ /*13028*/;
  assign _2988_ = ~q[6] /*13027*/;
  assign _2989_ = sum_18[12] & q[6] /*13026*/;
  assign _2990_ = m_18[12] & _2988_ /*13025*/;
  assign r_18[18] = _2990_ | _2989_ /*13024*/;
  assign _2991_ = ~q[6] /*13023*/;
  assign _2992_ = sum_18[13] & q[6] /*13022*/;
  assign _2993_ = m_18[13] & _2991_ /*13021*/;
  assign r_18[19] = _2993_ | _2992_ /*13020*/;
  assign _2994_ = ~q[6] /*13019*/;
  assign _2995_ = sum_18[14] & q[6] /*13018*/;
  assign _2996_ = m_18[14] & _2994_ /*13017*/;
  assign r_18[20] = _2996_ | _2995_ /*13016*/;
  assign _2997_ = ~q[6] /*13015*/;
  assign _2998_ = sum_18[15] & q[6] /*13014*/;
  assign _2999_ = m_18[15] & _2997_ /*13013*/;
  assign r_18[21] = _2999_ | _2998_ /*13012*/;
  assign _3000_ = ~q[6] /*13011*/;
  assign _3001_ = sum_18[16] & q[6] /*13010*/;
  assign _3002_ = m_18[16] & _3000_ /*13009*/;
  assign r_18[22] = _3002_ | _3001_ /*13008*/;
  assign _3003_ = ~q[6] /*13007*/;
  assign _3004_ = sum_18[17] & q[6] /*13006*/;
  assign _3005_ = m_18[17] & _3003_ /*13005*/;
  assign r_18[23] = _3005_ | _3004_ /*13004*/;
  assign _3006_ = ~q[6] /*13003*/;
  assign _3007_ = sum_18[18] & q[6] /*13002*/;
  assign _3008_ = m_18[18] & _3006_ /*13001*/;
  assign r_18[24] = _3008_ | _3007_ /*13000*/;
  assign _3009_ = ~q[6] /*12999*/;
  assign _3010_ = sum_18[19] & q[6] /*12998*/;
  assign _3011_ = m_18[19] & _3009_ /*12997*/;
  assign r_18[25] = _3011_ | _3010_ /*12996*/;
  assign _3012_ = ~q[6] /*12995*/;
  assign _3013_ = sum_18[20] & q[6] /*12994*/;
  assign _3014_ = m_18[20] & _3012_ /*12993*/;
  assign r_18[26] = _3014_ | _3013_ /*12992*/;
  assign _3015_ = ~q[6] /*12991*/;
  assign _3016_ = sum_18[21] & q[6] /*12990*/;
  assign _3017_ = m_18[21] & _3015_ /*12989*/;
  assign r_18[27] = _3017_ | _3016_ /*12988*/;
  assign _3018_ = ~q[6] /*12987*/;
  assign _3019_ = sum_18[22] & q[6] /*12986*/;
  assign _3020_ = m_18[22] & _3018_ /*12985*/;
  assign r_18[28] = _3020_ | _3019_ /*12984*/;
  assign _3021_ = ~q[6] /*12983*/;
  assign _3022_ = sum_18[23] & q[6] /*12982*/;
  assign _3023_ = m_18[23] & _3021_ /*12981*/;
  assign r_18[29] = _3023_ | _3022_ /*12980*/;
assign r_18[0]= r_17[0] /*12979*/;
assign r_18[1]= r_17[1] /*12978*/;
assign r_18[2]= r_17[2] /*12977*/;
assign r_18[3]= r_17[3] /*12976*/;
assign r_18[4]= r_17[4] /*12975*/;
assign r_18[5]= r_17[5] /*12974*/;
  assign inv_19[0] = ~div[0] /*12912*/;
  assign inv_19[1] = ~div[1] /*12911*/;
  assign inv_19[2] = ~div[2] /*12910*/;
  assign inv_19[3] = ~div[3] /*12909*/;
  assign inv_19[4] = ~div[4] /*12908*/;
  assign inv_19[5] = ~div[5] /*12907*/;
  assign inv_19[6] = ~div[6] /*12906*/;
  assign inv_19[7] = ~div[7] /*12905*/;
  assign inv_19[8] = ~div[8] /*12904*/;
  assign inv_19[9] = ~div[9] /*12903*/;
  assign inv_19[10] = ~div[10] /*12902*/;
  assign inv_19[11] = ~div[11] /*12901*/;
  assign inv_19[12] = ~div[12] /*12900*/;
  assign inv_19[13] = ~div[13] /*12899*/;
  assign inv_19[14] = ~div[14] /*12898*/;
  assign inv_19[15] = ~div[15] /*12897*/;
  assign inv_19[16] = ~div[16] /*12896*/;
  assign inv_19[17] = ~div[17] /*12895*/;
  assign inv_19[18] = ~div[18] /*12894*/;
  assign inv_19[19] = ~div[19] /*12893*/;
  assign inv_19[20] = ~div[20] /*12892*/;
  assign inv_19[21] = ~div[21] /*12891*/;
  assign inv_19[22] = ~div[22] /*12890*/;
assign inv_19[23] = oneWire /*12889*/;
  assign _3024_ = inv_19[0] ^ r_18[5] /*12887*/;
  assign sum_19[0] = _3024_ ^ oneWire /*12886*/;
  assign _3025_ = _3024_ & oneWire /*12885*/;
  assign _3026_ = inv_19[0] & r_18[5] /*12884*/;
  assign _3027_ = _3025_ | _3026_ /*12883*/;
  assign _3028_ = inv_19[1] ^ r_18[6] /*12882*/;
  assign sum_19[1] = _3028_ ^ _3027_ /*12881*/;
  assign _3029_ = _3028_ & _3027_ /*12880*/;
  assign _3030_ = inv_19[1] & r_18[6] /*12879*/;
  assign _3031_ = _3029_ | _3030_ /*12878*/;
  assign _3032_ = inv_19[2] ^ r_18[7] /*12876*/;
  assign sum_19[2] = _3032_ ^ _3031_ /*12875*/;
  assign _3033_ = _3032_ & _3031_ /*12874*/;
  assign _3034_ = inv_19[2] & r_18[7] /*12873*/;
  assign _3035_ = _3033_ | _3034_ /*12872*/;
  assign _3036_ = inv_19[3] ^ r_18[8] /*12870*/;
  assign sum_19[3] = _3036_ ^ _3035_ /*12869*/;
  assign _3037_ = _3036_ & _3035_ /*12868*/;
  assign _3038_ = inv_19[3] & r_18[8] /*12867*/;
  assign _3039_ = _3037_ | _3038_ /*12866*/;
  assign _3040_ = inv_19[4] ^ r_18[9] /*12864*/;
  assign sum_19[4] = _3040_ ^ _3039_ /*12863*/;
  assign _3041_ = _3040_ & _3039_ /*12862*/;
  assign _3042_ = inv_19[4] & r_18[9] /*12861*/;
  assign _3043_ = _3041_ | _3042_ /*12860*/;
  assign _3044_ = inv_19[5] ^ r_18[10] /*12858*/;
  assign sum_19[5] = _3044_ ^ _3043_ /*12857*/;
  assign _3045_ = _3044_ & _3043_ /*12856*/;
  assign _3046_ = inv_19[5] & r_18[10] /*12855*/;
  assign _3047_ = _3045_ | _3046_ /*12854*/;
  assign _3048_ = inv_19[6] ^ r_18[11] /*12852*/;
  assign sum_19[6] = _3048_ ^ _3047_ /*12851*/;
  assign _3049_ = _3048_ & _3047_ /*12850*/;
  assign _3050_ = inv_19[6] & r_18[11] /*12849*/;
  assign _3051_ = _3049_ | _3050_ /*12848*/;
  assign _3052_ = inv_19[7] ^ r_18[12] /*12846*/;
  assign sum_19[7] = _3052_ ^ _3051_ /*12845*/;
  assign _3053_ = _3052_ & _3051_ /*12844*/;
  assign _3054_ = inv_19[7] & r_18[12] /*12843*/;
  assign _3055_ = _3053_ | _3054_ /*12842*/;
  assign _3056_ = inv_19[8] ^ r_18[13] /*12840*/;
  assign sum_19[8] = _3056_ ^ _3055_ /*12839*/;
  assign _3057_ = _3056_ & _3055_ /*12838*/;
  assign _3058_ = inv_19[8] & r_18[13] /*12837*/;
  assign _3059_ = _3057_ | _3058_ /*12836*/;
  assign _3060_ = inv_19[9] ^ r_18[14] /*12834*/;
  assign sum_19[9] = _3060_ ^ _3059_ /*12833*/;
  assign _3061_ = _3060_ & _3059_ /*12832*/;
  assign _3062_ = inv_19[9] & r_18[14] /*12831*/;
  assign _3063_ = _3061_ | _3062_ /*12830*/;
  assign _3064_ = inv_19[10] ^ r_18[15] /*12828*/;
  assign sum_19[10] = _3064_ ^ _3063_ /*12827*/;
  assign _3065_ = _3064_ & _3063_ /*12826*/;
  assign _3066_ = inv_19[10] & r_18[15] /*12825*/;
  assign _3067_ = _3065_ | _3066_ /*12824*/;
  assign _3068_ = inv_19[11] ^ r_18[16] /*12822*/;
  assign sum_19[11] = _3068_ ^ _3067_ /*12821*/;
  assign _3069_ = _3068_ & _3067_ /*12820*/;
  assign _3070_ = inv_19[11] & r_18[16] /*12819*/;
  assign _3071_ = _3069_ | _3070_ /*12818*/;
  assign _3072_ = inv_19[12] ^ r_18[17] /*12816*/;
  assign sum_19[12] = _3072_ ^ _3071_ /*12815*/;
  assign _3073_ = _3072_ & _3071_ /*12814*/;
  assign _3074_ = inv_19[12] & r_18[17] /*12813*/;
  assign _3075_ = _3073_ | _3074_ /*12812*/;
  assign _3076_ = inv_19[13] ^ r_18[18] /*12810*/;
  assign sum_19[13] = _3076_ ^ _3075_ /*12809*/;
  assign _3077_ = _3076_ & _3075_ /*12808*/;
  assign _3078_ = inv_19[13] & r_18[18] /*12807*/;
  assign _3079_ = _3077_ | _3078_ /*12806*/;
  assign _3080_ = inv_19[14] ^ r_18[19] /*12804*/;
  assign sum_19[14] = _3080_ ^ _3079_ /*12803*/;
  assign _3081_ = _3080_ & _3079_ /*12802*/;
  assign _3082_ = inv_19[14] & r_18[19] /*12801*/;
  assign _3083_ = _3081_ | _3082_ /*12800*/;
  assign _3084_ = inv_19[15] ^ r_18[20] /*12798*/;
  assign sum_19[15] = _3084_ ^ _3083_ /*12797*/;
  assign _3085_ = _3084_ & _3083_ /*12796*/;
  assign _3086_ = inv_19[15] & r_18[20] /*12795*/;
  assign _3087_ = _3085_ | _3086_ /*12794*/;
  assign _3088_ = inv_19[16] ^ r_18[21] /*12792*/;
  assign sum_19[16] = _3088_ ^ _3087_ /*12791*/;
  assign _3089_ = _3088_ & _3087_ /*12790*/;
  assign _3090_ = inv_19[16] & r_18[21] /*12789*/;
  assign _3091_ = _3089_ | _3090_ /*12788*/;
  assign _3092_ = inv_19[17] ^ r_18[22] /*12786*/;
  assign sum_19[17] = _3092_ ^ _3091_ /*12785*/;
  assign _3093_ = _3092_ & _3091_ /*12784*/;
  assign _3094_ = inv_19[17] & r_18[22] /*12783*/;
  assign _3095_ = _3093_ | _3094_ /*12782*/;
  assign _3096_ = inv_19[18] ^ r_18[23] /*12780*/;
  assign sum_19[18] = _3096_ ^ _3095_ /*12779*/;
  assign _3097_ = _3096_ & _3095_ /*12778*/;
  assign _3098_ = inv_19[18] & r_18[23] /*12777*/;
  assign _3099_ = _3097_ | _3098_ /*12776*/;
  assign _3100_ = inv_19[19] ^ r_18[24] /*12774*/;
  assign sum_19[19] = _3100_ ^ _3099_ /*12773*/;
  assign _3101_ = _3100_ & _3099_ /*12772*/;
  assign _3102_ = inv_19[19] & r_18[24] /*12771*/;
  assign _3103_ = _3101_ | _3102_ /*12770*/;
  assign _3104_ = inv_19[20] ^ r_18[25] /*12768*/;
  assign sum_19[20] = _3104_ ^ _3103_ /*12767*/;
  assign _3105_ = _3104_ & _3103_ /*12766*/;
  assign _3106_ = inv_19[20] & r_18[25] /*12765*/;
  assign _3107_ = _3105_ | _3106_ /*12764*/;
  assign _3108_ = inv_19[21] ^ r_18[26] /*12762*/;
  assign sum_19[21] = _3108_ ^ _3107_ /*12761*/;
  assign _3109_ = _3108_ & _3107_ /*12760*/;
  assign _3110_ = inv_19[21] & r_18[26] /*12759*/;
  assign _3111_ = _3109_ | _3110_ /*12758*/;
  assign _3112_ = inv_19[22] ^ r_18[27] /*12756*/;
  assign sum_19[22] = _3112_ ^ _3111_ /*12755*/;
  assign _3113_ = _3112_ & _3111_ /*12754*/;
  assign _3114_ = inv_19[22] & r_18[27] /*12753*/;
  assign _3115_ = _3113_ | _3114_ /*12752*/;
  assign _3116_ = inv_19[23] ^ r_18[28] /*12750*/;
  assign sum_19[23] = _3116_ ^ _3115_ /*12749*/;
  assign _3117_ = _3116_ & _3115_ /*12748*/;
  assign _3118_ = inv_19[23] & r_18[28] /*12747*/;
  assign _3119_ = _3117_ | _3118_ /*12746*/;
  assign q[5] = ~sum_19[23] /*12765*/;
  assign m_19[0] = r_18[5] /*12764*/;
  assign m_19[1] = r_18[6] /*12763*/;
  assign m_19[2] = r_18[7] /*12762*/;
  assign m_19[3] = r_18[8] /*12761*/;
  assign m_19[4] = r_18[9] /*12760*/;
  assign m_19[5] = r_18[10] /*12759*/;
  assign m_19[6] = r_18[11] /*12758*/;
  assign m_19[7] = r_18[12] /*12757*/;
  assign m_19[8] = r_18[13] /*12756*/;
  assign m_19[9] = r_18[14] /*12755*/;
  assign m_19[10] = r_18[15] /*12754*/;
  assign m_19[11] = r_18[16] /*12753*/;
  assign m_19[12] = r_18[17] /*12752*/;
  assign m_19[13] = r_18[18] /*12751*/;
  assign m_19[14] = r_18[19] /*12750*/;
  assign m_19[15] = r_18[20] /*12749*/;
  assign m_19[16] = r_18[21] /*12748*/;
  assign m_19[17] = r_18[22] /*12747*/;
  assign m_19[18] = r_18[23] /*12746*/;
  assign m_19[19] = r_18[24] /*12745*/;
  assign m_19[20] = r_18[25] /*12744*/;
  assign m_19[21] = r_18[26] /*12743*/;
  assign m_19[22] = r_18[27] /*12742*/;
  assign m_19[23] = r_18[28] /*12741*/;
  assign _3120_ = ~q[5] /*12739*/;
  assign _3121_ = sum_19[0] & q[5] /*12738*/;
  assign _3122_ = m_19[0] & _3120_ /*12737*/;
  assign r_19[5] = _3122_ | _3121_ /*12736*/;
  assign _3123_ = ~q[5] /*12735*/;
  assign _3124_ = sum_19[1] & q[5] /*12734*/;
  assign _3125_ = m_19[1] & _3123_ /*12733*/;
  assign r_19[6] = _3125_ | _3124_ /*12732*/;
  assign _3126_ = ~q[5] /*12731*/;
  assign _3127_ = sum_19[2] & q[5] /*12730*/;
  assign _3128_ = m_19[2] & _3126_ /*12729*/;
  assign r_19[7] = _3128_ | _3127_ /*12728*/;
  assign _3129_ = ~q[5] /*12727*/;
  assign _3130_ = sum_19[3] & q[5] /*12726*/;
  assign _3131_ = m_19[3] & _3129_ /*12725*/;
  assign r_19[8] = _3131_ | _3130_ /*12724*/;
  assign _3132_ = ~q[5] /*12723*/;
  assign _3133_ = sum_19[4] & q[5] /*12722*/;
  assign _3134_ = m_19[4] & _3132_ /*12721*/;
  assign r_19[9] = _3134_ | _3133_ /*12720*/;
  assign _3135_ = ~q[5] /*12719*/;
  assign _3136_ = sum_19[5] & q[5] /*12718*/;
  assign _3137_ = m_19[5] & _3135_ /*12717*/;
  assign r_19[10] = _3137_ | _3136_ /*12716*/;
  assign _3138_ = ~q[5] /*12715*/;
  assign _3139_ = sum_19[6] & q[5] /*12714*/;
  assign _3140_ = m_19[6] & _3138_ /*12713*/;
  assign r_19[11] = _3140_ | _3139_ /*12712*/;
  assign _3141_ = ~q[5] /*12711*/;
  assign _3142_ = sum_19[7] & q[5] /*12710*/;
  assign _3143_ = m_19[7] & _3141_ /*12709*/;
  assign r_19[12] = _3143_ | _3142_ /*12708*/;
  assign _3144_ = ~q[5] /*12707*/;
  assign _3145_ = sum_19[8] & q[5] /*12706*/;
  assign _3146_ = m_19[8] & _3144_ /*12705*/;
  assign r_19[13] = _3146_ | _3145_ /*12704*/;
  assign _3147_ = ~q[5] /*12703*/;
  assign _3148_ = sum_19[9] & q[5] /*12702*/;
  assign _3149_ = m_19[9] & _3147_ /*12701*/;
  assign r_19[14] = _3149_ | _3148_ /*12700*/;
  assign _3150_ = ~q[5] /*12699*/;
  assign _3151_ = sum_19[10] & q[5] /*12698*/;
  assign _3152_ = m_19[10] & _3150_ /*12697*/;
  assign r_19[15] = _3152_ | _3151_ /*12696*/;
  assign _3153_ = ~q[5] /*12695*/;
  assign _3154_ = sum_19[11] & q[5] /*12694*/;
  assign _3155_ = m_19[11] & _3153_ /*12693*/;
  assign r_19[16] = _3155_ | _3154_ /*12692*/;
  assign _3156_ = ~q[5] /*12691*/;
  assign _3157_ = sum_19[12] & q[5] /*12690*/;
  assign _3158_ = m_19[12] & _3156_ /*12689*/;
  assign r_19[17] = _3158_ | _3157_ /*12688*/;
  assign _3159_ = ~q[5] /*12687*/;
  assign _3160_ = sum_19[13] & q[5] /*12686*/;
  assign _3161_ = m_19[13] & _3159_ /*12685*/;
  assign r_19[18] = _3161_ | _3160_ /*12684*/;
  assign _3162_ = ~q[5] /*12683*/;
  assign _3163_ = sum_19[14] & q[5] /*12682*/;
  assign _3164_ = m_19[14] & _3162_ /*12681*/;
  assign r_19[19] = _3164_ | _3163_ /*12680*/;
  assign _3165_ = ~q[5] /*12679*/;
  assign _3166_ = sum_19[15] & q[5] /*12678*/;
  assign _3167_ = m_19[15] & _3165_ /*12677*/;
  assign r_19[20] = _3167_ | _3166_ /*12676*/;
  assign _3168_ = ~q[5] /*12675*/;
  assign _3169_ = sum_19[16] & q[5] /*12674*/;
  assign _3170_ = m_19[16] & _3168_ /*12673*/;
  assign r_19[21] = _3170_ | _3169_ /*12672*/;
  assign _3171_ = ~q[5] /*12671*/;
  assign _3172_ = sum_19[17] & q[5] /*12670*/;
  assign _3173_ = m_19[17] & _3171_ /*12669*/;
  assign r_19[22] = _3173_ | _3172_ /*12668*/;
  assign _3174_ = ~q[5] /*12667*/;
  assign _3175_ = sum_19[18] & q[5] /*12666*/;
  assign _3176_ = m_19[18] & _3174_ /*12665*/;
  assign r_19[23] = _3176_ | _3175_ /*12664*/;
  assign _3177_ = ~q[5] /*12663*/;
  assign _3178_ = sum_19[19] & q[5] /*12662*/;
  assign _3179_ = m_19[19] & _3177_ /*12661*/;
  assign r_19[24] = _3179_ | _3178_ /*12660*/;
  assign _3180_ = ~q[5] /*12659*/;
  assign _3181_ = sum_19[20] & q[5] /*12658*/;
  assign _3182_ = m_19[20] & _3180_ /*12657*/;
  assign r_19[25] = _3182_ | _3181_ /*12656*/;
  assign _3183_ = ~q[5] /*12655*/;
  assign _3184_ = sum_19[21] & q[5] /*12654*/;
  assign _3185_ = m_19[21] & _3183_ /*12653*/;
  assign r_19[26] = _3185_ | _3184_ /*12652*/;
  assign _3186_ = ~q[5] /*12651*/;
  assign _3187_ = sum_19[22] & q[5] /*12650*/;
  assign _3188_ = m_19[22] & _3186_ /*12649*/;
  assign r_19[27] = _3188_ | _3187_ /*12648*/;
  assign _3189_ = ~q[5] /*12647*/;
  assign _3190_ = sum_19[23] & q[5] /*12646*/;
  assign _3191_ = m_19[23] & _3189_ /*12645*/;
  assign r_19[28] = _3191_ | _3190_ /*12644*/;
assign r_19[0]= r_18[0] /*12643*/;
assign r_19[1]= r_18[1] /*12642*/;
assign r_19[2]= r_18[2] /*12641*/;
assign r_19[3]= r_18[3] /*12640*/;
assign r_19[4]= r_18[4] /*12639*/;
  assign inv_20[0] = ~div[0] /*12576*/;
  assign inv_20[1] = ~div[1] /*12575*/;
  assign inv_20[2] = ~div[2] /*12574*/;
  assign inv_20[3] = ~div[3] /*12573*/;
  assign inv_20[4] = ~div[4] /*12572*/;
  assign inv_20[5] = ~div[5] /*12571*/;
  assign inv_20[6] = ~div[6] /*12570*/;
  assign inv_20[7] = ~div[7] /*12569*/;
  assign inv_20[8] = ~div[8] /*12568*/;
  assign inv_20[9] = ~div[9] /*12567*/;
  assign inv_20[10] = ~div[10] /*12566*/;
  assign inv_20[11] = ~div[11] /*12565*/;
  assign inv_20[12] = ~div[12] /*12564*/;
  assign inv_20[13] = ~div[13] /*12563*/;
  assign inv_20[14] = ~div[14] /*12562*/;
  assign inv_20[15] = ~div[15] /*12561*/;
  assign inv_20[16] = ~div[16] /*12560*/;
  assign inv_20[17] = ~div[17] /*12559*/;
  assign inv_20[18] = ~div[18] /*12558*/;
  assign inv_20[19] = ~div[19] /*12557*/;
  assign inv_20[20] = ~div[20] /*12556*/;
  assign inv_20[21] = ~div[21] /*12555*/;
  assign inv_20[22] = ~div[22] /*12554*/;
assign inv_20[23] = oneWire /*12553*/;
  assign _3192_ = inv_20[0] ^ r_19[4] /*12551*/;
  assign sum_20[0] = _3192_ ^ oneWire /*12550*/;
  assign _3193_ = _3192_ & oneWire /*12549*/;
  assign _3194_ = inv_20[0] & r_19[4] /*12548*/;
  assign _3195_ = _3193_ | _3194_ /*12547*/;
  assign _3196_ = inv_20[1] ^ r_19[5] /*12546*/;
  assign sum_20[1] = _3196_ ^ _3195_ /*12545*/;
  assign _3197_ = _3196_ & _3195_ /*12544*/;
  assign _3198_ = inv_20[1] & r_19[5] /*12543*/;
  assign _3199_ = _3197_ | _3198_ /*12542*/;
  assign _3200_ = inv_20[2] ^ r_19[6] /*12540*/;
  assign sum_20[2] = _3200_ ^ _3199_ /*12539*/;
  assign _3201_ = _3200_ & _3199_ /*12538*/;
  assign _3202_ = inv_20[2] & r_19[6] /*12537*/;
  assign _3203_ = _3201_ | _3202_ /*12536*/;
  assign _3204_ = inv_20[3] ^ r_19[7] /*12534*/;
  assign sum_20[3] = _3204_ ^ _3203_ /*12533*/;
  assign _3205_ = _3204_ & _3203_ /*12532*/;
  assign _3206_ = inv_20[3] & r_19[7] /*12531*/;
  assign _3207_ = _3205_ | _3206_ /*12530*/;
  assign _3208_ = inv_20[4] ^ r_19[8] /*12528*/;
  assign sum_20[4] = _3208_ ^ _3207_ /*12527*/;
  assign _3209_ = _3208_ & _3207_ /*12526*/;
  assign _3210_ = inv_20[4] & r_19[8] /*12525*/;
  assign _3211_ = _3209_ | _3210_ /*12524*/;
  assign _3212_ = inv_20[5] ^ r_19[9] /*12522*/;
  assign sum_20[5] = _3212_ ^ _3211_ /*12521*/;
  assign _3213_ = _3212_ & _3211_ /*12520*/;
  assign _3214_ = inv_20[5] & r_19[9] /*12519*/;
  assign _3215_ = _3213_ | _3214_ /*12518*/;
  assign _3216_ = inv_20[6] ^ r_19[10] /*12516*/;
  assign sum_20[6] = _3216_ ^ _3215_ /*12515*/;
  assign _3217_ = _3216_ & _3215_ /*12514*/;
  assign _3218_ = inv_20[6] & r_19[10] /*12513*/;
  assign _3219_ = _3217_ | _3218_ /*12512*/;
  assign _3220_ = inv_20[7] ^ r_19[11] /*12510*/;
  assign sum_20[7] = _3220_ ^ _3219_ /*12509*/;
  assign _3221_ = _3220_ & _3219_ /*12508*/;
  assign _3222_ = inv_20[7] & r_19[11] /*12507*/;
  assign _3223_ = _3221_ | _3222_ /*12506*/;
  assign _3224_ = inv_20[8] ^ r_19[12] /*12504*/;
  assign sum_20[8] = _3224_ ^ _3223_ /*12503*/;
  assign _3225_ = _3224_ & _3223_ /*12502*/;
  assign _3226_ = inv_20[8] & r_19[12] /*12501*/;
  assign _3227_ = _3225_ | _3226_ /*12500*/;
  assign _3228_ = inv_20[9] ^ r_19[13] /*12498*/;
  assign sum_20[9] = _3228_ ^ _3227_ /*12497*/;
  assign _3229_ = _3228_ & _3227_ /*12496*/;
  assign _3230_ = inv_20[9] & r_19[13] /*12495*/;
  assign _3231_ = _3229_ | _3230_ /*12494*/;
  assign _3232_ = inv_20[10] ^ r_19[14] /*12492*/;
  assign sum_20[10] = _3232_ ^ _3231_ /*12491*/;
  assign _3233_ = _3232_ & _3231_ /*12490*/;
  assign _3234_ = inv_20[10] & r_19[14] /*12489*/;
  assign _3235_ = _3233_ | _3234_ /*12488*/;
  assign _3236_ = inv_20[11] ^ r_19[15] /*12486*/;
  assign sum_20[11] = _3236_ ^ _3235_ /*12485*/;
  assign _3237_ = _3236_ & _3235_ /*12484*/;
  assign _3238_ = inv_20[11] & r_19[15] /*12483*/;
  assign _3239_ = _3237_ | _3238_ /*12482*/;
  assign _3240_ = inv_20[12] ^ r_19[16] /*12480*/;
  assign sum_20[12] = _3240_ ^ _3239_ /*12479*/;
  assign _3241_ = _3240_ & _3239_ /*12478*/;
  assign _3242_ = inv_20[12] & r_19[16] /*12477*/;
  assign _3243_ = _3241_ | _3242_ /*12476*/;
  assign _3244_ = inv_20[13] ^ r_19[17] /*12474*/;
  assign sum_20[13] = _3244_ ^ _3243_ /*12473*/;
  assign _3245_ = _3244_ & _3243_ /*12472*/;
  assign _3246_ = inv_20[13] & r_19[17] /*12471*/;
  assign _3247_ = _3245_ | _3246_ /*12470*/;
  assign _3248_ = inv_20[14] ^ r_19[18] /*12468*/;
  assign sum_20[14] = _3248_ ^ _3247_ /*12467*/;
  assign _3249_ = _3248_ & _3247_ /*12466*/;
  assign _3250_ = inv_20[14] & r_19[18] /*12465*/;
  assign _3251_ = _3249_ | _3250_ /*12464*/;
  assign _3252_ = inv_20[15] ^ r_19[19] /*12462*/;
  assign sum_20[15] = _3252_ ^ _3251_ /*12461*/;
  assign _3253_ = _3252_ & _3251_ /*12460*/;
  assign _3254_ = inv_20[15] & r_19[19] /*12459*/;
  assign _3255_ = _3253_ | _3254_ /*12458*/;
  assign _3256_ = inv_20[16] ^ r_19[20] /*12456*/;
  assign sum_20[16] = _3256_ ^ _3255_ /*12455*/;
  assign _3257_ = _3256_ & _3255_ /*12454*/;
  assign _3258_ = inv_20[16] & r_19[20] /*12453*/;
  assign _3259_ = _3257_ | _3258_ /*12452*/;
  assign _3260_ = inv_20[17] ^ r_19[21] /*12450*/;
  assign sum_20[17] = _3260_ ^ _3259_ /*12449*/;
  assign _3261_ = _3260_ & _3259_ /*12448*/;
  assign _3262_ = inv_20[17] & r_19[21] /*12447*/;
  assign _3263_ = _3261_ | _3262_ /*12446*/;
  assign _3264_ = inv_20[18] ^ r_19[22] /*12444*/;
  assign sum_20[18] = _3264_ ^ _3263_ /*12443*/;
  assign _3265_ = _3264_ & _3263_ /*12442*/;
  assign _3266_ = inv_20[18] & r_19[22] /*12441*/;
  assign _3267_ = _3265_ | _3266_ /*12440*/;
  assign _3268_ = inv_20[19] ^ r_19[23] /*12438*/;
  assign sum_20[19] = _3268_ ^ _3267_ /*12437*/;
  assign _3269_ = _3268_ & _3267_ /*12436*/;
  assign _3270_ = inv_20[19] & r_19[23] /*12435*/;
  assign _3271_ = _3269_ | _3270_ /*12434*/;
  assign _3272_ = inv_20[20] ^ r_19[24] /*12432*/;
  assign sum_20[20] = _3272_ ^ _3271_ /*12431*/;
  assign _3273_ = _3272_ & _3271_ /*12430*/;
  assign _3274_ = inv_20[20] & r_19[24] /*12429*/;
  assign _3275_ = _3273_ | _3274_ /*12428*/;
  assign _3276_ = inv_20[21] ^ r_19[25] /*12426*/;
  assign sum_20[21] = _3276_ ^ _3275_ /*12425*/;
  assign _3277_ = _3276_ & _3275_ /*12424*/;
  assign _3278_ = inv_20[21] & r_19[25] /*12423*/;
  assign _3279_ = _3277_ | _3278_ /*12422*/;
  assign _3280_ = inv_20[22] ^ r_19[26] /*12420*/;
  assign sum_20[22] = _3280_ ^ _3279_ /*12419*/;
  assign _3281_ = _3280_ & _3279_ /*12418*/;
  assign _3282_ = inv_20[22] & r_19[26] /*12417*/;
  assign _3283_ = _3281_ | _3282_ /*12416*/;
  assign _3284_ = inv_20[23] ^ r_19[27] /*12414*/;
  assign sum_20[23] = _3284_ ^ _3283_ /*12413*/;
  assign _3285_ = _3284_ & _3283_ /*12412*/;
  assign _3286_ = inv_20[23] & r_19[27] /*12411*/;
  assign _3287_ = _3285_ | _3286_ /*12410*/;
  assign q[4] = ~sum_20[23] /*12429*/;
  assign m_20[0] = r_19[4] /*12428*/;
  assign m_20[1] = r_19[5] /*12427*/;
  assign m_20[2] = r_19[6] /*12426*/;
  assign m_20[3] = r_19[7] /*12425*/;
  assign m_20[4] = r_19[8] /*12424*/;
  assign m_20[5] = r_19[9] /*12423*/;
  assign m_20[6] = r_19[10] /*12422*/;
  assign m_20[7] = r_19[11] /*12421*/;
  assign m_20[8] = r_19[12] /*12420*/;
  assign m_20[9] = r_19[13] /*12419*/;
  assign m_20[10] = r_19[14] /*12418*/;
  assign m_20[11] = r_19[15] /*12417*/;
  assign m_20[12] = r_19[16] /*12416*/;
  assign m_20[13] = r_19[17] /*12415*/;
  assign m_20[14] = r_19[18] /*12414*/;
  assign m_20[15] = r_19[19] /*12413*/;
  assign m_20[16] = r_19[20] /*12412*/;
  assign m_20[17] = r_19[21] /*12411*/;
  assign m_20[18] = r_19[22] /*12410*/;
  assign m_20[19] = r_19[23] /*12409*/;
  assign m_20[20] = r_19[24] /*12408*/;
  assign m_20[21] = r_19[25] /*12407*/;
  assign m_20[22] = r_19[26] /*12406*/;
  assign m_20[23] = r_19[27] /*12405*/;
  assign _3288_ = ~q[4] /*12403*/;
  assign _3289_ = sum_20[0] & q[4] /*12402*/;
  assign _3290_ = m_20[0] & _3288_ /*12401*/;
  assign r_20[4] = _3290_ | _3289_ /*12400*/;
  assign _3291_ = ~q[4] /*12399*/;
  assign _3292_ = sum_20[1] & q[4] /*12398*/;
  assign _3293_ = m_20[1] & _3291_ /*12397*/;
  assign r_20[5] = _3293_ | _3292_ /*12396*/;
  assign _3294_ = ~q[4] /*12395*/;
  assign _3295_ = sum_20[2] & q[4] /*12394*/;
  assign _3296_ = m_20[2] & _3294_ /*12393*/;
  assign r_20[6] = _3296_ | _3295_ /*12392*/;
  assign _3297_ = ~q[4] /*12391*/;
  assign _3298_ = sum_20[3] & q[4] /*12390*/;
  assign _3299_ = m_20[3] & _3297_ /*12389*/;
  assign r_20[7] = _3299_ | _3298_ /*12388*/;
  assign _3300_ = ~q[4] /*12387*/;
  assign _3301_ = sum_20[4] & q[4] /*12386*/;
  assign _3302_ = m_20[4] & _3300_ /*12385*/;
  assign r_20[8] = _3302_ | _3301_ /*12384*/;
  assign _3303_ = ~q[4] /*12383*/;
  assign _3304_ = sum_20[5] & q[4] /*12382*/;
  assign _3305_ = m_20[5] & _3303_ /*12381*/;
  assign r_20[9] = _3305_ | _3304_ /*12380*/;
  assign _3306_ = ~q[4] /*12379*/;
  assign _3307_ = sum_20[6] & q[4] /*12378*/;
  assign _3308_ = m_20[6] & _3306_ /*12377*/;
  assign r_20[10] = _3308_ | _3307_ /*12376*/;
  assign _3309_ = ~q[4] /*12375*/;
  assign _3310_ = sum_20[7] & q[4] /*12374*/;
  assign _3311_ = m_20[7] & _3309_ /*12373*/;
  assign r_20[11] = _3311_ | _3310_ /*12372*/;
  assign _3312_ = ~q[4] /*12371*/;
  assign _3313_ = sum_20[8] & q[4] /*12370*/;
  assign _3314_ = m_20[8] & _3312_ /*12369*/;
  assign r_20[12] = _3314_ | _3313_ /*12368*/;
  assign _3315_ = ~q[4] /*12367*/;
  assign _3316_ = sum_20[9] & q[4] /*12366*/;
  assign _3317_ = m_20[9] & _3315_ /*12365*/;
  assign r_20[13] = _3317_ | _3316_ /*12364*/;
  assign _3318_ = ~q[4] /*12363*/;
  assign _3319_ = sum_20[10] & q[4] /*12362*/;
  assign _3320_ = m_20[10] & _3318_ /*12361*/;
  assign r_20[14] = _3320_ | _3319_ /*12360*/;
  assign _3321_ = ~q[4] /*12359*/;
  assign _3322_ = sum_20[11] & q[4] /*12358*/;
  assign _3323_ = m_20[11] & _3321_ /*12357*/;
  assign r_20[15] = _3323_ | _3322_ /*12356*/;
  assign _3324_ = ~q[4] /*12355*/;
  assign _3325_ = sum_20[12] & q[4] /*12354*/;
  assign _3326_ = m_20[12] & _3324_ /*12353*/;
  assign r_20[16] = _3326_ | _3325_ /*12352*/;
  assign _3327_ = ~q[4] /*12351*/;
  assign _3328_ = sum_20[13] & q[4] /*12350*/;
  assign _3329_ = m_20[13] & _3327_ /*12349*/;
  assign r_20[17] = _3329_ | _3328_ /*12348*/;
  assign _3330_ = ~q[4] /*12347*/;
  assign _3331_ = sum_20[14] & q[4] /*12346*/;
  assign _3332_ = m_20[14] & _3330_ /*12345*/;
  assign r_20[18] = _3332_ | _3331_ /*12344*/;
  assign _3333_ = ~q[4] /*12343*/;
  assign _3334_ = sum_20[15] & q[4] /*12342*/;
  assign _3335_ = m_20[15] & _3333_ /*12341*/;
  assign r_20[19] = _3335_ | _3334_ /*12340*/;
  assign _3336_ = ~q[4] /*12339*/;
  assign _3337_ = sum_20[16] & q[4] /*12338*/;
  assign _3338_ = m_20[16] & _3336_ /*12337*/;
  assign r_20[20] = _3338_ | _3337_ /*12336*/;
  assign _3339_ = ~q[4] /*12335*/;
  assign _3340_ = sum_20[17] & q[4] /*12334*/;
  assign _3341_ = m_20[17] & _3339_ /*12333*/;
  assign r_20[21] = _3341_ | _3340_ /*12332*/;
  assign _3342_ = ~q[4] /*12331*/;
  assign _3343_ = sum_20[18] & q[4] /*12330*/;
  assign _3344_ = m_20[18] & _3342_ /*12329*/;
  assign r_20[22] = _3344_ | _3343_ /*12328*/;
  assign _3345_ = ~q[4] /*12327*/;
  assign _3346_ = sum_20[19] & q[4] /*12326*/;
  assign _3347_ = m_20[19] & _3345_ /*12325*/;
  assign r_20[23] = _3347_ | _3346_ /*12324*/;
  assign _3348_ = ~q[4] /*12323*/;
  assign _3349_ = sum_20[20] & q[4] /*12322*/;
  assign _3350_ = m_20[20] & _3348_ /*12321*/;
  assign r_20[24] = _3350_ | _3349_ /*12320*/;
  assign _3351_ = ~q[4] /*12319*/;
  assign _3352_ = sum_20[21] & q[4] /*12318*/;
  assign _3353_ = m_20[21] & _3351_ /*12317*/;
  assign r_20[25] = _3353_ | _3352_ /*12316*/;
  assign _3354_ = ~q[4] /*12315*/;
  assign _3355_ = sum_20[22] & q[4] /*12314*/;
  assign _3356_ = m_20[22] & _3354_ /*12313*/;
  assign r_20[26] = _3356_ | _3355_ /*12312*/;
  assign _3357_ = ~q[4] /*12311*/;
  assign _3358_ = sum_20[23] & q[4] /*12310*/;
  assign _3359_ = m_20[23] & _3357_ /*12309*/;
  assign r_20[27] = _3359_ | _3358_ /*12308*/;
assign r_20[0]= r_19[0] /*12307*/;
assign r_20[1]= r_19[1] /*12306*/;
assign r_20[2]= r_19[2] /*12305*/;
assign r_20[3]= r_19[3] /*12304*/;
  assign inv_21[0] = ~div[0] /*12240*/;
  assign inv_21[1] = ~div[1] /*12239*/;
  assign inv_21[2] = ~div[2] /*12238*/;
  assign inv_21[3] = ~div[3] /*12237*/;
  assign inv_21[4] = ~div[4] /*12236*/;
  assign inv_21[5] = ~div[5] /*12235*/;
  assign inv_21[6] = ~div[6] /*12234*/;
  assign inv_21[7] = ~div[7] /*12233*/;
  assign inv_21[8] = ~div[8] /*12232*/;
  assign inv_21[9] = ~div[9] /*12231*/;
  assign inv_21[10] = ~div[10] /*12230*/;
  assign inv_21[11] = ~div[11] /*12229*/;
  assign inv_21[12] = ~div[12] /*12228*/;
  assign inv_21[13] = ~div[13] /*12227*/;
  assign inv_21[14] = ~div[14] /*12226*/;
  assign inv_21[15] = ~div[15] /*12225*/;
  assign inv_21[16] = ~div[16] /*12224*/;
  assign inv_21[17] = ~div[17] /*12223*/;
  assign inv_21[18] = ~div[18] /*12222*/;
  assign inv_21[19] = ~div[19] /*12221*/;
  assign inv_21[20] = ~div[20] /*12220*/;
  assign inv_21[21] = ~div[21] /*12219*/;
  assign inv_21[22] = ~div[22] /*12218*/;
assign inv_21[23] = oneWire /*12217*/;
  assign _3360_ = inv_21[0] ^ r_20[3] /*12215*/;
  assign sum_21[0] = _3360_ ^ oneWire /*12214*/;
  assign _3361_ = _3360_ & oneWire /*12213*/;
  assign _3362_ = inv_21[0] & r_20[3] /*12212*/;
  assign _3363_ = _3361_ | _3362_ /*12211*/;
  assign _3364_ = inv_21[1] ^ r_20[4] /*12210*/;
  assign sum_21[1] = _3364_ ^ _3363_ /*12209*/;
  assign _3365_ = _3364_ & _3363_ /*12208*/;
  assign _3366_ = inv_21[1] & r_20[4] /*12207*/;
  assign _3367_ = _3365_ | _3366_ /*12206*/;
  assign _3368_ = inv_21[2] ^ r_20[5] /*12204*/;
  assign sum_21[2] = _3368_ ^ _3367_ /*12203*/;
  assign _3369_ = _3368_ & _3367_ /*12202*/;
  assign _3370_ = inv_21[2] & r_20[5] /*12201*/;
  assign _3371_ = _3369_ | _3370_ /*12200*/;
  assign _3372_ = inv_21[3] ^ r_20[6] /*12198*/;
  assign sum_21[3] = _3372_ ^ _3371_ /*12197*/;
  assign _3373_ = _3372_ & _3371_ /*12196*/;
  assign _3374_ = inv_21[3] & r_20[6] /*12195*/;
  assign _3375_ = _3373_ | _3374_ /*12194*/;
  assign _3376_ = inv_21[4] ^ r_20[7] /*12192*/;
  assign sum_21[4] = _3376_ ^ _3375_ /*12191*/;
  assign _3377_ = _3376_ & _3375_ /*12190*/;
  assign _3378_ = inv_21[4] & r_20[7] /*12189*/;
  assign _3379_ = _3377_ | _3378_ /*12188*/;
  assign _3380_ = inv_21[5] ^ r_20[8] /*12186*/;
  assign sum_21[5] = _3380_ ^ _3379_ /*12185*/;
  assign _3381_ = _3380_ & _3379_ /*12184*/;
  assign _3382_ = inv_21[5] & r_20[8] /*12183*/;
  assign _3383_ = _3381_ | _3382_ /*12182*/;
  assign _3384_ = inv_21[6] ^ r_20[9] /*12180*/;
  assign sum_21[6] = _3384_ ^ _3383_ /*12179*/;
  assign _3385_ = _3384_ & _3383_ /*12178*/;
  assign _3386_ = inv_21[6] & r_20[9] /*12177*/;
  assign _3387_ = _3385_ | _3386_ /*12176*/;
  assign _3388_ = inv_21[7] ^ r_20[10] /*12174*/;
  assign sum_21[7] = _3388_ ^ _3387_ /*12173*/;
  assign _3389_ = _3388_ & _3387_ /*12172*/;
  assign _3390_ = inv_21[7] & r_20[10] /*12171*/;
  assign _3391_ = _3389_ | _3390_ /*12170*/;
  assign _3392_ = inv_21[8] ^ r_20[11] /*12168*/;
  assign sum_21[8] = _3392_ ^ _3391_ /*12167*/;
  assign _3393_ = _3392_ & _3391_ /*12166*/;
  assign _3394_ = inv_21[8] & r_20[11] /*12165*/;
  assign _3395_ = _3393_ | _3394_ /*12164*/;
  assign _3396_ = inv_21[9] ^ r_20[12] /*12162*/;
  assign sum_21[9] = _3396_ ^ _3395_ /*12161*/;
  assign _3397_ = _3396_ & _3395_ /*12160*/;
  assign _3398_ = inv_21[9] & r_20[12] /*12159*/;
  assign _3399_ = _3397_ | _3398_ /*12158*/;
  assign _3400_ = inv_21[10] ^ r_20[13] /*12156*/;
  assign sum_21[10] = _3400_ ^ _3399_ /*12155*/;
  assign _3401_ = _3400_ & _3399_ /*12154*/;
  assign _3402_ = inv_21[10] & r_20[13] /*12153*/;
  assign _3403_ = _3401_ | _3402_ /*12152*/;
  assign _3404_ = inv_21[11] ^ r_20[14] /*12150*/;
  assign sum_21[11] = _3404_ ^ _3403_ /*12149*/;
  assign _3405_ = _3404_ & _3403_ /*12148*/;
  assign _3406_ = inv_21[11] & r_20[14] /*12147*/;
  assign _3407_ = _3405_ | _3406_ /*12146*/;
  assign _3408_ = inv_21[12] ^ r_20[15] /*12144*/;
  assign sum_21[12] = _3408_ ^ _3407_ /*12143*/;
  assign _3409_ = _3408_ & _3407_ /*12142*/;
  assign _3410_ = inv_21[12] & r_20[15] /*12141*/;
  assign _3411_ = _3409_ | _3410_ /*12140*/;
  assign _3412_ = inv_21[13] ^ r_20[16] /*12138*/;
  assign sum_21[13] = _3412_ ^ _3411_ /*12137*/;
  assign _3413_ = _3412_ & _3411_ /*12136*/;
  assign _3414_ = inv_21[13] & r_20[16] /*12135*/;
  assign _3415_ = _3413_ | _3414_ /*12134*/;
  assign _3416_ = inv_21[14] ^ r_20[17] /*12132*/;
  assign sum_21[14] = _3416_ ^ _3415_ /*12131*/;
  assign _3417_ = _3416_ & _3415_ /*12130*/;
  assign _3418_ = inv_21[14] & r_20[17] /*12129*/;
  assign _3419_ = _3417_ | _3418_ /*12128*/;
  assign _3420_ = inv_21[15] ^ r_20[18] /*12126*/;
  assign sum_21[15] = _3420_ ^ _3419_ /*12125*/;
  assign _3421_ = _3420_ & _3419_ /*12124*/;
  assign _3422_ = inv_21[15] & r_20[18] /*12123*/;
  assign _3423_ = _3421_ | _3422_ /*12122*/;
  assign _3424_ = inv_21[16] ^ r_20[19] /*12120*/;
  assign sum_21[16] = _3424_ ^ _3423_ /*12119*/;
  assign _3425_ = _3424_ & _3423_ /*12118*/;
  assign _3426_ = inv_21[16] & r_20[19] /*12117*/;
  assign _3427_ = _3425_ | _3426_ /*12116*/;
  assign _3428_ = inv_21[17] ^ r_20[20] /*12114*/;
  assign sum_21[17] = _3428_ ^ _3427_ /*12113*/;
  assign _3429_ = _3428_ & _3427_ /*12112*/;
  assign _3430_ = inv_21[17] & r_20[20] /*12111*/;
  assign _3431_ = _3429_ | _3430_ /*12110*/;
  assign _3432_ = inv_21[18] ^ r_20[21] /*12108*/;
  assign sum_21[18] = _3432_ ^ _3431_ /*12107*/;
  assign _3433_ = _3432_ & _3431_ /*12106*/;
  assign _3434_ = inv_21[18] & r_20[21] /*12105*/;
  assign _3435_ = _3433_ | _3434_ /*12104*/;
  assign _3436_ = inv_21[19] ^ r_20[22] /*12102*/;
  assign sum_21[19] = _3436_ ^ _3435_ /*12101*/;
  assign _3437_ = _3436_ & _3435_ /*12100*/;
  assign _3438_ = inv_21[19] & r_20[22] /*12099*/;
  assign _3439_ = _3437_ | _3438_ /*12098*/;
  assign _3440_ = inv_21[20] ^ r_20[23] /*12096*/;
  assign sum_21[20] = _3440_ ^ _3439_ /*12095*/;
  assign _3441_ = _3440_ & _3439_ /*12094*/;
  assign _3442_ = inv_21[20] & r_20[23] /*12093*/;
  assign _3443_ = _3441_ | _3442_ /*12092*/;
  assign _3444_ = inv_21[21] ^ r_20[24] /*12090*/;
  assign sum_21[21] = _3444_ ^ _3443_ /*12089*/;
  assign _3445_ = _3444_ & _3443_ /*12088*/;
  assign _3446_ = inv_21[21] & r_20[24] /*12087*/;
  assign _3447_ = _3445_ | _3446_ /*12086*/;
  assign _3448_ = inv_21[22] ^ r_20[25] /*12084*/;
  assign sum_21[22] = _3448_ ^ _3447_ /*12083*/;
  assign _3449_ = _3448_ & _3447_ /*12082*/;
  assign _3450_ = inv_21[22] & r_20[25] /*12081*/;
  assign _3451_ = _3449_ | _3450_ /*12080*/;
  assign _3452_ = inv_21[23] ^ r_20[26] /*12078*/;
  assign sum_21[23] = _3452_ ^ _3451_ /*12077*/;
  assign _3453_ = _3452_ & _3451_ /*12076*/;
  assign _3454_ = inv_21[23] & r_20[26] /*12075*/;
  assign _3455_ = _3453_ | _3454_ /*12074*/;
  assign q[3] = ~sum_21[23] /*12093*/;
  assign m_21[0] = r_20[3] /*12092*/;
  assign m_21[1] = r_20[4] /*12091*/;
  assign m_21[2] = r_20[5] /*12090*/;
  assign m_21[3] = r_20[6] /*12089*/;
  assign m_21[4] = r_20[7] /*12088*/;
  assign m_21[5] = r_20[8] /*12087*/;
  assign m_21[6] = r_20[9] /*12086*/;
  assign m_21[7] = r_20[10] /*12085*/;
  assign m_21[8] = r_20[11] /*12084*/;
  assign m_21[9] = r_20[12] /*12083*/;
  assign m_21[10] = r_20[13] /*12082*/;
  assign m_21[11] = r_20[14] /*12081*/;
  assign m_21[12] = r_20[15] /*12080*/;
  assign m_21[13] = r_20[16] /*12079*/;
  assign m_21[14] = r_20[17] /*12078*/;
  assign m_21[15] = r_20[18] /*12077*/;
  assign m_21[16] = r_20[19] /*12076*/;
  assign m_21[17] = r_20[20] /*12075*/;
  assign m_21[18] = r_20[21] /*12074*/;
  assign m_21[19] = r_20[22] /*12073*/;
  assign m_21[20] = r_20[23] /*12072*/;
  assign m_21[21] = r_20[24] /*12071*/;
  assign m_21[22] = r_20[25] /*12070*/;
  assign m_21[23] = r_20[26] /*12069*/;
  assign _3456_ = ~q[3] /*12067*/;
  assign _3457_ = sum_21[0] & q[3] /*12066*/;
  assign _3458_ = m_21[0] & _3456_ /*12065*/;
  assign r_21[3] = _3458_ | _3457_ /*12064*/;
  assign _3459_ = ~q[3] /*12063*/;
  assign _3460_ = sum_21[1] & q[3] /*12062*/;
  assign _3461_ = m_21[1] & _3459_ /*12061*/;
  assign r_21[4] = _3461_ | _3460_ /*12060*/;
  assign _3462_ = ~q[3] /*12059*/;
  assign _3463_ = sum_21[2] & q[3] /*12058*/;
  assign _3464_ = m_21[2] & _3462_ /*12057*/;
  assign r_21[5] = _3464_ | _3463_ /*12056*/;
  assign _3465_ = ~q[3] /*12055*/;
  assign _3466_ = sum_21[3] & q[3] /*12054*/;
  assign _3467_ = m_21[3] & _3465_ /*12053*/;
  assign r_21[6] = _3467_ | _3466_ /*12052*/;
  assign _3468_ = ~q[3] /*12051*/;
  assign _3469_ = sum_21[4] & q[3] /*12050*/;
  assign _3470_ = m_21[4] & _3468_ /*12049*/;
  assign r_21[7] = _3470_ | _3469_ /*12048*/;
  assign _3471_ = ~q[3] /*12047*/;
  assign _3472_ = sum_21[5] & q[3] /*12046*/;
  assign _3473_ = m_21[5] & _3471_ /*12045*/;
  assign r_21[8] = _3473_ | _3472_ /*12044*/;
  assign _3474_ = ~q[3] /*12043*/;
  assign _3475_ = sum_21[6] & q[3] /*12042*/;
  assign _3476_ = m_21[6] & _3474_ /*12041*/;
  assign r_21[9] = _3476_ | _3475_ /*12040*/;
  assign _3477_ = ~q[3] /*12039*/;
  assign _3478_ = sum_21[7] & q[3] /*12038*/;
  assign _3479_ = m_21[7] & _3477_ /*12037*/;
  assign r_21[10] = _3479_ | _3478_ /*12036*/;
  assign _3480_ = ~q[3] /*12035*/;
  assign _3481_ = sum_21[8] & q[3] /*12034*/;
  assign _3482_ = m_21[8] & _3480_ /*12033*/;
  assign r_21[11] = _3482_ | _3481_ /*12032*/;
  assign _3483_ = ~q[3] /*12031*/;
  assign _3484_ = sum_21[9] & q[3] /*12030*/;
  assign _3485_ = m_21[9] & _3483_ /*12029*/;
  assign r_21[12] = _3485_ | _3484_ /*12028*/;
  assign _3486_ = ~q[3] /*12027*/;
  assign _3487_ = sum_21[10] & q[3] /*12026*/;
  assign _3488_ = m_21[10] & _3486_ /*12025*/;
  assign r_21[13] = _3488_ | _3487_ /*12024*/;
  assign _3489_ = ~q[3] /*12023*/;
  assign _3490_ = sum_21[11] & q[3] /*12022*/;
  assign _3491_ = m_21[11] & _3489_ /*12021*/;
  assign r_21[14] = _3491_ | _3490_ /*12020*/;
  assign _3492_ = ~q[3] /*12019*/;
  assign _3493_ = sum_21[12] & q[3] /*12018*/;
  assign _3494_ = m_21[12] & _3492_ /*12017*/;
  assign r_21[15] = _3494_ | _3493_ /*12016*/;
  assign _3495_ = ~q[3] /*12015*/;
  assign _3496_ = sum_21[13] & q[3] /*12014*/;
  assign _3497_ = m_21[13] & _3495_ /*12013*/;
  assign r_21[16] = _3497_ | _3496_ /*12012*/;
  assign _3498_ = ~q[3] /*12011*/;
  assign _3499_ = sum_21[14] & q[3] /*12010*/;
  assign _3500_ = m_21[14] & _3498_ /*12009*/;
  assign r_21[17] = _3500_ | _3499_ /*12008*/;
  assign _3501_ = ~q[3] /*12007*/;
  assign _3502_ = sum_21[15] & q[3] /*12006*/;
  assign _3503_ = m_21[15] & _3501_ /*12005*/;
  assign r_21[18] = _3503_ | _3502_ /*12004*/;
  assign _3504_ = ~q[3] /*12003*/;
  assign _3505_ = sum_21[16] & q[3] /*12002*/;
  assign _3506_ = m_21[16] & _3504_ /*12001*/;
  assign r_21[19] = _3506_ | _3505_ /*12000*/;
  assign _3507_ = ~q[3] /*11999*/;
  assign _3508_ = sum_21[17] & q[3] /*11998*/;
  assign _3509_ = m_21[17] & _3507_ /*11997*/;
  assign r_21[20] = _3509_ | _3508_ /*11996*/;
  assign _3510_ = ~q[3] /*11995*/;
  assign _3511_ = sum_21[18] & q[3] /*11994*/;
  assign _3512_ = m_21[18] & _3510_ /*11993*/;
  assign r_21[21] = _3512_ | _3511_ /*11992*/;
  assign _3513_ = ~q[3] /*11991*/;
  assign _3514_ = sum_21[19] & q[3] /*11990*/;
  assign _3515_ = m_21[19] & _3513_ /*11989*/;
  assign r_21[22] = _3515_ | _3514_ /*11988*/;
  assign _3516_ = ~q[3] /*11987*/;
  assign _3517_ = sum_21[20] & q[3] /*11986*/;
  assign _3518_ = m_21[20] & _3516_ /*11985*/;
  assign r_21[23] = _3518_ | _3517_ /*11984*/;
  assign _3519_ = ~q[3] /*11983*/;
  assign _3520_ = sum_21[21] & q[3] /*11982*/;
  assign _3521_ = m_21[21] & _3519_ /*11981*/;
  assign r_21[24] = _3521_ | _3520_ /*11980*/;
  assign _3522_ = ~q[3] /*11979*/;
  assign _3523_ = sum_21[22] & q[3] /*11978*/;
  assign _3524_ = m_21[22] & _3522_ /*11977*/;
  assign r_21[25] = _3524_ | _3523_ /*11976*/;
  assign _3525_ = ~q[3] /*11975*/;
  assign _3526_ = sum_21[23] & q[3] /*11974*/;
  assign _3527_ = m_21[23] & _3525_ /*11973*/;
  assign r_21[26] = _3527_ | _3526_ /*11972*/;
assign r_21[0]= r_20[0] /*11971*/;
assign r_21[1]= r_20[1] /*11970*/;
assign r_21[2]= r_20[2] /*11969*/;
  assign inv_22[0] = ~div[0] /*11904*/;
  assign inv_22[1] = ~div[1] /*11903*/;
  assign inv_22[2] = ~div[2] /*11902*/;
  assign inv_22[3] = ~div[3] /*11901*/;
  assign inv_22[4] = ~div[4] /*11900*/;
  assign inv_22[5] = ~div[5] /*11899*/;
  assign inv_22[6] = ~div[6] /*11898*/;
  assign inv_22[7] = ~div[7] /*11897*/;
  assign inv_22[8] = ~div[8] /*11896*/;
  assign inv_22[9] = ~div[9] /*11895*/;
  assign inv_22[10] = ~div[10] /*11894*/;
  assign inv_22[11] = ~div[11] /*11893*/;
  assign inv_22[12] = ~div[12] /*11892*/;
  assign inv_22[13] = ~div[13] /*11891*/;
  assign inv_22[14] = ~div[14] /*11890*/;
  assign inv_22[15] = ~div[15] /*11889*/;
  assign inv_22[16] = ~div[16] /*11888*/;
  assign inv_22[17] = ~div[17] /*11887*/;
  assign inv_22[18] = ~div[18] /*11886*/;
  assign inv_22[19] = ~div[19] /*11885*/;
  assign inv_22[20] = ~div[20] /*11884*/;
  assign inv_22[21] = ~div[21] /*11883*/;
  assign inv_22[22] = ~div[22] /*11882*/;
assign inv_22[23] = oneWire /*11881*/;
  assign _3528_ = inv_22[0] ^ r_21[2] /*11879*/;
  assign sum_22[0] = _3528_ ^ oneWire /*11878*/;
  assign _3529_ = _3528_ & oneWire /*11877*/;
  assign _3530_ = inv_22[0] & r_21[2] /*11876*/;
  assign _3531_ = _3529_ | _3530_ /*11875*/;
  assign _3532_ = inv_22[1] ^ r_21[3] /*11874*/;
  assign sum_22[1] = _3532_ ^ _3531_ /*11873*/;
  assign _3533_ = _3532_ & _3531_ /*11872*/;
  assign _3534_ = inv_22[1] & r_21[3] /*11871*/;
  assign _3535_ = _3533_ | _3534_ /*11870*/;
  assign _3536_ = inv_22[2] ^ r_21[4] /*11868*/;
  assign sum_22[2] = _3536_ ^ _3535_ /*11867*/;
  assign _3537_ = _3536_ & _3535_ /*11866*/;
  assign _3538_ = inv_22[2] & r_21[4] /*11865*/;
  assign _3539_ = _3537_ | _3538_ /*11864*/;
  assign _3540_ = inv_22[3] ^ r_21[5] /*11862*/;
  assign sum_22[3] = _3540_ ^ _3539_ /*11861*/;
  assign _3541_ = _3540_ & _3539_ /*11860*/;
  assign _3542_ = inv_22[3] & r_21[5] /*11859*/;
  assign _3543_ = _3541_ | _3542_ /*11858*/;
  assign _3544_ = inv_22[4] ^ r_21[6] /*11856*/;
  assign sum_22[4] = _3544_ ^ _3543_ /*11855*/;
  assign _3545_ = _3544_ & _3543_ /*11854*/;
  assign _3546_ = inv_22[4] & r_21[6] /*11853*/;
  assign _3547_ = _3545_ | _3546_ /*11852*/;
  assign _3548_ = inv_22[5] ^ r_21[7] /*11850*/;
  assign sum_22[5] = _3548_ ^ _3547_ /*11849*/;
  assign _3549_ = _3548_ & _3547_ /*11848*/;
  assign _3550_ = inv_22[5] & r_21[7] /*11847*/;
  assign _3551_ = _3549_ | _3550_ /*11846*/;
  assign _3552_ = inv_22[6] ^ r_21[8] /*11844*/;
  assign sum_22[6] = _3552_ ^ _3551_ /*11843*/;
  assign _3553_ = _3552_ & _3551_ /*11842*/;
  assign _3554_ = inv_22[6] & r_21[8] /*11841*/;
  assign _3555_ = _3553_ | _3554_ /*11840*/;
  assign _3556_ = inv_22[7] ^ r_21[9] /*11838*/;
  assign sum_22[7] = _3556_ ^ _3555_ /*11837*/;
  assign _3557_ = _3556_ & _3555_ /*11836*/;
  assign _3558_ = inv_22[7] & r_21[9] /*11835*/;
  assign _3559_ = _3557_ | _3558_ /*11834*/;
  assign _3560_ = inv_22[8] ^ r_21[10] /*11832*/;
  assign sum_22[8] = _3560_ ^ _3559_ /*11831*/;
  assign _3561_ = _3560_ & _3559_ /*11830*/;
  assign _3562_ = inv_22[8] & r_21[10] /*11829*/;
  assign _3563_ = _3561_ | _3562_ /*11828*/;
  assign _3564_ = inv_22[9] ^ r_21[11] /*11826*/;
  assign sum_22[9] = _3564_ ^ _3563_ /*11825*/;
  assign _3565_ = _3564_ & _3563_ /*11824*/;
  assign _3566_ = inv_22[9] & r_21[11] /*11823*/;
  assign _3567_ = _3565_ | _3566_ /*11822*/;
  assign _3568_ = inv_22[10] ^ r_21[12] /*11820*/;
  assign sum_22[10] = _3568_ ^ _3567_ /*11819*/;
  assign _3569_ = _3568_ & _3567_ /*11818*/;
  assign _3570_ = inv_22[10] & r_21[12] /*11817*/;
  assign _3571_ = _3569_ | _3570_ /*11816*/;
  assign _3572_ = inv_22[11] ^ r_21[13] /*11814*/;
  assign sum_22[11] = _3572_ ^ _3571_ /*11813*/;
  assign _3573_ = _3572_ & _3571_ /*11812*/;
  assign _3574_ = inv_22[11] & r_21[13] /*11811*/;
  assign _3575_ = _3573_ | _3574_ /*11810*/;
  assign _3576_ = inv_22[12] ^ r_21[14] /*11808*/;
  assign sum_22[12] = _3576_ ^ _3575_ /*11807*/;
  assign _3577_ = _3576_ & _3575_ /*11806*/;
  assign _3578_ = inv_22[12] & r_21[14] /*11805*/;
  assign _3579_ = _3577_ | _3578_ /*11804*/;
  assign _3580_ = inv_22[13] ^ r_21[15] /*11802*/;
  assign sum_22[13] = _3580_ ^ _3579_ /*11801*/;
  assign _3581_ = _3580_ & _3579_ /*11800*/;
  assign _3582_ = inv_22[13] & r_21[15] /*11799*/;
  assign _3583_ = _3581_ | _3582_ /*11798*/;
  assign _3584_ = inv_22[14] ^ r_21[16] /*11796*/;
  assign sum_22[14] = _3584_ ^ _3583_ /*11795*/;
  assign _3585_ = _3584_ & _3583_ /*11794*/;
  assign _3586_ = inv_22[14] & r_21[16] /*11793*/;
  assign _3587_ = _3585_ | _3586_ /*11792*/;
  assign _3588_ = inv_22[15] ^ r_21[17] /*11790*/;
  assign sum_22[15] = _3588_ ^ _3587_ /*11789*/;
  assign _3589_ = _3588_ & _3587_ /*11788*/;
  assign _3590_ = inv_22[15] & r_21[17] /*11787*/;
  assign _3591_ = _3589_ | _3590_ /*11786*/;
  assign _3592_ = inv_22[16] ^ r_21[18] /*11784*/;
  assign sum_22[16] = _3592_ ^ _3591_ /*11783*/;
  assign _3593_ = _3592_ & _3591_ /*11782*/;
  assign _3594_ = inv_22[16] & r_21[18] /*11781*/;
  assign _3595_ = _3593_ | _3594_ /*11780*/;
  assign _3596_ = inv_22[17] ^ r_21[19] /*11778*/;
  assign sum_22[17] = _3596_ ^ _3595_ /*11777*/;
  assign _3597_ = _3596_ & _3595_ /*11776*/;
  assign _3598_ = inv_22[17] & r_21[19] /*11775*/;
  assign _3599_ = _3597_ | _3598_ /*11774*/;
  assign _3600_ = inv_22[18] ^ r_21[20] /*11772*/;
  assign sum_22[18] = _3600_ ^ _3599_ /*11771*/;
  assign _3601_ = _3600_ & _3599_ /*11770*/;
  assign _3602_ = inv_22[18] & r_21[20] /*11769*/;
  assign _3603_ = _3601_ | _3602_ /*11768*/;
  assign _3604_ = inv_22[19] ^ r_21[21] /*11766*/;
  assign sum_22[19] = _3604_ ^ _3603_ /*11765*/;
  assign _3605_ = _3604_ & _3603_ /*11764*/;
  assign _3606_ = inv_22[19] & r_21[21] /*11763*/;
  assign _3607_ = _3605_ | _3606_ /*11762*/;
  assign _3608_ = inv_22[20] ^ r_21[22] /*11760*/;
  assign sum_22[20] = _3608_ ^ _3607_ /*11759*/;
  assign _3609_ = _3608_ & _3607_ /*11758*/;
  assign _3610_ = inv_22[20] & r_21[22] /*11757*/;
  assign _3611_ = _3609_ | _3610_ /*11756*/;
  assign _3612_ = inv_22[21] ^ r_21[23] /*11754*/;
  assign sum_22[21] = _3612_ ^ _3611_ /*11753*/;
  assign _3613_ = _3612_ & _3611_ /*11752*/;
  assign _3614_ = inv_22[21] & r_21[23] /*11751*/;
  assign _3615_ = _3613_ | _3614_ /*11750*/;
  assign _3616_ = inv_22[22] ^ r_21[24] /*11748*/;
  assign sum_22[22] = _3616_ ^ _3615_ /*11747*/;
  assign _3617_ = _3616_ & _3615_ /*11746*/;
  assign _3618_ = inv_22[22] & r_21[24] /*11745*/;
  assign _3619_ = _3617_ | _3618_ /*11744*/;
  assign _3620_ = inv_22[23] ^ r_21[25] /*11742*/;
  assign sum_22[23] = _3620_ ^ _3619_ /*11741*/;
  assign _3621_ = _3620_ & _3619_ /*11740*/;
  assign _3622_ = inv_22[23] & r_21[25] /*11739*/;
  assign _3623_ = _3621_ | _3622_ /*11738*/;
  assign q[2] = ~sum_22[23] /*11757*/;
  assign m_22[0] = r_21[2] /*11756*/;
  assign m_22[1] = r_21[3] /*11755*/;
  assign m_22[2] = r_21[4] /*11754*/;
  assign m_22[3] = r_21[5] /*11753*/;
  assign m_22[4] = r_21[6] /*11752*/;
  assign m_22[5] = r_21[7] /*11751*/;
  assign m_22[6] = r_21[8] /*11750*/;
  assign m_22[7] = r_21[9] /*11749*/;
  assign m_22[8] = r_21[10] /*11748*/;
  assign m_22[9] = r_21[11] /*11747*/;
  assign m_22[10] = r_21[12] /*11746*/;
  assign m_22[11] = r_21[13] /*11745*/;
  assign m_22[12] = r_21[14] /*11744*/;
  assign m_22[13] = r_21[15] /*11743*/;
  assign m_22[14] = r_21[16] /*11742*/;
  assign m_22[15] = r_21[17] /*11741*/;
  assign m_22[16] = r_21[18] /*11740*/;
  assign m_22[17] = r_21[19] /*11739*/;
  assign m_22[18] = r_21[20] /*11738*/;
  assign m_22[19] = r_21[21] /*11737*/;
  assign m_22[20] = r_21[22] /*11736*/;
  assign m_22[21] = r_21[23] /*11735*/;
  assign m_22[22] = r_21[24] /*11734*/;
  assign m_22[23] = r_21[25] /*11733*/;
  assign _3624_ = ~q[2] /*11731*/;
  assign _3625_ = sum_22[0] & q[2] /*11730*/;
  assign _3626_ = m_22[0] & _3624_ /*11729*/;
  assign r_22[2] = _3626_ | _3625_ /*11728*/;
  assign _3627_ = ~q[2] /*11727*/;
  assign _3628_ = sum_22[1] & q[2] /*11726*/;
  assign _3629_ = m_22[1] & _3627_ /*11725*/;
  assign r_22[3] = _3629_ | _3628_ /*11724*/;
  assign _3630_ = ~q[2] /*11723*/;
  assign _3631_ = sum_22[2] & q[2] /*11722*/;
  assign _3632_ = m_22[2] & _3630_ /*11721*/;
  assign r_22[4] = _3632_ | _3631_ /*11720*/;
  assign _3633_ = ~q[2] /*11719*/;
  assign _3634_ = sum_22[3] & q[2] /*11718*/;
  assign _3635_ = m_22[3] & _3633_ /*11717*/;
  assign r_22[5] = _3635_ | _3634_ /*11716*/;
  assign _3636_ = ~q[2] /*11715*/;
  assign _3637_ = sum_22[4] & q[2] /*11714*/;
  assign _3638_ = m_22[4] & _3636_ /*11713*/;
  assign r_22[6] = _3638_ | _3637_ /*11712*/;
  assign _3639_ = ~q[2] /*11711*/;
  assign _3640_ = sum_22[5] & q[2] /*11710*/;
  assign _3641_ = m_22[5] & _3639_ /*11709*/;
  assign r_22[7] = _3641_ | _3640_ /*11708*/;
  assign _3642_ = ~q[2] /*11707*/;
  assign _3643_ = sum_22[6] & q[2] /*11706*/;
  assign _3644_ = m_22[6] & _3642_ /*11705*/;
  assign r_22[8] = _3644_ | _3643_ /*11704*/;
  assign _3645_ = ~q[2] /*11703*/;
  assign _3646_ = sum_22[7] & q[2] /*11702*/;
  assign _3647_ = m_22[7] & _3645_ /*11701*/;
  assign r_22[9] = _3647_ | _3646_ /*11700*/;
  assign _3648_ = ~q[2] /*11699*/;
  assign _3649_ = sum_22[8] & q[2] /*11698*/;
  assign _3650_ = m_22[8] & _3648_ /*11697*/;
  assign r_22[10] = _3650_ | _3649_ /*11696*/;
  assign _3651_ = ~q[2] /*11695*/;
  assign _3652_ = sum_22[9] & q[2] /*11694*/;
  assign _3653_ = m_22[9] & _3651_ /*11693*/;
  assign r_22[11] = _3653_ | _3652_ /*11692*/;
  assign _3654_ = ~q[2] /*11691*/;
  assign _3655_ = sum_22[10] & q[2] /*11690*/;
  assign _3656_ = m_22[10] & _3654_ /*11689*/;
  assign r_22[12] = _3656_ | _3655_ /*11688*/;
  assign _3657_ = ~q[2] /*11687*/;
  assign _3658_ = sum_22[11] & q[2] /*11686*/;
  assign _3659_ = m_22[11] & _3657_ /*11685*/;
  assign r_22[13] = _3659_ | _3658_ /*11684*/;
  assign _3660_ = ~q[2] /*11683*/;
  assign _3661_ = sum_22[12] & q[2] /*11682*/;
  assign _3662_ = m_22[12] & _3660_ /*11681*/;
  assign r_22[14] = _3662_ | _3661_ /*11680*/;
  assign _3663_ = ~q[2] /*11679*/;
  assign _3664_ = sum_22[13] & q[2] /*11678*/;
  assign _3665_ = m_22[13] & _3663_ /*11677*/;
  assign r_22[15] = _3665_ | _3664_ /*11676*/;
  assign _3666_ = ~q[2] /*11675*/;
  assign _3667_ = sum_22[14] & q[2] /*11674*/;
  assign _3668_ = m_22[14] & _3666_ /*11673*/;
  assign r_22[16] = _3668_ | _3667_ /*11672*/;
  assign _3669_ = ~q[2] /*11671*/;
  assign _3670_ = sum_22[15] & q[2] /*11670*/;
  assign _3671_ = m_22[15] & _3669_ /*11669*/;
  assign r_22[17] = _3671_ | _3670_ /*11668*/;
  assign _3672_ = ~q[2] /*11667*/;
  assign _3673_ = sum_22[16] & q[2] /*11666*/;
  assign _3674_ = m_22[16] & _3672_ /*11665*/;
  assign r_22[18] = _3674_ | _3673_ /*11664*/;
  assign _3675_ = ~q[2] /*11663*/;
  assign _3676_ = sum_22[17] & q[2] /*11662*/;
  assign _3677_ = m_22[17] & _3675_ /*11661*/;
  assign r_22[19] = _3677_ | _3676_ /*11660*/;
  assign _3678_ = ~q[2] /*11659*/;
  assign _3679_ = sum_22[18] & q[2] /*11658*/;
  assign _3680_ = m_22[18] & _3678_ /*11657*/;
  assign r_22[20] = _3680_ | _3679_ /*11656*/;
  assign _3681_ = ~q[2] /*11655*/;
  assign _3682_ = sum_22[19] & q[2] /*11654*/;
  assign _3683_ = m_22[19] & _3681_ /*11653*/;
  assign r_22[21] = _3683_ | _3682_ /*11652*/;
  assign _3684_ = ~q[2] /*11651*/;
  assign _3685_ = sum_22[20] & q[2] /*11650*/;
  assign _3686_ = m_22[20] & _3684_ /*11649*/;
  assign r_22[22] = _3686_ | _3685_ /*11648*/;
  assign _3687_ = ~q[2] /*11647*/;
  assign _3688_ = sum_22[21] & q[2] /*11646*/;
  assign _3689_ = m_22[21] & _3687_ /*11645*/;
  assign r_22[23] = _3689_ | _3688_ /*11644*/;
  assign _3690_ = ~q[2] /*11643*/;
  assign _3691_ = sum_22[22] & q[2] /*11642*/;
  assign _3692_ = m_22[22] & _3690_ /*11641*/;
  assign r_22[24] = _3692_ | _3691_ /*11640*/;
  assign _3693_ = ~q[2] /*11639*/;
  assign _3694_ = sum_22[23] & q[2] /*11638*/;
  assign _3695_ = m_22[23] & _3693_ /*11637*/;
  assign r_22[25] = _3695_ | _3694_ /*11636*/;
assign r_22[0]= r_21[0] /*11635*/;
assign r_22[1]= r_21[1] /*11634*/;
  assign inv_23[0] = ~div[0] /*11568*/;
  assign inv_23[1] = ~div[1] /*11567*/;
  assign inv_23[2] = ~div[2] /*11566*/;
  assign inv_23[3] = ~div[3] /*11565*/;
  assign inv_23[4] = ~div[4] /*11564*/;
  assign inv_23[5] = ~div[5] /*11563*/;
  assign inv_23[6] = ~div[6] /*11562*/;
  assign inv_23[7] = ~div[7] /*11561*/;
  assign inv_23[8] = ~div[8] /*11560*/;
  assign inv_23[9] = ~div[9] /*11559*/;
  assign inv_23[10] = ~div[10] /*11558*/;
  assign inv_23[11] = ~div[11] /*11557*/;
  assign inv_23[12] = ~div[12] /*11556*/;
  assign inv_23[13] = ~div[13] /*11555*/;
  assign inv_23[14] = ~div[14] /*11554*/;
  assign inv_23[15] = ~div[15] /*11553*/;
  assign inv_23[16] = ~div[16] /*11552*/;
  assign inv_23[17] = ~div[17] /*11551*/;
  assign inv_23[18] = ~div[18] /*11550*/;
  assign inv_23[19] = ~div[19] /*11549*/;
  assign inv_23[20] = ~div[20] /*11548*/;
  assign inv_23[21] = ~div[21] /*11547*/;
  assign inv_23[22] = ~div[22] /*11546*/;
assign inv_23[23] = oneWire /*11545*/;
  assign _3696_ = inv_23[0] ^ r_22[1] /*11543*/;
  assign sum_23[0] = _3696_ ^ oneWire /*11542*/;
  assign _3697_ = _3696_ & oneWire /*11541*/;
  assign _3698_ = inv_23[0] & r_22[1] /*11540*/;
  assign _3699_ = _3697_ | _3698_ /*11539*/;
  assign _3700_ = inv_23[1] ^ r_22[2] /*11538*/;
  assign sum_23[1] = _3700_ ^ _3699_ /*11537*/;
  assign _3701_ = _3700_ & _3699_ /*11536*/;
  assign _3702_ = inv_23[1] & r_22[2] /*11535*/;
  assign _3703_ = _3701_ | _3702_ /*11534*/;
  assign _3704_ = inv_23[2] ^ r_22[3] /*11532*/;
  assign sum_23[2] = _3704_ ^ _3703_ /*11531*/;
  assign _3705_ = _3704_ & _3703_ /*11530*/;
  assign _3706_ = inv_23[2] & r_22[3] /*11529*/;
  assign _3707_ = _3705_ | _3706_ /*11528*/;
  assign _3708_ = inv_23[3] ^ r_22[4] /*11526*/;
  assign sum_23[3] = _3708_ ^ _3707_ /*11525*/;
  assign _3709_ = _3708_ & _3707_ /*11524*/;
  assign _3710_ = inv_23[3] & r_22[4] /*11523*/;
  assign _3711_ = _3709_ | _3710_ /*11522*/;
  assign _3712_ = inv_23[4] ^ r_22[5] /*11520*/;
  assign sum_23[4] = _3712_ ^ _3711_ /*11519*/;
  assign _3713_ = _3712_ & _3711_ /*11518*/;
  assign _3714_ = inv_23[4] & r_22[5] /*11517*/;
  assign _3715_ = _3713_ | _3714_ /*11516*/;
  assign _3716_ = inv_23[5] ^ r_22[6] /*11514*/;
  assign sum_23[5] = _3716_ ^ _3715_ /*11513*/;
  assign _3717_ = _3716_ & _3715_ /*11512*/;
  assign _3718_ = inv_23[5] & r_22[6] /*11511*/;
  assign _3719_ = _3717_ | _3718_ /*11510*/;
  assign _3720_ = inv_23[6] ^ r_22[7] /*11508*/;
  assign sum_23[6] = _3720_ ^ _3719_ /*11507*/;
  assign _3721_ = _3720_ & _3719_ /*11506*/;
  assign _3722_ = inv_23[6] & r_22[7] /*11505*/;
  assign _3723_ = _3721_ | _3722_ /*11504*/;
  assign _3724_ = inv_23[7] ^ r_22[8] /*11502*/;
  assign sum_23[7] = _3724_ ^ _3723_ /*11501*/;
  assign _3725_ = _3724_ & _3723_ /*11500*/;
  assign _3726_ = inv_23[7] & r_22[8] /*11499*/;
  assign _3727_ = _3725_ | _3726_ /*11498*/;
  assign _3728_ = inv_23[8] ^ r_22[9] /*11496*/;
  assign sum_23[8] = _3728_ ^ _3727_ /*11495*/;
  assign _3729_ = _3728_ & _3727_ /*11494*/;
  assign _3730_ = inv_23[8] & r_22[9] /*11493*/;
  assign _3731_ = _3729_ | _3730_ /*11492*/;
  assign _3732_ = inv_23[9] ^ r_22[10] /*11490*/;
  assign sum_23[9] = _3732_ ^ _3731_ /*11489*/;
  assign _3733_ = _3732_ & _3731_ /*11488*/;
  assign _3734_ = inv_23[9] & r_22[10] /*11487*/;
  assign _3735_ = _3733_ | _3734_ /*11486*/;
  assign _3736_ = inv_23[10] ^ r_22[11] /*11484*/;
  assign sum_23[10] = _3736_ ^ _3735_ /*11483*/;
  assign _3737_ = _3736_ & _3735_ /*11482*/;
  assign _3738_ = inv_23[10] & r_22[11] /*11481*/;
  assign _3739_ = _3737_ | _3738_ /*11480*/;
  assign _3740_ = inv_23[11] ^ r_22[12] /*11478*/;
  assign sum_23[11] = _3740_ ^ _3739_ /*11477*/;
  assign _3741_ = _3740_ & _3739_ /*11476*/;
  assign _3742_ = inv_23[11] & r_22[12] /*11475*/;
  assign _3743_ = _3741_ | _3742_ /*11474*/;
  assign _3744_ = inv_23[12] ^ r_22[13] /*11472*/;
  assign sum_23[12] = _3744_ ^ _3743_ /*11471*/;
  assign _3745_ = _3744_ & _3743_ /*11470*/;
  assign _3746_ = inv_23[12] & r_22[13] /*11469*/;
  assign _3747_ = _3745_ | _3746_ /*11468*/;
  assign _3748_ = inv_23[13] ^ r_22[14] /*11466*/;
  assign sum_23[13] = _3748_ ^ _3747_ /*11465*/;
  assign _3749_ = _3748_ & _3747_ /*11464*/;
  assign _3750_ = inv_23[13] & r_22[14] /*11463*/;
  assign _3751_ = _3749_ | _3750_ /*11462*/;
  assign _3752_ = inv_23[14] ^ r_22[15] /*11460*/;
  assign sum_23[14] = _3752_ ^ _3751_ /*11459*/;
  assign _3753_ = _3752_ & _3751_ /*11458*/;
  assign _3754_ = inv_23[14] & r_22[15] /*11457*/;
  assign _3755_ = _3753_ | _3754_ /*11456*/;
  assign _3756_ = inv_23[15] ^ r_22[16] /*11454*/;
  assign sum_23[15] = _3756_ ^ _3755_ /*11453*/;
  assign _3757_ = _3756_ & _3755_ /*11452*/;
  assign _3758_ = inv_23[15] & r_22[16] /*11451*/;
  assign _3759_ = _3757_ | _3758_ /*11450*/;
  assign _3760_ = inv_23[16] ^ r_22[17] /*11448*/;
  assign sum_23[16] = _3760_ ^ _3759_ /*11447*/;
  assign _3761_ = _3760_ & _3759_ /*11446*/;
  assign _3762_ = inv_23[16] & r_22[17] /*11445*/;
  assign _3763_ = _3761_ | _3762_ /*11444*/;
  assign _3764_ = inv_23[17] ^ r_22[18] /*11442*/;
  assign sum_23[17] = _3764_ ^ _3763_ /*11441*/;
  assign _3765_ = _3764_ & _3763_ /*11440*/;
  assign _3766_ = inv_23[17] & r_22[18] /*11439*/;
  assign _3767_ = _3765_ | _3766_ /*11438*/;
  assign _3768_ = inv_23[18] ^ r_22[19] /*11436*/;
  assign sum_23[18] = _3768_ ^ _3767_ /*11435*/;
  assign _3769_ = _3768_ & _3767_ /*11434*/;
  assign _3770_ = inv_23[18] & r_22[19] /*11433*/;
  assign _3771_ = _3769_ | _3770_ /*11432*/;
  assign _3772_ = inv_23[19] ^ r_22[20] /*11430*/;
  assign sum_23[19] = _3772_ ^ _3771_ /*11429*/;
  assign _3773_ = _3772_ & _3771_ /*11428*/;
  assign _3774_ = inv_23[19] & r_22[20] /*11427*/;
  assign _3775_ = _3773_ | _3774_ /*11426*/;
  assign _3776_ = inv_23[20] ^ r_22[21] /*11424*/;
  assign sum_23[20] = _3776_ ^ _3775_ /*11423*/;
  assign _3777_ = _3776_ & _3775_ /*11422*/;
  assign _3778_ = inv_23[20] & r_22[21] /*11421*/;
  assign _3779_ = _3777_ | _3778_ /*11420*/;
  assign _3780_ = inv_23[21] ^ r_22[22] /*11418*/;
  assign sum_23[21] = _3780_ ^ _3779_ /*11417*/;
  assign _3781_ = _3780_ & _3779_ /*11416*/;
  assign _3782_ = inv_23[21] & r_22[22] /*11415*/;
  assign _3783_ = _3781_ | _3782_ /*11414*/;
  assign _3784_ = inv_23[22] ^ r_22[23] /*11412*/;
  assign sum_23[22] = _3784_ ^ _3783_ /*11411*/;
  assign _3785_ = _3784_ & _3783_ /*11410*/;
  assign _3786_ = inv_23[22] & r_22[23] /*11409*/;
  assign _3787_ = _3785_ | _3786_ /*11408*/;
  assign _3788_ = inv_23[23] ^ r_22[24] /*11406*/;
  assign sum_23[23] = _3788_ ^ _3787_ /*11405*/;
  assign _3789_ = _3788_ & _3787_ /*11404*/;
  assign _3790_ = inv_23[23] & r_22[24] /*11403*/;
  assign _3791_ = _3789_ | _3790_ /*11402*/;
  assign q[1] = ~sum_23[23] /*11421*/;
  assign m_23[0] = r_22[1] /*11420*/;
  assign m_23[1] = r_22[2] /*11419*/;
  assign m_23[2] = r_22[3] /*11418*/;
  assign m_23[3] = r_22[4] /*11417*/;
  assign m_23[4] = r_22[5] /*11416*/;
  assign m_23[5] = r_22[6] /*11415*/;
  assign m_23[6] = r_22[7] /*11414*/;
  assign m_23[7] = r_22[8] /*11413*/;
  assign m_23[8] = r_22[9] /*11412*/;
  assign m_23[9] = r_22[10] /*11411*/;
  assign m_23[10] = r_22[11] /*11410*/;
  assign m_23[11] = r_22[12] /*11409*/;
  assign m_23[12] = r_22[13] /*11408*/;
  assign m_23[13] = r_22[14] /*11407*/;
  assign m_23[14] = r_22[15] /*11406*/;
  assign m_23[15] = r_22[16] /*11405*/;
  assign m_23[16] = r_22[17] /*11404*/;
  assign m_23[17] = r_22[18] /*11403*/;
  assign m_23[18] = r_22[19] /*11402*/;
  assign m_23[19] = r_22[20] /*11401*/;
  assign m_23[20] = r_22[21] /*11400*/;
  assign m_23[21] = r_22[22] /*11399*/;
  assign m_23[22] = r_22[23] /*11398*/;
  assign m_23[23] = r_22[24] /*11397*/;
  assign _3792_ = ~q[1] /*11395*/;
  assign _3793_ = sum_23[0] & q[1] /*11394*/;
  assign _3794_ = m_23[0] & _3792_ /*11393*/;
  assign r_23[1] = _3794_ | _3793_ /*11392*/;
  assign _3795_ = ~q[1] /*11391*/;
  assign _3796_ = sum_23[1] & q[1] /*11390*/;
  assign _3797_ = m_23[1] & _3795_ /*11389*/;
  assign r_23[2] = _3797_ | _3796_ /*11388*/;
  assign _3798_ = ~q[1] /*11387*/;
  assign _3799_ = sum_23[2] & q[1] /*11386*/;
  assign _3800_ = m_23[2] & _3798_ /*11385*/;
  assign r_23[3] = _3800_ | _3799_ /*11384*/;
  assign _3801_ = ~q[1] /*11383*/;
  assign _3802_ = sum_23[3] & q[1] /*11382*/;
  assign _3803_ = m_23[3] & _3801_ /*11381*/;
  assign r_23[4] = _3803_ | _3802_ /*11380*/;
  assign _3804_ = ~q[1] /*11379*/;
  assign _3805_ = sum_23[4] & q[1] /*11378*/;
  assign _3806_ = m_23[4] & _3804_ /*11377*/;
  assign r_23[5] = _3806_ | _3805_ /*11376*/;
  assign _3807_ = ~q[1] /*11375*/;
  assign _3808_ = sum_23[5] & q[1] /*11374*/;
  assign _3809_ = m_23[5] & _3807_ /*11373*/;
  assign r_23[6] = _3809_ | _3808_ /*11372*/;
  assign _3810_ = ~q[1] /*11371*/;
  assign _3811_ = sum_23[6] & q[1] /*11370*/;
  assign _3812_ = m_23[6] & _3810_ /*11369*/;
  assign r_23[7] = _3812_ | _3811_ /*11368*/;
  assign _3813_ = ~q[1] /*11367*/;
  assign _3814_ = sum_23[7] & q[1] /*11366*/;
  assign _3815_ = m_23[7] & _3813_ /*11365*/;
  assign r_23[8] = _3815_ | _3814_ /*11364*/;
  assign _3816_ = ~q[1] /*11363*/;
  assign _3817_ = sum_23[8] & q[1] /*11362*/;
  assign _3818_ = m_23[8] & _3816_ /*11361*/;
  assign r_23[9] = _3818_ | _3817_ /*11360*/;
  assign _3819_ = ~q[1] /*11359*/;
  assign _3820_ = sum_23[9] & q[1] /*11358*/;
  assign _3821_ = m_23[9] & _3819_ /*11357*/;
  assign r_23[10] = _3821_ | _3820_ /*11356*/;
  assign _3822_ = ~q[1] /*11355*/;
  assign _3823_ = sum_23[10] & q[1] /*11354*/;
  assign _3824_ = m_23[10] & _3822_ /*11353*/;
  assign r_23[11] = _3824_ | _3823_ /*11352*/;
  assign _3825_ = ~q[1] /*11351*/;
  assign _3826_ = sum_23[11] & q[1] /*11350*/;
  assign _3827_ = m_23[11] & _3825_ /*11349*/;
  assign r_23[12] = _3827_ | _3826_ /*11348*/;
  assign _3828_ = ~q[1] /*11347*/;
  assign _3829_ = sum_23[12] & q[1] /*11346*/;
  assign _3830_ = m_23[12] & _3828_ /*11345*/;
  assign r_23[13] = _3830_ | _3829_ /*11344*/;
  assign _3831_ = ~q[1] /*11343*/;
  assign _3832_ = sum_23[13] & q[1] /*11342*/;
  assign _3833_ = m_23[13] & _3831_ /*11341*/;
  assign r_23[14] = _3833_ | _3832_ /*11340*/;
  assign _3834_ = ~q[1] /*11339*/;
  assign _3835_ = sum_23[14] & q[1] /*11338*/;
  assign _3836_ = m_23[14] & _3834_ /*11337*/;
  assign r_23[15] = _3836_ | _3835_ /*11336*/;
  assign _3837_ = ~q[1] /*11335*/;
  assign _3838_ = sum_23[15] & q[1] /*11334*/;
  assign _3839_ = m_23[15] & _3837_ /*11333*/;
  assign r_23[16] = _3839_ | _3838_ /*11332*/;
  assign _3840_ = ~q[1] /*11331*/;
  assign _3841_ = sum_23[16] & q[1] /*11330*/;
  assign _3842_ = m_23[16] & _3840_ /*11329*/;
  assign r_23[17] = _3842_ | _3841_ /*11328*/;
  assign _3843_ = ~q[1] /*11327*/;
  assign _3844_ = sum_23[17] & q[1] /*11326*/;
  assign _3845_ = m_23[17] & _3843_ /*11325*/;
  assign r_23[18] = _3845_ | _3844_ /*11324*/;
  assign _3846_ = ~q[1] /*11323*/;
  assign _3847_ = sum_23[18] & q[1] /*11322*/;
  assign _3848_ = m_23[18] & _3846_ /*11321*/;
  assign r_23[19] = _3848_ | _3847_ /*11320*/;
  assign _3849_ = ~q[1] /*11319*/;
  assign _3850_ = sum_23[19] & q[1] /*11318*/;
  assign _3851_ = m_23[19] & _3849_ /*11317*/;
  assign r_23[20] = _3851_ | _3850_ /*11316*/;
  assign _3852_ = ~q[1] /*11315*/;
  assign _3853_ = sum_23[20] & q[1] /*11314*/;
  assign _3854_ = m_23[20] & _3852_ /*11313*/;
  assign r_23[21] = _3854_ | _3853_ /*11312*/;
  assign _3855_ = ~q[1] /*11311*/;
  assign _3856_ = sum_23[21] & q[1] /*11310*/;
  assign _3857_ = m_23[21] & _3855_ /*11309*/;
  assign r_23[22] = _3857_ | _3856_ /*11308*/;
  assign _3858_ = ~q[1] /*11307*/;
  assign _3859_ = sum_23[22] & q[1] /*11306*/;
  assign _3860_ = m_23[22] & _3858_ /*11305*/;
  assign r_23[23] = _3860_ | _3859_ /*11304*/;
  assign _3861_ = ~q[1] /*11303*/;
  assign _3862_ = sum_23[23] & q[1] /*11302*/;
  assign _3863_ = m_23[23] & _3861_ /*11301*/;
  assign r_23[24] = _3863_ | _3862_ /*11300*/;
assign r_23[0]= r_22[0] /*11299*/;
  assign inv_24[0] = ~div[0] /*11232*/;
  assign inv_24[1] = ~div[1] /*11231*/;
  assign inv_24[2] = ~div[2] /*11230*/;
  assign inv_24[3] = ~div[3] /*11229*/;
  assign inv_24[4] = ~div[4] /*11228*/;
  assign inv_24[5] = ~div[5] /*11227*/;
  assign inv_24[6] = ~div[6] /*11226*/;
  assign inv_24[7] = ~div[7] /*11225*/;
  assign inv_24[8] = ~div[8] /*11224*/;
  assign inv_24[9] = ~div[9] /*11223*/;
  assign inv_24[10] = ~div[10] /*11222*/;
  assign inv_24[11] = ~div[11] /*11221*/;
  assign inv_24[12] = ~div[12] /*11220*/;
  assign inv_24[13] = ~div[13] /*11219*/;
  assign inv_24[14] = ~div[14] /*11218*/;
  assign inv_24[15] = ~div[15] /*11217*/;
  assign inv_24[16] = ~div[16] /*11216*/;
  assign inv_24[17] = ~div[17] /*11215*/;
  assign inv_24[18] = ~div[18] /*11214*/;
  assign inv_24[19] = ~div[19] /*11213*/;
  assign inv_24[20] = ~div[20] /*11212*/;
  assign inv_24[21] = ~div[21] /*11211*/;
  assign inv_24[22] = ~div[22] /*11210*/;
assign inv_24[23] = oneWire /*11209*/;
  assign _3864_ = inv_24[0] ^ r_23[0] /*11207*/;
  assign sum_24[0] = _3864_ ^ oneWire /*11206*/;
  assign _3865_ = _3864_ & oneWire /*11205*/;
  assign _3866_ = inv_24[0] & r_23[0] /*11204*/;
  assign _3867_ = _3865_ | _3866_ /*11203*/;
  assign _3868_ = inv_24[1] ^ r_23[1] /*11202*/;
  assign sum_24[1] = _3868_ ^ _3867_ /*11201*/;
  assign _3869_ = _3868_ & _3867_ /*11200*/;
  assign _3870_ = inv_24[1] & r_23[1] /*11199*/;
  assign _3871_ = _3869_ | _3870_ /*11198*/;
  assign _3872_ = inv_24[2] ^ r_23[2] /*11196*/;
  assign sum_24[2] = _3872_ ^ _3871_ /*11195*/;
  assign _3873_ = _3872_ & _3871_ /*11194*/;
  assign _3874_ = inv_24[2] & r_23[2] /*11193*/;
  assign _3875_ = _3873_ | _3874_ /*11192*/;
  assign _3876_ = inv_24[3] ^ r_23[3] /*11190*/;
  assign sum_24[3] = _3876_ ^ _3875_ /*11189*/;
  assign _3877_ = _3876_ & _3875_ /*11188*/;
  assign _3878_ = inv_24[3] & r_23[3] /*11187*/;
  assign _3879_ = _3877_ | _3878_ /*11186*/;
  assign _3880_ = inv_24[4] ^ r_23[4] /*11184*/;
  assign sum_24[4] = _3880_ ^ _3879_ /*11183*/;
  assign _3881_ = _3880_ & _3879_ /*11182*/;
  assign _3882_ = inv_24[4] & r_23[4] /*11181*/;
  assign _3883_ = _3881_ | _3882_ /*11180*/;
  assign _3884_ = inv_24[5] ^ r_23[5] /*11178*/;
  assign sum_24[5] = _3884_ ^ _3883_ /*11177*/;
  assign _3885_ = _3884_ & _3883_ /*11176*/;
  assign _3886_ = inv_24[5] & r_23[5] /*11175*/;
  assign _3887_ = _3885_ | _3886_ /*11174*/;
  assign _3888_ = inv_24[6] ^ r_23[6] /*11172*/;
  assign sum_24[6] = _3888_ ^ _3887_ /*11171*/;
  assign _3889_ = _3888_ & _3887_ /*11170*/;
  assign _3890_ = inv_24[6] & r_23[6] /*11169*/;
  assign _3891_ = _3889_ | _3890_ /*11168*/;
  assign _3892_ = inv_24[7] ^ r_23[7] /*11166*/;
  assign sum_24[7] = _3892_ ^ _3891_ /*11165*/;
  assign _3893_ = _3892_ & _3891_ /*11164*/;
  assign _3894_ = inv_24[7] & r_23[7] /*11163*/;
  assign _3895_ = _3893_ | _3894_ /*11162*/;
  assign _3896_ = inv_24[8] ^ r_23[8] /*11160*/;
  assign sum_24[8] = _3896_ ^ _3895_ /*11159*/;
  assign _3897_ = _3896_ & _3895_ /*11158*/;
  assign _3898_ = inv_24[8] & r_23[8] /*11157*/;
  assign _3899_ = _3897_ | _3898_ /*11156*/;
  assign _3900_ = inv_24[9] ^ r_23[9] /*11154*/;
  assign sum_24[9] = _3900_ ^ _3899_ /*11153*/;
  assign _3901_ = _3900_ & _3899_ /*11152*/;
  assign _3902_ = inv_24[9] & r_23[9] /*11151*/;
  assign _3903_ = _3901_ | _3902_ /*11150*/;
  assign _3904_ = inv_24[10] ^ r_23[10] /*11148*/;
  assign sum_24[10] = _3904_ ^ _3903_ /*11147*/;
  assign _3905_ = _3904_ & _3903_ /*11146*/;
  assign _3906_ = inv_24[10] & r_23[10] /*11145*/;
  assign _3907_ = _3905_ | _3906_ /*11144*/;
  assign _3908_ = inv_24[11] ^ r_23[11] /*11142*/;
  assign sum_24[11] = _3908_ ^ _3907_ /*11141*/;
  assign _3909_ = _3908_ & _3907_ /*11140*/;
  assign _3910_ = inv_24[11] & r_23[11] /*11139*/;
  assign _3911_ = _3909_ | _3910_ /*11138*/;
  assign _3912_ = inv_24[12] ^ r_23[12] /*11136*/;
  assign sum_24[12] = _3912_ ^ _3911_ /*11135*/;
  assign _3913_ = _3912_ & _3911_ /*11134*/;
  assign _3914_ = inv_24[12] & r_23[12] /*11133*/;
  assign _3915_ = _3913_ | _3914_ /*11132*/;
  assign _3916_ = inv_24[13] ^ r_23[13] /*11130*/;
  assign sum_24[13] = _3916_ ^ _3915_ /*11129*/;
  assign _3917_ = _3916_ & _3915_ /*11128*/;
  assign _3918_ = inv_24[13] & r_23[13] /*11127*/;
  assign _3919_ = _3917_ | _3918_ /*11126*/;
  assign _3920_ = inv_24[14] ^ r_23[14] /*11124*/;
  assign sum_24[14] = _3920_ ^ _3919_ /*11123*/;
  assign _3921_ = _3920_ & _3919_ /*11122*/;
  assign _3922_ = inv_24[14] & r_23[14] /*11121*/;
  assign _3923_ = _3921_ | _3922_ /*11120*/;
  assign _3924_ = inv_24[15] ^ r_23[15] /*11118*/;
  assign sum_24[15] = _3924_ ^ _3923_ /*11117*/;
  assign _3925_ = _3924_ & _3923_ /*11116*/;
  assign _3926_ = inv_24[15] & r_23[15] /*11115*/;
  assign _3927_ = _3925_ | _3926_ /*11114*/;
  assign _3928_ = inv_24[16] ^ r_23[16] /*11112*/;
  assign sum_24[16] = _3928_ ^ _3927_ /*11111*/;
  assign _3929_ = _3928_ & _3927_ /*11110*/;
  assign _3930_ = inv_24[16] & r_23[16] /*11109*/;
  assign _3931_ = _3929_ | _3930_ /*11108*/;
  assign _3932_ = inv_24[17] ^ r_23[17] /*11106*/;
  assign sum_24[17] = _3932_ ^ _3931_ /*11105*/;
  assign _3933_ = _3932_ & _3931_ /*11104*/;
  assign _3934_ = inv_24[17] & r_23[17] /*11103*/;
  assign _3935_ = _3933_ | _3934_ /*11102*/;
  assign _3936_ = inv_24[18] ^ r_23[18] /*11100*/;
  assign sum_24[18] = _3936_ ^ _3935_ /*11099*/;
  assign _3937_ = _3936_ & _3935_ /*11098*/;
  assign _3938_ = inv_24[18] & r_23[18] /*11097*/;
  assign _3939_ = _3937_ | _3938_ /*11096*/;
  assign _3940_ = inv_24[19] ^ r_23[19] /*11094*/;
  assign sum_24[19] = _3940_ ^ _3939_ /*11093*/;
  assign _3941_ = _3940_ & _3939_ /*11092*/;
  assign _3942_ = inv_24[19] & r_23[19] /*11091*/;
  assign _3943_ = _3941_ | _3942_ /*11090*/;
  assign _3944_ = inv_24[20] ^ r_23[20] /*11088*/;
  assign sum_24[20] = _3944_ ^ _3943_ /*11087*/;
  assign _3945_ = _3944_ & _3943_ /*11086*/;
  assign _3946_ = inv_24[20] & r_23[20] /*11085*/;
  assign _3947_ = _3945_ | _3946_ /*11084*/;
  assign _3948_ = inv_24[21] ^ r_23[21] /*11082*/;
  assign sum_24[21] = _3948_ ^ _3947_ /*11081*/;
  assign _3949_ = _3948_ & _3947_ /*11080*/;
  assign _3950_ = inv_24[21] & r_23[21] /*11079*/;
  assign _3951_ = _3949_ | _3950_ /*11078*/;
  assign _3952_ = inv_24[22] ^ r_23[22] /*11076*/;
  assign sum_24[22] = _3952_ ^ _3951_ /*11075*/;
  assign _3953_ = _3952_ & _3951_ /*11074*/;
  assign _3954_ = inv_24[22] & r_23[22] /*11073*/;
  assign _3955_ = _3953_ | _3954_ /*11072*/;
  assign _3956_ = inv_24[23] ^ r_23[23] /*11070*/;
  assign sum_24[23] = _3956_ ^ _3955_ /*11069*/;
  assign _3957_ = _3956_ & _3955_ /*11068*/;
  assign _3958_ = inv_24[23] & r_23[23] /*11067*/;
  assign _3959_ = _3957_ | _3958_ /*11066*/;
  assign q[0] = ~sum_24[23] /*11085*/;
  assign m_24[0] = r_23[0] /*11084*/;
  assign m_24[1] = r_23[1] /*11083*/;
  assign m_24[2] = r_23[2] /*11082*/;
  assign m_24[3] = r_23[3] /*11081*/;
  assign m_24[4] = r_23[4] /*11080*/;
  assign m_24[5] = r_23[5] /*11079*/;
  assign m_24[6] = r_23[6] /*11078*/;
  assign m_24[7] = r_23[7] /*11077*/;
  assign m_24[8] = r_23[8] /*11076*/;
  assign m_24[9] = r_23[9] /*11075*/;
  assign m_24[10] = r_23[10] /*11074*/;
  assign m_24[11] = r_23[11] /*11073*/;
  assign m_24[12] = r_23[12] /*11072*/;
  assign m_24[13] = r_23[13] /*11071*/;
  assign m_24[14] = r_23[14] /*11070*/;
  assign m_24[15] = r_23[15] /*11069*/;
  assign m_24[16] = r_23[16] /*11068*/;
  assign m_24[17] = r_23[17] /*11067*/;
  assign m_24[18] = r_23[18] /*11066*/;
  assign m_24[19] = r_23[19] /*11065*/;
  assign m_24[20] = r_23[20] /*11064*/;
  assign m_24[21] = r_23[21] /*11063*/;
  assign m_24[22] = r_23[22] /*11062*/;
  assign m_24[23] = r_23[23] /*11061*/;
  assign _3960_ = ~q[0] /*11059*/;
  assign _3961_ = sum_24[0] & q[0] /*11058*/;
  assign _3962_ = m_24[0] & _3960_ /*11057*/;
  assign r_24[0] = _3962_ | _3961_ /*11056*/;
  assign _3963_ = ~q[0] /*11055*/;
  assign _3964_ = sum_24[1] & q[0] /*11054*/;
  assign _3965_ = m_24[1] & _3963_ /*11053*/;
  assign r_24[1] = _3965_ | _3964_ /*11052*/;
  assign _3966_ = ~q[0] /*11051*/;
  assign _3967_ = sum_24[2] & q[0] /*11050*/;
  assign _3968_ = m_24[2] & _3966_ /*11049*/;
  assign r_24[2] = _3968_ | _3967_ /*11048*/;
  assign _3969_ = ~q[0] /*11047*/;
  assign _3970_ = sum_24[3] & q[0] /*11046*/;
  assign _3971_ = m_24[3] & _3969_ /*11045*/;
  assign r_24[3] = _3971_ | _3970_ /*11044*/;
  assign _3972_ = ~q[0] /*11043*/;
  assign _3973_ = sum_24[4] & q[0] /*11042*/;
  assign _3974_ = m_24[4] & _3972_ /*11041*/;
  assign r_24[4] = _3974_ | _3973_ /*11040*/;
  assign _3975_ = ~q[0] /*11039*/;
  assign _3976_ = sum_24[5] & q[0] /*11038*/;
  assign _3977_ = m_24[5] & _3975_ /*11037*/;
  assign r_24[5] = _3977_ | _3976_ /*11036*/;
  assign _3978_ = ~q[0] /*11035*/;
  assign _3979_ = sum_24[6] & q[0] /*11034*/;
  assign _3980_ = m_24[6] & _3978_ /*11033*/;
  assign r_24[6] = _3980_ | _3979_ /*11032*/;
  assign _3981_ = ~q[0] /*11031*/;
  assign _3982_ = sum_24[7] & q[0] /*11030*/;
  assign _3983_ = m_24[7] & _3981_ /*11029*/;
  assign r_24[7] = _3983_ | _3982_ /*11028*/;
  assign _3984_ = ~q[0] /*11027*/;
  assign _3985_ = sum_24[8] & q[0] /*11026*/;
  assign _3986_ = m_24[8] & _3984_ /*11025*/;
  assign r_24[8] = _3986_ | _3985_ /*11024*/;
  assign _3987_ = ~q[0] /*11023*/;
  assign _3988_ = sum_24[9] & q[0] /*11022*/;
  assign _3989_ = m_24[9] & _3987_ /*11021*/;
  assign r_24[9] = _3989_ | _3988_ /*11020*/;
  assign _3990_ = ~q[0] /*11019*/;
  assign _3991_ = sum_24[10] & q[0] /*11018*/;
  assign _3992_ = m_24[10] & _3990_ /*11017*/;
  assign r_24[10] = _3992_ | _3991_ /*11016*/;
  assign _3993_ = ~q[0] /*11015*/;
  assign _3994_ = sum_24[11] & q[0] /*11014*/;
  assign _3995_ = m_24[11] & _3993_ /*11013*/;
  assign r_24[11] = _3995_ | _3994_ /*11012*/;
  assign _3996_ = ~q[0] /*11011*/;
  assign _3997_ = sum_24[12] & q[0] /*11010*/;
  assign _3998_ = m_24[12] & _3996_ /*11009*/;
  assign r_24[12] = _3998_ | _3997_ /*11008*/;
  assign _3999_ = ~q[0] /*11007*/;
  assign _4000_ = sum_24[13] & q[0] /*11006*/;
  assign _4001_ = m_24[13] & _3999_ /*11005*/;
  assign r_24[13] = _4001_ | _4000_ /*11004*/;
  assign _4002_ = ~q[0] /*11003*/;
  assign _4003_ = sum_24[14] & q[0] /*11002*/;
  assign _4004_ = m_24[14] & _4002_ /*11001*/;
  assign r_24[14] = _4004_ | _4003_ /*11000*/;
  assign _4005_ = ~q[0] /*10999*/;
  assign _4006_ = sum_24[15] & q[0] /*10998*/;
  assign _4007_ = m_24[15] & _4005_ /*10997*/;
  assign r_24[15] = _4007_ | _4006_ /*10996*/;
  assign _4008_ = ~q[0] /*10995*/;
  assign _4009_ = sum_24[16] & q[0] /*10994*/;
  assign _4010_ = m_24[16] & _4008_ /*10993*/;
  assign r_24[16] = _4010_ | _4009_ /*10992*/;
  assign _4011_ = ~q[0] /*10991*/;
  assign _4012_ = sum_24[17] & q[0] /*10990*/;
  assign _4013_ = m_24[17] & _4011_ /*10989*/;
  assign r_24[17] = _4013_ | _4012_ /*10988*/;
  assign _4014_ = ~q[0] /*10987*/;
  assign _4015_ = sum_24[18] & q[0] /*10986*/;
  assign _4016_ = m_24[18] & _4014_ /*10985*/;
  assign r_24[18] = _4016_ | _4015_ /*10984*/;
  assign _4017_ = ~q[0] /*10983*/;
  assign _4018_ = sum_24[19] & q[0] /*10982*/;
  assign _4019_ = m_24[19] & _4017_ /*10981*/;
  assign r_24[19] = _4019_ | _4018_ /*10980*/;
  assign _4020_ = ~q[0] /*10979*/;
  assign _4021_ = sum_24[20] & q[0] /*10978*/;
  assign _4022_ = m_24[20] & _4020_ /*10977*/;
  assign r_24[20] = _4022_ | _4021_ /*10976*/;
  assign _4023_ = ~q[0] /*10975*/;
  assign _4024_ = sum_24[21] & q[0] /*10974*/;
  assign _4025_ = m_24[21] & _4023_ /*10973*/;
  assign r_24[21] = _4025_ | _4024_ /*10972*/;
  assign _4026_ = ~q[0] /*10971*/;
  assign _4027_ = sum_24[22] & q[0] /*10970*/;
  assign _4028_ = m_24[22] & _4026_ /*10969*/;
  assign r_24[22] = _4028_ | _4027_ /*10968*/;
  assign _4029_ = ~q[0] /*10967*/;
  assign _4030_ = sum_24[23] & q[0] /*10966*/;
  assign _4031_ = m_24[23] & _4029_ /*10965*/;
  assign r_24[23] = _4031_ | _4030_ /*10964*/;
  assign rout[0] = r_24[0] /*0*/;
  assign rout[1] = r_24[1] /*1*/;
  assign rout[2] = r_24[2] /*2*/;
  assign rout[3] = r_24[3] /*3*/;
  assign rout[4] = r_24[4] /*4*/;
  assign rout[5] = r_24[5] /*5*/;
  assign rout[6] = r_24[6] /*6*/;
  assign rout[7] = r_24[7] /*7*/;
  assign rout[8] = r_24[8] /*8*/;
  assign rout[9] = r_24[9] /*9*/;
  assign rout[10] = r_24[10] /*10*/;
  assign rout[11] = r_24[11] /*11*/;
  assign rout[12] = r_24[12] /*12*/;
  assign rout[13] = r_24[13] /*13*/;
  assign rout[14] = r_24[14] /*14*/;
  assign rout[15] = r_24[15] /*15*/;
  assign rout[16] = r_24[16] /*16*/;
  assign rout[17] = r_24[17] /*17*/;
  assign rout[18] = r_24[18] /*18*/;
  assign rout[19] = r_24[19] /*19*/;
  assign rout[20] = r_24[20] /*20*/;
  assign rout[21] = r_24[21] /*21*/;
  assign rout[22] = r_24[22] /*22*/;
  assign rout[23] = r_24[23] /*23*/;
endmodule