module divider(R_0, D, Q, R_n1);
input [61:0] R_0;
input [30:0] D;
output [31:0] Q;
output [30:0] R_n1;
wire _0_;
wire _1_;
wire _2_;
wire _3_;
wire _4_;
wire _5_;
wire _6_;
wire _7_;
wire _8_;
wire _9_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
wire _29_;
wire _30_;
wire _31_;
wire _32_;
wire _33_;
wire _34_;
wire _35_;
wire _36_;
wire _37_;
wire _38_;
wire _39_;
wire _40_;
wire _41_;
wire _42_;
wire _43_;
wire _44_;
wire _45_;
wire _46_;
wire _47_;
wire _48_;
wire _49_;
wire _50_;
wire _51_;
wire _52_;
wire _53_;
wire _54_;
wire _55_;
wire _56_;
wire _57_;
wire _58_;
wire _59_;
wire _60_;
wire _61_;
wire _62_;
wire _63_;
wire _64_;
wire _65_;
wire _66_;
wire _67_;
wire _68_;
wire _69_;
wire _70_;
wire _71_;
wire _72_;
wire _73_;
wire _74_;
wire _75_;
wire _76_;
wire _77_;
wire _78_;
wire _79_;
wire _80_;
wire _81_;
wire _82_;
wire _83_;
wire _84_;
wire _85_;
wire _86_;
wire _87_;
wire _88_;
wire _89_;
wire _90_;
wire _91_;
wire _92_;
wire _93_;
wire _94_;
wire _95_;
wire _96_;
wire _97_;
wire _98_;
wire _99_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
wire _255_;
wire _256_;
wire _257_;
wire _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire _267_;
wire _268_;
wire _269_;
wire _270_;
wire _271_;
wire _272_;
wire _273_;
wire _274_;
wire _275_;
wire _276_;
wire _277_;
wire _278_;
wire _279_;
wire _280_;
wire _281_;
wire _282_;
wire _283_;
wire _284_;
wire _285_;
wire _286_;
wire _287_;
wire _288_;
wire _289_;
wire _290_;
wire _291_;
wire _292_;
wire _293_;
wire _294_;
wire _295_;
wire _296_;
wire _297_;
wire _298_;
wire _299_;
wire _300_;
wire _301_;
wire _302_;
wire _303_;
wire _304_;
wire _305_;
wire _306_;
wire _307_;
wire _308_;
wire _309_;
wire _310_;
wire _311_;
wire _312_;
wire _313_;
wire _314_;
wire _315_;
wire _316_;
wire _317_;
wire _318_;
wire _319_;
wire _320_;
wire _321_;
wire _322_;
wire _323_;
wire _324_;
wire _325_;
wire _326_;
wire _327_;
wire _328_;
wire _329_;
wire _330_;
wire _331_;
wire _332_;
wire _333_;
wire _334_;
wire _335_;
wire _336_;
wire _337_;
wire _338_;
wire _339_;
wire _340_;
wire _341_;
wire _342_;
wire _343_;
wire _344_;
wire _345_;
wire _346_;
wire _347_;
wire _348_;
wire _349_;
wire _350_;
wire _351_;
wire _352_;
wire _353_;
wire _354_;
wire _355_;
wire _356_;
wire _357_;
wire _358_;
wire _359_;
wire _360_;
wire _361_;
wire _362_;
wire _363_;
wire _364_;
wire _365_;
wire _366_;
wire _367_;
wire _368_;
wire _369_;
wire _370_;
wire _371_;
wire _372_;
wire _373_;
wire _374_;
wire _375_;
wire _376_;
wire _377_;
wire _378_;
wire _379_;
wire _380_;
wire _381_;
wire _382_;
wire _383_;
wire _384_;
wire _385_;
wire _386_;
wire _387_;
wire _388_;
wire _389_;
wire _390_;
wire _391_;
wire _392_;
wire _393_;
wire _394_;
wire _395_;
wire _396_;
wire _397_;
wire _398_;
wire _399_;
wire _400_;
wire _401_;
wire _402_;
wire _403_;
wire _404_;
wire _405_;
wire _406_;
wire _407_;
wire _408_;
wire _409_;
wire _410_;
wire _411_;
wire _412_;
wire _413_;
wire _414_;
wire _415_;
wire _416_;
wire _417_;
wire _418_;
wire _419_;
wire _420_;
wire _421_;
wire _422_;
wire _423_;
wire _424_;
wire _425_;
wire _426_;
wire _427_;
wire _428_;
wire _429_;
wire _430_;
wire _431_;
wire _432_;
wire _433_;
wire _434_;
wire _435_;
wire _436_;
wire _437_;
wire _438_;
wire _439_;
wire _440_;
wire _441_;
wire _442_;
wire _443_;
wire _444_;
wire _445_;
wire _446_;
wire _447_;
wire _448_;
wire _449_;
wire _450_;
wire _451_;
wire _452_;
wire _453_;
wire _454_;
wire _455_;
wire _456_;
wire _457_;
wire _458_;
wire _459_;
wire _460_;
wire _461_;
wire _462_;
wire _463_;
wire _464_;
wire _465_;
wire _466_;
wire _467_;
wire _468_;
wire _469_;
wire _470_;
wire _471_;
wire _472_;
wire _473_;
wire _474_;
wire _475_;
wire _476_;
wire _477_;
wire _478_;
wire _479_;
wire _480_;
wire _481_;
wire _482_;
wire _483_;
wire _484_;
wire _485_;
wire _486_;
wire _487_;
wire _488_;
wire _489_;
wire _490_;
wire _491_;
wire _492_;
wire _493_;
wire _494_;
wire _495_;
wire _496_;
wire _497_;
wire _498_;
wire _499_;
wire _500_;
wire _501_;
wire _502_;
wire _503_;
wire _504_;
wire _505_;
wire _506_;
wire _507_;
wire _508_;
wire _509_;
wire _510_;
wire _511_;
wire _512_;
wire _513_;
wire _514_;
wire _515_;
wire _516_;
wire _517_;
wire _518_;
wire _519_;
wire _520_;
wire _521_;
wire _522_;
wire _523_;
wire _524_;
wire _525_;
wire _526_;
wire _527_;
wire _528_;
wire _529_;
wire _530_;
wire _531_;
wire _532_;
wire _533_;
wire _534_;
wire _535_;
wire _536_;
wire _537_;
wire _538_;
wire _539_;
wire _540_;
wire _541_;
wire _542_;
wire _543_;
wire _544_;
wire _545_;
wire _546_;
wire _547_;
wire _548_;
wire _549_;
wire _550_;
wire _551_;
wire _552_;
wire _553_;
wire _554_;
wire _555_;
wire _556_;
wire _557_;
wire _558_;
wire _559_;
wire _560_;
wire _561_;
wire _562_;
wire _563_;
wire _564_;
wire _565_;
wire _566_;
wire _567_;
wire _568_;
wire _569_;
wire _570_;
wire _571_;
wire _572_;
wire _573_;
wire _574_;
wire _575_;
wire _576_;
wire _577_;
wire _578_;
wire _579_;
wire _580_;
wire _581_;
wire _582_;
wire _583_;
wire _584_;
wire _585_;
wire _586_;
wire _587_;
wire _588_;
wire _589_;
wire _590_;
wire _591_;
wire _592_;
wire _593_;
wire _594_;
wire _595_;
wire _596_;
wire _597_;
wire _598_;
wire _599_;
wire _600_;
wire _601_;
wire _602_;
wire _603_;
wire _604_;
wire _605_;
wire _606_;
wire _607_;
wire _608_;
wire _609_;
wire _610_;
wire _611_;
wire _612_;
wire _613_;
wire _614_;
wire _615_;
wire _616_;
wire _617_;
wire _618_;
wire _619_;
wire _620_;
wire _621_;
wire _622_;
wire _623_;
wire _624_;
wire _625_;
wire _626_;
wire _627_;
wire _628_;
wire _629_;
wire _630_;
wire _631_;
wire _632_;
wire _633_;
wire _634_;
wire _635_;
wire _636_;
wire _637_;
wire _638_;
wire _639_;
wire _640_;
wire _641_;
wire _642_;
wire _643_;
wire _644_;
wire _645_;
wire _646_;
wire _647_;
wire _648_;
wire _649_;
wire _650_;
wire _651_;
wire _652_;
wire _653_;
wire _654_;
wire _655_;
wire _656_;
wire _657_;
wire _658_;
wire _659_;
wire _660_;
wire _661_;
wire _662_;
wire _663_;
wire _664_;
wire _665_;
wire _666_;
wire _667_;
wire _668_;
wire _669_;
wire _670_;
wire _671_;
wire _672_;
wire _673_;
wire _674_;
wire _675_;
wire _676_;
wire _677_;
wire _678_;
wire _679_;
wire _680_;
wire _681_;
wire _682_;
wire _683_;
wire _684_;
wire _685_;
wire _686_;
wire _687_;
wire _688_;
wire _689_;
wire _690_;
wire _691_;
wire _692_;
wire _693_;
wire _694_;
wire _695_;
wire _696_;
wire _697_;
wire _698_;
wire _699_;
wire _700_;
wire _701_;
wire _702_;
wire _703_;
wire _704_;
wire _705_;
wire _706_;
wire _707_;
wire _708_;
wire _709_;
wire _710_;
wire _711_;
wire _712_;
wire _713_;
wire _714_;
wire _715_;
wire _716_;
wire _717_;
wire _718_;
wire _719_;
wire _720_;
wire _721_;
wire _722_;
wire _723_;
wire _724_;
wire _725_;
wire _726_;
wire _727_;
wire _728_;
wire _729_;
wire _730_;
wire _731_;
wire _732_;
wire _733_;
wire _734_;
wire _735_;
wire _736_;
wire _737_;
wire _738_;
wire _739_;
wire _740_;
wire _741_;
wire _742_;
wire _743_;
wire _744_;
wire _745_;
wire _746_;
wire _747_;
wire _748_;
wire _749_;
wire _750_;
wire _751_;
wire _752_;
wire _753_;
wire _754_;
wire _755_;
wire _756_;
wire _757_;
wire _758_;
wire _759_;
wire _760_;
wire _761_;
wire _762_;
wire _763_;
wire _764_;
wire _765_;
wire _766_;
wire _767_;
wire _768_;
wire _769_;
wire _770_;
wire _771_;
wire _772_;
wire _773_;
wire _774_;
wire _775_;
wire _776_;
wire _777_;
wire _778_;
wire _779_;
wire _780_;
wire _781_;
wire _782_;
wire _783_;
wire _784_;
wire _785_;
wire _786_;
wire _787_;
wire _788_;
wire _789_;
wire _790_;
wire _791_;
wire _792_;
wire _793_;
wire _794_;
wire _795_;
wire _796_;
wire _797_;
wire _798_;
wire _799_;
wire _800_;
wire _801_;
wire _802_;
wire _803_;
wire _804_;
wire _805_;
wire _806_;
wire _807_;
wire _808_;
wire _809_;
wire _810_;
wire _811_;
wire _812_;
wire _813_;
wire _814_;
wire _815_;
wire _816_;
wire _817_;
wire _818_;
wire _819_;
wire _820_;
wire _821_;
wire _822_;
wire _823_;
wire _824_;
wire _825_;
wire _826_;
wire _827_;
wire _828_;
wire _829_;
wire _830_;
wire _831_;
wire _832_;
wire _833_;
wire _834_;
wire _835_;
wire _836_;
wire _837_;
wire _838_;
wire _839_;
wire _840_;
wire _841_;
wire _842_;
wire _843_;
wire _844_;
wire _845_;
wire _846_;
wire _847_;
wire _848_;
wire _849_;
wire _850_;
wire _851_;
wire _852_;
wire _853_;
wire _854_;
wire _855_;
wire _856_;
wire _857_;
wire _858_;
wire _859_;
wire _860_;
wire _861_;
wire _862_;
wire _863_;
wire _864_;
wire _865_;
wire _866_;
wire _867_;
wire _868_;
wire _869_;
wire _870_;
wire _871_;
wire _872_;
wire _873_;
wire _874_;
wire _875_;
wire _876_;
wire _877_;
wire _878_;
wire _879_;
wire _880_;
wire _881_;
wire _882_;
wire _883_;
wire _884_;
wire _885_;
wire _886_;
wire _887_;
wire _888_;
wire _889_;
wire _890_;
wire _891_;
wire _892_;
wire _893_;
wire _894_;
wire _895_;
wire _896_;
wire _897_;
wire _898_;
wire _899_;
wire _900_;
wire _901_;
wire _902_;
wire _903_;
wire _904_;
wire _905_;
wire _906_;
wire _907_;
wire _908_;
wire _909_;
wire _910_;
wire _911_;
wire _912_;
wire _913_;
wire _914_;
wire _915_;
wire _916_;
wire _917_;
wire _918_;
wire _919_;
wire _920_;
wire _921_;
wire _922_;
wire _923_;
wire _924_;
wire _925_;
wire _926_;
wire _927_;
wire _928_;
wire _929_;
wire _930_;
wire _931_;
wire _932_;
wire _933_;
wire _934_;
wire _935_;
wire _936_;
wire _937_;
wire _938_;
wire _939_;
wire _940_;
wire _941_;
wire _942_;
wire _943_;
wire _944_;
wire _945_;
wire _946_;
wire _947_;
wire _948_;
wire _949_;
wire _950_;
wire _951_;
wire _952_;
wire _953_;
wire _954_;
wire _955_;
wire _956_;
wire _957_;
wire _958_;
wire _959_;
wire _960_;
wire _961_;
wire _962_;
wire _963_;
wire _964_;
wire _965_;
wire _966_;
wire _967_;
wire _968_;
wire _969_;
wire _970_;
wire _971_;
wire _972_;
wire _973_;
wire _974_;
wire _975_;
wire _976_;
wire _977_;
wire _978_;
wire _979_;
wire _980_;
wire _981_;
wire _982_;
wire _983_;
wire _984_;
wire _985_;
wire _986_;
wire _987_;
wire _988_;
wire _989_;
wire _990_;
wire _991_;
wire _992_;
wire _993_;
wire _994_;
wire _995_;
wire _996_;
wire _997_;
wire _998_;
wire _999_;
wire _1000_;
wire _1001_;
wire _1002_;
wire _1003_;
wire _1004_;
wire _1005_;
wire _1006_;
wire _1007_;
wire _1008_;
wire _1009_;
wire _1010_;
wire _1011_;
wire _1012_;
wire _1013_;
wire _1014_;
wire _1015_;
wire _1016_;
wire _1017_;
wire _1018_;
wire _1019_;
wire _1020_;
wire _1021_;
wire _1022_;
wire _1023_;
wire _1024_;
wire _1025_;
wire _1026_;
wire _1027_;
wire _1028_;
wire _1029_;
wire _1030_;
wire _1031_;
wire _1032_;
wire _1033_;
wire _1034_;
wire _1035_;
wire _1036_;
wire _1037_;
wire _1038_;
wire _1039_;
wire _1040_;
wire _1041_;
wire _1042_;
wire _1043_;
wire _1044_;
wire _1045_;
wire _1046_;
wire _1047_;
wire _1048_;
wire _1049_;
wire _1050_;
wire _1051_;
wire _1052_;
wire _1053_;
wire _1054_;
wire _1055_;
wire _1056_;
wire _1057_;
wire _1058_;
wire _1059_;
wire _1060_;
wire _1061_;
wire _1062_;
wire _1063_;
wire _1064_;
wire _1065_;
wire _1066_;
wire _1067_;
wire _1068_;
wire _1069_;
wire _1070_;
wire _1071_;
wire _1072_;
wire _1073_;
wire _1074_;
wire _1075_;
wire _1076_;
wire _1077_;
wire _1078_;
wire _1079_;
wire _1080_;
wire _1081_;
wire _1082_;
wire _1083_;
wire _1084_;
wire _1085_;
wire _1086_;
wire _1087_;
wire _1088_;
wire _1089_;
wire _1090_;
wire _1091_;
wire _1092_;
wire _1093_;
wire _1094_;
wire _1095_;
wire _1096_;
wire _1097_;
wire _1098_;
wire _1099_;
wire _1100_;
wire _1101_;
wire _1102_;
wire _1103_;
wire _1104_;
wire _1105_;
wire _1106_;
wire _1107_;
wire _1108_;
wire _1109_;
wire _1110_;
wire _1111_;
wire _1112_;
wire _1113_;
wire _1114_;
wire _1115_;
wire _1116_;
wire _1117_;
wire _1118_;
wire _1119_;
wire _1120_;
wire _1121_;
wire _1122_;
wire _1123_;
wire _1124_;
wire _1125_;
wire _1126_;
wire _1127_;
wire _1128_;
wire _1129_;
wire _1130_;
wire _1131_;
wire _1132_;
wire _1133_;
wire _1134_;
wire _1135_;
wire _1136_;
wire _1137_;
wire _1138_;
wire _1139_;
wire _1140_;
wire _1141_;
wire _1142_;
wire _1143_;
wire _1144_;
wire _1145_;
wire _1146_;
wire _1147_;
wire _1148_;
wire _1149_;
wire _1150_;
wire _1151_;
wire _1152_;
wire _1153_;
wire _1154_;
wire _1155_;
wire _1156_;
wire _1157_;
wire _1158_;
wire _1159_;
wire _1160_;
wire _1161_;
wire _1162_;
wire _1163_;
wire _1164_;
wire _1165_;
wire _1166_;
wire _1167_;
wire _1168_;
wire _1169_;
wire _1170_;
wire _1171_;
wire _1172_;
wire _1173_;
wire _1174_;
wire _1175_;
wire _1176_;
wire _1177_;
wire _1178_;
wire _1179_;
wire _1180_;
wire _1181_;
wire _1182_;
wire _1183_;
wire _1184_;
wire _1185_;
wire _1186_;
wire _1187_;
wire _1188_;
wire _1189_;
wire _1190_;
wire _1191_;
wire _1192_;
wire _1193_;
wire _1194_;
wire _1195_;
wire _1196_;
wire _1197_;
wire _1198_;
wire _1199_;
wire _1200_;
wire _1201_;
wire _1202_;
wire _1203_;
wire _1204_;
wire _1205_;
wire _1206_;
wire _1207_;
wire _1208_;
wire _1209_;
wire _1210_;
wire _1211_;
wire _1212_;
wire _1213_;
wire _1214_;
wire _1215_;
wire _1216_;
wire _1217_;
wire _1218_;
wire _1219_;
wire _1220_;
wire _1221_;
wire _1222_;
wire _1223_;
wire _1224_;
wire _1225_;
wire _1226_;
wire _1227_;
wire _1228_;
wire _1229_;
wire _1230_;
wire _1231_;
wire _1232_;
wire _1233_;
wire _1234_;
wire _1235_;
wire _1236_;
wire _1237_;
wire _1238_;
wire _1239_;
wire _1240_;
wire _1241_;
wire _1242_;
wire _1243_;
wire _1244_;
wire _1245_;
wire _1246_;
wire _1247_;
wire _1248_;
wire _1249_;
wire _1250_;
wire _1251_;
wire _1252_;
wire _1253_;
wire _1254_;
wire _1255_;
wire _1256_;
wire _1257_;
wire _1258_;
wire _1259_;
wire _1260_;
wire _1261_;
wire _1262_;
wire _1263_;
wire _1264_;
wire _1265_;
wire _1266_;
wire _1267_;
wire _1268_;
wire _1269_;
wire _1270_;
wire _1271_;
wire _1272_;
wire _1273_;
wire _1274_;
wire _1275_;
wire _1276_;
wire _1277_;
wire _1278_;
wire _1279_;
wire _1280_;
wire _1281_;
wire _1282_;
wire _1283_;
wire _1284_;
wire _1285_;
wire _1286_;
wire _1287_;
wire _1288_;
wire _1289_;
wire _1290_;
wire _1291_;
wire _1292_;
wire _1293_;
wire _1294_;
wire _1295_;
wire _1296_;
wire _1297_;
wire _1298_;
wire _1299_;
wire _1300_;
wire _1301_;
wire _1302_;
wire _1303_;
wire _1304_;
wire _1305_;
wire _1306_;
wire _1307_;
wire _1308_;
wire _1309_;
wire _1310_;
wire _1311_;
wire _1312_;
wire _1313_;
wire _1314_;
wire _1315_;
wire _1316_;
wire _1317_;
wire _1318_;
wire _1319_;
wire _1320_;
wire _1321_;
wire _1322_;
wire _1323_;
wire _1324_;
wire _1325_;
wire _1326_;
wire _1327_;
wire _1328_;
wire _1329_;
wire _1330_;
wire _1331_;
wire _1332_;
wire _1333_;
wire _1334_;
wire _1335_;
wire _1336_;
wire _1337_;
wire _1338_;
wire _1339_;
wire _1340_;
wire _1341_;
wire _1342_;
wire _1343_;
wire _1344_;
wire _1345_;
wire _1346_;
wire _1347_;
wire _1348_;
wire _1349_;
wire _1350_;
wire _1351_;
wire _1352_;
wire _1353_;
wire _1354_;
wire _1355_;
wire _1356_;
wire _1357_;
wire _1358_;
wire _1359_;
wire _1360_;
wire _1361_;
wire _1362_;
wire _1363_;
wire _1364_;
wire _1365_;
wire _1366_;
wire _1367_;
wire _1368_;
wire _1369_;
wire _1370_;
wire _1371_;
wire _1372_;
wire _1373_;
wire _1374_;
wire _1375_;
wire _1376_;
wire _1377_;
wire _1378_;
wire _1379_;
wire _1380_;
wire _1381_;
wire _1382_;
wire _1383_;
wire _1384_;
wire _1385_;
wire _1386_;
wire _1387_;
wire _1388_;
wire _1389_;
wire _1390_;
wire _1391_;
wire _1392_;
wire _1393_;
wire _1394_;
wire _1395_;
wire _1396_;
wire _1397_;
wire _1398_;
wire _1399_;
wire _1400_;
wire _1401_;
wire _1402_;
wire _1403_;
wire _1404_;
wire _1405_;
wire _1406_;
wire _1407_;
wire _1408_;
wire _1409_;
wire _1410_;
wire _1411_;
wire _1412_;
wire _1413_;
wire _1414_;
wire _1415_;
wire _1416_;
wire _1417_;
wire _1418_;
wire _1419_;
wire _1420_;
wire _1421_;
wire _1422_;
wire _1423_;
wire _1424_;
wire _1425_;
wire _1426_;
wire _1427_;
wire _1428_;
wire _1429_;
wire _1430_;
wire _1431_;
wire _1432_;
wire _1433_;
wire _1434_;
wire _1435_;
wire _1436_;
wire _1437_;
wire _1438_;
wire _1439_;
wire _1440_;
wire _1441_;
wire _1442_;
wire _1443_;
wire _1444_;
wire _1445_;
wire _1446_;
wire _1447_;
wire _1448_;
wire _1449_;
wire _1450_;
wire _1451_;
wire _1452_;
wire _1453_;
wire _1454_;
wire _1455_;
wire _1456_;
wire _1457_;
wire _1458_;
wire _1459_;
wire _1460_;
wire _1461_;
wire _1462_;
wire _1463_;
wire _1464_;
wire _1465_;
wire _1466_;
wire _1467_;
wire _1468_;
wire _1469_;
wire _1470_;
wire _1471_;
wire _1472_;
wire _1473_;
wire _1474_;
wire _1475_;
wire _1476_;
wire _1477_;
wire _1478_;
wire _1479_;
wire _1480_;
wire _1481_;
wire _1482_;
wire _1483_;
wire _1484_;
wire _1485_;
wire _1486_;
wire _1487_;
wire _1488_;
wire _1489_;
wire _1490_;
wire _1491_;
wire _1492_;
wire _1493_;
wire _1494_;
wire _1495_;
wire _1496_;
wire _1497_;
wire _1498_;
wire _1499_;
wire _1500_;
wire _1501_;
wire _1502_;
wire _1503_;
wire _1504_;
wire _1505_;
wire _1506_;
wire _1507_;
wire _1508_;
wire _1509_;
wire _1510_;
wire _1511_;
wire _1512_;
wire _1513_;
wire _1514_;
wire _1515_;
wire _1516_;
wire _1517_;
wire _1518_;
wire _1519_;
wire _1520_;
wire _1521_;
wire _1522_;
wire _1523_;
wire _1524_;
wire _1525_;
wire _1526_;
wire _1527_;
wire _1528_;
wire _1529_;
wire _1530_;
wire _1531_;
wire _1532_;
wire _1533_;
wire _1534_;
wire _1535_;
wire _1536_;
wire _1537_;
wire _1538_;
wire _1539_;
wire _1540_;
wire _1541_;
wire _1542_;
wire _1543_;
wire _1544_;
wire _1545_;
wire _1546_;
wire _1547_;
wire _1548_;
wire _1549_;
wire _1550_;
wire _1551_;
wire _1552_;
wire _1553_;
wire _1554_;
wire _1555_;
wire _1556_;
wire _1557_;
wire _1558_;
wire _1559_;
wire _1560_;
wire _1561_;
wire _1562_;
wire _1563_;
wire _1564_;
wire _1565_;
wire _1566_;
wire _1567_;
wire _1568_;
wire _1569_;
wire _1570_;
wire _1571_;
wire _1572_;
wire _1573_;
wire _1574_;
wire _1575_;
wire _1576_;
wire _1577_;
wire _1578_;
wire _1579_;
wire _1580_;
wire _1581_;
wire _1582_;
wire _1583_;
wire _1584_;
wire _1585_;
wire _1586_;
wire _1587_;
wire _1588_;
wire _1589_;
wire _1590_;
wire _1591_;
wire _1592_;
wire _1593_;
wire _1594_;
wire _1595_;
wire _1596_;
wire _1597_;
wire _1598_;
wire _1599_;
wire _1600_;
wire _1601_;
wire _1602_;
wire _1603_;
wire _1604_;
wire _1605_;
wire _1606_;
wire _1607_;
wire _1608_;
wire _1609_;
wire _1610_;
wire _1611_;
wire _1612_;
wire _1613_;
wire _1614_;
wire _1615_;
wire _1616_;
wire _1617_;
wire _1618_;
wire _1619_;
wire _1620_;
wire _1621_;
wire _1622_;
wire _1623_;
wire _1624_;
wire _1625_;
wire _1626_;
wire _1627_;
wire _1628_;
wire _1629_;
wire _1630_;
wire _1631_;
wire _1632_;
wire _1633_;
wire _1634_;
wire _1635_;
wire _1636_;
wire _1637_;
wire _1638_;
wire _1639_;
wire _1640_;
wire _1641_;
wire _1642_;
wire _1643_;
wire _1644_;
wire _1645_;
wire _1646_;
wire _1647_;
wire _1648_;
wire _1649_;
wire _1650_;
wire _1651_;
wire _1652_;
wire _1653_;
wire _1654_;
wire _1655_;
wire _1656_;
wire _1657_;
wire _1658_;
wire _1659_;
wire _1660_;
wire _1661_;
wire _1662_;
wire _1663_;
wire _1664_;
wire _1665_;
wire _1666_;
wire _1667_;
wire _1668_;
wire _1669_;
wire _1670_;
wire _1671_;
wire _1672_;
wire _1673_;
wire _1674_;
wire _1675_;
wire _1676_;
wire _1677_;
wire _1678_;
wire _1679_;
wire _1680_;
wire _1681_;
wire _1682_;
wire _1683_;
wire _1684_;
wire _1685_;
wire _1686_;
wire _1687_;
wire _1688_;
wire _1689_;
wire _1690_;
wire _1691_;
wire _1692_;
wire _1693_;
wire _1694_;
wire _1695_;
wire _1696_;
wire _1697_;
wire _1698_;
wire _1699_;
wire _1700_;
wire _1701_;
wire _1702_;
wire _1703_;
wire _1704_;
wire _1705_;
wire _1706_;
wire _1707_;
wire _1708_;
wire _1709_;
wire _1710_;
wire _1711_;
wire _1712_;
wire _1713_;
wire _1714_;
wire _1715_;
wire _1716_;
wire _1717_;
wire _1718_;
wire _1719_;
wire _1720_;
wire _1721_;
wire _1722_;
wire _1723_;
wire _1724_;
wire _1725_;
wire _1726_;
wire _1727_;
wire _1728_;
wire _1729_;
wire _1730_;
wire _1731_;
wire _1732_;
wire _1733_;
wire _1734_;
wire _1735_;
wire _1736_;
wire _1737_;
wire _1738_;
wire _1739_;
wire _1740_;
wire _1741_;
wire _1742_;
wire _1743_;
wire _1744_;
wire _1745_;
wire _1746_;
wire _1747_;
wire _1748_;
wire _1749_;
wire _1750_;
wire _1751_;
wire _1752_;
wire _1753_;
wire _1754_;
wire _1755_;
wire _1756_;
wire _1757_;
wire _1758_;
wire _1759_;
wire _1760_;
wire _1761_;
wire _1762_;
wire _1763_;
wire _1764_;
wire _1765_;
wire _1766_;
wire _1767_;
wire _1768_;
wire _1769_;
wire _1770_;
wire _1771_;
wire _1772_;
wire _1773_;
wire _1774_;
wire _1775_;
wire _1776_;
wire _1777_;
wire _1778_;
wire _1779_;
wire _1780_;
wire _1781_;
wire _1782_;
wire _1783_;
wire _1784_;
wire _1785_;
wire _1786_;
wire _1787_;
wire _1788_;
wire _1789_;
wire _1790_;
wire _1791_;
wire _1792_;
wire _1793_;
wire _1794_;
wire _1795_;
wire _1796_;
wire _1797_;
wire _1798_;
wire _1799_;
wire _1800_;
wire _1801_;
wire _1802_;
wire _1803_;
wire _1804_;
wire _1805_;
wire _1806_;
wire _1807_;
wire _1808_;
wire _1809_;
wire _1810_;
wire _1811_;
wire _1812_;
wire _1813_;
wire _1814_;
wire _1815_;
wire _1816_;
wire _1817_;
wire _1818_;
wire _1819_;
wire _1820_;
wire _1821_;
wire _1822_;
wire _1823_;
wire _1824_;
wire _1825_;
wire _1826_;
wire _1827_;
wire _1828_;
wire _1829_;
wire _1830_;
wire _1831_;
wire _1832_;
wire _1833_;
wire _1834_;
wire _1835_;
wire _1836_;
wire _1837_;
wire _1838_;
wire _1839_;
wire _1840_;
wire _1841_;
wire _1842_;
wire _1843_;
wire _1844_;
wire _1845_;
wire _1846_;
wire _1847_;
wire _1848_;
wire _1849_;
wire _1850_;
wire _1851_;
wire _1852_;
wire _1853_;
wire _1854_;
wire _1855_;
wire _1856_;
wire _1857_;
wire _1858_;
wire _1859_;
wire _1860_;
wire _1861_;
wire _1862_;
wire _1863_;
wire _1864_;
wire _1865_;
wire _1866_;
wire _1867_;
wire _1868_;
wire _1869_;
wire _1870_;
wire _1871_;
wire _1872_;
wire _1873_;
wire _1874_;
wire _1875_;
wire _1876_;
wire _1877_;
wire _1878_;
wire _1879_;
wire _1880_;
wire _1881_;
wire _1882_;
wire _1883_;
wire _1884_;
wire _1885_;
wire _1886_;
wire _1887_;
wire _1888_;
wire _1889_;
wire _1890_;
wire _1891_;
wire _1892_;
wire _1893_;
wire _1894_;
wire _1895_;
wire _1896_;
wire _1897_;
wire _1898_;
wire _1899_;
wire _1900_;
wire _1901_;
wire _1902_;
wire _1903_;
wire _1904_;
wire _1905_;
wire _1906_;
wire _1907_;
wire _1908_;
wire _1909_;
wire _1910_;
wire _1911_;
wire _1912_;
wire _1913_;
wire _1914_;
wire _1915_;
wire _1916_;
wire _1917_;
wire _1918_;
wire _1919_;
wire _1920_;
wire _1921_;
wire _1922_;
wire _1923_;
wire _1924_;
wire _1925_;
wire _1926_;
wire _1927_;
wire _1928_;
wire _1929_;
wire _1930_;
wire _1931_;
wire _1932_;
wire _1933_;
wire _1934_;
wire _1935_;
wire _1936_;
wire _1937_;
wire _1938_;
wire _1939_;
wire _1940_;
wire _1941_;
wire _1942_;
wire _1943_;
wire _1944_;
wire _1945_;
wire _1946_;
wire _1947_;
wire _1948_;
wire _1949_;
wire _1950_;
wire _1951_;
wire _1952_;
wire _1953_;
wire _1954_;
wire _1955_;
wire _1956_;
wire _1957_;
wire _1958_;
wire _1959_;
wire _1960_;
wire _1961_;
wire _1962_;
wire _1963_;
wire _1964_;
wire _1965_;
wire _1966_;
wire _1967_;
wire _1968_;
wire _1969_;
wire _1970_;
wire _1971_;
wire _1972_;
wire _1973_;
wire _1974_;
wire _1975_;
wire _1976_;
wire _1977_;
wire _1978_;
wire _1979_;
wire _1980_;
wire _1981_;
wire _1982_;
wire _1983_;
wire _1984_;
wire _1985_;
wire _1986_;
wire _1987_;
wire _1988_;
wire _1989_;
wire _1990_;
wire _1991_;
wire _1992_;
wire _1993_;
wire _1994_;
wire _1995_;
wire _1996_;
wire _1997_;
wire _1998_;
wire _1999_;
wire _2000_;
wire _2001_;
wire _2002_;
wire _2003_;
wire _2004_;
wire _2005_;
wire _2006_;
wire _2007_;
wire _2008_;
wire _2009_;
wire _2010_;
wire _2011_;
wire _2012_;
wire _2013_;
wire _2014_;
wire _2015_;
wire _2016_;
wire _2017_;
wire _2018_;
wire _2019_;
wire _2020_;
wire _2021_;
wire _2022_;
wire _2023_;
wire _2024_;
wire _2025_;
wire _2026_;
wire _2027_;
wire _2028_;
wire _2029_;
wire _2030_;
wire _2031_;
wire _2032_;
wire _2033_;
wire _2034_;
wire _2035_;
wire _2036_;
wire _2037_;
wire _2038_;
wire _2039_;
wire _2040_;
wire _2041_;
wire _2042_;
wire _2043_;
wire _2044_;
wire _2045_;
wire _2046_;
wire _2047_;
wire _2048_;
wire _2049_;
wire _2050_;
wire _2051_;
wire _2052_;
wire _2053_;
wire _2054_;
wire _2055_;
wire _2056_;
wire _2057_;
wire _2058_;
wire _2059_;
wire _2060_;
wire _2061_;
wire _2062_;
wire _2063_;
wire _2064_;
wire _2065_;
wire _2066_;
wire _2067_;
wire _2068_;
wire _2069_;
wire _2070_;
wire _2071_;
wire _2072_;
wire _2073_;
wire _2074_;
wire _2075_;
wire _2076_;
wire _2077_;
wire _2078_;
wire _2079_;
wire _2080_;
wire _2081_;
wire _2082_;
wire _2083_;
wire _2084_;
wire _2085_;
wire _2086_;
wire _2087_;
wire _2088_;
wire _2089_;
wire _2090_;
wire _2091_;
wire _2092_;
wire _2093_;
wire _2094_;
wire _2095_;
wire _2096_;
wire _2097_;
wire _2098_;
wire _2099_;
wire _2100_;
wire _2101_;
wire _2102_;
wire _2103_;
wire _2104_;
wire _2105_;
wire _2106_;
wire _2107_;
wire _2108_;
wire _2109_;
wire _2110_;
wire _2111_;
wire _2112_;
wire _2113_;
wire _2114_;
wire _2115_;
wire _2116_;
wire _2117_;
wire _2118_;
wire _2119_;
wire _2120_;
wire _2121_;
wire _2122_;
wire _2123_;
wire _2124_;
wire _2125_;
wire _2126_;
wire _2127_;
wire _2128_;
wire _2129_;
wire _2130_;
wire _2131_;
wire _2132_;
wire _2133_;
wire _2134_;
wire _2135_;
wire _2136_;
wire _2137_;
wire _2138_;
wire _2139_;
wire _2140_;
wire _2141_;
wire _2142_;
wire _2143_;
wire _2144_;
wire _2145_;
wire _2146_;
wire _2147_;
wire _2148_;
wire _2149_;
wire _2150_;
wire _2151_;
wire _2152_;
wire _2153_;
wire _2154_;
wire _2155_;
wire _2156_;
wire _2157_;
wire _2158_;
wire _2159_;
wire _2160_;
wire _2161_;
wire _2162_;
wire _2163_;
wire _2164_;
wire _2165_;
wire _2166_;
wire _2167_;
wire _2168_;
wire _2169_;
wire _2170_;
wire _2171_;
wire _2172_;
wire _2173_;
wire _2174_;
wire _2175_;
wire _2176_;
wire _2177_;
wire _2178_;
wire _2179_;
wire _2180_;
wire _2181_;
wire _2182_;
wire _2183_;
wire _2184_;
wire _2185_;
wire _2186_;
wire _2187_;
wire _2188_;
wire _2189_;
wire _2190_;
wire _2191_;
wire _2192_;
wire _2193_;
wire _2194_;
wire _2195_;
wire _2196_;
wire _2197_;
wire _2198_;
wire _2199_;
wire _2200_;
wire _2201_;
wire _2202_;
wire _2203_;
wire _2204_;
wire _2205_;
wire _2206_;
wire _2207_;
wire _2208_;
wire _2209_;
wire _2210_;
wire _2211_;
wire _2212_;
wire _2213_;
wire _2214_;
wire _2215_;
wire _2216_;
wire _2217_;
wire _2218_;
wire _2219_;
wire _2220_;
wire _2221_;
wire _2222_;
wire _2223_;
wire _2224_;
wire _2225_;
wire _2226_;
wire _2227_;
wire _2228_;
wire _2229_;
wire _2230_;
wire _2231_;
wire _2232_;
wire _2233_;
wire _2234_;
wire _2235_;
wire _2236_;
wire _2237_;
wire _2238_;
wire _2239_;
wire _2240_;
wire _2241_;
wire _2242_;
wire _2243_;
wire _2244_;
wire _2245_;
wire _2246_;
wire _2247_;
wire _2248_;
wire _2249_;
wire _2250_;
wire _2251_;
wire _2252_;
wire _2253_;
wire _2254_;
wire _2255_;
wire _2256_;
wire _2257_;
wire _2258_;
wire _2259_;
wire _2260_;
wire _2261_;
wire _2262_;
wire _2263_;
wire _2264_;
wire _2265_;
wire _2266_;
wire _2267_;
wire _2268_;
wire _2269_;
wire _2270_;
wire _2271_;
wire _2272_;
wire _2273_;
wire _2274_;
wire _2275_;
wire _2276_;
wire _2277_;
wire _2278_;
wire _2279_;
wire _2280_;
wire _2281_;
wire _2282_;
wire _2283_;
wire _2284_;
wire _2285_;
wire _2286_;
wire _2287_;
wire _2288_;
wire _2289_;
wire _2290_;
wire _2291_;
wire _2292_;
wire _2293_;
wire _2294_;
wire _2295_;
wire _2296_;
wire _2297_;
wire _2298_;
wire _2299_;
wire _2300_;
wire _2301_;
wire _2302_;
wire _2303_;
wire _2304_;
wire _2305_;
wire _2306_;
wire _2307_;
wire _2308_;
wire _2309_;
wire _2310_;
wire _2311_;
wire _2312_;
wire _2313_;
wire _2314_;
wire _2315_;
wire _2316_;
wire _2317_;
wire _2318_;
wire _2319_;
wire _2320_;
wire _2321_;
wire _2322_;
wire _2323_;
wire _2324_;
wire _2325_;
wire _2326_;
wire _2327_;
wire _2328_;
wire _2329_;
wire _2330_;
wire _2331_;
wire _2332_;
wire _2333_;
wire _2334_;
wire _2335_;
wire _2336_;
wire _2337_;
wire _2338_;
wire _2339_;
wire _2340_;
wire _2341_;
wire _2342_;
wire _2343_;
wire _2344_;
wire _2345_;
wire _2346_;
wire _2347_;
wire _2348_;
wire _2349_;
wire _2350_;
wire _2351_;
wire _2352_;
wire _2353_;
wire _2354_;
wire _2355_;
wire _2356_;
wire _2357_;
wire _2358_;
wire _2359_;
wire _2360_;
wire _2361_;
wire _2362_;
wire _2363_;
wire _2364_;
wire _2365_;
wire _2366_;
wire _2367_;
wire _2368_;
wire _2369_;
wire _2370_;
wire _2371_;
wire _2372_;
wire _2373_;
wire _2374_;
wire _2375_;
wire _2376_;
wire _2377_;
wire _2378_;
wire _2379_;
wire _2380_;
wire _2381_;
wire _2382_;
wire _2383_;
wire _2384_;
wire _2385_;
wire _2386_;
wire _2387_;
wire _2388_;
wire _2389_;
wire _2390_;
wire _2391_;
wire _2392_;
wire _2393_;
wire _2394_;
wire _2395_;
wire _2396_;
wire _2397_;
wire _2398_;
wire _2399_;
wire _2400_;
wire _2401_;
wire _2402_;
wire _2403_;
wire _2404_;
wire _2405_;
wire _2406_;
wire _2407_;
wire _2408_;
wire _2409_;
wire _2410_;
wire _2411_;
wire _2412_;
wire _2413_;
wire _2414_;
wire _2415_;
wire _2416_;
wire _2417_;
wire _2418_;
wire _2419_;
wire _2420_;
wire _2421_;
wire _2422_;
wire _2423_;
wire _2424_;
wire _2425_;
wire _2426_;
wire _2427_;
wire _2428_;
wire _2429_;
wire _2430_;
wire _2431_;
wire _2432_;
wire _2433_;
wire _2434_;
wire _2435_;
wire _2436_;
wire _2437_;
wire _2438_;
wire _2439_;
wire _2440_;
wire _2441_;
wire _2442_;
wire _2443_;
wire _2444_;
wire _2445_;
wire _2446_;
wire _2447_;
wire _2448_;
wire _2449_;
wire _2450_;
wire _2451_;
wire _2452_;
wire _2453_;
wire _2454_;
wire _2455_;
wire _2456_;
wire _2457_;
wire _2458_;
wire _2459_;
wire _2460_;
wire _2461_;
wire _2462_;
wire _2463_;
wire _2464_;
wire _2465_;
wire _2466_;
wire _2467_;
wire _2468_;
wire _2469_;
wire _2470_;
wire _2471_;
wire _2472_;
wire _2473_;
wire _2474_;
wire _2475_;
wire _2476_;
wire _2477_;
wire _2478_;
wire _2479_;
wire _2480_;
wire _2481_;
wire _2482_;
wire _2483_;
wire _2484_;
wire _2485_;
wire _2486_;
wire _2487_;
wire _2488_;
wire _2489_;
wire _2490_;
wire _2491_;
wire _2492_;
wire _2493_;
wire _2494_;
wire _2495_;
wire _2496_;
wire _2497_;
wire _2498_;
wire _2499_;
wire _2500_;
wire _2501_;
wire _2502_;
wire _2503_;
wire _2504_;
wire _2505_;
wire _2506_;
wire _2507_;
wire _2508_;
wire _2509_;
wire _2510_;
wire _2511_;
wire _2512_;
wire _2513_;
wire _2514_;
wire _2515_;
wire _2516_;
wire _2517_;
wire _2518_;
wire _2519_;
wire _2520_;
wire _2521_;
wire _2522_;
wire _2523_;
wire _2524_;
wire _2525_;
wire _2526_;
wire _2527_;
wire _2528_;
wire _2529_;
wire _2530_;
wire _2531_;
wire _2532_;
wire _2533_;
wire _2534_;
wire _2535_;
wire _2536_;
wire _2537_;
wire _2538_;
wire _2539_;
wire _2540_;
wire _2541_;
wire _2542_;
wire _2543_;
wire _2544_;
wire _2545_;
wire _2546_;
wire _2547_;
wire _2548_;
wire _2549_;
wire _2550_;
wire _2551_;
wire _2552_;
wire _2553_;
wire _2554_;
wire _2555_;
wire _2556_;
wire _2557_;
wire _2558_;
wire _2559_;
wire _2560_;
wire _2561_;
wire _2562_;
wire _2563_;
wire _2564_;
wire _2565_;
wire _2566_;
wire _2567_;
wire _2568_;
wire _2569_;
wire _2570_;
wire _2571_;
wire _2572_;
wire _2573_;
wire _2574_;
wire _2575_;
wire _2576_;
wire _2577_;
wire _2578_;
wire _2579_;
wire _2580_;
wire _2581_;
wire _2582_;
wire _2583_;
wire _2584_;
wire _2585_;
wire _2586_;
wire _2587_;
wire _2588_;
wire _2589_;
wire _2590_;
wire _2591_;
wire _2592_;
wire _2593_;
wire _2594_;
wire _2595_;
wire _2596_;
wire _2597_;
wire _2598_;
wire _2599_;
wire _2600_;
wire _2601_;
wire _2602_;
wire _2603_;
wire _2604_;
wire _2605_;
wire _2606_;
wire _2607_;
wire _2608_;
wire _2609_;
wire _2610_;
wire _2611_;
wire _2612_;
wire _2613_;
wire _2614_;
wire _2615_;
wire _2616_;
wire _2617_;
wire _2618_;
wire _2619_;
wire _2620_;
wire _2621_;
wire _2622_;
wire _2623_;
wire _2624_;
wire _2625_;
wire _2626_;
wire _2627_;
wire _2628_;
wire _2629_;
wire _2630_;
wire _2631_;
wire _2632_;
wire _2633_;
wire _2634_;
wire _2635_;
wire _2636_;
wire _2637_;
wire _2638_;
wire _2639_;
wire _2640_;
wire _2641_;
wire _2642_;
wire _2643_;
wire _2644_;
wire _2645_;
wire _2646_;
wire _2647_;
wire _2648_;
wire _2649_;
wire _2650_;
wire _2651_;
wire _2652_;
wire _2653_;
wire _2654_;
wire _2655_;
wire _2656_;
wire _2657_;
wire _2658_;
wire _2659_;
wire _2660_;
wire _2661_;
wire _2662_;
wire _2663_;
wire _2664_;
wire _2665_;
wire _2666_;
wire _2667_;
wire _2668_;
wire _2669_;
wire _2670_;
wire _2671_;
wire _2672_;
wire _2673_;
wire _2674_;
wire _2675_;
wire _2676_;
wire _2677_;
wire _2678_;
wire _2679_;
wire _2680_;
wire _2681_;
wire _2682_;
wire _2683_;
wire _2684_;
wire _2685_;
wire _2686_;
wire _2687_;
wire _2688_;
wire _2689_;
wire _2690_;
wire _2691_;
wire _2692_;
wire _2693_;
wire _2694_;
wire _2695_;
wire _2696_;
wire _2697_;
wire _2698_;
wire _2699_;
wire _2700_;
wire _2701_;
wire _2702_;
wire _2703_;
wire _2704_;
wire _2705_;
wire _2706_;
wire _2707_;
wire _2708_;
wire _2709_;
wire _2710_;
wire _2711_;
wire _2712_;
wire _2713_;
wire _2714_;
wire _2715_;
wire _2716_;
wire _2717_;
wire _2718_;
wire _2719_;
wire _2720_;
wire _2721_;
wire _2722_;
wire _2723_;
wire _2724_;
wire _2725_;
wire _2726_;
wire _2727_;
wire _2728_;
wire _2729_;
wire _2730_;
wire _2731_;
wire _2732_;
wire _2733_;
wire _2734_;
wire _2735_;
wire _2736_;
wire _2737_;
wire _2738_;
wire _2739_;
wire _2740_;
wire _2741_;
wire _2742_;
wire _2743_;
wire _2744_;
wire _2745_;
wire _2746_;
wire _2747_;
wire _2748_;
wire _2749_;
wire _2750_;
wire _2751_;
wire _2752_;
wire _2753_;
wire _2754_;
wire _2755_;
wire _2756_;
wire _2757_;
wire _2758_;
wire _2759_;
wire _2760_;
wire _2761_;
wire _2762_;
wire _2763_;
wire _2764_;
wire _2765_;
wire _2766_;
wire _2767_;
wire _2768_;
wire _2769_;
wire _2770_;
wire _2771_;
wire _2772_;
wire _2773_;
wire _2774_;
wire _2775_;
wire _2776_;
wire _2777_;
wire _2778_;
wire _2779_;
wire _2780_;
wire _2781_;
wire _2782_;
wire _2783_;
wire _2784_;
wire _2785_;
wire _2786_;
wire _2787_;
wire _2788_;
wire _2789_;
wire _2790_;
wire _2791_;
wire _2792_;
wire _2793_;
wire _2794_;
wire _2795_;
wire _2796_;
wire _2797_;
wire _2798_;
wire _2799_;
wire _2800_;
wire _2801_;
wire _2802_;
wire _2803_;
wire _2804_;
wire _2805_;
wire _2806_;
wire _2807_;
wire _2808_;
wire _2809_;
wire _2810_;
wire _2811_;
wire _2812_;
wire _2813_;
wire _2814_;
wire _2815_;
wire _2816_;
wire _2817_;
wire _2818_;
wire _2819_;
wire _2820_;
wire _2821_;
wire _2822_;
wire _2823_;
wire _2824_;
wire _2825_;
wire _2826_;
wire _2827_;
wire _2828_;
wire _2829_;
wire _2830_;
wire _2831_;
wire _2832_;
wire _2833_;
wire _2834_;
wire _2835_;
wire _2836_;
wire _2837_;
wire _2838_;
wire _2839_;
wire _2840_;
wire _2841_;
wire _2842_;
wire _2843_;
wire _2844_;
wire _2845_;
wire _2846_;
wire _2847_;
wire _2848_;
wire _2849_;
wire _2850_;
wire _2851_;
wire _2852_;
wire _2853_;
wire _2854_;
wire _2855_;
wire _2856_;
wire _2857_;
wire _2858_;
wire _2859_;
wire _2860_;
wire _2861_;
wire _2862_;
wire _2863_;
wire _2864_;
wire _2865_;
wire _2866_;
wire _2867_;
wire _2868_;
wire _2869_;
wire _2870_;
wire _2871_;
wire _2872_;
wire _2873_;
wire _2874_;
wire _2875_;
wire _2876_;
wire _2877_;
wire _2878_;
wire _2879_;
wire _2880_;
wire _2881_;
wire _2882_;
wire _2883_;
wire _2884_;
wire _2885_;
wire _2886_;
wire _2887_;
wire _2888_;
wire _2889_;
wire _2890_;
wire _2891_;
wire _2892_;
wire _2893_;
wire _2894_;
wire _2895_;
wire _2896_;
wire _2897_;
wire _2898_;
wire _2899_;
wire _2900_;
wire _2901_;
wire _2902_;
wire _2903_;
wire _2904_;
wire _2905_;
wire _2906_;
wire _2907_;
wire _2908_;
wire _2909_;
wire _2910_;
wire _2911_;
wire _2912_;
wire _2913_;
wire _2914_;
wire _2915_;
wire _2916_;
wire _2917_;
wire _2918_;
wire _2919_;
wire _2920_;
wire _2921_;
wire _2922_;
wire _2923_;
wire _2924_;
wire _2925_;
wire _2926_;
wire _2927_;
wire _2928_;
wire _2929_;
wire _2930_;
wire _2931_;
wire _2932_;
wire _2933_;
wire _2934_;
wire _2935_;
wire _2936_;
wire _2937_;
wire _2938_;
wire _2939_;
wire _2940_;
wire _2941_;
wire _2942_;
wire _2943_;
wire _2944_;
wire _2945_;
wire _2946_;
wire _2947_;
wire _2948_;
wire _2949_;
wire _2950_;
wire _2951_;
wire _2952_;
wire _2953_;
wire _2954_;
wire _2955_;
wire _2956_;
wire _2957_;
wire _2958_;
wire _2959_;
wire _2960_;
wire _2961_;
wire _2962_;
wire _2963_;
wire _2964_;
wire _2965_;
wire _2966_;
wire _2967_;
wire _2968_;
wire _2969_;
wire _2970_;
wire _2971_;
wire _2972_;
wire _2973_;
wire _2974_;
wire _2975_;
wire _2976_;
wire _2977_;
wire _2978_;
wire _2979_;
wire _2980_;
wire _2981_;
wire _2982_;
wire _2983_;
wire _2984_;
wire _2985_;
wire _2986_;
wire _2987_;
wire _2988_;
wire _2989_;
wire _2990_;
wire _2991_;
wire _2992_;
wire _2993_;
wire _2994_;
wire _2995_;
wire _2996_;
wire _2997_;
wire _2998_;
wire _2999_;
wire _3000_;
wire _3001_;
wire _3002_;
wire _3003_;
wire _3004_;
wire _3005_;
wire _3006_;
wire _3007_;
wire _3008_;
wire _3009_;
wire _3010_;
wire _3011_;
wire _3012_;
wire _3013_;
wire _3014_;
wire _3015_;
wire _3016_;
wire _3017_;
wire _3018_;
wire _3019_;
wire _3020_;
wire _3021_;
wire _3022_;
wire _3023_;
wire _3024_;
wire _3025_;
wire _3026_;
wire _3027_;
wire _3028_;
wire _3029_;
wire _3030_;
wire _3031_;
wire _3032_;
wire _3033_;
wire _3034_;
wire _3035_;
wire _3036_;
wire _3037_;
wire _3038_;
wire _3039_;
wire _3040_;
wire _3041_;
wire _3042_;
wire _3043_;
wire _3044_;
wire _3045_;
wire _3046_;
wire _3047_;
wire _3048_;
wire _3049_;
wire _3050_;
wire _3051_;
wire _3052_;
wire _3053_;
wire _3054_;
wire _3055_;
wire _3056_;
wire _3057_;
wire _3058_;
wire _3059_;
wire _3060_;
wire _3061_;
wire _3062_;
wire _3063_;
wire _3064_;
wire _3065_;
wire _3066_;
wire _3067_;
wire _3068_;
wire _3069_;
wire _3070_;
wire _3071_;
wire _3072_;
wire _3073_;
wire _3074_;
wire _3075_;
wire _3076_;
wire _3077_;
wire _3078_;
wire _3079_;
wire _3080_;
wire _3081_;
wire _3082_;
wire _3083_;
wire _3084_;
wire _3085_;
wire _3086_;
wire _3087_;
wire _3088_;
wire _3089_;
wire _3090_;
wire _3091_;
wire _3092_;
wire _3093_;
wire _3094_;
wire _3095_;
wire _3096_;
wire _3097_;
wire _3098_;
wire _3099_;
wire _3100_;
wire _3101_;
wire _3102_;
wire _3103_;
wire _3104_;
wire _3105_;
wire _3106_;
wire _3107_;
wire _3108_;
wire _3109_;
wire _3110_;
wire _3111_;
wire _3112_;
wire _3113_;
wire _3114_;
wire _3115_;
wire _3116_;
wire _3117_;
wire _3118_;
wire _3119_;
wire _3120_;
wire _3121_;
wire _3122_;
wire _3123_;
wire _3124_;
wire _3125_;
wire _3126_;
wire _3127_;
wire _3128_;
wire _3129_;
wire _3130_;
wire _3131_;
wire _3132_;
wire _3133_;
wire _3134_;
wire _3135_;
wire _3136_;
wire _3137_;
wire _3138_;
wire _3139_;
wire _3140_;
wire _3141_;
wire _3142_;
wire _3143_;
wire _3144_;
wire _3145_;
wire _3146_;
wire _3147_;
wire _3148_;
wire _3149_;
wire _3150_;
wire _3151_;
wire _3152_;
wire _3153_;
wire _3154_;
wire _3155_;
wire _3156_;
wire _3157_;
wire _3158_;
wire _3159_;
wire _3160_;
wire _3161_;
wire _3162_;
wire _3163_;
wire _3164_;
wire _3165_;
wire _3166_;
wire _3167_;
wire _3168_;
wire _3169_;
wire _3170_;
wire _3171_;
wire _3172_;
wire _3173_;
wire _3174_;
wire _3175_;
wire _3176_;
wire _3177_;
wire _3178_;
wire _3179_;
wire _3180_;
wire _3181_;
wire _3182_;
wire _3183_;
wire _3184_;
wire _3185_;
wire _3186_;
wire _3187_;
wire _3188_;
wire _3189_;
wire _3190_;
wire _3191_;
wire _3192_;
wire _3193_;
wire _3194_;
wire _3195_;
wire _3196_;
wire _3197_;
wire _3198_;
wire _3199_;
wire _3200_;
wire _3201_;
wire _3202_;
wire _3203_;
wire _3204_;
wire _3205_;
wire _3206_;
wire _3207_;
wire _3208_;
wire _3209_;
wire _3210_;
wire _3211_;
wire _3212_;
wire _3213_;
wire _3214_;
wire _3215_;
wire _3216_;
wire _3217_;
wire _3218_;
wire _3219_;
wire _3220_;
wire _3221_;
wire _3222_;
wire _3223_;
wire _3224_;
wire _3225_;
wire _3226_;
wire _3227_;
wire _3228_;
wire _3229_;
wire _3230_;
wire _3231_;
wire _3232_;
wire _3233_;
wire _3234_;
wire _3235_;
wire _3236_;
wire _3237_;
wire _3238_;
wire _3239_;
wire _3240_;
wire _3241_;
wire _3242_;
wire _3243_;
wire _3244_;
wire _3245_;
wire _3246_;
wire _3247_;
wire _3248_;
wire _3249_;
wire _3250_;
wire _3251_;
wire _3252_;
wire _3253_;
wire _3254_;
wire _3255_;
wire _3256_;
wire _3257_;
wire _3258_;
wire _3259_;
wire _3260_;
wire _3261_;
wire _3262_;
wire _3263_;
wire _3264_;
wire _3265_;
wire _3266_;
wire _3267_;
wire _3268_;
wire _3269_;
wire _3270_;
wire _3271_;
wire _3272_;
wire _3273_;
wire _3274_;
wire _3275_;
wire _3276_;
wire _3277_;
wire _3278_;
wire _3279_;
wire _3280_;
wire _3281_;
wire _3282_;
wire _3283_;
wire _3284_;
wire _3285_;
wire _3286_;
wire _3287_;
wire _3288_;
wire _3289_;
wire _3290_;
wire _3291_;
wire _3292_;
wire _3293_;
wire _3294_;
wire _3295_;
wire _3296_;
wire _3297_;
wire _3298_;
wire _3299_;
wire _3300_;
wire _3301_;
wire _3302_;
wire _3303_;
wire _3304_;
wire _3305_;
wire _3306_;
wire _3307_;
wire _3308_;
wire _3309_;
wire _3310_;
wire _3311_;
wire _3312_;
wire _3313_;
wire _3314_;
wire _3315_;
wire _3316_;
wire _3317_;
wire _3318_;
wire _3319_;
wire _3320_;
wire _3321_;
wire _3322_;
wire _3323_;
wire _3324_;
wire _3325_;
wire _3326_;
wire _3327_;
wire _3328_;
wire _3329_;
wire _3330_;
wire _3331_;
wire _3332_;
wire _3333_;
wire _3334_;
wire _3335_;
wire _3336_;
wire _3337_;
wire _3338_;
wire _3339_;
wire _3340_;
wire _3341_;
wire _3342_;
wire _3343_;
wire _3344_;
wire _3345_;
wire _3346_;
wire _3347_;
wire _3348_;
wire _3349_;
wire _3350_;
wire _3351_;
wire _3352_;
wire _3353_;
wire _3354_;
wire _3355_;
wire _3356_;
wire _3357_;
wire _3358_;
wire _3359_;
wire _3360_;
wire _3361_;
wire _3362_;
wire _3363_;
wire _3364_;
wire _3365_;
wire _3366_;
wire _3367_;
wire _3368_;
wire _3369_;
wire _3370_;
wire _3371_;
wire _3372_;
wire _3373_;
wire _3374_;
wire _3375_;
wire _3376_;
wire _3377_;
wire _3378_;
wire _3379_;
wire _3380_;
wire _3381_;
wire _3382_;
wire _3383_;
wire _3384_;
wire _3385_;
wire _3386_;
wire _3387_;
wire _3388_;
wire _3389_;
wire _3390_;
wire _3391_;
wire _3392_;
wire _3393_;
wire _3394_;
wire _3395_;
wire _3396_;
wire _3397_;
wire _3398_;
wire _3399_;
wire _3400_;
wire _3401_;
wire _3402_;
wire _3403_;
wire _3404_;
wire _3405_;
wire _3406_;
wire _3407_;
wire _3408_;
wire _3409_;
wire _3410_;
wire _3411_;
wire _3412_;
wire _3413_;
wire _3414_;
wire _3415_;
wire _3416_;
wire _3417_;
wire _3418_;
wire _3419_;
wire _3420_;
wire _3421_;
wire _3422_;
wire _3423_;
wire _3424_;
wire _3425_;
wire _3426_;
wire _3427_;
wire _3428_;
wire _3429_;
wire _3430_;
wire _3431_;
wire _3432_;
wire _3433_;
wire _3434_;
wire _3435_;
wire _3436_;
wire _3437_;
wire _3438_;
wire _3439_;
wire _3440_;
wire _3441_;
wire _3442_;
wire _3443_;
wire _3444_;
wire _3445_;
wire _3446_;
wire _3447_;
wire _3448_;
wire _3449_;
wire _3450_;
wire _3451_;
wire _3452_;
wire _3453_;
wire _3454_;
wire _3455_;
wire _3456_;
wire _3457_;
wire _3458_;
wire _3459_;
wire _3460_;
wire _3461_;
wire _3462_;
wire _3463_;
wire _3464_;
wire _3465_;
wire _3466_;
wire _3467_;
wire _3468_;
wire _3469_;
wire _3470_;
wire _3471_;
wire _3472_;
wire _3473_;
wire _3474_;
wire _3475_;
wire _3476_;
wire _3477_;
wire _3478_;
wire _3479_;
wire _3480_;
wire _3481_;
wire _3482_;
wire _3483_;
wire _3484_;
wire _3485_;
wire _3486_;
wire _3487_;
wire _3488_;
wire _3489_;
wire _3490_;
wire _3491_;
wire _3492_;
wire _3493_;
wire _3494_;
wire _3495_;
wire _3496_;
wire _3497_;
wire _3498_;
wire _3499_;
wire _3500_;
wire _3501_;
wire _3502_;
wire _3503_;
wire _3504_;
wire _3505_;
wire _3506_;
wire _3507_;
wire _3508_;
wire _3509_;
wire _3510_;
wire _3511_;
wire _3512_;
wire _3513_;
wire _3514_;
wire _3515_;
wire _3516_;
wire _3517_;
wire _3518_;
wire _3519_;
wire _3520_;
wire _3521_;
wire _3522_;
wire _3523_;
wire _3524_;
wire _3525_;
wire _3526_;
wire _3527_;
wire _3528_;
wire _3529_;
wire _3530_;
wire _3531_;
wire _3532_;
wire _3533_;
wire _3534_;
wire _3535_;
wire _3536_;
wire _3537_;
wire _3538_;
wire _3539_;
wire _3540_;
wire _3541_;
wire _3542_;
wire _3543_;
wire _3544_;
wire _3545_;
wire _3546_;
wire _3547_;
wire _3548_;
wire _3549_;
wire _3550_;
wire _3551_;
wire _3552_;
wire _3553_;
wire _3554_;
wire _3555_;
wire _3556_;
wire _3557_;
wire _3558_;
wire _3559_;
wire _3560_;
wire _3561_;
wire _3562_;
wire _3563_;
wire _3564_;
wire _3565_;
wire _3566_;
wire _3567_;
wire _3568_;
wire _3569_;
wire _3570_;
wire _3571_;
wire _3572_;
wire _3573_;
wire _3574_;
wire _3575_;
wire _3576_;
wire _3577_;
wire _3578_;
wire _3579_;
wire _3580_;
wire _3581_;
wire _3582_;
wire _3583_;
wire _3584_;
wire _3585_;
wire _3586_;
wire _3587_;
wire _3588_;
wire _3589_;
wire _3590_;
wire _3591_;
wire _3592_;
wire _3593_;
wire _3594_;
wire _3595_;
wire _3596_;
wire _3597_;
wire _3598_;
wire _3599_;
wire _3600_;
wire _3601_;
wire _3602_;
wire _3603_;
wire _3604_;
wire _3605_;
wire _3606_;
wire _3607_;
wire _3608_;
wire _3609_;
wire _3610_;
wire _3611_;
wire _3612_;
wire _3613_;
wire _3614_;
wire _3615_;
wire _3616_;
wire _3617_;
wire _3618_;
wire _3619_;
wire _3620_;
wire _3621_;
wire _3622_;
wire _3623_;
wire _3624_;
wire _3625_;
wire _3626_;
wire _3627_;
wire _3628_;
wire _3629_;
wire _3630_;
wire _3631_;
wire _3632_;
wire _3633_;
wire _3634_;
wire _3635_;
wire _3636_;
wire _3637_;
wire _3638_;
wire _3639_;
wire _3640_;
wire _3641_;
wire _3642_;
wire _3643_;
wire _3644_;
wire _3645_;
wire _3646_;
wire _3647_;
wire _3648_;
wire _3649_;
wire _3650_;
wire _3651_;
wire _3652_;
wire _3653_;
wire _3654_;
wire _3655_;
wire _3656_;
wire _3657_;
wire _3658_;
wire _3659_;
wire _3660_;
wire _3661_;
wire _3662_;
wire _3663_;
wire _3664_;
wire _3665_;
wire _3666_;
wire _3667_;
wire _3668_;
wire _3669_;
wire _3670_;
wire _3671_;
wire _3672_;
wire _3673_;
wire _3674_;
wire _3675_;
wire _3676_;
wire _3677_;
wire _3678_;
wire _3679_;
wire _3680_;
wire _3681_;
wire _3682_;
wire _3683_;
wire _3684_;
wire _3685_;
wire _3686_;
wire _3687_;
wire _3688_;
wire _3689_;
wire _3690_;
wire _3691_;
wire _3692_;
wire _3693_;
wire _3694_;
wire _3695_;
wire _3696_;
wire _3697_;
wire _3698_;
wire _3699_;
wire _3700_;
wire _3701_;
wire _3702_;
wire _3703_;
wire _3704_;
wire _3705_;
wire _3706_;
wire _3707_;
wire _3708_;
wire _3709_;
wire _3710_;
wire _3711_;
wire _3712_;
wire _3713_;
wire _3714_;
wire _3715_;
wire _3716_;
wire _3717_;
wire _3718_;
wire _3719_;
wire _3720_;
wire _3721_;
wire _3722_;
wire _3723_;
wire _3724_;
wire _3725_;
wire _3726_;
wire _3727_;
wire _3728_;
wire _3729_;
wire _3730_;
wire _3731_;
wire _3732_;
wire _3733_;
wire _3734_;
wire _3735_;
wire _3736_;
wire _3737_;
wire _3738_;
wire _3739_;
wire _3740_;
wire _3741_;
wire _3742_;
wire _3743_;
wire _3744_;
wire _3745_;
wire _3746_;
wire _3747_;
wire _3748_;
wire _3749_;
wire _3750_;
wire _3751_;
wire _3752_;
wire _3753_;
wire _3754_;
wire _3755_;
wire _3756_;
wire _3757_;
wire _3758_;
wire _3759_;
wire _3760_;
wire _3761_;
wire _3762_;
wire _3763_;
wire _3764_;
wire _3765_;
wire _3766_;
wire _3767_;
wire _3768_;
wire _3769_;
wire _3770_;
wire _3771_;
wire _3772_;
wire _3773_;
wire _3774_;
wire _3775_;
wire _3776_;
wire _3777_;
wire _3778_;
wire _3779_;
wire _3780_;
wire _3781_;
wire _3782_;
wire _3783_;
wire _3784_;
wire _3785_;
wire _3786_;
wire _3787_;
wire _3788_;
wire _3789_;
wire _3790_;
wire _3791_;
wire _3792_;
wire _3793_;
wire _3794_;
wire _3795_;
wire _3796_;
wire _3797_;
wire _3798_;
wire _3799_;
wire _3800_;
wire _3801_;
wire _3802_;
wire _3803_;
wire _3804_;
wire _3805_;
wire _3806_;
wire _3807_;
wire _3808_;
wire _3809_;
wire _3810_;
wire _3811_;
wire _3812_;
wire _3813_;
wire _3814_;
wire _3815_;
wire _3816_;
wire _3817_;
wire _3818_;
wire _3819_;
wire _3820_;
wire _3821_;
wire _3822_;
wire _3823_;
wire _3824_;
wire _3825_;
wire _3826_;
wire _3827_;
wire _3828_;
wire _3829_;
wire _3830_;
wire _3831_;
wire _3832_;
wire _3833_;
wire _3834_;
wire _3835_;
wire _3836_;
wire _3837_;
wire _3838_;
wire _3839_;
wire _3840_;
wire _3841_;
wire _3842_;
wire _3843_;
wire _3844_;
wire _3845_;
wire _3846_;
wire _3847_;
wire _3848_;
wire _3849_;
wire _3850_;
wire _3851_;
wire _3852_;
wire _3853_;
wire _3854_;
wire _3855_;
wire _3856_;
wire _3857_;
wire _3858_;
wire _3859_;
wire _3860_;
wire _3861_;
wire _3862_;
wire _3863_;
wire _3864_;
wire _3865_;
wire _3866_;
wire _3867_;
wire _3868_;
wire _3869_;
wire _3870_;
wire _3871_;
wire _3872_;
wire _3873_;
wire _3874_;
wire _3875_;
wire _3876_;
wire _3877_;
wire _3878_;
wire _3879_;
wire _3880_;
wire _3881_;
wire _3882_;
wire _3883_;
wire _3884_;
wire _3885_;
wire _3886_;
wire _3887_;
wire _3888_;
wire _3889_;
wire _3890_;
wire _3891_;
wire _3892_;
wire _3893_;
wire _3894_;
wire _3895_;
wire _3896_;
wire _3897_;
wire _3898_;
wire _3899_;
wire _3900_;
wire _3901_;
wire _3902_;
wire _3903_;
wire _3904_;
wire _3905_;
wire _3906_;
wire _3907_;
wire _3908_;
wire _3909_;
wire _3910_;
wire _3911_;
wire _3912_;
wire _3913_;
wire _3914_;
wire _3915_;
wire _3916_;
wire _3917_;
wire _3918_;
wire _3919_;
wire _3920_;
wire _3921_;
wire _3922_;
wire _3923_;
wire _3924_;
wire _3925_;
wire _3926_;
wire _3927_;
wire _3928_;
wire _3929_;
wire _3930_;
wire _3931_;
wire _3932_;
wire _3933_;
wire _3934_;
wire _3935_;
wire _3936_;
wire _3937_;
wire _3938_;
wire _3939_;
wire _3940_;
wire _3941_;
wire _3942_;
wire _3943_;
wire _3944_;
wire _3945_;
wire _3946_;
wire _3947_;
wire _3948_;
wire _3949_;
wire _3950_;
wire _3951_;
wire _3952_;
wire _3953_;
wire _3954_;
wire _3955_;
wire _3956_;
wire _3957_;
wire _3958_;
wire _3959_;
wire _3960_;
wire _3961_;
wire _3962_;
wire _3963_;
wire _3964_;
wire _3965_;
wire _3966_;
wire _3967_;
wire _3968_;
wire _3969_;
wire _3970_;
wire _3971_;
wire _3972_;
wire _3973_;
wire _3974_;
wire _3975_;
wire _3976_;
wire _3977_;
wire _3978_;
wire _3979_;
wire _3980_;
wire _3981_;
wire _3982_;
wire _3983_;
wire _3984_;
wire _3985_;
wire _3986_;
wire _3987_;
wire _3988_;
wire _3989_;
wire _3990_;
wire _3991_;
wire _3992_;
wire _3993_;
wire _3994_;
wire _3995_;
wire _3996_;
wire _3997_;
wire _3998_;
wire _3999_;
wire _4000_;
wire _4001_;
wire _4002_;
wire _4003_;
wire _4004_;
wire _4005_;
wire _4006_;
wire _4007_;
wire _4008_;
wire _4009_;
wire _4010_;
wire _4011_;
wire _4012_;
wire _4013_;
wire _4014_;
wire _4015_;
wire _4016_;
wire _4017_;
wire _4018_;
wire _4019_;
wire _4020_;
wire _4021_;
wire _4022_;
wire _4023_;
wire _4024_;
wire _4025_;
wire _4026_;
wire _4027_;
wire _4028_;
wire _4029_;
wire _4030_;
wire _4031_;
wire _4032_;
wire _4033_;
wire _4034_;
wire _4035_;
wire _4036_;
wire _4037_;
wire _4038_;
wire _4039_;
wire _4040_;
wire _4041_;
wire _4042_;
wire _4043_;
wire _4044_;
wire _4045_;
wire _4046_;
wire _4047_;
wire _4048_;
wire _4049_;
wire _4050_;
wire _4051_;
wire _4052_;
wire _4053_;
wire _4054_;
wire _4055_;
wire _4056_;
wire _4057_;
wire _4058_;
wire _4059_;
wire _4060_;
wire _4061_;
wire _4062_;
wire _4063_;
wire _4064_;
wire _4065_;
wire _4066_;
wire _4067_;
wire _4068_;
wire _4069_;
wire _4070_;
wire _4071_;
wire _4072_;
wire _4073_;
wire _4074_;
wire _4075_;
wire _4076_;
wire _4077_;
wire _4078_;
wire _4079_;
wire _4080_;
wire _4081_;
wire _4082_;
wire _4083_;
wire _4084_;
wire _4085_;
wire _4086_;
wire _4087_;
wire _4088_;
wire _4089_;
wire _4090_;
wire _4091_;
wire _4092_;
wire _4093_;
wire _4094_;
wire _4095_;
wire _4096_;
wire _4097_;
wire _4098_;
wire _4099_;
wire _4100_;
wire _4101_;
wire _4102_;
wire _4103_;
wire _4104_;
wire _4105_;
wire _4106_;
wire _4107_;
wire _4108_;
wire _4109_;
wire _4110_;
wire _4111_;
wire _4112_;
wire _4113_;
wire _4114_;
wire _4115_;
wire _4116_;
wire _4117_;
wire _4118_;
wire _4119_;
wire _4120_;
wire _4121_;
wire _4122_;
wire _4123_;
wire _4124_;
wire _4125_;
wire _4126_;
wire _4127_;
wire _4128_;
wire _4129_;
wire _4130_;
wire _4131_;
wire _4132_;
wire _4133_;
wire _4134_;
wire _4135_;
wire _4136_;
wire _4137_;
wire _4138_;
wire _4139_;
wire _4140_;
wire _4141_;
wire _4142_;
wire _4143_;
wire _4144_;
wire _4145_;
wire _4146_;
wire _4147_;
wire _4148_;
wire _4149_;
wire _4150_;
wire _4151_;
wire _4152_;
wire _4153_;
wire _4154_;
wire _4155_;
wire _4156_;
wire _4157_;
wire _4158_;
wire _4159_;
wire _4160_;
wire _4161_;
wire _4162_;
wire _4163_;
wire _4164_;
wire _4165_;
wire _4166_;
wire _4167_;
wire _4168_;
wire _4169_;
wire _4170_;
wire _4171_;
wire _4172_;
wire _4173_;
wire _4174_;
wire _4175_;
wire _4176_;
wire _4177_;
wire _4178_;
wire _4179_;
wire _4180_;
wire _4181_;
wire _4182_;
wire _4183_;
wire _4184_;
wire _4185_;
wire _4186_;
wire _4187_;
wire _4188_;
wire _4189_;
wire _4190_;
wire _4191_;
wire _4192_;
wire _4193_;
wire _4194_;
wire _4195_;
wire _4196_;
wire _4197_;
wire _4198_;
wire _4199_;
wire _4200_;
wire _4201_;
wire _4202_;
wire _4203_;
wire _4204_;
wire _4205_;
wire _4206_;
wire _4207_;
wire _4208_;
wire _4209_;
wire _4210_;
wire _4211_;
wire _4212_;
wire _4213_;
wire _4214_;
wire _4215_;
wire _4216_;
wire _4217_;
wire _4218_;
wire _4219_;
wire _4220_;
wire _4221_;
wire _4222_;
wire _4223_;
wire _4224_;
wire _4225_;
wire _4226_;
wire _4227_;
wire _4228_;
wire _4229_;
wire _4230_;
wire _4231_;
wire _4232_;
wire _4233_;
wire _4234_;
wire _4235_;
wire _4236_;
wire _4237_;
wire _4238_;
wire _4239_;
wire _4240_;
wire _4241_;
wire _4242_;
wire _4243_;
wire _4244_;
wire _4245_;
wire _4246_;
wire _4247_;
wire _4248_;
wire _4249_;
wire _4250_;
wire _4251_;
wire _4252_;
wire _4253_;
wire _4254_;
wire _4255_;
wire _4256_;
wire _4257_;
wire _4258_;
wire _4259_;
wire _4260_;
wire _4261_;
wire _4262_;
wire _4263_;
wire _4264_;
wire _4265_;
wire _4266_;
wire _4267_;
wire _4268_;
wire _4269_;
wire _4270_;
wire _4271_;
wire _4272_;
wire _4273_;
wire _4274_;
wire _4275_;
wire _4276_;
wire _4277_;
wire _4278_;
wire _4279_;
wire _4280_;
wire _4281_;
wire _4282_;
wire _4283_;
wire _4284_;
wire _4285_;
wire _4286_;
wire _4287_;
wire _4288_;
wire _4289_;
wire _4290_;
wire _4291_;
wire _4292_;
wire _4293_;
wire _4294_;
wire _4295_;
wire _4296_;
wire _4297_;
wire _4298_;
wire _4299_;
wire _4300_;
wire _4301_;
wire _4302_;
wire _4303_;
wire _4304_;
wire _4305_;
wire _4306_;
wire _4307_;
wire _4308_;
wire _4309_;
wire _4310_;
wire _4311_;
wire _4312_;
wire _4313_;
wire _4314_;
wire _4315_;
wire _4316_;
wire _4317_;
wire _4318_;
wire _4319_;
wire _4320_;
wire _4321_;
wire _4322_;
wire _4323_;
wire _4324_;
wire _4325_;
wire _4326_;
wire _4327_;
wire _4328_;
wire _4329_;
wire _4330_;
wire _4331_;
wire _4332_;
wire _4333_;
wire _4334_;
wire _4335_;
wire _4336_;
wire _4337_;
wire _4338_;
wire _4339_;
wire _4340_;
wire _4341_;
wire _4342_;
wire _4343_;
wire _4344_;
wire _4345_;
wire _4346_;
wire _4347_;
wire _4348_;
wire _4349_;
wire _4350_;
wire _4351_;
wire _4352_;
wire _4353_;
wire _4354_;
wire _4355_;
wire _4356_;
wire _4357_;
wire _4358_;
wire _4359_;
wire _4360_;
wire _4361_;
wire _4362_;
wire _4363_;
wire _4364_;
wire _4365_;
wire _4366_;
wire _4367_;
wire _4368_;
wire _4369_;
wire _4370_;
wire _4371_;
wire _4372_;
wire _4373_;
wire _4374_;
wire _4375_;
wire _4376_;
wire _4377_;
wire _4378_;
wire _4379_;
wire _4380_;
wire _4381_;
wire _4382_;
wire _4383_;
wire _4384_;
wire _4385_;
wire _4386_;
wire _4387_;
wire _4388_;
wire _4389_;
wire _4390_;
wire _4391_;
wire _4392_;
wire _4393_;
wire _4394_;
wire _4395_;
wire _4396_;
wire _4397_;
wire _4398_;
wire _4399_;
wire _4400_;
wire _4401_;
wire _4402_;
wire _4403_;
wire _4404_;
wire _4405_;
wire _4406_;
wire _4407_;
wire _4408_;
wire _4409_;
wire _4410_;
wire _4411_;
wire _4412_;
wire _4413_;
wire _4414_;
wire _4415_;
wire _4416_;
wire _4417_;
wire _4418_;
wire _4419_;
wire _4420_;
wire _4421_;
wire _4422_;
wire _4423_;
wire _4424_;
wire _4425_;
wire _4426_;
wire _4427_;
wire _4428_;
wire _4429_;
wire _4430_;
wire _4431_;
wire _4432_;
wire _4433_;
wire _4434_;
wire _4435_;
wire _4436_;
wire _4437_;
wire _4438_;
wire _4439_;
wire _4440_;
wire _4441_;
wire _4442_;
wire _4443_;
wire _4444_;
wire _4445_;
wire _4446_;
wire _4447_;
wire _4448_;
wire _4449_;
wire _4450_;
wire _4451_;
wire _4452_;
wire _4453_;
wire _4454_;
wire _4455_;
wire _4456_;
wire _4457_;
wire _4458_;
wire _4459_;
wire _4460_;
wire _4461_;
wire _4462_;
wire _4463_;
wire _4464_;
wire _4465_;
wire _4466_;
wire _4467_;
wire _4468_;
wire _4469_;
wire _4470_;
wire _4471_;
wire _4472_;
wire _4473_;
wire _4474_;
wire _4475_;
wire _4476_;
wire _4477_;
wire _4478_;
wire _4479_;
wire _4480_;
wire _4481_;
wire _4482_;
wire _4483_;
wire _4484_;
wire _4485_;
wire _4486_;
wire _4487_;
wire _4488_;
wire _4489_;
wire _4490_;
wire _4491_;
wire _4492_;
wire _4493_;
wire _4494_;
wire _4495_;
wire _4496_;
wire _4497_;
wire _4498_;
wire _4499_;
wire _4500_;
wire _4501_;
wire _4502_;
wire _4503_;
wire _4504_;
wire _4505_;
wire _4506_;
wire _4507_;
wire _4508_;
wire _4509_;
wire _4510_;
wire _4511_;
wire _4512_;
wire _4513_;
wire _4514_;
wire _4515_;
wire _4516_;
wire _4517_;
wire _4518_;
wire _4519_;
wire _4520_;
wire _4521_;
wire _4522_;
wire _4523_;
wire _4524_;
wire _4525_;
wire _4526_;
wire _4527_;
wire _4528_;
wire _4529_;
wire _4530_;
wire _4531_;
wire _4532_;
wire _4533_;
wire _4534_;
wire _4535_;
wire _4536_;
wire _4537_;
wire _4538_;
wire _4539_;
wire _4540_;
wire _4541_;
wire _4542_;
wire _4543_;
wire _4544_;
wire _4545_;
wire _4546_;
wire _4547_;
wire _4548_;
wire _4549_;
wire _4550_;
wire _4551_;
wire _4552_;
wire _4553_;
wire _4554_;
wire _4555_;
wire _4556_;
wire _4557_;
wire _4558_;
wire _4559_;
wire _4560_;
wire _4561_;
wire _4562_;
wire _4563_;
wire _4564_;
wire _4565_;
wire _4566_;
wire _4567_;
wire _4568_;
wire _4569_;
wire _4570_;
wire _4571_;
wire _4572_;
wire _4573_;
wire _4574_;
wire _4575_;
wire _4576_;
wire _4577_;
wire _4578_;
wire _4579_;
wire _4580_;
wire _4581_;
wire _4582_;
wire _4583_;
wire _4584_;
wire _4585_;
wire _4586_;
wire _4587_;
wire _4588_;
wire _4589_;
wire _4590_;
wire _4591_;
wire _4592_;
wire _4593_;
wire _4594_;
wire _4595_;
wire _4596_;
wire _4597_;
wire _4598_;
wire _4599_;
wire _4600_;
wire _4601_;
wire _4602_;
wire _4603_;
wire _4604_;
wire _4605_;
wire _4606_;
wire _4607_;
wire _4608_;
wire _4609_;
wire _4610_;
wire _4611_;
wire _4612_;
wire _4613_;
wire _4614_;
wire _4615_;
wire _4616_;
wire _4617_;
wire _4618_;
wire _4619_;
wire _4620_;
wire _4621_;
wire _4622_;
wire _4623_;
wire _4624_;
wire _4625_;
wire _4626_;
wire _4627_;
wire _4628_;
wire _4629_;
wire _4630_;
wire _4631_;
wire _4632_;
wire _4633_;
wire _4634_;
wire _4635_;
wire _4636_;
wire _4637_;
wire _4638_;
wire _4639_;
wire _4640_;
wire _4641_;
wire _4642_;
wire _4643_;
wire _4644_;
wire _4645_;
wire _4646_;
wire _4647_;
wire _4648_;
wire _4649_;
wire _4650_;
wire _4651_;
wire _4652_;
wire _4653_;
wire _4654_;
wire _4655_;
wire _4656_;
wire _4657_;
wire _4658_;
wire _4659_;
wire _4660_;
wire _4661_;
wire _4662_;
wire _4663_;
wire _4664_;
wire _4665_;
wire _4666_;
wire _4667_;
wire _4668_;
wire _4669_;
wire _4670_;
wire _4671_;
wire _4672_;
wire _4673_;
wire _4674_;
wire _4675_;
wire _4676_;
wire _4677_;
wire _4678_;
wire _4679_;
wire _4680_;
wire _4681_;
wire _4682_;
wire _4683_;
wire _4684_;
wire _4685_;
wire _4686_;
wire _4687_;
wire _4688_;
wire _4689_;
wire _4690_;
wire _4691_;
wire _4692_;
wire _4693_;
wire _4694_;
wire _4695_;
wire _4696_;
wire _4697_;
wire _4698_;
wire _4699_;
wire _4700_;
wire _4701_;
wire _4702_;
wire _4703_;
wire _4704_;
wire _4705_;
wire _4706_;
wire _4707_;
wire _4708_;
wire _4709_;
wire _4710_;
wire _4711_;
wire _4712_;
wire _4713_;
wire _4714_;
wire _4715_;
wire _4716_;
wire _4717_;
wire _4718_;
wire _4719_;
wire _4720_;
wire _4721_;
wire _4722_;
wire _4723_;
wire _4724_;
wire _4725_;
wire _4726_;
wire _4727_;
wire _4728_;
wire _4729_;
wire _4730_;
wire _4731_;
wire _4732_;
wire _4733_;
wire _4734_;
wire _4735_;
wire _4736_;
wire _4737_;
wire _4738_;
wire _4739_;
wire _4740_;
wire _4741_;
wire _4742_;
wire _4743_;
wire _4744_;
wire _4745_;
wire _4746_;
wire _4747_;
wire _4748_;
wire _4749_;
wire _4750_;
wire _4751_;
wire _4752_;
wire _4753_;
wire _4754_;
wire _4755_;
wire _4756_;
wire _4757_;
wire _4758_;
wire _4759_;
wire _4760_;
wire _4761_;
wire _4762_;
wire _4763_;
wire _4764_;
wire _4765_;
wire _4766_;
wire _4767_;
wire _4768_;
wire _4769_;
wire _4770_;
wire _4771_;
wire _4772_;
wire _4773_;
wire _4774_;
wire _4775_;
wire _4776_;
wire _4777_;
wire _4778_;
wire _4779_;
wire _4780_;
wire _4781_;
wire _4782_;
wire _4783_;
wire _4784_;
wire _4785_;
wire _4786_;
wire _4787_;
wire _4788_;
wire _4789_;
wire _4790_;
wire _4791_;
wire _4792_;
wire _4793_;
wire _4794_;
wire _4795_;
wire _4796_;
wire _4797_;
wire _4798_;
wire _4799_;
wire _4800_;
wire _4801_;
wire _4802_;
wire _4803_;
wire _4804_;
wire _4805_;
wire _4806_;
wire _4807_;
wire _4808_;
wire _4809_;
wire _4810_;
wire _4811_;
wire _4812_;
wire _4813_;
wire _4814_;
wire _4815_;
wire _4816_;
wire _4817_;
wire _4818_;
wire _4819_;
wire _4820_;
wire _4821_;
wire _4822_;
wire _4823_;
wire _4824_;
wire _4825_;
wire _4826_;
wire _4827_;
wire _4828_;
wire _4829_;
wire _4830_;
wire _4831_;
wire _4832_;
wire _4833_;
wire _4834_;
wire _4835_;
wire _4836_;
wire _4837_;
wire _4838_;
wire _4839_;
wire _4840_;
wire _4841_;
wire _4842_;
wire _4843_;
wire _4844_;
wire _4845_;
wire _4846_;
wire _4847_;
wire _4848_;
wire _4849_;
wire _4850_;
wire _4851_;
wire _4852_;
wire _4853_;
wire _4854_;
wire _4855_;
wire _4856_;
wire _4857_;
wire _4858_;
wire _4859_;
wire _4860_;
wire _4861_;
wire _4862_;
wire _4863_;
wire _4864_;
wire _4865_;
wire _4866_;
wire _4867_;
wire _4868_;
wire _4869_;
wire _4870_;
wire _4871_;
wire _4872_;
wire _4873_;
wire _4874_;
wire _4875_;
wire _4876_;
wire _4877_;
wire _4878_;
wire _4879_;
wire _4880_;
wire _4881_;
wire _4882_;
wire _4883_;
wire _4884_;
wire _4885_;
wire _4886_;
wire _4887_;
wire _4888_;
wire _4889_;
wire _4890_;
wire _4891_;
wire _4892_;
wire _4893_;
wire _4894_;
wire _4895_;
wire _4896_;
wire _4897_;
wire _4898_;
wire _4899_;
wire _4900_;
wire _4901_;
wire _4902_;
wire _4903_;
wire _4904_;
wire _4905_;
wire _4906_;
wire _4907_;
wire _4908_;
wire _4909_;
wire _4910_;
wire _4911_;
wire _4912_;
wire _4913_;
wire _4914_;
wire _4915_;
wire _4916_;
wire _4917_;
wire _4918_;
wire _4919_;
wire _4920_;
wire _4921_;
wire _4922_;
wire _4923_;
wire _4924_;
wire _4925_;
wire _4926_;
wire _4927_;
wire _4928_;
wire _4929_;
wire _4930_;
wire _4931_;
wire _4932_;
wire _4933_;
wire _4934_;
wire _4935_;
wire _4936_;
wire _4937_;
wire _4938_;
wire _4939_;
wire _4940_;
wire _4941_;
wire _4942_;
wire _4943_;
wire _4944_;
wire _4945_;
wire _4946_;
wire _4947_;
wire _4948_;
wire _4949_;
wire _4950_;
wire _4951_;
wire _4952_;
wire _4953_;
wire _4954_;
wire _4955_;
wire _4956_;
wire _4957_;
wire _4958_;
wire _4959_;
wire _4960_;
wire _4961_;
wire _4962_;
wire _4963_;
wire _4964_;
wire _4965_;
wire _4966_;
wire _4967_;
wire _4968_;
wire _4969_;
wire _4970_;
wire _4971_;
wire _4972_;
wire _4973_;
wire _4974_;
wire _4975_;
wire _4976_;
wire _4977_;
wire _4978_;
wire _4979_;
wire _4980_;
wire _4981_;
wire _4982_;
wire _4983_;
wire _4984_;
wire _4985_;
wire _4986_;
wire _4987_;
wire _4988_;
wire _4989_;
wire _4990_;
wire _4991_;
wire _4992_;
wire _4993_;
wire _4994_;
wire _4995_;
wire _4996_;
wire _4997_;
wire _4998_;
wire _4999_;
wire _5000_;
wire _5001_;
wire _5002_;
wire _5003_;
wire _5004_;
wire _5005_;
wire _5006_;
wire _5007_;
wire _5008_;
wire _5009_;
wire _5010_;
wire _5011_;
wire _5012_;
wire _5013_;
wire _5014_;
wire _5015_;
wire _5016_;
wire _5017_;
wire _5018_;
wire _5019_;
wire _5020_;
wire _5021_;
wire _5022_;
wire _5023_;
wire _5024_;
wire _5025_;
wire _5026_;
wire _5027_;
wire _5028_;
wire _5029_;
wire _5030_;
wire _5031_;
wire _5032_;
wire _5033_;
wire _5034_;
wire _5035_;
wire _5036_;
wire _5037_;
wire _5038_;
wire _5039_;
wire _5040_;
wire _5041_;
wire _5042_;
wire _5043_;
wire _5044_;
wire _5045_;
wire _5046_;
wire _5047_;
wire _5048_;
wire _5049_;
wire _5050_;
wire _5051_;
wire _5052_;
wire _5053_;
wire _5054_;
wire _5055_;
wire _5056_;
wire _5057_;
wire _5058_;
wire _5059_;
wire _5060_;
wire _5061_;
wire _5062_;
wire _5063_;
wire _5064_;
wire _5065_;
wire _5066_;
wire _5067_;
wire _5068_;
wire _5069_;
wire _5070_;
wire _5071_;
wire _5072_;
wire _5073_;
wire _5074_;
wire _5075_;
wire _5076_;
wire _5077_;
wire _5078_;
wire _5079_;
wire _5080_;
wire _5081_;
wire _5082_;
wire _5083_;
wire _5084_;
wire _5085_;
wire _5086_;
wire _5087_;
wire _5088_;
wire _5089_;
wire _5090_;
wire _5091_;
wire _5092_;
wire _5093_;
wire _5094_;
wire _5095_;
wire _5096_;
wire _5097_;
wire _5098_;
wire _5099_;
wire _5100_;
wire _5101_;
wire _5102_;
wire _5103_;
wire _5104_;
wire _5105_;
wire _5106_;
wire _5107_;
wire _5108_;
wire _5109_;
wire _5110_;
wire _5111_;
wire _5112_;
wire _5113_;
wire _5114_;
wire _5115_;
wire _5116_;
wire _5117_;
wire _5118_;
wire _5119_;
wire _5120_;
wire _5121_;
wire _5122_;
wire _5123_;
wire _5124_;
wire _5125_;
wire _5126_;
wire _5127_;
wire _5128_;
wire _5129_;
wire _5130_;
wire _5131_;
wire _5132_;
wire _5133_;
wire _5134_;
wire _5135_;
wire _5136_;
wire _5137_;
wire _5138_;
wire _5139_;
wire _5140_;
wire _5141_;
wire _5142_;
wire _5143_;
wire _5144_;
wire _5145_;
wire _5146_;
wire _5147_;
wire _5148_;
wire _5149_;
wire _5150_;
wire _5151_;
wire _5152_;
wire _5153_;
wire _5154_;
wire _5155_;
wire _5156_;
wire _5157_;
wire _5158_;
wire _5159_;
wire _5160_;
wire _5161_;
wire _5162_;
wire _5163_;
wire _5164_;
wire _5165_;
wire _5166_;
wire _5167_;
wire _5168_;
wire _5169_;
wire _5170_;
wire _5171_;
wire _5172_;
wire _5173_;
wire _5174_;
wire _5175_;
wire _5176_;
wire _5177_;
wire _5178_;
wire _5179_;
wire _5180_;
wire _5181_;
wire _5182_;
wire _5183_;
wire _5184_;
wire _5185_;
wire _5186_;
wire _5187_;
wire _5188_;
wire _5189_;
wire _5190_;
wire _5191_;
wire _5192_;
wire _5193_;
wire _5194_;
wire _5195_;
wire _5196_;
wire _5197_;
wire _5198_;
wire _5199_;
wire _5200_;
wire _5201_;
wire _5202_;
wire _5203_;
wire _5204_;
wire _5205_;
wire _5206_;
wire _5207_;
wire _5208_;
wire _5209_;
wire _5210_;
wire _5211_;
wire _5212_;
wire _5213_;
wire _5214_;
wire _5215_;
wire _5216_;
wire _5217_;
wire _5218_;
wire _5219_;
wire _5220_;
wire _5221_;
wire _5222_;
wire _5223_;
wire _5224_;
wire _5225_;
wire _5226_;
wire _5227_;
wire _5228_;
wire _5229_;
wire _5230_;
wire _5231_;
wire _5232_;
wire _5233_;
wire _5234_;
wire _5235_;
wire _5236_;
wire _5237_;
wire _5238_;
wire _5239_;
wire _5240_;
wire _5241_;
wire _5242_;
wire _5243_;
wire _5244_;
wire _5245_;
wire _5246_;
wire _5247_;
wire _5248_;
wire _5249_;
wire _5250_;
wire _5251_;
wire _5252_;
wire _5253_;
wire _5254_;
wire _5255_;
wire _5256_;
wire _5257_;
wire _5258_;
wire _5259_;
wire _5260_;
wire _5261_;
wire _5262_;
wire _5263_;
wire _5264_;
wire _5265_;
wire _5266_;
wire _5267_;
wire _5268_;
wire _5269_;
wire _5270_;
wire _5271_;
wire _5272_;
wire _5273_;
wire _5274_;
wire _5275_;
wire _5276_;
wire _5277_;
wire _5278_;
wire _5279_;
wire _5280_;
wire _5281_;
wire _5282_;
wire _5283_;
wire _5284_;
wire _5285_;
wire _5286_;
wire _5287_;
wire _5288_;
wire _5289_;
wire _5290_;
wire _5291_;
wire _5292_;
wire _5293_;
wire _5294_;
wire _5295_;
wire _5296_;
wire _5297_;
wire _5298_;
wire _5299_;
wire _5300_;
wire _5301_;
wire _5302_;
wire _5303_;
wire _5304_;
wire _5305_;
wire _5306_;
wire _5307_;
wire _5308_;
wire _5309_;
wire _5310_;
wire _5311_;
wire _5312_;
wire _5313_;
wire _5314_;
wire _5315_;
wire _5316_;
wire _5317_;
wire _5318_;
wire _5319_;
wire _5320_;
wire _5321_;
wire _5322_;
wire _5323_;
wire _5324_;
wire _5325_;
wire _5326_;
wire _5327_;
wire _5328_;
wire _5329_;
wire _5330_;
wire _5331_;
wire _5332_;
wire _5333_;
wire _5334_;
wire _5335_;
wire _5336_;
wire _5337_;
wire _5338_;
wire _5339_;
wire _5340_;
wire _5341_;
wire _5342_;
wire _5343_;
wire _5344_;
wire _5345_;
wire _5346_;
wire _5347_;
wire _5348_;
wire _5349_;
wire _5350_;
wire _5351_;
wire _5352_;
wire _5353_;
wire _5354_;
wire _5355_;
wire _5356_;
wire _5357_;
wire _5358_;
wire _5359_;
wire _5360_;
wire _5361_;
wire _5362_;
wire _5363_;
wire _5364_;
wire _5365_;
wire _5366_;
wire _5367_;
wire _5368_;
wire _5369_;
wire _5370_;
wire _5371_;
wire _5372_;
wire _5373_;
wire _5374_;
wire _5375_;
wire _5376_;
wire _5377_;
wire _5378_;
wire _5379_;
wire _5380_;
wire _5381_;
wire _5382_;
wire _5383_;
wire _5384_;
wire _5385_;
wire _5386_;
wire _5387_;
wire _5388_;
wire _5389_;
wire _5390_;
wire _5391_;
wire _5392_;
wire _5393_;
wire _5394_;
wire _5395_;
wire _5396_;
wire _5397_;
wire _5398_;
wire _5399_;
wire _5400_;
wire _5401_;
wire _5402_;
wire _5403_;
wire _5404_;
wire _5405_;
wire _5406_;
wire _5407_;
wire _5408_;
wire _5409_;
wire _5410_;
wire _5411_;
wire _5412_;
wire _5413_;
wire _5414_;
wire _5415_;
wire _5416_;
wire _5417_;
wire _5418_;
wire _5419_;
wire _5420_;
wire _5421_;
wire _5422_;
wire _5423_;
wire _5424_;
wire _5425_;
wire _5426_;
wire _5427_;
wire _5428_;
wire _5429_;
wire _5430_;
wire _5431_;
wire _5432_;
wire _5433_;
wire _5434_;
wire _5435_;
wire _5436_;
wire _5437_;
wire _5438_;
wire _5439_;
wire _5440_;
wire _5441_;
wire _5442_;
wire _5443_;
wire _5444_;
wire _5445_;
wire _5446_;
wire _5447_;
wire _5448_;
wire _5449_;
wire _5450_;
wire _5451_;
wire _5452_;
wire _5453_;
wire _5454_;
wire _5455_;
wire _5456_;
wire _5457_;
wire _5458_;
wire _5459_;
wire _5460_;
wire _5461_;
wire _5462_;
wire _5463_;
wire _5464_;
wire _5465_;
wire _5466_;
wire _5467_;
wire _5468_;
wire _5469_;
wire _5470_;
wire _5471_;
wire _5472_;
wire _5473_;
wire _5474_;
wire _5475_;
wire _5476_;
wire _5477_;
wire _5478_;
wire _5479_;
wire _5480_;
wire _5481_;
wire _5482_;
wire _5483_;
wire _5484_;
wire _5485_;
wire _5486_;
wire _5487_;
wire _5488_;
wire _5489_;
wire _5490_;
wire _5491_;
wire _5492_;
wire _5493_;
wire _5494_;
wire _5495_;
wire _5496_;
wire _5497_;
wire _5498_;
wire _5499_;
wire _5500_;
wire _5501_;
wire _5502_;
wire _5503_;
wire _5504_;
wire _5505_;
wire _5506_;
wire _5507_;
wire _5508_;
wire _5509_;
wire _5510_;
wire _5511_;
wire _5512_;
wire _5513_;
wire _5514_;
wire _5515_;
wire _5516_;
wire _5517_;
wire _5518_;
wire _5519_;
wire _5520_;
wire _5521_;
wire _5522_;
wire _5523_;
wire _5524_;
wire _5525_;
wire _5526_;
wire _5527_;
wire _5528_;
wire _5529_;
wire _5530_;
wire _5531_;
wire _5532_;
wire _5533_;
wire _5534_;
wire _5535_;
wire _5536_;
wire _5537_;
wire _5538_;
wire _5539_;
wire _5540_;
wire _5541_;
wire _5542_;
wire _5543_;
wire _5544_;
wire _5545_;
wire _5546_;
wire _5547_;
wire _5548_;
wire _5549_;
wire _5550_;
wire _5551_;
wire _5552_;
wire _5553_;
wire _5554_;
wire _5555_;
wire _5556_;
wire _5557_;
wire _5558_;
wire _5559_;
wire _5560_;
wire _5561_;
wire _5562_;
wire _5563_;
wire _5564_;
wire _5565_;
wire _5566_;
wire _5567_;
wire _5568_;
wire _5569_;
wire _5570_;
wire _5571_;
wire _5572_;
wire _5573_;
wire _5574_;
wire _5575_;
wire _5576_;
wire _5577_;
wire _5578_;
wire _5579_;
wire _5580_;
wire _5581_;
wire _5582_;
wire _5583_;
wire _5584_;
wire _5585_;
wire _5586_;
wire _5587_;
wire _5588_;
wire _5589_;
wire _5590_;
wire _5591_;
wire _5592_;
wire _5593_;
wire _5594_;
wire _5595_;
wire _5596_;
wire _5597_;
wire _5598_;
wire _5599_;
wire _5600_;
wire _5601_;
wire _5602_;
wire _5603_;
wire _5604_;
wire _5605_;
wire _5606_;
wire _5607_;
wire _5608_;
wire _5609_;
wire _5610_;
wire _5611_;
wire _5612_;
wire _5613_;
wire _5614_;
wire _5615_;
wire _5616_;
wire _5617_;
wire _5618_;
wire _5619_;
wire _5620_;
wire _5621_;
wire _5622_;
wire _5623_;
wire _5624_;
wire _5625_;
wire _5626_;
wire _5627_;
wire _5628_;
wire _5629_;
wire _5630_;
wire _5631_;
wire _5632_;
wire _5633_;
wire _5634_;
wire _5635_;
wire _5636_;
wire _5637_;
wire _5638_;
wire _5639_;
wire _5640_;
wire _5641_;
wire _5642_;
wire _5643_;
wire _5644_;
wire _5645_;
wire _5646_;
wire _5647_;
wire _5648_;
wire _5649_;
wire _5650_;
wire _5651_;
wire _5652_;
wire _5653_;
wire _5654_;
wire _5655_;
wire _5656_;
wire _5657_;
wire _5658_;
wire _5659_;
wire _5660_;
wire _5661_;
wire _5662_;
wire _5663_;
wire _5664_;
wire _5665_;
wire _5666_;
wire _5667_;
wire _5668_;
wire _5669_;
wire _5670_;
wire _5671_;
wire _5672_;
wire _5673_;
wire _5674_;
wire _5675_;
wire _5676_;
wire _5677_;
wire _5678_;
wire _5679_;
wire _5680_;
wire _5681_;
wire _5682_;
wire _5683_;
wire _5684_;
wire _5685_;
wire _5686_;
wire _5687_;
wire _5688_;
wire _5689_;
wire _5690_;
wire _5691_;
wire _5692_;
wire _5693_;
wire _5694_;
wire _5695_;
wire _5696_;
wire _5697_;
wire _5698_;
wire _5699_;
wire _5700_;
wire _5701_;
wire _5702_;
wire _5703_;
wire _5704_;
wire _5705_;
wire _5706_;
wire _5707_;
wire _5708_;
wire _5709_;
wire _5710_;
wire _5711_;
wire _5712_;
wire _5713_;
wire _5714_;
wire _5715_;
wire _5716_;
wire _5717_;
wire _5718_;
wire _5719_;
wire _5720_;
wire _5721_;
wire _5722_;
wire _5723_;
wire _5724_;
wire _5725_;
wire _5726_;
wire _5727_;
wire _5728_;
wire _5729_;
wire _5730_;
wire _5731_;
wire _5732_;
wire _5733_;
wire _5734_;
wire _5735_;
wire _5736_;
wire _5737_;
wire _5738_;
wire _5739_;
wire _5740_;
wire _5741_;
wire _5742_;
wire _5743_;
wire _5744_;
wire _5745_;
wire _5746_;
wire _5747_;
wire _5748_;
wire _5749_;
wire _5750_;
wire _5751_;
wire _5752_;
wire _5753_;
wire _5754_;
wire _5755_;
wire _5756_;
wire _5757_;
wire _5758_;
wire _5759_;
wire _5760_;
wire _5761_;
wire _5762_;
wire _5763_;
wire _5764_;
wire _5765_;
wire _5766_;
wire _5767_;
wire _5768_;
wire _5769_;
wire _5770_;
wire _5771_;
wire _5772_;
wire _5773_;
wire _5774_;
wire _5775_;
wire _5776_;
wire _5777_;
wire _5778_;
wire _5779_;
wire _5780_;
wire _5781_;
wire _5782_;
wire _5783_;
wire _5784_;
wire _5785_;
wire _5786_;
wire _5787_;
wire _5788_;
wire _5789_;
wire _5790_;
wire _5791_;
wire _5792_;
wire _5793_;
wire _5794_;
wire _5795_;
wire _5796_;
wire _5797_;
wire _5798_;
wire _5799_;
wire _5800_;
wire _5801_;
wire _5802_;
wire _5803_;
wire _5804_;
wire _5805_;
wire _5806_;
wire _5807_;
wire _5808_;
wire _5809_;
wire _5810_;
wire _5811_;
wire _5812_;
wire _5813_;
wire _5814_;
wire _5815_;
wire _5816_;
wire _5817_;
wire _5818_;
wire _5819_;
wire _5820_;
wire _5821_;
wire _5822_;
wire _5823_;
wire _5824_;
wire _5825_;
wire _5826_;
wire _5827_;
wire _5828_;
wire _5829_;
wire _5830_;
wire _5831_;
wire _5832_;
wire _5833_;
wire _5834_;
wire _5835_;
wire _5836_;
wire _5837_;
wire _5838_;
wire _5839_;
wire _5840_;
wire _5841_;
wire _5842_;
wire _5843_;
wire _5844_;
wire _5845_;
wire _5846_;
wire _5847_;
wire _5848_;
wire _5849_;
wire _5850_;
wire _5851_;
wire _5852_;
wire _5853_;
wire _5854_;
wire _5855_;
wire _5856_;
wire _5857_;
wire _5858_;
wire _5859_;
wire _5860_;
wire _5861_;
wire _5862_;
wire _5863_;
wire _5864_;
wire _5865_;
wire _5866_;
wire _5867_;
wire _5868_;
wire _5869_;
wire _5870_;
wire _5871_;
wire _5872_;
wire _5873_;
wire _5874_;
wire _5875_;
wire _5876_;
wire _5877_;
wire _5878_;
wire _5879_;
wire _5880_;
wire _5881_;
wire _5882_;
wire _5883_;
wire _5884_;
wire _5885_;
wire _5886_;
wire _5887_;
wire _5888_;
wire _5889_;
wire _5890_;
wire _5891_;
wire _5892_;
wire _5893_;
wire _5894_;
wire _5895_;
wire _5896_;
wire _5897_;
wire _5898_;
wire _5899_;
wire _5900_;
wire _5901_;
wire _5902_;
wire _5903_;
wire _5904_;
wire _5905_;
wire _5906_;
wire _5907_;
wire _5908_;
wire _5909_;
wire _5910_;
wire _5911_;
wire _5912_;
wire _5913_;
wire _5914_;
wire _5915_;
wire _5916_;
wire _5917_;
wire _5918_;
wire _5919_;
wire _5920_;
wire _5921_;
wire _5922_;
wire _5923_;
wire _5924_;
wire _5925_;
wire _5926_;
wire _5927_;
wire _5928_;
wire _5929_;
wire _5930_;
wire _5931_;
wire _5932_;
wire _5933_;
wire _5934_;
wire _5935_;
wire _5936_;
wire _5937_;
wire _5938_;
wire _5939_;
wire _5940_;
wire _5941_;
wire _5942_;
wire _5943_;
wire _5944_;
wire _5945_;
wire _5946_;
wire _5947_;
wire _5948_;
wire _5949_;
wire _5950_;
wire _5951_;
wire _5952_;
wire _5953_;
wire _5954_;
wire _5955_;
wire _5956_;
wire _5957_;
wire _5958_;
wire _5959_;
wire _5960_;
wire _5961_;
wire _5962_;
wire _5963_;
wire _5964_;
wire _5965_;
wire _5966_;
wire _5967_;
wire _5968_;
wire _5969_;
wire _5970_;
wire _5971_;
wire _5972_;
wire _5973_;
wire _5974_;
wire _5975_;
wire _5976_;
wire _5977_;
wire _5978_;
wire _5979_;
wire _5980_;
wire _5981_;
wire _5982_;
wire _5983_;
wire _5984_;
wire _5985_;
wire _5986_;
wire _5987_;
wire _5988_;
wire _5989_;
wire _5990_;
wire _5991_;
wire _5992_;
wire _5993_;
wire _5994_;
wire _5995_;
wire _5996_;
wire _5997_;
wire _5998_;
wire _5999_;
wire _6000_;
wire _6001_;
wire _6002_;
wire _6003_;
wire _6004_;
wire _6005_;
wire _6006_;
wire _6007_;
wire _6008_;
wire _6009_;
wire _6010_;
wire _6011_;
wire _6012_;
wire _6013_;
wire _6014_;
wire _6015_;
wire _6016_;
wire _6017_;
wire _6018_;
wire _6019_;
wire _6020_;
wire _6021_;
wire _6022_;
wire _6023_;
wire _6024_;
wire _6025_;
wire _6026_;
wire _6027_;
wire _6028_;
wire _6029_;
wire _6030_;
wire _6031_;
wire _6032_;
wire _6033_;
wire _6034_;
wire _6035_;
wire _6036_;
wire _6037_;
wire _6038_;
wire _6039_;
wire _6040_;
wire _6041_;
wire _6042_;
wire _6043_;
wire _6044_;
wire _6045_;
wire _6046_;
wire _6047_;
wire _6048_;
wire _6049_;
wire _6050_;
wire _6051_;
wire _6052_;
wire _6053_;
wire _6054_;
wire _6055_;
wire _6056_;
wire _6057_;
wire _6058_;
wire _6059_;
wire _6060_;
wire _6061_;
wire _6062_;
wire _6063_;
wire _6064_;
wire _6065_;
wire _6066_;
wire _6067_;
wire _6068_;
wire _6069_;
wire _6070_;
wire _6071_;
wire _6072_;
wire _6073_;
wire _6074_;
wire _6075_;
wire _6076_;
wire _6077_;
wire _6078_;
wire _6079_;
wire _6080_;
wire _6081_;
wire _6082_;
wire _6083_;
wire _6084_;
wire _6085_;
wire _6086_;
wire _6087_;
wire _6088_;
wire _6089_;
wire _6090_;
wire _6091_;
wire _6092_;
wire _6093_;
wire _6094_;
wire _6095_;
wire _6096_;
wire _6097_;
wire _6098_;
wire _6099_;
wire _6100_;
wire _6101_;
wire _6102_;
wire _6103_;
wire _6104_;
wire _6105_;
wire _6106_;
wire _6107_;
wire _6108_;
wire _6109_;
wire _6110_;
wire _6111_;
wire _6112_;
wire _6113_;
wire _6114_;
wire _6115_;
wire _6116_;
wire _6117_;
wire _6118_;
wire _6119_;
wire _6120_;
wire _6121_;
wire _6122_;
wire _6123_;
wire _6124_;
wire _6125_;
wire _6126_;
wire _6127_;
wire _6128_;
wire _6129_;
wire _6130_;
wire _6131_;
wire _6132_;
wire _6133_;
wire _6134_;
wire _6135_;
wire _6136_;
wire _6137_;
wire _6138_;
wire _6139_;
wire _6140_;
wire _6141_;
wire _6142_;
wire _6143_;
wire _6144_;
wire _6145_;
wire _6146_;
wire _6147_;
wire _6148_;
wire _6149_;
wire _6150_;
wire _6151_;
wire _6152_;
wire _6153_;
wire _6154_;
wire _6155_;
wire _6156_;
wire _6157_;
wire _6158_;
wire _6159_;
wire _6160_;
wire _6161_;
wire _6162_;
wire _6163_;
wire _6164_;
wire _6165_;
wire _6166_;
wire _6167_;
wire _6168_;
wire _6169_;
wire _6170_;
wire _6171_;
wire _6172_;
wire _6173_;
wire _6174_;
wire _6175_;
wire _6176_;
wire _6177_;
wire _6178_;
wire _6179_;
wire _6180_;
wire _6181_;
wire _6182_;
wire _6183_;
wire _6184_;
wire _6185_;
wire _6186_;
wire _6187_;
wire _6188_;
wire _6189_;
wire _6190_;
wire _6191_;
wire _6192_;
wire _6193_;
wire _6194_;
wire _6195_;
wire _6196_;
wire _6197_;
wire _6198_;
wire _6199_;
wire _6200_;
wire _6201_;
wire _6202_;
wire _6203_;
wire _6204_;
wire _6205_;
wire _6206_;
wire _6207_;
wire _6208_;
wire _6209_;
wire _6210_;
wire _6211_;
wire _6212_;
wire _6213_;
wire _6214_;
wire _6215_;
wire _6216_;
wire _6217_;
wire _6218_;
wire _6219_;
wire _6220_;
wire _6221_;
wire _6222_;
wire _6223_;
wire _6224_;
wire _6225_;
wire _6226_;
wire _6227_;
wire _6228_;
wire _6229_;
wire _6230_;
wire _6231_;
wire _6232_;
wire _6233_;
wire _6234_;
wire _6235_;
wire _6236_;
wire _6237_;
wire _6238_;
wire _6239_;
wire _6240_;
wire _6241_;
wire _6242_;
wire _6243_;
wire _6244_;
wire _6245_;
wire _6246_;
wire _6247_;
wire _6248_;
wire _6249_;
wire _6250_;
wire _6251_;
wire _6252_;
wire _6253_;
wire _6254_;
wire _6255_;
wire _6256_;
wire _6257_;
wire _6258_;
wire _6259_;
wire _6260_;
wire _6261_;
wire _6262_;
wire _6263_;
wire _6264_;
wire _6265_;
wire _6266_;
wire _6267_;
wire _6268_;
wire _6269_;
wire _6270_;
wire _6271_;
wire _6272_;
wire _6273_;
wire _6274_;
wire _6275_;
wire _6276_;
wire _6277_;
wire _6278_;
wire _6279_;
wire _6280_;
wire _6281_;
wire _6282_;
wire _6283_;
wire _6284_;
wire _6285_;
wire _6286_;
wire _6287_;
wire _6288_;
wire _6289_;
wire _6290_;
wire _6291_;
wire _6292_;
wire _6293_;
wire _6294_;
wire _6295_;
wire _6296_;
wire _6297_;
wire _6298_;
wire _6299_;
wire _6300_;
wire _6301_;
wire _6302_;
wire _6303_;
wire _6304_;
wire _6305_;
wire _6306_;
wire _6307_;
wire _6308_;
wire _6309_;
wire _6310_;
wire _6311_;
wire _6312_;
wire _6313_;
wire _6314_;
wire _6315_;
wire _6316_;
wire _6317_;
wire _6318_;
wire _6319_;
wire _6320_;
wire _6321_;
wire _6322_;
wire _6323_;
wire _6324_;
wire _6325_;
wire _6326_;
wire _6327_;
wire _6328_;
wire _6329_;
wire _6330_;
wire _6331_;
wire _6332_;
wire _6333_;
wire _6334_;
wire _6335_;
wire _6336_;
wire _6337_;
wire _6338_;
wire _6339_;
wire _6340_;
wire _6341_;
wire _6342_;
wire _6343_;
wire _6344_;
wire _6345_;
wire _6346_;
wire _6347_;
wire _6348_;
wire _6349_;
wire _6350_;
wire _6351_;
wire _6352_;
wire _6353_;
wire _6354_;
wire _6355_;
wire _6356_;
wire _6357_;
wire _6358_;
wire _6359_;
wire _6360_;
wire _6361_;
wire _6362_;
wire _6363_;
wire _6364_;
wire _6365_;
wire _6366_;
wire _6367_;
wire _6368_;
wire _6369_;
wire _6370_;
wire _6371_;
wire _6372_;
wire _6373_;
wire _6374_;
wire _6375_;
wire _6376_;
wire _6377_;
wire _6378_;
wire _6379_;
wire _6380_;
wire _6381_;
wire _6382_;
wire _6383_;
wire _6384_;
wire _6385_;
wire _6386_;
wire _6387_;
wire _6388_;
wire _6389_;
wire _6390_;
wire _6391_;
wire _6392_;
wire _6393_;
wire _6394_;
wire _6395_;
wire _6396_;
wire _6397_;
wire _6398_;
wire _6399_;
wire _6400_;
wire _6401_;
wire _6402_;
wire _6403_;
wire _6404_;
wire _6405_;
wire _6406_;
wire _6407_;
wire _6408_;
wire _6409_;
wire _6410_;
wire _6411_;
wire _6412_;
wire _6413_;
wire _6414_;
wire _6415_;
wire _6416_;
wire _6417_;
wire _6418_;
wire _6419_;
wire _6420_;
wire _6421_;
wire _6422_;
wire _6423_;
wire _6424_;
wire _6425_;
wire _6426_;
wire _6427_;
wire _6428_;
wire _6429_;
wire _6430_;
wire _6431_;
wire _6432_;
wire _6433_;
wire _6434_;
wire _6435_;
wire _6436_;
wire _6437_;
wire _6438_;
wire _6439_;
wire _6440_;
wire _6441_;
wire _6442_;
wire _6443_;
wire _6444_;
wire _6445_;
wire _6446_;
wire _6447_;
wire _6448_;
wire _6449_;
wire _6450_;
wire _6451_;
wire _6452_;
wire _6453_;
wire _6454_;
wire _6455_;
wire _6456_;
wire _6457_;
wire _6458_;
wire _6459_;
wire _6460_;
wire _6461_;
wire _6462_;
wire _6463_;
wire _6464_;
wire _6465_;
wire _6466_;
wire _6467_;
wire _6468_;
wire _6469_;
wire _6470_;
wire _6471_;
wire _6472_;
wire _6473_;
wire _6474_;
wire _6475_;
wire _6476_;
wire _6477_;
wire _6478_;
wire _6479_;
wire _6480_;
wire _6481_;
wire _6482_;
wire _6483_;
wire _6484_;
wire _6485_;
wire _6486_;
wire _6487_;
wire _6488_;
wire _6489_;
wire _6490_;
wire _6491_;
wire _6492_;
wire _6493_;
wire _6494_;
wire _6495_;
wire _6496_;
wire _6497_;
wire _6498_;
wire _6499_;
wire _6500_;
wire _6501_;
wire _6502_;
wire _6503_;
wire _6504_;
wire _6505_;
wire _6506_;
wire _6507_;
wire _6508_;
wire _6509_;
wire _6510_;
wire _6511_;
wire _6512_;
wire _6513_;
wire _6514_;
wire _6515_;
wire _6516_;
wire _6517_;
wire _6518_;
wire _6519_;
wire _6520_;
wire _6521_;
wire _6522_;
wire _6523_;
wire _6524_;
wire _6525_;
wire _6526_;
wire _6527_;
wire _6528_;
wire _6529_;
wire _6530_;
wire _6531_;
wire _6532_;
wire _6533_;
wire _6534_;
wire _6535_;
wire _6536_;
wire _6537_;
wire _6538_;
wire _6539_;
wire _6540_;
wire _6541_;
wire _6542_;
wire _6543_;
wire _6544_;
wire _6545_;
wire _6546_;
wire _6547_;
wire _6548_;
wire _6549_;
wire _6550_;
wire _6551_;
wire _6552_;
wire _6553_;
wire _6554_;
wire _6555_;
wire _6556_;
wire _6557_;
wire _6558_;
wire _6559_;
wire _6560_;
wire _6561_;
wire _6562_;
wire _6563_;
wire _6564_;
wire _6565_;
wire _6566_;
wire _6567_;
wire _6568_;
wire _6569_;
wire _6570_;
wire _6571_;
wire _6572_;
wire _6573_;
wire _6574_;
wire _6575_;
wire _6576_;
wire _6577_;
wire _6578_;
wire _6579_;
wire _6580_;
wire _6581_;
wire _6582_;
wire _6583_;
wire _6584_;
wire _6585_;
wire _6586_;
wire _6587_;
wire _6588_;
wire _6589_;
wire _6590_;
wire _6591_;
wire _6592_;
wire _6593_;
wire _6594_;
wire _6595_;
wire _6596_;
wire _6597_;
wire _6598_;
wire _6599_;
wire _6600_;
wire _6601_;
wire _6602_;
wire _6603_;
wire _6604_;
wire _6605_;
wire _6606_;
wire _6607_;
wire _6608_;
wire _6609_;
wire _6610_;
wire _6611_;
wire _6612_;
wire _6613_;
wire _6614_;
wire _6615_;
wire _6616_;
wire _6617_;
wire _6618_;
wire _6619_;
wire _6620_;
wire _6621_;
wire _6622_;
wire _6623_;
wire _6624_;
wire _6625_;
wire _6626_;
wire _6627_;
wire _6628_;
wire _6629_;
wire _6630_;
wire _6631_;
wire _6632_;
wire _6633_;
wire _6634_;
wire _6635_;
wire _6636_;
wire _6637_;
wire _6638_;
wire _6639_;
wire _6640_;
wire _6641_;
wire _6642_;
wire _6643_;
wire _6644_;
wire _6645_;
wire _6646_;
wire _6647_;
wire _6648_;
wire _6649_;
wire _6650_;
wire _6651_;
wire _6652_;
wire _6653_;
wire _6654_;
wire _6655_;
wire _6656_;
wire _6657_;
wire _6658_;
wire _6659_;
wire _6660_;
wire _6661_;
wire _6662_;
wire _6663_;
wire _6664_;
wire _6665_;
wire _6666_;
wire _6667_;
wire _6668_;
wire _6669_;
wire _6670_;
wire _6671_;
wire _6672_;
wire _6673_;
wire _6674_;
wire _6675_;
wire _6676_;
wire _6677_;
wire _6678_;
wire _6679_;
wire _6680_;
wire _6681_;
wire _6682_;
wire _6683_;
wire _6684_;
wire _6685_;
wire _6686_;
wire _6687_;
wire _6688_;
wire _6689_;
wire _6690_;
wire _6691_;
wire _6692_;
wire _6693_;
wire _6694_;
wire _6695_;
wire _6696_;
wire _6697_;
wire _6698_;
wire _6699_;
wire _6700_;
wire _6701_;
wire _6702_;
wire _6703_;
wire _6704_;
wire _6705_;
wire _6706_;
wire _6707_;
wire _6708_;
wire _6709_;
wire _6710_;
wire _6711_;
wire _6712_;
wire _6713_;
wire _6714_;
wire _6715_;
wire _6716_;
wire _6717_;
wire _6718_;
wire _6719_;
wire _6720_;
wire _6721_;
wire _6722_;
wire _6723_;
wire _6724_;
wire _6725_;
wire _6726_;
wire _6727_;
wire _6728_;
wire _6729_;
wire _6730_;
wire _6731_;
wire _6732_;
wire _6733_;
wire _6734_;
wire _6735_;
wire _6736_;
wire _6737_;
wire _6738_;
wire _6739_;
wire _6740_;
wire _6741_;
wire _6742_;
wire _6743_;
wire _6744_;
wire _6745_;
wire _6746_;
wire _6747_;
wire _6748_;
wire _6749_;
wire _6750_;
wire _6751_;
wire _6752_;
wire _6753_;
wire _6754_;
wire _6755_;
wire _6756_;
wire _6757_;
wire _6758_;
wire _6759_;
wire _6760_;
wire _6761_;
wire _6762_;
wire _6763_;
wire _6764_;
wire _6765_;
wire _6766_;
wire _6767_;
wire _6768_;
wire _6769_;
wire _6770_;
wire _6771_;
wire _6772_;
wire _6773_;
wire _6774_;
wire _6775_;
wire _6776_;
wire _6777_;
wire _6778_;
wire _6779_;
wire _6780_;
wire _6781_;
wire _6782_;
wire _6783_;
wire _6784_;
wire _6785_;
wire _6786_;
wire _6787_;
wire _6788_;
wire _6789_;
wire _6790_;
wire _6791_;
wire _6792_;
wire _6793_;
wire _6794_;
wire _6795_;
wire _6796_;
wire _6797_;
wire _6798_;
wire _6799_;
wire _6800_;
wire _6801_;
wire _6802_;
wire _6803_;
wire _6804_;
wire _6805_;
wire _6806_;
wire _6807_;
wire _6808_;
wire _6809_;
wire _6810_;
wire _6811_;
wire _6812_;
wire _6813_;
wire _6814_;
wire _6815_;
wire _6816_;
wire _6817_;
wire _6818_;
wire _6819_;
wire _6820_;
wire _6821_;
wire _6822_;
wire _6823_;
wire _6824_;
wire _6825_;
wire _6826_;
wire _6827_;
wire _6828_;
wire _6829_;
wire _6830_;
wire _6831_;
wire _6832_;
wire _6833_;
wire _6834_;
wire _6835_;
wire _6836_;
wire _6837_;
wire _6838_;
wire _6839_;
wire _6840_;
wire _6841_;
wire _6842_;
wire _6843_;
wire _6844_;
wire _6845_;
wire _6846_;
wire _6847_;
wire _6848_;
wire _6849_;
wire _6850_;
wire _6851_;
wire _6852_;
wire _6853_;
wire _6854_;
wire _6855_;
wire _6856_;
wire _6857_;
wire _6858_;
wire _6859_;
wire _6860_;
wire _6861_;
wire _6862_;
wire _6863_;
wire _6864_;
wire _6865_;
wire _6866_;
wire _6867_;
wire _6868_;
wire _6869_;
wire _6870_;
wire _6871_;
wire _6872_;
wire _6873_;
wire _6874_;
wire _6875_;
wire _6876_;
wire _6877_;
wire _6878_;
wire _6879_;
wire _6880_;
wire _6881_;
wire _6882_;
wire _6883_;
wire _6884_;
wire _6885_;
wire _6886_;
wire _6887_;
wire _6888_;
wire _6889_;
wire _6890_;
wire _6891_;
wire _6892_;
wire _6893_;
wire _6894_;
wire _6895_;
wire _6896_;
wire _6897_;
wire _6898_;
wire _6899_;
wire _6900_;
wire _6901_;
wire _6902_;
wire _6903_;
wire _6904_;
wire _6905_;
wire _6906_;
wire _6907_;
wire _6908_;
wire _6909_;
wire _6910_;
wire _6911_;
wire _6912_;
wire _6913_;
wire _6914_;
wire _6915_;
wire _6916_;
wire _6917_;
wire _6918_;
wire _6919_;
wire _6920_;
wire _6921_;
wire _6922_;
wire _6923_;
wire _6924_;
wire _6925_;
wire _6926_;
wire _6927_;
wire _6928_;
wire _6929_;
wire _6930_;
wire _6931_;
wire _6932_;
wire _6933_;
wire _6934_;
wire _6935_;
wire _6936_;
wire _6937_;
wire _6938_;
wire _6939_;
wire _6940_;
wire _6941_;
wire _6942_;
wire _6943_;
wire _6944_;
wire _6945_;
wire _6946_;
wire _6947_;
wire _6948_;
wire _6949_;
wire _6950_;
wire _6951_;
wire _6952_;
wire _6953_;
wire _6954_;
wire _6955_;
wire _6956_;
wire _6957_;
wire _6958_;
wire _6959_;
wire _6960_;
wire _6961_;
wire _6962_;
wire _6963_;
wire _6964_;
wire _6965_;
wire _6966_;
wire _6967_;
wire _6968_;
wire _6969_;
wire _6970_;
wire _6971_;
wire _6972_;
wire _6973_;
wire _6974_;
wire _6975_;
wire _6976_;
wire _6977_;
wire _6978_;
wire _6979_;
wire _6980_;
wire _6981_;
wire _6982_;
wire _6983_;
wire _6984_;
wire _6985_;
wire _6986_;
wire _6987_;
wire _6988_;
wire _6989_;
wire _6990_;
wire _6991_;
wire _6992_;
wire _6993_;
wire _6994_;
wire _6995_;
wire _6996_;
wire _6997_;
wire _6998_;
wire _6999_;
wire _7000_;
wire _7001_;
wire _7002_;
wire _7003_;
wire _7004_;
wire _7005_;
wire _7006_;
wire _7007_;
wire _7008_;
wire _7009_;
wire _7010_;
wire _7011_;
wire _7012_;
wire _7013_;
wire _7014_;
wire _7015_;
wire _7016_;
wire _7017_;
wire _7018_;
wire _7019_;
wire _7020_;
wire _7021_;
wire _7022_;
wire _7023_;
wire _7024_;
wire _7025_;
wire _7026_;
wire _7027_;
wire _7028_;
wire _7029_;
wire _7030_;
wire _7031_;
wire _7032_;
wire _7033_;
wire _7034_;
wire _7035_;
wire _7036_;
wire _7037_;
wire _7038_;
wire _7039_;
wire _7040_;
wire _7041_;
wire _7042_;
wire _7043_;
wire _7044_;
wire _7045_;
wire _7046_;
wire _7047_;
wire _7048_;
wire _7049_;
wire _7050_;
wire _7051_;
wire _7052_;
wire _7053_;
wire _7054_;
wire _7055_;
wire _7056_;
wire _7057_;
wire _7058_;
wire _7059_;
wire _7060_;
wire _7061_;
wire _7062_;
wire _7063_;
wire _7064_;
wire _7065_;
wire _7066_;
wire _7067_;
wire _7068_;
wire _7069_;
wire _7070_;
wire _7071_;
wire _7072_;
wire _7073_;
wire _7074_;
wire _7075_;
wire _7076_;
wire _7077_;
wire _7078_;
wire _7079_;
wire _7080_;
wire _7081_;
wire _7082_;
wire _7083_;
wire _7084_;
wire _7085_;
wire _7086_;
wire _7087_;
wire _7088_;
wire _7089_;
wire _7090_;
wire _7091_;
wire _7092_;
wire _7093_;
wire _7094_;
wire _7095_;
wire _7096_;
wire _7097_;
wire _7098_;
wire _7099_;
wire _7100_;
wire _7101_;
wire _7102_;
wire _7103_;
wire _7104_;
wire _7105_;
wire _7106_;
wire _7107_;
wire _7108_;
wire _7109_;
wire _7110_;
wire _7111_;
wire _7112_;
wire _7113_;
wire _7114_;
wire _7115_;
wire _7116_;
wire _7117_;
wire _7118_;
wire _7119_;
wire _7120_;
wire _7121_;
wire _7122_;
wire _7123_;
wire _7124_;
wire _7125_;
wire _7126_;
wire _7127_;
wire _7128_;
wire _7129_;
wire _7130_;
wire _7131_;
wire _7132_;
wire _7133_;
wire _7134_;
wire _7135_;
wire _7136_;
wire _7137_;
wire _7138_;
wire _7139_;
wire _7140_;
wire _7141_;
wire _7142_;
wire _7143_;
wire _7144_;
wire _7145_;
wire _7146_;
wire _7147_;
wire _7148_;
wire _7149_;
wire _7150_;
wire _7151_;
wire _7152_;
wire _7153_;
wire _7154_;
wire _7155_;
wire _7156_;
wire _7157_;
wire _7158_;
wire _7159_;
wire _7160_;
wire _7161_;
wire _7162_;
wire _7163_;
wire _7164_;
wire _7165_;
wire _7166_;
wire _7167_;
wire _7168_;
wire _7169_;
wire _7170_;
wire _7171_;
wire _7172_;
wire _7173_;
wire _7174_;
wire _7175_;
wire _7176_;
wire _7177_;
wire _7178_;
wire _7179_;
wire _7180_;
wire _7181_;
wire _7182_;
wire _7183_;
wire _7184_;
wire _7185_;
wire _7186_;
wire _7187_;
wire _7188_;
wire _7189_;
wire _7190_;
wire _7191_;
wire _7192_;
wire _7193_;
wire _7194_;
wire _7195_;
wire _7196_;
wire _7197_;
wire _7198_;
wire _7199_;
wire _7200_;
wire _7201_;
wire _7202_;
wire _7203_;
wire _7204_;
wire _7205_;
wire _7206_;
wire _7207_;
wire _7208_;
wire _7209_;
wire _7210_;
wire _7211_;
wire _7212_;
wire _7213_;
wire _7214_;
wire _7215_;
wire _7216_;
wire _7217_;
wire _7218_;
wire _7219_;
wire _7220_;
wire _7221_;
wire _7222_;
wire _7223_;
wire _7224_;
wire _7225_;
wire _7226_;
wire _7227_;
wire _7228_;
wire _7229_;
wire _7230_;
wire _7231_;
wire _7232_;
wire _7233_;
wire _7234_;
wire _7235_;
wire _7236_;
wire _7237_;
wire _7238_;
wire _7239_;
wire _7240_;
wire _7241_;
wire _7242_;
wire _7243_;
wire _7244_;
wire _7245_;
wire _7246_;
wire _7247_;
wire _7248_;
wire _7249_;
wire _7250_;
wire _7251_;
wire _7252_;
wire _7253_;
wire _7254_;
wire _7255_;
wire _7256_;
wire _7257_;
wire _7258_;
wire _7259_;
wire _7260_;
wire _7261_;
wire _7262_;
wire _7263_;
wire _7264_;
wire _7265_;
wire _7266_;
wire _7267_;
wire _7268_;
wire _7269_;
wire _7270_;
wire _7271_;
wire _7272_;
wire _7273_;
wire _7274_;
wire _7275_;
wire _7276_;
wire _7277_;
wire _7278_;
wire _7279_;
wire _7280_;
wire _7281_;
wire _7282_;
wire _7283_;
wire _7284_;
wire _7285_;
wire _7286_;
wire _7287_;
wire _7288_;
wire _7289_;
wire _7290_;
wire _7291_;
wire _7292_;
wire _7293_;
wire _7294_;
wire _7295_;
wire _7296_;
wire _7297_;
wire _7298_;
wire _7299_;
wire _7300_;
wire _7301_;
wire _7302_;
wire _7303_;
wire _7304_;
wire _7305_;
wire _7306_;
wire _7307_;
wire _7308_;
wire _7309_;
wire _7310_;
wire _7311_;
wire _7312_;
wire _7313_;
wire _7314_;
wire _7315_;
wire _7316_;
wire _7317_;
wire _7318_;
wire _7319_;
wire _7320_;
wire _7321_;
wire _7322_;
wire _7323_;
wire _7324_;
wire _7325_;
wire _7326_;
wire _7327_;
wire _7328_;
wire _7329_;
wire _7330_;
wire _7331_;
wire _7332_;
wire _7333_;
wire _7334_;
wire _7335_;
wire _7336_;
wire _7337_;
wire _7338_;
wire _7339_;
wire _7340_;
wire _7341_;
wire _7342_;
wire _7343_;
wire _7344_;
wire _7345_;
wire _7346_;
wire _7347_;
wire _7348_;
wire _7349_;
wire _7350_;
wire _7351_;
wire _7352_;
wire _7353_;
wire _7354_;
wire _7355_;
wire _7356_;
wire _7357_;
wire _7358_;
wire _7359_;
wire _7360_;
wire _7361_;
wire _7362_;
wire _7363_;
wire _7364_;
wire _7365_;
wire _7366_;
wire _7367_;
wire _7368_;
wire _7369_;
wire _7370_;
wire _7371_;
wire _7372_;
wire _7373_;
wire _7374_;
wire _7375_;
wire _7376_;
wire _7377_;
wire _7378_;
wire _7379_;
wire _7380_;
wire _7381_;
wire _7382_;
wire _7383_;
wire _7384_;
wire _7385_;
wire _7386_;
wire _7387_;
wire _7388_;
wire _7389_;
wire _7390_;
wire _7391_;
wire _7392_;
wire _7393_;
wire _7394_;
wire _7395_;
wire _7396_;
wire _7397_;
wire _7398_;
wire _7399_;
wire _7400_;
wire _7401_;
wire _7402_;
wire _7403_;
wire _7404_;
wire _7405_;
wire _7406_;
wire _7407_;
wire _7408_;
wire _7409_;
wire _7410_;
wire _7411_;
wire _7412_;
wire _7413_;
wire _7414_;
wire _7415_;
wire _7416_;
wire _7417_;
wire _7418_;
wire _7419_;
wire _7420_;
wire _7421_;
wire _7422_;
wire _7423_;
wire _7424_;
wire _7425_;
wire _7426_;
wire _7427_;
wire _7428_;
wire _7429_;
wire _7430_;
wire _7431_;
wire _7432_;
wire _7433_;
wire _7434_;
wire _7435_;
wire _7436_;
wire _7437_;
wire _7438_;
wire _7439_;
wire _7440_;
wire _7441_;
wire _7442_;
wire _7443_;
wire _7444_;
wire _7445_;
wire _7446_;
wire _7447_;
wire _7448_;
wire _7449_;
wire _7450_;
wire _7451_;
wire _7452_;
wire _7453_;
wire _7454_;
wire _7455_;
wire _7456_;
wire _7457_;
wire _7458_;
wire _7459_;
wire _7460_;
wire _7461_;
wire _7462_;
wire _7463_;
wire _7464_;
wire _7465_;
wire _7466_;
wire _7467_;
wire _7468_;
wire _7469_;
wire _7470_;
wire _7471_;
wire _7472_;
wire _7473_;
wire _7474_;
wire _7475_;
wire _7476_;
wire _7477_;
wire _7478_;
wire _7479_;
wire _7480_;
wire _7481_;
wire _7482_;
wire _7483_;
wire _7484_;
wire _7485_;
wire _7486_;
wire _7487_;
wire _7488_;
wire _7489_;
wire _7490_;
wire _7491_;
wire _7492_;
wire _7493_;
wire _7494_;
wire _7495_;
wire _7496_;
wire _7497_;
wire _7498_;
wire _7499_;
wire _7500_;
wire _7501_;
wire _7502_;
wire _7503_;
wire _7504_;
wire _7505_;
wire _7506_;
wire _7507_;
wire _7508_;
wire _7509_;
wire _7510_;
wire _7511_;
wire _7512_;
wire _7513_;
wire _7514_;
wire _7515_;
wire _7516_;
wire _7517_;
wire _7518_;
wire _7519_;
wire _7520_;
wire _7521_;
wire _7522_;
wire _7523_;
wire _7524_;
wire _7525_;
wire _7526_;
wire _7527_;
wire _7528_;
wire _7529_;
wire _7530_;
wire _7531_;
wire _7532_;
wire _7533_;
wire _7534_;
wire _7535_;
wire _7536_;
wire _7537_;
wire _7538_;
wire _7539_;
wire _7540_;
wire _7541_;
wire _7542_;
wire _7543_;
wire _7544_;
wire _7545_;
wire _7546_;
wire _7547_;
wire _7548_;
wire _7549_;
wire _7550_;
wire _7551_;
wire _7552_;
wire _7553_;
wire _7554_;
wire _7555_;
wire _7556_;
wire _7557_;
wire _7558_;
wire _7559_;
wire _7560_;
wire _7561_;
wire _7562_;
wire _7563_;
wire _7564_;
wire _7565_;
wire _7566_;
wire _7567_;
wire _7568_;
wire _7569_;
wire _7570_;
wire _7571_;
wire _7572_;
wire _7573_;
wire _7574_;
wire _7575_;
wire _7576_;
wire _7577_;
wire _7578_;
wire _7579_;
wire _7580_;
wire _7581_;
wire _7582_;
wire _7583_;
wire _7584_;
wire _7585_;
wire _7586_;
wire _7587_;
wire _7588_;
wire _7589_;
wire _7590_;
wire _7591_;
wire _7592_;
wire _7593_;
wire _7594_;
wire _7595_;
wire _7596_;
wire _7597_;
wire _7598_;
wire _7599_;
wire _7600_;
wire _7601_;
wire _7602_;
wire _7603_;
wire _7604_;
wire _7605_;
wire _7606_;
wire _7607_;
wire _7608_;
wire _7609_;
wire _7610_;
wire _7611_;
wire _7612_;
wire _7613_;
wire _7614_;
wire _7615_;
wire _7616_;
wire _7617_;
wire _7618_;
wire _7619_;
wire _7620_;
wire _7621_;
wire _7622_;
wire _7623_;
wire _7624_;
wire _7625_;
wire _7626_;
wire _7627_;
wire _7628_;
wire _7629_;
wire _7630_;
wire _7631_;
wire _7632_;
wire _7633_;
wire _7634_;
wire _7635_;
wire _7636_;
wire _7637_;
wire _7638_;
wire _7639_;
wire _7640_;
wire _7641_;
wire _7642_;
wire _7643_;
wire _7644_;
wire _7645_;
wire _7646_;
wire _7647_;
wire _7648_;
wire _7649_;
wire _7650_;
wire _7651_;
wire _7652_;
wire _7653_;
wire _7654_;
wire _7655_;
wire _7656_;
wire _7657_;
wire _7658_;
wire _7659_;
wire _7660_;
wire _7661_;
wire _7662_;
wire _7663_;
wire _7664_;
wire _7665_;
wire _7666_;
wire _7667_;
wire _7668_;
wire _7669_;
wire _7670_;
wire _7671_;
wire _7672_;
wire _7673_;
wire _7674_;
wire _7675_;
wire _7676_;
wire _7677_;
wire _7678_;
wire _7679_;
wire _7680_;
wire _7681_;
wire _7682_;
wire _7683_;
wire _7684_;
wire _7685_;
wire _7686_;
wire _7687_;
wire _7688_;
wire _7689_;
wire _7690_;
wire _7691_;
wire _7692_;
wire _7693_;
wire _7694_;
wire _7695_;
wire _7696_;
wire _7697_;
wire _7698_;
wire _7699_;
wire _7700_;
wire _7701_;
wire _7702_;
wire _7703_;
wire _7704_;
wire _7705_;
wire _7706_;
wire _7707_;
wire _7708_;
wire _7709_;
wire _7710_;
wire _7711_;
wire _7712_;
wire _7713_;
wire _7714_;
wire _7715_;
wire _7716_;
wire _7717_;
wire _7718_;
wire _7719_;
wire _7720_;
wire _7721_;
wire _7722_;
wire _7723_;
wire _7724_;
wire _7725_;
wire _7726_;
wire _7727_;
wire _7728_;
wire _7729_;
wire _7730_;
wire _7731_;
wire _7732_;
wire _7733_;
wire _7734_;
wire _7735_;
wire _7736_;
wire _7737_;
wire _7738_;
wire _7739_;
wire _7740_;
wire _7741_;
wire _7742_;
wire _7743_;
wire _7744_;
wire _7745_;
wire _7746_;
wire _7747_;
wire _7748_;
wire _7749_;
wire _7750_;
wire _7751_;
wire _7752_;
wire _7753_;
wire _7754_;
wire _7755_;
wire _7756_;
wire _7757_;
wire _7758_;
wire _7759_;
wire _7760_;
wire _7761_;
wire _7762_;
wire _7763_;
wire _7764_;
wire _7765_;
wire _7766_;
wire _7767_;
wire _7768_;
wire _7769_;
wire _7770_;
wire _7771_;
wire _7772_;
wire _7773_;
wire _7774_;
wire _7775_;
wire _7776_;
wire _7777_;
wire _7778_;
wire _7779_;
wire _7780_;
wire _7781_;
wire _7782_;
wire _7783_;
wire _7784_;
wire _7785_;
wire _7786_;
wire _7787_;
wire _7788_;
wire _7789_;
wire _7790_;
wire _7791_;
wire _7792_;
wire _7793_;
wire _7794_;
wire _7795_;
wire _7796_;
wire _7797_;
wire _7798_;
wire _7799_;
wire _7800_;
wire _7801_;
wire _7802_;
wire _7803_;
wire _7804_;
wire _7805_;
wire _7806_;
wire _7807_;
wire _7808_;
wire _7809_;
wire _7810_;
wire _7811_;
wire _7812_;
wire _7813_;
wire _7814_;
wire _7815_;
wire _7816_;
wire _7817_;
wire _7818_;
wire _7819_;
wire _7820_;
wire _7821_;
wire _7822_;
wire _7823_;
wire _7824_;
wire _7825_;
wire _7826_;
wire _7827_;
wire _7828_;
wire _7829_;
wire _7830_;
wire _7831_;
wire _7832_;
wire _7833_;
wire _7834_;
wire _7835_;
wire _7836_;
wire _7837_;
wire _7838_;
wire _7839_;
wire _7840_;
wire _7841_;
wire _7842_;
wire _7843_;
wire _7844_;
wire _7845_;
wire _7846_;
wire _7847_;
wire _7848_;
wire _7849_;
wire _7850_;
wire _7851_;
wire _7852_;
wire _7853_;
wire _7854_;
wire _7855_;
wire _7856_;
wire _7857_;
wire _7858_;
wire _7859_;
wire _7860_;
wire _7861_;
wire _7862_;
wire _7863_;
wire _7864_;
wire _7865_;
wire _7866_;
wire _7867_;
wire _7868_;
wire _7869_;
wire _7870_;
wire _7871_;
wire _7872_;
wire _7873_;
wire _7874_;
wire _7875_;
wire _7876_;
wire _7877_;
wire _7878_;
wire _7879_;
wire _7880_;
wire _7881_;
wire _7882_;
wire _7883_;
wire _7884_;
wire _7885_;
wire _7886_;
wire _7887_;
wire _7888_;
wire _7889_;
wire _7890_;
wire _7891_;
wire _7892_;
wire _7893_;
wire _7894_;
wire _7895_;
wire _7896_;
wire _7897_;
wire _7898_;
wire _7899_;
wire _7900_;
wire _7901_;
wire _7902_;
wire _7903_;
wire _7904_;
wire _7905_;
wire _7906_;
wire _7907_;
wire _7908_;
wire _7909_;
wire _7910_;
wire _7911_;
wire _7912_;
wire _7913_;
wire _7914_;
wire _7915_;
wire _7916_;
wire _7917_;
wire _7918_;
wire _7919_;
wire _7920_;
wire _7921_;
wire _7922_;
wire _7923_;
wire _7924_;
wire _7925_;
wire _7926_;
wire _7927_;
wire _7928_;
wire _7929_;
wire _7930_;
wire _7931_;
wire _7932_;
wire _7933_;
wire _7934_;
wire _7935_;
wire _7936_;
wire _7937_;
wire _7938_;
wire _7939_;
wire _7940_;
wire _7941_;
wire _7942_;
wire _7943_;
wire _7944_;
wire _7945_;
wire _7946_;
wire _7947_;
wire _7948_;
wire _7949_;
wire _7950_;
wire _7951_;
wire _7952_;
wire _7953_;
wire _7954_;
wire _7955_;
wire _7956_;
wire _7957_;
wire _7958_;
wire _7959_;
wire _7960_;
wire _7961_;
wire _7962_;
wire _7963_;
wire _7964_;
wire _7965_;
wire _7966_;
wire _7967_;
wire _7968_;
wire _7969_;
wire _7970_;
wire _7971_;
wire _7972_;
wire _7973_;
wire _7974_;
wire _7975_;
wire _7976_;
wire _7977_;
wire _7978_;
wire _7979_;
wire _7980_;
wire _7981_;
wire _7982_;
wire _7983_;
wire _7984_;
wire _7985_;
wire _7986_;
wire _7987_;
wire _7988_;
wire _7989_;
wire _7990_;
wire _7991_;
wire _7992_;
wire _7993_;
wire _7994_;
wire _7995_;
wire _7996_;
wire _7997_;
wire _7998_;
wire _7999_;
wire _8000_;
wire _8001_;
wire _8002_;
wire _8003_;
wire _8004_;
wire _8005_;
wire _8006_;
wire _8007_;
wire _8008_;
wire _8009_;
wire _8010_;
wire _8011_;
wire _8012_;
wire _8013_;
wire _8014_;
wire _8015_;
wire _8016_;
wire _8017_;
wire _8018_;
wire _8019_;
wire _8020_;
wire _8021_;
wire _8022_;
wire _8023_;
wire _8024_;
wire _8025_;
wire _8026_;
wire _8027_;
wire _8028_;
wire _8029_;
wire _8030_;
wire _8031_;
wire _8032_;
wire _8033_;
wire _8034_;
wire _8035_;
wire _8036_;
wire _8037_;
wire _8038_;
wire _8039_;
wire _8040_;
wire _8041_;
wire _8042_;
wire _8043_;
wire _8044_;
wire _8045_;
wire _8046_;
wire _8047_;
wire _8048_;
wire _8049_;
wire _8050_;
wire _8051_;
wire _8052_;
wire _8053_;
wire _8054_;
wire _8055_;
wire _8056_;
wire _8057_;
wire _8058_;
wire _8059_;
wire _8060_;
wire _8061_;
wire _8062_;
wire _8063_;
wire _8064_;
wire _8065_;
wire _8066_;
wire _8067_;
wire _8068_;
wire _8069_;
wire _8070_;
wire _8071_;
wire _8072_;
wire _8073_;
wire _8074_;
wire _8075_;
wire _8076_;
wire _8077_;
wire _8078_;
wire _8079_;
wire _8080_;
wire _8081_;
wire _8082_;
wire _8083_;
wire _8084_;
wire _8085_;
wire _8086_;
wire _8087_;
wire _8088_;
wire _8089_;
wire _8090_;
wire _8091_;
wire _8092_;
wire _8093_;
wire _8094_;
wire _8095_;
wire _8096_;
wire _8097_;
wire _8098_;
wire _8099_;
wire _8100_;
wire _8101_;
wire _8102_;
wire _8103_;
wire _8104_;
wire _8105_;
wire _8106_;
wire _8107_;
wire _8108_;
wire _8109_;
wire _8110_;
wire _8111_;
wire _8112_;
wire _8113_;
wire _8114_;
wire _8115_;
wire _8116_;
wire _8117_;
wire _8118_;
wire _8119_;
wire _8120_;
wire _8121_;
wire _8122_;
wire _8123_;
wire _8124_;
wire _8125_;
wire _8126_;
wire _8127_;
wire _8128_;
wire _8129_;
wire _8130_;
wire _8131_;
wire _8132_;
wire _8133_;
wire _8134_;
wire _8135_;
wire _8136_;
wire _8137_;
wire _8138_;
wire _8139_;
wire _8140_;
wire _8141_;
wire _8142_;
wire _8143_;
wire _8144_;
wire _8145_;
wire _8146_;
wire _8147_;
wire _8148_;
wire _8149_;
wire _8150_;
wire _8151_;
wire _8152_;
wire _8153_;
wire _8154_;
wire _8155_;
wire _8156_;
wire _8157_;
wire _8158_;
wire _8159_;
wire _8160_;
wire _8161_;
wire _8162_;
wire _8163_;
wire _8164_;
wire _8165_;
wire _8166_;
wire _8167_;
wire _8168_;
wire _8169_;
wire _8170_;
wire _8171_;
wire _8172_;
wire _8173_;
wire _8174_;
wire _8175_;
wire _8176_;
wire _8177_;
wire _8178_;
wire _8179_;
wire _8180_;
wire _8181_;
wire _8182_;
wire _8183_;
wire _8184_;
wire _8185_;
wire _8186_;
wire _8187_;
wire _8188_;
wire _8189_;
wire _8190_;
wire _8191_;
wire _8192_;
wire _8193_;
wire _8194_;
wire _8195_;
wire _8196_;
wire _8197_;
wire _8198_;
wire _8199_;
wire _8200_;
wire _8201_;
wire _8202_;
wire _8203_;
wire _8204_;
wire _8205_;
wire _8206_;
wire _8207_;
wire _8208_;
wire _8209_;
wire _8210_;
wire _8211_;
wire _8212_;
wire _8213_;
wire _8214_;
wire _8215_;
wire _8216_;
wire _8217_;
wire _8218_;
wire _8219_;
wire _8220_;
wire _8221_;
wire _8222_;
wire _8223_;
wire _8224_;
wire _8225_;
wire _8226_;
wire _8227_;
wire _8228_;
wire _8229_;
wire _8230_;
wire _8231_;
wire _8232_;
wire _8233_;
wire _8234_;
wire _8235_;
wire _8236_;
wire _8237_;
wire _8238_;
wire _8239_;
wire _8240_;
wire _8241_;
wire _8242_;
wire _8243_;
wire _8244_;
wire _8245_;
wire _8246_;
wire _8247_;
wire _8248_;
wire _8249_;
wire _8250_;
wire _8251_;
wire _8252_;
wire _8253_;
wire _8254_;
wire _8255_;
wire _8256_;
wire _8257_;
wire _8258_;
wire _8259_;
wire _8260_;
wire _8261_;
wire _8262_;
wire _8263_;
wire _8264_;
wire _8265_;
wire _8266_;
wire _8267_;
wire _8268_;
wire _8269_;
wire _8270_;
wire _8271_;
wire _8272_;
wire _8273_;
wire _8274_;
wire _8275_;
wire _8276_;
wire _8277_;
wire _8278_;
wire _8279_;
wire _8280_;
wire _8281_;
wire _8282_;
wire _8283_;
wire _8284_;
wire _8285_;
wire _8286_;
wire _8287_;
wire _8288_;
wire _8289_;
wire _8290_;
wire _8291_;
wire _8292_;
wire _8293_;
wire _8294_;
wire _8295_;
wire _8296_;
wire _8297_;
wire _8298_;
wire _8299_;
wire _8300_;
wire _8301_;
wire _8302_;
wire _8303_;
wire _8304_;
wire _8305_;
wire _8306_;
wire _8307_;
wire _8308_;
wire _8309_;
wire _8310_;
wire _8311_;
wire _8312_;
wire _8313_;
wire _8314_;
wire _8315_;
wire _8316_;
wire _8317_;
wire _8318_;
wire _8319_;
wire _8320_;
wire _8321_;
wire _8322_;
wire _8323_;
wire _8324_;
wire _8325_;
wire _8326_;
wire _8327_;
wire _8328_;
wire _8329_;
wire _8330_;
wire _8331_;
wire _8332_;
wire _8333_;
wire _8334_;
wire _8335_;
wire _8336_;
wire _8337_;
wire _8338_;
wire _8339_;
wire _8340_;
wire _8341_;
wire _8342_;
wire _8343_;
wire _8344_;
wire _8345_;
wire _8346_;
wire _8347_;
wire _8348_;
wire _8349_;
wire _8350_;
wire _8351_;
wire _8352_;
wire _8353_;
wire _8354_;
wire _8355_;
wire _8356_;
wire _8357_;
wire _8358_;
wire _8359_;
wire _8360_;
wire _8361_;
wire _8362_;
wire _8363_;
wire _8364_;
wire _8365_;
wire _8366_;
wire _8367_;
wire _8368_;
wire _8369_;
wire _8370_;
wire _8371_;
wire _8372_;
wire _8373_;
wire _8374_;
wire _8375_;
wire _8376_;
wire _8377_;
wire _8378_;
wire _8379_;
wire _8380_;
wire _8381_;
wire _8382_;
wire _8383_;
wire _8384_;
wire _8385_;
wire _8386_;
wire _8387_;
wire _8388_;
wire _8389_;
wire _8390_;
wire _8391_;
wire _8392_;
wire _8393_;
wire _8394_;
wire _8395_;
wire _8396_;
wire _8397_;
wire _8398_;
wire _8399_;
wire _8400_;
wire _8401_;
wire _8402_;
wire _8403_;
wire _8404_;
wire _8405_;
wire _8406_;
wire _8407_;
wire _8408_;
wire _8409_;
wire _8410_;
wire _8411_;
wire _8412_;
wire _8413_;
wire _8414_;
wire _8415_;
wire _8416_;
wire _8417_;
wire _8418_;
wire _8419_;
wire _8420_;
wire _8421_;
wire _8422_;
wire _8423_;
wire _8424_;
wire _8425_;
wire _8426_;
wire _8427_;
wire _8428_;
wire _8429_;
wire _8430_;
wire _8431_;
wire _8432_;
wire _8433_;
wire _8434_;
wire _8435_;
wire _8436_;
wire _8437_;
wire _8438_;
wire _8439_;
wire _8440_;
wire _8441_;
wire _8442_;
wire _8443_;
wire _8444_;
wire _8445_;
wire _8446_;
wire _8447_;
wire _8448_;
wire _8449_;
wire _8450_;
wire _8451_;
wire _8452_;
wire _8453_;
wire _8454_;
wire _8455_;
wire _8456_;
wire _8457_;
wire _8458_;
wire _8459_;
wire _8460_;
wire _8461_;
wire _8462_;
wire _8463_;
wire _8464_;
wire _8465_;
wire _8466_;
wire _8467_;
wire _8468_;
wire _8469_;
wire _8470_;
wire _8471_;
wire _8472_;
wire _8473_;
wire _8474_;
wire _8475_;
wire _8476_;
wire _8477_;
wire _8478_;
wire _8479_;
wire _8480_;
wire _8481_;
wire _8482_;
wire _8483_;
wire _8484_;
wire _8485_;
wire _8486_;
wire _8487_;
wire _8488_;
wire _8489_;
wire _8490_;
wire _8491_;
wire _8492_;
wire _8493_;
wire _8494_;
wire _8495_;
wire _8496_;
wire _8497_;
wire _8498_;
wire _8499_;
wire _8500_;
wire _8501_;
wire _8502_;
wire _8503_;
wire _8504_;
wire _8505_;
wire _8506_;
wire _8507_;
wire _8508_;
wire _8509_;
wire _8510_;
wire _8511_;
wire _8512_;
wire _8513_;
wire _8514_;
wire _8515_;
wire _8516_;
wire _8517_;
wire _8518_;
wire _8519_;
wire _8520_;
wire _8521_;
wire _8522_;
wire _8523_;
wire _8524_;
wire _8525_;
wire _8526_;
wire _8527_;
wire _8528_;
wire _8529_;
wire _8530_;
wire _8531_;
wire _8532_;
wire _8533_;
wire _8534_;
wire _8535_;
wire _8536_;
wire _8537_;
wire _8538_;
wire _8539_;
wire _8540_;
wire _8541_;
wire _8542_;
wire _8543_;
wire _8544_;
wire _8545_;
wire _8546_;
wire _8547_;
wire _8548_;
wire _8549_;
wire _8550_;
wire _8551_;
wire _8552_;
wire _8553_;
wire _8554_;
wire _8555_;
wire _8556_;
wire _8557_;
wire _8558_;
wire _8559_;
wire _8560_;
wire _8561_;
wire _8562_;
wire _8563_;
wire _8564_;
wire _8565_;
wire _8566_;
wire _8567_;
wire _8568_;
wire _8569_;
wire _8570_;
wire _8571_;
wire _8572_;
wire _8573_;
wire _8574_;
wire _8575_;
wire _8576_;
wire _8577_;
wire _8578_;
wire _8579_;
wire _8580_;
wire _8581_;
wire _8582_;
wire _8583_;
wire _8584_;
wire _8585_;
wire _8586_;
wire _8587_;
wire _8588_;
wire _8589_;
wire _8590_;
wire _8591_;
wire _8592_;
wire _8593_;
wire _8594_;
wire _8595_;
wire _8596_;
wire _8597_;
wire _8598_;
wire _8599_;
wire _8600_;
wire _8601_;
wire _8602_;
wire _8603_;
wire _8604_;
wire _8605_;
wire _8606_;
wire _8607_;
wire _8608_;
wire _8609_;
wire _8610_;
wire _8611_;
wire _8612_;
wire _8613_;
wire _8614_;
wire _8615_;
wire _8616_;
wire _8617_;
wire _8618_;
wire _8619_;
wire _8620_;
wire _8621_;
wire _8622_;
wire _8623_;
wire _8624_;
wire _8625_;
wire _8626_;
wire _8627_;
wire _8628_;
wire _8629_;
wire _8630_;
wire _8631_;
wire _8632_;
wire _8633_;
wire _8634_;
wire _8635_;
wire _8636_;
wire _8637_;
wire _8638_;
wire _8639_;
wire _8640_;
wire _8641_;
wire _8642_;
wire _8643_;
wire _8644_;
wire _8645_;
wire _8646_;
wire _8647_;
wire _8648_;
wire _8649_;
wire _8650_;
wire _8651_;
wire _8652_;
wire _8653_;
wire _8654_;
wire _8655_;
wire _8656_;
wire _8657_;
wire _8658_;
wire _8659_;
wire _8660_;
wire _8661_;
wire _8662_;
wire _8663_;
wire _8664_;
wire _8665_;
wire _8666_;
wire _8667_;
wire _8668_;
wire _8669_;
wire _8670_;
wire _8671_;
wire _8672_;
wire _8673_;
wire _8674_;
wire _8675_;
wire _8676_;
wire _8677_;
wire _8678_;
wire _8679_;
wire _8680_;
wire _8681_;
wire _8682_;
wire _8683_;
wire _8684_;
wire _8685_;
wire _8686_;
wire _8687_;
wire _8688_;
wire _8689_;
wire _8690_;
wire _8691_;
wire _8692_;
wire _8693_;
wire _8694_;
wire _8695_;
wire _8696_;
wire _8697_;
wire _8698_;
wire _8699_;
wire _8700_;
wire _8701_;
wire _8702_;
wire _8703_;
wire _8704_;
wire _8705_;
wire _8706_;
wire _8707_;
wire _8708_;
wire _8709_;
wire _8710_;
wire _8711_;
wire _8712_;
wire _8713_;
wire _8714_;
wire _8715_;
wire _8716_;
wire _8717_;
wire _8718_;
wire _8719_;
wire _8720_;
wire _8721_;
wire _8722_;
wire _8723_;
wire _8724_;
wire _8725_;
wire _8726_;
wire _8727_;
wire _8728_;
wire _8729_;
wire _8730_;
wire _8731_;
wire _8732_;
wire _8733_;
wire _8734_;
wire _8735_;
wire _8736_;
wire _8737_;
wire _8738_;
wire _8739_;
wire _8740_;
wire _8741_;
wire _8742_;
wire _8743_;
wire _8744_;
wire _8745_;
wire _8746_;
wire _8747_;
wire _8748_;
wire _8749_;
wire _8750_;
wire _8751_;
wire _8752_;
wire _8753_;
wire _8754_;
wire _8755_;
wire _8756_;
wire _8757_;
wire _8758_;
wire _8759_;
wire _8760_;
wire _8761_;
wire _8762_;
wire _8763_;
wire _8764_;
wire _8765_;
wire _8766_;
wire _8767_;
wire _8768_;
wire _8769_;
wire _8770_;
wire _8771_;
wire _8772_;
wire _8773_;
wire _8774_;
wire _8775_;
wire _8776_;
wire _8777_;
wire _8778_;
wire _8779_;
wire _8780_;
wire _8781_;
wire _8782_;
wire _8783_;
wire _8784_;
wire _8785_;
wire _8786_;
wire _8787_;
wire _8788_;
wire _8789_;
wire _8790_;
wire _8791_;
wire _8792_;
wire _8793_;
wire _8794_;
wire _8795_;
wire _8796_;
wire _8797_;
wire _8798_;
wire _8799_;
wire _8800_;
wire _8801_;
wire _8802_;
wire _8803_;
wire _8804_;
wire _8805_;
wire _8806_;
wire _8807_;
wire _8808_;
wire _8809_;
wire _8810_;
wire _8811_;
wire _8812_;
wire _8813_;
wire _8814_;
wire _8815_;
wire _8816_;
wire _8817_;
wire _8818_;
wire _8819_;
wire _8820_;
wire _8821_;
wire _8822_;
wire _8823_;
wire _8824_;
wire _8825_;
wire _8826_;
wire _8827_;
wire _8828_;
wire _8829_;
wire _8830_;
wire _8831_;
wire _8832_;
wire _8833_;
wire _8834_;
wire _8835_;
wire _8836_;
wire _8837_;
wire _8838_;
wire _8839_;
wire _8840_;
wire _8841_;
wire _8842_;
wire _8843_;
wire _8844_;
wire _8845_;
wire _8846_;
wire _8847_;
wire _8848_;
wire _8849_;
wire _8850_;
wire _8851_;
wire _8852_;
wire _8853_;
wire _8854_;
wire _8855_;
wire _8856_;
wire _8857_;
wire _8858_;
wire _8859_;
wire _8860_;
wire _8861_;
wire _8862_;
wire _8863_;
wire _8864_;
wire _8865_;
wire _8866_;
wire _8867_;
wire _8868_;
wire _8869_;
wire _8870_;
wire _8871_;
wire _8872_;
wire _8873_;
wire _8874_;
wire _8875_;
wire _8876_;
wire _8877_;
wire _8878_;
wire _8879_;
wire _8880_;
wire _8881_;
wire _8882_;
wire _8883_;
wire _8884_;
wire _8885_;
wire _8886_;
wire _8887_;
wire _8888_;
wire _8889_;
wire _8890_;
wire _8891_;
wire _8892_;
wire _8893_;
wire _8894_;
wire _8895_;
wire _8896_;
wire _8897_;
wire _8898_;
wire _8899_;
wire _8900_;
wire _8901_;
wire _8902_;
wire _8903_;
wire _8904_;
wire _8905_;
wire _8906_;
wire _8907_;
wire _8908_;
wire _8909_;
wire _8910_;
wire _8911_;
wire _8912_;
wire _8913_;
wire _8914_;
wire _8915_;
wire _8916_;
wire _8917_;
wire _8918_;
wire _8919_;
wire _8920_;
wire _8921_;
wire _8922_;
wire _8923_;
wire _8924_;
wire _8925_;
wire _8926_;
wire _8927_;
wire _8928_;
wire _8929_;
wire _8930_;
wire _8931_;
wire _8932_;
wire _8933_;
wire _8934_;
wire _8935_;
wire _8936_;
wire _8937_;
wire _8938_;
wire _8939_;
wire _8940_;
wire _8941_;
wire _8942_;
wire _8943_;
wire _8944_;
wire _8945_;
wire _8946_;
wire _8947_;
wire _8948_;
wire _8949_;
wire _8950_;
wire _8951_;
wire _8952_;
wire _8953_;
wire _8954_;
wire _8955_;
wire _8956_;
wire _8957_;
wire _8958_;
wire _8959_;
wire _8960_;
wire _8961_;
wire _8962_;
wire _8963_;
wire _8964_;
wire _8965_;
wire _8966_;
wire _8967_;
wire _8968_;
wire _8969_;
wire _8970_;
wire _8971_;
wire _8972_;
wire _8973_;
wire _8974_;
wire _8975_;
wire _8976_;
wire _8977_;
wire _8978_;
wire _8979_;
wire _8980_;
wire _8981_;
wire _8982_;
wire _8983_;
wire _8984_;
wire _8985_;
wire _8986_;
wire _8987_;
wire _8988_;
wire _8989_;
wire _8990_;
wire _8991_;
wire _8992_;
wire _8993_;
wire _8994_;
wire _8995_;
wire _8996_;
wire _8997_;
wire _8998_;
wire _8999_;
wire _9000_;
wire _9001_;
wire _9002_;
wire _9003_;
wire _9004_;
wire _9005_;
wire _9006_;
wire _9007_;
wire _9008_;
wire _9009_;
wire _9010_;
wire _9011_;
wire _9012_;
wire _9013_;
wire _9014_;
wire _9015_;
wire _9016_;
wire _9017_;
wire _9018_;
wire _9019_;
wire _9020_;
wire _9021_;
wire _9022_;
wire _9023_;
wire _9024_;
wire _9025_;
wire _9026_;
wire _9027_;
wire _9028_;
wire _9029_;
wire _9030_;
wire _9031_;
wire _9032_;
wire _9033_;
wire _9034_;
wire _9035_;
wire _9036_;
wire _9037_;
wire _9038_;
wire _9039_;
wire _9040_;
wire _9041_;
wire _9042_;
wire _9043_;
wire _9044_;
wire _9045_;
wire _9046_;
wire _9047_;
wire _9048_;
wire _9049_;
wire _9050_;
wire _9051_;
wire _9052_;
wire _9053_;
wire _9054_;
wire _9055_;
wire _9056_;
wire _9057_;
wire _9058_;
wire _9059_;
wire _9060_;
wire _9061_;
wire _9062_;
wire _9063_;
wire _9064_;
wire _9065_;
wire _9066_;
wire _9067_;
wire _9068_;
wire _9069_;
wire _9070_;
wire _9071_;
wire _9072_;
wire _9073_;
wire _9074_;
wire _9075_;
wire _9076_;
wire _9077_;
wire _9078_;
wire _9079_;
wire _9080_;
wire _9081_;
wire _9082_;
wire _9083_;
wire _9084_;
wire _9085_;
wire _9086_;
wire _9087_;
wire _9088_;
wire _9089_;
wire _9090_;
wire _9091_;
wire _9092_;
wire _9093_;
wire _9094_;
wire _9095_;
wire _9096_;
wire _9097_;
wire _9098_;
wire _9099_;
wire _9100_;
wire _9101_;
wire _9102_;
wire _9103_;
wire _9104_;
wire _9105_;
wire _9106_;
wire _9107_;
wire _9108_;
wire _9109_;
wire _9110_;
wire _9111_;
wire _9112_;
wire _9113_;
wire _9114_;
wire _9115_;
wire _9116_;
wire _9117_;
wire _9118_;
wire _9119_;
wire _9120_;
wire _9121_;
wire _9122_;
wire _9123_;
wire _9124_;
wire _9125_;
wire _9126_;
wire _9127_;
wire _9128_;
wire _9129_;
wire _9130_;
wire _9131_;
wire _9132_;
wire _9133_;
wire _9134_;
wire _9135_;
wire _9136_;
wire _9137_;
wire _9138_;
wire _9139_;
wire _9140_;
wire _9141_;
wire _9142_;
wire _9143_;
wire _9144_;
wire _9145_;
wire _9146_;
wire _9147_;
wire _9148_;
wire _9149_;
wire _9150_;
wire _9151_;
wire _9152_;
wire _9153_;
wire _9154_;
wire _9155_;
wire _9156_;
wire _9157_;
wire _9158_;
wire _9159_;
wire _9160_;
wire _9161_;
wire _9162_;
wire _9163_;
wire _9164_;
wire _9165_;
wire _9166_;
wire _9167_;
wire _9168_;
wire _9169_;
wire _9170_;
wire _9171_;
wire _9172_;
wire _9173_;
wire _9174_;
wire _9175_;
wire _9176_;
wire _9177_;
wire _9178_;
wire _9179_;
wire _9180_;
wire _9181_;
wire _9182_;
wire _9183_;
wire _9184_;
wire _9185_;
wire _9186_;
wire _9187_;
wire _9188_;
wire _9189_;
wire _9190_;
wire _9191_;
wire _9192_;
wire _9193_;
wire _9194_;
wire _9195_;
wire _9196_;
wire _9197_;
wire _9198_;
wire _9199_;
wire _9200_;
wire _9201_;
wire _9202_;
wire _9203_;
wire _9204_;
wire _9205_;
wire _9206_;
wire _9207_;
wire _9208_;
wire _9209_;
wire _9210_;
wire _9211_;
wire _9212_;
wire _9213_;
wire _9214_;
wire _9215_;
wire _9216_;
wire _9217_;
wire _9218_;
wire _9219_;
wire _9220_;
wire _9221_;
wire _9222_;
wire _9223_;
wire _9224_;
wire _9225_;
wire _9226_;
wire _9227_;
wire _9228_;
wire _9229_;
wire _9230_;
wire _9231_;
wire _9232_;
wire _9233_;
wire _9234_;
wire _9235_;
wire _9236_;
wire _9237_;
wire _9238_;
wire _9239_;
wire _9240_;
wire _9241_;
wire _9242_;
wire _9243_;
wire _9244_;
wire _9245_;
wire _9246_;
wire _9247_;
wire _9248_;
wire _9249_;
wire _9250_;
wire _9251_;
wire _9252_;
wire _9253_;
wire _9254_;
wire _9255_;
wire _9256_;
wire _9257_;
wire _9258_;
wire _9259_;
wire _9260_;
wire _9261_;
wire _9262_;
wire _9263_;
wire _9264_;
wire _9265_;
wire _9266_;
wire _9267_;
wire _9268_;
wire _9269_;
wire _9270_;
wire _9271_;
wire _9272_;
wire _9273_;
wire _9274_;
wire _9275_;
wire _9276_;
wire _9277_;
wire _9278_;
wire _9279_;
wire _9280_;
wire _9281_;
wire _9282_;
wire _9283_;
wire _9284_;
wire _9285_;
wire _9286_;
wire _9287_;
wire _9288_;
wire _9289_;
wire _9290_;
wire _9291_;
wire _9292_;
wire _9293_;
wire _9294_;
wire _9295_;
wire _9296_;
wire _9297_;
wire _9298_;
wire _9299_;
wire _9300_;
wire _9301_;
wire _9302_;
wire _9303_;
wire _9304_;
wire _9305_;
wire _9306_;
wire _9307_;
wire _9308_;
wire _9309_;
wire _9310_;
wire _9311_;
wire _9312_;
wire _9313_;
wire _9314_;
wire _9315_;
wire _9316_;
wire _9317_;
wire _9318_;
wire _9319_;
wire _9320_;
wire _9321_;
wire _9322_;
wire _9323_;
wire _9324_;
wire _9325_;
wire _9326_;
wire _9327_;
wire _9328_;
wire _9329_;
wire _9330_;
wire _9331_;
wire _9332_;
wire _9333_;
wire _9334_;
wire _9335_;
wire _9336_;
wire _9337_;
wire _9338_;
wire _9339_;
wire _9340_;
wire _9341_;
wire _9342_;
wire _9343_;
wire _9344_;
wire _9345_;
wire _9346_;
wire _9347_;
wire _9348_;
wire _9349_;
wire _9350_;
wire _9351_;
wire _9352_;
wire _9353_;
wire _9354_;
wire _9355_;
wire _9356_;
wire _9357_;
wire _9358_;
wire _9359_;
wire _9360_;
wire _9361_;
wire _9362_;
wire _9363_;
wire _9364_;
wire _9365_;
wire _9366_;
wire _9367_;
wire _9368_;
wire _9369_;
wire _9370_;
wire _9371_;
wire _9372_;
wire _9373_;
wire _9374_;
wire _9375_;
wire _9376_;
wire _9377_;
wire _9378_;
wire _9379_;
wire _9380_;
wire _9381_;
wire _9382_;
wire _9383_;
wire _9384_;
wire _9385_;
wire _9386_;
wire _9387_;
wire _9388_;
wire _9389_;
wire _9390_;
wire _9391_;
wire _9392_;
wire _9393_;
wire _9394_;
wire _9395_;
wire _9396_;
wire _9397_;
wire _9398_;
wire _9399_;
wire _9400_;
wire _9401_;
wire _9402_;
wire _9403_;
wire _9404_;
wire _9405_;
wire _9406_;
wire _9407_;
wire _9408_;
wire _9409_;
wire _9410_;
wire _9411_;
wire _9412_;
wire _9413_;
wire _9414_;
wire _9415_;
wire _9416_;
wire _9417_;
wire _9418_;
wire _9419_;
wire _9420_;
wire _9421_;
wire _9422_;
wire _9423_;
wire _9424_;
wire _9425_;
wire _9426_;
wire _9427_;
wire _9428_;
wire _9429_;
wire _9430_;
wire _9431_;
wire _9432_;
wire _9433_;
wire _9434_;
wire _9435_;
wire _9436_;
wire _9437_;
wire _9438_;
wire _9439_;
wire _9440_;
wire _9441_;
wire _9442_;
wire _9443_;
wire _9444_;
wire _9445_;
wire _9446_;
wire _9447_;
wire _9448_;
wire _9449_;
wire _9450_;
wire _9451_;
wire _9452_;
wire _9453_;
wire _9454_;
wire _9455_;
wire _9456_;
wire _9457_;
wire _9458_;
wire _9459_;
wire _9460_;
wire _9461_;
wire _9462_;
wire _9463_;
wire _9464_;
wire _9465_;
wire _9466_;
wire _9467_;
wire _9468_;
wire _9469_;
wire _9470_;
wire _9471_;
wire _9472_;
wire _9473_;
wire _9474_;
wire _9475_;
wire _9476_;
wire _9477_;
wire _9478_;
wire _9479_;
wire _9480_;
wire _9481_;
wire _9482_;
wire _9483_;
wire _9484_;
wire _9485_;
wire _9486_;
wire _9487_;
wire _9488_;
wire _9489_;
wire _9490_;
wire _9491_;
wire _9492_;
wire _9493_;
wire _9494_;
wire _9495_;
wire _9496_;
wire _9497_;
wire _9498_;
wire _9499_;
wire _9500_;
wire _9501_;
wire _9502_;
wire _9503_;
wire _9504_;
wire _9505_;
wire _9506_;
wire _9507_;
wire _9508_;
wire _9509_;
wire _9510_;
wire _9511_;
wire _9512_;
wire _9513_;
wire _9514_;
wire _9515_;
wire _9516_;
wire _9517_;
wire _9518_;
wire _9519_;
wire _9520_;
wire _9521_;
wire _9522_;
wire _9523_;
wire _9524_;
wire _9525_;
wire _9526_;
wire _9527_;
wire _9528_;
wire _9529_;
wire _9530_;
wire _9531_;
wire _9532_;
wire _9533_;
wire _9534_;
wire _9535_;
wire _9536_;
wire _9537_;
wire _9538_;
wire _9539_;
wire _9540_;
wire _9541_;
wire _9542_;
wire _9543_;
wire _9544_;
wire _9545_;
wire _9546_;
wire _9547_;
wire _9548_;
wire _9549_;
wire _9550_;
wire _9551_;
wire _9552_;
wire _9553_;
wire _9554_;
wire _9555_;
wire _9556_;
wire _9557_;
wire _9558_;
wire _9559_;
wire _9560_;
wire _9561_;
wire _9562_;
wire _9563_;
wire _9564_;
wire _9565_;
wire _9566_;
wire _9567_;
wire _9568_;
wire _9569_;
wire _9570_;
wire _9571_;
wire _9572_;
wire _9573_;
wire _9574_;
wire _9575_;
wire _9576_;
wire _9577_;
wire _9578_;
wire _9579_;
wire _9580_;
wire _9581_;
wire _9582_;
wire _9583_;
wire _9584_;
wire _9585_;
wire _9586_;
wire _9587_;
wire _9588_;
wire _9589_;
wire _9590_;
wire _9591_;
wire _9592_;
wire _9593_;
wire _9594_;
wire _9595_;
wire _9596_;
wire _9597_;
wire _9598_;
wire _9599_;
wire _9600_;
wire _9601_;
wire _9602_;
wire _9603_;
wire _9604_;
wire _9605_;
wire _9606_;
wire _9607_;
wire _9608_;
wire _9609_;
wire _9610_;
wire _9611_;
wire _9612_;
wire _9613_;
wire _9614_;
wire _9615_;
wire _9616_;
wire _9617_;
wire _9618_;
wire _9619_;
wire _9620_;
wire _9621_;
wire _9622_;
wire _9623_;
wire _9624_;
wire _9625_;
wire _9626_;
wire _9627_;
wire _9628_;
wire _9629_;
wire _9630_;
wire _9631_;
wire _9632_;
wire _9633_;
wire _9634_;
wire _9635_;
wire _9636_;
wire _9637_;
wire _9638_;
wire _9639_;
wire _9640_;
wire _9641_;
wire _9642_;
wire _9643_;
wire _9644_;
wire _9645_;
wire _9646_;
wire _9647_;
wire _9648_;
wire _9649_;
wire _9650_;
wire _9651_;
wire _9652_;
wire _9653_;
wire _9654_;
wire _9655_;
wire _9656_;
wire _9657_;
wire _9658_;
wire _9659_;
wire _9660_;
wire _9661_;
wire _9662_;
wire _9663_;
wire _9664_;
wire _9665_;
wire _9666_;
wire _9667_;
wire _9668_;
wire _9669_;
wire _9670_;
wire _9671_;
wire _9672_;
wire _9673_;
wire _9674_;
wire _9675_;
wire _9676_;
wire _9677_;
wire _9678_;
wire _9679_;
wire _9680_;
wire _9681_;
wire _9682_;
wire _9683_;
wire _9684_;
wire _9685_;
wire _9686_;
wire _9687_;
wire _9688_;
wire _9689_;
wire _9690_;
wire _9691_;
wire _9692_;
wire _9693_;
wire _9694_;
wire _9695_;
wire _9696_;
wire _9697_;
wire _9698_;
wire _9699_;
wire _9700_;
wire _9701_;
wire _9702_;
wire _9703_;
wire _9704_;
wire _9705_;
wire _9706_;
wire _9707_;
wire _9708_;
wire _9709_;
wire _9710_;
wire _9711_;
wire _9712_;
wire _9713_;
wire _9714_;
wire _9715_;
wire _9716_;
wire _9717_;
wire _9718_;
wire _9719_;
wire _9720_;
wire _9721_;
wire _9722_;
wire _9723_;
wire _9724_;
wire _9725_;
wire _9726_;
wire _9727_;
wire _9728_;
wire _9729_;
wire _9730_;
wire _9731_;
wire _9732_;
wire _9733_;
wire _9734_;
wire _9735_;
wire _9736_;
wire _9737_;
wire _9738_;
wire _9739_;
wire _9740_;
wire _9741_;
wire _9742_;
wire _9743_;
wire _9744_;
wire _9745_;
wire _9746_;
wire _9747_;
wire _9748_;
wire _9749_;
wire _9750_;
wire _9751_;
wire _9752_;
wire _9753_;
wire _9754_;
wire _9755_;
wire _9756_;
wire _9757_;
wire _9758_;
wire _9759_;
wire _9760_;
wire _9761_;
wire _9762_;
wire _9763_;
wire _9764_;
wire _9765_;
wire _9766_;
wire _9767_;
wire _9768_;
wire _9769_;
wire _9770_;
wire _9771_;
wire _9772_;
wire _9773_;
wire _9774_;
wire _9775_;
wire _9776_;
wire _9777_;
wire _9778_;
wire _9779_;
wire _9780_;
wire _9781_;
wire _9782_;
wire _9783_;
wire _9784_;
wire _9785_;
wire _9786_;
wire _9787_;
wire _9788_;
wire _9789_;
wire _9790_;
wire _9791_;
wire _9792_;
wire _9793_;
wire _9794_;
wire _9795_;
wire _9796_;
wire _9797_;
wire _9798_;
wire _9799_;
wire _9800_;
wire _9801_;
wire _9802_;
wire _9803_;
wire _9804_;
wire _9805_;
wire _9806_;
wire _9807_;
wire _9808_;
wire _9809_;
wire _9810_;
wire _9811_;
wire _9812_;
wire _9813_;
wire _9814_;
wire _9815_;
wire _9816_;
wire _9817_;
wire _9818_;
wire _9819_;
wire _9820_;
wire _9821_;
wire _9822_;
wire _9823_;
wire _9824_;
wire _9825_;
wire _9826_;
wire _9827_;
wire _9828_;
wire _9829_;
wire _9830_;
wire _9831_;
wire _9832_;
wire _9833_;
wire _9834_;
wire _9835_;
wire _9836_;
wire _9837_;
wire _9838_;
wire _9839_;
wire _9840_;
wire _9841_;
wire _9842_;
wire _9843_;
wire _9844_;
wire _9845_;
wire _9846_;
wire _9847_;
wire _9848_;
wire _9849_;
wire _9850_;
wire _9851_;
wire _9852_;
wire _9853_;
wire _9854_;
wire _9855_;
wire _9856_;
wire _9857_;
wire _9858_;
wire _9859_;
wire _9860_;
wire _9861_;
wire _9862_;
wire _9863_;
wire _9864_;
wire _9865_;
wire _9866_;
wire _9867_;
wire _9868_;
wire _9869_;
wire _9870_;
wire _9871_;
wire _9872_;
wire _9873_;
wire _9874_;
wire _9875_;
wire _9876_;
wire _9877_;
wire _9878_;
wire _9879_;
wire _9880_;
wire _9881_;
wire _9882_;
wire _9883_;
wire _9884_;
wire _9885_;
wire _9886_;
wire _9887_;
wire _9888_;
wire _9889_;
wire _9890_;
wire _9891_;
wire _9892_;
wire _9893_;
wire _9894_;
wire _9895_;
wire _9896_;
wire _9897_;
wire _9898_;
wire _9899_;
wire _9900_;
wire _9901_;
wire _9902_;
wire _9903_;
wire _9904_;
wire _9905_;
wire _9906_;
wire _9907_;
wire _9908_;
wire _9909_;
wire _9910_;
wire _9911_;
wire _9912_;
wire _9913_;
wire _9914_;
wire _9915_;
wire _9916_;
wire _9917_;
wire _9918_;
wire _9919_;
wire _9920_;
wire _9921_;
wire _9922_;
wire _9923_;
wire _9924_;
wire _9925_;
wire _9926_;
wire _9927_;
wire _9928_;
wire _9929_;
wire _9930_;
wire _9931_;
wire _9932_;
wire _9933_;
wire _9934_;
wire _9935_;
wire _9936_;
wire _9937_;
wire _9938_;
wire _9939_;
wire _9940_;
wire _9941_;
wire _9942_;
wire _9943_;
wire _9944_;
wire _9945_;
wire _9946_;
wire _9947_;
wire _9948_;
wire _9949_;
wire _9950_;
wire _9951_;
wire _9952_;
wire _9953_;
wire _9954_;
wire _9955_;
wire _9956_;
wire _9957_;
wire _9958_;
wire _9959_;
wire _9960_;
wire _9961_;
wire _9962_;
wire _9963_;
wire _9964_;
wire _9965_;
wire _9966_;
wire _9967_;
wire _9968_;
wire _9969_;
wire _9970_;
wire _9971_;
wire _9972_;
wire _9973_;
wire _9974_;
wire _9975_;
wire _9976_;
wire _9977_;
wire _9978_;
wire _9979_;
wire _9980_;
wire _9981_;
wire _9982_;
wire _9983_;
wire _9984_;
wire _9985_;
wire _9986_;
wire _9987_;
wire _9988_;
wire _9989_;
wire _9990_;
wire _9991_;
wire _9992_;
wire _9993_;
wire _9994_;
wire _9995_;
wire _9996_;
wire _9997_;
wire _9998_;
wire _9999_;
wire _10000_;
wire _10001_;
wire _10002_;
wire _10003_;
wire _10004_;
wire _10005_;
wire _10006_;
wire _10007_;
wire _10008_;
wire _10009_;
wire _10010_;
wire _10011_;
wire _10012_;
wire _10013_;
wire _10014_;
wire _10015_;
wire _10016_;
wire _10017_;
wire _10018_;
wire _10019_;
wire _10020_;
wire _10021_;
wire _10022_;
wire _10023_;
wire _10024_;
wire _10025_;
wire _10026_;
wire _10027_;
wire _10028_;
wire _10029_;
wire _10030_;
wire _10031_;
wire _10032_;
wire _10033_;
wire _10034_;
wire _10035_;
wire _10036_;
wire _10037_;
wire _10038_;
wire _10039_;
wire _10040_;
wire _10041_;
wire _10042_;
wire _10043_;
wire _10044_;
wire _10045_;
wire _10046_;
wire _10047_;
wire _10048_;
wire _10049_;
wire _10050_;
wire _10051_;
wire _10052_;
wire _10053_;
wire _10054_;
wire _10055_;
wire _10056_;
wire _10057_;
wire _10058_;
wire _10059_;
wire _10060_;
wire _10061_;
wire _10062_;
wire _10063_;
wire _10064_;
wire _10065_;
wire _10066_;
wire _10067_;
wire _10068_;
wire _10069_;
wire _10070_;
wire _10071_;
wire _10072_;
wire _10073_;
wire _10074_;
wire _10075_;
wire _10076_;
wire _10077_;
wire _10078_;
wire _10079_;
wire _10080_;
wire _10081_;
wire _10082_;
wire _10083_;
wire _10084_;
wire _10085_;
wire _10086_;
wire _10087_;
wire _10088_;
wire _10089_;
wire _10090_;
wire _10091_;
wire _10092_;
wire _10093_;
wire _10094_;
wire _10095_;
wire _10096_;
wire _10097_;
wire _10098_;
wire _10099_;
wire _10100_;
wire _10101_;
wire _10102_;
wire _10103_;
wire _10104_;
wire _10105_;
wire _10106_;
wire _10107_;
wire _10108_;
wire _10109_;
wire _10110_;
wire _10111_;
wire _10112_;
wire _10113_;
wire _10114_;
wire _10115_;
wire _10116_;
wire _10117_;
wire _10118_;
wire _10119_;
wire _10120_;
wire _10121_;
wire _10122_;
wire _10123_;
wire _10124_;
wire _10125_;
wire _10126_;
wire _10127_;
wire _10128_;
wire _10129_;
wire _10130_;
wire _10131_;
wire _10132_;
wire _10133_;
wire _10134_;
wire _10135_;
wire _10136_;
wire _10137_;
wire _10138_;
wire _10139_;
wire _10140_;
wire _10141_;
wire _10142_;
wire _10143_;
wire _10144_;
wire _10145_;
wire _10146_;
wire _10147_;
wire _10148_;
wire _10149_;
wire _10150_;
wire _10151_;
wire _10152_;
wire _10153_;
wire _10154_;
wire _10155_;
wire _10156_;
wire _10157_;
wire _10158_;
wire _10159_;
wire _10160_;
wire _10161_;
wire _10162_;
wire _10163_;
wire _10164_;
wire _10165_;
wire _10166_;
wire _10167_;
wire _10168_;
wire _10169_;
wire _10170_;
wire _10171_;
wire _10172_;
wire _10173_;
wire _10174_;
wire _10175_;
wire _10176_;
wire _10177_;
wire _10178_;
wire _10179_;
wire _10180_;
wire _10181_;
wire _10182_;
wire _10183_;
wire _10184_;
wire _10185_;
wire _10186_;
wire _10187_;
wire _10188_;
wire _10189_;
wire _10190_;
wire _10191_;
wire _10192_;
wire _10193_;
wire _10194_;
wire _10195_;
wire _10196_;
wire _10197_;
wire _10198_;
wire _10199_;
wire _10200_;
wire _10201_;
wire _10202_;
wire _10203_;
wire _10204_;
wire _10205_;
wire _10206_;
wire _10207_;
wire _10208_;
wire _10209_;
wire _10210_;
wire _10211_;
wire _10212_;
wire _10213_;
wire _10214_;
wire _10215_;
wire _10216_;
wire _10217_;
wire _10218_;
wire _10219_;
wire _10220_;
wire _10221_;
wire _10222_;
wire _10223_;
wire _10224_;
wire _10225_;
wire _10226_;
wire _10227_;
wire _10228_;
wire _10229_;
wire _10230_;
wire _10231_;
wire _10232_;
wire _10233_;
wire _10234_;
wire _10235_;
wire _10236_;
wire _10237_;
wire _10238_;
wire _10239_;
wire _10240_;
wire _10241_;
wire _10242_;
wire _10243_;
wire _10244_;
wire _10245_;
wire _10246_;
wire _10247_;
wire _10248_;
wire _10249_;
wire _10250_;
wire _10251_;
wire _10252_;
wire _10253_;
wire _10254_;
wire _10255_;
wire _10256_;
wire _10257_;
wire _10258_;
wire _10259_;
wire _10260_;
wire _10261_;
wire _10262_;
wire _10263_;
wire _10264_;
wire _10265_;
wire _10266_;
wire _10267_;
wire _10268_;
wire _10269_;
wire _10270_;
wire _10271_;
wire _10272_;
wire _10273_;
wire _10274_;
wire _10275_;
wire _10276_;
wire _10277_;
wire _10278_;
wire _10279_;
wire _10280_;
wire _10281_;
wire _10282_;
wire _10283_;
wire _10284_;
wire _10285_;
wire _10286_;
wire _10287_;
wire _10288_;
wire _10289_;
wire _10290_;
wire _10291_;
wire _10292_;
wire _10293_;
wire _10294_;
wire _10295_;
wire _10296_;
wire _10297_;
wire _10298_;
wire _10299_;
wire _10300_;
wire _10301_;
wire _10302_;
wire _10303_;
wire _10304_;
wire _10305_;
wire _10306_;
wire _10307_;
wire _10308_;
wire _10309_;
wire _10310_;
wire _10311_;
wire _10312_;
wire _10313_;
wire _10314_;
wire _10315_;
wire _10316_;
wire _10317_;
wire _10318_;
wire _10319_;
wire _10320_;
wire _10321_;
wire _10322_;
wire _10323_;
wire _10324_;
wire _10325_;
wire _10326_;
wire _10327_;
wire _10328_;
wire _10329_;
wire _10330_;
wire _10331_;
wire _10332_;
wire _10333_;
wire _10334_;
wire _10335_;
wire _10336_;
wire _10337_;
wire _10338_;
wire _10339_;
wire _10340_;
wire _10341_;
wire _10342_;
wire _10343_;
wire _10344_;
wire _10345_;
wire _10346_;
wire _10347_;
wire _10348_;
wire _10349_;
wire _10350_;
wire _10351_;
wire _10352_;
wire _10353_;
wire _10354_;
wire _10355_;
wire _10356_;
wire _10357_;
wire _10358_;
wire _10359_;
wire _10360_;
wire _10361_;
wire _10362_;
wire _10363_;
wire _10364_;
wire _10365_;
wire _10366_;
wire _10367_;
wire _10368_;
wire _10369_;
wire _10370_;
wire _10371_;
wire _10372_;
wire _10373_;
wire _10374_;
wire _10375_;
wire _10376_;
wire _10377_;
wire _10378_;
wire _10379_;
wire _10380_;
wire _10381_;
wire _10382_;
wire _10383_;
wire _10384_;
wire _10385_;
wire _10386_;
wire _10387_;
wire _10388_;
wire _10389_;
wire _10390_;
wire _10391_;
wire _10392_;
wire _10393_;
wire _10394_;
wire _10395_;
wire _10396_;
wire _10397_;
wire _10398_;
wire _10399_;
wire _10400_;
wire _10401_;
wire _10402_;
wire _10403_;
wire _10404_;
wire _10405_;
wire _10406_;
wire _10407_;
wire _10408_;
wire _10409_;
wire _10410_;
wire _10411_;
wire _10412_;
wire _10413_;
wire _10414_;
wire _10415_;
wire _10416_;
wire _10417_;
wire _10418_;
wire _10419_;
wire _10420_;
wire _10421_;
wire _10422_;
wire _10423_;
wire _10424_;
wire _10425_;
wire _10426_;
wire _10427_;
wire _10428_;
wire _10429_;
wire _10430_;
wire _10431_;
wire _10432_;
wire _10433_;
wire _10434_;
wire _10435_;
wire _10436_;
wire _10437_;
wire _10438_;
wire _10439_;
wire _10440_;
wire _10441_;
wire _10442_;
wire _10443_;
wire _10444_;
wire _10445_;
wire _10446_;
wire _10447_;
wire _10448_;
wire _10449_;
wire _10450_;
wire _10451_;
wire _10452_;
wire _10453_;
wire _10454_;
wire _10455_;
wire _10456_;
wire _10457_;
wire _10458_;
wire _10459_;
wire _10460_;
wire _10461_;
wire _10462_;
wire _10463_;
wire _10464_;
wire _10465_;
wire _10466_;
wire _10467_;
wire _10468_;
wire _10469_;
wire _10470_;
wire _10471_;
wire _10472_;
wire _10473_;
wire _10474_;
wire _10475_;
wire _10476_;
wire _10477_;
wire _10478_;
wire _10479_;
wire _10480_;
wire _10481_;
wire _10482_;
wire _10483_;
wire _10484_;
wire _10485_;
wire _10486_;
wire _10487_;
wire _10488_;
wire _10489_;
wire _10490_;
wire _10491_;
wire _10492_;
wire _10493_;
wire _10494_;
wire _10495_;
wire _10496_;
wire _10497_;
wire _10498_;
wire _10499_;
wire _10500_;
wire _10501_;
wire _10502_;
wire _10503_;
wire _10504_;
wire _10505_;
wire _10506_;
wire _10507_;
wire _10508_;
wire _10509_;
wire _10510_;
wire _10511_;
wire _10512_;
wire _10513_;
wire _10514_;
wire _10515_;
wire _10516_;
wire _10517_;
wire _10518_;
wire _10519_;
wire _10520_;
wire _10521_;
wire _10522_;
wire _10523_;
wire _10524_;
wire _10525_;
wire _10526_;
wire _10527_;
wire _10528_;
wire _10529_;
wire _10530_;
wire _10531_;
wire _10532_;
wire _10533_;
wire _10534_;
wire _10535_;
wire _10536_;
wire _10537_;
wire _10538_;
wire _10539_;
wire _10540_;
wire _10541_;
wire _10542_;
wire _10543_;
wire _10544_;
wire _10545_;
wire _10546_;
wire _10547_;
wire _10548_;
wire _10549_;
wire _10550_;
wire _10551_;
wire _10552_;
wire _10553_;
wire _10554_;
wire _10555_;
wire _10556_;
wire _10557_;
wire _10558_;
wire _10559_;
wire _10560_;
wire _10561_;
wire _10562_;
wire _10563_;
wire _10564_;
wire _10565_;
wire _10566_;
wire _10567_;
wire _10568_;
wire _10569_;
wire _10570_;
wire _10571_;
wire _10572_;
wire _10573_;
wire _10574_;
wire _10575_;
wire _10576_;
wire _10577_;
wire _10578_;
wire _10579_;
wire _10580_;
wire _10581_;
wire _10582_;
wire _10583_;
wire _10584_;
wire _10585_;
wire _10586_;
wire _10587_;
wire _10588_;
wire _10589_;
wire _10590_;
wire _10591_;
wire _10592_;
wire _10593_;
wire _10594_;
wire _10595_;
wire _10596_;
wire _10597_;
wire _10598_;
wire _10599_;
wire _10600_;
wire _10601_;
wire _10602_;
wire _10603_;
wire _10604_;
wire _10605_;
wire _10606_;
wire _10607_;
wire _10608_;
wire _10609_;
wire _10610_;
wire _10611_;
wire _10612_;
wire _10613_;
wire _10614_;
wire _10615_;
wire _10616_;
wire _10617_;
wire _10618_;
wire _10619_;
wire _10620_;
wire _10621_;
wire _10622_;
wire _10623_;
wire _10624_;
wire _10625_;
wire _10626_;
wire _10627_;
wire _10628_;
wire _10629_;
wire _10630_;
wire _10631_;
wire _10632_;
wire _10633_;
wire _10634_;
wire _10635_;
wire _10636_;
wire _10637_;
wire _10638_;
wire _10639_;
wire _10640_;
wire _10641_;
wire _10642_;
wire _10643_;
wire _10644_;
wire _10645_;
wire _10646_;
wire _10647_;
wire _10648_;
wire _10649_;
wire _10650_;
wire _10651_;
wire _10652_;
wire _10653_;
wire _10654_;
wire _10655_;
wire _10656_;
wire _10657_;
wire _10658_;
wire _10659_;
wire _10660_;
wire _10661_;
wire _10662_;
wire _10663_;
wire _10664_;
wire _10665_;
wire _10666_;
wire _10667_;
wire _10668_;
wire _10669_;
wire _10670_;
wire _10671_;
wire _10672_;
wire _10673_;
wire _10674_;
wire _10675_;
wire _10676_;
wire _10677_;
wire _10678_;
wire _10679_;
wire _10680_;
wire _10681_;
wire _10682_;
wire _10683_;
wire _10684_;
wire _10685_;
wire _10686_;
wire _10687_;
wire _10688_;
wire _10689_;
wire _10690_;
wire _10691_;
wire _10692_;
wire _10693_;
wire _10694_;
wire _10695_;
wire _10696_;
wire _10697_;
wire _10698_;
wire _10699_;
wire _10700_;
wire _10701_;
wire _10702_;
wire _10703_;
wire _10704_;
wire _10705_;
wire _10706_;
wire _10707_;
wire _10708_;
wire _10709_;
wire _10710_;
wire _10711_;
wire _10712_;
wire _10713_;
wire _10714_;
wire _10715_;
wire _10716_;
wire _10717_;
wire _10718_;
wire _10719_;
wire _10720_;
wire _10721_;
wire _10722_;
wire _10723_;
wire _10724_;
wire _10725_;
wire _10726_;
wire _10727_;
wire _10728_;
wire _10729_;
wire _10730_;
wire _10731_;
wire _10732_;
wire _10733_;
wire _10734_;
wire _10735_;
wire _10736_;
wire _10737_;
wire _10738_;
wire _10739_;
wire _10740_;
wire _10741_;
wire _10742_;
wire _10743_;
wire _10744_;
wire _10745_;
wire _10746_;
wire _10747_;
wire _10748_;
wire _10749_;
wire _10750_;
wire _10751_;
wire _10752_;
wire _10753_;
wire _10754_;
wire _10755_;
wire _10756_;
wire _10757_;
wire _10758_;
wire _10759_;
wire _10760_;
wire _10761_;
wire _10762_;
wire _10763_;
wire _10764_;
wire _10765_;
wire _10766_;
wire _10767_;
wire _10768_;
wire _10769_;
wire _10770_;
wire _10771_;
wire _10772_;
wire _10773_;
wire _10774_;
wire _10775_;
wire _10776_;
wire _10777_;
wire _10778_;
wire _10779_;
wire _10780_;
wire _10781_;
wire _10782_;
wire _10783_;
wire _10784_;
wire _10785_;
wire _10786_;
wire _10787_;
wire _10788_;
wire _10789_;
wire _10790_;
wire _10791_;
wire _10792_;
wire _10793_;
wire _10794_;
wire _10795_;
wire _10796_;
wire _10797_;
wire _10798_;
wire _10799_;
wire _10800_;
wire _10801_;
wire _10802_;
wire _10803_;
wire _10804_;
wire _10805_;
wire _10806_;
wire _10807_;
wire _10808_;
wire _10809_;
wire _10810_;
wire _10811_;
wire _10812_;
wire _10813_;
wire _10814_;
wire _10815_;
wire _10816_;
wire _10817_;
wire _10818_;
wire _10819_;
wire _10820_;
wire _10821_;
wire _10822_;
wire _10823_;
wire _10824_;
wire _10825_;
wire _10826_;
wire _10827_;
wire _10828_;
wire _10829_;
wire _10830_;
wire _10831_;
wire _10832_;
wire _10833_;
wire _10834_;
wire _10835_;
wire _10836_;
wire _10837_;
wire _10838_;
wire _10839_;
wire _10840_;
wire _10841_;
wire _10842_;
wire _10843_;
wire _10844_;
wire _10845_;
wire _10846_;
wire _10847_;
wire _10848_;
wire _10849_;
wire _10850_;
wire _10851_;
wire _10852_;
wire _10853_;
wire _10854_;
wire _10855_;
wire _10856_;
wire _10857_;
wire _10858_;
wire _10859_;
wire _10860_;
wire _10861_;
wire _10862_;
wire _10863_;
wire _10864_;
wire _10865_;
wire _10866_;
wire _10867_;
wire _10868_;
wire _10869_;
wire _10870_;
wire _10871_;
wire _10872_;
wire _10873_;
wire _10874_;
wire _10875_;
wire _10876_;
wire _10877_;
wire _10878_;
wire _10879_;
wire _10880_;
wire _10881_;
wire _10882_;
wire _10883_;
wire _10884_;
wire _10885_;
wire _10886_;
wire _10887_;
wire _10888_;
wire _10889_;
wire _10890_;
wire _10891_;
wire _10892_;
wire _10893_;
wire _10894_;
wire _10895_;
wire _10896_;
wire _10897_;
wire _10898_;
wire _10899_;
wire _10900_;
wire _10901_;
wire _10902_;
wire _10903_;
wire _10904_;
wire _10905_;
wire _10906_;
wire _10907_;
wire _10908_;
wire _10909_;
wire _10910_;
wire _10911_;
wire _10912_;
wire _10913_;
wire _10914_;
wire _10915_;
wire _10916_;
wire _10917_;
wire _10918_;
wire _10919_;
wire _10920_;
wire _10921_;
wire _10922_;
wire _10923_;
wire _10924_;
wire _10925_;
wire _10926_;
wire _10927_;
wire _10928_;
wire _10929_;
wire _10930_;
wire _10931_;
wire _10932_;
wire _10933_;
wire _10934_;
wire _10935_;
wire _10936_;
wire _10937_;
wire _10938_;
wire _10939_;
wire _10940_;
wire _10941_;
wire _10942_;
wire _10943_;
wire _10944_;
wire _10945_;
wire _10946_;
wire _10947_;
wire _10948_;
wire _10949_;
wire _10950_;
wire _10951_;
wire _10952_;
wire _10953_;
wire _10954_;
wire _10955_;
wire _10956_;
wire _10957_;
wire _10958_;
wire _10959_;
wire _10960_;
wire _10961_;
wire _10962_;
wire _10963_;
wire _10964_;
wire _10965_;
wire _10966_;
wire _10967_;
wire _10968_;
wire _10969_;
wire _10970_;
wire _10971_;
wire _10972_;
wire _10973_;
wire _10974_;
wire _10975_;
wire _10976_;
wire _10977_;
wire _10978_;
wire _10979_;
wire _10980_;
wire _10981_;
wire _10982_;
wire _10983_;
wire _10984_;
wire _10985_;
wire _10986_;
wire _10987_;
wire _10988_;
wire _10989_;
wire _10990_;
wire _10991_;
wire _10992_;
wire _10993_;
wire _10994_;
wire _10995_;
wire _10996_;
wire _10997_;
wire _10998_;
wire _10999_;
wire _11000_;
wire _11001_;
wire _11002_;
wire _11003_;
wire _11004_;
wire _11005_;
wire _11006_;
wire _11007_;
wire _11008_;
wire _11009_;
wire _11010_;
wire _11011_;
wire _11012_;
wire _11013_;
wire _11014_;
wire _11015_;
wire _11016_;
wire _11017_;
wire _11018_;
wire _11019_;
wire _11020_;
wire _11021_;
wire _11022_;
wire _11023_;
wire _11024_;
wire _11025_;
wire _11026_;
wire _11027_;
wire _11028_;
wire _11029_;
wire _11030_;
wire _11031_;
wire _11032_;
wire _11033_;
wire _11034_;
wire _11035_;
wire _11036_;
wire _11037_;
wire _11038_;
wire _11039_;
wire _11040_;
wire _11041_;
wire _11042_;
wire _11043_;
wire _11044_;
wire _11045_;
wire _11046_;
wire _11047_;
wire _11048_;
wire _11049_;
wire _11050_;
wire _11051_;
wire _11052_;
wire _11053_;
wire _11054_;
wire _11055_;
wire _11056_;
wire _11057_;
wire _11058_;
wire _11059_;
wire _11060_;
wire _11061_;
wire _11062_;
wire _11063_;
wire _11064_;
wire _11065_;
wire _11066_;
wire _11067_;
wire _11068_;
wire _11069_;
wire _11070_;
wire _11071_;
wire _11072_;
wire _11073_;
wire _11074_;
wire _11075_;
wire _11076_;
wire _11077_;
wire _11078_;
wire _11079_;
wire _11080_;
wire _11081_;
wire _11082_;
wire _11083_;
wire _11084_;
wire _11085_;
wire _11086_;
wire _11087_;
wire _11088_;
wire _11089_;
wire _11090_;
wire _11091_;
wire _11092_;
wire _11093_;
wire _11094_;
wire _11095_;
wire _11096_;
wire _11097_;
wire _11098_;
wire _11099_;
wire _11100_;
wire _11101_;
wire _11102_;
wire _11103_;
wire _11104_;
wire _11105_;
wire _11106_;
wire _11107_;
wire _11108_;
wire _11109_;
wire _11110_;
wire _11111_;
wire _11112_;
wire _11113_;
wire _11114_;
wire _11115_;
wire _11116_;
wire _11117_;
wire _11118_;
wire _11119_;
wire _11120_;
wire _11121_;
wire _11122_;
wire _11123_;
wire _11124_;
wire _11125_;
wire _11126_;
wire _11127_;
wire _11128_;
wire _11129_;
wire _11130_;
wire _11131_;
wire _11132_;
wire _11133_;
wire _11134_;
wire _11135_;
wire _11136_;
wire _11137_;
wire _11138_;
wire _11139_;
wire _11140_;
wire _11141_;
wire _11142_;
wire _11143_;
wire _11144_;
wire _11145_;
wire _11146_;
wire _11147_;
wire _11148_;
wire _11149_;
wire _11150_;
wire _11151_;
wire _11152_;
wire _11153_;
wire _11154_;
wire _11155_;
wire _11156_;
wire _11157_;
wire _11158_;
wire _11159_;
wire _11160_;
wire _11161_;
wire _11162_;
wire _11163_;
wire _11164_;
wire _11165_;
wire _11166_;
wire _11167_;
wire _11168_;
wire _11169_;
wire _11170_;
wire _11171_;
wire _11172_;
wire _11173_;
wire _11174_;
wire _11175_;
wire _11176_;
wire _11177_;
wire _11178_;
wire _11179_;
wire _11180_;
wire _11181_;
wire _11182_;
wire _11183_;
wire _11184_;
wire _11185_;
wire _11186_;
wire _11187_;
wire _11188_;
wire _11189_;
wire _11190_;
wire _11191_;
wire _11192_;
wire _11193_;
wire _11194_;
wire _11195_;
wire _11196_;
wire _11197_;
wire _11198_;
wire _11199_;
wire _11200_;
wire _11201_;
wire _11202_;
wire _11203_;
wire _11204_;
wire _11205_;
wire _11206_;
wire _11207_;
wire _11208_;
wire _11209_;
wire _11210_;
wire _11211_;
wire _11212_;
wire _11213_;
wire _11214_;
wire _11215_;
wire _11216_;
wire _11217_;
wire _11218_;
wire _11219_;
wire _11220_;
wire _11221_;
wire _11222_;
wire _11223_;
wire _11224_;
wire _11225_;
wire _11226_;
wire _11227_;
wire _11228_;
wire _11229_;
wire _11230_;
wire _11231_;
wire _11232_;
wire _11233_;
wire _11234_;
wire _11235_;
wire _11236_;
wire _11237_;
wire _11238_;
wire _11239_;
wire _11240_;
wire _11241_;
wire _11242_;
wire _11243_;
wire _11244_;
wire _11245_;
wire _11246_;
wire _11247_;
wire _11248_;
wire _11249_;
wire _11250_;
wire _11251_;
wire _11252_;
wire _11253_;
wire _11254_;
wire _11255_;
wire _11256_;
wire _11257_;
wire _11258_;
wire _11259_;
wire _11260_;
wire _11261_;
wire _11262_;
wire _11263_;
wire _11264_;
wire _11265_;
wire _11266_;
wire _11267_;
wire _11268_;
wire _11269_;
wire _11270_;
wire _11271_;
wire _11272_;
wire _11273_;
wire _11274_;
wire _11275_;
wire _11276_;
wire _11277_;
wire _11278_;
wire _11279_;
wire _11280_;
wire _11281_;
wire _11282_;
wire _11283_;
wire _11284_;
wire _11285_;
wire _11286_;
wire _11287_;
wire _11288_;
wire _11289_;
wire _11290_;
wire _11291_;
wire _11292_;
wire _11293_;
wire _11294_;
wire _11295_;
wire _11296_;
wire _11297_;
wire _11298_;
wire _11299_;
wire _11300_;
wire _11301_;
wire _11302_;
wire _11303_;
wire _11304_;
wire _11305_;
wire _11306_;
wire _11307_;
wire _11308_;
wire _11309_;
wire _11310_;
wire _11311_;
wire _11312_;
wire _11313_;
wire _11314_;
wire _11315_;
wire _11316_;
wire _11317_;
wire _11318_;
wire _11319_;
wire _11320_;
wire _11321_;
wire _11322_;
wire _11323_;
wire _11324_;
wire _11325_;
wire _11326_;
wire _11327_;
wire _11328_;
wire _11329_;
wire _11330_;
wire _11331_;
wire _11332_;
wire _11333_;
wire _11334_;
wire _11335_;
wire _11336_;
wire _11337_;
wire _11338_;
wire _11339_;
wire _11340_;
wire _11341_;
wire _11342_;
wire _11343_;
wire _11344_;
wire _11345_;
wire _11346_;
wire _11347_;
wire _11348_;
wire _11349_;
wire _11350_;
wire _11351_;
wire _11352_;
wire _11353_;
wire _11354_;
wire _11355_;
wire _11356_;
wire _11357_;
wire _11358_;
wire _11359_;
wire _11360_;
wire _11361_;
wire _11362_;
wire _11363_;
wire _11364_;
wire _11365_;
wire _11366_;
wire _11367_;
wire _11368_;
wire _11369_;
wire _11370_;
wire _11371_;
wire _11372_;
wire _11373_;
wire _11374_;
wire _11375_;
wire _11376_;
wire _11377_;
wire _11378_;
wire _11379_;
wire _11380_;
wire _11381_;
wire _11382_;
wire _11383_;
wire _11384_;
wire _11385_;
wire _11386_;
wire _11387_;
wire _11388_;
wire _11389_;
wire _11390_;
wire _11391_;
wire _11392_;
wire _11393_;
wire _11394_;
wire _11395_;
wire _11396_;
wire _11397_;
wire _11398_;
wire _11399_;
wire _11400_;
wire _11401_;
wire _11402_;
wire _11403_;
wire _11404_;
wire _11405_;
wire _11406_;
wire _11407_;
wire _11408_;
wire _11409_;
wire _11410_;
wire _11411_;
wire _11412_;
wire _11413_;
wire _11414_;
wire _11415_;
wire _11416_;
wire _11417_;
wire _11418_;
wire _11419_;
wire _11420_;
wire _11421_;
wire _11422_;
wire _11423_;
wire _11424_;
wire _11425_;
wire _11426_;
wire _11427_;
wire _11428_;
wire _11429_;
wire _11430_;
wire _11431_;
wire _11432_;
wire _11433_;
wire _11434_;
wire _11435_;
wire _11436_;
wire _11437_;
wire _11438_;
wire _11439_;
wire _11440_;
wire _11441_;
wire _11442_;
wire _11443_;
wire _11444_;
wire _11445_;
wire _11446_;
wire _11447_;
wire _11448_;
wire _11449_;
wire _11450_;
wire _11451_;
wire _11452_;
wire _11453_;
wire _11454_;
wire _11455_;
wire _11456_;
wire _11457_;
wire _11458_;
wire _11459_;
wire _11460_;
wire _11461_;
wire _11462_;
wire _11463_;
wire _11464_;
wire _11465_;
wire _11466_;
wire _11467_;
wire _11468_;
wire _11469_;
wire _11470_;
wire _11471_;
wire _11472_;
wire _11473_;
wire _11474_;
wire _11475_;
wire _11476_;
wire _11477_;
wire _11478_;
wire _11479_;
wire _11480_;
wire _11481_;
wire _11482_;
wire _11483_;
wire _11484_;
wire _11485_;
wire _11486_;
wire _11487_;
wire _11488_;
wire _11489_;
wire _11490_;
wire _11491_;
wire _11492_;
wire _11493_;
wire _11494_;
wire _11495_;
wire _11496_;
wire _11497_;
wire _11498_;
wire _11499_;
wire _11500_;
wire _11501_;
wire _11502_;
wire _11503_;
wire _11504_;
wire _11505_;
wire _11506_;
wire _11507_;
wire _11508_;
wire _11509_;
wire _11510_;
wire _11511_;
wire _11512_;
wire _11513_;
wire _11514_;
wire _11515_;
wire _11516_;
wire _11517_;
wire _11518_;
wire _11519_;
wire _11520_;
wire _11521_;
wire _11522_;
wire _11523_;
wire _11524_;
wire _11525_;
wire _11526_;
wire _11527_;
wire _11528_;
wire _11529_;
wire _11530_;
wire _11531_;
wire _11532_;
wire _11533_;
wire _11534_;
wire _11535_;
wire _11536_;
wire _11537_;
wire _11538_;
wire _11539_;
wire _11540_;
wire _11541_;
wire _11542_;
wire _11543_;
wire _11544_;
wire _11545_;
wire _11546_;
wire _11547_;
wire _11548_;
wire _11549_;
wire _11550_;
wire _11551_;
wire _11552_;
wire _11553_;
wire _11554_;
wire _11555_;
wire _11556_;
wire _11557_;
wire _11558_;
wire _11559_;
wire _11560_;
wire _11561_;
wire _11562_;
wire _11563_;
wire _11564_;
wire _11565_;
wire _11566_;
wire _11567_;
wire _11568_;
wire _11569_;
wire _11570_;
wire _11571_;
wire _11572_;
wire _11573_;
wire _11574_;
wire _11575_;
wire _11576_;
wire _11577_;
wire _11578_;
wire _11579_;
wire _11580_;
wire _11581_;
wire _11582_;
wire _11583_;
wire _11584_;
wire _11585_;
wire _11586_;
wire _11587_;
wire _11588_;
wire _11589_;
wire _11590_;
wire _11591_;
wire _11592_;
wire _11593_;
wire _11594_;
wire _11595_;
wire _11596_;
wire _11597_;
wire _11598_;
wire _11599_;
wire _11600_;
wire _11601_;
wire _11602_;
wire _11603_;
wire _11604_;
wire _11605_;
wire _11606_;
wire _11607_;
wire _11608_;
wire _11609_;
wire _11610_;
wire _11611_;
wire _11612_;
wire _11613_;
wire _11614_;
wire _11615_;
wire _11616_;
wire _11617_;
wire _11618_;
wire _11619_;
wire _11620_;
wire _11621_;
wire _11622_;
wire _11623_;
wire _11624_;
wire _11625_;
wire _11626_;
wire _11627_;
wire _11628_;
wire _11629_;
wire _11630_;
wire _11631_;
wire _11632_;
wire _11633_;
wire _11634_;
wire _11635_;
wire _11636_;
wire _11637_;
wire _11638_;
wire _11639_;
wire _11640_;
wire _11641_;
wire _11642_;
wire _11643_;
wire _11644_;
wire _11645_;
wire _11646_;
wire _11647_;
wire _11648_;
wire _11649_;
wire _11650_;
wire _11651_;
wire _11652_;
wire _11653_;
wire _11654_;
wire _11655_;
wire _11656_;
wire _11657_;
wire _11658_;
wire _11659_;
wire _11660_;
wire _11661_;
wire _11662_;
wire _11663_;
wire _11664_;
wire _11665_;
wire _11666_;
wire _11667_;
wire _11668_;
wire _11669_;
wire _11670_;
wire _11671_;
wire _11672_;
wire _11673_;
wire _11674_;
wire _11675_;
wire _11676_;
wire _11677_;
wire _11678_;
wire _11679_;
wire _11680_;
wire _11681_;
wire _11682_;
wire _11683_;
wire _11684_;
wire _11685_;
wire _11686_;
wire _11687_;
wire _11688_;
wire _11689_;
wire _11690_;
wire _11691_;
wire _11692_;
wire _11693_;
wire _11694_;
wire _11695_;
wire _11696_;
wire _11697_;
wire _11698_;
wire _11699_;
wire _11700_;
wire _11701_;
wire _11702_;
wire _11703_;
wire _11704_;
wire _11705_;
wire _11706_;
wire _11707_;
wire _11708_;
wire _11709_;
wire _11710_;
wire _11711_;
wire _11712_;
wire _11713_;
wire _11714_;
wire _11715_;
wire _11716_;
wire _11717_;
wire _11718_;
wire _11719_;
wire _11720_;
wire _11721_;
wire _11722_;
wire _11723_;
wire _11724_;
wire _11725_;
wire _11726_;
wire _11727_;
wire _11728_;
wire _11729_;
wire _11730_;
wire _11731_;
wire _11732_;
wire _11733_;
wire _11734_;
wire _11735_;
wire _11736_;
wire _11737_;
wire _11738_;
wire _11739_;
wire _11740_;
wire _11741_;
wire _11742_;
wire _11743_;
wire _11744_;
wire _11745_;
wire _11746_;
wire _11747_;
wire _11748_;
wire _11749_;
wire _11750_;
wire _11751_;
wire _11752_;
wire _11753_;
wire _11754_;
wire _11755_;
wire _11756_;
wire _11757_;
wire _11758_;
wire _11759_;
wire _11760_;
wire _11761_;
wire _11762_;
wire _11763_;
wire _11764_;
wire _11765_;
wire _11766_;
wire _11767_;
wire _11768_;
wire _11769_;
wire _11770_;
wire _11771_;
wire _11772_;
wire _11773_;
wire _11774_;
wire _11775_;
wire _11776_;
wire _11777_;
wire _11778_;
wire _11779_;
wire _11780_;
wire _11781_;
wire _11782_;
wire _11783_;
wire _11784_;
wire _11785_;
wire _11786_;
wire _11787_;
wire _11788_;
wire _11789_;
wire _11790_;
wire _11791_;
wire _11792_;
wire _11793_;
wire _11794_;
wire _11795_;
wire _11796_;
wire _11797_;
wire _11798_;
wire _11799_;
wire _11800_;
wire _11801_;
wire _11802_;
wire _11803_;
wire _11804_;
wire _11805_;
wire _11806_;
wire _11807_;
wire _11808_;
wire _11809_;
wire _11810_;
wire _11811_;
wire _11812_;
wire _11813_;
wire _11814_;
wire _11815_;
wire _11816_;
wire _11817_;
wire _11818_;
wire _11819_;
wire _11820_;
wire _11821_;
wire _11822_;
wire _11823_;
wire _11824_;
wire _11825_;
wire _11826_;
wire _11827_;
wire _11828_;
wire _11829_;
wire _11830_;
wire _11831_;
wire _11832_;
wire _11833_;
wire _11834_;
wire _11835_;
wire _11836_;
wire _11837_;
wire _11838_;
wire _11839_;
wire _11840_;
wire _11841_;
wire _11842_;
wire _11843_;
wire _11844_;
wire _11845_;
wire _11846_;
wire _11847_;
wire _11848_;
wire _11849_;
wire _11850_;
wire _11851_;
wire _11852_;
wire _11853_;
wire _11854_;
wire _11855_;
wire _11856_;
wire _11857_;
wire _11858_;
wire _11859_;
wire _11860_;
wire _11861_;
wire _11862_;
wire _11863_;
wire _11864_;
wire _11865_;
wire _11866_;
wire _11867_;
wire _11868_;
wire _11869_;
wire _11870_;
wire _11871_;
wire _11872_;
wire _11873_;
wire _11874_;
wire _11875_;
wire _11876_;
wire _11877_;
wire _11878_;
wire _11879_;
wire _11880_;
wire _11881_;
wire _11882_;
wire _11883_;
wire _11884_;
wire _11885_;
wire _11886_;
wire _11887_;
wire _11888_;
wire _11889_;
wire _11890_;
wire _11891_;
wire _11892_;
wire _11893_;
wire _11894_;
wire _11895_;
wire _11896_;
wire _11897_;
wire _11898_;
wire _11899_;
wire _11900_;
wire _11901_;
wire _11902_;
wire _11903_;
wire _11904_;
wire _11905_;
wire _11906_;
wire _11907_;
wire _11908_;
wire _11909_;
wire _11910_;
wire _11911_;
wire _11912_;
wire _11913_;
wire _11914_;
wire _11915_;
wire _11916_;
wire _11917_;
wire _11918_;
wire _11919_;
wire _11920_;
wire _11921_;
wire _11922_;
wire _11923_;
wire _11924_;
wire _11925_;
wire _11926_;
wire _11927_;
wire _11928_;
wire _11929_;
wire _11930_;
wire _11931_;
wire _11932_;
wire _11933_;
wire _11934_;
wire _11935_;
wire _11936_;
wire _11937_;
wire _11938_;
wire _11939_;
wire _11940_;
wire _11941_;
wire _11942_;
wire _11943_;
wire _11944_;
wire _11945_;
wire _11946_;
wire _11947_;
wire _11948_;
wire _11949_;
wire _11950_;
wire _11951_;
wire _11952_;
wire _11953_;
wire _11954_;
wire _11955_;
wire _11956_;
wire _11957_;
wire _11958_;
wire _11959_;
wire _11960_;
wire _11961_;
wire _11962_;
wire _11963_;
wire _11964_;
wire _11965_;
wire _11966_;
wire _11967_;
wire _11968_;
wire _11969_;
wire _11970_;
wire _11971_;
wire _11972_;
wire _11973_;
wire _11974_;
wire _11975_;
wire _11976_;
wire _11977_;
wire _11978_;
wire _11979_;
wire _11980_;
wire _11981_;
wire _11982_;
wire _11983_;
wire _11984_;
wire _11985_;
wire _11986_;
wire _11987_;
wire _11988_;
wire _11989_;
wire _11990_;
wire _11991_;
wire _11992_;
wire _11993_;
wire _11994_;
wire _11995_;
wire _11996_;
wire _11997_;
wire _11998_;
wire _11999_;
wire _12000_;
wire _12001_;
wire _12002_;
wire _12003_;
wire _12004_;
wire _12005_;
wire _12006_;
wire _12007_;
wire _12008_;
wire _12009_;
wire _12010_;
wire _12011_;
wire _12012_;
wire _12013_;
wire _12014_;
wire _12015_;
wire _12016_;
wire _12017_;
wire _12018_;
wire _12019_;
wire _12020_;
wire _12021_;
wire _12022_;
wire _12023_;
wire _12024_;
wire _12025_;
wire _12026_;
wire _12027_;
wire _12028_;
wire _12029_;
wire _12030_;
wire _12031_;
wire _12032_;
wire _12033_;
wire _12034_;
wire _12035_;
wire _12036_;
wire _12037_;
wire _12038_;
wire _12039_;
wire _12040_;
wire _12041_;
wire _12042_;
wire _12043_;
wire _12044_;
wire _12045_;
wire _12046_;
wire _12047_;
wire _12048_;
wire _12049_;
wire _12050_;
wire _12051_;
wire _12052_;
wire _12053_;
wire _12054_;
wire _12055_;
wire _12056_;
wire _12057_;
wire _12058_;
wire _12059_;
wire _12060_;
wire _12061_;
wire _12062_;
wire _12063_;
wire _12064_;
wire _12065_;
wire _12066_;
wire _12067_;
wire _12068_;
wire _12069_;
wire _12070_;
wire _12071_;
wire _12072_;
wire _12073_;
wire _12074_;
wire _12075_;
wire _12076_;
wire _12077_;
wire _12078_;
wire _12079_;
wire _12080_;
wire _12081_;
wire _12082_;
wire _12083_;
wire _12084_;
wire _12085_;
wire _12086_;
wire _12087_;
wire _12088_;
wire _12089_;
wire _12090_;
wire _12091_;
wire _12092_;
wire _12093_;
wire _12094_;
wire _12095_;
wire _12096_;
wire _12097_;
wire _12098_;
wire _12099_;
wire _12100_;
wire _12101_;
wire _12102_;
wire _12103_;
wire _12104_;
wire _12105_;
wire _12106_;
wire _12107_;
wire _12108_;
wire _12109_;
wire _12110_;
wire _12111_;
wire _12112_;
wire _12113_;
wire _12114_;
wire _12115_;
wire _12116_;
wire _12117_;
wire _12118_;
wire _12119_;
wire _12120_;
wire _12121_;
wire _12122_;
wire _12123_;
wire _12124_;
wire _12125_;
wire _12126_;
wire _12127_;
wire _12128_;
wire _12129_;
wire _12130_;
wire _12131_;
wire _12132_;
wire _12133_;
wire _12134_;
wire _12135_;
wire _12136_;
wire _12137_;
wire _12138_;
wire _12139_;
wire _12140_;
wire _12141_;
wire _12142_;
wire _12143_;
wire _12144_;
wire _12145_;
wire _12146_;
wire _12147_;
wire _12148_;
wire _12149_;
wire _12150_;
wire _12151_;
wire _12152_;
wire _12153_;
wire _12154_;
wire _12155_;
wire _12156_;
wire _12157_;
wire _12158_;
wire _12159_;
wire _12160_;
wire _12161_;
wire _12162_;
wire _12163_;
wire _12164_;
wire _12165_;
wire _12166_;
wire _12167_;
wire _12168_;
wire _12169_;
wire _12170_;
wire _12171_;
wire _12172_;
wire _12173_;
wire _12174_;
wire _12175_;
wire _12176_;
wire _12177_;
wire _12178_;
wire _12179_;
wire _12180_;
wire _12181_;
wire _12182_;
wire _12183_;
wire _12184_;
wire _12185_;
wire _12186_;
wire _12187_;
wire _12188_;
wire _12189_;
wire _12190_;
wire _12191_;
wire _12192_;
wire _12193_;
wire _12194_;
wire _12195_;
wire _12196_;
wire _12197_;
wire _12198_;
wire _12199_;
wire _12200_;
wire _12201_;
wire _12202_;
wire _12203_;
wire _12204_;
wire _12205_;
wire _12206_;
wire _12207_;
wire _12208_;
wire _12209_;
wire _12210_;
wire _12211_;
wire _12212_;
wire _12213_;
wire _12214_;
wire _12215_;
wire _12216_;
wire _12217_;
wire _12218_;
wire _12219_;
wire _12220_;
wire _12221_;
wire _12222_;
wire _12223_;
wire _12224_;
wire _12225_;
wire _12226_;
wire _12227_;
wire _12228_;
wire _12229_;
wire _12230_;
wire _12231_;
wire _12232_;
wire _12233_;
wire _12234_;
wire _12235_;
wire _12236_;
wire _12237_;
wire _12238_;
wire _12239_;
wire _12240_;
wire _12241_;
wire _12242_;
wire _12243_;
wire _12244_;
wire _12245_;
wire _12246_;
wire _12247_;
wire _12248_;
wire _12249_;
wire _12250_;
wire _12251_;
wire _12252_;
wire _12253_;
wire _12254_;
wire _12255_;
wire _12256_;
wire _12257_;
wire _12258_;
wire _12259_;
wire _12260_;
wire _12261_;
wire _12262_;
wire _12263_;
wire _12264_;
wire _12265_;
wire _12266_;
wire _12267_;
wire _12268_;
wire _12269_;
wire _12270_;
wire _12271_;
wire _12272_;
wire _12273_;
wire _12274_;
wire _12275_;
wire _12276_;
wire _12277_;
wire _12278_;
wire _12279_;
wire _12280_;
wire _12281_;
wire _12282_;
wire _12283_;
wire _12284_;
wire _12285_;
wire _12286_;
wire _12287_;
wire _12288_;
wire _12289_;
wire _12290_;
wire _12291_;
wire _12292_;
wire _12293_;
wire _12294_;
wire _12295_;
wire _12296_;
wire _12297_;
wire _12298_;
wire _12299_;
wire _12300_;
wire _12301_;
wire _12302_;
wire _12303_;
wire _12304_;
wire _12305_;
wire _12306_;
wire _12307_;
wire _12308_;
wire _12309_;
wire _12310_;
wire _12311_;
wire _12312_;
wire _12313_;
wire _12314_;
wire _12315_;
wire _12316_;
wire _12317_;
wire _12318_;
wire _12319_;
wire _12320_;
wire _12321_;
wire _12322_;
wire _12323_;
wire _12324_;
wire _12325_;
wire _12326_;
wire _12327_;
wire _12328_;
wire _12329_;
wire _12330_;
wire _12331_;
wire _12332_;
wire _12333_;
wire _12334_;
wire _12335_;
wire _12336_;
wire _12337_;
wire _12338_;
wire _12339_;
wire _12340_;
wire _12341_;
wire _12342_;
wire _12343_;
wire _12344_;
wire _12345_;
wire _12346_;
wire _12347_;
wire _12348_;
wire _12349_;
wire _12350_;
wire _12351_;
wire _12352_;
wire _12353_;
wire _12354_;
wire _12355_;
wire _12356_;
wire _12357_;
wire _12358_;
wire _12359_;
wire _12360_;
wire _12361_;
wire _12362_;
wire _12363_;
wire _12364_;
wire _12365_;
wire _12366_;
wire _12367_;
wire _12368_;
wire _12369_;
wire _12370_;
wire _12371_;
wire _12372_;
wire _12373_;
wire _12374_;
wire _12375_;
wire _12376_;
wire _12377_;
wire _12378_;
wire _12379_;
wire _12380_;
wire _12381_;
wire _12382_;
wire _12383_;
wire _12384_;
wire _12385_;
wire _12386_;
wire _12387_;
wire _12388_;
wire _12389_;
wire _12390_;
wire _12391_;
wire _12392_;
wire _12393_;
wire _12394_;
wire _12395_;
wire _12396_;
wire _12397_;
wire _12398_;
wire _12399_;
wire _12400_;
wire _12401_;
wire _12402_;
wire _12403_;
wire _12404_;
wire _12405_;
wire _12406_;
wire _12407_;
wire _12408_;
wire _12409_;
wire _12410_;
wire _12411_;
wire _12412_;
wire _12413_;
wire _12414_;
wire _12415_;
wire _12416_;
wire _12417_;
wire _12418_;
wire _12419_;
wire _12420_;
wire _12421_;
wire _12422_;
wire _12423_;
wire _12424_;
wire _12425_;
wire _12426_;
wire _12427_;
wire _12428_;
wire _12429_;
wire _12430_;
wire _12431_;
wire _12432_;
wire _12433_;
wire _12434_;
wire _12435_;
wire _12436_;
wire _12437_;
wire _12438_;
wire _12439_;
wire _12440_;
wire _12441_;
wire _12442_;
wire _12443_;
wire _12444_;
wire _12445_;
wire _12446_;
wire _12447_;
wire _12448_;
wire _12449_;
wire _12450_;
wire _12451_;
wire _12452_;
wire _12453_;
wire _12454_;
wire _12455_;
wire _12456_;
wire _12457_;
wire _12458_;
wire _12459_;
wire _12460_;
wire _12461_;
wire _12462_;
wire _12463_;
wire _12464_;
wire _12465_;
wire _12466_;
wire _12467_;
wire _12468_;
wire _12469_;
wire _12470_;
wire _12471_;
wire _12472_;
wire _12473_;
wire _12474_;
wire _12475_;
wire _12476_;
wire _12477_;
wire _12478_;
wire _12479_;
wire _12480_;
wire _12481_;
wire _12482_;
wire _12483_;
wire _12484_;
wire _12485_;
wire _12486_;
wire _12487_;
wire _12488_;
wire _12489_;
wire _12490_;
wire _12491_;
wire _12492_;
wire _12493_;
wire _12494_;
wire _12495_;
wire _12496_;
wire _12497_;
wire _12498_;
wire _12499_;
wire _12500_;
wire _12501_;
wire _12502_;
wire _12503_;
wire _12504_;
wire _12505_;
wire _12506_;
wire _12507_;
wire _12508_;
wire _12509_;
wire _12510_;
wire _12511_;
wire _12512_;
wire _12513_;
wire _12514_;
wire _12515_;
wire _12516_;
wire _12517_;
wire _12518_;
wire _12519_;
wire _12520_;
wire _12521_;
wire _12522_;
wire _12523_;
wire _12524_;
wire _12525_;
wire _12526_;
wire _12527_;
wire _12528_;
wire _12529_;
wire _12530_;
wire _12531_;
wire _12532_;
wire _12533_;
wire _12534_;
wire _12535_;
wire _12536_;
wire _12537_;
wire _12538_;
wire _12539_;
wire _12540_;
wire _12541_;
wire _12542_;
wire _12543_;
wire _12544_;
wire _12545_;
wire _12546_;
wire _12547_;
wire _12548_;
wire _12549_;
wire _12550_;
wire _12551_;
wire _12552_;
wire _12553_;
wire _12554_;
wire _12555_;
wire _12556_;
wire _12557_;
wire _12558_;
wire _12559_;
wire _12560_;
wire _12561_;
wire _12562_;
wire _12563_;
wire _12564_;
wire _12565_;
wire _12566_;
wire _12567_;
wire _12568_;
wire _12569_;
wire _12570_;
wire _12571_;
wire _12572_;
wire _12573_;
wire _12574_;
wire _12575_;
wire _12576_;
wire _12577_;
wire _12578_;
wire _12579_;
wire _12580_;
wire _12581_;
wire _12582_;
wire _12583_;
wire _12584_;
wire _12585_;
wire _12586_;
wire _12587_;
wire _12588_;
wire _12589_;
wire _12590_;
wire _12591_;
wire _12592_;
wire _12593_;
wire _12594_;
wire _12595_;
wire _12596_;
wire _12597_;
wire _12598_;
wire _12599_;
wire _12600_;
wire _12601_;
wire _12602_;
wire _12603_;
wire _12604_;
wire _12605_;
wire _12606_;
wire _12607_;
wire _12608_;
wire _12609_;
wire _12610_;
wire _12611_;
wire _12612_;
wire _12613_;
wire _12614_;
wire _12615_;
wire _12616_;
wire _12617_;
wire _12618_;
wire _12619_;
wire _12620_;
wire _12621_;
wire _12622_;
wire _12623_;
wire _12624_;
wire _12625_;
wire _12626_;
wire _12627_;
wire _12628_;
wire _12629_;
wire _12630_;
wire _12631_;
wire _12632_;
wire _12633_;
wire _12634_;
wire _12635_;
wire _12636_;
wire _12637_;
wire _12638_;
wire _12639_;
wire _12640_;
wire _12641_;
wire _12642_;
wire _12643_;
wire _12644_;
wire _12645_;
wire _12646_;
wire _12647_;
wire _12648_;
wire _12649_;
wire _12650_;
wire _12651_;
wire _12652_;
wire _12653_;
wire _12654_;
wire _12655_;
wire _12656_;
wire _12657_;
wire _12658_;
wire _12659_;
wire _12660_;
wire _12661_;
wire _12662_;
wire _12663_;
wire _12664_;
wire _12665_;
wire _12666_;
wire _12667_;
wire _12668_;
wire _12669_;
wire _12670_;
wire _12671_;
wire _12672_;
wire _12673_;
wire _12674_;
wire _12675_;
wire _12676_;
wire _12677_;
wire _12678_;
wire _12679_;
wire _12680_;
wire _12681_;
wire _12682_;
wire _12683_;
wire _12684_;
wire _12685_;
wire _12686_;
wire _12687_;
wire _12688_;
wire _12689_;
wire _12690_;
wire _12691_;
wire _12692_;
wire _12693_;
wire _12694_;
wire _12695_;
wire _12696_;
wire _12697_;
wire _12698_;
wire _12699_;
wire _12700_;
wire _12701_;
wire _12702_;
wire _12703_;
wire _12704_;
wire _12705_;
wire _12706_;
wire _12707_;
wire _12708_;
wire _12709_;
wire _12710_;
wire _12711_;
wire _12712_;
wire _12713_;
wire _12714_;
wire _12715_;
wire _12716_;
wire _12717_;
wire _12718_;
wire _12719_;
wire _12720_;
wire _12721_;
wire _12722_;
wire _12723_;
wire _12724_;
wire _12725_;
wire _12726_;
wire _12727_;
wire _12728_;
wire _12729_;
wire _12730_;
wire _12731_;
wire _12732_;
wire _12733_;
wire _12734_;
wire _12735_;
wire _12736_;
wire _12737_;
wire _12738_;
wire _12739_;
wire _12740_;
wire _12741_;
wire _12742_;
wire _12743_;
wire _12744_;
wire _12745_;
wire _12746_;
wire _12747_;
wire _12748_;
wire _12749_;
wire _12750_;
wire _12751_;
wire _12752_;
wire _12753_;
wire _12754_;
wire _12755_;
wire _12756_;
wire _12757_;
wire _12758_;
wire _12759_;
wire _12760_;
wire _12761_;
wire _12762_;
wire _12763_;
wire _12764_;
wire _12765_;
wire _12766_;
wire _12767_;
wire _12768_;
wire _12769_;
wire _12770_;
wire _12771_;
wire _12772_;
wire _12773_;
wire _12774_;
wire _12775_;
wire _12776_;
wire _12777_;
wire _12778_;
wire _12779_;
wire _12780_;
wire _12781_;
wire _12782_;
wire _12783_;
wire _12784_;
wire _12785_;
wire _12786_;
wire _12787_;
wire _12788_;
wire _12789_;
wire _12790_;
wire _12791_;
wire _12792_;
wire _12793_;
wire _12794_;
wire _12795_;
wire _12796_;
wire _12797_;
wire _12798_;
wire _12799_;
wire _12800_;
wire _12801_;
wire _12802_;
wire _12803_;
wire _12804_;
wire _12805_;
wire _12806_;
wire _12807_;
wire _12808_;
wire _12809_;
wire _12810_;
wire _12811_;
wire _12812_;
wire _12813_;
wire _12814_;
wire _12815_;
wire _12816_;
wire _12817_;
wire _12818_;
wire _12819_;
wire _12820_;
wire _12821_;
wire _12822_;
wire _12823_;
wire _12824_;
wire _12825_;
wire _12826_;
wire _12827_;
wire _12828_;
wire _12829_;
wire _12830_;
wire _12831_;
wire _12832_;
wire _12833_;
wire _12834_;
wire _12835_;
wire _12836_;
wire _12837_;
wire _12838_;
wire _12839_;
wire _12840_;
wire _12841_;
wire _12842_;
wire _12843_;
wire _12844_;
wire _12845_;
wire _12846_;
wire _12847_;
wire _12848_;
wire _12849_;
wire _12850_;
wire _12851_;
wire _12852_;
wire _12853_;
wire _12854_;
wire _12855_;
wire _12856_;
wire _12857_;
wire _12858_;
wire _12859_;
wire _12860_;
wire _12861_;
wire _12862_;
wire _12863_;
wire _12864_;
wire _12865_;
wire _12866_;
wire _12867_;
wire _12868_;
wire _12869_;
wire _12870_;
wire _12871_;
wire _12872_;
wire _12873_;
wire _12874_;
wire _12875_;
wire _12876_;
wire _12877_;
wire _12878_;
wire _12879_;
wire _12880_;
wire _12881_;
wire _12882_;
wire _12883_;
wire _12884_;
wire _12885_;
wire _12886_;
wire _12887_;
wire _12888_;
wire _12889_;
wire _12890_;
wire _12891_;
wire _12892_;
wire _12893_;
wire _12894_;
wire _12895_;
wire _12896_;
wire _12897_;
wire _12898_;
wire _12899_;
wire _12900_;
wire _12901_;
wire _12902_;
wire _12903_;
wire _12904_;
wire _12905_;
wire _12906_;
wire _12907_;
wire _12908_;
wire _12909_;
wire _12910_;
wire _12911_;
wire _12912_;
wire _12913_;
wire _12914_;
wire _12915_;
wire _12916_;
wire _12917_;
wire _12918_;
wire _12919_;
wire _12920_;
wire _12921_;
wire _12922_;
wire _12923_;
wire _12924_;
wire _12925_;
wire _12926_;
wire _12927_;
wire _12928_;
wire _12929_;
wire _12930_;
wire _12931_;
wire _12932_;
wire _12933_;
wire _12934_;
wire _12935_;
wire _12936_;
wire _12937_;
wire _12938_;
wire _12939_;
wire _12940_;
wire _12941_;
wire _12942_;
wire _12943_;
wire _12944_;
wire _12945_;
wire _12946_;
wire _12947_;
wire _12948_;
wire _12949_;
wire _12950_;
wire _12951_;
wire _12952_;
wire _12953_;
wire _12954_;
wire _12955_;
wire _12956_;
wire _12957_;
wire _12958_;
wire _12959_;
wire _12960_;
wire _12961_;
wire _12962_;
wire _12963_;
wire _12964_;
wire _12965_;
wire _12966_;
wire _12967_;
wire _12968_;
wire _12969_;
wire _12970_;
wire _12971_;
wire _12972_;
wire _12973_;
wire _12974_;
wire _12975_;
wire _12976_;
wire _12977_;
wire _12978_;
wire _12979_;
wire _12980_;
wire _12981_;
wire _12982_;
wire _12983_;
wire _12984_;
wire _12985_;
wire _12986_;
wire _12987_;
wire _12988_;
wire _12989_;
wire _12990_;
wire _12991_;
wire _12992_;
wire _12993_;
wire _12994_;
wire _12995_;
wire _12996_;
wire _12997_;
wire _12998_;
wire _12999_;
wire _13000_;
wire _13001_;
wire _13002_;
wire _13003_;
wire _13004_;
wire _13005_;
wire _13006_;
wire _13007_;
wire _13008_;
wire _13009_;
wire _13010_;
wire _13011_;
wire _13012_;
wire _13013_;
wire _13014_;
wire _13015_;
wire _13016_;
wire _13017_;
wire _13018_;
wire _13019_;
wire _13020_;
wire _13021_;
wire _13022_;
wire _13023_;
wire _13024_;
wire _13025_;
wire _13026_;
wire _13027_;
wire _13028_;
wire _13029_;
wire _13030_;
wire _13031_;
wire _13032_;
wire _13033_;
wire _13034_;
wire _13035_;
wire _13036_;
wire _13037_;
wire _13038_;
wire _13039_;
wire _13040_;
wire _13041_;
wire _13042_;
wire _13043_;
wire _13044_;
wire _13045_;
wire _13046_;
wire _13047_;
wire _13048_;
wire _13049_;
wire _13050_;
wire _13051_;
wire _13052_;
wire _13053_;
wire _13054_;
wire _13055_;
wire _13056_;
wire _13057_;
wire _13058_;
wire _13059_;
wire _13060_;
wire _13061_;
wire _13062_;
wire _13063_;
wire _13064_;
wire _13065_;
wire _13066_;
wire _13067_;
wire _13068_;
wire _13069_;
wire _13070_;
wire _13071_;
wire _13072_;
wire _13073_;
wire _13074_;
wire _13075_;
wire _13076_;
wire _13077_;
wire _13078_;
wire _13079_;
wire _13080_;
wire _13081_;
wire _13082_;
wire _13083_;
wire _13084_;
wire _13085_;
wire _13086_;
wire _13087_;
wire _13088_;
wire _13089_;
wire _13090_;
wire _13091_;
wire _13092_;
wire _13093_;
wire _13094_;
wire _13095_;
wire _13096_;
wire _13097_;
wire _13098_;
wire _13099_;
wire _13100_;
wire _13101_;
wire _13102_;
wire _13103_;
wire _13104_;
wire _13105_;
wire _13106_;
wire _13107_;
wire _13108_;
wire _13109_;
wire _13110_;
wire _13111_;
wire _13112_;
wire _13113_;
wire _13114_;
wire _13115_;
wire _13116_;
wire _13117_;
wire _13118_;
wire _13119_;
wire _13120_;
wire _13121_;
wire _13122_;
wire _13123_;
wire _13124_;
wire _13125_;
wire _13126_;
wire _13127_;
wire _13128_;
wire _13129_;
wire _13130_;
wire _13131_;
wire _13132_;
wire _13133_;
wire _13134_;
wire _13135_;
wire _13136_;
wire _13137_;
wire _13138_;
wire _13139_;
wire _13140_;
wire _13141_;
wire _13142_;
wire _13143_;
wire _13144_;
wire _13145_;
wire _13146_;
wire _13147_;
wire _13148_;
wire _13149_;
wire _13150_;
wire _13151_;
wire _13152_;
wire _13153_;
wire _13154_;
wire _13155_;
wire _13156_;
wire _13157_;
wire _13158_;
wire _13159_;
wire _13160_;
wire _13161_;
wire _13162_;
wire _13163_;
wire _13164_;
wire _13165_;
wire _13166_;
wire _13167_;
wire _13168_;
wire _13169_;
wire _13170_;
wire _13171_;
wire _13172_;
wire _13173_;
wire _13174_;
wire _13175_;
wire _13176_;
wire _13177_;
wire _13178_;
wire _13179_;
wire _13180_;
wire _13181_;
wire _13182_;
wire _13183_;
wire _13184_;
wire _13185_;
wire _13186_;
wire _13187_;
wire _13188_;
wire _13189_;
wire _13190_;
wire _13191_;
wire _13192_;
wire _13193_;
wire _13194_;
wire _13195_;
wire _13196_;
wire _13197_;
wire _13198_;
wire _13199_;
wire _13200_;
wire _13201_;
wire _13202_;
wire _13203_;
wire _13204_;
wire _13205_;
wire _13206_;
wire _13207_;
wire _13208_;
wire _13209_;
wire _13210_;
wire _13211_;
wire _13212_;
wire _13213_;
wire _13214_;
wire _13215_;
wire _13216_;
wire _13217_;
wire _13218_;
wire _13219_;
wire _13220_;
wire _13221_;
wire _13222_;
wire _13223_;
wire _13224_;
wire _13225_;
wire _13226_;
wire _13227_;
wire _13228_;
wire _13229_;
wire _13230_;
wire _13231_;
wire _13232_;
wire _13233_;
wire _13234_;
wire _13235_;
wire _13236_;
wire _13237_;
wire _13238_;
wire _13239_;
wire _13240_;
wire _13241_;
wire _13242_;
wire _13243_;
wire _13244_;
wire _13245_;
wire _13246_;
wire _13247_;
wire _13248_;
wire _13249_;
wire _13250_;
wire _13251_;
wire _13252_;
wire _13253_;
wire _13254_;
wire _13255_;
wire _13256_;
wire _13257_;
wire _13258_;
wire _13259_;
wire _13260_;
wire _13261_;
wire _13262_;
wire _13263_;
wire _13264_;
wire _13265_;
wire _13266_;
wire _13267_;
wire _13268_;
wire _13269_;
wire _13270_;
wire _13271_;
wire _13272_;
wire _13273_;
wire _13274_;
wire _13275_;
wire _13276_;
wire _13277_;
wire _13278_;
wire _13279_;
wire _13280_;
wire _13281_;
wire _13282_;
wire _13283_;
wire _13284_;
wire _13285_;
wire _13286_;
wire _13287_;
wire _13288_;
wire _13289_;
wire _13290_;
wire _13291_;
wire _13292_;
wire _13293_;
wire _13294_;
wire _13295_;
wire _13296_;
wire _13297_;
wire _13298_;
wire _13299_;
wire _13300_;
wire _13301_;
wire _13302_;
wire _13303_;
wire _13304_;
wire _13305_;
wire _13306_;
wire _13307_;
wire _13308_;
wire _13309_;
wire _13310_;
wire _13311_;
wire _13312_;
wire _13313_;
wire _13314_;
wire _13315_;
wire _13316_;
wire _13317_;
wire _13318_;
wire _13319_;
wire _13320_;
wire _13321_;
wire _13322_;
wire _13323_;
wire _13324_;
wire _13325_;
wire _13326_;
wire _13327_;
wire _13328_;
wire _13329_;
wire _13330_;
wire _13331_;
wire _13332_;
wire _13333_;
wire _13334_;
wire _13335_;
wire _13336_;
wire _13337_;
wire _13338_;
wire _13339_;
wire _13340_;
wire _13341_;
wire _13342_;
wire _13343_;
wire _13344_;
wire _13345_;
wire _13346_;
wire _13347_;
wire _13348_;
wire _13349_;
wire _13350_;
wire _13351_;
wire _13352_;
wire _13353_;
wire _13354_;
wire _13355_;
wire _13356_;
wire _13357_;
wire _13358_;
wire _13359_;
wire _13360_;
wire _13361_;
wire _13362_;
wire _13363_;
wire _13364_;
wire _13365_;
wire _13366_;
wire _13367_;
wire _13368_;
wire _13369_;
wire _13370_;
wire _13371_;
wire _13372_;
wire _13373_;
wire _13374_;
wire _13375_;
wire _13376_;
wire _13377_;
wire _13378_;
wire _13379_;
wire _13380_;
wire _13381_;
wire _13382_;
wire _13383_;
wire _13384_;
wire _13385_;
wire _13386_;
wire _13387_;
wire _13388_;
wire _13389_;
wire _13390_;
wire _13391_;
wire _13392_;
wire _13393_;
wire _13394_;
wire _13395_;
wire _13396_;
wire _13397_;
wire _13398_;
wire _13399_;
wire _13400_;
wire _13401_;
wire _13402_;
wire _13403_;
wire _13404_;
wire _13405_;
wire _13406_;
wire _13407_;
wire _13408_;
wire _13409_;
wire _13410_;
wire _13411_;
wire _13412_;
wire _13413_;
wire _13414_;
wire _13415_;
wire _13416_;
wire _13417_;
wire _13418_;
wire _13419_;
wire _13420_;
wire _13421_;
wire _13422_;
wire _13423_;
wire _13424_;
wire _13425_;
wire _13426_;
wire _13427_;
wire _13428_;
wire _13429_;
wire _13430_;
wire _13431_;
wire _13432_;
wire _13433_;
wire _13434_;
wire _13435_;
wire _13436_;
wire _13437_;
wire _13438_;
wire _13439_;
wire _13440_;
wire _13441_;
wire _13442_;
wire _13443_;
wire _13444_;
wire _13445_;
wire _13446_;
wire _13447_;
wire _13448_;
wire _13449_;
wire _13450_;
wire _13451_;
wire _13452_;
wire _13453_;
wire _13454_;
wire _13455_;
wire _13456_;
wire _13457_;
wire _13458_;
wire _13459_;
wire _13460_;
wire _13461_;
wire _13462_;
wire _13463_;
wire _13464_;
wire _13465_;
wire _13466_;
wire _13467_;
wire _13468_;
wire _13469_;
wire _13470_;
wire _13471_;
wire _13472_;
wire _13473_;
wire _13474_;
wire _13475_;
wire _13476_;
wire _13477_;
wire _13478_;
wire _13479_;
wire _13480_;
wire _13481_;
wire _13482_;
wire _13483_;
wire _13484_;
wire _13485_;
wire _13486_;
wire _13487_;
wire _13488_;
wire _13489_;
wire _13490_;
wire _13491_;
wire _13492_;
wire _13493_;
wire _13494_;
wire _13495_;
wire _13496_;
wire _13497_;
wire _13498_;
wire _13499_;
wire _13500_;
wire _13501_;
wire _13502_;
wire _13503_;
wire _13504_;
wire _13505_;
wire _13506_;
wire _13507_;
wire _13508_;
wire _13509_;
wire _13510_;
wire _13511_;
wire _13512_;
wire _13513_;
wire _13514_;
wire _13515_;
wire _13516_;
wire _13517_;
wire _13518_;
wire _13519_;
wire _13520_;
wire _13521_;
wire _13522_;
wire _13523_;
wire _13524_;
wire _13525_;
wire _13526_;
wire _13527_;
wire _13528_;
wire _13529_;
wire _13530_;
wire _13531_;
wire _13532_;
wire _13533_;
wire _13534_;
wire _13535_;
wire _13536_;
wire _13537_;
wire _13538_;
wire _13539_;
wire _13540_;
wire _13541_;
wire _13542_;
wire _13543_;
wire _13544_;
wire _13545_;
wire _13546_;
wire _13547_;
wire _13548_;
wire _13549_;
wire _13550_;
wire _13551_;
wire _13552_;
wire _13553_;
wire _13554_;
wire _13555_;
wire _13556_;
wire _13557_;
wire _13558_;
wire _13559_;
wire _13560_;
wire _13561_;
wire _13562_;
wire _13563_;
wire _13564_;
wire _13565_;
wire _13566_;
wire _13567_;
wire _13568_;
wire _13569_;
wire _13570_;
wire _13571_;
wire _13572_;
wire _13573_;
wire _13574_;
wire _13575_;
wire _13576_;
wire _13577_;
wire _13578_;
wire _13579_;
wire _13580_;
wire _13581_;
wire _13582_;
wire _13583_;
wire _13584_;
wire _13585_;
wire _13586_;
wire _13587_;
wire _13588_;
wire _13589_;
wire _13590_;
wire _13591_;
wire _13592_;
wire _13593_;
wire _13594_;
wire _13595_;
wire _13596_;
wire _13597_;
wire _13598_;
wire _13599_;
wire _13600_;
wire _13601_;
wire _13602_;
wire _13603_;
wire _13604_;
wire _13605_;
wire _13606_;
wire _13607_;
wire _13608_;
wire _13609_;
wire _13610_;
wire _13611_;
wire _13612_;
wire _13613_;
wire _13614_;
wire _13615_;
wire _13616_;
wire _13617_;
wire _13618_;
wire _13619_;
wire _13620_;
wire _13621_;
wire _13622_;
wire _13623_;
wire _13624_;
wire _13625_;
wire _13626_;
wire _13627_;
wire _13628_;
wire _13629_;
wire _13630_;
wire _13631_;
wire _13632_;
wire _13633_;
wire _13634_;
wire _13635_;
wire _13636_;
wire _13637_;
wire _13638_;
wire _13639_;
wire _13640_;
wire _13641_;
wire _13642_;
wire _13643_;
wire _13644_;
wire _13645_;
wire _13646_;
wire _13647_;
wire _13648_;
wire _13649_;
wire _13650_;
wire _13651_;
wire _13652_;
wire _13653_;
wire _13654_;
wire _13655_;
wire _13656_;
wire _13657_;
wire _13658_;
wire _13659_;
wire _13660_;
wire _13661_;
wire _13662_;
wire _13663_;
wire _13664_;
wire _13665_;
wire _13666_;
wire _13667_;
wire _13668_;
wire _13669_;
wire _13670_;
wire _13671_;
wire _13672_;
wire _13673_;
wire _13674_;
wire _13675_;
wire _13676_;
wire _13677_;
wire _13678_;
wire _13679_;
wire _13680_;
wire _13681_;
wire _13682_;
wire _13683_;
wire _13684_;
wire _13685_;
wire _13686_;
wire _13687_;
wire _13688_;
wire _13689_;
wire _13690_;
wire _13691_;
wire _13692_;
wire _13693_;
wire _13694_;
wire _13695_;
wire _13696_;
wire _13697_;
wire _13698_;
wire _13699_;
wire _13700_;
wire _13701_;
wire _13702_;
wire _13703_;
wire _13704_;
wire _13705_;
wire _13706_;
wire _13707_;
wire _13708_;
wire _13709_;
wire _13710_;
wire _13711_;
wire _13712_;
wire _13713_;
wire _13714_;
wire _13715_;
wire _13716_;
wire _13717_;
wire _13718_;
wire _13719_;
wire _13720_;
wire _13721_;
wire _13722_;
wire _13723_;
wire _13724_;
wire _13725_;
wire _13726_;
wire _13727_;
wire _13728_;
wire _13729_;
wire _13730_;
wire _13731_;
wire _13732_;
wire _13733_;
wire _13734_;
wire _13735_;
wire _13736_;
wire _13737_;
wire _13738_;
wire _13739_;
wire _13740_;
wire _13741_;
wire _13742_;
wire _13743_;
wire _13744_;
wire _13745_;
wire _13746_;
wire _13747_;
wire _13748_;
wire _13749_;
wire _13750_;
wire _13751_;
wire _13752_;
wire _13753_;
wire _13754_;
wire _13755_;
wire _13756_;
wire _13757_;
wire _13758_;
wire _13759_;
wire _13760_;
wire _13761_;
wire _13762_;
wire _13763_;
wire _13764_;
wire _13765_;
wire _13766_;
wire _13767_;
wire _13768_;
wire _13769_;
wire _13770_;
wire _13771_;
wire _13772_;
wire _13773_;
wire _13774_;
wire _13775_;
wire _13776_;
wire _13777_;
wire _13778_;
wire _13779_;
wire _13780_;
wire _13781_;
wire _13782_;
wire _13783_;
wire _13784_;
wire _13785_;
wire _13786_;
wire _13787_;
wire _13788_;
wire _13789_;
wire _13790_;
wire _13791_;
wire _13792_;
wire _13793_;
wire _13794_;
wire _13795_;
wire _13796_;
wire _13797_;
wire _13798_;
wire _13799_;
wire _13800_;
wire _13801_;
wire _13802_;
wire _13803_;
wire _13804_;
wire _13805_;
wire _13806_;
wire _13807_;
wire _13808_;
wire _13809_;
wire _13810_;
wire _13811_;
wire _13812_;
wire _13813_;
wire _13814_;
wire _13815_;
wire _13816_;
wire _13817_;
wire _13818_;
wire _13819_;
wire _13820_;
wire _13821_;
wire _13822_;
wire _13823_;
wire _13824_;
wire _13825_;
wire _13826_;
wire _13827_;
wire _13828_;
wire _13829_;
wire _13830_;
wire _13831_;
wire _13832_;
wire _13833_;
wire _13834_;
wire _13835_;
wire _13836_;
wire _13837_;
wire _13838_;
wire _13839_;
wire _13840_;
wire _13841_;
wire _13842_;
wire _13843_;
wire _13844_;
wire _13845_;
wire _13846_;
wire _13847_;
wire _13848_;
wire _13849_;
wire _13850_;
wire _13851_;
wire _13852_;
wire _13853_;
wire _13854_;
wire _13855_;
wire _13856_;
wire _13857_;
wire _13858_;
wire _13859_;
wire _13860_;
wire _13861_;
wire _13862_;
wire _13863_;
wire _13864_;
wire _13865_;
wire _13866_;
wire _13867_;
wire _13868_;
wire _13869_;
wire _13870_;
wire _13871_;
wire _13872_;
wire _13873_;
wire _13874_;
wire _13875_;
wire _13876_;
wire _13877_;
wire _13878_;
wire _13879_;
wire _13880_;
wire _13881_;
wire _13882_;
wire _13883_;
wire _13884_;
wire _13885_;
wire _13886_;
wire _13887_;
wire _13888_;
wire _13889_;
wire _13890_;
wire _13891_;
wire _13892_;
wire _13893_;
wire _13894_;
wire _13895_;
wire _13896_;
wire _13897_;
wire _13898_;
wire _13899_;
wire _13900_;
wire _13901_;
wire _13902_;
wire _13903_;
wire _13904_;
wire _13905_;
wire _13906_;
wire _13907_;
wire _13908_;
wire _13909_;
wire _13910_;
wire _13911_;
wire _13912_;
wire _13913_;
wire _13914_;
wire _13915_;
wire _13916_;
wire _13917_;
wire _13918_;
wire _13919_;
wire _13920_;
wire _13921_;
wire _13922_;
wire _13923_;
wire _13924_;
wire _13925_;
wire _13926_;
wire _13927_;
wire _13928_;
wire _13929_;
wire _13930_;
wire _13931_;
wire _13932_;
wire _13933_;
wire _13934_;
wire _13935_;
wire _13936_;
wire _13937_;
wire _13938_;
wire _13939_;
wire _13940_;
wire _13941_;
wire _13942_;
wire _13943_;
wire _13944_;
wire _13945_;
wire _13946_;
wire _13947_;
wire _13948_;
wire _13949_;
wire _13950_;
wire _13951_;
wire _13952_;
wire _13953_;
wire _13954_;
wire _13955_;
wire _13956_;
wire _13957_;
wire _13958_;
wire _13959_;
wire _13960_;
wire _13961_;
wire _13962_;
wire _13963_;
wire _13964_;
wire _13965_;
wire _13966_;
wire _13967_;
wire _13968_;
wire _13969_;
wire _13970_;
wire _13971_;
wire _13972_;
wire _13973_;
wire _13974_;
wire _13975_;
wire _13976_;
wire _13977_;
wire _13978_;
wire _13979_;
wire _13980_;
wire _13981_;
wire _13982_;
wire _13983_;
wire _13984_;
wire _13985_;
wire _13986_;
wire _13987_;
wire _13988_;
wire _13989_;
wire _13990_;
wire _13991_;
wire _13992_;
wire _13993_;
wire _13994_;
wire _13995_;
wire _13996_;
wire _13997_;
wire _13998_;
wire _13999_;
wire _14000_;
wire _14001_;
wire _14002_;
wire _14003_;
wire _14004_;
wire _14005_;
wire _14006_;
wire _14007_;
wire _14008_;
wire _14009_;
wire _14010_;
wire _14011_;
wire _14012_;
wire _14013_;
wire _14014_;
wire _14015_;
wire _14016_;
wire _14017_;
wire _14018_;
wire _14019_;
wire _14020_;
wire _14021_;
wire _14022_;
wire _14023_;
wire _14024_;
wire _14025_;
wire _14026_;
wire _14027_;
wire _14028_;
wire _14029_;
wire _14030_;
wire _14031_;
wire _14032_;
wire _14033_;
wire _14034_;
wire _14035_;
wire _14036_;
wire _14037_;
wire _14038_;
wire _14039_;
wire _14040_;
wire _14041_;
wire _14042_;
wire _14043_;
wire _14044_;
wire _14045_;
wire _14046_;
wire _14047_;
wire _14048_;
wire _14049_;
wire _14050_;
wire _14051_;
wire _14052_;
wire _14053_;
wire _14054_;
wire _14055_;
wire _14056_;
wire _14057_;
wire _14058_;
wire _14059_;
wire _14060_;
wire _14061_;
wire _14062_;
wire _14063_;
wire _14064_;
wire _14065_;
wire _14066_;
wire _14067_;
wire _14068_;
wire _14069_;
wire _14070_;
wire _14071_;
wire _14072_;
wire _14073_;
wire _14074_;
wire _14075_;
wire _14076_;
wire _14077_;
wire _14078_;
wire _14079_;
wire _14080_;
wire _14081_;
wire _14082_;
wire _14083_;
wire _14084_;
wire _14085_;
wire _14086_;
wire _14087_;
wire _14088_;
wire _14089_;
wire _14090_;
wire _14091_;
wire _14092_;
wire _14093_;
wire _14094_;
wire _14095_;
wire _14096_;
wire _14097_;
wire _14098_;
wire _14099_;
wire _14100_;
wire _14101_;
wire _14102_;
wire _14103_;
wire _14104_;
wire _14105_;
wire _14106_;
wire _14107_;
wire _14108_;
wire _14109_;
wire _14110_;
wire _14111_;
wire _14112_;
wire _14113_;
wire _14114_;
wire _14115_;
wire _14116_;
wire _14117_;
wire _14118_;
wire _14119_;
wire _14120_;
wire _14121_;
wire _14122_;
wire _14123_;
wire _14124_;
wire _14125_;
wire _14126_;
wire _14127_;
wire _14128_;
wire _14129_;
wire _14130_;
wire _14131_;
wire _14132_;
wire _14133_;
wire _14134_;
wire _14135_;
wire _14136_;
wire _14137_;
wire _14138_;
wire _14139_;
wire _14140_;
wire _14141_;
wire _14142_;
wire _14143_;
wire _14144_;
wire _14145_;
wire _14146_;
wire _14147_;
wire _14148_;
wire _14149_;
wire _14150_;
wire _14151_;
wire _14152_;
wire _14153_;
wire _14154_;
wire _14155_;
wire _14156_;
wire _14157_;
wire _14158_;
wire _14159_;
wire _14160_;
wire _14161_;
wire _14162_;
wire _14163_;
wire _14164_;
wire _14165_;
wire _14166_;
wire _14167_;
wire _14168_;
wire _14169_;
wire _14170_;
wire _14171_;
wire _14172_;
wire _14173_;
wire _14174_;
wire _14175_;
wire _14176_;
wire _14177_;
wire _14178_;
wire _14179_;
wire _14180_;
wire _14181_;
wire _14182_;
wire _14183_;
wire _14184_;
wire _14185_;
wire _14186_;
wire _14187_;
wire _14188_;
wire _14189_;
wire _14190_;
wire _14191_;
wire _14192_;
wire _14193_;
wire _14194_;
wire _14195_;
wire _14196_;
wire _14197_;
wire _14198_;
wire _14199_;
wire _14200_;
wire _14201_;
wire _14202_;
wire _14203_;
wire _14204_;
wire _14205_;
wire _14206_;
wire _14207_;
wire _14208_;
wire _14209_;
wire _14210_;
wire _14211_;
wire _14212_;
wire _14213_;
wire _14214_;
wire _14215_;
wire _14216_;
wire _14217_;
wire _14218_;
wire _14219_;
wire _14220_;
wire _14221_;
wire _14222_;
wire _14223_;
wire _14224_;
wire _14225_;
wire _14226_;
wire _14227_;
wire _14228_;
wire _14229_;
wire _14230_;
wire _14231_;
wire _14232_;
wire _14233_;
wire _14234_;
wire _14235_;
wire _14236_;
wire _14237_;
wire _14238_;
wire _14239_;
wire _14240_;
wire _14241_;
wire _14242_;
wire _14243_;
wire _14244_;
wire _14245_;
wire _14246_;
wire _14247_;
wire _14248_;
wire _14249_;
wire _14250_;
wire _14251_;
wire _14252_;
wire _14253_;
wire _14254_;
wire _14255_;
wire _14256_;
wire _14257_;
wire _14258_;
wire _14259_;
wire _14260_;
wire _14261_;
wire _14262_;
wire _14263_;
wire _14264_;
wire _14265_;
wire _14266_;
wire _14267_;
wire _14268_;
wire _14269_;
wire _14270_;
wire _14271_;
wire _14272_;
wire _14273_;
wire _14274_;
wire _14275_;
wire _14276_;
wire _14277_;
wire _14278_;
wire _14279_;
wire _14280_;
wire _14281_;
wire _14282_;
wire _14283_;
wire _14284_;
wire _14285_;
wire _14286_;
wire _14287_;
wire _14288_;
wire _14289_;
wire _14290_;
wire _14291_;
wire _14292_;
wire _14293_;
wire _14294_;
wire _14295_;
wire _14296_;
wire _14297_;
wire _14298_;
wire _14299_;
wire _14300_;
wire _14301_;
wire _14302_;
wire _14303_;
wire _14304_;
wire _14305_;
wire _14306_;
wire _14307_;
wire _14308_;
wire _14309_;
wire _14310_;
wire _14311_;
wire _14312_;
wire _14313_;
wire _14314_;
wire _14315_;
wire _14316_;
wire _14317_;
wire _14318_;
wire _14319_;
wire _14320_;
wire _14321_;
wire _14322_;
wire _14323_;
wire _14324_;
wire _14325_;
wire _14326_;
wire _14327_;
wire _14328_;
wire _14329_;
wire _14330_;
wire _14331_;
wire _14332_;
wire _14333_;
wire _14334_;
wire _14335_;
wire _14336_;
wire _14337_;
wire _14338_;
wire _14339_;
wire _14340_;
wire _14341_;
wire _14342_;
wire _14343_;
wire _14344_;
wire _14345_;
wire _14346_;
wire _14347_;
wire _14348_;
wire _14349_;
wire _14350_;
wire _14351_;
wire _14352_;
wire _14353_;
wire _14354_;
wire _14355_;
wire _14356_;
wire _14357_;
wire _14358_;
wire _14359_;
wire _14360_;
wire _14361_;
wire _14362_;
wire _14363_;
wire _14364_;
wire _14365_;
wire _14366_;
wire _14367_;
wire _14368_;
wire _14369_;
wire _14370_;
wire _14371_;
wire _14372_;
wire _14373_;
wire _14374_;
wire _14375_;
wire _14376_;
wire _14377_;
wire _14378_;
wire _14379_;
wire _14380_;
wire _14381_;
wire _14382_;
wire _14383_;
wire _14384_;
wire _14385_;
wire _14386_;
wire _14387_;
wire _14388_;
wire _14389_;
wire _14390_;
wire _14391_;
wire _14392_;
wire _14393_;
wire _14394_;
wire _14395_;
wire _14396_;
wire _14397_;
wire _14398_;
wire _14399_;
wire _14400_;
wire _14401_;
wire _14402_;
wire _14403_;
wire _14404_;
wire _14405_;
wire _14406_;
wire _14407_;
wire _14408_;
wire _14409_;
wire _14410_;
wire _14411_;
wire _14412_;
wire _14413_;
wire _14414_;
wire _14415_;
wire _14416_;
wire _14417_;
wire _14418_;
wire _14419_;
wire _14420_;
wire _14421_;
wire _14422_;
wire _14423_;
wire _14424_;
wire _14425_;
wire _14426_;
wire _14427_;
wire _14428_;
wire _14429_;
wire _14430_;
wire _14431_;
wire _14432_;
wire _14433_;
wire _14434_;
wire _14435_;
wire _14436_;
wire _14437_;
wire _14438_;
wire _14439_;
wire _14440_;
wire _14441_;
wire _14442_;
wire _14443_;
wire _14444_;
wire _14445_;
wire _14446_;
wire _14447_;
wire _14448_;
wire _14449_;
wire _14450_;
wire _14451_;
wire _14452_;
wire _14453_;
wire _14454_;
wire _14455_;
wire _14456_;
wire _14457_;
wire _14458_;
wire _14459_;
wire _14460_;
wire _14461_;
wire _14462_;
wire _14463_;
wire _14464_;
wire _14465_;
wire _14466_;
wire _14467_;
wire _14468_;
wire _14469_;
wire _14470_;
wire _14471_;
wire _14472_;
wire _14473_;
wire _14474_;
wire _14475_;
wire _14476_;
wire _14477_;
wire _14478_;
wire _14479_;
wire _14480_;
wire _14481_;
wire _14482_;
wire _14483_;
wire _14484_;
wire _14485_;
wire _14486_;
wire _14487_;
wire _14488_;
wire _14489_;
wire _14490_;
wire _14491_;
wire _14492_;
wire _14493_;
wire _14494_;
wire _14495_;
wire _14496_;
wire _14497_;
wire _14498_;
wire _14499_;
wire _14500_;
wire _14501_;
wire _14502_;
wire _14503_;
wire _14504_;
wire _14505_;
wire _14506_;
wire _14507_;
wire _14508_;
wire _14509_;
wire _14510_;
wire _14511_;
wire _14512_;
wire _14513_;
wire _14514_;
wire _14515_;
wire _14516_;
wire _14517_;
wire _14518_;
wire _14519_;
wire _14520_;
wire _14521_;
wire _14522_;
wire _14523_;
wire _14524_;
wire _14525_;
wire _14526_;
wire _14527_;
wire _14528_;
wire _14529_;
wire _14530_;
wire _14531_;
wire _14532_;
wire _14533_;
wire _14534_;
wire _14535_;
wire _14536_;
wire _14537_;
wire _14538_;
wire _14539_;
wire _14540_;
wire _14541_;
wire _14542_;
wire _14543_;
wire _14544_;
wire _14545_;
wire _14546_;
wire _14547_;
wire _14548_;
wire _14549_;
wire _14550_;
wire _14551_;
wire _14552_;
wire _14553_;
wire _14554_;
wire _14555_;
wire _14556_;
wire _14557_;
wire _14558_;
wire _14559_;
wire _14560_;
wire _14561_;
wire _14562_;
wire _14563_;
wire _14564_;
wire _14565_;
wire _14566_;
wire _14567_;
wire _14568_;
wire _14569_;
wire _14570_;
wire _14571_;
wire _14572_;
wire _14573_;
wire _14574_;
wire _14575_;
wire _14576_;
wire _14577_;
wire _14578_;
wire _14579_;
wire _14580_;
wire _14581_;
wire _14582_;
wire _14583_;
wire _14584_;
wire _14585_;
wire _14586_;
wire _14587_;
wire _14588_;
wire _14589_;
wire _14590_;
wire _14591_;
wire _14592_;
wire _14593_;
wire _14594_;
wire _14595_;
wire _14596_;
wire _14597_;
wire _14598_;
wire _14599_;
wire _14600_;
wire _14601_;
wire _14602_;
wire _14603_;
wire _14604_;
wire _14605_;
wire _14606_;
wire _14607_;
wire _14608_;
wire _14609_;
wire _14610_;
wire _14611_;
wire _14612_;
wire _14613_;
wire _14614_;
wire _14615_;
wire _14616_;
wire _14617_;
wire _14618_;
wire _14619_;
wire _14620_;
wire _14621_;
wire _14622_;
wire _14623_;
wire _14624_;
wire _14625_;
wire _14626_;
wire _14627_;
wire _14628_;
wire _14629_;
wire _14630_;
wire _14631_;
wire _14632_;
wire _14633_;
wire _14634_;
wire _14635_;
wire _14636_;
wire _14637_;
wire _14638_;
wire _14639_;
wire _14640_;
wire _14641_;
wire _14642_;
wire _14643_;
wire _14644_;
wire _14645_;
wire _14646_;
wire _14647_;
wire _14648_;
wire _14649_;
wire _14650_;
wire _14651_;
wire _14652_;
wire _14653_;
wire _14654_;
wire _14655_;
wire _14656_;
wire _14657_;
wire _14658_;
wire _14659_;
wire _14660_;
wire _14661_;
wire _14662_;
wire _14663_;
wire _14664_;
wire _14665_;
wire _14666_;
wire _14667_;
wire _14668_;
wire _14669_;
wire _14670_;
wire _14671_;
wire _14672_;
wire _14673_;
wire _14674_;
wire _14675_;
wire _14676_;
wire _14677_;
wire _14678_;
wire _14679_;
wire _14680_;
wire _14681_;
wire _14682_;
wire _14683_;
wire _14684_;
wire _14685_;
wire _14686_;
wire _14687_;
wire _14688_;
wire _14689_;
wire _14690_;
wire _14691_;
wire _14692_;
wire _14693_;
wire _14694_;
wire _14695_;
wire _14696_;
wire _14697_;
wire _14698_;
wire _14699_;
wire _14700_;
wire _14701_;
wire _14702_;
wire _14703_;
wire _14704_;
wire _14705_;
wire _14706_;
wire _14707_;
wire _14708_;
wire _14709_;
wire _14710_;
wire _14711_;
wire _14712_;
wire _14713_;
wire _14714_;
wire _14715_;
wire _14716_;
wire _14717_;
wire _14718_;
wire _14719_;
wire _14720_;
wire _14721_;
wire _14722_;
wire _14723_;
wire _14724_;
wire _14725_;
wire _14726_;
wire _14727_;
wire _14728_;
wire _14729_;
wire _14730_;
wire _14731_;
wire _14732_;
wire _14733_;
wire _14734_;
wire _14735_;
wire _14736_;
wire _14737_;
wire _14738_;
wire _14739_;
wire _14740_;
wire _14741_;
wire _14742_;
wire _14743_;
wire _14744_;
wire _14745_;
wire _14746_;
wire _14747_;
wire _14748_;
wire _14749_;
wire _14750_;
wire _14751_;
wire _14752_;
wire _14753_;
wire _14754_;
wire _14755_;
wire _14756_;
wire _14757_;
wire _14758_;
wire _14759_;
wire _14760_;
wire _14761_;
wire _14762_;
wire _14763_;
wire _14764_;
wire _14765_;
wire _14766_;
wire _14767_;
wire _14768_;
wire _14769_;
wire _14770_;
wire _14771_;
wire _14772_;
wire _14773_;
wire _14774_;
wire _14775_;
wire _14776_;
wire _14777_;
wire _14778_;
wire _14779_;
wire _14780_;
wire _14781_;
wire _14782_;
wire _14783_;
wire _14784_;
wire _14785_;
wire _14786_;
wire _14787_;
wire _14788_;
wire _14789_;
wire _14790_;
wire _14791_;
wire _14792_;
wire _14793_;
wire _14794_;
wire _14795_;
wire _14796_;
wire _14797_;
wire _14798_;
wire _14799_;
wire _14800_;
wire _14801_;
wire _14802_;
wire _14803_;
wire _14804_;
wire _14805_;
wire _14806_;
wire _14807_;
wire _14808_;
wire _14809_;
wire _14810_;
wire _14811_;
wire _14812_;
wire _14813_;
wire _14814_;
wire _14815_;
wire _14816_;
wire _14817_;
wire _14818_;
wire _14819_;
wire _14820_;
wire _14821_;
wire _14822_;
wire _14823_;
wire _14824_;
wire _14825_;
wire _14826_;
wire _14827_;
wire _14828_;
wire _14829_;
wire _14830_;
wire _14831_;
wire _14832_;
wire _14833_;
wire _14834_;
wire _14835_;
wire _14836_;
wire _14837_;
wire _14838_;
wire _14839_;
wire _14840_;
wire _14841_;
wire _14842_;
wire _14843_;
wire _14844_;
wire _14845_;
wire _14846_;
wire _14847_;
wire _14848_;
wire _14849_;
wire _14850_;
wire _14851_;
wire _14852_;
wire _14853_;
wire _14854_;
wire _14855_;
wire _14856_;
wire _14857_;
wire _14858_;
wire _14859_;
wire _14860_;
wire _14861_;
wire _14862_;
wire _14863_;
wire _14864_;
wire _14865_;
wire _14866_;
wire _14867_;
wire _14868_;
wire _14869_;
wire _14870_;
wire _14871_;
wire _14872_;
wire _14873_;
wire _14874_;
wire _14875_;
wire _14876_;
wire _14877_;
wire _14878_;
wire _14879_;
wire _14880_;
wire _14881_;
wire _14882_;
wire _14883_;
wire _14884_;
wire _14885_;
wire _14886_;
wire _14887_;
wire _14888_;
wire _14889_;
wire _14890_;
wire _14891_;
wire _14892_;
wire _14893_;
wire _14894_;
wire _14895_;
wire _14896_;
wire _14897_;
wire _14898_;
wire _14899_;
wire _14900_;
wire _14901_;
wire _14902_;
wire _14903_;
wire _14904_;
wire _14905_;
wire _14906_;
wire _14907_;
wire _14908_;
wire _14909_;
wire _14910_;
wire _14911_;
wire _14912_;
wire _14913_;
wire _14914_;
wire _14915_;
wire _14916_;
wire _14917_;
wire _14918_;
wire _14919_;
wire _14920_;
wire _14921_;
wire _14922_;
wire _14923_;
wire _14924_;
wire _14925_;
wire _14926_;
wire _14927_;
wire _14928_;
wire _14929_;
wire _14930_;
wire _14931_;
wire _14932_;
wire _14933_;
wire _14934_;
wire _14935_;
wire _14936_;
wire _14937_;
wire _14938_;
wire _14939_;
wire _14940_;
wire _14941_;
wire _14942_;
wire _14943_;
wire _14944_;
wire _14945_;
wire _14946_;
wire _14947_;
wire _14948_;
wire _14949_;
wire _14950_;
wire _14951_;
wire _14952_;
wire _14953_;
wire _14954_;
wire _14955_;
wire _14956_;
wire _14957_;
wire _14958_;
wire _14959_;
wire _14960_;
wire _14961_;
wire _14962_;
wire _14963_;
wire _14964_;
wire _14965_;
wire _14966_;
wire _14967_;
wire _14968_;
wire _14969_;
wire _14970_;
wire _14971_;
wire _14972_;
wire _14973_;
wire _14974_;
wire _14975_;
wire _14976_;
wire _14977_;
wire _14978_;
wire _14979_;
wire _14980_;
wire _14981_;
wire _14982_;
wire _14983_;
wire _14984_;
wire _14985_;
wire _14986_;
wire _14987_;
wire _14988_;
wire _14989_;
wire _14990_;
wire _14991_;
wire _14992_;
wire _14993_;
wire _14994_;
wire _14995_;
wire _14996_;
wire _14997_;
wire _14998_;
wire _14999_;
wire _15000_;
wire _15001_;
wire _15002_;
wire _15003_;
wire _15004_;
wire _15005_;
wire _15006_;
wire _15007_;
wire _15008_;
wire _15009_;
wire _15010_;
wire _15011_;
wire _15012_;
wire _15013_;
wire _15014_;
wire _15015_;
wire _15016_;
wire _15017_;
wire _15018_;
wire _15019_;
wire _15020_;
wire _15021_;
wire _15022_;
wire _15023_;
wire _15024_;
wire _15025_;
wire _15026_;
wire _15027_;
wire _15028_;
wire _15029_;
wire _15030_;
wire _15031_;
wire _15032_;
wire _15033_;
wire _15034_;
wire _15035_;
wire _15036_;
wire _15037_;
wire _15038_;
wire _15039_;
wire _15040_;
wire _15041_;
wire _15042_;
wire _15043_;
wire _15044_;
wire _15045_;
wire _15046_;
wire _15047_;
wire _15048_;
wire _15049_;
wire _15050_;
wire _15051_;
wire _15052_;
wire _15053_;
wire _15054_;
wire _15055_;
wire _15056_;
wire _15057_;
wire _15058_;
wire _15059_;
wire _15060_;
wire _15061_;
wire _15062_;
wire _15063_;
wire _15064_;
wire _15065_;
wire _15066_;
wire _15067_;
wire _15068_;
wire _15069_;
wire _15070_;
wire _15071_;
wire _15072_;
wire _15073_;
wire _15074_;
wire _15075_;
wire _15076_;
wire _15077_;
wire _15078_;
wire _15079_;
wire _15080_;
wire _15081_;
wire _15082_;
wire _15083_;
wire _15084_;
wire _15085_;
wire _15086_;
wire _15087_;
wire _15088_;
wire _15089_;
wire _15090_;
wire _15091_;
wire _15092_;
wire _15093_;
wire _15094_;
wire _15095_;
wire _15096_;
wire _15097_;
wire _15098_;
wire _15099_;
wire _15100_;
wire _15101_;
wire _15102_;
wire _15103_;
wire _15104_;
wire _15105_;
wire _15106_;
wire _15107_;
wire _15108_;
wire _15109_;
wire _15110_;
wire _15111_;
wire _15112_;
wire _15113_;
wire _15114_;
wire _15115_;
wire _15116_;
wire _15117_;
wire _15118_;
wire _15119_;
wire _15120_;
wire _15121_;
wire _15122_;
wire _15123_;
wire _15124_;
wire _15125_;
wire _15126_;
wire _15127_;
wire _15128_;
wire _15129_;
wire _15130_;
wire _15131_;
wire _15132_;
wire _15133_;
wire _15134_;
wire _15135_;
wire _15136_;
wire _15137_;
wire _15138_;
wire _15139_;
wire _15140_;
wire _15141_;
wire _15142_;
wire _15143_;
wire _15144_;
wire _15145_;
wire _15146_;
wire _15147_;
wire _15148_;
wire _15149_;
wire _15150_;
wire _15151_;
wire _15152_;
wire _15153_;
wire _15154_;
wire _15155_;
wire _15156_;
wire _15157_;
wire _15158_;
wire _15159_;
wire _15160_;
wire _15161_;
wire _15162_;
wire _15163_;
wire _15164_;
wire _15165_;
wire _15166_;
wire _15167_;
wire _15168_;
wire _15169_;
wire _15170_;
wire _15171_;
wire _15172_;
wire _15173_;
wire _15174_;
wire _15175_;
wire _15176_;
wire _15177_;
wire _15178_;
wire _15179_;
wire _15180_;
wire _15181_;
wire _15182_;
wire _15183_;
wire _15184_;
wire _15185_;
wire _15186_;
wire _15187_;
wire _15188_;
wire _15189_;
wire _15190_;
wire _15191_;
wire _15192_;
wire _15193_;
wire _15194_;
wire _15195_;
wire _15196_;
wire _15197_;
wire _15198_;
wire _15199_;
wire _15200_;
wire _15201_;
wire _15202_;
wire _15203_;
wire _15204_;
wire _15205_;
wire _15206_;
wire _15207_;
wire _15208_;
wire _15209_;
wire _15210_;
wire _15211_;
wire _15212_;
wire _15213_;
wire _15214_;
wire _15215_;
wire _15216_;
wire _15217_;
wire _15218_;
wire _15219_;
wire _15220_;
wire _15221_;
wire _15222_;
wire _15223_;
wire _15224_;
wire _15225_;
wire _15226_;
wire _15227_;
wire _15228_;
wire _15229_;
wire _15230_;
wire _15231_;
wire _15232_;
wire _15233_;
wire _15234_;
wire _15235_;
wire _15236_;
wire _15237_;
wire _15238_;
wire _15239_;
wire _15240_;
wire _15241_;
wire _15242_;
wire _15243_;
wire _15244_;
wire _15245_;
wire _15246_;
wire _15247_;
wire _15248_;
wire _15249_;
wire _15250_;
wire _15251_;
wire _15252_;
wire _15253_;
wire _15254_;
wire _15255_;
wire _15256_;
wire _15257_;
wire _15258_;
wire _15259_;
wire _15260_;
wire _15261_;
wire _15262_;
wire _15263_;
wire _15264_;
wire _15265_;
wire _15266_;
wire _15267_;
wire _15268_;
wire _15269_;
wire _15270_;
wire _15271_;
wire _15272_;
wire _15273_;
wire _15274_;
wire _15275_;
wire _15276_;
wire _15277_;
wire _15278_;
wire _15279_;
wire _15280_;
wire _15281_;
wire _15282_;
wire _15283_;
wire _15284_;
wire _15285_;
wire _15286_;
wire _15287_;
wire _15288_;
wire _15289_;
wire _15290_;
wire _15291_;
wire _15292_;
wire _15293_;
wire _15294_;
wire _15295_;
wire _15296_;
wire _15297_;
wire _15298_;
wire _15299_;
wire _15300_;
wire _15301_;
wire _15302_;
wire _15303_;
wire _15304_;
wire _15305_;
wire _15306_;
wire _15307_;
wire _15308_;
wire _15309_;
wire _15310_;
wire _15311_;
wire _15312_;
wire _15313_;
wire _15314_;
wire _15315_;
wire _15316_;
wire _15317_;
wire _15318_;
wire _15319_;
wire _15320_;
wire _15321_;
wire _15322_;
wire _15323_;
wire _15324_;
wire _15325_;
wire _15326_;
wire _15327_;
wire _15328_;
wire _15329_;
wire _15330_;
wire _15331_;
wire _15332_;
wire _15333_;
wire _15334_;
wire _15335_;
wire _15336_;
wire _15337_;
wire _15338_;
wire _15339_;
wire _15340_;
wire _15341_;
wire _15342_;
wire _15343_;
wire _15344_;
wire _15345_;
wire _15346_;
wire _15347_;
wire _15348_;
wire _15349_;
wire _15350_;
wire _15351_;
wire _15352_;
wire _15353_;
wire _15354_;
wire _15355_;
wire _15356_;
wire _15357_;
wire _15358_;
wire _15359_;
wire _15360_;
wire _15361_;
wire _15362_;
wire _15363_;
wire _15364_;
wire _15365_;
wire _15366_;
wire _15367_;
wire _15368_;
wire _15369_;
wire _15370_;
wire _15371_;
wire _15372_;
wire _15373_;
wire _15374_;
wire _15375_;
wire _15376_;
wire _15377_;
wire _15378_;
wire _15379_;
wire _15380_;
wire _15381_;
wire _15382_;
wire _15383_;
wire _15384_;
wire _15385_;
wire _15386_;
wire _15387_;
wire _15388_;
wire _15389_;
wire _15390_;
wire _15391_;
wire _15392_;
wire _15393_;
wire _15394_;
wire _15395_;
wire _15396_;
wire _15397_;
wire _15398_;
wire _15399_;
wire _15400_;
wire _15401_;
wire _15402_;
wire _15403_;
wire _15404_;
wire _15405_;
wire _15406_;
wire _15407_;
wire _15408_;
wire _15409_;
wire _15410_;
wire _15411_;
wire _15412_;
wire _15413_;
wire _15414_;
wire _15415_;
wire _15416_;
wire _15417_;
wire _15418_;
wire _15419_;
wire _15420_;
wire _15421_;
wire _15422_;
wire _15423_;
wire _15424_;
wire _15425_;
wire _15426_;
wire _15427_;
wire _15428_;
wire _15429_;
wire _15430_;
wire _15431_;
wire _15432_;
wire _15433_;
wire _15434_;
wire _15435_;
wire _15436_;
wire _15437_;
wire _15438_;
wire _15439_;
wire _15440_;
wire _15441_;
wire _15442_;
wire _15443_;
wire _15444_;
wire _15445_;
wire _15446_;
wire _15447_;
wire _15448_;
wire _15449_;
wire _15450_;
wire _15451_;
wire _15452_;
wire _15453_;
wire _15454_;
wire _15455_;
wire _15456_;
wire _15457_;
wire _15458_;
wire _15459_;
wire _15460_;
wire _15461_;
wire _15462_;
wire _15463_;
wire _15464_;
wire _15465_;
wire _15466_;
wire _15467_;
wire _15468_;
wire _15469_;
wire _15470_;
wire _15471_;
wire _15472_;
wire _15473_;
wire _15474_;
wire _15475_;
wire _15476_;
wire _15477_;
wire _15478_;
wire _15479_;
wire _15480_;
wire _15481_;
wire _15482_;
wire _15483_;
wire _15484_;
wire _15485_;
wire _15486_;
wire _15487_;
wire _15488_;
wire _15489_;
wire _15490_;
wire _15491_;
wire _15492_;
wire _15493_;
wire _15494_;
wire _15495_;
wire _15496_;
wire _15497_;
wire _15498_;
wire _15499_;
wire _15500_;
wire _15501_;
wire _15502_;
wire _15503_;
wire _15504_;
wire _15505_;
wire _15506_;
wire _15507_;
wire _15508_;
wire _15509_;
wire _15510_;
wire _15511_;
wire _15512_;
wire _15513_;
wire _15514_;
wire _15515_;
wire _15516_;
wire _15517_;
wire _15518_;
wire _15519_;
wire _15520_;
wire _15521_;
wire _15522_;
wire _15523_;
wire _15524_;
wire _15525_;
wire _15526_;
wire _15527_;
wire _15528_;
wire _15529_;
wire _15530_;
wire _15531_;
wire _15532_;
wire _15533_;
wire _15534_;
wire _15535_;
wire _15536_;
wire _15537_;
wire _15538_;
wire _15539_;
wire _15540_;
wire _15541_;
wire _15542_;
wire _15543_;
wire _15544_;
wire _15545_;
wire _15546_;
wire _15547_;
wire _15548_;
wire _15549_;
wire _15550_;
wire _15551_;
wire _15552_;
wire _15553_;
wire _15554_;
wire _15555_;
wire _15556_;
wire _15557_;
wire _15558_;
wire _15559_;
wire _15560_;
wire _15561_;
wire _15562_;
wire _15563_;
wire _15564_;
wire _15565_;
wire _15566_;
wire _15567_;
wire _15568_;
wire _15569_;
wire _15570_;
wire _15571_;
wire _15572_;
wire _15573_;
wire _15574_;
wire _15575_;
wire _15576_;
wire _15577_;
wire _15578_;
wire _15579_;
wire _15580_;
wire _15581_;
wire _15582_;
wire _15583_;
wire _15584_;
wire _15585_;
wire _15586_;
wire _15587_;
wire _15588_;
wire _15589_;
wire _15590_;
wire _15591_;
wire _15592_;
wire _15593_;
wire _15594_;
wire _15595_;
wire _15596_;
wire _15597_;
wire _15598_;
wire _15599_;
wire _15600_;
wire _15601_;
wire _15602_;
wire _15603_;
wire _15604_;
wire _15605_;
wire _15606_;
wire _15607_;
wire _15608_;
wire _15609_;
wire _15610_;
wire _15611_;
wire _15612_;
wire _15613_;
wire _15614_;
wire _15615_;
wire _15616_;
wire _15617_;
wire _15618_;
wire _15619_;
wire _15620_;
wire _15621_;
wire _15622_;
wire _15623_;
wire _15624_;
wire _15625_;
wire _15626_;
wire _15627_;
wire _15628_;
wire _15629_;
wire _15630_;
wire _15631_;
wire _15632_;
wire _15633_;
wire _15634_;
wire _15635_;
wire _15636_;
wire _15637_;
wire _15638_;
wire _15639_;
wire _15640_;
wire _15641_;
wire _15642_;
wire _15643_;
wire _15644_;
wire _15645_;
wire _15646_;
wire _15647_;
wire _15648_;
wire _15649_;
wire _15650_;
wire _15651_;
wire _15652_;
wire _15653_;
wire _15654_;
wire _15655_;
wire _15656_;
wire _15657_;
wire _15658_;
wire _15659_;
wire _15660_;
wire _15661_;
wire _15662_;
wire _15663_;
wire _15664_;
wire _15665_;
wire _15666_;
wire _15667_;
wire _15668_;
wire _15669_;
wire _15670_;
wire _15671_;
wire _15672_;
wire _15673_;
wire _15674_;
wire _15675_;
wire _15676_;
wire _15677_;
wire _15678_;
wire _15679_;
wire _15680_;
wire _15681_;
wire _15682_;
wire _15683_;
wire _15684_;
wire _15685_;
wire _15686_;
wire _15687_;
wire _15688_;
wire _15689_;
wire _15690_;
wire _15691_;
wire _15692_;
wire _15693_;
wire _15694_;
wire _15695_;
wire _15696_;
wire _15697_;
wire _15698_;
wire _15699_;
wire _15700_;
wire _15701_;
wire _15702_;
wire _15703_;
wire _15704_;
wire _15705_;
wire _15706_;
wire _15707_;
wire _15708_;
wire _15709_;
wire _15710_;
wire _15711_;
wire _15712_;
wire _15713_;
wire _15714_;
wire _15715_;
wire _15716_;
wire _15717_;
wire _15718_;
wire _15719_;
wire _15720_;
wire _15721_;
wire _15722_;
wire _15723_;
wire _15724_;
wire _15725_;
wire _15726_;
wire _15727_;
wire _15728_;
wire _15729_;
wire _15730_;
wire _15731_;
wire _15732_;
wire _15733_;
wire _15734_;
wire _15735_;
wire _15736_;
wire _15737_;
wire _15738_;
wire _15739_;
wire _15740_;
wire _15741_;
wire _15742_;
wire _15743_;
wire _15744_;
wire _15745_;
wire _15746_;
wire _15747_;
wire _15748_;
wire _15749_;
wire _15750_;
wire _15751_;
wire _15752_;
wire _15753_;
wire _15754_;
wire _15755_;
wire _15756_;
wire _15757_;
wire _15758_;
wire _15759_;
wire _15760_;
wire _15761_;
wire _15762_;
wire _15763_;
wire _15764_;
wire _15765_;
wire _15766_;
wire _15767_;
wire _15768_;
wire _15769_;
wire _15770_;
wire _15771_;
wire _15772_;
wire _15773_;
wire _15774_;
wire _15775_;
wire _15776_;
wire _15777_;
wire _15778_;
wire _15779_;
wire _15780_;
wire _15781_;
wire _15782_;
wire _15783_;
wire _15784_;
wire _15785_;
wire _15786_;
wire _15787_;
wire _15788_;
wire _15789_;
wire _15790_;
wire _15791_;
wire _15792_;
wire _15793_;
wire _15794_;
wire _15795_;
wire _15796_;
wire _15797_;
wire _15798_;
wire _15799_;
wire _15800_;
wire _15801_;
wire _15802_;
wire _15803_;
wire _15804_;
wire _15805_;
wire _15806_;
wire _15807_;
wire _15808_;
wire _15809_;
wire _15810_;
wire _15811_;
wire _15812_;
wire _15813_;
wire _15814_;
wire _15815_;
wire _15816_;
wire _15817_;
wire _15818_;
wire _15819_;
wire _15820_;
wire _15821_;
wire _15822_;
wire _15823_;
wire _15824_;
wire _15825_;
wire _15826_;
wire _15827_;
wire _15828_;
wire _15829_;
wire _15830_;
wire _15831_;
wire _15832_;
wire _15833_;
wire _15834_;
wire _15835_;
wire _15836_;
wire _15837_;
wire _15838_;
wire _15839_;
wire _15840_;
wire _15841_;
wire _15842_;
wire _15843_;
wire _15844_;
wire _15845_;
wire _15846_;
wire _15847_;
wire _15848_;
wire _15849_;
wire _15850_;
wire _15851_;
wire _15852_;
wire _15853_;
wire _15854_;
wire _15855_;
wire _15856_;
wire _15857_;
wire _15858_;
wire _15859_;
wire _15860_;
wire _15861_;
wire _15862_;
wire _15863_;
wire _15864_;
wire _15865_;
wire _15866_;
wire _15867_;
wire _15868_;
wire _15869_;
wire _15870_;
wire _15871_;
wire _15872_;
wire _15873_;
wire _15874_;
wire _15875_;
wire _15876_;
wire _15877_;
wire _15878_;
wire _15879_;
wire _15880_;
wire _15881_;
wire _15882_;
wire _15883_;
wire _15884_;
wire _15885_;
wire _15886_;
wire _15887_;
wire _15888_;
wire _15889_;
wire _15890_;
wire _15891_;
wire _15892_;
wire _15893_;
wire _15894_;
wire _15895_;
wire _15896_;
wire _15897_;
wire _15898_;
wire _15899_;
wire _15900_;
wire _15901_;
wire _15902_;
wire _15903_;
wire _15904_;
wire _15905_;
wire _15906_;
wire _15907_;
wire _15908_;
wire _15909_;
wire _15910_;
wire _15911_;
wire _15912_;
wire _15913_;
wire _15914_;
wire _15915_;
wire _15916_;
wire _15917_;
wire _15918_;
wire _15919_;
wire _15920_;
wire _15921_;
wire _15922_;
wire _15923_;
wire _15924_;
wire _15925_;
wire _15926_;
wire _15927_;
wire _15928_;
wire _15929_;
wire _15930_;
wire _15931_;
wire _15932_;
wire _15933_;
wire _15934_;
wire _15935_;
wire _15936_;
wire _15937_;
wire _15938_;
wire _15939_;
wire _15940_;
wire _15941_;
wire _15942_;
wire _15943_;
wire _15944_;
wire _15945_;
wire _15946_;
wire _15947_;
wire _15948_;
wire _15949_;
wire _15950_;
wire _15951_;
wire _15952_;
wire _15953_;
wire _15954_;
wire _15955_;
wire _15956_;
wire _15957_;
wire _15958_;
wire _15959_;
wire _15960_;
wire _15961_;
wire _15962_;
wire _15963_;
wire _15964_;
wire _15965_;
wire _15966_;
wire _15967_;
wire _15968_;
wire _15969_;
wire _15970_;
wire _15971_;
wire _15972_;
wire _15973_;
wire _15974_;
wire _15975_;
wire _15976_;
wire _15977_;
wire _15978_;
wire _15979_;
wire _15980_;
wire _15981_;
wire _15982_;
wire _15983_;
wire _15984_;
wire _15985_;
wire _15986_;
wire _15987_;
wire _15988_;
wire _15989_;
wire _15990_;
wire _15991_;
wire _15992_;
wire _15993_;
wire _15994_;
wire _15995_;
wire _15996_;
wire _15997_;
wire _15998_;
wire _15999_;
wire _16000_;
wire _16001_;
wire _16002_;
wire _16003_;
wire _16004_;
wire _16005_;
wire _16006_;
wire _16007_;
wire _16008_;
wire _16009_;
wire _16010_;
wire _16011_;
wire _16012_;
wire _16013_;
wire _16014_;
wire _16015_;
wire _16016_;
wire _16017_;
wire _16018_;
wire _16019_;
wire _16020_;
wire _16021_;
wire _16022_;
wire _16023_;
wire _16024_;
wire _16025_;
wire _16026_;
wire _16027_;
wire _16028_;
wire _16029_;
wire _16030_;
wire _16031_;
wire _16032_;
wire _16033_;
wire _16034_;
wire _16035_;
wire _16036_;
wire _16037_;
wire _16038_;
wire _16039_;
wire _16040_;
wire _16041_;
wire _16042_;
wire _16043_;
wire _16044_;
wire _16045_;
wire _16046_;
wire _16047_;
wire _16048_;
wire _16049_;
wire _16050_;
wire _16051_;
wire _16052_;
wire _16053_;
wire _16054_;
wire _16055_;
wire _16056_;
wire _16057_;
wire _16058_;
wire _16059_;
wire _16060_;
wire _16061_;
wire _16062_;
wire _16063_;
wire _16064_;
wire _16065_;
wire _16066_;
wire _16067_;
wire _16068_;
wire _16069_;
wire _16070_;
wire _16071_;
wire _16072_;
wire _16073_;
wire _16074_;
wire _16075_;
wire _16076_;
wire _16077_;
wire _16078_;
wire _16079_;
wire _16080_;
wire _16081_;
wire _16082_;
wire _16083_;
wire _16084_;
wire _16085_;
wire _16086_;
wire _16087_;
wire _16088_;
wire _16089_;
wire _16090_;
wire _16091_;
wire _16092_;
wire _16093_;
wire _16094_;
wire _16095_;
wire _16096_;
wire _16097_;
wire _16098_;
wire _16099_;
wire _16100_;
wire _16101_;
wire _16102_;
wire _16103_;
wire _16104_;
wire _16105_;
wire _16106_;
wire _16107_;
wire _16108_;
wire _16109_;
wire _16110_;
wire _16111_;
wire _16112_;
wire _16113_;
wire _16114_;
wire _16115_;
wire _16116_;
wire _16117_;
wire _16118_;
wire _16119_;
wire _16120_;
wire _16121_;
wire _16122_;
wire _16123_;
wire _16124_;
wire _16125_;
wire _16126_;
wire _16127_;
wire _16128_;
wire _16129_;
wire _16130_;
wire _16131_;
wire _16132_;
wire _16133_;
wire _16134_;
wire _16135_;
wire _16136_;
wire _16137_;
wire _16138_;
wire _16139_;
wire _16140_;
wire _16141_;
wire _16142_;
wire _16143_;
wire _16144_;
wire _16145_;
wire _16146_;
wire _16147_;
wire _16148_;
wire _16149_;
wire _16150_;
wire _16151_;
wire _16152_;
wire _16153_;
wire _16154_;
wire _16155_;
wire _16156_;
wire _16157_;
wire _16158_;
wire _16159_;
wire _16160_;
wire _16161_;
wire _16162_;
wire _16163_;
wire _16164_;
wire _16165_;
wire _16166_;
wire _16167_;
wire _16168_;
wire _16169_;
wire _16170_;
wire _16171_;
wire _16172_;
wire _16173_;
wire _16174_;
wire _16175_;
wire _16176_;
wire _16177_;
wire _16178_;
wire _16179_;
wire _16180_;
wire _16181_;
wire _16182_;
wire _16183_;
wire _16184_;
wire _16185_;
wire _16186_;
wire _16187_;
wire _16188_;
wire _16189_;
wire _16190_;
wire _16191_;
wire _16192_;
wire _16193_;
wire _16194_;
wire _16195_;
wire _16196_;
wire _16197_;
wire _16198_;
wire _16199_;
wire _16200_;
wire _16201_;
wire _16202_;
wire _16203_;
wire _16204_;
wire _16205_;
wire _16206_;
wire _16207_;
wire _16208_;
wire _16209_;
wire _16210_;
wire _16211_;
wire _16212_;
wire _16213_;
wire _16214_;
wire _16215_;
wire _16216_;
wire _16217_;
wire _16218_;
wire _16219_;
wire _16220_;
wire _16221_;
wire _16222_;
wire _16223_;
wire _16224_;
wire _16225_;
wire _16226_;
wire _16227_;
wire _16228_;
wire _16229_;
wire _16230_;
wire _16231_;
wire _16232_;
wire _16233_;
wire _16234_;
wire _16235_;
wire _16236_;
wire _16237_;
wire _16238_;
wire _16239_;
wire _16240_;
wire _16241_;
wire _16242_;
wire _16243_;
wire _16244_;
wire _16245_;
wire _16246_;
wire _16247_;
wire _16248_;
wire _16249_;
wire _16250_;
wire _16251_;
wire _16252_;
wire _16253_;
wire _16254_;
wire _16255_;
wire _16256_;
wire _16257_;
wire _16258_;
wire _16259_;
wire _16260_;
wire _16261_;
wire _16262_;
wire _16263_;
wire _16264_;
wire _16265_;
wire _16266_;
wire _16267_;
wire _16268_;
wire _16269_;
wire _16270_;
wire _16271_;
wire _16272_;
wire _16273_;
wire _16274_;
wire _16275_;
wire _16276_;
wire _16277_;
wire _16278_;
wire _16279_;
wire _16280_;
wire _16281_;
wire _16282_;
wire _16283_;
wire _16284_;
wire _16285_;
wire _16286_;
wire _16287_;
wire _16288_;
wire _16289_;
wire _16290_;
wire _16291_;
wire _16292_;
wire _16293_;
wire _16294_;
wire _16295_;
wire _16296_;
wire _16297_;
wire _16298_;
wire _16299_;
wire _16300_;
wire _16301_;
wire _16302_;
wire _16303_;
wire _16304_;
wire _16305_;
wire _16306_;
wire _16307_;
wire _16308_;
wire _16309_;
wire _16310_;
wire _16311_;
wire _16312_;
wire _16313_;
wire _16314_;
wire _16315_;
wire _16316_;
wire _16317_;
wire _16318_;
wire _16319_;
wire _16320_;
wire _16321_;
wire _16322_;
wire _16323_;
wire _16324_;
wire _16325_;
wire _16326_;
wire _16327_;
wire _16328_;
wire _16329_;
wire _16330_;
wire _16331_;
wire _16332_;
wire _16333_;
wire _16334_;
wire _16335_;
wire _16336_;
wire _16337_;
wire _16338_;
wire _16339_;
wire _16340_;
wire _16341_;
wire _16342_;
wire _16343_;
wire _16344_;
wire _16345_;
wire _16346_;
wire _16347_;
wire _16348_;
wire _16349_;
wire _16350_;
wire _16351_;
wire _16352_;
wire _16353_;
wire _16354_;
wire _16355_;
wire _16356_;
wire _16357_;
wire _16358_;
wire _16359_;
wire _16360_;
wire _16361_;
wire _16362_;
wire _16363_;
wire _16364_;
wire _16365_;
wire _16366_;
wire _16367_;
wire _16368_;
wire _16369_;
wire _16370_;
wire _16371_;
wire _16372_;
wire _16373_;
wire _16374_;
wire _16375_;
wire _16376_;
wire _16377_;
wire _16378_;
wire _16379_;
wire _16380_;
wire _16381_;
wire _16382_;
wire _16383_;
wire _16384_;
wire _16385_;
wire _16386_;
wire _16387_;
wire _16388_;
wire _16389_;
wire _16390_;
wire _16391_;
wire _16392_;
wire _16393_;
wire _16394_;
wire _16395_;
wire _16396_;
wire _16397_;
wire _16398_;
wire _16399_;
wire _16400_;
wire _16401_;
wire _16402_;
wire _16403_;
wire _16404_;
wire _16405_;
wire _16406_;
wire _16407_;
wire _16408_;
wire _16409_;
wire _16410_;
wire _16411_;
wire _16412_;
wire _16413_;
wire _16414_;
wire _16415_;
wire _16416_;
wire _16417_;
wire _16418_;
wire _16419_;
wire _16420_;
wire _16421_;
wire _16422_;
wire _16423_;
wire _16424_;
wire _16425_;
wire _16426_;
wire _16427_;
wire _16428_;
wire _16429_;
wire _16430_;
wire _16431_;
wire _16432_;
wire _16433_;
wire _16434_;
wire _16435_;
wire _16436_;
wire _16437_;
wire _16438_;
wire _16439_;
wire _16440_;
wire _16441_;
wire _16442_;
wire _16443_;
wire _16444_;
wire _16445_;
wire _16446_;
wire _16447_;
wire _16448_;
wire _16449_;
wire _16450_;
wire _16451_;
wire _16452_;
wire _16453_;
wire _16454_;
wire _16455_;
wire _16456_;
wire _16457_;
wire _16458_;
wire _16459_;
wire _16460_;
wire _16461_;
wire _16462_;
wire _16463_;
wire _16464_;
wire _16465_;
wire _16466_;
wire _16467_;
wire _16468_;
wire _16469_;
wire _16470_;
wire _16471_;
wire _16472_;
wire _16473_;
wire _16474_;
wire _16475_;
wire _16476_;
wire _16477_;
wire _16478_;
wire _16479_;
wire _16480_;
wire _16481_;
wire _16482_;
wire _16483_;
wire _16484_;
wire _16485_;
wire _16486_;
wire _16487_;
wire _16488_;
wire _16489_;
wire _16490_;
wire _16491_;
wire _16492_;
wire _16493_;
wire _16494_;
wire _16495_;
wire _16496_;
wire _16497_;
wire _16498_;
wire _16499_;
wire _16500_;
wire _16501_;
wire _16502_;
wire _16503_;
wire _16504_;
wire _16505_;
wire _16506_;
wire _16507_;
wire _16508_;
wire _16509_;
wire _16510_;
wire _16511_;
wire _16512_;
wire _16513_;
wire _16514_;
wire _16515_;
wire _16516_;
wire _16517_;
wire _16518_;
wire _16519_;
wire _16520_;
wire _16521_;
wire _16522_;
wire _16523_;
wire _16524_;
wire _16525_;
wire _16526_;
wire _16527_;
wire _16528_;
wire _16529_;
wire _16530_;
wire _16531_;
wire _16532_;
wire _16533_;
wire _16534_;
wire _16535_;
wire _16536_;
wire _16537_;
wire _16538_;
wire _16539_;
wire _16540_;
wire _16541_;
wire _16542_;
wire _16543_;
wire _16544_;
wire _16545_;
wire _16546_;
wire _16547_;
wire _16548_;
wire _16549_;
wire _16550_;
wire _16551_;
wire _16552_;
wire _16553_;
wire _16554_;
wire _16555_;
wire _16556_;
wire _16557_;
wire _16558_;
wire _16559_;
wire _16560_;
wire _16561_;
wire _16562_;
wire _16563_;
wire _16564_;
wire _16565_;
wire _16566_;
wire _16567_;
wire _16568_;
wire _16569_;
wire _16570_;
wire _16571_;
wire _16572_;
wire _16573_;
wire _16574_;
wire _16575_;
wire _16576_;
wire _16577_;
wire _16578_;
wire _16579_;
wire _16580_;
wire _16581_;
wire _16582_;
wire _16583_;
wire _16584_;
wire _16585_;
wire _16586_;
wire _16587_;
wire _16588_;
wire _16589_;
wire _16590_;
wire _16591_;
wire _16592_;
wire _16593_;
wire _16594_;
wire _16595_;
wire _16596_;
wire _16597_;
wire _16598_;
wire _16599_;
wire _16600_;
wire _16601_;
wire _16602_;
wire _16603_;
wire _16604_;
wire _16605_;
wire _16606_;
wire _16607_;
wire _16608_;
wire _16609_;
wire _16610_;
wire _16611_;
wire _16612_;
wire _16613_;
wire _16614_;
wire _16615_;
wire _16616_;
wire _16617_;
wire _16618_;
wire _16619_;
wire _16620_;
wire _16621_;
wire _16622_;
wire _16623_;
wire _16624_;
wire _16625_;
wire _16626_;
wire _16627_;
wire _16628_;
wire _16629_;
wire _16630_;
wire _16631_;
wire _16632_;
wire _16633_;
wire _16634_;
wire _16635_;
wire _16636_;
wire _16637_;
wire _16638_;
wire _16639_;
wire _16640_;
wire _16641_;
wire _16642_;
wire _16643_;
wire _16644_;
wire _16645_;
wire _16646_;
wire _16647_;
wire _16648_;
wire _16649_;
wire _16650_;
wire _16651_;
wire _16652_;
wire _16653_;
wire _16654_;
wire _16655_;
wire _16656_;
wire _16657_;
wire _16658_;
wire _16659_;
wire _16660_;
wire _16661_;
wire _16662_;
wire _16663_;
wire _16664_;
wire _16665_;
wire _16666_;
wire _16667_;
wire _16668_;
wire _16669_;
wire _16670_;
wire _16671_;
wire _16672_;
wire _16673_;
wire _16674_;
wire _16675_;
wire _16676_;
wire _16677_;
wire _16678_;
wire _16679_;
wire _16680_;
wire _16681_;
wire _16682_;
wire _16683_;
wire _16684_;
wire _16685_;
wire _16686_;
wire _16687_;
wire _16688_;
wire _16689_;
wire _16690_;
wire _16691_;
wire _16692_;
wire _16693_;
wire _16694_;
wire _16695_;
wire _16696_;
wire _16697_;
wire _16698_;
wire _16699_;
wire _16700_;
wire _16701_;
wire _16702_;
wire _16703_;
wire _16704_;
wire _16705_;
wire _16706_;
wire _16707_;
wire _16708_;
wire _16709_;
wire _16710_;
wire _16711_;
wire _16712_;
wire _16713_;
wire _16714_;
wire _16715_;
wire _16716_;
wire _16717_;
wire _16718_;
wire _16719_;
wire _16720_;
wire _16721_;
wire _16722_;
wire _16723_;
wire _16724_;
wire _16725_;
wire _16726_;
wire _16727_;
wire _16728_;
wire _16729_;
wire _16730_;
wire _16731_;
wire _16732_;
wire _16733_;
wire _16734_;
wire _16735_;
wire _16736_;
wire _16737_;
wire _16738_;
wire _16739_;
wire _16740_;
wire _16741_;
wire _16742_;
wire _16743_;
wire _16744_;
wire _16745_;
wire _16746_;
wire _16747_;
wire _16748_;
wire _16749_;
wire _16750_;
wire _16751_;
wire _16752_;
wire _16753_;
wire _16754_;
wire _16755_;
wire _16756_;
wire _16757_;
wire _16758_;
wire _16759_;
wire _16760_;
wire _16761_;
wire _16762_;
wire _16763_;
wire _16764_;
wire _16765_;
wire _16766_;
wire _16767_;
wire _16768_;
wire _16769_;
wire _16770_;
wire _16771_;
wire _16772_;
wire _16773_;
wire _16774_;
wire _16775_;
wire _16776_;
wire _16777_;
wire _16778_;
wire _16779_;
wire _16780_;
wire _16781_;
wire _16782_;
wire _16783_;
wire _16784_;
wire _16785_;
wire _16786_;
wire _16787_;
wire _16788_;
wire _16789_;
wire _16790_;
wire _16791_;
wire _16792_;
wire _16793_;
wire _16794_;
wire _16795_;
wire _16796_;
wire _16797_;
wire _16798_;
wire _16799_;
wire _16800_;
wire _16801_;
wire _16802_;
wire _16803_;
wire _16804_;
wire _16805_;
wire _16806_;
wire _16807_;
wire _16808_;
wire _16809_;
wire _16810_;
wire _16811_;
wire _16812_;
wire _16813_;
wire _16814_;
wire _16815_;
wire _16816_;
wire _16817_;
wire _16818_;
wire _16819_;
wire _16820_;
wire _16821_;
wire _16822_;
wire _16823_;
wire _16824_;
wire _16825_;
wire _16826_;
wire _16827_;
wire _16828_;
wire _16829_;
wire _16830_;
wire _16831_;
wire _16832_;
wire _16833_;
wire _16834_;
wire _16835_;
wire _16836_;
wire _16837_;
wire _16838_;
wire _16839_;
wire _16840_;
wire _16841_;
wire _16842_;
wire _16843_;
wire _16844_;
wire _16845_;
wire _16846_;
wire _16847_;
wire _16848_;
wire _16849_;
wire _16850_;
wire _16851_;
wire _16852_;
wire _16853_;
wire _16854_;
wire _16855_;
wire _16856_;
wire _16857_;
wire _16858_;
wire _16859_;
wire _16860_;
wire _16861_;
wire _16862_;
wire _16863_;
wire _16864_;
wire _16865_;
wire _16866_;
wire _16867_;
wire _16868_;
wire _16869_;
wire _16870_;
wire _16871_;
wire _16872_;
wire _16873_;
wire _16874_;
wire _16875_;
wire _16876_;
wire _16877_;
wire _16878_;
wire _16879_;
wire _16880_;
wire _16881_;
wire _16882_;
wire _16883_;
wire _16884_;
wire _16885_;
wire _16886_;
wire _16887_;
wire _16888_;
wire _16889_;
wire _16890_;
wire _16891_;
wire _16892_;
wire _16893_;
wire _16894_;
wire _16895_;
wire _16896_;
wire _16897_;
wire _16898_;
wire _16899_;
wire _16900_;
wire _16901_;
wire _16902_;
wire _16903_;
wire _16904_;
wire _16905_;
wire _16906_;
wire _16907_;
wire _16908_;
wire _16909_;
wire _16910_;
wire _16911_;
wire _16912_;
wire _16913_;
wire _16914_;
wire _16915_;
wire _16916_;
wire _16917_;
wire _16918_;
wire _16919_;
wire _16920_;
wire _16921_;
wire _16922_;
wire _16923_;
wire _16924_;
wire _16925_;
wire _16926_;
wire _16927_;
wire _16928_;
wire _16929_;
wire _16930_;
wire _16931_;
wire _16932_;
wire _16933_;
wire _16934_;
wire _16935_;
wire _16936_;
wire _16937_;
wire _16938_;
wire _16939_;
wire _16940_;
wire _16941_;
wire _16942_;
wire _16943_;
wire _16944_;
wire _16945_;
wire _16946_;
wire _16947_;
wire _16948_;
wire _16949_;
wire _16950_;
wire _16951_;
wire _16952_;
wire _16953_;
wire _16954_;
wire _16955_;
wire _16956_;
wire _16957_;
wire _16958_;
wire _16959_;
wire _16960_;
wire _16961_;
wire _16962_;
wire _16963_;
wire _16964_;
wire _16965_;
wire _16966_;
wire _16967_;
wire _16968_;
wire _16969_;
wire _16970_;
wire _16971_;
wire _16972_;
wire _16973_;
wire _16974_;
wire _16975_;
wire _16976_;
wire _16977_;
wire _16978_;
wire _16979_;
wire _16980_;
wire _16981_;
wire _16982_;
wire _16983_;
wire _16984_;
wire _16985_;
wire _16986_;
wire _16987_;
wire _16988_;
wire _16989_;
wire _16990_;
wire _16991_;
wire _16992_;
wire _16993_;
wire _16994_;
wire _16995_;
wire _16996_;
wire _16997_;
wire _16998_;
wire _16999_;
wire _17000_;
wire _17001_;
wire _17002_;
wire _17003_;
wire _17004_;
wire _17005_;
wire _17006_;
wire _17007_;
wire _17008_;
wire _17009_;
wire _17010_;
wire _17011_;
wire _17012_;
wire _17013_;
wire _17014_;
wire _17015_;
wire _17016_;
wire _17017_;
wire _17018_;
wire _17019_;
wire _17020_;
wire _17021_;
wire _17022_;
wire _17023_;
wire _17024_;
wire _17025_;
wire _17026_;
wire _17027_;
wire _17028_;
wire _17029_;
wire _17030_;
wire _17031_;
wire _17032_;
wire _17033_;
wire _17034_;
wire _17035_;
wire _17036_;
wire _17037_;
wire _17038_;
wire _17039_;
wire _17040_;
wire _17041_;
wire _17042_;
wire _17043_;
wire _17044_;
wire _17045_;
wire _17046_;
wire _17047_;
wire _17048_;
wire _17049_;
wire _17050_;
wire _17051_;
wire _17052_;
wire _17053_;
wire _17054_;
wire _17055_;
wire _17056_;
wire _17057_;
wire _17058_;
wire _17059_;
wire _17060_;
wire _17061_;
wire _17062_;
wire _17063_;
wire _17064_;
wire _17065_;
wire _17066_;
wire _17067_;
wire _17068_;
wire _17069_;
wire _17070_;
wire _17071_;
wire _17072_;
wire _17073_;
wire _17074_;
wire _17075_;
wire _17076_;
wire _17077_;
wire _17078_;
wire _17079_;
wire _17080_;
wire _17081_;
wire _17082_;
wire _17083_;
wire _17084_;
wire _17085_;
wire _17086_;
wire _17087_;
wire _17088_;
wire _17089_;
wire _17090_;
wire _17091_;
wire _17092_;
wire _17093_;
wire _17094_;
wire _17095_;
wire _17096_;
wire _17097_;
wire _17098_;
wire _17099_;
wire _17100_;
wire _17101_;
wire _17102_;
wire _17103_;
wire _17104_;
wire _17105_;
wire _17106_;
wire _17107_;
wire _17108_;
wire _17109_;
wire _17110_;
wire _17111_;
wire _17112_;
wire _17113_;
wire _17114_;
wire _17115_;
wire _17116_;
wire _17117_;
wire _17118_;
wire _17119_;
wire _17120_;
wire _17121_;
wire _17122_;
wire _17123_;
wire _17124_;
wire _17125_;
wire _17126_;
wire _17127_;
wire _17128_;
wire _17129_;
wire _17130_;
wire _17131_;
wire _17132_;
wire _17133_;
wire _17134_;
wire _17135_;
wire _17136_;
wire _17137_;
wire _17138_;
wire _17139_;
wire _17140_;
wire _17141_;
wire _17142_;
wire _17143_;
wire _17144_;
wire _17145_;
wire _17146_;
wire _17147_;
wire _17148_;
wire _17149_;
wire _17150_;
wire _17151_;
wire _17152_;
wire _17153_;
wire _17154_;
wire _17155_;
wire _17156_;
wire _17157_;
wire _17158_;
wire _17159_;
wire _17160_;
wire _17161_;
wire _17162_;
wire _17163_;
wire _17164_;
wire _17165_;
wire _17166_;
wire _17167_;
wire _17168_;
wire _17169_;
wire _17170_;
wire _17171_;
wire _17172_;
wire _17173_;
wire _17174_;
wire _17175_;
wire _17176_;
wire _17177_;
wire _17178_;
wire _17179_;
wire _17180_;
wire _17181_;
wire _17182_;
wire _17183_;
wire _17184_;
wire _17185_;
wire _17186_;
wire _17187_;
wire _17188_;
wire _17189_;
wire _17190_;
wire _17191_;
wire _17192_;
wire _17193_;
wire _17194_;
wire _17195_;
wire _17196_;
wire _17197_;
wire _17198_;
wire _17199_;
wire _17200_;
wire _17201_;
wire _17202_;
wire _17203_;
wire _17204_;
wire _17205_;
wire _17206_;
wire _17207_;
wire _17208_;
wire _17209_;
wire _17210_;
wire _17211_;
wire _17212_;
wire _17213_;
wire _17214_;
wire _17215_;
wire _17216_;
wire _17217_;
wire _17218_;
wire _17219_;
wire _17220_;
wire _17221_;
wire _17222_;
wire _17223_;
wire _17224_;
wire _17225_;
wire _17226_;
wire _17227_;
wire _17228_;
wire _17229_;
wire _17230_;
wire _17231_;
wire _17232_;
wire _17233_;
wire _17234_;
wire _17235_;
wire _17236_;
wire _17237_;
wire _17238_;
wire _17239_;
wire _17240_;
wire _17241_;
wire _17242_;
wire _17243_;
wire _17244_;
wire _17245_;
wire _17246_;
wire _17247_;
wire _17248_;
wire _17249_;
wire _17250_;
wire _17251_;
wire _17252_;
wire _17253_;
wire _17254_;
wire _17255_;
wire _17256_;
wire _17257_;
wire _17258_;
wire _17259_;
wire _17260_;
wire _17261_;
wire _17262_;
wire _17263_;
wire _17264_;
wire _17265_;
wire _17266_;
wire _17267_;
wire _17268_;
wire _17269_;
wire _17270_;
wire _17271_;
wire _17272_;
wire _17273_;
wire _17274_;
wire _17275_;
wire _17276_;
wire _17277_;
wire _17278_;
wire _17279_;
wire _17280_;
wire _17281_;
wire _17282_;
wire _17283_;
wire _17284_;
wire _17285_;
wire _17286_;
wire _17287_;
wire _17288_;
wire _17289_;
wire _17290_;
wire _17291_;
wire _17292_;
wire _17293_;
wire _17294_;
wire _17295_;
wire _17296_;
wire _17297_;
wire _17298_;
wire _17299_;
wire _17300_;
wire _17301_;
wire _17302_;
wire _17303_;
wire _17304_;
wire _17305_;
wire _17306_;
wire _17307_;
wire _17308_;
wire _17309_;
wire _17310_;
wire _17311_;
wire _17312_;
wire _17313_;
wire _17314_;
wire _17315_;
wire _17316_;
wire _17317_;
wire _17318_;
wire _17319_;
wire _17320_;
wire _17321_;
wire _17322_;
wire _17323_;
wire _17324_;
wire _17325_;
wire _17326_;
wire _17327_;
wire _17328_;
wire _17329_;
wire _17330_;
wire _17331_;
wire _17332_;
wire _17333_;
wire _17334_;
wire _17335_;
wire _17336_;
wire _17337_;
wire _17338_;
wire _17339_;
wire _17340_;
wire _17341_;
wire _17342_;
wire _17343_;
wire _17344_;
wire _17345_;
wire _17346_;
wire _17347_;
wire _17348_;
wire _17349_;
wire _17350_;
wire _17351_;
wire _17352_;
wire _17353_;
wire _17354_;
wire _17355_;
wire _17356_;
wire _17357_;
wire _17358_;
wire _17359_;
wire _17360_;
wire _17361_;
wire _17362_;
wire _17363_;
wire _17364_;
wire _17365_;
wire _17366_;
wire _17367_;
wire _17368_;
wire _17369_;
wire _17370_;
wire _17371_;
wire _17372_;
wire _17373_;
wire _17374_;
wire _17375_;
wire _17376_;
wire _17377_;
wire _17378_;
wire _17379_;
wire _17380_;
wire _17381_;
wire _17382_;
wire _17383_;
wire _17384_;
wire _17385_;
wire _17386_;
wire _17387_;
wire _17388_;
wire _17389_;
wire _17390_;
wire _17391_;
wire _17392_;
wire _17393_;
wire _17394_;
wire _17395_;
wire _17396_;
wire _17397_;
wire _17398_;
wire _17399_;
wire _17400_;
wire _17401_;
wire _17402_;
wire _17403_;
wire _17404_;
wire _17405_;
wire _17406_;
wire _17407_;
wire _17408_;
wire _17409_;
wire _17410_;
wire _17411_;
wire _17412_;
wire _17413_;
wire _17414_;
wire _17415_;
wire _17416_;
wire _17417_;
wire _17418_;
wire _17419_;
wire _17420_;
wire _17421_;
wire _17422_;
wire _17423_;
wire _17424_;
wire _17425_;
wire _17426_;
wire _17427_;
wire _17428_;
wire _17429_;
wire _17430_;
wire _17431_;
wire _17432_;
wire _17433_;
wire _17434_;
wire _17435_;
wire _17436_;
wire _17437_;
wire _17438_;
wire _17439_;
wire _17440_;
wire _17441_;
wire _17442_;
wire _17443_;
wire _17444_;
wire _17445_;
wire _17446_;
wire _17447_;
wire _17448_;
wire _17449_;
wire _17450_;
wire _17451_;
wire _17452_;
wire _17453_;
wire _17454_;
wire _17455_;
wire _17456_;
wire _17457_;
wire _17458_;
wire _17459_;
wire _17460_;
wire _17461_;
wire _17462_;
wire _17463_;
wire _17464_;
wire _17465_;
wire _17466_;
wire _17467_;
wire _17468_;
wire _17469_;
wire _17470_;
wire _17471_;
wire _17472_;
wire _17473_;
wire _17474_;
wire _17475_;
wire _17476_;
wire _17477_;
wire _17478_;
wire _17479_;
wire _17480_;
wire _17481_;
wire _17482_;
wire _17483_;
wire _17484_;
wire _17485_;
wire _17486_;
wire _17487_;
wire _17488_;
wire _17489_;
wire _17490_;
wire _17491_;
wire _17492_;
wire _17493_;
wire _17494_;
wire _17495_;
wire _17496_;
wire _17497_;
wire _17498_;
wire _17499_;
wire _17500_;
wire _17501_;
wire _17502_;
wire _17503_;
wire _17504_;
wire _17505_;
wire _17506_;
wire _17507_;
wire _17508_;
wire _17509_;
wire _17510_;
wire _17511_;
wire _17512_;
wire _17513_;
wire _17514_;
wire _17515_;
wire _17516_;
wire _17517_;
wire _17518_;
wire _17519_;
wire _17520_;
wire _17521_;
wire _17522_;
wire _17523_;
wire _17524_;
wire _17525_;
wire _17526_;
wire _17527_;
wire _17528_;
wire _17529_;
wire _17530_;
wire _17531_;
wire _17532_;
wire _17533_;
wire _17534_;
wire _17535_;
wire _17536_;
wire _17537_;
wire _17538_;
wire _17539_;
wire _17540_;
wire _17541_;
wire _17542_;
wire _17543_;
wire _17544_;
wire _17545_;
wire _17546_;
wire _17547_;
wire _17548_;
wire _17549_;
wire _17550_;
wire _17551_;
wire _17552_;
wire _17553_;
wire _17554_;
wire _17555_;
wire _17556_;
wire _17557_;
wire _17558_;
wire _17559_;
wire _17560_;
wire _17561_;
wire _17562_;
wire _17563_;
wire _17564_;
wire _17565_;
wire _17566_;
wire _17567_;
wire _17568_;
wire _17569_;
wire _17570_;
wire _17571_;
wire _17572_;
wire _17573_;
wire _17574_;
wire _17575_;
wire _17576_;
wire _17577_;
wire _17578_;
wire _17579_;
wire _17580_;
wire _17581_;
wire _17582_;
wire _17583_;
wire _17584_;
wire _17585_;
wire _17586_;
wire _17587_;
wire _17588_;
wire _17589_;
wire _17590_;
wire _17591_;
wire _17592_;
wire _17593_;
wire _17594_;
wire _17595_;
wire _17596_;
wire _17597_;
wire _17598_;
wire _17599_;
wire _17600_;
wire _17601_;
wire _17602_;
wire _17603_;
wire _17604_;
wire _17605_;
wire _17606_;
wire _17607_;
wire _17608_;
wire _17609_;
wire _17610_;
wire _17611_;
wire _17612_;
wire _17613_;
wire _17614_;
wire _17615_;
wire _17616_;
wire _17617_;
wire _17618_;
wire _17619_;
wire _17620_;
wire _17621_;
wire _17622_;
wire _17623_;
wire _17624_;
wire _17625_;
wire _17626_;
wire _17627_;
wire _17628_;
wire _17629_;
wire _17630_;
wire _17631_;
wire _17632_;
wire _17633_;
wire _17634_;
wire _17635_;
wire _17636_;
wire _17637_;
wire _17638_;
wire _17639_;
wire _17640_;
wire _17641_;
wire _17642_;
wire _17643_;
wire _17644_;
wire _17645_;
wire _17646_;
wire _17647_;
wire _17648_;
wire _17649_;
wire _17650_;
wire _17651_;
wire _17652_;
wire _17653_;
wire _17654_;
wire _17655_;
wire _17656_;
wire _17657_;
wire _17658_;
wire _17659_;
wire _17660_;
wire _17661_;
wire _17662_;
wire _17663_;
wire _17664_;
wire _17665_;
wire _17666_;
wire _17667_;
wire _17668_;
wire _17669_;
wire _17670_;
wire _17671_;
wire _17672_;
wire _17673_;
wire _17674_;
wire _17675_;
wire _17676_;
wire _17677_;
wire _17678_;
wire _17679_;
wire _17680_;
wire _17681_;
wire _17682_;
wire _17683_;
wire _17684_;
wire _17685_;
wire _17686_;
wire _17687_;
wire _17688_;
wire _17689_;
wire _17690_;
wire _17691_;
wire _17692_;
wire _17693_;
wire _17694_;
wire _17695_;
wire _17696_;
wire _17697_;
wire _17698_;
wire _17699_;
wire _17700_;
wire _17701_;
wire _17702_;
wire _17703_;
wire _17704_;
wire _17705_;
wire _17706_;
wire _17707_;
wire _17708_;
wire _17709_;
wire _17710_;
wire _17711_;
wire _17712_;
wire _17713_;
wire _17714_;
wire _17715_;
wire _17716_;
wire _17717_;
wire _17718_;
wire _17719_;
wire _17720_;
wire _17721_;
wire _17722_;
wire _17723_;
wire _17724_;
wire _17725_;
wire _17726_;
wire _17727_;
wire _17728_;
wire _17729_;
wire _17730_;
wire _17731_;
wire _17732_;
wire _17733_;
wire _17734_;
wire _17735_;
wire _17736_;
wire _17737_;
wire _17738_;
wire _17739_;
wire _17740_;
wire _17741_;
wire _17742_;
wire _17743_;
wire _17744_;
wire _17745_;
wire _17746_;
wire _17747_;
wire _17748_;
wire _17749_;
wire _17750_;
wire _17751_;
wire _17752_;
wire _17753_;
wire _17754_;
wire _17755_;
wire _17756_;
wire _17757_;
wire _17758_;
wire _17759_;
wire _17760_;
wire _17761_;
wire _17762_;
wire _17763_;
wire _17764_;
wire _17765_;
wire _17766_;
wire _17767_;
wire _17768_;
wire _17769_;
wire _17770_;
wire _17771_;
wire _17772_;
wire _17773_;
wire _17774_;
wire _17775_;
wire _17776_;
wire _17777_;
wire _17778_;
wire _17779_;
wire _17780_;
wire _17781_;
wire _17782_;
wire _17783_;
wire _17784_;
wire _17785_;
wire _17786_;
wire _17787_;
wire _17788_;
wire _17789_;
wire _17790_;
wire _17791_;
wire _17792_;
wire _17793_;
wire _17794_;
wire _17795_;
wire _17796_;
wire _17797_;
wire _17798_;
wire _17799_;
wire _17800_;
wire _17801_;
wire _17802_;
wire _17803_;
wire _17804_;
wire _17805_;
wire _17806_;
wire _17807_;
wire _17808_;
wire _17809_;
wire _17810_;
wire _17811_;
wire _17812_;
wire _17813_;
wire _17814_;
wire _17815_;
wire _17816_;
wire _17817_;
wire _17818_;
wire _17819_;
wire _17820_;
wire _17821_;
wire _17822_;
wire _17823_;
wire _17824_;
wire _17825_;
wire _17826_;
wire _17827_;
wire _17828_;
wire _17829_;
wire _17830_;
wire _17831_;
wire _17832_;
wire _17833_;
wire _17834_;
wire _17835_;
wire _17836_;
wire _17837_;
wire _17838_;
wire _17839_;
wire _17840_;
wire _17841_;
wire _17842_;
wire _17843_;
wire _17844_;
wire _17845_;
wire _17846_;
wire _17847_;
wire _17848_;
wire _17849_;
wire _17850_;
wire _17851_;
wire _17852_;
wire _17853_;
wire _17854_;
wire _17855_;
wire _17856_;
wire _17857_;
wire _17858_;
wire _17859_;
wire _17860_;
wire _17861_;
wire _17862_;
wire _17863_;
wire _17864_;
wire _17865_;
wire _17866_;
wire _17867_;
wire _17868_;
wire _17869_;
wire _17870_;
wire _17871_;
wire _17872_;
wire _17873_;
wire _17874_;
wire _17875_;
wire _17876_;
wire _17877_;
wire _17878_;
wire _17879_;
wire _17880_;
wire _17881_;
wire _17882_;
wire _17883_;
wire _17884_;
wire _17885_;
wire _17886_;
wire _17887_;
wire _17888_;
wire _17889_;
wire _17890_;
wire _17891_;
wire _17892_;
wire _17893_;
wire _17894_;
wire _17895_;
wire _17896_;
wire _17897_;
wire _17898_;
wire _17899_;
wire _17900_;
wire _17901_;
wire _17902_;
wire _17903_;
wire _17904_;
wire _17905_;
wire _17906_;
wire _17907_;
wire _17908_;
wire _17909_;
wire _17910_;
wire _17911_;
wire _17912_;
wire _17913_;
wire _17914_;
wire _17915_;
wire _17916_;
wire _17917_;
wire _17918_;
wire _17919_;
wire _17920_;
wire _17921_;
wire _17922_;
wire _17923_;
wire _17924_;
wire _17925_;
wire _17926_;
wire _17927_;
wire _17928_;
wire _17929_;
wire _17930_;
wire _17931_;
wire _17932_;
wire _17933_;
wire _17934_;
wire _17935_;
wire _17936_;
wire _17937_;
wire _17938_;
wire _17939_;
wire _17940_;
wire _17941_;
wire _17942_;
wire _17943_;
wire _17944_;
wire _17945_;
wire _17946_;
wire _17947_;
wire _17948_;
wire _17949_;
wire _17950_;
wire _17951_;
wire _17952_;
wire _17953_;
wire _17954_;
wire _17955_;
wire _17956_;
wire _17957_;
wire _17958_;
wire _17959_;
wire _17960_;
wire _17961_;
wire _17962_;
wire _17963_;
wire _17964_;
wire _17965_;
wire _17966_;
wire _17967_;
wire _17968_;
wire _17969_;
wire _17970_;
wire _17971_;
wire _17972_;
wire _17973_;
wire _17974_;
wire _17975_;
wire _17976_;
wire _17977_;
wire _17978_;
wire _17979_;
wire _17980_;
wire _17981_;
wire _17982_;
wire _17983_;
wire _17984_;
wire _17985_;
wire _17986_;
wire _17987_;
wire _17988_;
wire _17989_;
wire _17990_;
wire _17991_;
wire _17992_;
wire _17993_;
wire _17994_;
wire _17995_;
wire _17996_;
wire _17997_;
wire _17998_;
wire _17999_;
wire _18000_;
wire _18001_;
wire _18002_;
wire _18003_;
wire _18004_;
wire _18005_;
wire _18006_;
wire _18007_;
wire _18008_;
wire _18009_;
wire _18010_;
wire _18011_;
wire _18012_;
wire _18013_;
wire _18014_;
wire _18015_;
wire _18016_;
wire _18017_;
wire _18018_;
wire _18019_;
wire _18020_;
wire _18021_;
wire _18022_;
wire _18023_;
wire _18024_;
wire _18025_;
wire _18026_;
wire _18027_;
wire _18028_;
wire _18029_;
wire _18030_;
wire _18031_;
wire _18032_;
wire _18033_;
wire _18034_;
wire _18035_;
wire _18036_;
wire _18037_;
wire _18038_;
wire _18039_;
wire _18040_;
wire _18041_;
wire _18042_;
wire _18043_;
wire _18044_;
wire _18045_;
wire _18046_;
wire _18047_;
wire _18048_;
wire _18049_;
wire _18050_;
wire _18051_;
wire _18052_;
wire _18053_;
wire _18054_;
wire _18055_;
wire _18056_;
wire _18057_;
wire _18058_;
wire _18059_;
wire _18060_;
wire _18061_;
wire _18062_;
wire _18063_;
wire _18064_;
wire _18065_;
wire _18066_;
wire _18067_;
wire _18068_;
wire _18069_;
wire _18070_;
wire _18071_;
wire _18072_;
wire _18073_;
wire _18074_;
wire _18075_;
wire _18076_;
wire _18077_;
wire _18078_;
wire _18079_;
wire _18080_;
wire _18081_;
wire _18082_;
wire _18083_;
wire _18084_;
wire _18085_;
wire _18086_;
wire _18087_;
wire _18088_;
wire _18089_;
wire _18090_;
wire _18091_;
wire _18092_;
wire _18093_;
wire _18094_;
wire _18095_;
wire _18096_;
wire _18097_;
wire _18098_;
wire _18099_;
wire _18100_;
wire _18101_;
wire _18102_;
wire _18103_;
wire _18104_;
wire _18105_;
wire _18106_;
wire _18107_;
wire _18108_;
wire _18109_;
wire _18110_;
wire _18111_;
wire _18112_;
wire _18113_;
wire _18114_;
wire _18115_;
wire _18116_;
wire _18117_;
wire _18118_;
wire _18119_;
wire _18120_;
wire _18121_;
wire _18122_;
wire _18123_;
wire _18124_;
wire _18125_;
wire _18126_;
wire _18127_;
wire _18128_;
wire _18129_;
wire _18130_;
wire _18131_;
wire _18132_;
wire _18133_;
wire _18134_;
wire _18135_;
wire _18136_;
wire _18137_;
wire _18138_;
wire _18139_;
wire _18140_;
wire _18141_;
wire _18142_;
wire _18143_;
wire _18144_;
wire _18145_;
wire _18146_;
wire _18147_;
wire _18148_;
wire _18149_;
wire _18150_;
wire _18151_;
wire _18152_;
wire _18153_;
wire _18154_;
wire _18155_;
wire _18156_;
wire _18157_;
wire _18158_;
wire _18159_;
wire _18160_;
wire _18161_;
wire _18162_;
wire _18163_;
wire _18164_;
wire _18165_;
wire _18166_;
wire _18167_;
wire _18168_;
wire _18169_;
wire _18170_;
wire _18171_;
wire _18172_;
wire _18173_;
wire _18174_;
wire _18175_;
wire _18176_;
wire _18177_;
wire _18178_;
wire _18179_;
wire _18180_;
wire _18181_;
wire _18182_;
wire _18183_;
wire _18184_;
wire _18185_;
wire _18186_;
wire _18187_;
wire _18188_;
wire _18189_;
wire _18190_;
wire _18191_;
wire _18192_;
wire _18193_;
wire _18194_;
wire _18195_;
wire _18196_;
wire _18197_;
wire _18198_;
wire _18199_;
wire _18200_;
wire _18201_;
wire _18202_;
wire _18203_;
wire _18204_;
wire _18205_;
wire _18206_;
wire _18207_;
wire _18208_;
wire _18209_;
wire _18210_;
wire _18211_;
wire _18212_;
wire _18213_;
wire _18214_;
wire _18215_;
wire _18216_;
wire _18217_;
wire _18218_;
wire _18219_;
wire _18220_;
wire _18221_;
wire _18222_;
wire _18223_;
wire _18224_;
wire _18225_;
wire _18226_;
wire _18227_;
wire _18228_;
wire _18229_;
wire _18230_;
wire _18231_;
wire _18232_;
wire _18233_;
wire _18234_;
wire _18235_;
wire _18236_;
wire _18237_;
wire _18238_;
wire _18239_;
wire _18240_;
wire _18241_;
wire _18242_;
wire _18243_;
wire _18244_;
wire _18245_;
wire _18246_;
wire _18247_;
wire _18248_;
wire _18249_;
wire _18250_;
wire _18251_;
wire _18252_;
wire _18253_;
wire _18254_;
wire _18255_;
wire _18256_;
wire _18257_;
wire _18258_;
wire _18259_;
wire _18260_;
wire _18261_;
wire _18262_;
wire _18263_;
wire _18264_;
wire _18265_;
wire _18266_;
wire _18267_;
wire _18268_;
wire _18269_;
wire _18270_;
wire _18271_;
wire _18272_;
wire _18273_;
wire _18274_;
wire _18275_;
wire _18276_;
wire _18277_;
wire _18278_;
wire _18279_;
wire _18280_;
wire _18281_;
wire _18282_;
wire _18283_;
wire _18284_;
wire _18285_;
wire _18286_;
wire _18287_;
wire _18288_;
wire _18289_;
wire _18290_;
wire _18291_;
wire _18292_;
wire _18293_;
wire _18294_;
wire _18295_;
wire _18296_;
wire _18297_;
wire _18298_;
wire _18299_;
wire _18300_;
wire _18301_;
wire _18302_;
wire _18303_;
wire _18304_;
wire _18305_;
wire _18306_;
wire _18307_;
wire _18308_;
wire _18309_;
wire _18310_;
wire _18311_;
wire _18312_;
wire _18313_;
wire _18314_;
wire _18315_;
wire _18316_;
wire _18317_;
wire _18318_;
wire _18319_;
wire _18320_;
wire _18321_;
wire _18322_;
wire _18323_;
wire _18324_;
wire _18325_;
wire _18326_;
wire _18327_;
wire _18328_;
wire _18329_;
wire _18330_;
wire _18331_;
wire _18332_;
wire _18333_;
wire _18334_;
wire _18335_;
wire _18336_;
wire _18337_;
wire _18338_;
wire _18339_;
wire _18340_;
wire _18341_;
wire _18342_;
wire _18343_;
wire _18344_;
wire _18345_;
wire _18346_;
wire _18347_;
wire _18348_;
wire _18349_;
wire _18350_;
wire _18351_;
wire _18352_;
wire _18353_;
wire _18354_;
wire _18355_;
wire _18356_;
wire _18357_;
wire _18358_;
wire _18359_;
wire _18360_;
wire _18361_;
wire _18362_;
wire _18363_;
wire _18364_;
wire _18365_;
wire _18366_;
wire _18367_;
wire _18368_;
wire _18369_;
wire _18370_;
wire _18371_;
wire _18372_;
wire _18373_;
wire _18374_;
wire _18375_;
wire _18376_;
wire _18377_;
wire _18378_;
wire _18379_;
wire _18380_;
wire _18381_;
wire _18382_;
wire _18383_;
wire _18384_;
wire _18385_;
wire _18386_;
wire _18387_;
wire _18388_;
wire _18389_;
wire _18390_;
wire _18391_;
wire _18392_;
wire _18393_;
wire _18394_;
wire _18395_;
wire _18396_;
wire _18397_;
wire _18398_;
wire _18399_;
wire _18400_;
wire _18401_;
wire _18402_;
wire _18403_;
wire _18404_;
wire _18405_;
wire _18406_;
wire _18407_;
wire _18408_;
wire _18409_;
wire _18410_;
wire _18411_;
wire _18412_;
wire _18413_;
wire _18414_;
wire _18415_;
wire _18416_;
wire _18417_;
wire _18418_;
wire _18419_;
wire _18420_;
wire _18421_;
wire _18422_;
wire _18423_;
wire _18424_;
wire _18425_;
wire _18426_;
wire _18427_;
wire _18428_;
wire _18429_;
wire _18430_;
wire _18431_;
wire _18432_;
wire _18433_;
wire _18434_;
wire _18435_;
wire _18436_;
wire _18437_;
wire _18438_;
wire _18439_;
wire _18440_;
wire _18441_;
wire _18442_;
wire _18443_;
wire _18444_;
wire _18445_;
wire _18446_;
wire _18447_;
wire _18448_;
wire _18449_;
wire _18450_;
wire _18451_;
wire _18452_;
wire _18453_;
wire _18454_;
wire _18455_;
wire _18456_;
wire _18457_;
wire _18458_;
wire _18459_;
wire _18460_;
wire _18461_;
wire _18462_;
wire _18463_;
wire _18464_;
wire _18465_;
wire _18466_;
wire _18467_;
wire _18468_;
wire _18469_;
wire _18470_;
wire _18471_;
wire _18472_;
wire _18473_;
wire _18474_;
wire _18475_;
wire _18476_;
wire _18477_;
wire _18478_;
wire _18479_;
wire _18480_;
wire _18481_;
wire _18482_;
wire _18483_;
wire _18484_;
wire _18485_;
wire _18486_;
wire _18487_;
wire _18488_;
wire _18489_;
wire _18490_;
wire _18491_;
wire _18492_;
wire _18493_;
wire _18494_;
wire _18495_;
wire _18496_;
wire _18497_;
wire _18498_;
wire _18499_;
wire _18500_;
wire _18501_;
wire _18502_;
wire _18503_;
wire _18504_;
wire _18505_;
wire _18506_;
wire _18507_;
wire _18508_;
wire _18509_;
wire _18510_;
wire _18511_;
wire _18512_;
wire _18513_;
wire _18514_;
wire _18515_;
wire _18516_;
wire _18517_;
wire _18518_;
wire _18519_;
wire _18520_;
wire _18521_;
wire _18522_;
wire _18523_;
wire _18524_;
wire _18525_;
wire _18526_;
wire _18527_;
wire _18528_;
wire _18529_;
wire _18530_;
wire _18531_;
wire _18532_;
wire _18533_;
wire _18534_;
wire _18535_;
wire _18536_;
wire _18537_;
wire _18538_;
wire _18539_;
wire _18540_;
wire _18541_;
wire _18542_;
wire _18543_;
wire _18544_;
wire _18545_;
wire _18546_;
wire _18547_;
wire _18548_;
wire _18549_;
wire _18550_;
wire _18551_;
wire _18552_;
wire _18553_;
wire _18554_;
wire _18555_;
wire _18556_;
wire _18557_;
wire _18558_;
wire _18559_;
wire _18560_;
wire _18561_;
wire _18562_;
wire _18563_;
wire _18564_;
wire _18565_;
wire _18566_;
wire _18567_;
wire _18568_;
wire _18569_;
wire _18570_;
wire _18571_;
wire _18572_;
wire _18573_;
wire _18574_;
wire _18575_;
wire _18576_;
wire _18577_;
wire _18578_;
wire _18579_;
wire _18580_;
wire _18581_;
wire _18582_;
wire _18583_;
wire _18584_;
wire _18585_;
wire _18586_;
wire _18587_;
wire _18588_;
wire _18589_;
wire _18590_;
wire _18591_;
wire _18592_;
wire _18593_;
wire _18594_;
wire _18595_;
wire _18596_;
wire _18597_;
wire _18598_;
wire _18599_;
wire _18600_;
wire _18601_;
wire _18602_;
wire _18603_;
wire _18604_;
wire _18605_;
wire _18606_;
wire _18607_;
wire _18608_;
wire _18609_;
wire _18610_;
wire _18611_;
wire _18612_;
wire _18613_;
wire _18614_;
wire _18615_;
wire _18616_;
wire _18617_;
wire _18618_;
wire _18619_;
wire _18620_;
wire _18621_;
wire _18622_;
wire _18623_;
wire _18624_;
wire _18625_;
wire _18626_;
wire _18627_;
wire _18628_;
wire _18629_;
wire _18630_;
wire _18631_;
wire _18632_;
wire _18633_;
wire _18634_;
wire _18635_;
wire _18636_;
wire _18637_;
wire _18638_;
wire _18639_;
wire _18640_;
wire _18641_;
wire _18642_;
wire _18643_;
wire _18644_;
wire _18645_;
wire _18646_;
wire _18647_;
wire _18648_;
wire _18649_;
wire _18650_;
wire _18651_;
wire _18652_;
wire _18653_;
wire _18654_;
wire _18655_;
wire _18656_;
wire _18657_;
wire _18658_;
wire _18659_;
wire _18660_;
wire _18661_;
wire _18662_;
wire _18663_;
wire _18664_;
wire _18665_;
wire _18666_;
wire _18667_;
wire _18668_;
wire _18669_;
wire _18670_;
wire _18671_;
wire _18672_;
wire _18673_;
wire _18674_;
wire _18675_;
wire _18676_;
wire _18677_;
wire _18678_;
wire _18679_;
wire _18680_;
wire _18681_;
wire _18682_;
wire _18683_;
wire _18684_;
wire _18685_;
wire _18686_;
wire _18687_;
wire _18688_;
wire _18689_;
wire _18690_;
wire _18691_;
wire _18692_;
wire _18693_;
wire _18694_;
wire _18695_;
wire _18696_;
wire _18697_;
wire _18698_;
wire _18699_;
wire _18700_;
wire _18701_;
wire _18702_;
wire _18703_;
wire _18704_;
wire _18705_;
wire _18706_;
wire _18707_;
wire _18708_;
wire _18709_;
wire _18710_;
wire _18711_;
wire _18712_;
wire _18713_;
wire _18714_;
wire _18715_;
wire _18716_;
wire _18717_;
wire _18718_;
wire _18719_;
wire _18720_;
wire _18721_;
wire _18722_;
wire _18723_;
wire _18724_;
wire _18725_;
wire _18726_;
wire _18727_;
wire _18728_;
wire _18729_;
wire _18730_;
wire _18731_;
wire _18732_;
wire _18733_;
wire _18734_;
wire _18735_;
wire _18736_;
wire _18737_;
wire _18738_;
wire _18739_;
wire _18740_;
wire _18741_;
wire _18742_;
wire _18743_;
wire _18744_;
wire _18745_;
wire _18746_;
wire _18747_;
wire _18748_;
wire _18749_;
wire _18750_;
wire _18751_;
wire _18752_;
wire _18753_;
wire _18754_;
wire _18755_;
wire _18756_;
wire _18757_;
wire _18758_;
wire _18759_;
wire _18760_;
wire _18761_;
wire _18762_;
wire _18763_;
wire _18764_;
wire _18765_;
wire _18766_;
wire _18767_;
wire _18768_;
wire _18769_;
wire _18770_;
wire _18771_;
wire _18772_;
wire _18773_;
wire _18774_;
wire _18775_;
wire _18776_;
wire _18777_;
wire _18778_;
wire _18779_;
wire _18780_;
wire _18781_;
wire _18782_;
wire _18783_;
wire _18784_;
wire _18785_;
wire _18786_;
wire _18787_;
wire _18788_;
wire _18789_;
wire _18790_;
wire _18791_;
wire _18792_;
wire _18793_;
wire _18794_;
wire _18795_;
wire _18796_;
wire _18797_;
wire _18798_;
wire _18799_;
wire _18800_;
wire _18801_;
wire _18802_;
wire _18803_;
wire _18804_;
wire _18805_;
wire _18806_;
wire _18807_;
wire _18808_;
wire _18809_;
wire _18810_;
wire _18811_;
wire _18812_;
wire _18813_;
wire _18814_;
wire _18815_;
wire _18816_;
wire _18817_;
wire _18818_;
wire _18819_;
wire _18820_;
wire _18821_;
wire _18822_;
wire _18823_;
wire _18824_;
wire _18825_;
wire _18826_;
wire _18827_;
wire _18828_;
wire _18829_;
wire _18830_;
wire _18831_;
wire _18832_;
wire _18833_;
wire _18834_;
wire _18835_;
wire _18836_;
wire _18837_;
wire _18838_;
wire _18839_;
wire _18840_;
wire _18841_;
wire _18842_;
wire _18843_;
wire _18844_;
wire _18845_;
wire _18846_;
wire _18847_;
wire _18848_;
wire _18849_;
wire _18850_;
wire _18851_;
wire _18852_;
wire _18853_;
wire _18854_;
wire _18855_;
wire _18856_;
wire _18857_;
wire _18858_;
wire _18859_;
wire _18860_;
wire _18861_;
wire _18862_;
wire _18863_;
wire _18864_;
wire _18865_;
wire _18866_;
wire _18867_;
wire _18868_;
wire _18869_;
wire _18870_;
wire _18871_;
wire _18872_;
wire _18873_;
wire _18874_;
wire _18875_;
wire _18876_;
wire _18877_;
wire _18878_;
wire _18879_;
wire _18880_;
wire _18881_;
wire _18882_;
wire _18883_;
wire _18884_;
wire _18885_;
wire _18886_;
wire _18887_;
wire _18888_;
wire _18889_;
wire _18890_;
wire _18891_;
wire _18892_;
wire _18893_;
wire _18894_;
wire _18895_;
wire _18896_;
wire _18897_;
wire _18898_;
wire _18899_;
wire _18900_;
wire _18901_;
wire _18902_;
wire _18903_;
wire _18904_;
wire _18905_;
wire _18906_;
wire _18907_;
wire _18908_;
wire _18909_;
wire _18910_;
wire _18911_;
wire _18912_;
wire _18913_;
wire _18914_;
wire _18915_;
wire _18916_;
wire _18917_;
wire _18918_;
wire _18919_;
wire _18920_;
wire _18921_;
wire _18922_;
wire _18923_;
wire _18924_;
wire _18925_;
wire _18926_;
wire _18927_;
wire _18928_;
wire _18929_;
wire _18930_;
wire _18931_;
wire _18932_;
wire _18933_;
wire _18934_;
wire _18935_;
wire _18936_;
wire _18937_;
wire _18938_;
wire _18939_;
wire _18940_;
wire _18941_;
wire _18942_;
wire _18943_;
wire _18944_;
wire _18945_;
wire _18946_;
wire _18947_;
wire _18948_;
wire _18949_;
wire _18950_;
wire _18951_;
wire _18952_;
wire _18953_;
wire _18954_;
wire _18955_;
wire _18956_;
wire _18957_;
wire _18958_;
wire _18959_;
wire _18960_;
wire _18961_;
wire _18962_;
wire _18963_;
wire _18964_;
wire _18965_;
wire _18966_;
wire _18967_;
wire _18968_;
wire _18969_;
wire _18970_;
wire _18971_;
wire _18972_;
wire _18973_;
wire _18974_;
wire _18975_;
wire _18976_;
wire _18977_;
wire _18978_;
wire _18979_;
wire _18980_;
wire _18981_;
wire _18982_;
wire _18983_;
wire _18984_;
wire _18985_;
wire _18986_;
wire _18987_;
wire _18988_;
wire _18989_;
wire _18990_;
wire _18991_;
wire _18992_;
wire _18993_;
wire _18994_;
wire _18995_;
wire _18996_;
wire _18997_;
wire _18998_;
wire _18999_;
wire _19000_;
wire _19001_;
wire _19002_;
wire _19003_;
wire _19004_;
wire _19005_;
wire _19006_;
wire _19007_;
wire _19008_;
wire _19009_;
wire _19010_;
wire _19011_;
wire _19012_;
wire _19013_;
wire _19014_;
wire _19015_;
wire _19016_;
wire _19017_;
wire _19018_;
wire _19019_;
wire _19020_;
wire _19021_;
wire _19022_;
wire _19023_;
wire _19024_;
wire _19025_;
wire _19026_;
wire _19027_;
wire _19028_;
wire _19029_;
wire _19030_;
wire _19031_;
wire _19032_;
wire _19033_;
wire _19034_;
wire _19035_;
wire _19036_;
wire _19037_;
wire _19038_;
wire _19039_;
wire _19040_;
wire _19041_;
wire _19042_;
wire _19043_;
wire _19044_;
wire _19045_;
wire _19046_;
wire _19047_;
wire _19048_;
wire _19049_;
wire _19050_;
wire _19051_;
wire _19052_;
wire _19053_;
wire _19054_;
wire _19055_;
wire _19056_;
wire _19057_;
wire _19058_;
wire _19059_;
wire _19060_;
wire _19061_;
wire _19062_;
wire _19063_;
wire _19064_;
wire _19065_;
wire _19066_;
wire _19067_;
wire _19068_;
wire _19069_;
wire _19070_;
wire _19071_;
wire _19072_;
wire _19073_;
wire _19074_;
wire _19075_;
wire _19076_;
wire _19077_;
wire _19078_;
wire _19079_;
wire _19080_;
wire _19081_;
wire _19082_;
wire _19083_;
wire _19084_;
wire _19085_;
wire _19086_;
wire _19087_;
wire _19088_;
wire _19089_;
wire _19090_;
wire _19091_;
wire _19092_;
wire _19093_;
wire _19094_;
wire _19095_;
wire _19096_;
wire _19097_;
wire _19098_;
wire _19099_;
wire _19100_;
wire _19101_;
wire _19102_;
wire _19103_;
wire _19104_;
wire _19105_;
wire _19106_;
wire _19107_;
wire _19108_;
wire _19109_;
wire _19110_;
wire _19111_;
wire _19112_;
wire _19113_;
wire _19114_;
wire _19115_;
wire _19116_;
wire _19117_;
wire _19118_;
wire _19119_;
wire _19120_;
wire _19121_;
wire _19122_;
wire _19123_;
wire _19124_;
wire _19125_;
wire _19126_;
wire _19127_;
wire _19128_;
wire _19129_;
wire _19130_;
wire _19131_;
wire _19132_;
wire _19133_;
wire _19134_;
wire _19135_;
wire _19136_;
wire _19137_;
wire _19138_;
wire _19139_;
wire _19140_;
wire _19141_;
wire _19142_;
wire _19143_;
wire _19144_;
wire _19145_;
wire _19146_;
wire _19147_;
wire _19148_;
wire _19149_;
wire _19150_;
wire _19151_;
wire _19152_;
wire _19153_;
wire _19154_;
wire _19155_;
wire _19156_;
wire _19157_;
wire _19158_;
wire _19159_;
wire _19160_;
wire _19161_;
wire _19162_;
wire _19163_;
wire _19164_;
wire _19165_;
wire _19166_;
wire _19167_;
wire _19168_;
wire _19169_;
wire _19170_;
wire _19171_;
wire _19172_;
wire _19173_;
wire _19174_;
wire _19175_;
wire _19176_;
wire _19177_;
wire _19178_;
wire _19179_;
wire _19180_;
wire _19181_;
wire _19182_;
wire _19183_;
wire _19184_;
wire _19185_;
wire _19186_;
wire _19187_;
wire _19188_;
wire _19189_;
wire _19190_;
wire _19191_;
wire _19192_;
wire _19193_;
wire _19194_;
wire _19195_;
wire _19196_;
wire _19197_;
wire _19198_;
wire _19199_;
wire _19200_;
wire _19201_;
wire _19202_;
wire _19203_;
wire _19204_;
wire _19205_;
wire _19206_;
wire _19207_;
wire _19208_;
wire _19209_;
wire _19210_;
wire _19211_;
wire _19212_;
wire _19213_;
wire _19214_;
wire _19215_;
wire _19216_;
wire _19217_;
wire _19218_;
wire _19219_;
wire _19220_;
wire _19221_;
wire _19222_;
wire _19223_;
wire _19224_;
wire _19225_;
wire _19226_;
wire _19227_;
wire _19228_;
wire _19229_;
wire _19230_;
wire _19231_;
wire _19232_;
wire _19233_;
wire _19234_;
wire _19235_;
wire _19236_;
wire _19237_;
wire _19238_;
wire _19239_;
wire _19240_;
wire _19241_;
wire _19242_;
wire _19243_;
wire _19244_;
wire _19245_;
wire _19246_;
wire _19247_;
wire _19248_;
wire _19249_;
wire _19250_;
wire _19251_;
wire _19252_;
wire _19253_;
wire _19254_;
wire _19255_;
wire _19256_;
wire _19257_;
wire _19258_;
wire _19259_;
wire _19260_;
wire _19261_;
wire _19262_;
wire _19263_;
wire _19264_;
wire _19265_;
wire _19266_;
wire _19267_;
wire _19268_;
wire _19269_;
wire _19270_;
wire _19271_;
wire _19272_;
wire _19273_;
wire _19274_;
wire _19275_;
wire _19276_;
wire _19277_;
wire _19278_;
wire _19279_;
wire _19280_;
wire _19281_;
wire _19282_;
wire _19283_;
wire _19284_;
wire _19285_;
wire _19286_;
wire _19287_;
wire _19288_;
wire _19289_;
wire _19290_;
wire _19291_;
wire _19292_;
wire _19293_;
wire _19294_;
wire _19295_;
wire _19296_;
wire _19297_;
wire _19298_;
wire _19299_;
wire _19300_;
wire _19301_;
wire _19302_;
wire _19303_;
wire _19304_;
wire _19305_;
wire _19306_;
wire _19307_;
wire _19308_;
wire _19309_;
wire _19310_;
wire _19311_;
wire _19312_;
wire _19313_;
wire _19314_;
wire _19315_;
wire _19316_;
wire _19317_;
wire _19318_;
wire _19319_;
wire _19320_;
wire _19321_;
wire _19322_;
wire _19323_;
wire _19324_;
wire _19325_;
wire _19326_;
wire _19327_;
wire _19328_;
wire _19329_;
wire _19330_;
wire _19331_;
wire _19332_;
wire _19333_;
wire _19334_;
wire _19335_;
wire _19336_;
wire _19337_;
wire _19338_;
wire _19339_;
wire _19340_;
wire _19341_;
wire _19342_;
wire _19343_;
wire _19344_;
wire _19345_;
wire _19346_;
wire _19347_;
wire _19348_;
wire _19349_;
wire _19350_;
wire _19351_;
wire _19352_;
wire _19353_;
wire _19354_;
wire _19355_;
wire _19356_;
wire _19357_;
wire _19358_;
wire _19359_;
wire _19360_;
wire _19361_;
wire _19362_;
wire _19363_;
wire _19364_;
wire _19365_;
wire _19366_;
wire _19367_;
wire _19368_;
wire _19369_;
wire _19370_;
wire _19371_;
wire _19372_;
wire _19373_;
wire _19374_;
wire _19375_;
wire _19376_;
wire _19377_;
wire _19378_;
wire _19379_;
wire _19380_;
wire _19381_;
wire _19382_;
wire _19383_;
wire _19384_;
wire _19385_;
wire _19386_;
wire _19387_;
wire _19388_;
wire _19389_;
wire _19390_;
wire _19391_;
wire _19392_;
wire _19393_;
wire _19394_;
wire _19395_;
wire _19396_;
wire _19397_;
wire _19398_;
wire _19399_;
wire _19400_;
wire _19401_;
wire _19402_;
wire _19403_;
wire _19404_;
wire _19405_;
wire _19406_;
wire _19407_;
wire _19408_;
wire _19409_;
wire _19410_;
wire _19411_;
wire _19412_;
wire _19413_;
wire _19414_;
wire _19415_;
wire _19416_;
wire _19417_;
wire _19418_;
wire _19419_;
wire _19420_;
wire _19421_;
wire _19422_;
wire _19423_;
wire _19424_;
wire _19425_;
wire _19426_;
wire _19427_;
wire _19428_;
wire _19429_;
wire _19430_;
wire _19431_;
wire _19432_;
wire _19433_;
wire _19434_;
wire _19435_;
wire _19436_;
wire _19437_;
wire _19438_;
wire _19439_;
wire _19440_;
wire _19441_;
wire _19442_;
wire _19443_;
wire _19444_;
wire _19445_;
wire _19446_;
wire _19447_;
wire _19448_;
wire _19449_;
wire _19450_;
wire _19451_;
wire _19452_;
wire _19453_;
wire _19454_;
wire _19455_;
wire _19456_;
wire _19457_;
wire _19458_;
wire _19459_;
wire _19460_;
wire _19461_;
wire _19462_;
wire _19463_;
wire _19464_;
wire _19465_;
wire _19466_;
wire _19467_;
wire _19468_;
wire _19469_;
wire _19470_;
wire _19471_;
wire _19472_;
wire _19473_;
wire _19474_;
wire _19475_;
wire _19476_;
wire _19477_;
wire _19478_;
wire _19479_;
wire _19480_;
wire _19481_;
wire _19482_;
wire _19483_;
wire _19484_;
wire _19485_;
wire _19486_;
wire _19487_;
wire _19488_;
wire _19489_;
wire _19490_;
wire _19491_;
wire _19492_;
wire _19493_;
wire _19494_;
wire _19495_;
wire _19496_;
wire _19497_;
wire _19498_;
wire _19499_;
wire _19500_;
wire _19501_;
wire _19502_;
wire _19503_;
wire _19504_;
wire _19505_;
wire _19506_;
wire _19507_;
wire _19508_;
wire _19509_;
wire _19510_;
wire _19511_;
wire _19512_;
wire _19513_;
wire _19514_;
wire _19515_;
wire _19516_;
wire _19517_;
wire _19518_;
wire _19519_;
wire _19520_;
wire _19521_;
wire _19522_;
wire _19523_;
wire _19524_;
wire _19525_;
wire _19526_;
wire _19527_;
wire _19528_;
wire _19529_;
wire _19530_;
wire _19531_;
wire _19532_;
wire _19533_;
wire _19534_;
wire _19535_;
wire _19536_;
wire _19537_;
wire _19538_;
wire _19539_;
wire _19540_;
wire _19541_;
wire _19542_;
wire _19543_;
wire _19544_;
wire _19545_;
wire _19546_;
wire _19547_;
wire _19548_;
wire _19549_;
wire _19550_;
wire _19551_;
wire _19552_;
wire _19553_;
wire _19554_;
wire _19555_;
wire _19556_;
wire _19557_;
wire _19558_;
wire _19559_;
wire _19560_;
wire _19561_;
wire _19562_;
wire _19563_;
wire _19564_;
wire _19565_;
wire _19566_;
wire _19567_;
wire _19568_;
wire _19569_;
wire _19570_;
wire _19571_;
wire _19572_;
wire _19573_;
wire _19574_;
wire _19575_;
wire _19576_;
wire _19577_;
wire _19578_;
wire _19579_;
wire _19580_;
wire _19581_;
wire _19582_;
wire _19583_;
wire _19584_;
wire _19585_;
wire _19586_;
wire _19587_;
wire _19588_;
wire _19589_;
wire _19590_;
wire _19591_;
wire _19592_;
wire _19593_;
wire _19594_;
wire _19595_;
wire _19596_;
wire _19597_;
wire _19598_;
wire _19599_;
wire _19600_;
wire _19601_;
wire _19602_;
wire _19603_;
wire _19604_;
wire _19605_;
wire _19606_;
wire _19607_;
wire _19608_;
wire _19609_;
wire _19610_;
wire _19611_;
wire _19612_;
wire _19613_;
wire _19614_;
wire _19615_;
wire _19616_;
wire _19617_;
wire _19618_;
wire _19619_;
wire _19620_;
wire _19621_;
wire _19622_;
wire _19623_;
wire _19624_;
wire _19625_;
wire _19626_;
wire _19627_;
wire _19628_;
wire _19629_;
wire _19630_;
wire _19631_;
wire _19632_;
wire _19633_;
wire _19634_;
wire _19635_;
wire _19636_;
wire _19637_;
wire _19638_;
wire _19639_;
wire _19640_;
wire _19641_;
wire _19642_;
wire _19643_;
wire _19644_;
wire _19645_;
wire _19646_;
wire _19647_;
wire _19648_;
wire _19649_;
wire _19650_;
wire _19651_;
wire _19652_;
wire _19653_;
wire _19654_;
wire _19655_;
wire _19656_;
wire _19657_;
wire _19658_;
wire _19659_;
wire _19660_;
wire _19661_;
wire _19662_;
wire _19663_;
wire _19664_;
wire _19665_;
wire _19666_;
wire _19667_;
wire _19668_;
wire _19669_;
wire _19670_;
wire _19671_;
wire _19672_;
wire _19673_;
wire _19674_;
wire _19675_;
wire _19676_;
wire _19677_;
wire _19678_;
wire _19679_;
wire _19680_;
wire _19681_;
wire _19682_;
wire _19683_;
wire _19684_;
wire _19685_;
wire _19686_;
wire _19687_;
wire _19688_;
wire _19689_;
wire _19690_;
wire _19691_;
wire _19692_;
wire _19693_;
wire _19694_;
wire _19695_;
wire _19696_;
wire _19697_;
wire _19698_;
wire _19699_;
wire _19700_;
wire _19701_;
wire _19702_;
wire _19703_;
wire _19704_;
wire _19705_;
wire _19706_;
wire _19707_;
wire _19708_;
wire _19709_;
wire _19710_;
wire _19711_;
wire _19712_;
wire _19713_;
wire _19714_;
wire _19715_;
wire _19716_;
wire _19717_;
wire _19718_;
wire _19719_;
wire _19720_;
wire _19721_;
wire _19722_;
wire _19723_;
wire _19724_;
wire _19725_;
wire _19726_;
wire _19727_;
wire _19728_;
wire _19729_;
wire _19730_;
wire _19731_;
wire _19732_;
wire _19733_;
wire _19734_;
wire _19735_;
wire _19736_;
wire _19737_;
wire _19738_;
wire _19739_;
wire _19740_;
wire _19741_;
wire _19742_;
wire _19743_;
wire _19744_;
wire _19745_;
wire _19746_;
wire _19747_;
wire _19748_;
wire _19749_;
wire _19750_;
wire _19751_;
wire _19752_;
wire _19753_;
wire _19754_;
wire _19755_;
wire _19756_;
wire _19757_;
wire _19758_;
wire _19759_;
wire _19760_;
wire _19761_;
wire _19762_;
wire _19763_;
wire _19764_;
wire _19765_;
wire _19766_;
wire _19767_;
wire _19768_;
wire _19769_;
wire _19770_;
wire _19771_;
wire _19772_;
wire _19773_;
wire _19774_;
wire _19775_;
wire _19776_;
wire _19777_;
wire _19778_;
wire _19779_;
wire _19780_;
wire _19781_;
wire _19782_;
wire _19783_;
wire _19784_;
wire _19785_;
wire _19786_;
wire _19787_;
wire _19788_;
wire _19789_;
wire _19790_;
wire _19791_;
wire _19792_;
wire _19793_;
wire _19794_;
wire _19795_;
wire _19796_;
wire _19797_;
wire _19798_;
wire _19799_;
wire _19800_;
wire _19801_;
wire _19802_;
wire _19803_;
wire _19804_;
wire _19805_;
wire _19806_;
wire _19807_;
wire _19808_;
wire _19809_;
wire _19810_;
wire _19811_;
wire _19812_;
wire _19813_;
wire _19814_;
wire _19815_;
wire _19816_;
wire _19817_;
wire _19818_;
wire _19819_;
wire _19820_;
wire _19821_;
wire _19822_;
wire _19823_;
wire _19824_;
wire _19825_;
wire _19826_;
wire _19827_;
wire _19828_;
wire _19829_;
wire _19830_;
wire _19831_;
wire _19832_;
wire _19833_;
wire _19834_;
wire _19835_;
wire _19836_;
wire _19837_;
wire _19838_;
wire _19839_;
wire _19840_;
wire _19841_;
wire _19842_;
wire _19843_;
wire _19844_;
wire _19845_;
wire _19846_;
wire _19847_;
wire _19848_;
wire _19849_;
wire _19850_;
wire _19851_;
wire _19852_;
wire _19853_;
wire _19854_;
wire _19855_;
wire _19856_;
wire _19857_;
wire _19858_;
wire _19859_;
wire _19860_;
wire _19861_;
wire _19862_;
wire _19863_;
wire _19864_;
wire _19865_;
wire _19866_;
wire _19867_;
wire _19868_;
wire _19869_;
wire _19870_;
wire _19871_;
wire _19872_;
wire _19873_;
wire _19874_;
wire _19875_;
wire _19876_;
wire _19877_;
wire _19878_;
wire _19879_;
wire _19880_;
wire _19881_;
wire _19882_;
wire _19883_;
wire _19884_;
wire _19885_;
wire _19886_;
wire _19887_;
wire _19888_;
wire _19889_;
wire _19890_;
wire _19891_;
wire _19892_;
wire _19893_;
wire _19894_;
wire _19895_;
wire _19896_;
wire _19897_;
wire _19898_;
wire _19899_;
wire _19900_;
wire _19901_;
wire _19902_;
wire _19903_;
wire _19904_;
wire _19905_;
wire _19906_;
wire _19907_;
wire _19908_;
wire _19909_;
wire _19910_;
wire _19911_;
wire _19912_;
wire _19913_;
wire _19914_;
wire _19915_;
wire _19916_;
wire _19917_;
wire _19918_;
wire _19919_;
wire _19920_;
wire _19921_;
wire _19922_;
wire _19923_;
wire _19924_;
wire _19925_;
wire _19926_;
wire _19927_;
wire _19928_;
wire _19929_;
wire _19930_;
wire _19931_;
wire _19932_;
wire _19933_;
wire _19934_;
wire _19935_;
wire _19936_;
wire _19937_;
wire _19938_;
wire _19939_;
wire _19940_;
wire _19941_;
wire _19942_;
wire _19943_;
wire _19944_;
wire _19945_;
wire _19946_;
wire _19947_;
wire _19948_;
wire _19949_;
wire _19950_;
wire _19951_;
wire _19952_;
wire _19953_;
wire _19954_;
wire _19955_;
wire _19956_;
wire _19957_;
wire _19958_;
wire _19959_;
wire _19960_;
wire _19961_;
wire _19962_;
wire _19963_;
wire _19964_;
wire _19965_;
wire _19966_;
wire _19967_;
wire _19968_;
wire _19969_;
wire _19970_;
wire _19971_;
wire _19972_;
wire _19973_;
wire _19974_;
wire _19975_;
wire _19976_;
wire _19977_;
wire _19978_;
wire _19979_;
wire _19980_;
wire _19981_;
wire _19982_;
wire _19983_;
wire _19984_;
wire _19985_;
wire _19986_;
wire _19987_;
wire _19988_;
wire _19989_;
wire _19990_;
wire _19991_;
wire _19992_;
wire _19993_;
wire _19994_;
wire _19995_;
wire _19996_;
wire _19997_;
wire _19998_;
wire _19999_;
wire _20000_;
wire _20001_;
wire _20002_;
wire _20003_;
wire _20004_;
wire _20005_;
wire _20006_;
wire _20007_;
wire _20008_;
wire _20009_;
wire _20010_;
wire _20011_;
wire _20012_;
wire _20013_;
wire _20014_;
wire _20015_;
wire _20016_;
wire _20017_;
wire _20018_;
wire _20019_;
wire _20020_;
wire _20021_;
wire _20022_;
wire _20023_;
wire _20024_;
wire _20025_;
wire _20026_;
wire _20027_;
wire _20028_;
wire _20029_;
wire _20030_;
wire _20031_;
wire _20032_;
wire _20033_;
wire _20034_;
wire _20035_;
wire _20036_;
wire _20037_;
wire _20038_;
wire _20039_;
wire _20040_;
wire _20041_;
wire _20042_;
wire _20043_;
wire _20044_;
wire _20045_;
wire _20046_;
wire _20047_;
wire _20048_;
wire _20049_;
wire _20050_;
wire _20051_;
wire _20052_;
wire _20053_;
wire _20054_;
wire _20055_;
wire _20056_;
wire _20057_;
wire _20058_;
wire _20059_;
wire _20060_;
wire _20061_;
wire _20062_;
wire _20063_;
wire _20064_;
wire _20065_;
wire _20066_;
wire _20067_;
wire _20068_;
wire _20069_;
wire _20070_;
wire _20071_;
wire _20072_;
wire _20073_;
wire _20074_;
wire _20075_;
wire _20076_;
wire _20077_;
wire _20078_;
wire _20079_;
wire _20080_;
wire _20081_;
wire _20082_;
wire _20083_;
wire _20084_;
wire _20085_;
wire _20086_;
wire _20087_;
wire _20088_;
wire _20089_;
wire _20090_;
wire _20091_;
wire _20092_;
wire _20093_;
wire _20094_;
wire _20095_;
wire _20096_;
wire _20097_;
wire _20098_;
wire _20099_;
wire _20100_;
wire _20101_;
wire _20102_;
wire _20103_;
wire _20104_;
wire _20105_;
wire _20106_;
wire _20107_;
wire _20108_;
wire _20109_;
wire _20110_;
wire _20111_;
wire _20112_;
wire _20113_;
wire _20114_;
wire _20115_;
wire _20116_;
wire _20117_;
wire _20118_;
wire _20119_;
wire _20120_;
wire _20121_;
wire _20122_;
wire _20123_;
wire _20124_;
wire _20125_;
wire _20126_;
wire _20127_;
wire _20128_;
wire _20129_;
wire _20130_;
wire _20131_;
wire _20132_;
wire _20133_;
wire _20134_;
wire _20135_;
wire _20136_;
wire _20137_;
wire _20138_;
wire _20139_;
wire _20140_;
wire _20141_;
wire _20142_;
wire _20143_;
wire _20144_;
wire _20145_;
wire _20146_;
wire _20147_;
wire _20148_;
wire _20149_;
wire _20150_;
wire _20151_;
wire _20152_;
wire _20153_;
wire _20154_;
wire _20155_;
wire _20156_;
wire _20157_;
wire _20158_;
wire _20159_;
wire _20160_;
wire _20161_;
wire _20162_;
wire _20163_;
wire _20164_;
wire _20165_;
wire _20166_;
wire _20167_;
wire _20168_;
wire _20169_;
wire _20170_;
wire _20171_;
wire _20172_;
wire _20173_;
wire _20174_;
wire _20175_;
wire _20176_;
wire _20177_;
wire _20178_;
wire _20179_;
wire _20180_;
wire _20181_;
wire _20182_;
wire _20183_;
wire _20184_;
wire _20185_;
wire _20186_;
wire _20187_;
wire _20188_;
wire _20189_;
wire _20190_;
wire _20191_;
wire _20192_;
wire _20193_;
wire _20194_;
wire _20195_;
wire _20196_;
wire _20197_;
wire _20198_;
wire _20199_;
wire _20200_;
wire _20201_;
wire _20202_;
wire _20203_;
wire _20204_;
wire _20205_;
wire _20206_;
wire _20207_;
wire _20208_;
wire _20209_;
wire _20210_;
wire _20211_;
wire _20212_;
wire _20213_;
wire _20214_;
wire _20215_;
wire _20216_;
wire _20217_;
wire _20218_;
wire _20219_;
wire _20220_;
wire _20221_;
wire _20222_;
wire _20223_;
wire _20224_;
wire _20225_;
wire _20226_;
wire _20227_;
wire _20228_;
wire _20229_;
wire _20230_;
wire _20231_;
wire _20232_;
wire _20233_;
wire _20234_;
wire _20235_;
wire _20236_;
wire _20237_;
wire _20238_;
wire _20239_;
wire _20240_;
wire _20241_;
wire _20242_;
wire _20243_;
wire _20244_;
wire _20245_;
wire _20246_;
wire _20247_;
wire _20248_;
wire _20249_;
wire _20250_;
wire _20251_;
wire _20252_;
wire _20253_;
wire _20254_;
wire _20255_;
wire _20256_;
wire _20257_;
wire _20258_;
wire _20259_;
wire _20260_;
wire _20261_;
wire _20262_;
wire _20263_;
wire _20264_;
wire _20265_;
wire _20266_;
wire _20267_;
wire _20268_;
wire _20269_;
wire _20270_;
wire _20271_;
wire _20272_;
wire _20273_;
wire _20274_;
wire _20275_;
wire _20276_;
wire _20277_;
wire _20278_;
wire _20279_;
wire _20280_;
wire _20281_;
wire _20282_;
wire _20283_;
wire _20284_;
wire _20285_;
wire _20286_;
wire _20287_;
wire _20288_;
wire _20289_;
wire _20290_;
wire _20291_;
wire _20292_;
wire _20293_;
wire _20294_;
wire _20295_;
wire _20296_;
wire _20297_;
wire _20298_;
wire _20299_;
wire _20300_;
wire _20301_;
wire _20302_;
wire _20303_;
wire _20304_;
wire _20305_;
wire _20306_;
wire _20307_;
wire _20308_;
wire _20309_;
wire _20310_;
wire _20311_;
wire _20312_;
wire _20313_;
wire _20314_;
wire _20315_;
wire _20316_;
wire _20317_;
wire _20318_;
wire _20319_;
wire _20320_;
wire _20321_;
wire _20322_;
wire _20323_;
wire _20324_;
wire _20325_;
wire _20326_;
wire _20327_;
wire _20328_;
wire _20329_;
wire _20330_;
wire _20331_;
wire _20332_;
wire _20333_;
wire _20334_;
wire _20335_;
wire _20336_;
wire _20337_;
wire _20338_;
wire _20339_;
wire _20340_;
wire _20341_;
wire _20342_;
wire _20343_;
wire _20344_;
wire _20345_;
wire _20346_;
wire _20347_;
wire _20348_;
wire _20349_;
wire _20350_;
wire _20351_;
wire _20352_;
wire _20353_;
wire _20354_;
wire _20355_;
wire _20356_;
wire _20357_;
wire _20358_;
wire _20359_;
wire _20360_;
wire _20361_;
wire _20362_;
wire _20363_;
wire _20364_;
wire _20365_;
wire _20366_;
wire _20367_;
wire _20368_;
wire _20369_;
wire _20370_;
wire _20371_;
wire _20372_;
wire _20373_;
wire _20374_;
wire _20375_;
wire _20376_;
wire _20377_;
wire _20378_;
wire _20379_;
wire _20380_;
wire _20381_;
wire _20382_;
wire _20383_;
wire _20384_;
wire _20385_;
wire _20386_;
wire _20387_;
wire _20388_;
wire _20389_;
wire _20390_;
wire _20391_;
wire _20392_;
wire _20393_;
wire _20394_;
wire _20395_;
wire _20396_;
wire _20397_;
wire _20398_;
wire _20399_;
wire _20400_;
wire _20401_;
wire _20402_;
wire _20403_;
wire _20404_;
wire _20405_;
wire _20406_;
wire _20407_;
wire _20408_;
wire _20409_;
wire _20410_;
wire _20411_;
wire _20412_;
wire _20413_;
wire _20414_;
wire _20415_;
wire _20416_;
wire _20417_;
wire _20418_;
wire _20419_;
wire _20420_;
wire _20421_;
wire _20422_;
wire _20423_;
wire _20424_;
wire _20425_;
wire _20426_;
wire _20427_;
wire _20428_;
wire _20429_;
wire _20430_;
wire _20431_;
wire _20432_;
wire _20433_;
wire _20434_;
wire _20435_;
wire _20436_;
wire _20437_;
wire _20438_;
wire _20439_;
wire _20440_;
wire _20441_;
wire _20442_;
wire _20443_;
wire _20444_;
wire _20445_;
wire _20446_;
wire _20447_;
wire _20448_;
wire _20449_;
wire _20450_;
wire _20451_;
wire _20452_;
wire _20453_;
wire _20454_;
wire _20455_;
wire _20456_;
wire _20457_;
wire _20458_;
wire _20459_;
wire _20460_;
wire _20461_;
wire _20462_;
wire _20463_;
wire _20464_;
wire _20465_;
wire _20466_;
wire _20467_;
wire _20468_;
wire _20469_;
wire _20470_;
wire _20471_;
wire _20472_;
wire _20473_;
wire _20474_;
wire _20475_;
wire _20476_;
wire _20477_;
wire _20478_;
wire _20479_;
wire _20480_;
wire _20481_;
wire _20482_;
wire _20483_;
wire _20484_;
wire _20485_;
wire _20486_;
wire _20487_;
wire _20488_;
wire _20489_;
wire _20490_;
wire _20491_;
wire _20492_;
wire _20493_;
wire _20494_;
wire _20495_;
wire _20496_;
wire _20497_;
wire _20498_;
wire _20499_;
wire _20500_;
wire _20501_;
wire _20502_;
wire _20503_;
wire _20504_;
wire _20505_;
wire _20506_;
wire _20507_;
wire _20508_;
wire _20509_;
wire _20510_;
wire _20511_;
wire _20512_;
wire _20513_;
wire _20514_;
wire _20515_;
wire _20516_;
wire _20517_;
wire _20518_;
wire _20519_;
wire _20520_;
wire _20521_;
wire _20522_;
wire _20523_;
wire _20524_;
wire _20525_;
wire _20526_;
wire _20527_;
wire _20528_;
wire _20529_;
wire _20530_;
wire _20531_;
wire _20532_;
wire _20533_;
wire _20534_;
wire _20535_;
wire _20536_;
wire _20537_;
wire _20538_;
wire _20539_;
wire _20540_;
wire _20541_;
wire _20542_;
wire _20543_;
wire _20544_;
wire _20545_;
wire _20546_;
wire _20547_;
wire _20548_;
wire _20549_;
wire _20550_;
wire _20551_;
wire _20552_;
wire _20553_;
wire _20554_;
wire _20555_;
wire _20556_;
wire _20557_;
wire _20558_;
wire _20559_;
wire _20560_;
wire _20561_;
wire _20562_;
wire _20563_;
wire _20564_;
wire _20565_;
wire _20566_;
wire _20567_;
wire _20568_;
wire _20569_;
wire _20570_;
wire _20571_;
wire _20572_;
wire _20573_;
wire _20574_;
wire _20575_;
wire _20576_;
wire _20577_;
wire _20578_;
wire _20579_;
wire _20580_;
wire _20581_;
wire _20582_;
wire _20583_;
wire _20584_;
wire _20585_;
wire _20586_;
wire _20587_;
wire _20588_;
wire _20589_;
wire _20590_;
wire _20591_;
wire _20592_;
wire _20593_;
wire _20594_;
wire _20595_;
wire _20596_;
wire _20597_;
wire _20598_;
wire _20599_;
wire _20600_;
wire _20601_;
wire _20602_;
wire _20603_;
wire _20604_;
wire _20605_;
wire _20606_;
wire _20607_;
wire _20608_;
wire _20609_;
wire _20610_;
wire _20611_;
wire _20612_;
wire _20613_;
wire _20614_;
wire _20615_;
wire _20616_;
wire _20617_;
wire _20618_;
wire _20619_;
wire _20620_;
wire _20621_;
wire _20622_;
wire _20623_;
wire _20624_;
wire _20625_;
wire _20626_;
wire _20627_;
wire _20628_;
wire _20629_;
wire _20630_;
wire _20631_;
wire _20632_;
wire _20633_;
wire _20634_;
wire _20635_;
wire _20636_;
wire _20637_;
wire _20638_;
wire _20639_;
wire _20640_;
wire _20641_;
wire _20642_;
wire _20643_;
wire _20644_;
wire _20645_;
wire _20646_;
wire _20647_;
wire _20648_;
wire _20649_;
wire _20650_;
wire _20651_;
wire _20652_;
wire _20653_;
wire _20654_;
wire _20655_;
wire _20656_;
wire _20657_;
wire _20658_;
wire _20659_;
wire _20660_;
wire _20661_;
wire _20662_;
wire _20663_;
wire _20664_;
wire _20665_;
wire _20666_;
wire _20667_;
wire _20668_;
wire _20669_;
wire _20670_;
wire _20671_;
wire _20672_;
wire _20673_;
wire _20674_;
wire _20675_;
wire _20676_;
wire _20677_;
wire _20678_;
wire _20679_;
wire _20680_;
wire _20681_;
wire _20682_;
wire _20683_;
wire _20684_;
wire _20685_;
wire _20686_;
wire _20687_;
wire _20688_;
wire _20689_;
wire _20690_;
wire _20691_;
wire _20692_;
wire _20693_;
wire _20694_;
wire _20695_;
wire _20696_;
wire _20697_;
wire _20698_;
wire _20699_;
wire _20700_;
wire _20701_;
wire _20702_;
wire _20703_;
wire _20704_;
wire _20705_;
wire _20706_;
wire _20707_;
wire _20708_;
wire _20709_;
wire _20710_;
wire _20711_;
wire _20712_;
wire _20713_;
wire _20714_;
wire _20715_;
wire _20716_;
wire _20717_;
wire _20718_;
wire _20719_;
wire _20720_;
wire _20721_;
wire _20722_;
wire _20723_;
wire _20724_;
wire _20725_;
wire _20726_;
wire _20727_;
wire _20728_;
wire _20729_;
wire _20730_;
wire _20731_;
wire _20732_;
wire _20733_;
wire _20734_;
wire _20735_;
wire _20736_;
wire _20737_;
wire _20738_;
wire _20739_;
wire _20740_;
wire _20741_;
wire _20742_;
wire _20743_;
wire _20744_;
wire _20745_;
wire _20746_;
wire _20747_;
wire _20748_;
wire _20749_;
wire _20750_;
wire _20751_;
wire _20752_;
wire _20753_;
wire _20754_;
wire _20755_;
wire _20756_;
wire _20757_;
wire _20758_;
wire _20759_;
wire _20760_;
wire _20761_;
wire _20762_;
wire _20763_;
wire _20764_;
wire _20765_;
wire _20766_;
wire _20767_;
wire _20768_;
wire _20769_;
wire _20770_;
wire _20771_;
wire _20772_;
wire _20773_;
wire _20774_;
wire _20775_;
wire _20776_;
wire _20777_;
wire _20778_;
wire _20779_;
wire _20780_;
wire _20781_;
wire _20782_;
wire _20783_;
wire _20784_;
wire _20785_;
wire _20786_;
wire _20787_;
wire _20788_;
wire _20789_;
wire _20790_;
wire _20791_;
wire _20792_;
wire _20793_;
wire _20794_;
wire _20795_;
wire _20796_;
wire _20797_;
wire _20798_;
wire _20799_;
wire _20800_;
wire _20801_;
wire _20802_;
wire _20803_;
wire _20804_;
wire _20805_;
wire _20806_;
wire _20807_;
wire _20808_;
wire _20809_;
wire _20810_;
wire _20811_;
wire _20812_;
wire _20813_;
wire _20814_;
wire _20815_;
wire _20816_;
wire _20817_;
wire _20818_;
wire _20819_;
wire _20820_;
wire _20821_;
wire _20822_;
wire _20823_;
wire _20824_;
wire _20825_;
wire _20826_;
wire _20827_;
wire _20828_;
wire _20829_;
wire _20830_;
wire _20831_;
wire _20832_;
wire _20833_;
wire _20834_;
wire _20835_;
wire _20836_;
wire _20837_;
wire _20838_;
wire _20839_;
wire _20840_;
wire _20841_;
wire _20842_;
wire _20843_;
wire _20844_;
wire _20845_;
wire _20846_;
wire _20847_;
wire _20848_;
wire _20849_;
wire _20850_;
wire _20851_;
wire _20852_;
wire _20853_;
wire _20854_;
wire _20855_;
wire _20856_;
wire _20857_;
wire _20858_;
wire _20859_;
wire _20860_;
wire _20861_;
wire _20862_;
wire _20863_;
wire _20864_;
wire _20865_;
wire _20866_;
wire _20867_;
wire _20868_;
wire _20869_;
wire _20870_;
wire _20871_;
wire _20872_;
wire _20873_;
wire _20874_;
wire _20875_;
wire _20876_;
wire _20877_;
wire _20878_;
wire _20879_;
wire _20880_;
wire _20881_;
wire _20882_;
wire _20883_;
wire _20884_;
wire _20885_;
wire _20886_;
wire _20887_;
wire _20888_;
wire _20889_;
wire _20890_;
wire _20891_;
wire _20892_;
wire _20893_;
wire _20894_;
wire _20895_;
wire _20896_;
wire _20897_;
wire _20898_;
wire _20899_;
wire _20900_;
wire _20901_;
wire _20902_;
wire _20903_;
wire _20904_;
wire _20905_;
wire _20906_;
wire _20907_;
wire _20908_;
wire _20909_;
wire _20910_;
wire _20911_;
wire _20912_;
wire _20913_;
wire _20914_;
wire _20915_;
wire _20916_;
wire _20917_;
wire _20918_;
wire _20919_;
wire _20920_;
wire _20921_;
wire _20922_;
wire _20923_;
wire _20924_;
wire _20925_;
wire _20926_;
wire _20927_;
wire _20928_;
wire _20929_;
wire _20930_;
wire _20931_;
wire _20932_;
wire _20933_;
wire _20934_;
wire _20935_;
wire _20936_;
wire _20937_;
wire _20938_;
wire _20939_;
wire _20940_;
wire _20941_;
wire _20942_;
wire _20943_;
wire _20944_;
wire _20945_;
wire _20946_;
wire _20947_;
wire _20948_;
wire _20949_;
wire _20950_;
wire _20951_;
wire _20952_;
wire _20953_;
wire _20954_;
wire _20955_;
wire _20956_;
wire _20957_;
wire _20958_;
wire _20959_;
wire _20960_;
wire _20961_;
wire _20962_;
wire _20963_;
wire _20964_;
wire _20965_;
wire _20966_;
wire _20967_;
wire _20968_;
wire _20969_;
wire _20970_;
wire _20971_;
wire _20972_;
wire _20973_;
wire _20974_;
wire _20975_;
wire _20976_;
wire _20977_;
wire _20978_;
wire _20979_;
wire _20980_;
wire _20981_;
wire _20982_;
wire _20983_;
wire _20984_;
wire _20985_;
wire _20986_;
wire _20987_;
wire _20988_;
wire _20989_;
wire _20990_;
wire _20991_;
wire _20992_;
wire _20993_;
wire _20994_;
wire _20995_;
wire _20996_;
wire _20997_;
wire _20998_;
wire _20999_;
wire _21000_;
wire _21001_;
wire _21002_;
wire _21003_;
wire _21004_;
wire _21005_;
wire _21006_;
wire _21007_;
wire _21008_;
wire _21009_;
wire _21010_;
wire _21011_;
wire _21012_;
wire _21013_;
wire _21014_;
wire _21015_;
wire _21016_;
wire _21017_;
wire _21018_;
wire _21019_;
wire _21020_;
wire _21021_;
wire _21022_;
wire _21023_;
wire _21024_;
wire _21025_;
wire _21026_;
wire _21027_;
wire _21028_;
wire _21029_;
wire _21030_;
wire _21031_;
wire _21032_;
wire _21033_;
wire _21034_;
wire _21035_;
wire _21036_;
wire _21037_;
wire _21038_;
wire _21039_;
wire _21040_;
wire _21041_;
wire _21042_;
wire _21043_;
wire _21044_;
wire _21045_;
wire _21046_;
wire _21047_;
wire _21048_;
wire _21049_;
wire _21050_;
wire _21051_;
wire _21052_;
wire _21053_;
wire _21054_;
wire _21055_;
wire _21056_;
wire _21057_;
wire _21058_;
wire _21059_;
wire _21060_;
wire _21061_;
wire _21062_;
wire _21063_;
wire _21064_;
wire _21065_;
wire _21066_;
wire _21067_;
wire _21068_;
wire _21069_;
wire _21070_;
wire _21071_;
wire _21072_;
wire _21073_;
wire _21074_;
wire _21075_;
wire _21076_;
wire _21077_;
wire _21078_;
wire _21079_;
wire _21080_;
wire _21081_;
wire _21082_;
wire _21083_;
wire _21084_;
wire _21085_;
wire _21086_;
wire _21087_;
wire _21088_;
wire _21089_;
wire _21090_;
wire _21091_;
wire _21092_;
wire _21093_;
wire _21094_;
wire _21095_;
wire _21096_;
wire _21097_;
wire _21098_;
wire _21099_;
wire _21100_;
wire _21101_;
wire _21102_;
wire _21103_;
wire _21104_;
wire _21105_;
wire zeroWire;
wire oneWire;
assign zeroWire = 1'b0 /*25202*/;
assign oneWire = 1'b1 /*25202*/;
assign _37_ = ~D[0] /*25008*/;
assign _34_ = R_0[31] & _37_ /*25004*/;
assign _35_ = R_0[31] ^ _37_ /*25007*/;
assign _36_ = oneWire & _35_ /*25005*/;
assign _0_ = oneWire ^ _35_ /*25006*/;
assign _33_ = _34_ | _36_ /*25003*/;
assign _42_ = ~D[1] /*25002*/;
assign _39_ = R_0[32] & _42_ /*24998*/;
assign _40_ = R_0[32] ^ _42_ /*25001*/;
assign _41_ = _33_ & _40_ /*24999*/;
assign _1_ = _33_ ^ _40_ /*25000*/;
assign _38_ = _39_ | _41_ /*24997*/;
assign _47_ = ~D[2] /*24996*/;
assign _44_ = R_0[33] & _47_ /*24992*/;
assign _45_ = R_0[33] ^ _47_ /*24995*/;
assign _46_ = _38_ & _45_ /*24993*/;
assign _2_ = _38_ ^ _45_ /*24994*/;
assign _43_ = _44_ | _46_ /*24991*/;
assign _52_ = ~D[3] /*24990*/;
assign _49_ = R_0[34] & _52_ /*24986*/;
assign _50_ = R_0[34] ^ _52_ /*24989*/;
assign _51_ = _43_ & _50_ /*24987*/;
assign _3_ = _43_ ^ _50_ /*24988*/;
assign _48_ = _49_ | _51_ /*24985*/;
assign _57_ = ~D[4] /*24984*/;
assign _54_ = R_0[35] & _57_ /*24980*/;
assign _55_ = R_0[35] ^ _57_ /*24983*/;
assign _56_ = _48_ & _55_ /*24981*/;
assign _4_ = _48_ ^ _55_ /*24982*/;
assign _53_ = _54_ | _56_ /*24979*/;
assign _62_ = ~D[5] /*24978*/;
assign _59_ = R_0[36] & _62_ /*24974*/;
assign _60_ = R_0[36] ^ _62_ /*24977*/;
assign _61_ = _53_ & _60_ /*24975*/;
assign _5_ = _53_ ^ _60_ /*24976*/;
assign _58_ = _59_ | _61_ /*24973*/;
assign _67_ = ~D[6] /*24972*/;
assign _64_ = R_0[37] & _67_ /*24968*/;
assign _65_ = R_0[37] ^ _67_ /*24971*/;
assign _66_ = _58_ & _65_ /*24969*/;
assign _6_ = _58_ ^ _65_ /*24970*/;
assign _63_ = _64_ | _66_ /*24967*/;
assign _72_ = ~D[7] /*24966*/;
assign _69_ = R_0[38] & _72_ /*24962*/;
assign _70_ = R_0[38] ^ _72_ /*24965*/;
assign _71_ = _63_ & _70_ /*24963*/;
assign _7_ = _63_ ^ _70_ /*24964*/;
assign _68_ = _69_ | _71_ /*24961*/;
assign _77_ = ~D[8] /*24960*/;
assign _74_ = R_0[39] & _77_ /*24956*/;
assign _75_ = R_0[39] ^ _77_ /*24959*/;
assign _76_ = _68_ & _75_ /*24957*/;
assign _8_ = _68_ ^ _75_ /*24958*/;
assign _73_ = _74_ | _76_ /*24955*/;
assign _82_ = ~D[9] /*24954*/;
assign _79_ = R_0[40] & _82_ /*24950*/;
assign _80_ = R_0[40] ^ _82_ /*24953*/;
assign _81_ = _73_ & _80_ /*24951*/;
assign _9_ = _73_ ^ _80_ /*24952*/;
assign _78_ = _79_ | _81_ /*24949*/;
assign _87_ = ~D[10] /*24948*/;
assign _84_ = R_0[41] & _87_ /*24944*/;
assign _85_ = R_0[41] ^ _87_ /*24947*/;
assign _86_ = _78_ & _85_ /*24945*/;
assign _10_ = _78_ ^ _85_ /*24946*/;
assign _83_ = _84_ | _86_ /*24943*/;
assign _92_ = ~D[11] /*24942*/;
assign _89_ = R_0[42] & _92_ /*24938*/;
assign _90_ = R_0[42] ^ _92_ /*24941*/;
assign _91_ = _83_ & _90_ /*24939*/;
assign _11_ = _83_ ^ _90_ /*24940*/;
assign _88_ = _89_ | _91_ /*24937*/;
assign _97_ = ~D[12] /*24936*/;
assign _94_ = R_0[43] & _97_ /*24932*/;
assign _95_ = R_0[43] ^ _97_ /*24935*/;
assign _96_ = _88_ & _95_ /*24933*/;
assign _12_ = _88_ ^ _95_ /*24934*/;
assign _93_ = _94_ | _96_ /*24931*/;
assign _102_ = ~D[13] /*24930*/;
assign _99_ = R_0[44] & _102_ /*24926*/;
assign _100_ = R_0[44] ^ _102_ /*24929*/;
assign _101_ = _93_ & _100_ /*24927*/;
assign _13_ = _93_ ^ _100_ /*24928*/;
assign _98_ = _99_ | _101_ /*24925*/;
assign _107_ = ~D[14] /*24924*/;
assign _104_ = R_0[45] & _107_ /*24920*/;
assign _105_ = R_0[45] ^ _107_ /*24923*/;
assign _106_ = _98_ & _105_ /*24921*/;
assign _14_ = _98_ ^ _105_ /*24922*/;
assign _103_ = _104_ | _106_ /*24919*/;
assign _112_ = ~D[15] /*24918*/;
assign _109_ = R_0[46] & _112_ /*24914*/;
assign _110_ = R_0[46] ^ _112_ /*24917*/;
assign _111_ = _103_ & _110_ /*24915*/;
assign _15_ = _103_ ^ _110_ /*24916*/;
assign _108_ = _109_ | _111_ /*24913*/;
assign _117_ = ~D[16] /*24912*/;
assign _114_ = R_0[47] & _117_ /*24908*/;
assign _115_ = R_0[47] ^ _117_ /*24911*/;
assign _116_ = _108_ & _115_ /*24909*/;
assign _16_ = _108_ ^ _115_ /*24910*/;
assign _113_ = _114_ | _116_ /*24907*/;
assign _122_ = ~D[17] /*24906*/;
assign _119_ = R_0[48] & _122_ /*24902*/;
assign _120_ = R_0[48] ^ _122_ /*24905*/;
assign _121_ = _113_ & _120_ /*24903*/;
assign _17_ = _113_ ^ _120_ /*24904*/;
assign _118_ = _119_ | _121_ /*24901*/;
assign _127_ = ~D[18] /*24900*/;
assign _124_ = R_0[49] & _127_ /*24896*/;
assign _125_ = R_0[49] ^ _127_ /*24899*/;
assign _126_ = _118_ & _125_ /*24897*/;
assign _18_ = _118_ ^ _125_ /*24898*/;
assign _123_ = _124_ | _126_ /*24895*/;
assign _132_ = ~D[19] /*24894*/;
assign _129_ = R_0[50] & _132_ /*24890*/;
assign _130_ = R_0[50] ^ _132_ /*24893*/;
assign _131_ = _123_ & _130_ /*24891*/;
assign _19_ = _123_ ^ _130_ /*24892*/;
assign _128_ = _129_ | _131_ /*24889*/;
assign _137_ = ~D[20] /*24888*/;
assign _134_ = R_0[51] & _137_ /*24884*/;
assign _135_ = R_0[51] ^ _137_ /*24887*/;
assign _136_ = _128_ & _135_ /*24885*/;
assign _20_ = _128_ ^ _135_ /*24886*/;
assign _133_ = _134_ | _136_ /*24883*/;
assign _142_ = ~D[21] /*24882*/;
assign _139_ = R_0[52] & _142_ /*24878*/;
assign _140_ = R_0[52] ^ _142_ /*24881*/;
assign _141_ = _133_ & _140_ /*24879*/;
assign _21_ = _133_ ^ _140_ /*24880*/;
assign _138_ = _139_ | _141_ /*24877*/;
assign _147_ = ~D[22] /*24876*/;
assign _144_ = R_0[53] & _147_ /*24872*/;
assign _145_ = R_0[53] ^ _147_ /*24875*/;
assign _146_ = _138_ & _145_ /*24873*/;
assign _22_ = _138_ ^ _145_ /*24874*/;
assign _143_ = _144_ | _146_ /*24871*/;
assign _152_ = ~D[23] /*24870*/;
assign _149_ = R_0[54] & _152_ /*24866*/;
assign _150_ = R_0[54] ^ _152_ /*24869*/;
assign _151_ = _143_ & _150_ /*24867*/;
assign _23_ = _143_ ^ _150_ /*24868*/;
assign _148_ = _149_ | _151_ /*24865*/;
assign _157_ = ~D[24] /*24864*/;
assign _154_ = R_0[55] & _157_ /*24860*/;
assign _155_ = R_0[55] ^ _157_ /*24863*/;
assign _156_ = _148_ & _155_ /*24861*/;
assign _24_ = _148_ ^ _155_ /*24862*/;
assign _153_ = _154_ | _156_ /*24859*/;
assign _162_ = ~D[25] /*24858*/;
assign _159_ = R_0[56] & _162_ /*24854*/;
assign _160_ = R_0[56] ^ _162_ /*24857*/;
assign _161_ = _153_ & _160_ /*24855*/;
assign _25_ = _153_ ^ _160_ /*24856*/;
assign _158_ = _159_ | _161_ /*24853*/;
assign _167_ = ~D[26] /*24852*/;
assign _164_ = R_0[57] & _167_ /*24848*/;
assign _165_ = R_0[57] ^ _167_ /*24851*/;
assign _166_ = _158_ & _165_ /*24849*/;
assign _26_ = _158_ ^ _165_ /*24850*/;
assign _163_ = _164_ | _166_ /*24847*/;
assign _172_ = ~D[27] /*24846*/;
assign _169_ = R_0[58] & _172_ /*24842*/;
assign _170_ = R_0[58] ^ _172_ /*24845*/;
assign _171_ = _163_ & _170_ /*24843*/;
assign _27_ = _163_ ^ _170_ /*24844*/;
assign _168_ = _169_ | _171_ /*24841*/;
assign _177_ = ~D[28] /*24840*/;
assign _174_ = R_0[59] & _177_ /*24836*/;
assign _175_ = R_0[59] ^ _177_ /*24839*/;
assign _176_ = _168_ & _175_ /*24837*/;
assign _28_ = _168_ ^ _175_ /*24838*/;
assign _173_ = _174_ | _176_ /*24835*/;
assign _182_ = ~D[29] /*24834*/;
assign _179_ = R_0[60] & _182_ /*24830*/;
assign _180_ = R_0[60] ^ _182_ /*24833*/;
assign _181_ = _173_ & _180_ /*24831*/;
assign _29_ = _173_ ^ _180_ /*24832*/;
assign _178_ = _179_ | _181_ /*24829*/;
assign _187_ = ~D[30] /*24828*/;
assign _184_ = R_0[61] & _187_ /*24824*/;
assign _185_ = R_0[61] ^ _187_ /*24827*/;
assign _186_ = _178_ & _185_ /*24825*/;
assign _30_ = _178_ ^ _185_ /*24826*/;
assign _183_ = _184_ | _186_ /*24823*/;
assign _188_ = zeroWire & oneWire /*24818*/;
assign _189_ = zeroWire ^ oneWire /*24821*/;
assign _190_ = _183_ & _189_ /*24819*/;
assign _31_ = _183_ ^ _189_ /*24820*/;
assign Q[31] = _188_ | _190_ /*24817*/;
assign _227_ = ~Q[31] /*24625*/;
assign _226_ = _227_ & D[0] /*24624*/;
assign _229_ = _0_ & _226_ /*24619*/;
assign _230_ = _0_ ^ _226_ /*24622*/;
assign _231_ = zeroWire & _230_ /*24620*/;
assign _193_ = zeroWire ^ _230_ /*24621*/;
assign _228_ = _229_ | _231_ /*24618*/;
assign _233_ = ~Q[31] /*24617*/;
assign _232_ = _233_ & D[1] /*24616*/;
assign _235_ = _1_ & _232_ /*24611*/;
assign _236_ = _1_ ^ _232_ /*24614*/;
assign _237_ = _228_ & _236_ /*24612*/;
assign _194_ = _228_ ^ _236_ /*24613*/;
assign _234_ = _235_ | _237_ /*24610*/;
assign _239_ = ~Q[31] /*24609*/;
assign _238_ = _239_ & D[2] /*24608*/;
assign _241_ = _2_ & _238_ /*24603*/;
assign _242_ = _2_ ^ _238_ /*24606*/;
assign _243_ = _234_ & _242_ /*24604*/;
assign _195_ = _234_ ^ _242_ /*24605*/;
assign _240_ = _241_ | _243_ /*24602*/;
assign _245_ = ~Q[31] /*24601*/;
assign _244_ = _245_ & D[3] /*24600*/;
assign _247_ = _3_ & _244_ /*24595*/;
assign _248_ = _3_ ^ _244_ /*24598*/;
assign _249_ = _240_ & _248_ /*24596*/;
assign _196_ = _240_ ^ _248_ /*24597*/;
assign _246_ = _247_ | _249_ /*24594*/;
assign _251_ = ~Q[31] /*24593*/;
assign _250_ = _251_ & D[4] /*24592*/;
assign _253_ = _4_ & _250_ /*24587*/;
assign _254_ = _4_ ^ _250_ /*24590*/;
assign _255_ = _246_ & _254_ /*24588*/;
assign _197_ = _246_ ^ _254_ /*24589*/;
assign _252_ = _253_ | _255_ /*24586*/;
assign _257_ = ~Q[31] /*24585*/;
assign _256_ = _257_ & D[5] /*24584*/;
assign _259_ = _5_ & _256_ /*24579*/;
assign _260_ = _5_ ^ _256_ /*24582*/;
assign _261_ = _252_ & _260_ /*24580*/;
assign _198_ = _252_ ^ _260_ /*24581*/;
assign _258_ = _259_ | _261_ /*24578*/;
assign _263_ = ~Q[31] /*24577*/;
assign _262_ = _263_ & D[6] /*24576*/;
assign _265_ = _6_ & _262_ /*24571*/;
assign _266_ = _6_ ^ _262_ /*24574*/;
assign _267_ = _258_ & _266_ /*24572*/;
assign _199_ = _258_ ^ _266_ /*24573*/;
assign _264_ = _265_ | _267_ /*24570*/;
assign _269_ = ~Q[31] /*24569*/;
assign _268_ = _269_ & D[7] /*24568*/;
assign _271_ = _7_ & _268_ /*24563*/;
assign _272_ = _7_ ^ _268_ /*24566*/;
assign _273_ = _264_ & _272_ /*24564*/;
assign _200_ = _264_ ^ _272_ /*24565*/;
assign _270_ = _271_ | _273_ /*24562*/;
assign _275_ = ~Q[31] /*24561*/;
assign _274_ = _275_ & D[8] /*24560*/;
assign _277_ = _8_ & _274_ /*24555*/;
assign _278_ = _8_ ^ _274_ /*24558*/;
assign _279_ = _270_ & _278_ /*24556*/;
assign _201_ = _270_ ^ _278_ /*24557*/;
assign _276_ = _277_ | _279_ /*24554*/;
assign _281_ = ~Q[31] /*24553*/;
assign _280_ = _281_ & D[9] /*24552*/;
assign _283_ = _9_ & _280_ /*24547*/;
assign _284_ = _9_ ^ _280_ /*24550*/;
assign _285_ = _276_ & _284_ /*24548*/;
assign _202_ = _276_ ^ _284_ /*24549*/;
assign _282_ = _283_ | _285_ /*24546*/;
assign _287_ = ~Q[31] /*24545*/;
assign _286_ = _287_ & D[10] /*24544*/;
assign _289_ = _10_ & _286_ /*24539*/;
assign _290_ = _10_ ^ _286_ /*24542*/;
assign _291_ = _282_ & _290_ /*24540*/;
assign _203_ = _282_ ^ _290_ /*24541*/;
assign _288_ = _289_ | _291_ /*24538*/;
assign _293_ = ~Q[31] /*24537*/;
assign _292_ = _293_ & D[11] /*24536*/;
assign _295_ = _11_ & _292_ /*24531*/;
assign _296_ = _11_ ^ _292_ /*24534*/;
assign _297_ = _288_ & _296_ /*24532*/;
assign _204_ = _288_ ^ _296_ /*24533*/;
assign _294_ = _295_ | _297_ /*24530*/;
assign _299_ = ~Q[31] /*24529*/;
assign _298_ = _299_ & D[12] /*24528*/;
assign _301_ = _12_ & _298_ /*24523*/;
assign _302_ = _12_ ^ _298_ /*24526*/;
assign _303_ = _294_ & _302_ /*24524*/;
assign _205_ = _294_ ^ _302_ /*24525*/;
assign _300_ = _301_ | _303_ /*24522*/;
assign _305_ = ~Q[31] /*24521*/;
assign _304_ = _305_ & D[13] /*24520*/;
assign _307_ = _13_ & _304_ /*24515*/;
assign _308_ = _13_ ^ _304_ /*24518*/;
assign _309_ = _300_ & _308_ /*24516*/;
assign _206_ = _300_ ^ _308_ /*24517*/;
assign _306_ = _307_ | _309_ /*24514*/;
assign _311_ = ~Q[31] /*24513*/;
assign _310_ = _311_ & D[14] /*24512*/;
assign _313_ = _14_ & _310_ /*24507*/;
assign _314_ = _14_ ^ _310_ /*24510*/;
assign _315_ = _306_ & _314_ /*24508*/;
assign _207_ = _306_ ^ _314_ /*24509*/;
assign _312_ = _313_ | _315_ /*24506*/;
assign _317_ = ~Q[31] /*24505*/;
assign _316_ = _317_ & D[15] /*24504*/;
assign _319_ = _15_ & _316_ /*24499*/;
assign _320_ = _15_ ^ _316_ /*24502*/;
assign _321_ = _312_ & _320_ /*24500*/;
assign _208_ = _312_ ^ _320_ /*24501*/;
assign _318_ = _319_ | _321_ /*24498*/;
assign _323_ = ~Q[31] /*24497*/;
assign _322_ = _323_ & D[16] /*24496*/;
assign _325_ = _16_ & _322_ /*24491*/;
assign _326_ = _16_ ^ _322_ /*24494*/;
assign _327_ = _318_ & _326_ /*24492*/;
assign _209_ = _318_ ^ _326_ /*24493*/;
assign _324_ = _325_ | _327_ /*24490*/;
assign _329_ = ~Q[31] /*24489*/;
assign _328_ = _329_ & D[17] /*24488*/;
assign _331_ = _17_ & _328_ /*24483*/;
assign _332_ = _17_ ^ _328_ /*24486*/;
assign _333_ = _324_ & _332_ /*24484*/;
assign _210_ = _324_ ^ _332_ /*24485*/;
assign _330_ = _331_ | _333_ /*24482*/;
assign _335_ = ~Q[31] /*24481*/;
assign _334_ = _335_ & D[18] /*24480*/;
assign _337_ = _18_ & _334_ /*24475*/;
assign _338_ = _18_ ^ _334_ /*24478*/;
assign _339_ = _330_ & _338_ /*24476*/;
assign _211_ = _330_ ^ _338_ /*24477*/;
assign _336_ = _337_ | _339_ /*24474*/;
assign _341_ = ~Q[31] /*24473*/;
assign _340_ = _341_ & D[19] /*24472*/;
assign _343_ = _19_ & _340_ /*24467*/;
assign _344_ = _19_ ^ _340_ /*24470*/;
assign _345_ = _336_ & _344_ /*24468*/;
assign _212_ = _336_ ^ _344_ /*24469*/;
assign _342_ = _343_ | _345_ /*24466*/;
assign _347_ = ~Q[31] /*24465*/;
assign _346_ = _347_ & D[20] /*24464*/;
assign _349_ = _20_ & _346_ /*24459*/;
assign _350_ = _20_ ^ _346_ /*24462*/;
assign _351_ = _342_ & _350_ /*24460*/;
assign _213_ = _342_ ^ _350_ /*24461*/;
assign _348_ = _349_ | _351_ /*24458*/;
assign _353_ = ~Q[31] /*24457*/;
assign _352_ = _353_ & D[21] /*24456*/;
assign _355_ = _21_ & _352_ /*24451*/;
assign _356_ = _21_ ^ _352_ /*24454*/;
assign _357_ = _348_ & _356_ /*24452*/;
assign _214_ = _348_ ^ _356_ /*24453*/;
assign _354_ = _355_ | _357_ /*24450*/;
assign _359_ = ~Q[31] /*24449*/;
assign _358_ = _359_ & D[22] /*24448*/;
assign _361_ = _22_ & _358_ /*24443*/;
assign _362_ = _22_ ^ _358_ /*24446*/;
assign _363_ = _354_ & _362_ /*24444*/;
assign _215_ = _354_ ^ _362_ /*24445*/;
assign _360_ = _361_ | _363_ /*24442*/;
assign _365_ = ~Q[31] /*24441*/;
assign _364_ = _365_ & D[23] /*24440*/;
assign _367_ = _23_ & _364_ /*24435*/;
assign _368_ = _23_ ^ _364_ /*24438*/;
assign _369_ = _360_ & _368_ /*24436*/;
assign _216_ = _360_ ^ _368_ /*24437*/;
assign _366_ = _367_ | _369_ /*24434*/;
assign _371_ = ~Q[31] /*24433*/;
assign _370_ = _371_ & D[24] /*24432*/;
assign _373_ = _24_ & _370_ /*24427*/;
assign _374_ = _24_ ^ _370_ /*24430*/;
assign _375_ = _366_ & _374_ /*24428*/;
assign _217_ = _366_ ^ _374_ /*24429*/;
assign _372_ = _373_ | _375_ /*24426*/;
assign _377_ = ~Q[31] /*24425*/;
assign _376_ = _377_ & D[25] /*24424*/;
assign _379_ = _25_ & _376_ /*24419*/;
assign _380_ = _25_ ^ _376_ /*24422*/;
assign _381_ = _372_ & _380_ /*24420*/;
assign _218_ = _372_ ^ _380_ /*24421*/;
assign _378_ = _379_ | _381_ /*24418*/;
assign _383_ = ~Q[31] /*24417*/;
assign _382_ = _383_ & D[26] /*24416*/;
assign _385_ = _26_ & _382_ /*24411*/;
assign _386_ = _26_ ^ _382_ /*24414*/;
assign _387_ = _378_ & _386_ /*24412*/;
assign _219_ = _378_ ^ _386_ /*24413*/;
assign _384_ = _385_ | _387_ /*24410*/;
assign _389_ = ~Q[31] /*24409*/;
assign _388_ = _389_ & D[27] /*24408*/;
assign _391_ = _27_ & _388_ /*24403*/;
assign _392_ = _27_ ^ _388_ /*24406*/;
assign _393_ = _384_ & _392_ /*24404*/;
assign _220_ = _384_ ^ _392_ /*24405*/;
assign _390_ = _391_ | _393_ /*24402*/;
assign _395_ = ~Q[31] /*24401*/;
assign _394_ = _395_ & D[28] /*24400*/;
assign _397_ = _28_ & _394_ /*24395*/;
assign _398_ = _28_ ^ _394_ /*24398*/;
assign _399_ = _390_ & _398_ /*24396*/;
assign _221_ = _390_ ^ _398_ /*24397*/;
assign _396_ = _397_ | _399_ /*24394*/;
assign _401_ = ~Q[31] /*24393*/;
assign _400_ = _401_ & D[29] /*24392*/;
assign _403_ = _29_ & _400_ /*24387*/;
assign _404_ = _29_ ^ _400_ /*24390*/;
assign _405_ = _396_ & _404_ /*24388*/;
assign _222_ = _396_ ^ _404_ /*24389*/;
assign _402_ = _403_ | _405_ /*24386*/;
assign _407_ = ~Q[31] /*24385*/;
assign _406_ = _407_ & D[30] /*24384*/;
assign _409_ = _30_ & _406_ /*24379*/;
assign _410_ = _30_ ^ _406_ /*24382*/;
assign _411_ = _402_ & _410_ /*24380*/;
assign _223_ = _402_ ^ _410_ /*24381*/;
assign _408_ = _409_ | _411_ /*24378*/;
assign _413_ = ~Q[31] /*24377*/;
assign _412_ = _413_ & zeroWire /*24376*/;
assign _414_ = _31_ ^ _412_ /*24374*/;
assign _224_ = _414_ ^ _408_ /*24373*/;
assign _453_ = ~D[0] /*24247*/;
assign _450_ = R_0[30] & _453_ /*24243*/;
assign _451_ = R_0[30] ^ _453_ /*24246*/;
assign _452_ = oneWire & _451_ /*24244*/;
assign _417_ = oneWire ^ _451_ /*24245*/;
assign _449_ = _450_ | _452_ /*24242*/;
assign _458_ = ~D[1] /*24241*/;
assign _455_ = _193_ & _458_ /*24237*/;
assign _456_ = _193_ ^ _458_ /*24240*/;
assign _457_ = _449_ & _456_ /*24238*/;
assign _418_ = _449_ ^ _456_ /*24239*/;
assign _454_ = _455_ | _457_ /*24236*/;
assign _463_ = ~D[2] /*24235*/;
assign _460_ = _194_ & _463_ /*24231*/;
assign _461_ = _194_ ^ _463_ /*24234*/;
assign _462_ = _454_ & _461_ /*24232*/;
assign _419_ = _454_ ^ _461_ /*24233*/;
assign _459_ = _460_ | _462_ /*24230*/;
assign _468_ = ~D[3] /*24229*/;
assign _465_ = _195_ & _468_ /*24225*/;
assign _466_ = _195_ ^ _468_ /*24228*/;
assign _467_ = _459_ & _466_ /*24226*/;
assign _420_ = _459_ ^ _466_ /*24227*/;
assign _464_ = _465_ | _467_ /*24224*/;
assign _473_ = ~D[4] /*24223*/;
assign _470_ = _196_ & _473_ /*24219*/;
assign _471_ = _196_ ^ _473_ /*24222*/;
assign _472_ = _464_ & _471_ /*24220*/;
assign _421_ = _464_ ^ _471_ /*24221*/;
assign _469_ = _470_ | _472_ /*24218*/;
assign _478_ = ~D[5] /*24217*/;
assign _475_ = _197_ & _478_ /*24213*/;
assign _476_ = _197_ ^ _478_ /*24216*/;
assign _477_ = _469_ & _476_ /*24214*/;
assign _422_ = _469_ ^ _476_ /*24215*/;
assign _474_ = _475_ | _477_ /*24212*/;
assign _483_ = ~D[6] /*24211*/;
assign _480_ = _198_ & _483_ /*24207*/;
assign _481_ = _198_ ^ _483_ /*24210*/;
assign _482_ = _474_ & _481_ /*24208*/;
assign _423_ = _474_ ^ _481_ /*24209*/;
assign _479_ = _480_ | _482_ /*24206*/;
assign _488_ = ~D[7] /*24205*/;
assign _485_ = _199_ & _488_ /*24201*/;
assign _486_ = _199_ ^ _488_ /*24204*/;
assign _487_ = _479_ & _486_ /*24202*/;
assign _424_ = _479_ ^ _486_ /*24203*/;
assign _484_ = _485_ | _487_ /*24200*/;
assign _493_ = ~D[8] /*24199*/;
assign _490_ = _200_ & _493_ /*24195*/;
assign _491_ = _200_ ^ _493_ /*24198*/;
assign _492_ = _484_ & _491_ /*24196*/;
assign _425_ = _484_ ^ _491_ /*24197*/;
assign _489_ = _490_ | _492_ /*24194*/;
assign _498_ = ~D[9] /*24193*/;
assign _495_ = _201_ & _498_ /*24189*/;
assign _496_ = _201_ ^ _498_ /*24192*/;
assign _497_ = _489_ & _496_ /*24190*/;
assign _426_ = _489_ ^ _496_ /*24191*/;
assign _494_ = _495_ | _497_ /*24188*/;
assign _503_ = ~D[10] /*24187*/;
assign _500_ = _202_ & _503_ /*24183*/;
assign _501_ = _202_ ^ _503_ /*24186*/;
assign _502_ = _494_ & _501_ /*24184*/;
assign _427_ = _494_ ^ _501_ /*24185*/;
assign _499_ = _500_ | _502_ /*24182*/;
assign _508_ = ~D[11] /*24181*/;
assign _505_ = _203_ & _508_ /*24177*/;
assign _506_ = _203_ ^ _508_ /*24180*/;
assign _507_ = _499_ & _506_ /*24178*/;
assign _428_ = _499_ ^ _506_ /*24179*/;
assign _504_ = _505_ | _507_ /*24176*/;
assign _513_ = ~D[12] /*24175*/;
assign _510_ = _204_ & _513_ /*24171*/;
assign _511_ = _204_ ^ _513_ /*24174*/;
assign _512_ = _504_ & _511_ /*24172*/;
assign _429_ = _504_ ^ _511_ /*24173*/;
assign _509_ = _510_ | _512_ /*24170*/;
assign _518_ = ~D[13] /*24169*/;
assign _515_ = _205_ & _518_ /*24165*/;
assign _516_ = _205_ ^ _518_ /*24168*/;
assign _517_ = _509_ & _516_ /*24166*/;
assign _430_ = _509_ ^ _516_ /*24167*/;
assign _514_ = _515_ | _517_ /*24164*/;
assign _523_ = ~D[14] /*24163*/;
assign _520_ = _206_ & _523_ /*24159*/;
assign _521_ = _206_ ^ _523_ /*24162*/;
assign _522_ = _514_ & _521_ /*24160*/;
assign _431_ = _514_ ^ _521_ /*24161*/;
assign _519_ = _520_ | _522_ /*24158*/;
assign _528_ = ~D[15] /*24157*/;
assign _525_ = _207_ & _528_ /*24153*/;
assign _526_ = _207_ ^ _528_ /*24156*/;
assign _527_ = _519_ & _526_ /*24154*/;
assign _432_ = _519_ ^ _526_ /*24155*/;
assign _524_ = _525_ | _527_ /*24152*/;
assign _533_ = ~D[16] /*24151*/;
assign _530_ = _208_ & _533_ /*24147*/;
assign _531_ = _208_ ^ _533_ /*24150*/;
assign _532_ = _524_ & _531_ /*24148*/;
assign _433_ = _524_ ^ _531_ /*24149*/;
assign _529_ = _530_ | _532_ /*24146*/;
assign _538_ = ~D[17] /*24145*/;
assign _535_ = _209_ & _538_ /*24141*/;
assign _536_ = _209_ ^ _538_ /*24144*/;
assign _537_ = _529_ & _536_ /*24142*/;
assign _434_ = _529_ ^ _536_ /*24143*/;
assign _534_ = _535_ | _537_ /*24140*/;
assign _543_ = ~D[18] /*24139*/;
assign _540_ = _210_ & _543_ /*24135*/;
assign _541_ = _210_ ^ _543_ /*24138*/;
assign _542_ = _534_ & _541_ /*24136*/;
assign _435_ = _534_ ^ _541_ /*24137*/;
assign _539_ = _540_ | _542_ /*24134*/;
assign _548_ = ~D[19] /*24133*/;
assign _545_ = _211_ & _548_ /*24129*/;
assign _546_ = _211_ ^ _548_ /*24132*/;
assign _547_ = _539_ & _546_ /*24130*/;
assign _436_ = _539_ ^ _546_ /*24131*/;
assign _544_ = _545_ | _547_ /*24128*/;
assign _553_ = ~D[20] /*24127*/;
assign _550_ = _212_ & _553_ /*24123*/;
assign _551_ = _212_ ^ _553_ /*24126*/;
assign _552_ = _544_ & _551_ /*24124*/;
assign _437_ = _544_ ^ _551_ /*24125*/;
assign _549_ = _550_ | _552_ /*24122*/;
assign _558_ = ~D[21] /*24121*/;
assign _555_ = _213_ & _558_ /*24117*/;
assign _556_ = _213_ ^ _558_ /*24120*/;
assign _557_ = _549_ & _556_ /*24118*/;
assign _438_ = _549_ ^ _556_ /*24119*/;
assign _554_ = _555_ | _557_ /*24116*/;
assign _563_ = ~D[22] /*24115*/;
assign _560_ = _214_ & _563_ /*24111*/;
assign _561_ = _214_ ^ _563_ /*24114*/;
assign _562_ = _554_ & _561_ /*24112*/;
assign _439_ = _554_ ^ _561_ /*24113*/;
assign _559_ = _560_ | _562_ /*24110*/;
assign _568_ = ~D[23] /*24109*/;
assign _565_ = _215_ & _568_ /*24105*/;
assign _566_ = _215_ ^ _568_ /*24108*/;
assign _567_ = _559_ & _566_ /*24106*/;
assign _440_ = _559_ ^ _566_ /*24107*/;
assign _564_ = _565_ | _567_ /*24104*/;
assign _573_ = ~D[24] /*24103*/;
assign _570_ = _216_ & _573_ /*24099*/;
assign _571_ = _216_ ^ _573_ /*24102*/;
assign _572_ = _564_ & _571_ /*24100*/;
assign _441_ = _564_ ^ _571_ /*24101*/;
assign _569_ = _570_ | _572_ /*24098*/;
assign _578_ = ~D[25] /*24097*/;
assign _575_ = _217_ & _578_ /*24093*/;
assign _576_ = _217_ ^ _578_ /*24096*/;
assign _577_ = _569_ & _576_ /*24094*/;
assign _442_ = _569_ ^ _576_ /*24095*/;
assign _574_ = _575_ | _577_ /*24092*/;
assign _583_ = ~D[26] /*24091*/;
assign _580_ = _218_ & _583_ /*24087*/;
assign _581_ = _218_ ^ _583_ /*24090*/;
assign _582_ = _574_ & _581_ /*24088*/;
assign _443_ = _574_ ^ _581_ /*24089*/;
assign _579_ = _580_ | _582_ /*24086*/;
assign _588_ = ~D[27] /*24085*/;
assign _585_ = _219_ & _588_ /*24081*/;
assign _586_ = _219_ ^ _588_ /*24084*/;
assign _587_ = _579_ & _586_ /*24082*/;
assign _444_ = _579_ ^ _586_ /*24083*/;
assign _584_ = _585_ | _587_ /*24080*/;
assign _593_ = ~D[28] /*24079*/;
assign _590_ = _220_ & _593_ /*24075*/;
assign _591_ = _220_ ^ _593_ /*24078*/;
assign _592_ = _584_ & _591_ /*24076*/;
assign _445_ = _584_ ^ _591_ /*24077*/;
assign _589_ = _590_ | _592_ /*24074*/;
assign _598_ = ~D[29] /*24073*/;
assign _595_ = _221_ & _598_ /*24069*/;
assign _596_ = _221_ ^ _598_ /*24072*/;
assign _597_ = _589_ & _596_ /*24070*/;
assign _446_ = _589_ ^ _596_ /*24071*/;
assign _594_ = _595_ | _597_ /*24068*/;
assign _603_ = ~D[30] /*24067*/;
assign _600_ = _222_ & _603_ /*24063*/;
assign _601_ = _222_ ^ _603_ /*24066*/;
assign _602_ = _594_ & _601_ /*24064*/;
assign _447_ = _594_ ^ _601_ /*24065*/;
assign _599_ = _600_ | _602_ /*24062*/;
assign _604_ = _223_ & oneWire /*24057*/;
assign _605_ = _223_ ^ oneWire /*24060*/;
assign _606_ = _599_ & _605_ /*24058*/;
assign _448_ = _599_ ^ _605_ /*24059*/;
assign Q[30] = _604_ | _606_ /*24056*/;
assign _675_ = ~Q[30] /*23863*/;
assign _674_ = _675_ & D[0] /*23862*/;
assign _677_ = _417_ & _674_ /*23857*/;
assign _678_ = _417_ ^ _674_ /*23860*/;
assign _679_ = zeroWire & _678_ /*23858*/;
assign _641_ = zeroWire ^ _678_ /*23859*/;
assign _676_ = _677_ | _679_ /*23856*/;
assign _681_ = ~Q[30] /*23855*/;
assign _680_ = _681_ & D[1] /*23854*/;
assign _683_ = _418_ & _680_ /*23849*/;
assign _684_ = _418_ ^ _680_ /*23852*/;
assign _685_ = _676_ & _684_ /*23850*/;
assign _642_ = _676_ ^ _684_ /*23851*/;
assign _682_ = _683_ | _685_ /*23848*/;
assign _687_ = ~Q[30] /*23847*/;
assign _686_ = _687_ & D[2] /*23846*/;
assign _689_ = _419_ & _686_ /*23841*/;
assign _690_ = _419_ ^ _686_ /*23844*/;
assign _691_ = _682_ & _690_ /*23842*/;
assign _643_ = _682_ ^ _690_ /*23843*/;
assign _688_ = _689_ | _691_ /*23840*/;
assign _693_ = ~Q[30] /*23839*/;
assign _692_ = _693_ & D[3] /*23838*/;
assign _695_ = _420_ & _692_ /*23833*/;
assign _696_ = _420_ ^ _692_ /*23836*/;
assign _697_ = _688_ & _696_ /*23834*/;
assign _644_ = _688_ ^ _696_ /*23835*/;
assign _694_ = _695_ | _697_ /*23832*/;
assign _699_ = ~Q[30] /*23831*/;
assign _698_ = _699_ & D[4] /*23830*/;
assign _701_ = _421_ & _698_ /*23825*/;
assign _702_ = _421_ ^ _698_ /*23828*/;
assign _703_ = _694_ & _702_ /*23826*/;
assign _645_ = _694_ ^ _702_ /*23827*/;
assign _700_ = _701_ | _703_ /*23824*/;
assign _705_ = ~Q[30] /*23823*/;
assign _704_ = _705_ & D[5] /*23822*/;
assign _707_ = _422_ & _704_ /*23817*/;
assign _708_ = _422_ ^ _704_ /*23820*/;
assign _709_ = _700_ & _708_ /*23818*/;
assign _646_ = _700_ ^ _708_ /*23819*/;
assign _706_ = _707_ | _709_ /*23816*/;
assign _711_ = ~Q[30] /*23815*/;
assign _710_ = _711_ & D[6] /*23814*/;
assign _713_ = _423_ & _710_ /*23809*/;
assign _714_ = _423_ ^ _710_ /*23812*/;
assign _715_ = _706_ & _714_ /*23810*/;
assign _647_ = _706_ ^ _714_ /*23811*/;
assign _712_ = _713_ | _715_ /*23808*/;
assign _717_ = ~Q[30] /*23807*/;
assign _716_ = _717_ & D[7] /*23806*/;
assign _719_ = _424_ & _716_ /*23801*/;
assign _720_ = _424_ ^ _716_ /*23804*/;
assign _721_ = _712_ & _720_ /*23802*/;
assign _648_ = _712_ ^ _720_ /*23803*/;
assign _718_ = _719_ | _721_ /*23800*/;
assign _723_ = ~Q[30] /*23799*/;
assign _722_ = _723_ & D[8] /*23798*/;
assign _725_ = _425_ & _722_ /*23793*/;
assign _726_ = _425_ ^ _722_ /*23796*/;
assign _727_ = _718_ & _726_ /*23794*/;
assign _649_ = _718_ ^ _726_ /*23795*/;
assign _724_ = _725_ | _727_ /*23792*/;
assign _729_ = ~Q[30] /*23791*/;
assign _728_ = _729_ & D[9] /*23790*/;
assign _731_ = _426_ & _728_ /*23785*/;
assign _732_ = _426_ ^ _728_ /*23788*/;
assign _733_ = _724_ & _732_ /*23786*/;
assign _650_ = _724_ ^ _732_ /*23787*/;
assign _730_ = _731_ | _733_ /*23784*/;
assign _735_ = ~Q[30] /*23783*/;
assign _734_ = _735_ & D[10] /*23782*/;
assign _737_ = _427_ & _734_ /*23777*/;
assign _738_ = _427_ ^ _734_ /*23780*/;
assign _739_ = _730_ & _738_ /*23778*/;
assign _651_ = _730_ ^ _738_ /*23779*/;
assign _736_ = _737_ | _739_ /*23776*/;
assign _741_ = ~Q[30] /*23775*/;
assign _740_ = _741_ & D[11] /*23774*/;
assign _743_ = _428_ & _740_ /*23769*/;
assign _744_ = _428_ ^ _740_ /*23772*/;
assign _745_ = _736_ & _744_ /*23770*/;
assign _652_ = _736_ ^ _744_ /*23771*/;
assign _742_ = _743_ | _745_ /*23768*/;
assign _747_ = ~Q[30] /*23767*/;
assign _746_ = _747_ & D[12] /*23766*/;
assign _749_ = _429_ & _746_ /*23761*/;
assign _750_ = _429_ ^ _746_ /*23764*/;
assign _751_ = _742_ & _750_ /*23762*/;
assign _653_ = _742_ ^ _750_ /*23763*/;
assign _748_ = _749_ | _751_ /*23760*/;
assign _753_ = ~Q[30] /*23759*/;
assign _752_ = _753_ & D[13] /*23758*/;
assign _755_ = _430_ & _752_ /*23753*/;
assign _756_ = _430_ ^ _752_ /*23756*/;
assign _757_ = _748_ & _756_ /*23754*/;
assign _654_ = _748_ ^ _756_ /*23755*/;
assign _754_ = _755_ | _757_ /*23752*/;
assign _759_ = ~Q[30] /*23751*/;
assign _758_ = _759_ & D[14] /*23750*/;
assign _761_ = _431_ & _758_ /*23745*/;
assign _762_ = _431_ ^ _758_ /*23748*/;
assign _763_ = _754_ & _762_ /*23746*/;
assign _655_ = _754_ ^ _762_ /*23747*/;
assign _760_ = _761_ | _763_ /*23744*/;
assign _765_ = ~Q[30] /*23743*/;
assign _764_ = _765_ & D[15] /*23742*/;
assign _767_ = _432_ & _764_ /*23737*/;
assign _768_ = _432_ ^ _764_ /*23740*/;
assign _769_ = _760_ & _768_ /*23738*/;
assign _656_ = _760_ ^ _768_ /*23739*/;
assign _766_ = _767_ | _769_ /*23736*/;
assign _771_ = ~Q[30] /*23735*/;
assign _770_ = _771_ & D[16] /*23734*/;
assign _773_ = _433_ & _770_ /*23729*/;
assign _774_ = _433_ ^ _770_ /*23732*/;
assign _775_ = _766_ & _774_ /*23730*/;
assign _657_ = _766_ ^ _774_ /*23731*/;
assign _772_ = _773_ | _775_ /*23728*/;
assign _777_ = ~Q[30] /*23727*/;
assign _776_ = _777_ & D[17] /*23726*/;
assign _779_ = _434_ & _776_ /*23721*/;
assign _780_ = _434_ ^ _776_ /*23724*/;
assign _781_ = _772_ & _780_ /*23722*/;
assign _658_ = _772_ ^ _780_ /*23723*/;
assign _778_ = _779_ | _781_ /*23720*/;
assign _783_ = ~Q[30] /*23719*/;
assign _782_ = _783_ & D[18] /*23718*/;
assign _785_ = _435_ & _782_ /*23713*/;
assign _786_ = _435_ ^ _782_ /*23716*/;
assign _787_ = _778_ & _786_ /*23714*/;
assign _659_ = _778_ ^ _786_ /*23715*/;
assign _784_ = _785_ | _787_ /*23712*/;
assign _789_ = ~Q[30] /*23711*/;
assign _788_ = _789_ & D[19] /*23710*/;
assign _791_ = _436_ & _788_ /*23705*/;
assign _792_ = _436_ ^ _788_ /*23708*/;
assign _793_ = _784_ & _792_ /*23706*/;
assign _660_ = _784_ ^ _792_ /*23707*/;
assign _790_ = _791_ | _793_ /*23704*/;
assign _795_ = ~Q[30] /*23703*/;
assign _794_ = _795_ & D[20] /*23702*/;
assign _797_ = _437_ & _794_ /*23697*/;
assign _798_ = _437_ ^ _794_ /*23700*/;
assign _799_ = _790_ & _798_ /*23698*/;
assign _661_ = _790_ ^ _798_ /*23699*/;
assign _796_ = _797_ | _799_ /*23696*/;
assign _801_ = ~Q[30] /*23695*/;
assign _800_ = _801_ & D[21] /*23694*/;
assign _803_ = _438_ & _800_ /*23689*/;
assign _804_ = _438_ ^ _800_ /*23692*/;
assign _805_ = _796_ & _804_ /*23690*/;
assign _662_ = _796_ ^ _804_ /*23691*/;
assign _802_ = _803_ | _805_ /*23688*/;
assign _807_ = ~Q[30] /*23687*/;
assign _806_ = _807_ & D[22] /*23686*/;
assign _809_ = _439_ & _806_ /*23681*/;
assign _810_ = _439_ ^ _806_ /*23684*/;
assign _811_ = _802_ & _810_ /*23682*/;
assign _663_ = _802_ ^ _810_ /*23683*/;
assign _808_ = _809_ | _811_ /*23680*/;
assign _813_ = ~Q[30] /*23679*/;
assign _812_ = _813_ & D[23] /*23678*/;
assign _815_ = _440_ & _812_ /*23673*/;
assign _816_ = _440_ ^ _812_ /*23676*/;
assign _817_ = _808_ & _816_ /*23674*/;
assign _664_ = _808_ ^ _816_ /*23675*/;
assign _814_ = _815_ | _817_ /*23672*/;
assign _819_ = ~Q[30] /*23671*/;
assign _818_ = _819_ & D[24] /*23670*/;
assign _821_ = _441_ & _818_ /*23665*/;
assign _822_ = _441_ ^ _818_ /*23668*/;
assign _823_ = _814_ & _822_ /*23666*/;
assign _665_ = _814_ ^ _822_ /*23667*/;
assign _820_ = _821_ | _823_ /*23664*/;
assign _825_ = ~Q[30] /*23663*/;
assign _824_ = _825_ & D[25] /*23662*/;
assign _827_ = _442_ & _824_ /*23657*/;
assign _828_ = _442_ ^ _824_ /*23660*/;
assign _829_ = _820_ & _828_ /*23658*/;
assign _666_ = _820_ ^ _828_ /*23659*/;
assign _826_ = _827_ | _829_ /*23656*/;
assign _831_ = ~Q[30] /*23655*/;
assign _830_ = _831_ & D[26] /*23654*/;
assign _833_ = _443_ & _830_ /*23649*/;
assign _834_ = _443_ ^ _830_ /*23652*/;
assign _835_ = _826_ & _834_ /*23650*/;
assign _667_ = _826_ ^ _834_ /*23651*/;
assign _832_ = _833_ | _835_ /*23648*/;
assign _837_ = ~Q[30] /*23647*/;
assign _836_ = _837_ & D[27] /*23646*/;
assign _839_ = _444_ & _836_ /*23641*/;
assign _840_ = _444_ ^ _836_ /*23644*/;
assign _841_ = _832_ & _840_ /*23642*/;
assign _668_ = _832_ ^ _840_ /*23643*/;
assign _838_ = _839_ | _841_ /*23640*/;
assign _843_ = ~Q[30] /*23639*/;
assign _842_ = _843_ & D[28] /*23638*/;
assign _845_ = _445_ & _842_ /*23633*/;
assign _846_ = _445_ ^ _842_ /*23636*/;
assign _847_ = _838_ & _846_ /*23634*/;
assign _669_ = _838_ ^ _846_ /*23635*/;
assign _844_ = _845_ | _847_ /*23632*/;
assign _849_ = ~Q[30] /*23631*/;
assign _848_ = _849_ & D[29] /*23630*/;
assign _851_ = _446_ & _848_ /*23625*/;
assign _852_ = _446_ ^ _848_ /*23628*/;
assign _853_ = _844_ & _852_ /*23626*/;
assign _670_ = _844_ ^ _852_ /*23627*/;
assign _850_ = _851_ | _853_ /*23624*/;
assign _855_ = ~Q[30] /*23623*/;
assign _854_ = _855_ & D[30] /*23622*/;
assign _857_ = _447_ & _854_ /*23617*/;
assign _858_ = _447_ ^ _854_ /*23620*/;
assign _859_ = _850_ & _858_ /*23618*/;
assign _671_ = _850_ ^ _858_ /*23619*/;
assign _856_ = _857_ | _859_ /*23616*/;
assign _861_ = ~Q[30] /*23615*/;
assign _860_ = _861_ & zeroWire /*23614*/;
assign _862_ = _448_ ^ _860_ /*23612*/;
assign _672_ = _862_ ^ _856_ /*23611*/;
assign _901_ = ~D[0] /*23485*/;
assign _898_ = R_0[29] & _901_ /*23481*/;
assign _899_ = R_0[29] ^ _901_ /*23484*/;
assign _900_ = oneWire & _899_ /*23482*/;
assign _865_ = oneWire ^ _899_ /*23483*/;
assign _897_ = _898_ | _900_ /*23480*/;
assign _906_ = ~D[1] /*23479*/;
assign _903_ = _641_ & _906_ /*23475*/;
assign _904_ = _641_ ^ _906_ /*23478*/;
assign _905_ = _897_ & _904_ /*23476*/;
assign _866_ = _897_ ^ _904_ /*23477*/;
assign _902_ = _903_ | _905_ /*23474*/;
assign _911_ = ~D[2] /*23473*/;
assign _908_ = _642_ & _911_ /*23469*/;
assign _909_ = _642_ ^ _911_ /*23472*/;
assign _910_ = _902_ & _909_ /*23470*/;
assign _867_ = _902_ ^ _909_ /*23471*/;
assign _907_ = _908_ | _910_ /*23468*/;
assign _916_ = ~D[3] /*23467*/;
assign _913_ = _643_ & _916_ /*23463*/;
assign _914_ = _643_ ^ _916_ /*23466*/;
assign _915_ = _907_ & _914_ /*23464*/;
assign _868_ = _907_ ^ _914_ /*23465*/;
assign _912_ = _913_ | _915_ /*23462*/;
assign _921_ = ~D[4] /*23461*/;
assign _918_ = _644_ & _921_ /*23457*/;
assign _919_ = _644_ ^ _921_ /*23460*/;
assign _920_ = _912_ & _919_ /*23458*/;
assign _869_ = _912_ ^ _919_ /*23459*/;
assign _917_ = _918_ | _920_ /*23456*/;
assign _926_ = ~D[5] /*23455*/;
assign _923_ = _645_ & _926_ /*23451*/;
assign _924_ = _645_ ^ _926_ /*23454*/;
assign _925_ = _917_ & _924_ /*23452*/;
assign _870_ = _917_ ^ _924_ /*23453*/;
assign _922_ = _923_ | _925_ /*23450*/;
assign _931_ = ~D[6] /*23449*/;
assign _928_ = _646_ & _931_ /*23445*/;
assign _929_ = _646_ ^ _931_ /*23448*/;
assign _930_ = _922_ & _929_ /*23446*/;
assign _871_ = _922_ ^ _929_ /*23447*/;
assign _927_ = _928_ | _930_ /*23444*/;
assign _936_ = ~D[7] /*23443*/;
assign _933_ = _647_ & _936_ /*23439*/;
assign _934_ = _647_ ^ _936_ /*23442*/;
assign _935_ = _927_ & _934_ /*23440*/;
assign _872_ = _927_ ^ _934_ /*23441*/;
assign _932_ = _933_ | _935_ /*23438*/;
assign _941_ = ~D[8] /*23437*/;
assign _938_ = _648_ & _941_ /*23433*/;
assign _939_ = _648_ ^ _941_ /*23436*/;
assign _940_ = _932_ & _939_ /*23434*/;
assign _873_ = _932_ ^ _939_ /*23435*/;
assign _937_ = _938_ | _940_ /*23432*/;
assign _946_ = ~D[9] /*23431*/;
assign _943_ = _649_ & _946_ /*23427*/;
assign _944_ = _649_ ^ _946_ /*23430*/;
assign _945_ = _937_ & _944_ /*23428*/;
assign _874_ = _937_ ^ _944_ /*23429*/;
assign _942_ = _943_ | _945_ /*23426*/;
assign _951_ = ~D[10] /*23425*/;
assign _948_ = _650_ & _951_ /*23421*/;
assign _949_ = _650_ ^ _951_ /*23424*/;
assign _950_ = _942_ & _949_ /*23422*/;
assign _875_ = _942_ ^ _949_ /*23423*/;
assign _947_ = _948_ | _950_ /*23420*/;
assign _956_ = ~D[11] /*23419*/;
assign _953_ = _651_ & _956_ /*23415*/;
assign _954_ = _651_ ^ _956_ /*23418*/;
assign _955_ = _947_ & _954_ /*23416*/;
assign _876_ = _947_ ^ _954_ /*23417*/;
assign _952_ = _953_ | _955_ /*23414*/;
assign _961_ = ~D[12] /*23413*/;
assign _958_ = _652_ & _961_ /*23409*/;
assign _959_ = _652_ ^ _961_ /*23412*/;
assign _960_ = _952_ & _959_ /*23410*/;
assign _877_ = _952_ ^ _959_ /*23411*/;
assign _957_ = _958_ | _960_ /*23408*/;
assign _966_ = ~D[13] /*23407*/;
assign _963_ = _653_ & _966_ /*23403*/;
assign _964_ = _653_ ^ _966_ /*23406*/;
assign _965_ = _957_ & _964_ /*23404*/;
assign _878_ = _957_ ^ _964_ /*23405*/;
assign _962_ = _963_ | _965_ /*23402*/;
assign _971_ = ~D[14] /*23401*/;
assign _968_ = _654_ & _971_ /*23397*/;
assign _969_ = _654_ ^ _971_ /*23400*/;
assign _970_ = _962_ & _969_ /*23398*/;
assign _879_ = _962_ ^ _969_ /*23399*/;
assign _967_ = _968_ | _970_ /*23396*/;
assign _976_ = ~D[15] /*23395*/;
assign _973_ = _655_ & _976_ /*23391*/;
assign _974_ = _655_ ^ _976_ /*23394*/;
assign _975_ = _967_ & _974_ /*23392*/;
assign _880_ = _967_ ^ _974_ /*23393*/;
assign _972_ = _973_ | _975_ /*23390*/;
assign _981_ = ~D[16] /*23389*/;
assign _978_ = _656_ & _981_ /*23385*/;
assign _979_ = _656_ ^ _981_ /*23388*/;
assign _980_ = _972_ & _979_ /*23386*/;
assign _881_ = _972_ ^ _979_ /*23387*/;
assign _977_ = _978_ | _980_ /*23384*/;
assign _986_ = ~D[17] /*23383*/;
assign _983_ = _657_ & _986_ /*23379*/;
assign _984_ = _657_ ^ _986_ /*23382*/;
assign _985_ = _977_ & _984_ /*23380*/;
assign _882_ = _977_ ^ _984_ /*23381*/;
assign _982_ = _983_ | _985_ /*23378*/;
assign _991_ = ~D[18] /*23377*/;
assign _988_ = _658_ & _991_ /*23373*/;
assign _989_ = _658_ ^ _991_ /*23376*/;
assign _990_ = _982_ & _989_ /*23374*/;
assign _883_ = _982_ ^ _989_ /*23375*/;
assign _987_ = _988_ | _990_ /*23372*/;
assign _996_ = ~D[19] /*23371*/;
assign _993_ = _659_ & _996_ /*23367*/;
assign _994_ = _659_ ^ _996_ /*23370*/;
assign _995_ = _987_ & _994_ /*23368*/;
assign _884_ = _987_ ^ _994_ /*23369*/;
assign _992_ = _993_ | _995_ /*23366*/;
assign _1001_ = ~D[20] /*23365*/;
assign _998_ = _660_ & _1001_ /*23361*/;
assign _999_ = _660_ ^ _1001_ /*23364*/;
assign _1000_ = _992_ & _999_ /*23362*/;
assign _885_ = _992_ ^ _999_ /*23363*/;
assign _997_ = _998_ | _1000_ /*23360*/;
assign _1006_ = ~D[21] /*23359*/;
assign _1003_ = _661_ & _1006_ /*23355*/;
assign _1004_ = _661_ ^ _1006_ /*23358*/;
assign _1005_ = _997_ & _1004_ /*23356*/;
assign _886_ = _997_ ^ _1004_ /*23357*/;
assign _1002_ = _1003_ | _1005_ /*23354*/;
assign _1011_ = ~D[22] /*23353*/;
assign _1008_ = _662_ & _1011_ /*23349*/;
assign _1009_ = _662_ ^ _1011_ /*23352*/;
assign _1010_ = _1002_ & _1009_ /*23350*/;
assign _887_ = _1002_ ^ _1009_ /*23351*/;
assign _1007_ = _1008_ | _1010_ /*23348*/;
assign _1016_ = ~D[23] /*23347*/;
assign _1013_ = _663_ & _1016_ /*23343*/;
assign _1014_ = _663_ ^ _1016_ /*23346*/;
assign _1015_ = _1007_ & _1014_ /*23344*/;
assign _888_ = _1007_ ^ _1014_ /*23345*/;
assign _1012_ = _1013_ | _1015_ /*23342*/;
assign _1021_ = ~D[24] /*23341*/;
assign _1018_ = _664_ & _1021_ /*23337*/;
assign _1019_ = _664_ ^ _1021_ /*23340*/;
assign _1020_ = _1012_ & _1019_ /*23338*/;
assign _889_ = _1012_ ^ _1019_ /*23339*/;
assign _1017_ = _1018_ | _1020_ /*23336*/;
assign _1026_ = ~D[25] /*23335*/;
assign _1023_ = _665_ & _1026_ /*23331*/;
assign _1024_ = _665_ ^ _1026_ /*23334*/;
assign _1025_ = _1017_ & _1024_ /*23332*/;
assign _890_ = _1017_ ^ _1024_ /*23333*/;
assign _1022_ = _1023_ | _1025_ /*23330*/;
assign _1031_ = ~D[26] /*23329*/;
assign _1028_ = _666_ & _1031_ /*23325*/;
assign _1029_ = _666_ ^ _1031_ /*23328*/;
assign _1030_ = _1022_ & _1029_ /*23326*/;
assign _891_ = _1022_ ^ _1029_ /*23327*/;
assign _1027_ = _1028_ | _1030_ /*23324*/;
assign _1036_ = ~D[27] /*23323*/;
assign _1033_ = _667_ & _1036_ /*23319*/;
assign _1034_ = _667_ ^ _1036_ /*23322*/;
assign _1035_ = _1027_ & _1034_ /*23320*/;
assign _892_ = _1027_ ^ _1034_ /*23321*/;
assign _1032_ = _1033_ | _1035_ /*23318*/;
assign _1041_ = ~D[28] /*23317*/;
assign _1038_ = _668_ & _1041_ /*23313*/;
assign _1039_ = _668_ ^ _1041_ /*23316*/;
assign _1040_ = _1032_ & _1039_ /*23314*/;
assign _893_ = _1032_ ^ _1039_ /*23315*/;
assign _1037_ = _1038_ | _1040_ /*23312*/;
assign _1046_ = ~D[29] /*23311*/;
assign _1043_ = _669_ & _1046_ /*23307*/;
assign _1044_ = _669_ ^ _1046_ /*23310*/;
assign _1045_ = _1037_ & _1044_ /*23308*/;
assign _894_ = _1037_ ^ _1044_ /*23309*/;
assign _1042_ = _1043_ | _1045_ /*23306*/;
assign _1051_ = ~D[30] /*23305*/;
assign _1048_ = _670_ & _1051_ /*23301*/;
assign _1049_ = _670_ ^ _1051_ /*23304*/;
assign _1050_ = _1042_ & _1049_ /*23302*/;
assign _895_ = _1042_ ^ _1049_ /*23303*/;
assign _1047_ = _1048_ | _1050_ /*23300*/;
assign _1052_ = _671_ & oneWire /*23295*/;
assign _1053_ = _671_ ^ oneWire /*23298*/;
assign _1054_ = _1047_ & _1053_ /*23296*/;
assign _896_ = _1047_ ^ _1053_ /*23297*/;
assign Q[29] = _1052_ | _1054_ /*23294*/;
assign _1123_ = ~Q[29] /*23101*/;
assign _1122_ = _1123_ & D[0] /*23100*/;
assign _1125_ = _865_ & _1122_ /*23095*/;
assign _1126_ = _865_ ^ _1122_ /*23098*/;
assign _1127_ = zeroWire & _1126_ /*23096*/;
assign _1089_ = zeroWire ^ _1126_ /*23097*/;
assign _1124_ = _1125_ | _1127_ /*23094*/;
assign _1129_ = ~Q[29] /*23093*/;
assign _1128_ = _1129_ & D[1] /*23092*/;
assign _1131_ = _866_ & _1128_ /*23087*/;
assign _1132_ = _866_ ^ _1128_ /*23090*/;
assign _1133_ = _1124_ & _1132_ /*23088*/;
assign _1090_ = _1124_ ^ _1132_ /*23089*/;
assign _1130_ = _1131_ | _1133_ /*23086*/;
assign _1135_ = ~Q[29] /*23085*/;
assign _1134_ = _1135_ & D[2] /*23084*/;
assign _1137_ = _867_ & _1134_ /*23079*/;
assign _1138_ = _867_ ^ _1134_ /*23082*/;
assign _1139_ = _1130_ & _1138_ /*23080*/;
assign _1091_ = _1130_ ^ _1138_ /*23081*/;
assign _1136_ = _1137_ | _1139_ /*23078*/;
assign _1141_ = ~Q[29] /*23077*/;
assign _1140_ = _1141_ & D[3] /*23076*/;
assign _1143_ = _868_ & _1140_ /*23071*/;
assign _1144_ = _868_ ^ _1140_ /*23074*/;
assign _1145_ = _1136_ & _1144_ /*23072*/;
assign _1092_ = _1136_ ^ _1144_ /*23073*/;
assign _1142_ = _1143_ | _1145_ /*23070*/;
assign _1147_ = ~Q[29] /*23069*/;
assign _1146_ = _1147_ & D[4] /*23068*/;
assign _1149_ = _869_ & _1146_ /*23063*/;
assign _1150_ = _869_ ^ _1146_ /*23066*/;
assign _1151_ = _1142_ & _1150_ /*23064*/;
assign _1093_ = _1142_ ^ _1150_ /*23065*/;
assign _1148_ = _1149_ | _1151_ /*23062*/;
assign _1153_ = ~Q[29] /*23061*/;
assign _1152_ = _1153_ & D[5] /*23060*/;
assign _1155_ = _870_ & _1152_ /*23055*/;
assign _1156_ = _870_ ^ _1152_ /*23058*/;
assign _1157_ = _1148_ & _1156_ /*23056*/;
assign _1094_ = _1148_ ^ _1156_ /*23057*/;
assign _1154_ = _1155_ | _1157_ /*23054*/;
assign _1159_ = ~Q[29] /*23053*/;
assign _1158_ = _1159_ & D[6] /*23052*/;
assign _1161_ = _871_ & _1158_ /*23047*/;
assign _1162_ = _871_ ^ _1158_ /*23050*/;
assign _1163_ = _1154_ & _1162_ /*23048*/;
assign _1095_ = _1154_ ^ _1162_ /*23049*/;
assign _1160_ = _1161_ | _1163_ /*23046*/;
assign _1165_ = ~Q[29] /*23045*/;
assign _1164_ = _1165_ & D[7] /*23044*/;
assign _1167_ = _872_ & _1164_ /*23039*/;
assign _1168_ = _872_ ^ _1164_ /*23042*/;
assign _1169_ = _1160_ & _1168_ /*23040*/;
assign _1096_ = _1160_ ^ _1168_ /*23041*/;
assign _1166_ = _1167_ | _1169_ /*23038*/;
assign _1171_ = ~Q[29] /*23037*/;
assign _1170_ = _1171_ & D[8] /*23036*/;
assign _1173_ = _873_ & _1170_ /*23031*/;
assign _1174_ = _873_ ^ _1170_ /*23034*/;
assign _1175_ = _1166_ & _1174_ /*23032*/;
assign _1097_ = _1166_ ^ _1174_ /*23033*/;
assign _1172_ = _1173_ | _1175_ /*23030*/;
assign _1177_ = ~Q[29] /*23029*/;
assign _1176_ = _1177_ & D[9] /*23028*/;
assign _1179_ = _874_ & _1176_ /*23023*/;
assign _1180_ = _874_ ^ _1176_ /*23026*/;
assign _1181_ = _1172_ & _1180_ /*23024*/;
assign _1098_ = _1172_ ^ _1180_ /*23025*/;
assign _1178_ = _1179_ | _1181_ /*23022*/;
assign _1183_ = ~Q[29] /*23021*/;
assign _1182_ = _1183_ & D[10] /*23020*/;
assign _1185_ = _875_ & _1182_ /*23015*/;
assign _1186_ = _875_ ^ _1182_ /*23018*/;
assign _1187_ = _1178_ & _1186_ /*23016*/;
assign _1099_ = _1178_ ^ _1186_ /*23017*/;
assign _1184_ = _1185_ | _1187_ /*23014*/;
assign _1189_ = ~Q[29] /*23013*/;
assign _1188_ = _1189_ & D[11] /*23012*/;
assign _1191_ = _876_ & _1188_ /*23007*/;
assign _1192_ = _876_ ^ _1188_ /*23010*/;
assign _1193_ = _1184_ & _1192_ /*23008*/;
assign _1100_ = _1184_ ^ _1192_ /*23009*/;
assign _1190_ = _1191_ | _1193_ /*23006*/;
assign _1195_ = ~Q[29] /*23005*/;
assign _1194_ = _1195_ & D[12] /*23004*/;
assign _1197_ = _877_ & _1194_ /*22999*/;
assign _1198_ = _877_ ^ _1194_ /*23002*/;
assign _1199_ = _1190_ & _1198_ /*23000*/;
assign _1101_ = _1190_ ^ _1198_ /*23001*/;
assign _1196_ = _1197_ | _1199_ /*22998*/;
assign _1201_ = ~Q[29] /*22997*/;
assign _1200_ = _1201_ & D[13] /*22996*/;
assign _1203_ = _878_ & _1200_ /*22991*/;
assign _1204_ = _878_ ^ _1200_ /*22994*/;
assign _1205_ = _1196_ & _1204_ /*22992*/;
assign _1102_ = _1196_ ^ _1204_ /*22993*/;
assign _1202_ = _1203_ | _1205_ /*22990*/;
assign _1207_ = ~Q[29] /*22989*/;
assign _1206_ = _1207_ & D[14] /*22988*/;
assign _1209_ = _879_ & _1206_ /*22983*/;
assign _1210_ = _879_ ^ _1206_ /*22986*/;
assign _1211_ = _1202_ & _1210_ /*22984*/;
assign _1103_ = _1202_ ^ _1210_ /*22985*/;
assign _1208_ = _1209_ | _1211_ /*22982*/;
assign _1213_ = ~Q[29] /*22981*/;
assign _1212_ = _1213_ & D[15] /*22980*/;
assign _1215_ = _880_ & _1212_ /*22975*/;
assign _1216_ = _880_ ^ _1212_ /*22978*/;
assign _1217_ = _1208_ & _1216_ /*22976*/;
assign _1104_ = _1208_ ^ _1216_ /*22977*/;
assign _1214_ = _1215_ | _1217_ /*22974*/;
assign _1219_ = ~Q[29] /*22973*/;
assign _1218_ = _1219_ & D[16] /*22972*/;
assign _1221_ = _881_ & _1218_ /*22967*/;
assign _1222_ = _881_ ^ _1218_ /*22970*/;
assign _1223_ = _1214_ & _1222_ /*22968*/;
assign _1105_ = _1214_ ^ _1222_ /*22969*/;
assign _1220_ = _1221_ | _1223_ /*22966*/;
assign _1225_ = ~Q[29] /*22965*/;
assign _1224_ = _1225_ & D[17] /*22964*/;
assign _1227_ = _882_ & _1224_ /*22959*/;
assign _1228_ = _882_ ^ _1224_ /*22962*/;
assign _1229_ = _1220_ & _1228_ /*22960*/;
assign _1106_ = _1220_ ^ _1228_ /*22961*/;
assign _1226_ = _1227_ | _1229_ /*22958*/;
assign _1231_ = ~Q[29] /*22957*/;
assign _1230_ = _1231_ & D[18] /*22956*/;
assign _1233_ = _883_ & _1230_ /*22951*/;
assign _1234_ = _883_ ^ _1230_ /*22954*/;
assign _1235_ = _1226_ & _1234_ /*22952*/;
assign _1107_ = _1226_ ^ _1234_ /*22953*/;
assign _1232_ = _1233_ | _1235_ /*22950*/;
assign _1237_ = ~Q[29] /*22949*/;
assign _1236_ = _1237_ & D[19] /*22948*/;
assign _1239_ = _884_ & _1236_ /*22943*/;
assign _1240_ = _884_ ^ _1236_ /*22946*/;
assign _1241_ = _1232_ & _1240_ /*22944*/;
assign _1108_ = _1232_ ^ _1240_ /*22945*/;
assign _1238_ = _1239_ | _1241_ /*22942*/;
assign _1243_ = ~Q[29] /*22941*/;
assign _1242_ = _1243_ & D[20] /*22940*/;
assign _1245_ = _885_ & _1242_ /*22935*/;
assign _1246_ = _885_ ^ _1242_ /*22938*/;
assign _1247_ = _1238_ & _1246_ /*22936*/;
assign _1109_ = _1238_ ^ _1246_ /*22937*/;
assign _1244_ = _1245_ | _1247_ /*22934*/;
assign _1249_ = ~Q[29] /*22933*/;
assign _1248_ = _1249_ & D[21] /*22932*/;
assign _1251_ = _886_ & _1248_ /*22927*/;
assign _1252_ = _886_ ^ _1248_ /*22930*/;
assign _1253_ = _1244_ & _1252_ /*22928*/;
assign _1110_ = _1244_ ^ _1252_ /*22929*/;
assign _1250_ = _1251_ | _1253_ /*22926*/;
assign _1255_ = ~Q[29] /*22925*/;
assign _1254_ = _1255_ & D[22] /*22924*/;
assign _1257_ = _887_ & _1254_ /*22919*/;
assign _1258_ = _887_ ^ _1254_ /*22922*/;
assign _1259_ = _1250_ & _1258_ /*22920*/;
assign _1111_ = _1250_ ^ _1258_ /*22921*/;
assign _1256_ = _1257_ | _1259_ /*22918*/;
assign _1261_ = ~Q[29] /*22917*/;
assign _1260_ = _1261_ & D[23] /*22916*/;
assign _1263_ = _888_ & _1260_ /*22911*/;
assign _1264_ = _888_ ^ _1260_ /*22914*/;
assign _1265_ = _1256_ & _1264_ /*22912*/;
assign _1112_ = _1256_ ^ _1264_ /*22913*/;
assign _1262_ = _1263_ | _1265_ /*22910*/;
assign _1267_ = ~Q[29] /*22909*/;
assign _1266_ = _1267_ & D[24] /*22908*/;
assign _1269_ = _889_ & _1266_ /*22903*/;
assign _1270_ = _889_ ^ _1266_ /*22906*/;
assign _1271_ = _1262_ & _1270_ /*22904*/;
assign _1113_ = _1262_ ^ _1270_ /*22905*/;
assign _1268_ = _1269_ | _1271_ /*22902*/;
assign _1273_ = ~Q[29] /*22901*/;
assign _1272_ = _1273_ & D[25] /*22900*/;
assign _1275_ = _890_ & _1272_ /*22895*/;
assign _1276_ = _890_ ^ _1272_ /*22898*/;
assign _1277_ = _1268_ & _1276_ /*22896*/;
assign _1114_ = _1268_ ^ _1276_ /*22897*/;
assign _1274_ = _1275_ | _1277_ /*22894*/;
assign _1279_ = ~Q[29] /*22893*/;
assign _1278_ = _1279_ & D[26] /*22892*/;
assign _1281_ = _891_ & _1278_ /*22887*/;
assign _1282_ = _891_ ^ _1278_ /*22890*/;
assign _1283_ = _1274_ & _1282_ /*22888*/;
assign _1115_ = _1274_ ^ _1282_ /*22889*/;
assign _1280_ = _1281_ | _1283_ /*22886*/;
assign _1285_ = ~Q[29] /*22885*/;
assign _1284_ = _1285_ & D[27] /*22884*/;
assign _1287_ = _892_ & _1284_ /*22879*/;
assign _1288_ = _892_ ^ _1284_ /*22882*/;
assign _1289_ = _1280_ & _1288_ /*22880*/;
assign _1116_ = _1280_ ^ _1288_ /*22881*/;
assign _1286_ = _1287_ | _1289_ /*22878*/;
assign _1291_ = ~Q[29] /*22877*/;
assign _1290_ = _1291_ & D[28] /*22876*/;
assign _1293_ = _893_ & _1290_ /*22871*/;
assign _1294_ = _893_ ^ _1290_ /*22874*/;
assign _1295_ = _1286_ & _1294_ /*22872*/;
assign _1117_ = _1286_ ^ _1294_ /*22873*/;
assign _1292_ = _1293_ | _1295_ /*22870*/;
assign _1297_ = ~Q[29] /*22869*/;
assign _1296_ = _1297_ & D[29] /*22868*/;
assign _1299_ = _894_ & _1296_ /*22863*/;
assign _1300_ = _894_ ^ _1296_ /*22866*/;
assign _1301_ = _1292_ & _1300_ /*22864*/;
assign _1118_ = _1292_ ^ _1300_ /*22865*/;
assign _1298_ = _1299_ | _1301_ /*22862*/;
assign _1303_ = ~Q[29] /*22861*/;
assign _1302_ = _1303_ & D[30] /*22860*/;
assign _1305_ = _895_ & _1302_ /*22855*/;
assign _1306_ = _895_ ^ _1302_ /*22858*/;
assign _1307_ = _1298_ & _1306_ /*22856*/;
assign _1119_ = _1298_ ^ _1306_ /*22857*/;
assign _1304_ = _1305_ | _1307_ /*22854*/;
assign _1309_ = ~Q[29] /*22853*/;
assign _1308_ = _1309_ & zeroWire /*22852*/;
assign _1310_ = _896_ ^ _1308_ /*22850*/;
assign _1120_ = _1310_ ^ _1304_ /*22849*/;
assign _1349_ = ~D[0] /*22723*/;
assign _1346_ = R_0[28] & _1349_ /*22719*/;
assign _1347_ = R_0[28] ^ _1349_ /*22722*/;
assign _1348_ = oneWire & _1347_ /*22720*/;
assign _1313_ = oneWire ^ _1347_ /*22721*/;
assign _1345_ = _1346_ | _1348_ /*22718*/;
assign _1354_ = ~D[1] /*22717*/;
assign _1351_ = _1089_ & _1354_ /*22713*/;
assign _1352_ = _1089_ ^ _1354_ /*22716*/;
assign _1353_ = _1345_ & _1352_ /*22714*/;
assign _1314_ = _1345_ ^ _1352_ /*22715*/;
assign _1350_ = _1351_ | _1353_ /*22712*/;
assign _1359_ = ~D[2] /*22711*/;
assign _1356_ = _1090_ & _1359_ /*22707*/;
assign _1357_ = _1090_ ^ _1359_ /*22710*/;
assign _1358_ = _1350_ & _1357_ /*22708*/;
assign _1315_ = _1350_ ^ _1357_ /*22709*/;
assign _1355_ = _1356_ | _1358_ /*22706*/;
assign _1364_ = ~D[3] /*22705*/;
assign _1361_ = _1091_ & _1364_ /*22701*/;
assign _1362_ = _1091_ ^ _1364_ /*22704*/;
assign _1363_ = _1355_ & _1362_ /*22702*/;
assign _1316_ = _1355_ ^ _1362_ /*22703*/;
assign _1360_ = _1361_ | _1363_ /*22700*/;
assign _1369_ = ~D[4] /*22699*/;
assign _1366_ = _1092_ & _1369_ /*22695*/;
assign _1367_ = _1092_ ^ _1369_ /*22698*/;
assign _1368_ = _1360_ & _1367_ /*22696*/;
assign _1317_ = _1360_ ^ _1367_ /*22697*/;
assign _1365_ = _1366_ | _1368_ /*22694*/;
assign _1374_ = ~D[5] /*22693*/;
assign _1371_ = _1093_ & _1374_ /*22689*/;
assign _1372_ = _1093_ ^ _1374_ /*22692*/;
assign _1373_ = _1365_ & _1372_ /*22690*/;
assign _1318_ = _1365_ ^ _1372_ /*22691*/;
assign _1370_ = _1371_ | _1373_ /*22688*/;
assign _1379_ = ~D[6] /*22687*/;
assign _1376_ = _1094_ & _1379_ /*22683*/;
assign _1377_ = _1094_ ^ _1379_ /*22686*/;
assign _1378_ = _1370_ & _1377_ /*22684*/;
assign _1319_ = _1370_ ^ _1377_ /*22685*/;
assign _1375_ = _1376_ | _1378_ /*22682*/;
assign _1384_ = ~D[7] /*22681*/;
assign _1381_ = _1095_ & _1384_ /*22677*/;
assign _1382_ = _1095_ ^ _1384_ /*22680*/;
assign _1383_ = _1375_ & _1382_ /*22678*/;
assign _1320_ = _1375_ ^ _1382_ /*22679*/;
assign _1380_ = _1381_ | _1383_ /*22676*/;
assign _1389_ = ~D[8] /*22675*/;
assign _1386_ = _1096_ & _1389_ /*22671*/;
assign _1387_ = _1096_ ^ _1389_ /*22674*/;
assign _1388_ = _1380_ & _1387_ /*22672*/;
assign _1321_ = _1380_ ^ _1387_ /*22673*/;
assign _1385_ = _1386_ | _1388_ /*22670*/;
assign _1394_ = ~D[9] /*22669*/;
assign _1391_ = _1097_ & _1394_ /*22665*/;
assign _1392_ = _1097_ ^ _1394_ /*22668*/;
assign _1393_ = _1385_ & _1392_ /*22666*/;
assign _1322_ = _1385_ ^ _1392_ /*22667*/;
assign _1390_ = _1391_ | _1393_ /*22664*/;
assign _1399_ = ~D[10] /*22663*/;
assign _1396_ = _1098_ & _1399_ /*22659*/;
assign _1397_ = _1098_ ^ _1399_ /*22662*/;
assign _1398_ = _1390_ & _1397_ /*22660*/;
assign _1323_ = _1390_ ^ _1397_ /*22661*/;
assign _1395_ = _1396_ | _1398_ /*22658*/;
assign _1404_ = ~D[11] /*22657*/;
assign _1401_ = _1099_ & _1404_ /*22653*/;
assign _1402_ = _1099_ ^ _1404_ /*22656*/;
assign _1403_ = _1395_ & _1402_ /*22654*/;
assign _1324_ = _1395_ ^ _1402_ /*22655*/;
assign _1400_ = _1401_ | _1403_ /*22652*/;
assign _1409_ = ~D[12] /*22651*/;
assign _1406_ = _1100_ & _1409_ /*22647*/;
assign _1407_ = _1100_ ^ _1409_ /*22650*/;
assign _1408_ = _1400_ & _1407_ /*22648*/;
assign _1325_ = _1400_ ^ _1407_ /*22649*/;
assign _1405_ = _1406_ | _1408_ /*22646*/;
assign _1414_ = ~D[13] /*22645*/;
assign _1411_ = _1101_ & _1414_ /*22641*/;
assign _1412_ = _1101_ ^ _1414_ /*22644*/;
assign _1413_ = _1405_ & _1412_ /*22642*/;
assign _1326_ = _1405_ ^ _1412_ /*22643*/;
assign _1410_ = _1411_ | _1413_ /*22640*/;
assign _1419_ = ~D[14] /*22639*/;
assign _1416_ = _1102_ & _1419_ /*22635*/;
assign _1417_ = _1102_ ^ _1419_ /*22638*/;
assign _1418_ = _1410_ & _1417_ /*22636*/;
assign _1327_ = _1410_ ^ _1417_ /*22637*/;
assign _1415_ = _1416_ | _1418_ /*22634*/;
assign _1424_ = ~D[15] /*22633*/;
assign _1421_ = _1103_ & _1424_ /*22629*/;
assign _1422_ = _1103_ ^ _1424_ /*22632*/;
assign _1423_ = _1415_ & _1422_ /*22630*/;
assign _1328_ = _1415_ ^ _1422_ /*22631*/;
assign _1420_ = _1421_ | _1423_ /*22628*/;
assign _1429_ = ~D[16] /*22627*/;
assign _1426_ = _1104_ & _1429_ /*22623*/;
assign _1427_ = _1104_ ^ _1429_ /*22626*/;
assign _1428_ = _1420_ & _1427_ /*22624*/;
assign _1329_ = _1420_ ^ _1427_ /*22625*/;
assign _1425_ = _1426_ | _1428_ /*22622*/;
assign _1434_ = ~D[17] /*22621*/;
assign _1431_ = _1105_ & _1434_ /*22617*/;
assign _1432_ = _1105_ ^ _1434_ /*22620*/;
assign _1433_ = _1425_ & _1432_ /*22618*/;
assign _1330_ = _1425_ ^ _1432_ /*22619*/;
assign _1430_ = _1431_ | _1433_ /*22616*/;
assign _1439_ = ~D[18] /*22615*/;
assign _1436_ = _1106_ & _1439_ /*22611*/;
assign _1437_ = _1106_ ^ _1439_ /*22614*/;
assign _1438_ = _1430_ & _1437_ /*22612*/;
assign _1331_ = _1430_ ^ _1437_ /*22613*/;
assign _1435_ = _1436_ | _1438_ /*22610*/;
assign _1444_ = ~D[19] /*22609*/;
assign _1441_ = _1107_ & _1444_ /*22605*/;
assign _1442_ = _1107_ ^ _1444_ /*22608*/;
assign _1443_ = _1435_ & _1442_ /*22606*/;
assign _1332_ = _1435_ ^ _1442_ /*22607*/;
assign _1440_ = _1441_ | _1443_ /*22604*/;
assign _1449_ = ~D[20] /*22603*/;
assign _1446_ = _1108_ & _1449_ /*22599*/;
assign _1447_ = _1108_ ^ _1449_ /*22602*/;
assign _1448_ = _1440_ & _1447_ /*22600*/;
assign _1333_ = _1440_ ^ _1447_ /*22601*/;
assign _1445_ = _1446_ | _1448_ /*22598*/;
assign _1454_ = ~D[21] /*22597*/;
assign _1451_ = _1109_ & _1454_ /*22593*/;
assign _1452_ = _1109_ ^ _1454_ /*22596*/;
assign _1453_ = _1445_ & _1452_ /*22594*/;
assign _1334_ = _1445_ ^ _1452_ /*22595*/;
assign _1450_ = _1451_ | _1453_ /*22592*/;
assign _1459_ = ~D[22] /*22591*/;
assign _1456_ = _1110_ & _1459_ /*22587*/;
assign _1457_ = _1110_ ^ _1459_ /*22590*/;
assign _1458_ = _1450_ & _1457_ /*22588*/;
assign _1335_ = _1450_ ^ _1457_ /*22589*/;
assign _1455_ = _1456_ | _1458_ /*22586*/;
assign _1464_ = ~D[23] /*22585*/;
assign _1461_ = _1111_ & _1464_ /*22581*/;
assign _1462_ = _1111_ ^ _1464_ /*22584*/;
assign _1463_ = _1455_ & _1462_ /*22582*/;
assign _1336_ = _1455_ ^ _1462_ /*22583*/;
assign _1460_ = _1461_ | _1463_ /*22580*/;
assign _1469_ = ~D[24] /*22579*/;
assign _1466_ = _1112_ & _1469_ /*22575*/;
assign _1467_ = _1112_ ^ _1469_ /*22578*/;
assign _1468_ = _1460_ & _1467_ /*22576*/;
assign _1337_ = _1460_ ^ _1467_ /*22577*/;
assign _1465_ = _1466_ | _1468_ /*22574*/;
assign _1474_ = ~D[25] /*22573*/;
assign _1471_ = _1113_ & _1474_ /*22569*/;
assign _1472_ = _1113_ ^ _1474_ /*22572*/;
assign _1473_ = _1465_ & _1472_ /*22570*/;
assign _1338_ = _1465_ ^ _1472_ /*22571*/;
assign _1470_ = _1471_ | _1473_ /*22568*/;
assign _1479_ = ~D[26] /*22567*/;
assign _1476_ = _1114_ & _1479_ /*22563*/;
assign _1477_ = _1114_ ^ _1479_ /*22566*/;
assign _1478_ = _1470_ & _1477_ /*22564*/;
assign _1339_ = _1470_ ^ _1477_ /*22565*/;
assign _1475_ = _1476_ | _1478_ /*22562*/;
assign _1484_ = ~D[27] /*22561*/;
assign _1481_ = _1115_ & _1484_ /*22557*/;
assign _1482_ = _1115_ ^ _1484_ /*22560*/;
assign _1483_ = _1475_ & _1482_ /*22558*/;
assign _1340_ = _1475_ ^ _1482_ /*22559*/;
assign _1480_ = _1481_ | _1483_ /*22556*/;
assign _1489_ = ~D[28] /*22555*/;
assign _1486_ = _1116_ & _1489_ /*22551*/;
assign _1487_ = _1116_ ^ _1489_ /*22554*/;
assign _1488_ = _1480_ & _1487_ /*22552*/;
assign _1341_ = _1480_ ^ _1487_ /*22553*/;
assign _1485_ = _1486_ | _1488_ /*22550*/;
assign _1494_ = ~D[29] /*22549*/;
assign _1491_ = _1117_ & _1494_ /*22545*/;
assign _1492_ = _1117_ ^ _1494_ /*22548*/;
assign _1493_ = _1485_ & _1492_ /*22546*/;
assign _1342_ = _1485_ ^ _1492_ /*22547*/;
assign _1490_ = _1491_ | _1493_ /*22544*/;
assign _1499_ = ~D[30] /*22543*/;
assign _1496_ = _1118_ & _1499_ /*22539*/;
assign _1497_ = _1118_ ^ _1499_ /*22542*/;
assign _1498_ = _1490_ & _1497_ /*22540*/;
assign _1343_ = _1490_ ^ _1497_ /*22541*/;
assign _1495_ = _1496_ | _1498_ /*22538*/;
assign _1500_ = _1119_ & oneWire /*22533*/;
assign _1501_ = _1119_ ^ oneWire /*22536*/;
assign _1502_ = _1495_ & _1501_ /*22534*/;
assign _1344_ = _1495_ ^ _1501_ /*22535*/;
assign Q[28] = _1500_ | _1502_ /*22532*/;
assign _1571_ = ~Q[28] /*22339*/;
assign _1570_ = _1571_ & D[0] /*22338*/;
assign _1573_ = _1313_ & _1570_ /*22333*/;
assign _1574_ = _1313_ ^ _1570_ /*22336*/;
assign _1575_ = zeroWire & _1574_ /*22334*/;
assign _1537_ = zeroWire ^ _1574_ /*22335*/;
assign _1572_ = _1573_ | _1575_ /*22332*/;
assign _1577_ = ~Q[28] /*22331*/;
assign _1576_ = _1577_ & D[1] /*22330*/;
assign _1579_ = _1314_ & _1576_ /*22325*/;
assign _1580_ = _1314_ ^ _1576_ /*22328*/;
assign _1581_ = _1572_ & _1580_ /*22326*/;
assign _1538_ = _1572_ ^ _1580_ /*22327*/;
assign _1578_ = _1579_ | _1581_ /*22324*/;
assign _1583_ = ~Q[28] /*22323*/;
assign _1582_ = _1583_ & D[2] /*22322*/;
assign _1585_ = _1315_ & _1582_ /*22317*/;
assign _1586_ = _1315_ ^ _1582_ /*22320*/;
assign _1587_ = _1578_ & _1586_ /*22318*/;
assign _1539_ = _1578_ ^ _1586_ /*22319*/;
assign _1584_ = _1585_ | _1587_ /*22316*/;
assign _1589_ = ~Q[28] /*22315*/;
assign _1588_ = _1589_ & D[3] /*22314*/;
assign _1591_ = _1316_ & _1588_ /*22309*/;
assign _1592_ = _1316_ ^ _1588_ /*22312*/;
assign _1593_ = _1584_ & _1592_ /*22310*/;
assign _1540_ = _1584_ ^ _1592_ /*22311*/;
assign _1590_ = _1591_ | _1593_ /*22308*/;
assign _1595_ = ~Q[28] /*22307*/;
assign _1594_ = _1595_ & D[4] /*22306*/;
assign _1597_ = _1317_ & _1594_ /*22301*/;
assign _1598_ = _1317_ ^ _1594_ /*22304*/;
assign _1599_ = _1590_ & _1598_ /*22302*/;
assign _1541_ = _1590_ ^ _1598_ /*22303*/;
assign _1596_ = _1597_ | _1599_ /*22300*/;
assign _1601_ = ~Q[28] /*22299*/;
assign _1600_ = _1601_ & D[5] /*22298*/;
assign _1603_ = _1318_ & _1600_ /*22293*/;
assign _1604_ = _1318_ ^ _1600_ /*22296*/;
assign _1605_ = _1596_ & _1604_ /*22294*/;
assign _1542_ = _1596_ ^ _1604_ /*22295*/;
assign _1602_ = _1603_ | _1605_ /*22292*/;
assign _1607_ = ~Q[28] /*22291*/;
assign _1606_ = _1607_ & D[6] /*22290*/;
assign _1609_ = _1319_ & _1606_ /*22285*/;
assign _1610_ = _1319_ ^ _1606_ /*22288*/;
assign _1611_ = _1602_ & _1610_ /*22286*/;
assign _1543_ = _1602_ ^ _1610_ /*22287*/;
assign _1608_ = _1609_ | _1611_ /*22284*/;
assign _1613_ = ~Q[28] /*22283*/;
assign _1612_ = _1613_ & D[7] /*22282*/;
assign _1615_ = _1320_ & _1612_ /*22277*/;
assign _1616_ = _1320_ ^ _1612_ /*22280*/;
assign _1617_ = _1608_ & _1616_ /*22278*/;
assign _1544_ = _1608_ ^ _1616_ /*22279*/;
assign _1614_ = _1615_ | _1617_ /*22276*/;
assign _1619_ = ~Q[28] /*22275*/;
assign _1618_ = _1619_ & D[8] /*22274*/;
assign _1621_ = _1321_ & _1618_ /*22269*/;
assign _1622_ = _1321_ ^ _1618_ /*22272*/;
assign _1623_ = _1614_ & _1622_ /*22270*/;
assign _1545_ = _1614_ ^ _1622_ /*22271*/;
assign _1620_ = _1621_ | _1623_ /*22268*/;
assign _1625_ = ~Q[28] /*22267*/;
assign _1624_ = _1625_ & D[9] /*22266*/;
assign _1627_ = _1322_ & _1624_ /*22261*/;
assign _1628_ = _1322_ ^ _1624_ /*22264*/;
assign _1629_ = _1620_ & _1628_ /*22262*/;
assign _1546_ = _1620_ ^ _1628_ /*22263*/;
assign _1626_ = _1627_ | _1629_ /*22260*/;
assign _1631_ = ~Q[28] /*22259*/;
assign _1630_ = _1631_ & D[10] /*22258*/;
assign _1633_ = _1323_ & _1630_ /*22253*/;
assign _1634_ = _1323_ ^ _1630_ /*22256*/;
assign _1635_ = _1626_ & _1634_ /*22254*/;
assign _1547_ = _1626_ ^ _1634_ /*22255*/;
assign _1632_ = _1633_ | _1635_ /*22252*/;
assign _1637_ = ~Q[28] /*22251*/;
assign _1636_ = _1637_ & D[11] /*22250*/;
assign _1639_ = _1324_ & _1636_ /*22245*/;
assign _1640_ = _1324_ ^ _1636_ /*22248*/;
assign _1641_ = _1632_ & _1640_ /*22246*/;
assign _1548_ = _1632_ ^ _1640_ /*22247*/;
assign _1638_ = _1639_ | _1641_ /*22244*/;
assign _1643_ = ~Q[28] /*22243*/;
assign _1642_ = _1643_ & D[12] /*22242*/;
assign _1645_ = _1325_ & _1642_ /*22237*/;
assign _1646_ = _1325_ ^ _1642_ /*22240*/;
assign _1647_ = _1638_ & _1646_ /*22238*/;
assign _1549_ = _1638_ ^ _1646_ /*22239*/;
assign _1644_ = _1645_ | _1647_ /*22236*/;
assign _1649_ = ~Q[28] /*22235*/;
assign _1648_ = _1649_ & D[13] /*22234*/;
assign _1651_ = _1326_ & _1648_ /*22229*/;
assign _1652_ = _1326_ ^ _1648_ /*22232*/;
assign _1653_ = _1644_ & _1652_ /*22230*/;
assign _1550_ = _1644_ ^ _1652_ /*22231*/;
assign _1650_ = _1651_ | _1653_ /*22228*/;
assign _1655_ = ~Q[28] /*22227*/;
assign _1654_ = _1655_ & D[14] /*22226*/;
assign _1657_ = _1327_ & _1654_ /*22221*/;
assign _1658_ = _1327_ ^ _1654_ /*22224*/;
assign _1659_ = _1650_ & _1658_ /*22222*/;
assign _1551_ = _1650_ ^ _1658_ /*22223*/;
assign _1656_ = _1657_ | _1659_ /*22220*/;
assign _1661_ = ~Q[28] /*22219*/;
assign _1660_ = _1661_ & D[15] /*22218*/;
assign _1663_ = _1328_ & _1660_ /*22213*/;
assign _1664_ = _1328_ ^ _1660_ /*22216*/;
assign _1665_ = _1656_ & _1664_ /*22214*/;
assign _1552_ = _1656_ ^ _1664_ /*22215*/;
assign _1662_ = _1663_ | _1665_ /*22212*/;
assign _1667_ = ~Q[28] /*22211*/;
assign _1666_ = _1667_ & D[16] /*22210*/;
assign _1669_ = _1329_ & _1666_ /*22205*/;
assign _1670_ = _1329_ ^ _1666_ /*22208*/;
assign _1671_ = _1662_ & _1670_ /*22206*/;
assign _1553_ = _1662_ ^ _1670_ /*22207*/;
assign _1668_ = _1669_ | _1671_ /*22204*/;
assign _1673_ = ~Q[28] /*22203*/;
assign _1672_ = _1673_ & D[17] /*22202*/;
assign _1675_ = _1330_ & _1672_ /*22197*/;
assign _1676_ = _1330_ ^ _1672_ /*22200*/;
assign _1677_ = _1668_ & _1676_ /*22198*/;
assign _1554_ = _1668_ ^ _1676_ /*22199*/;
assign _1674_ = _1675_ | _1677_ /*22196*/;
assign _1679_ = ~Q[28] /*22195*/;
assign _1678_ = _1679_ & D[18] /*22194*/;
assign _1681_ = _1331_ & _1678_ /*22189*/;
assign _1682_ = _1331_ ^ _1678_ /*22192*/;
assign _1683_ = _1674_ & _1682_ /*22190*/;
assign _1555_ = _1674_ ^ _1682_ /*22191*/;
assign _1680_ = _1681_ | _1683_ /*22188*/;
assign _1685_ = ~Q[28] /*22187*/;
assign _1684_ = _1685_ & D[19] /*22186*/;
assign _1687_ = _1332_ & _1684_ /*22181*/;
assign _1688_ = _1332_ ^ _1684_ /*22184*/;
assign _1689_ = _1680_ & _1688_ /*22182*/;
assign _1556_ = _1680_ ^ _1688_ /*22183*/;
assign _1686_ = _1687_ | _1689_ /*22180*/;
assign _1691_ = ~Q[28] /*22179*/;
assign _1690_ = _1691_ & D[20] /*22178*/;
assign _1693_ = _1333_ & _1690_ /*22173*/;
assign _1694_ = _1333_ ^ _1690_ /*22176*/;
assign _1695_ = _1686_ & _1694_ /*22174*/;
assign _1557_ = _1686_ ^ _1694_ /*22175*/;
assign _1692_ = _1693_ | _1695_ /*22172*/;
assign _1697_ = ~Q[28] /*22171*/;
assign _1696_ = _1697_ & D[21] /*22170*/;
assign _1699_ = _1334_ & _1696_ /*22165*/;
assign _1700_ = _1334_ ^ _1696_ /*22168*/;
assign _1701_ = _1692_ & _1700_ /*22166*/;
assign _1558_ = _1692_ ^ _1700_ /*22167*/;
assign _1698_ = _1699_ | _1701_ /*22164*/;
assign _1703_ = ~Q[28] /*22163*/;
assign _1702_ = _1703_ & D[22] /*22162*/;
assign _1705_ = _1335_ & _1702_ /*22157*/;
assign _1706_ = _1335_ ^ _1702_ /*22160*/;
assign _1707_ = _1698_ & _1706_ /*22158*/;
assign _1559_ = _1698_ ^ _1706_ /*22159*/;
assign _1704_ = _1705_ | _1707_ /*22156*/;
assign _1709_ = ~Q[28] /*22155*/;
assign _1708_ = _1709_ & D[23] /*22154*/;
assign _1711_ = _1336_ & _1708_ /*22149*/;
assign _1712_ = _1336_ ^ _1708_ /*22152*/;
assign _1713_ = _1704_ & _1712_ /*22150*/;
assign _1560_ = _1704_ ^ _1712_ /*22151*/;
assign _1710_ = _1711_ | _1713_ /*22148*/;
assign _1715_ = ~Q[28] /*22147*/;
assign _1714_ = _1715_ & D[24] /*22146*/;
assign _1717_ = _1337_ & _1714_ /*22141*/;
assign _1718_ = _1337_ ^ _1714_ /*22144*/;
assign _1719_ = _1710_ & _1718_ /*22142*/;
assign _1561_ = _1710_ ^ _1718_ /*22143*/;
assign _1716_ = _1717_ | _1719_ /*22140*/;
assign _1721_ = ~Q[28] /*22139*/;
assign _1720_ = _1721_ & D[25] /*22138*/;
assign _1723_ = _1338_ & _1720_ /*22133*/;
assign _1724_ = _1338_ ^ _1720_ /*22136*/;
assign _1725_ = _1716_ & _1724_ /*22134*/;
assign _1562_ = _1716_ ^ _1724_ /*22135*/;
assign _1722_ = _1723_ | _1725_ /*22132*/;
assign _1727_ = ~Q[28] /*22131*/;
assign _1726_ = _1727_ & D[26] /*22130*/;
assign _1729_ = _1339_ & _1726_ /*22125*/;
assign _1730_ = _1339_ ^ _1726_ /*22128*/;
assign _1731_ = _1722_ & _1730_ /*22126*/;
assign _1563_ = _1722_ ^ _1730_ /*22127*/;
assign _1728_ = _1729_ | _1731_ /*22124*/;
assign _1733_ = ~Q[28] /*22123*/;
assign _1732_ = _1733_ & D[27] /*22122*/;
assign _1735_ = _1340_ & _1732_ /*22117*/;
assign _1736_ = _1340_ ^ _1732_ /*22120*/;
assign _1737_ = _1728_ & _1736_ /*22118*/;
assign _1564_ = _1728_ ^ _1736_ /*22119*/;
assign _1734_ = _1735_ | _1737_ /*22116*/;
assign _1739_ = ~Q[28] /*22115*/;
assign _1738_ = _1739_ & D[28] /*22114*/;
assign _1741_ = _1341_ & _1738_ /*22109*/;
assign _1742_ = _1341_ ^ _1738_ /*22112*/;
assign _1743_ = _1734_ & _1742_ /*22110*/;
assign _1565_ = _1734_ ^ _1742_ /*22111*/;
assign _1740_ = _1741_ | _1743_ /*22108*/;
assign _1745_ = ~Q[28] /*22107*/;
assign _1744_ = _1745_ & D[29] /*22106*/;
assign _1747_ = _1342_ & _1744_ /*22101*/;
assign _1748_ = _1342_ ^ _1744_ /*22104*/;
assign _1749_ = _1740_ & _1748_ /*22102*/;
assign _1566_ = _1740_ ^ _1748_ /*22103*/;
assign _1746_ = _1747_ | _1749_ /*22100*/;
assign _1751_ = ~Q[28] /*22099*/;
assign _1750_ = _1751_ & D[30] /*22098*/;
assign _1753_ = _1343_ & _1750_ /*22093*/;
assign _1754_ = _1343_ ^ _1750_ /*22096*/;
assign _1755_ = _1746_ & _1754_ /*22094*/;
assign _1567_ = _1746_ ^ _1754_ /*22095*/;
assign _1752_ = _1753_ | _1755_ /*22092*/;
assign _1757_ = ~Q[28] /*22091*/;
assign _1756_ = _1757_ & zeroWire /*22090*/;
assign _1758_ = _1344_ ^ _1756_ /*22088*/;
assign _1568_ = _1758_ ^ _1752_ /*22087*/;
assign _1797_ = ~D[0] /*21961*/;
assign _1794_ = R_0[27] & _1797_ /*21957*/;
assign _1795_ = R_0[27] ^ _1797_ /*21960*/;
assign _1796_ = oneWire & _1795_ /*21958*/;
assign _1761_ = oneWire ^ _1795_ /*21959*/;
assign _1793_ = _1794_ | _1796_ /*21956*/;
assign _1802_ = ~D[1] /*21955*/;
assign _1799_ = _1537_ & _1802_ /*21951*/;
assign _1800_ = _1537_ ^ _1802_ /*21954*/;
assign _1801_ = _1793_ & _1800_ /*21952*/;
assign _1762_ = _1793_ ^ _1800_ /*21953*/;
assign _1798_ = _1799_ | _1801_ /*21950*/;
assign _1807_ = ~D[2] /*21949*/;
assign _1804_ = _1538_ & _1807_ /*21945*/;
assign _1805_ = _1538_ ^ _1807_ /*21948*/;
assign _1806_ = _1798_ & _1805_ /*21946*/;
assign _1763_ = _1798_ ^ _1805_ /*21947*/;
assign _1803_ = _1804_ | _1806_ /*21944*/;
assign _1812_ = ~D[3] /*21943*/;
assign _1809_ = _1539_ & _1812_ /*21939*/;
assign _1810_ = _1539_ ^ _1812_ /*21942*/;
assign _1811_ = _1803_ & _1810_ /*21940*/;
assign _1764_ = _1803_ ^ _1810_ /*21941*/;
assign _1808_ = _1809_ | _1811_ /*21938*/;
assign _1817_ = ~D[4] /*21937*/;
assign _1814_ = _1540_ & _1817_ /*21933*/;
assign _1815_ = _1540_ ^ _1817_ /*21936*/;
assign _1816_ = _1808_ & _1815_ /*21934*/;
assign _1765_ = _1808_ ^ _1815_ /*21935*/;
assign _1813_ = _1814_ | _1816_ /*21932*/;
assign _1822_ = ~D[5] /*21931*/;
assign _1819_ = _1541_ & _1822_ /*21927*/;
assign _1820_ = _1541_ ^ _1822_ /*21930*/;
assign _1821_ = _1813_ & _1820_ /*21928*/;
assign _1766_ = _1813_ ^ _1820_ /*21929*/;
assign _1818_ = _1819_ | _1821_ /*21926*/;
assign _1827_ = ~D[6] /*21925*/;
assign _1824_ = _1542_ & _1827_ /*21921*/;
assign _1825_ = _1542_ ^ _1827_ /*21924*/;
assign _1826_ = _1818_ & _1825_ /*21922*/;
assign _1767_ = _1818_ ^ _1825_ /*21923*/;
assign _1823_ = _1824_ | _1826_ /*21920*/;
assign _1832_ = ~D[7] /*21919*/;
assign _1829_ = _1543_ & _1832_ /*21915*/;
assign _1830_ = _1543_ ^ _1832_ /*21918*/;
assign _1831_ = _1823_ & _1830_ /*21916*/;
assign _1768_ = _1823_ ^ _1830_ /*21917*/;
assign _1828_ = _1829_ | _1831_ /*21914*/;
assign _1837_ = ~D[8] /*21913*/;
assign _1834_ = _1544_ & _1837_ /*21909*/;
assign _1835_ = _1544_ ^ _1837_ /*21912*/;
assign _1836_ = _1828_ & _1835_ /*21910*/;
assign _1769_ = _1828_ ^ _1835_ /*21911*/;
assign _1833_ = _1834_ | _1836_ /*21908*/;
assign _1842_ = ~D[9] /*21907*/;
assign _1839_ = _1545_ & _1842_ /*21903*/;
assign _1840_ = _1545_ ^ _1842_ /*21906*/;
assign _1841_ = _1833_ & _1840_ /*21904*/;
assign _1770_ = _1833_ ^ _1840_ /*21905*/;
assign _1838_ = _1839_ | _1841_ /*21902*/;
assign _1847_ = ~D[10] /*21901*/;
assign _1844_ = _1546_ & _1847_ /*21897*/;
assign _1845_ = _1546_ ^ _1847_ /*21900*/;
assign _1846_ = _1838_ & _1845_ /*21898*/;
assign _1771_ = _1838_ ^ _1845_ /*21899*/;
assign _1843_ = _1844_ | _1846_ /*21896*/;
assign _1852_ = ~D[11] /*21895*/;
assign _1849_ = _1547_ & _1852_ /*21891*/;
assign _1850_ = _1547_ ^ _1852_ /*21894*/;
assign _1851_ = _1843_ & _1850_ /*21892*/;
assign _1772_ = _1843_ ^ _1850_ /*21893*/;
assign _1848_ = _1849_ | _1851_ /*21890*/;
assign _1857_ = ~D[12] /*21889*/;
assign _1854_ = _1548_ & _1857_ /*21885*/;
assign _1855_ = _1548_ ^ _1857_ /*21888*/;
assign _1856_ = _1848_ & _1855_ /*21886*/;
assign _1773_ = _1848_ ^ _1855_ /*21887*/;
assign _1853_ = _1854_ | _1856_ /*21884*/;
assign _1862_ = ~D[13] /*21883*/;
assign _1859_ = _1549_ & _1862_ /*21879*/;
assign _1860_ = _1549_ ^ _1862_ /*21882*/;
assign _1861_ = _1853_ & _1860_ /*21880*/;
assign _1774_ = _1853_ ^ _1860_ /*21881*/;
assign _1858_ = _1859_ | _1861_ /*21878*/;
assign _1867_ = ~D[14] /*21877*/;
assign _1864_ = _1550_ & _1867_ /*21873*/;
assign _1865_ = _1550_ ^ _1867_ /*21876*/;
assign _1866_ = _1858_ & _1865_ /*21874*/;
assign _1775_ = _1858_ ^ _1865_ /*21875*/;
assign _1863_ = _1864_ | _1866_ /*21872*/;
assign _1872_ = ~D[15] /*21871*/;
assign _1869_ = _1551_ & _1872_ /*21867*/;
assign _1870_ = _1551_ ^ _1872_ /*21870*/;
assign _1871_ = _1863_ & _1870_ /*21868*/;
assign _1776_ = _1863_ ^ _1870_ /*21869*/;
assign _1868_ = _1869_ | _1871_ /*21866*/;
assign _1877_ = ~D[16] /*21865*/;
assign _1874_ = _1552_ & _1877_ /*21861*/;
assign _1875_ = _1552_ ^ _1877_ /*21864*/;
assign _1876_ = _1868_ & _1875_ /*21862*/;
assign _1777_ = _1868_ ^ _1875_ /*21863*/;
assign _1873_ = _1874_ | _1876_ /*21860*/;
assign _1882_ = ~D[17] /*21859*/;
assign _1879_ = _1553_ & _1882_ /*21855*/;
assign _1880_ = _1553_ ^ _1882_ /*21858*/;
assign _1881_ = _1873_ & _1880_ /*21856*/;
assign _1778_ = _1873_ ^ _1880_ /*21857*/;
assign _1878_ = _1879_ | _1881_ /*21854*/;
assign _1887_ = ~D[18] /*21853*/;
assign _1884_ = _1554_ & _1887_ /*21849*/;
assign _1885_ = _1554_ ^ _1887_ /*21852*/;
assign _1886_ = _1878_ & _1885_ /*21850*/;
assign _1779_ = _1878_ ^ _1885_ /*21851*/;
assign _1883_ = _1884_ | _1886_ /*21848*/;
assign _1892_ = ~D[19] /*21847*/;
assign _1889_ = _1555_ & _1892_ /*21843*/;
assign _1890_ = _1555_ ^ _1892_ /*21846*/;
assign _1891_ = _1883_ & _1890_ /*21844*/;
assign _1780_ = _1883_ ^ _1890_ /*21845*/;
assign _1888_ = _1889_ | _1891_ /*21842*/;
assign _1897_ = ~D[20] /*21841*/;
assign _1894_ = _1556_ & _1897_ /*21837*/;
assign _1895_ = _1556_ ^ _1897_ /*21840*/;
assign _1896_ = _1888_ & _1895_ /*21838*/;
assign _1781_ = _1888_ ^ _1895_ /*21839*/;
assign _1893_ = _1894_ | _1896_ /*21836*/;
assign _1902_ = ~D[21] /*21835*/;
assign _1899_ = _1557_ & _1902_ /*21831*/;
assign _1900_ = _1557_ ^ _1902_ /*21834*/;
assign _1901_ = _1893_ & _1900_ /*21832*/;
assign _1782_ = _1893_ ^ _1900_ /*21833*/;
assign _1898_ = _1899_ | _1901_ /*21830*/;
assign _1907_ = ~D[22] /*21829*/;
assign _1904_ = _1558_ & _1907_ /*21825*/;
assign _1905_ = _1558_ ^ _1907_ /*21828*/;
assign _1906_ = _1898_ & _1905_ /*21826*/;
assign _1783_ = _1898_ ^ _1905_ /*21827*/;
assign _1903_ = _1904_ | _1906_ /*21824*/;
assign _1912_ = ~D[23] /*21823*/;
assign _1909_ = _1559_ & _1912_ /*21819*/;
assign _1910_ = _1559_ ^ _1912_ /*21822*/;
assign _1911_ = _1903_ & _1910_ /*21820*/;
assign _1784_ = _1903_ ^ _1910_ /*21821*/;
assign _1908_ = _1909_ | _1911_ /*21818*/;
assign _1917_ = ~D[24] /*21817*/;
assign _1914_ = _1560_ & _1917_ /*21813*/;
assign _1915_ = _1560_ ^ _1917_ /*21816*/;
assign _1916_ = _1908_ & _1915_ /*21814*/;
assign _1785_ = _1908_ ^ _1915_ /*21815*/;
assign _1913_ = _1914_ | _1916_ /*21812*/;
assign _1922_ = ~D[25] /*21811*/;
assign _1919_ = _1561_ & _1922_ /*21807*/;
assign _1920_ = _1561_ ^ _1922_ /*21810*/;
assign _1921_ = _1913_ & _1920_ /*21808*/;
assign _1786_ = _1913_ ^ _1920_ /*21809*/;
assign _1918_ = _1919_ | _1921_ /*21806*/;
assign _1927_ = ~D[26] /*21805*/;
assign _1924_ = _1562_ & _1927_ /*21801*/;
assign _1925_ = _1562_ ^ _1927_ /*21804*/;
assign _1926_ = _1918_ & _1925_ /*21802*/;
assign _1787_ = _1918_ ^ _1925_ /*21803*/;
assign _1923_ = _1924_ | _1926_ /*21800*/;
assign _1932_ = ~D[27] /*21799*/;
assign _1929_ = _1563_ & _1932_ /*21795*/;
assign _1930_ = _1563_ ^ _1932_ /*21798*/;
assign _1931_ = _1923_ & _1930_ /*21796*/;
assign _1788_ = _1923_ ^ _1930_ /*21797*/;
assign _1928_ = _1929_ | _1931_ /*21794*/;
assign _1937_ = ~D[28] /*21793*/;
assign _1934_ = _1564_ & _1937_ /*21789*/;
assign _1935_ = _1564_ ^ _1937_ /*21792*/;
assign _1936_ = _1928_ & _1935_ /*21790*/;
assign _1789_ = _1928_ ^ _1935_ /*21791*/;
assign _1933_ = _1934_ | _1936_ /*21788*/;
assign _1942_ = ~D[29] /*21787*/;
assign _1939_ = _1565_ & _1942_ /*21783*/;
assign _1940_ = _1565_ ^ _1942_ /*21786*/;
assign _1941_ = _1933_ & _1940_ /*21784*/;
assign _1790_ = _1933_ ^ _1940_ /*21785*/;
assign _1938_ = _1939_ | _1941_ /*21782*/;
assign _1947_ = ~D[30] /*21781*/;
assign _1944_ = _1566_ & _1947_ /*21777*/;
assign _1945_ = _1566_ ^ _1947_ /*21780*/;
assign _1946_ = _1938_ & _1945_ /*21778*/;
assign _1791_ = _1938_ ^ _1945_ /*21779*/;
assign _1943_ = _1944_ | _1946_ /*21776*/;
assign _1948_ = _1567_ & oneWire /*21771*/;
assign _1949_ = _1567_ ^ oneWire /*21774*/;
assign _1950_ = _1943_ & _1949_ /*21772*/;
assign _1792_ = _1943_ ^ _1949_ /*21773*/;
assign Q[27] = _1948_ | _1950_ /*21770*/;
assign _2019_ = ~Q[27] /*21577*/;
assign _2018_ = _2019_ & D[0] /*21576*/;
assign _2021_ = _1761_ & _2018_ /*21571*/;
assign _2022_ = _1761_ ^ _2018_ /*21574*/;
assign _2023_ = zeroWire & _2022_ /*21572*/;
assign _1985_ = zeroWire ^ _2022_ /*21573*/;
assign _2020_ = _2021_ | _2023_ /*21570*/;
assign _2025_ = ~Q[27] /*21569*/;
assign _2024_ = _2025_ & D[1] /*21568*/;
assign _2027_ = _1762_ & _2024_ /*21563*/;
assign _2028_ = _1762_ ^ _2024_ /*21566*/;
assign _2029_ = _2020_ & _2028_ /*21564*/;
assign _1986_ = _2020_ ^ _2028_ /*21565*/;
assign _2026_ = _2027_ | _2029_ /*21562*/;
assign _2031_ = ~Q[27] /*21561*/;
assign _2030_ = _2031_ & D[2] /*21560*/;
assign _2033_ = _1763_ & _2030_ /*21555*/;
assign _2034_ = _1763_ ^ _2030_ /*21558*/;
assign _2035_ = _2026_ & _2034_ /*21556*/;
assign _1987_ = _2026_ ^ _2034_ /*21557*/;
assign _2032_ = _2033_ | _2035_ /*21554*/;
assign _2037_ = ~Q[27] /*21553*/;
assign _2036_ = _2037_ & D[3] /*21552*/;
assign _2039_ = _1764_ & _2036_ /*21547*/;
assign _2040_ = _1764_ ^ _2036_ /*21550*/;
assign _2041_ = _2032_ & _2040_ /*21548*/;
assign _1988_ = _2032_ ^ _2040_ /*21549*/;
assign _2038_ = _2039_ | _2041_ /*21546*/;
assign _2043_ = ~Q[27] /*21545*/;
assign _2042_ = _2043_ & D[4] /*21544*/;
assign _2045_ = _1765_ & _2042_ /*21539*/;
assign _2046_ = _1765_ ^ _2042_ /*21542*/;
assign _2047_ = _2038_ & _2046_ /*21540*/;
assign _1989_ = _2038_ ^ _2046_ /*21541*/;
assign _2044_ = _2045_ | _2047_ /*21538*/;
assign _2049_ = ~Q[27] /*21537*/;
assign _2048_ = _2049_ & D[5] /*21536*/;
assign _2051_ = _1766_ & _2048_ /*21531*/;
assign _2052_ = _1766_ ^ _2048_ /*21534*/;
assign _2053_ = _2044_ & _2052_ /*21532*/;
assign _1990_ = _2044_ ^ _2052_ /*21533*/;
assign _2050_ = _2051_ | _2053_ /*21530*/;
assign _2055_ = ~Q[27] /*21529*/;
assign _2054_ = _2055_ & D[6] /*21528*/;
assign _2057_ = _1767_ & _2054_ /*21523*/;
assign _2058_ = _1767_ ^ _2054_ /*21526*/;
assign _2059_ = _2050_ & _2058_ /*21524*/;
assign _1991_ = _2050_ ^ _2058_ /*21525*/;
assign _2056_ = _2057_ | _2059_ /*21522*/;
assign _2061_ = ~Q[27] /*21521*/;
assign _2060_ = _2061_ & D[7] /*21520*/;
assign _2063_ = _1768_ & _2060_ /*21515*/;
assign _2064_ = _1768_ ^ _2060_ /*21518*/;
assign _2065_ = _2056_ & _2064_ /*21516*/;
assign _1992_ = _2056_ ^ _2064_ /*21517*/;
assign _2062_ = _2063_ | _2065_ /*21514*/;
assign _2067_ = ~Q[27] /*21513*/;
assign _2066_ = _2067_ & D[8] /*21512*/;
assign _2069_ = _1769_ & _2066_ /*21507*/;
assign _2070_ = _1769_ ^ _2066_ /*21510*/;
assign _2071_ = _2062_ & _2070_ /*21508*/;
assign _1993_ = _2062_ ^ _2070_ /*21509*/;
assign _2068_ = _2069_ | _2071_ /*21506*/;
assign _2073_ = ~Q[27] /*21505*/;
assign _2072_ = _2073_ & D[9] /*21504*/;
assign _2075_ = _1770_ & _2072_ /*21499*/;
assign _2076_ = _1770_ ^ _2072_ /*21502*/;
assign _2077_ = _2068_ & _2076_ /*21500*/;
assign _1994_ = _2068_ ^ _2076_ /*21501*/;
assign _2074_ = _2075_ | _2077_ /*21498*/;
assign _2079_ = ~Q[27] /*21497*/;
assign _2078_ = _2079_ & D[10] /*21496*/;
assign _2081_ = _1771_ & _2078_ /*21491*/;
assign _2082_ = _1771_ ^ _2078_ /*21494*/;
assign _2083_ = _2074_ & _2082_ /*21492*/;
assign _1995_ = _2074_ ^ _2082_ /*21493*/;
assign _2080_ = _2081_ | _2083_ /*21490*/;
assign _2085_ = ~Q[27] /*21489*/;
assign _2084_ = _2085_ & D[11] /*21488*/;
assign _2087_ = _1772_ & _2084_ /*21483*/;
assign _2088_ = _1772_ ^ _2084_ /*21486*/;
assign _2089_ = _2080_ & _2088_ /*21484*/;
assign _1996_ = _2080_ ^ _2088_ /*21485*/;
assign _2086_ = _2087_ | _2089_ /*21482*/;
assign _2091_ = ~Q[27] /*21481*/;
assign _2090_ = _2091_ & D[12] /*21480*/;
assign _2093_ = _1773_ & _2090_ /*21475*/;
assign _2094_ = _1773_ ^ _2090_ /*21478*/;
assign _2095_ = _2086_ & _2094_ /*21476*/;
assign _1997_ = _2086_ ^ _2094_ /*21477*/;
assign _2092_ = _2093_ | _2095_ /*21474*/;
assign _2097_ = ~Q[27] /*21473*/;
assign _2096_ = _2097_ & D[13] /*21472*/;
assign _2099_ = _1774_ & _2096_ /*21467*/;
assign _2100_ = _1774_ ^ _2096_ /*21470*/;
assign _2101_ = _2092_ & _2100_ /*21468*/;
assign _1998_ = _2092_ ^ _2100_ /*21469*/;
assign _2098_ = _2099_ | _2101_ /*21466*/;
assign _2103_ = ~Q[27] /*21465*/;
assign _2102_ = _2103_ & D[14] /*21464*/;
assign _2105_ = _1775_ & _2102_ /*21459*/;
assign _2106_ = _1775_ ^ _2102_ /*21462*/;
assign _2107_ = _2098_ & _2106_ /*21460*/;
assign _1999_ = _2098_ ^ _2106_ /*21461*/;
assign _2104_ = _2105_ | _2107_ /*21458*/;
assign _2109_ = ~Q[27] /*21457*/;
assign _2108_ = _2109_ & D[15] /*21456*/;
assign _2111_ = _1776_ & _2108_ /*21451*/;
assign _2112_ = _1776_ ^ _2108_ /*21454*/;
assign _2113_ = _2104_ & _2112_ /*21452*/;
assign _2000_ = _2104_ ^ _2112_ /*21453*/;
assign _2110_ = _2111_ | _2113_ /*21450*/;
assign _2115_ = ~Q[27] /*21449*/;
assign _2114_ = _2115_ & D[16] /*21448*/;
assign _2117_ = _1777_ & _2114_ /*21443*/;
assign _2118_ = _1777_ ^ _2114_ /*21446*/;
assign _2119_ = _2110_ & _2118_ /*21444*/;
assign _2001_ = _2110_ ^ _2118_ /*21445*/;
assign _2116_ = _2117_ | _2119_ /*21442*/;
assign _2121_ = ~Q[27] /*21441*/;
assign _2120_ = _2121_ & D[17] /*21440*/;
assign _2123_ = _1778_ & _2120_ /*21435*/;
assign _2124_ = _1778_ ^ _2120_ /*21438*/;
assign _2125_ = _2116_ & _2124_ /*21436*/;
assign _2002_ = _2116_ ^ _2124_ /*21437*/;
assign _2122_ = _2123_ | _2125_ /*21434*/;
assign _2127_ = ~Q[27] /*21433*/;
assign _2126_ = _2127_ & D[18] /*21432*/;
assign _2129_ = _1779_ & _2126_ /*21427*/;
assign _2130_ = _1779_ ^ _2126_ /*21430*/;
assign _2131_ = _2122_ & _2130_ /*21428*/;
assign _2003_ = _2122_ ^ _2130_ /*21429*/;
assign _2128_ = _2129_ | _2131_ /*21426*/;
assign _2133_ = ~Q[27] /*21425*/;
assign _2132_ = _2133_ & D[19] /*21424*/;
assign _2135_ = _1780_ & _2132_ /*21419*/;
assign _2136_ = _1780_ ^ _2132_ /*21422*/;
assign _2137_ = _2128_ & _2136_ /*21420*/;
assign _2004_ = _2128_ ^ _2136_ /*21421*/;
assign _2134_ = _2135_ | _2137_ /*21418*/;
assign _2139_ = ~Q[27] /*21417*/;
assign _2138_ = _2139_ & D[20] /*21416*/;
assign _2141_ = _1781_ & _2138_ /*21411*/;
assign _2142_ = _1781_ ^ _2138_ /*21414*/;
assign _2143_ = _2134_ & _2142_ /*21412*/;
assign _2005_ = _2134_ ^ _2142_ /*21413*/;
assign _2140_ = _2141_ | _2143_ /*21410*/;
assign _2145_ = ~Q[27] /*21409*/;
assign _2144_ = _2145_ & D[21] /*21408*/;
assign _2147_ = _1782_ & _2144_ /*21403*/;
assign _2148_ = _1782_ ^ _2144_ /*21406*/;
assign _2149_ = _2140_ & _2148_ /*21404*/;
assign _2006_ = _2140_ ^ _2148_ /*21405*/;
assign _2146_ = _2147_ | _2149_ /*21402*/;
assign _2151_ = ~Q[27] /*21401*/;
assign _2150_ = _2151_ & D[22] /*21400*/;
assign _2153_ = _1783_ & _2150_ /*21395*/;
assign _2154_ = _1783_ ^ _2150_ /*21398*/;
assign _2155_ = _2146_ & _2154_ /*21396*/;
assign _2007_ = _2146_ ^ _2154_ /*21397*/;
assign _2152_ = _2153_ | _2155_ /*21394*/;
assign _2157_ = ~Q[27] /*21393*/;
assign _2156_ = _2157_ & D[23] /*21392*/;
assign _2159_ = _1784_ & _2156_ /*21387*/;
assign _2160_ = _1784_ ^ _2156_ /*21390*/;
assign _2161_ = _2152_ & _2160_ /*21388*/;
assign _2008_ = _2152_ ^ _2160_ /*21389*/;
assign _2158_ = _2159_ | _2161_ /*21386*/;
assign _2163_ = ~Q[27] /*21385*/;
assign _2162_ = _2163_ & D[24] /*21384*/;
assign _2165_ = _1785_ & _2162_ /*21379*/;
assign _2166_ = _1785_ ^ _2162_ /*21382*/;
assign _2167_ = _2158_ & _2166_ /*21380*/;
assign _2009_ = _2158_ ^ _2166_ /*21381*/;
assign _2164_ = _2165_ | _2167_ /*21378*/;
assign _2169_ = ~Q[27] /*21377*/;
assign _2168_ = _2169_ & D[25] /*21376*/;
assign _2171_ = _1786_ & _2168_ /*21371*/;
assign _2172_ = _1786_ ^ _2168_ /*21374*/;
assign _2173_ = _2164_ & _2172_ /*21372*/;
assign _2010_ = _2164_ ^ _2172_ /*21373*/;
assign _2170_ = _2171_ | _2173_ /*21370*/;
assign _2175_ = ~Q[27] /*21369*/;
assign _2174_ = _2175_ & D[26] /*21368*/;
assign _2177_ = _1787_ & _2174_ /*21363*/;
assign _2178_ = _1787_ ^ _2174_ /*21366*/;
assign _2179_ = _2170_ & _2178_ /*21364*/;
assign _2011_ = _2170_ ^ _2178_ /*21365*/;
assign _2176_ = _2177_ | _2179_ /*21362*/;
assign _2181_ = ~Q[27] /*21361*/;
assign _2180_ = _2181_ & D[27] /*21360*/;
assign _2183_ = _1788_ & _2180_ /*21355*/;
assign _2184_ = _1788_ ^ _2180_ /*21358*/;
assign _2185_ = _2176_ & _2184_ /*21356*/;
assign _2012_ = _2176_ ^ _2184_ /*21357*/;
assign _2182_ = _2183_ | _2185_ /*21354*/;
assign _2187_ = ~Q[27] /*21353*/;
assign _2186_ = _2187_ & D[28] /*21352*/;
assign _2189_ = _1789_ & _2186_ /*21347*/;
assign _2190_ = _1789_ ^ _2186_ /*21350*/;
assign _2191_ = _2182_ & _2190_ /*21348*/;
assign _2013_ = _2182_ ^ _2190_ /*21349*/;
assign _2188_ = _2189_ | _2191_ /*21346*/;
assign _2193_ = ~Q[27] /*21345*/;
assign _2192_ = _2193_ & D[29] /*21344*/;
assign _2195_ = _1790_ & _2192_ /*21339*/;
assign _2196_ = _1790_ ^ _2192_ /*21342*/;
assign _2197_ = _2188_ & _2196_ /*21340*/;
assign _2014_ = _2188_ ^ _2196_ /*21341*/;
assign _2194_ = _2195_ | _2197_ /*21338*/;
assign _2199_ = ~Q[27] /*21337*/;
assign _2198_ = _2199_ & D[30] /*21336*/;
assign _2201_ = _1791_ & _2198_ /*21331*/;
assign _2202_ = _1791_ ^ _2198_ /*21334*/;
assign _2203_ = _2194_ & _2202_ /*21332*/;
assign _2015_ = _2194_ ^ _2202_ /*21333*/;
assign _2200_ = _2201_ | _2203_ /*21330*/;
assign _2205_ = ~Q[27] /*21329*/;
assign _2204_ = _2205_ & zeroWire /*21328*/;
assign _2206_ = _1792_ ^ _2204_ /*21326*/;
assign _2016_ = _2206_ ^ _2200_ /*21325*/;
assign _2245_ = ~D[0] /*21199*/;
assign _2242_ = R_0[26] & _2245_ /*21195*/;
assign _2243_ = R_0[26] ^ _2245_ /*21198*/;
assign _2244_ = oneWire & _2243_ /*21196*/;
assign _2209_ = oneWire ^ _2243_ /*21197*/;
assign _2241_ = _2242_ | _2244_ /*21194*/;
assign _2250_ = ~D[1] /*21193*/;
assign _2247_ = _1985_ & _2250_ /*21189*/;
assign _2248_ = _1985_ ^ _2250_ /*21192*/;
assign _2249_ = _2241_ & _2248_ /*21190*/;
assign _2210_ = _2241_ ^ _2248_ /*21191*/;
assign _2246_ = _2247_ | _2249_ /*21188*/;
assign _2255_ = ~D[2] /*21187*/;
assign _2252_ = _1986_ & _2255_ /*21183*/;
assign _2253_ = _1986_ ^ _2255_ /*21186*/;
assign _2254_ = _2246_ & _2253_ /*21184*/;
assign _2211_ = _2246_ ^ _2253_ /*21185*/;
assign _2251_ = _2252_ | _2254_ /*21182*/;
assign _2260_ = ~D[3] /*21181*/;
assign _2257_ = _1987_ & _2260_ /*21177*/;
assign _2258_ = _1987_ ^ _2260_ /*21180*/;
assign _2259_ = _2251_ & _2258_ /*21178*/;
assign _2212_ = _2251_ ^ _2258_ /*21179*/;
assign _2256_ = _2257_ | _2259_ /*21176*/;
assign _2265_ = ~D[4] /*21175*/;
assign _2262_ = _1988_ & _2265_ /*21171*/;
assign _2263_ = _1988_ ^ _2265_ /*21174*/;
assign _2264_ = _2256_ & _2263_ /*21172*/;
assign _2213_ = _2256_ ^ _2263_ /*21173*/;
assign _2261_ = _2262_ | _2264_ /*21170*/;
assign _2270_ = ~D[5] /*21169*/;
assign _2267_ = _1989_ & _2270_ /*21165*/;
assign _2268_ = _1989_ ^ _2270_ /*21168*/;
assign _2269_ = _2261_ & _2268_ /*21166*/;
assign _2214_ = _2261_ ^ _2268_ /*21167*/;
assign _2266_ = _2267_ | _2269_ /*21164*/;
assign _2275_ = ~D[6] /*21163*/;
assign _2272_ = _1990_ & _2275_ /*21159*/;
assign _2273_ = _1990_ ^ _2275_ /*21162*/;
assign _2274_ = _2266_ & _2273_ /*21160*/;
assign _2215_ = _2266_ ^ _2273_ /*21161*/;
assign _2271_ = _2272_ | _2274_ /*21158*/;
assign _2280_ = ~D[7] /*21157*/;
assign _2277_ = _1991_ & _2280_ /*21153*/;
assign _2278_ = _1991_ ^ _2280_ /*21156*/;
assign _2279_ = _2271_ & _2278_ /*21154*/;
assign _2216_ = _2271_ ^ _2278_ /*21155*/;
assign _2276_ = _2277_ | _2279_ /*21152*/;
assign _2285_ = ~D[8] /*21151*/;
assign _2282_ = _1992_ & _2285_ /*21147*/;
assign _2283_ = _1992_ ^ _2285_ /*21150*/;
assign _2284_ = _2276_ & _2283_ /*21148*/;
assign _2217_ = _2276_ ^ _2283_ /*21149*/;
assign _2281_ = _2282_ | _2284_ /*21146*/;
assign _2290_ = ~D[9] /*21145*/;
assign _2287_ = _1993_ & _2290_ /*21141*/;
assign _2288_ = _1993_ ^ _2290_ /*21144*/;
assign _2289_ = _2281_ & _2288_ /*21142*/;
assign _2218_ = _2281_ ^ _2288_ /*21143*/;
assign _2286_ = _2287_ | _2289_ /*21140*/;
assign _2295_ = ~D[10] /*21139*/;
assign _2292_ = _1994_ & _2295_ /*21135*/;
assign _2293_ = _1994_ ^ _2295_ /*21138*/;
assign _2294_ = _2286_ & _2293_ /*21136*/;
assign _2219_ = _2286_ ^ _2293_ /*21137*/;
assign _2291_ = _2292_ | _2294_ /*21134*/;
assign _2300_ = ~D[11] /*21133*/;
assign _2297_ = _1995_ & _2300_ /*21129*/;
assign _2298_ = _1995_ ^ _2300_ /*21132*/;
assign _2299_ = _2291_ & _2298_ /*21130*/;
assign _2220_ = _2291_ ^ _2298_ /*21131*/;
assign _2296_ = _2297_ | _2299_ /*21128*/;
assign _2305_ = ~D[12] /*21127*/;
assign _2302_ = _1996_ & _2305_ /*21123*/;
assign _2303_ = _1996_ ^ _2305_ /*21126*/;
assign _2304_ = _2296_ & _2303_ /*21124*/;
assign _2221_ = _2296_ ^ _2303_ /*21125*/;
assign _2301_ = _2302_ | _2304_ /*21122*/;
assign _2310_ = ~D[13] /*21121*/;
assign _2307_ = _1997_ & _2310_ /*21117*/;
assign _2308_ = _1997_ ^ _2310_ /*21120*/;
assign _2309_ = _2301_ & _2308_ /*21118*/;
assign _2222_ = _2301_ ^ _2308_ /*21119*/;
assign _2306_ = _2307_ | _2309_ /*21116*/;
assign _2315_ = ~D[14] /*21115*/;
assign _2312_ = _1998_ & _2315_ /*21111*/;
assign _2313_ = _1998_ ^ _2315_ /*21114*/;
assign _2314_ = _2306_ & _2313_ /*21112*/;
assign _2223_ = _2306_ ^ _2313_ /*21113*/;
assign _2311_ = _2312_ | _2314_ /*21110*/;
assign _2320_ = ~D[15] /*21109*/;
assign _2317_ = _1999_ & _2320_ /*21105*/;
assign _2318_ = _1999_ ^ _2320_ /*21108*/;
assign _2319_ = _2311_ & _2318_ /*21106*/;
assign _2224_ = _2311_ ^ _2318_ /*21107*/;
assign _2316_ = _2317_ | _2319_ /*21104*/;
assign _2325_ = ~D[16] /*21103*/;
assign _2322_ = _2000_ & _2325_ /*21099*/;
assign _2323_ = _2000_ ^ _2325_ /*21102*/;
assign _2324_ = _2316_ & _2323_ /*21100*/;
assign _2225_ = _2316_ ^ _2323_ /*21101*/;
assign _2321_ = _2322_ | _2324_ /*21098*/;
assign _2330_ = ~D[17] /*21097*/;
assign _2327_ = _2001_ & _2330_ /*21093*/;
assign _2328_ = _2001_ ^ _2330_ /*21096*/;
assign _2329_ = _2321_ & _2328_ /*21094*/;
assign _2226_ = _2321_ ^ _2328_ /*21095*/;
assign _2326_ = _2327_ | _2329_ /*21092*/;
assign _2335_ = ~D[18] /*21091*/;
assign _2332_ = _2002_ & _2335_ /*21087*/;
assign _2333_ = _2002_ ^ _2335_ /*21090*/;
assign _2334_ = _2326_ & _2333_ /*21088*/;
assign _2227_ = _2326_ ^ _2333_ /*21089*/;
assign _2331_ = _2332_ | _2334_ /*21086*/;
assign _2340_ = ~D[19] /*21085*/;
assign _2337_ = _2003_ & _2340_ /*21081*/;
assign _2338_ = _2003_ ^ _2340_ /*21084*/;
assign _2339_ = _2331_ & _2338_ /*21082*/;
assign _2228_ = _2331_ ^ _2338_ /*21083*/;
assign _2336_ = _2337_ | _2339_ /*21080*/;
assign _2345_ = ~D[20] /*21079*/;
assign _2342_ = _2004_ & _2345_ /*21075*/;
assign _2343_ = _2004_ ^ _2345_ /*21078*/;
assign _2344_ = _2336_ & _2343_ /*21076*/;
assign _2229_ = _2336_ ^ _2343_ /*21077*/;
assign _2341_ = _2342_ | _2344_ /*21074*/;
assign _2350_ = ~D[21] /*21073*/;
assign _2347_ = _2005_ & _2350_ /*21069*/;
assign _2348_ = _2005_ ^ _2350_ /*21072*/;
assign _2349_ = _2341_ & _2348_ /*21070*/;
assign _2230_ = _2341_ ^ _2348_ /*21071*/;
assign _2346_ = _2347_ | _2349_ /*21068*/;
assign _2355_ = ~D[22] /*21067*/;
assign _2352_ = _2006_ & _2355_ /*21063*/;
assign _2353_ = _2006_ ^ _2355_ /*21066*/;
assign _2354_ = _2346_ & _2353_ /*21064*/;
assign _2231_ = _2346_ ^ _2353_ /*21065*/;
assign _2351_ = _2352_ | _2354_ /*21062*/;
assign _2360_ = ~D[23] /*21061*/;
assign _2357_ = _2007_ & _2360_ /*21057*/;
assign _2358_ = _2007_ ^ _2360_ /*21060*/;
assign _2359_ = _2351_ & _2358_ /*21058*/;
assign _2232_ = _2351_ ^ _2358_ /*21059*/;
assign _2356_ = _2357_ | _2359_ /*21056*/;
assign _2365_ = ~D[24] /*21055*/;
assign _2362_ = _2008_ & _2365_ /*21051*/;
assign _2363_ = _2008_ ^ _2365_ /*21054*/;
assign _2364_ = _2356_ & _2363_ /*21052*/;
assign _2233_ = _2356_ ^ _2363_ /*21053*/;
assign _2361_ = _2362_ | _2364_ /*21050*/;
assign _2370_ = ~D[25] /*21049*/;
assign _2367_ = _2009_ & _2370_ /*21045*/;
assign _2368_ = _2009_ ^ _2370_ /*21048*/;
assign _2369_ = _2361_ & _2368_ /*21046*/;
assign _2234_ = _2361_ ^ _2368_ /*21047*/;
assign _2366_ = _2367_ | _2369_ /*21044*/;
assign _2375_ = ~D[26] /*21043*/;
assign _2372_ = _2010_ & _2375_ /*21039*/;
assign _2373_ = _2010_ ^ _2375_ /*21042*/;
assign _2374_ = _2366_ & _2373_ /*21040*/;
assign _2235_ = _2366_ ^ _2373_ /*21041*/;
assign _2371_ = _2372_ | _2374_ /*21038*/;
assign _2380_ = ~D[27] /*21037*/;
assign _2377_ = _2011_ & _2380_ /*21033*/;
assign _2378_ = _2011_ ^ _2380_ /*21036*/;
assign _2379_ = _2371_ & _2378_ /*21034*/;
assign _2236_ = _2371_ ^ _2378_ /*21035*/;
assign _2376_ = _2377_ | _2379_ /*21032*/;
assign _2385_ = ~D[28] /*21031*/;
assign _2382_ = _2012_ & _2385_ /*21027*/;
assign _2383_ = _2012_ ^ _2385_ /*21030*/;
assign _2384_ = _2376_ & _2383_ /*21028*/;
assign _2237_ = _2376_ ^ _2383_ /*21029*/;
assign _2381_ = _2382_ | _2384_ /*21026*/;
assign _2390_ = ~D[29] /*21025*/;
assign _2387_ = _2013_ & _2390_ /*21021*/;
assign _2388_ = _2013_ ^ _2390_ /*21024*/;
assign _2389_ = _2381_ & _2388_ /*21022*/;
assign _2238_ = _2381_ ^ _2388_ /*21023*/;
assign _2386_ = _2387_ | _2389_ /*21020*/;
assign _2395_ = ~D[30] /*21019*/;
assign _2392_ = _2014_ & _2395_ /*21015*/;
assign _2393_ = _2014_ ^ _2395_ /*21018*/;
assign _2394_ = _2386_ & _2393_ /*21016*/;
assign _2239_ = _2386_ ^ _2393_ /*21017*/;
assign _2391_ = _2392_ | _2394_ /*21014*/;
assign _2396_ = _2015_ & oneWire /*21009*/;
assign _2397_ = _2015_ ^ oneWire /*21012*/;
assign _2398_ = _2391_ & _2397_ /*21010*/;
assign _2240_ = _2391_ ^ _2397_ /*21011*/;
assign Q[26] = _2396_ | _2398_ /*21008*/;
assign _2467_ = ~Q[26] /*20815*/;
assign _2466_ = _2467_ & D[0] /*20814*/;
assign _2469_ = _2209_ & _2466_ /*20809*/;
assign _2470_ = _2209_ ^ _2466_ /*20812*/;
assign _2471_ = zeroWire & _2470_ /*20810*/;
assign _2433_ = zeroWire ^ _2470_ /*20811*/;
assign _2468_ = _2469_ | _2471_ /*20808*/;
assign _2473_ = ~Q[26] /*20807*/;
assign _2472_ = _2473_ & D[1] /*20806*/;
assign _2475_ = _2210_ & _2472_ /*20801*/;
assign _2476_ = _2210_ ^ _2472_ /*20804*/;
assign _2477_ = _2468_ & _2476_ /*20802*/;
assign _2434_ = _2468_ ^ _2476_ /*20803*/;
assign _2474_ = _2475_ | _2477_ /*20800*/;
assign _2479_ = ~Q[26] /*20799*/;
assign _2478_ = _2479_ & D[2] /*20798*/;
assign _2481_ = _2211_ & _2478_ /*20793*/;
assign _2482_ = _2211_ ^ _2478_ /*20796*/;
assign _2483_ = _2474_ & _2482_ /*20794*/;
assign _2435_ = _2474_ ^ _2482_ /*20795*/;
assign _2480_ = _2481_ | _2483_ /*20792*/;
assign _2485_ = ~Q[26] /*20791*/;
assign _2484_ = _2485_ & D[3] /*20790*/;
assign _2487_ = _2212_ & _2484_ /*20785*/;
assign _2488_ = _2212_ ^ _2484_ /*20788*/;
assign _2489_ = _2480_ & _2488_ /*20786*/;
assign _2436_ = _2480_ ^ _2488_ /*20787*/;
assign _2486_ = _2487_ | _2489_ /*20784*/;
assign _2491_ = ~Q[26] /*20783*/;
assign _2490_ = _2491_ & D[4] /*20782*/;
assign _2493_ = _2213_ & _2490_ /*20777*/;
assign _2494_ = _2213_ ^ _2490_ /*20780*/;
assign _2495_ = _2486_ & _2494_ /*20778*/;
assign _2437_ = _2486_ ^ _2494_ /*20779*/;
assign _2492_ = _2493_ | _2495_ /*20776*/;
assign _2497_ = ~Q[26] /*20775*/;
assign _2496_ = _2497_ & D[5] /*20774*/;
assign _2499_ = _2214_ & _2496_ /*20769*/;
assign _2500_ = _2214_ ^ _2496_ /*20772*/;
assign _2501_ = _2492_ & _2500_ /*20770*/;
assign _2438_ = _2492_ ^ _2500_ /*20771*/;
assign _2498_ = _2499_ | _2501_ /*20768*/;
assign _2503_ = ~Q[26] /*20767*/;
assign _2502_ = _2503_ & D[6] /*20766*/;
assign _2505_ = _2215_ & _2502_ /*20761*/;
assign _2506_ = _2215_ ^ _2502_ /*20764*/;
assign _2507_ = _2498_ & _2506_ /*20762*/;
assign _2439_ = _2498_ ^ _2506_ /*20763*/;
assign _2504_ = _2505_ | _2507_ /*20760*/;
assign _2509_ = ~Q[26] /*20759*/;
assign _2508_ = _2509_ & D[7] /*20758*/;
assign _2511_ = _2216_ & _2508_ /*20753*/;
assign _2512_ = _2216_ ^ _2508_ /*20756*/;
assign _2513_ = _2504_ & _2512_ /*20754*/;
assign _2440_ = _2504_ ^ _2512_ /*20755*/;
assign _2510_ = _2511_ | _2513_ /*20752*/;
assign _2515_ = ~Q[26] /*20751*/;
assign _2514_ = _2515_ & D[8] /*20750*/;
assign _2517_ = _2217_ & _2514_ /*20745*/;
assign _2518_ = _2217_ ^ _2514_ /*20748*/;
assign _2519_ = _2510_ & _2518_ /*20746*/;
assign _2441_ = _2510_ ^ _2518_ /*20747*/;
assign _2516_ = _2517_ | _2519_ /*20744*/;
assign _2521_ = ~Q[26] /*20743*/;
assign _2520_ = _2521_ & D[9] /*20742*/;
assign _2523_ = _2218_ & _2520_ /*20737*/;
assign _2524_ = _2218_ ^ _2520_ /*20740*/;
assign _2525_ = _2516_ & _2524_ /*20738*/;
assign _2442_ = _2516_ ^ _2524_ /*20739*/;
assign _2522_ = _2523_ | _2525_ /*20736*/;
assign _2527_ = ~Q[26] /*20735*/;
assign _2526_ = _2527_ & D[10] /*20734*/;
assign _2529_ = _2219_ & _2526_ /*20729*/;
assign _2530_ = _2219_ ^ _2526_ /*20732*/;
assign _2531_ = _2522_ & _2530_ /*20730*/;
assign _2443_ = _2522_ ^ _2530_ /*20731*/;
assign _2528_ = _2529_ | _2531_ /*20728*/;
assign _2533_ = ~Q[26] /*20727*/;
assign _2532_ = _2533_ & D[11] /*20726*/;
assign _2535_ = _2220_ & _2532_ /*20721*/;
assign _2536_ = _2220_ ^ _2532_ /*20724*/;
assign _2537_ = _2528_ & _2536_ /*20722*/;
assign _2444_ = _2528_ ^ _2536_ /*20723*/;
assign _2534_ = _2535_ | _2537_ /*20720*/;
assign _2539_ = ~Q[26] /*20719*/;
assign _2538_ = _2539_ & D[12] /*20718*/;
assign _2541_ = _2221_ & _2538_ /*20713*/;
assign _2542_ = _2221_ ^ _2538_ /*20716*/;
assign _2543_ = _2534_ & _2542_ /*20714*/;
assign _2445_ = _2534_ ^ _2542_ /*20715*/;
assign _2540_ = _2541_ | _2543_ /*20712*/;
assign _2545_ = ~Q[26] /*20711*/;
assign _2544_ = _2545_ & D[13] /*20710*/;
assign _2547_ = _2222_ & _2544_ /*20705*/;
assign _2548_ = _2222_ ^ _2544_ /*20708*/;
assign _2549_ = _2540_ & _2548_ /*20706*/;
assign _2446_ = _2540_ ^ _2548_ /*20707*/;
assign _2546_ = _2547_ | _2549_ /*20704*/;
assign _2551_ = ~Q[26] /*20703*/;
assign _2550_ = _2551_ & D[14] /*20702*/;
assign _2553_ = _2223_ & _2550_ /*20697*/;
assign _2554_ = _2223_ ^ _2550_ /*20700*/;
assign _2555_ = _2546_ & _2554_ /*20698*/;
assign _2447_ = _2546_ ^ _2554_ /*20699*/;
assign _2552_ = _2553_ | _2555_ /*20696*/;
assign _2557_ = ~Q[26] /*20695*/;
assign _2556_ = _2557_ & D[15] /*20694*/;
assign _2559_ = _2224_ & _2556_ /*20689*/;
assign _2560_ = _2224_ ^ _2556_ /*20692*/;
assign _2561_ = _2552_ & _2560_ /*20690*/;
assign _2448_ = _2552_ ^ _2560_ /*20691*/;
assign _2558_ = _2559_ | _2561_ /*20688*/;
assign _2563_ = ~Q[26] /*20687*/;
assign _2562_ = _2563_ & D[16] /*20686*/;
assign _2565_ = _2225_ & _2562_ /*20681*/;
assign _2566_ = _2225_ ^ _2562_ /*20684*/;
assign _2567_ = _2558_ & _2566_ /*20682*/;
assign _2449_ = _2558_ ^ _2566_ /*20683*/;
assign _2564_ = _2565_ | _2567_ /*20680*/;
assign _2569_ = ~Q[26] /*20679*/;
assign _2568_ = _2569_ & D[17] /*20678*/;
assign _2571_ = _2226_ & _2568_ /*20673*/;
assign _2572_ = _2226_ ^ _2568_ /*20676*/;
assign _2573_ = _2564_ & _2572_ /*20674*/;
assign _2450_ = _2564_ ^ _2572_ /*20675*/;
assign _2570_ = _2571_ | _2573_ /*20672*/;
assign _2575_ = ~Q[26] /*20671*/;
assign _2574_ = _2575_ & D[18] /*20670*/;
assign _2577_ = _2227_ & _2574_ /*20665*/;
assign _2578_ = _2227_ ^ _2574_ /*20668*/;
assign _2579_ = _2570_ & _2578_ /*20666*/;
assign _2451_ = _2570_ ^ _2578_ /*20667*/;
assign _2576_ = _2577_ | _2579_ /*20664*/;
assign _2581_ = ~Q[26] /*20663*/;
assign _2580_ = _2581_ & D[19] /*20662*/;
assign _2583_ = _2228_ & _2580_ /*20657*/;
assign _2584_ = _2228_ ^ _2580_ /*20660*/;
assign _2585_ = _2576_ & _2584_ /*20658*/;
assign _2452_ = _2576_ ^ _2584_ /*20659*/;
assign _2582_ = _2583_ | _2585_ /*20656*/;
assign _2587_ = ~Q[26] /*20655*/;
assign _2586_ = _2587_ & D[20] /*20654*/;
assign _2589_ = _2229_ & _2586_ /*20649*/;
assign _2590_ = _2229_ ^ _2586_ /*20652*/;
assign _2591_ = _2582_ & _2590_ /*20650*/;
assign _2453_ = _2582_ ^ _2590_ /*20651*/;
assign _2588_ = _2589_ | _2591_ /*20648*/;
assign _2593_ = ~Q[26] /*20647*/;
assign _2592_ = _2593_ & D[21] /*20646*/;
assign _2595_ = _2230_ & _2592_ /*20641*/;
assign _2596_ = _2230_ ^ _2592_ /*20644*/;
assign _2597_ = _2588_ & _2596_ /*20642*/;
assign _2454_ = _2588_ ^ _2596_ /*20643*/;
assign _2594_ = _2595_ | _2597_ /*20640*/;
assign _2599_ = ~Q[26] /*20639*/;
assign _2598_ = _2599_ & D[22] /*20638*/;
assign _2601_ = _2231_ & _2598_ /*20633*/;
assign _2602_ = _2231_ ^ _2598_ /*20636*/;
assign _2603_ = _2594_ & _2602_ /*20634*/;
assign _2455_ = _2594_ ^ _2602_ /*20635*/;
assign _2600_ = _2601_ | _2603_ /*20632*/;
assign _2605_ = ~Q[26] /*20631*/;
assign _2604_ = _2605_ & D[23] /*20630*/;
assign _2607_ = _2232_ & _2604_ /*20625*/;
assign _2608_ = _2232_ ^ _2604_ /*20628*/;
assign _2609_ = _2600_ & _2608_ /*20626*/;
assign _2456_ = _2600_ ^ _2608_ /*20627*/;
assign _2606_ = _2607_ | _2609_ /*20624*/;
assign _2611_ = ~Q[26] /*20623*/;
assign _2610_ = _2611_ & D[24] /*20622*/;
assign _2613_ = _2233_ & _2610_ /*20617*/;
assign _2614_ = _2233_ ^ _2610_ /*20620*/;
assign _2615_ = _2606_ & _2614_ /*20618*/;
assign _2457_ = _2606_ ^ _2614_ /*20619*/;
assign _2612_ = _2613_ | _2615_ /*20616*/;
assign _2617_ = ~Q[26] /*20615*/;
assign _2616_ = _2617_ & D[25] /*20614*/;
assign _2619_ = _2234_ & _2616_ /*20609*/;
assign _2620_ = _2234_ ^ _2616_ /*20612*/;
assign _2621_ = _2612_ & _2620_ /*20610*/;
assign _2458_ = _2612_ ^ _2620_ /*20611*/;
assign _2618_ = _2619_ | _2621_ /*20608*/;
assign _2623_ = ~Q[26] /*20607*/;
assign _2622_ = _2623_ & D[26] /*20606*/;
assign _2625_ = _2235_ & _2622_ /*20601*/;
assign _2626_ = _2235_ ^ _2622_ /*20604*/;
assign _2627_ = _2618_ & _2626_ /*20602*/;
assign _2459_ = _2618_ ^ _2626_ /*20603*/;
assign _2624_ = _2625_ | _2627_ /*20600*/;
assign _2629_ = ~Q[26] /*20599*/;
assign _2628_ = _2629_ & D[27] /*20598*/;
assign _2631_ = _2236_ & _2628_ /*20593*/;
assign _2632_ = _2236_ ^ _2628_ /*20596*/;
assign _2633_ = _2624_ & _2632_ /*20594*/;
assign _2460_ = _2624_ ^ _2632_ /*20595*/;
assign _2630_ = _2631_ | _2633_ /*20592*/;
assign _2635_ = ~Q[26] /*20591*/;
assign _2634_ = _2635_ & D[28] /*20590*/;
assign _2637_ = _2237_ & _2634_ /*20585*/;
assign _2638_ = _2237_ ^ _2634_ /*20588*/;
assign _2639_ = _2630_ & _2638_ /*20586*/;
assign _2461_ = _2630_ ^ _2638_ /*20587*/;
assign _2636_ = _2637_ | _2639_ /*20584*/;
assign _2641_ = ~Q[26] /*20583*/;
assign _2640_ = _2641_ & D[29] /*20582*/;
assign _2643_ = _2238_ & _2640_ /*20577*/;
assign _2644_ = _2238_ ^ _2640_ /*20580*/;
assign _2645_ = _2636_ & _2644_ /*20578*/;
assign _2462_ = _2636_ ^ _2644_ /*20579*/;
assign _2642_ = _2643_ | _2645_ /*20576*/;
assign _2647_ = ~Q[26] /*20575*/;
assign _2646_ = _2647_ & D[30] /*20574*/;
assign _2649_ = _2239_ & _2646_ /*20569*/;
assign _2650_ = _2239_ ^ _2646_ /*20572*/;
assign _2651_ = _2642_ & _2650_ /*20570*/;
assign _2463_ = _2642_ ^ _2650_ /*20571*/;
assign _2648_ = _2649_ | _2651_ /*20568*/;
assign _2653_ = ~Q[26] /*20567*/;
assign _2652_ = _2653_ & zeroWire /*20566*/;
assign _2654_ = _2240_ ^ _2652_ /*20564*/;
assign _2464_ = _2654_ ^ _2648_ /*20563*/;
assign _2693_ = ~D[0] /*20437*/;
assign _2690_ = R_0[25] & _2693_ /*20433*/;
assign _2691_ = R_0[25] ^ _2693_ /*20436*/;
assign _2692_ = oneWire & _2691_ /*20434*/;
assign _2657_ = oneWire ^ _2691_ /*20435*/;
assign _2689_ = _2690_ | _2692_ /*20432*/;
assign _2698_ = ~D[1] /*20431*/;
assign _2695_ = _2433_ & _2698_ /*20427*/;
assign _2696_ = _2433_ ^ _2698_ /*20430*/;
assign _2697_ = _2689_ & _2696_ /*20428*/;
assign _2658_ = _2689_ ^ _2696_ /*20429*/;
assign _2694_ = _2695_ | _2697_ /*20426*/;
assign _2703_ = ~D[2] /*20425*/;
assign _2700_ = _2434_ & _2703_ /*20421*/;
assign _2701_ = _2434_ ^ _2703_ /*20424*/;
assign _2702_ = _2694_ & _2701_ /*20422*/;
assign _2659_ = _2694_ ^ _2701_ /*20423*/;
assign _2699_ = _2700_ | _2702_ /*20420*/;
assign _2708_ = ~D[3] /*20419*/;
assign _2705_ = _2435_ & _2708_ /*20415*/;
assign _2706_ = _2435_ ^ _2708_ /*20418*/;
assign _2707_ = _2699_ & _2706_ /*20416*/;
assign _2660_ = _2699_ ^ _2706_ /*20417*/;
assign _2704_ = _2705_ | _2707_ /*20414*/;
assign _2713_ = ~D[4] /*20413*/;
assign _2710_ = _2436_ & _2713_ /*20409*/;
assign _2711_ = _2436_ ^ _2713_ /*20412*/;
assign _2712_ = _2704_ & _2711_ /*20410*/;
assign _2661_ = _2704_ ^ _2711_ /*20411*/;
assign _2709_ = _2710_ | _2712_ /*20408*/;
assign _2718_ = ~D[5] /*20407*/;
assign _2715_ = _2437_ & _2718_ /*20403*/;
assign _2716_ = _2437_ ^ _2718_ /*20406*/;
assign _2717_ = _2709_ & _2716_ /*20404*/;
assign _2662_ = _2709_ ^ _2716_ /*20405*/;
assign _2714_ = _2715_ | _2717_ /*20402*/;
assign _2723_ = ~D[6] /*20401*/;
assign _2720_ = _2438_ & _2723_ /*20397*/;
assign _2721_ = _2438_ ^ _2723_ /*20400*/;
assign _2722_ = _2714_ & _2721_ /*20398*/;
assign _2663_ = _2714_ ^ _2721_ /*20399*/;
assign _2719_ = _2720_ | _2722_ /*20396*/;
assign _2728_ = ~D[7] /*20395*/;
assign _2725_ = _2439_ & _2728_ /*20391*/;
assign _2726_ = _2439_ ^ _2728_ /*20394*/;
assign _2727_ = _2719_ & _2726_ /*20392*/;
assign _2664_ = _2719_ ^ _2726_ /*20393*/;
assign _2724_ = _2725_ | _2727_ /*20390*/;
assign _2733_ = ~D[8] /*20389*/;
assign _2730_ = _2440_ & _2733_ /*20385*/;
assign _2731_ = _2440_ ^ _2733_ /*20388*/;
assign _2732_ = _2724_ & _2731_ /*20386*/;
assign _2665_ = _2724_ ^ _2731_ /*20387*/;
assign _2729_ = _2730_ | _2732_ /*20384*/;
assign _2738_ = ~D[9] /*20383*/;
assign _2735_ = _2441_ & _2738_ /*20379*/;
assign _2736_ = _2441_ ^ _2738_ /*20382*/;
assign _2737_ = _2729_ & _2736_ /*20380*/;
assign _2666_ = _2729_ ^ _2736_ /*20381*/;
assign _2734_ = _2735_ | _2737_ /*20378*/;
assign _2743_ = ~D[10] /*20377*/;
assign _2740_ = _2442_ & _2743_ /*20373*/;
assign _2741_ = _2442_ ^ _2743_ /*20376*/;
assign _2742_ = _2734_ & _2741_ /*20374*/;
assign _2667_ = _2734_ ^ _2741_ /*20375*/;
assign _2739_ = _2740_ | _2742_ /*20372*/;
assign _2748_ = ~D[11] /*20371*/;
assign _2745_ = _2443_ & _2748_ /*20367*/;
assign _2746_ = _2443_ ^ _2748_ /*20370*/;
assign _2747_ = _2739_ & _2746_ /*20368*/;
assign _2668_ = _2739_ ^ _2746_ /*20369*/;
assign _2744_ = _2745_ | _2747_ /*20366*/;
assign _2753_ = ~D[12] /*20365*/;
assign _2750_ = _2444_ & _2753_ /*20361*/;
assign _2751_ = _2444_ ^ _2753_ /*20364*/;
assign _2752_ = _2744_ & _2751_ /*20362*/;
assign _2669_ = _2744_ ^ _2751_ /*20363*/;
assign _2749_ = _2750_ | _2752_ /*20360*/;
assign _2758_ = ~D[13] /*20359*/;
assign _2755_ = _2445_ & _2758_ /*20355*/;
assign _2756_ = _2445_ ^ _2758_ /*20358*/;
assign _2757_ = _2749_ & _2756_ /*20356*/;
assign _2670_ = _2749_ ^ _2756_ /*20357*/;
assign _2754_ = _2755_ | _2757_ /*20354*/;
assign _2763_ = ~D[14] /*20353*/;
assign _2760_ = _2446_ & _2763_ /*20349*/;
assign _2761_ = _2446_ ^ _2763_ /*20352*/;
assign _2762_ = _2754_ & _2761_ /*20350*/;
assign _2671_ = _2754_ ^ _2761_ /*20351*/;
assign _2759_ = _2760_ | _2762_ /*20348*/;
assign _2768_ = ~D[15] /*20347*/;
assign _2765_ = _2447_ & _2768_ /*20343*/;
assign _2766_ = _2447_ ^ _2768_ /*20346*/;
assign _2767_ = _2759_ & _2766_ /*20344*/;
assign _2672_ = _2759_ ^ _2766_ /*20345*/;
assign _2764_ = _2765_ | _2767_ /*20342*/;
assign _2773_ = ~D[16] /*20341*/;
assign _2770_ = _2448_ & _2773_ /*20337*/;
assign _2771_ = _2448_ ^ _2773_ /*20340*/;
assign _2772_ = _2764_ & _2771_ /*20338*/;
assign _2673_ = _2764_ ^ _2771_ /*20339*/;
assign _2769_ = _2770_ | _2772_ /*20336*/;
assign _2778_ = ~D[17] /*20335*/;
assign _2775_ = _2449_ & _2778_ /*20331*/;
assign _2776_ = _2449_ ^ _2778_ /*20334*/;
assign _2777_ = _2769_ & _2776_ /*20332*/;
assign _2674_ = _2769_ ^ _2776_ /*20333*/;
assign _2774_ = _2775_ | _2777_ /*20330*/;
assign _2783_ = ~D[18] /*20329*/;
assign _2780_ = _2450_ & _2783_ /*20325*/;
assign _2781_ = _2450_ ^ _2783_ /*20328*/;
assign _2782_ = _2774_ & _2781_ /*20326*/;
assign _2675_ = _2774_ ^ _2781_ /*20327*/;
assign _2779_ = _2780_ | _2782_ /*20324*/;
assign _2788_ = ~D[19] /*20323*/;
assign _2785_ = _2451_ & _2788_ /*20319*/;
assign _2786_ = _2451_ ^ _2788_ /*20322*/;
assign _2787_ = _2779_ & _2786_ /*20320*/;
assign _2676_ = _2779_ ^ _2786_ /*20321*/;
assign _2784_ = _2785_ | _2787_ /*20318*/;
assign _2793_ = ~D[20] /*20317*/;
assign _2790_ = _2452_ & _2793_ /*20313*/;
assign _2791_ = _2452_ ^ _2793_ /*20316*/;
assign _2792_ = _2784_ & _2791_ /*20314*/;
assign _2677_ = _2784_ ^ _2791_ /*20315*/;
assign _2789_ = _2790_ | _2792_ /*20312*/;
assign _2798_ = ~D[21] /*20311*/;
assign _2795_ = _2453_ & _2798_ /*20307*/;
assign _2796_ = _2453_ ^ _2798_ /*20310*/;
assign _2797_ = _2789_ & _2796_ /*20308*/;
assign _2678_ = _2789_ ^ _2796_ /*20309*/;
assign _2794_ = _2795_ | _2797_ /*20306*/;
assign _2803_ = ~D[22] /*20305*/;
assign _2800_ = _2454_ & _2803_ /*20301*/;
assign _2801_ = _2454_ ^ _2803_ /*20304*/;
assign _2802_ = _2794_ & _2801_ /*20302*/;
assign _2679_ = _2794_ ^ _2801_ /*20303*/;
assign _2799_ = _2800_ | _2802_ /*20300*/;
assign _2808_ = ~D[23] /*20299*/;
assign _2805_ = _2455_ & _2808_ /*20295*/;
assign _2806_ = _2455_ ^ _2808_ /*20298*/;
assign _2807_ = _2799_ & _2806_ /*20296*/;
assign _2680_ = _2799_ ^ _2806_ /*20297*/;
assign _2804_ = _2805_ | _2807_ /*20294*/;
assign _2813_ = ~D[24] /*20293*/;
assign _2810_ = _2456_ & _2813_ /*20289*/;
assign _2811_ = _2456_ ^ _2813_ /*20292*/;
assign _2812_ = _2804_ & _2811_ /*20290*/;
assign _2681_ = _2804_ ^ _2811_ /*20291*/;
assign _2809_ = _2810_ | _2812_ /*20288*/;
assign _2818_ = ~D[25] /*20287*/;
assign _2815_ = _2457_ & _2818_ /*20283*/;
assign _2816_ = _2457_ ^ _2818_ /*20286*/;
assign _2817_ = _2809_ & _2816_ /*20284*/;
assign _2682_ = _2809_ ^ _2816_ /*20285*/;
assign _2814_ = _2815_ | _2817_ /*20282*/;
assign _2823_ = ~D[26] /*20281*/;
assign _2820_ = _2458_ & _2823_ /*20277*/;
assign _2821_ = _2458_ ^ _2823_ /*20280*/;
assign _2822_ = _2814_ & _2821_ /*20278*/;
assign _2683_ = _2814_ ^ _2821_ /*20279*/;
assign _2819_ = _2820_ | _2822_ /*20276*/;
assign _2828_ = ~D[27] /*20275*/;
assign _2825_ = _2459_ & _2828_ /*20271*/;
assign _2826_ = _2459_ ^ _2828_ /*20274*/;
assign _2827_ = _2819_ & _2826_ /*20272*/;
assign _2684_ = _2819_ ^ _2826_ /*20273*/;
assign _2824_ = _2825_ | _2827_ /*20270*/;
assign _2833_ = ~D[28] /*20269*/;
assign _2830_ = _2460_ & _2833_ /*20265*/;
assign _2831_ = _2460_ ^ _2833_ /*20268*/;
assign _2832_ = _2824_ & _2831_ /*20266*/;
assign _2685_ = _2824_ ^ _2831_ /*20267*/;
assign _2829_ = _2830_ | _2832_ /*20264*/;
assign _2838_ = ~D[29] /*20263*/;
assign _2835_ = _2461_ & _2838_ /*20259*/;
assign _2836_ = _2461_ ^ _2838_ /*20262*/;
assign _2837_ = _2829_ & _2836_ /*20260*/;
assign _2686_ = _2829_ ^ _2836_ /*20261*/;
assign _2834_ = _2835_ | _2837_ /*20258*/;
assign _2843_ = ~D[30] /*20257*/;
assign _2840_ = _2462_ & _2843_ /*20253*/;
assign _2841_ = _2462_ ^ _2843_ /*20256*/;
assign _2842_ = _2834_ & _2841_ /*20254*/;
assign _2687_ = _2834_ ^ _2841_ /*20255*/;
assign _2839_ = _2840_ | _2842_ /*20252*/;
assign _2844_ = _2463_ & oneWire /*20247*/;
assign _2845_ = _2463_ ^ oneWire /*20250*/;
assign _2846_ = _2839_ & _2845_ /*20248*/;
assign _2688_ = _2839_ ^ _2845_ /*20249*/;
assign Q[25] = _2844_ | _2846_ /*20246*/;
assign _2915_ = ~Q[25] /*20053*/;
assign _2914_ = _2915_ & D[0] /*20052*/;
assign _2917_ = _2657_ & _2914_ /*20047*/;
assign _2918_ = _2657_ ^ _2914_ /*20050*/;
assign _2919_ = zeroWire & _2918_ /*20048*/;
assign _2881_ = zeroWire ^ _2918_ /*20049*/;
assign _2916_ = _2917_ | _2919_ /*20046*/;
assign _2921_ = ~Q[25] /*20045*/;
assign _2920_ = _2921_ & D[1] /*20044*/;
assign _2923_ = _2658_ & _2920_ /*20039*/;
assign _2924_ = _2658_ ^ _2920_ /*20042*/;
assign _2925_ = _2916_ & _2924_ /*20040*/;
assign _2882_ = _2916_ ^ _2924_ /*20041*/;
assign _2922_ = _2923_ | _2925_ /*20038*/;
assign _2927_ = ~Q[25] /*20037*/;
assign _2926_ = _2927_ & D[2] /*20036*/;
assign _2929_ = _2659_ & _2926_ /*20031*/;
assign _2930_ = _2659_ ^ _2926_ /*20034*/;
assign _2931_ = _2922_ & _2930_ /*20032*/;
assign _2883_ = _2922_ ^ _2930_ /*20033*/;
assign _2928_ = _2929_ | _2931_ /*20030*/;
assign _2933_ = ~Q[25] /*20029*/;
assign _2932_ = _2933_ & D[3] /*20028*/;
assign _2935_ = _2660_ & _2932_ /*20023*/;
assign _2936_ = _2660_ ^ _2932_ /*20026*/;
assign _2937_ = _2928_ & _2936_ /*20024*/;
assign _2884_ = _2928_ ^ _2936_ /*20025*/;
assign _2934_ = _2935_ | _2937_ /*20022*/;
assign _2939_ = ~Q[25] /*20021*/;
assign _2938_ = _2939_ & D[4] /*20020*/;
assign _2941_ = _2661_ & _2938_ /*20015*/;
assign _2942_ = _2661_ ^ _2938_ /*20018*/;
assign _2943_ = _2934_ & _2942_ /*20016*/;
assign _2885_ = _2934_ ^ _2942_ /*20017*/;
assign _2940_ = _2941_ | _2943_ /*20014*/;
assign _2945_ = ~Q[25] /*20013*/;
assign _2944_ = _2945_ & D[5] /*20012*/;
assign _2947_ = _2662_ & _2944_ /*20007*/;
assign _2948_ = _2662_ ^ _2944_ /*20010*/;
assign _2949_ = _2940_ & _2948_ /*20008*/;
assign _2886_ = _2940_ ^ _2948_ /*20009*/;
assign _2946_ = _2947_ | _2949_ /*20006*/;
assign _2951_ = ~Q[25] /*20005*/;
assign _2950_ = _2951_ & D[6] /*20004*/;
assign _2953_ = _2663_ & _2950_ /*19999*/;
assign _2954_ = _2663_ ^ _2950_ /*20002*/;
assign _2955_ = _2946_ & _2954_ /*20000*/;
assign _2887_ = _2946_ ^ _2954_ /*20001*/;
assign _2952_ = _2953_ | _2955_ /*19998*/;
assign _2957_ = ~Q[25] /*19997*/;
assign _2956_ = _2957_ & D[7] /*19996*/;
assign _2959_ = _2664_ & _2956_ /*19991*/;
assign _2960_ = _2664_ ^ _2956_ /*19994*/;
assign _2961_ = _2952_ & _2960_ /*19992*/;
assign _2888_ = _2952_ ^ _2960_ /*19993*/;
assign _2958_ = _2959_ | _2961_ /*19990*/;
assign _2963_ = ~Q[25] /*19989*/;
assign _2962_ = _2963_ & D[8] /*19988*/;
assign _2965_ = _2665_ & _2962_ /*19983*/;
assign _2966_ = _2665_ ^ _2962_ /*19986*/;
assign _2967_ = _2958_ & _2966_ /*19984*/;
assign _2889_ = _2958_ ^ _2966_ /*19985*/;
assign _2964_ = _2965_ | _2967_ /*19982*/;
assign _2969_ = ~Q[25] /*19981*/;
assign _2968_ = _2969_ & D[9] /*19980*/;
assign _2971_ = _2666_ & _2968_ /*19975*/;
assign _2972_ = _2666_ ^ _2968_ /*19978*/;
assign _2973_ = _2964_ & _2972_ /*19976*/;
assign _2890_ = _2964_ ^ _2972_ /*19977*/;
assign _2970_ = _2971_ | _2973_ /*19974*/;
assign _2975_ = ~Q[25] /*19973*/;
assign _2974_ = _2975_ & D[10] /*19972*/;
assign _2977_ = _2667_ & _2974_ /*19967*/;
assign _2978_ = _2667_ ^ _2974_ /*19970*/;
assign _2979_ = _2970_ & _2978_ /*19968*/;
assign _2891_ = _2970_ ^ _2978_ /*19969*/;
assign _2976_ = _2977_ | _2979_ /*19966*/;
assign _2981_ = ~Q[25] /*19965*/;
assign _2980_ = _2981_ & D[11] /*19964*/;
assign _2983_ = _2668_ & _2980_ /*19959*/;
assign _2984_ = _2668_ ^ _2980_ /*19962*/;
assign _2985_ = _2976_ & _2984_ /*19960*/;
assign _2892_ = _2976_ ^ _2984_ /*19961*/;
assign _2982_ = _2983_ | _2985_ /*19958*/;
assign _2987_ = ~Q[25] /*19957*/;
assign _2986_ = _2987_ & D[12] /*19956*/;
assign _2989_ = _2669_ & _2986_ /*19951*/;
assign _2990_ = _2669_ ^ _2986_ /*19954*/;
assign _2991_ = _2982_ & _2990_ /*19952*/;
assign _2893_ = _2982_ ^ _2990_ /*19953*/;
assign _2988_ = _2989_ | _2991_ /*19950*/;
assign _2993_ = ~Q[25] /*19949*/;
assign _2992_ = _2993_ & D[13] /*19948*/;
assign _2995_ = _2670_ & _2992_ /*19943*/;
assign _2996_ = _2670_ ^ _2992_ /*19946*/;
assign _2997_ = _2988_ & _2996_ /*19944*/;
assign _2894_ = _2988_ ^ _2996_ /*19945*/;
assign _2994_ = _2995_ | _2997_ /*19942*/;
assign _2999_ = ~Q[25] /*19941*/;
assign _2998_ = _2999_ & D[14] /*19940*/;
assign _3001_ = _2671_ & _2998_ /*19935*/;
assign _3002_ = _2671_ ^ _2998_ /*19938*/;
assign _3003_ = _2994_ & _3002_ /*19936*/;
assign _2895_ = _2994_ ^ _3002_ /*19937*/;
assign _3000_ = _3001_ | _3003_ /*19934*/;
assign _3005_ = ~Q[25] /*19933*/;
assign _3004_ = _3005_ & D[15] /*19932*/;
assign _3007_ = _2672_ & _3004_ /*19927*/;
assign _3008_ = _2672_ ^ _3004_ /*19930*/;
assign _3009_ = _3000_ & _3008_ /*19928*/;
assign _2896_ = _3000_ ^ _3008_ /*19929*/;
assign _3006_ = _3007_ | _3009_ /*19926*/;
assign _3011_ = ~Q[25] /*19925*/;
assign _3010_ = _3011_ & D[16] /*19924*/;
assign _3013_ = _2673_ & _3010_ /*19919*/;
assign _3014_ = _2673_ ^ _3010_ /*19922*/;
assign _3015_ = _3006_ & _3014_ /*19920*/;
assign _2897_ = _3006_ ^ _3014_ /*19921*/;
assign _3012_ = _3013_ | _3015_ /*19918*/;
assign _3017_ = ~Q[25] /*19917*/;
assign _3016_ = _3017_ & D[17] /*19916*/;
assign _3019_ = _2674_ & _3016_ /*19911*/;
assign _3020_ = _2674_ ^ _3016_ /*19914*/;
assign _3021_ = _3012_ & _3020_ /*19912*/;
assign _2898_ = _3012_ ^ _3020_ /*19913*/;
assign _3018_ = _3019_ | _3021_ /*19910*/;
assign _3023_ = ~Q[25] /*19909*/;
assign _3022_ = _3023_ & D[18] /*19908*/;
assign _3025_ = _2675_ & _3022_ /*19903*/;
assign _3026_ = _2675_ ^ _3022_ /*19906*/;
assign _3027_ = _3018_ & _3026_ /*19904*/;
assign _2899_ = _3018_ ^ _3026_ /*19905*/;
assign _3024_ = _3025_ | _3027_ /*19902*/;
assign _3029_ = ~Q[25] /*19901*/;
assign _3028_ = _3029_ & D[19] /*19900*/;
assign _3031_ = _2676_ & _3028_ /*19895*/;
assign _3032_ = _2676_ ^ _3028_ /*19898*/;
assign _3033_ = _3024_ & _3032_ /*19896*/;
assign _2900_ = _3024_ ^ _3032_ /*19897*/;
assign _3030_ = _3031_ | _3033_ /*19894*/;
assign _3035_ = ~Q[25] /*19893*/;
assign _3034_ = _3035_ & D[20] /*19892*/;
assign _3037_ = _2677_ & _3034_ /*19887*/;
assign _3038_ = _2677_ ^ _3034_ /*19890*/;
assign _3039_ = _3030_ & _3038_ /*19888*/;
assign _2901_ = _3030_ ^ _3038_ /*19889*/;
assign _3036_ = _3037_ | _3039_ /*19886*/;
assign _3041_ = ~Q[25] /*19885*/;
assign _3040_ = _3041_ & D[21] /*19884*/;
assign _3043_ = _2678_ & _3040_ /*19879*/;
assign _3044_ = _2678_ ^ _3040_ /*19882*/;
assign _3045_ = _3036_ & _3044_ /*19880*/;
assign _2902_ = _3036_ ^ _3044_ /*19881*/;
assign _3042_ = _3043_ | _3045_ /*19878*/;
assign _3047_ = ~Q[25] /*19877*/;
assign _3046_ = _3047_ & D[22] /*19876*/;
assign _3049_ = _2679_ & _3046_ /*19871*/;
assign _3050_ = _2679_ ^ _3046_ /*19874*/;
assign _3051_ = _3042_ & _3050_ /*19872*/;
assign _2903_ = _3042_ ^ _3050_ /*19873*/;
assign _3048_ = _3049_ | _3051_ /*19870*/;
assign _3053_ = ~Q[25] /*19869*/;
assign _3052_ = _3053_ & D[23] /*19868*/;
assign _3055_ = _2680_ & _3052_ /*19863*/;
assign _3056_ = _2680_ ^ _3052_ /*19866*/;
assign _3057_ = _3048_ & _3056_ /*19864*/;
assign _2904_ = _3048_ ^ _3056_ /*19865*/;
assign _3054_ = _3055_ | _3057_ /*19862*/;
assign _3059_ = ~Q[25] /*19861*/;
assign _3058_ = _3059_ & D[24] /*19860*/;
assign _3061_ = _2681_ & _3058_ /*19855*/;
assign _3062_ = _2681_ ^ _3058_ /*19858*/;
assign _3063_ = _3054_ & _3062_ /*19856*/;
assign _2905_ = _3054_ ^ _3062_ /*19857*/;
assign _3060_ = _3061_ | _3063_ /*19854*/;
assign _3065_ = ~Q[25] /*19853*/;
assign _3064_ = _3065_ & D[25] /*19852*/;
assign _3067_ = _2682_ & _3064_ /*19847*/;
assign _3068_ = _2682_ ^ _3064_ /*19850*/;
assign _3069_ = _3060_ & _3068_ /*19848*/;
assign _2906_ = _3060_ ^ _3068_ /*19849*/;
assign _3066_ = _3067_ | _3069_ /*19846*/;
assign _3071_ = ~Q[25] /*19845*/;
assign _3070_ = _3071_ & D[26] /*19844*/;
assign _3073_ = _2683_ & _3070_ /*19839*/;
assign _3074_ = _2683_ ^ _3070_ /*19842*/;
assign _3075_ = _3066_ & _3074_ /*19840*/;
assign _2907_ = _3066_ ^ _3074_ /*19841*/;
assign _3072_ = _3073_ | _3075_ /*19838*/;
assign _3077_ = ~Q[25] /*19837*/;
assign _3076_ = _3077_ & D[27] /*19836*/;
assign _3079_ = _2684_ & _3076_ /*19831*/;
assign _3080_ = _2684_ ^ _3076_ /*19834*/;
assign _3081_ = _3072_ & _3080_ /*19832*/;
assign _2908_ = _3072_ ^ _3080_ /*19833*/;
assign _3078_ = _3079_ | _3081_ /*19830*/;
assign _3083_ = ~Q[25] /*19829*/;
assign _3082_ = _3083_ & D[28] /*19828*/;
assign _3085_ = _2685_ & _3082_ /*19823*/;
assign _3086_ = _2685_ ^ _3082_ /*19826*/;
assign _3087_ = _3078_ & _3086_ /*19824*/;
assign _2909_ = _3078_ ^ _3086_ /*19825*/;
assign _3084_ = _3085_ | _3087_ /*19822*/;
assign _3089_ = ~Q[25] /*19821*/;
assign _3088_ = _3089_ & D[29] /*19820*/;
assign _3091_ = _2686_ & _3088_ /*19815*/;
assign _3092_ = _2686_ ^ _3088_ /*19818*/;
assign _3093_ = _3084_ & _3092_ /*19816*/;
assign _2910_ = _3084_ ^ _3092_ /*19817*/;
assign _3090_ = _3091_ | _3093_ /*19814*/;
assign _3095_ = ~Q[25] /*19813*/;
assign _3094_ = _3095_ & D[30] /*19812*/;
assign _3097_ = _2687_ & _3094_ /*19807*/;
assign _3098_ = _2687_ ^ _3094_ /*19810*/;
assign _3099_ = _3090_ & _3098_ /*19808*/;
assign _2911_ = _3090_ ^ _3098_ /*19809*/;
assign _3096_ = _3097_ | _3099_ /*19806*/;
assign _3101_ = ~Q[25] /*19805*/;
assign _3100_ = _3101_ & zeroWire /*19804*/;
assign _3102_ = _2688_ ^ _3100_ /*19802*/;
assign _2912_ = _3102_ ^ _3096_ /*19801*/;
assign _3141_ = ~D[0] /*19675*/;
assign _3138_ = R_0[24] & _3141_ /*19671*/;
assign _3139_ = R_0[24] ^ _3141_ /*19674*/;
assign _3140_ = oneWire & _3139_ /*19672*/;
assign _3105_ = oneWire ^ _3139_ /*19673*/;
assign _3137_ = _3138_ | _3140_ /*19670*/;
assign _3146_ = ~D[1] /*19669*/;
assign _3143_ = _2881_ & _3146_ /*19665*/;
assign _3144_ = _2881_ ^ _3146_ /*19668*/;
assign _3145_ = _3137_ & _3144_ /*19666*/;
assign _3106_ = _3137_ ^ _3144_ /*19667*/;
assign _3142_ = _3143_ | _3145_ /*19664*/;
assign _3151_ = ~D[2] /*19663*/;
assign _3148_ = _2882_ & _3151_ /*19659*/;
assign _3149_ = _2882_ ^ _3151_ /*19662*/;
assign _3150_ = _3142_ & _3149_ /*19660*/;
assign _3107_ = _3142_ ^ _3149_ /*19661*/;
assign _3147_ = _3148_ | _3150_ /*19658*/;
assign _3156_ = ~D[3] /*19657*/;
assign _3153_ = _2883_ & _3156_ /*19653*/;
assign _3154_ = _2883_ ^ _3156_ /*19656*/;
assign _3155_ = _3147_ & _3154_ /*19654*/;
assign _3108_ = _3147_ ^ _3154_ /*19655*/;
assign _3152_ = _3153_ | _3155_ /*19652*/;
assign _3161_ = ~D[4] /*19651*/;
assign _3158_ = _2884_ & _3161_ /*19647*/;
assign _3159_ = _2884_ ^ _3161_ /*19650*/;
assign _3160_ = _3152_ & _3159_ /*19648*/;
assign _3109_ = _3152_ ^ _3159_ /*19649*/;
assign _3157_ = _3158_ | _3160_ /*19646*/;
assign _3166_ = ~D[5] /*19645*/;
assign _3163_ = _2885_ & _3166_ /*19641*/;
assign _3164_ = _2885_ ^ _3166_ /*19644*/;
assign _3165_ = _3157_ & _3164_ /*19642*/;
assign _3110_ = _3157_ ^ _3164_ /*19643*/;
assign _3162_ = _3163_ | _3165_ /*19640*/;
assign _3171_ = ~D[6] /*19639*/;
assign _3168_ = _2886_ & _3171_ /*19635*/;
assign _3169_ = _2886_ ^ _3171_ /*19638*/;
assign _3170_ = _3162_ & _3169_ /*19636*/;
assign _3111_ = _3162_ ^ _3169_ /*19637*/;
assign _3167_ = _3168_ | _3170_ /*19634*/;
assign _3176_ = ~D[7] /*19633*/;
assign _3173_ = _2887_ & _3176_ /*19629*/;
assign _3174_ = _2887_ ^ _3176_ /*19632*/;
assign _3175_ = _3167_ & _3174_ /*19630*/;
assign _3112_ = _3167_ ^ _3174_ /*19631*/;
assign _3172_ = _3173_ | _3175_ /*19628*/;
assign _3181_ = ~D[8] /*19627*/;
assign _3178_ = _2888_ & _3181_ /*19623*/;
assign _3179_ = _2888_ ^ _3181_ /*19626*/;
assign _3180_ = _3172_ & _3179_ /*19624*/;
assign _3113_ = _3172_ ^ _3179_ /*19625*/;
assign _3177_ = _3178_ | _3180_ /*19622*/;
assign _3186_ = ~D[9] /*19621*/;
assign _3183_ = _2889_ & _3186_ /*19617*/;
assign _3184_ = _2889_ ^ _3186_ /*19620*/;
assign _3185_ = _3177_ & _3184_ /*19618*/;
assign _3114_ = _3177_ ^ _3184_ /*19619*/;
assign _3182_ = _3183_ | _3185_ /*19616*/;
assign _3191_ = ~D[10] /*19615*/;
assign _3188_ = _2890_ & _3191_ /*19611*/;
assign _3189_ = _2890_ ^ _3191_ /*19614*/;
assign _3190_ = _3182_ & _3189_ /*19612*/;
assign _3115_ = _3182_ ^ _3189_ /*19613*/;
assign _3187_ = _3188_ | _3190_ /*19610*/;
assign _3196_ = ~D[11] /*19609*/;
assign _3193_ = _2891_ & _3196_ /*19605*/;
assign _3194_ = _2891_ ^ _3196_ /*19608*/;
assign _3195_ = _3187_ & _3194_ /*19606*/;
assign _3116_ = _3187_ ^ _3194_ /*19607*/;
assign _3192_ = _3193_ | _3195_ /*19604*/;
assign _3201_ = ~D[12] /*19603*/;
assign _3198_ = _2892_ & _3201_ /*19599*/;
assign _3199_ = _2892_ ^ _3201_ /*19602*/;
assign _3200_ = _3192_ & _3199_ /*19600*/;
assign _3117_ = _3192_ ^ _3199_ /*19601*/;
assign _3197_ = _3198_ | _3200_ /*19598*/;
assign _3206_ = ~D[13] /*19597*/;
assign _3203_ = _2893_ & _3206_ /*19593*/;
assign _3204_ = _2893_ ^ _3206_ /*19596*/;
assign _3205_ = _3197_ & _3204_ /*19594*/;
assign _3118_ = _3197_ ^ _3204_ /*19595*/;
assign _3202_ = _3203_ | _3205_ /*19592*/;
assign _3211_ = ~D[14] /*19591*/;
assign _3208_ = _2894_ & _3211_ /*19587*/;
assign _3209_ = _2894_ ^ _3211_ /*19590*/;
assign _3210_ = _3202_ & _3209_ /*19588*/;
assign _3119_ = _3202_ ^ _3209_ /*19589*/;
assign _3207_ = _3208_ | _3210_ /*19586*/;
assign _3216_ = ~D[15] /*19585*/;
assign _3213_ = _2895_ & _3216_ /*19581*/;
assign _3214_ = _2895_ ^ _3216_ /*19584*/;
assign _3215_ = _3207_ & _3214_ /*19582*/;
assign _3120_ = _3207_ ^ _3214_ /*19583*/;
assign _3212_ = _3213_ | _3215_ /*19580*/;
assign _3221_ = ~D[16] /*19579*/;
assign _3218_ = _2896_ & _3221_ /*19575*/;
assign _3219_ = _2896_ ^ _3221_ /*19578*/;
assign _3220_ = _3212_ & _3219_ /*19576*/;
assign _3121_ = _3212_ ^ _3219_ /*19577*/;
assign _3217_ = _3218_ | _3220_ /*19574*/;
assign _3226_ = ~D[17] /*19573*/;
assign _3223_ = _2897_ & _3226_ /*19569*/;
assign _3224_ = _2897_ ^ _3226_ /*19572*/;
assign _3225_ = _3217_ & _3224_ /*19570*/;
assign _3122_ = _3217_ ^ _3224_ /*19571*/;
assign _3222_ = _3223_ | _3225_ /*19568*/;
assign _3231_ = ~D[18] /*19567*/;
assign _3228_ = _2898_ & _3231_ /*19563*/;
assign _3229_ = _2898_ ^ _3231_ /*19566*/;
assign _3230_ = _3222_ & _3229_ /*19564*/;
assign _3123_ = _3222_ ^ _3229_ /*19565*/;
assign _3227_ = _3228_ | _3230_ /*19562*/;
assign _3236_ = ~D[19] /*19561*/;
assign _3233_ = _2899_ & _3236_ /*19557*/;
assign _3234_ = _2899_ ^ _3236_ /*19560*/;
assign _3235_ = _3227_ & _3234_ /*19558*/;
assign _3124_ = _3227_ ^ _3234_ /*19559*/;
assign _3232_ = _3233_ | _3235_ /*19556*/;
assign _3241_ = ~D[20] /*19555*/;
assign _3238_ = _2900_ & _3241_ /*19551*/;
assign _3239_ = _2900_ ^ _3241_ /*19554*/;
assign _3240_ = _3232_ & _3239_ /*19552*/;
assign _3125_ = _3232_ ^ _3239_ /*19553*/;
assign _3237_ = _3238_ | _3240_ /*19550*/;
assign _3246_ = ~D[21] /*19549*/;
assign _3243_ = _2901_ & _3246_ /*19545*/;
assign _3244_ = _2901_ ^ _3246_ /*19548*/;
assign _3245_ = _3237_ & _3244_ /*19546*/;
assign _3126_ = _3237_ ^ _3244_ /*19547*/;
assign _3242_ = _3243_ | _3245_ /*19544*/;
assign _3251_ = ~D[22] /*19543*/;
assign _3248_ = _2902_ & _3251_ /*19539*/;
assign _3249_ = _2902_ ^ _3251_ /*19542*/;
assign _3250_ = _3242_ & _3249_ /*19540*/;
assign _3127_ = _3242_ ^ _3249_ /*19541*/;
assign _3247_ = _3248_ | _3250_ /*19538*/;
assign _3256_ = ~D[23] /*19537*/;
assign _3253_ = _2903_ & _3256_ /*19533*/;
assign _3254_ = _2903_ ^ _3256_ /*19536*/;
assign _3255_ = _3247_ & _3254_ /*19534*/;
assign _3128_ = _3247_ ^ _3254_ /*19535*/;
assign _3252_ = _3253_ | _3255_ /*19532*/;
assign _3261_ = ~D[24] /*19531*/;
assign _3258_ = _2904_ & _3261_ /*19527*/;
assign _3259_ = _2904_ ^ _3261_ /*19530*/;
assign _3260_ = _3252_ & _3259_ /*19528*/;
assign _3129_ = _3252_ ^ _3259_ /*19529*/;
assign _3257_ = _3258_ | _3260_ /*19526*/;
assign _3266_ = ~D[25] /*19525*/;
assign _3263_ = _2905_ & _3266_ /*19521*/;
assign _3264_ = _2905_ ^ _3266_ /*19524*/;
assign _3265_ = _3257_ & _3264_ /*19522*/;
assign _3130_ = _3257_ ^ _3264_ /*19523*/;
assign _3262_ = _3263_ | _3265_ /*19520*/;
assign _3271_ = ~D[26] /*19519*/;
assign _3268_ = _2906_ & _3271_ /*19515*/;
assign _3269_ = _2906_ ^ _3271_ /*19518*/;
assign _3270_ = _3262_ & _3269_ /*19516*/;
assign _3131_ = _3262_ ^ _3269_ /*19517*/;
assign _3267_ = _3268_ | _3270_ /*19514*/;
assign _3276_ = ~D[27] /*19513*/;
assign _3273_ = _2907_ & _3276_ /*19509*/;
assign _3274_ = _2907_ ^ _3276_ /*19512*/;
assign _3275_ = _3267_ & _3274_ /*19510*/;
assign _3132_ = _3267_ ^ _3274_ /*19511*/;
assign _3272_ = _3273_ | _3275_ /*19508*/;
assign _3281_ = ~D[28] /*19507*/;
assign _3278_ = _2908_ & _3281_ /*19503*/;
assign _3279_ = _2908_ ^ _3281_ /*19506*/;
assign _3280_ = _3272_ & _3279_ /*19504*/;
assign _3133_ = _3272_ ^ _3279_ /*19505*/;
assign _3277_ = _3278_ | _3280_ /*19502*/;
assign _3286_ = ~D[29] /*19501*/;
assign _3283_ = _2909_ & _3286_ /*19497*/;
assign _3284_ = _2909_ ^ _3286_ /*19500*/;
assign _3285_ = _3277_ & _3284_ /*19498*/;
assign _3134_ = _3277_ ^ _3284_ /*19499*/;
assign _3282_ = _3283_ | _3285_ /*19496*/;
assign _3291_ = ~D[30] /*19495*/;
assign _3288_ = _2910_ & _3291_ /*19491*/;
assign _3289_ = _2910_ ^ _3291_ /*19494*/;
assign _3290_ = _3282_ & _3289_ /*19492*/;
assign _3135_ = _3282_ ^ _3289_ /*19493*/;
assign _3287_ = _3288_ | _3290_ /*19490*/;
assign _3292_ = _2911_ & oneWire /*19485*/;
assign _3293_ = _2911_ ^ oneWire /*19488*/;
assign _3294_ = _3287_ & _3293_ /*19486*/;
assign _3136_ = _3287_ ^ _3293_ /*19487*/;
assign Q[24] = _3292_ | _3294_ /*19484*/;
assign _3363_ = ~Q[24] /*19291*/;
assign _3362_ = _3363_ & D[0] /*19290*/;
assign _3365_ = _3105_ & _3362_ /*19285*/;
assign _3366_ = _3105_ ^ _3362_ /*19288*/;
assign _3367_ = zeroWire & _3366_ /*19286*/;
assign _3329_ = zeroWire ^ _3366_ /*19287*/;
assign _3364_ = _3365_ | _3367_ /*19284*/;
assign _3369_ = ~Q[24] /*19283*/;
assign _3368_ = _3369_ & D[1] /*19282*/;
assign _3371_ = _3106_ & _3368_ /*19277*/;
assign _3372_ = _3106_ ^ _3368_ /*19280*/;
assign _3373_ = _3364_ & _3372_ /*19278*/;
assign _3330_ = _3364_ ^ _3372_ /*19279*/;
assign _3370_ = _3371_ | _3373_ /*19276*/;
assign _3375_ = ~Q[24] /*19275*/;
assign _3374_ = _3375_ & D[2] /*19274*/;
assign _3377_ = _3107_ & _3374_ /*19269*/;
assign _3378_ = _3107_ ^ _3374_ /*19272*/;
assign _3379_ = _3370_ & _3378_ /*19270*/;
assign _3331_ = _3370_ ^ _3378_ /*19271*/;
assign _3376_ = _3377_ | _3379_ /*19268*/;
assign _3381_ = ~Q[24] /*19267*/;
assign _3380_ = _3381_ & D[3] /*19266*/;
assign _3383_ = _3108_ & _3380_ /*19261*/;
assign _3384_ = _3108_ ^ _3380_ /*19264*/;
assign _3385_ = _3376_ & _3384_ /*19262*/;
assign _3332_ = _3376_ ^ _3384_ /*19263*/;
assign _3382_ = _3383_ | _3385_ /*19260*/;
assign _3387_ = ~Q[24] /*19259*/;
assign _3386_ = _3387_ & D[4] /*19258*/;
assign _3389_ = _3109_ & _3386_ /*19253*/;
assign _3390_ = _3109_ ^ _3386_ /*19256*/;
assign _3391_ = _3382_ & _3390_ /*19254*/;
assign _3333_ = _3382_ ^ _3390_ /*19255*/;
assign _3388_ = _3389_ | _3391_ /*19252*/;
assign _3393_ = ~Q[24] /*19251*/;
assign _3392_ = _3393_ & D[5] /*19250*/;
assign _3395_ = _3110_ & _3392_ /*19245*/;
assign _3396_ = _3110_ ^ _3392_ /*19248*/;
assign _3397_ = _3388_ & _3396_ /*19246*/;
assign _3334_ = _3388_ ^ _3396_ /*19247*/;
assign _3394_ = _3395_ | _3397_ /*19244*/;
assign _3399_ = ~Q[24] /*19243*/;
assign _3398_ = _3399_ & D[6] /*19242*/;
assign _3401_ = _3111_ & _3398_ /*19237*/;
assign _3402_ = _3111_ ^ _3398_ /*19240*/;
assign _3403_ = _3394_ & _3402_ /*19238*/;
assign _3335_ = _3394_ ^ _3402_ /*19239*/;
assign _3400_ = _3401_ | _3403_ /*19236*/;
assign _3405_ = ~Q[24] /*19235*/;
assign _3404_ = _3405_ & D[7] /*19234*/;
assign _3407_ = _3112_ & _3404_ /*19229*/;
assign _3408_ = _3112_ ^ _3404_ /*19232*/;
assign _3409_ = _3400_ & _3408_ /*19230*/;
assign _3336_ = _3400_ ^ _3408_ /*19231*/;
assign _3406_ = _3407_ | _3409_ /*19228*/;
assign _3411_ = ~Q[24] /*19227*/;
assign _3410_ = _3411_ & D[8] /*19226*/;
assign _3413_ = _3113_ & _3410_ /*19221*/;
assign _3414_ = _3113_ ^ _3410_ /*19224*/;
assign _3415_ = _3406_ & _3414_ /*19222*/;
assign _3337_ = _3406_ ^ _3414_ /*19223*/;
assign _3412_ = _3413_ | _3415_ /*19220*/;
assign _3417_ = ~Q[24] /*19219*/;
assign _3416_ = _3417_ & D[9] /*19218*/;
assign _3419_ = _3114_ & _3416_ /*19213*/;
assign _3420_ = _3114_ ^ _3416_ /*19216*/;
assign _3421_ = _3412_ & _3420_ /*19214*/;
assign _3338_ = _3412_ ^ _3420_ /*19215*/;
assign _3418_ = _3419_ | _3421_ /*19212*/;
assign _3423_ = ~Q[24] /*19211*/;
assign _3422_ = _3423_ & D[10] /*19210*/;
assign _3425_ = _3115_ & _3422_ /*19205*/;
assign _3426_ = _3115_ ^ _3422_ /*19208*/;
assign _3427_ = _3418_ & _3426_ /*19206*/;
assign _3339_ = _3418_ ^ _3426_ /*19207*/;
assign _3424_ = _3425_ | _3427_ /*19204*/;
assign _3429_ = ~Q[24] /*19203*/;
assign _3428_ = _3429_ & D[11] /*19202*/;
assign _3431_ = _3116_ & _3428_ /*19197*/;
assign _3432_ = _3116_ ^ _3428_ /*19200*/;
assign _3433_ = _3424_ & _3432_ /*19198*/;
assign _3340_ = _3424_ ^ _3432_ /*19199*/;
assign _3430_ = _3431_ | _3433_ /*19196*/;
assign _3435_ = ~Q[24] /*19195*/;
assign _3434_ = _3435_ & D[12] /*19194*/;
assign _3437_ = _3117_ & _3434_ /*19189*/;
assign _3438_ = _3117_ ^ _3434_ /*19192*/;
assign _3439_ = _3430_ & _3438_ /*19190*/;
assign _3341_ = _3430_ ^ _3438_ /*19191*/;
assign _3436_ = _3437_ | _3439_ /*19188*/;
assign _3441_ = ~Q[24] /*19187*/;
assign _3440_ = _3441_ & D[13] /*19186*/;
assign _3443_ = _3118_ & _3440_ /*19181*/;
assign _3444_ = _3118_ ^ _3440_ /*19184*/;
assign _3445_ = _3436_ & _3444_ /*19182*/;
assign _3342_ = _3436_ ^ _3444_ /*19183*/;
assign _3442_ = _3443_ | _3445_ /*19180*/;
assign _3447_ = ~Q[24] /*19179*/;
assign _3446_ = _3447_ & D[14] /*19178*/;
assign _3449_ = _3119_ & _3446_ /*19173*/;
assign _3450_ = _3119_ ^ _3446_ /*19176*/;
assign _3451_ = _3442_ & _3450_ /*19174*/;
assign _3343_ = _3442_ ^ _3450_ /*19175*/;
assign _3448_ = _3449_ | _3451_ /*19172*/;
assign _3453_ = ~Q[24] /*19171*/;
assign _3452_ = _3453_ & D[15] /*19170*/;
assign _3455_ = _3120_ & _3452_ /*19165*/;
assign _3456_ = _3120_ ^ _3452_ /*19168*/;
assign _3457_ = _3448_ & _3456_ /*19166*/;
assign _3344_ = _3448_ ^ _3456_ /*19167*/;
assign _3454_ = _3455_ | _3457_ /*19164*/;
assign _3459_ = ~Q[24] /*19163*/;
assign _3458_ = _3459_ & D[16] /*19162*/;
assign _3461_ = _3121_ & _3458_ /*19157*/;
assign _3462_ = _3121_ ^ _3458_ /*19160*/;
assign _3463_ = _3454_ & _3462_ /*19158*/;
assign _3345_ = _3454_ ^ _3462_ /*19159*/;
assign _3460_ = _3461_ | _3463_ /*19156*/;
assign _3465_ = ~Q[24] /*19155*/;
assign _3464_ = _3465_ & D[17] /*19154*/;
assign _3467_ = _3122_ & _3464_ /*19149*/;
assign _3468_ = _3122_ ^ _3464_ /*19152*/;
assign _3469_ = _3460_ & _3468_ /*19150*/;
assign _3346_ = _3460_ ^ _3468_ /*19151*/;
assign _3466_ = _3467_ | _3469_ /*19148*/;
assign _3471_ = ~Q[24] /*19147*/;
assign _3470_ = _3471_ & D[18] /*19146*/;
assign _3473_ = _3123_ & _3470_ /*19141*/;
assign _3474_ = _3123_ ^ _3470_ /*19144*/;
assign _3475_ = _3466_ & _3474_ /*19142*/;
assign _3347_ = _3466_ ^ _3474_ /*19143*/;
assign _3472_ = _3473_ | _3475_ /*19140*/;
assign _3477_ = ~Q[24] /*19139*/;
assign _3476_ = _3477_ & D[19] /*19138*/;
assign _3479_ = _3124_ & _3476_ /*19133*/;
assign _3480_ = _3124_ ^ _3476_ /*19136*/;
assign _3481_ = _3472_ & _3480_ /*19134*/;
assign _3348_ = _3472_ ^ _3480_ /*19135*/;
assign _3478_ = _3479_ | _3481_ /*19132*/;
assign _3483_ = ~Q[24] /*19131*/;
assign _3482_ = _3483_ & D[20] /*19130*/;
assign _3485_ = _3125_ & _3482_ /*19125*/;
assign _3486_ = _3125_ ^ _3482_ /*19128*/;
assign _3487_ = _3478_ & _3486_ /*19126*/;
assign _3349_ = _3478_ ^ _3486_ /*19127*/;
assign _3484_ = _3485_ | _3487_ /*19124*/;
assign _3489_ = ~Q[24] /*19123*/;
assign _3488_ = _3489_ & D[21] /*19122*/;
assign _3491_ = _3126_ & _3488_ /*19117*/;
assign _3492_ = _3126_ ^ _3488_ /*19120*/;
assign _3493_ = _3484_ & _3492_ /*19118*/;
assign _3350_ = _3484_ ^ _3492_ /*19119*/;
assign _3490_ = _3491_ | _3493_ /*19116*/;
assign _3495_ = ~Q[24] /*19115*/;
assign _3494_ = _3495_ & D[22] /*19114*/;
assign _3497_ = _3127_ & _3494_ /*19109*/;
assign _3498_ = _3127_ ^ _3494_ /*19112*/;
assign _3499_ = _3490_ & _3498_ /*19110*/;
assign _3351_ = _3490_ ^ _3498_ /*19111*/;
assign _3496_ = _3497_ | _3499_ /*19108*/;
assign _3501_ = ~Q[24] /*19107*/;
assign _3500_ = _3501_ & D[23] /*19106*/;
assign _3503_ = _3128_ & _3500_ /*19101*/;
assign _3504_ = _3128_ ^ _3500_ /*19104*/;
assign _3505_ = _3496_ & _3504_ /*19102*/;
assign _3352_ = _3496_ ^ _3504_ /*19103*/;
assign _3502_ = _3503_ | _3505_ /*19100*/;
assign _3507_ = ~Q[24] /*19099*/;
assign _3506_ = _3507_ & D[24] /*19098*/;
assign _3509_ = _3129_ & _3506_ /*19093*/;
assign _3510_ = _3129_ ^ _3506_ /*19096*/;
assign _3511_ = _3502_ & _3510_ /*19094*/;
assign _3353_ = _3502_ ^ _3510_ /*19095*/;
assign _3508_ = _3509_ | _3511_ /*19092*/;
assign _3513_ = ~Q[24] /*19091*/;
assign _3512_ = _3513_ & D[25] /*19090*/;
assign _3515_ = _3130_ & _3512_ /*19085*/;
assign _3516_ = _3130_ ^ _3512_ /*19088*/;
assign _3517_ = _3508_ & _3516_ /*19086*/;
assign _3354_ = _3508_ ^ _3516_ /*19087*/;
assign _3514_ = _3515_ | _3517_ /*19084*/;
assign _3519_ = ~Q[24] /*19083*/;
assign _3518_ = _3519_ & D[26] /*19082*/;
assign _3521_ = _3131_ & _3518_ /*19077*/;
assign _3522_ = _3131_ ^ _3518_ /*19080*/;
assign _3523_ = _3514_ & _3522_ /*19078*/;
assign _3355_ = _3514_ ^ _3522_ /*19079*/;
assign _3520_ = _3521_ | _3523_ /*19076*/;
assign _3525_ = ~Q[24] /*19075*/;
assign _3524_ = _3525_ & D[27] /*19074*/;
assign _3527_ = _3132_ & _3524_ /*19069*/;
assign _3528_ = _3132_ ^ _3524_ /*19072*/;
assign _3529_ = _3520_ & _3528_ /*19070*/;
assign _3356_ = _3520_ ^ _3528_ /*19071*/;
assign _3526_ = _3527_ | _3529_ /*19068*/;
assign _3531_ = ~Q[24] /*19067*/;
assign _3530_ = _3531_ & D[28] /*19066*/;
assign _3533_ = _3133_ & _3530_ /*19061*/;
assign _3534_ = _3133_ ^ _3530_ /*19064*/;
assign _3535_ = _3526_ & _3534_ /*19062*/;
assign _3357_ = _3526_ ^ _3534_ /*19063*/;
assign _3532_ = _3533_ | _3535_ /*19060*/;
assign _3537_ = ~Q[24] /*19059*/;
assign _3536_ = _3537_ & D[29] /*19058*/;
assign _3539_ = _3134_ & _3536_ /*19053*/;
assign _3540_ = _3134_ ^ _3536_ /*19056*/;
assign _3541_ = _3532_ & _3540_ /*19054*/;
assign _3358_ = _3532_ ^ _3540_ /*19055*/;
assign _3538_ = _3539_ | _3541_ /*19052*/;
assign _3543_ = ~Q[24] /*19051*/;
assign _3542_ = _3543_ & D[30] /*19050*/;
assign _3545_ = _3135_ & _3542_ /*19045*/;
assign _3546_ = _3135_ ^ _3542_ /*19048*/;
assign _3547_ = _3538_ & _3546_ /*19046*/;
assign _3359_ = _3538_ ^ _3546_ /*19047*/;
assign _3544_ = _3545_ | _3547_ /*19044*/;
assign _3549_ = ~Q[24] /*19043*/;
assign _3548_ = _3549_ & zeroWire /*19042*/;
assign _3550_ = _3136_ ^ _3548_ /*19040*/;
assign _3360_ = _3550_ ^ _3544_ /*19039*/;
assign _3589_ = ~D[0] /*18913*/;
assign _3586_ = R_0[23] & _3589_ /*18909*/;
assign _3587_ = R_0[23] ^ _3589_ /*18912*/;
assign _3588_ = oneWire & _3587_ /*18910*/;
assign _3553_ = oneWire ^ _3587_ /*18911*/;
assign _3585_ = _3586_ | _3588_ /*18908*/;
assign _3594_ = ~D[1] /*18907*/;
assign _3591_ = _3329_ & _3594_ /*18903*/;
assign _3592_ = _3329_ ^ _3594_ /*18906*/;
assign _3593_ = _3585_ & _3592_ /*18904*/;
assign _3554_ = _3585_ ^ _3592_ /*18905*/;
assign _3590_ = _3591_ | _3593_ /*18902*/;
assign _3599_ = ~D[2] /*18901*/;
assign _3596_ = _3330_ & _3599_ /*18897*/;
assign _3597_ = _3330_ ^ _3599_ /*18900*/;
assign _3598_ = _3590_ & _3597_ /*18898*/;
assign _3555_ = _3590_ ^ _3597_ /*18899*/;
assign _3595_ = _3596_ | _3598_ /*18896*/;
assign _3604_ = ~D[3] /*18895*/;
assign _3601_ = _3331_ & _3604_ /*18891*/;
assign _3602_ = _3331_ ^ _3604_ /*18894*/;
assign _3603_ = _3595_ & _3602_ /*18892*/;
assign _3556_ = _3595_ ^ _3602_ /*18893*/;
assign _3600_ = _3601_ | _3603_ /*18890*/;
assign _3609_ = ~D[4] /*18889*/;
assign _3606_ = _3332_ & _3609_ /*18885*/;
assign _3607_ = _3332_ ^ _3609_ /*18888*/;
assign _3608_ = _3600_ & _3607_ /*18886*/;
assign _3557_ = _3600_ ^ _3607_ /*18887*/;
assign _3605_ = _3606_ | _3608_ /*18884*/;
assign _3614_ = ~D[5] /*18883*/;
assign _3611_ = _3333_ & _3614_ /*18879*/;
assign _3612_ = _3333_ ^ _3614_ /*18882*/;
assign _3613_ = _3605_ & _3612_ /*18880*/;
assign _3558_ = _3605_ ^ _3612_ /*18881*/;
assign _3610_ = _3611_ | _3613_ /*18878*/;
assign _3619_ = ~D[6] /*18877*/;
assign _3616_ = _3334_ & _3619_ /*18873*/;
assign _3617_ = _3334_ ^ _3619_ /*18876*/;
assign _3618_ = _3610_ & _3617_ /*18874*/;
assign _3559_ = _3610_ ^ _3617_ /*18875*/;
assign _3615_ = _3616_ | _3618_ /*18872*/;
assign _3624_ = ~D[7] /*18871*/;
assign _3621_ = _3335_ & _3624_ /*18867*/;
assign _3622_ = _3335_ ^ _3624_ /*18870*/;
assign _3623_ = _3615_ & _3622_ /*18868*/;
assign _3560_ = _3615_ ^ _3622_ /*18869*/;
assign _3620_ = _3621_ | _3623_ /*18866*/;
assign _3629_ = ~D[8] /*18865*/;
assign _3626_ = _3336_ & _3629_ /*18861*/;
assign _3627_ = _3336_ ^ _3629_ /*18864*/;
assign _3628_ = _3620_ & _3627_ /*18862*/;
assign _3561_ = _3620_ ^ _3627_ /*18863*/;
assign _3625_ = _3626_ | _3628_ /*18860*/;
assign _3634_ = ~D[9] /*18859*/;
assign _3631_ = _3337_ & _3634_ /*18855*/;
assign _3632_ = _3337_ ^ _3634_ /*18858*/;
assign _3633_ = _3625_ & _3632_ /*18856*/;
assign _3562_ = _3625_ ^ _3632_ /*18857*/;
assign _3630_ = _3631_ | _3633_ /*18854*/;
assign _3639_ = ~D[10] /*18853*/;
assign _3636_ = _3338_ & _3639_ /*18849*/;
assign _3637_ = _3338_ ^ _3639_ /*18852*/;
assign _3638_ = _3630_ & _3637_ /*18850*/;
assign _3563_ = _3630_ ^ _3637_ /*18851*/;
assign _3635_ = _3636_ | _3638_ /*18848*/;
assign _3644_ = ~D[11] /*18847*/;
assign _3641_ = _3339_ & _3644_ /*18843*/;
assign _3642_ = _3339_ ^ _3644_ /*18846*/;
assign _3643_ = _3635_ & _3642_ /*18844*/;
assign _3564_ = _3635_ ^ _3642_ /*18845*/;
assign _3640_ = _3641_ | _3643_ /*18842*/;
assign _3649_ = ~D[12] /*18841*/;
assign _3646_ = _3340_ & _3649_ /*18837*/;
assign _3647_ = _3340_ ^ _3649_ /*18840*/;
assign _3648_ = _3640_ & _3647_ /*18838*/;
assign _3565_ = _3640_ ^ _3647_ /*18839*/;
assign _3645_ = _3646_ | _3648_ /*18836*/;
assign _3654_ = ~D[13] /*18835*/;
assign _3651_ = _3341_ & _3654_ /*18831*/;
assign _3652_ = _3341_ ^ _3654_ /*18834*/;
assign _3653_ = _3645_ & _3652_ /*18832*/;
assign _3566_ = _3645_ ^ _3652_ /*18833*/;
assign _3650_ = _3651_ | _3653_ /*18830*/;
assign _3659_ = ~D[14] /*18829*/;
assign _3656_ = _3342_ & _3659_ /*18825*/;
assign _3657_ = _3342_ ^ _3659_ /*18828*/;
assign _3658_ = _3650_ & _3657_ /*18826*/;
assign _3567_ = _3650_ ^ _3657_ /*18827*/;
assign _3655_ = _3656_ | _3658_ /*18824*/;
assign _3664_ = ~D[15] /*18823*/;
assign _3661_ = _3343_ & _3664_ /*18819*/;
assign _3662_ = _3343_ ^ _3664_ /*18822*/;
assign _3663_ = _3655_ & _3662_ /*18820*/;
assign _3568_ = _3655_ ^ _3662_ /*18821*/;
assign _3660_ = _3661_ | _3663_ /*18818*/;
assign _3669_ = ~D[16] /*18817*/;
assign _3666_ = _3344_ & _3669_ /*18813*/;
assign _3667_ = _3344_ ^ _3669_ /*18816*/;
assign _3668_ = _3660_ & _3667_ /*18814*/;
assign _3569_ = _3660_ ^ _3667_ /*18815*/;
assign _3665_ = _3666_ | _3668_ /*18812*/;
assign _3674_ = ~D[17] /*18811*/;
assign _3671_ = _3345_ & _3674_ /*18807*/;
assign _3672_ = _3345_ ^ _3674_ /*18810*/;
assign _3673_ = _3665_ & _3672_ /*18808*/;
assign _3570_ = _3665_ ^ _3672_ /*18809*/;
assign _3670_ = _3671_ | _3673_ /*18806*/;
assign _3679_ = ~D[18] /*18805*/;
assign _3676_ = _3346_ & _3679_ /*18801*/;
assign _3677_ = _3346_ ^ _3679_ /*18804*/;
assign _3678_ = _3670_ & _3677_ /*18802*/;
assign _3571_ = _3670_ ^ _3677_ /*18803*/;
assign _3675_ = _3676_ | _3678_ /*18800*/;
assign _3684_ = ~D[19] /*18799*/;
assign _3681_ = _3347_ & _3684_ /*18795*/;
assign _3682_ = _3347_ ^ _3684_ /*18798*/;
assign _3683_ = _3675_ & _3682_ /*18796*/;
assign _3572_ = _3675_ ^ _3682_ /*18797*/;
assign _3680_ = _3681_ | _3683_ /*18794*/;
assign _3689_ = ~D[20] /*18793*/;
assign _3686_ = _3348_ & _3689_ /*18789*/;
assign _3687_ = _3348_ ^ _3689_ /*18792*/;
assign _3688_ = _3680_ & _3687_ /*18790*/;
assign _3573_ = _3680_ ^ _3687_ /*18791*/;
assign _3685_ = _3686_ | _3688_ /*18788*/;
assign _3694_ = ~D[21] /*18787*/;
assign _3691_ = _3349_ & _3694_ /*18783*/;
assign _3692_ = _3349_ ^ _3694_ /*18786*/;
assign _3693_ = _3685_ & _3692_ /*18784*/;
assign _3574_ = _3685_ ^ _3692_ /*18785*/;
assign _3690_ = _3691_ | _3693_ /*18782*/;
assign _3699_ = ~D[22] /*18781*/;
assign _3696_ = _3350_ & _3699_ /*18777*/;
assign _3697_ = _3350_ ^ _3699_ /*18780*/;
assign _3698_ = _3690_ & _3697_ /*18778*/;
assign _3575_ = _3690_ ^ _3697_ /*18779*/;
assign _3695_ = _3696_ | _3698_ /*18776*/;
assign _3704_ = ~D[23] /*18775*/;
assign _3701_ = _3351_ & _3704_ /*18771*/;
assign _3702_ = _3351_ ^ _3704_ /*18774*/;
assign _3703_ = _3695_ & _3702_ /*18772*/;
assign _3576_ = _3695_ ^ _3702_ /*18773*/;
assign _3700_ = _3701_ | _3703_ /*18770*/;
assign _3709_ = ~D[24] /*18769*/;
assign _3706_ = _3352_ & _3709_ /*18765*/;
assign _3707_ = _3352_ ^ _3709_ /*18768*/;
assign _3708_ = _3700_ & _3707_ /*18766*/;
assign _3577_ = _3700_ ^ _3707_ /*18767*/;
assign _3705_ = _3706_ | _3708_ /*18764*/;
assign _3714_ = ~D[25] /*18763*/;
assign _3711_ = _3353_ & _3714_ /*18759*/;
assign _3712_ = _3353_ ^ _3714_ /*18762*/;
assign _3713_ = _3705_ & _3712_ /*18760*/;
assign _3578_ = _3705_ ^ _3712_ /*18761*/;
assign _3710_ = _3711_ | _3713_ /*18758*/;
assign _3719_ = ~D[26] /*18757*/;
assign _3716_ = _3354_ & _3719_ /*18753*/;
assign _3717_ = _3354_ ^ _3719_ /*18756*/;
assign _3718_ = _3710_ & _3717_ /*18754*/;
assign _3579_ = _3710_ ^ _3717_ /*18755*/;
assign _3715_ = _3716_ | _3718_ /*18752*/;
assign _3724_ = ~D[27] /*18751*/;
assign _3721_ = _3355_ & _3724_ /*18747*/;
assign _3722_ = _3355_ ^ _3724_ /*18750*/;
assign _3723_ = _3715_ & _3722_ /*18748*/;
assign _3580_ = _3715_ ^ _3722_ /*18749*/;
assign _3720_ = _3721_ | _3723_ /*18746*/;
assign _3729_ = ~D[28] /*18745*/;
assign _3726_ = _3356_ & _3729_ /*18741*/;
assign _3727_ = _3356_ ^ _3729_ /*18744*/;
assign _3728_ = _3720_ & _3727_ /*18742*/;
assign _3581_ = _3720_ ^ _3727_ /*18743*/;
assign _3725_ = _3726_ | _3728_ /*18740*/;
assign _3734_ = ~D[29] /*18739*/;
assign _3731_ = _3357_ & _3734_ /*18735*/;
assign _3732_ = _3357_ ^ _3734_ /*18738*/;
assign _3733_ = _3725_ & _3732_ /*18736*/;
assign _3582_ = _3725_ ^ _3732_ /*18737*/;
assign _3730_ = _3731_ | _3733_ /*18734*/;
assign _3739_ = ~D[30] /*18733*/;
assign _3736_ = _3358_ & _3739_ /*18729*/;
assign _3737_ = _3358_ ^ _3739_ /*18732*/;
assign _3738_ = _3730_ & _3737_ /*18730*/;
assign _3583_ = _3730_ ^ _3737_ /*18731*/;
assign _3735_ = _3736_ | _3738_ /*18728*/;
assign _3740_ = _3359_ & oneWire /*18723*/;
assign _3741_ = _3359_ ^ oneWire /*18726*/;
assign _3742_ = _3735_ & _3741_ /*18724*/;
assign _3584_ = _3735_ ^ _3741_ /*18725*/;
assign Q[23] = _3740_ | _3742_ /*18722*/;
assign _3811_ = ~Q[23] /*18529*/;
assign _3810_ = _3811_ & D[0] /*18528*/;
assign _3813_ = _3553_ & _3810_ /*18523*/;
assign _3814_ = _3553_ ^ _3810_ /*18526*/;
assign _3815_ = zeroWire & _3814_ /*18524*/;
assign _3777_ = zeroWire ^ _3814_ /*18525*/;
assign _3812_ = _3813_ | _3815_ /*18522*/;
assign _3817_ = ~Q[23] /*18521*/;
assign _3816_ = _3817_ & D[1] /*18520*/;
assign _3819_ = _3554_ & _3816_ /*18515*/;
assign _3820_ = _3554_ ^ _3816_ /*18518*/;
assign _3821_ = _3812_ & _3820_ /*18516*/;
assign _3778_ = _3812_ ^ _3820_ /*18517*/;
assign _3818_ = _3819_ | _3821_ /*18514*/;
assign _3823_ = ~Q[23] /*18513*/;
assign _3822_ = _3823_ & D[2] /*18512*/;
assign _3825_ = _3555_ & _3822_ /*18507*/;
assign _3826_ = _3555_ ^ _3822_ /*18510*/;
assign _3827_ = _3818_ & _3826_ /*18508*/;
assign _3779_ = _3818_ ^ _3826_ /*18509*/;
assign _3824_ = _3825_ | _3827_ /*18506*/;
assign _3829_ = ~Q[23] /*18505*/;
assign _3828_ = _3829_ & D[3] /*18504*/;
assign _3831_ = _3556_ & _3828_ /*18499*/;
assign _3832_ = _3556_ ^ _3828_ /*18502*/;
assign _3833_ = _3824_ & _3832_ /*18500*/;
assign _3780_ = _3824_ ^ _3832_ /*18501*/;
assign _3830_ = _3831_ | _3833_ /*18498*/;
assign _3835_ = ~Q[23] /*18497*/;
assign _3834_ = _3835_ & D[4] /*18496*/;
assign _3837_ = _3557_ & _3834_ /*18491*/;
assign _3838_ = _3557_ ^ _3834_ /*18494*/;
assign _3839_ = _3830_ & _3838_ /*18492*/;
assign _3781_ = _3830_ ^ _3838_ /*18493*/;
assign _3836_ = _3837_ | _3839_ /*18490*/;
assign _3841_ = ~Q[23] /*18489*/;
assign _3840_ = _3841_ & D[5] /*18488*/;
assign _3843_ = _3558_ & _3840_ /*18483*/;
assign _3844_ = _3558_ ^ _3840_ /*18486*/;
assign _3845_ = _3836_ & _3844_ /*18484*/;
assign _3782_ = _3836_ ^ _3844_ /*18485*/;
assign _3842_ = _3843_ | _3845_ /*18482*/;
assign _3847_ = ~Q[23] /*18481*/;
assign _3846_ = _3847_ & D[6] /*18480*/;
assign _3849_ = _3559_ & _3846_ /*18475*/;
assign _3850_ = _3559_ ^ _3846_ /*18478*/;
assign _3851_ = _3842_ & _3850_ /*18476*/;
assign _3783_ = _3842_ ^ _3850_ /*18477*/;
assign _3848_ = _3849_ | _3851_ /*18474*/;
assign _3853_ = ~Q[23] /*18473*/;
assign _3852_ = _3853_ & D[7] /*18472*/;
assign _3855_ = _3560_ & _3852_ /*18467*/;
assign _3856_ = _3560_ ^ _3852_ /*18470*/;
assign _3857_ = _3848_ & _3856_ /*18468*/;
assign _3784_ = _3848_ ^ _3856_ /*18469*/;
assign _3854_ = _3855_ | _3857_ /*18466*/;
assign _3859_ = ~Q[23] /*18465*/;
assign _3858_ = _3859_ & D[8] /*18464*/;
assign _3861_ = _3561_ & _3858_ /*18459*/;
assign _3862_ = _3561_ ^ _3858_ /*18462*/;
assign _3863_ = _3854_ & _3862_ /*18460*/;
assign _3785_ = _3854_ ^ _3862_ /*18461*/;
assign _3860_ = _3861_ | _3863_ /*18458*/;
assign _3865_ = ~Q[23] /*18457*/;
assign _3864_ = _3865_ & D[9] /*18456*/;
assign _3867_ = _3562_ & _3864_ /*18451*/;
assign _3868_ = _3562_ ^ _3864_ /*18454*/;
assign _3869_ = _3860_ & _3868_ /*18452*/;
assign _3786_ = _3860_ ^ _3868_ /*18453*/;
assign _3866_ = _3867_ | _3869_ /*18450*/;
assign _3871_ = ~Q[23] /*18449*/;
assign _3870_ = _3871_ & D[10] /*18448*/;
assign _3873_ = _3563_ & _3870_ /*18443*/;
assign _3874_ = _3563_ ^ _3870_ /*18446*/;
assign _3875_ = _3866_ & _3874_ /*18444*/;
assign _3787_ = _3866_ ^ _3874_ /*18445*/;
assign _3872_ = _3873_ | _3875_ /*18442*/;
assign _3877_ = ~Q[23] /*18441*/;
assign _3876_ = _3877_ & D[11] /*18440*/;
assign _3879_ = _3564_ & _3876_ /*18435*/;
assign _3880_ = _3564_ ^ _3876_ /*18438*/;
assign _3881_ = _3872_ & _3880_ /*18436*/;
assign _3788_ = _3872_ ^ _3880_ /*18437*/;
assign _3878_ = _3879_ | _3881_ /*18434*/;
assign _3883_ = ~Q[23] /*18433*/;
assign _3882_ = _3883_ & D[12] /*18432*/;
assign _3885_ = _3565_ & _3882_ /*18427*/;
assign _3886_ = _3565_ ^ _3882_ /*18430*/;
assign _3887_ = _3878_ & _3886_ /*18428*/;
assign _3789_ = _3878_ ^ _3886_ /*18429*/;
assign _3884_ = _3885_ | _3887_ /*18426*/;
assign _3889_ = ~Q[23] /*18425*/;
assign _3888_ = _3889_ & D[13] /*18424*/;
assign _3891_ = _3566_ & _3888_ /*18419*/;
assign _3892_ = _3566_ ^ _3888_ /*18422*/;
assign _3893_ = _3884_ & _3892_ /*18420*/;
assign _3790_ = _3884_ ^ _3892_ /*18421*/;
assign _3890_ = _3891_ | _3893_ /*18418*/;
assign _3895_ = ~Q[23] /*18417*/;
assign _3894_ = _3895_ & D[14] /*18416*/;
assign _3897_ = _3567_ & _3894_ /*18411*/;
assign _3898_ = _3567_ ^ _3894_ /*18414*/;
assign _3899_ = _3890_ & _3898_ /*18412*/;
assign _3791_ = _3890_ ^ _3898_ /*18413*/;
assign _3896_ = _3897_ | _3899_ /*18410*/;
assign _3901_ = ~Q[23] /*18409*/;
assign _3900_ = _3901_ & D[15] /*18408*/;
assign _3903_ = _3568_ & _3900_ /*18403*/;
assign _3904_ = _3568_ ^ _3900_ /*18406*/;
assign _3905_ = _3896_ & _3904_ /*18404*/;
assign _3792_ = _3896_ ^ _3904_ /*18405*/;
assign _3902_ = _3903_ | _3905_ /*18402*/;
assign _3907_ = ~Q[23] /*18401*/;
assign _3906_ = _3907_ & D[16] /*18400*/;
assign _3909_ = _3569_ & _3906_ /*18395*/;
assign _3910_ = _3569_ ^ _3906_ /*18398*/;
assign _3911_ = _3902_ & _3910_ /*18396*/;
assign _3793_ = _3902_ ^ _3910_ /*18397*/;
assign _3908_ = _3909_ | _3911_ /*18394*/;
assign _3913_ = ~Q[23] /*18393*/;
assign _3912_ = _3913_ & D[17] /*18392*/;
assign _3915_ = _3570_ & _3912_ /*18387*/;
assign _3916_ = _3570_ ^ _3912_ /*18390*/;
assign _3917_ = _3908_ & _3916_ /*18388*/;
assign _3794_ = _3908_ ^ _3916_ /*18389*/;
assign _3914_ = _3915_ | _3917_ /*18386*/;
assign _3919_ = ~Q[23] /*18385*/;
assign _3918_ = _3919_ & D[18] /*18384*/;
assign _3921_ = _3571_ & _3918_ /*18379*/;
assign _3922_ = _3571_ ^ _3918_ /*18382*/;
assign _3923_ = _3914_ & _3922_ /*18380*/;
assign _3795_ = _3914_ ^ _3922_ /*18381*/;
assign _3920_ = _3921_ | _3923_ /*18378*/;
assign _3925_ = ~Q[23] /*18377*/;
assign _3924_ = _3925_ & D[19] /*18376*/;
assign _3927_ = _3572_ & _3924_ /*18371*/;
assign _3928_ = _3572_ ^ _3924_ /*18374*/;
assign _3929_ = _3920_ & _3928_ /*18372*/;
assign _3796_ = _3920_ ^ _3928_ /*18373*/;
assign _3926_ = _3927_ | _3929_ /*18370*/;
assign _3931_ = ~Q[23] /*18369*/;
assign _3930_ = _3931_ & D[20] /*18368*/;
assign _3933_ = _3573_ & _3930_ /*18363*/;
assign _3934_ = _3573_ ^ _3930_ /*18366*/;
assign _3935_ = _3926_ & _3934_ /*18364*/;
assign _3797_ = _3926_ ^ _3934_ /*18365*/;
assign _3932_ = _3933_ | _3935_ /*18362*/;
assign _3937_ = ~Q[23] /*18361*/;
assign _3936_ = _3937_ & D[21] /*18360*/;
assign _3939_ = _3574_ & _3936_ /*18355*/;
assign _3940_ = _3574_ ^ _3936_ /*18358*/;
assign _3941_ = _3932_ & _3940_ /*18356*/;
assign _3798_ = _3932_ ^ _3940_ /*18357*/;
assign _3938_ = _3939_ | _3941_ /*18354*/;
assign _3943_ = ~Q[23] /*18353*/;
assign _3942_ = _3943_ & D[22] /*18352*/;
assign _3945_ = _3575_ & _3942_ /*18347*/;
assign _3946_ = _3575_ ^ _3942_ /*18350*/;
assign _3947_ = _3938_ & _3946_ /*18348*/;
assign _3799_ = _3938_ ^ _3946_ /*18349*/;
assign _3944_ = _3945_ | _3947_ /*18346*/;
assign _3949_ = ~Q[23] /*18345*/;
assign _3948_ = _3949_ & D[23] /*18344*/;
assign _3951_ = _3576_ & _3948_ /*18339*/;
assign _3952_ = _3576_ ^ _3948_ /*18342*/;
assign _3953_ = _3944_ & _3952_ /*18340*/;
assign _3800_ = _3944_ ^ _3952_ /*18341*/;
assign _3950_ = _3951_ | _3953_ /*18338*/;
assign _3955_ = ~Q[23] /*18337*/;
assign _3954_ = _3955_ & D[24] /*18336*/;
assign _3957_ = _3577_ & _3954_ /*18331*/;
assign _3958_ = _3577_ ^ _3954_ /*18334*/;
assign _3959_ = _3950_ & _3958_ /*18332*/;
assign _3801_ = _3950_ ^ _3958_ /*18333*/;
assign _3956_ = _3957_ | _3959_ /*18330*/;
assign _3961_ = ~Q[23] /*18329*/;
assign _3960_ = _3961_ & D[25] /*18328*/;
assign _3963_ = _3578_ & _3960_ /*18323*/;
assign _3964_ = _3578_ ^ _3960_ /*18326*/;
assign _3965_ = _3956_ & _3964_ /*18324*/;
assign _3802_ = _3956_ ^ _3964_ /*18325*/;
assign _3962_ = _3963_ | _3965_ /*18322*/;
assign _3967_ = ~Q[23] /*18321*/;
assign _3966_ = _3967_ & D[26] /*18320*/;
assign _3969_ = _3579_ & _3966_ /*18315*/;
assign _3970_ = _3579_ ^ _3966_ /*18318*/;
assign _3971_ = _3962_ & _3970_ /*18316*/;
assign _3803_ = _3962_ ^ _3970_ /*18317*/;
assign _3968_ = _3969_ | _3971_ /*18314*/;
assign _3973_ = ~Q[23] /*18313*/;
assign _3972_ = _3973_ & D[27] /*18312*/;
assign _3975_ = _3580_ & _3972_ /*18307*/;
assign _3976_ = _3580_ ^ _3972_ /*18310*/;
assign _3977_ = _3968_ & _3976_ /*18308*/;
assign _3804_ = _3968_ ^ _3976_ /*18309*/;
assign _3974_ = _3975_ | _3977_ /*18306*/;
assign _3979_ = ~Q[23] /*18305*/;
assign _3978_ = _3979_ & D[28] /*18304*/;
assign _3981_ = _3581_ & _3978_ /*18299*/;
assign _3982_ = _3581_ ^ _3978_ /*18302*/;
assign _3983_ = _3974_ & _3982_ /*18300*/;
assign _3805_ = _3974_ ^ _3982_ /*18301*/;
assign _3980_ = _3981_ | _3983_ /*18298*/;
assign _3985_ = ~Q[23] /*18297*/;
assign _3984_ = _3985_ & D[29] /*18296*/;
assign _3987_ = _3582_ & _3984_ /*18291*/;
assign _3988_ = _3582_ ^ _3984_ /*18294*/;
assign _3989_ = _3980_ & _3988_ /*18292*/;
assign _3806_ = _3980_ ^ _3988_ /*18293*/;
assign _3986_ = _3987_ | _3989_ /*18290*/;
assign _3991_ = ~Q[23] /*18289*/;
assign _3990_ = _3991_ & D[30] /*18288*/;
assign _3993_ = _3583_ & _3990_ /*18283*/;
assign _3994_ = _3583_ ^ _3990_ /*18286*/;
assign _3995_ = _3986_ & _3994_ /*18284*/;
assign _3807_ = _3986_ ^ _3994_ /*18285*/;
assign _3992_ = _3993_ | _3995_ /*18282*/;
assign _3997_ = ~Q[23] /*18281*/;
assign _3996_ = _3997_ & zeroWire /*18280*/;
assign _3998_ = _3584_ ^ _3996_ /*18278*/;
assign _3808_ = _3998_ ^ _3992_ /*18277*/;
assign _4037_ = ~D[0] /*18151*/;
assign _4034_ = R_0[22] & _4037_ /*18147*/;
assign _4035_ = R_0[22] ^ _4037_ /*18150*/;
assign _4036_ = oneWire & _4035_ /*18148*/;
assign _4001_ = oneWire ^ _4035_ /*18149*/;
assign _4033_ = _4034_ | _4036_ /*18146*/;
assign _4042_ = ~D[1] /*18145*/;
assign _4039_ = _3777_ & _4042_ /*18141*/;
assign _4040_ = _3777_ ^ _4042_ /*18144*/;
assign _4041_ = _4033_ & _4040_ /*18142*/;
assign _4002_ = _4033_ ^ _4040_ /*18143*/;
assign _4038_ = _4039_ | _4041_ /*18140*/;
assign _4047_ = ~D[2] /*18139*/;
assign _4044_ = _3778_ & _4047_ /*18135*/;
assign _4045_ = _3778_ ^ _4047_ /*18138*/;
assign _4046_ = _4038_ & _4045_ /*18136*/;
assign _4003_ = _4038_ ^ _4045_ /*18137*/;
assign _4043_ = _4044_ | _4046_ /*18134*/;
assign _4052_ = ~D[3] /*18133*/;
assign _4049_ = _3779_ & _4052_ /*18129*/;
assign _4050_ = _3779_ ^ _4052_ /*18132*/;
assign _4051_ = _4043_ & _4050_ /*18130*/;
assign _4004_ = _4043_ ^ _4050_ /*18131*/;
assign _4048_ = _4049_ | _4051_ /*18128*/;
assign _4057_ = ~D[4] /*18127*/;
assign _4054_ = _3780_ & _4057_ /*18123*/;
assign _4055_ = _3780_ ^ _4057_ /*18126*/;
assign _4056_ = _4048_ & _4055_ /*18124*/;
assign _4005_ = _4048_ ^ _4055_ /*18125*/;
assign _4053_ = _4054_ | _4056_ /*18122*/;
assign _4062_ = ~D[5] /*18121*/;
assign _4059_ = _3781_ & _4062_ /*18117*/;
assign _4060_ = _3781_ ^ _4062_ /*18120*/;
assign _4061_ = _4053_ & _4060_ /*18118*/;
assign _4006_ = _4053_ ^ _4060_ /*18119*/;
assign _4058_ = _4059_ | _4061_ /*18116*/;
assign _4067_ = ~D[6] /*18115*/;
assign _4064_ = _3782_ & _4067_ /*18111*/;
assign _4065_ = _3782_ ^ _4067_ /*18114*/;
assign _4066_ = _4058_ & _4065_ /*18112*/;
assign _4007_ = _4058_ ^ _4065_ /*18113*/;
assign _4063_ = _4064_ | _4066_ /*18110*/;
assign _4072_ = ~D[7] /*18109*/;
assign _4069_ = _3783_ & _4072_ /*18105*/;
assign _4070_ = _3783_ ^ _4072_ /*18108*/;
assign _4071_ = _4063_ & _4070_ /*18106*/;
assign _4008_ = _4063_ ^ _4070_ /*18107*/;
assign _4068_ = _4069_ | _4071_ /*18104*/;
assign _4077_ = ~D[8] /*18103*/;
assign _4074_ = _3784_ & _4077_ /*18099*/;
assign _4075_ = _3784_ ^ _4077_ /*18102*/;
assign _4076_ = _4068_ & _4075_ /*18100*/;
assign _4009_ = _4068_ ^ _4075_ /*18101*/;
assign _4073_ = _4074_ | _4076_ /*18098*/;
assign _4082_ = ~D[9] /*18097*/;
assign _4079_ = _3785_ & _4082_ /*18093*/;
assign _4080_ = _3785_ ^ _4082_ /*18096*/;
assign _4081_ = _4073_ & _4080_ /*18094*/;
assign _4010_ = _4073_ ^ _4080_ /*18095*/;
assign _4078_ = _4079_ | _4081_ /*18092*/;
assign _4087_ = ~D[10] /*18091*/;
assign _4084_ = _3786_ & _4087_ /*18087*/;
assign _4085_ = _3786_ ^ _4087_ /*18090*/;
assign _4086_ = _4078_ & _4085_ /*18088*/;
assign _4011_ = _4078_ ^ _4085_ /*18089*/;
assign _4083_ = _4084_ | _4086_ /*18086*/;
assign _4092_ = ~D[11] /*18085*/;
assign _4089_ = _3787_ & _4092_ /*18081*/;
assign _4090_ = _3787_ ^ _4092_ /*18084*/;
assign _4091_ = _4083_ & _4090_ /*18082*/;
assign _4012_ = _4083_ ^ _4090_ /*18083*/;
assign _4088_ = _4089_ | _4091_ /*18080*/;
assign _4097_ = ~D[12] /*18079*/;
assign _4094_ = _3788_ & _4097_ /*18075*/;
assign _4095_ = _3788_ ^ _4097_ /*18078*/;
assign _4096_ = _4088_ & _4095_ /*18076*/;
assign _4013_ = _4088_ ^ _4095_ /*18077*/;
assign _4093_ = _4094_ | _4096_ /*18074*/;
assign _4102_ = ~D[13] /*18073*/;
assign _4099_ = _3789_ & _4102_ /*18069*/;
assign _4100_ = _3789_ ^ _4102_ /*18072*/;
assign _4101_ = _4093_ & _4100_ /*18070*/;
assign _4014_ = _4093_ ^ _4100_ /*18071*/;
assign _4098_ = _4099_ | _4101_ /*18068*/;
assign _4107_ = ~D[14] /*18067*/;
assign _4104_ = _3790_ & _4107_ /*18063*/;
assign _4105_ = _3790_ ^ _4107_ /*18066*/;
assign _4106_ = _4098_ & _4105_ /*18064*/;
assign _4015_ = _4098_ ^ _4105_ /*18065*/;
assign _4103_ = _4104_ | _4106_ /*18062*/;
assign _4112_ = ~D[15] /*18061*/;
assign _4109_ = _3791_ & _4112_ /*18057*/;
assign _4110_ = _3791_ ^ _4112_ /*18060*/;
assign _4111_ = _4103_ & _4110_ /*18058*/;
assign _4016_ = _4103_ ^ _4110_ /*18059*/;
assign _4108_ = _4109_ | _4111_ /*18056*/;
assign _4117_ = ~D[16] /*18055*/;
assign _4114_ = _3792_ & _4117_ /*18051*/;
assign _4115_ = _3792_ ^ _4117_ /*18054*/;
assign _4116_ = _4108_ & _4115_ /*18052*/;
assign _4017_ = _4108_ ^ _4115_ /*18053*/;
assign _4113_ = _4114_ | _4116_ /*18050*/;
assign _4122_ = ~D[17] /*18049*/;
assign _4119_ = _3793_ & _4122_ /*18045*/;
assign _4120_ = _3793_ ^ _4122_ /*18048*/;
assign _4121_ = _4113_ & _4120_ /*18046*/;
assign _4018_ = _4113_ ^ _4120_ /*18047*/;
assign _4118_ = _4119_ | _4121_ /*18044*/;
assign _4127_ = ~D[18] /*18043*/;
assign _4124_ = _3794_ & _4127_ /*18039*/;
assign _4125_ = _3794_ ^ _4127_ /*18042*/;
assign _4126_ = _4118_ & _4125_ /*18040*/;
assign _4019_ = _4118_ ^ _4125_ /*18041*/;
assign _4123_ = _4124_ | _4126_ /*18038*/;
assign _4132_ = ~D[19] /*18037*/;
assign _4129_ = _3795_ & _4132_ /*18033*/;
assign _4130_ = _3795_ ^ _4132_ /*18036*/;
assign _4131_ = _4123_ & _4130_ /*18034*/;
assign _4020_ = _4123_ ^ _4130_ /*18035*/;
assign _4128_ = _4129_ | _4131_ /*18032*/;
assign _4137_ = ~D[20] /*18031*/;
assign _4134_ = _3796_ & _4137_ /*18027*/;
assign _4135_ = _3796_ ^ _4137_ /*18030*/;
assign _4136_ = _4128_ & _4135_ /*18028*/;
assign _4021_ = _4128_ ^ _4135_ /*18029*/;
assign _4133_ = _4134_ | _4136_ /*18026*/;
assign _4142_ = ~D[21] /*18025*/;
assign _4139_ = _3797_ & _4142_ /*18021*/;
assign _4140_ = _3797_ ^ _4142_ /*18024*/;
assign _4141_ = _4133_ & _4140_ /*18022*/;
assign _4022_ = _4133_ ^ _4140_ /*18023*/;
assign _4138_ = _4139_ | _4141_ /*18020*/;
assign _4147_ = ~D[22] /*18019*/;
assign _4144_ = _3798_ & _4147_ /*18015*/;
assign _4145_ = _3798_ ^ _4147_ /*18018*/;
assign _4146_ = _4138_ & _4145_ /*18016*/;
assign _4023_ = _4138_ ^ _4145_ /*18017*/;
assign _4143_ = _4144_ | _4146_ /*18014*/;
assign _4152_ = ~D[23] /*18013*/;
assign _4149_ = _3799_ & _4152_ /*18009*/;
assign _4150_ = _3799_ ^ _4152_ /*18012*/;
assign _4151_ = _4143_ & _4150_ /*18010*/;
assign _4024_ = _4143_ ^ _4150_ /*18011*/;
assign _4148_ = _4149_ | _4151_ /*18008*/;
assign _4157_ = ~D[24] /*18007*/;
assign _4154_ = _3800_ & _4157_ /*18003*/;
assign _4155_ = _3800_ ^ _4157_ /*18006*/;
assign _4156_ = _4148_ & _4155_ /*18004*/;
assign _4025_ = _4148_ ^ _4155_ /*18005*/;
assign _4153_ = _4154_ | _4156_ /*18002*/;
assign _4162_ = ~D[25] /*18001*/;
assign _4159_ = _3801_ & _4162_ /*17997*/;
assign _4160_ = _3801_ ^ _4162_ /*18000*/;
assign _4161_ = _4153_ & _4160_ /*17998*/;
assign _4026_ = _4153_ ^ _4160_ /*17999*/;
assign _4158_ = _4159_ | _4161_ /*17996*/;
assign _4167_ = ~D[26] /*17995*/;
assign _4164_ = _3802_ & _4167_ /*17991*/;
assign _4165_ = _3802_ ^ _4167_ /*17994*/;
assign _4166_ = _4158_ & _4165_ /*17992*/;
assign _4027_ = _4158_ ^ _4165_ /*17993*/;
assign _4163_ = _4164_ | _4166_ /*17990*/;
assign _4172_ = ~D[27] /*17989*/;
assign _4169_ = _3803_ & _4172_ /*17985*/;
assign _4170_ = _3803_ ^ _4172_ /*17988*/;
assign _4171_ = _4163_ & _4170_ /*17986*/;
assign _4028_ = _4163_ ^ _4170_ /*17987*/;
assign _4168_ = _4169_ | _4171_ /*17984*/;
assign _4177_ = ~D[28] /*17983*/;
assign _4174_ = _3804_ & _4177_ /*17979*/;
assign _4175_ = _3804_ ^ _4177_ /*17982*/;
assign _4176_ = _4168_ & _4175_ /*17980*/;
assign _4029_ = _4168_ ^ _4175_ /*17981*/;
assign _4173_ = _4174_ | _4176_ /*17978*/;
assign _4182_ = ~D[29] /*17977*/;
assign _4179_ = _3805_ & _4182_ /*17973*/;
assign _4180_ = _3805_ ^ _4182_ /*17976*/;
assign _4181_ = _4173_ & _4180_ /*17974*/;
assign _4030_ = _4173_ ^ _4180_ /*17975*/;
assign _4178_ = _4179_ | _4181_ /*17972*/;
assign _4187_ = ~D[30] /*17971*/;
assign _4184_ = _3806_ & _4187_ /*17967*/;
assign _4185_ = _3806_ ^ _4187_ /*17970*/;
assign _4186_ = _4178_ & _4185_ /*17968*/;
assign _4031_ = _4178_ ^ _4185_ /*17969*/;
assign _4183_ = _4184_ | _4186_ /*17966*/;
assign _4188_ = _3807_ & oneWire /*17961*/;
assign _4189_ = _3807_ ^ oneWire /*17964*/;
assign _4190_ = _4183_ & _4189_ /*17962*/;
assign _4032_ = _4183_ ^ _4189_ /*17963*/;
assign Q[22] = _4188_ | _4190_ /*17960*/;
assign _4259_ = ~Q[22] /*17767*/;
assign _4258_ = _4259_ & D[0] /*17766*/;
assign _4261_ = _4001_ & _4258_ /*17761*/;
assign _4262_ = _4001_ ^ _4258_ /*17764*/;
assign _4263_ = zeroWire & _4262_ /*17762*/;
assign _4225_ = zeroWire ^ _4262_ /*17763*/;
assign _4260_ = _4261_ | _4263_ /*17760*/;
assign _4265_ = ~Q[22] /*17759*/;
assign _4264_ = _4265_ & D[1] /*17758*/;
assign _4267_ = _4002_ & _4264_ /*17753*/;
assign _4268_ = _4002_ ^ _4264_ /*17756*/;
assign _4269_ = _4260_ & _4268_ /*17754*/;
assign _4226_ = _4260_ ^ _4268_ /*17755*/;
assign _4266_ = _4267_ | _4269_ /*17752*/;
assign _4271_ = ~Q[22] /*17751*/;
assign _4270_ = _4271_ & D[2] /*17750*/;
assign _4273_ = _4003_ & _4270_ /*17745*/;
assign _4274_ = _4003_ ^ _4270_ /*17748*/;
assign _4275_ = _4266_ & _4274_ /*17746*/;
assign _4227_ = _4266_ ^ _4274_ /*17747*/;
assign _4272_ = _4273_ | _4275_ /*17744*/;
assign _4277_ = ~Q[22] /*17743*/;
assign _4276_ = _4277_ & D[3] /*17742*/;
assign _4279_ = _4004_ & _4276_ /*17737*/;
assign _4280_ = _4004_ ^ _4276_ /*17740*/;
assign _4281_ = _4272_ & _4280_ /*17738*/;
assign _4228_ = _4272_ ^ _4280_ /*17739*/;
assign _4278_ = _4279_ | _4281_ /*17736*/;
assign _4283_ = ~Q[22] /*17735*/;
assign _4282_ = _4283_ & D[4] /*17734*/;
assign _4285_ = _4005_ & _4282_ /*17729*/;
assign _4286_ = _4005_ ^ _4282_ /*17732*/;
assign _4287_ = _4278_ & _4286_ /*17730*/;
assign _4229_ = _4278_ ^ _4286_ /*17731*/;
assign _4284_ = _4285_ | _4287_ /*17728*/;
assign _4289_ = ~Q[22] /*17727*/;
assign _4288_ = _4289_ & D[5] /*17726*/;
assign _4291_ = _4006_ & _4288_ /*17721*/;
assign _4292_ = _4006_ ^ _4288_ /*17724*/;
assign _4293_ = _4284_ & _4292_ /*17722*/;
assign _4230_ = _4284_ ^ _4292_ /*17723*/;
assign _4290_ = _4291_ | _4293_ /*17720*/;
assign _4295_ = ~Q[22] /*17719*/;
assign _4294_ = _4295_ & D[6] /*17718*/;
assign _4297_ = _4007_ & _4294_ /*17713*/;
assign _4298_ = _4007_ ^ _4294_ /*17716*/;
assign _4299_ = _4290_ & _4298_ /*17714*/;
assign _4231_ = _4290_ ^ _4298_ /*17715*/;
assign _4296_ = _4297_ | _4299_ /*17712*/;
assign _4301_ = ~Q[22] /*17711*/;
assign _4300_ = _4301_ & D[7] /*17710*/;
assign _4303_ = _4008_ & _4300_ /*17705*/;
assign _4304_ = _4008_ ^ _4300_ /*17708*/;
assign _4305_ = _4296_ & _4304_ /*17706*/;
assign _4232_ = _4296_ ^ _4304_ /*17707*/;
assign _4302_ = _4303_ | _4305_ /*17704*/;
assign _4307_ = ~Q[22] /*17703*/;
assign _4306_ = _4307_ & D[8] /*17702*/;
assign _4309_ = _4009_ & _4306_ /*17697*/;
assign _4310_ = _4009_ ^ _4306_ /*17700*/;
assign _4311_ = _4302_ & _4310_ /*17698*/;
assign _4233_ = _4302_ ^ _4310_ /*17699*/;
assign _4308_ = _4309_ | _4311_ /*17696*/;
assign _4313_ = ~Q[22] /*17695*/;
assign _4312_ = _4313_ & D[9] /*17694*/;
assign _4315_ = _4010_ & _4312_ /*17689*/;
assign _4316_ = _4010_ ^ _4312_ /*17692*/;
assign _4317_ = _4308_ & _4316_ /*17690*/;
assign _4234_ = _4308_ ^ _4316_ /*17691*/;
assign _4314_ = _4315_ | _4317_ /*17688*/;
assign _4319_ = ~Q[22] /*17687*/;
assign _4318_ = _4319_ & D[10] /*17686*/;
assign _4321_ = _4011_ & _4318_ /*17681*/;
assign _4322_ = _4011_ ^ _4318_ /*17684*/;
assign _4323_ = _4314_ & _4322_ /*17682*/;
assign _4235_ = _4314_ ^ _4322_ /*17683*/;
assign _4320_ = _4321_ | _4323_ /*17680*/;
assign _4325_ = ~Q[22] /*17679*/;
assign _4324_ = _4325_ & D[11] /*17678*/;
assign _4327_ = _4012_ & _4324_ /*17673*/;
assign _4328_ = _4012_ ^ _4324_ /*17676*/;
assign _4329_ = _4320_ & _4328_ /*17674*/;
assign _4236_ = _4320_ ^ _4328_ /*17675*/;
assign _4326_ = _4327_ | _4329_ /*17672*/;
assign _4331_ = ~Q[22] /*17671*/;
assign _4330_ = _4331_ & D[12] /*17670*/;
assign _4333_ = _4013_ & _4330_ /*17665*/;
assign _4334_ = _4013_ ^ _4330_ /*17668*/;
assign _4335_ = _4326_ & _4334_ /*17666*/;
assign _4237_ = _4326_ ^ _4334_ /*17667*/;
assign _4332_ = _4333_ | _4335_ /*17664*/;
assign _4337_ = ~Q[22] /*17663*/;
assign _4336_ = _4337_ & D[13] /*17662*/;
assign _4339_ = _4014_ & _4336_ /*17657*/;
assign _4340_ = _4014_ ^ _4336_ /*17660*/;
assign _4341_ = _4332_ & _4340_ /*17658*/;
assign _4238_ = _4332_ ^ _4340_ /*17659*/;
assign _4338_ = _4339_ | _4341_ /*17656*/;
assign _4343_ = ~Q[22] /*17655*/;
assign _4342_ = _4343_ & D[14] /*17654*/;
assign _4345_ = _4015_ & _4342_ /*17649*/;
assign _4346_ = _4015_ ^ _4342_ /*17652*/;
assign _4347_ = _4338_ & _4346_ /*17650*/;
assign _4239_ = _4338_ ^ _4346_ /*17651*/;
assign _4344_ = _4345_ | _4347_ /*17648*/;
assign _4349_ = ~Q[22] /*17647*/;
assign _4348_ = _4349_ & D[15] /*17646*/;
assign _4351_ = _4016_ & _4348_ /*17641*/;
assign _4352_ = _4016_ ^ _4348_ /*17644*/;
assign _4353_ = _4344_ & _4352_ /*17642*/;
assign _4240_ = _4344_ ^ _4352_ /*17643*/;
assign _4350_ = _4351_ | _4353_ /*17640*/;
assign _4355_ = ~Q[22] /*17639*/;
assign _4354_ = _4355_ & D[16] /*17638*/;
assign _4357_ = _4017_ & _4354_ /*17633*/;
assign _4358_ = _4017_ ^ _4354_ /*17636*/;
assign _4359_ = _4350_ & _4358_ /*17634*/;
assign _4241_ = _4350_ ^ _4358_ /*17635*/;
assign _4356_ = _4357_ | _4359_ /*17632*/;
assign _4361_ = ~Q[22] /*17631*/;
assign _4360_ = _4361_ & D[17] /*17630*/;
assign _4363_ = _4018_ & _4360_ /*17625*/;
assign _4364_ = _4018_ ^ _4360_ /*17628*/;
assign _4365_ = _4356_ & _4364_ /*17626*/;
assign _4242_ = _4356_ ^ _4364_ /*17627*/;
assign _4362_ = _4363_ | _4365_ /*17624*/;
assign _4367_ = ~Q[22] /*17623*/;
assign _4366_ = _4367_ & D[18] /*17622*/;
assign _4369_ = _4019_ & _4366_ /*17617*/;
assign _4370_ = _4019_ ^ _4366_ /*17620*/;
assign _4371_ = _4362_ & _4370_ /*17618*/;
assign _4243_ = _4362_ ^ _4370_ /*17619*/;
assign _4368_ = _4369_ | _4371_ /*17616*/;
assign _4373_ = ~Q[22] /*17615*/;
assign _4372_ = _4373_ & D[19] /*17614*/;
assign _4375_ = _4020_ & _4372_ /*17609*/;
assign _4376_ = _4020_ ^ _4372_ /*17612*/;
assign _4377_ = _4368_ & _4376_ /*17610*/;
assign _4244_ = _4368_ ^ _4376_ /*17611*/;
assign _4374_ = _4375_ | _4377_ /*17608*/;
assign _4379_ = ~Q[22] /*17607*/;
assign _4378_ = _4379_ & D[20] /*17606*/;
assign _4381_ = _4021_ & _4378_ /*17601*/;
assign _4382_ = _4021_ ^ _4378_ /*17604*/;
assign _4383_ = _4374_ & _4382_ /*17602*/;
assign _4245_ = _4374_ ^ _4382_ /*17603*/;
assign _4380_ = _4381_ | _4383_ /*17600*/;
assign _4385_ = ~Q[22] /*17599*/;
assign _4384_ = _4385_ & D[21] /*17598*/;
assign _4387_ = _4022_ & _4384_ /*17593*/;
assign _4388_ = _4022_ ^ _4384_ /*17596*/;
assign _4389_ = _4380_ & _4388_ /*17594*/;
assign _4246_ = _4380_ ^ _4388_ /*17595*/;
assign _4386_ = _4387_ | _4389_ /*17592*/;
assign _4391_ = ~Q[22] /*17591*/;
assign _4390_ = _4391_ & D[22] /*17590*/;
assign _4393_ = _4023_ & _4390_ /*17585*/;
assign _4394_ = _4023_ ^ _4390_ /*17588*/;
assign _4395_ = _4386_ & _4394_ /*17586*/;
assign _4247_ = _4386_ ^ _4394_ /*17587*/;
assign _4392_ = _4393_ | _4395_ /*17584*/;
assign _4397_ = ~Q[22] /*17583*/;
assign _4396_ = _4397_ & D[23] /*17582*/;
assign _4399_ = _4024_ & _4396_ /*17577*/;
assign _4400_ = _4024_ ^ _4396_ /*17580*/;
assign _4401_ = _4392_ & _4400_ /*17578*/;
assign _4248_ = _4392_ ^ _4400_ /*17579*/;
assign _4398_ = _4399_ | _4401_ /*17576*/;
assign _4403_ = ~Q[22] /*17575*/;
assign _4402_ = _4403_ & D[24] /*17574*/;
assign _4405_ = _4025_ & _4402_ /*17569*/;
assign _4406_ = _4025_ ^ _4402_ /*17572*/;
assign _4407_ = _4398_ & _4406_ /*17570*/;
assign _4249_ = _4398_ ^ _4406_ /*17571*/;
assign _4404_ = _4405_ | _4407_ /*17568*/;
assign _4409_ = ~Q[22] /*17567*/;
assign _4408_ = _4409_ & D[25] /*17566*/;
assign _4411_ = _4026_ & _4408_ /*17561*/;
assign _4412_ = _4026_ ^ _4408_ /*17564*/;
assign _4413_ = _4404_ & _4412_ /*17562*/;
assign _4250_ = _4404_ ^ _4412_ /*17563*/;
assign _4410_ = _4411_ | _4413_ /*17560*/;
assign _4415_ = ~Q[22] /*17559*/;
assign _4414_ = _4415_ & D[26] /*17558*/;
assign _4417_ = _4027_ & _4414_ /*17553*/;
assign _4418_ = _4027_ ^ _4414_ /*17556*/;
assign _4419_ = _4410_ & _4418_ /*17554*/;
assign _4251_ = _4410_ ^ _4418_ /*17555*/;
assign _4416_ = _4417_ | _4419_ /*17552*/;
assign _4421_ = ~Q[22] /*17551*/;
assign _4420_ = _4421_ & D[27] /*17550*/;
assign _4423_ = _4028_ & _4420_ /*17545*/;
assign _4424_ = _4028_ ^ _4420_ /*17548*/;
assign _4425_ = _4416_ & _4424_ /*17546*/;
assign _4252_ = _4416_ ^ _4424_ /*17547*/;
assign _4422_ = _4423_ | _4425_ /*17544*/;
assign _4427_ = ~Q[22] /*17543*/;
assign _4426_ = _4427_ & D[28] /*17542*/;
assign _4429_ = _4029_ & _4426_ /*17537*/;
assign _4430_ = _4029_ ^ _4426_ /*17540*/;
assign _4431_ = _4422_ & _4430_ /*17538*/;
assign _4253_ = _4422_ ^ _4430_ /*17539*/;
assign _4428_ = _4429_ | _4431_ /*17536*/;
assign _4433_ = ~Q[22] /*17535*/;
assign _4432_ = _4433_ & D[29] /*17534*/;
assign _4435_ = _4030_ & _4432_ /*17529*/;
assign _4436_ = _4030_ ^ _4432_ /*17532*/;
assign _4437_ = _4428_ & _4436_ /*17530*/;
assign _4254_ = _4428_ ^ _4436_ /*17531*/;
assign _4434_ = _4435_ | _4437_ /*17528*/;
assign _4439_ = ~Q[22] /*17527*/;
assign _4438_ = _4439_ & D[30] /*17526*/;
assign _4441_ = _4031_ & _4438_ /*17521*/;
assign _4442_ = _4031_ ^ _4438_ /*17524*/;
assign _4443_ = _4434_ & _4442_ /*17522*/;
assign _4255_ = _4434_ ^ _4442_ /*17523*/;
assign _4440_ = _4441_ | _4443_ /*17520*/;
assign _4445_ = ~Q[22] /*17519*/;
assign _4444_ = _4445_ & zeroWire /*17518*/;
assign _4446_ = _4032_ ^ _4444_ /*17516*/;
assign _4256_ = _4446_ ^ _4440_ /*17515*/;
assign _4485_ = ~D[0] /*17389*/;
assign _4482_ = R_0[21] & _4485_ /*17385*/;
assign _4483_ = R_0[21] ^ _4485_ /*17388*/;
assign _4484_ = oneWire & _4483_ /*17386*/;
assign _4449_ = oneWire ^ _4483_ /*17387*/;
assign _4481_ = _4482_ | _4484_ /*17384*/;
assign _4490_ = ~D[1] /*17383*/;
assign _4487_ = _4225_ & _4490_ /*17379*/;
assign _4488_ = _4225_ ^ _4490_ /*17382*/;
assign _4489_ = _4481_ & _4488_ /*17380*/;
assign _4450_ = _4481_ ^ _4488_ /*17381*/;
assign _4486_ = _4487_ | _4489_ /*17378*/;
assign _4495_ = ~D[2] /*17377*/;
assign _4492_ = _4226_ & _4495_ /*17373*/;
assign _4493_ = _4226_ ^ _4495_ /*17376*/;
assign _4494_ = _4486_ & _4493_ /*17374*/;
assign _4451_ = _4486_ ^ _4493_ /*17375*/;
assign _4491_ = _4492_ | _4494_ /*17372*/;
assign _4500_ = ~D[3] /*17371*/;
assign _4497_ = _4227_ & _4500_ /*17367*/;
assign _4498_ = _4227_ ^ _4500_ /*17370*/;
assign _4499_ = _4491_ & _4498_ /*17368*/;
assign _4452_ = _4491_ ^ _4498_ /*17369*/;
assign _4496_ = _4497_ | _4499_ /*17366*/;
assign _4505_ = ~D[4] /*17365*/;
assign _4502_ = _4228_ & _4505_ /*17361*/;
assign _4503_ = _4228_ ^ _4505_ /*17364*/;
assign _4504_ = _4496_ & _4503_ /*17362*/;
assign _4453_ = _4496_ ^ _4503_ /*17363*/;
assign _4501_ = _4502_ | _4504_ /*17360*/;
assign _4510_ = ~D[5] /*17359*/;
assign _4507_ = _4229_ & _4510_ /*17355*/;
assign _4508_ = _4229_ ^ _4510_ /*17358*/;
assign _4509_ = _4501_ & _4508_ /*17356*/;
assign _4454_ = _4501_ ^ _4508_ /*17357*/;
assign _4506_ = _4507_ | _4509_ /*17354*/;
assign _4515_ = ~D[6] /*17353*/;
assign _4512_ = _4230_ & _4515_ /*17349*/;
assign _4513_ = _4230_ ^ _4515_ /*17352*/;
assign _4514_ = _4506_ & _4513_ /*17350*/;
assign _4455_ = _4506_ ^ _4513_ /*17351*/;
assign _4511_ = _4512_ | _4514_ /*17348*/;
assign _4520_ = ~D[7] /*17347*/;
assign _4517_ = _4231_ & _4520_ /*17343*/;
assign _4518_ = _4231_ ^ _4520_ /*17346*/;
assign _4519_ = _4511_ & _4518_ /*17344*/;
assign _4456_ = _4511_ ^ _4518_ /*17345*/;
assign _4516_ = _4517_ | _4519_ /*17342*/;
assign _4525_ = ~D[8] /*17341*/;
assign _4522_ = _4232_ & _4525_ /*17337*/;
assign _4523_ = _4232_ ^ _4525_ /*17340*/;
assign _4524_ = _4516_ & _4523_ /*17338*/;
assign _4457_ = _4516_ ^ _4523_ /*17339*/;
assign _4521_ = _4522_ | _4524_ /*17336*/;
assign _4530_ = ~D[9] /*17335*/;
assign _4527_ = _4233_ & _4530_ /*17331*/;
assign _4528_ = _4233_ ^ _4530_ /*17334*/;
assign _4529_ = _4521_ & _4528_ /*17332*/;
assign _4458_ = _4521_ ^ _4528_ /*17333*/;
assign _4526_ = _4527_ | _4529_ /*17330*/;
assign _4535_ = ~D[10] /*17329*/;
assign _4532_ = _4234_ & _4535_ /*17325*/;
assign _4533_ = _4234_ ^ _4535_ /*17328*/;
assign _4534_ = _4526_ & _4533_ /*17326*/;
assign _4459_ = _4526_ ^ _4533_ /*17327*/;
assign _4531_ = _4532_ | _4534_ /*17324*/;
assign _4540_ = ~D[11] /*17323*/;
assign _4537_ = _4235_ & _4540_ /*17319*/;
assign _4538_ = _4235_ ^ _4540_ /*17322*/;
assign _4539_ = _4531_ & _4538_ /*17320*/;
assign _4460_ = _4531_ ^ _4538_ /*17321*/;
assign _4536_ = _4537_ | _4539_ /*17318*/;
assign _4545_ = ~D[12] /*17317*/;
assign _4542_ = _4236_ & _4545_ /*17313*/;
assign _4543_ = _4236_ ^ _4545_ /*17316*/;
assign _4544_ = _4536_ & _4543_ /*17314*/;
assign _4461_ = _4536_ ^ _4543_ /*17315*/;
assign _4541_ = _4542_ | _4544_ /*17312*/;
assign _4550_ = ~D[13] /*17311*/;
assign _4547_ = _4237_ & _4550_ /*17307*/;
assign _4548_ = _4237_ ^ _4550_ /*17310*/;
assign _4549_ = _4541_ & _4548_ /*17308*/;
assign _4462_ = _4541_ ^ _4548_ /*17309*/;
assign _4546_ = _4547_ | _4549_ /*17306*/;
assign _4555_ = ~D[14] /*17305*/;
assign _4552_ = _4238_ & _4555_ /*17301*/;
assign _4553_ = _4238_ ^ _4555_ /*17304*/;
assign _4554_ = _4546_ & _4553_ /*17302*/;
assign _4463_ = _4546_ ^ _4553_ /*17303*/;
assign _4551_ = _4552_ | _4554_ /*17300*/;
assign _4560_ = ~D[15] /*17299*/;
assign _4557_ = _4239_ & _4560_ /*17295*/;
assign _4558_ = _4239_ ^ _4560_ /*17298*/;
assign _4559_ = _4551_ & _4558_ /*17296*/;
assign _4464_ = _4551_ ^ _4558_ /*17297*/;
assign _4556_ = _4557_ | _4559_ /*17294*/;
assign _4565_ = ~D[16] /*17293*/;
assign _4562_ = _4240_ & _4565_ /*17289*/;
assign _4563_ = _4240_ ^ _4565_ /*17292*/;
assign _4564_ = _4556_ & _4563_ /*17290*/;
assign _4465_ = _4556_ ^ _4563_ /*17291*/;
assign _4561_ = _4562_ | _4564_ /*17288*/;
assign _4570_ = ~D[17] /*17287*/;
assign _4567_ = _4241_ & _4570_ /*17283*/;
assign _4568_ = _4241_ ^ _4570_ /*17286*/;
assign _4569_ = _4561_ & _4568_ /*17284*/;
assign _4466_ = _4561_ ^ _4568_ /*17285*/;
assign _4566_ = _4567_ | _4569_ /*17282*/;
assign _4575_ = ~D[18] /*17281*/;
assign _4572_ = _4242_ & _4575_ /*17277*/;
assign _4573_ = _4242_ ^ _4575_ /*17280*/;
assign _4574_ = _4566_ & _4573_ /*17278*/;
assign _4467_ = _4566_ ^ _4573_ /*17279*/;
assign _4571_ = _4572_ | _4574_ /*17276*/;
assign _4580_ = ~D[19] /*17275*/;
assign _4577_ = _4243_ & _4580_ /*17271*/;
assign _4578_ = _4243_ ^ _4580_ /*17274*/;
assign _4579_ = _4571_ & _4578_ /*17272*/;
assign _4468_ = _4571_ ^ _4578_ /*17273*/;
assign _4576_ = _4577_ | _4579_ /*17270*/;
assign _4585_ = ~D[20] /*17269*/;
assign _4582_ = _4244_ & _4585_ /*17265*/;
assign _4583_ = _4244_ ^ _4585_ /*17268*/;
assign _4584_ = _4576_ & _4583_ /*17266*/;
assign _4469_ = _4576_ ^ _4583_ /*17267*/;
assign _4581_ = _4582_ | _4584_ /*17264*/;
assign _4590_ = ~D[21] /*17263*/;
assign _4587_ = _4245_ & _4590_ /*17259*/;
assign _4588_ = _4245_ ^ _4590_ /*17262*/;
assign _4589_ = _4581_ & _4588_ /*17260*/;
assign _4470_ = _4581_ ^ _4588_ /*17261*/;
assign _4586_ = _4587_ | _4589_ /*17258*/;
assign _4595_ = ~D[22] /*17257*/;
assign _4592_ = _4246_ & _4595_ /*17253*/;
assign _4593_ = _4246_ ^ _4595_ /*17256*/;
assign _4594_ = _4586_ & _4593_ /*17254*/;
assign _4471_ = _4586_ ^ _4593_ /*17255*/;
assign _4591_ = _4592_ | _4594_ /*17252*/;
assign _4600_ = ~D[23] /*17251*/;
assign _4597_ = _4247_ & _4600_ /*17247*/;
assign _4598_ = _4247_ ^ _4600_ /*17250*/;
assign _4599_ = _4591_ & _4598_ /*17248*/;
assign _4472_ = _4591_ ^ _4598_ /*17249*/;
assign _4596_ = _4597_ | _4599_ /*17246*/;
assign _4605_ = ~D[24] /*17245*/;
assign _4602_ = _4248_ & _4605_ /*17241*/;
assign _4603_ = _4248_ ^ _4605_ /*17244*/;
assign _4604_ = _4596_ & _4603_ /*17242*/;
assign _4473_ = _4596_ ^ _4603_ /*17243*/;
assign _4601_ = _4602_ | _4604_ /*17240*/;
assign _4610_ = ~D[25] /*17239*/;
assign _4607_ = _4249_ & _4610_ /*17235*/;
assign _4608_ = _4249_ ^ _4610_ /*17238*/;
assign _4609_ = _4601_ & _4608_ /*17236*/;
assign _4474_ = _4601_ ^ _4608_ /*17237*/;
assign _4606_ = _4607_ | _4609_ /*17234*/;
assign _4615_ = ~D[26] /*17233*/;
assign _4612_ = _4250_ & _4615_ /*17229*/;
assign _4613_ = _4250_ ^ _4615_ /*17232*/;
assign _4614_ = _4606_ & _4613_ /*17230*/;
assign _4475_ = _4606_ ^ _4613_ /*17231*/;
assign _4611_ = _4612_ | _4614_ /*17228*/;
assign _4620_ = ~D[27] /*17227*/;
assign _4617_ = _4251_ & _4620_ /*17223*/;
assign _4618_ = _4251_ ^ _4620_ /*17226*/;
assign _4619_ = _4611_ & _4618_ /*17224*/;
assign _4476_ = _4611_ ^ _4618_ /*17225*/;
assign _4616_ = _4617_ | _4619_ /*17222*/;
assign _4625_ = ~D[28] /*17221*/;
assign _4622_ = _4252_ & _4625_ /*17217*/;
assign _4623_ = _4252_ ^ _4625_ /*17220*/;
assign _4624_ = _4616_ & _4623_ /*17218*/;
assign _4477_ = _4616_ ^ _4623_ /*17219*/;
assign _4621_ = _4622_ | _4624_ /*17216*/;
assign _4630_ = ~D[29] /*17215*/;
assign _4627_ = _4253_ & _4630_ /*17211*/;
assign _4628_ = _4253_ ^ _4630_ /*17214*/;
assign _4629_ = _4621_ & _4628_ /*17212*/;
assign _4478_ = _4621_ ^ _4628_ /*17213*/;
assign _4626_ = _4627_ | _4629_ /*17210*/;
assign _4635_ = ~D[30] /*17209*/;
assign _4632_ = _4254_ & _4635_ /*17205*/;
assign _4633_ = _4254_ ^ _4635_ /*17208*/;
assign _4634_ = _4626_ & _4633_ /*17206*/;
assign _4479_ = _4626_ ^ _4633_ /*17207*/;
assign _4631_ = _4632_ | _4634_ /*17204*/;
assign _4636_ = _4255_ & oneWire /*17199*/;
assign _4637_ = _4255_ ^ oneWire /*17202*/;
assign _4638_ = _4631_ & _4637_ /*17200*/;
assign _4480_ = _4631_ ^ _4637_ /*17201*/;
assign Q[21] = _4636_ | _4638_ /*17198*/;
assign _4707_ = ~Q[21] /*17005*/;
assign _4706_ = _4707_ & D[0] /*17004*/;
assign _4709_ = _4449_ & _4706_ /*16999*/;
assign _4710_ = _4449_ ^ _4706_ /*17002*/;
assign _4711_ = zeroWire & _4710_ /*17000*/;
assign _4673_ = zeroWire ^ _4710_ /*17001*/;
assign _4708_ = _4709_ | _4711_ /*16998*/;
assign _4713_ = ~Q[21] /*16997*/;
assign _4712_ = _4713_ & D[1] /*16996*/;
assign _4715_ = _4450_ & _4712_ /*16991*/;
assign _4716_ = _4450_ ^ _4712_ /*16994*/;
assign _4717_ = _4708_ & _4716_ /*16992*/;
assign _4674_ = _4708_ ^ _4716_ /*16993*/;
assign _4714_ = _4715_ | _4717_ /*16990*/;
assign _4719_ = ~Q[21] /*16989*/;
assign _4718_ = _4719_ & D[2] /*16988*/;
assign _4721_ = _4451_ & _4718_ /*16983*/;
assign _4722_ = _4451_ ^ _4718_ /*16986*/;
assign _4723_ = _4714_ & _4722_ /*16984*/;
assign _4675_ = _4714_ ^ _4722_ /*16985*/;
assign _4720_ = _4721_ | _4723_ /*16982*/;
assign _4725_ = ~Q[21] /*16981*/;
assign _4724_ = _4725_ & D[3] /*16980*/;
assign _4727_ = _4452_ & _4724_ /*16975*/;
assign _4728_ = _4452_ ^ _4724_ /*16978*/;
assign _4729_ = _4720_ & _4728_ /*16976*/;
assign _4676_ = _4720_ ^ _4728_ /*16977*/;
assign _4726_ = _4727_ | _4729_ /*16974*/;
assign _4731_ = ~Q[21] /*16973*/;
assign _4730_ = _4731_ & D[4] /*16972*/;
assign _4733_ = _4453_ & _4730_ /*16967*/;
assign _4734_ = _4453_ ^ _4730_ /*16970*/;
assign _4735_ = _4726_ & _4734_ /*16968*/;
assign _4677_ = _4726_ ^ _4734_ /*16969*/;
assign _4732_ = _4733_ | _4735_ /*16966*/;
assign _4737_ = ~Q[21] /*16965*/;
assign _4736_ = _4737_ & D[5] /*16964*/;
assign _4739_ = _4454_ & _4736_ /*16959*/;
assign _4740_ = _4454_ ^ _4736_ /*16962*/;
assign _4741_ = _4732_ & _4740_ /*16960*/;
assign _4678_ = _4732_ ^ _4740_ /*16961*/;
assign _4738_ = _4739_ | _4741_ /*16958*/;
assign _4743_ = ~Q[21] /*16957*/;
assign _4742_ = _4743_ & D[6] /*16956*/;
assign _4745_ = _4455_ & _4742_ /*16951*/;
assign _4746_ = _4455_ ^ _4742_ /*16954*/;
assign _4747_ = _4738_ & _4746_ /*16952*/;
assign _4679_ = _4738_ ^ _4746_ /*16953*/;
assign _4744_ = _4745_ | _4747_ /*16950*/;
assign _4749_ = ~Q[21] /*16949*/;
assign _4748_ = _4749_ & D[7] /*16948*/;
assign _4751_ = _4456_ & _4748_ /*16943*/;
assign _4752_ = _4456_ ^ _4748_ /*16946*/;
assign _4753_ = _4744_ & _4752_ /*16944*/;
assign _4680_ = _4744_ ^ _4752_ /*16945*/;
assign _4750_ = _4751_ | _4753_ /*16942*/;
assign _4755_ = ~Q[21] /*16941*/;
assign _4754_ = _4755_ & D[8] /*16940*/;
assign _4757_ = _4457_ & _4754_ /*16935*/;
assign _4758_ = _4457_ ^ _4754_ /*16938*/;
assign _4759_ = _4750_ & _4758_ /*16936*/;
assign _4681_ = _4750_ ^ _4758_ /*16937*/;
assign _4756_ = _4757_ | _4759_ /*16934*/;
assign _4761_ = ~Q[21] /*16933*/;
assign _4760_ = _4761_ & D[9] /*16932*/;
assign _4763_ = _4458_ & _4760_ /*16927*/;
assign _4764_ = _4458_ ^ _4760_ /*16930*/;
assign _4765_ = _4756_ & _4764_ /*16928*/;
assign _4682_ = _4756_ ^ _4764_ /*16929*/;
assign _4762_ = _4763_ | _4765_ /*16926*/;
assign _4767_ = ~Q[21] /*16925*/;
assign _4766_ = _4767_ & D[10] /*16924*/;
assign _4769_ = _4459_ & _4766_ /*16919*/;
assign _4770_ = _4459_ ^ _4766_ /*16922*/;
assign _4771_ = _4762_ & _4770_ /*16920*/;
assign _4683_ = _4762_ ^ _4770_ /*16921*/;
assign _4768_ = _4769_ | _4771_ /*16918*/;
assign _4773_ = ~Q[21] /*16917*/;
assign _4772_ = _4773_ & D[11] /*16916*/;
assign _4775_ = _4460_ & _4772_ /*16911*/;
assign _4776_ = _4460_ ^ _4772_ /*16914*/;
assign _4777_ = _4768_ & _4776_ /*16912*/;
assign _4684_ = _4768_ ^ _4776_ /*16913*/;
assign _4774_ = _4775_ | _4777_ /*16910*/;
assign _4779_ = ~Q[21] /*16909*/;
assign _4778_ = _4779_ & D[12] /*16908*/;
assign _4781_ = _4461_ & _4778_ /*16903*/;
assign _4782_ = _4461_ ^ _4778_ /*16906*/;
assign _4783_ = _4774_ & _4782_ /*16904*/;
assign _4685_ = _4774_ ^ _4782_ /*16905*/;
assign _4780_ = _4781_ | _4783_ /*16902*/;
assign _4785_ = ~Q[21] /*16901*/;
assign _4784_ = _4785_ & D[13] /*16900*/;
assign _4787_ = _4462_ & _4784_ /*16895*/;
assign _4788_ = _4462_ ^ _4784_ /*16898*/;
assign _4789_ = _4780_ & _4788_ /*16896*/;
assign _4686_ = _4780_ ^ _4788_ /*16897*/;
assign _4786_ = _4787_ | _4789_ /*16894*/;
assign _4791_ = ~Q[21] /*16893*/;
assign _4790_ = _4791_ & D[14] /*16892*/;
assign _4793_ = _4463_ & _4790_ /*16887*/;
assign _4794_ = _4463_ ^ _4790_ /*16890*/;
assign _4795_ = _4786_ & _4794_ /*16888*/;
assign _4687_ = _4786_ ^ _4794_ /*16889*/;
assign _4792_ = _4793_ | _4795_ /*16886*/;
assign _4797_ = ~Q[21] /*16885*/;
assign _4796_ = _4797_ & D[15] /*16884*/;
assign _4799_ = _4464_ & _4796_ /*16879*/;
assign _4800_ = _4464_ ^ _4796_ /*16882*/;
assign _4801_ = _4792_ & _4800_ /*16880*/;
assign _4688_ = _4792_ ^ _4800_ /*16881*/;
assign _4798_ = _4799_ | _4801_ /*16878*/;
assign _4803_ = ~Q[21] /*16877*/;
assign _4802_ = _4803_ & D[16] /*16876*/;
assign _4805_ = _4465_ & _4802_ /*16871*/;
assign _4806_ = _4465_ ^ _4802_ /*16874*/;
assign _4807_ = _4798_ & _4806_ /*16872*/;
assign _4689_ = _4798_ ^ _4806_ /*16873*/;
assign _4804_ = _4805_ | _4807_ /*16870*/;
assign _4809_ = ~Q[21] /*16869*/;
assign _4808_ = _4809_ & D[17] /*16868*/;
assign _4811_ = _4466_ & _4808_ /*16863*/;
assign _4812_ = _4466_ ^ _4808_ /*16866*/;
assign _4813_ = _4804_ & _4812_ /*16864*/;
assign _4690_ = _4804_ ^ _4812_ /*16865*/;
assign _4810_ = _4811_ | _4813_ /*16862*/;
assign _4815_ = ~Q[21] /*16861*/;
assign _4814_ = _4815_ & D[18] /*16860*/;
assign _4817_ = _4467_ & _4814_ /*16855*/;
assign _4818_ = _4467_ ^ _4814_ /*16858*/;
assign _4819_ = _4810_ & _4818_ /*16856*/;
assign _4691_ = _4810_ ^ _4818_ /*16857*/;
assign _4816_ = _4817_ | _4819_ /*16854*/;
assign _4821_ = ~Q[21] /*16853*/;
assign _4820_ = _4821_ & D[19] /*16852*/;
assign _4823_ = _4468_ & _4820_ /*16847*/;
assign _4824_ = _4468_ ^ _4820_ /*16850*/;
assign _4825_ = _4816_ & _4824_ /*16848*/;
assign _4692_ = _4816_ ^ _4824_ /*16849*/;
assign _4822_ = _4823_ | _4825_ /*16846*/;
assign _4827_ = ~Q[21] /*16845*/;
assign _4826_ = _4827_ & D[20] /*16844*/;
assign _4829_ = _4469_ & _4826_ /*16839*/;
assign _4830_ = _4469_ ^ _4826_ /*16842*/;
assign _4831_ = _4822_ & _4830_ /*16840*/;
assign _4693_ = _4822_ ^ _4830_ /*16841*/;
assign _4828_ = _4829_ | _4831_ /*16838*/;
assign _4833_ = ~Q[21] /*16837*/;
assign _4832_ = _4833_ & D[21] /*16836*/;
assign _4835_ = _4470_ & _4832_ /*16831*/;
assign _4836_ = _4470_ ^ _4832_ /*16834*/;
assign _4837_ = _4828_ & _4836_ /*16832*/;
assign _4694_ = _4828_ ^ _4836_ /*16833*/;
assign _4834_ = _4835_ | _4837_ /*16830*/;
assign _4839_ = ~Q[21] /*16829*/;
assign _4838_ = _4839_ & D[22] /*16828*/;
assign _4841_ = _4471_ & _4838_ /*16823*/;
assign _4842_ = _4471_ ^ _4838_ /*16826*/;
assign _4843_ = _4834_ & _4842_ /*16824*/;
assign _4695_ = _4834_ ^ _4842_ /*16825*/;
assign _4840_ = _4841_ | _4843_ /*16822*/;
assign _4845_ = ~Q[21] /*16821*/;
assign _4844_ = _4845_ & D[23] /*16820*/;
assign _4847_ = _4472_ & _4844_ /*16815*/;
assign _4848_ = _4472_ ^ _4844_ /*16818*/;
assign _4849_ = _4840_ & _4848_ /*16816*/;
assign _4696_ = _4840_ ^ _4848_ /*16817*/;
assign _4846_ = _4847_ | _4849_ /*16814*/;
assign _4851_ = ~Q[21] /*16813*/;
assign _4850_ = _4851_ & D[24] /*16812*/;
assign _4853_ = _4473_ & _4850_ /*16807*/;
assign _4854_ = _4473_ ^ _4850_ /*16810*/;
assign _4855_ = _4846_ & _4854_ /*16808*/;
assign _4697_ = _4846_ ^ _4854_ /*16809*/;
assign _4852_ = _4853_ | _4855_ /*16806*/;
assign _4857_ = ~Q[21] /*16805*/;
assign _4856_ = _4857_ & D[25] /*16804*/;
assign _4859_ = _4474_ & _4856_ /*16799*/;
assign _4860_ = _4474_ ^ _4856_ /*16802*/;
assign _4861_ = _4852_ & _4860_ /*16800*/;
assign _4698_ = _4852_ ^ _4860_ /*16801*/;
assign _4858_ = _4859_ | _4861_ /*16798*/;
assign _4863_ = ~Q[21] /*16797*/;
assign _4862_ = _4863_ & D[26] /*16796*/;
assign _4865_ = _4475_ & _4862_ /*16791*/;
assign _4866_ = _4475_ ^ _4862_ /*16794*/;
assign _4867_ = _4858_ & _4866_ /*16792*/;
assign _4699_ = _4858_ ^ _4866_ /*16793*/;
assign _4864_ = _4865_ | _4867_ /*16790*/;
assign _4869_ = ~Q[21] /*16789*/;
assign _4868_ = _4869_ & D[27] /*16788*/;
assign _4871_ = _4476_ & _4868_ /*16783*/;
assign _4872_ = _4476_ ^ _4868_ /*16786*/;
assign _4873_ = _4864_ & _4872_ /*16784*/;
assign _4700_ = _4864_ ^ _4872_ /*16785*/;
assign _4870_ = _4871_ | _4873_ /*16782*/;
assign _4875_ = ~Q[21] /*16781*/;
assign _4874_ = _4875_ & D[28] /*16780*/;
assign _4877_ = _4477_ & _4874_ /*16775*/;
assign _4878_ = _4477_ ^ _4874_ /*16778*/;
assign _4879_ = _4870_ & _4878_ /*16776*/;
assign _4701_ = _4870_ ^ _4878_ /*16777*/;
assign _4876_ = _4877_ | _4879_ /*16774*/;
assign _4881_ = ~Q[21] /*16773*/;
assign _4880_ = _4881_ & D[29] /*16772*/;
assign _4883_ = _4478_ & _4880_ /*16767*/;
assign _4884_ = _4478_ ^ _4880_ /*16770*/;
assign _4885_ = _4876_ & _4884_ /*16768*/;
assign _4702_ = _4876_ ^ _4884_ /*16769*/;
assign _4882_ = _4883_ | _4885_ /*16766*/;
assign _4887_ = ~Q[21] /*16765*/;
assign _4886_ = _4887_ & D[30] /*16764*/;
assign _4889_ = _4479_ & _4886_ /*16759*/;
assign _4890_ = _4479_ ^ _4886_ /*16762*/;
assign _4891_ = _4882_ & _4890_ /*16760*/;
assign _4703_ = _4882_ ^ _4890_ /*16761*/;
assign _4888_ = _4889_ | _4891_ /*16758*/;
assign _4893_ = ~Q[21] /*16757*/;
assign _4892_ = _4893_ & zeroWire /*16756*/;
assign _4894_ = _4480_ ^ _4892_ /*16754*/;
assign _4704_ = _4894_ ^ _4888_ /*16753*/;
assign _4933_ = ~D[0] /*16627*/;
assign _4930_ = R_0[20] & _4933_ /*16623*/;
assign _4931_ = R_0[20] ^ _4933_ /*16626*/;
assign _4932_ = oneWire & _4931_ /*16624*/;
assign _4897_ = oneWire ^ _4931_ /*16625*/;
assign _4929_ = _4930_ | _4932_ /*16622*/;
assign _4938_ = ~D[1] /*16621*/;
assign _4935_ = _4673_ & _4938_ /*16617*/;
assign _4936_ = _4673_ ^ _4938_ /*16620*/;
assign _4937_ = _4929_ & _4936_ /*16618*/;
assign _4898_ = _4929_ ^ _4936_ /*16619*/;
assign _4934_ = _4935_ | _4937_ /*16616*/;
assign _4943_ = ~D[2] /*16615*/;
assign _4940_ = _4674_ & _4943_ /*16611*/;
assign _4941_ = _4674_ ^ _4943_ /*16614*/;
assign _4942_ = _4934_ & _4941_ /*16612*/;
assign _4899_ = _4934_ ^ _4941_ /*16613*/;
assign _4939_ = _4940_ | _4942_ /*16610*/;
assign _4948_ = ~D[3] /*16609*/;
assign _4945_ = _4675_ & _4948_ /*16605*/;
assign _4946_ = _4675_ ^ _4948_ /*16608*/;
assign _4947_ = _4939_ & _4946_ /*16606*/;
assign _4900_ = _4939_ ^ _4946_ /*16607*/;
assign _4944_ = _4945_ | _4947_ /*16604*/;
assign _4953_ = ~D[4] /*16603*/;
assign _4950_ = _4676_ & _4953_ /*16599*/;
assign _4951_ = _4676_ ^ _4953_ /*16602*/;
assign _4952_ = _4944_ & _4951_ /*16600*/;
assign _4901_ = _4944_ ^ _4951_ /*16601*/;
assign _4949_ = _4950_ | _4952_ /*16598*/;
assign _4958_ = ~D[5] /*16597*/;
assign _4955_ = _4677_ & _4958_ /*16593*/;
assign _4956_ = _4677_ ^ _4958_ /*16596*/;
assign _4957_ = _4949_ & _4956_ /*16594*/;
assign _4902_ = _4949_ ^ _4956_ /*16595*/;
assign _4954_ = _4955_ | _4957_ /*16592*/;
assign _4963_ = ~D[6] /*16591*/;
assign _4960_ = _4678_ & _4963_ /*16587*/;
assign _4961_ = _4678_ ^ _4963_ /*16590*/;
assign _4962_ = _4954_ & _4961_ /*16588*/;
assign _4903_ = _4954_ ^ _4961_ /*16589*/;
assign _4959_ = _4960_ | _4962_ /*16586*/;
assign _4968_ = ~D[7] /*16585*/;
assign _4965_ = _4679_ & _4968_ /*16581*/;
assign _4966_ = _4679_ ^ _4968_ /*16584*/;
assign _4967_ = _4959_ & _4966_ /*16582*/;
assign _4904_ = _4959_ ^ _4966_ /*16583*/;
assign _4964_ = _4965_ | _4967_ /*16580*/;
assign _4973_ = ~D[8] /*16579*/;
assign _4970_ = _4680_ & _4973_ /*16575*/;
assign _4971_ = _4680_ ^ _4973_ /*16578*/;
assign _4972_ = _4964_ & _4971_ /*16576*/;
assign _4905_ = _4964_ ^ _4971_ /*16577*/;
assign _4969_ = _4970_ | _4972_ /*16574*/;
assign _4978_ = ~D[9] /*16573*/;
assign _4975_ = _4681_ & _4978_ /*16569*/;
assign _4976_ = _4681_ ^ _4978_ /*16572*/;
assign _4977_ = _4969_ & _4976_ /*16570*/;
assign _4906_ = _4969_ ^ _4976_ /*16571*/;
assign _4974_ = _4975_ | _4977_ /*16568*/;
assign _4983_ = ~D[10] /*16567*/;
assign _4980_ = _4682_ & _4983_ /*16563*/;
assign _4981_ = _4682_ ^ _4983_ /*16566*/;
assign _4982_ = _4974_ & _4981_ /*16564*/;
assign _4907_ = _4974_ ^ _4981_ /*16565*/;
assign _4979_ = _4980_ | _4982_ /*16562*/;
assign _4988_ = ~D[11] /*16561*/;
assign _4985_ = _4683_ & _4988_ /*16557*/;
assign _4986_ = _4683_ ^ _4988_ /*16560*/;
assign _4987_ = _4979_ & _4986_ /*16558*/;
assign _4908_ = _4979_ ^ _4986_ /*16559*/;
assign _4984_ = _4985_ | _4987_ /*16556*/;
assign _4993_ = ~D[12] /*16555*/;
assign _4990_ = _4684_ & _4993_ /*16551*/;
assign _4991_ = _4684_ ^ _4993_ /*16554*/;
assign _4992_ = _4984_ & _4991_ /*16552*/;
assign _4909_ = _4984_ ^ _4991_ /*16553*/;
assign _4989_ = _4990_ | _4992_ /*16550*/;
assign _4998_ = ~D[13] /*16549*/;
assign _4995_ = _4685_ & _4998_ /*16545*/;
assign _4996_ = _4685_ ^ _4998_ /*16548*/;
assign _4997_ = _4989_ & _4996_ /*16546*/;
assign _4910_ = _4989_ ^ _4996_ /*16547*/;
assign _4994_ = _4995_ | _4997_ /*16544*/;
assign _5003_ = ~D[14] /*16543*/;
assign _5000_ = _4686_ & _5003_ /*16539*/;
assign _5001_ = _4686_ ^ _5003_ /*16542*/;
assign _5002_ = _4994_ & _5001_ /*16540*/;
assign _4911_ = _4994_ ^ _5001_ /*16541*/;
assign _4999_ = _5000_ | _5002_ /*16538*/;
assign _5008_ = ~D[15] /*16537*/;
assign _5005_ = _4687_ & _5008_ /*16533*/;
assign _5006_ = _4687_ ^ _5008_ /*16536*/;
assign _5007_ = _4999_ & _5006_ /*16534*/;
assign _4912_ = _4999_ ^ _5006_ /*16535*/;
assign _5004_ = _5005_ | _5007_ /*16532*/;
assign _5013_ = ~D[16] /*16531*/;
assign _5010_ = _4688_ & _5013_ /*16527*/;
assign _5011_ = _4688_ ^ _5013_ /*16530*/;
assign _5012_ = _5004_ & _5011_ /*16528*/;
assign _4913_ = _5004_ ^ _5011_ /*16529*/;
assign _5009_ = _5010_ | _5012_ /*16526*/;
assign _5018_ = ~D[17] /*16525*/;
assign _5015_ = _4689_ & _5018_ /*16521*/;
assign _5016_ = _4689_ ^ _5018_ /*16524*/;
assign _5017_ = _5009_ & _5016_ /*16522*/;
assign _4914_ = _5009_ ^ _5016_ /*16523*/;
assign _5014_ = _5015_ | _5017_ /*16520*/;
assign _5023_ = ~D[18] /*16519*/;
assign _5020_ = _4690_ & _5023_ /*16515*/;
assign _5021_ = _4690_ ^ _5023_ /*16518*/;
assign _5022_ = _5014_ & _5021_ /*16516*/;
assign _4915_ = _5014_ ^ _5021_ /*16517*/;
assign _5019_ = _5020_ | _5022_ /*16514*/;
assign _5028_ = ~D[19] /*16513*/;
assign _5025_ = _4691_ & _5028_ /*16509*/;
assign _5026_ = _4691_ ^ _5028_ /*16512*/;
assign _5027_ = _5019_ & _5026_ /*16510*/;
assign _4916_ = _5019_ ^ _5026_ /*16511*/;
assign _5024_ = _5025_ | _5027_ /*16508*/;
assign _5033_ = ~D[20] /*16507*/;
assign _5030_ = _4692_ & _5033_ /*16503*/;
assign _5031_ = _4692_ ^ _5033_ /*16506*/;
assign _5032_ = _5024_ & _5031_ /*16504*/;
assign _4917_ = _5024_ ^ _5031_ /*16505*/;
assign _5029_ = _5030_ | _5032_ /*16502*/;
assign _5038_ = ~D[21] /*16501*/;
assign _5035_ = _4693_ & _5038_ /*16497*/;
assign _5036_ = _4693_ ^ _5038_ /*16500*/;
assign _5037_ = _5029_ & _5036_ /*16498*/;
assign _4918_ = _5029_ ^ _5036_ /*16499*/;
assign _5034_ = _5035_ | _5037_ /*16496*/;
assign _5043_ = ~D[22] /*16495*/;
assign _5040_ = _4694_ & _5043_ /*16491*/;
assign _5041_ = _4694_ ^ _5043_ /*16494*/;
assign _5042_ = _5034_ & _5041_ /*16492*/;
assign _4919_ = _5034_ ^ _5041_ /*16493*/;
assign _5039_ = _5040_ | _5042_ /*16490*/;
assign _5048_ = ~D[23] /*16489*/;
assign _5045_ = _4695_ & _5048_ /*16485*/;
assign _5046_ = _4695_ ^ _5048_ /*16488*/;
assign _5047_ = _5039_ & _5046_ /*16486*/;
assign _4920_ = _5039_ ^ _5046_ /*16487*/;
assign _5044_ = _5045_ | _5047_ /*16484*/;
assign _5053_ = ~D[24] /*16483*/;
assign _5050_ = _4696_ & _5053_ /*16479*/;
assign _5051_ = _4696_ ^ _5053_ /*16482*/;
assign _5052_ = _5044_ & _5051_ /*16480*/;
assign _4921_ = _5044_ ^ _5051_ /*16481*/;
assign _5049_ = _5050_ | _5052_ /*16478*/;
assign _5058_ = ~D[25] /*16477*/;
assign _5055_ = _4697_ & _5058_ /*16473*/;
assign _5056_ = _4697_ ^ _5058_ /*16476*/;
assign _5057_ = _5049_ & _5056_ /*16474*/;
assign _4922_ = _5049_ ^ _5056_ /*16475*/;
assign _5054_ = _5055_ | _5057_ /*16472*/;
assign _5063_ = ~D[26] /*16471*/;
assign _5060_ = _4698_ & _5063_ /*16467*/;
assign _5061_ = _4698_ ^ _5063_ /*16470*/;
assign _5062_ = _5054_ & _5061_ /*16468*/;
assign _4923_ = _5054_ ^ _5061_ /*16469*/;
assign _5059_ = _5060_ | _5062_ /*16466*/;
assign _5068_ = ~D[27] /*16465*/;
assign _5065_ = _4699_ & _5068_ /*16461*/;
assign _5066_ = _4699_ ^ _5068_ /*16464*/;
assign _5067_ = _5059_ & _5066_ /*16462*/;
assign _4924_ = _5059_ ^ _5066_ /*16463*/;
assign _5064_ = _5065_ | _5067_ /*16460*/;
assign _5073_ = ~D[28] /*16459*/;
assign _5070_ = _4700_ & _5073_ /*16455*/;
assign _5071_ = _4700_ ^ _5073_ /*16458*/;
assign _5072_ = _5064_ & _5071_ /*16456*/;
assign _4925_ = _5064_ ^ _5071_ /*16457*/;
assign _5069_ = _5070_ | _5072_ /*16454*/;
assign _5078_ = ~D[29] /*16453*/;
assign _5075_ = _4701_ & _5078_ /*16449*/;
assign _5076_ = _4701_ ^ _5078_ /*16452*/;
assign _5077_ = _5069_ & _5076_ /*16450*/;
assign _4926_ = _5069_ ^ _5076_ /*16451*/;
assign _5074_ = _5075_ | _5077_ /*16448*/;
assign _5083_ = ~D[30] /*16447*/;
assign _5080_ = _4702_ & _5083_ /*16443*/;
assign _5081_ = _4702_ ^ _5083_ /*16446*/;
assign _5082_ = _5074_ & _5081_ /*16444*/;
assign _4927_ = _5074_ ^ _5081_ /*16445*/;
assign _5079_ = _5080_ | _5082_ /*16442*/;
assign _5084_ = _4703_ & oneWire /*16437*/;
assign _5085_ = _4703_ ^ oneWire /*16440*/;
assign _5086_ = _5079_ & _5085_ /*16438*/;
assign _4928_ = _5079_ ^ _5085_ /*16439*/;
assign Q[20] = _5084_ | _5086_ /*16436*/;
assign _5155_ = ~Q[20] /*16243*/;
assign _5154_ = _5155_ & D[0] /*16242*/;
assign _5157_ = _4897_ & _5154_ /*16237*/;
assign _5158_ = _4897_ ^ _5154_ /*16240*/;
assign _5159_ = zeroWire & _5158_ /*16238*/;
assign _5121_ = zeroWire ^ _5158_ /*16239*/;
assign _5156_ = _5157_ | _5159_ /*16236*/;
assign _5161_ = ~Q[20] /*16235*/;
assign _5160_ = _5161_ & D[1] /*16234*/;
assign _5163_ = _4898_ & _5160_ /*16229*/;
assign _5164_ = _4898_ ^ _5160_ /*16232*/;
assign _5165_ = _5156_ & _5164_ /*16230*/;
assign _5122_ = _5156_ ^ _5164_ /*16231*/;
assign _5162_ = _5163_ | _5165_ /*16228*/;
assign _5167_ = ~Q[20] /*16227*/;
assign _5166_ = _5167_ & D[2] /*16226*/;
assign _5169_ = _4899_ & _5166_ /*16221*/;
assign _5170_ = _4899_ ^ _5166_ /*16224*/;
assign _5171_ = _5162_ & _5170_ /*16222*/;
assign _5123_ = _5162_ ^ _5170_ /*16223*/;
assign _5168_ = _5169_ | _5171_ /*16220*/;
assign _5173_ = ~Q[20] /*16219*/;
assign _5172_ = _5173_ & D[3] /*16218*/;
assign _5175_ = _4900_ & _5172_ /*16213*/;
assign _5176_ = _4900_ ^ _5172_ /*16216*/;
assign _5177_ = _5168_ & _5176_ /*16214*/;
assign _5124_ = _5168_ ^ _5176_ /*16215*/;
assign _5174_ = _5175_ | _5177_ /*16212*/;
assign _5179_ = ~Q[20] /*16211*/;
assign _5178_ = _5179_ & D[4] /*16210*/;
assign _5181_ = _4901_ & _5178_ /*16205*/;
assign _5182_ = _4901_ ^ _5178_ /*16208*/;
assign _5183_ = _5174_ & _5182_ /*16206*/;
assign _5125_ = _5174_ ^ _5182_ /*16207*/;
assign _5180_ = _5181_ | _5183_ /*16204*/;
assign _5185_ = ~Q[20] /*16203*/;
assign _5184_ = _5185_ & D[5] /*16202*/;
assign _5187_ = _4902_ & _5184_ /*16197*/;
assign _5188_ = _4902_ ^ _5184_ /*16200*/;
assign _5189_ = _5180_ & _5188_ /*16198*/;
assign _5126_ = _5180_ ^ _5188_ /*16199*/;
assign _5186_ = _5187_ | _5189_ /*16196*/;
assign _5191_ = ~Q[20] /*16195*/;
assign _5190_ = _5191_ & D[6] /*16194*/;
assign _5193_ = _4903_ & _5190_ /*16189*/;
assign _5194_ = _4903_ ^ _5190_ /*16192*/;
assign _5195_ = _5186_ & _5194_ /*16190*/;
assign _5127_ = _5186_ ^ _5194_ /*16191*/;
assign _5192_ = _5193_ | _5195_ /*16188*/;
assign _5197_ = ~Q[20] /*16187*/;
assign _5196_ = _5197_ & D[7] /*16186*/;
assign _5199_ = _4904_ & _5196_ /*16181*/;
assign _5200_ = _4904_ ^ _5196_ /*16184*/;
assign _5201_ = _5192_ & _5200_ /*16182*/;
assign _5128_ = _5192_ ^ _5200_ /*16183*/;
assign _5198_ = _5199_ | _5201_ /*16180*/;
assign _5203_ = ~Q[20] /*16179*/;
assign _5202_ = _5203_ & D[8] /*16178*/;
assign _5205_ = _4905_ & _5202_ /*16173*/;
assign _5206_ = _4905_ ^ _5202_ /*16176*/;
assign _5207_ = _5198_ & _5206_ /*16174*/;
assign _5129_ = _5198_ ^ _5206_ /*16175*/;
assign _5204_ = _5205_ | _5207_ /*16172*/;
assign _5209_ = ~Q[20] /*16171*/;
assign _5208_ = _5209_ & D[9] /*16170*/;
assign _5211_ = _4906_ & _5208_ /*16165*/;
assign _5212_ = _4906_ ^ _5208_ /*16168*/;
assign _5213_ = _5204_ & _5212_ /*16166*/;
assign _5130_ = _5204_ ^ _5212_ /*16167*/;
assign _5210_ = _5211_ | _5213_ /*16164*/;
assign _5215_ = ~Q[20] /*16163*/;
assign _5214_ = _5215_ & D[10] /*16162*/;
assign _5217_ = _4907_ & _5214_ /*16157*/;
assign _5218_ = _4907_ ^ _5214_ /*16160*/;
assign _5219_ = _5210_ & _5218_ /*16158*/;
assign _5131_ = _5210_ ^ _5218_ /*16159*/;
assign _5216_ = _5217_ | _5219_ /*16156*/;
assign _5221_ = ~Q[20] /*16155*/;
assign _5220_ = _5221_ & D[11] /*16154*/;
assign _5223_ = _4908_ & _5220_ /*16149*/;
assign _5224_ = _4908_ ^ _5220_ /*16152*/;
assign _5225_ = _5216_ & _5224_ /*16150*/;
assign _5132_ = _5216_ ^ _5224_ /*16151*/;
assign _5222_ = _5223_ | _5225_ /*16148*/;
assign _5227_ = ~Q[20] /*16147*/;
assign _5226_ = _5227_ & D[12] /*16146*/;
assign _5229_ = _4909_ & _5226_ /*16141*/;
assign _5230_ = _4909_ ^ _5226_ /*16144*/;
assign _5231_ = _5222_ & _5230_ /*16142*/;
assign _5133_ = _5222_ ^ _5230_ /*16143*/;
assign _5228_ = _5229_ | _5231_ /*16140*/;
assign _5233_ = ~Q[20] /*16139*/;
assign _5232_ = _5233_ & D[13] /*16138*/;
assign _5235_ = _4910_ & _5232_ /*16133*/;
assign _5236_ = _4910_ ^ _5232_ /*16136*/;
assign _5237_ = _5228_ & _5236_ /*16134*/;
assign _5134_ = _5228_ ^ _5236_ /*16135*/;
assign _5234_ = _5235_ | _5237_ /*16132*/;
assign _5239_ = ~Q[20] /*16131*/;
assign _5238_ = _5239_ & D[14] /*16130*/;
assign _5241_ = _4911_ & _5238_ /*16125*/;
assign _5242_ = _4911_ ^ _5238_ /*16128*/;
assign _5243_ = _5234_ & _5242_ /*16126*/;
assign _5135_ = _5234_ ^ _5242_ /*16127*/;
assign _5240_ = _5241_ | _5243_ /*16124*/;
assign _5245_ = ~Q[20] /*16123*/;
assign _5244_ = _5245_ & D[15] /*16122*/;
assign _5247_ = _4912_ & _5244_ /*16117*/;
assign _5248_ = _4912_ ^ _5244_ /*16120*/;
assign _5249_ = _5240_ & _5248_ /*16118*/;
assign _5136_ = _5240_ ^ _5248_ /*16119*/;
assign _5246_ = _5247_ | _5249_ /*16116*/;
assign _5251_ = ~Q[20] /*16115*/;
assign _5250_ = _5251_ & D[16] /*16114*/;
assign _5253_ = _4913_ & _5250_ /*16109*/;
assign _5254_ = _4913_ ^ _5250_ /*16112*/;
assign _5255_ = _5246_ & _5254_ /*16110*/;
assign _5137_ = _5246_ ^ _5254_ /*16111*/;
assign _5252_ = _5253_ | _5255_ /*16108*/;
assign _5257_ = ~Q[20] /*16107*/;
assign _5256_ = _5257_ & D[17] /*16106*/;
assign _5259_ = _4914_ & _5256_ /*16101*/;
assign _5260_ = _4914_ ^ _5256_ /*16104*/;
assign _5261_ = _5252_ & _5260_ /*16102*/;
assign _5138_ = _5252_ ^ _5260_ /*16103*/;
assign _5258_ = _5259_ | _5261_ /*16100*/;
assign _5263_ = ~Q[20] /*16099*/;
assign _5262_ = _5263_ & D[18] /*16098*/;
assign _5265_ = _4915_ & _5262_ /*16093*/;
assign _5266_ = _4915_ ^ _5262_ /*16096*/;
assign _5267_ = _5258_ & _5266_ /*16094*/;
assign _5139_ = _5258_ ^ _5266_ /*16095*/;
assign _5264_ = _5265_ | _5267_ /*16092*/;
assign _5269_ = ~Q[20] /*16091*/;
assign _5268_ = _5269_ & D[19] /*16090*/;
assign _5271_ = _4916_ & _5268_ /*16085*/;
assign _5272_ = _4916_ ^ _5268_ /*16088*/;
assign _5273_ = _5264_ & _5272_ /*16086*/;
assign _5140_ = _5264_ ^ _5272_ /*16087*/;
assign _5270_ = _5271_ | _5273_ /*16084*/;
assign _5275_ = ~Q[20] /*16083*/;
assign _5274_ = _5275_ & D[20] /*16082*/;
assign _5277_ = _4917_ & _5274_ /*16077*/;
assign _5278_ = _4917_ ^ _5274_ /*16080*/;
assign _5279_ = _5270_ & _5278_ /*16078*/;
assign _5141_ = _5270_ ^ _5278_ /*16079*/;
assign _5276_ = _5277_ | _5279_ /*16076*/;
assign _5281_ = ~Q[20] /*16075*/;
assign _5280_ = _5281_ & D[21] /*16074*/;
assign _5283_ = _4918_ & _5280_ /*16069*/;
assign _5284_ = _4918_ ^ _5280_ /*16072*/;
assign _5285_ = _5276_ & _5284_ /*16070*/;
assign _5142_ = _5276_ ^ _5284_ /*16071*/;
assign _5282_ = _5283_ | _5285_ /*16068*/;
assign _5287_ = ~Q[20] /*16067*/;
assign _5286_ = _5287_ & D[22] /*16066*/;
assign _5289_ = _4919_ & _5286_ /*16061*/;
assign _5290_ = _4919_ ^ _5286_ /*16064*/;
assign _5291_ = _5282_ & _5290_ /*16062*/;
assign _5143_ = _5282_ ^ _5290_ /*16063*/;
assign _5288_ = _5289_ | _5291_ /*16060*/;
assign _5293_ = ~Q[20] /*16059*/;
assign _5292_ = _5293_ & D[23] /*16058*/;
assign _5295_ = _4920_ & _5292_ /*16053*/;
assign _5296_ = _4920_ ^ _5292_ /*16056*/;
assign _5297_ = _5288_ & _5296_ /*16054*/;
assign _5144_ = _5288_ ^ _5296_ /*16055*/;
assign _5294_ = _5295_ | _5297_ /*16052*/;
assign _5299_ = ~Q[20] /*16051*/;
assign _5298_ = _5299_ & D[24] /*16050*/;
assign _5301_ = _4921_ & _5298_ /*16045*/;
assign _5302_ = _4921_ ^ _5298_ /*16048*/;
assign _5303_ = _5294_ & _5302_ /*16046*/;
assign _5145_ = _5294_ ^ _5302_ /*16047*/;
assign _5300_ = _5301_ | _5303_ /*16044*/;
assign _5305_ = ~Q[20] /*16043*/;
assign _5304_ = _5305_ & D[25] /*16042*/;
assign _5307_ = _4922_ & _5304_ /*16037*/;
assign _5308_ = _4922_ ^ _5304_ /*16040*/;
assign _5309_ = _5300_ & _5308_ /*16038*/;
assign _5146_ = _5300_ ^ _5308_ /*16039*/;
assign _5306_ = _5307_ | _5309_ /*16036*/;
assign _5311_ = ~Q[20] /*16035*/;
assign _5310_ = _5311_ & D[26] /*16034*/;
assign _5313_ = _4923_ & _5310_ /*16029*/;
assign _5314_ = _4923_ ^ _5310_ /*16032*/;
assign _5315_ = _5306_ & _5314_ /*16030*/;
assign _5147_ = _5306_ ^ _5314_ /*16031*/;
assign _5312_ = _5313_ | _5315_ /*16028*/;
assign _5317_ = ~Q[20] /*16027*/;
assign _5316_ = _5317_ & D[27] /*16026*/;
assign _5319_ = _4924_ & _5316_ /*16021*/;
assign _5320_ = _4924_ ^ _5316_ /*16024*/;
assign _5321_ = _5312_ & _5320_ /*16022*/;
assign _5148_ = _5312_ ^ _5320_ /*16023*/;
assign _5318_ = _5319_ | _5321_ /*16020*/;
assign _5323_ = ~Q[20] /*16019*/;
assign _5322_ = _5323_ & D[28] /*16018*/;
assign _5325_ = _4925_ & _5322_ /*16013*/;
assign _5326_ = _4925_ ^ _5322_ /*16016*/;
assign _5327_ = _5318_ & _5326_ /*16014*/;
assign _5149_ = _5318_ ^ _5326_ /*16015*/;
assign _5324_ = _5325_ | _5327_ /*16012*/;
assign _5329_ = ~Q[20] /*16011*/;
assign _5328_ = _5329_ & D[29] /*16010*/;
assign _5331_ = _4926_ & _5328_ /*16005*/;
assign _5332_ = _4926_ ^ _5328_ /*16008*/;
assign _5333_ = _5324_ & _5332_ /*16006*/;
assign _5150_ = _5324_ ^ _5332_ /*16007*/;
assign _5330_ = _5331_ | _5333_ /*16004*/;
assign _5335_ = ~Q[20] /*16003*/;
assign _5334_ = _5335_ & D[30] /*16002*/;
assign _5337_ = _4927_ & _5334_ /*15997*/;
assign _5338_ = _4927_ ^ _5334_ /*16000*/;
assign _5339_ = _5330_ & _5338_ /*15998*/;
assign _5151_ = _5330_ ^ _5338_ /*15999*/;
assign _5336_ = _5337_ | _5339_ /*15996*/;
assign _5341_ = ~Q[20] /*15995*/;
assign _5340_ = _5341_ & zeroWire /*15994*/;
assign _5342_ = _4928_ ^ _5340_ /*15992*/;
assign _5152_ = _5342_ ^ _5336_ /*15991*/;
assign _5381_ = ~D[0] /*15865*/;
assign _5378_ = R_0[19] & _5381_ /*15861*/;
assign _5379_ = R_0[19] ^ _5381_ /*15864*/;
assign _5380_ = oneWire & _5379_ /*15862*/;
assign _5345_ = oneWire ^ _5379_ /*15863*/;
assign _5377_ = _5378_ | _5380_ /*15860*/;
assign _5386_ = ~D[1] /*15859*/;
assign _5383_ = _5121_ & _5386_ /*15855*/;
assign _5384_ = _5121_ ^ _5386_ /*15858*/;
assign _5385_ = _5377_ & _5384_ /*15856*/;
assign _5346_ = _5377_ ^ _5384_ /*15857*/;
assign _5382_ = _5383_ | _5385_ /*15854*/;
assign _5391_ = ~D[2] /*15853*/;
assign _5388_ = _5122_ & _5391_ /*15849*/;
assign _5389_ = _5122_ ^ _5391_ /*15852*/;
assign _5390_ = _5382_ & _5389_ /*15850*/;
assign _5347_ = _5382_ ^ _5389_ /*15851*/;
assign _5387_ = _5388_ | _5390_ /*15848*/;
assign _5396_ = ~D[3] /*15847*/;
assign _5393_ = _5123_ & _5396_ /*15843*/;
assign _5394_ = _5123_ ^ _5396_ /*15846*/;
assign _5395_ = _5387_ & _5394_ /*15844*/;
assign _5348_ = _5387_ ^ _5394_ /*15845*/;
assign _5392_ = _5393_ | _5395_ /*15842*/;
assign _5401_ = ~D[4] /*15841*/;
assign _5398_ = _5124_ & _5401_ /*15837*/;
assign _5399_ = _5124_ ^ _5401_ /*15840*/;
assign _5400_ = _5392_ & _5399_ /*15838*/;
assign _5349_ = _5392_ ^ _5399_ /*15839*/;
assign _5397_ = _5398_ | _5400_ /*15836*/;
assign _5406_ = ~D[5] /*15835*/;
assign _5403_ = _5125_ & _5406_ /*15831*/;
assign _5404_ = _5125_ ^ _5406_ /*15834*/;
assign _5405_ = _5397_ & _5404_ /*15832*/;
assign _5350_ = _5397_ ^ _5404_ /*15833*/;
assign _5402_ = _5403_ | _5405_ /*15830*/;
assign _5411_ = ~D[6] /*15829*/;
assign _5408_ = _5126_ & _5411_ /*15825*/;
assign _5409_ = _5126_ ^ _5411_ /*15828*/;
assign _5410_ = _5402_ & _5409_ /*15826*/;
assign _5351_ = _5402_ ^ _5409_ /*15827*/;
assign _5407_ = _5408_ | _5410_ /*15824*/;
assign _5416_ = ~D[7] /*15823*/;
assign _5413_ = _5127_ & _5416_ /*15819*/;
assign _5414_ = _5127_ ^ _5416_ /*15822*/;
assign _5415_ = _5407_ & _5414_ /*15820*/;
assign _5352_ = _5407_ ^ _5414_ /*15821*/;
assign _5412_ = _5413_ | _5415_ /*15818*/;
assign _5421_ = ~D[8] /*15817*/;
assign _5418_ = _5128_ & _5421_ /*15813*/;
assign _5419_ = _5128_ ^ _5421_ /*15816*/;
assign _5420_ = _5412_ & _5419_ /*15814*/;
assign _5353_ = _5412_ ^ _5419_ /*15815*/;
assign _5417_ = _5418_ | _5420_ /*15812*/;
assign _5426_ = ~D[9] /*15811*/;
assign _5423_ = _5129_ & _5426_ /*15807*/;
assign _5424_ = _5129_ ^ _5426_ /*15810*/;
assign _5425_ = _5417_ & _5424_ /*15808*/;
assign _5354_ = _5417_ ^ _5424_ /*15809*/;
assign _5422_ = _5423_ | _5425_ /*15806*/;
assign _5431_ = ~D[10] /*15805*/;
assign _5428_ = _5130_ & _5431_ /*15801*/;
assign _5429_ = _5130_ ^ _5431_ /*15804*/;
assign _5430_ = _5422_ & _5429_ /*15802*/;
assign _5355_ = _5422_ ^ _5429_ /*15803*/;
assign _5427_ = _5428_ | _5430_ /*15800*/;
assign _5436_ = ~D[11] /*15799*/;
assign _5433_ = _5131_ & _5436_ /*15795*/;
assign _5434_ = _5131_ ^ _5436_ /*15798*/;
assign _5435_ = _5427_ & _5434_ /*15796*/;
assign _5356_ = _5427_ ^ _5434_ /*15797*/;
assign _5432_ = _5433_ | _5435_ /*15794*/;
assign _5441_ = ~D[12] /*15793*/;
assign _5438_ = _5132_ & _5441_ /*15789*/;
assign _5439_ = _5132_ ^ _5441_ /*15792*/;
assign _5440_ = _5432_ & _5439_ /*15790*/;
assign _5357_ = _5432_ ^ _5439_ /*15791*/;
assign _5437_ = _5438_ | _5440_ /*15788*/;
assign _5446_ = ~D[13] /*15787*/;
assign _5443_ = _5133_ & _5446_ /*15783*/;
assign _5444_ = _5133_ ^ _5446_ /*15786*/;
assign _5445_ = _5437_ & _5444_ /*15784*/;
assign _5358_ = _5437_ ^ _5444_ /*15785*/;
assign _5442_ = _5443_ | _5445_ /*15782*/;
assign _5451_ = ~D[14] /*15781*/;
assign _5448_ = _5134_ & _5451_ /*15777*/;
assign _5449_ = _5134_ ^ _5451_ /*15780*/;
assign _5450_ = _5442_ & _5449_ /*15778*/;
assign _5359_ = _5442_ ^ _5449_ /*15779*/;
assign _5447_ = _5448_ | _5450_ /*15776*/;
assign _5456_ = ~D[15] /*15775*/;
assign _5453_ = _5135_ & _5456_ /*15771*/;
assign _5454_ = _5135_ ^ _5456_ /*15774*/;
assign _5455_ = _5447_ & _5454_ /*15772*/;
assign _5360_ = _5447_ ^ _5454_ /*15773*/;
assign _5452_ = _5453_ | _5455_ /*15770*/;
assign _5461_ = ~D[16] /*15769*/;
assign _5458_ = _5136_ & _5461_ /*15765*/;
assign _5459_ = _5136_ ^ _5461_ /*15768*/;
assign _5460_ = _5452_ & _5459_ /*15766*/;
assign _5361_ = _5452_ ^ _5459_ /*15767*/;
assign _5457_ = _5458_ | _5460_ /*15764*/;
assign _5466_ = ~D[17] /*15763*/;
assign _5463_ = _5137_ & _5466_ /*15759*/;
assign _5464_ = _5137_ ^ _5466_ /*15762*/;
assign _5465_ = _5457_ & _5464_ /*15760*/;
assign _5362_ = _5457_ ^ _5464_ /*15761*/;
assign _5462_ = _5463_ | _5465_ /*15758*/;
assign _5471_ = ~D[18] /*15757*/;
assign _5468_ = _5138_ & _5471_ /*15753*/;
assign _5469_ = _5138_ ^ _5471_ /*15756*/;
assign _5470_ = _5462_ & _5469_ /*15754*/;
assign _5363_ = _5462_ ^ _5469_ /*15755*/;
assign _5467_ = _5468_ | _5470_ /*15752*/;
assign _5476_ = ~D[19] /*15751*/;
assign _5473_ = _5139_ & _5476_ /*15747*/;
assign _5474_ = _5139_ ^ _5476_ /*15750*/;
assign _5475_ = _5467_ & _5474_ /*15748*/;
assign _5364_ = _5467_ ^ _5474_ /*15749*/;
assign _5472_ = _5473_ | _5475_ /*15746*/;
assign _5481_ = ~D[20] /*15745*/;
assign _5478_ = _5140_ & _5481_ /*15741*/;
assign _5479_ = _5140_ ^ _5481_ /*15744*/;
assign _5480_ = _5472_ & _5479_ /*15742*/;
assign _5365_ = _5472_ ^ _5479_ /*15743*/;
assign _5477_ = _5478_ | _5480_ /*15740*/;
assign _5486_ = ~D[21] /*15739*/;
assign _5483_ = _5141_ & _5486_ /*15735*/;
assign _5484_ = _5141_ ^ _5486_ /*15738*/;
assign _5485_ = _5477_ & _5484_ /*15736*/;
assign _5366_ = _5477_ ^ _5484_ /*15737*/;
assign _5482_ = _5483_ | _5485_ /*15734*/;
assign _5491_ = ~D[22] /*15733*/;
assign _5488_ = _5142_ & _5491_ /*15729*/;
assign _5489_ = _5142_ ^ _5491_ /*15732*/;
assign _5490_ = _5482_ & _5489_ /*15730*/;
assign _5367_ = _5482_ ^ _5489_ /*15731*/;
assign _5487_ = _5488_ | _5490_ /*15728*/;
assign _5496_ = ~D[23] /*15727*/;
assign _5493_ = _5143_ & _5496_ /*15723*/;
assign _5494_ = _5143_ ^ _5496_ /*15726*/;
assign _5495_ = _5487_ & _5494_ /*15724*/;
assign _5368_ = _5487_ ^ _5494_ /*15725*/;
assign _5492_ = _5493_ | _5495_ /*15722*/;
assign _5501_ = ~D[24] /*15721*/;
assign _5498_ = _5144_ & _5501_ /*15717*/;
assign _5499_ = _5144_ ^ _5501_ /*15720*/;
assign _5500_ = _5492_ & _5499_ /*15718*/;
assign _5369_ = _5492_ ^ _5499_ /*15719*/;
assign _5497_ = _5498_ | _5500_ /*15716*/;
assign _5506_ = ~D[25] /*15715*/;
assign _5503_ = _5145_ & _5506_ /*15711*/;
assign _5504_ = _5145_ ^ _5506_ /*15714*/;
assign _5505_ = _5497_ & _5504_ /*15712*/;
assign _5370_ = _5497_ ^ _5504_ /*15713*/;
assign _5502_ = _5503_ | _5505_ /*15710*/;
assign _5511_ = ~D[26] /*15709*/;
assign _5508_ = _5146_ & _5511_ /*15705*/;
assign _5509_ = _5146_ ^ _5511_ /*15708*/;
assign _5510_ = _5502_ & _5509_ /*15706*/;
assign _5371_ = _5502_ ^ _5509_ /*15707*/;
assign _5507_ = _5508_ | _5510_ /*15704*/;
assign _5516_ = ~D[27] /*15703*/;
assign _5513_ = _5147_ & _5516_ /*15699*/;
assign _5514_ = _5147_ ^ _5516_ /*15702*/;
assign _5515_ = _5507_ & _5514_ /*15700*/;
assign _5372_ = _5507_ ^ _5514_ /*15701*/;
assign _5512_ = _5513_ | _5515_ /*15698*/;
assign _5521_ = ~D[28] /*15697*/;
assign _5518_ = _5148_ & _5521_ /*15693*/;
assign _5519_ = _5148_ ^ _5521_ /*15696*/;
assign _5520_ = _5512_ & _5519_ /*15694*/;
assign _5373_ = _5512_ ^ _5519_ /*15695*/;
assign _5517_ = _5518_ | _5520_ /*15692*/;
assign _5526_ = ~D[29] /*15691*/;
assign _5523_ = _5149_ & _5526_ /*15687*/;
assign _5524_ = _5149_ ^ _5526_ /*15690*/;
assign _5525_ = _5517_ & _5524_ /*15688*/;
assign _5374_ = _5517_ ^ _5524_ /*15689*/;
assign _5522_ = _5523_ | _5525_ /*15686*/;
assign _5531_ = ~D[30] /*15685*/;
assign _5528_ = _5150_ & _5531_ /*15681*/;
assign _5529_ = _5150_ ^ _5531_ /*15684*/;
assign _5530_ = _5522_ & _5529_ /*15682*/;
assign _5375_ = _5522_ ^ _5529_ /*15683*/;
assign _5527_ = _5528_ | _5530_ /*15680*/;
assign _5532_ = _5151_ & oneWire /*15675*/;
assign _5533_ = _5151_ ^ oneWire /*15678*/;
assign _5534_ = _5527_ & _5533_ /*15676*/;
assign _5376_ = _5527_ ^ _5533_ /*15677*/;
assign Q[19] = _5532_ | _5534_ /*15674*/;
assign _5603_ = ~Q[19] /*15481*/;
assign _5602_ = _5603_ & D[0] /*15480*/;
assign _5605_ = _5345_ & _5602_ /*15475*/;
assign _5606_ = _5345_ ^ _5602_ /*15478*/;
assign _5607_ = zeroWire & _5606_ /*15476*/;
assign _5569_ = zeroWire ^ _5606_ /*15477*/;
assign _5604_ = _5605_ | _5607_ /*15474*/;
assign _5609_ = ~Q[19] /*15473*/;
assign _5608_ = _5609_ & D[1] /*15472*/;
assign _5611_ = _5346_ & _5608_ /*15467*/;
assign _5612_ = _5346_ ^ _5608_ /*15470*/;
assign _5613_ = _5604_ & _5612_ /*15468*/;
assign _5570_ = _5604_ ^ _5612_ /*15469*/;
assign _5610_ = _5611_ | _5613_ /*15466*/;
assign _5615_ = ~Q[19] /*15465*/;
assign _5614_ = _5615_ & D[2] /*15464*/;
assign _5617_ = _5347_ & _5614_ /*15459*/;
assign _5618_ = _5347_ ^ _5614_ /*15462*/;
assign _5619_ = _5610_ & _5618_ /*15460*/;
assign _5571_ = _5610_ ^ _5618_ /*15461*/;
assign _5616_ = _5617_ | _5619_ /*15458*/;
assign _5621_ = ~Q[19] /*15457*/;
assign _5620_ = _5621_ & D[3] /*15456*/;
assign _5623_ = _5348_ & _5620_ /*15451*/;
assign _5624_ = _5348_ ^ _5620_ /*15454*/;
assign _5625_ = _5616_ & _5624_ /*15452*/;
assign _5572_ = _5616_ ^ _5624_ /*15453*/;
assign _5622_ = _5623_ | _5625_ /*15450*/;
assign _5627_ = ~Q[19] /*15449*/;
assign _5626_ = _5627_ & D[4] /*15448*/;
assign _5629_ = _5349_ & _5626_ /*15443*/;
assign _5630_ = _5349_ ^ _5626_ /*15446*/;
assign _5631_ = _5622_ & _5630_ /*15444*/;
assign _5573_ = _5622_ ^ _5630_ /*15445*/;
assign _5628_ = _5629_ | _5631_ /*15442*/;
assign _5633_ = ~Q[19] /*15441*/;
assign _5632_ = _5633_ & D[5] /*15440*/;
assign _5635_ = _5350_ & _5632_ /*15435*/;
assign _5636_ = _5350_ ^ _5632_ /*15438*/;
assign _5637_ = _5628_ & _5636_ /*15436*/;
assign _5574_ = _5628_ ^ _5636_ /*15437*/;
assign _5634_ = _5635_ | _5637_ /*15434*/;
assign _5639_ = ~Q[19] /*15433*/;
assign _5638_ = _5639_ & D[6] /*15432*/;
assign _5641_ = _5351_ & _5638_ /*15427*/;
assign _5642_ = _5351_ ^ _5638_ /*15430*/;
assign _5643_ = _5634_ & _5642_ /*15428*/;
assign _5575_ = _5634_ ^ _5642_ /*15429*/;
assign _5640_ = _5641_ | _5643_ /*15426*/;
assign _5645_ = ~Q[19] /*15425*/;
assign _5644_ = _5645_ & D[7] /*15424*/;
assign _5647_ = _5352_ & _5644_ /*15419*/;
assign _5648_ = _5352_ ^ _5644_ /*15422*/;
assign _5649_ = _5640_ & _5648_ /*15420*/;
assign _5576_ = _5640_ ^ _5648_ /*15421*/;
assign _5646_ = _5647_ | _5649_ /*15418*/;
assign _5651_ = ~Q[19] /*15417*/;
assign _5650_ = _5651_ & D[8] /*15416*/;
assign _5653_ = _5353_ & _5650_ /*15411*/;
assign _5654_ = _5353_ ^ _5650_ /*15414*/;
assign _5655_ = _5646_ & _5654_ /*15412*/;
assign _5577_ = _5646_ ^ _5654_ /*15413*/;
assign _5652_ = _5653_ | _5655_ /*15410*/;
assign _5657_ = ~Q[19] /*15409*/;
assign _5656_ = _5657_ & D[9] /*15408*/;
assign _5659_ = _5354_ & _5656_ /*15403*/;
assign _5660_ = _5354_ ^ _5656_ /*15406*/;
assign _5661_ = _5652_ & _5660_ /*15404*/;
assign _5578_ = _5652_ ^ _5660_ /*15405*/;
assign _5658_ = _5659_ | _5661_ /*15402*/;
assign _5663_ = ~Q[19] /*15401*/;
assign _5662_ = _5663_ & D[10] /*15400*/;
assign _5665_ = _5355_ & _5662_ /*15395*/;
assign _5666_ = _5355_ ^ _5662_ /*15398*/;
assign _5667_ = _5658_ & _5666_ /*15396*/;
assign _5579_ = _5658_ ^ _5666_ /*15397*/;
assign _5664_ = _5665_ | _5667_ /*15394*/;
assign _5669_ = ~Q[19] /*15393*/;
assign _5668_ = _5669_ & D[11] /*15392*/;
assign _5671_ = _5356_ & _5668_ /*15387*/;
assign _5672_ = _5356_ ^ _5668_ /*15390*/;
assign _5673_ = _5664_ & _5672_ /*15388*/;
assign _5580_ = _5664_ ^ _5672_ /*15389*/;
assign _5670_ = _5671_ | _5673_ /*15386*/;
assign _5675_ = ~Q[19] /*15385*/;
assign _5674_ = _5675_ & D[12] /*15384*/;
assign _5677_ = _5357_ & _5674_ /*15379*/;
assign _5678_ = _5357_ ^ _5674_ /*15382*/;
assign _5679_ = _5670_ & _5678_ /*15380*/;
assign _5581_ = _5670_ ^ _5678_ /*15381*/;
assign _5676_ = _5677_ | _5679_ /*15378*/;
assign _5681_ = ~Q[19] /*15377*/;
assign _5680_ = _5681_ & D[13] /*15376*/;
assign _5683_ = _5358_ & _5680_ /*15371*/;
assign _5684_ = _5358_ ^ _5680_ /*15374*/;
assign _5685_ = _5676_ & _5684_ /*15372*/;
assign _5582_ = _5676_ ^ _5684_ /*15373*/;
assign _5682_ = _5683_ | _5685_ /*15370*/;
assign _5687_ = ~Q[19] /*15369*/;
assign _5686_ = _5687_ & D[14] /*15368*/;
assign _5689_ = _5359_ & _5686_ /*15363*/;
assign _5690_ = _5359_ ^ _5686_ /*15366*/;
assign _5691_ = _5682_ & _5690_ /*15364*/;
assign _5583_ = _5682_ ^ _5690_ /*15365*/;
assign _5688_ = _5689_ | _5691_ /*15362*/;
assign _5693_ = ~Q[19] /*15361*/;
assign _5692_ = _5693_ & D[15] /*15360*/;
assign _5695_ = _5360_ & _5692_ /*15355*/;
assign _5696_ = _5360_ ^ _5692_ /*15358*/;
assign _5697_ = _5688_ & _5696_ /*15356*/;
assign _5584_ = _5688_ ^ _5696_ /*15357*/;
assign _5694_ = _5695_ | _5697_ /*15354*/;
assign _5699_ = ~Q[19] /*15353*/;
assign _5698_ = _5699_ & D[16] /*15352*/;
assign _5701_ = _5361_ & _5698_ /*15347*/;
assign _5702_ = _5361_ ^ _5698_ /*15350*/;
assign _5703_ = _5694_ & _5702_ /*15348*/;
assign _5585_ = _5694_ ^ _5702_ /*15349*/;
assign _5700_ = _5701_ | _5703_ /*15346*/;
assign _5705_ = ~Q[19] /*15345*/;
assign _5704_ = _5705_ & D[17] /*15344*/;
assign _5707_ = _5362_ & _5704_ /*15339*/;
assign _5708_ = _5362_ ^ _5704_ /*15342*/;
assign _5709_ = _5700_ & _5708_ /*15340*/;
assign _5586_ = _5700_ ^ _5708_ /*15341*/;
assign _5706_ = _5707_ | _5709_ /*15338*/;
assign _5711_ = ~Q[19] /*15337*/;
assign _5710_ = _5711_ & D[18] /*15336*/;
assign _5713_ = _5363_ & _5710_ /*15331*/;
assign _5714_ = _5363_ ^ _5710_ /*15334*/;
assign _5715_ = _5706_ & _5714_ /*15332*/;
assign _5587_ = _5706_ ^ _5714_ /*15333*/;
assign _5712_ = _5713_ | _5715_ /*15330*/;
assign _5717_ = ~Q[19] /*15329*/;
assign _5716_ = _5717_ & D[19] /*15328*/;
assign _5719_ = _5364_ & _5716_ /*15323*/;
assign _5720_ = _5364_ ^ _5716_ /*15326*/;
assign _5721_ = _5712_ & _5720_ /*15324*/;
assign _5588_ = _5712_ ^ _5720_ /*15325*/;
assign _5718_ = _5719_ | _5721_ /*15322*/;
assign _5723_ = ~Q[19] /*15321*/;
assign _5722_ = _5723_ & D[20] /*15320*/;
assign _5725_ = _5365_ & _5722_ /*15315*/;
assign _5726_ = _5365_ ^ _5722_ /*15318*/;
assign _5727_ = _5718_ & _5726_ /*15316*/;
assign _5589_ = _5718_ ^ _5726_ /*15317*/;
assign _5724_ = _5725_ | _5727_ /*15314*/;
assign _5729_ = ~Q[19] /*15313*/;
assign _5728_ = _5729_ & D[21] /*15312*/;
assign _5731_ = _5366_ & _5728_ /*15307*/;
assign _5732_ = _5366_ ^ _5728_ /*15310*/;
assign _5733_ = _5724_ & _5732_ /*15308*/;
assign _5590_ = _5724_ ^ _5732_ /*15309*/;
assign _5730_ = _5731_ | _5733_ /*15306*/;
assign _5735_ = ~Q[19] /*15305*/;
assign _5734_ = _5735_ & D[22] /*15304*/;
assign _5737_ = _5367_ & _5734_ /*15299*/;
assign _5738_ = _5367_ ^ _5734_ /*15302*/;
assign _5739_ = _5730_ & _5738_ /*15300*/;
assign _5591_ = _5730_ ^ _5738_ /*15301*/;
assign _5736_ = _5737_ | _5739_ /*15298*/;
assign _5741_ = ~Q[19] /*15297*/;
assign _5740_ = _5741_ & D[23] /*15296*/;
assign _5743_ = _5368_ & _5740_ /*15291*/;
assign _5744_ = _5368_ ^ _5740_ /*15294*/;
assign _5745_ = _5736_ & _5744_ /*15292*/;
assign _5592_ = _5736_ ^ _5744_ /*15293*/;
assign _5742_ = _5743_ | _5745_ /*15290*/;
assign _5747_ = ~Q[19] /*15289*/;
assign _5746_ = _5747_ & D[24] /*15288*/;
assign _5749_ = _5369_ & _5746_ /*15283*/;
assign _5750_ = _5369_ ^ _5746_ /*15286*/;
assign _5751_ = _5742_ & _5750_ /*15284*/;
assign _5593_ = _5742_ ^ _5750_ /*15285*/;
assign _5748_ = _5749_ | _5751_ /*15282*/;
assign _5753_ = ~Q[19] /*15281*/;
assign _5752_ = _5753_ & D[25] /*15280*/;
assign _5755_ = _5370_ & _5752_ /*15275*/;
assign _5756_ = _5370_ ^ _5752_ /*15278*/;
assign _5757_ = _5748_ & _5756_ /*15276*/;
assign _5594_ = _5748_ ^ _5756_ /*15277*/;
assign _5754_ = _5755_ | _5757_ /*15274*/;
assign _5759_ = ~Q[19] /*15273*/;
assign _5758_ = _5759_ & D[26] /*15272*/;
assign _5761_ = _5371_ & _5758_ /*15267*/;
assign _5762_ = _5371_ ^ _5758_ /*15270*/;
assign _5763_ = _5754_ & _5762_ /*15268*/;
assign _5595_ = _5754_ ^ _5762_ /*15269*/;
assign _5760_ = _5761_ | _5763_ /*15266*/;
assign _5765_ = ~Q[19] /*15265*/;
assign _5764_ = _5765_ & D[27] /*15264*/;
assign _5767_ = _5372_ & _5764_ /*15259*/;
assign _5768_ = _5372_ ^ _5764_ /*15262*/;
assign _5769_ = _5760_ & _5768_ /*15260*/;
assign _5596_ = _5760_ ^ _5768_ /*15261*/;
assign _5766_ = _5767_ | _5769_ /*15258*/;
assign _5771_ = ~Q[19] /*15257*/;
assign _5770_ = _5771_ & D[28] /*15256*/;
assign _5773_ = _5373_ & _5770_ /*15251*/;
assign _5774_ = _5373_ ^ _5770_ /*15254*/;
assign _5775_ = _5766_ & _5774_ /*15252*/;
assign _5597_ = _5766_ ^ _5774_ /*15253*/;
assign _5772_ = _5773_ | _5775_ /*15250*/;
assign _5777_ = ~Q[19] /*15249*/;
assign _5776_ = _5777_ & D[29] /*15248*/;
assign _5779_ = _5374_ & _5776_ /*15243*/;
assign _5780_ = _5374_ ^ _5776_ /*15246*/;
assign _5781_ = _5772_ & _5780_ /*15244*/;
assign _5598_ = _5772_ ^ _5780_ /*15245*/;
assign _5778_ = _5779_ | _5781_ /*15242*/;
assign _5783_ = ~Q[19] /*15241*/;
assign _5782_ = _5783_ & D[30] /*15240*/;
assign _5785_ = _5375_ & _5782_ /*15235*/;
assign _5786_ = _5375_ ^ _5782_ /*15238*/;
assign _5787_ = _5778_ & _5786_ /*15236*/;
assign _5599_ = _5778_ ^ _5786_ /*15237*/;
assign _5784_ = _5785_ | _5787_ /*15234*/;
assign _5789_ = ~Q[19] /*15233*/;
assign _5788_ = _5789_ & zeroWire /*15232*/;
assign _5790_ = _5376_ ^ _5788_ /*15230*/;
assign _5600_ = _5790_ ^ _5784_ /*15229*/;
assign _5829_ = ~D[0] /*15103*/;
assign _5826_ = R_0[18] & _5829_ /*15099*/;
assign _5827_ = R_0[18] ^ _5829_ /*15102*/;
assign _5828_ = oneWire & _5827_ /*15100*/;
assign _5793_ = oneWire ^ _5827_ /*15101*/;
assign _5825_ = _5826_ | _5828_ /*15098*/;
assign _5834_ = ~D[1] /*15097*/;
assign _5831_ = _5569_ & _5834_ /*15093*/;
assign _5832_ = _5569_ ^ _5834_ /*15096*/;
assign _5833_ = _5825_ & _5832_ /*15094*/;
assign _5794_ = _5825_ ^ _5832_ /*15095*/;
assign _5830_ = _5831_ | _5833_ /*15092*/;
assign _5839_ = ~D[2] /*15091*/;
assign _5836_ = _5570_ & _5839_ /*15087*/;
assign _5837_ = _5570_ ^ _5839_ /*15090*/;
assign _5838_ = _5830_ & _5837_ /*15088*/;
assign _5795_ = _5830_ ^ _5837_ /*15089*/;
assign _5835_ = _5836_ | _5838_ /*15086*/;
assign _5844_ = ~D[3] /*15085*/;
assign _5841_ = _5571_ & _5844_ /*15081*/;
assign _5842_ = _5571_ ^ _5844_ /*15084*/;
assign _5843_ = _5835_ & _5842_ /*15082*/;
assign _5796_ = _5835_ ^ _5842_ /*15083*/;
assign _5840_ = _5841_ | _5843_ /*15080*/;
assign _5849_ = ~D[4] /*15079*/;
assign _5846_ = _5572_ & _5849_ /*15075*/;
assign _5847_ = _5572_ ^ _5849_ /*15078*/;
assign _5848_ = _5840_ & _5847_ /*15076*/;
assign _5797_ = _5840_ ^ _5847_ /*15077*/;
assign _5845_ = _5846_ | _5848_ /*15074*/;
assign _5854_ = ~D[5] /*15073*/;
assign _5851_ = _5573_ & _5854_ /*15069*/;
assign _5852_ = _5573_ ^ _5854_ /*15072*/;
assign _5853_ = _5845_ & _5852_ /*15070*/;
assign _5798_ = _5845_ ^ _5852_ /*15071*/;
assign _5850_ = _5851_ | _5853_ /*15068*/;
assign _5859_ = ~D[6] /*15067*/;
assign _5856_ = _5574_ & _5859_ /*15063*/;
assign _5857_ = _5574_ ^ _5859_ /*15066*/;
assign _5858_ = _5850_ & _5857_ /*15064*/;
assign _5799_ = _5850_ ^ _5857_ /*15065*/;
assign _5855_ = _5856_ | _5858_ /*15062*/;
assign _5864_ = ~D[7] /*15061*/;
assign _5861_ = _5575_ & _5864_ /*15057*/;
assign _5862_ = _5575_ ^ _5864_ /*15060*/;
assign _5863_ = _5855_ & _5862_ /*15058*/;
assign _5800_ = _5855_ ^ _5862_ /*15059*/;
assign _5860_ = _5861_ | _5863_ /*15056*/;
assign _5869_ = ~D[8] /*15055*/;
assign _5866_ = _5576_ & _5869_ /*15051*/;
assign _5867_ = _5576_ ^ _5869_ /*15054*/;
assign _5868_ = _5860_ & _5867_ /*15052*/;
assign _5801_ = _5860_ ^ _5867_ /*15053*/;
assign _5865_ = _5866_ | _5868_ /*15050*/;
assign _5874_ = ~D[9] /*15049*/;
assign _5871_ = _5577_ & _5874_ /*15045*/;
assign _5872_ = _5577_ ^ _5874_ /*15048*/;
assign _5873_ = _5865_ & _5872_ /*15046*/;
assign _5802_ = _5865_ ^ _5872_ /*15047*/;
assign _5870_ = _5871_ | _5873_ /*15044*/;
assign _5879_ = ~D[10] /*15043*/;
assign _5876_ = _5578_ & _5879_ /*15039*/;
assign _5877_ = _5578_ ^ _5879_ /*15042*/;
assign _5878_ = _5870_ & _5877_ /*15040*/;
assign _5803_ = _5870_ ^ _5877_ /*15041*/;
assign _5875_ = _5876_ | _5878_ /*15038*/;
assign _5884_ = ~D[11] /*15037*/;
assign _5881_ = _5579_ & _5884_ /*15033*/;
assign _5882_ = _5579_ ^ _5884_ /*15036*/;
assign _5883_ = _5875_ & _5882_ /*15034*/;
assign _5804_ = _5875_ ^ _5882_ /*15035*/;
assign _5880_ = _5881_ | _5883_ /*15032*/;
assign _5889_ = ~D[12] /*15031*/;
assign _5886_ = _5580_ & _5889_ /*15027*/;
assign _5887_ = _5580_ ^ _5889_ /*15030*/;
assign _5888_ = _5880_ & _5887_ /*15028*/;
assign _5805_ = _5880_ ^ _5887_ /*15029*/;
assign _5885_ = _5886_ | _5888_ /*15026*/;
assign _5894_ = ~D[13] /*15025*/;
assign _5891_ = _5581_ & _5894_ /*15021*/;
assign _5892_ = _5581_ ^ _5894_ /*15024*/;
assign _5893_ = _5885_ & _5892_ /*15022*/;
assign _5806_ = _5885_ ^ _5892_ /*15023*/;
assign _5890_ = _5891_ | _5893_ /*15020*/;
assign _5899_ = ~D[14] /*15019*/;
assign _5896_ = _5582_ & _5899_ /*15015*/;
assign _5897_ = _5582_ ^ _5899_ /*15018*/;
assign _5898_ = _5890_ & _5897_ /*15016*/;
assign _5807_ = _5890_ ^ _5897_ /*15017*/;
assign _5895_ = _5896_ | _5898_ /*15014*/;
assign _5904_ = ~D[15] /*15013*/;
assign _5901_ = _5583_ & _5904_ /*15009*/;
assign _5902_ = _5583_ ^ _5904_ /*15012*/;
assign _5903_ = _5895_ & _5902_ /*15010*/;
assign _5808_ = _5895_ ^ _5902_ /*15011*/;
assign _5900_ = _5901_ | _5903_ /*15008*/;
assign _5909_ = ~D[16] /*15007*/;
assign _5906_ = _5584_ & _5909_ /*15003*/;
assign _5907_ = _5584_ ^ _5909_ /*15006*/;
assign _5908_ = _5900_ & _5907_ /*15004*/;
assign _5809_ = _5900_ ^ _5907_ /*15005*/;
assign _5905_ = _5906_ | _5908_ /*15002*/;
assign _5914_ = ~D[17] /*15001*/;
assign _5911_ = _5585_ & _5914_ /*14997*/;
assign _5912_ = _5585_ ^ _5914_ /*15000*/;
assign _5913_ = _5905_ & _5912_ /*14998*/;
assign _5810_ = _5905_ ^ _5912_ /*14999*/;
assign _5910_ = _5911_ | _5913_ /*14996*/;
assign _5919_ = ~D[18] /*14995*/;
assign _5916_ = _5586_ & _5919_ /*14991*/;
assign _5917_ = _5586_ ^ _5919_ /*14994*/;
assign _5918_ = _5910_ & _5917_ /*14992*/;
assign _5811_ = _5910_ ^ _5917_ /*14993*/;
assign _5915_ = _5916_ | _5918_ /*14990*/;
assign _5924_ = ~D[19] /*14989*/;
assign _5921_ = _5587_ & _5924_ /*14985*/;
assign _5922_ = _5587_ ^ _5924_ /*14988*/;
assign _5923_ = _5915_ & _5922_ /*14986*/;
assign _5812_ = _5915_ ^ _5922_ /*14987*/;
assign _5920_ = _5921_ | _5923_ /*14984*/;
assign _5929_ = ~D[20] /*14983*/;
assign _5926_ = _5588_ & _5929_ /*14979*/;
assign _5927_ = _5588_ ^ _5929_ /*14982*/;
assign _5928_ = _5920_ & _5927_ /*14980*/;
assign _5813_ = _5920_ ^ _5927_ /*14981*/;
assign _5925_ = _5926_ | _5928_ /*14978*/;
assign _5934_ = ~D[21] /*14977*/;
assign _5931_ = _5589_ & _5934_ /*14973*/;
assign _5932_ = _5589_ ^ _5934_ /*14976*/;
assign _5933_ = _5925_ & _5932_ /*14974*/;
assign _5814_ = _5925_ ^ _5932_ /*14975*/;
assign _5930_ = _5931_ | _5933_ /*14972*/;
assign _5939_ = ~D[22] /*14971*/;
assign _5936_ = _5590_ & _5939_ /*14967*/;
assign _5937_ = _5590_ ^ _5939_ /*14970*/;
assign _5938_ = _5930_ & _5937_ /*14968*/;
assign _5815_ = _5930_ ^ _5937_ /*14969*/;
assign _5935_ = _5936_ | _5938_ /*14966*/;
assign _5944_ = ~D[23] /*14965*/;
assign _5941_ = _5591_ & _5944_ /*14961*/;
assign _5942_ = _5591_ ^ _5944_ /*14964*/;
assign _5943_ = _5935_ & _5942_ /*14962*/;
assign _5816_ = _5935_ ^ _5942_ /*14963*/;
assign _5940_ = _5941_ | _5943_ /*14960*/;
assign _5949_ = ~D[24] /*14959*/;
assign _5946_ = _5592_ & _5949_ /*14955*/;
assign _5947_ = _5592_ ^ _5949_ /*14958*/;
assign _5948_ = _5940_ & _5947_ /*14956*/;
assign _5817_ = _5940_ ^ _5947_ /*14957*/;
assign _5945_ = _5946_ | _5948_ /*14954*/;
assign _5954_ = ~D[25] /*14953*/;
assign _5951_ = _5593_ & _5954_ /*14949*/;
assign _5952_ = _5593_ ^ _5954_ /*14952*/;
assign _5953_ = _5945_ & _5952_ /*14950*/;
assign _5818_ = _5945_ ^ _5952_ /*14951*/;
assign _5950_ = _5951_ | _5953_ /*14948*/;
assign _5959_ = ~D[26] /*14947*/;
assign _5956_ = _5594_ & _5959_ /*14943*/;
assign _5957_ = _5594_ ^ _5959_ /*14946*/;
assign _5958_ = _5950_ & _5957_ /*14944*/;
assign _5819_ = _5950_ ^ _5957_ /*14945*/;
assign _5955_ = _5956_ | _5958_ /*14942*/;
assign _5964_ = ~D[27] /*14941*/;
assign _5961_ = _5595_ & _5964_ /*14937*/;
assign _5962_ = _5595_ ^ _5964_ /*14940*/;
assign _5963_ = _5955_ & _5962_ /*14938*/;
assign _5820_ = _5955_ ^ _5962_ /*14939*/;
assign _5960_ = _5961_ | _5963_ /*14936*/;
assign _5969_ = ~D[28] /*14935*/;
assign _5966_ = _5596_ & _5969_ /*14931*/;
assign _5967_ = _5596_ ^ _5969_ /*14934*/;
assign _5968_ = _5960_ & _5967_ /*14932*/;
assign _5821_ = _5960_ ^ _5967_ /*14933*/;
assign _5965_ = _5966_ | _5968_ /*14930*/;
assign _5974_ = ~D[29] /*14929*/;
assign _5971_ = _5597_ & _5974_ /*14925*/;
assign _5972_ = _5597_ ^ _5974_ /*14928*/;
assign _5973_ = _5965_ & _5972_ /*14926*/;
assign _5822_ = _5965_ ^ _5972_ /*14927*/;
assign _5970_ = _5971_ | _5973_ /*14924*/;
assign _5979_ = ~D[30] /*14923*/;
assign _5976_ = _5598_ & _5979_ /*14919*/;
assign _5977_ = _5598_ ^ _5979_ /*14922*/;
assign _5978_ = _5970_ & _5977_ /*14920*/;
assign _5823_ = _5970_ ^ _5977_ /*14921*/;
assign _5975_ = _5976_ | _5978_ /*14918*/;
assign _5980_ = _5599_ & oneWire /*14913*/;
assign _5981_ = _5599_ ^ oneWire /*14916*/;
assign _5982_ = _5975_ & _5981_ /*14914*/;
assign _5824_ = _5975_ ^ _5981_ /*14915*/;
assign Q[18] = _5980_ | _5982_ /*14912*/;
assign _6051_ = ~Q[18] /*14719*/;
assign _6050_ = _6051_ & D[0] /*14718*/;
assign _6053_ = _5793_ & _6050_ /*14713*/;
assign _6054_ = _5793_ ^ _6050_ /*14716*/;
assign _6055_ = zeroWire & _6054_ /*14714*/;
assign _6017_ = zeroWire ^ _6054_ /*14715*/;
assign _6052_ = _6053_ | _6055_ /*14712*/;
assign _6057_ = ~Q[18] /*14711*/;
assign _6056_ = _6057_ & D[1] /*14710*/;
assign _6059_ = _5794_ & _6056_ /*14705*/;
assign _6060_ = _5794_ ^ _6056_ /*14708*/;
assign _6061_ = _6052_ & _6060_ /*14706*/;
assign _6018_ = _6052_ ^ _6060_ /*14707*/;
assign _6058_ = _6059_ | _6061_ /*14704*/;
assign _6063_ = ~Q[18] /*14703*/;
assign _6062_ = _6063_ & D[2] /*14702*/;
assign _6065_ = _5795_ & _6062_ /*14697*/;
assign _6066_ = _5795_ ^ _6062_ /*14700*/;
assign _6067_ = _6058_ & _6066_ /*14698*/;
assign _6019_ = _6058_ ^ _6066_ /*14699*/;
assign _6064_ = _6065_ | _6067_ /*14696*/;
assign _6069_ = ~Q[18] /*14695*/;
assign _6068_ = _6069_ & D[3] /*14694*/;
assign _6071_ = _5796_ & _6068_ /*14689*/;
assign _6072_ = _5796_ ^ _6068_ /*14692*/;
assign _6073_ = _6064_ & _6072_ /*14690*/;
assign _6020_ = _6064_ ^ _6072_ /*14691*/;
assign _6070_ = _6071_ | _6073_ /*14688*/;
assign _6075_ = ~Q[18] /*14687*/;
assign _6074_ = _6075_ & D[4] /*14686*/;
assign _6077_ = _5797_ & _6074_ /*14681*/;
assign _6078_ = _5797_ ^ _6074_ /*14684*/;
assign _6079_ = _6070_ & _6078_ /*14682*/;
assign _6021_ = _6070_ ^ _6078_ /*14683*/;
assign _6076_ = _6077_ | _6079_ /*14680*/;
assign _6081_ = ~Q[18] /*14679*/;
assign _6080_ = _6081_ & D[5] /*14678*/;
assign _6083_ = _5798_ & _6080_ /*14673*/;
assign _6084_ = _5798_ ^ _6080_ /*14676*/;
assign _6085_ = _6076_ & _6084_ /*14674*/;
assign _6022_ = _6076_ ^ _6084_ /*14675*/;
assign _6082_ = _6083_ | _6085_ /*14672*/;
assign _6087_ = ~Q[18] /*14671*/;
assign _6086_ = _6087_ & D[6] /*14670*/;
assign _6089_ = _5799_ & _6086_ /*14665*/;
assign _6090_ = _5799_ ^ _6086_ /*14668*/;
assign _6091_ = _6082_ & _6090_ /*14666*/;
assign _6023_ = _6082_ ^ _6090_ /*14667*/;
assign _6088_ = _6089_ | _6091_ /*14664*/;
assign _6093_ = ~Q[18] /*14663*/;
assign _6092_ = _6093_ & D[7] /*14662*/;
assign _6095_ = _5800_ & _6092_ /*14657*/;
assign _6096_ = _5800_ ^ _6092_ /*14660*/;
assign _6097_ = _6088_ & _6096_ /*14658*/;
assign _6024_ = _6088_ ^ _6096_ /*14659*/;
assign _6094_ = _6095_ | _6097_ /*14656*/;
assign _6099_ = ~Q[18] /*14655*/;
assign _6098_ = _6099_ & D[8] /*14654*/;
assign _6101_ = _5801_ & _6098_ /*14649*/;
assign _6102_ = _5801_ ^ _6098_ /*14652*/;
assign _6103_ = _6094_ & _6102_ /*14650*/;
assign _6025_ = _6094_ ^ _6102_ /*14651*/;
assign _6100_ = _6101_ | _6103_ /*14648*/;
assign _6105_ = ~Q[18] /*14647*/;
assign _6104_ = _6105_ & D[9] /*14646*/;
assign _6107_ = _5802_ & _6104_ /*14641*/;
assign _6108_ = _5802_ ^ _6104_ /*14644*/;
assign _6109_ = _6100_ & _6108_ /*14642*/;
assign _6026_ = _6100_ ^ _6108_ /*14643*/;
assign _6106_ = _6107_ | _6109_ /*14640*/;
assign _6111_ = ~Q[18] /*14639*/;
assign _6110_ = _6111_ & D[10] /*14638*/;
assign _6113_ = _5803_ & _6110_ /*14633*/;
assign _6114_ = _5803_ ^ _6110_ /*14636*/;
assign _6115_ = _6106_ & _6114_ /*14634*/;
assign _6027_ = _6106_ ^ _6114_ /*14635*/;
assign _6112_ = _6113_ | _6115_ /*14632*/;
assign _6117_ = ~Q[18] /*14631*/;
assign _6116_ = _6117_ & D[11] /*14630*/;
assign _6119_ = _5804_ & _6116_ /*14625*/;
assign _6120_ = _5804_ ^ _6116_ /*14628*/;
assign _6121_ = _6112_ & _6120_ /*14626*/;
assign _6028_ = _6112_ ^ _6120_ /*14627*/;
assign _6118_ = _6119_ | _6121_ /*14624*/;
assign _6123_ = ~Q[18] /*14623*/;
assign _6122_ = _6123_ & D[12] /*14622*/;
assign _6125_ = _5805_ & _6122_ /*14617*/;
assign _6126_ = _5805_ ^ _6122_ /*14620*/;
assign _6127_ = _6118_ & _6126_ /*14618*/;
assign _6029_ = _6118_ ^ _6126_ /*14619*/;
assign _6124_ = _6125_ | _6127_ /*14616*/;
assign _6129_ = ~Q[18] /*14615*/;
assign _6128_ = _6129_ & D[13] /*14614*/;
assign _6131_ = _5806_ & _6128_ /*14609*/;
assign _6132_ = _5806_ ^ _6128_ /*14612*/;
assign _6133_ = _6124_ & _6132_ /*14610*/;
assign _6030_ = _6124_ ^ _6132_ /*14611*/;
assign _6130_ = _6131_ | _6133_ /*14608*/;
assign _6135_ = ~Q[18] /*14607*/;
assign _6134_ = _6135_ & D[14] /*14606*/;
assign _6137_ = _5807_ & _6134_ /*14601*/;
assign _6138_ = _5807_ ^ _6134_ /*14604*/;
assign _6139_ = _6130_ & _6138_ /*14602*/;
assign _6031_ = _6130_ ^ _6138_ /*14603*/;
assign _6136_ = _6137_ | _6139_ /*14600*/;
assign _6141_ = ~Q[18] /*14599*/;
assign _6140_ = _6141_ & D[15] /*14598*/;
assign _6143_ = _5808_ & _6140_ /*14593*/;
assign _6144_ = _5808_ ^ _6140_ /*14596*/;
assign _6145_ = _6136_ & _6144_ /*14594*/;
assign _6032_ = _6136_ ^ _6144_ /*14595*/;
assign _6142_ = _6143_ | _6145_ /*14592*/;
assign _6147_ = ~Q[18] /*14591*/;
assign _6146_ = _6147_ & D[16] /*14590*/;
assign _6149_ = _5809_ & _6146_ /*14585*/;
assign _6150_ = _5809_ ^ _6146_ /*14588*/;
assign _6151_ = _6142_ & _6150_ /*14586*/;
assign _6033_ = _6142_ ^ _6150_ /*14587*/;
assign _6148_ = _6149_ | _6151_ /*14584*/;
assign _6153_ = ~Q[18] /*14583*/;
assign _6152_ = _6153_ & D[17] /*14582*/;
assign _6155_ = _5810_ & _6152_ /*14577*/;
assign _6156_ = _5810_ ^ _6152_ /*14580*/;
assign _6157_ = _6148_ & _6156_ /*14578*/;
assign _6034_ = _6148_ ^ _6156_ /*14579*/;
assign _6154_ = _6155_ | _6157_ /*14576*/;
assign _6159_ = ~Q[18] /*14575*/;
assign _6158_ = _6159_ & D[18] /*14574*/;
assign _6161_ = _5811_ & _6158_ /*14569*/;
assign _6162_ = _5811_ ^ _6158_ /*14572*/;
assign _6163_ = _6154_ & _6162_ /*14570*/;
assign _6035_ = _6154_ ^ _6162_ /*14571*/;
assign _6160_ = _6161_ | _6163_ /*14568*/;
assign _6165_ = ~Q[18] /*14567*/;
assign _6164_ = _6165_ & D[19] /*14566*/;
assign _6167_ = _5812_ & _6164_ /*14561*/;
assign _6168_ = _5812_ ^ _6164_ /*14564*/;
assign _6169_ = _6160_ & _6168_ /*14562*/;
assign _6036_ = _6160_ ^ _6168_ /*14563*/;
assign _6166_ = _6167_ | _6169_ /*14560*/;
assign _6171_ = ~Q[18] /*14559*/;
assign _6170_ = _6171_ & D[20] /*14558*/;
assign _6173_ = _5813_ & _6170_ /*14553*/;
assign _6174_ = _5813_ ^ _6170_ /*14556*/;
assign _6175_ = _6166_ & _6174_ /*14554*/;
assign _6037_ = _6166_ ^ _6174_ /*14555*/;
assign _6172_ = _6173_ | _6175_ /*14552*/;
assign _6177_ = ~Q[18] /*14551*/;
assign _6176_ = _6177_ & D[21] /*14550*/;
assign _6179_ = _5814_ & _6176_ /*14545*/;
assign _6180_ = _5814_ ^ _6176_ /*14548*/;
assign _6181_ = _6172_ & _6180_ /*14546*/;
assign _6038_ = _6172_ ^ _6180_ /*14547*/;
assign _6178_ = _6179_ | _6181_ /*14544*/;
assign _6183_ = ~Q[18] /*14543*/;
assign _6182_ = _6183_ & D[22] /*14542*/;
assign _6185_ = _5815_ & _6182_ /*14537*/;
assign _6186_ = _5815_ ^ _6182_ /*14540*/;
assign _6187_ = _6178_ & _6186_ /*14538*/;
assign _6039_ = _6178_ ^ _6186_ /*14539*/;
assign _6184_ = _6185_ | _6187_ /*14536*/;
assign _6189_ = ~Q[18] /*14535*/;
assign _6188_ = _6189_ & D[23] /*14534*/;
assign _6191_ = _5816_ & _6188_ /*14529*/;
assign _6192_ = _5816_ ^ _6188_ /*14532*/;
assign _6193_ = _6184_ & _6192_ /*14530*/;
assign _6040_ = _6184_ ^ _6192_ /*14531*/;
assign _6190_ = _6191_ | _6193_ /*14528*/;
assign _6195_ = ~Q[18] /*14527*/;
assign _6194_ = _6195_ & D[24] /*14526*/;
assign _6197_ = _5817_ & _6194_ /*14521*/;
assign _6198_ = _5817_ ^ _6194_ /*14524*/;
assign _6199_ = _6190_ & _6198_ /*14522*/;
assign _6041_ = _6190_ ^ _6198_ /*14523*/;
assign _6196_ = _6197_ | _6199_ /*14520*/;
assign _6201_ = ~Q[18] /*14519*/;
assign _6200_ = _6201_ & D[25] /*14518*/;
assign _6203_ = _5818_ & _6200_ /*14513*/;
assign _6204_ = _5818_ ^ _6200_ /*14516*/;
assign _6205_ = _6196_ & _6204_ /*14514*/;
assign _6042_ = _6196_ ^ _6204_ /*14515*/;
assign _6202_ = _6203_ | _6205_ /*14512*/;
assign _6207_ = ~Q[18] /*14511*/;
assign _6206_ = _6207_ & D[26] /*14510*/;
assign _6209_ = _5819_ & _6206_ /*14505*/;
assign _6210_ = _5819_ ^ _6206_ /*14508*/;
assign _6211_ = _6202_ & _6210_ /*14506*/;
assign _6043_ = _6202_ ^ _6210_ /*14507*/;
assign _6208_ = _6209_ | _6211_ /*14504*/;
assign _6213_ = ~Q[18] /*14503*/;
assign _6212_ = _6213_ & D[27] /*14502*/;
assign _6215_ = _5820_ & _6212_ /*14497*/;
assign _6216_ = _5820_ ^ _6212_ /*14500*/;
assign _6217_ = _6208_ & _6216_ /*14498*/;
assign _6044_ = _6208_ ^ _6216_ /*14499*/;
assign _6214_ = _6215_ | _6217_ /*14496*/;
assign _6219_ = ~Q[18] /*14495*/;
assign _6218_ = _6219_ & D[28] /*14494*/;
assign _6221_ = _5821_ & _6218_ /*14489*/;
assign _6222_ = _5821_ ^ _6218_ /*14492*/;
assign _6223_ = _6214_ & _6222_ /*14490*/;
assign _6045_ = _6214_ ^ _6222_ /*14491*/;
assign _6220_ = _6221_ | _6223_ /*14488*/;
assign _6225_ = ~Q[18] /*14487*/;
assign _6224_ = _6225_ & D[29] /*14486*/;
assign _6227_ = _5822_ & _6224_ /*14481*/;
assign _6228_ = _5822_ ^ _6224_ /*14484*/;
assign _6229_ = _6220_ & _6228_ /*14482*/;
assign _6046_ = _6220_ ^ _6228_ /*14483*/;
assign _6226_ = _6227_ | _6229_ /*14480*/;
assign _6231_ = ~Q[18] /*14479*/;
assign _6230_ = _6231_ & D[30] /*14478*/;
assign _6233_ = _5823_ & _6230_ /*14473*/;
assign _6234_ = _5823_ ^ _6230_ /*14476*/;
assign _6235_ = _6226_ & _6234_ /*14474*/;
assign _6047_ = _6226_ ^ _6234_ /*14475*/;
assign _6232_ = _6233_ | _6235_ /*14472*/;
assign _6237_ = ~Q[18] /*14471*/;
assign _6236_ = _6237_ & zeroWire /*14470*/;
assign _6238_ = _5824_ ^ _6236_ /*14468*/;
assign _6048_ = _6238_ ^ _6232_ /*14467*/;
assign _6277_ = ~D[0] /*14341*/;
assign _6274_ = R_0[17] & _6277_ /*14337*/;
assign _6275_ = R_0[17] ^ _6277_ /*14340*/;
assign _6276_ = oneWire & _6275_ /*14338*/;
assign _6241_ = oneWire ^ _6275_ /*14339*/;
assign _6273_ = _6274_ | _6276_ /*14336*/;
assign _6282_ = ~D[1] /*14335*/;
assign _6279_ = _6017_ & _6282_ /*14331*/;
assign _6280_ = _6017_ ^ _6282_ /*14334*/;
assign _6281_ = _6273_ & _6280_ /*14332*/;
assign _6242_ = _6273_ ^ _6280_ /*14333*/;
assign _6278_ = _6279_ | _6281_ /*14330*/;
assign _6287_ = ~D[2] /*14329*/;
assign _6284_ = _6018_ & _6287_ /*14325*/;
assign _6285_ = _6018_ ^ _6287_ /*14328*/;
assign _6286_ = _6278_ & _6285_ /*14326*/;
assign _6243_ = _6278_ ^ _6285_ /*14327*/;
assign _6283_ = _6284_ | _6286_ /*14324*/;
assign _6292_ = ~D[3] /*14323*/;
assign _6289_ = _6019_ & _6292_ /*14319*/;
assign _6290_ = _6019_ ^ _6292_ /*14322*/;
assign _6291_ = _6283_ & _6290_ /*14320*/;
assign _6244_ = _6283_ ^ _6290_ /*14321*/;
assign _6288_ = _6289_ | _6291_ /*14318*/;
assign _6297_ = ~D[4] /*14317*/;
assign _6294_ = _6020_ & _6297_ /*14313*/;
assign _6295_ = _6020_ ^ _6297_ /*14316*/;
assign _6296_ = _6288_ & _6295_ /*14314*/;
assign _6245_ = _6288_ ^ _6295_ /*14315*/;
assign _6293_ = _6294_ | _6296_ /*14312*/;
assign _6302_ = ~D[5] /*14311*/;
assign _6299_ = _6021_ & _6302_ /*14307*/;
assign _6300_ = _6021_ ^ _6302_ /*14310*/;
assign _6301_ = _6293_ & _6300_ /*14308*/;
assign _6246_ = _6293_ ^ _6300_ /*14309*/;
assign _6298_ = _6299_ | _6301_ /*14306*/;
assign _6307_ = ~D[6] /*14305*/;
assign _6304_ = _6022_ & _6307_ /*14301*/;
assign _6305_ = _6022_ ^ _6307_ /*14304*/;
assign _6306_ = _6298_ & _6305_ /*14302*/;
assign _6247_ = _6298_ ^ _6305_ /*14303*/;
assign _6303_ = _6304_ | _6306_ /*14300*/;
assign _6312_ = ~D[7] /*14299*/;
assign _6309_ = _6023_ & _6312_ /*14295*/;
assign _6310_ = _6023_ ^ _6312_ /*14298*/;
assign _6311_ = _6303_ & _6310_ /*14296*/;
assign _6248_ = _6303_ ^ _6310_ /*14297*/;
assign _6308_ = _6309_ | _6311_ /*14294*/;
assign _6317_ = ~D[8] /*14293*/;
assign _6314_ = _6024_ & _6317_ /*14289*/;
assign _6315_ = _6024_ ^ _6317_ /*14292*/;
assign _6316_ = _6308_ & _6315_ /*14290*/;
assign _6249_ = _6308_ ^ _6315_ /*14291*/;
assign _6313_ = _6314_ | _6316_ /*14288*/;
assign _6322_ = ~D[9] /*14287*/;
assign _6319_ = _6025_ & _6322_ /*14283*/;
assign _6320_ = _6025_ ^ _6322_ /*14286*/;
assign _6321_ = _6313_ & _6320_ /*14284*/;
assign _6250_ = _6313_ ^ _6320_ /*14285*/;
assign _6318_ = _6319_ | _6321_ /*14282*/;
assign _6327_ = ~D[10] /*14281*/;
assign _6324_ = _6026_ & _6327_ /*14277*/;
assign _6325_ = _6026_ ^ _6327_ /*14280*/;
assign _6326_ = _6318_ & _6325_ /*14278*/;
assign _6251_ = _6318_ ^ _6325_ /*14279*/;
assign _6323_ = _6324_ | _6326_ /*14276*/;
assign _6332_ = ~D[11] /*14275*/;
assign _6329_ = _6027_ & _6332_ /*14271*/;
assign _6330_ = _6027_ ^ _6332_ /*14274*/;
assign _6331_ = _6323_ & _6330_ /*14272*/;
assign _6252_ = _6323_ ^ _6330_ /*14273*/;
assign _6328_ = _6329_ | _6331_ /*14270*/;
assign _6337_ = ~D[12] /*14269*/;
assign _6334_ = _6028_ & _6337_ /*14265*/;
assign _6335_ = _6028_ ^ _6337_ /*14268*/;
assign _6336_ = _6328_ & _6335_ /*14266*/;
assign _6253_ = _6328_ ^ _6335_ /*14267*/;
assign _6333_ = _6334_ | _6336_ /*14264*/;
assign _6342_ = ~D[13] /*14263*/;
assign _6339_ = _6029_ & _6342_ /*14259*/;
assign _6340_ = _6029_ ^ _6342_ /*14262*/;
assign _6341_ = _6333_ & _6340_ /*14260*/;
assign _6254_ = _6333_ ^ _6340_ /*14261*/;
assign _6338_ = _6339_ | _6341_ /*14258*/;
assign _6347_ = ~D[14] /*14257*/;
assign _6344_ = _6030_ & _6347_ /*14253*/;
assign _6345_ = _6030_ ^ _6347_ /*14256*/;
assign _6346_ = _6338_ & _6345_ /*14254*/;
assign _6255_ = _6338_ ^ _6345_ /*14255*/;
assign _6343_ = _6344_ | _6346_ /*14252*/;
assign _6352_ = ~D[15] /*14251*/;
assign _6349_ = _6031_ & _6352_ /*14247*/;
assign _6350_ = _6031_ ^ _6352_ /*14250*/;
assign _6351_ = _6343_ & _6350_ /*14248*/;
assign _6256_ = _6343_ ^ _6350_ /*14249*/;
assign _6348_ = _6349_ | _6351_ /*14246*/;
assign _6357_ = ~D[16] /*14245*/;
assign _6354_ = _6032_ & _6357_ /*14241*/;
assign _6355_ = _6032_ ^ _6357_ /*14244*/;
assign _6356_ = _6348_ & _6355_ /*14242*/;
assign _6257_ = _6348_ ^ _6355_ /*14243*/;
assign _6353_ = _6354_ | _6356_ /*14240*/;
assign _6362_ = ~D[17] /*14239*/;
assign _6359_ = _6033_ & _6362_ /*14235*/;
assign _6360_ = _6033_ ^ _6362_ /*14238*/;
assign _6361_ = _6353_ & _6360_ /*14236*/;
assign _6258_ = _6353_ ^ _6360_ /*14237*/;
assign _6358_ = _6359_ | _6361_ /*14234*/;
assign _6367_ = ~D[18] /*14233*/;
assign _6364_ = _6034_ & _6367_ /*14229*/;
assign _6365_ = _6034_ ^ _6367_ /*14232*/;
assign _6366_ = _6358_ & _6365_ /*14230*/;
assign _6259_ = _6358_ ^ _6365_ /*14231*/;
assign _6363_ = _6364_ | _6366_ /*14228*/;
assign _6372_ = ~D[19] /*14227*/;
assign _6369_ = _6035_ & _6372_ /*14223*/;
assign _6370_ = _6035_ ^ _6372_ /*14226*/;
assign _6371_ = _6363_ & _6370_ /*14224*/;
assign _6260_ = _6363_ ^ _6370_ /*14225*/;
assign _6368_ = _6369_ | _6371_ /*14222*/;
assign _6377_ = ~D[20] /*14221*/;
assign _6374_ = _6036_ & _6377_ /*14217*/;
assign _6375_ = _6036_ ^ _6377_ /*14220*/;
assign _6376_ = _6368_ & _6375_ /*14218*/;
assign _6261_ = _6368_ ^ _6375_ /*14219*/;
assign _6373_ = _6374_ | _6376_ /*14216*/;
assign _6382_ = ~D[21] /*14215*/;
assign _6379_ = _6037_ & _6382_ /*14211*/;
assign _6380_ = _6037_ ^ _6382_ /*14214*/;
assign _6381_ = _6373_ & _6380_ /*14212*/;
assign _6262_ = _6373_ ^ _6380_ /*14213*/;
assign _6378_ = _6379_ | _6381_ /*14210*/;
assign _6387_ = ~D[22] /*14209*/;
assign _6384_ = _6038_ & _6387_ /*14205*/;
assign _6385_ = _6038_ ^ _6387_ /*14208*/;
assign _6386_ = _6378_ & _6385_ /*14206*/;
assign _6263_ = _6378_ ^ _6385_ /*14207*/;
assign _6383_ = _6384_ | _6386_ /*14204*/;
assign _6392_ = ~D[23] /*14203*/;
assign _6389_ = _6039_ & _6392_ /*14199*/;
assign _6390_ = _6039_ ^ _6392_ /*14202*/;
assign _6391_ = _6383_ & _6390_ /*14200*/;
assign _6264_ = _6383_ ^ _6390_ /*14201*/;
assign _6388_ = _6389_ | _6391_ /*14198*/;
assign _6397_ = ~D[24] /*14197*/;
assign _6394_ = _6040_ & _6397_ /*14193*/;
assign _6395_ = _6040_ ^ _6397_ /*14196*/;
assign _6396_ = _6388_ & _6395_ /*14194*/;
assign _6265_ = _6388_ ^ _6395_ /*14195*/;
assign _6393_ = _6394_ | _6396_ /*14192*/;
assign _6402_ = ~D[25] /*14191*/;
assign _6399_ = _6041_ & _6402_ /*14187*/;
assign _6400_ = _6041_ ^ _6402_ /*14190*/;
assign _6401_ = _6393_ & _6400_ /*14188*/;
assign _6266_ = _6393_ ^ _6400_ /*14189*/;
assign _6398_ = _6399_ | _6401_ /*14186*/;
assign _6407_ = ~D[26] /*14185*/;
assign _6404_ = _6042_ & _6407_ /*14181*/;
assign _6405_ = _6042_ ^ _6407_ /*14184*/;
assign _6406_ = _6398_ & _6405_ /*14182*/;
assign _6267_ = _6398_ ^ _6405_ /*14183*/;
assign _6403_ = _6404_ | _6406_ /*14180*/;
assign _6412_ = ~D[27] /*14179*/;
assign _6409_ = _6043_ & _6412_ /*14175*/;
assign _6410_ = _6043_ ^ _6412_ /*14178*/;
assign _6411_ = _6403_ & _6410_ /*14176*/;
assign _6268_ = _6403_ ^ _6410_ /*14177*/;
assign _6408_ = _6409_ | _6411_ /*14174*/;
assign _6417_ = ~D[28] /*14173*/;
assign _6414_ = _6044_ & _6417_ /*14169*/;
assign _6415_ = _6044_ ^ _6417_ /*14172*/;
assign _6416_ = _6408_ & _6415_ /*14170*/;
assign _6269_ = _6408_ ^ _6415_ /*14171*/;
assign _6413_ = _6414_ | _6416_ /*14168*/;
assign _6422_ = ~D[29] /*14167*/;
assign _6419_ = _6045_ & _6422_ /*14163*/;
assign _6420_ = _6045_ ^ _6422_ /*14166*/;
assign _6421_ = _6413_ & _6420_ /*14164*/;
assign _6270_ = _6413_ ^ _6420_ /*14165*/;
assign _6418_ = _6419_ | _6421_ /*14162*/;
assign _6427_ = ~D[30] /*14161*/;
assign _6424_ = _6046_ & _6427_ /*14157*/;
assign _6425_ = _6046_ ^ _6427_ /*14160*/;
assign _6426_ = _6418_ & _6425_ /*14158*/;
assign _6271_ = _6418_ ^ _6425_ /*14159*/;
assign _6423_ = _6424_ | _6426_ /*14156*/;
assign _6428_ = _6047_ & oneWire /*14151*/;
assign _6429_ = _6047_ ^ oneWire /*14154*/;
assign _6430_ = _6423_ & _6429_ /*14152*/;
assign _6272_ = _6423_ ^ _6429_ /*14153*/;
assign Q[17] = _6428_ | _6430_ /*14150*/;
assign _6499_ = ~Q[17] /*13957*/;
assign _6498_ = _6499_ & D[0] /*13956*/;
assign _6501_ = _6241_ & _6498_ /*13951*/;
assign _6502_ = _6241_ ^ _6498_ /*13954*/;
assign _6503_ = zeroWire & _6502_ /*13952*/;
assign _6465_ = zeroWire ^ _6502_ /*13953*/;
assign _6500_ = _6501_ | _6503_ /*13950*/;
assign _6505_ = ~Q[17] /*13949*/;
assign _6504_ = _6505_ & D[1] /*13948*/;
assign _6507_ = _6242_ & _6504_ /*13943*/;
assign _6508_ = _6242_ ^ _6504_ /*13946*/;
assign _6509_ = _6500_ & _6508_ /*13944*/;
assign _6466_ = _6500_ ^ _6508_ /*13945*/;
assign _6506_ = _6507_ | _6509_ /*13942*/;
assign _6511_ = ~Q[17] /*13941*/;
assign _6510_ = _6511_ & D[2] /*13940*/;
assign _6513_ = _6243_ & _6510_ /*13935*/;
assign _6514_ = _6243_ ^ _6510_ /*13938*/;
assign _6515_ = _6506_ & _6514_ /*13936*/;
assign _6467_ = _6506_ ^ _6514_ /*13937*/;
assign _6512_ = _6513_ | _6515_ /*13934*/;
assign _6517_ = ~Q[17] /*13933*/;
assign _6516_ = _6517_ & D[3] /*13932*/;
assign _6519_ = _6244_ & _6516_ /*13927*/;
assign _6520_ = _6244_ ^ _6516_ /*13930*/;
assign _6521_ = _6512_ & _6520_ /*13928*/;
assign _6468_ = _6512_ ^ _6520_ /*13929*/;
assign _6518_ = _6519_ | _6521_ /*13926*/;
assign _6523_ = ~Q[17] /*13925*/;
assign _6522_ = _6523_ & D[4] /*13924*/;
assign _6525_ = _6245_ & _6522_ /*13919*/;
assign _6526_ = _6245_ ^ _6522_ /*13922*/;
assign _6527_ = _6518_ & _6526_ /*13920*/;
assign _6469_ = _6518_ ^ _6526_ /*13921*/;
assign _6524_ = _6525_ | _6527_ /*13918*/;
assign _6529_ = ~Q[17] /*13917*/;
assign _6528_ = _6529_ & D[5] /*13916*/;
assign _6531_ = _6246_ & _6528_ /*13911*/;
assign _6532_ = _6246_ ^ _6528_ /*13914*/;
assign _6533_ = _6524_ & _6532_ /*13912*/;
assign _6470_ = _6524_ ^ _6532_ /*13913*/;
assign _6530_ = _6531_ | _6533_ /*13910*/;
assign _6535_ = ~Q[17] /*13909*/;
assign _6534_ = _6535_ & D[6] /*13908*/;
assign _6537_ = _6247_ & _6534_ /*13903*/;
assign _6538_ = _6247_ ^ _6534_ /*13906*/;
assign _6539_ = _6530_ & _6538_ /*13904*/;
assign _6471_ = _6530_ ^ _6538_ /*13905*/;
assign _6536_ = _6537_ | _6539_ /*13902*/;
assign _6541_ = ~Q[17] /*13901*/;
assign _6540_ = _6541_ & D[7] /*13900*/;
assign _6543_ = _6248_ & _6540_ /*13895*/;
assign _6544_ = _6248_ ^ _6540_ /*13898*/;
assign _6545_ = _6536_ & _6544_ /*13896*/;
assign _6472_ = _6536_ ^ _6544_ /*13897*/;
assign _6542_ = _6543_ | _6545_ /*13894*/;
assign _6547_ = ~Q[17] /*13893*/;
assign _6546_ = _6547_ & D[8] /*13892*/;
assign _6549_ = _6249_ & _6546_ /*13887*/;
assign _6550_ = _6249_ ^ _6546_ /*13890*/;
assign _6551_ = _6542_ & _6550_ /*13888*/;
assign _6473_ = _6542_ ^ _6550_ /*13889*/;
assign _6548_ = _6549_ | _6551_ /*13886*/;
assign _6553_ = ~Q[17] /*13885*/;
assign _6552_ = _6553_ & D[9] /*13884*/;
assign _6555_ = _6250_ & _6552_ /*13879*/;
assign _6556_ = _6250_ ^ _6552_ /*13882*/;
assign _6557_ = _6548_ & _6556_ /*13880*/;
assign _6474_ = _6548_ ^ _6556_ /*13881*/;
assign _6554_ = _6555_ | _6557_ /*13878*/;
assign _6559_ = ~Q[17] /*13877*/;
assign _6558_ = _6559_ & D[10] /*13876*/;
assign _6561_ = _6251_ & _6558_ /*13871*/;
assign _6562_ = _6251_ ^ _6558_ /*13874*/;
assign _6563_ = _6554_ & _6562_ /*13872*/;
assign _6475_ = _6554_ ^ _6562_ /*13873*/;
assign _6560_ = _6561_ | _6563_ /*13870*/;
assign _6565_ = ~Q[17] /*13869*/;
assign _6564_ = _6565_ & D[11] /*13868*/;
assign _6567_ = _6252_ & _6564_ /*13863*/;
assign _6568_ = _6252_ ^ _6564_ /*13866*/;
assign _6569_ = _6560_ & _6568_ /*13864*/;
assign _6476_ = _6560_ ^ _6568_ /*13865*/;
assign _6566_ = _6567_ | _6569_ /*13862*/;
assign _6571_ = ~Q[17] /*13861*/;
assign _6570_ = _6571_ & D[12] /*13860*/;
assign _6573_ = _6253_ & _6570_ /*13855*/;
assign _6574_ = _6253_ ^ _6570_ /*13858*/;
assign _6575_ = _6566_ & _6574_ /*13856*/;
assign _6477_ = _6566_ ^ _6574_ /*13857*/;
assign _6572_ = _6573_ | _6575_ /*13854*/;
assign _6577_ = ~Q[17] /*13853*/;
assign _6576_ = _6577_ & D[13] /*13852*/;
assign _6579_ = _6254_ & _6576_ /*13847*/;
assign _6580_ = _6254_ ^ _6576_ /*13850*/;
assign _6581_ = _6572_ & _6580_ /*13848*/;
assign _6478_ = _6572_ ^ _6580_ /*13849*/;
assign _6578_ = _6579_ | _6581_ /*13846*/;
assign _6583_ = ~Q[17] /*13845*/;
assign _6582_ = _6583_ & D[14] /*13844*/;
assign _6585_ = _6255_ & _6582_ /*13839*/;
assign _6586_ = _6255_ ^ _6582_ /*13842*/;
assign _6587_ = _6578_ & _6586_ /*13840*/;
assign _6479_ = _6578_ ^ _6586_ /*13841*/;
assign _6584_ = _6585_ | _6587_ /*13838*/;
assign _6589_ = ~Q[17] /*13837*/;
assign _6588_ = _6589_ & D[15] /*13836*/;
assign _6591_ = _6256_ & _6588_ /*13831*/;
assign _6592_ = _6256_ ^ _6588_ /*13834*/;
assign _6593_ = _6584_ & _6592_ /*13832*/;
assign _6480_ = _6584_ ^ _6592_ /*13833*/;
assign _6590_ = _6591_ | _6593_ /*13830*/;
assign _6595_ = ~Q[17] /*13829*/;
assign _6594_ = _6595_ & D[16] /*13828*/;
assign _6597_ = _6257_ & _6594_ /*13823*/;
assign _6598_ = _6257_ ^ _6594_ /*13826*/;
assign _6599_ = _6590_ & _6598_ /*13824*/;
assign _6481_ = _6590_ ^ _6598_ /*13825*/;
assign _6596_ = _6597_ | _6599_ /*13822*/;
assign _6601_ = ~Q[17] /*13821*/;
assign _6600_ = _6601_ & D[17] /*13820*/;
assign _6603_ = _6258_ & _6600_ /*13815*/;
assign _6604_ = _6258_ ^ _6600_ /*13818*/;
assign _6605_ = _6596_ & _6604_ /*13816*/;
assign _6482_ = _6596_ ^ _6604_ /*13817*/;
assign _6602_ = _6603_ | _6605_ /*13814*/;
assign _6607_ = ~Q[17] /*13813*/;
assign _6606_ = _6607_ & D[18] /*13812*/;
assign _6609_ = _6259_ & _6606_ /*13807*/;
assign _6610_ = _6259_ ^ _6606_ /*13810*/;
assign _6611_ = _6602_ & _6610_ /*13808*/;
assign _6483_ = _6602_ ^ _6610_ /*13809*/;
assign _6608_ = _6609_ | _6611_ /*13806*/;
assign _6613_ = ~Q[17] /*13805*/;
assign _6612_ = _6613_ & D[19] /*13804*/;
assign _6615_ = _6260_ & _6612_ /*13799*/;
assign _6616_ = _6260_ ^ _6612_ /*13802*/;
assign _6617_ = _6608_ & _6616_ /*13800*/;
assign _6484_ = _6608_ ^ _6616_ /*13801*/;
assign _6614_ = _6615_ | _6617_ /*13798*/;
assign _6619_ = ~Q[17] /*13797*/;
assign _6618_ = _6619_ & D[20] /*13796*/;
assign _6621_ = _6261_ & _6618_ /*13791*/;
assign _6622_ = _6261_ ^ _6618_ /*13794*/;
assign _6623_ = _6614_ & _6622_ /*13792*/;
assign _6485_ = _6614_ ^ _6622_ /*13793*/;
assign _6620_ = _6621_ | _6623_ /*13790*/;
assign _6625_ = ~Q[17] /*13789*/;
assign _6624_ = _6625_ & D[21] /*13788*/;
assign _6627_ = _6262_ & _6624_ /*13783*/;
assign _6628_ = _6262_ ^ _6624_ /*13786*/;
assign _6629_ = _6620_ & _6628_ /*13784*/;
assign _6486_ = _6620_ ^ _6628_ /*13785*/;
assign _6626_ = _6627_ | _6629_ /*13782*/;
assign _6631_ = ~Q[17] /*13781*/;
assign _6630_ = _6631_ & D[22] /*13780*/;
assign _6633_ = _6263_ & _6630_ /*13775*/;
assign _6634_ = _6263_ ^ _6630_ /*13778*/;
assign _6635_ = _6626_ & _6634_ /*13776*/;
assign _6487_ = _6626_ ^ _6634_ /*13777*/;
assign _6632_ = _6633_ | _6635_ /*13774*/;
assign _6637_ = ~Q[17] /*13773*/;
assign _6636_ = _6637_ & D[23] /*13772*/;
assign _6639_ = _6264_ & _6636_ /*13767*/;
assign _6640_ = _6264_ ^ _6636_ /*13770*/;
assign _6641_ = _6632_ & _6640_ /*13768*/;
assign _6488_ = _6632_ ^ _6640_ /*13769*/;
assign _6638_ = _6639_ | _6641_ /*13766*/;
assign _6643_ = ~Q[17] /*13765*/;
assign _6642_ = _6643_ & D[24] /*13764*/;
assign _6645_ = _6265_ & _6642_ /*13759*/;
assign _6646_ = _6265_ ^ _6642_ /*13762*/;
assign _6647_ = _6638_ & _6646_ /*13760*/;
assign _6489_ = _6638_ ^ _6646_ /*13761*/;
assign _6644_ = _6645_ | _6647_ /*13758*/;
assign _6649_ = ~Q[17] /*13757*/;
assign _6648_ = _6649_ & D[25] /*13756*/;
assign _6651_ = _6266_ & _6648_ /*13751*/;
assign _6652_ = _6266_ ^ _6648_ /*13754*/;
assign _6653_ = _6644_ & _6652_ /*13752*/;
assign _6490_ = _6644_ ^ _6652_ /*13753*/;
assign _6650_ = _6651_ | _6653_ /*13750*/;
assign _6655_ = ~Q[17] /*13749*/;
assign _6654_ = _6655_ & D[26] /*13748*/;
assign _6657_ = _6267_ & _6654_ /*13743*/;
assign _6658_ = _6267_ ^ _6654_ /*13746*/;
assign _6659_ = _6650_ & _6658_ /*13744*/;
assign _6491_ = _6650_ ^ _6658_ /*13745*/;
assign _6656_ = _6657_ | _6659_ /*13742*/;
assign _6661_ = ~Q[17] /*13741*/;
assign _6660_ = _6661_ & D[27] /*13740*/;
assign _6663_ = _6268_ & _6660_ /*13735*/;
assign _6664_ = _6268_ ^ _6660_ /*13738*/;
assign _6665_ = _6656_ & _6664_ /*13736*/;
assign _6492_ = _6656_ ^ _6664_ /*13737*/;
assign _6662_ = _6663_ | _6665_ /*13734*/;
assign _6667_ = ~Q[17] /*13733*/;
assign _6666_ = _6667_ & D[28] /*13732*/;
assign _6669_ = _6269_ & _6666_ /*13727*/;
assign _6670_ = _6269_ ^ _6666_ /*13730*/;
assign _6671_ = _6662_ & _6670_ /*13728*/;
assign _6493_ = _6662_ ^ _6670_ /*13729*/;
assign _6668_ = _6669_ | _6671_ /*13726*/;
assign _6673_ = ~Q[17] /*13725*/;
assign _6672_ = _6673_ & D[29] /*13724*/;
assign _6675_ = _6270_ & _6672_ /*13719*/;
assign _6676_ = _6270_ ^ _6672_ /*13722*/;
assign _6677_ = _6668_ & _6676_ /*13720*/;
assign _6494_ = _6668_ ^ _6676_ /*13721*/;
assign _6674_ = _6675_ | _6677_ /*13718*/;
assign _6679_ = ~Q[17] /*13717*/;
assign _6678_ = _6679_ & D[30] /*13716*/;
assign _6681_ = _6271_ & _6678_ /*13711*/;
assign _6682_ = _6271_ ^ _6678_ /*13714*/;
assign _6683_ = _6674_ & _6682_ /*13712*/;
assign _6495_ = _6674_ ^ _6682_ /*13713*/;
assign _6680_ = _6681_ | _6683_ /*13710*/;
assign _6685_ = ~Q[17] /*13709*/;
assign _6684_ = _6685_ & zeroWire /*13708*/;
assign _6686_ = _6272_ ^ _6684_ /*13706*/;
assign _6496_ = _6686_ ^ _6680_ /*13705*/;
assign _6725_ = ~D[0] /*13579*/;
assign _6722_ = R_0[16] & _6725_ /*13575*/;
assign _6723_ = R_0[16] ^ _6725_ /*13578*/;
assign _6724_ = oneWire & _6723_ /*13576*/;
assign _6689_ = oneWire ^ _6723_ /*13577*/;
assign _6721_ = _6722_ | _6724_ /*13574*/;
assign _6730_ = ~D[1] /*13573*/;
assign _6727_ = _6465_ & _6730_ /*13569*/;
assign _6728_ = _6465_ ^ _6730_ /*13572*/;
assign _6729_ = _6721_ & _6728_ /*13570*/;
assign _6690_ = _6721_ ^ _6728_ /*13571*/;
assign _6726_ = _6727_ | _6729_ /*13568*/;
assign _6735_ = ~D[2] /*13567*/;
assign _6732_ = _6466_ & _6735_ /*13563*/;
assign _6733_ = _6466_ ^ _6735_ /*13566*/;
assign _6734_ = _6726_ & _6733_ /*13564*/;
assign _6691_ = _6726_ ^ _6733_ /*13565*/;
assign _6731_ = _6732_ | _6734_ /*13562*/;
assign _6740_ = ~D[3] /*13561*/;
assign _6737_ = _6467_ & _6740_ /*13557*/;
assign _6738_ = _6467_ ^ _6740_ /*13560*/;
assign _6739_ = _6731_ & _6738_ /*13558*/;
assign _6692_ = _6731_ ^ _6738_ /*13559*/;
assign _6736_ = _6737_ | _6739_ /*13556*/;
assign _6745_ = ~D[4] /*13555*/;
assign _6742_ = _6468_ & _6745_ /*13551*/;
assign _6743_ = _6468_ ^ _6745_ /*13554*/;
assign _6744_ = _6736_ & _6743_ /*13552*/;
assign _6693_ = _6736_ ^ _6743_ /*13553*/;
assign _6741_ = _6742_ | _6744_ /*13550*/;
assign _6750_ = ~D[5] /*13549*/;
assign _6747_ = _6469_ & _6750_ /*13545*/;
assign _6748_ = _6469_ ^ _6750_ /*13548*/;
assign _6749_ = _6741_ & _6748_ /*13546*/;
assign _6694_ = _6741_ ^ _6748_ /*13547*/;
assign _6746_ = _6747_ | _6749_ /*13544*/;
assign _6755_ = ~D[6] /*13543*/;
assign _6752_ = _6470_ & _6755_ /*13539*/;
assign _6753_ = _6470_ ^ _6755_ /*13542*/;
assign _6754_ = _6746_ & _6753_ /*13540*/;
assign _6695_ = _6746_ ^ _6753_ /*13541*/;
assign _6751_ = _6752_ | _6754_ /*13538*/;
assign _6760_ = ~D[7] /*13537*/;
assign _6757_ = _6471_ & _6760_ /*13533*/;
assign _6758_ = _6471_ ^ _6760_ /*13536*/;
assign _6759_ = _6751_ & _6758_ /*13534*/;
assign _6696_ = _6751_ ^ _6758_ /*13535*/;
assign _6756_ = _6757_ | _6759_ /*13532*/;
assign _6765_ = ~D[8] /*13531*/;
assign _6762_ = _6472_ & _6765_ /*13527*/;
assign _6763_ = _6472_ ^ _6765_ /*13530*/;
assign _6764_ = _6756_ & _6763_ /*13528*/;
assign _6697_ = _6756_ ^ _6763_ /*13529*/;
assign _6761_ = _6762_ | _6764_ /*13526*/;
assign _6770_ = ~D[9] /*13525*/;
assign _6767_ = _6473_ & _6770_ /*13521*/;
assign _6768_ = _6473_ ^ _6770_ /*13524*/;
assign _6769_ = _6761_ & _6768_ /*13522*/;
assign _6698_ = _6761_ ^ _6768_ /*13523*/;
assign _6766_ = _6767_ | _6769_ /*13520*/;
assign _6775_ = ~D[10] /*13519*/;
assign _6772_ = _6474_ & _6775_ /*13515*/;
assign _6773_ = _6474_ ^ _6775_ /*13518*/;
assign _6774_ = _6766_ & _6773_ /*13516*/;
assign _6699_ = _6766_ ^ _6773_ /*13517*/;
assign _6771_ = _6772_ | _6774_ /*13514*/;
assign _6780_ = ~D[11] /*13513*/;
assign _6777_ = _6475_ & _6780_ /*13509*/;
assign _6778_ = _6475_ ^ _6780_ /*13512*/;
assign _6779_ = _6771_ & _6778_ /*13510*/;
assign _6700_ = _6771_ ^ _6778_ /*13511*/;
assign _6776_ = _6777_ | _6779_ /*13508*/;
assign _6785_ = ~D[12] /*13507*/;
assign _6782_ = _6476_ & _6785_ /*13503*/;
assign _6783_ = _6476_ ^ _6785_ /*13506*/;
assign _6784_ = _6776_ & _6783_ /*13504*/;
assign _6701_ = _6776_ ^ _6783_ /*13505*/;
assign _6781_ = _6782_ | _6784_ /*13502*/;
assign _6790_ = ~D[13] /*13501*/;
assign _6787_ = _6477_ & _6790_ /*13497*/;
assign _6788_ = _6477_ ^ _6790_ /*13500*/;
assign _6789_ = _6781_ & _6788_ /*13498*/;
assign _6702_ = _6781_ ^ _6788_ /*13499*/;
assign _6786_ = _6787_ | _6789_ /*13496*/;
assign _6795_ = ~D[14] /*13495*/;
assign _6792_ = _6478_ & _6795_ /*13491*/;
assign _6793_ = _6478_ ^ _6795_ /*13494*/;
assign _6794_ = _6786_ & _6793_ /*13492*/;
assign _6703_ = _6786_ ^ _6793_ /*13493*/;
assign _6791_ = _6792_ | _6794_ /*13490*/;
assign _6800_ = ~D[15] /*13489*/;
assign _6797_ = _6479_ & _6800_ /*13485*/;
assign _6798_ = _6479_ ^ _6800_ /*13488*/;
assign _6799_ = _6791_ & _6798_ /*13486*/;
assign _6704_ = _6791_ ^ _6798_ /*13487*/;
assign _6796_ = _6797_ | _6799_ /*13484*/;
assign _6805_ = ~D[16] /*13483*/;
assign _6802_ = _6480_ & _6805_ /*13479*/;
assign _6803_ = _6480_ ^ _6805_ /*13482*/;
assign _6804_ = _6796_ & _6803_ /*13480*/;
assign _6705_ = _6796_ ^ _6803_ /*13481*/;
assign _6801_ = _6802_ | _6804_ /*13478*/;
assign _6810_ = ~D[17] /*13477*/;
assign _6807_ = _6481_ & _6810_ /*13473*/;
assign _6808_ = _6481_ ^ _6810_ /*13476*/;
assign _6809_ = _6801_ & _6808_ /*13474*/;
assign _6706_ = _6801_ ^ _6808_ /*13475*/;
assign _6806_ = _6807_ | _6809_ /*13472*/;
assign _6815_ = ~D[18] /*13471*/;
assign _6812_ = _6482_ & _6815_ /*13467*/;
assign _6813_ = _6482_ ^ _6815_ /*13470*/;
assign _6814_ = _6806_ & _6813_ /*13468*/;
assign _6707_ = _6806_ ^ _6813_ /*13469*/;
assign _6811_ = _6812_ | _6814_ /*13466*/;
assign _6820_ = ~D[19] /*13465*/;
assign _6817_ = _6483_ & _6820_ /*13461*/;
assign _6818_ = _6483_ ^ _6820_ /*13464*/;
assign _6819_ = _6811_ & _6818_ /*13462*/;
assign _6708_ = _6811_ ^ _6818_ /*13463*/;
assign _6816_ = _6817_ | _6819_ /*13460*/;
assign _6825_ = ~D[20] /*13459*/;
assign _6822_ = _6484_ & _6825_ /*13455*/;
assign _6823_ = _6484_ ^ _6825_ /*13458*/;
assign _6824_ = _6816_ & _6823_ /*13456*/;
assign _6709_ = _6816_ ^ _6823_ /*13457*/;
assign _6821_ = _6822_ | _6824_ /*13454*/;
assign _6830_ = ~D[21] /*13453*/;
assign _6827_ = _6485_ & _6830_ /*13449*/;
assign _6828_ = _6485_ ^ _6830_ /*13452*/;
assign _6829_ = _6821_ & _6828_ /*13450*/;
assign _6710_ = _6821_ ^ _6828_ /*13451*/;
assign _6826_ = _6827_ | _6829_ /*13448*/;
assign _6835_ = ~D[22] /*13447*/;
assign _6832_ = _6486_ & _6835_ /*13443*/;
assign _6833_ = _6486_ ^ _6835_ /*13446*/;
assign _6834_ = _6826_ & _6833_ /*13444*/;
assign _6711_ = _6826_ ^ _6833_ /*13445*/;
assign _6831_ = _6832_ | _6834_ /*13442*/;
assign _6840_ = ~D[23] /*13441*/;
assign _6837_ = _6487_ & _6840_ /*13437*/;
assign _6838_ = _6487_ ^ _6840_ /*13440*/;
assign _6839_ = _6831_ & _6838_ /*13438*/;
assign _6712_ = _6831_ ^ _6838_ /*13439*/;
assign _6836_ = _6837_ | _6839_ /*13436*/;
assign _6845_ = ~D[24] /*13435*/;
assign _6842_ = _6488_ & _6845_ /*13431*/;
assign _6843_ = _6488_ ^ _6845_ /*13434*/;
assign _6844_ = _6836_ & _6843_ /*13432*/;
assign _6713_ = _6836_ ^ _6843_ /*13433*/;
assign _6841_ = _6842_ | _6844_ /*13430*/;
assign _6850_ = ~D[25] /*13429*/;
assign _6847_ = _6489_ & _6850_ /*13425*/;
assign _6848_ = _6489_ ^ _6850_ /*13428*/;
assign _6849_ = _6841_ & _6848_ /*13426*/;
assign _6714_ = _6841_ ^ _6848_ /*13427*/;
assign _6846_ = _6847_ | _6849_ /*13424*/;
assign _6855_ = ~D[26] /*13423*/;
assign _6852_ = _6490_ & _6855_ /*13419*/;
assign _6853_ = _6490_ ^ _6855_ /*13422*/;
assign _6854_ = _6846_ & _6853_ /*13420*/;
assign _6715_ = _6846_ ^ _6853_ /*13421*/;
assign _6851_ = _6852_ | _6854_ /*13418*/;
assign _6860_ = ~D[27] /*13417*/;
assign _6857_ = _6491_ & _6860_ /*13413*/;
assign _6858_ = _6491_ ^ _6860_ /*13416*/;
assign _6859_ = _6851_ & _6858_ /*13414*/;
assign _6716_ = _6851_ ^ _6858_ /*13415*/;
assign _6856_ = _6857_ | _6859_ /*13412*/;
assign _6865_ = ~D[28] /*13411*/;
assign _6862_ = _6492_ & _6865_ /*13407*/;
assign _6863_ = _6492_ ^ _6865_ /*13410*/;
assign _6864_ = _6856_ & _6863_ /*13408*/;
assign _6717_ = _6856_ ^ _6863_ /*13409*/;
assign _6861_ = _6862_ | _6864_ /*13406*/;
assign _6870_ = ~D[29] /*13405*/;
assign _6867_ = _6493_ & _6870_ /*13401*/;
assign _6868_ = _6493_ ^ _6870_ /*13404*/;
assign _6869_ = _6861_ & _6868_ /*13402*/;
assign _6718_ = _6861_ ^ _6868_ /*13403*/;
assign _6866_ = _6867_ | _6869_ /*13400*/;
assign _6875_ = ~D[30] /*13399*/;
assign _6872_ = _6494_ & _6875_ /*13395*/;
assign _6873_ = _6494_ ^ _6875_ /*13398*/;
assign _6874_ = _6866_ & _6873_ /*13396*/;
assign _6719_ = _6866_ ^ _6873_ /*13397*/;
assign _6871_ = _6872_ | _6874_ /*13394*/;
assign _6876_ = _6495_ & oneWire /*13389*/;
assign _6877_ = _6495_ ^ oneWire /*13392*/;
assign _6878_ = _6871_ & _6877_ /*13390*/;
assign _6720_ = _6871_ ^ _6877_ /*13391*/;
assign Q[16] = _6876_ | _6878_ /*13388*/;
assign _6947_ = ~Q[16] /*13195*/;
assign _6946_ = _6947_ & D[0] /*13194*/;
assign _6949_ = _6689_ & _6946_ /*13189*/;
assign _6950_ = _6689_ ^ _6946_ /*13192*/;
assign _6951_ = zeroWire & _6950_ /*13190*/;
assign _6913_ = zeroWire ^ _6950_ /*13191*/;
assign _6948_ = _6949_ | _6951_ /*13188*/;
assign _6953_ = ~Q[16] /*13187*/;
assign _6952_ = _6953_ & D[1] /*13186*/;
assign _6955_ = _6690_ & _6952_ /*13181*/;
assign _6956_ = _6690_ ^ _6952_ /*13184*/;
assign _6957_ = _6948_ & _6956_ /*13182*/;
assign _6914_ = _6948_ ^ _6956_ /*13183*/;
assign _6954_ = _6955_ | _6957_ /*13180*/;
assign _6959_ = ~Q[16] /*13179*/;
assign _6958_ = _6959_ & D[2] /*13178*/;
assign _6961_ = _6691_ & _6958_ /*13173*/;
assign _6962_ = _6691_ ^ _6958_ /*13176*/;
assign _6963_ = _6954_ & _6962_ /*13174*/;
assign _6915_ = _6954_ ^ _6962_ /*13175*/;
assign _6960_ = _6961_ | _6963_ /*13172*/;
assign _6965_ = ~Q[16] /*13171*/;
assign _6964_ = _6965_ & D[3] /*13170*/;
assign _6967_ = _6692_ & _6964_ /*13165*/;
assign _6968_ = _6692_ ^ _6964_ /*13168*/;
assign _6969_ = _6960_ & _6968_ /*13166*/;
assign _6916_ = _6960_ ^ _6968_ /*13167*/;
assign _6966_ = _6967_ | _6969_ /*13164*/;
assign _6971_ = ~Q[16] /*13163*/;
assign _6970_ = _6971_ & D[4] /*13162*/;
assign _6973_ = _6693_ & _6970_ /*13157*/;
assign _6974_ = _6693_ ^ _6970_ /*13160*/;
assign _6975_ = _6966_ & _6974_ /*13158*/;
assign _6917_ = _6966_ ^ _6974_ /*13159*/;
assign _6972_ = _6973_ | _6975_ /*13156*/;
assign _6977_ = ~Q[16] /*13155*/;
assign _6976_ = _6977_ & D[5] /*13154*/;
assign _6979_ = _6694_ & _6976_ /*13149*/;
assign _6980_ = _6694_ ^ _6976_ /*13152*/;
assign _6981_ = _6972_ & _6980_ /*13150*/;
assign _6918_ = _6972_ ^ _6980_ /*13151*/;
assign _6978_ = _6979_ | _6981_ /*13148*/;
assign _6983_ = ~Q[16] /*13147*/;
assign _6982_ = _6983_ & D[6] /*13146*/;
assign _6985_ = _6695_ & _6982_ /*13141*/;
assign _6986_ = _6695_ ^ _6982_ /*13144*/;
assign _6987_ = _6978_ & _6986_ /*13142*/;
assign _6919_ = _6978_ ^ _6986_ /*13143*/;
assign _6984_ = _6985_ | _6987_ /*13140*/;
assign _6989_ = ~Q[16] /*13139*/;
assign _6988_ = _6989_ & D[7] /*13138*/;
assign _6991_ = _6696_ & _6988_ /*13133*/;
assign _6992_ = _6696_ ^ _6988_ /*13136*/;
assign _6993_ = _6984_ & _6992_ /*13134*/;
assign _6920_ = _6984_ ^ _6992_ /*13135*/;
assign _6990_ = _6991_ | _6993_ /*13132*/;
assign _6995_ = ~Q[16] /*13131*/;
assign _6994_ = _6995_ & D[8] /*13130*/;
assign _6997_ = _6697_ & _6994_ /*13125*/;
assign _6998_ = _6697_ ^ _6994_ /*13128*/;
assign _6999_ = _6990_ & _6998_ /*13126*/;
assign _6921_ = _6990_ ^ _6998_ /*13127*/;
assign _6996_ = _6997_ | _6999_ /*13124*/;
assign _7001_ = ~Q[16] /*13123*/;
assign _7000_ = _7001_ & D[9] /*13122*/;
assign _7003_ = _6698_ & _7000_ /*13117*/;
assign _7004_ = _6698_ ^ _7000_ /*13120*/;
assign _7005_ = _6996_ & _7004_ /*13118*/;
assign _6922_ = _6996_ ^ _7004_ /*13119*/;
assign _7002_ = _7003_ | _7005_ /*13116*/;
assign _7007_ = ~Q[16] /*13115*/;
assign _7006_ = _7007_ & D[10] /*13114*/;
assign _7009_ = _6699_ & _7006_ /*13109*/;
assign _7010_ = _6699_ ^ _7006_ /*13112*/;
assign _7011_ = _7002_ & _7010_ /*13110*/;
assign _6923_ = _7002_ ^ _7010_ /*13111*/;
assign _7008_ = _7009_ | _7011_ /*13108*/;
assign _7013_ = ~Q[16] /*13107*/;
assign _7012_ = _7013_ & D[11] /*13106*/;
assign _7015_ = _6700_ & _7012_ /*13101*/;
assign _7016_ = _6700_ ^ _7012_ /*13104*/;
assign _7017_ = _7008_ & _7016_ /*13102*/;
assign _6924_ = _7008_ ^ _7016_ /*13103*/;
assign _7014_ = _7015_ | _7017_ /*13100*/;
assign _7019_ = ~Q[16] /*13099*/;
assign _7018_ = _7019_ & D[12] /*13098*/;
assign _7021_ = _6701_ & _7018_ /*13093*/;
assign _7022_ = _6701_ ^ _7018_ /*13096*/;
assign _7023_ = _7014_ & _7022_ /*13094*/;
assign _6925_ = _7014_ ^ _7022_ /*13095*/;
assign _7020_ = _7021_ | _7023_ /*13092*/;
assign _7025_ = ~Q[16] /*13091*/;
assign _7024_ = _7025_ & D[13] /*13090*/;
assign _7027_ = _6702_ & _7024_ /*13085*/;
assign _7028_ = _6702_ ^ _7024_ /*13088*/;
assign _7029_ = _7020_ & _7028_ /*13086*/;
assign _6926_ = _7020_ ^ _7028_ /*13087*/;
assign _7026_ = _7027_ | _7029_ /*13084*/;
assign _7031_ = ~Q[16] /*13083*/;
assign _7030_ = _7031_ & D[14] /*13082*/;
assign _7033_ = _6703_ & _7030_ /*13077*/;
assign _7034_ = _6703_ ^ _7030_ /*13080*/;
assign _7035_ = _7026_ & _7034_ /*13078*/;
assign _6927_ = _7026_ ^ _7034_ /*13079*/;
assign _7032_ = _7033_ | _7035_ /*13076*/;
assign _7037_ = ~Q[16] /*13075*/;
assign _7036_ = _7037_ & D[15] /*13074*/;
assign _7039_ = _6704_ & _7036_ /*13069*/;
assign _7040_ = _6704_ ^ _7036_ /*13072*/;
assign _7041_ = _7032_ & _7040_ /*13070*/;
assign _6928_ = _7032_ ^ _7040_ /*13071*/;
assign _7038_ = _7039_ | _7041_ /*13068*/;
assign _7043_ = ~Q[16] /*13067*/;
assign _7042_ = _7043_ & D[16] /*13066*/;
assign _7045_ = _6705_ & _7042_ /*13061*/;
assign _7046_ = _6705_ ^ _7042_ /*13064*/;
assign _7047_ = _7038_ & _7046_ /*13062*/;
assign _6929_ = _7038_ ^ _7046_ /*13063*/;
assign _7044_ = _7045_ | _7047_ /*13060*/;
assign _7049_ = ~Q[16] /*13059*/;
assign _7048_ = _7049_ & D[17] /*13058*/;
assign _7051_ = _6706_ & _7048_ /*13053*/;
assign _7052_ = _6706_ ^ _7048_ /*13056*/;
assign _7053_ = _7044_ & _7052_ /*13054*/;
assign _6930_ = _7044_ ^ _7052_ /*13055*/;
assign _7050_ = _7051_ | _7053_ /*13052*/;
assign _7055_ = ~Q[16] /*13051*/;
assign _7054_ = _7055_ & D[18] /*13050*/;
assign _7057_ = _6707_ & _7054_ /*13045*/;
assign _7058_ = _6707_ ^ _7054_ /*13048*/;
assign _7059_ = _7050_ & _7058_ /*13046*/;
assign _6931_ = _7050_ ^ _7058_ /*13047*/;
assign _7056_ = _7057_ | _7059_ /*13044*/;
assign _7061_ = ~Q[16] /*13043*/;
assign _7060_ = _7061_ & D[19] /*13042*/;
assign _7063_ = _6708_ & _7060_ /*13037*/;
assign _7064_ = _6708_ ^ _7060_ /*13040*/;
assign _7065_ = _7056_ & _7064_ /*13038*/;
assign _6932_ = _7056_ ^ _7064_ /*13039*/;
assign _7062_ = _7063_ | _7065_ /*13036*/;
assign _7067_ = ~Q[16] /*13035*/;
assign _7066_ = _7067_ & D[20] /*13034*/;
assign _7069_ = _6709_ & _7066_ /*13029*/;
assign _7070_ = _6709_ ^ _7066_ /*13032*/;
assign _7071_ = _7062_ & _7070_ /*13030*/;
assign _6933_ = _7062_ ^ _7070_ /*13031*/;
assign _7068_ = _7069_ | _7071_ /*13028*/;
assign _7073_ = ~Q[16] /*13027*/;
assign _7072_ = _7073_ & D[21] /*13026*/;
assign _7075_ = _6710_ & _7072_ /*13021*/;
assign _7076_ = _6710_ ^ _7072_ /*13024*/;
assign _7077_ = _7068_ & _7076_ /*13022*/;
assign _6934_ = _7068_ ^ _7076_ /*13023*/;
assign _7074_ = _7075_ | _7077_ /*13020*/;
assign _7079_ = ~Q[16] /*13019*/;
assign _7078_ = _7079_ & D[22] /*13018*/;
assign _7081_ = _6711_ & _7078_ /*13013*/;
assign _7082_ = _6711_ ^ _7078_ /*13016*/;
assign _7083_ = _7074_ & _7082_ /*13014*/;
assign _6935_ = _7074_ ^ _7082_ /*13015*/;
assign _7080_ = _7081_ | _7083_ /*13012*/;
assign _7085_ = ~Q[16] /*13011*/;
assign _7084_ = _7085_ & D[23] /*13010*/;
assign _7087_ = _6712_ & _7084_ /*13005*/;
assign _7088_ = _6712_ ^ _7084_ /*13008*/;
assign _7089_ = _7080_ & _7088_ /*13006*/;
assign _6936_ = _7080_ ^ _7088_ /*13007*/;
assign _7086_ = _7087_ | _7089_ /*13004*/;
assign _7091_ = ~Q[16] /*13003*/;
assign _7090_ = _7091_ & D[24] /*13002*/;
assign _7093_ = _6713_ & _7090_ /*12997*/;
assign _7094_ = _6713_ ^ _7090_ /*13000*/;
assign _7095_ = _7086_ & _7094_ /*12998*/;
assign _6937_ = _7086_ ^ _7094_ /*12999*/;
assign _7092_ = _7093_ | _7095_ /*12996*/;
assign _7097_ = ~Q[16] /*12995*/;
assign _7096_ = _7097_ & D[25] /*12994*/;
assign _7099_ = _6714_ & _7096_ /*12989*/;
assign _7100_ = _6714_ ^ _7096_ /*12992*/;
assign _7101_ = _7092_ & _7100_ /*12990*/;
assign _6938_ = _7092_ ^ _7100_ /*12991*/;
assign _7098_ = _7099_ | _7101_ /*12988*/;
assign _7103_ = ~Q[16] /*12987*/;
assign _7102_ = _7103_ & D[26] /*12986*/;
assign _7105_ = _6715_ & _7102_ /*12981*/;
assign _7106_ = _6715_ ^ _7102_ /*12984*/;
assign _7107_ = _7098_ & _7106_ /*12982*/;
assign _6939_ = _7098_ ^ _7106_ /*12983*/;
assign _7104_ = _7105_ | _7107_ /*12980*/;
assign _7109_ = ~Q[16] /*12979*/;
assign _7108_ = _7109_ & D[27] /*12978*/;
assign _7111_ = _6716_ & _7108_ /*12973*/;
assign _7112_ = _6716_ ^ _7108_ /*12976*/;
assign _7113_ = _7104_ & _7112_ /*12974*/;
assign _6940_ = _7104_ ^ _7112_ /*12975*/;
assign _7110_ = _7111_ | _7113_ /*12972*/;
assign _7115_ = ~Q[16] /*12971*/;
assign _7114_ = _7115_ & D[28] /*12970*/;
assign _7117_ = _6717_ & _7114_ /*12965*/;
assign _7118_ = _6717_ ^ _7114_ /*12968*/;
assign _7119_ = _7110_ & _7118_ /*12966*/;
assign _6941_ = _7110_ ^ _7118_ /*12967*/;
assign _7116_ = _7117_ | _7119_ /*12964*/;
assign _7121_ = ~Q[16] /*12963*/;
assign _7120_ = _7121_ & D[29] /*12962*/;
assign _7123_ = _6718_ & _7120_ /*12957*/;
assign _7124_ = _6718_ ^ _7120_ /*12960*/;
assign _7125_ = _7116_ & _7124_ /*12958*/;
assign _6942_ = _7116_ ^ _7124_ /*12959*/;
assign _7122_ = _7123_ | _7125_ /*12956*/;
assign _7127_ = ~Q[16] /*12955*/;
assign _7126_ = _7127_ & D[30] /*12954*/;
assign _7129_ = _6719_ & _7126_ /*12949*/;
assign _7130_ = _6719_ ^ _7126_ /*12952*/;
assign _7131_ = _7122_ & _7130_ /*12950*/;
assign _6943_ = _7122_ ^ _7130_ /*12951*/;
assign _7128_ = _7129_ | _7131_ /*12948*/;
assign _7133_ = ~Q[16] /*12947*/;
assign _7132_ = _7133_ & zeroWire /*12946*/;
assign _7134_ = _6720_ ^ _7132_ /*12944*/;
assign _6944_ = _7134_ ^ _7128_ /*12943*/;
assign _7173_ = ~D[0] /*12817*/;
assign _7170_ = R_0[15] & _7173_ /*12813*/;
assign _7171_ = R_0[15] ^ _7173_ /*12816*/;
assign _7172_ = oneWire & _7171_ /*12814*/;
assign _7137_ = oneWire ^ _7171_ /*12815*/;
assign _7169_ = _7170_ | _7172_ /*12812*/;
assign _7178_ = ~D[1] /*12811*/;
assign _7175_ = _6913_ & _7178_ /*12807*/;
assign _7176_ = _6913_ ^ _7178_ /*12810*/;
assign _7177_ = _7169_ & _7176_ /*12808*/;
assign _7138_ = _7169_ ^ _7176_ /*12809*/;
assign _7174_ = _7175_ | _7177_ /*12806*/;
assign _7183_ = ~D[2] /*12805*/;
assign _7180_ = _6914_ & _7183_ /*12801*/;
assign _7181_ = _6914_ ^ _7183_ /*12804*/;
assign _7182_ = _7174_ & _7181_ /*12802*/;
assign _7139_ = _7174_ ^ _7181_ /*12803*/;
assign _7179_ = _7180_ | _7182_ /*12800*/;
assign _7188_ = ~D[3] /*12799*/;
assign _7185_ = _6915_ & _7188_ /*12795*/;
assign _7186_ = _6915_ ^ _7188_ /*12798*/;
assign _7187_ = _7179_ & _7186_ /*12796*/;
assign _7140_ = _7179_ ^ _7186_ /*12797*/;
assign _7184_ = _7185_ | _7187_ /*12794*/;
assign _7193_ = ~D[4] /*12793*/;
assign _7190_ = _6916_ & _7193_ /*12789*/;
assign _7191_ = _6916_ ^ _7193_ /*12792*/;
assign _7192_ = _7184_ & _7191_ /*12790*/;
assign _7141_ = _7184_ ^ _7191_ /*12791*/;
assign _7189_ = _7190_ | _7192_ /*12788*/;
assign _7198_ = ~D[5] /*12787*/;
assign _7195_ = _6917_ & _7198_ /*12783*/;
assign _7196_ = _6917_ ^ _7198_ /*12786*/;
assign _7197_ = _7189_ & _7196_ /*12784*/;
assign _7142_ = _7189_ ^ _7196_ /*12785*/;
assign _7194_ = _7195_ | _7197_ /*12782*/;
assign _7203_ = ~D[6] /*12781*/;
assign _7200_ = _6918_ & _7203_ /*12777*/;
assign _7201_ = _6918_ ^ _7203_ /*12780*/;
assign _7202_ = _7194_ & _7201_ /*12778*/;
assign _7143_ = _7194_ ^ _7201_ /*12779*/;
assign _7199_ = _7200_ | _7202_ /*12776*/;
assign _7208_ = ~D[7] /*12775*/;
assign _7205_ = _6919_ & _7208_ /*12771*/;
assign _7206_ = _6919_ ^ _7208_ /*12774*/;
assign _7207_ = _7199_ & _7206_ /*12772*/;
assign _7144_ = _7199_ ^ _7206_ /*12773*/;
assign _7204_ = _7205_ | _7207_ /*12770*/;
assign _7213_ = ~D[8] /*12769*/;
assign _7210_ = _6920_ & _7213_ /*12765*/;
assign _7211_ = _6920_ ^ _7213_ /*12768*/;
assign _7212_ = _7204_ & _7211_ /*12766*/;
assign _7145_ = _7204_ ^ _7211_ /*12767*/;
assign _7209_ = _7210_ | _7212_ /*12764*/;
assign _7218_ = ~D[9] /*12763*/;
assign _7215_ = _6921_ & _7218_ /*12759*/;
assign _7216_ = _6921_ ^ _7218_ /*12762*/;
assign _7217_ = _7209_ & _7216_ /*12760*/;
assign _7146_ = _7209_ ^ _7216_ /*12761*/;
assign _7214_ = _7215_ | _7217_ /*12758*/;
assign _7223_ = ~D[10] /*12757*/;
assign _7220_ = _6922_ & _7223_ /*12753*/;
assign _7221_ = _6922_ ^ _7223_ /*12756*/;
assign _7222_ = _7214_ & _7221_ /*12754*/;
assign _7147_ = _7214_ ^ _7221_ /*12755*/;
assign _7219_ = _7220_ | _7222_ /*12752*/;
assign _7228_ = ~D[11] /*12751*/;
assign _7225_ = _6923_ & _7228_ /*12747*/;
assign _7226_ = _6923_ ^ _7228_ /*12750*/;
assign _7227_ = _7219_ & _7226_ /*12748*/;
assign _7148_ = _7219_ ^ _7226_ /*12749*/;
assign _7224_ = _7225_ | _7227_ /*12746*/;
assign _7233_ = ~D[12] /*12745*/;
assign _7230_ = _6924_ & _7233_ /*12741*/;
assign _7231_ = _6924_ ^ _7233_ /*12744*/;
assign _7232_ = _7224_ & _7231_ /*12742*/;
assign _7149_ = _7224_ ^ _7231_ /*12743*/;
assign _7229_ = _7230_ | _7232_ /*12740*/;
assign _7238_ = ~D[13] /*12739*/;
assign _7235_ = _6925_ & _7238_ /*12735*/;
assign _7236_ = _6925_ ^ _7238_ /*12738*/;
assign _7237_ = _7229_ & _7236_ /*12736*/;
assign _7150_ = _7229_ ^ _7236_ /*12737*/;
assign _7234_ = _7235_ | _7237_ /*12734*/;
assign _7243_ = ~D[14] /*12733*/;
assign _7240_ = _6926_ & _7243_ /*12729*/;
assign _7241_ = _6926_ ^ _7243_ /*12732*/;
assign _7242_ = _7234_ & _7241_ /*12730*/;
assign _7151_ = _7234_ ^ _7241_ /*12731*/;
assign _7239_ = _7240_ | _7242_ /*12728*/;
assign _7248_ = ~D[15] /*12727*/;
assign _7245_ = _6927_ & _7248_ /*12723*/;
assign _7246_ = _6927_ ^ _7248_ /*12726*/;
assign _7247_ = _7239_ & _7246_ /*12724*/;
assign _7152_ = _7239_ ^ _7246_ /*12725*/;
assign _7244_ = _7245_ | _7247_ /*12722*/;
assign _7253_ = ~D[16] /*12721*/;
assign _7250_ = _6928_ & _7253_ /*12717*/;
assign _7251_ = _6928_ ^ _7253_ /*12720*/;
assign _7252_ = _7244_ & _7251_ /*12718*/;
assign _7153_ = _7244_ ^ _7251_ /*12719*/;
assign _7249_ = _7250_ | _7252_ /*12716*/;
assign _7258_ = ~D[17] /*12715*/;
assign _7255_ = _6929_ & _7258_ /*12711*/;
assign _7256_ = _6929_ ^ _7258_ /*12714*/;
assign _7257_ = _7249_ & _7256_ /*12712*/;
assign _7154_ = _7249_ ^ _7256_ /*12713*/;
assign _7254_ = _7255_ | _7257_ /*12710*/;
assign _7263_ = ~D[18] /*12709*/;
assign _7260_ = _6930_ & _7263_ /*12705*/;
assign _7261_ = _6930_ ^ _7263_ /*12708*/;
assign _7262_ = _7254_ & _7261_ /*12706*/;
assign _7155_ = _7254_ ^ _7261_ /*12707*/;
assign _7259_ = _7260_ | _7262_ /*12704*/;
assign _7268_ = ~D[19] /*12703*/;
assign _7265_ = _6931_ & _7268_ /*12699*/;
assign _7266_ = _6931_ ^ _7268_ /*12702*/;
assign _7267_ = _7259_ & _7266_ /*12700*/;
assign _7156_ = _7259_ ^ _7266_ /*12701*/;
assign _7264_ = _7265_ | _7267_ /*12698*/;
assign _7273_ = ~D[20] /*12697*/;
assign _7270_ = _6932_ & _7273_ /*12693*/;
assign _7271_ = _6932_ ^ _7273_ /*12696*/;
assign _7272_ = _7264_ & _7271_ /*12694*/;
assign _7157_ = _7264_ ^ _7271_ /*12695*/;
assign _7269_ = _7270_ | _7272_ /*12692*/;
assign _7278_ = ~D[21] /*12691*/;
assign _7275_ = _6933_ & _7278_ /*12687*/;
assign _7276_ = _6933_ ^ _7278_ /*12690*/;
assign _7277_ = _7269_ & _7276_ /*12688*/;
assign _7158_ = _7269_ ^ _7276_ /*12689*/;
assign _7274_ = _7275_ | _7277_ /*12686*/;
assign _7283_ = ~D[22] /*12685*/;
assign _7280_ = _6934_ & _7283_ /*12681*/;
assign _7281_ = _6934_ ^ _7283_ /*12684*/;
assign _7282_ = _7274_ & _7281_ /*12682*/;
assign _7159_ = _7274_ ^ _7281_ /*12683*/;
assign _7279_ = _7280_ | _7282_ /*12680*/;
assign _7288_ = ~D[23] /*12679*/;
assign _7285_ = _6935_ & _7288_ /*12675*/;
assign _7286_ = _6935_ ^ _7288_ /*12678*/;
assign _7287_ = _7279_ & _7286_ /*12676*/;
assign _7160_ = _7279_ ^ _7286_ /*12677*/;
assign _7284_ = _7285_ | _7287_ /*12674*/;
assign _7293_ = ~D[24] /*12673*/;
assign _7290_ = _6936_ & _7293_ /*12669*/;
assign _7291_ = _6936_ ^ _7293_ /*12672*/;
assign _7292_ = _7284_ & _7291_ /*12670*/;
assign _7161_ = _7284_ ^ _7291_ /*12671*/;
assign _7289_ = _7290_ | _7292_ /*12668*/;
assign _7298_ = ~D[25] /*12667*/;
assign _7295_ = _6937_ & _7298_ /*12663*/;
assign _7296_ = _6937_ ^ _7298_ /*12666*/;
assign _7297_ = _7289_ & _7296_ /*12664*/;
assign _7162_ = _7289_ ^ _7296_ /*12665*/;
assign _7294_ = _7295_ | _7297_ /*12662*/;
assign _7303_ = ~D[26] /*12661*/;
assign _7300_ = _6938_ & _7303_ /*12657*/;
assign _7301_ = _6938_ ^ _7303_ /*12660*/;
assign _7302_ = _7294_ & _7301_ /*12658*/;
assign _7163_ = _7294_ ^ _7301_ /*12659*/;
assign _7299_ = _7300_ | _7302_ /*12656*/;
assign _7308_ = ~D[27] /*12655*/;
assign _7305_ = _6939_ & _7308_ /*12651*/;
assign _7306_ = _6939_ ^ _7308_ /*12654*/;
assign _7307_ = _7299_ & _7306_ /*12652*/;
assign _7164_ = _7299_ ^ _7306_ /*12653*/;
assign _7304_ = _7305_ | _7307_ /*12650*/;
assign _7313_ = ~D[28] /*12649*/;
assign _7310_ = _6940_ & _7313_ /*12645*/;
assign _7311_ = _6940_ ^ _7313_ /*12648*/;
assign _7312_ = _7304_ & _7311_ /*12646*/;
assign _7165_ = _7304_ ^ _7311_ /*12647*/;
assign _7309_ = _7310_ | _7312_ /*12644*/;
assign _7318_ = ~D[29] /*12643*/;
assign _7315_ = _6941_ & _7318_ /*12639*/;
assign _7316_ = _6941_ ^ _7318_ /*12642*/;
assign _7317_ = _7309_ & _7316_ /*12640*/;
assign _7166_ = _7309_ ^ _7316_ /*12641*/;
assign _7314_ = _7315_ | _7317_ /*12638*/;
assign _7323_ = ~D[30] /*12637*/;
assign _7320_ = _6942_ & _7323_ /*12633*/;
assign _7321_ = _6942_ ^ _7323_ /*12636*/;
assign _7322_ = _7314_ & _7321_ /*12634*/;
assign _7167_ = _7314_ ^ _7321_ /*12635*/;
assign _7319_ = _7320_ | _7322_ /*12632*/;
assign _7324_ = _6943_ & oneWire /*12627*/;
assign _7325_ = _6943_ ^ oneWire /*12630*/;
assign _7326_ = _7319_ & _7325_ /*12628*/;
assign _7168_ = _7319_ ^ _7325_ /*12629*/;
assign Q[15] = _7324_ | _7326_ /*12626*/;
assign _7395_ = ~Q[15] /*12433*/;
assign _7394_ = _7395_ & D[0] /*12432*/;
assign _7397_ = _7137_ & _7394_ /*12427*/;
assign _7398_ = _7137_ ^ _7394_ /*12430*/;
assign _7399_ = zeroWire & _7398_ /*12428*/;
assign _7361_ = zeroWire ^ _7398_ /*12429*/;
assign _7396_ = _7397_ | _7399_ /*12426*/;
assign _7401_ = ~Q[15] /*12425*/;
assign _7400_ = _7401_ & D[1] /*12424*/;
assign _7403_ = _7138_ & _7400_ /*12419*/;
assign _7404_ = _7138_ ^ _7400_ /*12422*/;
assign _7405_ = _7396_ & _7404_ /*12420*/;
assign _7362_ = _7396_ ^ _7404_ /*12421*/;
assign _7402_ = _7403_ | _7405_ /*12418*/;
assign _7407_ = ~Q[15] /*12417*/;
assign _7406_ = _7407_ & D[2] /*12416*/;
assign _7409_ = _7139_ & _7406_ /*12411*/;
assign _7410_ = _7139_ ^ _7406_ /*12414*/;
assign _7411_ = _7402_ & _7410_ /*12412*/;
assign _7363_ = _7402_ ^ _7410_ /*12413*/;
assign _7408_ = _7409_ | _7411_ /*12410*/;
assign _7413_ = ~Q[15] /*12409*/;
assign _7412_ = _7413_ & D[3] /*12408*/;
assign _7415_ = _7140_ & _7412_ /*12403*/;
assign _7416_ = _7140_ ^ _7412_ /*12406*/;
assign _7417_ = _7408_ & _7416_ /*12404*/;
assign _7364_ = _7408_ ^ _7416_ /*12405*/;
assign _7414_ = _7415_ | _7417_ /*12402*/;
assign _7419_ = ~Q[15] /*12401*/;
assign _7418_ = _7419_ & D[4] /*12400*/;
assign _7421_ = _7141_ & _7418_ /*12395*/;
assign _7422_ = _7141_ ^ _7418_ /*12398*/;
assign _7423_ = _7414_ & _7422_ /*12396*/;
assign _7365_ = _7414_ ^ _7422_ /*12397*/;
assign _7420_ = _7421_ | _7423_ /*12394*/;
assign _7425_ = ~Q[15] /*12393*/;
assign _7424_ = _7425_ & D[5] /*12392*/;
assign _7427_ = _7142_ & _7424_ /*12387*/;
assign _7428_ = _7142_ ^ _7424_ /*12390*/;
assign _7429_ = _7420_ & _7428_ /*12388*/;
assign _7366_ = _7420_ ^ _7428_ /*12389*/;
assign _7426_ = _7427_ | _7429_ /*12386*/;
assign _7431_ = ~Q[15] /*12385*/;
assign _7430_ = _7431_ & D[6] /*12384*/;
assign _7433_ = _7143_ & _7430_ /*12379*/;
assign _7434_ = _7143_ ^ _7430_ /*12382*/;
assign _7435_ = _7426_ & _7434_ /*12380*/;
assign _7367_ = _7426_ ^ _7434_ /*12381*/;
assign _7432_ = _7433_ | _7435_ /*12378*/;
assign _7437_ = ~Q[15] /*12377*/;
assign _7436_ = _7437_ & D[7] /*12376*/;
assign _7439_ = _7144_ & _7436_ /*12371*/;
assign _7440_ = _7144_ ^ _7436_ /*12374*/;
assign _7441_ = _7432_ & _7440_ /*12372*/;
assign _7368_ = _7432_ ^ _7440_ /*12373*/;
assign _7438_ = _7439_ | _7441_ /*12370*/;
assign _7443_ = ~Q[15] /*12369*/;
assign _7442_ = _7443_ & D[8] /*12368*/;
assign _7445_ = _7145_ & _7442_ /*12363*/;
assign _7446_ = _7145_ ^ _7442_ /*12366*/;
assign _7447_ = _7438_ & _7446_ /*12364*/;
assign _7369_ = _7438_ ^ _7446_ /*12365*/;
assign _7444_ = _7445_ | _7447_ /*12362*/;
assign _7449_ = ~Q[15] /*12361*/;
assign _7448_ = _7449_ & D[9] /*12360*/;
assign _7451_ = _7146_ & _7448_ /*12355*/;
assign _7452_ = _7146_ ^ _7448_ /*12358*/;
assign _7453_ = _7444_ & _7452_ /*12356*/;
assign _7370_ = _7444_ ^ _7452_ /*12357*/;
assign _7450_ = _7451_ | _7453_ /*12354*/;
assign _7455_ = ~Q[15] /*12353*/;
assign _7454_ = _7455_ & D[10] /*12352*/;
assign _7457_ = _7147_ & _7454_ /*12347*/;
assign _7458_ = _7147_ ^ _7454_ /*12350*/;
assign _7459_ = _7450_ & _7458_ /*12348*/;
assign _7371_ = _7450_ ^ _7458_ /*12349*/;
assign _7456_ = _7457_ | _7459_ /*12346*/;
assign _7461_ = ~Q[15] /*12345*/;
assign _7460_ = _7461_ & D[11] /*12344*/;
assign _7463_ = _7148_ & _7460_ /*12339*/;
assign _7464_ = _7148_ ^ _7460_ /*12342*/;
assign _7465_ = _7456_ & _7464_ /*12340*/;
assign _7372_ = _7456_ ^ _7464_ /*12341*/;
assign _7462_ = _7463_ | _7465_ /*12338*/;
assign _7467_ = ~Q[15] /*12337*/;
assign _7466_ = _7467_ & D[12] /*12336*/;
assign _7469_ = _7149_ & _7466_ /*12331*/;
assign _7470_ = _7149_ ^ _7466_ /*12334*/;
assign _7471_ = _7462_ & _7470_ /*12332*/;
assign _7373_ = _7462_ ^ _7470_ /*12333*/;
assign _7468_ = _7469_ | _7471_ /*12330*/;
assign _7473_ = ~Q[15] /*12329*/;
assign _7472_ = _7473_ & D[13] /*12328*/;
assign _7475_ = _7150_ & _7472_ /*12323*/;
assign _7476_ = _7150_ ^ _7472_ /*12326*/;
assign _7477_ = _7468_ & _7476_ /*12324*/;
assign _7374_ = _7468_ ^ _7476_ /*12325*/;
assign _7474_ = _7475_ | _7477_ /*12322*/;
assign _7479_ = ~Q[15] /*12321*/;
assign _7478_ = _7479_ & D[14] /*12320*/;
assign _7481_ = _7151_ & _7478_ /*12315*/;
assign _7482_ = _7151_ ^ _7478_ /*12318*/;
assign _7483_ = _7474_ & _7482_ /*12316*/;
assign _7375_ = _7474_ ^ _7482_ /*12317*/;
assign _7480_ = _7481_ | _7483_ /*12314*/;
assign _7485_ = ~Q[15] /*12313*/;
assign _7484_ = _7485_ & D[15] /*12312*/;
assign _7487_ = _7152_ & _7484_ /*12307*/;
assign _7488_ = _7152_ ^ _7484_ /*12310*/;
assign _7489_ = _7480_ & _7488_ /*12308*/;
assign _7376_ = _7480_ ^ _7488_ /*12309*/;
assign _7486_ = _7487_ | _7489_ /*12306*/;
assign _7491_ = ~Q[15] /*12305*/;
assign _7490_ = _7491_ & D[16] /*12304*/;
assign _7493_ = _7153_ & _7490_ /*12299*/;
assign _7494_ = _7153_ ^ _7490_ /*12302*/;
assign _7495_ = _7486_ & _7494_ /*12300*/;
assign _7377_ = _7486_ ^ _7494_ /*12301*/;
assign _7492_ = _7493_ | _7495_ /*12298*/;
assign _7497_ = ~Q[15] /*12297*/;
assign _7496_ = _7497_ & D[17] /*12296*/;
assign _7499_ = _7154_ & _7496_ /*12291*/;
assign _7500_ = _7154_ ^ _7496_ /*12294*/;
assign _7501_ = _7492_ & _7500_ /*12292*/;
assign _7378_ = _7492_ ^ _7500_ /*12293*/;
assign _7498_ = _7499_ | _7501_ /*12290*/;
assign _7503_ = ~Q[15] /*12289*/;
assign _7502_ = _7503_ & D[18] /*12288*/;
assign _7505_ = _7155_ & _7502_ /*12283*/;
assign _7506_ = _7155_ ^ _7502_ /*12286*/;
assign _7507_ = _7498_ & _7506_ /*12284*/;
assign _7379_ = _7498_ ^ _7506_ /*12285*/;
assign _7504_ = _7505_ | _7507_ /*12282*/;
assign _7509_ = ~Q[15] /*12281*/;
assign _7508_ = _7509_ & D[19] /*12280*/;
assign _7511_ = _7156_ & _7508_ /*12275*/;
assign _7512_ = _7156_ ^ _7508_ /*12278*/;
assign _7513_ = _7504_ & _7512_ /*12276*/;
assign _7380_ = _7504_ ^ _7512_ /*12277*/;
assign _7510_ = _7511_ | _7513_ /*12274*/;
assign _7515_ = ~Q[15] /*12273*/;
assign _7514_ = _7515_ & D[20] /*12272*/;
assign _7517_ = _7157_ & _7514_ /*12267*/;
assign _7518_ = _7157_ ^ _7514_ /*12270*/;
assign _7519_ = _7510_ & _7518_ /*12268*/;
assign _7381_ = _7510_ ^ _7518_ /*12269*/;
assign _7516_ = _7517_ | _7519_ /*12266*/;
assign _7521_ = ~Q[15] /*12265*/;
assign _7520_ = _7521_ & D[21] /*12264*/;
assign _7523_ = _7158_ & _7520_ /*12259*/;
assign _7524_ = _7158_ ^ _7520_ /*12262*/;
assign _7525_ = _7516_ & _7524_ /*12260*/;
assign _7382_ = _7516_ ^ _7524_ /*12261*/;
assign _7522_ = _7523_ | _7525_ /*12258*/;
assign _7527_ = ~Q[15] /*12257*/;
assign _7526_ = _7527_ & D[22] /*12256*/;
assign _7529_ = _7159_ & _7526_ /*12251*/;
assign _7530_ = _7159_ ^ _7526_ /*12254*/;
assign _7531_ = _7522_ & _7530_ /*12252*/;
assign _7383_ = _7522_ ^ _7530_ /*12253*/;
assign _7528_ = _7529_ | _7531_ /*12250*/;
assign _7533_ = ~Q[15] /*12249*/;
assign _7532_ = _7533_ & D[23] /*12248*/;
assign _7535_ = _7160_ & _7532_ /*12243*/;
assign _7536_ = _7160_ ^ _7532_ /*12246*/;
assign _7537_ = _7528_ & _7536_ /*12244*/;
assign _7384_ = _7528_ ^ _7536_ /*12245*/;
assign _7534_ = _7535_ | _7537_ /*12242*/;
assign _7539_ = ~Q[15] /*12241*/;
assign _7538_ = _7539_ & D[24] /*12240*/;
assign _7541_ = _7161_ & _7538_ /*12235*/;
assign _7542_ = _7161_ ^ _7538_ /*12238*/;
assign _7543_ = _7534_ & _7542_ /*12236*/;
assign _7385_ = _7534_ ^ _7542_ /*12237*/;
assign _7540_ = _7541_ | _7543_ /*12234*/;
assign _7545_ = ~Q[15] /*12233*/;
assign _7544_ = _7545_ & D[25] /*12232*/;
assign _7547_ = _7162_ & _7544_ /*12227*/;
assign _7548_ = _7162_ ^ _7544_ /*12230*/;
assign _7549_ = _7540_ & _7548_ /*12228*/;
assign _7386_ = _7540_ ^ _7548_ /*12229*/;
assign _7546_ = _7547_ | _7549_ /*12226*/;
assign _7551_ = ~Q[15] /*12225*/;
assign _7550_ = _7551_ & D[26] /*12224*/;
assign _7553_ = _7163_ & _7550_ /*12219*/;
assign _7554_ = _7163_ ^ _7550_ /*12222*/;
assign _7555_ = _7546_ & _7554_ /*12220*/;
assign _7387_ = _7546_ ^ _7554_ /*12221*/;
assign _7552_ = _7553_ | _7555_ /*12218*/;
assign _7557_ = ~Q[15] /*12217*/;
assign _7556_ = _7557_ & D[27] /*12216*/;
assign _7559_ = _7164_ & _7556_ /*12211*/;
assign _7560_ = _7164_ ^ _7556_ /*12214*/;
assign _7561_ = _7552_ & _7560_ /*12212*/;
assign _7388_ = _7552_ ^ _7560_ /*12213*/;
assign _7558_ = _7559_ | _7561_ /*12210*/;
assign _7563_ = ~Q[15] /*12209*/;
assign _7562_ = _7563_ & D[28] /*12208*/;
assign _7565_ = _7165_ & _7562_ /*12203*/;
assign _7566_ = _7165_ ^ _7562_ /*12206*/;
assign _7567_ = _7558_ & _7566_ /*12204*/;
assign _7389_ = _7558_ ^ _7566_ /*12205*/;
assign _7564_ = _7565_ | _7567_ /*12202*/;
assign _7569_ = ~Q[15] /*12201*/;
assign _7568_ = _7569_ & D[29] /*12200*/;
assign _7571_ = _7166_ & _7568_ /*12195*/;
assign _7572_ = _7166_ ^ _7568_ /*12198*/;
assign _7573_ = _7564_ & _7572_ /*12196*/;
assign _7390_ = _7564_ ^ _7572_ /*12197*/;
assign _7570_ = _7571_ | _7573_ /*12194*/;
assign _7575_ = ~Q[15] /*12193*/;
assign _7574_ = _7575_ & D[30] /*12192*/;
assign _7577_ = _7167_ & _7574_ /*12187*/;
assign _7578_ = _7167_ ^ _7574_ /*12190*/;
assign _7579_ = _7570_ & _7578_ /*12188*/;
assign _7391_ = _7570_ ^ _7578_ /*12189*/;
assign _7576_ = _7577_ | _7579_ /*12186*/;
assign _7581_ = ~Q[15] /*12185*/;
assign _7580_ = _7581_ & zeroWire /*12184*/;
assign _7582_ = _7168_ ^ _7580_ /*12182*/;
assign _7392_ = _7582_ ^ _7576_ /*12181*/;
assign _7621_ = ~D[0] /*12055*/;
assign _7618_ = R_0[14] & _7621_ /*12051*/;
assign _7619_ = R_0[14] ^ _7621_ /*12054*/;
assign _7620_ = oneWire & _7619_ /*12052*/;
assign _7585_ = oneWire ^ _7619_ /*12053*/;
assign _7617_ = _7618_ | _7620_ /*12050*/;
assign _7626_ = ~D[1] /*12049*/;
assign _7623_ = _7361_ & _7626_ /*12045*/;
assign _7624_ = _7361_ ^ _7626_ /*12048*/;
assign _7625_ = _7617_ & _7624_ /*12046*/;
assign _7586_ = _7617_ ^ _7624_ /*12047*/;
assign _7622_ = _7623_ | _7625_ /*12044*/;
assign _7631_ = ~D[2] /*12043*/;
assign _7628_ = _7362_ & _7631_ /*12039*/;
assign _7629_ = _7362_ ^ _7631_ /*12042*/;
assign _7630_ = _7622_ & _7629_ /*12040*/;
assign _7587_ = _7622_ ^ _7629_ /*12041*/;
assign _7627_ = _7628_ | _7630_ /*12038*/;
assign _7636_ = ~D[3] /*12037*/;
assign _7633_ = _7363_ & _7636_ /*12033*/;
assign _7634_ = _7363_ ^ _7636_ /*12036*/;
assign _7635_ = _7627_ & _7634_ /*12034*/;
assign _7588_ = _7627_ ^ _7634_ /*12035*/;
assign _7632_ = _7633_ | _7635_ /*12032*/;
assign _7641_ = ~D[4] /*12031*/;
assign _7638_ = _7364_ & _7641_ /*12027*/;
assign _7639_ = _7364_ ^ _7641_ /*12030*/;
assign _7640_ = _7632_ & _7639_ /*12028*/;
assign _7589_ = _7632_ ^ _7639_ /*12029*/;
assign _7637_ = _7638_ | _7640_ /*12026*/;
assign _7646_ = ~D[5] /*12025*/;
assign _7643_ = _7365_ & _7646_ /*12021*/;
assign _7644_ = _7365_ ^ _7646_ /*12024*/;
assign _7645_ = _7637_ & _7644_ /*12022*/;
assign _7590_ = _7637_ ^ _7644_ /*12023*/;
assign _7642_ = _7643_ | _7645_ /*12020*/;
assign _7651_ = ~D[6] /*12019*/;
assign _7648_ = _7366_ & _7651_ /*12015*/;
assign _7649_ = _7366_ ^ _7651_ /*12018*/;
assign _7650_ = _7642_ & _7649_ /*12016*/;
assign _7591_ = _7642_ ^ _7649_ /*12017*/;
assign _7647_ = _7648_ | _7650_ /*12014*/;
assign _7656_ = ~D[7] /*12013*/;
assign _7653_ = _7367_ & _7656_ /*12009*/;
assign _7654_ = _7367_ ^ _7656_ /*12012*/;
assign _7655_ = _7647_ & _7654_ /*12010*/;
assign _7592_ = _7647_ ^ _7654_ /*12011*/;
assign _7652_ = _7653_ | _7655_ /*12008*/;
assign _7661_ = ~D[8] /*12007*/;
assign _7658_ = _7368_ & _7661_ /*12003*/;
assign _7659_ = _7368_ ^ _7661_ /*12006*/;
assign _7660_ = _7652_ & _7659_ /*12004*/;
assign _7593_ = _7652_ ^ _7659_ /*12005*/;
assign _7657_ = _7658_ | _7660_ /*12002*/;
assign _7666_ = ~D[9] /*12001*/;
assign _7663_ = _7369_ & _7666_ /*11997*/;
assign _7664_ = _7369_ ^ _7666_ /*12000*/;
assign _7665_ = _7657_ & _7664_ /*11998*/;
assign _7594_ = _7657_ ^ _7664_ /*11999*/;
assign _7662_ = _7663_ | _7665_ /*11996*/;
assign _7671_ = ~D[10] /*11995*/;
assign _7668_ = _7370_ & _7671_ /*11991*/;
assign _7669_ = _7370_ ^ _7671_ /*11994*/;
assign _7670_ = _7662_ & _7669_ /*11992*/;
assign _7595_ = _7662_ ^ _7669_ /*11993*/;
assign _7667_ = _7668_ | _7670_ /*11990*/;
assign _7676_ = ~D[11] /*11989*/;
assign _7673_ = _7371_ & _7676_ /*11985*/;
assign _7674_ = _7371_ ^ _7676_ /*11988*/;
assign _7675_ = _7667_ & _7674_ /*11986*/;
assign _7596_ = _7667_ ^ _7674_ /*11987*/;
assign _7672_ = _7673_ | _7675_ /*11984*/;
assign _7681_ = ~D[12] /*11983*/;
assign _7678_ = _7372_ & _7681_ /*11979*/;
assign _7679_ = _7372_ ^ _7681_ /*11982*/;
assign _7680_ = _7672_ & _7679_ /*11980*/;
assign _7597_ = _7672_ ^ _7679_ /*11981*/;
assign _7677_ = _7678_ | _7680_ /*11978*/;
assign _7686_ = ~D[13] /*11977*/;
assign _7683_ = _7373_ & _7686_ /*11973*/;
assign _7684_ = _7373_ ^ _7686_ /*11976*/;
assign _7685_ = _7677_ & _7684_ /*11974*/;
assign _7598_ = _7677_ ^ _7684_ /*11975*/;
assign _7682_ = _7683_ | _7685_ /*11972*/;
assign _7691_ = ~D[14] /*11971*/;
assign _7688_ = _7374_ & _7691_ /*11967*/;
assign _7689_ = _7374_ ^ _7691_ /*11970*/;
assign _7690_ = _7682_ & _7689_ /*11968*/;
assign _7599_ = _7682_ ^ _7689_ /*11969*/;
assign _7687_ = _7688_ | _7690_ /*11966*/;
assign _7696_ = ~D[15] /*11965*/;
assign _7693_ = _7375_ & _7696_ /*11961*/;
assign _7694_ = _7375_ ^ _7696_ /*11964*/;
assign _7695_ = _7687_ & _7694_ /*11962*/;
assign _7600_ = _7687_ ^ _7694_ /*11963*/;
assign _7692_ = _7693_ | _7695_ /*11960*/;
assign _7701_ = ~D[16] /*11959*/;
assign _7698_ = _7376_ & _7701_ /*11955*/;
assign _7699_ = _7376_ ^ _7701_ /*11958*/;
assign _7700_ = _7692_ & _7699_ /*11956*/;
assign _7601_ = _7692_ ^ _7699_ /*11957*/;
assign _7697_ = _7698_ | _7700_ /*11954*/;
assign _7706_ = ~D[17] /*11953*/;
assign _7703_ = _7377_ & _7706_ /*11949*/;
assign _7704_ = _7377_ ^ _7706_ /*11952*/;
assign _7705_ = _7697_ & _7704_ /*11950*/;
assign _7602_ = _7697_ ^ _7704_ /*11951*/;
assign _7702_ = _7703_ | _7705_ /*11948*/;
assign _7711_ = ~D[18] /*11947*/;
assign _7708_ = _7378_ & _7711_ /*11943*/;
assign _7709_ = _7378_ ^ _7711_ /*11946*/;
assign _7710_ = _7702_ & _7709_ /*11944*/;
assign _7603_ = _7702_ ^ _7709_ /*11945*/;
assign _7707_ = _7708_ | _7710_ /*11942*/;
assign _7716_ = ~D[19] /*11941*/;
assign _7713_ = _7379_ & _7716_ /*11937*/;
assign _7714_ = _7379_ ^ _7716_ /*11940*/;
assign _7715_ = _7707_ & _7714_ /*11938*/;
assign _7604_ = _7707_ ^ _7714_ /*11939*/;
assign _7712_ = _7713_ | _7715_ /*11936*/;
assign _7721_ = ~D[20] /*11935*/;
assign _7718_ = _7380_ & _7721_ /*11931*/;
assign _7719_ = _7380_ ^ _7721_ /*11934*/;
assign _7720_ = _7712_ & _7719_ /*11932*/;
assign _7605_ = _7712_ ^ _7719_ /*11933*/;
assign _7717_ = _7718_ | _7720_ /*11930*/;
assign _7726_ = ~D[21] /*11929*/;
assign _7723_ = _7381_ & _7726_ /*11925*/;
assign _7724_ = _7381_ ^ _7726_ /*11928*/;
assign _7725_ = _7717_ & _7724_ /*11926*/;
assign _7606_ = _7717_ ^ _7724_ /*11927*/;
assign _7722_ = _7723_ | _7725_ /*11924*/;
assign _7731_ = ~D[22] /*11923*/;
assign _7728_ = _7382_ & _7731_ /*11919*/;
assign _7729_ = _7382_ ^ _7731_ /*11922*/;
assign _7730_ = _7722_ & _7729_ /*11920*/;
assign _7607_ = _7722_ ^ _7729_ /*11921*/;
assign _7727_ = _7728_ | _7730_ /*11918*/;
assign _7736_ = ~D[23] /*11917*/;
assign _7733_ = _7383_ & _7736_ /*11913*/;
assign _7734_ = _7383_ ^ _7736_ /*11916*/;
assign _7735_ = _7727_ & _7734_ /*11914*/;
assign _7608_ = _7727_ ^ _7734_ /*11915*/;
assign _7732_ = _7733_ | _7735_ /*11912*/;
assign _7741_ = ~D[24] /*11911*/;
assign _7738_ = _7384_ & _7741_ /*11907*/;
assign _7739_ = _7384_ ^ _7741_ /*11910*/;
assign _7740_ = _7732_ & _7739_ /*11908*/;
assign _7609_ = _7732_ ^ _7739_ /*11909*/;
assign _7737_ = _7738_ | _7740_ /*11906*/;
assign _7746_ = ~D[25] /*11905*/;
assign _7743_ = _7385_ & _7746_ /*11901*/;
assign _7744_ = _7385_ ^ _7746_ /*11904*/;
assign _7745_ = _7737_ & _7744_ /*11902*/;
assign _7610_ = _7737_ ^ _7744_ /*11903*/;
assign _7742_ = _7743_ | _7745_ /*11900*/;
assign _7751_ = ~D[26] /*11899*/;
assign _7748_ = _7386_ & _7751_ /*11895*/;
assign _7749_ = _7386_ ^ _7751_ /*11898*/;
assign _7750_ = _7742_ & _7749_ /*11896*/;
assign _7611_ = _7742_ ^ _7749_ /*11897*/;
assign _7747_ = _7748_ | _7750_ /*11894*/;
assign _7756_ = ~D[27] /*11893*/;
assign _7753_ = _7387_ & _7756_ /*11889*/;
assign _7754_ = _7387_ ^ _7756_ /*11892*/;
assign _7755_ = _7747_ & _7754_ /*11890*/;
assign _7612_ = _7747_ ^ _7754_ /*11891*/;
assign _7752_ = _7753_ | _7755_ /*11888*/;
assign _7761_ = ~D[28] /*11887*/;
assign _7758_ = _7388_ & _7761_ /*11883*/;
assign _7759_ = _7388_ ^ _7761_ /*11886*/;
assign _7760_ = _7752_ & _7759_ /*11884*/;
assign _7613_ = _7752_ ^ _7759_ /*11885*/;
assign _7757_ = _7758_ | _7760_ /*11882*/;
assign _7766_ = ~D[29] /*11881*/;
assign _7763_ = _7389_ & _7766_ /*11877*/;
assign _7764_ = _7389_ ^ _7766_ /*11880*/;
assign _7765_ = _7757_ & _7764_ /*11878*/;
assign _7614_ = _7757_ ^ _7764_ /*11879*/;
assign _7762_ = _7763_ | _7765_ /*11876*/;
assign _7771_ = ~D[30] /*11875*/;
assign _7768_ = _7390_ & _7771_ /*11871*/;
assign _7769_ = _7390_ ^ _7771_ /*11874*/;
assign _7770_ = _7762_ & _7769_ /*11872*/;
assign _7615_ = _7762_ ^ _7769_ /*11873*/;
assign _7767_ = _7768_ | _7770_ /*11870*/;
assign _7772_ = _7391_ & oneWire /*11865*/;
assign _7773_ = _7391_ ^ oneWire /*11868*/;
assign _7774_ = _7767_ & _7773_ /*11866*/;
assign _7616_ = _7767_ ^ _7773_ /*11867*/;
assign Q[14] = _7772_ | _7774_ /*11864*/;
assign _7843_ = ~Q[14] /*11671*/;
assign _7842_ = _7843_ & D[0] /*11670*/;
assign _7845_ = _7585_ & _7842_ /*11665*/;
assign _7846_ = _7585_ ^ _7842_ /*11668*/;
assign _7847_ = zeroWire & _7846_ /*11666*/;
assign _7809_ = zeroWire ^ _7846_ /*11667*/;
assign _7844_ = _7845_ | _7847_ /*11664*/;
assign _7849_ = ~Q[14] /*11663*/;
assign _7848_ = _7849_ & D[1] /*11662*/;
assign _7851_ = _7586_ & _7848_ /*11657*/;
assign _7852_ = _7586_ ^ _7848_ /*11660*/;
assign _7853_ = _7844_ & _7852_ /*11658*/;
assign _7810_ = _7844_ ^ _7852_ /*11659*/;
assign _7850_ = _7851_ | _7853_ /*11656*/;
assign _7855_ = ~Q[14] /*11655*/;
assign _7854_ = _7855_ & D[2] /*11654*/;
assign _7857_ = _7587_ & _7854_ /*11649*/;
assign _7858_ = _7587_ ^ _7854_ /*11652*/;
assign _7859_ = _7850_ & _7858_ /*11650*/;
assign _7811_ = _7850_ ^ _7858_ /*11651*/;
assign _7856_ = _7857_ | _7859_ /*11648*/;
assign _7861_ = ~Q[14] /*11647*/;
assign _7860_ = _7861_ & D[3] /*11646*/;
assign _7863_ = _7588_ & _7860_ /*11641*/;
assign _7864_ = _7588_ ^ _7860_ /*11644*/;
assign _7865_ = _7856_ & _7864_ /*11642*/;
assign _7812_ = _7856_ ^ _7864_ /*11643*/;
assign _7862_ = _7863_ | _7865_ /*11640*/;
assign _7867_ = ~Q[14] /*11639*/;
assign _7866_ = _7867_ & D[4] /*11638*/;
assign _7869_ = _7589_ & _7866_ /*11633*/;
assign _7870_ = _7589_ ^ _7866_ /*11636*/;
assign _7871_ = _7862_ & _7870_ /*11634*/;
assign _7813_ = _7862_ ^ _7870_ /*11635*/;
assign _7868_ = _7869_ | _7871_ /*11632*/;
assign _7873_ = ~Q[14] /*11631*/;
assign _7872_ = _7873_ & D[5] /*11630*/;
assign _7875_ = _7590_ & _7872_ /*11625*/;
assign _7876_ = _7590_ ^ _7872_ /*11628*/;
assign _7877_ = _7868_ & _7876_ /*11626*/;
assign _7814_ = _7868_ ^ _7876_ /*11627*/;
assign _7874_ = _7875_ | _7877_ /*11624*/;
assign _7879_ = ~Q[14] /*11623*/;
assign _7878_ = _7879_ & D[6] /*11622*/;
assign _7881_ = _7591_ & _7878_ /*11617*/;
assign _7882_ = _7591_ ^ _7878_ /*11620*/;
assign _7883_ = _7874_ & _7882_ /*11618*/;
assign _7815_ = _7874_ ^ _7882_ /*11619*/;
assign _7880_ = _7881_ | _7883_ /*11616*/;
assign _7885_ = ~Q[14] /*11615*/;
assign _7884_ = _7885_ & D[7] /*11614*/;
assign _7887_ = _7592_ & _7884_ /*11609*/;
assign _7888_ = _7592_ ^ _7884_ /*11612*/;
assign _7889_ = _7880_ & _7888_ /*11610*/;
assign _7816_ = _7880_ ^ _7888_ /*11611*/;
assign _7886_ = _7887_ | _7889_ /*11608*/;
assign _7891_ = ~Q[14] /*11607*/;
assign _7890_ = _7891_ & D[8] /*11606*/;
assign _7893_ = _7593_ & _7890_ /*11601*/;
assign _7894_ = _7593_ ^ _7890_ /*11604*/;
assign _7895_ = _7886_ & _7894_ /*11602*/;
assign _7817_ = _7886_ ^ _7894_ /*11603*/;
assign _7892_ = _7893_ | _7895_ /*11600*/;
assign _7897_ = ~Q[14] /*11599*/;
assign _7896_ = _7897_ & D[9] /*11598*/;
assign _7899_ = _7594_ & _7896_ /*11593*/;
assign _7900_ = _7594_ ^ _7896_ /*11596*/;
assign _7901_ = _7892_ & _7900_ /*11594*/;
assign _7818_ = _7892_ ^ _7900_ /*11595*/;
assign _7898_ = _7899_ | _7901_ /*11592*/;
assign _7903_ = ~Q[14] /*11591*/;
assign _7902_ = _7903_ & D[10] /*11590*/;
assign _7905_ = _7595_ & _7902_ /*11585*/;
assign _7906_ = _7595_ ^ _7902_ /*11588*/;
assign _7907_ = _7898_ & _7906_ /*11586*/;
assign _7819_ = _7898_ ^ _7906_ /*11587*/;
assign _7904_ = _7905_ | _7907_ /*11584*/;
assign _7909_ = ~Q[14] /*11583*/;
assign _7908_ = _7909_ & D[11] /*11582*/;
assign _7911_ = _7596_ & _7908_ /*11577*/;
assign _7912_ = _7596_ ^ _7908_ /*11580*/;
assign _7913_ = _7904_ & _7912_ /*11578*/;
assign _7820_ = _7904_ ^ _7912_ /*11579*/;
assign _7910_ = _7911_ | _7913_ /*11576*/;
assign _7915_ = ~Q[14] /*11575*/;
assign _7914_ = _7915_ & D[12] /*11574*/;
assign _7917_ = _7597_ & _7914_ /*11569*/;
assign _7918_ = _7597_ ^ _7914_ /*11572*/;
assign _7919_ = _7910_ & _7918_ /*11570*/;
assign _7821_ = _7910_ ^ _7918_ /*11571*/;
assign _7916_ = _7917_ | _7919_ /*11568*/;
assign _7921_ = ~Q[14] /*11567*/;
assign _7920_ = _7921_ & D[13] /*11566*/;
assign _7923_ = _7598_ & _7920_ /*11561*/;
assign _7924_ = _7598_ ^ _7920_ /*11564*/;
assign _7925_ = _7916_ & _7924_ /*11562*/;
assign _7822_ = _7916_ ^ _7924_ /*11563*/;
assign _7922_ = _7923_ | _7925_ /*11560*/;
assign _7927_ = ~Q[14] /*11559*/;
assign _7926_ = _7927_ & D[14] /*11558*/;
assign _7929_ = _7599_ & _7926_ /*11553*/;
assign _7930_ = _7599_ ^ _7926_ /*11556*/;
assign _7931_ = _7922_ & _7930_ /*11554*/;
assign _7823_ = _7922_ ^ _7930_ /*11555*/;
assign _7928_ = _7929_ | _7931_ /*11552*/;
assign _7933_ = ~Q[14] /*11551*/;
assign _7932_ = _7933_ & D[15] /*11550*/;
assign _7935_ = _7600_ & _7932_ /*11545*/;
assign _7936_ = _7600_ ^ _7932_ /*11548*/;
assign _7937_ = _7928_ & _7936_ /*11546*/;
assign _7824_ = _7928_ ^ _7936_ /*11547*/;
assign _7934_ = _7935_ | _7937_ /*11544*/;
assign _7939_ = ~Q[14] /*11543*/;
assign _7938_ = _7939_ & D[16] /*11542*/;
assign _7941_ = _7601_ & _7938_ /*11537*/;
assign _7942_ = _7601_ ^ _7938_ /*11540*/;
assign _7943_ = _7934_ & _7942_ /*11538*/;
assign _7825_ = _7934_ ^ _7942_ /*11539*/;
assign _7940_ = _7941_ | _7943_ /*11536*/;
assign _7945_ = ~Q[14] /*11535*/;
assign _7944_ = _7945_ & D[17] /*11534*/;
assign _7947_ = _7602_ & _7944_ /*11529*/;
assign _7948_ = _7602_ ^ _7944_ /*11532*/;
assign _7949_ = _7940_ & _7948_ /*11530*/;
assign _7826_ = _7940_ ^ _7948_ /*11531*/;
assign _7946_ = _7947_ | _7949_ /*11528*/;
assign _7951_ = ~Q[14] /*11527*/;
assign _7950_ = _7951_ & D[18] /*11526*/;
assign _7953_ = _7603_ & _7950_ /*11521*/;
assign _7954_ = _7603_ ^ _7950_ /*11524*/;
assign _7955_ = _7946_ & _7954_ /*11522*/;
assign _7827_ = _7946_ ^ _7954_ /*11523*/;
assign _7952_ = _7953_ | _7955_ /*11520*/;
assign _7957_ = ~Q[14] /*11519*/;
assign _7956_ = _7957_ & D[19] /*11518*/;
assign _7959_ = _7604_ & _7956_ /*11513*/;
assign _7960_ = _7604_ ^ _7956_ /*11516*/;
assign _7961_ = _7952_ & _7960_ /*11514*/;
assign _7828_ = _7952_ ^ _7960_ /*11515*/;
assign _7958_ = _7959_ | _7961_ /*11512*/;
assign _7963_ = ~Q[14] /*11511*/;
assign _7962_ = _7963_ & D[20] /*11510*/;
assign _7965_ = _7605_ & _7962_ /*11505*/;
assign _7966_ = _7605_ ^ _7962_ /*11508*/;
assign _7967_ = _7958_ & _7966_ /*11506*/;
assign _7829_ = _7958_ ^ _7966_ /*11507*/;
assign _7964_ = _7965_ | _7967_ /*11504*/;
assign _7969_ = ~Q[14] /*11503*/;
assign _7968_ = _7969_ & D[21] /*11502*/;
assign _7971_ = _7606_ & _7968_ /*11497*/;
assign _7972_ = _7606_ ^ _7968_ /*11500*/;
assign _7973_ = _7964_ & _7972_ /*11498*/;
assign _7830_ = _7964_ ^ _7972_ /*11499*/;
assign _7970_ = _7971_ | _7973_ /*11496*/;
assign _7975_ = ~Q[14] /*11495*/;
assign _7974_ = _7975_ & D[22] /*11494*/;
assign _7977_ = _7607_ & _7974_ /*11489*/;
assign _7978_ = _7607_ ^ _7974_ /*11492*/;
assign _7979_ = _7970_ & _7978_ /*11490*/;
assign _7831_ = _7970_ ^ _7978_ /*11491*/;
assign _7976_ = _7977_ | _7979_ /*11488*/;
assign _7981_ = ~Q[14] /*11487*/;
assign _7980_ = _7981_ & D[23] /*11486*/;
assign _7983_ = _7608_ & _7980_ /*11481*/;
assign _7984_ = _7608_ ^ _7980_ /*11484*/;
assign _7985_ = _7976_ & _7984_ /*11482*/;
assign _7832_ = _7976_ ^ _7984_ /*11483*/;
assign _7982_ = _7983_ | _7985_ /*11480*/;
assign _7987_ = ~Q[14] /*11479*/;
assign _7986_ = _7987_ & D[24] /*11478*/;
assign _7989_ = _7609_ & _7986_ /*11473*/;
assign _7990_ = _7609_ ^ _7986_ /*11476*/;
assign _7991_ = _7982_ & _7990_ /*11474*/;
assign _7833_ = _7982_ ^ _7990_ /*11475*/;
assign _7988_ = _7989_ | _7991_ /*11472*/;
assign _7993_ = ~Q[14] /*11471*/;
assign _7992_ = _7993_ & D[25] /*11470*/;
assign _7995_ = _7610_ & _7992_ /*11465*/;
assign _7996_ = _7610_ ^ _7992_ /*11468*/;
assign _7997_ = _7988_ & _7996_ /*11466*/;
assign _7834_ = _7988_ ^ _7996_ /*11467*/;
assign _7994_ = _7995_ | _7997_ /*11464*/;
assign _7999_ = ~Q[14] /*11463*/;
assign _7998_ = _7999_ & D[26] /*11462*/;
assign _8001_ = _7611_ & _7998_ /*11457*/;
assign _8002_ = _7611_ ^ _7998_ /*11460*/;
assign _8003_ = _7994_ & _8002_ /*11458*/;
assign _7835_ = _7994_ ^ _8002_ /*11459*/;
assign _8000_ = _8001_ | _8003_ /*11456*/;
assign _8005_ = ~Q[14] /*11455*/;
assign _8004_ = _8005_ & D[27] /*11454*/;
assign _8007_ = _7612_ & _8004_ /*11449*/;
assign _8008_ = _7612_ ^ _8004_ /*11452*/;
assign _8009_ = _8000_ & _8008_ /*11450*/;
assign _7836_ = _8000_ ^ _8008_ /*11451*/;
assign _8006_ = _8007_ | _8009_ /*11448*/;
assign _8011_ = ~Q[14] /*11447*/;
assign _8010_ = _8011_ & D[28] /*11446*/;
assign _8013_ = _7613_ & _8010_ /*11441*/;
assign _8014_ = _7613_ ^ _8010_ /*11444*/;
assign _8015_ = _8006_ & _8014_ /*11442*/;
assign _7837_ = _8006_ ^ _8014_ /*11443*/;
assign _8012_ = _8013_ | _8015_ /*11440*/;
assign _8017_ = ~Q[14] /*11439*/;
assign _8016_ = _8017_ & D[29] /*11438*/;
assign _8019_ = _7614_ & _8016_ /*11433*/;
assign _8020_ = _7614_ ^ _8016_ /*11436*/;
assign _8021_ = _8012_ & _8020_ /*11434*/;
assign _7838_ = _8012_ ^ _8020_ /*11435*/;
assign _8018_ = _8019_ | _8021_ /*11432*/;
assign _8023_ = ~Q[14] /*11431*/;
assign _8022_ = _8023_ & D[30] /*11430*/;
assign _8025_ = _7615_ & _8022_ /*11425*/;
assign _8026_ = _7615_ ^ _8022_ /*11428*/;
assign _8027_ = _8018_ & _8026_ /*11426*/;
assign _7839_ = _8018_ ^ _8026_ /*11427*/;
assign _8024_ = _8025_ | _8027_ /*11424*/;
assign _8029_ = ~Q[14] /*11423*/;
assign _8028_ = _8029_ & zeroWire /*11422*/;
assign _8030_ = _7616_ ^ _8028_ /*11420*/;
assign _7840_ = _8030_ ^ _8024_ /*11419*/;
assign _8069_ = ~D[0] /*11293*/;
assign _8066_ = R_0[13] & _8069_ /*11289*/;
assign _8067_ = R_0[13] ^ _8069_ /*11292*/;
assign _8068_ = oneWire & _8067_ /*11290*/;
assign _8033_ = oneWire ^ _8067_ /*11291*/;
assign _8065_ = _8066_ | _8068_ /*11288*/;
assign _8074_ = ~D[1] /*11287*/;
assign _8071_ = _7809_ & _8074_ /*11283*/;
assign _8072_ = _7809_ ^ _8074_ /*11286*/;
assign _8073_ = _8065_ & _8072_ /*11284*/;
assign _8034_ = _8065_ ^ _8072_ /*11285*/;
assign _8070_ = _8071_ | _8073_ /*11282*/;
assign _8079_ = ~D[2] /*11281*/;
assign _8076_ = _7810_ & _8079_ /*11277*/;
assign _8077_ = _7810_ ^ _8079_ /*11280*/;
assign _8078_ = _8070_ & _8077_ /*11278*/;
assign _8035_ = _8070_ ^ _8077_ /*11279*/;
assign _8075_ = _8076_ | _8078_ /*11276*/;
assign _8084_ = ~D[3] /*11275*/;
assign _8081_ = _7811_ & _8084_ /*11271*/;
assign _8082_ = _7811_ ^ _8084_ /*11274*/;
assign _8083_ = _8075_ & _8082_ /*11272*/;
assign _8036_ = _8075_ ^ _8082_ /*11273*/;
assign _8080_ = _8081_ | _8083_ /*11270*/;
assign _8089_ = ~D[4] /*11269*/;
assign _8086_ = _7812_ & _8089_ /*11265*/;
assign _8087_ = _7812_ ^ _8089_ /*11268*/;
assign _8088_ = _8080_ & _8087_ /*11266*/;
assign _8037_ = _8080_ ^ _8087_ /*11267*/;
assign _8085_ = _8086_ | _8088_ /*11264*/;
assign _8094_ = ~D[5] /*11263*/;
assign _8091_ = _7813_ & _8094_ /*11259*/;
assign _8092_ = _7813_ ^ _8094_ /*11262*/;
assign _8093_ = _8085_ & _8092_ /*11260*/;
assign _8038_ = _8085_ ^ _8092_ /*11261*/;
assign _8090_ = _8091_ | _8093_ /*11258*/;
assign _8099_ = ~D[6] /*11257*/;
assign _8096_ = _7814_ & _8099_ /*11253*/;
assign _8097_ = _7814_ ^ _8099_ /*11256*/;
assign _8098_ = _8090_ & _8097_ /*11254*/;
assign _8039_ = _8090_ ^ _8097_ /*11255*/;
assign _8095_ = _8096_ | _8098_ /*11252*/;
assign _8104_ = ~D[7] /*11251*/;
assign _8101_ = _7815_ & _8104_ /*11247*/;
assign _8102_ = _7815_ ^ _8104_ /*11250*/;
assign _8103_ = _8095_ & _8102_ /*11248*/;
assign _8040_ = _8095_ ^ _8102_ /*11249*/;
assign _8100_ = _8101_ | _8103_ /*11246*/;
assign _8109_ = ~D[8] /*11245*/;
assign _8106_ = _7816_ & _8109_ /*11241*/;
assign _8107_ = _7816_ ^ _8109_ /*11244*/;
assign _8108_ = _8100_ & _8107_ /*11242*/;
assign _8041_ = _8100_ ^ _8107_ /*11243*/;
assign _8105_ = _8106_ | _8108_ /*11240*/;
assign _8114_ = ~D[9] /*11239*/;
assign _8111_ = _7817_ & _8114_ /*11235*/;
assign _8112_ = _7817_ ^ _8114_ /*11238*/;
assign _8113_ = _8105_ & _8112_ /*11236*/;
assign _8042_ = _8105_ ^ _8112_ /*11237*/;
assign _8110_ = _8111_ | _8113_ /*11234*/;
assign _8119_ = ~D[10] /*11233*/;
assign _8116_ = _7818_ & _8119_ /*11229*/;
assign _8117_ = _7818_ ^ _8119_ /*11232*/;
assign _8118_ = _8110_ & _8117_ /*11230*/;
assign _8043_ = _8110_ ^ _8117_ /*11231*/;
assign _8115_ = _8116_ | _8118_ /*11228*/;
assign _8124_ = ~D[11] /*11227*/;
assign _8121_ = _7819_ & _8124_ /*11223*/;
assign _8122_ = _7819_ ^ _8124_ /*11226*/;
assign _8123_ = _8115_ & _8122_ /*11224*/;
assign _8044_ = _8115_ ^ _8122_ /*11225*/;
assign _8120_ = _8121_ | _8123_ /*11222*/;
assign _8129_ = ~D[12] /*11221*/;
assign _8126_ = _7820_ & _8129_ /*11217*/;
assign _8127_ = _7820_ ^ _8129_ /*11220*/;
assign _8128_ = _8120_ & _8127_ /*11218*/;
assign _8045_ = _8120_ ^ _8127_ /*11219*/;
assign _8125_ = _8126_ | _8128_ /*11216*/;
assign _8134_ = ~D[13] /*11215*/;
assign _8131_ = _7821_ & _8134_ /*11211*/;
assign _8132_ = _7821_ ^ _8134_ /*11214*/;
assign _8133_ = _8125_ & _8132_ /*11212*/;
assign _8046_ = _8125_ ^ _8132_ /*11213*/;
assign _8130_ = _8131_ | _8133_ /*11210*/;
assign _8139_ = ~D[14] /*11209*/;
assign _8136_ = _7822_ & _8139_ /*11205*/;
assign _8137_ = _7822_ ^ _8139_ /*11208*/;
assign _8138_ = _8130_ & _8137_ /*11206*/;
assign _8047_ = _8130_ ^ _8137_ /*11207*/;
assign _8135_ = _8136_ | _8138_ /*11204*/;
assign _8144_ = ~D[15] /*11203*/;
assign _8141_ = _7823_ & _8144_ /*11199*/;
assign _8142_ = _7823_ ^ _8144_ /*11202*/;
assign _8143_ = _8135_ & _8142_ /*11200*/;
assign _8048_ = _8135_ ^ _8142_ /*11201*/;
assign _8140_ = _8141_ | _8143_ /*11198*/;
assign _8149_ = ~D[16] /*11197*/;
assign _8146_ = _7824_ & _8149_ /*11193*/;
assign _8147_ = _7824_ ^ _8149_ /*11196*/;
assign _8148_ = _8140_ & _8147_ /*11194*/;
assign _8049_ = _8140_ ^ _8147_ /*11195*/;
assign _8145_ = _8146_ | _8148_ /*11192*/;
assign _8154_ = ~D[17] /*11191*/;
assign _8151_ = _7825_ & _8154_ /*11187*/;
assign _8152_ = _7825_ ^ _8154_ /*11190*/;
assign _8153_ = _8145_ & _8152_ /*11188*/;
assign _8050_ = _8145_ ^ _8152_ /*11189*/;
assign _8150_ = _8151_ | _8153_ /*11186*/;
assign _8159_ = ~D[18] /*11185*/;
assign _8156_ = _7826_ & _8159_ /*11181*/;
assign _8157_ = _7826_ ^ _8159_ /*11184*/;
assign _8158_ = _8150_ & _8157_ /*11182*/;
assign _8051_ = _8150_ ^ _8157_ /*11183*/;
assign _8155_ = _8156_ | _8158_ /*11180*/;
assign _8164_ = ~D[19] /*11179*/;
assign _8161_ = _7827_ & _8164_ /*11175*/;
assign _8162_ = _7827_ ^ _8164_ /*11178*/;
assign _8163_ = _8155_ & _8162_ /*11176*/;
assign _8052_ = _8155_ ^ _8162_ /*11177*/;
assign _8160_ = _8161_ | _8163_ /*11174*/;
assign _8169_ = ~D[20] /*11173*/;
assign _8166_ = _7828_ & _8169_ /*11169*/;
assign _8167_ = _7828_ ^ _8169_ /*11172*/;
assign _8168_ = _8160_ & _8167_ /*11170*/;
assign _8053_ = _8160_ ^ _8167_ /*11171*/;
assign _8165_ = _8166_ | _8168_ /*11168*/;
assign _8174_ = ~D[21] /*11167*/;
assign _8171_ = _7829_ & _8174_ /*11163*/;
assign _8172_ = _7829_ ^ _8174_ /*11166*/;
assign _8173_ = _8165_ & _8172_ /*11164*/;
assign _8054_ = _8165_ ^ _8172_ /*11165*/;
assign _8170_ = _8171_ | _8173_ /*11162*/;
assign _8179_ = ~D[22] /*11161*/;
assign _8176_ = _7830_ & _8179_ /*11157*/;
assign _8177_ = _7830_ ^ _8179_ /*11160*/;
assign _8178_ = _8170_ & _8177_ /*11158*/;
assign _8055_ = _8170_ ^ _8177_ /*11159*/;
assign _8175_ = _8176_ | _8178_ /*11156*/;
assign _8184_ = ~D[23] /*11155*/;
assign _8181_ = _7831_ & _8184_ /*11151*/;
assign _8182_ = _7831_ ^ _8184_ /*11154*/;
assign _8183_ = _8175_ & _8182_ /*11152*/;
assign _8056_ = _8175_ ^ _8182_ /*11153*/;
assign _8180_ = _8181_ | _8183_ /*11150*/;
assign _8189_ = ~D[24] /*11149*/;
assign _8186_ = _7832_ & _8189_ /*11145*/;
assign _8187_ = _7832_ ^ _8189_ /*11148*/;
assign _8188_ = _8180_ & _8187_ /*11146*/;
assign _8057_ = _8180_ ^ _8187_ /*11147*/;
assign _8185_ = _8186_ | _8188_ /*11144*/;
assign _8194_ = ~D[25] /*11143*/;
assign _8191_ = _7833_ & _8194_ /*11139*/;
assign _8192_ = _7833_ ^ _8194_ /*11142*/;
assign _8193_ = _8185_ & _8192_ /*11140*/;
assign _8058_ = _8185_ ^ _8192_ /*11141*/;
assign _8190_ = _8191_ | _8193_ /*11138*/;
assign _8199_ = ~D[26] /*11137*/;
assign _8196_ = _7834_ & _8199_ /*11133*/;
assign _8197_ = _7834_ ^ _8199_ /*11136*/;
assign _8198_ = _8190_ & _8197_ /*11134*/;
assign _8059_ = _8190_ ^ _8197_ /*11135*/;
assign _8195_ = _8196_ | _8198_ /*11132*/;
assign _8204_ = ~D[27] /*11131*/;
assign _8201_ = _7835_ & _8204_ /*11127*/;
assign _8202_ = _7835_ ^ _8204_ /*11130*/;
assign _8203_ = _8195_ & _8202_ /*11128*/;
assign _8060_ = _8195_ ^ _8202_ /*11129*/;
assign _8200_ = _8201_ | _8203_ /*11126*/;
assign _8209_ = ~D[28] /*11125*/;
assign _8206_ = _7836_ & _8209_ /*11121*/;
assign _8207_ = _7836_ ^ _8209_ /*11124*/;
assign _8208_ = _8200_ & _8207_ /*11122*/;
assign _8061_ = _8200_ ^ _8207_ /*11123*/;
assign _8205_ = _8206_ | _8208_ /*11120*/;
assign _8214_ = ~D[29] /*11119*/;
assign _8211_ = _7837_ & _8214_ /*11115*/;
assign _8212_ = _7837_ ^ _8214_ /*11118*/;
assign _8213_ = _8205_ & _8212_ /*11116*/;
assign _8062_ = _8205_ ^ _8212_ /*11117*/;
assign _8210_ = _8211_ | _8213_ /*11114*/;
assign _8219_ = ~D[30] /*11113*/;
assign _8216_ = _7838_ & _8219_ /*11109*/;
assign _8217_ = _7838_ ^ _8219_ /*11112*/;
assign _8218_ = _8210_ & _8217_ /*11110*/;
assign _8063_ = _8210_ ^ _8217_ /*11111*/;
assign _8215_ = _8216_ | _8218_ /*11108*/;
assign _8220_ = _7839_ & oneWire /*11103*/;
assign _8221_ = _7839_ ^ oneWire /*11106*/;
assign _8222_ = _8215_ & _8221_ /*11104*/;
assign _8064_ = _8215_ ^ _8221_ /*11105*/;
assign Q[13] = _8220_ | _8222_ /*11102*/;
assign _8291_ = ~Q[13] /*10909*/;
assign _8290_ = _8291_ & D[0] /*10908*/;
assign _8293_ = _8033_ & _8290_ /*10903*/;
assign _8294_ = _8033_ ^ _8290_ /*10906*/;
assign _8295_ = zeroWire & _8294_ /*10904*/;
assign _8257_ = zeroWire ^ _8294_ /*10905*/;
assign _8292_ = _8293_ | _8295_ /*10902*/;
assign _8297_ = ~Q[13] /*10901*/;
assign _8296_ = _8297_ & D[1] /*10900*/;
assign _8299_ = _8034_ & _8296_ /*10895*/;
assign _8300_ = _8034_ ^ _8296_ /*10898*/;
assign _8301_ = _8292_ & _8300_ /*10896*/;
assign _8258_ = _8292_ ^ _8300_ /*10897*/;
assign _8298_ = _8299_ | _8301_ /*10894*/;
assign _8303_ = ~Q[13] /*10893*/;
assign _8302_ = _8303_ & D[2] /*10892*/;
assign _8305_ = _8035_ & _8302_ /*10887*/;
assign _8306_ = _8035_ ^ _8302_ /*10890*/;
assign _8307_ = _8298_ & _8306_ /*10888*/;
assign _8259_ = _8298_ ^ _8306_ /*10889*/;
assign _8304_ = _8305_ | _8307_ /*10886*/;
assign _8309_ = ~Q[13] /*10885*/;
assign _8308_ = _8309_ & D[3] /*10884*/;
assign _8311_ = _8036_ & _8308_ /*10879*/;
assign _8312_ = _8036_ ^ _8308_ /*10882*/;
assign _8313_ = _8304_ & _8312_ /*10880*/;
assign _8260_ = _8304_ ^ _8312_ /*10881*/;
assign _8310_ = _8311_ | _8313_ /*10878*/;
assign _8315_ = ~Q[13] /*10877*/;
assign _8314_ = _8315_ & D[4] /*10876*/;
assign _8317_ = _8037_ & _8314_ /*10871*/;
assign _8318_ = _8037_ ^ _8314_ /*10874*/;
assign _8319_ = _8310_ & _8318_ /*10872*/;
assign _8261_ = _8310_ ^ _8318_ /*10873*/;
assign _8316_ = _8317_ | _8319_ /*10870*/;
assign _8321_ = ~Q[13] /*10869*/;
assign _8320_ = _8321_ & D[5] /*10868*/;
assign _8323_ = _8038_ & _8320_ /*10863*/;
assign _8324_ = _8038_ ^ _8320_ /*10866*/;
assign _8325_ = _8316_ & _8324_ /*10864*/;
assign _8262_ = _8316_ ^ _8324_ /*10865*/;
assign _8322_ = _8323_ | _8325_ /*10862*/;
assign _8327_ = ~Q[13] /*10861*/;
assign _8326_ = _8327_ & D[6] /*10860*/;
assign _8329_ = _8039_ & _8326_ /*10855*/;
assign _8330_ = _8039_ ^ _8326_ /*10858*/;
assign _8331_ = _8322_ & _8330_ /*10856*/;
assign _8263_ = _8322_ ^ _8330_ /*10857*/;
assign _8328_ = _8329_ | _8331_ /*10854*/;
assign _8333_ = ~Q[13] /*10853*/;
assign _8332_ = _8333_ & D[7] /*10852*/;
assign _8335_ = _8040_ & _8332_ /*10847*/;
assign _8336_ = _8040_ ^ _8332_ /*10850*/;
assign _8337_ = _8328_ & _8336_ /*10848*/;
assign _8264_ = _8328_ ^ _8336_ /*10849*/;
assign _8334_ = _8335_ | _8337_ /*10846*/;
assign _8339_ = ~Q[13] /*10845*/;
assign _8338_ = _8339_ & D[8] /*10844*/;
assign _8341_ = _8041_ & _8338_ /*10839*/;
assign _8342_ = _8041_ ^ _8338_ /*10842*/;
assign _8343_ = _8334_ & _8342_ /*10840*/;
assign _8265_ = _8334_ ^ _8342_ /*10841*/;
assign _8340_ = _8341_ | _8343_ /*10838*/;
assign _8345_ = ~Q[13] /*10837*/;
assign _8344_ = _8345_ & D[9] /*10836*/;
assign _8347_ = _8042_ & _8344_ /*10831*/;
assign _8348_ = _8042_ ^ _8344_ /*10834*/;
assign _8349_ = _8340_ & _8348_ /*10832*/;
assign _8266_ = _8340_ ^ _8348_ /*10833*/;
assign _8346_ = _8347_ | _8349_ /*10830*/;
assign _8351_ = ~Q[13] /*10829*/;
assign _8350_ = _8351_ & D[10] /*10828*/;
assign _8353_ = _8043_ & _8350_ /*10823*/;
assign _8354_ = _8043_ ^ _8350_ /*10826*/;
assign _8355_ = _8346_ & _8354_ /*10824*/;
assign _8267_ = _8346_ ^ _8354_ /*10825*/;
assign _8352_ = _8353_ | _8355_ /*10822*/;
assign _8357_ = ~Q[13] /*10821*/;
assign _8356_ = _8357_ & D[11] /*10820*/;
assign _8359_ = _8044_ & _8356_ /*10815*/;
assign _8360_ = _8044_ ^ _8356_ /*10818*/;
assign _8361_ = _8352_ & _8360_ /*10816*/;
assign _8268_ = _8352_ ^ _8360_ /*10817*/;
assign _8358_ = _8359_ | _8361_ /*10814*/;
assign _8363_ = ~Q[13] /*10813*/;
assign _8362_ = _8363_ & D[12] /*10812*/;
assign _8365_ = _8045_ & _8362_ /*10807*/;
assign _8366_ = _8045_ ^ _8362_ /*10810*/;
assign _8367_ = _8358_ & _8366_ /*10808*/;
assign _8269_ = _8358_ ^ _8366_ /*10809*/;
assign _8364_ = _8365_ | _8367_ /*10806*/;
assign _8369_ = ~Q[13] /*10805*/;
assign _8368_ = _8369_ & D[13] /*10804*/;
assign _8371_ = _8046_ & _8368_ /*10799*/;
assign _8372_ = _8046_ ^ _8368_ /*10802*/;
assign _8373_ = _8364_ & _8372_ /*10800*/;
assign _8270_ = _8364_ ^ _8372_ /*10801*/;
assign _8370_ = _8371_ | _8373_ /*10798*/;
assign _8375_ = ~Q[13] /*10797*/;
assign _8374_ = _8375_ & D[14] /*10796*/;
assign _8377_ = _8047_ & _8374_ /*10791*/;
assign _8378_ = _8047_ ^ _8374_ /*10794*/;
assign _8379_ = _8370_ & _8378_ /*10792*/;
assign _8271_ = _8370_ ^ _8378_ /*10793*/;
assign _8376_ = _8377_ | _8379_ /*10790*/;
assign _8381_ = ~Q[13] /*10789*/;
assign _8380_ = _8381_ & D[15] /*10788*/;
assign _8383_ = _8048_ & _8380_ /*10783*/;
assign _8384_ = _8048_ ^ _8380_ /*10786*/;
assign _8385_ = _8376_ & _8384_ /*10784*/;
assign _8272_ = _8376_ ^ _8384_ /*10785*/;
assign _8382_ = _8383_ | _8385_ /*10782*/;
assign _8387_ = ~Q[13] /*10781*/;
assign _8386_ = _8387_ & D[16] /*10780*/;
assign _8389_ = _8049_ & _8386_ /*10775*/;
assign _8390_ = _8049_ ^ _8386_ /*10778*/;
assign _8391_ = _8382_ & _8390_ /*10776*/;
assign _8273_ = _8382_ ^ _8390_ /*10777*/;
assign _8388_ = _8389_ | _8391_ /*10774*/;
assign _8393_ = ~Q[13] /*10773*/;
assign _8392_ = _8393_ & D[17] /*10772*/;
assign _8395_ = _8050_ & _8392_ /*10767*/;
assign _8396_ = _8050_ ^ _8392_ /*10770*/;
assign _8397_ = _8388_ & _8396_ /*10768*/;
assign _8274_ = _8388_ ^ _8396_ /*10769*/;
assign _8394_ = _8395_ | _8397_ /*10766*/;
assign _8399_ = ~Q[13] /*10765*/;
assign _8398_ = _8399_ & D[18] /*10764*/;
assign _8401_ = _8051_ & _8398_ /*10759*/;
assign _8402_ = _8051_ ^ _8398_ /*10762*/;
assign _8403_ = _8394_ & _8402_ /*10760*/;
assign _8275_ = _8394_ ^ _8402_ /*10761*/;
assign _8400_ = _8401_ | _8403_ /*10758*/;
assign _8405_ = ~Q[13] /*10757*/;
assign _8404_ = _8405_ & D[19] /*10756*/;
assign _8407_ = _8052_ & _8404_ /*10751*/;
assign _8408_ = _8052_ ^ _8404_ /*10754*/;
assign _8409_ = _8400_ & _8408_ /*10752*/;
assign _8276_ = _8400_ ^ _8408_ /*10753*/;
assign _8406_ = _8407_ | _8409_ /*10750*/;
assign _8411_ = ~Q[13] /*10749*/;
assign _8410_ = _8411_ & D[20] /*10748*/;
assign _8413_ = _8053_ & _8410_ /*10743*/;
assign _8414_ = _8053_ ^ _8410_ /*10746*/;
assign _8415_ = _8406_ & _8414_ /*10744*/;
assign _8277_ = _8406_ ^ _8414_ /*10745*/;
assign _8412_ = _8413_ | _8415_ /*10742*/;
assign _8417_ = ~Q[13] /*10741*/;
assign _8416_ = _8417_ & D[21] /*10740*/;
assign _8419_ = _8054_ & _8416_ /*10735*/;
assign _8420_ = _8054_ ^ _8416_ /*10738*/;
assign _8421_ = _8412_ & _8420_ /*10736*/;
assign _8278_ = _8412_ ^ _8420_ /*10737*/;
assign _8418_ = _8419_ | _8421_ /*10734*/;
assign _8423_ = ~Q[13] /*10733*/;
assign _8422_ = _8423_ & D[22] /*10732*/;
assign _8425_ = _8055_ & _8422_ /*10727*/;
assign _8426_ = _8055_ ^ _8422_ /*10730*/;
assign _8427_ = _8418_ & _8426_ /*10728*/;
assign _8279_ = _8418_ ^ _8426_ /*10729*/;
assign _8424_ = _8425_ | _8427_ /*10726*/;
assign _8429_ = ~Q[13] /*10725*/;
assign _8428_ = _8429_ & D[23] /*10724*/;
assign _8431_ = _8056_ & _8428_ /*10719*/;
assign _8432_ = _8056_ ^ _8428_ /*10722*/;
assign _8433_ = _8424_ & _8432_ /*10720*/;
assign _8280_ = _8424_ ^ _8432_ /*10721*/;
assign _8430_ = _8431_ | _8433_ /*10718*/;
assign _8435_ = ~Q[13] /*10717*/;
assign _8434_ = _8435_ & D[24] /*10716*/;
assign _8437_ = _8057_ & _8434_ /*10711*/;
assign _8438_ = _8057_ ^ _8434_ /*10714*/;
assign _8439_ = _8430_ & _8438_ /*10712*/;
assign _8281_ = _8430_ ^ _8438_ /*10713*/;
assign _8436_ = _8437_ | _8439_ /*10710*/;
assign _8441_ = ~Q[13] /*10709*/;
assign _8440_ = _8441_ & D[25] /*10708*/;
assign _8443_ = _8058_ & _8440_ /*10703*/;
assign _8444_ = _8058_ ^ _8440_ /*10706*/;
assign _8445_ = _8436_ & _8444_ /*10704*/;
assign _8282_ = _8436_ ^ _8444_ /*10705*/;
assign _8442_ = _8443_ | _8445_ /*10702*/;
assign _8447_ = ~Q[13] /*10701*/;
assign _8446_ = _8447_ & D[26] /*10700*/;
assign _8449_ = _8059_ & _8446_ /*10695*/;
assign _8450_ = _8059_ ^ _8446_ /*10698*/;
assign _8451_ = _8442_ & _8450_ /*10696*/;
assign _8283_ = _8442_ ^ _8450_ /*10697*/;
assign _8448_ = _8449_ | _8451_ /*10694*/;
assign _8453_ = ~Q[13] /*10693*/;
assign _8452_ = _8453_ & D[27] /*10692*/;
assign _8455_ = _8060_ & _8452_ /*10687*/;
assign _8456_ = _8060_ ^ _8452_ /*10690*/;
assign _8457_ = _8448_ & _8456_ /*10688*/;
assign _8284_ = _8448_ ^ _8456_ /*10689*/;
assign _8454_ = _8455_ | _8457_ /*10686*/;
assign _8459_ = ~Q[13] /*10685*/;
assign _8458_ = _8459_ & D[28] /*10684*/;
assign _8461_ = _8061_ & _8458_ /*10679*/;
assign _8462_ = _8061_ ^ _8458_ /*10682*/;
assign _8463_ = _8454_ & _8462_ /*10680*/;
assign _8285_ = _8454_ ^ _8462_ /*10681*/;
assign _8460_ = _8461_ | _8463_ /*10678*/;
assign _8465_ = ~Q[13] /*10677*/;
assign _8464_ = _8465_ & D[29] /*10676*/;
assign _8467_ = _8062_ & _8464_ /*10671*/;
assign _8468_ = _8062_ ^ _8464_ /*10674*/;
assign _8469_ = _8460_ & _8468_ /*10672*/;
assign _8286_ = _8460_ ^ _8468_ /*10673*/;
assign _8466_ = _8467_ | _8469_ /*10670*/;
assign _8471_ = ~Q[13] /*10669*/;
assign _8470_ = _8471_ & D[30] /*10668*/;
assign _8473_ = _8063_ & _8470_ /*10663*/;
assign _8474_ = _8063_ ^ _8470_ /*10666*/;
assign _8475_ = _8466_ & _8474_ /*10664*/;
assign _8287_ = _8466_ ^ _8474_ /*10665*/;
assign _8472_ = _8473_ | _8475_ /*10662*/;
assign _8477_ = ~Q[13] /*10661*/;
assign _8476_ = _8477_ & zeroWire /*10660*/;
assign _8478_ = _8064_ ^ _8476_ /*10658*/;
assign _8288_ = _8478_ ^ _8472_ /*10657*/;
assign _8517_ = ~D[0] /*10531*/;
assign _8514_ = R_0[12] & _8517_ /*10527*/;
assign _8515_ = R_0[12] ^ _8517_ /*10530*/;
assign _8516_ = oneWire & _8515_ /*10528*/;
assign _8481_ = oneWire ^ _8515_ /*10529*/;
assign _8513_ = _8514_ | _8516_ /*10526*/;
assign _8522_ = ~D[1] /*10525*/;
assign _8519_ = _8257_ & _8522_ /*10521*/;
assign _8520_ = _8257_ ^ _8522_ /*10524*/;
assign _8521_ = _8513_ & _8520_ /*10522*/;
assign _8482_ = _8513_ ^ _8520_ /*10523*/;
assign _8518_ = _8519_ | _8521_ /*10520*/;
assign _8527_ = ~D[2] /*10519*/;
assign _8524_ = _8258_ & _8527_ /*10515*/;
assign _8525_ = _8258_ ^ _8527_ /*10518*/;
assign _8526_ = _8518_ & _8525_ /*10516*/;
assign _8483_ = _8518_ ^ _8525_ /*10517*/;
assign _8523_ = _8524_ | _8526_ /*10514*/;
assign _8532_ = ~D[3] /*10513*/;
assign _8529_ = _8259_ & _8532_ /*10509*/;
assign _8530_ = _8259_ ^ _8532_ /*10512*/;
assign _8531_ = _8523_ & _8530_ /*10510*/;
assign _8484_ = _8523_ ^ _8530_ /*10511*/;
assign _8528_ = _8529_ | _8531_ /*10508*/;
assign _8537_ = ~D[4] /*10507*/;
assign _8534_ = _8260_ & _8537_ /*10503*/;
assign _8535_ = _8260_ ^ _8537_ /*10506*/;
assign _8536_ = _8528_ & _8535_ /*10504*/;
assign _8485_ = _8528_ ^ _8535_ /*10505*/;
assign _8533_ = _8534_ | _8536_ /*10502*/;
assign _8542_ = ~D[5] /*10501*/;
assign _8539_ = _8261_ & _8542_ /*10497*/;
assign _8540_ = _8261_ ^ _8542_ /*10500*/;
assign _8541_ = _8533_ & _8540_ /*10498*/;
assign _8486_ = _8533_ ^ _8540_ /*10499*/;
assign _8538_ = _8539_ | _8541_ /*10496*/;
assign _8547_ = ~D[6] /*10495*/;
assign _8544_ = _8262_ & _8547_ /*10491*/;
assign _8545_ = _8262_ ^ _8547_ /*10494*/;
assign _8546_ = _8538_ & _8545_ /*10492*/;
assign _8487_ = _8538_ ^ _8545_ /*10493*/;
assign _8543_ = _8544_ | _8546_ /*10490*/;
assign _8552_ = ~D[7] /*10489*/;
assign _8549_ = _8263_ & _8552_ /*10485*/;
assign _8550_ = _8263_ ^ _8552_ /*10488*/;
assign _8551_ = _8543_ & _8550_ /*10486*/;
assign _8488_ = _8543_ ^ _8550_ /*10487*/;
assign _8548_ = _8549_ | _8551_ /*10484*/;
assign _8557_ = ~D[8] /*10483*/;
assign _8554_ = _8264_ & _8557_ /*10479*/;
assign _8555_ = _8264_ ^ _8557_ /*10482*/;
assign _8556_ = _8548_ & _8555_ /*10480*/;
assign _8489_ = _8548_ ^ _8555_ /*10481*/;
assign _8553_ = _8554_ | _8556_ /*10478*/;
assign _8562_ = ~D[9] /*10477*/;
assign _8559_ = _8265_ & _8562_ /*10473*/;
assign _8560_ = _8265_ ^ _8562_ /*10476*/;
assign _8561_ = _8553_ & _8560_ /*10474*/;
assign _8490_ = _8553_ ^ _8560_ /*10475*/;
assign _8558_ = _8559_ | _8561_ /*10472*/;
assign _8567_ = ~D[10] /*10471*/;
assign _8564_ = _8266_ & _8567_ /*10467*/;
assign _8565_ = _8266_ ^ _8567_ /*10470*/;
assign _8566_ = _8558_ & _8565_ /*10468*/;
assign _8491_ = _8558_ ^ _8565_ /*10469*/;
assign _8563_ = _8564_ | _8566_ /*10466*/;
assign _8572_ = ~D[11] /*10465*/;
assign _8569_ = _8267_ & _8572_ /*10461*/;
assign _8570_ = _8267_ ^ _8572_ /*10464*/;
assign _8571_ = _8563_ & _8570_ /*10462*/;
assign _8492_ = _8563_ ^ _8570_ /*10463*/;
assign _8568_ = _8569_ | _8571_ /*10460*/;
assign _8577_ = ~D[12] /*10459*/;
assign _8574_ = _8268_ & _8577_ /*10455*/;
assign _8575_ = _8268_ ^ _8577_ /*10458*/;
assign _8576_ = _8568_ & _8575_ /*10456*/;
assign _8493_ = _8568_ ^ _8575_ /*10457*/;
assign _8573_ = _8574_ | _8576_ /*10454*/;
assign _8582_ = ~D[13] /*10453*/;
assign _8579_ = _8269_ & _8582_ /*10449*/;
assign _8580_ = _8269_ ^ _8582_ /*10452*/;
assign _8581_ = _8573_ & _8580_ /*10450*/;
assign _8494_ = _8573_ ^ _8580_ /*10451*/;
assign _8578_ = _8579_ | _8581_ /*10448*/;
assign _8587_ = ~D[14] /*10447*/;
assign _8584_ = _8270_ & _8587_ /*10443*/;
assign _8585_ = _8270_ ^ _8587_ /*10446*/;
assign _8586_ = _8578_ & _8585_ /*10444*/;
assign _8495_ = _8578_ ^ _8585_ /*10445*/;
assign _8583_ = _8584_ | _8586_ /*10442*/;
assign _8592_ = ~D[15] /*10441*/;
assign _8589_ = _8271_ & _8592_ /*10437*/;
assign _8590_ = _8271_ ^ _8592_ /*10440*/;
assign _8591_ = _8583_ & _8590_ /*10438*/;
assign _8496_ = _8583_ ^ _8590_ /*10439*/;
assign _8588_ = _8589_ | _8591_ /*10436*/;
assign _8597_ = ~D[16] /*10435*/;
assign _8594_ = _8272_ & _8597_ /*10431*/;
assign _8595_ = _8272_ ^ _8597_ /*10434*/;
assign _8596_ = _8588_ & _8595_ /*10432*/;
assign _8497_ = _8588_ ^ _8595_ /*10433*/;
assign _8593_ = _8594_ | _8596_ /*10430*/;
assign _8602_ = ~D[17] /*10429*/;
assign _8599_ = _8273_ & _8602_ /*10425*/;
assign _8600_ = _8273_ ^ _8602_ /*10428*/;
assign _8601_ = _8593_ & _8600_ /*10426*/;
assign _8498_ = _8593_ ^ _8600_ /*10427*/;
assign _8598_ = _8599_ | _8601_ /*10424*/;
assign _8607_ = ~D[18] /*10423*/;
assign _8604_ = _8274_ & _8607_ /*10419*/;
assign _8605_ = _8274_ ^ _8607_ /*10422*/;
assign _8606_ = _8598_ & _8605_ /*10420*/;
assign _8499_ = _8598_ ^ _8605_ /*10421*/;
assign _8603_ = _8604_ | _8606_ /*10418*/;
assign _8612_ = ~D[19] /*10417*/;
assign _8609_ = _8275_ & _8612_ /*10413*/;
assign _8610_ = _8275_ ^ _8612_ /*10416*/;
assign _8611_ = _8603_ & _8610_ /*10414*/;
assign _8500_ = _8603_ ^ _8610_ /*10415*/;
assign _8608_ = _8609_ | _8611_ /*10412*/;
assign _8617_ = ~D[20] /*10411*/;
assign _8614_ = _8276_ & _8617_ /*10407*/;
assign _8615_ = _8276_ ^ _8617_ /*10410*/;
assign _8616_ = _8608_ & _8615_ /*10408*/;
assign _8501_ = _8608_ ^ _8615_ /*10409*/;
assign _8613_ = _8614_ | _8616_ /*10406*/;
assign _8622_ = ~D[21] /*10405*/;
assign _8619_ = _8277_ & _8622_ /*10401*/;
assign _8620_ = _8277_ ^ _8622_ /*10404*/;
assign _8621_ = _8613_ & _8620_ /*10402*/;
assign _8502_ = _8613_ ^ _8620_ /*10403*/;
assign _8618_ = _8619_ | _8621_ /*10400*/;
assign _8627_ = ~D[22] /*10399*/;
assign _8624_ = _8278_ & _8627_ /*10395*/;
assign _8625_ = _8278_ ^ _8627_ /*10398*/;
assign _8626_ = _8618_ & _8625_ /*10396*/;
assign _8503_ = _8618_ ^ _8625_ /*10397*/;
assign _8623_ = _8624_ | _8626_ /*10394*/;
assign _8632_ = ~D[23] /*10393*/;
assign _8629_ = _8279_ & _8632_ /*10389*/;
assign _8630_ = _8279_ ^ _8632_ /*10392*/;
assign _8631_ = _8623_ & _8630_ /*10390*/;
assign _8504_ = _8623_ ^ _8630_ /*10391*/;
assign _8628_ = _8629_ | _8631_ /*10388*/;
assign _8637_ = ~D[24] /*10387*/;
assign _8634_ = _8280_ & _8637_ /*10383*/;
assign _8635_ = _8280_ ^ _8637_ /*10386*/;
assign _8636_ = _8628_ & _8635_ /*10384*/;
assign _8505_ = _8628_ ^ _8635_ /*10385*/;
assign _8633_ = _8634_ | _8636_ /*10382*/;
assign _8642_ = ~D[25] /*10381*/;
assign _8639_ = _8281_ & _8642_ /*10377*/;
assign _8640_ = _8281_ ^ _8642_ /*10380*/;
assign _8641_ = _8633_ & _8640_ /*10378*/;
assign _8506_ = _8633_ ^ _8640_ /*10379*/;
assign _8638_ = _8639_ | _8641_ /*10376*/;
assign _8647_ = ~D[26] /*10375*/;
assign _8644_ = _8282_ & _8647_ /*10371*/;
assign _8645_ = _8282_ ^ _8647_ /*10374*/;
assign _8646_ = _8638_ & _8645_ /*10372*/;
assign _8507_ = _8638_ ^ _8645_ /*10373*/;
assign _8643_ = _8644_ | _8646_ /*10370*/;
assign _8652_ = ~D[27] /*10369*/;
assign _8649_ = _8283_ & _8652_ /*10365*/;
assign _8650_ = _8283_ ^ _8652_ /*10368*/;
assign _8651_ = _8643_ & _8650_ /*10366*/;
assign _8508_ = _8643_ ^ _8650_ /*10367*/;
assign _8648_ = _8649_ | _8651_ /*10364*/;
assign _8657_ = ~D[28] /*10363*/;
assign _8654_ = _8284_ & _8657_ /*10359*/;
assign _8655_ = _8284_ ^ _8657_ /*10362*/;
assign _8656_ = _8648_ & _8655_ /*10360*/;
assign _8509_ = _8648_ ^ _8655_ /*10361*/;
assign _8653_ = _8654_ | _8656_ /*10358*/;
assign _8662_ = ~D[29] /*10357*/;
assign _8659_ = _8285_ & _8662_ /*10353*/;
assign _8660_ = _8285_ ^ _8662_ /*10356*/;
assign _8661_ = _8653_ & _8660_ /*10354*/;
assign _8510_ = _8653_ ^ _8660_ /*10355*/;
assign _8658_ = _8659_ | _8661_ /*10352*/;
assign _8667_ = ~D[30] /*10351*/;
assign _8664_ = _8286_ & _8667_ /*10347*/;
assign _8665_ = _8286_ ^ _8667_ /*10350*/;
assign _8666_ = _8658_ & _8665_ /*10348*/;
assign _8511_ = _8658_ ^ _8665_ /*10349*/;
assign _8663_ = _8664_ | _8666_ /*10346*/;
assign _8668_ = _8287_ & oneWire /*10341*/;
assign _8669_ = _8287_ ^ oneWire /*10344*/;
assign _8670_ = _8663_ & _8669_ /*10342*/;
assign _8512_ = _8663_ ^ _8669_ /*10343*/;
assign Q[12] = _8668_ | _8670_ /*10340*/;
assign _8739_ = ~Q[12] /*10147*/;
assign _8738_ = _8739_ & D[0] /*10146*/;
assign _8741_ = _8481_ & _8738_ /*10141*/;
assign _8742_ = _8481_ ^ _8738_ /*10144*/;
assign _8743_ = zeroWire & _8742_ /*10142*/;
assign _8705_ = zeroWire ^ _8742_ /*10143*/;
assign _8740_ = _8741_ | _8743_ /*10140*/;
assign _8745_ = ~Q[12] /*10139*/;
assign _8744_ = _8745_ & D[1] /*10138*/;
assign _8747_ = _8482_ & _8744_ /*10133*/;
assign _8748_ = _8482_ ^ _8744_ /*10136*/;
assign _8749_ = _8740_ & _8748_ /*10134*/;
assign _8706_ = _8740_ ^ _8748_ /*10135*/;
assign _8746_ = _8747_ | _8749_ /*10132*/;
assign _8751_ = ~Q[12] /*10131*/;
assign _8750_ = _8751_ & D[2] /*10130*/;
assign _8753_ = _8483_ & _8750_ /*10125*/;
assign _8754_ = _8483_ ^ _8750_ /*10128*/;
assign _8755_ = _8746_ & _8754_ /*10126*/;
assign _8707_ = _8746_ ^ _8754_ /*10127*/;
assign _8752_ = _8753_ | _8755_ /*10124*/;
assign _8757_ = ~Q[12] /*10123*/;
assign _8756_ = _8757_ & D[3] /*10122*/;
assign _8759_ = _8484_ & _8756_ /*10117*/;
assign _8760_ = _8484_ ^ _8756_ /*10120*/;
assign _8761_ = _8752_ & _8760_ /*10118*/;
assign _8708_ = _8752_ ^ _8760_ /*10119*/;
assign _8758_ = _8759_ | _8761_ /*10116*/;
assign _8763_ = ~Q[12] /*10115*/;
assign _8762_ = _8763_ & D[4] /*10114*/;
assign _8765_ = _8485_ & _8762_ /*10109*/;
assign _8766_ = _8485_ ^ _8762_ /*10112*/;
assign _8767_ = _8758_ & _8766_ /*10110*/;
assign _8709_ = _8758_ ^ _8766_ /*10111*/;
assign _8764_ = _8765_ | _8767_ /*10108*/;
assign _8769_ = ~Q[12] /*10107*/;
assign _8768_ = _8769_ & D[5] /*10106*/;
assign _8771_ = _8486_ & _8768_ /*10101*/;
assign _8772_ = _8486_ ^ _8768_ /*10104*/;
assign _8773_ = _8764_ & _8772_ /*10102*/;
assign _8710_ = _8764_ ^ _8772_ /*10103*/;
assign _8770_ = _8771_ | _8773_ /*10100*/;
assign _8775_ = ~Q[12] /*10099*/;
assign _8774_ = _8775_ & D[6] /*10098*/;
assign _8777_ = _8487_ & _8774_ /*10093*/;
assign _8778_ = _8487_ ^ _8774_ /*10096*/;
assign _8779_ = _8770_ & _8778_ /*10094*/;
assign _8711_ = _8770_ ^ _8778_ /*10095*/;
assign _8776_ = _8777_ | _8779_ /*10092*/;
assign _8781_ = ~Q[12] /*10091*/;
assign _8780_ = _8781_ & D[7] /*10090*/;
assign _8783_ = _8488_ & _8780_ /*10085*/;
assign _8784_ = _8488_ ^ _8780_ /*10088*/;
assign _8785_ = _8776_ & _8784_ /*10086*/;
assign _8712_ = _8776_ ^ _8784_ /*10087*/;
assign _8782_ = _8783_ | _8785_ /*10084*/;
assign _8787_ = ~Q[12] /*10083*/;
assign _8786_ = _8787_ & D[8] /*10082*/;
assign _8789_ = _8489_ & _8786_ /*10077*/;
assign _8790_ = _8489_ ^ _8786_ /*10080*/;
assign _8791_ = _8782_ & _8790_ /*10078*/;
assign _8713_ = _8782_ ^ _8790_ /*10079*/;
assign _8788_ = _8789_ | _8791_ /*10076*/;
assign _8793_ = ~Q[12] /*10075*/;
assign _8792_ = _8793_ & D[9] /*10074*/;
assign _8795_ = _8490_ & _8792_ /*10069*/;
assign _8796_ = _8490_ ^ _8792_ /*10072*/;
assign _8797_ = _8788_ & _8796_ /*10070*/;
assign _8714_ = _8788_ ^ _8796_ /*10071*/;
assign _8794_ = _8795_ | _8797_ /*10068*/;
assign _8799_ = ~Q[12] /*10067*/;
assign _8798_ = _8799_ & D[10] /*10066*/;
assign _8801_ = _8491_ & _8798_ /*10061*/;
assign _8802_ = _8491_ ^ _8798_ /*10064*/;
assign _8803_ = _8794_ & _8802_ /*10062*/;
assign _8715_ = _8794_ ^ _8802_ /*10063*/;
assign _8800_ = _8801_ | _8803_ /*10060*/;
assign _8805_ = ~Q[12] /*10059*/;
assign _8804_ = _8805_ & D[11] /*10058*/;
assign _8807_ = _8492_ & _8804_ /*10053*/;
assign _8808_ = _8492_ ^ _8804_ /*10056*/;
assign _8809_ = _8800_ & _8808_ /*10054*/;
assign _8716_ = _8800_ ^ _8808_ /*10055*/;
assign _8806_ = _8807_ | _8809_ /*10052*/;
assign _8811_ = ~Q[12] /*10051*/;
assign _8810_ = _8811_ & D[12] /*10050*/;
assign _8813_ = _8493_ & _8810_ /*10045*/;
assign _8814_ = _8493_ ^ _8810_ /*10048*/;
assign _8815_ = _8806_ & _8814_ /*10046*/;
assign _8717_ = _8806_ ^ _8814_ /*10047*/;
assign _8812_ = _8813_ | _8815_ /*10044*/;
assign _8817_ = ~Q[12] /*10043*/;
assign _8816_ = _8817_ & D[13] /*10042*/;
assign _8819_ = _8494_ & _8816_ /*10037*/;
assign _8820_ = _8494_ ^ _8816_ /*10040*/;
assign _8821_ = _8812_ & _8820_ /*10038*/;
assign _8718_ = _8812_ ^ _8820_ /*10039*/;
assign _8818_ = _8819_ | _8821_ /*10036*/;
assign _8823_ = ~Q[12] /*10035*/;
assign _8822_ = _8823_ & D[14] /*10034*/;
assign _8825_ = _8495_ & _8822_ /*10029*/;
assign _8826_ = _8495_ ^ _8822_ /*10032*/;
assign _8827_ = _8818_ & _8826_ /*10030*/;
assign _8719_ = _8818_ ^ _8826_ /*10031*/;
assign _8824_ = _8825_ | _8827_ /*10028*/;
assign _8829_ = ~Q[12] /*10027*/;
assign _8828_ = _8829_ & D[15] /*10026*/;
assign _8831_ = _8496_ & _8828_ /*10021*/;
assign _8832_ = _8496_ ^ _8828_ /*10024*/;
assign _8833_ = _8824_ & _8832_ /*10022*/;
assign _8720_ = _8824_ ^ _8832_ /*10023*/;
assign _8830_ = _8831_ | _8833_ /*10020*/;
assign _8835_ = ~Q[12] /*10019*/;
assign _8834_ = _8835_ & D[16] /*10018*/;
assign _8837_ = _8497_ & _8834_ /*10013*/;
assign _8838_ = _8497_ ^ _8834_ /*10016*/;
assign _8839_ = _8830_ & _8838_ /*10014*/;
assign _8721_ = _8830_ ^ _8838_ /*10015*/;
assign _8836_ = _8837_ | _8839_ /*10012*/;
assign _8841_ = ~Q[12] /*10011*/;
assign _8840_ = _8841_ & D[17] /*10010*/;
assign _8843_ = _8498_ & _8840_ /*10005*/;
assign _8844_ = _8498_ ^ _8840_ /*10008*/;
assign _8845_ = _8836_ & _8844_ /*10006*/;
assign _8722_ = _8836_ ^ _8844_ /*10007*/;
assign _8842_ = _8843_ | _8845_ /*10004*/;
assign _8847_ = ~Q[12] /*10003*/;
assign _8846_ = _8847_ & D[18] /*10002*/;
assign _8849_ = _8499_ & _8846_ /*9997*/;
assign _8850_ = _8499_ ^ _8846_ /*10000*/;
assign _8851_ = _8842_ & _8850_ /*9998*/;
assign _8723_ = _8842_ ^ _8850_ /*9999*/;
assign _8848_ = _8849_ | _8851_ /*9996*/;
assign _8853_ = ~Q[12] /*9995*/;
assign _8852_ = _8853_ & D[19] /*9994*/;
assign _8855_ = _8500_ & _8852_ /*9989*/;
assign _8856_ = _8500_ ^ _8852_ /*9992*/;
assign _8857_ = _8848_ & _8856_ /*9990*/;
assign _8724_ = _8848_ ^ _8856_ /*9991*/;
assign _8854_ = _8855_ | _8857_ /*9988*/;
assign _8859_ = ~Q[12] /*9987*/;
assign _8858_ = _8859_ & D[20] /*9986*/;
assign _8861_ = _8501_ & _8858_ /*9981*/;
assign _8862_ = _8501_ ^ _8858_ /*9984*/;
assign _8863_ = _8854_ & _8862_ /*9982*/;
assign _8725_ = _8854_ ^ _8862_ /*9983*/;
assign _8860_ = _8861_ | _8863_ /*9980*/;
assign _8865_ = ~Q[12] /*9979*/;
assign _8864_ = _8865_ & D[21] /*9978*/;
assign _8867_ = _8502_ & _8864_ /*9973*/;
assign _8868_ = _8502_ ^ _8864_ /*9976*/;
assign _8869_ = _8860_ & _8868_ /*9974*/;
assign _8726_ = _8860_ ^ _8868_ /*9975*/;
assign _8866_ = _8867_ | _8869_ /*9972*/;
assign _8871_ = ~Q[12] /*9971*/;
assign _8870_ = _8871_ & D[22] /*9970*/;
assign _8873_ = _8503_ & _8870_ /*9965*/;
assign _8874_ = _8503_ ^ _8870_ /*9968*/;
assign _8875_ = _8866_ & _8874_ /*9966*/;
assign _8727_ = _8866_ ^ _8874_ /*9967*/;
assign _8872_ = _8873_ | _8875_ /*9964*/;
assign _8877_ = ~Q[12] /*9963*/;
assign _8876_ = _8877_ & D[23] /*9962*/;
assign _8879_ = _8504_ & _8876_ /*9957*/;
assign _8880_ = _8504_ ^ _8876_ /*9960*/;
assign _8881_ = _8872_ & _8880_ /*9958*/;
assign _8728_ = _8872_ ^ _8880_ /*9959*/;
assign _8878_ = _8879_ | _8881_ /*9956*/;
assign _8883_ = ~Q[12] /*9955*/;
assign _8882_ = _8883_ & D[24] /*9954*/;
assign _8885_ = _8505_ & _8882_ /*9949*/;
assign _8886_ = _8505_ ^ _8882_ /*9952*/;
assign _8887_ = _8878_ & _8886_ /*9950*/;
assign _8729_ = _8878_ ^ _8886_ /*9951*/;
assign _8884_ = _8885_ | _8887_ /*9948*/;
assign _8889_ = ~Q[12] /*9947*/;
assign _8888_ = _8889_ & D[25] /*9946*/;
assign _8891_ = _8506_ & _8888_ /*9941*/;
assign _8892_ = _8506_ ^ _8888_ /*9944*/;
assign _8893_ = _8884_ & _8892_ /*9942*/;
assign _8730_ = _8884_ ^ _8892_ /*9943*/;
assign _8890_ = _8891_ | _8893_ /*9940*/;
assign _8895_ = ~Q[12] /*9939*/;
assign _8894_ = _8895_ & D[26] /*9938*/;
assign _8897_ = _8507_ & _8894_ /*9933*/;
assign _8898_ = _8507_ ^ _8894_ /*9936*/;
assign _8899_ = _8890_ & _8898_ /*9934*/;
assign _8731_ = _8890_ ^ _8898_ /*9935*/;
assign _8896_ = _8897_ | _8899_ /*9932*/;
assign _8901_ = ~Q[12] /*9931*/;
assign _8900_ = _8901_ & D[27] /*9930*/;
assign _8903_ = _8508_ & _8900_ /*9925*/;
assign _8904_ = _8508_ ^ _8900_ /*9928*/;
assign _8905_ = _8896_ & _8904_ /*9926*/;
assign _8732_ = _8896_ ^ _8904_ /*9927*/;
assign _8902_ = _8903_ | _8905_ /*9924*/;
assign _8907_ = ~Q[12] /*9923*/;
assign _8906_ = _8907_ & D[28] /*9922*/;
assign _8909_ = _8509_ & _8906_ /*9917*/;
assign _8910_ = _8509_ ^ _8906_ /*9920*/;
assign _8911_ = _8902_ & _8910_ /*9918*/;
assign _8733_ = _8902_ ^ _8910_ /*9919*/;
assign _8908_ = _8909_ | _8911_ /*9916*/;
assign _8913_ = ~Q[12] /*9915*/;
assign _8912_ = _8913_ & D[29] /*9914*/;
assign _8915_ = _8510_ & _8912_ /*9909*/;
assign _8916_ = _8510_ ^ _8912_ /*9912*/;
assign _8917_ = _8908_ & _8916_ /*9910*/;
assign _8734_ = _8908_ ^ _8916_ /*9911*/;
assign _8914_ = _8915_ | _8917_ /*9908*/;
assign _8919_ = ~Q[12] /*9907*/;
assign _8918_ = _8919_ & D[30] /*9906*/;
assign _8921_ = _8511_ & _8918_ /*9901*/;
assign _8922_ = _8511_ ^ _8918_ /*9904*/;
assign _8923_ = _8914_ & _8922_ /*9902*/;
assign _8735_ = _8914_ ^ _8922_ /*9903*/;
assign _8920_ = _8921_ | _8923_ /*9900*/;
assign _8925_ = ~Q[12] /*9899*/;
assign _8924_ = _8925_ & zeroWire /*9898*/;
assign _8926_ = _8512_ ^ _8924_ /*9896*/;
assign _8736_ = _8926_ ^ _8920_ /*9895*/;
assign _8965_ = ~D[0] /*9769*/;
assign _8962_ = R_0[11] & _8965_ /*9765*/;
assign _8963_ = R_0[11] ^ _8965_ /*9768*/;
assign _8964_ = oneWire & _8963_ /*9766*/;
assign _8929_ = oneWire ^ _8963_ /*9767*/;
assign _8961_ = _8962_ | _8964_ /*9764*/;
assign _8970_ = ~D[1] /*9763*/;
assign _8967_ = _8705_ & _8970_ /*9759*/;
assign _8968_ = _8705_ ^ _8970_ /*9762*/;
assign _8969_ = _8961_ & _8968_ /*9760*/;
assign _8930_ = _8961_ ^ _8968_ /*9761*/;
assign _8966_ = _8967_ | _8969_ /*9758*/;
assign _8975_ = ~D[2] /*9757*/;
assign _8972_ = _8706_ & _8975_ /*9753*/;
assign _8973_ = _8706_ ^ _8975_ /*9756*/;
assign _8974_ = _8966_ & _8973_ /*9754*/;
assign _8931_ = _8966_ ^ _8973_ /*9755*/;
assign _8971_ = _8972_ | _8974_ /*9752*/;
assign _8980_ = ~D[3] /*9751*/;
assign _8977_ = _8707_ & _8980_ /*9747*/;
assign _8978_ = _8707_ ^ _8980_ /*9750*/;
assign _8979_ = _8971_ & _8978_ /*9748*/;
assign _8932_ = _8971_ ^ _8978_ /*9749*/;
assign _8976_ = _8977_ | _8979_ /*9746*/;
assign _8985_ = ~D[4] /*9745*/;
assign _8982_ = _8708_ & _8985_ /*9741*/;
assign _8983_ = _8708_ ^ _8985_ /*9744*/;
assign _8984_ = _8976_ & _8983_ /*9742*/;
assign _8933_ = _8976_ ^ _8983_ /*9743*/;
assign _8981_ = _8982_ | _8984_ /*9740*/;
assign _8990_ = ~D[5] /*9739*/;
assign _8987_ = _8709_ & _8990_ /*9735*/;
assign _8988_ = _8709_ ^ _8990_ /*9738*/;
assign _8989_ = _8981_ & _8988_ /*9736*/;
assign _8934_ = _8981_ ^ _8988_ /*9737*/;
assign _8986_ = _8987_ | _8989_ /*9734*/;
assign _8995_ = ~D[6] /*9733*/;
assign _8992_ = _8710_ & _8995_ /*9729*/;
assign _8993_ = _8710_ ^ _8995_ /*9732*/;
assign _8994_ = _8986_ & _8993_ /*9730*/;
assign _8935_ = _8986_ ^ _8993_ /*9731*/;
assign _8991_ = _8992_ | _8994_ /*9728*/;
assign _9000_ = ~D[7] /*9727*/;
assign _8997_ = _8711_ & _9000_ /*9723*/;
assign _8998_ = _8711_ ^ _9000_ /*9726*/;
assign _8999_ = _8991_ & _8998_ /*9724*/;
assign _8936_ = _8991_ ^ _8998_ /*9725*/;
assign _8996_ = _8997_ | _8999_ /*9722*/;
assign _9005_ = ~D[8] /*9721*/;
assign _9002_ = _8712_ & _9005_ /*9717*/;
assign _9003_ = _8712_ ^ _9005_ /*9720*/;
assign _9004_ = _8996_ & _9003_ /*9718*/;
assign _8937_ = _8996_ ^ _9003_ /*9719*/;
assign _9001_ = _9002_ | _9004_ /*9716*/;
assign _9010_ = ~D[9] /*9715*/;
assign _9007_ = _8713_ & _9010_ /*9711*/;
assign _9008_ = _8713_ ^ _9010_ /*9714*/;
assign _9009_ = _9001_ & _9008_ /*9712*/;
assign _8938_ = _9001_ ^ _9008_ /*9713*/;
assign _9006_ = _9007_ | _9009_ /*9710*/;
assign _9015_ = ~D[10] /*9709*/;
assign _9012_ = _8714_ & _9015_ /*9705*/;
assign _9013_ = _8714_ ^ _9015_ /*9708*/;
assign _9014_ = _9006_ & _9013_ /*9706*/;
assign _8939_ = _9006_ ^ _9013_ /*9707*/;
assign _9011_ = _9012_ | _9014_ /*9704*/;
assign _9020_ = ~D[11] /*9703*/;
assign _9017_ = _8715_ & _9020_ /*9699*/;
assign _9018_ = _8715_ ^ _9020_ /*9702*/;
assign _9019_ = _9011_ & _9018_ /*9700*/;
assign _8940_ = _9011_ ^ _9018_ /*9701*/;
assign _9016_ = _9017_ | _9019_ /*9698*/;
assign _9025_ = ~D[12] /*9697*/;
assign _9022_ = _8716_ & _9025_ /*9693*/;
assign _9023_ = _8716_ ^ _9025_ /*9696*/;
assign _9024_ = _9016_ & _9023_ /*9694*/;
assign _8941_ = _9016_ ^ _9023_ /*9695*/;
assign _9021_ = _9022_ | _9024_ /*9692*/;
assign _9030_ = ~D[13] /*9691*/;
assign _9027_ = _8717_ & _9030_ /*9687*/;
assign _9028_ = _8717_ ^ _9030_ /*9690*/;
assign _9029_ = _9021_ & _9028_ /*9688*/;
assign _8942_ = _9021_ ^ _9028_ /*9689*/;
assign _9026_ = _9027_ | _9029_ /*9686*/;
assign _9035_ = ~D[14] /*9685*/;
assign _9032_ = _8718_ & _9035_ /*9681*/;
assign _9033_ = _8718_ ^ _9035_ /*9684*/;
assign _9034_ = _9026_ & _9033_ /*9682*/;
assign _8943_ = _9026_ ^ _9033_ /*9683*/;
assign _9031_ = _9032_ | _9034_ /*9680*/;
assign _9040_ = ~D[15] /*9679*/;
assign _9037_ = _8719_ & _9040_ /*9675*/;
assign _9038_ = _8719_ ^ _9040_ /*9678*/;
assign _9039_ = _9031_ & _9038_ /*9676*/;
assign _8944_ = _9031_ ^ _9038_ /*9677*/;
assign _9036_ = _9037_ | _9039_ /*9674*/;
assign _9045_ = ~D[16] /*9673*/;
assign _9042_ = _8720_ & _9045_ /*9669*/;
assign _9043_ = _8720_ ^ _9045_ /*9672*/;
assign _9044_ = _9036_ & _9043_ /*9670*/;
assign _8945_ = _9036_ ^ _9043_ /*9671*/;
assign _9041_ = _9042_ | _9044_ /*9668*/;
assign _9050_ = ~D[17] /*9667*/;
assign _9047_ = _8721_ & _9050_ /*9663*/;
assign _9048_ = _8721_ ^ _9050_ /*9666*/;
assign _9049_ = _9041_ & _9048_ /*9664*/;
assign _8946_ = _9041_ ^ _9048_ /*9665*/;
assign _9046_ = _9047_ | _9049_ /*9662*/;
assign _9055_ = ~D[18] /*9661*/;
assign _9052_ = _8722_ & _9055_ /*9657*/;
assign _9053_ = _8722_ ^ _9055_ /*9660*/;
assign _9054_ = _9046_ & _9053_ /*9658*/;
assign _8947_ = _9046_ ^ _9053_ /*9659*/;
assign _9051_ = _9052_ | _9054_ /*9656*/;
assign _9060_ = ~D[19] /*9655*/;
assign _9057_ = _8723_ & _9060_ /*9651*/;
assign _9058_ = _8723_ ^ _9060_ /*9654*/;
assign _9059_ = _9051_ & _9058_ /*9652*/;
assign _8948_ = _9051_ ^ _9058_ /*9653*/;
assign _9056_ = _9057_ | _9059_ /*9650*/;
assign _9065_ = ~D[20] /*9649*/;
assign _9062_ = _8724_ & _9065_ /*9645*/;
assign _9063_ = _8724_ ^ _9065_ /*9648*/;
assign _9064_ = _9056_ & _9063_ /*9646*/;
assign _8949_ = _9056_ ^ _9063_ /*9647*/;
assign _9061_ = _9062_ | _9064_ /*9644*/;
assign _9070_ = ~D[21] /*9643*/;
assign _9067_ = _8725_ & _9070_ /*9639*/;
assign _9068_ = _8725_ ^ _9070_ /*9642*/;
assign _9069_ = _9061_ & _9068_ /*9640*/;
assign _8950_ = _9061_ ^ _9068_ /*9641*/;
assign _9066_ = _9067_ | _9069_ /*9638*/;
assign _9075_ = ~D[22] /*9637*/;
assign _9072_ = _8726_ & _9075_ /*9633*/;
assign _9073_ = _8726_ ^ _9075_ /*9636*/;
assign _9074_ = _9066_ & _9073_ /*9634*/;
assign _8951_ = _9066_ ^ _9073_ /*9635*/;
assign _9071_ = _9072_ | _9074_ /*9632*/;
assign _9080_ = ~D[23] /*9631*/;
assign _9077_ = _8727_ & _9080_ /*9627*/;
assign _9078_ = _8727_ ^ _9080_ /*9630*/;
assign _9079_ = _9071_ & _9078_ /*9628*/;
assign _8952_ = _9071_ ^ _9078_ /*9629*/;
assign _9076_ = _9077_ | _9079_ /*9626*/;
assign _9085_ = ~D[24] /*9625*/;
assign _9082_ = _8728_ & _9085_ /*9621*/;
assign _9083_ = _8728_ ^ _9085_ /*9624*/;
assign _9084_ = _9076_ & _9083_ /*9622*/;
assign _8953_ = _9076_ ^ _9083_ /*9623*/;
assign _9081_ = _9082_ | _9084_ /*9620*/;
assign _9090_ = ~D[25] /*9619*/;
assign _9087_ = _8729_ & _9090_ /*9615*/;
assign _9088_ = _8729_ ^ _9090_ /*9618*/;
assign _9089_ = _9081_ & _9088_ /*9616*/;
assign _8954_ = _9081_ ^ _9088_ /*9617*/;
assign _9086_ = _9087_ | _9089_ /*9614*/;
assign _9095_ = ~D[26] /*9613*/;
assign _9092_ = _8730_ & _9095_ /*9609*/;
assign _9093_ = _8730_ ^ _9095_ /*9612*/;
assign _9094_ = _9086_ & _9093_ /*9610*/;
assign _8955_ = _9086_ ^ _9093_ /*9611*/;
assign _9091_ = _9092_ | _9094_ /*9608*/;
assign _9100_ = ~D[27] /*9607*/;
assign _9097_ = _8731_ & _9100_ /*9603*/;
assign _9098_ = _8731_ ^ _9100_ /*9606*/;
assign _9099_ = _9091_ & _9098_ /*9604*/;
assign _8956_ = _9091_ ^ _9098_ /*9605*/;
assign _9096_ = _9097_ | _9099_ /*9602*/;
assign _9105_ = ~D[28] /*9601*/;
assign _9102_ = _8732_ & _9105_ /*9597*/;
assign _9103_ = _8732_ ^ _9105_ /*9600*/;
assign _9104_ = _9096_ & _9103_ /*9598*/;
assign _8957_ = _9096_ ^ _9103_ /*9599*/;
assign _9101_ = _9102_ | _9104_ /*9596*/;
assign _9110_ = ~D[29] /*9595*/;
assign _9107_ = _8733_ & _9110_ /*9591*/;
assign _9108_ = _8733_ ^ _9110_ /*9594*/;
assign _9109_ = _9101_ & _9108_ /*9592*/;
assign _8958_ = _9101_ ^ _9108_ /*9593*/;
assign _9106_ = _9107_ | _9109_ /*9590*/;
assign _9115_ = ~D[30] /*9589*/;
assign _9112_ = _8734_ & _9115_ /*9585*/;
assign _9113_ = _8734_ ^ _9115_ /*9588*/;
assign _9114_ = _9106_ & _9113_ /*9586*/;
assign _8959_ = _9106_ ^ _9113_ /*9587*/;
assign _9111_ = _9112_ | _9114_ /*9584*/;
assign _9116_ = _8735_ & oneWire /*9579*/;
assign _9117_ = _8735_ ^ oneWire /*9582*/;
assign _9118_ = _9111_ & _9117_ /*9580*/;
assign _8960_ = _9111_ ^ _9117_ /*9581*/;
assign Q[11] = _9116_ | _9118_ /*9578*/;
assign _9187_ = ~Q[11] /*9385*/;
assign _9186_ = _9187_ & D[0] /*9384*/;
assign _9189_ = _8929_ & _9186_ /*9379*/;
assign _9190_ = _8929_ ^ _9186_ /*9382*/;
assign _9191_ = zeroWire & _9190_ /*9380*/;
assign _9153_ = zeroWire ^ _9190_ /*9381*/;
assign _9188_ = _9189_ | _9191_ /*9378*/;
assign _9193_ = ~Q[11] /*9377*/;
assign _9192_ = _9193_ & D[1] /*9376*/;
assign _9195_ = _8930_ & _9192_ /*9371*/;
assign _9196_ = _8930_ ^ _9192_ /*9374*/;
assign _9197_ = _9188_ & _9196_ /*9372*/;
assign _9154_ = _9188_ ^ _9196_ /*9373*/;
assign _9194_ = _9195_ | _9197_ /*9370*/;
assign _9199_ = ~Q[11] /*9369*/;
assign _9198_ = _9199_ & D[2] /*9368*/;
assign _9201_ = _8931_ & _9198_ /*9363*/;
assign _9202_ = _8931_ ^ _9198_ /*9366*/;
assign _9203_ = _9194_ & _9202_ /*9364*/;
assign _9155_ = _9194_ ^ _9202_ /*9365*/;
assign _9200_ = _9201_ | _9203_ /*9362*/;
assign _9205_ = ~Q[11] /*9361*/;
assign _9204_ = _9205_ & D[3] /*9360*/;
assign _9207_ = _8932_ & _9204_ /*9355*/;
assign _9208_ = _8932_ ^ _9204_ /*9358*/;
assign _9209_ = _9200_ & _9208_ /*9356*/;
assign _9156_ = _9200_ ^ _9208_ /*9357*/;
assign _9206_ = _9207_ | _9209_ /*9354*/;
assign _9211_ = ~Q[11] /*9353*/;
assign _9210_ = _9211_ & D[4] /*9352*/;
assign _9213_ = _8933_ & _9210_ /*9347*/;
assign _9214_ = _8933_ ^ _9210_ /*9350*/;
assign _9215_ = _9206_ & _9214_ /*9348*/;
assign _9157_ = _9206_ ^ _9214_ /*9349*/;
assign _9212_ = _9213_ | _9215_ /*9346*/;
assign _9217_ = ~Q[11] /*9345*/;
assign _9216_ = _9217_ & D[5] /*9344*/;
assign _9219_ = _8934_ & _9216_ /*9339*/;
assign _9220_ = _8934_ ^ _9216_ /*9342*/;
assign _9221_ = _9212_ & _9220_ /*9340*/;
assign _9158_ = _9212_ ^ _9220_ /*9341*/;
assign _9218_ = _9219_ | _9221_ /*9338*/;
assign _9223_ = ~Q[11] /*9337*/;
assign _9222_ = _9223_ & D[6] /*9336*/;
assign _9225_ = _8935_ & _9222_ /*9331*/;
assign _9226_ = _8935_ ^ _9222_ /*9334*/;
assign _9227_ = _9218_ & _9226_ /*9332*/;
assign _9159_ = _9218_ ^ _9226_ /*9333*/;
assign _9224_ = _9225_ | _9227_ /*9330*/;
assign _9229_ = ~Q[11] /*9329*/;
assign _9228_ = _9229_ & D[7] /*9328*/;
assign _9231_ = _8936_ & _9228_ /*9323*/;
assign _9232_ = _8936_ ^ _9228_ /*9326*/;
assign _9233_ = _9224_ & _9232_ /*9324*/;
assign _9160_ = _9224_ ^ _9232_ /*9325*/;
assign _9230_ = _9231_ | _9233_ /*9322*/;
assign _9235_ = ~Q[11] /*9321*/;
assign _9234_ = _9235_ & D[8] /*9320*/;
assign _9237_ = _8937_ & _9234_ /*9315*/;
assign _9238_ = _8937_ ^ _9234_ /*9318*/;
assign _9239_ = _9230_ & _9238_ /*9316*/;
assign _9161_ = _9230_ ^ _9238_ /*9317*/;
assign _9236_ = _9237_ | _9239_ /*9314*/;
assign _9241_ = ~Q[11] /*9313*/;
assign _9240_ = _9241_ & D[9] /*9312*/;
assign _9243_ = _8938_ & _9240_ /*9307*/;
assign _9244_ = _8938_ ^ _9240_ /*9310*/;
assign _9245_ = _9236_ & _9244_ /*9308*/;
assign _9162_ = _9236_ ^ _9244_ /*9309*/;
assign _9242_ = _9243_ | _9245_ /*9306*/;
assign _9247_ = ~Q[11] /*9305*/;
assign _9246_ = _9247_ & D[10] /*9304*/;
assign _9249_ = _8939_ & _9246_ /*9299*/;
assign _9250_ = _8939_ ^ _9246_ /*9302*/;
assign _9251_ = _9242_ & _9250_ /*9300*/;
assign _9163_ = _9242_ ^ _9250_ /*9301*/;
assign _9248_ = _9249_ | _9251_ /*9298*/;
assign _9253_ = ~Q[11] /*9297*/;
assign _9252_ = _9253_ & D[11] /*9296*/;
assign _9255_ = _8940_ & _9252_ /*9291*/;
assign _9256_ = _8940_ ^ _9252_ /*9294*/;
assign _9257_ = _9248_ & _9256_ /*9292*/;
assign _9164_ = _9248_ ^ _9256_ /*9293*/;
assign _9254_ = _9255_ | _9257_ /*9290*/;
assign _9259_ = ~Q[11] /*9289*/;
assign _9258_ = _9259_ & D[12] /*9288*/;
assign _9261_ = _8941_ & _9258_ /*9283*/;
assign _9262_ = _8941_ ^ _9258_ /*9286*/;
assign _9263_ = _9254_ & _9262_ /*9284*/;
assign _9165_ = _9254_ ^ _9262_ /*9285*/;
assign _9260_ = _9261_ | _9263_ /*9282*/;
assign _9265_ = ~Q[11] /*9281*/;
assign _9264_ = _9265_ & D[13] /*9280*/;
assign _9267_ = _8942_ & _9264_ /*9275*/;
assign _9268_ = _8942_ ^ _9264_ /*9278*/;
assign _9269_ = _9260_ & _9268_ /*9276*/;
assign _9166_ = _9260_ ^ _9268_ /*9277*/;
assign _9266_ = _9267_ | _9269_ /*9274*/;
assign _9271_ = ~Q[11] /*9273*/;
assign _9270_ = _9271_ & D[14] /*9272*/;
assign _9273_ = _8943_ & _9270_ /*9267*/;
assign _9274_ = _8943_ ^ _9270_ /*9270*/;
assign _9275_ = _9266_ & _9274_ /*9268*/;
assign _9167_ = _9266_ ^ _9274_ /*9269*/;
assign _9272_ = _9273_ | _9275_ /*9266*/;
assign _9277_ = ~Q[11] /*9265*/;
assign _9276_ = _9277_ & D[15] /*9264*/;
assign _9279_ = _8944_ & _9276_ /*9259*/;
assign _9280_ = _8944_ ^ _9276_ /*9262*/;
assign _9281_ = _9272_ & _9280_ /*9260*/;
assign _9168_ = _9272_ ^ _9280_ /*9261*/;
assign _9278_ = _9279_ | _9281_ /*9258*/;
assign _9283_ = ~Q[11] /*9257*/;
assign _9282_ = _9283_ & D[16] /*9256*/;
assign _9285_ = _8945_ & _9282_ /*9251*/;
assign _9286_ = _8945_ ^ _9282_ /*9254*/;
assign _9287_ = _9278_ & _9286_ /*9252*/;
assign _9169_ = _9278_ ^ _9286_ /*9253*/;
assign _9284_ = _9285_ | _9287_ /*9250*/;
assign _9289_ = ~Q[11] /*9249*/;
assign _9288_ = _9289_ & D[17] /*9248*/;
assign _9291_ = _8946_ & _9288_ /*9243*/;
assign _9292_ = _8946_ ^ _9288_ /*9246*/;
assign _9293_ = _9284_ & _9292_ /*9244*/;
assign _9170_ = _9284_ ^ _9292_ /*9245*/;
assign _9290_ = _9291_ | _9293_ /*9242*/;
assign _9295_ = ~Q[11] /*9241*/;
assign _9294_ = _9295_ & D[18] /*9240*/;
assign _9297_ = _8947_ & _9294_ /*9235*/;
assign _9298_ = _8947_ ^ _9294_ /*9238*/;
assign _9299_ = _9290_ & _9298_ /*9236*/;
assign _9171_ = _9290_ ^ _9298_ /*9237*/;
assign _9296_ = _9297_ | _9299_ /*9234*/;
assign _9301_ = ~Q[11] /*9233*/;
assign _9300_ = _9301_ & D[19] /*9232*/;
assign _9303_ = _8948_ & _9300_ /*9227*/;
assign _9304_ = _8948_ ^ _9300_ /*9230*/;
assign _9305_ = _9296_ & _9304_ /*9228*/;
assign _9172_ = _9296_ ^ _9304_ /*9229*/;
assign _9302_ = _9303_ | _9305_ /*9226*/;
assign _9307_ = ~Q[11] /*9225*/;
assign _9306_ = _9307_ & D[20] /*9224*/;
assign _9309_ = _8949_ & _9306_ /*9219*/;
assign _9310_ = _8949_ ^ _9306_ /*9222*/;
assign _9311_ = _9302_ & _9310_ /*9220*/;
assign _9173_ = _9302_ ^ _9310_ /*9221*/;
assign _9308_ = _9309_ | _9311_ /*9218*/;
assign _9313_ = ~Q[11] /*9217*/;
assign _9312_ = _9313_ & D[21] /*9216*/;
assign _9315_ = _8950_ & _9312_ /*9211*/;
assign _9316_ = _8950_ ^ _9312_ /*9214*/;
assign _9317_ = _9308_ & _9316_ /*9212*/;
assign _9174_ = _9308_ ^ _9316_ /*9213*/;
assign _9314_ = _9315_ | _9317_ /*9210*/;
assign _9319_ = ~Q[11] /*9209*/;
assign _9318_ = _9319_ & D[22] /*9208*/;
assign _9321_ = _8951_ & _9318_ /*9203*/;
assign _9322_ = _8951_ ^ _9318_ /*9206*/;
assign _9323_ = _9314_ & _9322_ /*9204*/;
assign _9175_ = _9314_ ^ _9322_ /*9205*/;
assign _9320_ = _9321_ | _9323_ /*9202*/;
assign _9325_ = ~Q[11] /*9201*/;
assign _9324_ = _9325_ & D[23] /*9200*/;
assign _9327_ = _8952_ & _9324_ /*9195*/;
assign _9328_ = _8952_ ^ _9324_ /*9198*/;
assign _9329_ = _9320_ & _9328_ /*9196*/;
assign _9176_ = _9320_ ^ _9328_ /*9197*/;
assign _9326_ = _9327_ | _9329_ /*9194*/;
assign _9331_ = ~Q[11] /*9193*/;
assign _9330_ = _9331_ & D[24] /*9192*/;
assign _9333_ = _8953_ & _9330_ /*9187*/;
assign _9334_ = _8953_ ^ _9330_ /*9190*/;
assign _9335_ = _9326_ & _9334_ /*9188*/;
assign _9177_ = _9326_ ^ _9334_ /*9189*/;
assign _9332_ = _9333_ | _9335_ /*9186*/;
assign _9337_ = ~Q[11] /*9185*/;
assign _9336_ = _9337_ & D[25] /*9184*/;
assign _9339_ = _8954_ & _9336_ /*9179*/;
assign _9340_ = _8954_ ^ _9336_ /*9182*/;
assign _9341_ = _9332_ & _9340_ /*9180*/;
assign _9178_ = _9332_ ^ _9340_ /*9181*/;
assign _9338_ = _9339_ | _9341_ /*9178*/;
assign _9343_ = ~Q[11] /*9177*/;
assign _9342_ = _9343_ & D[26] /*9176*/;
assign _9345_ = _8955_ & _9342_ /*9171*/;
assign _9346_ = _8955_ ^ _9342_ /*9174*/;
assign _9347_ = _9338_ & _9346_ /*9172*/;
assign _9179_ = _9338_ ^ _9346_ /*9173*/;
assign _9344_ = _9345_ | _9347_ /*9170*/;
assign _9349_ = ~Q[11] /*9169*/;
assign _9348_ = _9349_ & D[27] /*9168*/;
assign _9351_ = _8956_ & _9348_ /*9163*/;
assign _9352_ = _8956_ ^ _9348_ /*9166*/;
assign _9353_ = _9344_ & _9352_ /*9164*/;
assign _9180_ = _9344_ ^ _9352_ /*9165*/;
assign _9350_ = _9351_ | _9353_ /*9162*/;
assign _9355_ = ~Q[11] /*9161*/;
assign _9354_ = _9355_ & D[28] /*9160*/;
assign _9357_ = _8957_ & _9354_ /*9155*/;
assign _9358_ = _8957_ ^ _9354_ /*9158*/;
assign _9359_ = _9350_ & _9358_ /*9156*/;
assign _9181_ = _9350_ ^ _9358_ /*9157*/;
assign _9356_ = _9357_ | _9359_ /*9154*/;
assign _9361_ = ~Q[11] /*9153*/;
assign _9360_ = _9361_ & D[29] /*9152*/;
assign _9363_ = _8958_ & _9360_ /*9147*/;
assign _9364_ = _8958_ ^ _9360_ /*9150*/;
assign _9365_ = _9356_ & _9364_ /*9148*/;
assign _9182_ = _9356_ ^ _9364_ /*9149*/;
assign _9362_ = _9363_ | _9365_ /*9146*/;
assign _9367_ = ~Q[11] /*9145*/;
assign _9366_ = _9367_ & D[30] /*9144*/;
assign _9369_ = _8959_ & _9366_ /*9139*/;
assign _9370_ = _8959_ ^ _9366_ /*9142*/;
assign _9371_ = _9362_ & _9370_ /*9140*/;
assign _9183_ = _9362_ ^ _9370_ /*9141*/;
assign _9368_ = _9369_ | _9371_ /*9138*/;
assign _9373_ = ~Q[11] /*9137*/;
assign _9372_ = _9373_ & zeroWire /*9136*/;
assign _9374_ = _8960_ ^ _9372_ /*9134*/;
assign _9184_ = _9374_ ^ _9368_ /*9133*/;
assign _9413_ = ~D[0] /*9007*/;
assign _9410_ = R_0[10] & _9413_ /*9003*/;
assign _9411_ = R_0[10] ^ _9413_ /*9006*/;
assign _9412_ = oneWire & _9411_ /*9004*/;
assign _9377_ = oneWire ^ _9411_ /*9005*/;
assign _9409_ = _9410_ | _9412_ /*9002*/;
assign _9418_ = ~D[1] /*9001*/;
assign _9415_ = _9153_ & _9418_ /*8997*/;
assign _9416_ = _9153_ ^ _9418_ /*9000*/;
assign _9417_ = _9409_ & _9416_ /*8998*/;
assign _9378_ = _9409_ ^ _9416_ /*8999*/;
assign _9414_ = _9415_ | _9417_ /*8996*/;
assign _9423_ = ~D[2] /*8995*/;
assign _9420_ = _9154_ & _9423_ /*8991*/;
assign _9421_ = _9154_ ^ _9423_ /*8994*/;
assign _9422_ = _9414_ & _9421_ /*8992*/;
assign _9379_ = _9414_ ^ _9421_ /*8993*/;
assign _9419_ = _9420_ | _9422_ /*8990*/;
assign _9428_ = ~D[3] /*8989*/;
assign _9425_ = _9155_ & _9428_ /*8985*/;
assign _9426_ = _9155_ ^ _9428_ /*8988*/;
assign _9427_ = _9419_ & _9426_ /*8986*/;
assign _9380_ = _9419_ ^ _9426_ /*8987*/;
assign _9424_ = _9425_ | _9427_ /*8984*/;
assign _9433_ = ~D[4] /*8983*/;
assign _9430_ = _9156_ & _9433_ /*8979*/;
assign _9431_ = _9156_ ^ _9433_ /*8982*/;
assign _9432_ = _9424_ & _9431_ /*8980*/;
assign _9381_ = _9424_ ^ _9431_ /*8981*/;
assign _9429_ = _9430_ | _9432_ /*8978*/;
assign _9438_ = ~D[5] /*8977*/;
assign _9435_ = _9157_ & _9438_ /*8973*/;
assign _9436_ = _9157_ ^ _9438_ /*8976*/;
assign _9437_ = _9429_ & _9436_ /*8974*/;
assign _9382_ = _9429_ ^ _9436_ /*8975*/;
assign _9434_ = _9435_ | _9437_ /*8972*/;
assign _9443_ = ~D[6] /*8971*/;
assign _9440_ = _9158_ & _9443_ /*8967*/;
assign _9441_ = _9158_ ^ _9443_ /*8970*/;
assign _9442_ = _9434_ & _9441_ /*8968*/;
assign _9383_ = _9434_ ^ _9441_ /*8969*/;
assign _9439_ = _9440_ | _9442_ /*8966*/;
assign _9448_ = ~D[7] /*8965*/;
assign _9445_ = _9159_ & _9448_ /*8961*/;
assign _9446_ = _9159_ ^ _9448_ /*8964*/;
assign _9447_ = _9439_ & _9446_ /*8962*/;
assign _9384_ = _9439_ ^ _9446_ /*8963*/;
assign _9444_ = _9445_ | _9447_ /*8960*/;
assign _9453_ = ~D[8] /*8959*/;
assign _9450_ = _9160_ & _9453_ /*8955*/;
assign _9451_ = _9160_ ^ _9453_ /*8958*/;
assign _9452_ = _9444_ & _9451_ /*8956*/;
assign _9385_ = _9444_ ^ _9451_ /*8957*/;
assign _9449_ = _9450_ | _9452_ /*8954*/;
assign _9458_ = ~D[9] /*8953*/;
assign _9455_ = _9161_ & _9458_ /*8949*/;
assign _9456_ = _9161_ ^ _9458_ /*8952*/;
assign _9457_ = _9449_ & _9456_ /*8950*/;
assign _9386_ = _9449_ ^ _9456_ /*8951*/;
assign _9454_ = _9455_ | _9457_ /*8948*/;
assign _9463_ = ~D[10] /*8947*/;
assign _9460_ = _9162_ & _9463_ /*8943*/;
assign _9461_ = _9162_ ^ _9463_ /*8946*/;
assign _9462_ = _9454_ & _9461_ /*8944*/;
assign _9387_ = _9454_ ^ _9461_ /*8945*/;
assign _9459_ = _9460_ | _9462_ /*8942*/;
assign _9468_ = ~D[11] /*8941*/;
assign _9465_ = _9163_ & _9468_ /*8937*/;
assign _9466_ = _9163_ ^ _9468_ /*8940*/;
assign _9467_ = _9459_ & _9466_ /*8938*/;
assign _9388_ = _9459_ ^ _9466_ /*8939*/;
assign _9464_ = _9465_ | _9467_ /*8936*/;
assign _9473_ = ~D[12] /*8935*/;
assign _9470_ = _9164_ & _9473_ /*8931*/;
assign _9471_ = _9164_ ^ _9473_ /*8934*/;
assign _9472_ = _9464_ & _9471_ /*8932*/;
assign _9389_ = _9464_ ^ _9471_ /*8933*/;
assign _9469_ = _9470_ | _9472_ /*8930*/;
assign _9478_ = ~D[13] /*8929*/;
assign _9475_ = _9165_ & _9478_ /*8925*/;
assign _9476_ = _9165_ ^ _9478_ /*8928*/;
assign _9477_ = _9469_ & _9476_ /*8926*/;
assign _9390_ = _9469_ ^ _9476_ /*8927*/;
assign _9474_ = _9475_ | _9477_ /*8924*/;
assign _9483_ = ~D[14] /*8923*/;
assign _9480_ = _9166_ & _9483_ /*8919*/;
assign _9481_ = _9166_ ^ _9483_ /*8922*/;
assign _9482_ = _9474_ & _9481_ /*8920*/;
assign _9391_ = _9474_ ^ _9481_ /*8921*/;
assign _9479_ = _9480_ | _9482_ /*8918*/;
assign _9488_ = ~D[15] /*8917*/;
assign _9485_ = _9167_ & _9488_ /*8913*/;
assign _9486_ = _9167_ ^ _9488_ /*8916*/;
assign _9487_ = _9479_ & _9486_ /*8914*/;
assign _9392_ = _9479_ ^ _9486_ /*8915*/;
assign _9484_ = _9485_ | _9487_ /*8912*/;
assign _9493_ = ~D[16] /*8911*/;
assign _9490_ = _9168_ & _9493_ /*8907*/;
assign _9491_ = _9168_ ^ _9493_ /*8910*/;
assign _9492_ = _9484_ & _9491_ /*8908*/;
assign _9393_ = _9484_ ^ _9491_ /*8909*/;
assign _9489_ = _9490_ | _9492_ /*8906*/;
assign _9498_ = ~D[17] /*8905*/;
assign _9495_ = _9169_ & _9498_ /*8901*/;
assign _9496_ = _9169_ ^ _9498_ /*8904*/;
assign _9497_ = _9489_ & _9496_ /*8902*/;
assign _9394_ = _9489_ ^ _9496_ /*8903*/;
assign _9494_ = _9495_ | _9497_ /*8900*/;
assign _9503_ = ~D[18] /*8899*/;
assign _9500_ = _9170_ & _9503_ /*8895*/;
assign _9501_ = _9170_ ^ _9503_ /*8898*/;
assign _9502_ = _9494_ & _9501_ /*8896*/;
assign _9395_ = _9494_ ^ _9501_ /*8897*/;
assign _9499_ = _9500_ | _9502_ /*8894*/;
assign _9508_ = ~D[19] /*8893*/;
assign _9505_ = _9171_ & _9508_ /*8889*/;
assign _9506_ = _9171_ ^ _9508_ /*8892*/;
assign _9507_ = _9499_ & _9506_ /*8890*/;
assign _9396_ = _9499_ ^ _9506_ /*8891*/;
assign _9504_ = _9505_ | _9507_ /*8888*/;
assign _9513_ = ~D[20] /*8887*/;
assign _9510_ = _9172_ & _9513_ /*8883*/;
assign _9511_ = _9172_ ^ _9513_ /*8886*/;
assign _9512_ = _9504_ & _9511_ /*8884*/;
assign _9397_ = _9504_ ^ _9511_ /*8885*/;
assign _9509_ = _9510_ | _9512_ /*8882*/;
assign _9518_ = ~D[21] /*8881*/;
assign _9515_ = _9173_ & _9518_ /*8877*/;
assign _9516_ = _9173_ ^ _9518_ /*8880*/;
assign _9517_ = _9509_ & _9516_ /*8878*/;
assign _9398_ = _9509_ ^ _9516_ /*8879*/;
assign _9514_ = _9515_ | _9517_ /*8876*/;
assign _9523_ = ~D[22] /*8875*/;
assign _9520_ = _9174_ & _9523_ /*8871*/;
assign _9521_ = _9174_ ^ _9523_ /*8874*/;
assign _9522_ = _9514_ & _9521_ /*8872*/;
assign _9399_ = _9514_ ^ _9521_ /*8873*/;
assign _9519_ = _9520_ | _9522_ /*8870*/;
assign _9528_ = ~D[23] /*8869*/;
assign _9525_ = _9175_ & _9528_ /*8865*/;
assign _9526_ = _9175_ ^ _9528_ /*8868*/;
assign _9527_ = _9519_ & _9526_ /*8866*/;
assign _9400_ = _9519_ ^ _9526_ /*8867*/;
assign _9524_ = _9525_ | _9527_ /*8864*/;
assign _9533_ = ~D[24] /*8863*/;
assign _9530_ = _9176_ & _9533_ /*8859*/;
assign _9531_ = _9176_ ^ _9533_ /*8862*/;
assign _9532_ = _9524_ & _9531_ /*8860*/;
assign _9401_ = _9524_ ^ _9531_ /*8861*/;
assign _9529_ = _9530_ | _9532_ /*8858*/;
assign _9538_ = ~D[25] /*8857*/;
assign _9535_ = _9177_ & _9538_ /*8853*/;
assign _9536_ = _9177_ ^ _9538_ /*8856*/;
assign _9537_ = _9529_ & _9536_ /*8854*/;
assign _9402_ = _9529_ ^ _9536_ /*8855*/;
assign _9534_ = _9535_ | _9537_ /*8852*/;
assign _9543_ = ~D[26] /*8851*/;
assign _9540_ = _9178_ & _9543_ /*8847*/;
assign _9541_ = _9178_ ^ _9543_ /*8850*/;
assign _9542_ = _9534_ & _9541_ /*8848*/;
assign _9403_ = _9534_ ^ _9541_ /*8849*/;
assign _9539_ = _9540_ | _9542_ /*8846*/;
assign _9548_ = ~D[27] /*8845*/;
assign _9545_ = _9179_ & _9548_ /*8841*/;
assign _9546_ = _9179_ ^ _9548_ /*8844*/;
assign _9547_ = _9539_ & _9546_ /*8842*/;
assign _9404_ = _9539_ ^ _9546_ /*8843*/;
assign _9544_ = _9545_ | _9547_ /*8840*/;
assign _9553_ = ~D[28] /*8839*/;
assign _9550_ = _9180_ & _9553_ /*8835*/;
assign _9551_ = _9180_ ^ _9553_ /*8838*/;
assign _9552_ = _9544_ & _9551_ /*8836*/;
assign _9405_ = _9544_ ^ _9551_ /*8837*/;
assign _9549_ = _9550_ | _9552_ /*8834*/;
assign _9558_ = ~D[29] /*8833*/;
assign _9555_ = _9181_ & _9558_ /*8829*/;
assign _9556_ = _9181_ ^ _9558_ /*8832*/;
assign _9557_ = _9549_ & _9556_ /*8830*/;
assign _9406_ = _9549_ ^ _9556_ /*8831*/;
assign _9554_ = _9555_ | _9557_ /*8828*/;
assign _9563_ = ~D[30] /*8827*/;
assign _9560_ = _9182_ & _9563_ /*8823*/;
assign _9561_ = _9182_ ^ _9563_ /*8826*/;
assign _9562_ = _9554_ & _9561_ /*8824*/;
assign _9407_ = _9554_ ^ _9561_ /*8825*/;
assign _9559_ = _9560_ | _9562_ /*8822*/;
assign _9564_ = _9183_ & oneWire /*8817*/;
assign _9565_ = _9183_ ^ oneWire /*8820*/;
assign _9566_ = _9559_ & _9565_ /*8818*/;
assign _9408_ = _9559_ ^ _9565_ /*8819*/;
assign Q[10] = _9564_ | _9566_ /*8816*/;
assign _9635_ = ~Q[10] /*8623*/;
assign _9634_ = _9635_ & D[0] /*8622*/;
assign _9637_ = _9377_ & _9634_ /*8617*/;
assign _9638_ = _9377_ ^ _9634_ /*8620*/;
assign _9639_ = zeroWire & _9638_ /*8618*/;
assign _9601_ = zeroWire ^ _9638_ /*8619*/;
assign _9636_ = _9637_ | _9639_ /*8616*/;
assign _9641_ = ~Q[10] /*8615*/;
assign _9640_ = _9641_ & D[1] /*8614*/;
assign _9643_ = _9378_ & _9640_ /*8609*/;
assign _9644_ = _9378_ ^ _9640_ /*8612*/;
assign _9645_ = _9636_ & _9644_ /*8610*/;
assign _9602_ = _9636_ ^ _9644_ /*8611*/;
assign _9642_ = _9643_ | _9645_ /*8608*/;
assign _9647_ = ~Q[10] /*8607*/;
assign _9646_ = _9647_ & D[2] /*8606*/;
assign _9649_ = _9379_ & _9646_ /*8601*/;
assign _9650_ = _9379_ ^ _9646_ /*8604*/;
assign _9651_ = _9642_ & _9650_ /*8602*/;
assign _9603_ = _9642_ ^ _9650_ /*8603*/;
assign _9648_ = _9649_ | _9651_ /*8600*/;
assign _9653_ = ~Q[10] /*8599*/;
assign _9652_ = _9653_ & D[3] /*8598*/;
assign _9655_ = _9380_ & _9652_ /*8593*/;
assign _9656_ = _9380_ ^ _9652_ /*8596*/;
assign _9657_ = _9648_ & _9656_ /*8594*/;
assign _9604_ = _9648_ ^ _9656_ /*8595*/;
assign _9654_ = _9655_ | _9657_ /*8592*/;
assign _9659_ = ~Q[10] /*8591*/;
assign _9658_ = _9659_ & D[4] /*8590*/;
assign _9661_ = _9381_ & _9658_ /*8585*/;
assign _9662_ = _9381_ ^ _9658_ /*8588*/;
assign _9663_ = _9654_ & _9662_ /*8586*/;
assign _9605_ = _9654_ ^ _9662_ /*8587*/;
assign _9660_ = _9661_ | _9663_ /*8584*/;
assign _9665_ = ~Q[10] /*8583*/;
assign _9664_ = _9665_ & D[5] /*8582*/;
assign _9667_ = _9382_ & _9664_ /*8577*/;
assign _9668_ = _9382_ ^ _9664_ /*8580*/;
assign _9669_ = _9660_ & _9668_ /*8578*/;
assign _9606_ = _9660_ ^ _9668_ /*8579*/;
assign _9666_ = _9667_ | _9669_ /*8576*/;
assign _9671_ = ~Q[10] /*8575*/;
assign _9670_ = _9671_ & D[6] /*8574*/;
assign _9673_ = _9383_ & _9670_ /*8569*/;
assign _9674_ = _9383_ ^ _9670_ /*8572*/;
assign _9675_ = _9666_ & _9674_ /*8570*/;
assign _9607_ = _9666_ ^ _9674_ /*8571*/;
assign _9672_ = _9673_ | _9675_ /*8568*/;
assign _9677_ = ~Q[10] /*8567*/;
assign _9676_ = _9677_ & D[7] /*8566*/;
assign _9679_ = _9384_ & _9676_ /*8561*/;
assign _9680_ = _9384_ ^ _9676_ /*8564*/;
assign _9681_ = _9672_ & _9680_ /*8562*/;
assign _9608_ = _9672_ ^ _9680_ /*8563*/;
assign _9678_ = _9679_ | _9681_ /*8560*/;
assign _9683_ = ~Q[10] /*8559*/;
assign _9682_ = _9683_ & D[8] /*8558*/;
assign _9685_ = _9385_ & _9682_ /*8553*/;
assign _9686_ = _9385_ ^ _9682_ /*8556*/;
assign _9687_ = _9678_ & _9686_ /*8554*/;
assign _9609_ = _9678_ ^ _9686_ /*8555*/;
assign _9684_ = _9685_ | _9687_ /*8552*/;
assign _9689_ = ~Q[10] /*8551*/;
assign _9688_ = _9689_ & D[9] /*8550*/;
assign _9691_ = _9386_ & _9688_ /*8545*/;
assign _9692_ = _9386_ ^ _9688_ /*8548*/;
assign _9693_ = _9684_ & _9692_ /*8546*/;
assign _9610_ = _9684_ ^ _9692_ /*8547*/;
assign _9690_ = _9691_ | _9693_ /*8544*/;
assign _9695_ = ~Q[10] /*8543*/;
assign _9694_ = _9695_ & D[10] /*8542*/;
assign _9697_ = _9387_ & _9694_ /*8537*/;
assign _9698_ = _9387_ ^ _9694_ /*8540*/;
assign _9699_ = _9690_ & _9698_ /*8538*/;
assign _9611_ = _9690_ ^ _9698_ /*8539*/;
assign _9696_ = _9697_ | _9699_ /*8536*/;
assign _9701_ = ~Q[10] /*8535*/;
assign _9700_ = _9701_ & D[11] /*8534*/;
assign _9703_ = _9388_ & _9700_ /*8529*/;
assign _9704_ = _9388_ ^ _9700_ /*8532*/;
assign _9705_ = _9696_ & _9704_ /*8530*/;
assign _9612_ = _9696_ ^ _9704_ /*8531*/;
assign _9702_ = _9703_ | _9705_ /*8528*/;
assign _9707_ = ~Q[10] /*8527*/;
assign _9706_ = _9707_ & D[12] /*8526*/;
assign _9709_ = _9389_ & _9706_ /*8521*/;
assign _9710_ = _9389_ ^ _9706_ /*8524*/;
assign _9711_ = _9702_ & _9710_ /*8522*/;
assign _9613_ = _9702_ ^ _9710_ /*8523*/;
assign _9708_ = _9709_ | _9711_ /*8520*/;
assign _9713_ = ~Q[10] /*8519*/;
assign _9712_ = _9713_ & D[13] /*8518*/;
assign _9715_ = _9390_ & _9712_ /*8513*/;
assign _9716_ = _9390_ ^ _9712_ /*8516*/;
assign _9717_ = _9708_ & _9716_ /*8514*/;
assign _9614_ = _9708_ ^ _9716_ /*8515*/;
assign _9714_ = _9715_ | _9717_ /*8512*/;
assign _9719_ = ~Q[10] /*8511*/;
assign _9718_ = _9719_ & D[14] /*8510*/;
assign _9721_ = _9391_ & _9718_ /*8505*/;
assign _9722_ = _9391_ ^ _9718_ /*8508*/;
assign _9723_ = _9714_ & _9722_ /*8506*/;
assign _9615_ = _9714_ ^ _9722_ /*8507*/;
assign _9720_ = _9721_ | _9723_ /*8504*/;
assign _9725_ = ~Q[10] /*8503*/;
assign _9724_ = _9725_ & D[15] /*8502*/;
assign _9727_ = _9392_ & _9724_ /*8497*/;
assign _9728_ = _9392_ ^ _9724_ /*8500*/;
assign _9729_ = _9720_ & _9728_ /*8498*/;
assign _9616_ = _9720_ ^ _9728_ /*8499*/;
assign _9726_ = _9727_ | _9729_ /*8496*/;
assign _9731_ = ~Q[10] /*8495*/;
assign _9730_ = _9731_ & D[16] /*8494*/;
assign _9733_ = _9393_ & _9730_ /*8489*/;
assign _9734_ = _9393_ ^ _9730_ /*8492*/;
assign _9735_ = _9726_ & _9734_ /*8490*/;
assign _9617_ = _9726_ ^ _9734_ /*8491*/;
assign _9732_ = _9733_ | _9735_ /*8488*/;
assign _9737_ = ~Q[10] /*8487*/;
assign _9736_ = _9737_ & D[17] /*8486*/;
assign _9739_ = _9394_ & _9736_ /*8481*/;
assign _9740_ = _9394_ ^ _9736_ /*8484*/;
assign _9741_ = _9732_ & _9740_ /*8482*/;
assign _9618_ = _9732_ ^ _9740_ /*8483*/;
assign _9738_ = _9739_ | _9741_ /*8480*/;
assign _9743_ = ~Q[10] /*8479*/;
assign _9742_ = _9743_ & D[18] /*8478*/;
assign _9745_ = _9395_ & _9742_ /*8473*/;
assign _9746_ = _9395_ ^ _9742_ /*8476*/;
assign _9747_ = _9738_ & _9746_ /*8474*/;
assign _9619_ = _9738_ ^ _9746_ /*8475*/;
assign _9744_ = _9745_ | _9747_ /*8472*/;
assign _9749_ = ~Q[10] /*8471*/;
assign _9748_ = _9749_ & D[19] /*8470*/;
assign _9751_ = _9396_ & _9748_ /*8465*/;
assign _9752_ = _9396_ ^ _9748_ /*8468*/;
assign _9753_ = _9744_ & _9752_ /*8466*/;
assign _9620_ = _9744_ ^ _9752_ /*8467*/;
assign _9750_ = _9751_ | _9753_ /*8464*/;
assign _9755_ = ~Q[10] /*8463*/;
assign _9754_ = _9755_ & D[20] /*8462*/;
assign _9757_ = _9397_ & _9754_ /*8457*/;
assign _9758_ = _9397_ ^ _9754_ /*8460*/;
assign _9759_ = _9750_ & _9758_ /*8458*/;
assign _9621_ = _9750_ ^ _9758_ /*8459*/;
assign _9756_ = _9757_ | _9759_ /*8456*/;
assign _9761_ = ~Q[10] /*8455*/;
assign _9760_ = _9761_ & D[21] /*8454*/;
assign _9763_ = _9398_ & _9760_ /*8449*/;
assign _9764_ = _9398_ ^ _9760_ /*8452*/;
assign _9765_ = _9756_ & _9764_ /*8450*/;
assign _9622_ = _9756_ ^ _9764_ /*8451*/;
assign _9762_ = _9763_ | _9765_ /*8448*/;
assign _9767_ = ~Q[10] /*8447*/;
assign _9766_ = _9767_ & D[22] /*8446*/;
assign _9769_ = _9399_ & _9766_ /*8441*/;
assign _9770_ = _9399_ ^ _9766_ /*8444*/;
assign _9771_ = _9762_ & _9770_ /*8442*/;
assign _9623_ = _9762_ ^ _9770_ /*8443*/;
assign _9768_ = _9769_ | _9771_ /*8440*/;
assign _9773_ = ~Q[10] /*8439*/;
assign _9772_ = _9773_ & D[23] /*8438*/;
assign _9775_ = _9400_ & _9772_ /*8433*/;
assign _9776_ = _9400_ ^ _9772_ /*8436*/;
assign _9777_ = _9768_ & _9776_ /*8434*/;
assign _9624_ = _9768_ ^ _9776_ /*8435*/;
assign _9774_ = _9775_ | _9777_ /*8432*/;
assign _9779_ = ~Q[10] /*8431*/;
assign _9778_ = _9779_ & D[24] /*8430*/;
assign _9781_ = _9401_ & _9778_ /*8425*/;
assign _9782_ = _9401_ ^ _9778_ /*8428*/;
assign _9783_ = _9774_ & _9782_ /*8426*/;
assign _9625_ = _9774_ ^ _9782_ /*8427*/;
assign _9780_ = _9781_ | _9783_ /*8424*/;
assign _9785_ = ~Q[10] /*8423*/;
assign _9784_ = _9785_ & D[25] /*8422*/;
assign _9787_ = _9402_ & _9784_ /*8417*/;
assign _9788_ = _9402_ ^ _9784_ /*8420*/;
assign _9789_ = _9780_ & _9788_ /*8418*/;
assign _9626_ = _9780_ ^ _9788_ /*8419*/;
assign _9786_ = _9787_ | _9789_ /*8416*/;
assign _9791_ = ~Q[10] /*8415*/;
assign _9790_ = _9791_ & D[26] /*8414*/;
assign _9793_ = _9403_ & _9790_ /*8409*/;
assign _9794_ = _9403_ ^ _9790_ /*8412*/;
assign _9795_ = _9786_ & _9794_ /*8410*/;
assign _9627_ = _9786_ ^ _9794_ /*8411*/;
assign _9792_ = _9793_ | _9795_ /*8408*/;
assign _9797_ = ~Q[10] /*8407*/;
assign _9796_ = _9797_ & D[27] /*8406*/;
assign _9799_ = _9404_ & _9796_ /*8401*/;
assign _9800_ = _9404_ ^ _9796_ /*8404*/;
assign _9801_ = _9792_ & _9800_ /*8402*/;
assign _9628_ = _9792_ ^ _9800_ /*8403*/;
assign _9798_ = _9799_ | _9801_ /*8400*/;
assign _9803_ = ~Q[10] /*8399*/;
assign _9802_ = _9803_ & D[28] /*8398*/;
assign _9805_ = _9405_ & _9802_ /*8393*/;
assign _9806_ = _9405_ ^ _9802_ /*8396*/;
assign _9807_ = _9798_ & _9806_ /*8394*/;
assign _9629_ = _9798_ ^ _9806_ /*8395*/;
assign _9804_ = _9805_ | _9807_ /*8392*/;
assign _9809_ = ~Q[10] /*8391*/;
assign _9808_ = _9809_ & D[29] /*8390*/;
assign _9811_ = _9406_ & _9808_ /*8385*/;
assign _9812_ = _9406_ ^ _9808_ /*8388*/;
assign _9813_ = _9804_ & _9812_ /*8386*/;
assign _9630_ = _9804_ ^ _9812_ /*8387*/;
assign _9810_ = _9811_ | _9813_ /*8384*/;
assign _9815_ = ~Q[10] /*8383*/;
assign _9814_ = _9815_ & D[30] /*8382*/;
assign _9817_ = _9407_ & _9814_ /*8377*/;
assign _9818_ = _9407_ ^ _9814_ /*8380*/;
assign _9819_ = _9810_ & _9818_ /*8378*/;
assign _9631_ = _9810_ ^ _9818_ /*8379*/;
assign _9816_ = _9817_ | _9819_ /*8376*/;
assign _9821_ = ~Q[10] /*8375*/;
assign _9820_ = _9821_ & zeroWire /*8374*/;
assign _9822_ = _9408_ ^ _9820_ /*8372*/;
assign _9632_ = _9822_ ^ _9816_ /*8371*/;
assign _9861_ = ~D[0] /*8245*/;
assign _9858_ = R_0[9] & _9861_ /*8241*/;
assign _9859_ = R_0[9] ^ _9861_ /*8244*/;
assign _9860_ = oneWire & _9859_ /*8242*/;
assign _9825_ = oneWire ^ _9859_ /*8243*/;
assign _9857_ = _9858_ | _9860_ /*8240*/;
assign _9866_ = ~D[1] /*8239*/;
assign _9863_ = _9601_ & _9866_ /*8235*/;
assign _9864_ = _9601_ ^ _9866_ /*8238*/;
assign _9865_ = _9857_ & _9864_ /*8236*/;
assign _9826_ = _9857_ ^ _9864_ /*8237*/;
assign _9862_ = _9863_ | _9865_ /*8234*/;
assign _9871_ = ~D[2] /*8233*/;
assign _9868_ = _9602_ & _9871_ /*8229*/;
assign _9869_ = _9602_ ^ _9871_ /*8232*/;
assign _9870_ = _9862_ & _9869_ /*8230*/;
assign _9827_ = _9862_ ^ _9869_ /*8231*/;
assign _9867_ = _9868_ | _9870_ /*8228*/;
assign _9876_ = ~D[3] /*8227*/;
assign _9873_ = _9603_ & _9876_ /*8223*/;
assign _9874_ = _9603_ ^ _9876_ /*8226*/;
assign _9875_ = _9867_ & _9874_ /*8224*/;
assign _9828_ = _9867_ ^ _9874_ /*8225*/;
assign _9872_ = _9873_ | _9875_ /*8222*/;
assign _9881_ = ~D[4] /*8221*/;
assign _9878_ = _9604_ & _9881_ /*8217*/;
assign _9879_ = _9604_ ^ _9881_ /*8220*/;
assign _9880_ = _9872_ & _9879_ /*8218*/;
assign _9829_ = _9872_ ^ _9879_ /*8219*/;
assign _9877_ = _9878_ | _9880_ /*8216*/;
assign _9886_ = ~D[5] /*8215*/;
assign _9883_ = _9605_ & _9886_ /*8211*/;
assign _9884_ = _9605_ ^ _9886_ /*8214*/;
assign _9885_ = _9877_ & _9884_ /*8212*/;
assign _9830_ = _9877_ ^ _9884_ /*8213*/;
assign _9882_ = _9883_ | _9885_ /*8210*/;
assign _9891_ = ~D[6] /*8209*/;
assign _9888_ = _9606_ & _9891_ /*8205*/;
assign _9889_ = _9606_ ^ _9891_ /*8208*/;
assign _9890_ = _9882_ & _9889_ /*8206*/;
assign _9831_ = _9882_ ^ _9889_ /*8207*/;
assign _9887_ = _9888_ | _9890_ /*8204*/;
assign _9896_ = ~D[7] /*8203*/;
assign _9893_ = _9607_ & _9896_ /*8199*/;
assign _9894_ = _9607_ ^ _9896_ /*8202*/;
assign _9895_ = _9887_ & _9894_ /*8200*/;
assign _9832_ = _9887_ ^ _9894_ /*8201*/;
assign _9892_ = _9893_ | _9895_ /*8198*/;
assign _9901_ = ~D[8] /*8197*/;
assign _9898_ = _9608_ & _9901_ /*8193*/;
assign _9899_ = _9608_ ^ _9901_ /*8196*/;
assign _9900_ = _9892_ & _9899_ /*8194*/;
assign _9833_ = _9892_ ^ _9899_ /*8195*/;
assign _9897_ = _9898_ | _9900_ /*8192*/;
assign _9906_ = ~D[9] /*8191*/;
assign _9903_ = _9609_ & _9906_ /*8187*/;
assign _9904_ = _9609_ ^ _9906_ /*8190*/;
assign _9905_ = _9897_ & _9904_ /*8188*/;
assign _9834_ = _9897_ ^ _9904_ /*8189*/;
assign _9902_ = _9903_ | _9905_ /*8186*/;
assign _9911_ = ~D[10] /*8185*/;
assign _9908_ = _9610_ & _9911_ /*8181*/;
assign _9909_ = _9610_ ^ _9911_ /*8184*/;
assign _9910_ = _9902_ & _9909_ /*8182*/;
assign _9835_ = _9902_ ^ _9909_ /*8183*/;
assign _9907_ = _9908_ | _9910_ /*8180*/;
assign _9916_ = ~D[11] /*8179*/;
assign _9913_ = _9611_ & _9916_ /*8175*/;
assign _9914_ = _9611_ ^ _9916_ /*8178*/;
assign _9915_ = _9907_ & _9914_ /*8176*/;
assign _9836_ = _9907_ ^ _9914_ /*8177*/;
assign _9912_ = _9913_ | _9915_ /*8174*/;
assign _9921_ = ~D[12] /*8173*/;
assign _9918_ = _9612_ & _9921_ /*8169*/;
assign _9919_ = _9612_ ^ _9921_ /*8172*/;
assign _9920_ = _9912_ & _9919_ /*8170*/;
assign _9837_ = _9912_ ^ _9919_ /*8171*/;
assign _9917_ = _9918_ | _9920_ /*8168*/;
assign _9926_ = ~D[13] /*8167*/;
assign _9923_ = _9613_ & _9926_ /*8163*/;
assign _9924_ = _9613_ ^ _9926_ /*8166*/;
assign _9925_ = _9917_ & _9924_ /*8164*/;
assign _9838_ = _9917_ ^ _9924_ /*8165*/;
assign _9922_ = _9923_ | _9925_ /*8162*/;
assign _9931_ = ~D[14] /*8161*/;
assign _9928_ = _9614_ & _9931_ /*8157*/;
assign _9929_ = _9614_ ^ _9931_ /*8160*/;
assign _9930_ = _9922_ & _9929_ /*8158*/;
assign _9839_ = _9922_ ^ _9929_ /*8159*/;
assign _9927_ = _9928_ | _9930_ /*8156*/;
assign _9936_ = ~D[15] /*8155*/;
assign _9933_ = _9615_ & _9936_ /*8151*/;
assign _9934_ = _9615_ ^ _9936_ /*8154*/;
assign _9935_ = _9927_ & _9934_ /*8152*/;
assign _9840_ = _9927_ ^ _9934_ /*8153*/;
assign _9932_ = _9933_ | _9935_ /*8150*/;
assign _9941_ = ~D[16] /*8149*/;
assign _9938_ = _9616_ & _9941_ /*8145*/;
assign _9939_ = _9616_ ^ _9941_ /*8148*/;
assign _9940_ = _9932_ & _9939_ /*8146*/;
assign _9841_ = _9932_ ^ _9939_ /*8147*/;
assign _9937_ = _9938_ | _9940_ /*8144*/;
assign _9946_ = ~D[17] /*8143*/;
assign _9943_ = _9617_ & _9946_ /*8139*/;
assign _9944_ = _9617_ ^ _9946_ /*8142*/;
assign _9945_ = _9937_ & _9944_ /*8140*/;
assign _9842_ = _9937_ ^ _9944_ /*8141*/;
assign _9942_ = _9943_ | _9945_ /*8138*/;
assign _9951_ = ~D[18] /*8137*/;
assign _9948_ = _9618_ & _9951_ /*8133*/;
assign _9949_ = _9618_ ^ _9951_ /*8136*/;
assign _9950_ = _9942_ & _9949_ /*8134*/;
assign _9843_ = _9942_ ^ _9949_ /*8135*/;
assign _9947_ = _9948_ | _9950_ /*8132*/;
assign _9956_ = ~D[19] /*8131*/;
assign _9953_ = _9619_ & _9956_ /*8127*/;
assign _9954_ = _9619_ ^ _9956_ /*8130*/;
assign _9955_ = _9947_ & _9954_ /*8128*/;
assign _9844_ = _9947_ ^ _9954_ /*8129*/;
assign _9952_ = _9953_ | _9955_ /*8126*/;
assign _9961_ = ~D[20] /*8125*/;
assign _9958_ = _9620_ & _9961_ /*8121*/;
assign _9959_ = _9620_ ^ _9961_ /*8124*/;
assign _9960_ = _9952_ & _9959_ /*8122*/;
assign _9845_ = _9952_ ^ _9959_ /*8123*/;
assign _9957_ = _9958_ | _9960_ /*8120*/;
assign _9966_ = ~D[21] /*8119*/;
assign _9963_ = _9621_ & _9966_ /*8115*/;
assign _9964_ = _9621_ ^ _9966_ /*8118*/;
assign _9965_ = _9957_ & _9964_ /*8116*/;
assign _9846_ = _9957_ ^ _9964_ /*8117*/;
assign _9962_ = _9963_ | _9965_ /*8114*/;
assign _9971_ = ~D[22] /*8113*/;
assign _9968_ = _9622_ & _9971_ /*8109*/;
assign _9969_ = _9622_ ^ _9971_ /*8112*/;
assign _9970_ = _9962_ & _9969_ /*8110*/;
assign _9847_ = _9962_ ^ _9969_ /*8111*/;
assign _9967_ = _9968_ | _9970_ /*8108*/;
assign _9976_ = ~D[23] /*8107*/;
assign _9973_ = _9623_ & _9976_ /*8103*/;
assign _9974_ = _9623_ ^ _9976_ /*8106*/;
assign _9975_ = _9967_ & _9974_ /*8104*/;
assign _9848_ = _9967_ ^ _9974_ /*8105*/;
assign _9972_ = _9973_ | _9975_ /*8102*/;
assign _9981_ = ~D[24] /*8101*/;
assign _9978_ = _9624_ & _9981_ /*8097*/;
assign _9979_ = _9624_ ^ _9981_ /*8100*/;
assign _9980_ = _9972_ & _9979_ /*8098*/;
assign _9849_ = _9972_ ^ _9979_ /*8099*/;
assign _9977_ = _9978_ | _9980_ /*8096*/;
assign _9986_ = ~D[25] /*8095*/;
assign _9983_ = _9625_ & _9986_ /*8091*/;
assign _9984_ = _9625_ ^ _9986_ /*8094*/;
assign _9985_ = _9977_ & _9984_ /*8092*/;
assign _9850_ = _9977_ ^ _9984_ /*8093*/;
assign _9982_ = _9983_ | _9985_ /*8090*/;
assign _9991_ = ~D[26] /*8089*/;
assign _9988_ = _9626_ & _9991_ /*8085*/;
assign _9989_ = _9626_ ^ _9991_ /*8088*/;
assign _9990_ = _9982_ & _9989_ /*8086*/;
assign _9851_ = _9982_ ^ _9989_ /*8087*/;
assign _9987_ = _9988_ | _9990_ /*8084*/;
assign _9996_ = ~D[27] /*8083*/;
assign _9993_ = _9627_ & _9996_ /*8079*/;
assign _9994_ = _9627_ ^ _9996_ /*8082*/;
assign _9995_ = _9987_ & _9994_ /*8080*/;
assign _9852_ = _9987_ ^ _9994_ /*8081*/;
assign _9992_ = _9993_ | _9995_ /*8078*/;
assign _10001_ = ~D[28] /*8077*/;
assign _9998_ = _9628_ & _10001_ /*8073*/;
assign _9999_ = _9628_ ^ _10001_ /*8076*/;
assign _10000_ = _9992_ & _9999_ /*8074*/;
assign _9853_ = _9992_ ^ _9999_ /*8075*/;
assign _9997_ = _9998_ | _10000_ /*8072*/;
assign _10006_ = ~D[29] /*8071*/;
assign _10003_ = _9629_ & _10006_ /*8067*/;
assign _10004_ = _9629_ ^ _10006_ /*8070*/;
assign _10005_ = _9997_ & _10004_ /*8068*/;
assign _9854_ = _9997_ ^ _10004_ /*8069*/;
assign _10002_ = _10003_ | _10005_ /*8066*/;
assign _10011_ = ~D[30] /*8065*/;
assign _10008_ = _9630_ & _10011_ /*8061*/;
assign _10009_ = _9630_ ^ _10011_ /*8064*/;
assign _10010_ = _10002_ & _10009_ /*8062*/;
assign _9855_ = _10002_ ^ _10009_ /*8063*/;
assign _10007_ = _10008_ | _10010_ /*8060*/;
assign _10012_ = _9631_ & oneWire /*8055*/;
assign _10013_ = _9631_ ^ oneWire /*8058*/;
assign _10014_ = _10007_ & _10013_ /*8056*/;
assign _9856_ = _10007_ ^ _10013_ /*8057*/;
assign Q[9] = _10012_ | _10014_ /*8054*/;
assign _10083_ = ~Q[9] /*7861*/;
assign _10082_ = _10083_ & D[0] /*7860*/;
assign _10085_ = _9825_ & _10082_ /*7855*/;
assign _10086_ = _9825_ ^ _10082_ /*7858*/;
assign _10087_ = zeroWire & _10086_ /*7856*/;
assign _10049_ = zeroWire ^ _10086_ /*7857*/;
assign _10084_ = _10085_ | _10087_ /*7854*/;
assign _10089_ = ~Q[9] /*7853*/;
assign _10088_ = _10089_ & D[1] /*7852*/;
assign _10091_ = _9826_ & _10088_ /*7847*/;
assign _10092_ = _9826_ ^ _10088_ /*7850*/;
assign _10093_ = _10084_ & _10092_ /*7848*/;
assign _10050_ = _10084_ ^ _10092_ /*7849*/;
assign _10090_ = _10091_ | _10093_ /*7846*/;
assign _10095_ = ~Q[9] /*7845*/;
assign _10094_ = _10095_ & D[2] /*7844*/;
assign _10097_ = _9827_ & _10094_ /*7839*/;
assign _10098_ = _9827_ ^ _10094_ /*7842*/;
assign _10099_ = _10090_ & _10098_ /*7840*/;
assign _10051_ = _10090_ ^ _10098_ /*7841*/;
assign _10096_ = _10097_ | _10099_ /*7838*/;
assign _10101_ = ~Q[9] /*7837*/;
assign _10100_ = _10101_ & D[3] /*7836*/;
assign _10103_ = _9828_ & _10100_ /*7831*/;
assign _10104_ = _9828_ ^ _10100_ /*7834*/;
assign _10105_ = _10096_ & _10104_ /*7832*/;
assign _10052_ = _10096_ ^ _10104_ /*7833*/;
assign _10102_ = _10103_ | _10105_ /*7830*/;
assign _10107_ = ~Q[9] /*7829*/;
assign _10106_ = _10107_ & D[4] /*7828*/;
assign _10109_ = _9829_ & _10106_ /*7823*/;
assign _10110_ = _9829_ ^ _10106_ /*7826*/;
assign _10111_ = _10102_ & _10110_ /*7824*/;
assign _10053_ = _10102_ ^ _10110_ /*7825*/;
assign _10108_ = _10109_ | _10111_ /*7822*/;
assign _10113_ = ~Q[9] /*7821*/;
assign _10112_ = _10113_ & D[5] /*7820*/;
assign _10115_ = _9830_ & _10112_ /*7815*/;
assign _10116_ = _9830_ ^ _10112_ /*7818*/;
assign _10117_ = _10108_ & _10116_ /*7816*/;
assign _10054_ = _10108_ ^ _10116_ /*7817*/;
assign _10114_ = _10115_ | _10117_ /*7814*/;
assign _10119_ = ~Q[9] /*7813*/;
assign _10118_ = _10119_ & D[6] /*7812*/;
assign _10121_ = _9831_ & _10118_ /*7807*/;
assign _10122_ = _9831_ ^ _10118_ /*7810*/;
assign _10123_ = _10114_ & _10122_ /*7808*/;
assign _10055_ = _10114_ ^ _10122_ /*7809*/;
assign _10120_ = _10121_ | _10123_ /*7806*/;
assign _10125_ = ~Q[9] /*7805*/;
assign _10124_ = _10125_ & D[7] /*7804*/;
assign _10127_ = _9832_ & _10124_ /*7799*/;
assign _10128_ = _9832_ ^ _10124_ /*7802*/;
assign _10129_ = _10120_ & _10128_ /*7800*/;
assign _10056_ = _10120_ ^ _10128_ /*7801*/;
assign _10126_ = _10127_ | _10129_ /*7798*/;
assign _10131_ = ~Q[9] /*7797*/;
assign _10130_ = _10131_ & D[8] /*7796*/;
assign _10133_ = _9833_ & _10130_ /*7791*/;
assign _10134_ = _9833_ ^ _10130_ /*7794*/;
assign _10135_ = _10126_ & _10134_ /*7792*/;
assign _10057_ = _10126_ ^ _10134_ /*7793*/;
assign _10132_ = _10133_ | _10135_ /*7790*/;
assign _10137_ = ~Q[9] /*7789*/;
assign _10136_ = _10137_ & D[9] /*7788*/;
assign _10139_ = _9834_ & _10136_ /*7783*/;
assign _10140_ = _9834_ ^ _10136_ /*7786*/;
assign _10141_ = _10132_ & _10140_ /*7784*/;
assign _10058_ = _10132_ ^ _10140_ /*7785*/;
assign _10138_ = _10139_ | _10141_ /*7782*/;
assign _10143_ = ~Q[9] /*7781*/;
assign _10142_ = _10143_ & D[10] /*7780*/;
assign _10145_ = _9835_ & _10142_ /*7775*/;
assign _10146_ = _9835_ ^ _10142_ /*7778*/;
assign _10147_ = _10138_ & _10146_ /*7776*/;
assign _10059_ = _10138_ ^ _10146_ /*7777*/;
assign _10144_ = _10145_ | _10147_ /*7774*/;
assign _10149_ = ~Q[9] /*7773*/;
assign _10148_ = _10149_ & D[11] /*7772*/;
assign _10151_ = _9836_ & _10148_ /*7767*/;
assign _10152_ = _9836_ ^ _10148_ /*7770*/;
assign _10153_ = _10144_ & _10152_ /*7768*/;
assign _10060_ = _10144_ ^ _10152_ /*7769*/;
assign _10150_ = _10151_ | _10153_ /*7766*/;
assign _10155_ = ~Q[9] /*7765*/;
assign _10154_ = _10155_ & D[12] /*7764*/;
assign _10157_ = _9837_ & _10154_ /*7759*/;
assign _10158_ = _9837_ ^ _10154_ /*7762*/;
assign _10159_ = _10150_ & _10158_ /*7760*/;
assign _10061_ = _10150_ ^ _10158_ /*7761*/;
assign _10156_ = _10157_ | _10159_ /*7758*/;
assign _10161_ = ~Q[9] /*7757*/;
assign _10160_ = _10161_ & D[13] /*7756*/;
assign _10163_ = _9838_ & _10160_ /*7751*/;
assign _10164_ = _9838_ ^ _10160_ /*7754*/;
assign _10165_ = _10156_ & _10164_ /*7752*/;
assign _10062_ = _10156_ ^ _10164_ /*7753*/;
assign _10162_ = _10163_ | _10165_ /*7750*/;
assign _10167_ = ~Q[9] /*7749*/;
assign _10166_ = _10167_ & D[14] /*7748*/;
assign _10169_ = _9839_ & _10166_ /*7743*/;
assign _10170_ = _9839_ ^ _10166_ /*7746*/;
assign _10171_ = _10162_ & _10170_ /*7744*/;
assign _10063_ = _10162_ ^ _10170_ /*7745*/;
assign _10168_ = _10169_ | _10171_ /*7742*/;
assign _10173_ = ~Q[9] /*7741*/;
assign _10172_ = _10173_ & D[15] /*7740*/;
assign _10175_ = _9840_ & _10172_ /*7735*/;
assign _10176_ = _9840_ ^ _10172_ /*7738*/;
assign _10177_ = _10168_ & _10176_ /*7736*/;
assign _10064_ = _10168_ ^ _10176_ /*7737*/;
assign _10174_ = _10175_ | _10177_ /*7734*/;
assign _10179_ = ~Q[9] /*7733*/;
assign _10178_ = _10179_ & D[16] /*7732*/;
assign _10181_ = _9841_ & _10178_ /*7727*/;
assign _10182_ = _9841_ ^ _10178_ /*7730*/;
assign _10183_ = _10174_ & _10182_ /*7728*/;
assign _10065_ = _10174_ ^ _10182_ /*7729*/;
assign _10180_ = _10181_ | _10183_ /*7726*/;
assign _10185_ = ~Q[9] /*7725*/;
assign _10184_ = _10185_ & D[17] /*7724*/;
assign _10187_ = _9842_ & _10184_ /*7719*/;
assign _10188_ = _9842_ ^ _10184_ /*7722*/;
assign _10189_ = _10180_ & _10188_ /*7720*/;
assign _10066_ = _10180_ ^ _10188_ /*7721*/;
assign _10186_ = _10187_ | _10189_ /*7718*/;
assign _10191_ = ~Q[9] /*7717*/;
assign _10190_ = _10191_ & D[18] /*7716*/;
assign _10193_ = _9843_ & _10190_ /*7711*/;
assign _10194_ = _9843_ ^ _10190_ /*7714*/;
assign _10195_ = _10186_ & _10194_ /*7712*/;
assign _10067_ = _10186_ ^ _10194_ /*7713*/;
assign _10192_ = _10193_ | _10195_ /*7710*/;
assign _10197_ = ~Q[9] /*7709*/;
assign _10196_ = _10197_ & D[19] /*7708*/;
assign _10199_ = _9844_ & _10196_ /*7703*/;
assign _10200_ = _9844_ ^ _10196_ /*7706*/;
assign _10201_ = _10192_ & _10200_ /*7704*/;
assign _10068_ = _10192_ ^ _10200_ /*7705*/;
assign _10198_ = _10199_ | _10201_ /*7702*/;
assign _10203_ = ~Q[9] /*7701*/;
assign _10202_ = _10203_ & D[20] /*7700*/;
assign _10205_ = _9845_ & _10202_ /*7695*/;
assign _10206_ = _9845_ ^ _10202_ /*7698*/;
assign _10207_ = _10198_ & _10206_ /*7696*/;
assign _10069_ = _10198_ ^ _10206_ /*7697*/;
assign _10204_ = _10205_ | _10207_ /*7694*/;
assign _10209_ = ~Q[9] /*7693*/;
assign _10208_ = _10209_ & D[21] /*7692*/;
assign _10211_ = _9846_ & _10208_ /*7687*/;
assign _10212_ = _9846_ ^ _10208_ /*7690*/;
assign _10213_ = _10204_ & _10212_ /*7688*/;
assign _10070_ = _10204_ ^ _10212_ /*7689*/;
assign _10210_ = _10211_ | _10213_ /*7686*/;
assign _10215_ = ~Q[9] /*7685*/;
assign _10214_ = _10215_ & D[22] /*7684*/;
assign _10217_ = _9847_ & _10214_ /*7679*/;
assign _10218_ = _9847_ ^ _10214_ /*7682*/;
assign _10219_ = _10210_ & _10218_ /*7680*/;
assign _10071_ = _10210_ ^ _10218_ /*7681*/;
assign _10216_ = _10217_ | _10219_ /*7678*/;
assign _10221_ = ~Q[9] /*7677*/;
assign _10220_ = _10221_ & D[23] /*7676*/;
assign _10223_ = _9848_ & _10220_ /*7671*/;
assign _10224_ = _9848_ ^ _10220_ /*7674*/;
assign _10225_ = _10216_ & _10224_ /*7672*/;
assign _10072_ = _10216_ ^ _10224_ /*7673*/;
assign _10222_ = _10223_ | _10225_ /*7670*/;
assign _10227_ = ~Q[9] /*7669*/;
assign _10226_ = _10227_ & D[24] /*7668*/;
assign _10229_ = _9849_ & _10226_ /*7663*/;
assign _10230_ = _9849_ ^ _10226_ /*7666*/;
assign _10231_ = _10222_ & _10230_ /*7664*/;
assign _10073_ = _10222_ ^ _10230_ /*7665*/;
assign _10228_ = _10229_ | _10231_ /*7662*/;
assign _10233_ = ~Q[9] /*7661*/;
assign _10232_ = _10233_ & D[25] /*7660*/;
assign _10235_ = _9850_ & _10232_ /*7655*/;
assign _10236_ = _9850_ ^ _10232_ /*7658*/;
assign _10237_ = _10228_ & _10236_ /*7656*/;
assign _10074_ = _10228_ ^ _10236_ /*7657*/;
assign _10234_ = _10235_ | _10237_ /*7654*/;
assign _10239_ = ~Q[9] /*7653*/;
assign _10238_ = _10239_ & D[26] /*7652*/;
assign _10241_ = _9851_ & _10238_ /*7647*/;
assign _10242_ = _9851_ ^ _10238_ /*7650*/;
assign _10243_ = _10234_ & _10242_ /*7648*/;
assign _10075_ = _10234_ ^ _10242_ /*7649*/;
assign _10240_ = _10241_ | _10243_ /*7646*/;
assign _10245_ = ~Q[9] /*7645*/;
assign _10244_ = _10245_ & D[27] /*7644*/;
assign _10247_ = _9852_ & _10244_ /*7639*/;
assign _10248_ = _9852_ ^ _10244_ /*7642*/;
assign _10249_ = _10240_ & _10248_ /*7640*/;
assign _10076_ = _10240_ ^ _10248_ /*7641*/;
assign _10246_ = _10247_ | _10249_ /*7638*/;
assign _10251_ = ~Q[9] /*7637*/;
assign _10250_ = _10251_ & D[28] /*7636*/;
assign _10253_ = _9853_ & _10250_ /*7631*/;
assign _10254_ = _9853_ ^ _10250_ /*7634*/;
assign _10255_ = _10246_ & _10254_ /*7632*/;
assign _10077_ = _10246_ ^ _10254_ /*7633*/;
assign _10252_ = _10253_ | _10255_ /*7630*/;
assign _10257_ = ~Q[9] /*7629*/;
assign _10256_ = _10257_ & D[29] /*7628*/;
assign _10259_ = _9854_ & _10256_ /*7623*/;
assign _10260_ = _9854_ ^ _10256_ /*7626*/;
assign _10261_ = _10252_ & _10260_ /*7624*/;
assign _10078_ = _10252_ ^ _10260_ /*7625*/;
assign _10258_ = _10259_ | _10261_ /*7622*/;
assign _10263_ = ~Q[9] /*7621*/;
assign _10262_ = _10263_ & D[30] /*7620*/;
assign _10265_ = _9855_ & _10262_ /*7615*/;
assign _10266_ = _9855_ ^ _10262_ /*7618*/;
assign _10267_ = _10258_ & _10266_ /*7616*/;
assign _10079_ = _10258_ ^ _10266_ /*7617*/;
assign _10264_ = _10265_ | _10267_ /*7614*/;
assign _10269_ = ~Q[9] /*7613*/;
assign _10268_ = _10269_ & zeroWire /*7612*/;
assign _10270_ = _9856_ ^ _10268_ /*7610*/;
assign _10080_ = _10270_ ^ _10264_ /*7609*/;
assign _10309_ = ~D[0] /*7483*/;
assign _10306_ = R_0[8] & _10309_ /*7479*/;
assign _10307_ = R_0[8] ^ _10309_ /*7482*/;
assign _10308_ = oneWire & _10307_ /*7480*/;
assign _10273_ = oneWire ^ _10307_ /*7481*/;
assign _10305_ = _10306_ | _10308_ /*7478*/;
assign _10314_ = ~D[1] /*7477*/;
assign _10311_ = _10049_ & _10314_ /*7473*/;
assign _10312_ = _10049_ ^ _10314_ /*7476*/;
assign _10313_ = _10305_ & _10312_ /*7474*/;
assign _10274_ = _10305_ ^ _10312_ /*7475*/;
assign _10310_ = _10311_ | _10313_ /*7472*/;
assign _10319_ = ~D[2] /*7471*/;
assign _10316_ = _10050_ & _10319_ /*7467*/;
assign _10317_ = _10050_ ^ _10319_ /*7470*/;
assign _10318_ = _10310_ & _10317_ /*7468*/;
assign _10275_ = _10310_ ^ _10317_ /*7469*/;
assign _10315_ = _10316_ | _10318_ /*7466*/;
assign _10324_ = ~D[3] /*7465*/;
assign _10321_ = _10051_ & _10324_ /*7461*/;
assign _10322_ = _10051_ ^ _10324_ /*7464*/;
assign _10323_ = _10315_ & _10322_ /*7462*/;
assign _10276_ = _10315_ ^ _10322_ /*7463*/;
assign _10320_ = _10321_ | _10323_ /*7460*/;
assign _10329_ = ~D[4] /*7459*/;
assign _10326_ = _10052_ & _10329_ /*7455*/;
assign _10327_ = _10052_ ^ _10329_ /*7458*/;
assign _10328_ = _10320_ & _10327_ /*7456*/;
assign _10277_ = _10320_ ^ _10327_ /*7457*/;
assign _10325_ = _10326_ | _10328_ /*7454*/;
assign _10334_ = ~D[5] /*7453*/;
assign _10331_ = _10053_ & _10334_ /*7449*/;
assign _10332_ = _10053_ ^ _10334_ /*7452*/;
assign _10333_ = _10325_ & _10332_ /*7450*/;
assign _10278_ = _10325_ ^ _10332_ /*7451*/;
assign _10330_ = _10331_ | _10333_ /*7448*/;
assign _10339_ = ~D[6] /*7447*/;
assign _10336_ = _10054_ & _10339_ /*7443*/;
assign _10337_ = _10054_ ^ _10339_ /*7446*/;
assign _10338_ = _10330_ & _10337_ /*7444*/;
assign _10279_ = _10330_ ^ _10337_ /*7445*/;
assign _10335_ = _10336_ | _10338_ /*7442*/;
assign _10344_ = ~D[7] /*7441*/;
assign _10341_ = _10055_ & _10344_ /*7437*/;
assign _10342_ = _10055_ ^ _10344_ /*7440*/;
assign _10343_ = _10335_ & _10342_ /*7438*/;
assign _10280_ = _10335_ ^ _10342_ /*7439*/;
assign _10340_ = _10341_ | _10343_ /*7436*/;
assign _10349_ = ~D[8] /*7435*/;
assign _10346_ = _10056_ & _10349_ /*7431*/;
assign _10347_ = _10056_ ^ _10349_ /*7434*/;
assign _10348_ = _10340_ & _10347_ /*7432*/;
assign _10281_ = _10340_ ^ _10347_ /*7433*/;
assign _10345_ = _10346_ | _10348_ /*7430*/;
assign _10354_ = ~D[9] /*7429*/;
assign _10351_ = _10057_ & _10354_ /*7425*/;
assign _10352_ = _10057_ ^ _10354_ /*7428*/;
assign _10353_ = _10345_ & _10352_ /*7426*/;
assign _10282_ = _10345_ ^ _10352_ /*7427*/;
assign _10350_ = _10351_ | _10353_ /*7424*/;
assign _10359_ = ~D[10] /*7423*/;
assign _10356_ = _10058_ & _10359_ /*7419*/;
assign _10357_ = _10058_ ^ _10359_ /*7422*/;
assign _10358_ = _10350_ & _10357_ /*7420*/;
assign _10283_ = _10350_ ^ _10357_ /*7421*/;
assign _10355_ = _10356_ | _10358_ /*7418*/;
assign _10364_ = ~D[11] /*7417*/;
assign _10361_ = _10059_ & _10364_ /*7413*/;
assign _10362_ = _10059_ ^ _10364_ /*7416*/;
assign _10363_ = _10355_ & _10362_ /*7414*/;
assign _10284_ = _10355_ ^ _10362_ /*7415*/;
assign _10360_ = _10361_ | _10363_ /*7412*/;
assign _10369_ = ~D[12] /*7411*/;
assign _10366_ = _10060_ & _10369_ /*7407*/;
assign _10367_ = _10060_ ^ _10369_ /*7410*/;
assign _10368_ = _10360_ & _10367_ /*7408*/;
assign _10285_ = _10360_ ^ _10367_ /*7409*/;
assign _10365_ = _10366_ | _10368_ /*7406*/;
assign _10374_ = ~D[13] /*7405*/;
assign _10371_ = _10061_ & _10374_ /*7401*/;
assign _10372_ = _10061_ ^ _10374_ /*7404*/;
assign _10373_ = _10365_ & _10372_ /*7402*/;
assign _10286_ = _10365_ ^ _10372_ /*7403*/;
assign _10370_ = _10371_ | _10373_ /*7400*/;
assign _10379_ = ~D[14] /*7399*/;
assign _10376_ = _10062_ & _10379_ /*7395*/;
assign _10377_ = _10062_ ^ _10379_ /*7398*/;
assign _10378_ = _10370_ & _10377_ /*7396*/;
assign _10287_ = _10370_ ^ _10377_ /*7397*/;
assign _10375_ = _10376_ | _10378_ /*7394*/;
assign _10384_ = ~D[15] /*7393*/;
assign _10381_ = _10063_ & _10384_ /*7389*/;
assign _10382_ = _10063_ ^ _10384_ /*7392*/;
assign _10383_ = _10375_ & _10382_ /*7390*/;
assign _10288_ = _10375_ ^ _10382_ /*7391*/;
assign _10380_ = _10381_ | _10383_ /*7388*/;
assign _10389_ = ~D[16] /*7387*/;
assign _10386_ = _10064_ & _10389_ /*7383*/;
assign _10387_ = _10064_ ^ _10389_ /*7386*/;
assign _10388_ = _10380_ & _10387_ /*7384*/;
assign _10289_ = _10380_ ^ _10387_ /*7385*/;
assign _10385_ = _10386_ | _10388_ /*7382*/;
assign _10394_ = ~D[17] /*7381*/;
assign _10391_ = _10065_ & _10394_ /*7377*/;
assign _10392_ = _10065_ ^ _10394_ /*7380*/;
assign _10393_ = _10385_ & _10392_ /*7378*/;
assign _10290_ = _10385_ ^ _10392_ /*7379*/;
assign _10390_ = _10391_ | _10393_ /*7376*/;
assign _10399_ = ~D[18] /*7375*/;
assign _10396_ = _10066_ & _10399_ /*7371*/;
assign _10397_ = _10066_ ^ _10399_ /*7374*/;
assign _10398_ = _10390_ & _10397_ /*7372*/;
assign _10291_ = _10390_ ^ _10397_ /*7373*/;
assign _10395_ = _10396_ | _10398_ /*7370*/;
assign _10404_ = ~D[19] /*7369*/;
assign _10401_ = _10067_ & _10404_ /*7365*/;
assign _10402_ = _10067_ ^ _10404_ /*7368*/;
assign _10403_ = _10395_ & _10402_ /*7366*/;
assign _10292_ = _10395_ ^ _10402_ /*7367*/;
assign _10400_ = _10401_ | _10403_ /*7364*/;
assign _10409_ = ~D[20] /*7363*/;
assign _10406_ = _10068_ & _10409_ /*7359*/;
assign _10407_ = _10068_ ^ _10409_ /*7362*/;
assign _10408_ = _10400_ & _10407_ /*7360*/;
assign _10293_ = _10400_ ^ _10407_ /*7361*/;
assign _10405_ = _10406_ | _10408_ /*7358*/;
assign _10414_ = ~D[21] /*7357*/;
assign _10411_ = _10069_ & _10414_ /*7353*/;
assign _10412_ = _10069_ ^ _10414_ /*7356*/;
assign _10413_ = _10405_ & _10412_ /*7354*/;
assign _10294_ = _10405_ ^ _10412_ /*7355*/;
assign _10410_ = _10411_ | _10413_ /*7352*/;
assign _10419_ = ~D[22] /*7351*/;
assign _10416_ = _10070_ & _10419_ /*7347*/;
assign _10417_ = _10070_ ^ _10419_ /*7350*/;
assign _10418_ = _10410_ & _10417_ /*7348*/;
assign _10295_ = _10410_ ^ _10417_ /*7349*/;
assign _10415_ = _10416_ | _10418_ /*7346*/;
assign _10424_ = ~D[23] /*7345*/;
assign _10421_ = _10071_ & _10424_ /*7341*/;
assign _10422_ = _10071_ ^ _10424_ /*7344*/;
assign _10423_ = _10415_ & _10422_ /*7342*/;
assign _10296_ = _10415_ ^ _10422_ /*7343*/;
assign _10420_ = _10421_ | _10423_ /*7340*/;
assign _10429_ = ~D[24] /*7339*/;
assign _10426_ = _10072_ & _10429_ /*7335*/;
assign _10427_ = _10072_ ^ _10429_ /*7338*/;
assign _10428_ = _10420_ & _10427_ /*7336*/;
assign _10297_ = _10420_ ^ _10427_ /*7337*/;
assign _10425_ = _10426_ | _10428_ /*7334*/;
assign _10434_ = ~D[25] /*7333*/;
assign _10431_ = _10073_ & _10434_ /*7329*/;
assign _10432_ = _10073_ ^ _10434_ /*7332*/;
assign _10433_ = _10425_ & _10432_ /*7330*/;
assign _10298_ = _10425_ ^ _10432_ /*7331*/;
assign _10430_ = _10431_ | _10433_ /*7328*/;
assign _10439_ = ~D[26] /*7327*/;
assign _10436_ = _10074_ & _10439_ /*7323*/;
assign _10437_ = _10074_ ^ _10439_ /*7326*/;
assign _10438_ = _10430_ & _10437_ /*7324*/;
assign _10299_ = _10430_ ^ _10437_ /*7325*/;
assign _10435_ = _10436_ | _10438_ /*7322*/;
assign _10444_ = ~D[27] /*7321*/;
assign _10441_ = _10075_ & _10444_ /*7317*/;
assign _10442_ = _10075_ ^ _10444_ /*7320*/;
assign _10443_ = _10435_ & _10442_ /*7318*/;
assign _10300_ = _10435_ ^ _10442_ /*7319*/;
assign _10440_ = _10441_ | _10443_ /*7316*/;
assign _10449_ = ~D[28] /*7315*/;
assign _10446_ = _10076_ & _10449_ /*7311*/;
assign _10447_ = _10076_ ^ _10449_ /*7314*/;
assign _10448_ = _10440_ & _10447_ /*7312*/;
assign _10301_ = _10440_ ^ _10447_ /*7313*/;
assign _10445_ = _10446_ | _10448_ /*7310*/;
assign _10454_ = ~D[29] /*7309*/;
assign _10451_ = _10077_ & _10454_ /*7305*/;
assign _10452_ = _10077_ ^ _10454_ /*7308*/;
assign _10453_ = _10445_ & _10452_ /*7306*/;
assign _10302_ = _10445_ ^ _10452_ /*7307*/;
assign _10450_ = _10451_ | _10453_ /*7304*/;
assign _10459_ = ~D[30] /*7303*/;
assign _10456_ = _10078_ & _10459_ /*7299*/;
assign _10457_ = _10078_ ^ _10459_ /*7302*/;
assign _10458_ = _10450_ & _10457_ /*7300*/;
assign _10303_ = _10450_ ^ _10457_ /*7301*/;
assign _10455_ = _10456_ | _10458_ /*7298*/;
assign _10460_ = _10079_ & oneWire /*7293*/;
assign _10461_ = _10079_ ^ oneWire /*7296*/;
assign _10462_ = _10455_ & _10461_ /*7294*/;
assign _10304_ = _10455_ ^ _10461_ /*7295*/;
assign Q[8] = _10460_ | _10462_ /*7292*/;
assign _10531_ = ~Q[8] /*7099*/;
assign _10530_ = _10531_ & D[0] /*7098*/;
assign _10533_ = _10273_ & _10530_ /*7093*/;
assign _10534_ = _10273_ ^ _10530_ /*7096*/;
assign _10535_ = zeroWire & _10534_ /*7094*/;
assign _10497_ = zeroWire ^ _10534_ /*7095*/;
assign _10532_ = _10533_ | _10535_ /*7092*/;
assign _10537_ = ~Q[8] /*7091*/;
assign _10536_ = _10537_ & D[1] /*7090*/;
assign _10539_ = _10274_ & _10536_ /*7085*/;
assign _10540_ = _10274_ ^ _10536_ /*7088*/;
assign _10541_ = _10532_ & _10540_ /*7086*/;
assign _10498_ = _10532_ ^ _10540_ /*7087*/;
assign _10538_ = _10539_ | _10541_ /*7084*/;
assign _10543_ = ~Q[8] /*7083*/;
assign _10542_ = _10543_ & D[2] /*7082*/;
assign _10545_ = _10275_ & _10542_ /*7077*/;
assign _10546_ = _10275_ ^ _10542_ /*7080*/;
assign _10547_ = _10538_ & _10546_ /*7078*/;
assign _10499_ = _10538_ ^ _10546_ /*7079*/;
assign _10544_ = _10545_ | _10547_ /*7076*/;
assign _10549_ = ~Q[8] /*7075*/;
assign _10548_ = _10549_ & D[3] /*7074*/;
assign _10551_ = _10276_ & _10548_ /*7069*/;
assign _10552_ = _10276_ ^ _10548_ /*7072*/;
assign _10553_ = _10544_ & _10552_ /*7070*/;
assign _10500_ = _10544_ ^ _10552_ /*7071*/;
assign _10550_ = _10551_ | _10553_ /*7068*/;
assign _10555_ = ~Q[8] /*7067*/;
assign _10554_ = _10555_ & D[4] /*7066*/;
assign _10557_ = _10277_ & _10554_ /*7061*/;
assign _10558_ = _10277_ ^ _10554_ /*7064*/;
assign _10559_ = _10550_ & _10558_ /*7062*/;
assign _10501_ = _10550_ ^ _10558_ /*7063*/;
assign _10556_ = _10557_ | _10559_ /*7060*/;
assign _10561_ = ~Q[8] /*7059*/;
assign _10560_ = _10561_ & D[5] /*7058*/;
assign _10563_ = _10278_ & _10560_ /*7053*/;
assign _10564_ = _10278_ ^ _10560_ /*7056*/;
assign _10565_ = _10556_ & _10564_ /*7054*/;
assign _10502_ = _10556_ ^ _10564_ /*7055*/;
assign _10562_ = _10563_ | _10565_ /*7052*/;
assign _10567_ = ~Q[8] /*7051*/;
assign _10566_ = _10567_ & D[6] /*7050*/;
assign _10569_ = _10279_ & _10566_ /*7045*/;
assign _10570_ = _10279_ ^ _10566_ /*7048*/;
assign _10571_ = _10562_ & _10570_ /*7046*/;
assign _10503_ = _10562_ ^ _10570_ /*7047*/;
assign _10568_ = _10569_ | _10571_ /*7044*/;
assign _10573_ = ~Q[8] /*7043*/;
assign _10572_ = _10573_ & D[7] /*7042*/;
assign _10575_ = _10280_ & _10572_ /*7037*/;
assign _10576_ = _10280_ ^ _10572_ /*7040*/;
assign _10577_ = _10568_ & _10576_ /*7038*/;
assign _10504_ = _10568_ ^ _10576_ /*7039*/;
assign _10574_ = _10575_ | _10577_ /*7036*/;
assign _10579_ = ~Q[8] /*7035*/;
assign _10578_ = _10579_ & D[8] /*7034*/;
assign _10581_ = _10281_ & _10578_ /*7029*/;
assign _10582_ = _10281_ ^ _10578_ /*7032*/;
assign _10583_ = _10574_ & _10582_ /*7030*/;
assign _10505_ = _10574_ ^ _10582_ /*7031*/;
assign _10580_ = _10581_ | _10583_ /*7028*/;
assign _10585_ = ~Q[8] /*7027*/;
assign _10584_ = _10585_ & D[9] /*7026*/;
assign _10587_ = _10282_ & _10584_ /*7021*/;
assign _10588_ = _10282_ ^ _10584_ /*7024*/;
assign _10589_ = _10580_ & _10588_ /*7022*/;
assign _10506_ = _10580_ ^ _10588_ /*7023*/;
assign _10586_ = _10587_ | _10589_ /*7020*/;
assign _10591_ = ~Q[8] /*7019*/;
assign _10590_ = _10591_ & D[10] /*7018*/;
assign _10593_ = _10283_ & _10590_ /*7013*/;
assign _10594_ = _10283_ ^ _10590_ /*7016*/;
assign _10595_ = _10586_ & _10594_ /*7014*/;
assign _10507_ = _10586_ ^ _10594_ /*7015*/;
assign _10592_ = _10593_ | _10595_ /*7012*/;
assign _10597_ = ~Q[8] /*7011*/;
assign _10596_ = _10597_ & D[11] /*7010*/;
assign _10599_ = _10284_ & _10596_ /*7005*/;
assign _10600_ = _10284_ ^ _10596_ /*7008*/;
assign _10601_ = _10592_ & _10600_ /*7006*/;
assign _10508_ = _10592_ ^ _10600_ /*7007*/;
assign _10598_ = _10599_ | _10601_ /*7004*/;
assign _10603_ = ~Q[8] /*7003*/;
assign _10602_ = _10603_ & D[12] /*7002*/;
assign _10605_ = _10285_ & _10602_ /*6997*/;
assign _10606_ = _10285_ ^ _10602_ /*7000*/;
assign _10607_ = _10598_ & _10606_ /*6998*/;
assign _10509_ = _10598_ ^ _10606_ /*6999*/;
assign _10604_ = _10605_ | _10607_ /*6996*/;
assign _10609_ = ~Q[8] /*6995*/;
assign _10608_ = _10609_ & D[13] /*6994*/;
assign _10611_ = _10286_ & _10608_ /*6989*/;
assign _10612_ = _10286_ ^ _10608_ /*6992*/;
assign _10613_ = _10604_ & _10612_ /*6990*/;
assign _10510_ = _10604_ ^ _10612_ /*6991*/;
assign _10610_ = _10611_ | _10613_ /*6988*/;
assign _10615_ = ~Q[8] /*6987*/;
assign _10614_ = _10615_ & D[14] /*6986*/;
assign _10617_ = _10287_ & _10614_ /*6981*/;
assign _10618_ = _10287_ ^ _10614_ /*6984*/;
assign _10619_ = _10610_ & _10618_ /*6982*/;
assign _10511_ = _10610_ ^ _10618_ /*6983*/;
assign _10616_ = _10617_ | _10619_ /*6980*/;
assign _10621_ = ~Q[8] /*6979*/;
assign _10620_ = _10621_ & D[15] /*6978*/;
assign _10623_ = _10288_ & _10620_ /*6973*/;
assign _10624_ = _10288_ ^ _10620_ /*6976*/;
assign _10625_ = _10616_ & _10624_ /*6974*/;
assign _10512_ = _10616_ ^ _10624_ /*6975*/;
assign _10622_ = _10623_ | _10625_ /*6972*/;
assign _10627_ = ~Q[8] /*6971*/;
assign _10626_ = _10627_ & D[16] /*6970*/;
assign _10629_ = _10289_ & _10626_ /*6965*/;
assign _10630_ = _10289_ ^ _10626_ /*6968*/;
assign _10631_ = _10622_ & _10630_ /*6966*/;
assign _10513_ = _10622_ ^ _10630_ /*6967*/;
assign _10628_ = _10629_ | _10631_ /*6964*/;
assign _10633_ = ~Q[8] /*6963*/;
assign _10632_ = _10633_ & D[17] /*6962*/;
assign _10635_ = _10290_ & _10632_ /*6957*/;
assign _10636_ = _10290_ ^ _10632_ /*6960*/;
assign _10637_ = _10628_ & _10636_ /*6958*/;
assign _10514_ = _10628_ ^ _10636_ /*6959*/;
assign _10634_ = _10635_ | _10637_ /*6956*/;
assign _10639_ = ~Q[8] /*6955*/;
assign _10638_ = _10639_ & D[18] /*6954*/;
assign _10641_ = _10291_ & _10638_ /*6949*/;
assign _10642_ = _10291_ ^ _10638_ /*6952*/;
assign _10643_ = _10634_ & _10642_ /*6950*/;
assign _10515_ = _10634_ ^ _10642_ /*6951*/;
assign _10640_ = _10641_ | _10643_ /*6948*/;
assign _10645_ = ~Q[8] /*6947*/;
assign _10644_ = _10645_ & D[19] /*6946*/;
assign _10647_ = _10292_ & _10644_ /*6941*/;
assign _10648_ = _10292_ ^ _10644_ /*6944*/;
assign _10649_ = _10640_ & _10648_ /*6942*/;
assign _10516_ = _10640_ ^ _10648_ /*6943*/;
assign _10646_ = _10647_ | _10649_ /*6940*/;
assign _10651_ = ~Q[8] /*6939*/;
assign _10650_ = _10651_ & D[20] /*6938*/;
assign _10653_ = _10293_ & _10650_ /*6933*/;
assign _10654_ = _10293_ ^ _10650_ /*6936*/;
assign _10655_ = _10646_ & _10654_ /*6934*/;
assign _10517_ = _10646_ ^ _10654_ /*6935*/;
assign _10652_ = _10653_ | _10655_ /*6932*/;
assign _10657_ = ~Q[8] /*6931*/;
assign _10656_ = _10657_ & D[21] /*6930*/;
assign _10659_ = _10294_ & _10656_ /*6925*/;
assign _10660_ = _10294_ ^ _10656_ /*6928*/;
assign _10661_ = _10652_ & _10660_ /*6926*/;
assign _10518_ = _10652_ ^ _10660_ /*6927*/;
assign _10658_ = _10659_ | _10661_ /*6924*/;
assign _10663_ = ~Q[8] /*6923*/;
assign _10662_ = _10663_ & D[22] /*6922*/;
assign _10665_ = _10295_ & _10662_ /*6917*/;
assign _10666_ = _10295_ ^ _10662_ /*6920*/;
assign _10667_ = _10658_ & _10666_ /*6918*/;
assign _10519_ = _10658_ ^ _10666_ /*6919*/;
assign _10664_ = _10665_ | _10667_ /*6916*/;
assign _10669_ = ~Q[8] /*6915*/;
assign _10668_ = _10669_ & D[23] /*6914*/;
assign _10671_ = _10296_ & _10668_ /*6909*/;
assign _10672_ = _10296_ ^ _10668_ /*6912*/;
assign _10673_ = _10664_ & _10672_ /*6910*/;
assign _10520_ = _10664_ ^ _10672_ /*6911*/;
assign _10670_ = _10671_ | _10673_ /*6908*/;
assign _10675_ = ~Q[8] /*6907*/;
assign _10674_ = _10675_ & D[24] /*6906*/;
assign _10677_ = _10297_ & _10674_ /*6901*/;
assign _10678_ = _10297_ ^ _10674_ /*6904*/;
assign _10679_ = _10670_ & _10678_ /*6902*/;
assign _10521_ = _10670_ ^ _10678_ /*6903*/;
assign _10676_ = _10677_ | _10679_ /*6900*/;
assign _10681_ = ~Q[8] /*6899*/;
assign _10680_ = _10681_ & D[25] /*6898*/;
assign _10683_ = _10298_ & _10680_ /*6893*/;
assign _10684_ = _10298_ ^ _10680_ /*6896*/;
assign _10685_ = _10676_ & _10684_ /*6894*/;
assign _10522_ = _10676_ ^ _10684_ /*6895*/;
assign _10682_ = _10683_ | _10685_ /*6892*/;
assign _10687_ = ~Q[8] /*6891*/;
assign _10686_ = _10687_ & D[26] /*6890*/;
assign _10689_ = _10299_ & _10686_ /*6885*/;
assign _10690_ = _10299_ ^ _10686_ /*6888*/;
assign _10691_ = _10682_ & _10690_ /*6886*/;
assign _10523_ = _10682_ ^ _10690_ /*6887*/;
assign _10688_ = _10689_ | _10691_ /*6884*/;
assign _10693_ = ~Q[8] /*6883*/;
assign _10692_ = _10693_ & D[27] /*6882*/;
assign _10695_ = _10300_ & _10692_ /*6877*/;
assign _10696_ = _10300_ ^ _10692_ /*6880*/;
assign _10697_ = _10688_ & _10696_ /*6878*/;
assign _10524_ = _10688_ ^ _10696_ /*6879*/;
assign _10694_ = _10695_ | _10697_ /*6876*/;
assign _10699_ = ~Q[8] /*6875*/;
assign _10698_ = _10699_ & D[28] /*6874*/;
assign _10701_ = _10301_ & _10698_ /*6869*/;
assign _10702_ = _10301_ ^ _10698_ /*6872*/;
assign _10703_ = _10694_ & _10702_ /*6870*/;
assign _10525_ = _10694_ ^ _10702_ /*6871*/;
assign _10700_ = _10701_ | _10703_ /*6868*/;
assign _10705_ = ~Q[8] /*6867*/;
assign _10704_ = _10705_ & D[29] /*6866*/;
assign _10707_ = _10302_ & _10704_ /*6861*/;
assign _10708_ = _10302_ ^ _10704_ /*6864*/;
assign _10709_ = _10700_ & _10708_ /*6862*/;
assign _10526_ = _10700_ ^ _10708_ /*6863*/;
assign _10706_ = _10707_ | _10709_ /*6860*/;
assign _10711_ = ~Q[8] /*6859*/;
assign _10710_ = _10711_ & D[30] /*6858*/;
assign _10713_ = _10303_ & _10710_ /*6853*/;
assign _10714_ = _10303_ ^ _10710_ /*6856*/;
assign _10715_ = _10706_ & _10714_ /*6854*/;
assign _10527_ = _10706_ ^ _10714_ /*6855*/;
assign _10712_ = _10713_ | _10715_ /*6852*/;
assign _10717_ = ~Q[8] /*6851*/;
assign _10716_ = _10717_ & zeroWire /*6850*/;
assign _10718_ = _10304_ ^ _10716_ /*6848*/;
assign _10528_ = _10718_ ^ _10712_ /*6847*/;
assign _10757_ = ~D[0] /*6721*/;
assign _10754_ = R_0[7] & _10757_ /*6717*/;
assign _10755_ = R_0[7] ^ _10757_ /*6720*/;
assign _10756_ = oneWire & _10755_ /*6718*/;
assign _10721_ = oneWire ^ _10755_ /*6719*/;
assign _10753_ = _10754_ | _10756_ /*6716*/;
assign _10762_ = ~D[1] /*6715*/;
assign _10759_ = _10497_ & _10762_ /*6711*/;
assign _10760_ = _10497_ ^ _10762_ /*6714*/;
assign _10761_ = _10753_ & _10760_ /*6712*/;
assign _10722_ = _10753_ ^ _10760_ /*6713*/;
assign _10758_ = _10759_ | _10761_ /*6710*/;
assign _10767_ = ~D[2] /*6709*/;
assign _10764_ = _10498_ & _10767_ /*6705*/;
assign _10765_ = _10498_ ^ _10767_ /*6708*/;
assign _10766_ = _10758_ & _10765_ /*6706*/;
assign _10723_ = _10758_ ^ _10765_ /*6707*/;
assign _10763_ = _10764_ | _10766_ /*6704*/;
assign _10772_ = ~D[3] /*6703*/;
assign _10769_ = _10499_ & _10772_ /*6699*/;
assign _10770_ = _10499_ ^ _10772_ /*6702*/;
assign _10771_ = _10763_ & _10770_ /*6700*/;
assign _10724_ = _10763_ ^ _10770_ /*6701*/;
assign _10768_ = _10769_ | _10771_ /*6698*/;
assign _10777_ = ~D[4] /*6697*/;
assign _10774_ = _10500_ & _10777_ /*6693*/;
assign _10775_ = _10500_ ^ _10777_ /*6696*/;
assign _10776_ = _10768_ & _10775_ /*6694*/;
assign _10725_ = _10768_ ^ _10775_ /*6695*/;
assign _10773_ = _10774_ | _10776_ /*6692*/;
assign _10782_ = ~D[5] /*6691*/;
assign _10779_ = _10501_ & _10782_ /*6687*/;
assign _10780_ = _10501_ ^ _10782_ /*6690*/;
assign _10781_ = _10773_ & _10780_ /*6688*/;
assign _10726_ = _10773_ ^ _10780_ /*6689*/;
assign _10778_ = _10779_ | _10781_ /*6686*/;
assign _10787_ = ~D[6] /*6685*/;
assign _10784_ = _10502_ & _10787_ /*6681*/;
assign _10785_ = _10502_ ^ _10787_ /*6684*/;
assign _10786_ = _10778_ & _10785_ /*6682*/;
assign _10727_ = _10778_ ^ _10785_ /*6683*/;
assign _10783_ = _10784_ | _10786_ /*6680*/;
assign _10792_ = ~D[7] /*6679*/;
assign _10789_ = _10503_ & _10792_ /*6675*/;
assign _10790_ = _10503_ ^ _10792_ /*6678*/;
assign _10791_ = _10783_ & _10790_ /*6676*/;
assign _10728_ = _10783_ ^ _10790_ /*6677*/;
assign _10788_ = _10789_ | _10791_ /*6674*/;
assign _10797_ = ~D[8] /*6673*/;
assign _10794_ = _10504_ & _10797_ /*6669*/;
assign _10795_ = _10504_ ^ _10797_ /*6672*/;
assign _10796_ = _10788_ & _10795_ /*6670*/;
assign _10729_ = _10788_ ^ _10795_ /*6671*/;
assign _10793_ = _10794_ | _10796_ /*6668*/;
assign _10802_ = ~D[9] /*6667*/;
assign _10799_ = _10505_ & _10802_ /*6663*/;
assign _10800_ = _10505_ ^ _10802_ /*6666*/;
assign _10801_ = _10793_ & _10800_ /*6664*/;
assign _10730_ = _10793_ ^ _10800_ /*6665*/;
assign _10798_ = _10799_ | _10801_ /*6662*/;
assign _10807_ = ~D[10] /*6661*/;
assign _10804_ = _10506_ & _10807_ /*6657*/;
assign _10805_ = _10506_ ^ _10807_ /*6660*/;
assign _10806_ = _10798_ & _10805_ /*6658*/;
assign _10731_ = _10798_ ^ _10805_ /*6659*/;
assign _10803_ = _10804_ | _10806_ /*6656*/;
assign _10812_ = ~D[11] /*6655*/;
assign _10809_ = _10507_ & _10812_ /*6651*/;
assign _10810_ = _10507_ ^ _10812_ /*6654*/;
assign _10811_ = _10803_ & _10810_ /*6652*/;
assign _10732_ = _10803_ ^ _10810_ /*6653*/;
assign _10808_ = _10809_ | _10811_ /*6650*/;
assign _10817_ = ~D[12] /*6649*/;
assign _10814_ = _10508_ & _10817_ /*6645*/;
assign _10815_ = _10508_ ^ _10817_ /*6648*/;
assign _10816_ = _10808_ & _10815_ /*6646*/;
assign _10733_ = _10808_ ^ _10815_ /*6647*/;
assign _10813_ = _10814_ | _10816_ /*6644*/;
assign _10822_ = ~D[13] /*6643*/;
assign _10819_ = _10509_ & _10822_ /*6639*/;
assign _10820_ = _10509_ ^ _10822_ /*6642*/;
assign _10821_ = _10813_ & _10820_ /*6640*/;
assign _10734_ = _10813_ ^ _10820_ /*6641*/;
assign _10818_ = _10819_ | _10821_ /*6638*/;
assign _10827_ = ~D[14] /*6637*/;
assign _10824_ = _10510_ & _10827_ /*6633*/;
assign _10825_ = _10510_ ^ _10827_ /*6636*/;
assign _10826_ = _10818_ & _10825_ /*6634*/;
assign _10735_ = _10818_ ^ _10825_ /*6635*/;
assign _10823_ = _10824_ | _10826_ /*6632*/;
assign _10832_ = ~D[15] /*6631*/;
assign _10829_ = _10511_ & _10832_ /*6627*/;
assign _10830_ = _10511_ ^ _10832_ /*6630*/;
assign _10831_ = _10823_ & _10830_ /*6628*/;
assign _10736_ = _10823_ ^ _10830_ /*6629*/;
assign _10828_ = _10829_ | _10831_ /*6626*/;
assign _10837_ = ~D[16] /*6625*/;
assign _10834_ = _10512_ & _10837_ /*6621*/;
assign _10835_ = _10512_ ^ _10837_ /*6624*/;
assign _10836_ = _10828_ & _10835_ /*6622*/;
assign _10737_ = _10828_ ^ _10835_ /*6623*/;
assign _10833_ = _10834_ | _10836_ /*6620*/;
assign _10842_ = ~D[17] /*6619*/;
assign _10839_ = _10513_ & _10842_ /*6615*/;
assign _10840_ = _10513_ ^ _10842_ /*6618*/;
assign _10841_ = _10833_ & _10840_ /*6616*/;
assign _10738_ = _10833_ ^ _10840_ /*6617*/;
assign _10838_ = _10839_ | _10841_ /*6614*/;
assign _10847_ = ~D[18] /*6613*/;
assign _10844_ = _10514_ & _10847_ /*6609*/;
assign _10845_ = _10514_ ^ _10847_ /*6612*/;
assign _10846_ = _10838_ & _10845_ /*6610*/;
assign _10739_ = _10838_ ^ _10845_ /*6611*/;
assign _10843_ = _10844_ | _10846_ /*6608*/;
assign _10852_ = ~D[19] /*6607*/;
assign _10849_ = _10515_ & _10852_ /*6603*/;
assign _10850_ = _10515_ ^ _10852_ /*6606*/;
assign _10851_ = _10843_ & _10850_ /*6604*/;
assign _10740_ = _10843_ ^ _10850_ /*6605*/;
assign _10848_ = _10849_ | _10851_ /*6602*/;
assign _10857_ = ~D[20] /*6601*/;
assign _10854_ = _10516_ & _10857_ /*6597*/;
assign _10855_ = _10516_ ^ _10857_ /*6600*/;
assign _10856_ = _10848_ & _10855_ /*6598*/;
assign _10741_ = _10848_ ^ _10855_ /*6599*/;
assign _10853_ = _10854_ | _10856_ /*6596*/;
assign _10862_ = ~D[21] /*6595*/;
assign _10859_ = _10517_ & _10862_ /*6591*/;
assign _10860_ = _10517_ ^ _10862_ /*6594*/;
assign _10861_ = _10853_ & _10860_ /*6592*/;
assign _10742_ = _10853_ ^ _10860_ /*6593*/;
assign _10858_ = _10859_ | _10861_ /*6590*/;
assign _10867_ = ~D[22] /*6589*/;
assign _10864_ = _10518_ & _10867_ /*6585*/;
assign _10865_ = _10518_ ^ _10867_ /*6588*/;
assign _10866_ = _10858_ & _10865_ /*6586*/;
assign _10743_ = _10858_ ^ _10865_ /*6587*/;
assign _10863_ = _10864_ | _10866_ /*6584*/;
assign _10872_ = ~D[23] /*6583*/;
assign _10869_ = _10519_ & _10872_ /*6579*/;
assign _10870_ = _10519_ ^ _10872_ /*6582*/;
assign _10871_ = _10863_ & _10870_ /*6580*/;
assign _10744_ = _10863_ ^ _10870_ /*6581*/;
assign _10868_ = _10869_ | _10871_ /*6578*/;
assign _10877_ = ~D[24] /*6577*/;
assign _10874_ = _10520_ & _10877_ /*6573*/;
assign _10875_ = _10520_ ^ _10877_ /*6576*/;
assign _10876_ = _10868_ & _10875_ /*6574*/;
assign _10745_ = _10868_ ^ _10875_ /*6575*/;
assign _10873_ = _10874_ | _10876_ /*6572*/;
assign _10882_ = ~D[25] /*6571*/;
assign _10879_ = _10521_ & _10882_ /*6567*/;
assign _10880_ = _10521_ ^ _10882_ /*6570*/;
assign _10881_ = _10873_ & _10880_ /*6568*/;
assign _10746_ = _10873_ ^ _10880_ /*6569*/;
assign _10878_ = _10879_ | _10881_ /*6566*/;
assign _10887_ = ~D[26] /*6565*/;
assign _10884_ = _10522_ & _10887_ /*6561*/;
assign _10885_ = _10522_ ^ _10887_ /*6564*/;
assign _10886_ = _10878_ & _10885_ /*6562*/;
assign _10747_ = _10878_ ^ _10885_ /*6563*/;
assign _10883_ = _10884_ | _10886_ /*6560*/;
assign _10892_ = ~D[27] /*6559*/;
assign _10889_ = _10523_ & _10892_ /*6555*/;
assign _10890_ = _10523_ ^ _10892_ /*6558*/;
assign _10891_ = _10883_ & _10890_ /*6556*/;
assign _10748_ = _10883_ ^ _10890_ /*6557*/;
assign _10888_ = _10889_ | _10891_ /*6554*/;
assign _10897_ = ~D[28] /*6553*/;
assign _10894_ = _10524_ & _10897_ /*6549*/;
assign _10895_ = _10524_ ^ _10897_ /*6552*/;
assign _10896_ = _10888_ & _10895_ /*6550*/;
assign _10749_ = _10888_ ^ _10895_ /*6551*/;
assign _10893_ = _10894_ | _10896_ /*6548*/;
assign _10902_ = ~D[29] /*6547*/;
assign _10899_ = _10525_ & _10902_ /*6543*/;
assign _10900_ = _10525_ ^ _10902_ /*6546*/;
assign _10901_ = _10893_ & _10900_ /*6544*/;
assign _10750_ = _10893_ ^ _10900_ /*6545*/;
assign _10898_ = _10899_ | _10901_ /*6542*/;
assign _10907_ = ~D[30] /*6541*/;
assign _10904_ = _10526_ & _10907_ /*6537*/;
assign _10905_ = _10526_ ^ _10907_ /*6540*/;
assign _10906_ = _10898_ & _10905_ /*6538*/;
assign _10751_ = _10898_ ^ _10905_ /*6539*/;
assign _10903_ = _10904_ | _10906_ /*6536*/;
assign _10908_ = _10527_ & oneWire /*6531*/;
assign _10909_ = _10527_ ^ oneWire /*6534*/;
assign _10910_ = _10903_ & _10909_ /*6532*/;
assign _10752_ = _10903_ ^ _10909_ /*6533*/;
assign Q[7] = _10908_ | _10910_ /*6530*/;
assign _10979_ = ~Q[7] /*6337*/;
assign _10978_ = _10979_ & D[0] /*6336*/;
assign _10981_ = _10721_ & _10978_ /*6331*/;
assign _10982_ = _10721_ ^ _10978_ /*6334*/;
assign _10983_ = zeroWire & _10982_ /*6332*/;
assign _10945_ = zeroWire ^ _10982_ /*6333*/;
assign _10980_ = _10981_ | _10983_ /*6330*/;
assign _10985_ = ~Q[7] /*6329*/;
assign _10984_ = _10985_ & D[1] /*6328*/;
assign _10987_ = _10722_ & _10984_ /*6323*/;
assign _10988_ = _10722_ ^ _10984_ /*6326*/;
assign _10989_ = _10980_ & _10988_ /*6324*/;
assign _10946_ = _10980_ ^ _10988_ /*6325*/;
assign _10986_ = _10987_ | _10989_ /*6322*/;
assign _10991_ = ~Q[7] /*6321*/;
assign _10990_ = _10991_ & D[2] /*6320*/;
assign _10993_ = _10723_ & _10990_ /*6315*/;
assign _10994_ = _10723_ ^ _10990_ /*6318*/;
assign _10995_ = _10986_ & _10994_ /*6316*/;
assign _10947_ = _10986_ ^ _10994_ /*6317*/;
assign _10992_ = _10993_ | _10995_ /*6314*/;
assign _10997_ = ~Q[7] /*6313*/;
assign _10996_ = _10997_ & D[3] /*6312*/;
assign _10999_ = _10724_ & _10996_ /*6307*/;
assign _11000_ = _10724_ ^ _10996_ /*6310*/;
assign _11001_ = _10992_ & _11000_ /*6308*/;
assign _10948_ = _10992_ ^ _11000_ /*6309*/;
assign _10998_ = _10999_ | _11001_ /*6306*/;
assign _11003_ = ~Q[7] /*6305*/;
assign _11002_ = _11003_ & D[4] /*6304*/;
assign _11005_ = _10725_ & _11002_ /*6299*/;
assign _11006_ = _10725_ ^ _11002_ /*6302*/;
assign _11007_ = _10998_ & _11006_ /*6300*/;
assign _10949_ = _10998_ ^ _11006_ /*6301*/;
assign _11004_ = _11005_ | _11007_ /*6298*/;
assign _11009_ = ~Q[7] /*6297*/;
assign _11008_ = _11009_ & D[5] /*6296*/;
assign _11011_ = _10726_ & _11008_ /*6291*/;
assign _11012_ = _10726_ ^ _11008_ /*6294*/;
assign _11013_ = _11004_ & _11012_ /*6292*/;
assign _10950_ = _11004_ ^ _11012_ /*6293*/;
assign _11010_ = _11011_ | _11013_ /*6290*/;
assign _11015_ = ~Q[7] /*6289*/;
assign _11014_ = _11015_ & D[6] /*6288*/;
assign _11017_ = _10727_ & _11014_ /*6283*/;
assign _11018_ = _10727_ ^ _11014_ /*6286*/;
assign _11019_ = _11010_ & _11018_ /*6284*/;
assign _10951_ = _11010_ ^ _11018_ /*6285*/;
assign _11016_ = _11017_ | _11019_ /*6282*/;
assign _11021_ = ~Q[7] /*6281*/;
assign _11020_ = _11021_ & D[7] /*6280*/;
assign _11023_ = _10728_ & _11020_ /*6275*/;
assign _11024_ = _10728_ ^ _11020_ /*6278*/;
assign _11025_ = _11016_ & _11024_ /*6276*/;
assign _10952_ = _11016_ ^ _11024_ /*6277*/;
assign _11022_ = _11023_ | _11025_ /*6274*/;
assign _11027_ = ~Q[7] /*6273*/;
assign _11026_ = _11027_ & D[8] /*6272*/;
assign _11029_ = _10729_ & _11026_ /*6267*/;
assign _11030_ = _10729_ ^ _11026_ /*6270*/;
assign _11031_ = _11022_ & _11030_ /*6268*/;
assign _10953_ = _11022_ ^ _11030_ /*6269*/;
assign _11028_ = _11029_ | _11031_ /*6266*/;
assign _11033_ = ~Q[7] /*6265*/;
assign _11032_ = _11033_ & D[9] /*6264*/;
assign _11035_ = _10730_ & _11032_ /*6259*/;
assign _11036_ = _10730_ ^ _11032_ /*6262*/;
assign _11037_ = _11028_ & _11036_ /*6260*/;
assign _10954_ = _11028_ ^ _11036_ /*6261*/;
assign _11034_ = _11035_ | _11037_ /*6258*/;
assign _11039_ = ~Q[7] /*6257*/;
assign _11038_ = _11039_ & D[10] /*6256*/;
assign _11041_ = _10731_ & _11038_ /*6251*/;
assign _11042_ = _10731_ ^ _11038_ /*6254*/;
assign _11043_ = _11034_ & _11042_ /*6252*/;
assign _10955_ = _11034_ ^ _11042_ /*6253*/;
assign _11040_ = _11041_ | _11043_ /*6250*/;
assign _11045_ = ~Q[7] /*6249*/;
assign _11044_ = _11045_ & D[11] /*6248*/;
assign _11047_ = _10732_ & _11044_ /*6243*/;
assign _11048_ = _10732_ ^ _11044_ /*6246*/;
assign _11049_ = _11040_ & _11048_ /*6244*/;
assign _10956_ = _11040_ ^ _11048_ /*6245*/;
assign _11046_ = _11047_ | _11049_ /*6242*/;
assign _11051_ = ~Q[7] /*6241*/;
assign _11050_ = _11051_ & D[12] /*6240*/;
assign _11053_ = _10733_ & _11050_ /*6235*/;
assign _11054_ = _10733_ ^ _11050_ /*6238*/;
assign _11055_ = _11046_ & _11054_ /*6236*/;
assign _10957_ = _11046_ ^ _11054_ /*6237*/;
assign _11052_ = _11053_ | _11055_ /*6234*/;
assign _11057_ = ~Q[7] /*6233*/;
assign _11056_ = _11057_ & D[13] /*6232*/;
assign _11059_ = _10734_ & _11056_ /*6227*/;
assign _11060_ = _10734_ ^ _11056_ /*6230*/;
assign _11061_ = _11052_ & _11060_ /*6228*/;
assign _10958_ = _11052_ ^ _11060_ /*6229*/;
assign _11058_ = _11059_ | _11061_ /*6226*/;
assign _11063_ = ~Q[7] /*6225*/;
assign _11062_ = _11063_ & D[14] /*6224*/;
assign _11065_ = _10735_ & _11062_ /*6219*/;
assign _11066_ = _10735_ ^ _11062_ /*6222*/;
assign _11067_ = _11058_ & _11066_ /*6220*/;
assign _10959_ = _11058_ ^ _11066_ /*6221*/;
assign _11064_ = _11065_ | _11067_ /*6218*/;
assign _11069_ = ~Q[7] /*6217*/;
assign _11068_ = _11069_ & D[15] /*6216*/;
assign _11071_ = _10736_ & _11068_ /*6211*/;
assign _11072_ = _10736_ ^ _11068_ /*6214*/;
assign _11073_ = _11064_ & _11072_ /*6212*/;
assign _10960_ = _11064_ ^ _11072_ /*6213*/;
assign _11070_ = _11071_ | _11073_ /*6210*/;
assign _11075_ = ~Q[7] /*6209*/;
assign _11074_ = _11075_ & D[16] /*6208*/;
assign _11077_ = _10737_ & _11074_ /*6203*/;
assign _11078_ = _10737_ ^ _11074_ /*6206*/;
assign _11079_ = _11070_ & _11078_ /*6204*/;
assign _10961_ = _11070_ ^ _11078_ /*6205*/;
assign _11076_ = _11077_ | _11079_ /*6202*/;
assign _11081_ = ~Q[7] /*6201*/;
assign _11080_ = _11081_ & D[17] /*6200*/;
assign _11083_ = _10738_ & _11080_ /*6195*/;
assign _11084_ = _10738_ ^ _11080_ /*6198*/;
assign _11085_ = _11076_ & _11084_ /*6196*/;
assign _10962_ = _11076_ ^ _11084_ /*6197*/;
assign _11082_ = _11083_ | _11085_ /*6194*/;
assign _11087_ = ~Q[7] /*6193*/;
assign _11086_ = _11087_ & D[18] /*6192*/;
assign _11089_ = _10739_ & _11086_ /*6187*/;
assign _11090_ = _10739_ ^ _11086_ /*6190*/;
assign _11091_ = _11082_ & _11090_ /*6188*/;
assign _10963_ = _11082_ ^ _11090_ /*6189*/;
assign _11088_ = _11089_ | _11091_ /*6186*/;
assign _11093_ = ~Q[7] /*6185*/;
assign _11092_ = _11093_ & D[19] /*6184*/;
assign _11095_ = _10740_ & _11092_ /*6179*/;
assign _11096_ = _10740_ ^ _11092_ /*6182*/;
assign _11097_ = _11088_ & _11096_ /*6180*/;
assign _10964_ = _11088_ ^ _11096_ /*6181*/;
assign _11094_ = _11095_ | _11097_ /*6178*/;
assign _11099_ = ~Q[7] /*6177*/;
assign _11098_ = _11099_ & D[20] /*6176*/;
assign _11101_ = _10741_ & _11098_ /*6171*/;
assign _11102_ = _10741_ ^ _11098_ /*6174*/;
assign _11103_ = _11094_ & _11102_ /*6172*/;
assign _10965_ = _11094_ ^ _11102_ /*6173*/;
assign _11100_ = _11101_ | _11103_ /*6170*/;
assign _11105_ = ~Q[7] /*6169*/;
assign _11104_ = _11105_ & D[21] /*6168*/;
assign _11107_ = _10742_ & _11104_ /*6163*/;
assign _11108_ = _10742_ ^ _11104_ /*6166*/;
assign _11109_ = _11100_ & _11108_ /*6164*/;
assign _10966_ = _11100_ ^ _11108_ /*6165*/;
assign _11106_ = _11107_ | _11109_ /*6162*/;
assign _11111_ = ~Q[7] /*6161*/;
assign _11110_ = _11111_ & D[22] /*6160*/;
assign _11113_ = _10743_ & _11110_ /*6155*/;
assign _11114_ = _10743_ ^ _11110_ /*6158*/;
assign _11115_ = _11106_ & _11114_ /*6156*/;
assign _10967_ = _11106_ ^ _11114_ /*6157*/;
assign _11112_ = _11113_ | _11115_ /*6154*/;
assign _11117_ = ~Q[7] /*6153*/;
assign _11116_ = _11117_ & D[23] /*6152*/;
assign _11119_ = _10744_ & _11116_ /*6147*/;
assign _11120_ = _10744_ ^ _11116_ /*6150*/;
assign _11121_ = _11112_ & _11120_ /*6148*/;
assign _10968_ = _11112_ ^ _11120_ /*6149*/;
assign _11118_ = _11119_ | _11121_ /*6146*/;
assign _11123_ = ~Q[7] /*6145*/;
assign _11122_ = _11123_ & D[24] /*6144*/;
assign _11125_ = _10745_ & _11122_ /*6139*/;
assign _11126_ = _10745_ ^ _11122_ /*6142*/;
assign _11127_ = _11118_ & _11126_ /*6140*/;
assign _10969_ = _11118_ ^ _11126_ /*6141*/;
assign _11124_ = _11125_ | _11127_ /*6138*/;
assign _11129_ = ~Q[7] /*6137*/;
assign _11128_ = _11129_ & D[25] /*6136*/;
assign _11131_ = _10746_ & _11128_ /*6131*/;
assign _11132_ = _10746_ ^ _11128_ /*6134*/;
assign _11133_ = _11124_ & _11132_ /*6132*/;
assign _10970_ = _11124_ ^ _11132_ /*6133*/;
assign _11130_ = _11131_ | _11133_ /*6130*/;
assign _11135_ = ~Q[7] /*6129*/;
assign _11134_ = _11135_ & D[26] /*6128*/;
assign _11137_ = _10747_ & _11134_ /*6123*/;
assign _11138_ = _10747_ ^ _11134_ /*6126*/;
assign _11139_ = _11130_ & _11138_ /*6124*/;
assign _10971_ = _11130_ ^ _11138_ /*6125*/;
assign _11136_ = _11137_ | _11139_ /*6122*/;
assign _11141_ = ~Q[7] /*6121*/;
assign _11140_ = _11141_ & D[27] /*6120*/;
assign _11143_ = _10748_ & _11140_ /*6115*/;
assign _11144_ = _10748_ ^ _11140_ /*6118*/;
assign _11145_ = _11136_ & _11144_ /*6116*/;
assign _10972_ = _11136_ ^ _11144_ /*6117*/;
assign _11142_ = _11143_ | _11145_ /*6114*/;
assign _11147_ = ~Q[7] /*6113*/;
assign _11146_ = _11147_ & D[28] /*6112*/;
assign _11149_ = _10749_ & _11146_ /*6107*/;
assign _11150_ = _10749_ ^ _11146_ /*6110*/;
assign _11151_ = _11142_ & _11150_ /*6108*/;
assign _10973_ = _11142_ ^ _11150_ /*6109*/;
assign _11148_ = _11149_ | _11151_ /*6106*/;
assign _11153_ = ~Q[7] /*6105*/;
assign _11152_ = _11153_ & D[29] /*6104*/;
assign _11155_ = _10750_ & _11152_ /*6099*/;
assign _11156_ = _10750_ ^ _11152_ /*6102*/;
assign _11157_ = _11148_ & _11156_ /*6100*/;
assign _10974_ = _11148_ ^ _11156_ /*6101*/;
assign _11154_ = _11155_ | _11157_ /*6098*/;
assign _11159_ = ~Q[7] /*6097*/;
assign _11158_ = _11159_ & D[30] /*6096*/;
assign _11161_ = _10751_ & _11158_ /*6091*/;
assign _11162_ = _10751_ ^ _11158_ /*6094*/;
assign _11163_ = _11154_ & _11162_ /*6092*/;
assign _10975_ = _11154_ ^ _11162_ /*6093*/;
assign _11160_ = _11161_ | _11163_ /*6090*/;
assign _11165_ = ~Q[7] /*6089*/;
assign _11164_ = _11165_ & zeroWire /*6088*/;
assign _11166_ = _10752_ ^ _11164_ /*6086*/;
assign _10976_ = _11166_ ^ _11160_ /*6085*/;
assign _11205_ = ~D[0] /*5959*/;
assign _11202_ = R_0[6] & _11205_ /*5955*/;
assign _11203_ = R_0[6] ^ _11205_ /*5958*/;
assign _11204_ = oneWire & _11203_ /*5956*/;
assign _11169_ = oneWire ^ _11203_ /*5957*/;
assign _11201_ = _11202_ | _11204_ /*5954*/;
assign _11210_ = ~D[1] /*5953*/;
assign _11207_ = _10945_ & _11210_ /*5949*/;
assign _11208_ = _10945_ ^ _11210_ /*5952*/;
assign _11209_ = _11201_ & _11208_ /*5950*/;
assign _11170_ = _11201_ ^ _11208_ /*5951*/;
assign _11206_ = _11207_ | _11209_ /*5948*/;
assign _11215_ = ~D[2] /*5947*/;
assign _11212_ = _10946_ & _11215_ /*5943*/;
assign _11213_ = _10946_ ^ _11215_ /*5946*/;
assign _11214_ = _11206_ & _11213_ /*5944*/;
assign _11171_ = _11206_ ^ _11213_ /*5945*/;
assign _11211_ = _11212_ | _11214_ /*5942*/;
assign _11220_ = ~D[3] /*5941*/;
assign _11217_ = _10947_ & _11220_ /*5937*/;
assign _11218_ = _10947_ ^ _11220_ /*5940*/;
assign _11219_ = _11211_ & _11218_ /*5938*/;
assign _11172_ = _11211_ ^ _11218_ /*5939*/;
assign _11216_ = _11217_ | _11219_ /*5936*/;
assign _11225_ = ~D[4] /*5935*/;
assign _11222_ = _10948_ & _11225_ /*5931*/;
assign _11223_ = _10948_ ^ _11225_ /*5934*/;
assign _11224_ = _11216_ & _11223_ /*5932*/;
assign _11173_ = _11216_ ^ _11223_ /*5933*/;
assign _11221_ = _11222_ | _11224_ /*5930*/;
assign _11230_ = ~D[5] /*5929*/;
assign _11227_ = _10949_ & _11230_ /*5925*/;
assign _11228_ = _10949_ ^ _11230_ /*5928*/;
assign _11229_ = _11221_ & _11228_ /*5926*/;
assign _11174_ = _11221_ ^ _11228_ /*5927*/;
assign _11226_ = _11227_ | _11229_ /*5924*/;
assign _11235_ = ~D[6] /*5923*/;
assign _11232_ = _10950_ & _11235_ /*5919*/;
assign _11233_ = _10950_ ^ _11235_ /*5922*/;
assign _11234_ = _11226_ & _11233_ /*5920*/;
assign _11175_ = _11226_ ^ _11233_ /*5921*/;
assign _11231_ = _11232_ | _11234_ /*5918*/;
assign _11240_ = ~D[7] /*5917*/;
assign _11237_ = _10951_ & _11240_ /*5913*/;
assign _11238_ = _10951_ ^ _11240_ /*5916*/;
assign _11239_ = _11231_ & _11238_ /*5914*/;
assign _11176_ = _11231_ ^ _11238_ /*5915*/;
assign _11236_ = _11237_ | _11239_ /*5912*/;
assign _11245_ = ~D[8] /*5911*/;
assign _11242_ = _10952_ & _11245_ /*5907*/;
assign _11243_ = _10952_ ^ _11245_ /*5910*/;
assign _11244_ = _11236_ & _11243_ /*5908*/;
assign _11177_ = _11236_ ^ _11243_ /*5909*/;
assign _11241_ = _11242_ | _11244_ /*5906*/;
assign _11250_ = ~D[9] /*5905*/;
assign _11247_ = _10953_ & _11250_ /*5901*/;
assign _11248_ = _10953_ ^ _11250_ /*5904*/;
assign _11249_ = _11241_ & _11248_ /*5902*/;
assign _11178_ = _11241_ ^ _11248_ /*5903*/;
assign _11246_ = _11247_ | _11249_ /*5900*/;
assign _11255_ = ~D[10] /*5899*/;
assign _11252_ = _10954_ & _11255_ /*5895*/;
assign _11253_ = _10954_ ^ _11255_ /*5898*/;
assign _11254_ = _11246_ & _11253_ /*5896*/;
assign _11179_ = _11246_ ^ _11253_ /*5897*/;
assign _11251_ = _11252_ | _11254_ /*5894*/;
assign _11260_ = ~D[11] /*5893*/;
assign _11257_ = _10955_ & _11260_ /*5889*/;
assign _11258_ = _10955_ ^ _11260_ /*5892*/;
assign _11259_ = _11251_ & _11258_ /*5890*/;
assign _11180_ = _11251_ ^ _11258_ /*5891*/;
assign _11256_ = _11257_ | _11259_ /*5888*/;
assign _11265_ = ~D[12] /*5887*/;
assign _11262_ = _10956_ & _11265_ /*5883*/;
assign _11263_ = _10956_ ^ _11265_ /*5886*/;
assign _11264_ = _11256_ & _11263_ /*5884*/;
assign _11181_ = _11256_ ^ _11263_ /*5885*/;
assign _11261_ = _11262_ | _11264_ /*5882*/;
assign _11270_ = ~D[13] /*5881*/;
assign _11267_ = _10957_ & _11270_ /*5877*/;
assign _11268_ = _10957_ ^ _11270_ /*5880*/;
assign _11269_ = _11261_ & _11268_ /*5878*/;
assign _11182_ = _11261_ ^ _11268_ /*5879*/;
assign _11266_ = _11267_ | _11269_ /*5876*/;
assign _11275_ = ~D[14] /*5875*/;
assign _11272_ = _10958_ & _11275_ /*5871*/;
assign _11273_ = _10958_ ^ _11275_ /*5874*/;
assign _11274_ = _11266_ & _11273_ /*5872*/;
assign _11183_ = _11266_ ^ _11273_ /*5873*/;
assign _11271_ = _11272_ | _11274_ /*5870*/;
assign _11280_ = ~D[15] /*5869*/;
assign _11277_ = _10959_ & _11280_ /*5865*/;
assign _11278_ = _10959_ ^ _11280_ /*5868*/;
assign _11279_ = _11271_ & _11278_ /*5866*/;
assign _11184_ = _11271_ ^ _11278_ /*5867*/;
assign _11276_ = _11277_ | _11279_ /*5864*/;
assign _11285_ = ~D[16] /*5863*/;
assign _11282_ = _10960_ & _11285_ /*5859*/;
assign _11283_ = _10960_ ^ _11285_ /*5862*/;
assign _11284_ = _11276_ & _11283_ /*5860*/;
assign _11185_ = _11276_ ^ _11283_ /*5861*/;
assign _11281_ = _11282_ | _11284_ /*5858*/;
assign _11290_ = ~D[17] /*5857*/;
assign _11287_ = _10961_ & _11290_ /*5853*/;
assign _11288_ = _10961_ ^ _11290_ /*5856*/;
assign _11289_ = _11281_ & _11288_ /*5854*/;
assign _11186_ = _11281_ ^ _11288_ /*5855*/;
assign _11286_ = _11287_ | _11289_ /*5852*/;
assign _11295_ = ~D[18] /*5851*/;
assign _11292_ = _10962_ & _11295_ /*5847*/;
assign _11293_ = _10962_ ^ _11295_ /*5850*/;
assign _11294_ = _11286_ & _11293_ /*5848*/;
assign _11187_ = _11286_ ^ _11293_ /*5849*/;
assign _11291_ = _11292_ | _11294_ /*5846*/;
assign _11300_ = ~D[19] /*5845*/;
assign _11297_ = _10963_ & _11300_ /*5841*/;
assign _11298_ = _10963_ ^ _11300_ /*5844*/;
assign _11299_ = _11291_ & _11298_ /*5842*/;
assign _11188_ = _11291_ ^ _11298_ /*5843*/;
assign _11296_ = _11297_ | _11299_ /*5840*/;
assign _11305_ = ~D[20] /*5839*/;
assign _11302_ = _10964_ & _11305_ /*5835*/;
assign _11303_ = _10964_ ^ _11305_ /*5838*/;
assign _11304_ = _11296_ & _11303_ /*5836*/;
assign _11189_ = _11296_ ^ _11303_ /*5837*/;
assign _11301_ = _11302_ | _11304_ /*5834*/;
assign _11310_ = ~D[21] /*5833*/;
assign _11307_ = _10965_ & _11310_ /*5829*/;
assign _11308_ = _10965_ ^ _11310_ /*5832*/;
assign _11309_ = _11301_ & _11308_ /*5830*/;
assign _11190_ = _11301_ ^ _11308_ /*5831*/;
assign _11306_ = _11307_ | _11309_ /*5828*/;
assign _11315_ = ~D[22] /*5827*/;
assign _11312_ = _10966_ & _11315_ /*5823*/;
assign _11313_ = _10966_ ^ _11315_ /*5826*/;
assign _11314_ = _11306_ & _11313_ /*5824*/;
assign _11191_ = _11306_ ^ _11313_ /*5825*/;
assign _11311_ = _11312_ | _11314_ /*5822*/;
assign _11320_ = ~D[23] /*5821*/;
assign _11317_ = _10967_ & _11320_ /*5817*/;
assign _11318_ = _10967_ ^ _11320_ /*5820*/;
assign _11319_ = _11311_ & _11318_ /*5818*/;
assign _11192_ = _11311_ ^ _11318_ /*5819*/;
assign _11316_ = _11317_ | _11319_ /*5816*/;
assign _11325_ = ~D[24] /*5815*/;
assign _11322_ = _10968_ & _11325_ /*5811*/;
assign _11323_ = _10968_ ^ _11325_ /*5814*/;
assign _11324_ = _11316_ & _11323_ /*5812*/;
assign _11193_ = _11316_ ^ _11323_ /*5813*/;
assign _11321_ = _11322_ | _11324_ /*5810*/;
assign _11330_ = ~D[25] /*5809*/;
assign _11327_ = _10969_ & _11330_ /*5805*/;
assign _11328_ = _10969_ ^ _11330_ /*5808*/;
assign _11329_ = _11321_ & _11328_ /*5806*/;
assign _11194_ = _11321_ ^ _11328_ /*5807*/;
assign _11326_ = _11327_ | _11329_ /*5804*/;
assign _11335_ = ~D[26] /*5803*/;
assign _11332_ = _10970_ & _11335_ /*5799*/;
assign _11333_ = _10970_ ^ _11335_ /*5802*/;
assign _11334_ = _11326_ & _11333_ /*5800*/;
assign _11195_ = _11326_ ^ _11333_ /*5801*/;
assign _11331_ = _11332_ | _11334_ /*5798*/;
assign _11340_ = ~D[27] /*5797*/;
assign _11337_ = _10971_ & _11340_ /*5793*/;
assign _11338_ = _10971_ ^ _11340_ /*5796*/;
assign _11339_ = _11331_ & _11338_ /*5794*/;
assign _11196_ = _11331_ ^ _11338_ /*5795*/;
assign _11336_ = _11337_ | _11339_ /*5792*/;
assign _11345_ = ~D[28] /*5791*/;
assign _11342_ = _10972_ & _11345_ /*5787*/;
assign _11343_ = _10972_ ^ _11345_ /*5790*/;
assign _11344_ = _11336_ & _11343_ /*5788*/;
assign _11197_ = _11336_ ^ _11343_ /*5789*/;
assign _11341_ = _11342_ | _11344_ /*5786*/;
assign _11350_ = ~D[29] /*5785*/;
assign _11347_ = _10973_ & _11350_ /*5781*/;
assign _11348_ = _10973_ ^ _11350_ /*5784*/;
assign _11349_ = _11341_ & _11348_ /*5782*/;
assign _11198_ = _11341_ ^ _11348_ /*5783*/;
assign _11346_ = _11347_ | _11349_ /*5780*/;
assign _11355_ = ~D[30] /*5779*/;
assign _11352_ = _10974_ & _11355_ /*5775*/;
assign _11353_ = _10974_ ^ _11355_ /*5778*/;
assign _11354_ = _11346_ & _11353_ /*5776*/;
assign _11199_ = _11346_ ^ _11353_ /*5777*/;
assign _11351_ = _11352_ | _11354_ /*5774*/;
assign _11356_ = _10975_ & oneWire /*5769*/;
assign _11357_ = _10975_ ^ oneWire /*5772*/;
assign _11358_ = _11351_ & _11357_ /*5770*/;
assign _11200_ = _11351_ ^ _11357_ /*5771*/;
assign Q[6] = _11356_ | _11358_ /*5768*/;
assign _11427_ = ~Q[6] /*5575*/;
assign _11426_ = _11427_ & D[0] /*5574*/;
assign _11429_ = _11169_ & _11426_ /*5569*/;
assign _11430_ = _11169_ ^ _11426_ /*5572*/;
assign _11431_ = zeroWire & _11430_ /*5570*/;
assign _11393_ = zeroWire ^ _11430_ /*5571*/;
assign _11428_ = _11429_ | _11431_ /*5568*/;
assign _11433_ = ~Q[6] /*5567*/;
assign _11432_ = _11433_ & D[1] /*5566*/;
assign _11435_ = _11170_ & _11432_ /*5561*/;
assign _11436_ = _11170_ ^ _11432_ /*5564*/;
assign _11437_ = _11428_ & _11436_ /*5562*/;
assign _11394_ = _11428_ ^ _11436_ /*5563*/;
assign _11434_ = _11435_ | _11437_ /*5560*/;
assign _11439_ = ~Q[6] /*5559*/;
assign _11438_ = _11439_ & D[2] /*5558*/;
assign _11441_ = _11171_ & _11438_ /*5553*/;
assign _11442_ = _11171_ ^ _11438_ /*5556*/;
assign _11443_ = _11434_ & _11442_ /*5554*/;
assign _11395_ = _11434_ ^ _11442_ /*5555*/;
assign _11440_ = _11441_ | _11443_ /*5552*/;
assign _11445_ = ~Q[6] /*5551*/;
assign _11444_ = _11445_ & D[3] /*5550*/;
assign _11447_ = _11172_ & _11444_ /*5545*/;
assign _11448_ = _11172_ ^ _11444_ /*5548*/;
assign _11449_ = _11440_ & _11448_ /*5546*/;
assign _11396_ = _11440_ ^ _11448_ /*5547*/;
assign _11446_ = _11447_ | _11449_ /*5544*/;
assign _11451_ = ~Q[6] /*5543*/;
assign _11450_ = _11451_ & D[4] /*5542*/;
assign _11453_ = _11173_ & _11450_ /*5537*/;
assign _11454_ = _11173_ ^ _11450_ /*5540*/;
assign _11455_ = _11446_ & _11454_ /*5538*/;
assign _11397_ = _11446_ ^ _11454_ /*5539*/;
assign _11452_ = _11453_ | _11455_ /*5536*/;
assign _11457_ = ~Q[6] /*5535*/;
assign _11456_ = _11457_ & D[5] /*5534*/;
assign _11459_ = _11174_ & _11456_ /*5529*/;
assign _11460_ = _11174_ ^ _11456_ /*5532*/;
assign _11461_ = _11452_ & _11460_ /*5530*/;
assign _11398_ = _11452_ ^ _11460_ /*5531*/;
assign _11458_ = _11459_ | _11461_ /*5528*/;
assign _11463_ = ~Q[6] /*5527*/;
assign _11462_ = _11463_ & D[6] /*5526*/;
assign _11465_ = _11175_ & _11462_ /*5521*/;
assign _11466_ = _11175_ ^ _11462_ /*5524*/;
assign _11467_ = _11458_ & _11466_ /*5522*/;
assign _11399_ = _11458_ ^ _11466_ /*5523*/;
assign _11464_ = _11465_ | _11467_ /*5520*/;
assign _11469_ = ~Q[6] /*5519*/;
assign _11468_ = _11469_ & D[7] /*5518*/;
assign _11471_ = _11176_ & _11468_ /*5513*/;
assign _11472_ = _11176_ ^ _11468_ /*5516*/;
assign _11473_ = _11464_ & _11472_ /*5514*/;
assign _11400_ = _11464_ ^ _11472_ /*5515*/;
assign _11470_ = _11471_ | _11473_ /*5512*/;
assign _11475_ = ~Q[6] /*5511*/;
assign _11474_ = _11475_ & D[8] /*5510*/;
assign _11477_ = _11177_ & _11474_ /*5505*/;
assign _11478_ = _11177_ ^ _11474_ /*5508*/;
assign _11479_ = _11470_ & _11478_ /*5506*/;
assign _11401_ = _11470_ ^ _11478_ /*5507*/;
assign _11476_ = _11477_ | _11479_ /*5504*/;
assign _11481_ = ~Q[6] /*5503*/;
assign _11480_ = _11481_ & D[9] /*5502*/;
assign _11483_ = _11178_ & _11480_ /*5497*/;
assign _11484_ = _11178_ ^ _11480_ /*5500*/;
assign _11485_ = _11476_ & _11484_ /*5498*/;
assign _11402_ = _11476_ ^ _11484_ /*5499*/;
assign _11482_ = _11483_ | _11485_ /*5496*/;
assign _11487_ = ~Q[6] /*5495*/;
assign _11486_ = _11487_ & D[10] /*5494*/;
assign _11489_ = _11179_ & _11486_ /*5489*/;
assign _11490_ = _11179_ ^ _11486_ /*5492*/;
assign _11491_ = _11482_ & _11490_ /*5490*/;
assign _11403_ = _11482_ ^ _11490_ /*5491*/;
assign _11488_ = _11489_ | _11491_ /*5488*/;
assign _11493_ = ~Q[6] /*5487*/;
assign _11492_ = _11493_ & D[11] /*5486*/;
assign _11495_ = _11180_ & _11492_ /*5481*/;
assign _11496_ = _11180_ ^ _11492_ /*5484*/;
assign _11497_ = _11488_ & _11496_ /*5482*/;
assign _11404_ = _11488_ ^ _11496_ /*5483*/;
assign _11494_ = _11495_ | _11497_ /*5480*/;
assign _11499_ = ~Q[6] /*5479*/;
assign _11498_ = _11499_ & D[12] /*5478*/;
assign _11501_ = _11181_ & _11498_ /*5473*/;
assign _11502_ = _11181_ ^ _11498_ /*5476*/;
assign _11503_ = _11494_ & _11502_ /*5474*/;
assign _11405_ = _11494_ ^ _11502_ /*5475*/;
assign _11500_ = _11501_ | _11503_ /*5472*/;
assign _11505_ = ~Q[6] /*5471*/;
assign _11504_ = _11505_ & D[13] /*5470*/;
assign _11507_ = _11182_ & _11504_ /*5465*/;
assign _11508_ = _11182_ ^ _11504_ /*5468*/;
assign _11509_ = _11500_ & _11508_ /*5466*/;
assign _11406_ = _11500_ ^ _11508_ /*5467*/;
assign _11506_ = _11507_ | _11509_ /*5464*/;
assign _11511_ = ~Q[6] /*5463*/;
assign _11510_ = _11511_ & D[14] /*5462*/;
assign _11513_ = _11183_ & _11510_ /*5457*/;
assign _11514_ = _11183_ ^ _11510_ /*5460*/;
assign _11515_ = _11506_ & _11514_ /*5458*/;
assign _11407_ = _11506_ ^ _11514_ /*5459*/;
assign _11512_ = _11513_ | _11515_ /*5456*/;
assign _11517_ = ~Q[6] /*5455*/;
assign _11516_ = _11517_ & D[15] /*5454*/;
assign _11519_ = _11184_ & _11516_ /*5449*/;
assign _11520_ = _11184_ ^ _11516_ /*5452*/;
assign _11521_ = _11512_ & _11520_ /*5450*/;
assign _11408_ = _11512_ ^ _11520_ /*5451*/;
assign _11518_ = _11519_ | _11521_ /*5448*/;
assign _11523_ = ~Q[6] /*5447*/;
assign _11522_ = _11523_ & D[16] /*5446*/;
assign _11525_ = _11185_ & _11522_ /*5441*/;
assign _11526_ = _11185_ ^ _11522_ /*5444*/;
assign _11527_ = _11518_ & _11526_ /*5442*/;
assign _11409_ = _11518_ ^ _11526_ /*5443*/;
assign _11524_ = _11525_ | _11527_ /*5440*/;
assign _11529_ = ~Q[6] /*5439*/;
assign _11528_ = _11529_ & D[17] /*5438*/;
assign _11531_ = _11186_ & _11528_ /*5433*/;
assign _11532_ = _11186_ ^ _11528_ /*5436*/;
assign _11533_ = _11524_ & _11532_ /*5434*/;
assign _11410_ = _11524_ ^ _11532_ /*5435*/;
assign _11530_ = _11531_ | _11533_ /*5432*/;
assign _11535_ = ~Q[6] /*5431*/;
assign _11534_ = _11535_ & D[18] /*5430*/;
assign _11537_ = _11187_ & _11534_ /*5425*/;
assign _11538_ = _11187_ ^ _11534_ /*5428*/;
assign _11539_ = _11530_ & _11538_ /*5426*/;
assign _11411_ = _11530_ ^ _11538_ /*5427*/;
assign _11536_ = _11537_ | _11539_ /*5424*/;
assign _11541_ = ~Q[6] /*5423*/;
assign _11540_ = _11541_ & D[19] /*5422*/;
assign _11543_ = _11188_ & _11540_ /*5417*/;
assign _11544_ = _11188_ ^ _11540_ /*5420*/;
assign _11545_ = _11536_ & _11544_ /*5418*/;
assign _11412_ = _11536_ ^ _11544_ /*5419*/;
assign _11542_ = _11543_ | _11545_ /*5416*/;
assign _11547_ = ~Q[6] /*5415*/;
assign _11546_ = _11547_ & D[20] /*5414*/;
assign _11549_ = _11189_ & _11546_ /*5409*/;
assign _11550_ = _11189_ ^ _11546_ /*5412*/;
assign _11551_ = _11542_ & _11550_ /*5410*/;
assign _11413_ = _11542_ ^ _11550_ /*5411*/;
assign _11548_ = _11549_ | _11551_ /*5408*/;
assign _11553_ = ~Q[6] /*5407*/;
assign _11552_ = _11553_ & D[21] /*5406*/;
assign _11555_ = _11190_ & _11552_ /*5401*/;
assign _11556_ = _11190_ ^ _11552_ /*5404*/;
assign _11557_ = _11548_ & _11556_ /*5402*/;
assign _11414_ = _11548_ ^ _11556_ /*5403*/;
assign _11554_ = _11555_ | _11557_ /*5400*/;
assign _11559_ = ~Q[6] /*5399*/;
assign _11558_ = _11559_ & D[22] /*5398*/;
assign _11561_ = _11191_ & _11558_ /*5393*/;
assign _11562_ = _11191_ ^ _11558_ /*5396*/;
assign _11563_ = _11554_ & _11562_ /*5394*/;
assign _11415_ = _11554_ ^ _11562_ /*5395*/;
assign _11560_ = _11561_ | _11563_ /*5392*/;
assign _11565_ = ~Q[6] /*5391*/;
assign _11564_ = _11565_ & D[23] /*5390*/;
assign _11567_ = _11192_ & _11564_ /*5385*/;
assign _11568_ = _11192_ ^ _11564_ /*5388*/;
assign _11569_ = _11560_ & _11568_ /*5386*/;
assign _11416_ = _11560_ ^ _11568_ /*5387*/;
assign _11566_ = _11567_ | _11569_ /*5384*/;
assign _11571_ = ~Q[6] /*5383*/;
assign _11570_ = _11571_ & D[24] /*5382*/;
assign _11573_ = _11193_ & _11570_ /*5377*/;
assign _11574_ = _11193_ ^ _11570_ /*5380*/;
assign _11575_ = _11566_ & _11574_ /*5378*/;
assign _11417_ = _11566_ ^ _11574_ /*5379*/;
assign _11572_ = _11573_ | _11575_ /*5376*/;
assign _11577_ = ~Q[6] /*5375*/;
assign _11576_ = _11577_ & D[25] /*5374*/;
assign _11579_ = _11194_ & _11576_ /*5369*/;
assign _11580_ = _11194_ ^ _11576_ /*5372*/;
assign _11581_ = _11572_ & _11580_ /*5370*/;
assign _11418_ = _11572_ ^ _11580_ /*5371*/;
assign _11578_ = _11579_ | _11581_ /*5368*/;
assign _11583_ = ~Q[6] /*5367*/;
assign _11582_ = _11583_ & D[26] /*5366*/;
assign _11585_ = _11195_ & _11582_ /*5361*/;
assign _11586_ = _11195_ ^ _11582_ /*5364*/;
assign _11587_ = _11578_ & _11586_ /*5362*/;
assign _11419_ = _11578_ ^ _11586_ /*5363*/;
assign _11584_ = _11585_ | _11587_ /*5360*/;
assign _11589_ = ~Q[6] /*5359*/;
assign _11588_ = _11589_ & D[27] /*5358*/;
assign _11591_ = _11196_ & _11588_ /*5353*/;
assign _11592_ = _11196_ ^ _11588_ /*5356*/;
assign _11593_ = _11584_ & _11592_ /*5354*/;
assign _11420_ = _11584_ ^ _11592_ /*5355*/;
assign _11590_ = _11591_ | _11593_ /*5352*/;
assign _11595_ = ~Q[6] /*5351*/;
assign _11594_ = _11595_ & D[28] /*5350*/;
assign _11597_ = _11197_ & _11594_ /*5345*/;
assign _11598_ = _11197_ ^ _11594_ /*5348*/;
assign _11599_ = _11590_ & _11598_ /*5346*/;
assign _11421_ = _11590_ ^ _11598_ /*5347*/;
assign _11596_ = _11597_ | _11599_ /*5344*/;
assign _11601_ = ~Q[6] /*5343*/;
assign _11600_ = _11601_ & D[29] /*5342*/;
assign _11603_ = _11198_ & _11600_ /*5337*/;
assign _11604_ = _11198_ ^ _11600_ /*5340*/;
assign _11605_ = _11596_ & _11604_ /*5338*/;
assign _11422_ = _11596_ ^ _11604_ /*5339*/;
assign _11602_ = _11603_ | _11605_ /*5336*/;
assign _11607_ = ~Q[6] /*5335*/;
assign _11606_ = _11607_ & D[30] /*5334*/;
assign _11609_ = _11199_ & _11606_ /*5329*/;
assign _11610_ = _11199_ ^ _11606_ /*5332*/;
assign _11611_ = _11602_ & _11610_ /*5330*/;
assign _11423_ = _11602_ ^ _11610_ /*5331*/;
assign _11608_ = _11609_ | _11611_ /*5328*/;
assign _11613_ = ~Q[6] /*5327*/;
assign _11612_ = _11613_ & zeroWire /*5326*/;
assign _11614_ = _11200_ ^ _11612_ /*5324*/;
assign _11424_ = _11614_ ^ _11608_ /*5323*/;
assign _11653_ = ~D[0] /*5197*/;
assign _11650_ = R_0[5] & _11653_ /*5193*/;
assign _11651_ = R_0[5] ^ _11653_ /*5196*/;
assign _11652_ = oneWire & _11651_ /*5194*/;
assign _11617_ = oneWire ^ _11651_ /*5195*/;
assign _11649_ = _11650_ | _11652_ /*5192*/;
assign _11658_ = ~D[1] /*5191*/;
assign _11655_ = _11393_ & _11658_ /*5187*/;
assign _11656_ = _11393_ ^ _11658_ /*5190*/;
assign _11657_ = _11649_ & _11656_ /*5188*/;
assign _11618_ = _11649_ ^ _11656_ /*5189*/;
assign _11654_ = _11655_ | _11657_ /*5186*/;
assign _11663_ = ~D[2] /*5185*/;
assign _11660_ = _11394_ & _11663_ /*5181*/;
assign _11661_ = _11394_ ^ _11663_ /*5184*/;
assign _11662_ = _11654_ & _11661_ /*5182*/;
assign _11619_ = _11654_ ^ _11661_ /*5183*/;
assign _11659_ = _11660_ | _11662_ /*5180*/;
assign _11668_ = ~D[3] /*5179*/;
assign _11665_ = _11395_ & _11668_ /*5175*/;
assign _11666_ = _11395_ ^ _11668_ /*5178*/;
assign _11667_ = _11659_ & _11666_ /*5176*/;
assign _11620_ = _11659_ ^ _11666_ /*5177*/;
assign _11664_ = _11665_ | _11667_ /*5174*/;
assign _11673_ = ~D[4] /*5173*/;
assign _11670_ = _11396_ & _11673_ /*5169*/;
assign _11671_ = _11396_ ^ _11673_ /*5172*/;
assign _11672_ = _11664_ & _11671_ /*5170*/;
assign _11621_ = _11664_ ^ _11671_ /*5171*/;
assign _11669_ = _11670_ | _11672_ /*5168*/;
assign _11678_ = ~D[5] /*5167*/;
assign _11675_ = _11397_ & _11678_ /*5163*/;
assign _11676_ = _11397_ ^ _11678_ /*5166*/;
assign _11677_ = _11669_ & _11676_ /*5164*/;
assign _11622_ = _11669_ ^ _11676_ /*5165*/;
assign _11674_ = _11675_ | _11677_ /*5162*/;
assign _11683_ = ~D[6] /*5161*/;
assign _11680_ = _11398_ & _11683_ /*5157*/;
assign _11681_ = _11398_ ^ _11683_ /*5160*/;
assign _11682_ = _11674_ & _11681_ /*5158*/;
assign _11623_ = _11674_ ^ _11681_ /*5159*/;
assign _11679_ = _11680_ | _11682_ /*5156*/;
assign _11688_ = ~D[7] /*5155*/;
assign _11685_ = _11399_ & _11688_ /*5151*/;
assign _11686_ = _11399_ ^ _11688_ /*5154*/;
assign _11687_ = _11679_ & _11686_ /*5152*/;
assign _11624_ = _11679_ ^ _11686_ /*5153*/;
assign _11684_ = _11685_ | _11687_ /*5150*/;
assign _11693_ = ~D[8] /*5149*/;
assign _11690_ = _11400_ & _11693_ /*5145*/;
assign _11691_ = _11400_ ^ _11693_ /*5148*/;
assign _11692_ = _11684_ & _11691_ /*5146*/;
assign _11625_ = _11684_ ^ _11691_ /*5147*/;
assign _11689_ = _11690_ | _11692_ /*5144*/;
assign _11698_ = ~D[9] /*5143*/;
assign _11695_ = _11401_ & _11698_ /*5139*/;
assign _11696_ = _11401_ ^ _11698_ /*5142*/;
assign _11697_ = _11689_ & _11696_ /*5140*/;
assign _11626_ = _11689_ ^ _11696_ /*5141*/;
assign _11694_ = _11695_ | _11697_ /*5138*/;
assign _11703_ = ~D[10] /*5137*/;
assign _11700_ = _11402_ & _11703_ /*5133*/;
assign _11701_ = _11402_ ^ _11703_ /*5136*/;
assign _11702_ = _11694_ & _11701_ /*5134*/;
assign _11627_ = _11694_ ^ _11701_ /*5135*/;
assign _11699_ = _11700_ | _11702_ /*5132*/;
assign _11708_ = ~D[11] /*5131*/;
assign _11705_ = _11403_ & _11708_ /*5127*/;
assign _11706_ = _11403_ ^ _11708_ /*5130*/;
assign _11707_ = _11699_ & _11706_ /*5128*/;
assign _11628_ = _11699_ ^ _11706_ /*5129*/;
assign _11704_ = _11705_ | _11707_ /*5126*/;
assign _11713_ = ~D[12] /*5125*/;
assign _11710_ = _11404_ & _11713_ /*5121*/;
assign _11711_ = _11404_ ^ _11713_ /*5124*/;
assign _11712_ = _11704_ & _11711_ /*5122*/;
assign _11629_ = _11704_ ^ _11711_ /*5123*/;
assign _11709_ = _11710_ | _11712_ /*5120*/;
assign _11718_ = ~D[13] /*5119*/;
assign _11715_ = _11405_ & _11718_ /*5115*/;
assign _11716_ = _11405_ ^ _11718_ /*5118*/;
assign _11717_ = _11709_ & _11716_ /*5116*/;
assign _11630_ = _11709_ ^ _11716_ /*5117*/;
assign _11714_ = _11715_ | _11717_ /*5114*/;
assign _11723_ = ~D[14] /*5113*/;
assign _11720_ = _11406_ & _11723_ /*5109*/;
assign _11721_ = _11406_ ^ _11723_ /*5112*/;
assign _11722_ = _11714_ & _11721_ /*5110*/;
assign _11631_ = _11714_ ^ _11721_ /*5111*/;
assign _11719_ = _11720_ | _11722_ /*5108*/;
assign _11728_ = ~D[15] /*5107*/;
assign _11725_ = _11407_ & _11728_ /*5103*/;
assign _11726_ = _11407_ ^ _11728_ /*5106*/;
assign _11727_ = _11719_ & _11726_ /*5104*/;
assign _11632_ = _11719_ ^ _11726_ /*5105*/;
assign _11724_ = _11725_ | _11727_ /*5102*/;
assign _11733_ = ~D[16] /*5101*/;
assign _11730_ = _11408_ & _11733_ /*5097*/;
assign _11731_ = _11408_ ^ _11733_ /*5100*/;
assign _11732_ = _11724_ & _11731_ /*5098*/;
assign _11633_ = _11724_ ^ _11731_ /*5099*/;
assign _11729_ = _11730_ | _11732_ /*5096*/;
assign _11738_ = ~D[17] /*5095*/;
assign _11735_ = _11409_ & _11738_ /*5091*/;
assign _11736_ = _11409_ ^ _11738_ /*5094*/;
assign _11737_ = _11729_ & _11736_ /*5092*/;
assign _11634_ = _11729_ ^ _11736_ /*5093*/;
assign _11734_ = _11735_ | _11737_ /*5090*/;
assign _11743_ = ~D[18] /*5089*/;
assign _11740_ = _11410_ & _11743_ /*5085*/;
assign _11741_ = _11410_ ^ _11743_ /*5088*/;
assign _11742_ = _11734_ & _11741_ /*5086*/;
assign _11635_ = _11734_ ^ _11741_ /*5087*/;
assign _11739_ = _11740_ | _11742_ /*5084*/;
assign _11748_ = ~D[19] /*5083*/;
assign _11745_ = _11411_ & _11748_ /*5079*/;
assign _11746_ = _11411_ ^ _11748_ /*5082*/;
assign _11747_ = _11739_ & _11746_ /*5080*/;
assign _11636_ = _11739_ ^ _11746_ /*5081*/;
assign _11744_ = _11745_ | _11747_ /*5078*/;
assign _11753_ = ~D[20] /*5077*/;
assign _11750_ = _11412_ & _11753_ /*5073*/;
assign _11751_ = _11412_ ^ _11753_ /*5076*/;
assign _11752_ = _11744_ & _11751_ /*5074*/;
assign _11637_ = _11744_ ^ _11751_ /*5075*/;
assign _11749_ = _11750_ | _11752_ /*5072*/;
assign _11758_ = ~D[21] /*5071*/;
assign _11755_ = _11413_ & _11758_ /*5067*/;
assign _11756_ = _11413_ ^ _11758_ /*5070*/;
assign _11757_ = _11749_ & _11756_ /*5068*/;
assign _11638_ = _11749_ ^ _11756_ /*5069*/;
assign _11754_ = _11755_ | _11757_ /*5066*/;
assign _11763_ = ~D[22] /*5065*/;
assign _11760_ = _11414_ & _11763_ /*5061*/;
assign _11761_ = _11414_ ^ _11763_ /*5064*/;
assign _11762_ = _11754_ & _11761_ /*5062*/;
assign _11639_ = _11754_ ^ _11761_ /*5063*/;
assign _11759_ = _11760_ | _11762_ /*5060*/;
assign _11768_ = ~D[23] /*5059*/;
assign _11765_ = _11415_ & _11768_ /*5055*/;
assign _11766_ = _11415_ ^ _11768_ /*5058*/;
assign _11767_ = _11759_ & _11766_ /*5056*/;
assign _11640_ = _11759_ ^ _11766_ /*5057*/;
assign _11764_ = _11765_ | _11767_ /*5054*/;
assign _11773_ = ~D[24] /*5053*/;
assign _11770_ = _11416_ & _11773_ /*5049*/;
assign _11771_ = _11416_ ^ _11773_ /*5052*/;
assign _11772_ = _11764_ & _11771_ /*5050*/;
assign _11641_ = _11764_ ^ _11771_ /*5051*/;
assign _11769_ = _11770_ | _11772_ /*5048*/;
assign _11778_ = ~D[25] /*5047*/;
assign _11775_ = _11417_ & _11778_ /*5043*/;
assign _11776_ = _11417_ ^ _11778_ /*5046*/;
assign _11777_ = _11769_ & _11776_ /*5044*/;
assign _11642_ = _11769_ ^ _11776_ /*5045*/;
assign _11774_ = _11775_ | _11777_ /*5042*/;
assign _11783_ = ~D[26] /*5041*/;
assign _11780_ = _11418_ & _11783_ /*5037*/;
assign _11781_ = _11418_ ^ _11783_ /*5040*/;
assign _11782_ = _11774_ & _11781_ /*5038*/;
assign _11643_ = _11774_ ^ _11781_ /*5039*/;
assign _11779_ = _11780_ | _11782_ /*5036*/;
assign _11788_ = ~D[27] /*5035*/;
assign _11785_ = _11419_ & _11788_ /*5031*/;
assign _11786_ = _11419_ ^ _11788_ /*5034*/;
assign _11787_ = _11779_ & _11786_ /*5032*/;
assign _11644_ = _11779_ ^ _11786_ /*5033*/;
assign _11784_ = _11785_ | _11787_ /*5030*/;
assign _11793_ = ~D[28] /*5029*/;
assign _11790_ = _11420_ & _11793_ /*5025*/;
assign _11791_ = _11420_ ^ _11793_ /*5028*/;
assign _11792_ = _11784_ & _11791_ /*5026*/;
assign _11645_ = _11784_ ^ _11791_ /*5027*/;
assign _11789_ = _11790_ | _11792_ /*5024*/;
assign _11798_ = ~D[29] /*5023*/;
assign _11795_ = _11421_ & _11798_ /*5019*/;
assign _11796_ = _11421_ ^ _11798_ /*5022*/;
assign _11797_ = _11789_ & _11796_ /*5020*/;
assign _11646_ = _11789_ ^ _11796_ /*5021*/;
assign _11794_ = _11795_ | _11797_ /*5018*/;
assign _11803_ = ~D[30] /*5017*/;
assign _11800_ = _11422_ & _11803_ /*5013*/;
assign _11801_ = _11422_ ^ _11803_ /*5016*/;
assign _11802_ = _11794_ & _11801_ /*5014*/;
assign _11647_ = _11794_ ^ _11801_ /*5015*/;
assign _11799_ = _11800_ | _11802_ /*5012*/;
assign _11804_ = _11423_ & oneWire /*5007*/;
assign _11805_ = _11423_ ^ oneWire /*5010*/;
assign _11806_ = _11799_ & _11805_ /*5008*/;
assign _11648_ = _11799_ ^ _11805_ /*5009*/;
assign Q[5] = _11804_ | _11806_ /*5006*/;
assign _11875_ = ~Q[5] /*4813*/;
assign _11874_ = _11875_ & D[0] /*4812*/;
assign _11877_ = _11617_ & _11874_ /*4807*/;
assign _11878_ = _11617_ ^ _11874_ /*4810*/;
assign _11879_ = zeroWire & _11878_ /*4808*/;
assign _11841_ = zeroWire ^ _11878_ /*4809*/;
assign _11876_ = _11877_ | _11879_ /*4806*/;
assign _11881_ = ~Q[5] /*4805*/;
assign _11880_ = _11881_ & D[1] /*4804*/;
assign _11883_ = _11618_ & _11880_ /*4799*/;
assign _11884_ = _11618_ ^ _11880_ /*4802*/;
assign _11885_ = _11876_ & _11884_ /*4800*/;
assign _11842_ = _11876_ ^ _11884_ /*4801*/;
assign _11882_ = _11883_ | _11885_ /*4798*/;
assign _11887_ = ~Q[5] /*4797*/;
assign _11886_ = _11887_ & D[2] /*4796*/;
assign _11889_ = _11619_ & _11886_ /*4791*/;
assign _11890_ = _11619_ ^ _11886_ /*4794*/;
assign _11891_ = _11882_ & _11890_ /*4792*/;
assign _11843_ = _11882_ ^ _11890_ /*4793*/;
assign _11888_ = _11889_ | _11891_ /*4790*/;
assign _11893_ = ~Q[5] /*4789*/;
assign _11892_ = _11893_ & D[3] /*4788*/;
assign _11895_ = _11620_ & _11892_ /*4783*/;
assign _11896_ = _11620_ ^ _11892_ /*4786*/;
assign _11897_ = _11888_ & _11896_ /*4784*/;
assign _11844_ = _11888_ ^ _11896_ /*4785*/;
assign _11894_ = _11895_ | _11897_ /*4782*/;
assign _11899_ = ~Q[5] /*4781*/;
assign _11898_ = _11899_ & D[4] /*4780*/;
assign _11901_ = _11621_ & _11898_ /*4775*/;
assign _11902_ = _11621_ ^ _11898_ /*4778*/;
assign _11903_ = _11894_ & _11902_ /*4776*/;
assign _11845_ = _11894_ ^ _11902_ /*4777*/;
assign _11900_ = _11901_ | _11903_ /*4774*/;
assign _11905_ = ~Q[5] /*4773*/;
assign _11904_ = _11905_ & D[5] /*4772*/;
assign _11907_ = _11622_ & _11904_ /*4767*/;
assign _11908_ = _11622_ ^ _11904_ /*4770*/;
assign _11909_ = _11900_ & _11908_ /*4768*/;
assign _11846_ = _11900_ ^ _11908_ /*4769*/;
assign _11906_ = _11907_ | _11909_ /*4766*/;
assign _11911_ = ~Q[5] /*4765*/;
assign _11910_ = _11911_ & D[6] /*4764*/;
assign _11913_ = _11623_ & _11910_ /*4759*/;
assign _11914_ = _11623_ ^ _11910_ /*4762*/;
assign _11915_ = _11906_ & _11914_ /*4760*/;
assign _11847_ = _11906_ ^ _11914_ /*4761*/;
assign _11912_ = _11913_ | _11915_ /*4758*/;
assign _11917_ = ~Q[5] /*4757*/;
assign _11916_ = _11917_ & D[7] /*4756*/;
assign _11919_ = _11624_ & _11916_ /*4751*/;
assign _11920_ = _11624_ ^ _11916_ /*4754*/;
assign _11921_ = _11912_ & _11920_ /*4752*/;
assign _11848_ = _11912_ ^ _11920_ /*4753*/;
assign _11918_ = _11919_ | _11921_ /*4750*/;
assign _11923_ = ~Q[5] /*4749*/;
assign _11922_ = _11923_ & D[8] /*4748*/;
assign _11925_ = _11625_ & _11922_ /*4743*/;
assign _11926_ = _11625_ ^ _11922_ /*4746*/;
assign _11927_ = _11918_ & _11926_ /*4744*/;
assign _11849_ = _11918_ ^ _11926_ /*4745*/;
assign _11924_ = _11925_ | _11927_ /*4742*/;
assign _11929_ = ~Q[5] /*4741*/;
assign _11928_ = _11929_ & D[9] /*4740*/;
assign _11931_ = _11626_ & _11928_ /*4735*/;
assign _11932_ = _11626_ ^ _11928_ /*4738*/;
assign _11933_ = _11924_ & _11932_ /*4736*/;
assign _11850_ = _11924_ ^ _11932_ /*4737*/;
assign _11930_ = _11931_ | _11933_ /*4734*/;
assign _11935_ = ~Q[5] /*4733*/;
assign _11934_ = _11935_ & D[10] /*4732*/;
assign _11937_ = _11627_ & _11934_ /*4727*/;
assign _11938_ = _11627_ ^ _11934_ /*4730*/;
assign _11939_ = _11930_ & _11938_ /*4728*/;
assign _11851_ = _11930_ ^ _11938_ /*4729*/;
assign _11936_ = _11937_ | _11939_ /*4726*/;
assign _11941_ = ~Q[5] /*4725*/;
assign _11940_ = _11941_ & D[11] /*4724*/;
assign _11943_ = _11628_ & _11940_ /*4719*/;
assign _11944_ = _11628_ ^ _11940_ /*4722*/;
assign _11945_ = _11936_ & _11944_ /*4720*/;
assign _11852_ = _11936_ ^ _11944_ /*4721*/;
assign _11942_ = _11943_ | _11945_ /*4718*/;
assign _11947_ = ~Q[5] /*4717*/;
assign _11946_ = _11947_ & D[12] /*4716*/;
assign _11949_ = _11629_ & _11946_ /*4711*/;
assign _11950_ = _11629_ ^ _11946_ /*4714*/;
assign _11951_ = _11942_ & _11950_ /*4712*/;
assign _11853_ = _11942_ ^ _11950_ /*4713*/;
assign _11948_ = _11949_ | _11951_ /*4710*/;
assign _11953_ = ~Q[5] /*4709*/;
assign _11952_ = _11953_ & D[13] /*4708*/;
assign _11955_ = _11630_ & _11952_ /*4703*/;
assign _11956_ = _11630_ ^ _11952_ /*4706*/;
assign _11957_ = _11948_ & _11956_ /*4704*/;
assign _11854_ = _11948_ ^ _11956_ /*4705*/;
assign _11954_ = _11955_ | _11957_ /*4702*/;
assign _11959_ = ~Q[5] /*4701*/;
assign _11958_ = _11959_ & D[14] /*4700*/;
assign _11961_ = _11631_ & _11958_ /*4695*/;
assign _11962_ = _11631_ ^ _11958_ /*4698*/;
assign _11963_ = _11954_ & _11962_ /*4696*/;
assign _11855_ = _11954_ ^ _11962_ /*4697*/;
assign _11960_ = _11961_ | _11963_ /*4694*/;
assign _11965_ = ~Q[5] /*4693*/;
assign _11964_ = _11965_ & D[15] /*4692*/;
assign _11967_ = _11632_ & _11964_ /*4687*/;
assign _11968_ = _11632_ ^ _11964_ /*4690*/;
assign _11969_ = _11960_ & _11968_ /*4688*/;
assign _11856_ = _11960_ ^ _11968_ /*4689*/;
assign _11966_ = _11967_ | _11969_ /*4686*/;
assign _11971_ = ~Q[5] /*4685*/;
assign _11970_ = _11971_ & D[16] /*4684*/;
assign _11973_ = _11633_ & _11970_ /*4679*/;
assign _11974_ = _11633_ ^ _11970_ /*4682*/;
assign _11975_ = _11966_ & _11974_ /*4680*/;
assign _11857_ = _11966_ ^ _11974_ /*4681*/;
assign _11972_ = _11973_ | _11975_ /*4678*/;
assign _11977_ = ~Q[5] /*4677*/;
assign _11976_ = _11977_ & D[17] /*4676*/;
assign _11979_ = _11634_ & _11976_ /*4671*/;
assign _11980_ = _11634_ ^ _11976_ /*4674*/;
assign _11981_ = _11972_ & _11980_ /*4672*/;
assign _11858_ = _11972_ ^ _11980_ /*4673*/;
assign _11978_ = _11979_ | _11981_ /*4670*/;
assign _11983_ = ~Q[5] /*4669*/;
assign _11982_ = _11983_ & D[18] /*4668*/;
assign _11985_ = _11635_ & _11982_ /*4663*/;
assign _11986_ = _11635_ ^ _11982_ /*4666*/;
assign _11987_ = _11978_ & _11986_ /*4664*/;
assign _11859_ = _11978_ ^ _11986_ /*4665*/;
assign _11984_ = _11985_ | _11987_ /*4662*/;
assign _11989_ = ~Q[5] /*4661*/;
assign _11988_ = _11989_ & D[19] /*4660*/;
assign _11991_ = _11636_ & _11988_ /*4655*/;
assign _11992_ = _11636_ ^ _11988_ /*4658*/;
assign _11993_ = _11984_ & _11992_ /*4656*/;
assign _11860_ = _11984_ ^ _11992_ /*4657*/;
assign _11990_ = _11991_ | _11993_ /*4654*/;
assign _11995_ = ~Q[5] /*4653*/;
assign _11994_ = _11995_ & D[20] /*4652*/;
assign _11997_ = _11637_ & _11994_ /*4647*/;
assign _11998_ = _11637_ ^ _11994_ /*4650*/;
assign _11999_ = _11990_ & _11998_ /*4648*/;
assign _11861_ = _11990_ ^ _11998_ /*4649*/;
assign _11996_ = _11997_ | _11999_ /*4646*/;
assign _12001_ = ~Q[5] /*4645*/;
assign _12000_ = _12001_ & D[21] /*4644*/;
assign _12003_ = _11638_ & _12000_ /*4639*/;
assign _12004_ = _11638_ ^ _12000_ /*4642*/;
assign _12005_ = _11996_ & _12004_ /*4640*/;
assign _11862_ = _11996_ ^ _12004_ /*4641*/;
assign _12002_ = _12003_ | _12005_ /*4638*/;
assign _12007_ = ~Q[5] /*4637*/;
assign _12006_ = _12007_ & D[22] /*4636*/;
assign _12009_ = _11639_ & _12006_ /*4631*/;
assign _12010_ = _11639_ ^ _12006_ /*4634*/;
assign _12011_ = _12002_ & _12010_ /*4632*/;
assign _11863_ = _12002_ ^ _12010_ /*4633*/;
assign _12008_ = _12009_ | _12011_ /*4630*/;
assign _12013_ = ~Q[5] /*4629*/;
assign _12012_ = _12013_ & D[23] /*4628*/;
assign _12015_ = _11640_ & _12012_ /*4623*/;
assign _12016_ = _11640_ ^ _12012_ /*4626*/;
assign _12017_ = _12008_ & _12016_ /*4624*/;
assign _11864_ = _12008_ ^ _12016_ /*4625*/;
assign _12014_ = _12015_ | _12017_ /*4622*/;
assign _12019_ = ~Q[5] /*4621*/;
assign _12018_ = _12019_ & D[24] /*4620*/;
assign _12021_ = _11641_ & _12018_ /*4615*/;
assign _12022_ = _11641_ ^ _12018_ /*4618*/;
assign _12023_ = _12014_ & _12022_ /*4616*/;
assign _11865_ = _12014_ ^ _12022_ /*4617*/;
assign _12020_ = _12021_ | _12023_ /*4614*/;
assign _12025_ = ~Q[5] /*4613*/;
assign _12024_ = _12025_ & D[25] /*4612*/;
assign _12027_ = _11642_ & _12024_ /*4607*/;
assign _12028_ = _11642_ ^ _12024_ /*4610*/;
assign _12029_ = _12020_ & _12028_ /*4608*/;
assign _11866_ = _12020_ ^ _12028_ /*4609*/;
assign _12026_ = _12027_ | _12029_ /*4606*/;
assign _12031_ = ~Q[5] /*4605*/;
assign _12030_ = _12031_ & D[26] /*4604*/;
assign _12033_ = _11643_ & _12030_ /*4599*/;
assign _12034_ = _11643_ ^ _12030_ /*4602*/;
assign _12035_ = _12026_ & _12034_ /*4600*/;
assign _11867_ = _12026_ ^ _12034_ /*4601*/;
assign _12032_ = _12033_ | _12035_ /*4598*/;
assign _12037_ = ~Q[5] /*4597*/;
assign _12036_ = _12037_ & D[27] /*4596*/;
assign _12039_ = _11644_ & _12036_ /*4591*/;
assign _12040_ = _11644_ ^ _12036_ /*4594*/;
assign _12041_ = _12032_ & _12040_ /*4592*/;
assign _11868_ = _12032_ ^ _12040_ /*4593*/;
assign _12038_ = _12039_ | _12041_ /*4590*/;
assign _12043_ = ~Q[5] /*4589*/;
assign _12042_ = _12043_ & D[28] /*4588*/;
assign _12045_ = _11645_ & _12042_ /*4583*/;
assign _12046_ = _11645_ ^ _12042_ /*4586*/;
assign _12047_ = _12038_ & _12046_ /*4584*/;
assign _11869_ = _12038_ ^ _12046_ /*4585*/;
assign _12044_ = _12045_ | _12047_ /*4582*/;
assign _12049_ = ~Q[5] /*4581*/;
assign _12048_ = _12049_ & D[29] /*4580*/;
assign _12051_ = _11646_ & _12048_ /*4575*/;
assign _12052_ = _11646_ ^ _12048_ /*4578*/;
assign _12053_ = _12044_ & _12052_ /*4576*/;
assign _11870_ = _12044_ ^ _12052_ /*4577*/;
assign _12050_ = _12051_ | _12053_ /*4574*/;
assign _12055_ = ~Q[5] /*4573*/;
assign _12054_ = _12055_ & D[30] /*4572*/;
assign _12057_ = _11647_ & _12054_ /*4567*/;
assign _12058_ = _11647_ ^ _12054_ /*4570*/;
assign _12059_ = _12050_ & _12058_ /*4568*/;
assign _11871_ = _12050_ ^ _12058_ /*4569*/;
assign _12056_ = _12057_ | _12059_ /*4566*/;
assign _12061_ = ~Q[5] /*4565*/;
assign _12060_ = _12061_ & zeroWire /*4564*/;
assign _12062_ = _11648_ ^ _12060_ /*4562*/;
assign _11872_ = _12062_ ^ _12056_ /*4561*/;
assign _12101_ = ~D[0] /*4435*/;
assign _12098_ = R_0[4] & _12101_ /*4431*/;
assign _12099_ = R_0[4] ^ _12101_ /*4434*/;
assign _12100_ = oneWire & _12099_ /*4432*/;
assign _12065_ = oneWire ^ _12099_ /*4433*/;
assign _12097_ = _12098_ | _12100_ /*4430*/;
assign _12106_ = ~D[1] /*4429*/;
assign _12103_ = _11841_ & _12106_ /*4425*/;
assign _12104_ = _11841_ ^ _12106_ /*4428*/;
assign _12105_ = _12097_ & _12104_ /*4426*/;
assign _12066_ = _12097_ ^ _12104_ /*4427*/;
assign _12102_ = _12103_ | _12105_ /*4424*/;
assign _12111_ = ~D[2] /*4423*/;
assign _12108_ = _11842_ & _12111_ /*4419*/;
assign _12109_ = _11842_ ^ _12111_ /*4422*/;
assign _12110_ = _12102_ & _12109_ /*4420*/;
assign _12067_ = _12102_ ^ _12109_ /*4421*/;
assign _12107_ = _12108_ | _12110_ /*4418*/;
assign _12116_ = ~D[3] /*4417*/;
assign _12113_ = _11843_ & _12116_ /*4413*/;
assign _12114_ = _11843_ ^ _12116_ /*4416*/;
assign _12115_ = _12107_ & _12114_ /*4414*/;
assign _12068_ = _12107_ ^ _12114_ /*4415*/;
assign _12112_ = _12113_ | _12115_ /*4412*/;
assign _12121_ = ~D[4] /*4411*/;
assign _12118_ = _11844_ & _12121_ /*4407*/;
assign _12119_ = _11844_ ^ _12121_ /*4410*/;
assign _12120_ = _12112_ & _12119_ /*4408*/;
assign _12069_ = _12112_ ^ _12119_ /*4409*/;
assign _12117_ = _12118_ | _12120_ /*4406*/;
assign _12126_ = ~D[5] /*4405*/;
assign _12123_ = _11845_ & _12126_ /*4401*/;
assign _12124_ = _11845_ ^ _12126_ /*4404*/;
assign _12125_ = _12117_ & _12124_ /*4402*/;
assign _12070_ = _12117_ ^ _12124_ /*4403*/;
assign _12122_ = _12123_ | _12125_ /*4400*/;
assign _12131_ = ~D[6] /*4399*/;
assign _12128_ = _11846_ & _12131_ /*4395*/;
assign _12129_ = _11846_ ^ _12131_ /*4398*/;
assign _12130_ = _12122_ & _12129_ /*4396*/;
assign _12071_ = _12122_ ^ _12129_ /*4397*/;
assign _12127_ = _12128_ | _12130_ /*4394*/;
assign _12136_ = ~D[7] /*4393*/;
assign _12133_ = _11847_ & _12136_ /*4389*/;
assign _12134_ = _11847_ ^ _12136_ /*4392*/;
assign _12135_ = _12127_ & _12134_ /*4390*/;
assign _12072_ = _12127_ ^ _12134_ /*4391*/;
assign _12132_ = _12133_ | _12135_ /*4388*/;
assign _12141_ = ~D[8] /*4387*/;
assign _12138_ = _11848_ & _12141_ /*4383*/;
assign _12139_ = _11848_ ^ _12141_ /*4386*/;
assign _12140_ = _12132_ & _12139_ /*4384*/;
assign _12073_ = _12132_ ^ _12139_ /*4385*/;
assign _12137_ = _12138_ | _12140_ /*4382*/;
assign _12146_ = ~D[9] /*4381*/;
assign _12143_ = _11849_ & _12146_ /*4377*/;
assign _12144_ = _11849_ ^ _12146_ /*4380*/;
assign _12145_ = _12137_ & _12144_ /*4378*/;
assign _12074_ = _12137_ ^ _12144_ /*4379*/;
assign _12142_ = _12143_ | _12145_ /*4376*/;
assign _12151_ = ~D[10] /*4375*/;
assign _12148_ = _11850_ & _12151_ /*4371*/;
assign _12149_ = _11850_ ^ _12151_ /*4374*/;
assign _12150_ = _12142_ & _12149_ /*4372*/;
assign _12075_ = _12142_ ^ _12149_ /*4373*/;
assign _12147_ = _12148_ | _12150_ /*4370*/;
assign _12156_ = ~D[11] /*4369*/;
assign _12153_ = _11851_ & _12156_ /*4365*/;
assign _12154_ = _11851_ ^ _12156_ /*4368*/;
assign _12155_ = _12147_ & _12154_ /*4366*/;
assign _12076_ = _12147_ ^ _12154_ /*4367*/;
assign _12152_ = _12153_ | _12155_ /*4364*/;
assign _12161_ = ~D[12] /*4363*/;
assign _12158_ = _11852_ & _12161_ /*4359*/;
assign _12159_ = _11852_ ^ _12161_ /*4362*/;
assign _12160_ = _12152_ & _12159_ /*4360*/;
assign _12077_ = _12152_ ^ _12159_ /*4361*/;
assign _12157_ = _12158_ | _12160_ /*4358*/;
assign _12166_ = ~D[13] /*4357*/;
assign _12163_ = _11853_ & _12166_ /*4353*/;
assign _12164_ = _11853_ ^ _12166_ /*4356*/;
assign _12165_ = _12157_ & _12164_ /*4354*/;
assign _12078_ = _12157_ ^ _12164_ /*4355*/;
assign _12162_ = _12163_ | _12165_ /*4352*/;
assign _12171_ = ~D[14] /*4351*/;
assign _12168_ = _11854_ & _12171_ /*4347*/;
assign _12169_ = _11854_ ^ _12171_ /*4350*/;
assign _12170_ = _12162_ & _12169_ /*4348*/;
assign _12079_ = _12162_ ^ _12169_ /*4349*/;
assign _12167_ = _12168_ | _12170_ /*4346*/;
assign _12176_ = ~D[15] /*4345*/;
assign _12173_ = _11855_ & _12176_ /*4341*/;
assign _12174_ = _11855_ ^ _12176_ /*4344*/;
assign _12175_ = _12167_ & _12174_ /*4342*/;
assign _12080_ = _12167_ ^ _12174_ /*4343*/;
assign _12172_ = _12173_ | _12175_ /*4340*/;
assign _12181_ = ~D[16] /*4339*/;
assign _12178_ = _11856_ & _12181_ /*4335*/;
assign _12179_ = _11856_ ^ _12181_ /*4338*/;
assign _12180_ = _12172_ & _12179_ /*4336*/;
assign _12081_ = _12172_ ^ _12179_ /*4337*/;
assign _12177_ = _12178_ | _12180_ /*4334*/;
assign _12186_ = ~D[17] /*4333*/;
assign _12183_ = _11857_ & _12186_ /*4329*/;
assign _12184_ = _11857_ ^ _12186_ /*4332*/;
assign _12185_ = _12177_ & _12184_ /*4330*/;
assign _12082_ = _12177_ ^ _12184_ /*4331*/;
assign _12182_ = _12183_ | _12185_ /*4328*/;
assign _12191_ = ~D[18] /*4327*/;
assign _12188_ = _11858_ & _12191_ /*4323*/;
assign _12189_ = _11858_ ^ _12191_ /*4326*/;
assign _12190_ = _12182_ & _12189_ /*4324*/;
assign _12083_ = _12182_ ^ _12189_ /*4325*/;
assign _12187_ = _12188_ | _12190_ /*4322*/;
assign _12196_ = ~D[19] /*4321*/;
assign _12193_ = _11859_ & _12196_ /*4317*/;
assign _12194_ = _11859_ ^ _12196_ /*4320*/;
assign _12195_ = _12187_ & _12194_ /*4318*/;
assign _12084_ = _12187_ ^ _12194_ /*4319*/;
assign _12192_ = _12193_ | _12195_ /*4316*/;
assign _12201_ = ~D[20] /*4315*/;
assign _12198_ = _11860_ & _12201_ /*4311*/;
assign _12199_ = _11860_ ^ _12201_ /*4314*/;
assign _12200_ = _12192_ & _12199_ /*4312*/;
assign _12085_ = _12192_ ^ _12199_ /*4313*/;
assign _12197_ = _12198_ | _12200_ /*4310*/;
assign _12206_ = ~D[21] /*4309*/;
assign _12203_ = _11861_ & _12206_ /*4305*/;
assign _12204_ = _11861_ ^ _12206_ /*4308*/;
assign _12205_ = _12197_ & _12204_ /*4306*/;
assign _12086_ = _12197_ ^ _12204_ /*4307*/;
assign _12202_ = _12203_ | _12205_ /*4304*/;
assign _12211_ = ~D[22] /*4303*/;
assign _12208_ = _11862_ & _12211_ /*4299*/;
assign _12209_ = _11862_ ^ _12211_ /*4302*/;
assign _12210_ = _12202_ & _12209_ /*4300*/;
assign _12087_ = _12202_ ^ _12209_ /*4301*/;
assign _12207_ = _12208_ | _12210_ /*4298*/;
assign _12216_ = ~D[23] /*4297*/;
assign _12213_ = _11863_ & _12216_ /*4293*/;
assign _12214_ = _11863_ ^ _12216_ /*4296*/;
assign _12215_ = _12207_ & _12214_ /*4294*/;
assign _12088_ = _12207_ ^ _12214_ /*4295*/;
assign _12212_ = _12213_ | _12215_ /*4292*/;
assign _12221_ = ~D[24] /*4291*/;
assign _12218_ = _11864_ & _12221_ /*4287*/;
assign _12219_ = _11864_ ^ _12221_ /*4290*/;
assign _12220_ = _12212_ & _12219_ /*4288*/;
assign _12089_ = _12212_ ^ _12219_ /*4289*/;
assign _12217_ = _12218_ | _12220_ /*4286*/;
assign _12226_ = ~D[25] /*4285*/;
assign _12223_ = _11865_ & _12226_ /*4281*/;
assign _12224_ = _11865_ ^ _12226_ /*4284*/;
assign _12225_ = _12217_ & _12224_ /*4282*/;
assign _12090_ = _12217_ ^ _12224_ /*4283*/;
assign _12222_ = _12223_ | _12225_ /*4280*/;
assign _12231_ = ~D[26] /*4279*/;
assign _12228_ = _11866_ & _12231_ /*4275*/;
assign _12229_ = _11866_ ^ _12231_ /*4278*/;
assign _12230_ = _12222_ & _12229_ /*4276*/;
assign _12091_ = _12222_ ^ _12229_ /*4277*/;
assign _12227_ = _12228_ | _12230_ /*4274*/;
assign _12236_ = ~D[27] /*4273*/;
assign _12233_ = _11867_ & _12236_ /*4269*/;
assign _12234_ = _11867_ ^ _12236_ /*4272*/;
assign _12235_ = _12227_ & _12234_ /*4270*/;
assign _12092_ = _12227_ ^ _12234_ /*4271*/;
assign _12232_ = _12233_ | _12235_ /*4268*/;
assign _12241_ = ~D[28] /*4267*/;
assign _12238_ = _11868_ & _12241_ /*4263*/;
assign _12239_ = _11868_ ^ _12241_ /*4266*/;
assign _12240_ = _12232_ & _12239_ /*4264*/;
assign _12093_ = _12232_ ^ _12239_ /*4265*/;
assign _12237_ = _12238_ | _12240_ /*4262*/;
assign _12246_ = ~D[29] /*4261*/;
assign _12243_ = _11869_ & _12246_ /*4257*/;
assign _12244_ = _11869_ ^ _12246_ /*4260*/;
assign _12245_ = _12237_ & _12244_ /*4258*/;
assign _12094_ = _12237_ ^ _12244_ /*4259*/;
assign _12242_ = _12243_ | _12245_ /*4256*/;
assign _12251_ = ~D[30] /*4255*/;
assign _12248_ = _11870_ & _12251_ /*4251*/;
assign _12249_ = _11870_ ^ _12251_ /*4254*/;
assign _12250_ = _12242_ & _12249_ /*4252*/;
assign _12095_ = _12242_ ^ _12249_ /*4253*/;
assign _12247_ = _12248_ | _12250_ /*4250*/;
assign _12252_ = _11871_ & oneWire /*4245*/;
assign _12253_ = _11871_ ^ oneWire /*4248*/;
assign _12254_ = _12247_ & _12253_ /*4246*/;
assign _12096_ = _12247_ ^ _12253_ /*4247*/;
assign Q[4] = _12252_ | _12254_ /*4244*/;
assign _12323_ = ~Q[4] /*4051*/;
assign _12322_ = _12323_ & D[0] /*4050*/;
assign _12325_ = _12065_ & _12322_ /*4045*/;
assign _12326_ = _12065_ ^ _12322_ /*4048*/;
assign _12327_ = zeroWire & _12326_ /*4046*/;
assign _12289_ = zeroWire ^ _12326_ /*4047*/;
assign _12324_ = _12325_ | _12327_ /*4044*/;
assign _12329_ = ~Q[4] /*4043*/;
assign _12328_ = _12329_ & D[1] /*4042*/;
assign _12331_ = _12066_ & _12328_ /*4037*/;
assign _12332_ = _12066_ ^ _12328_ /*4040*/;
assign _12333_ = _12324_ & _12332_ /*4038*/;
assign _12290_ = _12324_ ^ _12332_ /*4039*/;
assign _12330_ = _12331_ | _12333_ /*4036*/;
assign _12335_ = ~Q[4] /*4035*/;
assign _12334_ = _12335_ & D[2] /*4034*/;
assign _12337_ = _12067_ & _12334_ /*4029*/;
assign _12338_ = _12067_ ^ _12334_ /*4032*/;
assign _12339_ = _12330_ & _12338_ /*4030*/;
assign _12291_ = _12330_ ^ _12338_ /*4031*/;
assign _12336_ = _12337_ | _12339_ /*4028*/;
assign _12341_ = ~Q[4] /*4027*/;
assign _12340_ = _12341_ & D[3] /*4026*/;
assign _12343_ = _12068_ & _12340_ /*4021*/;
assign _12344_ = _12068_ ^ _12340_ /*4024*/;
assign _12345_ = _12336_ & _12344_ /*4022*/;
assign _12292_ = _12336_ ^ _12344_ /*4023*/;
assign _12342_ = _12343_ | _12345_ /*4020*/;
assign _12347_ = ~Q[4] /*4019*/;
assign _12346_ = _12347_ & D[4] /*4018*/;
assign _12349_ = _12069_ & _12346_ /*4013*/;
assign _12350_ = _12069_ ^ _12346_ /*4016*/;
assign _12351_ = _12342_ & _12350_ /*4014*/;
assign _12293_ = _12342_ ^ _12350_ /*4015*/;
assign _12348_ = _12349_ | _12351_ /*4012*/;
assign _12353_ = ~Q[4] /*4011*/;
assign _12352_ = _12353_ & D[5] /*4010*/;
assign _12355_ = _12070_ & _12352_ /*4005*/;
assign _12356_ = _12070_ ^ _12352_ /*4008*/;
assign _12357_ = _12348_ & _12356_ /*4006*/;
assign _12294_ = _12348_ ^ _12356_ /*4007*/;
assign _12354_ = _12355_ | _12357_ /*4004*/;
assign _12359_ = ~Q[4] /*4003*/;
assign _12358_ = _12359_ & D[6] /*4002*/;
assign _12361_ = _12071_ & _12358_ /*3997*/;
assign _12362_ = _12071_ ^ _12358_ /*4000*/;
assign _12363_ = _12354_ & _12362_ /*3998*/;
assign _12295_ = _12354_ ^ _12362_ /*3999*/;
assign _12360_ = _12361_ | _12363_ /*3996*/;
assign _12365_ = ~Q[4] /*3995*/;
assign _12364_ = _12365_ & D[7] /*3994*/;
assign _12367_ = _12072_ & _12364_ /*3989*/;
assign _12368_ = _12072_ ^ _12364_ /*3992*/;
assign _12369_ = _12360_ & _12368_ /*3990*/;
assign _12296_ = _12360_ ^ _12368_ /*3991*/;
assign _12366_ = _12367_ | _12369_ /*3988*/;
assign _12371_ = ~Q[4] /*3987*/;
assign _12370_ = _12371_ & D[8] /*3986*/;
assign _12373_ = _12073_ & _12370_ /*3981*/;
assign _12374_ = _12073_ ^ _12370_ /*3984*/;
assign _12375_ = _12366_ & _12374_ /*3982*/;
assign _12297_ = _12366_ ^ _12374_ /*3983*/;
assign _12372_ = _12373_ | _12375_ /*3980*/;
assign _12377_ = ~Q[4] /*3979*/;
assign _12376_ = _12377_ & D[9] /*3978*/;
assign _12379_ = _12074_ & _12376_ /*3973*/;
assign _12380_ = _12074_ ^ _12376_ /*3976*/;
assign _12381_ = _12372_ & _12380_ /*3974*/;
assign _12298_ = _12372_ ^ _12380_ /*3975*/;
assign _12378_ = _12379_ | _12381_ /*3972*/;
assign _12383_ = ~Q[4] /*3971*/;
assign _12382_ = _12383_ & D[10] /*3970*/;
assign _12385_ = _12075_ & _12382_ /*3965*/;
assign _12386_ = _12075_ ^ _12382_ /*3968*/;
assign _12387_ = _12378_ & _12386_ /*3966*/;
assign _12299_ = _12378_ ^ _12386_ /*3967*/;
assign _12384_ = _12385_ | _12387_ /*3964*/;
assign _12389_ = ~Q[4] /*3963*/;
assign _12388_ = _12389_ & D[11] /*3962*/;
assign _12391_ = _12076_ & _12388_ /*3957*/;
assign _12392_ = _12076_ ^ _12388_ /*3960*/;
assign _12393_ = _12384_ & _12392_ /*3958*/;
assign _12300_ = _12384_ ^ _12392_ /*3959*/;
assign _12390_ = _12391_ | _12393_ /*3956*/;
assign _12395_ = ~Q[4] /*3955*/;
assign _12394_ = _12395_ & D[12] /*3954*/;
assign _12397_ = _12077_ & _12394_ /*3949*/;
assign _12398_ = _12077_ ^ _12394_ /*3952*/;
assign _12399_ = _12390_ & _12398_ /*3950*/;
assign _12301_ = _12390_ ^ _12398_ /*3951*/;
assign _12396_ = _12397_ | _12399_ /*3948*/;
assign _12401_ = ~Q[4] /*3947*/;
assign _12400_ = _12401_ & D[13] /*3946*/;
assign _12403_ = _12078_ & _12400_ /*3941*/;
assign _12404_ = _12078_ ^ _12400_ /*3944*/;
assign _12405_ = _12396_ & _12404_ /*3942*/;
assign _12302_ = _12396_ ^ _12404_ /*3943*/;
assign _12402_ = _12403_ | _12405_ /*3940*/;
assign _12407_ = ~Q[4] /*3939*/;
assign _12406_ = _12407_ & D[14] /*3938*/;
assign _12409_ = _12079_ & _12406_ /*3933*/;
assign _12410_ = _12079_ ^ _12406_ /*3936*/;
assign _12411_ = _12402_ & _12410_ /*3934*/;
assign _12303_ = _12402_ ^ _12410_ /*3935*/;
assign _12408_ = _12409_ | _12411_ /*3932*/;
assign _12413_ = ~Q[4] /*3931*/;
assign _12412_ = _12413_ & D[15] /*3930*/;
assign _12415_ = _12080_ & _12412_ /*3925*/;
assign _12416_ = _12080_ ^ _12412_ /*3928*/;
assign _12417_ = _12408_ & _12416_ /*3926*/;
assign _12304_ = _12408_ ^ _12416_ /*3927*/;
assign _12414_ = _12415_ | _12417_ /*3924*/;
assign _12419_ = ~Q[4] /*3923*/;
assign _12418_ = _12419_ & D[16] /*3922*/;
assign _12421_ = _12081_ & _12418_ /*3917*/;
assign _12422_ = _12081_ ^ _12418_ /*3920*/;
assign _12423_ = _12414_ & _12422_ /*3918*/;
assign _12305_ = _12414_ ^ _12422_ /*3919*/;
assign _12420_ = _12421_ | _12423_ /*3916*/;
assign _12425_ = ~Q[4] /*3915*/;
assign _12424_ = _12425_ & D[17] /*3914*/;
assign _12427_ = _12082_ & _12424_ /*3909*/;
assign _12428_ = _12082_ ^ _12424_ /*3912*/;
assign _12429_ = _12420_ & _12428_ /*3910*/;
assign _12306_ = _12420_ ^ _12428_ /*3911*/;
assign _12426_ = _12427_ | _12429_ /*3908*/;
assign _12431_ = ~Q[4] /*3907*/;
assign _12430_ = _12431_ & D[18] /*3906*/;
assign _12433_ = _12083_ & _12430_ /*3901*/;
assign _12434_ = _12083_ ^ _12430_ /*3904*/;
assign _12435_ = _12426_ & _12434_ /*3902*/;
assign _12307_ = _12426_ ^ _12434_ /*3903*/;
assign _12432_ = _12433_ | _12435_ /*3900*/;
assign _12437_ = ~Q[4] /*3899*/;
assign _12436_ = _12437_ & D[19] /*3898*/;
assign _12439_ = _12084_ & _12436_ /*3893*/;
assign _12440_ = _12084_ ^ _12436_ /*3896*/;
assign _12441_ = _12432_ & _12440_ /*3894*/;
assign _12308_ = _12432_ ^ _12440_ /*3895*/;
assign _12438_ = _12439_ | _12441_ /*3892*/;
assign _12443_ = ~Q[4] /*3891*/;
assign _12442_ = _12443_ & D[20] /*3890*/;
assign _12445_ = _12085_ & _12442_ /*3885*/;
assign _12446_ = _12085_ ^ _12442_ /*3888*/;
assign _12447_ = _12438_ & _12446_ /*3886*/;
assign _12309_ = _12438_ ^ _12446_ /*3887*/;
assign _12444_ = _12445_ | _12447_ /*3884*/;
assign _12449_ = ~Q[4] /*3883*/;
assign _12448_ = _12449_ & D[21] /*3882*/;
assign _12451_ = _12086_ & _12448_ /*3877*/;
assign _12452_ = _12086_ ^ _12448_ /*3880*/;
assign _12453_ = _12444_ & _12452_ /*3878*/;
assign _12310_ = _12444_ ^ _12452_ /*3879*/;
assign _12450_ = _12451_ | _12453_ /*3876*/;
assign _12455_ = ~Q[4] /*3875*/;
assign _12454_ = _12455_ & D[22] /*3874*/;
assign _12457_ = _12087_ & _12454_ /*3869*/;
assign _12458_ = _12087_ ^ _12454_ /*3872*/;
assign _12459_ = _12450_ & _12458_ /*3870*/;
assign _12311_ = _12450_ ^ _12458_ /*3871*/;
assign _12456_ = _12457_ | _12459_ /*3868*/;
assign _12461_ = ~Q[4] /*3867*/;
assign _12460_ = _12461_ & D[23] /*3866*/;
assign _12463_ = _12088_ & _12460_ /*3861*/;
assign _12464_ = _12088_ ^ _12460_ /*3864*/;
assign _12465_ = _12456_ & _12464_ /*3862*/;
assign _12312_ = _12456_ ^ _12464_ /*3863*/;
assign _12462_ = _12463_ | _12465_ /*3860*/;
assign _12467_ = ~Q[4] /*3859*/;
assign _12466_ = _12467_ & D[24] /*3858*/;
assign _12469_ = _12089_ & _12466_ /*3853*/;
assign _12470_ = _12089_ ^ _12466_ /*3856*/;
assign _12471_ = _12462_ & _12470_ /*3854*/;
assign _12313_ = _12462_ ^ _12470_ /*3855*/;
assign _12468_ = _12469_ | _12471_ /*3852*/;
assign _12473_ = ~Q[4] /*3851*/;
assign _12472_ = _12473_ & D[25] /*3850*/;
assign _12475_ = _12090_ & _12472_ /*3845*/;
assign _12476_ = _12090_ ^ _12472_ /*3848*/;
assign _12477_ = _12468_ & _12476_ /*3846*/;
assign _12314_ = _12468_ ^ _12476_ /*3847*/;
assign _12474_ = _12475_ | _12477_ /*3844*/;
assign _12479_ = ~Q[4] /*3843*/;
assign _12478_ = _12479_ & D[26] /*3842*/;
assign _12481_ = _12091_ & _12478_ /*3837*/;
assign _12482_ = _12091_ ^ _12478_ /*3840*/;
assign _12483_ = _12474_ & _12482_ /*3838*/;
assign _12315_ = _12474_ ^ _12482_ /*3839*/;
assign _12480_ = _12481_ | _12483_ /*3836*/;
assign _12485_ = ~Q[4] /*3835*/;
assign _12484_ = _12485_ & D[27] /*3834*/;
assign _12487_ = _12092_ & _12484_ /*3829*/;
assign _12488_ = _12092_ ^ _12484_ /*3832*/;
assign _12489_ = _12480_ & _12488_ /*3830*/;
assign _12316_ = _12480_ ^ _12488_ /*3831*/;
assign _12486_ = _12487_ | _12489_ /*3828*/;
assign _12491_ = ~Q[4] /*3827*/;
assign _12490_ = _12491_ & D[28] /*3826*/;
assign _12493_ = _12093_ & _12490_ /*3821*/;
assign _12494_ = _12093_ ^ _12490_ /*3824*/;
assign _12495_ = _12486_ & _12494_ /*3822*/;
assign _12317_ = _12486_ ^ _12494_ /*3823*/;
assign _12492_ = _12493_ | _12495_ /*3820*/;
assign _12497_ = ~Q[4] /*3819*/;
assign _12496_ = _12497_ & D[29] /*3818*/;
assign _12499_ = _12094_ & _12496_ /*3813*/;
assign _12500_ = _12094_ ^ _12496_ /*3816*/;
assign _12501_ = _12492_ & _12500_ /*3814*/;
assign _12318_ = _12492_ ^ _12500_ /*3815*/;
assign _12498_ = _12499_ | _12501_ /*3812*/;
assign _12503_ = ~Q[4] /*3811*/;
assign _12502_ = _12503_ & D[30] /*3810*/;
assign _12505_ = _12095_ & _12502_ /*3805*/;
assign _12506_ = _12095_ ^ _12502_ /*3808*/;
assign _12507_ = _12498_ & _12506_ /*3806*/;
assign _12319_ = _12498_ ^ _12506_ /*3807*/;
assign _12504_ = _12505_ | _12507_ /*3804*/;
assign _12509_ = ~Q[4] /*3803*/;
assign _12508_ = _12509_ & zeroWire /*3802*/;
assign _12510_ = _12096_ ^ _12508_ /*3800*/;
assign _12320_ = _12510_ ^ _12504_ /*3799*/;
assign _12549_ = ~D[0] /*3673*/;
assign _12546_ = R_0[3] & _12549_ /*3669*/;
assign _12547_ = R_0[3] ^ _12549_ /*3672*/;
assign _12548_ = oneWire & _12547_ /*3670*/;
assign _12513_ = oneWire ^ _12547_ /*3671*/;
assign _12545_ = _12546_ | _12548_ /*3668*/;
assign _12554_ = ~D[1] /*3667*/;
assign _12551_ = _12289_ & _12554_ /*3663*/;
assign _12552_ = _12289_ ^ _12554_ /*3666*/;
assign _12553_ = _12545_ & _12552_ /*3664*/;
assign _12514_ = _12545_ ^ _12552_ /*3665*/;
assign _12550_ = _12551_ | _12553_ /*3662*/;
assign _12559_ = ~D[2] /*3661*/;
assign _12556_ = _12290_ & _12559_ /*3657*/;
assign _12557_ = _12290_ ^ _12559_ /*3660*/;
assign _12558_ = _12550_ & _12557_ /*3658*/;
assign _12515_ = _12550_ ^ _12557_ /*3659*/;
assign _12555_ = _12556_ | _12558_ /*3656*/;
assign _12564_ = ~D[3] /*3655*/;
assign _12561_ = _12291_ & _12564_ /*3651*/;
assign _12562_ = _12291_ ^ _12564_ /*3654*/;
assign _12563_ = _12555_ & _12562_ /*3652*/;
assign _12516_ = _12555_ ^ _12562_ /*3653*/;
assign _12560_ = _12561_ | _12563_ /*3650*/;
assign _12569_ = ~D[4] /*3649*/;
assign _12566_ = _12292_ & _12569_ /*3645*/;
assign _12567_ = _12292_ ^ _12569_ /*3648*/;
assign _12568_ = _12560_ & _12567_ /*3646*/;
assign _12517_ = _12560_ ^ _12567_ /*3647*/;
assign _12565_ = _12566_ | _12568_ /*3644*/;
assign _12574_ = ~D[5] /*3643*/;
assign _12571_ = _12293_ & _12574_ /*3639*/;
assign _12572_ = _12293_ ^ _12574_ /*3642*/;
assign _12573_ = _12565_ & _12572_ /*3640*/;
assign _12518_ = _12565_ ^ _12572_ /*3641*/;
assign _12570_ = _12571_ | _12573_ /*3638*/;
assign _12579_ = ~D[6] /*3637*/;
assign _12576_ = _12294_ & _12579_ /*3633*/;
assign _12577_ = _12294_ ^ _12579_ /*3636*/;
assign _12578_ = _12570_ & _12577_ /*3634*/;
assign _12519_ = _12570_ ^ _12577_ /*3635*/;
assign _12575_ = _12576_ | _12578_ /*3632*/;
assign _12584_ = ~D[7] /*3631*/;
assign _12581_ = _12295_ & _12584_ /*3627*/;
assign _12582_ = _12295_ ^ _12584_ /*3630*/;
assign _12583_ = _12575_ & _12582_ /*3628*/;
assign _12520_ = _12575_ ^ _12582_ /*3629*/;
assign _12580_ = _12581_ | _12583_ /*3626*/;
assign _12589_ = ~D[8] /*3625*/;
assign _12586_ = _12296_ & _12589_ /*3621*/;
assign _12587_ = _12296_ ^ _12589_ /*3624*/;
assign _12588_ = _12580_ & _12587_ /*3622*/;
assign _12521_ = _12580_ ^ _12587_ /*3623*/;
assign _12585_ = _12586_ | _12588_ /*3620*/;
assign _12594_ = ~D[9] /*3619*/;
assign _12591_ = _12297_ & _12594_ /*3615*/;
assign _12592_ = _12297_ ^ _12594_ /*3618*/;
assign _12593_ = _12585_ & _12592_ /*3616*/;
assign _12522_ = _12585_ ^ _12592_ /*3617*/;
assign _12590_ = _12591_ | _12593_ /*3614*/;
assign _12599_ = ~D[10] /*3613*/;
assign _12596_ = _12298_ & _12599_ /*3609*/;
assign _12597_ = _12298_ ^ _12599_ /*3612*/;
assign _12598_ = _12590_ & _12597_ /*3610*/;
assign _12523_ = _12590_ ^ _12597_ /*3611*/;
assign _12595_ = _12596_ | _12598_ /*3608*/;
assign _12604_ = ~D[11] /*3607*/;
assign _12601_ = _12299_ & _12604_ /*3603*/;
assign _12602_ = _12299_ ^ _12604_ /*3606*/;
assign _12603_ = _12595_ & _12602_ /*3604*/;
assign _12524_ = _12595_ ^ _12602_ /*3605*/;
assign _12600_ = _12601_ | _12603_ /*3602*/;
assign _12609_ = ~D[12] /*3601*/;
assign _12606_ = _12300_ & _12609_ /*3597*/;
assign _12607_ = _12300_ ^ _12609_ /*3600*/;
assign _12608_ = _12600_ & _12607_ /*3598*/;
assign _12525_ = _12600_ ^ _12607_ /*3599*/;
assign _12605_ = _12606_ | _12608_ /*3596*/;
assign _12614_ = ~D[13] /*3595*/;
assign _12611_ = _12301_ & _12614_ /*3591*/;
assign _12612_ = _12301_ ^ _12614_ /*3594*/;
assign _12613_ = _12605_ & _12612_ /*3592*/;
assign _12526_ = _12605_ ^ _12612_ /*3593*/;
assign _12610_ = _12611_ | _12613_ /*3590*/;
assign _12619_ = ~D[14] /*3589*/;
assign _12616_ = _12302_ & _12619_ /*3585*/;
assign _12617_ = _12302_ ^ _12619_ /*3588*/;
assign _12618_ = _12610_ & _12617_ /*3586*/;
assign _12527_ = _12610_ ^ _12617_ /*3587*/;
assign _12615_ = _12616_ | _12618_ /*3584*/;
assign _12624_ = ~D[15] /*3583*/;
assign _12621_ = _12303_ & _12624_ /*3579*/;
assign _12622_ = _12303_ ^ _12624_ /*3582*/;
assign _12623_ = _12615_ & _12622_ /*3580*/;
assign _12528_ = _12615_ ^ _12622_ /*3581*/;
assign _12620_ = _12621_ | _12623_ /*3578*/;
assign _12629_ = ~D[16] /*3577*/;
assign _12626_ = _12304_ & _12629_ /*3573*/;
assign _12627_ = _12304_ ^ _12629_ /*3576*/;
assign _12628_ = _12620_ & _12627_ /*3574*/;
assign _12529_ = _12620_ ^ _12627_ /*3575*/;
assign _12625_ = _12626_ | _12628_ /*3572*/;
assign _12634_ = ~D[17] /*3571*/;
assign _12631_ = _12305_ & _12634_ /*3567*/;
assign _12632_ = _12305_ ^ _12634_ /*3570*/;
assign _12633_ = _12625_ & _12632_ /*3568*/;
assign _12530_ = _12625_ ^ _12632_ /*3569*/;
assign _12630_ = _12631_ | _12633_ /*3566*/;
assign _12639_ = ~D[18] /*3565*/;
assign _12636_ = _12306_ & _12639_ /*3561*/;
assign _12637_ = _12306_ ^ _12639_ /*3564*/;
assign _12638_ = _12630_ & _12637_ /*3562*/;
assign _12531_ = _12630_ ^ _12637_ /*3563*/;
assign _12635_ = _12636_ | _12638_ /*3560*/;
assign _12644_ = ~D[19] /*3559*/;
assign _12641_ = _12307_ & _12644_ /*3555*/;
assign _12642_ = _12307_ ^ _12644_ /*3558*/;
assign _12643_ = _12635_ & _12642_ /*3556*/;
assign _12532_ = _12635_ ^ _12642_ /*3557*/;
assign _12640_ = _12641_ | _12643_ /*3554*/;
assign _12649_ = ~D[20] /*3553*/;
assign _12646_ = _12308_ & _12649_ /*3549*/;
assign _12647_ = _12308_ ^ _12649_ /*3552*/;
assign _12648_ = _12640_ & _12647_ /*3550*/;
assign _12533_ = _12640_ ^ _12647_ /*3551*/;
assign _12645_ = _12646_ | _12648_ /*3548*/;
assign _12654_ = ~D[21] /*3547*/;
assign _12651_ = _12309_ & _12654_ /*3543*/;
assign _12652_ = _12309_ ^ _12654_ /*3546*/;
assign _12653_ = _12645_ & _12652_ /*3544*/;
assign _12534_ = _12645_ ^ _12652_ /*3545*/;
assign _12650_ = _12651_ | _12653_ /*3542*/;
assign _12659_ = ~D[22] /*3541*/;
assign _12656_ = _12310_ & _12659_ /*3537*/;
assign _12657_ = _12310_ ^ _12659_ /*3540*/;
assign _12658_ = _12650_ & _12657_ /*3538*/;
assign _12535_ = _12650_ ^ _12657_ /*3539*/;
assign _12655_ = _12656_ | _12658_ /*3536*/;
assign _12664_ = ~D[23] /*3535*/;
assign _12661_ = _12311_ & _12664_ /*3531*/;
assign _12662_ = _12311_ ^ _12664_ /*3534*/;
assign _12663_ = _12655_ & _12662_ /*3532*/;
assign _12536_ = _12655_ ^ _12662_ /*3533*/;
assign _12660_ = _12661_ | _12663_ /*3530*/;
assign _12669_ = ~D[24] /*3529*/;
assign _12666_ = _12312_ & _12669_ /*3525*/;
assign _12667_ = _12312_ ^ _12669_ /*3528*/;
assign _12668_ = _12660_ & _12667_ /*3526*/;
assign _12537_ = _12660_ ^ _12667_ /*3527*/;
assign _12665_ = _12666_ | _12668_ /*3524*/;
assign _12674_ = ~D[25] /*3523*/;
assign _12671_ = _12313_ & _12674_ /*3519*/;
assign _12672_ = _12313_ ^ _12674_ /*3522*/;
assign _12673_ = _12665_ & _12672_ /*3520*/;
assign _12538_ = _12665_ ^ _12672_ /*3521*/;
assign _12670_ = _12671_ | _12673_ /*3518*/;
assign _12679_ = ~D[26] /*3517*/;
assign _12676_ = _12314_ & _12679_ /*3513*/;
assign _12677_ = _12314_ ^ _12679_ /*3516*/;
assign _12678_ = _12670_ & _12677_ /*3514*/;
assign _12539_ = _12670_ ^ _12677_ /*3515*/;
assign _12675_ = _12676_ | _12678_ /*3512*/;
assign _12684_ = ~D[27] /*3511*/;
assign _12681_ = _12315_ & _12684_ /*3507*/;
assign _12682_ = _12315_ ^ _12684_ /*3510*/;
assign _12683_ = _12675_ & _12682_ /*3508*/;
assign _12540_ = _12675_ ^ _12682_ /*3509*/;
assign _12680_ = _12681_ | _12683_ /*3506*/;
assign _12689_ = ~D[28] /*3505*/;
assign _12686_ = _12316_ & _12689_ /*3501*/;
assign _12687_ = _12316_ ^ _12689_ /*3504*/;
assign _12688_ = _12680_ & _12687_ /*3502*/;
assign _12541_ = _12680_ ^ _12687_ /*3503*/;
assign _12685_ = _12686_ | _12688_ /*3500*/;
assign _12694_ = ~D[29] /*3499*/;
assign _12691_ = _12317_ & _12694_ /*3495*/;
assign _12692_ = _12317_ ^ _12694_ /*3498*/;
assign _12693_ = _12685_ & _12692_ /*3496*/;
assign _12542_ = _12685_ ^ _12692_ /*3497*/;
assign _12690_ = _12691_ | _12693_ /*3494*/;
assign _12699_ = ~D[30] /*3493*/;
assign _12696_ = _12318_ & _12699_ /*3489*/;
assign _12697_ = _12318_ ^ _12699_ /*3492*/;
assign _12698_ = _12690_ & _12697_ /*3490*/;
assign _12543_ = _12690_ ^ _12697_ /*3491*/;
assign _12695_ = _12696_ | _12698_ /*3488*/;
assign _12700_ = _12319_ & oneWire /*3483*/;
assign _12701_ = _12319_ ^ oneWire /*3486*/;
assign _12702_ = _12695_ & _12701_ /*3484*/;
assign _12544_ = _12695_ ^ _12701_ /*3485*/;
assign Q[3] = _12700_ | _12702_ /*3482*/;
assign _12771_ = ~Q[3] /*3289*/;
assign _12770_ = _12771_ & D[0] /*3288*/;
assign _12773_ = _12513_ & _12770_ /*3283*/;
assign _12774_ = _12513_ ^ _12770_ /*3286*/;
assign _12775_ = zeroWire & _12774_ /*3284*/;
assign _12737_ = zeroWire ^ _12774_ /*3285*/;
assign _12772_ = _12773_ | _12775_ /*3282*/;
assign _12777_ = ~Q[3] /*3281*/;
assign _12776_ = _12777_ & D[1] /*3280*/;
assign _12779_ = _12514_ & _12776_ /*3275*/;
assign _12780_ = _12514_ ^ _12776_ /*3278*/;
assign _12781_ = _12772_ & _12780_ /*3276*/;
assign _12738_ = _12772_ ^ _12780_ /*3277*/;
assign _12778_ = _12779_ | _12781_ /*3274*/;
assign _12783_ = ~Q[3] /*3273*/;
assign _12782_ = _12783_ & D[2] /*3272*/;
assign _12785_ = _12515_ & _12782_ /*3267*/;
assign _12786_ = _12515_ ^ _12782_ /*3270*/;
assign _12787_ = _12778_ & _12786_ /*3268*/;
assign _12739_ = _12778_ ^ _12786_ /*3269*/;
assign _12784_ = _12785_ | _12787_ /*3266*/;
assign _12789_ = ~Q[3] /*3265*/;
assign _12788_ = _12789_ & D[3] /*3264*/;
assign _12791_ = _12516_ & _12788_ /*3259*/;
assign _12792_ = _12516_ ^ _12788_ /*3262*/;
assign _12793_ = _12784_ & _12792_ /*3260*/;
assign _12740_ = _12784_ ^ _12792_ /*3261*/;
assign _12790_ = _12791_ | _12793_ /*3258*/;
assign _12795_ = ~Q[3] /*3257*/;
assign _12794_ = _12795_ & D[4] /*3256*/;
assign _12797_ = _12517_ & _12794_ /*3251*/;
assign _12798_ = _12517_ ^ _12794_ /*3254*/;
assign _12799_ = _12790_ & _12798_ /*3252*/;
assign _12741_ = _12790_ ^ _12798_ /*3253*/;
assign _12796_ = _12797_ | _12799_ /*3250*/;
assign _12801_ = ~Q[3] /*3249*/;
assign _12800_ = _12801_ & D[5] /*3248*/;
assign _12803_ = _12518_ & _12800_ /*3243*/;
assign _12804_ = _12518_ ^ _12800_ /*3246*/;
assign _12805_ = _12796_ & _12804_ /*3244*/;
assign _12742_ = _12796_ ^ _12804_ /*3245*/;
assign _12802_ = _12803_ | _12805_ /*3242*/;
assign _12807_ = ~Q[3] /*3241*/;
assign _12806_ = _12807_ & D[6] /*3240*/;
assign _12809_ = _12519_ & _12806_ /*3235*/;
assign _12810_ = _12519_ ^ _12806_ /*3238*/;
assign _12811_ = _12802_ & _12810_ /*3236*/;
assign _12743_ = _12802_ ^ _12810_ /*3237*/;
assign _12808_ = _12809_ | _12811_ /*3234*/;
assign _12813_ = ~Q[3] /*3233*/;
assign _12812_ = _12813_ & D[7] /*3232*/;
assign _12815_ = _12520_ & _12812_ /*3227*/;
assign _12816_ = _12520_ ^ _12812_ /*3230*/;
assign _12817_ = _12808_ & _12816_ /*3228*/;
assign _12744_ = _12808_ ^ _12816_ /*3229*/;
assign _12814_ = _12815_ | _12817_ /*3226*/;
assign _12819_ = ~Q[3] /*3225*/;
assign _12818_ = _12819_ & D[8] /*3224*/;
assign _12821_ = _12521_ & _12818_ /*3219*/;
assign _12822_ = _12521_ ^ _12818_ /*3222*/;
assign _12823_ = _12814_ & _12822_ /*3220*/;
assign _12745_ = _12814_ ^ _12822_ /*3221*/;
assign _12820_ = _12821_ | _12823_ /*3218*/;
assign _12825_ = ~Q[3] /*3217*/;
assign _12824_ = _12825_ & D[9] /*3216*/;
assign _12827_ = _12522_ & _12824_ /*3211*/;
assign _12828_ = _12522_ ^ _12824_ /*3214*/;
assign _12829_ = _12820_ & _12828_ /*3212*/;
assign _12746_ = _12820_ ^ _12828_ /*3213*/;
assign _12826_ = _12827_ | _12829_ /*3210*/;
assign _12831_ = ~Q[3] /*3209*/;
assign _12830_ = _12831_ & D[10] /*3208*/;
assign _12833_ = _12523_ & _12830_ /*3203*/;
assign _12834_ = _12523_ ^ _12830_ /*3206*/;
assign _12835_ = _12826_ & _12834_ /*3204*/;
assign _12747_ = _12826_ ^ _12834_ /*3205*/;
assign _12832_ = _12833_ | _12835_ /*3202*/;
assign _12837_ = ~Q[3] /*3201*/;
assign _12836_ = _12837_ & D[11] /*3200*/;
assign _12839_ = _12524_ & _12836_ /*3195*/;
assign _12840_ = _12524_ ^ _12836_ /*3198*/;
assign _12841_ = _12832_ & _12840_ /*3196*/;
assign _12748_ = _12832_ ^ _12840_ /*3197*/;
assign _12838_ = _12839_ | _12841_ /*3194*/;
assign _12843_ = ~Q[3] /*3193*/;
assign _12842_ = _12843_ & D[12] /*3192*/;
assign _12845_ = _12525_ & _12842_ /*3187*/;
assign _12846_ = _12525_ ^ _12842_ /*3190*/;
assign _12847_ = _12838_ & _12846_ /*3188*/;
assign _12749_ = _12838_ ^ _12846_ /*3189*/;
assign _12844_ = _12845_ | _12847_ /*3186*/;
assign _12849_ = ~Q[3] /*3185*/;
assign _12848_ = _12849_ & D[13] /*3184*/;
assign _12851_ = _12526_ & _12848_ /*3179*/;
assign _12852_ = _12526_ ^ _12848_ /*3182*/;
assign _12853_ = _12844_ & _12852_ /*3180*/;
assign _12750_ = _12844_ ^ _12852_ /*3181*/;
assign _12850_ = _12851_ | _12853_ /*3178*/;
assign _12855_ = ~Q[3] /*3177*/;
assign _12854_ = _12855_ & D[14] /*3176*/;
assign _12857_ = _12527_ & _12854_ /*3171*/;
assign _12858_ = _12527_ ^ _12854_ /*3174*/;
assign _12859_ = _12850_ & _12858_ /*3172*/;
assign _12751_ = _12850_ ^ _12858_ /*3173*/;
assign _12856_ = _12857_ | _12859_ /*3170*/;
assign _12861_ = ~Q[3] /*3169*/;
assign _12860_ = _12861_ & D[15] /*3168*/;
assign _12863_ = _12528_ & _12860_ /*3163*/;
assign _12864_ = _12528_ ^ _12860_ /*3166*/;
assign _12865_ = _12856_ & _12864_ /*3164*/;
assign _12752_ = _12856_ ^ _12864_ /*3165*/;
assign _12862_ = _12863_ | _12865_ /*3162*/;
assign _12867_ = ~Q[3] /*3161*/;
assign _12866_ = _12867_ & D[16] /*3160*/;
assign _12869_ = _12529_ & _12866_ /*3155*/;
assign _12870_ = _12529_ ^ _12866_ /*3158*/;
assign _12871_ = _12862_ & _12870_ /*3156*/;
assign _12753_ = _12862_ ^ _12870_ /*3157*/;
assign _12868_ = _12869_ | _12871_ /*3154*/;
assign _12873_ = ~Q[3] /*3153*/;
assign _12872_ = _12873_ & D[17] /*3152*/;
assign _12875_ = _12530_ & _12872_ /*3147*/;
assign _12876_ = _12530_ ^ _12872_ /*3150*/;
assign _12877_ = _12868_ & _12876_ /*3148*/;
assign _12754_ = _12868_ ^ _12876_ /*3149*/;
assign _12874_ = _12875_ | _12877_ /*3146*/;
assign _12879_ = ~Q[3] /*3145*/;
assign _12878_ = _12879_ & D[18] /*3144*/;
assign _12881_ = _12531_ & _12878_ /*3139*/;
assign _12882_ = _12531_ ^ _12878_ /*3142*/;
assign _12883_ = _12874_ & _12882_ /*3140*/;
assign _12755_ = _12874_ ^ _12882_ /*3141*/;
assign _12880_ = _12881_ | _12883_ /*3138*/;
assign _12885_ = ~Q[3] /*3137*/;
assign _12884_ = _12885_ & D[19] /*3136*/;
assign _12887_ = _12532_ & _12884_ /*3131*/;
assign _12888_ = _12532_ ^ _12884_ /*3134*/;
assign _12889_ = _12880_ & _12888_ /*3132*/;
assign _12756_ = _12880_ ^ _12888_ /*3133*/;
assign _12886_ = _12887_ | _12889_ /*3130*/;
assign _12891_ = ~Q[3] /*3129*/;
assign _12890_ = _12891_ & D[20] /*3128*/;
assign _12893_ = _12533_ & _12890_ /*3123*/;
assign _12894_ = _12533_ ^ _12890_ /*3126*/;
assign _12895_ = _12886_ & _12894_ /*3124*/;
assign _12757_ = _12886_ ^ _12894_ /*3125*/;
assign _12892_ = _12893_ | _12895_ /*3122*/;
assign _12897_ = ~Q[3] /*3121*/;
assign _12896_ = _12897_ & D[21] /*3120*/;
assign _12899_ = _12534_ & _12896_ /*3115*/;
assign _12900_ = _12534_ ^ _12896_ /*3118*/;
assign _12901_ = _12892_ & _12900_ /*3116*/;
assign _12758_ = _12892_ ^ _12900_ /*3117*/;
assign _12898_ = _12899_ | _12901_ /*3114*/;
assign _12903_ = ~Q[3] /*3113*/;
assign _12902_ = _12903_ & D[22] /*3112*/;
assign _12905_ = _12535_ & _12902_ /*3107*/;
assign _12906_ = _12535_ ^ _12902_ /*3110*/;
assign _12907_ = _12898_ & _12906_ /*3108*/;
assign _12759_ = _12898_ ^ _12906_ /*3109*/;
assign _12904_ = _12905_ | _12907_ /*3106*/;
assign _12909_ = ~Q[3] /*3105*/;
assign _12908_ = _12909_ & D[23] /*3104*/;
assign _12911_ = _12536_ & _12908_ /*3099*/;
assign _12912_ = _12536_ ^ _12908_ /*3102*/;
assign _12913_ = _12904_ & _12912_ /*3100*/;
assign _12760_ = _12904_ ^ _12912_ /*3101*/;
assign _12910_ = _12911_ | _12913_ /*3098*/;
assign _12915_ = ~Q[3] /*3097*/;
assign _12914_ = _12915_ & D[24] /*3096*/;
assign _12917_ = _12537_ & _12914_ /*3091*/;
assign _12918_ = _12537_ ^ _12914_ /*3094*/;
assign _12919_ = _12910_ & _12918_ /*3092*/;
assign _12761_ = _12910_ ^ _12918_ /*3093*/;
assign _12916_ = _12917_ | _12919_ /*3090*/;
assign _12921_ = ~Q[3] /*3089*/;
assign _12920_ = _12921_ & D[25] /*3088*/;
assign _12923_ = _12538_ & _12920_ /*3083*/;
assign _12924_ = _12538_ ^ _12920_ /*3086*/;
assign _12925_ = _12916_ & _12924_ /*3084*/;
assign _12762_ = _12916_ ^ _12924_ /*3085*/;
assign _12922_ = _12923_ | _12925_ /*3082*/;
assign _12927_ = ~Q[3] /*3081*/;
assign _12926_ = _12927_ & D[26] /*3080*/;
assign _12929_ = _12539_ & _12926_ /*3075*/;
assign _12930_ = _12539_ ^ _12926_ /*3078*/;
assign _12931_ = _12922_ & _12930_ /*3076*/;
assign _12763_ = _12922_ ^ _12930_ /*3077*/;
assign _12928_ = _12929_ | _12931_ /*3074*/;
assign _12933_ = ~Q[3] /*3073*/;
assign _12932_ = _12933_ & D[27] /*3072*/;
assign _12935_ = _12540_ & _12932_ /*3067*/;
assign _12936_ = _12540_ ^ _12932_ /*3070*/;
assign _12937_ = _12928_ & _12936_ /*3068*/;
assign _12764_ = _12928_ ^ _12936_ /*3069*/;
assign _12934_ = _12935_ | _12937_ /*3066*/;
assign _12939_ = ~Q[3] /*3065*/;
assign _12938_ = _12939_ & D[28] /*3064*/;
assign _12941_ = _12541_ & _12938_ /*3059*/;
assign _12942_ = _12541_ ^ _12938_ /*3062*/;
assign _12943_ = _12934_ & _12942_ /*3060*/;
assign _12765_ = _12934_ ^ _12942_ /*3061*/;
assign _12940_ = _12941_ | _12943_ /*3058*/;
assign _12945_ = ~Q[3] /*3057*/;
assign _12944_ = _12945_ & D[29] /*3056*/;
assign _12947_ = _12542_ & _12944_ /*3051*/;
assign _12948_ = _12542_ ^ _12944_ /*3054*/;
assign _12949_ = _12940_ & _12948_ /*3052*/;
assign _12766_ = _12940_ ^ _12948_ /*3053*/;
assign _12946_ = _12947_ | _12949_ /*3050*/;
assign _12951_ = ~Q[3] /*3049*/;
assign _12950_ = _12951_ & D[30] /*3048*/;
assign _12953_ = _12543_ & _12950_ /*3043*/;
assign _12954_ = _12543_ ^ _12950_ /*3046*/;
assign _12955_ = _12946_ & _12954_ /*3044*/;
assign _12767_ = _12946_ ^ _12954_ /*3045*/;
assign _12952_ = _12953_ | _12955_ /*3042*/;
assign _12957_ = ~Q[3] /*3041*/;
assign _12956_ = _12957_ & zeroWire /*3040*/;
assign _12958_ = _12544_ ^ _12956_ /*3038*/;
assign _12768_ = _12958_ ^ _12952_ /*3037*/;
assign _12997_ = ~D[0] /*2911*/;
assign _12994_ = R_0[2] & _12997_ /*2907*/;
assign _12995_ = R_0[2] ^ _12997_ /*2910*/;
assign _12996_ = oneWire & _12995_ /*2908*/;
assign _12961_ = oneWire ^ _12995_ /*2909*/;
assign _12993_ = _12994_ | _12996_ /*2906*/;
assign _13002_ = ~D[1] /*2905*/;
assign _12999_ = _12737_ & _13002_ /*2901*/;
assign _13000_ = _12737_ ^ _13002_ /*2904*/;
assign _13001_ = _12993_ & _13000_ /*2902*/;
assign _12962_ = _12993_ ^ _13000_ /*2903*/;
assign _12998_ = _12999_ | _13001_ /*2900*/;
assign _13007_ = ~D[2] /*2899*/;
assign _13004_ = _12738_ & _13007_ /*2895*/;
assign _13005_ = _12738_ ^ _13007_ /*2898*/;
assign _13006_ = _12998_ & _13005_ /*2896*/;
assign _12963_ = _12998_ ^ _13005_ /*2897*/;
assign _13003_ = _13004_ | _13006_ /*2894*/;
assign _13012_ = ~D[3] /*2893*/;
assign _13009_ = _12739_ & _13012_ /*2889*/;
assign _13010_ = _12739_ ^ _13012_ /*2892*/;
assign _13011_ = _13003_ & _13010_ /*2890*/;
assign _12964_ = _13003_ ^ _13010_ /*2891*/;
assign _13008_ = _13009_ | _13011_ /*2888*/;
assign _13017_ = ~D[4] /*2887*/;
assign _13014_ = _12740_ & _13017_ /*2883*/;
assign _13015_ = _12740_ ^ _13017_ /*2886*/;
assign _13016_ = _13008_ & _13015_ /*2884*/;
assign _12965_ = _13008_ ^ _13015_ /*2885*/;
assign _13013_ = _13014_ | _13016_ /*2882*/;
assign _13022_ = ~D[5] /*2881*/;
assign _13019_ = _12741_ & _13022_ /*2877*/;
assign _13020_ = _12741_ ^ _13022_ /*2880*/;
assign _13021_ = _13013_ & _13020_ /*2878*/;
assign _12966_ = _13013_ ^ _13020_ /*2879*/;
assign _13018_ = _13019_ | _13021_ /*2876*/;
assign _13027_ = ~D[6] /*2875*/;
assign _13024_ = _12742_ & _13027_ /*2871*/;
assign _13025_ = _12742_ ^ _13027_ /*2874*/;
assign _13026_ = _13018_ & _13025_ /*2872*/;
assign _12967_ = _13018_ ^ _13025_ /*2873*/;
assign _13023_ = _13024_ | _13026_ /*2870*/;
assign _13032_ = ~D[7] /*2869*/;
assign _13029_ = _12743_ & _13032_ /*2865*/;
assign _13030_ = _12743_ ^ _13032_ /*2868*/;
assign _13031_ = _13023_ & _13030_ /*2866*/;
assign _12968_ = _13023_ ^ _13030_ /*2867*/;
assign _13028_ = _13029_ | _13031_ /*2864*/;
assign _13037_ = ~D[8] /*2863*/;
assign _13034_ = _12744_ & _13037_ /*2859*/;
assign _13035_ = _12744_ ^ _13037_ /*2862*/;
assign _13036_ = _13028_ & _13035_ /*2860*/;
assign _12969_ = _13028_ ^ _13035_ /*2861*/;
assign _13033_ = _13034_ | _13036_ /*2858*/;
assign _13042_ = ~D[9] /*2857*/;
assign _13039_ = _12745_ & _13042_ /*2853*/;
assign _13040_ = _12745_ ^ _13042_ /*2856*/;
assign _13041_ = _13033_ & _13040_ /*2854*/;
assign _12970_ = _13033_ ^ _13040_ /*2855*/;
assign _13038_ = _13039_ | _13041_ /*2852*/;
assign _13047_ = ~D[10] /*2851*/;
assign _13044_ = _12746_ & _13047_ /*2847*/;
assign _13045_ = _12746_ ^ _13047_ /*2850*/;
assign _13046_ = _13038_ & _13045_ /*2848*/;
assign _12971_ = _13038_ ^ _13045_ /*2849*/;
assign _13043_ = _13044_ | _13046_ /*2846*/;
assign _13052_ = ~D[11] /*2845*/;
assign _13049_ = _12747_ & _13052_ /*2841*/;
assign _13050_ = _12747_ ^ _13052_ /*2844*/;
assign _13051_ = _13043_ & _13050_ /*2842*/;
assign _12972_ = _13043_ ^ _13050_ /*2843*/;
assign _13048_ = _13049_ | _13051_ /*2840*/;
assign _13057_ = ~D[12] /*2839*/;
assign _13054_ = _12748_ & _13057_ /*2835*/;
assign _13055_ = _12748_ ^ _13057_ /*2838*/;
assign _13056_ = _13048_ & _13055_ /*2836*/;
assign _12973_ = _13048_ ^ _13055_ /*2837*/;
assign _13053_ = _13054_ | _13056_ /*2834*/;
assign _13062_ = ~D[13] /*2833*/;
assign _13059_ = _12749_ & _13062_ /*2829*/;
assign _13060_ = _12749_ ^ _13062_ /*2832*/;
assign _13061_ = _13053_ & _13060_ /*2830*/;
assign _12974_ = _13053_ ^ _13060_ /*2831*/;
assign _13058_ = _13059_ | _13061_ /*2828*/;
assign _13067_ = ~D[14] /*2827*/;
assign _13064_ = _12750_ & _13067_ /*2823*/;
assign _13065_ = _12750_ ^ _13067_ /*2826*/;
assign _13066_ = _13058_ & _13065_ /*2824*/;
assign _12975_ = _13058_ ^ _13065_ /*2825*/;
assign _13063_ = _13064_ | _13066_ /*2822*/;
assign _13072_ = ~D[15] /*2821*/;
assign _13069_ = _12751_ & _13072_ /*2817*/;
assign _13070_ = _12751_ ^ _13072_ /*2820*/;
assign _13071_ = _13063_ & _13070_ /*2818*/;
assign _12976_ = _13063_ ^ _13070_ /*2819*/;
assign _13068_ = _13069_ | _13071_ /*2816*/;
assign _13077_ = ~D[16] /*2815*/;
assign _13074_ = _12752_ & _13077_ /*2811*/;
assign _13075_ = _12752_ ^ _13077_ /*2814*/;
assign _13076_ = _13068_ & _13075_ /*2812*/;
assign _12977_ = _13068_ ^ _13075_ /*2813*/;
assign _13073_ = _13074_ | _13076_ /*2810*/;
assign _13082_ = ~D[17] /*2809*/;
assign _13079_ = _12753_ & _13082_ /*2805*/;
assign _13080_ = _12753_ ^ _13082_ /*2808*/;
assign _13081_ = _13073_ & _13080_ /*2806*/;
assign _12978_ = _13073_ ^ _13080_ /*2807*/;
assign _13078_ = _13079_ | _13081_ /*2804*/;
assign _13087_ = ~D[18] /*2803*/;
assign _13084_ = _12754_ & _13087_ /*2799*/;
assign _13085_ = _12754_ ^ _13087_ /*2802*/;
assign _13086_ = _13078_ & _13085_ /*2800*/;
assign _12979_ = _13078_ ^ _13085_ /*2801*/;
assign _13083_ = _13084_ | _13086_ /*2798*/;
assign _13092_ = ~D[19] /*2797*/;
assign _13089_ = _12755_ & _13092_ /*2793*/;
assign _13090_ = _12755_ ^ _13092_ /*2796*/;
assign _13091_ = _13083_ & _13090_ /*2794*/;
assign _12980_ = _13083_ ^ _13090_ /*2795*/;
assign _13088_ = _13089_ | _13091_ /*2792*/;
assign _13097_ = ~D[20] /*2791*/;
assign _13094_ = _12756_ & _13097_ /*2787*/;
assign _13095_ = _12756_ ^ _13097_ /*2790*/;
assign _13096_ = _13088_ & _13095_ /*2788*/;
assign _12981_ = _13088_ ^ _13095_ /*2789*/;
assign _13093_ = _13094_ | _13096_ /*2786*/;
assign _13102_ = ~D[21] /*2785*/;
assign _13099_ = _12757_ & _13102_ /*2781*/;
assign _13100_ = _12757_ ^ _13102_ /*2784*/;
assign _13101_ = _13093_ & _13100_ /*2782*/;
assign _12982_ = _13093_ ^ _13100_ /*2783*/;
assign _13098_ = _13099_ | _13101_ /*2780*/;
assign _13107_ = ~D[22] /*2779*/;
assign _13104_ = _12758_ & _13107_ /*2775*/;
assign _13105_ = _12758_ ^ _13107_ /*2778*/;
assign _13106_ = _13098_ & _13105_ /*2776*/;
assign _12983_ = _13098_ ^ _13105_ /*2777*/;
assign _13103_ = _13104_ | _13106_ /*2774*/;
assign _13112_ = ~D[23] /*2773*/;
assign _13109_ = _12759_ & _13112_ /*2769*/;
assign _13110_ = _12759_ ^ _13112_ /*2772*/;
assign _13111_ = _13103_ & _13110_ /*2770*/;
assign _12984_ = _13103_ ^ _13110_ /*2771*/;
assign _13108_ = _13109_ | _13111_ /*2768*/;
assign _13117_ = ~D[24] /*2767*/;
assign _13114_ = _12760_ & _13117_ /*2763*/;
assign _13115_ = _12760_ ^ _13117_ /*2766*/;
assign _13116_ = _13108_ & _13115_ /*2764*/;
assign _12985_ = _13108_ ^ _13115_ /*2765*/;
assign _13113_ = _13114_ | _13116_ /*2762*/;
assign _13122_ = ~D[25] /*2761*/;
assign _13119_ = _12761_ & _13122_ /*2757*/;
assign _13120_ = _12761_ ^ _13122_ /*2760*/;
assign _13121_ = _13113_ & _13120_ /*2758*/;
assign _12986_ = _13113_ ^ _13120_ /*2759*/;
assign _13118_ = _13119_ | _13121_ /*2756*/;
assign _13127_ = ~D[26] /*2755*/;
assign _13124_ = _12762_ & _13127_ /*2751*/;
assign _13125_ = _12762_ ^ _13127_ /*2754*/;
assign _13126_ = _13118_ & _13125_ /*2752*/;
assign _12987_ = _13118_ ^ _13125_ /*2753*/;
assign _13123_ = _13124_ | _13126_ /*2750*/;
assign _13132_ = ~D[27] /*2749*/;
assign _13129_ = _12763_ & _13132_ /*2745*/;
assign _13130_ = _12763_ ^ _13132_ /*2748*/;
assign _13131_ = _13123_ & _13130_ /*2746*/;
assign _12988_ = _13123_ ^ _13130_ /*2747*/;
assign _13128_ = _13129_ | _13131_ /*2744*/;
assign _13137_ = ~D[28] /*2743*/;
assign _13134_ = _12764_ & _13137_ /*2739*/;
assign _13135_ = _12764_ ^ _13137_ /*2742*/;
assign _13136_ = _13128_ & _13135_ /*2740*/;
assign _12989_ = _13128_ ^ _13135_ /*2741*/;
assign _13133_ = _13134_ | _13136_ /*2738*/;
assign _13142_ = ~D[29] /*2737*/;
assign _13139_ = _12765_ & _13142_ /*2733*/;
assign _13140_ = _12765_ ^ _13142_ /*2736*/;
assign _13141_ = _13133_ & _13140_ /*2734*/;
assign _12990_ = _13133_ ^ _13140_ /*2735*/;
assign _13138_ = _13139_ | _13141_ /*2732*/;
assign _13147_ = ~D[30] /*2731*/;
assign _13144_ = _12766_ & _13147_ /*2727*/;
assign _13145_ = _12766_ ^ _13147_ /*2730*/;
assign _13146_ = _13138_ & _13145_ /*2728*/;
assign _12991_ = _13138_ ^ _13145_ /*2729*/;
assign _13143_ = _13144_ | _13146_ /*2726*/;
assign _13148_ = _12767_ & oneWire /*2721*/;
assign _13149_ = _12767_ ^ oneWire /*2724*/;
assign _13150_ = _13143_ & _13149_ /*2722*/;
assign _12992_ = _13143_ ^ _13149_ /*2723*/;
assign Q[2] = _13148_ | _13150_ /*2720*/;
assign _13219_ = ~Q[2] /*2527*/;
assign _13218_ = _13219_ & D[0] /*2526*/;
assign _13221_ = _12961_ & _13218_ /*2521*/;
assign _13222_ = _12961_ ^ _13218_ /*2524*/;
assign _13223_ = zeroWire & _13222_ /*2522*/;
assign _13185_ = zeroWire ^ _13222_ /*2523*/;
assign _13220_ = _13221_ | _13223_ /*2520*/;
assign _13225_ = ~Q[2] /*2519*/;
assign _13224_ = _13225_ & D[1] /*2518*/;
assign _13227_ = _12962_ & _13224_ /*2513*/;
assign _13228_ = _12962_ ^ _13224_ /*2516*/;
assign _13229_ = _13220_ & _13228_ /*2514*/;
assign _13186_ = _13220_ ^ _13228_ /*2515*/;
assign _13226_ = _13227_ | _13229_ /*2512*/;
assign _13231_ = ~Q[2] /*2511*/;
assign _13230_ = _13231_ & D[2] /*2510*/;
assign _13233_ = _12963_ & _13230_ /*2505*/;
assign _13234_ = _12963_ ^ _13230_ /*2508*/;
assign _13235_ = _13226_ & _13234_ /*2506*/;
assign _13187_ = _13226_ ^ _13234_ /*2507*/;
assign _13232_ = _13233_ | _13235_ /*2504*/;
assign _13237_ = ~Q[2] /*2503*/;
assign _13236_ = _13237_ & D[3] /*2502*/;
assign _13239_ = _12964_ & _13236_ /*2497*/;
assign _13240_ = _12964_ ^ _13236_ /*2500*/;
assign _13241_ = _13232_ & _13240_ /*2498*/;
assign _13188_ = _13232_ ^ _13240_ /*2499*/;
assign _13238_ = _13239_ | _13241_ /*2496*/;
assign _13243_ = ~Q[2] /*2495*/;
assign _13242_ = _13243_ & D[4] /*2494*/;
assign _13245_ = _12965_ & _13242_ /*2489*/;
assign _13246_ = _12965_ ^ _13242_ /*2492*/;
assign _13247_ = _13238_ & _13246_ /*2490*/;
assign _13189_ = _13238_ ^ _13246_ /*2491*/;
assign _13244_ = _13245_ | _13247_ /*2488*/;
assign _13249_ = ~Q[2] /*2487*/;
assign _13248_ = _13249_ & D[5] /*2486*/;
assign _13251_ = _12966_ & _13248_ /*2481*/;
assign _13252_ = _12966_ ^ _13248_ /*2484*/;
assign _13253_ = _13244_ & _13252_ /*2482*/;
assign _13190_ = _13244_ ^ _13252_ /*2483*/;
assign _13250_ = _13251_ | _13253_ /*2480*/;
assign _13255_ = ~Q[2] /*2479*/;
assign _13254_ = _13255_ & D[6] /*2478*/;
assign _13257_ = _12967_ & _13254_ /*2473*/;
assign _13258_ = _12967_ ^ _13254_ /*2476*/;
assign _13259_ = _13250_ & _13258_ /*2474*/;
assign _13191_ = _13250_ ^ _13258_ /*2475*/;
assign _13256_ = _13257_ | _13259_ /*2472*/;
assign _13261_ = ~Q[2] /*2471*/;
assign _13260_ = _13261_ & D[7] /*2470*/;
assign _13263_ = _12968_ & _13260_ /*2465*/;
assign _13264_ = _12968_ ^ _13260_ /*2468*/;
assign _13265_ = _13256_ & _13264_ /*2466*/;
assign _13192_ = _13256_ ^ _13264_ /*2467*/;
assign _13262_ = _13263_ | _13265_ /*2464*/;
assign _13267_ = ~Q[2] /*2463*/;
assign _13266_ = _13267_ & D[8] /*2462*/;
assign _13269_ = _12969_ & _13266_ /*2457*/;
assign _13270_ = _12969_ ^ _13266_ /*2460*/;
assign _13271_ = _13262_ & _13270_ /*2458*/;
assign _13193_ = _13262_ ^ _13270_ /*2459*/;
assign _13268_ = _13269_ | _13271_ /*2456*/;
assign _13273_ = ~Q[2] /*2455*/;
assign _13272_ = _13273_ & D[9] /*2454*/;
assign _13275_ = _12970_ & _13272_ /*2449*/;
assign _13276_ = _12970_ ^ _13272_ /*2452*/;
assign _13277_ = _13268_ & _13276_ /*2450*/;
assign _13194_ = _13268_ ^ _13276_ /*2451*/;
assign _13274_ = _13275_ | _13277_ /*2448*/;
assign _13279_ = ~Q[2] /*2447*/;
assign _13278_ = _13279_ & D[10] /*2446*/;
assign _13281_ = _12971_ & _13278_ /*2441*/;
assign _13282_ = _12971_ ^ _13278_ /*2444*/;
assign _13283_ = _13274_ & _13282_ /*2442*/;
assign _13195_ = _13274_ ^ _13282_ /*2443*/;
assign _13280_ = _13281_ | _13283_ /*2440*/;
assign _13285_ = ~Q[2] /*2439*/;
assign _13284_ = _13285_ & D[11] /*2438*/;
assign _13287_ = _12972_ & _13284_ /*2433*/;
assign _13288_ = _12972_ ^ _13284_ /*2436*/;
assign _13289_ = _13280_ & _13288_ /*2434*/;
assign _13196_ = _13280_ ^ _13288_ /*2435*/;
assign _13286_ = _13287_ | _13289_ /*2432*/;
assign _13291_ = ~Q[2] /*2431*/;
assign _13290_ = _13291_ & D[12] /*2430*/;
assign _13293_ = _12973_ & _13290_ /*2425*/;
assign _13294_ = _12973_ ^ _13290_ /*2428*/;
assign _13295_ = _13286_ & _13294_ /*2426*/;
assign _13197_ = _13286_ ^ _13294_ /*2427*/;
assign _13292_ = _13293_ | _13295_ /*2424*/;
assign _13297_ = ~Q[2] /*2423*/;
assign _13296_ = _13297_ & D[13] /*2422*/;
assign _13299_ = _12974_ & _13296_ /*2417*/;
assign _13300_ = _12974_ ^ _13296_ /*2420*/;
assign _13301_ = _13292_ & _13300_ /*2418*/;
assign _13198_ = _13292_ ^ _13300_ /*2419*/;
assign _13298_ = _13299_ | _13301_ /*2416*/;
assign _13303_ = ~Q[2] /*2415*/;
assign _13302_ = _13303_ & D[14] /*2414*/;
assign _13305_ = _12975_ & _13302_ /*2409*/;
assign _13306_ = _12975_ ^ _13302_ /*2412*/;
assign _13307_ = _13298_ & _13306_ /*2410*/;
assign _13199_ = _13298_ ^ _13306_ /*2411*/;
assign _13304_ = _13305_ | _13307_ /*2408*/;
assign _13309_ = ~Q[2] /*2407*/;
assign _13308_ = _13309_ & D[15] /*2406*/;
assign _13311_ = _12976_ & _13308_ /*2401*/;
assign _13312_ = _12976_ ^ _13308_ /*2404*/;
assign _13313_ = _13304_ & _13312_ /*2402*/;
assign _13200_ = _13304_ ^ _13312_ /*2403*/;
assign _13310_ = _13311_ | _13313_ /*2400*/;
assign _13315_ = ~Q[2] /*2399*/;
assign _13314_ = _13315_ & D[16] /*2398*/;
assign _13317_ = _12977_ & _13314_ /*2393*/;
assign _13318_ = _12977_ ^ _13314_ /*2396*/;
assign _13319_ = _13310_ & _13318_ /*2394*/;
assign _13201_ = _13310_ ^ _13318_ /*2395*/;
assign _13316_ = _13317_ | _13319_ /*2392*/;
assign _13321_ = ~Q[2] /*2391*/;
assign _13320_ = _13321_ & D[17] /*2390*/;
assign _13323_ = _12978_ & _13320_ /*2385*/;
assign _13324_ = _12978_ ^ _13320_ /*2388*/;
assign _13325_ = _13316_ & _13324_ /*2386*/;
assign _13202_ = _13316_ ^ _13324_ /*2387*/;
assign _13322_ = _13323_ | _13325_ /*2384*/;
assign _13327_ = ~Q[2] /*2383*/;
assign _13326_ = _13327_ & D[18] /*2382*/;
assign _13329_ = _12979_ & _13326_ /*2377*/;
assign _13330_ = _12979_ ^ _13326_ /*2380*/;
assign _13331_ = _13322_ & _13330_ /*2378*/;
assign _13203_ = _13322_ ^ _13330_ /*2379*/;
assign _13328_ = _13329_ | _13331_ /*2376*/;
assign _13333_ = ~Q[2] /*2375*/;
assign _13332_ = _13333_ & D[19] /*2374*/;
assign _13335_ = _12980_ & _13332_ /*2369*/;
assign _13336_ = _12980_ ^ _13332_ /*2372*/;
assign _13337_ = _13328_ & _13336_ /*2370*/;
assign _13204_ = _13328_ ^ _13336_ /*2371*/;
assign _13334_ = _13335_ | _13337_ /*2368*/;
assign _13339_ = ~Q[2] /*2367*/;
assign _13338_ = _13339_ & D[20] /*2366*/;
assign _13341_ = _12981_ & _13338_ /*2361*/;
assign _13342_ = _12981_ ^ _13338_ /*2364*/;
assign _13343_ = _13334_ & _13342_ /*2362*/;
assign _13205_ = _13334_ ^ _13342_ /*2363*/;
assign _13340_ = _13341_ | _13343_ /*2360*/;
assign _13345_ = ~Q[2] /*2359*/;
assign _13344_ = _13345_ & D[21] /*2358*/;
assign _13347_ = _12982_ & _13344_ /*2353*/;
assign _13348_ = _12982_ ^ _13344_ /*2356*/;
assign _13349_ = _13340_ & _13348_ /*2354*/;
assign _13206_ = _13340_ ^ _13348_ /*2355*/;
assign _13346_ = _13347_ | _13349_ /*2352*/;
assign _13351_ = ~Q[2] /*2351*/;
assign _13350_ = _13351_ & D[22] /*2350*/;
assign _13353_ = _12983_ & _13350_ /*2345*/;
assign _13354_ = _12983_ ^ _13350_ /*2348*/;
assign _13355_ = _13346_ & _13354_ /*2346*/;
assign _13207_ = _13346_ ^ _13354_ /*2347*/;
assign _13352_ = _13353_ | _13355_ /*2344*/;
assign _13357_ = ~Q[2] /*2343*/;
assign _13356_ = _13357_ & D[23] /*2342*/;
assign _13359_ = _12984_ & _13356_ /*2337*/;
assign _13360_ = _12984_ ^ _13356_ /*2340*/;
assign _13361_ = _13352_ & _13360_ /*2338*/;
assign _13208_ = _13352_ ^ _13360_ /*2339*/;
assign _13358_ = _13359_ | _13361_ /*2336*/;
assign _13363_ = ~Q[2] /*2335*/;
assign _13362_ = _13363_ & D[24] /*2334*/;
assign _13365_ = _12985_ & _13362_ /*2329*/;
assign _13366_ = _12985_ ^ _13362_ /*2332*/;
assign _13367_ = _13358_ & _13366_ /*2330*/;
assign _13209_ = _13358_ ^ _13366_ /*2331*/;
assign _13364_ = _13365_ | _13367_ /*2328*/;
assign _13369_ = ~Q[2] /*2327*/;
assign _13368_ = _13369_ & D[25] /*2326*/;
assign _13371_ = _12986_ & _13368_ /*2321*/;
assign _13372_ = _12986_ ^ _13368_ /*2324*/;
assign _13373_ = _13364_ & _13372_ /*2322*/;
assign _13210_ = _13364_ ^ _13372_ /*2323*/;
assign _13370_ = _13371_ | _13373_ /*2320*/;
assign _13375_ = ~Q[2] /*2319*/;
assign _13374_ = _13375_ & D[26] /*2318*/;
assign _13377_ = _12987_ & _13374_ /*2313*/;
assign _13378_ = _12987_ ^ _13374_ /*2316*/;
assign _13379_ = _13370_ & _13378_ /*2314*/;
assign _13211_ = _13370_ ^ _13378_ /*2315*/;
assign _13376_ = _13377_ | _13379_ /*2312*/;
assign _13381_ = ~Q[2] /*2311*/;
assign _13380_ = _13381_ & D[27] /*2310*/;
assign _13383_ = _12988_ & _13380_ /*2305*/;
assign _13384_ = _12988_ ^ _13380_ /*2308*/;
assign _13385_ = _13376_ & _13384_ /*2306*/;
assign _13212_ = _13376_ ^ _13384_ /*2307*/;
assign _13382_ = _13383_ | _13385_ /*2304*/;
assign _13387_ = ~Q[2] /*2303*/;
assign _13386_ = _13387_ & D[28] /*2302*/;
assign _13389_ = _12989_ & _13386_ /*2297*/;
assign _13390_ = _12989_ ^ _13386_ /*2300*/;
assign _13391_ = _13382_ & _13390_ /*2298*/;
assign _13213_ = _13382_ ^ _13390_ /*2299*/;
assign _13388_ = _13389_ | _13391_ /*2296*/;
assign _13393_ = ~Q[2] /*2295*/;
assign _13392_ = _13393_ & D[29] /*2294*/;
assign _13395_ = _12990_ & _13392_ /*2289*/;
assign _13396_ = _12990_ ^ _13392_ /*2292*/;
assign _13397_ = _13388_ & _13396_ /*2290*/;
assign _13214_ = _13388_ ^ _13396_ /*2291*/;
assign _13394_ = _13395_ | _13397_ /*2288*/;
assign _13399_ = ~Q[2] /*2287*/;
assign _13398_ = _13399_ & D[30] /*2286*/;
assign _13401_ = _12991_ & _13398_ /*2281*/;
assign _13402_ = _12991_ ^ _13398_ /*2284*/;
assign _13403_ = _13394_ & _13402_ /*2282*/;
assign _13215_ = _13394_ ^ _13402_ /*2283*/;
assign _13400_ = _13401_ | _13403_ /*2280*/;
assign _13405_ = ~Q[2] /*2279*/;
assign _13404_ = _13405_ & zeroWire /*2278*/;
assign _13406_ = _12992_ ^ _13404_ /*2276*/;
assign _13216_ = _13406_ ^ _13400_ /*2275*/;
assign _13445_ = ~D[0] /*2149*/;
assign _13442_ = R_0[1] & _13445_ /*2145*/;
assign _13443_ = R_0[1] ^ _13445_ /*2148*/;
assign _13444_ = oneWire & _13443_ /*2146*/;
assign _13409_ = oneWire ^ _13443_ /*2147*/;
assign _13441_ = _13442_ | _13444_ /*2144*/;
assign _13450_ = ~D[1] /*2143*/;
assign _13447_ = _13185_ & _13450_ /*2139*/;
assign _13448_ = _13185_ ^ _13450_ /*2142*/;
assign _13449_ = _13441_ & _13448_ /*2140*/;
assign _13410_ = _13441_ ^ _13448_ /*2141*/;
assign _13446_ = _13447_ | _13449_ /*2138*/;
assign _13455_ = ~D[2] /*2137*/;
assign _13452_ = _13186_ & _13455_ /*2133*/;
assign _13453_ = _13186_ ^ _13455_ /*2136*/;
assign _13454_ = _13446_ & _13453_ /*2134*/;
assign _13411_ = _13446_ ^ _13453_ /*2135*/;
assign _13451_ = _13452_ | _13454_ /*2132*/;
assign _13460_ = ~D[3] /*2131*/;
assign _13457_ = _13187_ & _13460_ /*2127*/;
assign _13458_ = _13187_ ^ _13460_ /*2130*/;
assign _13459_ = _13451_ & _13458_ /*2128*/;
assign _13412_ = _13451_ ^ _13458_ /*2129*/;
assign _13456_ = _13457_ | _13459_ /*2126*/;
assign _13465_ = ~D[4] /*2125*/;
assign _13462_ = _13188_ & _13465_ /*2121*/;
assign _13463_ = _13188_ ^ _13465_ /*2124*/;
assign _13464_ = _13456_ & _13463_ /*2122*/;
assign _13413_ = _13456_ ^ _13463_ /*2123*/;
assign _13461_ = _13462_ | _13464_ /*2120*/;
assign _13470_ = ~D[5] /*2119*/;
assign _13467_ = _13189_ & _13470_ /*2115*/;
assign _13468_ = _13189_ ^ _13470_ /*2118*/;
assign _13469_ = _13461_ & _13468_ /*2116*/;
assign _13414_ = _13461_ ^ _13468_ /*2117*/;
assign _13466_ = _13467_ | _13469_ /*2114*/;
assign _13475_ = ~D[6] /*2113*/;
assign _13472_ = _13190_ & _13475_ /*2109*/;
assign _13473_ = _13190_ ^ _13475_ /*2112*/;
assign _13474_ = _13466_ & _13473_ /*2110*/;
assign _13415_ = _13466_ ^ _13473_ /*2111*/;
assign _13471_ = _13472_ | _13474_ /*2108*/;
assign _13480_ = ~D[7] /*2107*/;
assign _13477_ = _13191_ & _13480_ /*2103*/;
assign _13478_ = _13191_ ^ _13480_ /*2106*/;
assign _13479_ = _13471_ & _13478_ /*2104*/;
assign _13416_ = _13471_ ^ _13478_ /*2105*/;
assign _13476_ = _13477_ | _13479_ /*2102*/;
assign _13485_ = ~D[8] /*2101*/;
assign _13482_ = _13192_ & _13485_ /*2097*/;
assign _13483_ = _13192_ ^ _13485_ /*2100*/;
assign _13484_ = _13476_ & _13483_ /*2098*/;
assign _13417_ = _13476_ ^ _13483_ /*2099*/;
assign _13481_ = _13482_ | _13484_ /*2096*/;
assign _13490_ = ~D[9] /*2095*/;
assign _13487_ = _13193_ & _13490_ /*2091*/;
assign _13488_ = _13193_ ^ _13490_ /*2094*/;
assign _13489_ = _13481_ & _13488_ /*2092*/;
assign _13418_ = _13481_ ^ _13488_ /*2093*/;
assign _13486_ = _13487_ | _13489_ /*2090*/;
assign _13495_ = ~D[10] /*2089*/;
assign _13492_ = _13194_ & _13495_ /*2085*/;
assign _13493_ = _13194_ ^ _13495_ /*2088*/;
assign _13494_ = _13486_ & _13493_ /*2086*/;
assign _13419_ = _13486_ ^ _13493_ /*2087*/;
assign _13491_ = _13492_ | _13494_ /*2084*/;
assign _13500_ = ~D[11] /*2083*/;
assign _13497_ = _13195_ & _13500_ /*2079*/;
assign _13498_ = _13195_ ^ _13500_ /*2082*/;
assign _13499_ = _13491_ & _13498_ /*2080*/;
assign _13420_ = _13491_ ^ _13498_ /*2081*/;
assign _13496_ = _13497_ | _13499_ /*2078*/;
assign _13505_ = ~D[12] /*2077*/;
assign _13502_ = _13196_ & _13505_ /*2073*/;
assign _13503_ = _13196_ ^ _13505_ /*2076*/;
assign _13504_ = _13496_ & _13503_ /*2074*/;
assign _13421_ = _13496_ ^ _13503_ /*2075*/;
assign _13501_ = _13502_ | _13504_ /*2072*/;
assign _13510_ = ~D[13] /*2071*/;
assign _13507_ = _13197_ & _13510_ /*2067*/;
assign _13508_ = _13197_ ^ _13510_ /*2070*/;
assign _13509_ = _13501_ & _13508_ /*2068*/;
assign _13422_ = _13501_ ^ _13508_ /*2069*/;
assign _13506_ = _13507_ | _13509_ /*2066*/;
assign _13515_ = ~D[14] /*2065*/;
assign _13512_ = _13198_ & _13515_ /*2061*/;
assign _13513_ = _13198_ ^ _13515_ /*2064*/;
assign _13514_ = _13506_ & _13513_ /*2062*/;
assign _13423_ = _13506_ ^ _13513_ /*2063*/;
assign _13511_ = _13512_ | _13514_ /*2060*/;
assign _13520_ = ~D[15] /*2059*/;
assign _13517_ = _13199_ & _13520_ /*2055*/;
assign _13518_ = _13199_ ^ _13520_ /*2058*/;
assign _13519_ = _13511_ & _13518_ /*2056*/;
assign _13424_ = _13511_ ^ _13518_ /*2057*/;
assign _13516_ = _13517_ | _13519_ /*2054*/;
assign _13525_ = ~D[16] /*2053*/;
assign _13522_ = _13200_ & _13525_ /*2049*/;
assign _13523_ = _13200_ ^ _13525_ /*2052*/;
assign _13524_ = _13516_ & _13523_ /*2050*/;
assign _13425_ = _13516_ ^ _13523_ /*2051*/;
assign _13521_ = _13522_ | _13524_ /*2048*/;
assign _13530_ = ~D[17] /*2047*/;
assign _13527_ = _13201_ & _13530_ /*2043*/;
assign _13528_ = _13201_ ^ _13530_ /*2046*/;
assign _13529_ = _13521_ & _13528_ /*2044*/;
assign _13426_ = _13521_ ^ _13528_ /*2045*/;
assign _13526_ = _13527_ | _13529_ /*2042*/;
assign _13535_ = ~D[18] /*2041*/;
assign _13532_ = _13202_ & _13535_ /*2037*/;
assign _13533_ = _13202_ ^ _13535_ /*2040*/;
assign _13534_ = _13526_ & _13533_ /*2038*/;
assign _13427_ = _13526_ ^ _13533_ /*2039*/;
assign _13531_ = _13532_ | _13534_ /*2036*/;
assign _13540_ = ~D[19] /*2035*/;
assign _13537_ = _13203_ & _13540_ /*2031*/;
assign _13538_ = _13203_ ^ _13540_ /*2034*/;
assign _13539_ = _13531_ & _13538_ /*2032*/;
assign _13428_ = _13531_ ^ _13538_ /*2033*/;
assign _13536_ = _13537_ | _13539_ /*2030*/;
assign _13545_ = ~D[20] /*2029*/;
assign _13542_ = _13204_ & _13545_ /*2025*/;
assign _13543_ = _13204_ ^ _13545_ /*2028*/;
assign _13544_ = _13536_ & _13543_ /*2026*/;
assign _13429_ = _13536_ ^ _13543_ /*2027*/;
assign _13541_ = _13542_ | _13544_ /*2024*/;
assign _13550_ = ~D[21] /*2023*/;
assign _13547_ = _13205_ & _13550_ /*2019*/;
assign _13548_ = _13205_ ^ _13550_ /*2022*/;
assign _13549_ = _13541_ & _13548_ /*2020*/;
assign _13430_ = _13541_ ^ _13548_ /*2021*/;
assign _13546_ = _13547_ | _13549_ /*2018*/;
assign _13555_ = ~D[22] /*2017*/;
assign _13552_ = _13206_ & _13555_ /*2013*/;
assign _13553_ = _13206_ ^ _13555_ /*2016*/;
assign _13554_ = _13546_ & _13553_ /*2014*/;
assign _13431_ = _13546_ ^ _13553_ /*2015*/;
assign _13551_ = _13552_ | _13554_ /*2012*/;
assign _13560_ = ~D[23] /*2011*/;
assign _13557_ = _13207_ & _13560_ /*2007*/;
assign _13558_ = _13207_ ^ _13560_ /*2010*/;
assign _13559_ = _13551_ & _13558_ /*2008*/;
assign _13432_ = _13551_ ^ _13558_ /*2009*/;
assign _13556_ = _13557_ | _13559_ /*2006*/;
assign _13565_ = ~D[24] /*2005*/;
assign _13562_ = _13208_ & _13565_ /*2001*/;
assign _13563_ = _13208_ ^ _13565_ /*2004*/;
assign _13564_ = _13556_ & _13563_ /*2002*/;
assign _13433_ = _13556_ ^ _13563_ /*2003*/;
assign _13561_ = _13562_ | _13564_ /*2000*/;
assign _13570_ = ~D[25] /*1999*/;
assign _13567_ = _13209_ & _13570_ /*1995*/;
assign _13568_ = _13209_ ^ _13570_ /*1998*/;
assign _13569_ = _13561_ & _13568_ /*1996*/;
assign _13434_ = _13561_ ^ _13568_ /*1997*/;
assign _13566_ = _13567_ | _13569_ /*1994*/;
assign _13575_ = ~D[26] /*1993*/;
assign _13572_ = _13210_ & _13575_ /*1989*/;
assign _13573_ = _13210_ ^ _13575_ /*1992*/;
assign _13574_ = _13566_ & _13573_ /*1990*/;
assign _13435_ = _13566_ ^ _13573_ /*1991*/;
assign _13571_ = _13572_ | _13574_ /*1988*/;
assign _13580_ = ~D[27] /*1987*/;
assign _13577_ = _13211_ & _13580_ /*1983*/;
assign _13578_ = _13211_ ^ _13580_ /*1986*/;
assign _13579_ = _13571_ & _13578_ /*1984*/;
assign _13436_ = _13571_ ^ _13578_ /*1985*/;
assign _13576_ = _13577_ | _13579_ /*1982*/;
assign _13585_ = ~D[28] /*1981*/;
assign _13582_ = _13212_ & _13585_ /*1977*/;
assign _13583_ = _13212_ ^ _13585_ /*1980*/;
assign _13584_ = _13576_ & _13583_ /*1978*/;
assign _13437_ = _13576_ ^ _13583_ /*1979*/;
assign _13581_ = _13582_ | _13584_ /*1976*/;
assign _13590_ = ~D[29] /*1975*/;
assign _13587_ = _13213_ & _13590_ /*1971*/;
assign _13588_ = _13213_ ^ _13590_ /*1974*/;
assign _13589_ = _13581_ & _13588_ /*1972*/;
assign _13438_ = _13581_ ^ _13588_ /*1973*/;
assign _13586_ = _13587_ | _13589_ /*1970*/;
assign _13595_ = ~D[30] /*1969*/;
assign _13592_ = _13214_ & _13595_ /*1965*/;
assign _13593_ = _13214_ ^ _13595_ /*1968*/;
assign _13594_ = _13586_ & _13593_ /*1966*/;
assign _13439_ = _13586_ ^ _13593_ /*1967*/;
assign _13591_ = _13592_ | _13594_ /*1964*/;
assign _13596_ = _13215_ & oneWire /*1959*/;
assign _13597_ = _13215_ ^ oneWire /*1962*/;
assign _13598_ = _13591_ & _13597_ /*1960*/;
assign _13440_ = _13591_ ^ _13597_ /*1961*/;
assign Q[1] = _13596_ | _13598_ /*1958*/;
assign _13667_ = ~Q[1] /*1765*/;
assign _13666_ = _13667_ & D[0] /*1764*/;
assign _13669_ = _13409_ & _13666_ /*1759*/;
assign _13670_ = _13409_ ^ _13666_ /*1762*/;
assign _13671_ = zeroWire & _13670_ /*1760*/;
assign _13633_ = zeroWire ^ _13670_ /*1761*/;
assign _13668_ = _13669_ | _13671_ /*1758*/;
assign _13673_ = ~Q[1] /*1757*/;
assign _13672_ = _13673_ & D[1] /*1756*/;
assign _13675_ = _13410_ & _13672_ /*1751*/;
assign _13676_ = _13410_ ^ _13672_ /*1754*/;
assign _13677_ = _13668_ & _13676_ /*1752*/;
assign _13634_ = _13668_ ^ _13676_ /*1753*/;
assign _13674_ = _13675_ | _13677_ /*1750*/;
assign _13679_ = ~Q[1] /*1749*/;
assign _13678_ = _13679_ & D[2] /*1748*/;
assign _13681_ = _13411_ & _13678_ /*1743*/;
assign _13682_ = _13411_ ^ _13678_ /*1746*/;
assign _13683_ = _13674_ & _13682_ /*1744*/;
assign _13635_ = _13674_ ^ _13682_ /*1745*/;
assign _13680_ = _13681_ | _13683_ /*1742*/;
assign _13685_ = ~Q[1] /*1741*/;
assign _13684_ = _13685_ & D[3] /*1740*/;
assign _13687_ = _13412_ & _13684_ /*1735*/;
assign _13688_ = _13412_ ^ _13684_ /*1738*/;
assign _13689_ = _13680_ & _13688_ /*1736*/;
assign _13636_ = _13680_ ^ _13688_ /*1737*/;
assign _13686_ = _13687_ | _13689_ /*1734*/;
assign _13691_ = ~Q[1] /*1733*/;
assign _13690_ = _13691_ & D[4] /*1732*/;
assign _13693_ = _13413_ & _13690_ /*1727*/;
assign _13694_ = _13413_ ^ _13690_ /*1730*/;
assign _13695_ = _13686_ & _13694_ /*1728*/;
assign _13637_ = _13686_ ^ _13694_ /*1729*/;
assign _13692_ = _13693_ | _13695_ /*1726*/;
assign _13697_ = ~Q[1] /*1725*/;
assign _13696_ = _13697_ & D[5] /*1724*/;
assign _13699_ = _13414_ & _13696_ /*1719*/;
assign _13700_ = _13414_ ^ _13696_ /*1722*/;
assign _13701_ = _13692_ & _13700_ /*1720*/;
assign _13638_ = _13692_ ^ _13700_ /*1721*/;
assign _13698_ = _13699_ | _13701_ /*1718*/;
assign _13703_ = ~Q[1] /*1717*/;
assign _13702_ = _13703_ & D[6] /*1716*/;
assign _13705_ = _13415_ & _13702_ /*1711*/;
assign _13706_ = _13415_ ^ _13702_ /*1714*/;
assign _13707_ = _13698_ & _13706_ /*1712*/;
assign _13639_ = _13698_ ^ _13706_ /*1713*/;
assign _13704_ = _13705_ | _13707_ /*1710*/;
assign _13709_ = ~Q[1] /*1709*/;
assign _13708_ = _13709_ & D[7] /*1708*/;
assign _13711_ = _13416_ & _13708_ /*1703*/;
assign _13712_ = _13416_ ^ _13708_ /*1706*/;
assign _13713_ = _13704_ & _13712_ /*1704*/;
assign _13640_ = _13704_ ^ _13712_ /*1705*/;
assign _13710_ = _13711_ | _13713_ /*1702*/;
assign _13715_ = ~Q[1] /*1701*/;
assign _13714_ = _13715_ & D[8] /*1700*/;
assign _13717_ = _13417_ & _13714_ /*1695*/;
assign _13718_ = _13417_ ^ _13714_ /*1698*/;
assign _13719_ = _13710_ & _13718_ /*1696*/;
assign _13641_ = _13710_ ^ _13718_ /*1697*/;
assign _13716_ = _13717_ | _13719_ /*1694*/;
assign _13721_ = ~Q[1] /*1693*/;
assign _13720_ = _13721_ & D[9] /*1692*/;
assign _13723_ = _13418_ & _13720_ /*1687*/;
assign _13724_ = _13418_ ^ _13720_ /*1690*/;
assign _13725_ = _13716_ & _13724_ /*1688*/;
assign _13642_ = _13716_ ^ _13724_ /*1689*/;
assign _13722_ = _13723_ | _13725_ /*1686*/;
assign _13727_ = ~Q[1] /*1685*/;
assign _13726_ = _13727_ & D[10] /*1684*/;
assign _13729_ = _13419_ & _13726_ /*1679*/;
assign _13730_ = _13419_ ^ _13726_ /*1682*/;
assign _13731_ = _13722_ & _13730_ /*1680*/;
assign _13643_ = _13722_ ^ _13730_ /*1681*/;
assign _13728_ = _13729_ | _13731_ /*1678*/;
assign _13733_ = ~Q[1] /*1677*/;
assign _13732_ = _13733_ & D[11] /*1676*/;
assign _13735_ = _13420_ & _13732_ /*1671*/;
assign _13736_ = _13420_ ^ _13732_ /*1674*/;
assign _13737_ = _13728_ & _13736_ /*1672*/;
assign _13644_ = _13728_ ^ _13736_ /*1673*/;
assign _13734_ = _13735_ | _13737_ /*1670*/;
assign _13739_ = ~Q[1] /*1669*/;
assign _13738_ = _13739_ & D[12] /*1668*/;
assign _13741_ = _13421_ & _13738_ /*1663*/;
assign _13742_ = _13421_ ^ _13738_ /*1666*/;
assign _13743_ = _13734_ & _13742_ /*1664*/;
assign _13645_ = _13734_ ^ _13742_ /*1665*/;
assign _13740_ = _13741_ | _13743_ /*1662*/;
assign _13745_ = ~Q[1] /*1661*/;
assign _13744_ = _13745_ & D[13] /*1660*/;
assign _13747_ = _13422_ & _13744_ /*1655*/;
assign _13748_ = _13422_ ^ _13744_ /*1658*/;
assign _13749_ = _13740_ & _13748_ /*1656*/;
assign _13646_ = _13740_ ^ _13748_ /*1657*/;
assign _13746_ = _13747_ | _13749_ /*1654*/;
assign _13751_ = ~Q[1] /*1653*/;
assign _13750_ = _13751_ & D[14] /*1652*/;
assign _13753_ = _13423_ & _13750_ /*1647*/;
assign _13754_ = _13423_ ^ _13750_ /*1650*/;
assign _13755_ = _13746_ & _13754_ /*1648*/;
assign _13647_ = _13746_ ^ _13754_ /*1649*/;
assign _13752_ = _13753_ | _13755_ /*1646*/;
assign _13757_ = ~Q[1] /*1645*/;
assign _13756_ = _13757_ & D[15] /*1644*/;
assign _13759_ = _13424_ & _13756_ /*1639*/;
assign _13760_ = _13424_ ^ _13756_ /*1642*/;
assign _13761_ = _13752_ & _13760_ /*1640*/;
assign _13648_ = _13752_ ^ _13760_ /*1641*/;
assign _13758_ = _13759_ | _13761_ /*1638*/;
assign _13763_ = ~Q[1] /*1637*/;
assign _13762_ = _13763_ & D[16] /*1636*/;
assign _13765_ = _13425_ & _13762_ /*1631*/;
assign _13766_ = _13425_ ^ _13762_ /*1634*/;
assign _13767_ = _13758_ & _13766_ /*1632*/;
assign _13649_ = _13758_ ^ _13766_ /*1633*/;
assign _13764_ = _13765_ | _13767_ /*1630*/;
assign _13769_ = ~Q[1] /*1629*/;
assign _13768_ = _13769_ & D[17] /*1628*/;
assign _13771_ = _13426_ & _13768_ /*1623*/;
assign _13772_ = _13426_ ^ _13768_ /*1626*/;
assign _13773_ = _13764_ & _13772_ /*1624*/;
assign _13650_ = _13764_ ^ _13772_ /*1625*/;
assign _13770_ = _13771_ | _13773_ /*1622*/;
assign _13775_ = ~Q[1] /*1621*/;
assign _13774_ = _13775_ & D[18] /*1620*/;
assign _13777_ = _13427_ & _13774_ /*1615*/;
assign _13778_ = _13427_ ^ _13774_ /*1618*/;
assign _13779_ = _13770_ & _13778_ /*1616*/;
assign _13651_ = _13770_ ^ _13778_ /*1617*/;
assign _13776_ = _13777_ | _13779_ /*1614*/;
assign _13781_ = ~Q[1] /*1613*/;
assign _13780_ = _13781_ & D[19] /*1612*/;
assign _13783_ = _13428_ & _13780_ /*1607*/;
assign _13784_ = _13428_ ^ _13780_ /*1610*/;
assign _13785_ = _13776_ & _13784_ /*1608*/;
assign _13652_ = _13776_ ^ _13784_ /*1609*/;
assign _13782_ = _13783_ | _13785_ /*1606*/;
assign _13787_ = ~Q[1] /*1605*/;
assign _13786_ = _13787_ & D[20] /*1604*/;
assign _13789_ = _13429_ & _13786_ /*1599*/;
assign _13790_ = _13429_ ^ _13786_ /*1602*/;
assign _13791_ = _13782_ & _13790_ /*1600*/;
assign _13653_ = _13782_ ^ _13790_ /*1601*/;
assign _13788_ = _13789_ | _13791_ /*1598*/;
assign _13793_ = ~Q[1] /*1597*/;
assign _13792_ = _13793_ & D[21] /*1596*/;
assign _13795_ = _13430_ & _13792_ /*1591*/;
assign _13796_ = _13430_ ^ _13792_ /*1594*/;
assign _13797_ = _13788_ & _13796_ /*1592*/;
assign _13654_ = _13788_ ^ _13796_ /*1593*/;
assign _13794_ = _13795_ | _13797_ /*1590*/;
assign _13799_ = ~Q[1] /*1589*/;
assign _13798_ = _13799_ & D[22] /*1588*/;
assign _13801_ = _13431_ & _13798_ /*1583*/;
assign _13802_ = _13431_ ^ _13798_ /*1586*/;
assign _13803_ = _13794_ & _13802_ /*1584*/;
assign _13655_ = _13794_ ^ _13802_ /*1585*/;
assign _13800_ = _13801_ | _13803_ /*1582*/;
assign _13805_ = ~Q[1] /*1581*/;
assign _13804_ = _13805_ & D[23] /*1580*/;
assign _13807_ = _13432_ & _13804_ /*1575*/;
assign _13808_ = _13432_ ^ _13804_ /*1578*/;
assign _13809_ = _13800_ & _13808_ /*1576*/;
assign _13656_ = _13800_ ^ _13808_ /*1577*/;
assign _13806_ = _13807_ | _13809_ /*1574*/;
assign _13811_ = ~Q[1] /*1573*/;
assign _13810_ = _13811_ & D[24] /*1572*/;
assign _13813_ = _13433_ & _13810_ /*1567*/;
assign _13814_ = _13433_ ^ _13810_ /*1570*/;
assign _13815_ = _13806_ & _13814_ /*1568*/;
assign _13657_ = _13806_ ^ _13814_ /*1569*/;
assign _13812_ = _13813_ | _13815_ /*1566*/;
assign _13817_ = ~Q[1] /*1565*/;
assign _13816_ = _13817_ & D[25] /*1564*/;
assign _13819_ = _13434_ & _13816_ /*1559*/;
assign _13820_ = _13434_ ^ _13816_ /*1562*/;
assign _13821_ = _13812_ & _13820_ /*1560*/;
assign _13658_ = _13812_ ^ _13820_ /*1561*/;
assign _13818_ = _13819_ | _13821_ /*1558*/;
assign _13823_ = ~Q[1] /*1557*/;
assign _13822_ = _13823_ & D[26] /*1556*/;
assign _13825_ = _13435_ & _13822_ /*1551*/;
assign _13826_ = _13435_ ^ _13822_ /*1554*/;
assign _13827_ = _13818_ & _13826_ /*1552*/;
assign _13659_ = _13818_ ^ _13826_ /*1553*/;
assign _13824_ = _13825_ | _13827_ /*1550*/;
assign _13829_ = ~Q[1] /*1549*/;
assign _13828_ = _13829_ & D[27] /*1548*/;
assign _13831_ = _13436_ & _13828_ /*1543*/;
assign _13832_ = _13436_ ^ _13828_ /*1546*/;
assign _13833_ = _13824_ & _13832_ /*1544*/;
assign _13660_ = _13824_ ^ _13832_ /*1545*/;
assign _13830_ = _13831_ | _13833_ /*1542*/;
assign _13835_ = ~Q[1] /*1541*/;
assign _13834_ = _13835_ & D[28] /*1540*/;
assign _13837_ = _13437_ & _13834_ /*1535*/;
assign _13838_ = _13437_ ^ _13834_ /*1538*/;
assign _13839_ = _13830_ & _13838_ /*1536*/;
assign _13661_ = _13830_ ^ _13838_ /*1537*/;
assign _13836_ = _13837_ | _13839_ /*1534*/;
assign _13841_ = ~Q[1] /*1533*/;
assign _13840_ = _13841_ & D[29] /*1532*/;
assign _13843_ = _13438_ & _13840_ /*1527*/;
assign _13844_ = _13438_ ^ _13840_ /*1530*/;
assign _13845_ = _13836_ & _13844_ /*1528*/;
assign _13662_ = _13836_ ^ _13844_ /*1529*/;
assign _13842_ = _13843_ | _13845_ /*1526*/;
assign _13847_ = ~Q[1] /*1525*/;
assign _13846_ = _13847_ & D[30] /*1524*/;
assign _13849_ = _13439_ & _13846_ /*1519*/;
assign _13850_ = _13439_ ^ _13846_ /*1522*/;
assign _13851_ = _13842_ & _13850_ /*1520*/;
assign _13663_ = _13842_ ^ _13850_ /*1521*/;
assign _13848_ = _13849_ | _13851_ /*1518*/;
assign _13853_ = ~Q[1] /*1517*/;
assign _13852_ = _13853_ & zeroWire /*1516*/;
assign _13854_ = _13440_ ^ _13852_ /*1514*/;
assign _13664_ = _13854_ ^ _13848_ /*1513*/;
assign _13893_ = ~D[0] /*1387*/;
assign _13890_ = R_0[0] & _13893_ /*1383*/;
assign _13891_ = R_0[0] ^ _13893_ /*1386*/;
assign _13892_ = oneWire & _13891_ /*1384*/;
assign _13857_ = oneWire ^ _13891_ /*1385*/;
assign _13889_ = _13890_ | _13892_ /*1382*/;
assign _13898_ = ~D[1] /*1381*/;
assign _13895_ = _13633_ & _13898_ /*1377*/;
assign _13896_ = _13633_ ^ _13898_ /*1380*/;
assign _13897_ = _13889_ & _13896_ /*1378*/;
assign _13858_ = _13889_ ^ _13896_ /*1379*/;
assign _13894_ = _13895_ | _13897_ /*1376*/;
assign _13903_ = ~D[2] /*1375*/;
assign _13900_ = _13634_ & _13903_ /*1371*/;
assign _13901_ = _13634_ ^ _13903_ /*1374*/;
assign _13902_ = _13894_ & _13901_ /*1372*/;
assign _13859_ = _13894_ ^ _13901_ /*1373*/;
assign _13899_ = _13900_ | _13902_ /*1370*/;
assign _13908_ = ~D[3] /*1369*/;
assign _13905_ = _13635_ & _13908_ /*1365*/;
assign _13906_ = _13635_ ^ _13908_ /*1368*/;
assign _13907_ = _13899_ & _13906_ /*1366*/;
assign _13860_ = _13899_ ^ _13906_ /*1367*/;
assign _13904_ = _13905_ | _13907_ /*1364*/;
assign _13913_ = ~D[4] /*1363*/;
assign _13910_ = _13636_ & _13913_ /*1359*/;
assign _13911_ = _13636_ ^ _13913_ /*1362*/;
assign _13912_ = _13904_ & _13911_ /*1360*/;
assign _13861_ = _13904_ ^ _13911_ /*1361*/;
assign _13909_ = _13910_ | _13912_ /*1358*/;
assign _13918_ = ~D[5] /*1357*/;
assign _13915_ = _13637_ & _13918_ /*1353*/;
assign _13916_ = _13637_ ^ _13918_ /*1356*/;
assign _13917_ = _13909_ & _13916_ /*1354*/;
assign _13862_ = _13909_ ^ _13916_ /*1355*/;
assign _13914_ = _13915_ | _13917_ /*1352*/;
assign _13923_ = ~D[6] /*1351*/;
assign _13920_ = _13638_ & _13923_ /*1347*/;
assign _13921_ = _13638_ ^ _13923_ /*1350*/;
assign _13922_ = _13914_ & _13921_ /*1348*/;
assign _13863_ = _13914_ ^ _13921_ /*1349*/;
assign _13919_ = _13920_ | _13922_ /*1346*/;
assign _13928_ = ~D[7] /*1345*/;
assign _13925_ = _13639_ & _13928_ /*1341*/;
assign _13926_ = _13639_ ^ _13928_ /*1344*/;
assign _13927_ = _13919_ & _13926_ /*1342*/;
assign _13864_ = _13919_ ^ _13926_ /*1343*/;
assign _13924_ = _13925_ | _13927_ /*1340*/;
assign _13933_ = ~D[8] /*1339*/;
assign _13930_ = _13640_ & _13933_ /*1335*/;
assign _13931_ = _13640_ ^ _13933_ /*1338*/;
assign _13932_ = _13924_ & _13931_ /*1336*/;
assign _13865_ = _13924_ ^ _13931_ /*1337*/;
assign _13929_ = _13930_ | _13932_ /*1334*/;
assign _13938_ = ~D[9] /*1333*/;
assign _13935_ = _13641_ & _13938_ /*1329*/;
assign _13936_ = _13641_ ^ _13938_ /*1332*/;
assign _13937_ = _13929_ & _13936_ /*1330*/;
assign _13866_ = _13929_ ^ _13936_ /*1331*/;
assign _13934_ = _13935_ | _13937_ /*1328*/;
assign _13943_ = ~D[10] /*1327*/;
assign _13940_ = _13642_ & _13943_ /*1323*/;
assign _13941_ = _13642_ ^ _13943_ /*1326*/;
assign _13942_ = _13934_ & _13941_ /*1324*/;
assign _13867_ = _13934_ ^ _13941_ /*1325*/;
assign _13939_ = _13940_ | _13942_ /*1322*/;
assign _13948_ = ~D[11] /*1321*/;
assign _13945_ = _13643_ & _13948_ /*1317*/;
assign _13946_ = _13643_ ^ _13948_ /*1320*/;
assign _13947_ = _13939_ & _13946_ /*1318*/;
assign _13868_ = _13939_ ^ _13946_ /*1319*/;
assign _13944_ = _13945_ | _13947_ /*1316*/;
assign _13953_ = ~D[12] /*1315*/;
assign _13950_ = _13644_ & _13953_ /*1311*/;
assign _13951_ = _13644_ ^ _13953_ /*1314*/;
assign _13952_ = _13944_ & _13951_ /*1312*/;
assign _13869_ = _13944_ ^ _13951_ /*1313*/;
assign _13949_ = _13950_ | _13952_ /*1310*/;
assign _13958_ = ~D[13] /*1309*/;
assign _13955_ = _13645_ & _13958_ /*1305*/;
assign _13956_ = _13645_ ^ _13958_ /*1308*/;
assign _13957_ = _13949_ & _13956_ /*1306*/;
assign _13870_ = _13949_ ^ _13956_ /*1307*/;
assign _13954_ = _13955_ | _13957_ /*1304*/;
assign _13963_ = ~D[14] /*1303*/;
assign _13960_ = _13646_ & _13963_ /*1299*/;
assign _13961_ = _13646_ ^ _13963_ /*1302*/;
assign _13962_ = _13954_ & _13961_ /*1300*/;
assign _13871_ = _13954_ ^ _13961_ /*1301*/;
assign _13959_ = _13960_ | _13962_ /*1298*/;
assign _13968_ = ~D[15] /*1297*/;
assign _13965_ = _13647_ & _13968_ /*1293*/;
assign _13966_ = _13647_ ^ _13968_ /*1296*/;
assign _13967_ = _13959_ & _13966_ /*1294*/;
assign _13872_ = _13959_ ^ _13966_ /*1295*/;
assign _13964_ = _13965_ | _13967_ /*1292*/;
assign _13973_ = ~D[16] /*1291*/;
assign _13970_ = _13648_ & _13973_ /*1287*/;
assign _13971_ = _13648_ ^ _13973_ /*1290*/;
assign _13972_ = _13964_ & _13971_ /*1288*/;
assign _13873_ = _13964_ ^ _13971_ /*1289*/;
assign _13969_ = _13970_ | _13972_ /*1286*/;
assign _13978_ = ~D[17] /*1285*/;
assign _13975_ = _13649_ & _13978_ /*1281*/;
assign _13976_ = _13649_ ^ _13978_ /*1284*/;
assign _13977_ = _13969_ & _13976_ /*1282*/;
assign _13874_ = _13969_ ^ _13976_ /*1283*/;
assign _13974_ = _13975_ | _13977_ /*1280*/;
assign _13983_ = ~D[18] /*1279*/;
assign _13980_ = _13650_ & _13983_ /*1275*/;
assign _13981_ = _13650_ ^ _13983_ /*1278*/;
assign _13982_ = _13974_ & _13981_ /*1276*/;
assign _13875_ = _13974_ ^ _13981_ /*1277*/;
assign _13979_ = _13980_ | _13982_ /*1274*/;
assign _13988_ = ~D[19] /*1273*/;
assign _13985_ = _13651_ & _13988_ /*1269*/;
assign _13986_ = _13651_ ^ _13988_ /*1272*/;
assign _13987_ = _13979_ & _13986_ /*1270*/;
assign _13876_ = _13979_ ^ _13986_ /*1271*/;
assign _13984_ = _13985_ | _13987_ /*1268*/;
assign _13993_ = ~D[20] /*1267*/;
assign _13990_ = _13652_ & _13993_ /*1263*/;
assign _13991_ = _13652_ ^ _13993_ /*1266*/;
assign _13992_ = _13984_ & _13991_ /*1264*/;
assign _13877_ = _13984_ ^ _13991_ /*1265*/;
assign _13989_ = _13990_ | _13992_ /*1262*/;
assign _13998_ = ~D[21] /*1261*/;
assign _13995_ = _13653_ & _13998_ /*1257*/;
assign _13996_ = _13653_ ^ _13998_ /*1260*/;
assign _13997_ = _13989_ & _13996_ /*1258*/;
assign _13878_ = _13989_ ^ _13996_ /*1259*/;
assign _13994_ = _13995_ | _13997_ /*1256*/;
assign _14003_ = ~D[22] /*1255*/;
assign _14000_ = _13654_ & _14003_ /*1251*/;
assign _14001_ = _13654_ ^ _14003_ /*1254*/;
assign _14002_ = _13994_ & _14001_ /*1252*/;
assign _13879_ = _13994_ ^ _14001_ /*1253*/;
assign _13999_ = _14000_ | _14002_ /*1250*/;
assign _14008_ = ~D[23] /*1249*/;
assign _14005_ = _13655_ & _14008_ /*1245*/;
assign _14006_ = _13655_ ^ _14008_ /*1248*/;
assign _14007_ = _13999_ & _14006_ /*1246*/;
assign _13880_ = _13999_ ^ _14006_ /*1247*/;
assign _14004_ = _14005_ | _14007_ /*1244*/;
assign _14013_ = ~D[24] /*1243*/;
assign _14010_ = _13656_ & _14013_ /*1239*/;
assign _14011_ = _13656_ ^ _14013_ /*1242*/;
assign _14012_ = _14004_ & _14011_ /*1240*/;
assign _13881_ = _14004_ ^ _14011_ /*1241*/;
assign _14009_ = _14010_ | _14012_ /*1238*/;
assign _14018_ = ~D[25] /*1237*/;
assign _14015_ = _13657_ & _14018_ /*1233*/;
assign _14016_ = _13657_ ^ _14018_ /*1236*/;
assign _14017_ = _14009_ & _14016_ /*1234*/;
assign _13882_ = _14009_ ^ _14016_ /*1235*/;
assign _14014_ = _14015_ | _14017_ /*1232*/;
assign _14023_ = ~D[26] /*1231*/;
assign _14020_ = _13658_ & _14023_ /*1227*/;
assign _14021_ = _13658_ ^ _14023_ /*1230*/;
assign _14022_ = _14014_ & _14021_ /*1228*/;
assign _13883_ = _14014_ ^ _14021_ /*1229*/;
assign _14019_ = _14020_ | _14022_ /*1226*/;
assign _14028_ = ~D[27] /*1225*/;
assign _14025_ = _13659_ & _14028_ /*1221*/;
assign _14026_ = _13659_ ^ _14028_ /*1224*/;
assign _14027_ = _14019_ & _14026_ /*1222*/;
assign _13884_ = _14019_ ^ _14026_ /*1223*/;
assign _14024_ = _14025_ | _14027_ /*1220*/;
assign _14033_ = ~D[28] /*1219*/;
assign _14030_ = _13660_ & _14033_ /*1215*/;
assign _14031_ = _13660_ ^ _14033_ /*1218*/;
assign _14032_ = _14024_ & _14031_ /*1216*/;
assign _13885_ = _14024_ ^ _14031_ /*1217*/;
assign _14029_ = _14030_ | _14032_ /*1214*/;
assign _14038_ = ~D[29] /*1213*/;
assign _14035_ = _13661_ & _14038_ /*1209*/;
assign _14036_ = _13661_ ^ _14038_ /*1212*/;
assign _14037_ = _14029_ & _14036_ /*1210*/;
assign _13886_ = _14029_ ^ _14036_ /*1211*/;
assign _14034_ = _14035_ | _14037_ /*1208*/;
assign _14043_ = ~D[30] /*1207*/;
assign _14040_ = _13662_ & _14043_ /*1203*/;
assign _14041_ = _13662_ ^ _14043_ /*1206*/;
assign _14042_ = _14034_ & _14041_ /*1204*/;
assign _13887_ = _14034_ ^ _14041_ /*1205*/;
assign _14039_ = _14040_ | _14042_ /*1202*/;
assign _14044_ = _13663_ & oneWire /*1197*/;
assign _14045_ = _13663_ ^ oneWire /*1200*/;
assign _14046_ = _14039_ & _14045_ /*1198*/;
assign _13888_ = _14039_ ^ _14045_ /*1199*/;
assign Q[0] = _14044_ | _14046_ /*1196*/;
assign _14115_ = ~Q[0] /*1003*/;
assign _14114_ = _14115_ & D[0] /*1002*/;
assign _14117_ = _13857_ & _14114_ /*997*/;
assign _14118_ = _13857_ ^ _14114_ /*1000*/;
assign _14119_ = zeroWire & _14118_ /*998*/;
assign R_n1[0] = zeroWire ^ _14118_ /*999*/;
assign _14116_ = _14117_ | _14119_ /*996*/;
assign _14121_ = ~Q[0] /*995*/;
assign _14120_ = _14121_ & D[1] /*994*/;
assign _14123_ = _13858_ & _14120_ /*989*/;
assign _14124_ = _13858_ ^ _14120_ /*992*/;
assign _14125_ = _14116_ & _14124_ /*990*/;
assign R_n1[1] = _14116_ ^ _14124_ /*991*/;
assign _14122_ = _14123_ | _14125_ /*988*/;
assign _14127_ = ~Q[0] /*987*/;
assign _14126_ = _14127_ & D[2] /*986*/;
assign _14129_ = _13859_ & _14126_ /*981*/;
assign _14130_ = _13859_ ^ _14126_ /*984*/;
assign _14131_ = _14122_ & _14130_ /*982*/;
assign R_n1[2] = _14122_ ^ _14130_ /*983*/;
assign _14128_ = _14129_ | _14131_ /*980*/;
assign _14133_ = ~Q[0] /*979*/;
assign _14132_ = _14133_ & D[3] /*978*/;
assign _14135_ = _13860_ & _14132_ /*973*/;
assign _14136_ = _13860_ ^ _14132_ /*976*/;
assign _14137_ = _14128_ & _14136_ /*974*/;
assign R_n1[3] = _14128_ ^ _14136_ /*975*/;
assign _14134_ = _14135_ | _14137_ /*972*/;
assign _14139_ = ~Q[0] /*971*/;
assign _14138_ = _14139_ & D[4] /*970*/;
assign _14141_ = _13861_ & _14138_ /*965*/;
assign _14142_ = _13861_ ^ _14138_ /*968*/;
assign _14143_ = _14134_ & _14142_ /*966*/;
assign R_n1[4] = _14134_ ^ _14142_ /*967*/;
assign _14140_ = _14141_ | _14143_ /*964*/;
assign _14145_ = ~Q[0] /*963*/;
assign _14144_ = _14145_ & D[5] /*962*/;
assign _14147_ = _13862_ & _14144_ /*957*/;
assign _14148_ = _13862_ ^ _14144_ /*960*/;
assign _14149_ = _14140_ & _14148_ /*958*/;
assign R_n1[5] = _14140_ ^ _14148_ /*959*/;
assign _14146_ = _14147_ | _14149_ /*956*/;
assign _14151_ = ~Q[0] /*955*/;
assign _14150_ = _14151_ & D[6] /*954*/;
assign _14153_ = _13863_ & _14150_ /*949*/;
assign _14154_ = _13863_ ^ _14150_ /*952*/;
assign _14155_ = _14146_ & _14154_ /*950*/;
assign R_n1[6] = _14146_ ^ _14154_ /*951*/;
assign _14152_ = _14153_ | _14155_ /*948*/;
assign _14157_ = ~Q[0] /*947*/;
assign _14156_ = _14157_ & D[7] /*946*/;
assign _14159_ = _13864_ & _14156_ /*941*/;
assign _14160_ = _13864_ ^ _14156_ /*944*/;
assign _14161_ = _14152_ & _14160_ /*942*/;
assign R_n1[7] = _14152_ ^ _14160_ /*943*/;
assign _14158_ = _14159_ | _14161_ /*940*/;
assign _14163_ = ~Q[0] /*939*/;
assign _14162_ = _14163_ & D[8] /*938*/;
assign _14165_ = _13865_ & _14162_ /*933*/;
assign _14166_ = _13865_ ^ _14162_ /*936*/;
assign _14167_ = _14158_ & _14166_ /*934*/;
assign R_n1[8] = _14158_ ^ _14166_ /*935*/;
assign _14164_ = _14165_ | _14167_ /*932*/;
assign _14169_ = ~Q[0] /*931*/;
assign _14168_ = _14169_ & D[9] /*930*/;
assign _14171_ = _13866_ & _14168_ /*925*/;
assign _14172_ = _13866_ ^ _14168_ /*928*/;
assign _14173_ = _14164_ & _14172_ /*926*/;
assign R_n1[9] = _14164_ ^ _14172_ /*927*/;
assign _14170_ = _14171_ | _14173_ /*924*/;
assign _14175_ = ~Q[0] /*923*/;
assign _14174_ = _14175_ & D[10] /*922*/;
assign _14177_ = _13867_ & _14174_ /*917*/;
assign _14178_ = _13867_ ^ _14174_ /*920*/;
assign _14179_ = _14170_ & _14178_ /*918*/;
assign R_n1[10] = _14170_ ^ _14178_ /*919*/;
assign _14176_ = _14177_ | _14179_ /*916*/;
assign _14181_ = ~Q[0] /*915*/;
assign _14180_ = _14181_ & D[11] /*914*/;
assign _14183_ = _13868_ & _14180_ /*909*/;
assign _14184_ = _13868_ ^ _14180_ /*912*/;
assign _14185_ = _14176_ & _14184_ /*910*/;
assign R_n1[11] = _14176_ ^ _14184_ /*911*/;
assign _14182_ = _14183_ | _14185_ /*908*/;
assign _14187_ = ~Q[0] /*907*/;
assign _14186_ = _14187_ & D[12] /*906*/;
assign _14189_ = _13869_ & _14186_ /*901*/;
assign _14190_ = _13869_ ^ _14186_ /*904*/;
assign _14191_ = _14182_ & _14190_ /*902*/;
assign R_n1[12] = _14182_ ^ _14190_ /*903*/;
assign _14188_ = _14189_ | _14191_ /*900*/;
assign _14193_ = ~Q[0] /*899*/;
assign _14192_ = _14193_ & D[13] /*898*/;
assign _14195_ = _13870_ & _14192_ /*893*/;
assign _14196_ = _13870_ ^ _14192_ /*896*/;
assign _14197_ = _14188_ & _14196_ /*894*/;
assign R_n1[13] = _14188_ ^ _14196_ /*895*/;
assign _14194_ = _14195_ | _14197_ /*892*/;
assign _14199_ = ~Q[0] /*891*/;
assign _14198_ = _14199_ & D[14] /*890*/;
assign _14201_ = _13871_ & _14198_ /*885*/;
assign _14202_ = _13871_ ^ _14198_ /*888*/;
assign _14203_ = _14194_ & _14202_ /*886*/;
assign R_n1[14] = _14194_ ^ _14202_ /*887*/;
assign _14200_ = _14201_ | _14203_ /*884*/;
assign _14205_ = ~Q[0] /*883*/;
assign _14204_ = _14205_ & D[15] /*882*/;
assign _14207_ = _13872_ & _14204_ /*877*/;
assign _14208_ = _13872_ ^ _14204_ /*880*/;
assign _14209_ = _14200_ & _14208_ /*878*/;
assign R_n1[15] = _14200_ ^ _14208_ /*879*/;
assign _14206_ = _14207_ | _14209_ /*876*/;
assign _14211_ = ~Q[0] /*875*/;
assign _14210_ = _14211_ & D[16] /*874*/;
assign _14213_ = _13873_ & _14210_ /*869*/;
assign _14214_ = _13873_ ^ _14210_ /*872*/;
assign _14215_ = _14206_ & _14214_ /*870*/;
assign R_n1[16] = _14206_ ^ _14214_ /*871*/;
assign _14212_ = _14213_ | _14215_ /*868*/;
assign _14217_ = ~Q[0] /*867*/;
assign _14216_ = _14217_ & D[17] /*866*/;
assign _14219_ = _13874_ & _14216_ /*861*/;
assign _14220_ = _13874_ ^ _14216_ /*864*/;
assign _14221_ = _14212_ & _14220_ /*862*/;
assign R_n1[17] = _14212_ ^ _14220_ /*863*/;
assign _14218_ = _14219_ | _14221_ /*860*/;
assign _14223_ = ~Q[0] /*859*/;
assign _14222_ = _14223_ & D[18] /*858*/;
assign _14225_ = _13875_ & _14222_ /*853*/;
assign _14226_ = _13875_ ^ _14222_ /*856*/;
assign _14227_ = _14218_ & _14226_ /*854*/;
assign R_n1[18] = _14218_ ^ _14226_ /*855*/;
assign _14224_ = _14225_ | _14227_ /*852*/;
assign _14229_ = ~Q[0] /*851*/;
assign _14228_ = _14229_ & D[19] /*850*/;
assign _14231_ = _13876_ & _14228_ /*845*/;
assign _14232_ = _13876_ ^ _14228_ /*848*/;
assign _14233_ = _14224_ & _14232_ /*846*/;
assign R_n1[19] = _14224_ ^ _14232_ /*847*/;
assign _14230_ = _14231_ | _14233_ /*844*/;
assign _14235_ = ~Q[0] /*843*/;
assign _14234_ = _14235_ & D[20] /*842*/;
assign _14237_ = _13877_ & _14234_ /*837*/;
assign _14238_ = _13877_ ^ _14234_ /*840*/;
assign _14239_ = _14230_ & _14238_ /*838*/;
assign R_n1[20] = _14230_ ^ _14238_ /*839*/;
assign _14236_ = _14237_ | _14239_ /*836*/;
assign _14241_ = ~Q[0] /*835*/;
assign _14240_ = _14241_ & D[21] /*834*/;
assign _14243_ = _13878_ & _14240_ /*829*/;
assign _14244_ = _13878_ ^ _14240_ /*832*/;
assign _14245_ = _14236_ & _14244_ /*830*/;
assign R_n1[21] = _14236_ ^ _14244_ /*831*/;
assign _14242_ = _14243_ | _14245_ /*828*/;
assign _14247_ = ~Q[0] /*827*/;
assign _14246_ = _14247_ & D[22] /*826*/;
assign _14249_ = _13879_ & _14246_ /*821*/;
assign _14250_ = _13879_ ^ _14246_ /*824*/;
assign _14251_ = _14242_ & _14250_ /*822*/;
assign R_n1[22] = _14242_ ^ _14250_ /*823*/;
assign _14248_ = _14249_ | _14251_ /*820*/;
assign _14253_ = ~Q[0] /*819*/;
assign _14252_ = _14253_ & D[23] /*818*/;
assign _14255_ = _13880_ & _14252_ /*813*/;
assign _14256_ = _13880_ ^ _14252_ /*816*/;
assign _14257_ = _14248_ & _14256_ /*814*/;
assign R_n1[23] = _14248_ ^ _14256_ /*815*/;
assign _14254_ = _14255_ | _14257_ /*812*/;
assign _14259_ = ~Q[0] /*811*/;
assign _14258_ = _14259_ & D[24] /*810*/;
assign _14261_ = _13881_ & _14258_ /*805*/;
assign _14262_ = _13881_ ^ _14258_ /*808*/;
assign _14263_ = _14254_ & _14262_ /*806*/;
assign R_n1[24] = _14254_ ^ _14262_ /*807*/;
assign _14260_ = _14261_ | _14263_ /*804*/;
assign _14265_ = ~Q[0] /*803*/;
assign _14264_ = _14265_ & D[25] /*802*/;
assign _14267_ = _13882_ & _14264_ /*797*/;
assign _14268_ = _13882_ ^ _14264_ /*800*/;
assign _14269_ = _14260_ & _14268_ /*798*/;
assign R_n1[25] = _14260_ ^ _14268_ /*799*/;
assign _14266_ = _14267_ | _14269_ /*796*/;
assign _14271_ = ~Q[0] /*795*/;
assign _14270_ = _14271_ & D[26] /*794*/;
assign _14273_ = _13883_ & _14270_ /*789*/;
assign _14274_ = _13883_ ^ _14270_ /*792*/;
assign _14275_ = _14266_ & _14274_ /*790*/;
assign R_n1[26] = _14266_ ^ _14274_ /*791*/;
assign _14272_ = _14273_ | _14275_ /*788*/;
assign _14277_ = ~Q[0] /*787*/;
assign _14276_ = _14277_ & D[27] /*786*/;
assign _14279_ = _13884_ & _14276_ /*781*/;
assign _14280_ = _13884_ ^ _14276_ /*784*/;
assign _14281_ = _14272_ & _14280_ /*782*/;
assign R_n1[27] = _14272_ ^ _14280_ /*783*/;
assign _14278_ = _14279_ | _14281_ /*780*/;
assign _14283_ = ~Q[0] /*779*/;
assign _14282_ = _14283_ & D[28] /*778*/;
assign _14285_ = _13885_ & _14282_ /*773*/;
assign _14286_ = _13885_ ^ _14282_ /*776*/;
assign _14287_ = _14278_ & _14286_ /*774*/;
assign R_n1[28] = _14278_ ^ _14286_ /*775*/;
assign _14284_ = _14285_ | _14287_ /*772*/;
assign _14289_ = ~Q[0] /*771*/;
assign _14288_ = _14289_ & D[29] /*770*/;
assign _14291_ = _13886_ & _14288_ /*765*/;
assign _14292_ = _13886_ ^ _14288_ /*768*/;
assign _14293_ = _14284_ & _14292_ /*766*/;
assign R_n1[29] = _14284_ ^ _14292_ /*767*/;
assign _14290_ = _14291_ | _14293_ /*764*/;
assign _14295_ = ~Q[0] /*763*/;
assign _14294_ = _14295_ & D[30] /*762*/;
assign _14297_ = _13887_ & _14294_ /*757*/;
assign _14298_ = _13887_ ^ _14294_ /*760*/;
assign _14299_ = _14290_ & _14298_ /*758*/;
assign R_n1[30] = _14290_ ^ _14298_ /*759*/;
assign _14296_ = _14297_ | _14299_ /*756*/;
endmodule
