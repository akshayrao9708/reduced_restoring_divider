module divider(q, rout, rin, div);
  wire _0_;
  wire _1_;
  wire _2_;
  wire _3_;
  wire _4_;
  wire _5_;
  wire _6_;
  wire _7_;
  wire _8_;
  wire _9_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  wire _38_;
  wire _39_;
  wire _40_;
  wire _41_;
  wire _42_;
  wire _43_;
  wire _44_;
  wire _45_;
  wire _46_;
  wire _47_;
  wire _48_;
  wire _49_;
  wire _50_;
  wire _51_;
  wire _52_;
  wire _53_;
  wire _54_;
  wire _55_;
  wire _56_;
  wire _57_;
  wire _58_;
  wire _59_;
  wire _60_;
  wire _61_;
  wire _62_;
  wire _63_;
  wire _64_;
  wire _65_;
  wire _66_;
  wire _67_;
  wire _68_;
  wire _69_;
  wire _70_;
  wire _71_;
  wire _72_;
  wire _73_;
  wire _74_;
  wire _75_;
  wire _76_;
  wire _77_;
  wire _78_;
  wire _79_;
  wire _80_;
  wire _81_;
  wire _82_;
  wire _83_;
  wire _84_;
  wire _85_;
  wire _86_;
  wire _87_;
  wire _88_;
  wire _89_;
  wire _90_;
  wire _91_;
  wire _92_;
  wire _93_;
  wire _94_;
  wire _95_;
  wire _96_;
  wire _97_;
  wire _98_;
  wire _99_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire _304_;
  wire _305_;
  wire _306_;
  wire _307_;
  wire _308_;
  wire _309_;
  wire _310_;
  wire _311_;
  wire _312_;
  wire _313_;
  wire _314_;
  wire _315_;
  wire _316_;
  wire _317_;
  wire _318_;
  wire _319_;
  wire _320_;
  wire _321_;
  wire _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire _326_;
  wire _327_;
  wire _328_;
  wire _329_;
  wire _330_;
  wire _331_;
  wire _332_;
  wire _333_;
  wire _334_;
  wire _335_;
  wire _336_;
  wire _337_;
  wire _338_;
  wire _339_;
  wire _340_;
  wire _341_;
  wire _342_;
  wire _343_;
  wire _344_;
  wire _345_;
  wire _346_;
  wire _347_;
  wire _348_;
  wire _349_;
  wire _350_;
  wire _351_;
  wire _352_;
  wire _353_;
  wire _354_;
  wire _355_;
  wire _356_;
  wire _357_;
  wire _358_;
  wire _359_;
  wire _360_;
  wire _361_;
  wire _362_;
  wire _363_;
  wire _364_;
  wire _365_;
  wire _366_;
  wire _367_;
  wire _368_;
  wire _369_;
  wire _370_;
  wire _371_;
  wire _372_;
  wire _373_;
  wire _374_;
  wire _375_;
  wire _376_;
  wire _377_;
  wire _378_;
  wire _379_;
  wire _380_;
  wire _381_;
  wire _382_;
  wire _383_;
  wire _384_;
  wire _385_;
  wire _386_;
  wire _387_;
  wire _388_;
  wire _389_;
  wire _390_;
  wire _391_;
  wire _392_;
  wire _393_;
  wire _394_;
  wire _395_;
  wire _396_;
  wire _397_;
  wire _398_;
  wire _399_;
  wire _400_;
  wire _401_;
  wire _402_;
  wire _403_;
  wire _404_;
  wire _405_;
  wire _406_;
  wire _407_;
  wire _408_;
  wire _409_;
  wire _410_;
  wire _411_;
  wire _412_;
  wire _413_;
  wire _414_;
  wire _415_;
  wire _416_;
  wire _417_;
  wire _418_;
  wire _419_;
  wire _420_;
  wire _421_;
  wire _422_;
  wire _423_;
  wire _424_;
  wire _425_;
  wire _426_;
  wire _427_;
  wire _428_;
  wire _429_;
  wire _430_;
  wire _431_;
  wire _432_;
  wire _433_;
  wire _434_;
  wire _435_;
  wire _436_;
  wire _437_;
  wire _438_;
  wire _439_;
  wire _440_;
  wire _441_;
  wire _442_;
  wire _443_;
  wire _444_;
  wire _445_;
  wire _446_;
  wire _447_;
  wire _448_;
  wire _449_;
  wire _450_;
  wire _451_;
  wire _452_;
  wire _453_;
  wire _454_;
  wire _455_;
  wire _456_;
  wire _457_;
  wire _458_;
  wire _459_;
  wire _460_;
  wire _461_;
  wire _462_;
  wire _463_;
  wire _464_;
  wire _465_;
  wire _466_;
  wire _467_;
  wire _468_;
  wire _469_;
  wire _470_;
  wire _471_;
  wire _472_;
  wire _473_;
  wire _474_;
  wire _475_;
  wire _476_;
  wire _477_;
  wire _478_;
  wire _479_;
  wire _480_;
  wire _481_;
  wire _482_;
  wire _483_;
  wire _484_;
  wire _485_;
  wire _486_;
  wire _487_;
  wire _488_;
  wire _489_;
  wire _490_;
  wire _491_;
  wire _492_;
  wire _493_;
  wire _494_;
  wire _495_;
  wire _496_;
  wire _497_;
  wire _498_;
  wire _499_;
  wire _500_;
  wire _501_;
  wire _502_;
  wire _503_;
  wire _504_;
  wire _505_;
  wire _506_;
  wire _507_;
  wire _508_;
  wire _509_;
  wire _510_;
  wire _511_;
  wire _512_;
  wire _513_;
  wire _514_;
  wire _515_;
  wire _516_;
  wire _517_;
  wire _518_;
  wire _519_;
  wire _520_;
  wire _521_;
  wire _522_;
  wire _523_;
  wire _524_;
  wire _525_;
  wire _526_;
  wire _527_;
  wire _528_;
  wire _529_;
  wire _530_;
  wire _531_;
  wire _532_;
  wire _533_;
  wire _534_;
  wire _535_;
  wire _536_;
  wire _537_;
  wire _538_;
  wire _539_;
  wire _540_;
  wire _541_;
  wire _542_;
  wire _543_;
  wire _544_;
  wire _545_;
  wire _546_;
  wire _547_;
  wire _548_;
  wire _549_;
  wire _550_;
  wire _551_;
  wire _552_;
  wire _553_;
  wire _554_;
  wire _555_;
  wire _556_;
  wire _557_;
  wire _558_;
  wire _559_;
  wire _560_;
  wire _561_;
  wire _562_;
  wire _563_;
  wire _564_;
  wire _565_;
  wire _566_;
  wire _567_;
  wire _568_;
  wire _569_;
  wire _570_;
  wire _571_;
  wire _572_;
  wire _573_;
  wire _574_;
  wire _575_;
  wire _576_;
  wire _577_;
  wire _578_;
  wire _579_;
  wire _580_;
  wire _581_;
  wire _582_;
  wire _583_;
  wire _584_;
  wire _585_;
  wire _586_;
  wire _587_;
  wire _588_;
  wire _589_;
  wire _590_;
  wire _591_;
  wire _592_;
  wire _593_;
  wire _594_;
  wire _595_;
  wire _596_;
  wire _597_;
  wire _598_;
  wire _599_;
  wire _600_;
  wire _601_;
  wire _602_;
  wire _603_;
  wire _604_;
  wire _605_;
  wire _606_;
  wire _607_;
  wire _608_;
  wire _609_;
  wire _610_;
  wire _611_;
  wire _612_;
  wire _613_;
  wire _614_;
  wire _615_;
  wire _616_;
  wire _617_;
  wire _618_;
  wire _619_;
  wire _620_;
  wire _621_;
  wire _622_;
  wire _623_;
  wire _624_;
  wire _625_;
  wire _626_;
  wire _627_;
  wire _628_;
  wire _629_;
  wire _630_;
  wire _631_;
  wire _632_;
  wire _633_;
  wire _634_;
  wire _635_;
  wire _636_;
  wire _637_;
  wire _638_;
  wire _639_;
  wire _640_;
  wire _641_;
  wire _642_;
  wire _643_;
  wire _644_;
  wire _645_;
  wire _646_;
  wire _647_;
  wire _648_;
  wire _649_;
  wire _650_;
  wire _651_;
  wire _652_;
  wire _653_;
  wire _654_;
  wire _655_;
  wire _656_;
  wire _657_;
  wire _658_;
  wire _659_;
  wire _660_;
  wire _661_;
  wire _662_;
  wire _663_;
  wire _664_;
  wire _665_;
  wire _666_;
  wire _667_;
  wire _668_;
  wire _669_;
  wire _670_;
  wire _671_;
  wire _672_;
  wire _673_;
  wire _674_;
  wire _675_;
  wire _676_;
  wire _677_;
  wire _678_;
  wire _679_;
  wire _680_;
  wire _681_;
  wire _682_;
  wire _683_;
  wire _684_;
  wire _685_;
  wire _686_;
  wire _687_;
  wire _688_;
  wire _689_;
  wire _690_;
  wire _691_;
  wire _692_;
  wire _693_;
  wire _694_;
  wire _695_;
  wire _696_;
  wire _697_;
  wire _698_;
  wire _699_;
  wire _700_;
  wire _701_;
  wire _702_;
  wire _703_;
  wire _704_;
  wire _705_;
  wire _706_;
  wire _707_;
  wire _708_;
  wire _709_;
  wire _710_;
  wire _711_;
  wire _712_;
  wire _713_;
  wire _714_;
  wire _715_;
  wire _716_;
  wire _717_;
  wire _718_;
  wire _719_;
  wire _720_;
  wire _721_;
  wire _722_;
  wire _723_;
  wire _724_;
  wire _725_;
  wire _726_;
  wire _727_;
  wire _728_;
  wire _729_;
  wire _730_;
  wire _731_;
  wire _732_;
  wire _733_;
  wire _734_;
  wire _735_;
  wire _736_;
  wire _737_;
  wire _738_;
  wire _739_;
  wire _740_;
  wire _741_;
  wire _742_;
  wire _743_;
  wire _744_;
  wire _745_;
  wire _746_;
  wire _747_;
  wire _748_;
  wire _749_;
  wire _750_;
  wire _751_;
  wire _752_;
  wire _753_;
  wire _754_;
  wire _755_;
  wire _756_;
  wire _757_;
  wire _758_;
  wire _759_;
  wire _760_;
  wire _761_;
  wire _762_;
  wire _763_;
  wire _764_;
  wire _765_;
  wire _766_;
  wire _767_;
  wire _768_;
  wire _769_;
  wire _770_;
  wire _771_;
  wire _772_;
  wire _773_;
  wire _774_;
  wire _775_;
  wire _776_;
  wire _777_;
  wire _778_;
  wire _779_;
  wire _780_;
  wire _781_;
  wire _782_;
  wire _783_;
  wire _784_;
  wire _785_;
  wire _786_;
  wire _787_;
  wire _788_;
  wire _789_;
  wire _790_;
  wire _791_;
  wire _792_;
  wire _793_;
  wire _794_;
  wire _795_;
  wire _796_;
  wire _797_;
  wire _798_;
  wire _799_;
  wire _800_;
  wire _801_;
  wire _802_;
  wire _803_;
  wire _804_;
  wire _805_;
  wire _806_;
  wire _807_;
  wire _808_;
  wire _809_;
  wire _810_;
  wire _811_;
  wire _812_;
  wire _813_;
  wire _814_;
  wire _815_;
  wire _816_;
  wire _817_;
  wire _818_;
  wire _819_;
  wire _820_;
  wire _821_;
  wire _822_;
  wire _823_;
  wire _824_;
  wire _825_;
  wire _826_;
  wire _827_;
  wire _828_;
  wire _829_;
  wire _830_;
  wire _831_;
  wire _832_;
  wire _833_;
  wire _834_;
  wire _835_;
  wire _836_;
  wire _837_;
  wire _838_;
  wire _839_;
  wire _840_;
  wire _841_;
  wire _842_;
  wire _843_;
  wire _844_;
  wire _845_;
  wire _846_;
  wire _847_;
  wire _848_;
  wire _849_;
  wire _850_;
  wire _851_;
  wire _852_;
  wire _853_;
  wire _854_;
  wire _855_;
  wire _856_;
  wire _857_;
  wire _858_;
  wire _859_;
  wire _860_;
  wire _861_;
  wire _862_;
  wire _863_;
  wire _864_;
  wire _865_;
  wire _866_;
  wire _867_;
  wire _868_;
  wire _869_;
  wire _870_;
  wire _871_;
  wire _872_;
  wire _873_;
  wire _874_;
  wire _875_;
  wire _876_;
  wire _877_;
  wire _878_;
  wire _879_;
  wire _880_;
  wire _881_;
  wire _882_;
  wire _883_;
  wire _884_;
  wire _885_;
  wire _886_;
  wire _887_;
  wire _888_;
  wire _889_;
  wire _890_;
  wire _891_;
  wire _892_;
  wire _893_;
  wire _894_;
  wire _895_;
  wire _896_;
  wire _897_;
  wire _898_;
  wire _899_;
  wire _900_;
  wire _901_;
  wire _902_;
  wire _903_;
  wire _904_;
  wire _905_;
  wire _906_;
  wire _907_;
  wire _908_;
  wire _909_;
  wire _910_;
  wire _911_;
  wire _912_;
  wire _913_;
  wire _914_;
  wire _915_;
  wire _916_;
  wire _917_;
  wire _918_;
  wire _919_;
  wire _920_;
  wire _921_;
  wire _922_;
  wire _923_;
  wire _924_;
  wire _925_;
  wire _926_;
  wire _927_;
  wire _928_;
  wire _929_;
  wire _930_;
  wire _931_;
  wire _932_;
  wire _933_;
  wire _934_;
  wire _935_;
  wire _936_;
  wire _937_;
  wire _938_;
  wire _939_;
  wire _940_;
  wire _941_;
  wire _942_;
  wire _943_;
  wire _944_;
  wire _945_;
  wire _946_;
  wire _947_;
  wire _948_;
  wire _949_;
  wire _950_;
  wire _951_;
  wire _952_;
  wire _953_;
  wire _954_;
  wire _955_;
  wire _956_;
  wire _957_;
  wire _958_;
  wire _959_;
  wire _960_;
  wire _961_;
  wire _962_;
  wire _963_;
  wire _964_;
  wire _965_;
  wire _966_;
  wire _967_;
  wire _968_;
  wire _969_;
  wire _970_;
  wire _971_;
  wire _972_;
  wire _973_;
  wire _974_;
  wire _975_;
  wire _976_;
  wire _977_;
  wire _978_;
  wire _979_;
  wire _980_;
  wire _981_;
  wire _982_;
  wire _983_;
  wire _984_;
  wire _985_;
  wire _986_;
  wire _987_;
  wire _988_;
  wire _989_;
  wire _990_;
  wire _991_;
  wire _992_;
  wire _993_;
  wire _994_;
  wire _995_;
  wire _996_;
  wire _997_;
  wire _998_;
  wire _999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire _1601_;
  wire _1602_;
  wire _1603_;
  wire _1604_;
  wire _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire _1611_;
  wire _1612_;
  wire _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire _1629_;
  wire _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire _1720_;
  wire _1721_;
  wire _1722_;
  wire _1723_;
  wire _1724_;
  wire _1725_;
  wire _1726_;
  wire _1727_;
  wire _1728_;
  wire _1729_;
  wire _1730_;
  wire _1731_;
  wire _1732_;
  wire _1733_;
  wire _1734_;
  wire _1735_;
  wire _1736_;
  wire _1737_;
  wire _1738_;
  wire _1739_;
  wire _1740_;
  wire _1741_;
  wire _1742_;
  wire _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire _1751_;
  wire _1752_;
  wire _1753_;
  wire _1754_;
  wire _1755_;
  wire _1756_;
  wire _1757_;
  wire _1758_;
  wire _1759_;
  wire _1760_;
  wire _1761_;
  wire _1762_;
  wire _1763_;
  wire _1764_;
  wire _1765_;
  wire _1766_;
  wire _1767_;
  wire _1768_;
  wire _1769_;
  wire _1770_;
  wire _1771_;
  wire _1772_;
  wire _1773_;
  wire _1774_;
  wire _1775_;
  wire _1776_;
  wire _1777_;
  wire _1778_;
  wire _1779_;
  wire _1780_;
  wire _1781_;
  wire _1782_;
  wire _1783_;
  wire _1784_;
  wire _1785_;
  wire _1786_;
  wire _1787_;
  wire _1788_;
  wire _1789_;
  wire _1790_;
  wire _1791_;
  wire [30:0] r_0;
  wire [30:0] r_1;
  wire [15:0] m_1;
  wire [15:0] sum_1;
  wire [15:0] inv_1;
  wire [29:0] r_2;
  wire [15:0] m_2;
  wire [15:0] sum_2;
  wire [15:0] inv_2;
  wire [28:0] r_3;
  wire [15:0] m_3;
  wire [15:0] sum_3;
  wire [15:0] inv_3;
  wire [27:0] r_4;
  wire [15:0] m_4;
  wire [15:0] sum_4;
  wire [15:0] inv_4;
  wire [26:0] r_5;
  wire [15:0] m_5;
  wire [15:0] sum_5;
  wire [15:0] inv_5;
  wire [25:0] r_6;
  wire [15:0] m_6;
  wire [15:0] sum_6;
  wire [15:0] inv_6;
  wire [24:0] r_7;
  wire [15:0] m_7;
  wire [15:0] sum_7;
  wire [15:0] inv_7;
  wire [23:0] r_8;
  wire [15:0] m_8;
  wire [15:0] sum_8;
  wire [15:0] inv_8;
  wire [22:0] r_9;
  wire [15:0] m_9;
  wire [15:0] sum_9;
  wire [15:0] inv_9;
  wire [21:0] r_10;
  wire [15:0] m_10;
  wire [15:0] sum_10;
  wire [15:0] inv_10;
  wire [20:0] r_11;
  wire [15:0] m_11;
  wire [15:0] sum_11;
  wire [15:0] inv_11;
  wire [19:0] r_12;
  wire [15:0] m_12;
  wire [15:0] sum_12;
  wire [15:0] inv_12;
  wire [18:0] r_13;
  wire [15:0] m_13;
  wire [15:0] sum_13;
  wire [15:0] inv_13;
  wire [17:0] r_14;
  wire [15:0] m_14;
  wire [15:0] sum_14;
  wire [15:0] inv_14;
  wire [16:0] r_15;
  wire [15:0] m_15;
  wire [15:0] sum_15;
  wire [15:0] inv_15;
  wire [15:0] r_16;
  wire [15:0] m_16;
  wire [15:0] sum_16;
  wire [15:0] inv_16;
  wire zeroWire;
  wire oneWire;
  input [29:0] rin;
  input [14:0] div;
  output [15:0] q;
  output [15:0] rout;
  assign zeroWire = 1'b0 /*0*/;
  assign oneWire = 1'b1 /*0*/;
  assign r_0[0] = rin[0] /*6519*/;
  assign r_0[1] = rin[1] /*6518*/;
  assign r_0[2] = rin[2] /*6517*/;
  assign r_0[3] = rin[3] /*6516*/;
  assign r_0[4] = rin[4] /*6515*/;
  assign r_0[5] = rin[5] /*6514*/;
  assign r_0[6] = rin[6] /*6513*/;
  assign r_0[7] = rin[7] /*6512*/;
  assign r_0[8] = rin[8] /*6511*/;
  assign r_0[9] = rin[9] /*6510*/;
  assign r_0[10] = rin[10] /*6509*/;
  assign r_0[11] = rin[11] /*6508*/;
  assign r_0[12] = rin[12] /*6507*/;
  assign r_0[13] = rin[13] /*6506*/;
  assign r_0[14] = rin[14] /*6505*/;
  assign r_0[15] = rin[15] /*6504*/;
  assign r_0[16] = rin[16] /*6503*/;
  assign r_0[17] = rin[17] /*6502*/;
  assign r_0[18] = rin[18] /*6501*/;
  assign r_0[19] = rin[19] /*6500*/;
  assign r_0[20] = rin[20] /*6499*/;
  assign r_0[21] = rin[21] /*6498*/;
  assign r_0[22] = rin[22] /*6497*/;
  assign r_0[23] = rin[23] /*6496*/;
  assign r_0[24] = rin[24] /*6495*/;
  assign r_0[25] = rin[25] /*6494*/;
  assign r_0[26] = rin[26] /*6493*/;
  assign r_0[27] = rin[27] /*6492*/;
  assign r_0[28] = rin[28] /*6491*/;
  assign r_0[29] = rin[29] /*6490*/;
  assign r_0[30] = zeroWire /*6489*/;
  assign inv_1[0] = ~div[0] /*6488*/;
  assign inv_1[1] = ~div[1] /*6487*/;
  assign inv_1[2] = ~div[2] /*6486*/;
  assign inv_1[3] = ~div[3] /*6485*/;
  assign inv_1[4] = ~div[4] /*6484*/;
  assign inv_1[5] = ~div[5] /*6483*/;
  assign inv_1[6] = ~div[6] /*6482*/;
  assign inv_1[7] = ~div[7] /*6481*/;
  assign inv_1[8] = ~div[8] /*6480*/;
  assign inv_1[9] = ~div[9] /*6479*/;
  assign inv_1[10] = ~div[10] /*6478*/;
  assign inv_1[11] = ~div[11] /*6477*/;
  assign inv_1[12] = ~div[12] /*6476*/;
  assign inv_1[13] = ~div[13] /*6475*/;
  assign inv_1[14] = ~div[14] /*6474*/;
assign inv_1[15] = oneWire /*6473*/;
  assign _0_ = inv_1[0] ^ r_0[15] /*6471*/;
  assign sum_1[0] = _0_ ^ oneWire /*6470*/;
  assign _1_ = _0_ & oneWire /*6469*/;
  assign _2_ = inv_1[0] & r_0[15] /*6468*/;
  assign _3_ = _1_ | _2_ /*6467*/;
  assign _4_ = inv_1[1] ^ r_0[16] /*6466*/;
  assign sum_1[1] = _4_ ^ _3_ /*6465*/;
  assign _5_ = _4_ & _3_ /*6464*/;
  assign _6_ = inv_1[1] & r_0[16] /*6463*/;
  assign _7_ = _5_ | _6_ /*6462*/;
  assign _8_ = inv_1[2] ^ r_0[17] /*6460*/;
  assign sum_1[2] = _8_ ^ _7_ /*6459*/;
  assign _9_ = _8_ & _7_ /*6458*/;
  assign _10_ = inv_1[2] & r_0[17] /*6457*/;
  assign _11_ = _9_ | _10_ /*6456*/;
  assign _12_ = inv_1[3] ^ r_0[18] /*6454*/;
  assign sum_1[3] = _12_ ^ _11_ /*6453*/;
  assign _13_ = _12_ & _11_ /*6452*/;
  assign _14_ = inv_1[3] & r_0[18] /*6451*/;
  assign _15_ = _13_ | _14_ /*6450*/;
  assign _16_ = inv_1[4] ^ r_0[19] /*6448*/;
  assign sum_1[4] = _16_ ^ _15_ /*6447*/;
  assign _17_ = _16_ & _15_ /*6446*/;
  assign _18_ = inv_1[4] & r_0[19] /*6445*/;
  assign _19_ = _17_ | _18_ /*6444*/;
  assign _20_ = inv_1[5] ^ r_0[20] /*6442*/;
  assign sum_1[5] = _20_ ^ _19_ /*6441*/;
  assign _21_ = _20_ & _19_ /*6440*/;
  assign _22_ = inv_1[5] & r_0[20] /*6439*/;
  assign _23_ = _21_ | _22_ /*6438*/;
  assign _24_ = inv_1[6] ^ r_0[21] /*6436*/;
  assign sum_1[6] = _24_ ^ _23_ /*6435*/;
  assign _25_ = _24_ & _23_ /*6434*/;
  assign _26_ = inv_1[6] & r_0[21] /*6433*/;
  assign _27_ = _25_ | _26_ /*6432*/;
  assign _28_ = inv_1[7] ^ r_0[22] /*6430*/;
  assign sum_1[7] = _28_ ^ _27_ /*6429*/;
  assign _29_ = _28_ & _27_ /*6428*/;
  assign _30_ = inv_1[7] & r_0[22] /*6427*/;
  assign _31_ = _29_ | _30_ /*6426*/;
  assign _32_ = inv_1[8] ^ r_0[23] /*6424*/;
  assign sum_1[8] = _32_ ^ _31_ /*6423*/;
  assign _33_ = _32_ & _31_ /*6422*/;
  assign _34_ = inv_1[8] & r_0[23] /*6421*/;
  assign _35_ = _33_ | _34_ /*6420*/;
  assign _36_ = inv_1[9] ^ r_0[24] /*6418*/;
  assign sum_1[9] = _36_ ^ _35_ /*6417*/;
  assign _37_ = _36_ & _35_ /*6416*/;
  assign _38_ = inv_1[9] & r_0[24] /*6415*/;
  assign _39_ = _37_ | _38_ /*6414*/;
  assign _40_ = inv_1[10] ^ r_0[25] /*6412*/;
  assign sum_1[10] = _40_ ^ _39_ /*6411*/;
  assign _41_ = _40_ & _39_ /*6410*/;
  assign _42_ = inv_1[10] & r_0[25] /*6409*/;
  assign _43_ = _41_ | _42_ /*6408*/;
  assign _44_ = inv_1[11] ^ r_0[26] /*6406*/;
  assign sum_1[11] = _44_ ^ _43_ /*6405*/;
  assign _45_ = _44_ & _43_ /*6404*/;
  assign _46_ = inv_1[11] & r_0[26] /*6403*/;
  assign _47_ = _45_ | _46_ /*6402*/;
  assign _48_ = inv_1[12] ^ r_0[27] /*6400*/;
  assign sum_1[12] = _48_ ^ _47_ /*6399*/;
  assign _49_ = _48_ & _47_ /*6398*/;
  assign _50_ = inv_1[12] & r_0[27] /*6397*/;
  assign _51_ = _49_ | _50_ /*6396*/;
  assign _52_ = inv_1[13] ^ r_0[28] /*6394*/;
  assign sum_1[13] = _52_ ^ _51_ /*6393*/;
  assign _53_ = _52_ & _51_ /*6392*/;
  assign _54_ = inv_1[13] & r_0[28] /*6391*/;
  assign _55_ = _53_ | _54_ /*6390*/;
  assign _56_ = inv_1[14] ^ r_0[29] /*6388*/;
  assign sum_1[14] = _56_ ^ _55_ /*6387*/;
  assign _57_ = _56_ & _55_ /*6386*/;
  assign _58_ = inv_1[14] & r_0[29] /*6385*/;
  assign _59_ = _57_ | _58_ /*6384*/;
  assign _60_ = inv_1[15] ^ r_0[30] /*6382*/;
  assign sum_1[15] = _60_ ^ _59_ /*6381*/;
  assign _61_ = _60_ & _59_ /*6380*/;
  assign _62_ = inv_1[15] & r_0[30] /*6379*/;
  assign _63_ = _61_ | _62_ /*6378*/;
  assign q[15] = ~sum_1[15] /*6389*/;
  assign m_1[0] = r_0[15] /*6388*/;
  assign m_1[1] = r_0[16] /*6387*/;
  assign m_1[2] = r_0[17] /*6386*/;
  assign m_1[3] = r_0[18] /*6385*/;
  assign m_1[4] = r_0[19] /*6384*/;
  assign m_1[5] = r_0[20] /*6383*/;
  assign m_1[6] = r_0[21] /*6382*/;
  assign m_1[7] = r_0[22] /*6381*/;
  assign m_1[8] = r_0[23] /*6380*/;
  assign m_1[9] = r_0[24] /*6379*/;
  assign m_1[10] = r_0[25] /*6378*/;
  assign m_1[11] = r_0[26] /*6377*/;
  assign m_1[12] = r_0[27] /*6376*/;
  assign m_1[13] = r_0[28] /*6375*/;
  assign m_1[14] = r_0[29] /*6374*/;
  assign m_1[15] = r_0[30] /*6373*/;
  assign _64_ = ~q[15] /*6371*/;
  assign _65_ = sum_1[0] & q[15] /*6370*/;
  assign _66_ = m_1[0] & _64_ /*6369*/;
  assign r_1[15] = _66_ | _65_ /*6368*/;
  assign _67_ = ~q[15] /*6367*/;
  assign _68_ = sum_1[1] & q[15] /*6366*/;
  assign _69_ = m_1[1] & _67_ /*6365*/;
  assign r_1[16] = _69_ | _68_ /*6364*/;
  assign _70_ = ~q[15] /*6363*/;
  assign _71_ = sum_1[2] & q[15] /*6362*/;
  assign _72_ = m_1[2] & _70_ /*6361*/;
  assign r_1[17] = _72_ | _71_ /*6360*/;
  assign _73_ = ~q[15] /*6359*/;
  assign _74_ = sum_1[3] & q[15] /*6358*/;
  assign _75_ = m_1[3] & _73_ /*6357*/;
  assign r_1[18] = _75_ | _74_ /*6356*/;
  assign _76_ = ~q[15] /*6355*/;
  assign _77_ = sum_1[4] & q[15] /*6354*/;
  assign _78_ = m_1[4] & _76_ /*6353*/;
  assign r_1[19] = _78_ | _77_ /*6352*/;
  assign _79_ = ~q[15] /*6351*/;
  assign _80_ = sum_1[5] & q[15] /*6350*/;
  assign _81_ = m_1[5] & _79_ /*6349*/;
  assign r_1[20] = _81_ | _80_ /*6348*/;
  assign _82_ = ~q[15] /*6347*/;
  assign _83_ = sum_1[6] & q[15] /*6346*/;
  assign _84_ = m_1[6] & _82_ /*6345*/;
  assign r_1[21] = _84_ | _83_ /*6344*/;
  assign _85_ = ~q[15] /*6343*/;
  assign _86_ = sum_1[7] & q[15] /*6342*/;
  assign _87_ = m_1[7] & _85_ /*6341*/;
  assign r_1[22] = _87_ | _86_ /*6340*/;
  assign _88_ = ~q[15] /*6339*/;
  assign _89_ = sum_1[8] & q[15] /*6338*/;
  assign _90_ = m_1[8] & _88_ /*6337*/;
  assign r_1[23] = _90_ | _89_ /*6336*/;
  assign _91_ = ~q[15] /*6335*/;
  assign _92_ = sum_1[9] & q[15] /*6334*/;
  assign _93_ = m_1[9] & _91_ /*6333*/;
  assign r_1[24] = _93_ | _92_ /*6332*/;
  assign _94_ = ~q[15] /*6331*/;
  assign _95_ = sum_1[10] & q[15] /*6330*/;
  assign _96_ = m_1[10] & _94_ /*6329*/;
  assign r_1[25] = _96_ | _95_ /*6328*/;
  assign _97_ = ~q[15] /*6327*/;
  assign _98_ = sum_1[11] & q[15] /*6326*/;
  assign _99_ = m_1[11] & _97_ /*6325*/;
  assign r_1[26] = _99_ | _98_ /*6324*/;
  assign _100_ = ~q[15] /*6323*/;
  assign _101_ = sum_1[12] & q[15] /*6322*/;
  assign _102_ = m_1[12] & _100_ /*6321*/;
  assign r_1[27] = _102_ | _101_ /*6320*/;
  assign _103_ = ~q[15] /*6319*/;
  assign _104_ = sum_1[13] & q[15] /*6318*/;
  assign _105_ = m_1[13] & _103_ /*6317*/;
  assign r_1[28] = _105_ | _104_ /*6316*/;
  assign _106_ = ~q[15] /*6315*/;
  assign _107_ = sum_1[14] & q[15] /*6314*/;
  assign _108_ = m_1[14] & _106_ /*6313*/;
  assign r_1[29] = _108_ | _107_ /*6312*/;
  assign _109_ = ~q[15] /*6311*/;
  assign _110_ = sum_1[15] & q[15] /*6310*/;
  assign _111_ = m_1[15] & _109_ /*6309*/;
  assign r_1[30] = _111_ | _110_ /*6308*/;
assign r_1[0]= r_0[0] /*6307*/;
assign r_1[1]= r_0[1] /*6306*/;
assign r_1[2]= r_0[2] /*6305*/;
assign r_1[3]= r_0[3] /*6304*/;
assign r_1[4]= r_0[4] /*6303*/;
assign r_1[5]= r_0[5] /*6302*/;
assign r_1[6]= r_0[6] /*6301*/;
assign r_1[7]= r_0[7] /*6300*/;
assign r_1[8]= r_0[8] /*6299*/;
assign r_1[9]= r_0[9] /*6298*/;
assign r_1[10]= r_0[10] /*6297*/;
assign r_1[11]= r_0[11] /*6296*/;
assign r_1[12]= r_0[12] /*6295*/;
assign r_1[13]= r_0[13] /*6294*/;
assign r_1[14]= r_0[14] /*6293*/;
  assign inv_2[0] = ~div[0] /*6264*/;
  assign inv_2[1] = ~div[1] /*6263*/;
  assign inv_2[2] = ~div[2] /*6262*/;
  assign inv_2[3] = ~div[3] /*6261*/;
  assign inv_2[4] = ~div[4] /*6260*/;
  assign inv_2[5] = ~div[5] /*6259*/;
  assign inv_2[6] = ~div[6] /*6258*/;
  assign inv_2[7] = ~div[7] /*6257*/;
  assign inv_2[8] = ~div[8] /*6256*/;
  assign inv_2[9] = ~div[9] /*6255*/;
  assign inv_2[10] = ~div[10] /*6254*/;
  assign inv_2[11] = ~div[11] /*6253*/;
  assign inv_2[12] = ~div[12] /*6252*/;
  assign inv_2[13] = ~div[13] /*6251*/;
  assign inv_2[14] = ~div[14] /*6250*/;
assign inv_2[15] = oneWire /*6249*/;
  assign _112_ = inv_2[0] ^ r_1[14] /*6247*/;
  assign sum_2[0] = _112_ ^ oneWire /*6246*/;
  assign _113_ = _112_ & oneWire /*6245*/;
  assign _114_ = inv_2[0] & r_1[14] /*6244*/;
  assign _115_ = _113_ | _114_ /*6243*/;
  assign _116_ = inv_2[1] ^ r_1[15] /*6242*/;
  assign sum_2[1] = _116_ ^ _115_ /*6241*/;
  assign _117_ = _116_ & _115_ /*6240*/;
  assign _118_ = inv_2[1] & r_1[15] /*6239*/;
  assign _119_ = _117_ | _118_ /*6238*/;
  assign _120_ = inv_2[2] ^ r_1[16] /*6236*/;
  assign sum_2[2] = _120_ ^ _119_ /*6235*/;
  assign _121_ = _120_ & _119_ /*6234*/;
  assign _122_ = inv_2[2] & r_1[16] /*6233*/;
  assign _123_ = _121_ | _122_ /*6232*/;
  assign _124_ = inv_2[3] ^ r_1[17] /*6230*/;
  assign sum_2[3] = _124_ ^ _123_ /*6229*/;
  assign _125_ = _124_ & _123_ /*6228*/;
  assign _126_ = inv_2[3] & r_1[17] /*6227*/;
  assign _127_ = _125_ | _126_ /*6226*/;
  assign _128_ = inv_2[4] ^ r_1[18] /*6224*/;
  assign sum_2[4] = _128_ ^ _127_ /*6223*/;
  assign _129_ = _128_ & _127_ /*6222*/;
  assign _130_ = inv_2[4] & r_1[18] /*6221*/;
  assign _131_ = _129_ | _130_ /*6220*/;
  assign _132_ = inv_2[5] ^ r_1[19] /*6218*/;
  assign sum_2[5] = _132_ ^ _131_ /*6217*/;
  assign _133_ = _132_ & _131_ /*6216*/;
  assign _134_ = inv_2[5] & r_1[19] /*6215*/;
  assign _135_ = _133_ | _134_ /*6214*/;
  assign _136_ = inv_2[6] ^ r_1[20] /*6212*/;
  assign sum_2[6] = _136_ ^ _135_ /*6211*/;
  assign _137_ = _136_ & _135_ /*6210*/;
  assign _138_ = inv_2[6] & r_1[20] /*6209*/;
  assign _139_ = _137_ | _138_ /*6208*/;
  assign _140_ = inv_2[7] ^ r_1[21] /*6206*/;
  assign sum_2[7] = _140_ ^ _139_ /*6205*/;
  assign _141_ = _140_ & _139_ /*6204*/;
  assign _142_ = inv_2[7] & r_1[21] /*6203*/;
  assign _143_ = _141_ | _142_ /*6202*/;
  assign _144_ = inv_2[8] ^ r_1[22] /*6200*/;
  assign sum_2[8] = _144_ ^ _143_ /*6199*/;
  assign _145_ = _144_ & _143_ /*6198*/;
  assign _146_ = inv_2[8] & r_1[22] /*6197*/;
  assign _147_ = _145_ | _146_ /*6196*/;
  assign _148_ = inv_2[9] ^ r_1[23] /*6194*/;
  assign sum_2[9] = _148_ ^ _147_ /*6193*/;
  assign _149_ = _148_ & _147_ /*6192*/;
  assign _150_ = inv_2[9] & r_1[23] /*6191*/;
  assign _151_ = _149_ | _150_ /*6190*/;
  assign _152_ = inv_2[10] ^ r_1[24] /*6188*/;
  assign sum_2[10] = _152_ ^ _151_ /*6187*/;
  assign _153_ = _152_ & _151_ /*6186*/;
  assign _154_ = inv_2[10] & r_1[24] /*6185*/;
  assign _155_ = _153_ | _154_ /*6184*/;
  assign _156_ = inv_2[11] ^ r_1[25] /*6182*/;
  assign sum_2[11] = _156_ ^ _155_ /*6181*/;
  assign _157_ = _156_ & _155_ /*6180*/;
  assign _158_ = inv_2[11] & r_1[25] /*6179*/;
  assign _159_ = _157_ | _158_ /*6178*/;
  assign _160_ = inv_2[12] ^ r_1[26] /*6176*/;
  assign sum_2[12] = _160_ ^ _159_ /*6175*/;
  assign _161_ = _160_ & _159_ /*6174*/;
  assign _162_ = inv_2[12] & r_1[26] /*6173*/;
  assign _163_ = _161_ | _162_ /*6172*/;
  assign _164_ = inv_2[13] ^ r_1[27] /*6170*/;
  assign sum_2[13] = _164_ ^ _163_ /*6169*/;
  assign _165_ = _164_ & _163_ /*6168*/;
  assign _166_ = inv_2[13] & r_1[27] /*6167*/;
  assign _167_ = _165_ | _166_ /*6166*/;
  assign _168_ = inv_2[14] ^ r_1[28] /*6164*/;
  assign sum_2[14] = _168_ ^ _167_ /*6163*/;
  assign _169_ = _168_ & _167_ /*6162*/;
  assign _170_ = inv_2[14] & r_1[28] /*6161*/;
  assign _171_ = _169_ | _170_ /*6160*/;
  assign _172_ = inv_2[15] ^ r_1[29] /*6158*/;
  assign sum_2[15] = _172_ ^ _171_ /*6157*/;
  assign _173_ = _172_ & _171_ /*6156*/;
  assign _174_ = inv_2[15] & r_1[29] /*6155*/;
  assign _175_ = _173_ | _174_ /*6154*/;
  assign q[14] = ~sum_2[15] /*6165*/;
  assign m_2[0] = r_1[14] /*6164*/;
  assign m_2[1] = r_1[15] /*6163*/;
  assign m_2[2] = r_1[16] /*6162*/;
  assign m_2[3] = r_1[17] /*6161*/;
  assign m_2[4] = r_1[18] /*6160*/;
  assign m_2[5] = r_1[19] /*6159*/;
  assign m_2[6] = r_1[20] /*6158*/;
  assign m_2[7] = r_1[21] /*6157*/;
  assign m_2[8] = r_1[22] /*6156*/;
  assign m_2[9] = r_1[23] /*6155*/;
  assign m_2[10] = r_1[24] /*6154*/;
  assign m_2[11] = r_1[25] /*6153*/;
  assign m_2[12] = r_1[26] /*6152*/;
  assign m_2[13] = r_1[27] /*6151*/;
  assign m_2[14] = r_1[28] /*6150*/;
  assign m_2[15] = r_1[29] /*6149*/;
  assign _176_ = ~q[14] /*6147*/;
  assign _177_ = sum_2[0] & q[14] /*6146*/;
  assign _178_ = m_2[0] & _176_ /*6145*/;
  assign r_2[14] = _178_ | _177_ /*6144*/;
  assign _179_ = ~q[14] /*6143*/;
  assign _180_ = sum_2[1] & q[14] /*6142*/;
  assign _181_ = m_2[1] & _179_ /*6141*/;
  assign r_2[15] = _181_ | _180_ /*6140*/;
  assign _182_ = ~q[14] /*6139*/;
  assign _183_ = sum_2[2] & q[14] /*6138*/;
  assign _184_ = m_2[2] & _182_ /*6137*/;
  assign r_2[16] = _184_ | _183_ /*6136*/;
  assign _185_ = ~q[14] /*6135*/;
  assign _186_ = sum_2[3] & q[14] /*6134*/;
  assign _187_ = m_2[3] & _185_ /*6133*/;
  assign r_2[17] = _187_ | _186_ /*6132*/;
  assign _188_ = ~q[14] /*6131*/;
  assign _189_ = sum_2[4] & q[14] /*6130*/;
  assign _190_ = m_2[4] & _188_ /*6129*/;
  assign r_2[18] = _190_ | _189_ /*6128*/;
  assign _191_ = ~q[14] /*6127*/;
  assign _192_ = sum_2[5] & q[14] /*6126*/;
  assign _193_ = m_2[5] & _191_ /*6125*/;
  assign r_2[19] = _193_ | _192_ /*6124*/;
  assign _194_ = ~q[14] /*6123*/;
  assign _195_ = sum_2[6] & q[14] /*6122*/;
  assign _196_ = m_2[6] & _194_ /*6121*/;
  assign r_2[20] = _196_ | _195_ /*6120*/;
  assign _197_ = ~q[14] /*6119*/;
  assign _198_ = sum_2[7] & q[14] /*6118*/;
  assign _199_ = m_2[7] & _197_ /*6117*/;
  assign r_2[21] = _199_ | _198_ /*6116*/;
  assign _200_ = ~q[14] /*6115*/;
  assign _201_ = sum_2[8] & q[14] /*6114*/;
  assign _202_ = m_2[8] & _200_ /*6113*/;
  assign r_2[22] = _202_ | _201_ /*6112*/;
  assign _203_ = ~q[14] /*6111*/;
  assign _204_ = sum_2[9] & q[14] /*6110*/;
  assign _205_ = m_2[9] & _203_ /*6109*/;
  assign r_2[23] = _205_ | _204_ /*6108*/;
  assign _206_ = ~q[14] /*6107*/;
  assign _207_ = sum_2[10] & q[14] /*6106*/;
  assign _208_ = m_2[10] & _206_ /*6105*/;
  assign r_2[24] = _208_ | _207_ /*6104*/;
  assign _209_ = ~q[14] /*6103*/;
  assign _210_ = sum_2[11] & q[14] /*6102*/;
  assign _211_ = m_2[11] & _209_ /*6101*/;
  assign r_2[25] = _211_ | _210_ /*6100*/;
  assign _212_ = ~q[14] /*6099*/;
  assign _213_ = sum_2[12] & q[14] /*6098*/;
  assign _214_ = m_2[12] & _212_ /*6097*/;
  assign r_2[26] = _214_ | _213_ /*6096*/;
  assign _215_ = ~q[14] /*6095*/;
  assign _216_ = sum_2[13] & q[14] /*6094*/;
  assign _217_ = m_2[13] & _215_ /*6093*/;
  assign r_2[27] = _217_ | _216_ /*6092*/;
  assign _218_ = ~q[14] /*6091*/;
  assign _219_ = sum_2[14] & q[14] /*6090*/;
  assign _220_ = m_2[14] & _218_ /*6089*/;
  assign r_2[28] = _220_ | _219_ /*6088*/;
  assign _221_ = ~q[14] /*6087*/;
  assign _222_ = sum_2[15] & q[14] /*6086*/;
  assign _223_ = m_2[15] & _221_ /*6085*/;
  assign r_2[29] = _223_ | _222_ /*6084*/;
assign r_2[0]= r_1[0] /*6083*/;
assign r_2[1]= r_1[1] /*6082*/;
assign r_2[2]= r_1[2] /*6081*/;
assign r_2[3]= r_1[3] /*6080*/;
assign r_2[4]= r_1[4] /*6079*/;
assign r_2[5]= r_1[5] /*6078*/;
assign r_2[6]= r_1[6] /*6077*/;
assign r_2[7]= r_1[7] /*6076*/;
assign r_2[8]= r_1[8] /*6075*/;
assign r_2[9]= r_1[9] /*6074*/;
assign r_2[10]= r_1[10] /*6073*/;
assign r_2[11]= r_1[11] /*6072*/;
assign r_2[12]= r_1[12] /*6071*/;
assign r_2[13]= r_1[13] /*6070*/;
  assign inv_3[0] = ~div[0] /*6040*/;
  assign inv_3[1] = ~div[1] /*6039*/;
  assign inv_3[2] = ~div[2] /*6038*/;
  assign inv_3[3] = ~div[3] /*6037*/;
  assign inv_3[4] = ~div[4] /*6036*/;
  assign inv_3[5] = ~div[5] /*6035*/;
  assign inv_3[6] = ~div[6] /*6034*/;
  assign inv_3[7] = ~div[7] /*6033*/;
  assign inv_3[8] = ~div[8] /*6032*/;
  assign inv_3[9] = ~div[9] /*6031*/;
  assign inv_3[10] = ~div[10] /*6030*/;
  assign inv_3[11] = ~div[11] /*6029*/;
  assign inv_3[12] = ~div[12] /*6028*/;
  assign inv_3[13] = ~div[13] /*6027*/;
  assign inv_3[14] = ~div[14] /*6026*/;
assign inv_3[15] = oneWire /*6025*/;
  assign _224_ = inv_3[0] ^ r_2[13] /*6023*/;
  assign sum_3[0] = _224_ ^ oneWire /*6022*/;
  assign _225_ = _224_ & oneWire /*6021*/;
  assign _226_ = inv_3[0] & r_2[13] /*6020*/;
  assign _227_ = _225_ | _226_ /*6019*/;
  assign _228_ = inv_3[1] ^ r_2[14] /*6018*/;
  assign sum_3[1] = _228_ ^ _227_ /*6017*/;
  assign _229_ = _228_ & _227_ /*6016*/;
  assign _230_ = inv_3[1] & r_2[14] /*6015*/;
  assign _231_ = _229_ | _230_ /*6014*/;
  assign _232_ = inv_3[2] ^ r_2[15] /*6012*/;
  assign sum_3[2] = _232_ ^ _231_ /*6011*/;
  assign _233_ = _232_ & _231_ /*6010*/;
  assign _234_ = inv_3[2] & r_2[15] /*6009*/;
  assign _235_ = _233_ | _234_ /*6008*/;
  assign _236_ = inv_3[3] ^ r_2[16] /*6006*/;
  assign sum_3[3] = _236_ ^ _235_ /*6005*/;
  assign _237_ = _236_ & _235_ /*6004*/;
  assign _238_ = inv_3[3] & r_2[16] /*6003*/;
  assign _239_ = _237_ | _238_ /*6002*/;
  assign _240_ = inv_3[4] ^ r_2[17] /*6000*/;
  assign sum_3[4] = _240_ ^ _239_ /*5999*/;
  assign _241_ = _240_ & _239_ /*5998*/;
  assign _242_ = inv_3[4] & r_2[17] /*5997*/;
  assign _243_ = _241_ | _242_ /*5996*/;
  assign _244_ = inv_3[5] ^ r_2[18] /*5994*/;
  assign sum_3[5] = _244_ ^ _243_ /*5993*/;
  assign _245_ = _244_ & _243_ /*5992*/;
  assign _246_ = inv_3[5] & r_2[18] /*5991*/;
  assign _247_ = _245_ | _246_ /*5990*/;
  assign _248_ = inv_3[6] ^ r_2[19] /*5988*/;
  assign sum_3[6] = _248_ ^ _247_ /*5987*/;
  assign _249_ = _248_ & _247_ /*5986*/;
  assign _250_ = inv_3[6] & r_2[19] /*5985*/;
  assign _251_ = _249_ | _250_ /*5984*/;
  assign _252_ = inv_3[7] ^ r_2[20] /*5982*/;
  assign sum_3[7] = _252_ ^ _251_ /*5981*/;
  assign _253_ = _252_ & _251_ /*5980*/;
  assign _254_ = inv_3[7] & r_2[20] /*5979*/;
  assign _255_ = _253_ | _254_ /*5978*/;
  assign _256_ = inv_3[8] ^ r_2[21] /*5976*/;
  assign sum_3[8] = _256_ ^ _255_ /*5975*/;
  assign _257_ = _256_ & _255_ /*5974*/;
  assign _258_ = inv_3[8] & r_2[21] /*5973*/;
  assign _259_ = _257_ | _258_ /*5972*/;
  assign _260_ = inv_3[9] ^ r_2[22] /*5970*/;
  assign sum_3[9] = _260_ ^ _259_ /*5969*/;
  assign _261_ = _260_ & _259_ /*5968*/;
  assign _262_ = inv_3[9] & r_2[22] /*5967*/;
  assign _263_ = _261_ | _262_ /*5966*/;
  assign _264_ = inv_3[10] ^ r_2[23] /*5964*/;
  assign sum_3[10] = _264_ ^ _263_ /*5963*/;
  assign _265_ = _264_ & _263_ /*5962*/;
  assign _266_ = inv_3[10] & r_2[23] /*5961*/;
  assign _267_ = _265_ | _266_ /*5960*/;
  assign _268_ = inv_3[11] ^ r_2[24] /*5958*/;
  assign sum_3[11] = _268_ ^ _267_ /*5957*/;
  assign _269_ = _268_ & _267_ /*5956*/;
  assign _270_ = inv_3[11] & r_2[24] /*5955*/;
  assign _271_ = _269_ | _270_ /*5954*/;
  assign _272_ = inv_3[12] ^ r_2[25] /*5952*/;
  assign sum_3[12] = _272_ ^ _271_ /*5951*/;
  assign _273_ = _272_ & _271_ /*5950*/;
  assign _274_ = inv_3[12] & r_2[25] /*5949*/;
  assign _275_ = _273_ | _274_ /*5948*/;
  assign _276_ = inv_3[13] ^ r_2[26] /*5946*/;
  assign sum_3[13] = _276_ ^ _275_ /*5945*/;
  assign _277_ = _276_ & _275_ /*5944*/;
  assign _278_ = inv_3[13] & r_2[26] /*5943*/;
  assign _279_ = _277_ | _278_ /*5942*/;
  assign _280_ = inv_3[14] ^ r_2[27] /*5940*/;
  assign sum_3[14] = _280_ ^ _279_ /*5939*/;
  assign _281_ = _280_ & _279_ /*5938*/;
  assign _282_ = inv_3[14] & r_2[27] /*5937*/;
  assign _283_ = _281_ | _282_ /*5936*/;
  assign _284_ = inv_3[15] ^ r_2[28] /*5934*/;
  assign sum_3[15] = _284_ ^ _283_ /*5933*/;
  assign _285_ = _284_ & _283_ /*5932*/;
  assign _286_ = inv_3[15] & r_2[28] /*5931*/;
  assign _287_ = _285_ | _286_ /*5930*/;
  assign q[13] = ~sum_3[15] /*5941*/;
  assign m_3[0] = r_2[13] /*5940*/;
  assign m_3[1] = r_2[14] /*5939*/;
  assign m_3[2] = r_2[15] /*5938*/;
  assign m_3[3] = r_2[16] /*5937*/;
  assign m_3[4] = r_2[17] /*5936*/;
  assign m_3[5] = r_2[18] /*5935*/;
  assign m_3[6] = r_2[19] /*5934*/;
  assign m_3[7] = r_2[20] /*5933*/;
  assign m_3[8] = r_2[21] /*5932*/;
  assign m_3[9] = r_2[22] /*5931*/;
  assign m_3[10] = r_2[23] /*5930*/;
  assign m_3[11] = r_2[24] /*5929*/;
  assign m_3[12] = r_2[25] /*5928*/;
  assign m_3[13] = r_2[26] /*5927*/;
  assign m_3[14] = r_2[27] /*5926*/;
  assign m_3[15] = r_2[28] /*5925*/;
  assign _288_ = ~q[13] /*5923*/;
  assign _289_ = sum_3[0] & q[13] /*5922*/;
  assign _290_ = m_3[0] & _288_ /*5921*/;
  assign r_3[13] = _290_ | _289_ /*5920*/;
  assign _291_ = ~q[13] /*5919*/;
  assign _292_ = sum_3[1] & q[13] /*5918*/;
  assign _293_ = m_3[1] & _291_ /*5917*/;
  assign r_3[14] = _293_ | _292_ /*5916*/;
  assign _294_ = ~q[13] /*5915*/;
  assign _295_ = sum_3[2] & q[13] /*5914*/;
  assign _296_ = m_3[2] & _294_ /*5913*/;
  assign r_3[15] = _296_ | _295_ /*5912*/;
  assign _297_ = ~q[13] /*5911*/;
  assign _298_ = sum_3[3] & q[13] /*5910*/;
  assign _299_ = m_3[3] & _297_ /*5909*/;
  assign r_3[16] = _299_ | _298_ /*5908*/;
  assign _300_ = ~q[13] /*5907*/;
  assign _301_ = sum_3[4] & q[13] /*5906*/;
  assign _302_ = m_3[4] & _300_ /*5905*/;
  assign r_3[17] = _302_ | _301_ /*5904*/;
  assign _303_ = ~q[13] /*5903*/;
  assign _304_ = sum_3[5] & q[13] /*5902*/;
  assign _305_ = m_3[5] & _303_ /*5901*/;
  assign r_3[18] = _305_ | _304_ /*5900*/;
  assign _306_ = ~q[13] /*5899*/;
  assign _307_ = sum_3[6] & q[13] /*5898*/;
  assign _308_ = m_3[6] & _306_ /*5897*/;
  assign r_3[19] = _308_ | _307_ /*5896*/;
  assign _309_ = ~q[13] /*5895*/;
  assign _310_ = sum_3[7] & q[13] /*5894*/;
  assign _311_ = m_3[7] & _309_ /*5893*/;
  assign r_3[20] = _311_ | _310_ /*5892*/;
  assign _312_ = ~q[13] /*5891*/;
  assign _313_ = sum_3[8] & q[13] /*5890*/;
  assign _314_ = m_3[8] & _312_ /*5889*/;
  assign r_3[21] = _314_ | _313_ /*5888*/;
  assign _315_ = ~q[13] /*5887*/;
  assign _316_ = sum_3[9] & q[13] /*5886*/;
  assign _317_ = m_3[9] & _315_ /*5885*/;
  assign r_3[22] = _317_ | _316_ /*5884*/;
  assign _318_ = ~q[13] /*5883*/;
  assign _319_ = sum_3[10] & q[13] /*5882*/;
  assign _320_ = m_3[10] & _318_ /*5881*/;
  assign r_3[23] = _320_ | _319_ /*5880*/;
  assign _321_ = ~q[13] /*5879*/;
  assign _322_ = sum_3[11] & q[13] /*5878*/;
  assign _323_ = m_3[11] & _321_ /*5877*/;
  assign r_3[24] = _323_ | _322_ /*5876*/;
  assign _324_ = ~q[13] /*5875*/;
  assign _325_ = sum_3[12] & q[13] /*5874*/;
  assign _326_ = m_3[12] & _324_ /*5873*/;
  assign r_3[25] = _326_ | _325_ /*5872*/;
  assign _327_ = ~q[13] /*5871*/;
  assign _328_ = sum_3[13] & q[13] /*5870*/;
  assign _329_ = m_3[13] & _327_ /*5869*/;
  assign r_3[26] = _329_ | _328_ /*5868*/;
  assign _330_ = ~q[13] /*5867*/;
  assign _331_ = sum_3[14] & q[13] /*5866*/;
  assign _332_ = m_3[14] & _330_ /*5865*/;
  assign r_3[27] = _332_ | _331_ /*5864*/;
  assign _333_ = ~q[13] /*5863*/;
  assign _334_ = sum_3[15] & q[13] /*5862*/;
  assign _335_ = m_3[15] & _333_ /*5861*/;
  assign r_3[28] = _335_ | _334_ /*5860*/;
assign r_3[0]= r_2[0] /*5859*/;
assign r_3[1]= r_2[1] /*5858*/;
assign r_3[2]= r_2[2] /*5857*/;
assign r_3[3]= r_2[3] /*5856*/;
assign r_3[4]= r_2[4] /*5855*/;
assign r_3[5]= r_2[5] /*5854*/;
assign r_3[6]= r_2[6] /*5853*/;
assign r_3[7]= r_2[7] /*5852*/;
assign r_3[8]= r_2[8] /*5851*/;
assign r_3[9]= r_2[9] /*5850*/;
assign r_3[10]= r_2[10] /*5849*/;
assign r_3[11]= r_2[11] /*5848*/;
assign r_3[12]= r_2[12] /*5847*/;
  assign inv_4[0] = ~div[0] /*5816*/;
  assign inv_4[1] = ~div[1] /*5815*/;
  assign inv_4[2] = ~div[2] /*5814*/;
  assign inv_4[3] = ~div[3] /*5813*/;
  assign inv_4[4] = ~div[4] /*5812*/;
  assign inv_4[5] = ~div[5] /*5811*/;
  assign inv_4[6] = ~div[6] /*5810*/;
  assign inv_4[7] = ~div[7] /*5809*/;
  assign inv_4[8] = ~div[8] /*5808*/;
  assign inv_4[9] = ~div[9] /*5807*/;
  assign inv_4[10] = ~div[10] /*5806*/;
  assign inv_4[11] = ~div[11] /*5805*/;
  assign inv_4[12] = ~div[12] /*5804*/;
  assign inv_4[13] = ~div[13] /*5803*/;
  assign inv_4[14] = ~div[14] /*5802*/;
assign inv_4[15] = oneWire /*5801*/;
  assign _336_ = inv_4[0] ^ r_3[12] /*5799*/;
  assign sum_4[0] = _336_ ^ oneWire /*5798*/;
  assign _337_ = _336_ & oneWire /*5797*/;
  assign _338_ = inv_4[0] & r_3[12] /*5796*/;
  assign _339_ = _337_ | _338_ /*5795*/;
  assign _340_ = inv_4[1] ^ r_3[13] /*5794*/;
  assign sum_4[1] = _340_ ^ _339_ /*5793*/;
  assign _341_ = _340_ & _339_ /*5792*/;
  assign _342_ = inv_4[1] & r_3[13] /*5791*/;
  assign _343_ = _341_ | _342_ /*5790*/;
  assign _344_ = inv_4[2] ^ r_3[14] /*5788*/;
  assign sum_4[2] = _344_ ^ _343_ /*5787*/;
  assign _345_ = _344_ & _343_ /*5786*/;
  assign _346_ = inv_4[2] & r_3[14] /*5785*/;
  assign _347_ = _345_ | _346_ /*5784*/;
  assign _348_ = inv_4[3] ^ r_3[15] /*5782*/;
  assign sum_4[3] = _348_ ^ _347_ /*5781*/;
  assign _349_ = _348_ & _347_ /*5780*/;
  assign _350_ = inv_4[3] & r_3[15] /*5779*/;
  assign _351_ = _349_ | _350_ /*5778*/;
  assign _352_ = inv_4[4] ^ r_3[16] /*5776*/;
  assign sum_4[4] = _352_ ^ _351_ /*5775*/;
  assign _353_ = _352_ & _351_ /*5774*/;
  assign _354_ = inv_4[4] & r_3[16] /*5773*/;
  assign _355_ = _353_ | _354_ /*5772*/;
  assign _356_ = inv_4[5] ^ r_3[17] /*5770*/;
  assign sum_4[5] = _356_ ^ _355_ /*5769*/;
  assign _357_ = _356_ & _355_ /*5768*/;
  assign _358_ = inv_4[5] & r_3[17] /*5767*/;
  assign _359_ = _357_ | _358_ /*5766*/;
  assign _360_ = inv_4[6] ^ r_3[18] /*5764*/;
  assign sum_4[6] = _360_ ^ _359_ /*5763*/;
  assign _361_ = _360_ & _359_ /*5762*/;
  assign _362_ = inv_4[6] & r_3[18] /*5761*/;
  assign _363_ = _361_ | _362_ /*5760*/;
  assign _364_ = inv_4[7] ^ r_3[19] /*5758*/;
  assign sum_4[7] = _364_ ^ _363_ /*5757*/;
  assign _365_ = _364_ & _363_ /*5756*/;
  assign _366_ = inv_4[7] & r_3[19] /*5755*/;
  assign _367_ = _365_ | _366_ /*5754*/;
  assign _368_ = inv_4[8] ^ r_3[20] /*5752*/;
  assign sum_4[8] = _368_ ^ _367_ /*5751*/;
  assign _369_ = _368_ & _367_ /*5750*/;
  assign _370_ = inv_4[8] & r_3[20] /*5749*/;
  assign _371_ = _369_ | _370_ /*5748*/;
  assign _372_ = inv_4[9] ^ r_3[21] /*5746*/;
  assign sum_4[9] = _372_ ^ _371_ /*5745*/;
  assign _373_ = _372_ & _371_ /*5744*/;
  assign _374_ = inv_4[9] & r_3[21] /*5743*/;
  assign _375_ = _373_ | _374_ /*5742*/;
  assign _376_ = inv_4[10] ^ r_3[22] /*5740*/;
  assign sum_4[10] = _376_ ^ _375_ /*5739*/;
  assign _377_ = _376_ & _375_ /*5738*/;
  assign _378_ = inv_4[10] & r_3[22] /*5737*/;
  assign _379_ = _377_ | _378_ /*5736*/;
  assign _380_ = inv_4[11] ^ r_3[23] /*5734*/;
  assign sum_4[11] = _380_ ^ _379_ /*5733*/;
  assign _381_ = _380_ & _379_ /*5732*/;
  assign _382_ = inv_4[11] & r_3[23] /*5731*/;
  assign _383_ = _381_ | _382_ /*5730*/;
  assign _384_ = inv_4[12] ^ r_3[24] /*5728*/;
  assign sum_4[12] = _384_ ^ _383_ /*5727*/;
  assign _385_ = _384_ & _383_ /*5726*/;
  assign _386_ = inv_4[12] & r_3[24] /*5725*/;
  assign _387_ = _385_ | _386_ /*5724*/;
  assign _388_ = inv_4[13] ^ r_3[25] /*5722*/;
  assign sum_4[13] = _388_ ^ _387_ /*5721*/;
  assign _389_ = _388_ & _387_ /*5720*/;
  assign _390_ = inv_4[13] & r_3[25] /*5719*/;
  assign _391_ = _389_ | _390_ /*5718*/;
  assign _392_ = inv_4[14] ^ r_3[26] /*5716*/;
  assign sum_4[14] = _392_ ^ _391_ /*5715*/;
  assign _393_ = _392_ & _391_ /*5714*/;
  assign _394_ = inv_4[14] & r_3[26] /*5713*/;
  assign _395_ = _393_ | _394_ /*5712*/;
  assign _396_ = inv_4[15] ^ r_3[27] /*5710*/;
  assign sum_4[15] = _396_ ^ _395_ /*5709*/;
  assign _397_ = _396_ & _395_ /*5708*/;
  assign _398_ = inv_4[15] & r_3[27] /*5707*/;
  assign _399_ = _397_ | _398_ /*5706*/;
  assign q[12] = ~sum_4[15] /*5717*/;
  assign m_4[0] = r_3[12] /*5716*/;
  assign m_4[1] = r_3[13] /*5715*/;
  assign m_4[2] = r_3[14] /*5714*/;
  assign m_4[3] = r_3[15] /*5713*/;
  assign m_4[4] = r_3[16] /*5712*/;
  assign m_4[5] = r_3[17] /*5711*/;
  assign m_4[6] = r_3[18] /*5710*/;
  assign m_4[7] = r_3[19] /*5709*/;
  assign m_4[8] = r_3[20] /*5708*/;
  assign m_4[9] = r_3[21] /*5707*/;
  assign m_4[10] = r_3[22] /*5706*/;
  assign m_4[11] = r_3[23] /*5705*/;
  assign m_4[12] = r_3[24] /*5704*/;
  assign m_4[13] = r_3[25] /*5703*/;
  assign m_4[14] = r_3[26] /*5702*/;
  assign m_4[15] = r_3[27] /*5701*/;
  assign _400_ = ~q[12] /*5699*/;
  assign _401_ = sum_4[0] & q[12] /*5698*/;
  assign _402_ = m_4[0] & _400_ /*5697*/;
  assign r_4[12] = _402_ | _401_ /*5696*/;
  assign _403_ = ~q[12] /*5695*/;
  assign _404_ = sum_4[1] & q[12] /*5694*/;
  assign _405_ = m_4[1] & _403_ /*5693*/;
  assign r_4[13] = _405_ | _404_ /*5692*/;
  assign _406_ = ~q[12] /*5691*/;
  assign _407_ = sum_4[2] & q[12] /*5690*/;
  assign _408_ = m_4[2] & _406_ /*5689*/;
  assign r_4[14] = _408_ | _407_ /*5688*/;
  assign _409_ = ~q[12] /*5687*/;
  assign _410_ = sum_4[3] & q[12] /*5686*/;
  assign _411_ = m_4[3] & _409_ /*5685*/;
  assign r_4[15] = _411_ | _410_ /*5684*/;
  assign _412_ = ~q[12] /*5683*/;
  assign _413_ = sum_4[4] & q[12] /*5682*/;
  assign _414_ = m_4[4] & _412_ /*5681*/;
  assign r_4[16] = _414_ | _413_ /*5680*/;
  assign _415_ = ~q[12] /*5679*/;
  assign _416_ = sum_4[5] & q[12] /*5678*/;
  assign _417_ = m_4[5] & _415_ /*5677*/;
  assign r_4[17] = _417_ | _416_ /*5676*/;
  assign _418_ = ~q[12] /*5675*/;
  assign _419_ = sum_4[6] & q[12] /*5674*/;
  assign _420_ = m_4[6] & _418_ /*5673*/;
  assign r_4[18] = _420_ | _419_ /*5672*/;
  assign _421_ = ~q[12] /*5671*/;
  assign _422_ = sum_4[7] & q[12] /*5670*/;
  assign _423_ = m_4[7] & _421_ /*5669*/;
  assign r_4[19] = _423_ | _422_ /*5668*/;
  assign _424_ = ~q[12] /*5667*/;
  assign _425_ = sum_4[8] & q[12] /*5666*/;
  assign _426_ = m_4[8] & _424_ /*5665*/;
  assign r_4[20] = _426_ | _425_ /*5664*/;
  assign _427_ = ~q[12] /*5663*/;
  assign _428_ = sum_4[9] & q[12] /*5662*/;
  assign _429_ = m_4[9] & _427_ /*5661*/;
  assign r_4[21] = _429_ | _428_ /*5660*/;
  assign _430_ = ~q[12] /*5659*/;
  assign _431_ = sum_4[10] & q[12] /*5658*/;
  assign _432_ = m_4[10] & _430_ /*5657*/;
  assign r_4[22] = _432_ | _431_ /*5656*/;
  assign _433_ = ~q[12] /*5655*/;
  assign _434_ = sum_4[11] & q[12] /*5654*/;
  assign _435_ = m_4[11] & _433_ /*5653*/;
  assign r_4[23] = _435_ | _434_ /*5652*/;
  assign _436_ = ~q[12] /*5651*/;
  assign _437_ = sum_4[12] & q[12] /*5650*/;
  assign _438_ = m_4[12] & _436_ /*5649*/;
  assign r_4[24] = _438_ | _437_ /*5648*/;
  assign _439_ = ~q[12] /*5647*/;
  assign _440_ = sum_4[13] & q[12] /*5646*/;
  assign _441_ = m_4[13] & _439_ /*5645*/;
  assign r_4[25] = _441_ | _440_ /*5644*/;
  assign _442_ = ~q[12] /*5643*/;
  assign _443_ = sum_4[14] & q[12] /*5642*/;
  assign _444_ = m_4[14] & _442_ /*5641*/;
  assign r_4[26] = _444_ | _443_ /*5640*/;
  assign _445_ = ~q[12] /*5639*/;
  assign _446_ = sum_4[15] & q[12] /*5638*/;
  assign _447_ = m_4[15] & _445_ /*5637*/;
  assign r_4[27] = _447_ | _446_ /*5636*/;
assign r_4[0]= r_3[0] /*5635*/;
assign r_4[1]= r_3[1] /*5634*/;
assign r_4[2]= r_3[2] /*5633*/;
assign r_4[3]= r_3[3] /*5632*/;
assign r_4[4]= r_3[4] /*5631*/;
assign r_4[5]= r_3[5] /*5630*/;
assign r_4[6]= r_3[6] /*5629*/;
assign r_4[7]= r_3[7] /*5628*/;
assign r_4[8]= r_3[8] /*5627*/;
assign r_4[9]= r_3[9] /*5626*/;
assign r_4[10]= r_3[10] /*5625*/;
assign r_4[11]= r_3[11] /*5624*/;
  assign inv_5[0] = ~div[0] /*5592*/;
  assign inv_5[1] = ~div[1] /*5591*/;
  assign inv_5[2] = ~div[2] /*5590*/;
  assign inv_5[3] = ~div[3] /*5589*/;
  assign inv_5[4] = ~div[4] /*5588*/;
  assign inv_5[5] = ~div[5] /*5587*/;
  assign inv_5[6] = ~div[6] /*5586*/;
  assign inv_5[7] = ~div[7] /*5585*/;
  assign inv_5[8] = ~div[8] /*5584*/;
  assign inv_5[9] = ~div[9] /*5583*/;
  assign inv_5[10] = ~div[10] /*5582*/;
  assign inv_5[11] = ~div[11] /*5581*/;
  assign inv_5[12] = ~div[12] /*5580*/;
  assign inv_5[13] = ~div[13] /*5579*/;
  assign inv_5[14] = ~div[14] /*5578*/;
assign inv_5[15] = oneWire /*5577*/;
  assign _448_ = inv_5[0] ^ r_4[11] /*5575*/;
  assign sum_5[0] = _448_ ^ oneWire /*5574*/;
  assign _449_ = _448_ & oneWire /*5573*/;
  assign _450_ = inv_5[0] & r_4[11] /*5572*/;
  assign _451_ = _449_ | _450_ /*5571*/;
  assign _452_ = inv_5[1] ^ r_4[12] /*5570*/;
  assign sum_5[1] = _452_ ^ _451_ /*5569*/;
  assign _453_ = _452_ & _451_ /*5568*/;
  assign _454_ = inv_5[1] & r_4[12] /*5567*/;
  assign _455_ = _453_ | _454_ /*5566*/;
  assign _456_ = inv_5[2] ^ r_4[13] /*5564*/;
  assign sum_5[2] = _456_ ^ _455_ /*5563*/;
  assign _457_ = _456_ & _455_ /*5562*/;
  assign _458_ = inv_5[2] & r_4[13] /*5561*/;
  assign _459_ = _457_ | _458_ /*5560*/;
  assign _460_ = inv_5[3] ^ r_4[14] /*5558*/;
  assign sum_5[3] = _460_ ^ _459_ /*5557*/;
  assign _461_ = _460_ & _459_ /*5556*/;
  assign _462_ = inv_5[3] & r_4[14] /*5555*/;
  assign _463_ = _461_ | _462_ /*5554*/;
  assign _464_ = inv_5[4] ^ r_4[15] /*5552*/;
  assign sum_5[4] = _464_ ^ _463_ /*5551*/;
  assign _465_ = _464_ & _463_ /*5550*/;
  assign _466_ = inv_5[4] & r_4[15] /*5549*/;
  assign _467_ = _465_ | _466_ /*5548*/;
  assign _468_ = inv_5[5] ^ r_4[16] /*5546*/;
  assign sum_5[5] = _468_ ^ _467_ /*5545*/;
  assign _469_ = _468_ & _467_ /*5544*/;
  assign _470_ = inv_5[5] & r_4[16] /*5543*/;
  assign _471_ = _469_ | _470_ /*5542*/;
  assign _472_ = inv_5[6] ^ r_4[17] /*5540*/;
  assign sum_5[6] = _472_ ^ _471_ /*5539*/;
  assign _473_ = _472_ & _471_ /*5538*/;
  assign _474_ = inv_5[6] & r_4[17] /*5537*/;
  assign _475_ = _473_ | _474_ /*5536*/;
  assign _476_ = inv_5[7] ^ r_4[18] /*5534*/;
  assign sum_5[7] = _476_ ^ _475_ /*5533*/;
  assign _477_ = _476_ & _475_ /*5532*/;
  assign _478_ = inv_5[7] & r_4[18] /*5531*/;
  assign _479_ = _477_ | _478_ /*5530*/;
  assign _480_ = inv_5[8] ^ r_4[19] /*5528*/;
  assign sum_5[8] = _480_ ^ _479_ /*5527*/;
  assign _481_ = _480_ & _479_ /*5526*/;
  assign _482_ = inv_5[8] & r_4[19] /*5525*/;
  assign _483_ = _481_ | _482_ /*5524*/;
  assign _484_ = inv_5[9] ^ r_4[20] /*5522*/;
  assign sum_5[9] = _484_ ^ _483_ /*5521*/;
  assign _485_ = _484_ & _483_ /*5520*/;
  assign _486_ = inv_5[9] & r_4[20] /*5519*/;
  assign _487_ = _485_ | _486_ /*5518*/;
  assign _488_ = inv_5[10] ^ r_4[21] /*5516*/;
  assign sum_5[10] = _488_ ^ _487_ /*5515*/;
  assign _489_ = _488_ & _487_ /*5514*/;
  assign _490_ = inv_5[10] & r_4[21] /*5513*/;
  assign _491_ = _489_ | _490_ /*5512*/;
  assign _492_ = inv_5[11] ^ r_4[22] /*5510*/;
  assign sum_5[11] = _492_ ^ _491_ /*5509*/;
  assign _493_ = _492_ & _491_ /*5508*/;
  assign _494_ = inv_5[11] & r_4[22] /*5507*/;
  assign _495_ = _493_ | _494_ /*5506*/;
  assign _496_ = inv_5[12] ^ r_4[23] /*5504*/;
  assign sum_5[12] = _496_ ^ _495_ /*5503*/;
  assign _497_ = _496_ & _495_ /*5502*/;
  assign _498_ = inv_5[12] & r_4[23] /*5501*/;
  assign _499_ = _497_ | _498_ /*5500*/;
  assign _500_ = inv_5[13] ^ r_4[24] /*5498*/;
  assign sum_5[13] = _500_ ^ _499_ /*5497*/;
  assign _501_ = _500_ & _499_ /*5496*/;
  assign _502_ = inv_5[13] & r_4[24] /*5495*/;
  assign _503_ = _501_ | _502_ /*5494*/;
  assign _504_ = inv_5[14] ^ r_4[25] /*5492*/;
  assign sum_5[14] = _504_ ^ _503_ /*5491*/;
  assign _505_ = _504_ & _503_ /*5490*/;
  assign _506_ = inv_5[14] & r_4[25] /*5489*/;
  assign _507_ = _505_ | _506_ /*5488*/;
  assign _508_ = inv_5[15] ^ r_4[26] /*5486*/;
  assign sum_5[15] = _508_ ^ _507_ /*5485*/;
  assign _509_ = _508_ & _507_ /*5484*/;
  assign _510_ = inv_5[15] & r_4[26] /*5483*/;
  assign _511_ = _509_ | _510_ /*5482*/;
  assign q[11] = ~sum_5[15] /*5493*/;
  assign m_5[0] = r_4[11] /*5492*/;
  assign m_5[1] = r_4[12] /*5491*/;
  assign m_5[2] = r_4[13] /*5490*/;
  assign m_5[3] = r_4[14] /*5489*/;
  assign m_5[4] = r_4[15] /*5488*/;
  assign m_5[5] = r_4[16] /*5487*/;
  assign m_5[6] = r_4[17] /*5486*/;
  assign m_5[7] = r_4[18] /*5485*/;
  assign m_5[8] = r_4[19] /*5484*/;
  assign m_5[9] = r_4[20] /*5483*/;
  assign m_5[10] = r_4[21] /*5482*/;
  assign m_5[11] = r_4[22] /*5481*/;
  assign m_5[12] = r_4[23] /*5480*/;
  assign m_5[13] = r_4[24] /*5479*/;
  assign m_5[14] = r_4[25] /*5478*/;
  assign m_5[15] = r_4[26] /*5477*/;
  assign _512_ = ~q[11] /*5475*/;
  assign _513_ = sum_5[0] & q[11] /*5474*/;
  assign _514_ = m_5[0] & _512_ /*5473*/;
  assign r_5[11] = _514_ | _513_ /*5472*/;
  assign _515_ = ~q[11] /*5471*/;
  assign _516_ = sum_5[1] & q[11] /*5470*/;
  assign _517_ = m_5[1] & _515_ /*5469*/;
  assign r_5[12] = _517_ | _516_ /*5468*/;
  assign _518_ = ~q[11] /*5467*/;
  assign _519_ = sum_5[2] & q[11] /*5466*/;
  assign _520_ = m_5[2] & _518_ /*5465*/;
  assign r_5[13] = _520_ | _519_ /*5464*/;
  assign _521_ = ~q[11] /*5463*/;
  assign _522_ = sum_5[3] & q[11] /*5462*/;
  assign _523_ = m_5[3] & _521_ /*5461*/;
  assign r_5[14] = _523_ | _522_ /*5460*/;
  assign _524_ = ~q[11] /*5459*/;
  assign _525_ = sum_5[4] & q[11] /*5458*/;
  assign _526_ = m_5[4] & _524_ /*5457*/;
  assign r_5[15] = _526_ | _525_ /*5456*/;
  assign _527_ = ~q[11] /*5455*/;
  assign _528_ = sum_5[5] & q[11] /*5454*/;
  assign _529_ = m_5[5] & _527_ /*5453*/;
  assign r_5[16] = _529_ | _528_ /*5452*/;
  assign _530_ = ~q[11] /*5451*/;
  assign _531_ = sum_5[6] & q[11] /*5450*/;
  assign _532_ = m_5[6] & _530_ /*5449*/;
  assign r_5[17] = _532_ | _531_ /*5448*/;
  assign _533_ = ~q[11] /*5447*/;
  assign _534_ = sum_5[7] & q[11] /*5446*/;
  assign _535_ = m_5[7] & _533_ /*5445*/;
  assign r_5[18] = _535_ | _534_ /*5444*/;
  assign _536_ = ~q[11] /*5443*/;
  assign _537_ = sum_5[8] & q[11] /*5442*/;
  assign _538_ = m_5[8] & _536_ /*5441*/;
  assign r_5[19] = _538_ | _537_ /*5440*/;
  assign _539_ = ~q[11] /*5439*/;
  assign _540_ = sum_5[9] & q[11] /*5438*/;
  assign _541_ = m_5[9] & _539_ /*5437*/;
  assign r_5[20] = _541_ | _540_ /*5436*/;
  assign _542_ = ~q[11] /*5435*/;
  assign _543_ = sum_5[10] & q[11] /*5434*/;
  assign _544_ = m_5[10] & _542_ /*5433*/;
  assign r_5[21] = _544_ | _543_ /*5432*/;
  assign _545_ = ~q[11] /*5431*/;
  assign _546_ = sum_5[11] & q[11] /*5430*/;
  assign _547_ = m_5[11] & _545_ /*5429*/;
  assign r_5[22] = _547_ | _546_ /*5428*/;
  assign _548_ = ~q[11] /*5427*/;
  assign _549_ = sum_5[12] & q[11] /*5426*/;
  assign _550_ = m_5[12] & _548_ /*5425*/;
  assign r_5[23] = _550_ | _549_ /*5424*/;
  assign _551_ = ~q[11] /*5423*/;
  assign _552_ = sum_5[13] & q[11] /*5422*/;
  assign _553_ = m_5[13] & _551_ /*5421*/;
  assign r_5[24] = _553_ | _552_ /*5420*/;
  assign _554_ = ~q[11] /*5419*/;
  assign _555_ = sum_5[14] & q[11] /*5418*/;
  assign _556_ = m_5[14] & _554_ /*5417*/;
  assign r_5[25] = _556_ | _555_ /*5416*/;
  assign _557_ = ~q[11] /*5415*/;
  assign _558_ = sum_5[15] & q[11] /*5414*/;
  assign _559_ = m_5[15] & _557_ /*5413*/;
  assign r_5[26] = _559_ | _558_ /*5412*/;
assign r_5[0]= r_4[0] /*5411*/;
assign r_5[1]= r_4[1] /*5410*/;
assign r_5[2]= r_4[2] /*5409*/;
assign r_5[3]= r_4[3] /*5408*/;
assign r_5[4]= r_4[4] /*5407*/;
assign r_5[5]= r_4[5] /*5406*/;
assign r_5[6]= r_4[6] /*5405*/;
assign r_5[7]= r_4[7] /*5404*/;
assign r_5[8]= r_4[8] /*5403*/;
assign r_5[9]= r_4[9] /*5402*/;
assign r_5[10]= r_4[10] /*5401*/;
  assign inv_6[0] = ~div[0] /*5368*/;
  assign inv_6[1] = ~div[1] /*5367*/;
  assign inv_6[2] = ~div[2] /*5366*/;
  assign inv_6[3] = ~div[3] /*5365*/;
  assign inv_6[4] = ~div[4] /*5364*/;
  assign inv_6[5] = ~div[5] /*5363*/;
  assign inv_6[6] = ~div[6] /*5362*/;
  assign inv_6[7] = ~div[7] /*5361*/;
  assign inv_6[8] = ~div[8] /*5360*/;
  assign inv_6[9] = ~div[9] /*5359*/;
  assign inv_6[10] = ~div[10] /*5358*/;
  assign inv_6[11] = ~div[11] /*5357*/;
  assign inv_6[12] = ~div[12] /*5356*/;
  assign inv_6[13] = ~div[13] /*5355*/;
  assign inv_6[14] = ~div[14] /*5354*/;
assign inv_6[15] = oneWire /*5353*/;
  assign _560_ = inv_6[0] ^ r_5[10] /*5351*/;
  assign sum_6[0] = _560_ ^ oneWire /*5350*/;
  assign _561_ = _560_ & oneWire /*5349*/;
  assign _562_ = inv_6[0] & r_5[10] /*5348*/;
  assign _563_ = _561_ | _562_ /*5347*/;
  assign _564_ = inv_6[1] ^ r_5[11] /*5346*/;
  assign sum_6[1] = _564_ ^ _563_ /*5345*/;
  assign _565_ = _564_ & _563_ /*5344*/;
  assign _566_ = inv_6[1] & r_5[11] /*5343*/;
  assign _567_ = _565_ | _566_ /*5342*/;
  assign _568_ = inv_6[2] ^ r_5[12] /*5340*/;
  assign sum_6[2] = _568_ ^ _567_ /*5339*/;
  assign _569_ = _568_ & _567_ /*5338*/;
  assign _570_ = inv_6[2] & r_5[12] /*5337*/;
  assign _571_ = _569_ | _570_ /*5336*/;
  assign _572_ = inv_6[3] ^ r_5[13] /*5334*/;
  assign sum_6[3] = _572_ ^ _571_ /*5333*/;
  assign _573_ = _572_ & _571_ /*5332*/;
  assign _574_ = inv_6[3] & r_5[13] /*5331*/;
  assign _575_ = _573_ | _574_ /*5330*/;
  assign _576_ = inv_6[4] ^ r_5[14] /*5328*/;
  assign sum_6[4] = _576_ ^ _575_ /*5327*/;
  assign _577_ = _576_ & _575_ /*5326*/;
  assign _578_ = inv_6[4] & r_5[14] /*5325*/;
  assign _579_ = _577_ | _578_ /*5324*/;
  assign _580_ = inv_6[5] ^ r_5[15] /*5322*/;
  assign sum_6[5] = _580_ ^ _579_ /*5321*/;
  assign _581_ = _580_ & _579_ /*5320*/;
  assign _582_ = inv_6[5] & r_5[15] /*5319*/;
  assign _583_ = _581_ | _582_ /*5318*/;
  assign _584_ = inv_6[6] ^ r_5[16] /*5316*/;
  assign sum_6[6] = _584_ ^ _583_ /*5315*/;
  assign _585_ = _584_ & _583_ /*5314*/;
  assign _586_ = inv_6[6] & r_5[16] /*5313*/;
  assign _587_ = _585_ | _586_ /*5312*/;
  assign _588_ = inv_6[7] ^ r_5[17] /*5310*/;
  assign sum_6[7] = _588_ ^ _587_ /*5309*/;
  assign _589_ = _588_ & _587_ /*5308*/;
  assign _590_ = inv_6[7] & r_5[17] /*5307*/;
  assign _591_ = _589_ | _590_ /*5306*/;
  assign _592_ = inv_6[8] ^ r_5[18] /*5304*/;
  assign sum_6[8] = _592_ ^ _591_ /*5303*/;
  assign _593_ = _592_ & _591_ /*5302*/;
  assign _594_ = inv_6[8] & r_5[18] /*5301*/;
  assign _595_ = _593_ | _594_ /*5300*/;
  assign _596_ = inv_6[9] ^ r_5[19] /*5298*/;
  assign sum_6[9] = _596_ ^ _595_ /*5297*/;
  assign _597_ = _596_ & _595_ /*5296*/;
  assign _598_ = inv_6[9] & r_5[19] /*5295*/;
  assign _599_ = _597_ | _598_ /*5294*/;
  assign _600_ = inv_6[10] ^ r_5[20] /*5292*/;
  assign sum_6[10] = _600_ ^ _599_ /*5291*/;
  assign _601_ = _600_ & _599_ /*5290*/;
  assign _602_ = inv_6[10] & r_5[20] /*5289*/;
  assign _603_ = _601_ | _602_ /*5288*/;
  assign _604_ = inv_6[11] ^ r_5[21] /*5286*/;
  assign sum_6[11] = _604_ ^ _603_ /*5285*/;
  assign _605_ = _604_ & _603_ /*5284*/;
  assign _606_ = inv_6[11] & r_5[21] /*5283*/;
  assign _607_ = _605_ | _606_ /*5282*/;
  assign _608_ = inv_6[12] ^ r_5[22] /*5280*/;
  assign sum_6[12] = _608_ ^ _607_ /*5279*/;
  assign _609_ = _608_ & _607_ /*5278*/;
  assign _610_ = inv_6[12] & r_5[22] /*5277*/;
  assign _611_ = _609_ | _610_ /*5276*/;
  assign _612_ = inv_6[13] ^ r_5[23] /*5274*/;
  assign sum_6[13] = _612_ ^ _611_ /*5273*/;
  assign _613_ = _612_ & _611_ /*5272*/;
  assign _614_ = inv_6[13] & r_5[23] /*5271*/;
  assign _615_ = _613_ | _614_ /*5270*/;
  assign _616_ = inv_6[14] ^ r_5[24] /*5268*/;
  assign sum_6[14] = _616_ ^ _615_ /*5267*/;
  assign _617_ = _616_ & _615_ /*5266*/;
  assign _618_ = inv_6[14] & r_5[24] /*5265*/;
  assign _619_ = _617_ | _618_ /*5264*/;
  assign _620_ = inv_6[15] ^ r_5[25] /*5262*/;
  assign sum_6[15] = _620_ ^ _619_ /*5261*/;
  assign _621_ = _620_ & _619_ /*5260*/;
  assign _622_ = inv_6[15] & r_5[25] /*5259*/;
  assign _623_ = _621_ | _622_ /*5258*/;
  assign q[10] = ~sum_6[15] /*5269*/;
  assign m_6[0] = r_5[10] /*5268*/;
  assign m_6[1] = r_5[11] /*5267*/;
  assign m_6[2] = r_5[12] /*5266*/;
  assign m_6[3] = r_5[13] /*5265*/;
  assign m_6[4] = r_5[14] /*5264*/;
  assign m_6[5] = r_5[15] /*5263*/;
  assign m_6[6] = r_5[16] /*5262*/;
  assign m_6[7] = r_5[17] /*5261*/;
  assign m_6[8] = r_5[18] /*5260*/;
  assign m_6[9] = r_5[19] /*5259*/;
  assign m_6[10] = r_5[20] /*5258*/;
  assign m_6[11] = r_5[21] /*5257*/;
  assign m_6[12] = r_5[22] /*5256*/;
  assign m_6[13] = r_5[23] /*5255*/;
  assign m_6[14] = r_5[24] /*5254*/;
  assign m_6[15] = r_5[25] /*5253*/;
  assign _624_ = ~q[10] /*5251*/;
  assign _625_ = sum_6[0] & q[10] /*5250*/;
  assign _626_ = m_6[0] & _624_ /*5249*/;
  assign r_6[10] = _626_ | _625_ /*5248*/;
  assign _627_ = ~q[10] /*5247*/;
  assign _628_ = sum_6[1] & q[10] /*5246*/;
  assign _629_ = m_6[1] & _627_ /*5245*/;
  assign r_6[11] = _629_ | _628_ /*5244*/;
  assign _630_ = ~q[10] /*5243*/;
  assign _631_ = sum_6[2] & q[10] /*5242*/;
  assign _632_ = m_6[2] & _630_ /*5241*/;
  assign r_6[12] = _632_ | _631_ /*5240*/;
  assign _633_ = ~q[10] /*5239*/;
  assign _634_ = sum_6[3] & q[10] /*5238*/;
  assign _635_ = m_6[3] & _633_ /*5237*/;
  assign r_6[13] = _635_ | _634_ /*5236*/;
  assign _636_ = ~q[10] /*5235*/;
  assign _637_ = sum_6[4] & q[10] /*5234*/;
  assign _638_ = m_6[4] & _636_ /*5233*/;
  assign r_6[14] = _638_ | _637_ /*5232*/;
  assign _639_ = ~q[10] /*5231*/;
  assign _640_ = sum_6[5] & q[10] /*5230*/;
  assign _641_ = m_6[5] & _639_ /*5229*/;
  assign r_6[15] = _641_ | _640_ /*5228*/;
  assign _642_ = ~q[10] /*5227*/;
  assign _643_ = sum_6[6] & q[10] /*5226*/;
  assign _644_ = m_6[6] & _642_ /*5225*/;
  assign r_6[16] = _644_ | _643_ /*5224*/;
  assign _645_ = ~q[10] /*5223*/;
  assign _646_ = sum_6[7] & q[10] /*5222*/;
  assign _647_ = m_6[7] & _645_ /*5221*/;
  assign r_6[17] = _647_ | _646_ /*5220*/;
  assign _648_ = ~q[10] /*5219*/;
  assign _649_ = sum_6[8] & q[10] /*5218*/;
  assign _650_ = m_6[8] & _648_ /*5217*/;
  assign r_6[18] = _650_ | _649_ /*5216*/;
  assign _651_ = ~q[10] /*5215*/;
  assign _652_ = sum_6[9] & q[10] /*5214*/;
  assign _653_ = m_6[9] & _651_ /*5213*/;
  assign r_6[19] = _653_ | _652_ /*5212*/;
  assign _654_ = ~q[10] /*5211*/;
  assign _655_ = sum_6[10] & q[10] /*5210*/;
  assign _656_ = m_6[10] & _654_ /*5209*/;
  assign r_6[20] = _656_ | _655_ /*5208*/;
  assign _657_ = ~q[10] /*5207*/;
  assign _658_ = sum_6[11] & q[10] /*5206*/;
  assign _659_ = m_6[11] & _657_ /*5205*/;
  assign r_6[21] = _659_ | _658_ /*5204*/;
  assign _660_ = ~q[10] /*5203*/;
  assign _661_ = sum_6[12] & q[10] /*5202*/;
  assign _662_ = m_6[12] & _660_ /*5201*/;
  assign r_6[22] = _662_ | _661_ /*5200*/;
  assign _663_ = ~q[10] /*5199*/;
  assign _664_ = sum_6[13] & q[10] /*5198*/;
  assign _665_ = m_6[13] & _663_ /*5197*/;
  assign r_6[23] = _665_ | _664_ /*5196*/;
  assign _666_ = ~q[10] /*5195*/;
  assign _667_ = sum_6[14] & q[10] /*5194*/;
  assign _668_ = m_6[14] & _666_ /*5193*/;
  assign r_6[24] = _668_ | _667_ /*5192*/;
  assign _669_ = ~q[10] /*5191*/;
  assign _670_ = sum_6[15] & q[10] /*5190*/;
  assign _671_ = m_6[15] & _669_ /*5189*/;
  assign r_6[25] = _671_ | _670_ /*5188*/;
assign r_6[0]= r_5[0] /*5187*/;
assign r_6[1]= r_5[1] /*5186*/;
assign r_6[2]= r_5[2] /*5185*/;
assign r_6[3]= r_5[3] /*5184*/;
assign r_6[4]= r_5[4] /*5183*/;
assign r_6[5]= r_5[5] /*5182*/;
assign r_6[6]= r_5[6] /*5181*/;
assign r_6[7]= r_5[7] /*5180*/;
assign r_6[8]= r_5[8] /*5179*/;
assign r_6[9]= r_5[9] /*5178*/;
  assign inv_7[0] = ~div[0] /*5144*/;
  assign inv_7[1] = ~div[1] /*5143*/;
  assign inv_7[2] = ~div[2] /*5142*/;
  assign inv_7[3] = ~div[3] /*5141*/;
  assign inv_7[4] = ~div[4] /*5140*/;
  assign inv_7[5] = ~div[5] /*5139*/;
  assign inv_7[6] = ~div[6] /*5138*/;
  assign inv_7[7] = ~div[7] /*5137*/;
  assign inv_7[8] = ~div[8] /*5136*/;
  assign inv_7[9] = ~div[9] /*5135*/;
  assign inv_7[10] = ~div[10] /*5134*/;
  assign inv_7[11] = ~div[11] /*5133*/;
  assign inv_7[12] = ~div[12] /*5132*/;
  assign inv_7[13] = ~div[13] /*5131*/;
  assign inv_7[14] = ~div[14] /*5130*/;
assign inv_7[15] = oneWire /*5129*/;
  assign _672_ = inv_7[0] ^ r_6[9] /*5127*/;
  assign sum_7[0] = _672_ ^ oneWire /*5126*/;
  assign _673_ = _672_ & oneWire /*5125*/;
  assign _674_ = inv_7[0] & r_6[9] /*5124*/;
  assign _675_ = _673_ | _674_ /*5123*/;
  assign _676_ = inv_7[1] ^ r_6[10] /*5122*/;
  assign sum_7[1] = _676_ ^ _675_ /*5121*/;
  assign _677_ = _676_ & _675_ /*5120*/;
  assign _678_ = inv_7[1] & r_6[10] /*5119*/;
  assign _679_ = _677_ | _678_ /*5118*/;
  assign _680_ = inv_7[2] ^ r_6[11] /*5116*/;
  assign sum_7[2] = _680_ ^ _679_ /*5115*/;
  assign _681_ = _680_ & _679_ /*5114*/;
  assign _682_ = inv_7[2] & r_6[11] /*5113*/;
  assign _683_ = _681_ | _682_ /*5112*/;
  assign _684_ = inv_7[3] ^ r_6[12] /*5110*/;
  assign sum_7[3] = _684_ ^ _683_ /*5109*/;
  assign _685_ = _684_ & _683_ /*5108*/;
  assign _686_ = inv_7[3] & r_6[12] /*5107*/;
  assign _687_ = _685_ | _686_ /*5106*/;
  assign _688_ = inv_7[4] ^ r_6[13] /*5104*/;
  assign sum_7[4] = _688_ ^ _687_ /*5103*/;
  assign _689_ = _688_ & _687_ /*5102*/;
  assign _690_ = inv_7[4] & r_6[13] /*5101*/;
  assign _691_ = _689_ | _690_ /*5100*/;
  assign _692_ = inv_7[5] ^ r_6[14] /*5098*/;
  assign sum_7[5] = _692_ ^ _691_ /*5097*/;
  assign _693_ = _692_ & _691_ /*5096*/;
  assign _694_ = inv_7[5] & r_6[14] /*5095*/;
  assign _695_ = _693_ | _694_ /*5094*/;
  assign _696_ = inv_7[6] ^ r_6[15] /*5092*/;
  assign sum_7[6] = _696_ ^ _695_ /*5091*/;
  assign _697_ = _696_ & _695_ /*5090*/;
  assign _698_ = inv_7[6] & r_6[15] /*5089*/;
  assign _699_ = _697_ | _698_ /*5088*/;
  assign _700_ = inv_7[7] ^ r_6[16] /*5086*/;
  assign sum_7[7] = _700_ ^ _699_ /*5085*/;
  assign _701_ = _700_ & _699_ /*5084*/;
  assign _702_ = inv_7[7] & r_6[16] /*5083*/;
  assign _703_ = _701_ | _702_ /*5082*/;
  assign _704_ = inv_7[8] ^ r_6[17] /*5080*/;
  assign sum_7[8] = _704_ ^ _703_ /*5079*/;
  assign _705_ = _704_ & _703_ /*5078*/;
  assign _706_ = inv_7[8] & r_6[17] /*5077*/;
  assign _707_ = _705_ | _706_ /*5076*/;
  assign _708_ = inv_7[9] ^ r_6[18] /*5074*/;
  assign sum_7[9] = _708_ ^ _707_ /*5073*/;
  assign _709_ = _708_ & _707_ /*5072*/;
  assign _710_ = inv_7[9] & r_6[18] /*5071*/;
  assign _711_ = _709_ | _710_ /*5070*/;
  assign _712_ = inv_7[10] ^ r_6[19] /*5068*/;
  assign sum_7[10] = _712_ ^ _711_ /*5067*/;
  assign _713_ = _712_ & _711_ /*5066*/;
  assign _714_ = inv_7[10] & r_6[19] /*5065*/;
  assign _715_ = _713_ | _714_ /*5064*/;
  assign _716_ = inv_7[11] ^ r_6[20] /*5062*/;
  assign sum_7[11] = _716_ ^ _715_ /*5061*/;
  assign _717_ = _716_ & _715_ /*5060*/;
  assign _718_ = inv_7[11] & r_6[20] /*5059*/;
  assign _719_ = _717_ | _718_ /*5058*/;
  assign _720_ = inv_7[12] ^ r_6[21] /*5056*/;
  assign sum_7[12] = _720_ ^ _719_ /*5055*/;
  assign _721_ = _720_ & _719_ /*5054*/;
  assign _722_ = inv_7[12] & r_6[21] /*5053*/;
  assign _723_ = _721_ | _722_ /*5052*/;
  assign _724_ = inv_7[13] ^ r_6[22] /*5050*/;
  assign sum_7[13] = _724_ ^ _723_ /*5049*/;
  assign _725_ = _724_ & _723_ /*5048*/;
  assign _726_ = inv_7[13] & r_6[22] /*5047*/;
  assign _727_ = _725_ | _726_ /*5046*/;
  assign _728_ = inv_7[14] ^ r_6[23] /*5044*/;
  assign sum_7[14] = _728_ ^ _727_ /*5043*/;
  assign _729_ = _728_ & _727_ /*5042*/;
  assign _730_ = inv_7[14] & r_6[23] /*5041*/;
  assign _731_ = _729_ | _730_ /*5040*/;
  assign _732_ = inv_7[15] ^ r_6[24] /*5038*/;
  assign sum_7[15] = _732_ ^ _731_ /*5037*/;
  assign _733_ = _732_ & _731_ /*5036*/;
  assign _734_ = inv_7[15] & r_6[24] /*5035*/;
  assign _735_ = _733_ | _734_ /*5034*/;
  assign q[9] = ~sum_7[15] /*5045*/;
  assign m_7[0] = r_6[9] /*5044*/;
  assign m_7[1] = r_6[10] /*5043*/;
  assign m_7[2] = r_6[11] /*5042*/;
  assign m_7[3] = r_6[12] /*5041*/;
  assign m_7[4] = r_6[13] /*5040*/;
  assign m_7[5] = r_6[14] /*5039*/;
  assign m_7[6] = r_6[15] /*5038*/;
  assign m_7[7] = r_6[16] /*5037*/;
  assign m_7[8] = r_6[17] /*5036*/;
  assign m_7[9] = r_6[18] /*5035*/;
  assign m_7[10] = r_6[19] /*5034*/;
  assign m_7[11] = r_6[20] /*5033*/;
  assign m_7[12] = r_6[21] /*5032*/;
  assign m_7[13] = r_6[22] /*5031*/;
  assign m_7[14] = r_6[23] /*5030*/;
  assign m_7[15] = r_6[24] /*5029*/;
  assign _736_ = ~q[9] /*5027*/;
  assign _737_ = sum_7[0] & q[9] /*5026*/;
  assign _738_ = m_7[0] & _736_ /*5025*/;
  assign r_7[9] = _738_ | _737_ /*5024*/;
  assign _739_ = ~q[9] /*5023*/;
  assign _740_ = sum_7[1] & q[9] /*5022*/;
  assign _741_ = m_7[1] & _739_ /*5021*/;
  assign r_7[10] = _741_ | _740_ /*5020*/;
  assign _742_ = ~q[9] /*5019*/;
  assign _743_ = sum_7[2] & q[9] /*5018*/;
  assign _744_ = m_7[2] & _742_ /*5017*/;
  assign r_7[11] = _744_ | _743_ /*5016*/;
  assign _745_ = ~q[9] /*5015*/;
  assign _746_ = sum_7[3] & q[9] /*5014*/;
  assign _747_ = m_7[3] & _745_ /*5013*/;
  assign r_7[12] = _747_ | _746_ /*5012*/;
  assign _748_ = ~q[9] /*5011*/;
  assign _749_ = sum_7[4] & q[9] /*5010*/;
  assign _750_ = m_7[4] & _748_ /*5009*/;
  assign r_7[13] = _750_ | _749_ /*5008*/;
  assign _751_ = ~q[9] /*5007*/;
  assign _752_ = sum_7[5] & q[9] /*5006*/;
  assign _753_ = m_7[5] & _751_ /*5005*/;
  assign r_7[14] = _753_ | _752_ /*5004*/;
  assign _754_ = ~q[9] /*5003*/;
  assign _755_ = sum_7[6] & q[9] /*5002*/;
  assign _756_ = m_7[6] & _754_ /*5001*/;
  assign r_7[15] = _756_ | _755_ /*5000*/;
  assign _757_ = ~q[9] /*4999*/;
  assign _758_ = sum_7[7] & q[9] /*4998*/;
  assign _759_ = m_7[7] & _757_ /*4997*/;
  assign r_7[16] = _759_ | _758_ /*4996*/;
  assign _760_ = ~q[9] /*4995*/;
  assign _761_ = sum_7[8] & q[9] /*4994*/;
  assign _762_ = m_7[8] & _760_ /*4993*/;
  assign r_7[17] = _762_ | _761_ /*4992*/;
  assign _763_ = ~q[9] /*4991*/;
  assign _764_ = sum_7[9] & q[9] /*4990*/;
  assign _765_ = m_7[9] & _763_ /*4989*/;
  assign r_7[18] = _765_ | _764_ /*4988*/;
  assign _766_ = ~q[9] /*4987*/;
  assign _767_ = sum_7[10] & q[9] /*4986*/;
  assign _768_ = m_7[10] & _766_ /*4985*/;
  assign r_7[19] = _768_ | _767_ /*4984*/;
  assign _769_ = ~q[9] /*4983*/;
  assign _770_ = sum_7[11] & q[9] /*4982*/;
  assign _771_ = m_7[11] & _769_ /*4981*/;
  assign r_7[20] = _771_ | _770_ /*4980*/;
  assign _772_ = ~q[9] /*4979*/;
  assign _773_ = sum_7[12] & q[9] /*4978*/;
  assign _774_ = m_7[12] & _772_ /*4977*/;
  assign r_7[21] = _774_ | _773_ /*4976*/;
  assign _775_ = ~q[9] /*4975*/;
  assign _776_ = sum_7[13] & q[9] /*4974*/;
  assign _777_ = m_7[13] & _775_ /*4973*/;
  assign r_7[22] = _777_ | _776_ /*4972*/;
  assign _778_ = ~q[9] /*4971*/;
  assign _779_ = sum_7[14] & q[9] /*4970*/;
  assign _780_ = m_7[14] & _778_ /*4969*/;
  assign r_7[23] = _780_ | _779_ /*4968*/;
  assign _781_ = ~q[9] /*4967*/;
  assign _782_ = sum_7[15] & q[9] /*4966*/;
  assign _783_ = m_7[15] & _781_ /*4965*/;
  assign r_7[24] = _783_ | _782_ /*4964*/;
assign r_7[0]= r_6[0] /*4963*/;
assign r_7[1]= r_6[1] /*4962*/;
assign r_7[2]= r_6[2] /*4961*/;
assign r_7[3]= r_6[3] /*4960*/;
assign r_7[4]= r_6[4] /*4959*/;
assign r_7[5]= r_6[5] /*4958*/;
assign r_7[6]= r_6[6] /*4957*/;
assign r_7[7]= r_6[7] /*4956*/;
assign r_7[8]= r_6[8] /*4955*/;
  assign inv_8[0] = ~div[0] /*4920*/;
  assign inv_8[1] = ~div[1] /*4919*/;
  assign inv_8[2] = ~div[2] /*4918*/;
  assign inv_8[3] = ~div[3] /*4917*/;
  assign inv_8[4] = ~div[4] /*4916*/;
  assign inv_8[5] = ~div[5] /*4915*/;
  assign inv_8[6] = ~div[6] /*4914*/;
  assign inv_8[7] = ~div[7] /*4913*/;
  assign inv_8[8] = ~div[8] /*4912*/;
  assign inv_8[9] = ~div[9] /*4911*/;
  assign inv_8[10] = ~div[10] /*4910*/;
  assign inv_8[11] = ~div[11] /*4909*/;
  assign inv_8[12] = ~div[12] /*4908*/;
  assign inv_8[13] = ~div[13] /*4907*/;
  assign inv_8[14] = ~div[14] /*4906*/;
assign inv_8[15] = oneWire /*4905*/;
  assign _784_ = inv_8[0] ^ r_7[8] /*4903*/;
  assign sum_8[0] = _784_ ^ oneWire /*4902*/;
  assign _785_ = _784_ & oneWire /*4901*/;
  assign _786_ = inv_8[0] & r_7[8] /*4900*/;
  assign _787_ = _785_ | _786_ /*4899*/;
  assign _788_ = inv_8[1] ^ r_7[9] /*4898*/;
  assign sum_8[1] = _788_ ^ _787_ /*4897*/;
  assign _789_ = _788_ & _787_ /*4896*/;
  assign _790_ = inv_8[1] & r_7[9] /*4895*/;
  assign _791_ = _789_ | _790_ /*4894*/;
  assign _792_ = inv_8[2] ^ r_7[10] /*4892*/;
  assign sum_8[2] = _792_ ^ _791_ /*4891*/;
  assign _793_ = _792_ & _791_ /*4890*/;
  assign _794_ = inv_8[2] & r_7[10] /*4889*/;
  assign _795_ = _793_ | _794_ /*4888*/;
  assign _796_ = inv_8[3] ^ r_7[11] /*4886*/;
  assign sum_8[3] = _796_ ^ _795_ /*4885*/;
  assign _797_ = _796_ & _795_ /*4884*/;
  assign _798_ = inv_8[3] & r_7[11] /*4883*/;
  assign _799_ = _797_ | _798_ /*4882*/;
  assign _800_ = inv_8[4] ^ r_7[12] /*4880*/;
  assign sum_8[4] = _800_ ^ _799_ /*4879*/;
  assign _801_ = _800_ & _799_ /*4878*/;
  assign _802_ = inv_8[4] & r_7[12] /*4877*/;
  assign _803_ = _801_ | _802_ /*4876*/;
  assign _804_ = inv_8[5] ^ r_7[13] /*4874*/;
  assign sum_8[5] = _804_ ^ _803_ /*4873*/;
  assign _805_ = _804_ & _803_ /*4872*/;
  assign _806_ = inv_8[5] & r_7[13] /*4871*/;
  assign _807_ = _805_ | _806_ /*4870*/;
  assign _808_ = inv_8[6] ^ r_7[14] /*4868*/;
  assign sum_8[6] = _808_ ^ _807_ /*4867*/;
  assign _809_ = _808_ & _807_ /*4866*/;
  assign _810_ = inv_8[6] & r_7[14] /*4865*/;
  assign _811_ = _809_ | _810_ /*4864*/;
  assign _812_ = inv_8[7] ^ r_7[15] /*4862*/;
  assign sum_8[7] = _812_ ^ _811_ /*4861*/;
  assign _813_ = _812_ & _811_ /*4860*/;
  assign _814_ = inv_8[7] & r_7[15] /*4859*/;
  assign _815_ = _813_ | _814_ /*4858*/;
  assign _816_ = inv_8[8] ^ r_7[16] /*4856*/;
  assign sum_8[8] = _816_ ^ _815_ /*4855*/;
  assign _817_ = _816_ & _815_ /*4854*/;
  assign _818_ = inv_8[8] & r_7[16] /*4853*/;
  assign _819_ = _817_ | _818_ /*4852*/;
  assign _820_ = inv_8[9] ^ r_7[17] /*4850*/;
  assign sum_8[9] = _820_ ^ _819_ /*4849*/;
  assign _821_ = _820_ & _819_ /*4848*/;
  assign _822_ = inv_8[9] & r_7[17] /*4847*/;
  assign _823_ = _821_ | _822_ /*4846*/;
  assign _824_ = inv_8[10] ^ r_7[18] /*4844*/;
  assign sum_8[10] = _824_ ^ _823_ /*4843*/;
  assign _825_ = _824_ & _823_ /*4842*/;
  assign _826_ = inv_8[10] & r_7[18] /*4841*/;
  assign _827_ = _825_ | _826_ /*4840*/;
  assign _828_ = inv_8[11] ^ r_7[19] /*4838*/;
  assign sum_8[11] = _828_ ^ _827_ /*4837*/;
  assign _829_ = _828_ & _827_ /*4836*/;
  assign _830_ = inv_8[11] & r_7[19] /*4835*/;
  assign _831_ = _829_ | _830_ /*4834*/;
  assign _832_ = inv_8[12] ^ r_7[20] /*4832*/;
  assign sum_8[12] = _832_ ^ _831_ /*4831*/;
  assign _833_ = _832_ & _831_ /*4830*/;
  assign _834_ = inv_8[12] & r_7[20] /*4829*/;
  assign _835_ = _833_ | _834_ /*4828*/;
  assign _836_ = inv_8[13] ^ r_7[21] /*4826*/;
  assign sum_8[13] = _836_ ^ _835_ /*4825*/;
  assign _837_ = _836_ & _835_ /*4824*/;
  assign _838_ = inv_8[13] & r_7[21] /*4823*/;
  assign _839_ = _837_ | _838_ /*4822*/;
  assign _840_ = inv_8[14] ^ r_7[22] /*4820*/;
  assign sum_8[14] = _840_ ^ _839_ /*4819*/;
  assign _841_ = _840_ & _839_ /*4818*/;
  assign _842_ = inv_8[14] & r_7[22] /*4817*/;
  assign _843_ = _841_ | _842_ /*4816*/;
  assign _844_ = inv_8[15] ^ r_7[23] /*4814*/;
  assign sum_8[15] = _844_ ^ _843_ /*4813*/;
  assign _845_ = _844_ & _843_ /*4812*/;
  assign _846_ = inv_8[15] & r_7[23] /*4811*/;
  assign _847_ = _845_ | _846_ /*4810*/;
  assign q[8] = ~sum_8[15] /*4821*/;
  assign m_8[0] = r_7[8] /*4820*/;
  assign m_8[1] = r_7[9] /*4819*/;
  assign m_8[2] = r_7[10] /*4818*/;
  assign m_8[3] = r_7[11] /*4817*/;
  assign m_8[4] = r_7[12] /*4816*/;
  assign m_8[5] = r_7[13] /*4815*/;
  assign m_8[6] = r_7[14] /*4814*/;
  assign m_8[7] = r_7[15] /*4813*/;
  assign m_8[8] = r_7[16] /*4812*/;
  assign m_8[9] = r_7[17] /*4811*/;
  assign m_8[10] = r_7[18] /*4810*/;
  assign m_8[11] = r_7[19] /*4809*/;
  assign m_8[12] = r_7[20] /*4808*/;
  assign m_8[13] = r_7[21] /*4807*/;
  assign m_8[14] = r_7[22] /*4806*/;
  assign m_8[15] = r_7[23] /*4805*/;
  assign _848_ = ~q[8] /*4803*/;
  assign _849_ = sum_8[0] & q[8] /*4802*/;
  assign _850_ = m_8[0] & _848_ /*4801*/;
  assign r_8[8] = _850_ | _849_ /*4800*/;
  assign _851_ = ~q[8] /*4799*/;
  assign _852_ = sum_8[1] & q[8] /*4798*/;
  assign _853_ = m_8[1] & _851_ /*4797*/;
  assign r_8[9] = _853_ | _852_ /*4796*/;
  assign _854_ = ~q[8] /*4795*/;
  assign _855_ = sum_8[2] & q[8] /*4794*/;
  assign _856_ = m_8[2] & _854_ /*4793*/;
  assign r_8[10] = _856_ | _855_ /*4792*/;
  assign _857_ = ~q[8] /*4791*/;
  assign _858_ = sum_8[3] & q[8] /*4790*/;
  assign _859_ = m_8[3] & _857_ /*4789*/;
  assign r_8[11] = _859_ | _858_ /*4788*/;
  assign _860_ = ~q[8] /*4787*/;
  assign _861_ = sum_8[4] & q[8] /*4786*/;
  assign _862_ = m_8[4] & _860_ /*4785*/;
  assign r_8[12] = _862_ | _861_ /*4784*/;
  assign _863_ = ~q[8] /*4783*/;
  assign _864_ = sum_8[5] & q[8] /*4782*/;
  assign _865_ = m_8[5] & _863_ /*4781*/;
  assign r_8[13] = _865_ | _864_ /*4780*/;
  assign _866_ = ~q[8] /*4779*/;
  assign _867_ = sum_8[6] & q[8] /*4778*/;
  assign _868_ = m_8[6] & _866_ /*4777*/;
  assign r_8[14] = _868_ | _867_ /*4776*/;
  assign _869_ = ~q[8] /*4775*/;
  assign _870_ = sum_8[7] & q[8] /*4774*/;
  assign _871_ = m_8[7] & _869_ /*4773*/;
  assign r_8[15] = _871_ | _870_ /*4772*/;
  assign _872_ = ~q[8] /*4771*/;
  assign _873_ = sum_8[8] & q[8] /*4770*/;
  assign _874_ = m_8[8] & _872_ /*4769*/;
  assign r_8[16] = _874_ | _873_ /*4768*/;
  assign _875_ = ~q[8] /*4767*/;
  assign _876_ = sum_8[9] & q[8] /*4766*/;
  assign _877_ = m_8[9] & _875_ /*4765*/;
  assign r_8[17] = _877_ | _876_ /*4764*/;
  assign _878_ = ~q[8] /*4763*/;
  assign _879_ = sum_8[10] & q[8] /*4762*/;
  assign _880_ = m_8[10] & _878_ /*4761*/;
  assign r_8[18] = _880_ | _879_ /*4760*/;
  assign _881_ = ~q[8] /*4759*/;
  assign _882_ = sum_8[11] & q[8] /*4758*/;
  assign _883_ = m_8[11] & _881_ /*4757*/;
  assign r_8[19] = _883_ | _882_ /*4756*/;
  assign _884_ = ~q[8] /*4755*/;
  assign _885_ = sum_8[12] & q[8] /*4754*/;
  assign _886_ = m_8[12] & _884_ /*4753*/;
  assign r_8[20] = _886_ | _885_ /*4752*/;
  assign _887_ = ~q[8] /*4751*/;
  assign _888_ = sum_8[13] & q[8] /*4750*/;
  assign _889_ = m_8[13] & _887_ /*4749*/;
  assign r_8[21] = _889_ | _888_ /*4748*/;
  assign _890_ = ~q[8] /*4747*/;
  assign _891_ = sum_8[14] & q[8] /*4746*/;
  assign _892_ = m_8[14] & _890_ /*4745*/;
  assign r_8[22] = _892_ | _891_ /*4744*/;
  assign _893_ = ~q[8] /*4743*/;
  assign _894_ = sum_8[15] & q[8] /*4742*/;
  assign _895_ = m_8[15] & _893_ /*4741*/;
  assign r_8[23] = _895_ | _894_ /*4740*/;
assign r_8[0]= r_7[0] /*4739*/;
assign r_8[1]= r_7[1] /*4738*/;
assign r_8[2]= r_7[2] /*4737*/;
assign r_8[3]= r_7[3] /*4736*/;
assign r_8[4]= r_7[4] /*4735*/;
assign r_8[5]= r_7[5] /*4734*/;
assign r_8[6]= r_7[6] /*4733*/;
assign r_8[7]= r_7[7] /*4732*/;
  assign inv_9[0] = ~div[0] /*4696*/;
  assign inv_9[1] = ~div[1] /*4695*/;
  assign inv_9[2] = ~div[2] /*4694*/;
  assign inv_9[3] = ~div[3] /*4693*/;
  assign inv_9[4] = ~div[4] /*4692*/;
  assign inv_9[5] = ~div[5] /*4691*/;
  assign inv_9[6] = ~div[6] /*4690*/;
  assign inv_9[7] = ~div[7] /*4689*/;
  assign inv_9[8] = ~div[8] /*4688*/;
  assign inv_9[9] = ~div[9] /*4687*/;
  assign inv_9[10] = ~div[10] /*4686*/;
  assign inv_9[11] = ~div[11] /*4685*/;
  assign inv_9[12] = ~div[12] /*4684*/;
  assign inv_9[13] = ~div[13] /*4683*/;
  assign inv_9[14] = ~div[14] /*4682*/;
assign inv_9[15] = oneWire /*4681*/;
  assign _896_ = inv_9[0] ^ r_8[7] /*4679*/;
  assign sum_9[0] = _896_ ^ oneWire /*4678*/;
  assign _897_ = _896_ & oneWire /*4677*/;
  assign _898_ = inv_9[0] & r_8[7] /*4676*/;
  assign _899_ = _897_ | _898_ /*4675*/;
  assign _900_ = inv_9[1] ^ r_8[8] /*4674*/;
  assign sum_9[1] = _900_ ^ _899_ /*4673*/;
  assign _901_ = _900_ & _899_ /*4672*/;
  assign _902_ = inv_9[1] & r_8[8] /*4671*/;
  assign _903_ = _901_ | _902_ /*4670*/;
  assign _904_ = inv_9[2] ^ r_8[9] /*4668*/;
  assign sum_9[2] = _904_ ^ _903_ /*4667*/;
  assign _905_ = _904_ & _903_ /*4666*/;
  assign _906_ = inv_9[2] & r_8[9] /*4665*/;
  assign _907_ = _905_ | _906_ /*4664*/;
  assign _908_ = inv_9[3] ^ r_8[10] /*4662*/;
  assign sum_9[3] = _908_ ^ _907_ /*4661*/;
  assign _909_ = _908_ & _907_ /*4660*/;
  assign _910_ = inv_9[3] & r_8[10] /*4659*/;
  assign _911_ = _909_ | _910_ /*4658*/;
  assign _912_ = inv_9[4] ^ r_8[11] /*4656*/;
  assign sum_9[4] = _912_ ^ _911_ /*4655*/;
  assign _913_ = _912_ & _911_ /*4654*/;
  assign _914_ = inv_9[4] & r_8[11] /*4653*/;
  assign _915_ = _913_ | _914_ /*4652*/;
  assign _916_ = inv_9[5] ^ r_8[12] /*4650*/;
  assign sum_9[5] = _916_ ^ _915_ /*4649*/;
  assign _917_ = _916_ & _915_ /*4648*/;
  assign _918_ = inv_9[5] & r_8[12] /*4647*/;
  assign _919_ = _917_ | _918_ /*4646*/;
  assign _920_ = inv_9[6] ^ r_8[13] /*4644*/;
  assign sum_9[6] = _920_ ^ _919_ /*4643*/;
  assign _921_ = _920_ & _919_ /*4642*/;
  assign _922_ = inv_9[6] & r_8[13] /*4641*/;
  assign _923_ = _921_ | _922_ /*4640*/;
  assign _924_ = inv_9[7] ^ r_8[14] /*4638*/;
  assign sum_9[7] = _924_ ^ _923_ /*4637*/;
  assign _925_ = _924_ & _923_ /*4636*/;
  assign _926_ = inv_9[7] & r_8[14] /*4635*/;
  assign _927_ = _925_ | _926_ /*4634*/;
  assign _928_ = inv_9[8] ^ r_8[15] /*4632*/;
  assign sum_9[8] = _928_ ^ _927_ /*4631*/;
  assign _929_ = _928_ & _927_ /*4630*/;
  assign _930_ = inv_9[8] & r_8[15] /*4629*/;
  assign _931_ = _929_ | _930_ /*4628*/;
  assign _932_ = inv_9[9] ^ r_8[16] /*4626*/;
  assign sum_9[9] = _932_ ^ _931_ /*4625*/;
  assign _933_ = _932_ & _931_ /*4624*/;
  assign _934_ = inv_9[9] & r_8[16] /*4623*/;
  assign _935_ = _933_ | _934_ /*4622*/;
  assign _936_ = inv_9[10] ^ r_8[17] /*4620*/;
  assign sum_9[10] = _936_ ^ _935_ /*4619*/;
  assign _937_ = _936_ & _935_ /*4618*/;
  assign _938_ = inv_9[10] & r_8[17] /*4617*/;
  assign _939_ = _937_ | _938_ /*4616*/;
  assign _940_ = inv_9[11] ^ r_8[18] /*4614*/;
  assign sum_9[11] = _940_ ^ _939_ /*4613*/;
  assign _941_ = _940_ & _939_ /*4612*/;
  assign _942_ = inv_9[11] & r_8[18] /*4611*/;
  assign _943_ = _941_ | _942_ /*4610*/;
  assign _944_ = inv_9[12] ^ r_8[19] /*4608*/;
  assign sum_9[12] = _944_ ^ _943_ /*4607*/;
  assign _945_ = _944_ & _943_ /*4606*/;
  assign _946_ = inv_9[12] & r_8[19] /*4605*/;
  assign _947_ = _945_ | _946_ /*4604*/;
  assign _948_ = inv_9[13] ^ r_8[20] /*4602*/;
  assign sum_9[13] = _948_ ^ _947_ /*4601*/;
  assign _949_ = _948_ & _947_ /*4600*/;
  assign _950_ = inv_9[13] & r_8[20] /*4599*/;
  assign _951_ = _949_ | _950_ /*4598*/;
  assign _952_ = inv_9[14] ^ r_8[21] /*4596*/;
  assign sum_9[14] = _952_ ^ _951_ /*4595*/;
  assign _953_ = _952_ & _951_ /*4594*/;
  assign _954_ = inv_9[14] & r_8[21] /*4593*/;
  assign _955_ = _953_ | _954_ /*4592*/;
  assign _956_ = inv_9[15] ^ r_8[22] /*4590*/;
  assign sum_9[15] = _956_ ^ _955_ /*4589*/;
  assign _957_ = _956_ & _955_ /*4588*/;
  assign _958_ = inv_9[15] & r_8[22] /*4587*/;
  assign _959_ = _957_ | _958_ /*4586*/;
  assign q[7] = ~sum_9[15] /*4597*/;
  assign m_9[0] = r_8[7] /*4596*/;
  assign m_9[1] = r_8[8] /*4595*/;
  assign m_9[2] = r_8[9] /*4594*/;
  assign m_9[3] = r_8[10] /*4593*/;
  assign m_9[4] = r_8[11] /*4592*/;
  assign m_9[5] = r_8[12] /*4591*/;
  assign m_9[6] = r_8[13] /*4590*/;
  assign m_9[7] = r_8[14] /*4589*/;
  assign m_9[8] = r_8[15] /*4588*/;
  assign m_9[9] = r_8[16] /*4587*/;
  assign m_9[10] = r_8[17] /*4586*/;
  assign m_9[11] = r_8[18] /*4585*/;
  assign m_9[12] = r_8[19] /*4584*/;
  assign m_9[13] = r_8[20] /*4583*/;
  assign m_9[14] = r_8[21] /*4582*/;
  assign m_9[15] = r_8[22] /*4581*/;
  assign _960_ = ~q[7] /*4579*/;
  assign _961_ = sum_9[0] & q[7] /*4578*/;
  assign _962_ = m_9[0] & _960_ /*4577*/;
  assign r_9[7] = _962_ | _961_ /*4576*/;
  assign _963_ = ~q[7] /*4575*/;
  assign _964_ = sum_9[1] & q[7] /*4574*/;
  assign _965_ = m_9[1] & _963_ /*4573*/;
  assign r_9[8] = _965_ | _964_ /*4572*/;
  assign _966_ = ~q[7] /*4571*/;
  assign _967_ = sum_9[2] & q[7] /*4570*/;
  assign _968_ = m_9[2] & _966_ /*4569*/;
  assign r_9[9] = _968_ | _967_ /*4568*/;
  assign _969_ = ~q[7] /*4567*/;
  assign _970_ = sum_9[3] & q[7] /*4566*/;
  assign _971_ = m_9[3] & _969_ /*4565*/;
  assign r_9[10] = _971_ | _970_ /*4564*/;
  assign _972_ = ~q[7] /*4563*/;
  assign _973_ = sum_9[4] & q[7] /*4562*/;
  assign _974_ = m_9[4] & _972_ /*4561*/;
  assign r_9[11] = _974_ | _973_ /*4560*/;
  assign _975_ = ~q[7] /*4559*/;
  assign _976_ = sum_9[5] & q[7] /*4558*/;
  assign _977_ = m_9[5] & _975_ /*4557*/;
  assign r_9[12] = _977_ | _976_ /*4556*/;
  assign _978_ = ~q[7] /*4555*/;
  assign _979_ = sum_9[6] & q[7] /*4554*/;
  assign _980_ = m_9[6] & _978_ /*4553*/;
  assign r_9[13] = _980_ | _979_ /*4552*/;
  assign _981_ = ~q[7] /*4551*/;
  assign _982_ = sum_9[7] & q[7] /*4550*/;
  assign _983_ = m_9[7] & _981_ /*4549*/;
  assign r_9[14] = _983_ | _982_ /*4548*/;
  assign _984_ = ~q[7] /*4547*/;
  assign _985_ = sum_9[8] & q[7] /*4546*/;
  assign _986_ = m_9[8] & _984_ /*4545*/;
  assign r_9[15] = _986_ | _985_ /*4544*/;
  assign _987_ = ~q[7] /*4543*/;
  assign _988_ = sum_9[9] & q[7] /*4542*/;
  assign _989_ = m_9[9] & _987_ /*4541*/;
  assign r_9[16] = _989_ | _988_ /*4540*/;
  assign _990_ = ~q[7] /*4539*/;
  assign _991_ = sum_9[10] & q[7] /*4538*/;
  assign _992_ = m_9[10] & _990_ /*4537*/;
  assign r_9[17] = _992_ | _991_ /*4536*/;
  assign _993_ = ~q[7] /*4535*/;
  assign _994_ = sum_9[11] & q[7] /*4534*/;
  assign _995_ = m_9[11] & _993_ /*4533*/;
  assign r_9[18] = _995_ | _994_ /*4532*/;
  assign _996_ = ~q[7] /*4531*/;
  assign _997_ = sum_9[12] & q[7] /*4530*/;
  assign _998_ = m_9[12] & _996_ /*4529*/;
  assign r_9[19] = _998_ | _997_ /*4528*/;
  assign _999_ = ~q[7] /*4527*/;
  assign _1000_ = sum_9[13] & q[7] /*4526*/;
  assign _1001_ = m_9[13] & _999_ /*4525*/;
  assign r_9[20] = _1001_ | _1000_ /*4524*/;
  assign _1002_ = ~q[7] /*4523*/;
  assign _1003_ = sum_9[14] & q[7] /*4522*/;
  assign _1004_ = m_9[14] & _1002_ /*4521*/;
  assign r_9[21] = _1004_ | _1003_ /*4520*/;
  assign _1005_ = ~q[7] /*4519*/;
  assign _1006_ = sum_9[15] & q[7] /*4518*/;
  assign _1007_ = m_9[15] & _1005_ /*4517*/;
  assign r_9[22] = _1007_ | _1006_ /*4516*/;
assign r_9[0]= r_8[0] /*4515*/;
assign r_9[1]= r_8[1] /*4514*/;
assign r_9[2]= r_8[2] /*4513*/;
assign r_9[3]= r_8[3] /*4512*/;
assign r_9[4]= r_8[4] /*4511*/;
assign r_9[5]= r_8[5] /*4510*/;
assign r_9[6]= r_8[6] /*4509*/;
  assign inv_10[0] = ~div[0] /*4472*/;
  assign inv_10[1] = ~div[1] /*4471*/;
  assign inv_10[2] = ~div[2] /*4470*/;
  assign inv_10[3] = ~div[3] /*4469*/;
  assign inv_10[4] = ~div[4] /*4468*/;
  assign inv_10[5] = ~div[5] /*4467*/;
  assign inv_10[6] = ~div[6] /*4466*/;
  assign inv_10[7] = ~div[7] /*4465*/;
  assign inv_10[8] = ~div[8] /*4464*/;
  assign inv_10[9] = ~div[9] /*4463*/;
  assign inv_10[10] = ~div[10] /*4462*/;
  assign inv_10[11] = ~div[11] /*4461*/;
  assign inv_10[12] = ~div[12] /*4460*/;
  assign inv_10[13] = ~div[13] /*4459*/;
  assign inv_10[14] = ~div[14] /*4458*/;
assign inv_10[15] = oneWire /*4457*/;
  assign _1008_ = inv_10[0] ^ r_9[6] /*4455*/;
  assign sum_10[0] = _1008_ ^ oneWire /*4454*/;
  assign _1009_ = _1008_ & oneWire /*4453*/;
  assign _1010_ = inv_10[0] & r_9[6] /*4452*/;
  assign _1011_ = _1009_ | _1010_ /*4451*/;
  assign _1012_ = inv_10[1] ^ r_9[7] /*4450*/;
  assign sum_10[1] = _1012_ ^ _1011_ /*4449*/;
  assign _1013_ = _1012_ & _1011_ /*4448*/;
  assign _1014_ = inv_10[1] & r_9[7] /*4447*/;
  assign _1015_ = _1013_ | _1014_ /*4446*/;
  assign _1016_ = inv_10[2] ^ r_9[8] /*4444*/;
  assign sum_10[2] = _1016_ ^ _1015_ /*4443*/;
  assign _1017_ = _1016_ & _1015_ /*4442*/;
  assign _1018_ = inv_10[2] & r_9[8] /*4441*/;
  assign _1019_ = _1017_ | _1018_ /*4440*/;
  assign _1020_ = inv_10[3] ^ r_9[9] /*4438*/;
  assign sum_10[3] = _1020_ ^ _1019_ /*4437*/;
  assign _1021_ = _1020_ & _1019_ /*4436*/;
  assign _1022_ = inv_10[3] & r_9[9] /*4435*/;
  assign _1023_ = _1021_ | _1022_ /*4434*/;
  assign _1024_ = inv_10[4] ^ r_9[10] /*4432*/;
  assign sum_10[4] = _1024_ ^ _1023_ /*4431*/;
  assign _1025_ = _1024_ & _1023_ /*4430*/;
  assign _1026_ = inv_10[4] & r_9[10] /*4429*/;
  assign _1027_ = _1025_ | _1026_ /*4428*/;
  assign _1028_ = inv_10[5] ^ r_9[11] /*4426*/;
  assign sum_10[5] = _1028_ ^ _1027_ /*4425*/;
  assign _1029_ = _1028_ & _1027_ /*4424*/;
  assign _1030_ = inv_10[5] & r_9[11] /*4423*/;
  assign _1031_ = _1029_ | _1030_ /*4422*/;
  assign _1032_ = inv_10[6] ^ r_9[12] /*4420*/;
  assign sum_10[6] = _1032_ ^ _1031_ /*4419*/;
  assign _1033_ = _1032_ & _1031_ /*4418*/;
  assign _1034_ = inv_10[6] & r_9[12] /*4417*/;
  assign _1035_ = _1033_ | _1034_ /*4416*/;
  assign _1036_ = inv_10[7] ^ r_9[13] /*4414*/;
  assign sum_10[7] = _1036_ ^ _1035_ /*4413*/;
  assign _1037_ = _1036_ & _1035_ /*4412*/;
  assign _1038_ = inv_10[7] & r_9[13] /*4411*/;
  assign _1039_ = _1037_ | _1038_ /*4410*/;
  assign _1040_ = inv_10[8] ^ r_9[14] /*4408*/;
  assign sum_10[8] = _1040_ ^ _1039_ /*4407*/;
  assign _1041_ = _1040_ & _1039_ /*4406*/;
  assign _1042_ = inv_10[8] & r_9[14] /*4405*/;
  assign _1043_ = _1041_ | _1042_ /*4404*/;
  assign _1044_ = inv_10[9] ^ r_9[15] /*4402*/;
  assign sum_10[9] = _1044_ ^ _1043_ /*4401*/;
  assign _1045_ = _1044_ & _1043_ /*4400*/;
  assign _1046_ = inv_10[9] & r_9[15] /*4399*/;
  assign _1047_ = _1045_ | _1046_ /*4398*/;
  assign _1048_ = inv_10[10] ^ r_9[16] /*4396*/;
  assign sum_10[10] = _1048_ ^ _1047_ /*4395*/;
  assign _1049_ = _1048_ & _1047_ /*4394*/;
  assign _1050_ = inv_10[10] & r_9[16] /*4393*/;
  assign _1051_ = _1049_ | _1050_ /*4392*/;
  assign _1052_ = inv_10[11] ^ r_9[17] /*4390*/;
  assign sum_10[11] = _1052_ ^ _1051_ /*4389*/;
  assign _1053_ = _1052_ & _1051_ /*4388*/;
  assign _1054_ = inv_10[11] & r_9[17] /*4387*/;
  assign _1055_ = _1053_ | _1054_ /*4386*/;
  assign _1056_ = inv_10[12] ^ r_9[18] /*4384*/;
  assign sum_10[12] = _1056_ ^ _1055_ /*4383*/;
  assign _1057_ = _1056_ & _1055_ /*4382*/;
  assign _1058_ = inv_10[12] & r_9[18] /*4381*/;
  assign _1059_ = _1057_ | _1058_ /*4380*/;
  assign _1060_ = inv_10[13] ^ r_9[19] /*4378*/;
  assign sum_10[13] = _1060_ ^ _1059_ /*4377*/;
  assign _1061_ = _1060_ & _1059_ /*4376*/;
  assign _1062_ = inv_10[13] & r_9[19] /*4375*/;
  assign _1063_ = _1061_ | _1062_ /*4374*/;
  assign _1064_ = inv_10[14] ^ r_9[20] /*4372*/;
  assign sum_10[14] = _1064_ ^ _1063_ /*4371*/;
  assign _1065_ = _1064_ & _1063_ /*4370*/;
  assign _1066_ = inv_10[14] & r_9[20] /*4369*/;
  assign _1067_ = _1065_ | _1066_ /*4368*/;
  assign _1068_ = inv_10[15] ^ r_9[21] /*4366*/;
  assign sum_10[15] = _1068_ ^ _1067_ /*4365*/;
  assign _1069_ = _1068_ & _1067_ /*4364*/;
  assign _1070_ = inv_10[15] & r_9[21] /*4363*/;
  assign _1071_ = _1069_ | _1070_ /*4362*/;
  assign q[6] = ~sum_10[15] /*4373*/;
  assign m_10[0] = r_9[6] /*4372*/;
  assign m_10[1] = r_9[7] /*4371*/;
  assign m_10[2] = r_9[8] /*4370*/;
  assign m_10[3] = r_9[9] /*4369*/;
  assign m_10[4] = r_9[10] /*4368*/;
  assign m_10[5] = r_9[11] /*4367*/;
  assign m_10[6] = r_9[12] /*4366*/;
  assign m_10[7] = r_9[13] /*4365*/;
  assign m_10[8] = r_9[14] /*4364*/;
  assign m_10[9] = r_9[15] /*4363*/;
  assign m_10[10] = r_9[16] /*4362*/;
  assign m_10[11] = r_9[17] /*4361*/;
  assign m_10[12] = r_9[18] /*4360*/;
  assign m_10[13] = r_9[19] /*4359*/;
  assign m_10[14] = r_9[20] /*4358*/;
  assign m_10[15] = r_9[21] /*4357*/;
  assign _1072_ = ~q[6] /*4355*/;
  assign _1073_ = sum_10[0] & q[6] /*4354*/;
  assign _1074_ = m_10[0] & _1072_ /*4353*/;
  assign r_10[6] = _1074_ | _1073_ /*4352*/;
  assign _1075_ = ~q[6] /*4351*/;
  assign _1076_ = sum_10[1] & q[6] /*4350*/;
  assign _1077_ = m_10[1] & _1075_ /*4349*/;
  assign r_10[7] = _1077_ | _1076_ /*4348*/;
  assign _1078_ = ~q[6] /*4347*/;
  assign _1079_ = sum_10[2] & q[6] /*4346*/;
  assign _1080_ = m_10[2] & _1078_ /*4345*/;
  assign r_10[8] = _1080_ | _1079_ /*4344*/;
  assign _1081_ = ~q[6] /*4343*/;
  assign _1082_ = sum_10[3] & q[6] /*4342*/;
  assign _1083_ = m_10[3] & _1081_ /*4341*/;
  assign r_10[9] = _1083_ | _1082_ /*4340*/;
  assign _1084_ = ~q[6] /*4339*/;
  assign _1085_ = sum_10[4] & q[6] /*4338*/;
  assign _1086_ = m_10[4] & _1084_ /*4337*/;
  assign r_10[10] = _1086_ | _1085_ /*4336*/;
  assign _1087_ = ~q[6] /*4335*/;
  assign _1088_ = sum_10[5] & q[6] /*4334*/;
  assign _1089_ = m_10[5] & _1087_ /*4333*/;
  assign r_10[11] = _1089_ | _1088_ /*4332*/;
  assign _1090_ = ~q[6] /*4331*/;
  assign _1091_ = sum_10[6] & q[6] /*4330*/;
  assign _1092_ = m_10[6] & _1090_ /*4329*/;
  assign r_10[12] = _1092_ | _1091_ /*4328*/;
  assign _1093_ = ~q[6] /*4327*/;
  assign _1094_ = sum_10[7] & q[6] /*4326*/;
  assign _1095_ = m_10[7] & _1093_ /*4325*/;
  assign r_10[13] = _1095_ | _1094_ /*4324*/;
  assign _1096_ = ~q[6] /*4323*/;
  assign _1097_ = sum_10[8] & q[6] /*4322*/;
  assign _1098_ = m_10[8] & _1096_ /*4321*/;
  assign r_10[14] = _1098_ | _1097_ /*4320*/;
  assign _1099_ = ~q[6] /*4319*/;
  assign _1100_ = sum_10[9] & q[6] /*4318*/;
  assign _1101_ = m_10[9] & _1099_ /*4317*/;
  assign r_10[15] = _1101_ | _1100_ /*4316*/;
  assign _1102_ = ~q[6] /*4315*/;
  assign _1103_ = sum_10[10] & q[6] /*4314*/;
  assign _1104_ = m_10[10] & _1102_ /*4313*/;
  assign r_10[16] = _1104_ | _1103_ /*4312*/;
  assign _1105_ = ~q[6] /*4311*/;
  assign _1106_ = sum_10[11] & q[6] /*4310*/;
  assign _1107_ = m_10[11] & _1105_ /*4309*/;
  assign r_10[17] = _1107_ | _1106_ /*4308*/;
  assign _1108_ = ~q[6] /*4307*/;
  assign _1109_ = sum_10[12] & q[6] /*4306*/;
  assign _1110_ = m_10[12] & _1108_ /*4305*/;
  assign r_10[18] = _1110_ | _1109_ /*4304*/;
  assign _1111_ = ~q[6] /*4303*/;
  assign _1112_ = sum_10[13] & q[6] /*4302*/;
  assign _1113_ = m_10[13] & _1111_ /*4301*/;
  assign r_10[19] = _1113_ | _1112_ /*4300*/;
  assign _1114_ = ~q[6] /*4299*/;
  assign _1115_ = sum_10[14] & q[6] /*4298*/;
  assign _1116_ = m_10[14] & _1114_ /*4297*/;
  assign r_10[20] = _1116_ | _1115_ /*4296*/;
  assign _1117_ = ~q[6] /*4295*/;
  assign _1118_ = sum_10[15] & q[6] /*4294*/;
  assign _1119_ = m_10[15] & _1117_ /*4293*/;
  assign r_10[21] = _1119_ | _1118_ /*4292*/;
assign r_10[0]= r_9[0] /*4291*/;
assign r_10[1]= r_9[1] /*4290*/;
assign r_10[2]= r_9[2] /*4289*/;
assign r_10[3]= r_9[3] /*4288*/;
assign r_10[4]= r_9[4] /*4287*/;
assign r_10[5]= r_9[5] /*4286*/;
  assign inv_11[0] = ~div[0] /*4248*/;
  assign inv_11[1] = ~div[1] /*4247*/;
  assign inv_11[2] = ~div[2] /*4246*/;
  assign inv_11[3] = ~div[3] /*4245*/;
  assign inv_11[4] = ~div[4] /*4244*/;
  assign inv_11[5] = ~div[5] /*4243*/;
  assign inv_11[6] = ~div[6] /*4242*/;
  assign inv_11[7] = ~div[7] /*4241*/;
  assign inv_11[8] = ~div[8] /*4240*/;
  assign inv_11[9] = ~div[9] /*4239*/;
  assign inv_11[10] = ~div[10] /*4238*/;
  assign inv_11[11] = ~div[11] /*4237*/;
  assign inv_11[12] = ~div[12] /*4236*/;
  assign inv_11[13] = ~div[13] /*4235*/;
  assign inv_11[14] = ~div[14] /*4234*/;
assign inv_11[15] = oneWire /*4233*/;
  assign _1120_ = inv_11[0] ^ r_10[5] /*4231*/;
  assign sum_11[0] = _1120_ ^ oneWire /*4230*/;
  assign _1121_ = _1120_ & oneWire /*4229*/;
  assign _1122_ = inv_11[0] & r_10[5] /*4228*/;
  assign _1123_ = _1121_ | _1122_ /*4227*/;
  assign _1124_ = inv_11[1] ^ r_10[6] /*4226*/;
  assign sum_11[1] = _1124_ ^ _1123_ /*4225*/;
  assign _1125_ = _1124_ & _1123_ /*4224*/;
  assign _1126_ = inv_11[1] & r_10[6] /*4223*/;
  assign _1127_ = _1125_ | _1126_ /*4222*/;
  assign _1128_ = inv_11[2] ^ r_10[7] /*4220*/;
  assign sum_11[2] = _1128_ ^ _1127_ /*4219*/;
  assign _1129_ = _1128_ & _1127_ /*4218*/;
  assign _1130_ = inv_11[2] & r_10[7] /*4217*/;
  assign _1131_ = _1129_ | _1130_ /*4216*/;
  assign _1132_ = inv_11[3] ^ r_10[8] /*4214*/;
  assign sum_11[3] = _1132_ ^ _1131_ /*4213*/;
  assign _1133_ = _1132_ & _1131_ /*4212*/;
  assign _1134_ = inv_11[3] & r_10[8] /*4211*/;
  assign _1135_ = _1133_ | _1134_ /*4210*/;
  assign _1136_ = inv_11[4] ^ r_10[9] /*4208*/;
  assign sum_11[4] = _1136_ ^ _1135_ /*4207*/;
  assign _1137_ = _1136_ & _1135_ /*4206*/;
  assign _1138_ = inv_11[4] & r_10[9] /*4205*/;
  assign _1139_ = _1137_ | _1138_ /*4204*/;
  assign _1140_ = inv_11[5] ^ r_10[10] /*4202*/;
  assign sum_11[5] = _1140_ ^ _1139_ /*4201*/;
  assign _1141_ = _1140_ & _1139_ /*4200*/;
  assign _1142_ = inv_11[5] & r_10[10] /*4199*/;
  assign _1143_ = _1141_ | _1142_ /*4198*/;
  assign _1144_ = inv_11[6] ^ r_10[11] /*4196*/;
  assign sum_11[6] = _1144_ ^ _1143_ /*4195*/;
  assign _1145_ = _1144_ & _1143_ /*4194*/;
  assign _1146_ = inv_11[6] & r_10[11] /*4193*/;
  assign _1147_ = _1145_ | _1146_ /*4192*/;
  assign _1148_ = inv_11[7] ^ r_10[12] /*4190*/;
  assign sum_11[7] = _1148_ ^ _1147_ /*4189*/;
  assign _1149_ = _1148_ & _1147_ /*4188*/;
  assign _1150_ = inv_11[7] & r_10[12] /*4187*/;
  assign _1151_ = _1149_ | _1150_ /*4186*/;
  assign _1152_ = inv_11[8] ^ r_10[13] /*4184*/;
  assign sum_11[8] = _1152_ ^ _1151_ /*4183*/;
  assign _1153_ = _1152_ & _1151_ /*4182*/;
  assign _1154_ = inv_11[8] & r_10[13] /*4181*/;
  assign _1155_ = _1153_ | _1154_ /*4180*/;
  assign _1156_ = inv_11[9] ^ r_10[14] /*4178*/;
  assign sum_11[9] = _1156_ ^ _1155_ /*4177*/;
  assign _1157_ = _1156_ & _1155_ /*4176*/;
  assign _1158_ = inv_11[9] & r_10[14] /*4175*/;
  assign _1159_ = _1157_ | _1158_ /*4174*/;
  assign _1160_ = inv_11[10] ^ r_10[15] /*4172*/;
  assign sum_11[10] = _1160_ ^ _1159_ /*4171*/;
  assign _1161_ = _1160_ & _1159_ /*4170*/;
  assign _1162_ = inv_11[10] & r_10[15] /*4169*/;
  assign _1163_ = _1161_ | _1162_ /*4168*/;
  assign _1164_ = inv_11[11] ^ r_10[16] /*4166*/;
  assign sum_11[11] = _1164_ ^ _1163_ /*4165*/;
  assign _1165_ = _1164_ & _1163_ /*4164*/;
  assign _1166_ = inv_11[11] & r_10[16] /*4163*/;
  assign _1167_ = _1165_ | _1166_ /*4162*/;
  assign _1168_ = inv_11[12] ^ r_10[17] /*4160*/;
  assign sum_11[12] = _1168_ ^ _1167_ /*4159*/;
  assign _1169_ = _1168_ & _1167_ /*4158*/;
  assign _1170_ = inv_11[12] & r_10[17] /*4157*/;
  assign _1171_ = _1169_ | _1170_ /*4156*/;
  assign _1172_ = inv_11[13] ^ r_10[18] /*4154*/;
  assign sum_11[13] = _1172_ ^ _1171_ /*4153*/;
  assign _1173_ = _1172_ & _1171_ /*4152*/;
  assign _1174_ = inv_11[13] & r_10[18] /*4151*/;
  assign _1175_ = _1173_ | _1174_ /*4150*/;
  assign _1176_ = inv_11[14] ^ r_10[19] /*4148*/;
  assign sum_11[14] = _1176_ ^ _1175_ /*4147*/;
  assign _1177_ = _1176_ & _1175_ /*4146*/;
  assign _1178_ = inv_11[14] & r_10[19] /*4145*/;
  assign _1179_ = _1177_ | _1178_ /*4144*/;
  assign _1180_ = inv_11[15] ^ r_10[20] /*4142*/;
  assign sum_11[15] = _1180_ ^ _1179_ /*4141*/;
  assign _1181_ = _1180_ & _1179_ /*4140*/;
  assign _1182_ = inv_11[15] & r_10[20] /*4139*/;
  assign _1183_ = _1181_ | _1182_ /*4138*/;
  assign q[5] = ~sum_11[15] /*4149*/;
  assign m_11[0] = r_10[5] /*4148*/;
  assign m_11[1] = r_10[6] /*4147*/;
  assign m_11[2] = r_10[7] /*4146*/;
  assign m_11[3] = r_10[8] /*4145*/;
  assign m_11[4] = r_10[9] /*4144*/;
  assign m_11[5] = r_10[10] /*4143*/;
  assign m_11[6] = r_10[11] /*4142*/;
  assign m_11[7] = r_10[12] /*4141*/;
  assign m_11[8] = r_10[13] /*4140*/;
  assign m_11[9] = r_10[14] /*4139*/;
  assign m_11[10] = r_10[15] /*4138*/;
  assign m_11[11] = r_10[16] /*4137*/;
  assign m_11[12] = r_10[17] /*4136*/;
  assign m_11[13] = r_10[18] /*4135*/;
  assign m_11[14] = r_10[19] /*4134*/;
  assign m_11[15] = r_10[20] /*4133*/;
  assign _1184_ = ~q[5] /*4131*/;
  assign _1185_ = sum_11[0] & q[5] /*4130*/;
  assign _1186_ = m_11[0] & _1184_ /*4129*/;
  assign r_11[5] = _1186_ | _1185_ /*4128*/;
  assign _1187_ = ~q[5] /*4127*/;
  assign _1188_ = sum_11[1] & q[5] /*4126*/;
  assign _1189_ = m_11[1] & _1187_ /*4125*/;
  assign r_11[6] = _1189_ | _1188_ /*4124*/;
  assign _1190_ = ~q[5] /*4123*/;
  assign _1191_ = sum_11[2] & q[5] /*4122*/;
  assign _1192_ = m_11[2] & _1190_ /*4121*/;
  assign r_11[7] = _1192_ | _1191_ /*4120*/;
  assign _1193_ = ~q[5] /*4119*/;
  assign _1194_ = sum_11[3] & q[5] /*4118*/;
  assign _1195_ = m_11[3] & _1193_ /*4117*/;
  assign r_11[8] = _1195_ | _1194_ /*4116*/;
  assign _1196_ = ~q[5] /*4115*/;
  assign _1197_ = sum_11[4] & q[5] /*4114*/;
  assign _1198_ = m_11[4] & _1196_ /*4113*/;
  assign r_11[9] = _1198_ | _1197_ /*4112*/;
  assign _1199_ = ~q[5] /*4111*/;
  assign _1200_ = sum_11[5] & q[5] /*4110*/;
  assign _1201_ = m_11[5] & _1199_ /*4109*/;
  assign r_11[10] = _1201_ | _1200_ /*4108*/;
  assign _1202_ = ~q[5] /*4107*/;
  assign _1203_ = sum_11[6] & q[5] /*4106*/;
  assign _1204_ = m_11[6] & _1202_ /*4105*/;
  assign r_11[11] = _1204_ | _1203_ /*4104*/;
  assign _1205_ = ~q[5] /*4103*/;
  assign _1206_ = sum_11[7] & q[5] /*4102*/;
  assign _1207_ = m_11[7] & _1205_ /*4101*/;
  assign r_11[12] = _1207_ | _1206_ /*4100*/;
  assign _1208_ = ~q[5] /*4099*/;
  assign _1209_ = sum_11[8] & q[5] /*4098*/;
  assign _1210_ = m_11[8] & _1208_ /*4097*/;
  assign r_11[13] = _1210_ | _1209_ /*4096*/;
  assign _1211_ = ~q[5] /*4095*/;
  assign _1212_ = sum_11[9] & q[5] /*4094*/;
  assign _1213_ = m_11[9] & _1211_ /*4093*/;
  assign r_11[14] = _1213_ | _1212_ /*4092*/;
  assign _1214_ = ~q[5] /*4091*/;
  assign _1215_ = sum_11[10] & q[5] /*4090*/;
  assign _1216_ = m_11[10] & _1214_ /*4089*/;
  assign r_11[15] = _1216_ | _1215_ /*4088*/;
  assign _1217_ = ~q[5] /*4087*/;
  assign _1218_ = sum_11[11] & q[5] /*4086*/;
  assign _1219_ = m_11[11] & _1217_ /*4085*/;
  assign r_11[16] = _1219_ | _1218_ /*4084*/;
  assign _1220_ = ~q[5] /*4083*/;
  assign _1221_ = sum_11[12] & q[5] /*4082*/;
  assign _1222_ = m_11[12] & _1220_ /*4081*/;
  assign r_11[17] = _1222_ | _1221_ /*4080*/;
  assign _1223_ = ~q[5] /*4079*/;
  assign _1224_ = sum_11[13] & q[5] /*4078*/;
  assign _1225_ = m_11[13] & _1223_ /*4077*/;
  assign r_11[18] = _1225_ | _1224_ /*4076*/;
  assign _1226_ = ~q[5] /*4075*/;
  assign _1227_ = sum_11[14] & q[5] /*4074*/;
  assign _1228_ = m_11[14] & _1226_ /*4073*/;
  assign r_11[19] = _1228_ | _1227_ /*4072*/;
  assign _1229_ = ~q[5] /*4071*/;
  assign _1230_ = sum_11[15] & q[5] /*4070*/;
  assign _1231_ = m_11[15] & _1229_ /*4069*/;
  assign r_11[20] = _1231_ | _1230_ /*4068*/;
assign r_11[0]= r_10[0] /*4067*/;
assign r_11[1]= r_10[1] /*4066*/;
assign r_11[2]= r_10[2] /*4065*/;
assign r_11[3]= r_10[3] /*4064*/;
assign r_11[4]= r_10[4] /*4063*/;
  assign inv_12[0] = ~div[0] /*4024*/;
  assign inv_12[1] = ~div[1] /*4023*/;
  assign inv_12[2] = ~div[2] /*4022*/;
  assign inv_12[3] = ~div[3] /*4021*/;
  assign inv_12[4] = ~div[4] /*4020*/;
  assign inv_12[5] = ~div[5] /*4019*/;
  assign inv_12[6] = ~div[6] /*4018*/;
  assign inv_12[7] = ~div[7] /*4017*/;
  assign inv_12[8] = ~div[8] /*4016*/;
  assign inv_12[9] = ~div[9] /*4015*/;
  assign inv_12[10] = ~div[10] /*4014*/;
  assign inv_12[11] = ~div[11] /*4013*/;
  assign inv_12[12] = ~div[12] /*4012*/;
  assign inv_12[13] = ~div[13] /*4011*/;
  assign inv_12[14] = ~div[14] /*4010*/;
assign inv_12[15] = oneWire /*4009*/;
  assign _1232_ = inv_12[0] ^ r_11[4] /*4007*/;
  assign sum_12[0] = _1232_ ^ oneWire /*4006*/;
  assign _1233_ = _1232_ & oneWire /*4005*/;
  assign _1234_ = inv_12[0] & r_11[4] /*4004*/;
  assign _1235_ = _1233_ | _1234_ /*4003*/;
  assign _1236_ = inv_12[1] ^ r_11[5] /*4002*/;
  assign sum_12[1] = _1236_ ^ _1235_ /*4001*/;
  assign _1237_ = _1236_ & _1235_ /*4000*/;
  assign _1238_ = inv_12[1] & r_11[5] /*3999*/;
  assign _1239_ = _1237_ | _1238_ /*3998*/;
  assign _1240_ = inv_12[2] ^ r_11[6] /*3996*/;
  assign sum_12[2] = _1240_ ^ _1239_ /*3995*/;
  assign _1241_ = _1240_ & _1239_ /*3994*/;
  assign _1242_ = inv_12[2] & r_11[6] /*3993*/;
  assign _1243_ = _1241_ | _1242_ /*3992*/;
  assign _1244_ = inv_12[3] ^ r_11[7] /*3990*/;
  assign sum_12[3] = _1244_ ^ _1243_ /*3989*/;
  assign _1245_ = _1244_ & _1243_ /*3988*/;
  assign _1246_ = inv_12[3] & r_11[7] /*3987*/;
  assign _1247_ = _1245_ | _1246_ /*3986*/;
  assign _1248_ = inv_12[4] ^ r_11[8] /*3984*/;
  assign sum_12[4] = _1248_ ^ _1247_ /*3983*/;
  assign _1249_ = _1248_ & _1247_ /*3982*/;
  assign _1250_ = inv_12[4] & r_11[8] /*3981*/;
  assign _1251_ = _1249_ | _1250_ /*3980*/;
  assign _1252_ = inv_12[5] ^ r_11[9] /*3978*/;
  assign sum_12[5] = _1252_ ^ _1251_ /*3977*/;
  assign _1253_ = _1252_ & _1251_ /*3976*/;
  assign _1254_ = inv_12[5] & r_11[9] /*3975*/;
  assign _1255_ = _1253_ | _1254_ /*3974*/;
  assign _1256_ = inv_12[6] ^ r_11[10] /*3972*/;
  assign sum_12[6] = _1256_ ^ _1255_ /*3971*/;
  assign _1257_ = _1256_ & _1255_ /*3970*/;
  assign _1258_ = inv_12[6] & r_11[10] /*3969*/;
  assign _1259_ = _1257_ | _1258_ /*3968*/;
  assign _1260_ = inv_12[7] ^ r_11[11] /*3966*/;
  assign sum_12[7] = _1260_ ^ _1259_ /*3965*/;
  assign _1261_ = _1260_ & _1259_ /*3964*/;
  assign _1262_ = inv_12[7] & r_11[11] /*3963*/;
  assign _1263_ = _1261_ | _1262_ /*3962*/;
  assign _1264_ = inv_12[8] ^ r_11[12] /*3960*/;
  assign sum_12[8] = _1264_ ^ _1263_ /*3959*/;
  assign _1265_ = _1264_ & _1263_ /*3958*/;
  assign _1266_ = inv_12[8] & r_11[12] /*3957*/;
  assign _1267_ = _1265_ | _1266_ /*3956*/;
  assign _1268_ = inv_12[9] ^ r_11[13] /*3954*/;
  assign sum_12[9] = _1268_ ^ _1267_ /*3953*/;
  assign _1269_ = _1268_ & _1267_ /*3952*/;
  assign _1270_ = inv_12[9] & r_11[13] /*3951*/;
  assign _1271_ = _1269_ | _1270_ /*3950*/;
  assign _1272_ = inv_12[10] ^ r_11[14] /*3948*/;
  assign sum_12[10] = _1272_ ^ _1271_ /*3947*/;
  assign _1273_ = _1272_ & _1271_ /*3946*/;
  assign _1274_ = inv_12[10] & r_11[14] /*3945*/;
  assign _1275_ = _1273_ | _1274_ /*3944*/;
  assign _1276_ = inv_12[11] ^ r_11[15] /*3942*/;
  assign sum_12[11] = _1276_ ^ _1275_ /*3941*/;
  assign _1277_ = _1276_ & _1275_ /*3940*/;
  assign _1278_ = inv_12[11] & r_11[15] /*3939*/;
  assign _1279_ = _1277_ | _1278_ /*3938*/;
  assign _1280_ = inv_12[12] ^ r_11[16] /*3936*/;
  assign sum_12[12] = _1280_ ^ _1279_ /*3935*/;
  assign _1281_ = _1280_ & _1279_ /*3934*/;
  assign _1282_ = inv_12[12] & r_11[16] /*3933*/;
  assign _1283_ = _1281_ | _1282_ /*3932*/;
  assign _1284_ = inv_12[13] ^ r_11[17] /*3930*/;
  assign sum_12[13] = _1284_ ^ _1283_ /*3929*/;
  assign _1285_ = _1284_ & _1283_ /*3928*/;
  assign _1286_ = inv_12[13] & r_11[17] /*3927*/;
  assign _1287_ = _1285_ | _1286_ /*3926*/;
  assign _1288_ = inv_12[14] ^ r_11[18] /*3924*/;
  assign sum_12[14] = _1288_ ^ _1287_ /*3923*/;
  assign _1289_ = _1288_ & _1287_ /*3922*/;
  assign _1290_ = inv_12[14] & r_11[18] /*3921*/;
  assign _1291_ = _1289_ | _1290_ /*3920*/;
  assign _1292_ = inv_12[15] ^ r_11[19] /*3918*/;
  assign sum_12[15] = _1292_ ^ _1291_ /*3917*/;
  assign _1293_ = _1292_ & _1291_ /*3916*/;
  assign _1294_ = inv_12[15] & r_11[19] /*3915*/;
  assign _1295_ = _1293_ | _1294_ /*3914*/;
  assign q[4] = ~sum_12[15] /*3925*/;
  assign m_12[0] = r_11[4] /*3924*/;
  assign m_12[1] = r_11[5] /*3923*/;
  assign m_12[2] = r_11[6] /*3922*/;
  assign m_12[3] = r_11[7] /*3921*/;
  assign m_12[4] = r_11[8] /*3920*/;
  assign m_12[5] = r_11[9] /*3919*/;
  assign m_12[6] = r_11[10] /*3918*/;
  assign m_12[7] = r_11[11] /*3917*/;
  assign m_12[8] = r_11[12] /*3916*/;
  assign m_12[9] = r_11[13] /*3915*/;
  assign m_12[10] = r_11[14] /*3914*/;
  assign m_12[11] = r_11[15] /*3913*/;
  assign m_12[12] = r_11[16] /*3912*/;
  assign m_12[13] = r_11[17] /*3911*/;
  assign m_12[14] = r_11[18] /*3910*/;
  assign m_12[15] = r_11[19] /*3909*/;
  assign _1296_ = ~q[4] /*3907*/;
  assign _1297_ = sum_12[0] & q[4] /*3906*/;
  assign _1298_ = m_12[0] & _1296_ /*3905*/;
  assign r_12[4] = _1298_ | _1297_ /*3904*/;
  assign _1299_ = ~q[4] /*3903*/;
  assign _1300_ = sum_12[1] & q[4] /*3902*/;
  assign _1301_ = m_12[1] & _1299_ /*3901*/;
  assign r_12[5] = _1301_ | _1300_ /*3900*/;
  assign _1302_ = ~q[4] /*3899*/;
  assign _1303_ = sum_12[2] & q[4] /*3898*/;
  assign _1304_ = m_12[2] & _1302_ /*3897*/;
  assign r_12[6] = _1304_ | _1303_ /*3896*/;
  assign _1305_ = ~q[4] /*3895*/;
  assign _1306_ = sum_12[3] & q[4] /*3894*/;
  assign _1307_ = m_12[3] & _1305_ /*3893*/;
  assign r_12[7] = _1307_ | _1306_ /*3892*/;
  assign _1308_ = ~q[4] /*3891*/;
  assign _1309_ = sum_12[4] & q[4] /*3890*/;
  assign _1310_ = m_12[4] & _1308_ /*3889*/;
  assign r_12[8] = _1310_ | _1309_ /*3888*/;
  assign _1311_ = ~q[4] /*3887*/;
  assign _1312_ = sum_12[5] & q[4] /*3886*/;
  assign _1313_ = m_12[5] & _1311_ /*3885*/;
  assign r_12[9] = _1313_ | _1312_ /*3884*/;
  assign _1314_ = ~q[4] /*3883*/;
  assign _1315_ = sum_12[6] & q[4] /*3882*/;
  assign _1316_ = m_12[6] & _1314_ /*3881*/;
  assign r_12[10] = _1316_ | _1315_ /*3880*/;
  assign _1317_ = ~q[4] /*3879*/;
  assign _1318_ = sum_12[7] & q[4] /*3878*/;
  assign _1319_ = m_12[7] & _1317_ /*3877*/;
  assign r_12[11] = _1319_ | _1318_ /*3876*/;
  assign _1320_ = ~q[4] /*3875*/;
  assign _1321_ = sum_12[8] & q[4] /*3874*/;
  assign _1322_ = m_12[8] & _1320_ /*3873*/;
  assign r_12[12] = _1322_ | _1321_ /*3872*/;
  assign _1323_ = ~q[4] /*3871*/;
  assign _1324_ = sum_12[9] & q[4] /*3870*/;
  assign _1325_ = m_12[9] & _1323_ /*3869*/;
  assign r_12[13] = _1325_ | _1324_ /*3868*/;
  assign _1326_ = ~q[4] /*3867*/;
  assign _1327_ = sum_12[10] & q[4] /*3866*/;
  assign _1328_ = m_12[10] & _1326_ /*3865*/;
  assign r_12[14] = _1328_ | _1327_ /*3864*/;
  assign _1329_ = ~q[4] /*3863*/;
  assign _1330_ = sum_12[11] & q[4] /*3862*/;
  assign _1331_ = m_12[11] & _1329_ /*3861*/;
  assign r_12[15] = _1331_ | _1330_ /*3860*/;
  assign _1332_ = ~q[4] /*3859*/;
  assign _1333_ = sum_12[12] & q[4] /*3858*/;
  assign _1334_ = m_12[12] & _1332_ /*3857*/;
  assign r_12[16] = _1334_ | _1333_ /*3856*/;
  assign _1335_ = ~q[4] /*3855*/;
  assign _1336_ = sum_12[13] & q[4] /*3854*/;
  assign _1337_ = m_12[13] & _1335_ /*3853*/;
  assign r_12[17] = _1337_ | _1336_ /*3852*/;
  assign _1338_ = ~q[4] /*3851*/;
  assign _1339_ = sum_12[14] & q[4] /*3850*/;
  assign _1340_ = m_12[14] & _1338_ /*3849*/;
  assign r_12[18] = _1340_ | _1339_ /*3848*/;
  assign _1341_ = ~q[4] /*3847*/;
  assign _1342_ = sum_12[15] & q[4] /*3846*/;
  assign _1343_ = m_12[15] & _1341_ /*3845*/;
  assign r_12[19] = _1343_ | _1342_ /*3844*/;
assign r_12[0]= r_11[0] /*3843*/;
assign r_12[1]= r_11[1] /*3842*/;
assign r_12[2]= r_11[2] /*3841*/;
assign r_12[3]= r_11[3] /*3840*/;
  assign inv_13[0] = ~div[0] /*3800*/;
  assign inv_13[1] = ~div[1] /*3799*/;
  assign inv_13[2] = ~div[2] /*3798*/;
  assign inv_13[3] = ~div[3] /*3797*/;
  assign inv_13[4] = ~div[4] /*3796*/;
  assign inv_13[5] = ~div[5] /*3795*/;
  assign inv_13[6] = ~div[6] /*3794*/;
  assign inv_13[7] = ~div[7] /*3793*/;
  assign inv_13[8] = ~div[8] /*3792*/;
  assign inv_13[9] = ~div[9] /*3791*/;
  assign inv_13[10] = ~div[10] /*3790*/;
  assign inv_13[11] = ~div[11] /*3789*/;
  assign inv_13[12] = ~div[12] /*3788*/;
  assign inv_13[13] = ~div[13] /*3787*/;
  assign inv_13[14] = ~div[14] /*3786*/;
assign inv_13[15] = oneWire /*3785*/;
  assign _1344_ = inv_13[0] ^ r_12[3] /*3783*/;
  assign sum_13[0] = _1344_ ^ oneWire /*3782*/;
  assign _1345_ = _1344_ & oneWire /*3781*/;
  assign _1346_ = inv_13[0] & r_12[3] /*3780*/;
  assign _1347_ = _1345_ | _1346_ /*3779*/;
  assign _1348_ = inv_13[1] ^ r_12[4] /*3778*/;
  assign sum_13[1] = _1348_ ^ _1347_ /*3777*/;
  assign _1349_ = _1348_ & _1347_ /*3776*/;
  assign _1350_ = inv_13[1] & r_12[4] /*3775*/;
  assign _1351_ = _1349_ | _1350_ /*3774*/;
  assign _1352_ = inv_13[2] ^ r_12[5] /*3772*/;
  assign sum_13[2] = _1352_ ^ _1351_ /*3771*/;
  assign _1353_ = _1352_ & _1351_ /*3770*/;
  assign _1354_ = inv_13[2] & r_12[5] /*3769*/;
  assign _1355_ = _1353_ | _1354_ /*3768*/;
  assign _1356_ = inv_13[3] ^ r_12[6] /*3766*/;
  assign sum_13[3] = _1356_ ^ _1355_ /*3765*/;
  assign _1357_ = _1356_ & _1355_ /*3764*/;
  assign _1358_ = inv_13[3] & r_12[6] /*3763*/;
  assign _1359_ = _1357_ | _1358_ /*3762*/;
  assign _1360_ = inv_13[4] ^ r_12[7] /*3760*/;
  assign sum_13[4] = _1360_ ^ _1359_ /*3759*/;
  assign _1361_ = _1360_ & _1359_ /*3758*/;
  assign _1362_ = inv_13[4] & r_12[7] /*3757*/;
  assign _1363_ = _1361_ | _1362_ /*3756*/;
  assign _1364_ = inv_13[5] ^ r_12[8] /*3754*/;
  assign sum_13[5] = _1364_ ^ _1363_ /*3753*/;
  assign _1365_ = _1364_ & _1363_ /*3752*/;
  assign _1366_ = inv_13[5] & r_12[8] /*3751*/;
  assign _1367_ = _1365_ | _1366_ /*3750*/;
  assign _1368_ = inv_13[6] ^ r_12[9] /*3748*/;
  assign sum_13[6] = _1368_ ^ _1367_ /*3747*/;
  assign _1369_ = _1368_ & _1367_ /*3746*/;
  assign _1370_ = inv_13[6] & r_12[9] /*3745*/;
  assign _1371_ = _1369_ | _1370_ /*3744*/;
  assign _1372_ = inv_13[7] ^ r_12[10] /*3742*/;
  assign sum_13[7] = _1372_ ^ _1371_ /*3741*/;
  assign _1373_ = _1372_ & _1371_ /*3740*/;
  assign _1374_ = inv_13[7] & r_12[10] /*3739*/;
  assign _1375_ = _1373_ | _1374_ /*3738*/;
  assign _1376_ = inv_13[8] ^ r_12[11] /*3736*/;
  assign sum_13[8] = _1376_ ^ _1375_ /*3735*/;
  assign _1377_ = _1376_ & _1375_ /*3734*/;
  assign _1378_ = inv_13[8] & r_12[11] /*3733*/;
  assign _1379_ = _1377_ | _1378_ /*3732*/;
  assign _1380_ = inv_13[9] ^ r_12[12] /*3730*/;
  assign sum_13[9] = _1380_ ^ _1379_ /*3729*/;
  assign _1381_ = _1380_ & _1379_ /*3728*/;
  assign _1382_ = inv_13[9] & r_12[12] /*3727*/;
  assign _1383_ = _1381_ | _1382_ /*3726*/;
  assign _1384_ = inv_13[10] ^ r_12[13] /*3724*/;
  assign sum_13[10] = _1384_ ^ _1383_ /*3723*/;
  assign _1385_ = _1384_ & _1383_ /*3722*/;
  assign _1386_ = inv_13[10] & r_12[13] /*3721*/;
  assign _1387_ = _1385_ | _1386_ /*3720*/;
  assign _1388_ = inv_13[11] ^ r_12[14] /*3718*/;
  assign sum_13[11] = _1388_ ^ _1387_ /*3717*/;
  assign _1389_ = _1388_ & _1387_ /*3716*/;
  assign _1390_ = inv_13[11] & r_12[14] /*3715*/;
  assign _1391_ = _1389_ | _1390_ /*3714*/;
  assign _1392_ = inv_13[12] ^ r_12[15] /*3712*/;
  assign sum_13[12] = _1392_ ^ _1391_ /*3711*/;
  assign _1393_ = _1392_ & _1391_ /*3710*/;
  assign _1394_ = inv_13[12] & r_12[15] /*3709*/;
  assign _1395_ = _1393_ | _1394_ /*3708*/;
  assign _1396_ = inv_13[13] ^ r_12[16] /*3706*/;
  assign sum_13[13] = _1396_ ^ _1395_ /*3705*/;
  assign _1397_ = _1396_ & _1395_ /*3704*/;
  assign _1398_ = inv_13[13] & r_12[16] /*3703*/;
  assign _1399_ = _1397_ | _1398_ /*3702*/;
  assign _1400_ = inv_13[14] ^ r_12[17] /*3700*/;
  assign sum_13[14] = _1400_ ^ _1399_ /*3699*/;
  assign _1401_ = _1400_ & _1399_ /*3698*/;
  assign _1402_ = inv_13[14] & r_12[17] /*3697*/;
  assign _1403_ = _1401_ | _1402_ /*3696*/;
  assign _1404_ = inv_13[15] ^ r_12[18] /*3694*/;
  assign sum_13[15] = _1404_ ^ _1403_ /*3693*/;
  assign _1405_ = _1404_ & _1403_ /*3692*/;
  assign _1406_ = inv_13[15] & r_12[18] /*3691*/;
  assign _1407_ = _1405_ | _1406_ /*3690*/;
  assign q[3] = ~sum_13[15] /*3701*/;
  assign m_13[0] = r_12[3] /*3700*/;
  assign m_13[1] = r_12[4] /*3699*/;
  assign m_13[2] = r_12[5] /*3698*/;
  assign m_13[3] = r_12[6] /*3697*/;
  assign m_13[4] = r_12[7] /*3696*/;
  assign m_13[5] = r_12[8] /*3695*/;
  assign m_13[6] = r_12[9] /*3694*/;
  assign m_13[7] = r_12[10] /*3693*/;
  assign m_13[8] = r_12[11] /*3692*/;
  assign m_13[9] = r_12[12] /*3691*/;
  assign m_13[10] = r_12[13] /*3690*/;
  assign m_13[11] = r_12[14] /*3689*/;
  assign m_13[12] = r_12[15] /*3688*/;
  assign m_13[13] = r_12[16] /*3687*/;
  assign m_13[14] = r_12[17] /*3686*/;
  assign m_13[15] = r_12[18] /*3685*/;
  assign _1408_ = ~q[3] /*3683*/;
  assign _1409_ = sum_13[0] & q[3] /*3682*/;
  assign _1410_ = m_13[0] & _1408_ /*3681*/;
  assign r_13[3] = _1410_ | _1409_ /*3680*/;
  assign _1411_ = ~q[3] /*3679*/;
  assign _1412_ = sum_13[1] & q[3] /*3678*/;
  assign _1413_ = m_13[1] & _1411_ /*3677*/;
  assign r_13[4] = _1413_ | _1412_ /*3676*/;
  assign _1414_ = ~q[3] /*3675*/;
  assign _1415_ = sum_13[2] & q[3] /*3674*/;
  assign _1416_ = m_13[2] & _1414_ /*3673*/;
  assign r_13[5] = _1416_ | _1415_ /*3672*/;
  assign _1417_ = ~q[3] /*3671*/;
  assign _1418_ = sum_13[3] & q[3] /*3670*/;
  assign _1419_ = m_13[3] & _1417_ /*3669*/;
  assign r_13[6] = _1419_ | _1418_ /*3668*/;
  assign _1420_ = ~q[3] /*3667*/;
  assign _1421_ = sum_13[4] & q[3] /*3666*/;
  assign _1422_ = m_13[4] & _1420_ /*3665*/;
  assign r_13[7] = _1422_ | _1421_ /*3664*/;
  assign _1423_ = ~q[3] /*3663*/;
  assign _1424_ = sum_13[5] & q[3] /*3662*/;
  assign _1425_ = m_13[5] & _1423_ /*3661*/;
  assign r_13[8] = _1425_ | _1424_ /*3660*/;
  assign _1426_ = ~q[3] /*3659*/;
  assign _1427_ = sum_13[6] & q[3] /*3658*/;
  assign _1428_ = m_13[6] & _1426_ /*3657*/;
  assign r_13[9] = _1428_ | _1427_ /*3656*/;
  assign _1429_ = ~q[3] /*3655*/;
  assign _1430_ = sum_13[7] & q[3] /*3654*/;
  assign _1431_ = m_13[7] & _1429_ /*3653*/;
  assign r_13[10] = _1431_ | _1430_ /*3652*/;
  assign _1432_ = ~q[3] /*3651*/;
  assign _1433_ = sum_13[8] & q[3] /*3650*/;
  assign _1434_ = m_13[8] & _1432_ /*3649*/;
  assign r_13[11] = _1434_ | _1433_ /*3648*/;
  assign _1435_ = ~q[3] /*3647*/;
  assign _1436_ = sum_13[9] & q[3] /*3646*/;
  assign _1437_ = m_13[9] & _1435_ /*3645*/;
  assign r_13[12] = _1437_ | _1436_ /*3644*/;
  assign _1438_ = ~q[3] /*3643*/;
  assign _1439_ = sum_13[10] & q[3] /*3642*/;
  assign _1440_ = m_13[10] & _1438_ /*3641*/;
  assign r_13[13] = _1440_ | _1439_ /*3640*/;
  assign _1441_ = ~q[3] /*3639*/;
  assign _1442_ = sum_13[11] & q[3] /*3638*/;
  assign _1443_ = m_13[11] & _1441_ /*3637*/;
  assign r_13[14] = _1443_ | _1442_ /*3636*/;
  assign _1444_ = ~q[3] /*3635*/;
  assign _1445_ = sum_13[12] & q[3] /*3634*/;
  assign _1446_ = m_13[12] & _1444_ /*3633*/;
  assign r_13[15] = _1446_ | _1445_ /*3632*/;
  assign _1447_ = ~q[3] /*3631*/;
  assign _1448_ = sum_13[13] & q[3] /*3630*/;
  assign _1449_ = m_13[13] & _1447_ /*3629*/;
  assign r_13[16] = _1449_ | _1448_ /*3628*/;
  assign _1450_ = ~q[3] /*3627*/;
  assign _1451_ = sum_13[14] & q[3] /*3626*/;
  assign _1452_ = m_13[14] & _1450_ /*3625*/;
  assign r_13[17] = _1452_ | _1451_ /*3624*/;
  assign _1453_ = ~q[3] /*3623*/;
  assign _1454_ = sum_13[15] & q[3] /*3622*/;
  assign _1455_ = m_13[15] & _1453_ /*3621*/;
  assign r_13[18] = _1455_ | _1454_ /*3620*/;
assign r_13[0]= r_12[0] /*3619*/;
assign r_13[1]= r_12[1] /*3618*/;
assign r_13[2]= r_12[2] /*3617*/;
  assign inv_14[0] = ~div[0] /*3576*/;
  assign inv_14[1] = ~div[1] /*3575*/;
  assign inv_14[2] = ~div[2] /*3574*/;
  assign inv_14[3] = ~div[3] /*3573*/;
  assign inv_14[4] = ~div[4] /*3572*/;
  assign inv_14[5] = ~div[5] /*3571*/;
  assign inv_14[6] = ~div[6] /*3570*/;
  assign inv_14[7] = ~div[7] /*3569*/;
  assign inv_14[8] = ~div[8] /*3568*/;
  assign inv_14[9] = ~div[9] /*3567*/;
  assign inv_14[10] = ~div[10] /*3566*/;
  assign inv_14[11] = ~div[11] /*3565*/;
  assign inv_14[12] = ~div[12] /*3564*/;
  assign inv_14[13] = ~div[13] /*3563*/;
  assign inv_14[14] = ~div[14] /*3562*/;
assign inv_14[15] = oneWire /*3561*/;
  assign _1456_ = inv_14[0] ^ r_13[2] /*3559*/;
  assign sum_14[0] = _1456_ ^ oneWire /*3558*/;
  assign _1457_ = _1456_ & oneWire /*3557*/;
  assign _1458_ = inv_14[0] & r_13[2] /*3556*/;
  assign _1459_ = _1457_ | _1458_ /*3555*/;
  assign _1460_ = inv_14[1] ^ r_13[3] /*3554*/;
  assign sum_14[1] = _1460_ ^ _1459_ /*3553*/;
  assign _1461_ = _1460_ & _1459_ /*3552*/;
  assign _1462_ = inv_14[1] & r_13[3] /*3551*/;
  assign _1463_ = _1461_ | _1462_ /*3550*/;
  assign _1464_ = inv_14[2] ^ r_13[4] /*3548*/;
  assign sum_14[2] = _1464_ ^ _1463_ /*3547*/;
  assign _1465_ = _1464_ & _1463_ /*3546*/;
  assign _1466_ = inv_14[2] & r_13[4] /*3545*/;
  assign _1467_ = _1465_ | _1466_ /*3544*/;
  assign _1468_ = inv_14[3] ^ r_13[5] /*3542*/;
  assign sum_14[3] = _1468_ ^ _1467_ /*3541*/;
  assign _1469_ = _1468_ & _1467_ /*3540*/;
  assign _1470_ = inv_14[3] & r_13[5] /*3539*/;
  assign _1471_ = _1469_ | _1470_ /*3538*/;
  assign _1472_ = inv_14[4] ^ r_13[6] /*3536*/;
  assign sum_14[4] = _1472_ ^ _1471_ /*3535*/;
  assign _1473_ = _1472_ & _1471_ /*3534*/;
  assign _1474_ = inv_14[4] & r_13[6] /*3533*/;
  assign _1475_ = _1473_ | _1474_ /*3532*/;
  assign _1476_ = inv_14[5] ^ r_13[7] /*3530*/;
  assign sum_14[5] = _1476_ ^ _1475_ /*3529*/;
  assign _1477_ = _1476_ & _1475_ /*3528*/;
  assign _1478_ = inv_14[5] & r_13[7] /*3527*/;
  assign _1479_ = _1477_ | _1478_ /*3526*/;
  assign _1480_ = inv_14[6] ^ r_13[8] /*3524*/;
  assign sum_14[6] = _1480_ ^ _1479_ /*3523*/;
  assign _1481_ = _1480_ & _1479_ /*3522*/;
  assign _1482_ = inv_14[6] & r_13[8] /*3521*/;
  assign _1483_ = _1481_ | _1482_ /*3520*/;
  assign _1484_ = inv_14[7] ^ r_13[9] /*3518*/;
  assign sum_14[7] = _1484_ ^ _1483_ /*3517*/;
  assign _1485_ = _1484_ & _1483_ /*3516*/;
  assign _1486_ = inv_14[7] & r_13[9] /*3515*/;
  assign _1487_ = _1485_ | _1486_ /*3514*/;
  assign _1488_ = inv_14[8] ^ r_13[10] /*3512*/;
  assign sum_14[8] = _1488_ ^ _1487_ /*3511*/;
  assign _1489_ = _1488_ & _1487_ /*3510*/;
  assign _1490_ = inv_14[8] & r_13[10] /*3509*/;
  assign _1491_ = _1489_ | _1490_ /*3508*/;
  assign _1492_ = inv_14[9] ^ r_13[11] /*3506*/;
  assign sum_14[9] = _1492_ ^ _1491_ /*3505*/;
  assign _1493_ = _1492_ & _1491_ /*3504*/;
  assign _1494_ = inv_14[9] & r_13[11] /*3503*/;
  assign _1495_ = _1493_ | _1494_ /*3502*/;
  assign _1496_ = inv_14[10] ^ r_13[12] /*3500*/;
  assign sum_14[10] = _1496_ ^ _1495_ /*3499*/;
  assign _1497_ = _1496_ & _1495_ /*3498*/;
  assign _1498_ = inv_14[10] & r_13[12] /*3497*/;
  assign _1499_ = _1497_ | _1498_ /*3496*/;
  assign _1500_ = inv_14[11] ^ r_13[13] /*3494*/;
  assign sum_14[11] = _1500_ ^ _1499_ /*3493*/;
  assign _1501_ = _1500_ & _1499_ /*3492*/;
  assign _1502_ = inv_14[11] & r_13[13] /*3491*/;
  assign _1503_ = _1501_ | _1502_ /*3490*/;
  assign _1504_ = inv_14[12] ^ r_13[14] /*3488*/;
  assign sum_14[12] = _1504_ ^ _1503_ /*3487*/;
  assign _1505_ = _1504_ & _1503_ /*3486*/;
  assign _1506_ = inv_14[12] & r_13[14] /*3485*/;
  assign _1507_ = _1505_ | _1506_ /*3484*/;
  assign _1508_ = inv_14[13] ^ r_13[15] /*3482*/;
  assign sum_14[13] = _1508_ ^ _1507_ /*3481*/;
  assign _1509_ = _1508_ & _1507_ /*3480*/;
  assign _1510_ = inv_14[13] & r_13[15] /*3479*/;
  assign _1511_ = _1509_ | _1510_ /*3478*/;
  assign _1512_ = inv_14[14] ^ r_13[16] /*3476*/;
  assign sum_14[14] = _1512_ ^ _1511_ /*3475*/;
  assign _1513_ = _1512_ & _1511_ /*3474*/;
  assign _1514_ = inv_14[14] & r_13[16] /*3473*/;
  assign _1515_ = _1513_ | _1514_ /*3472*/;
  assign _1516_ = inv_14[15] ^ r_13[17] /*3470*/;
  assign sum_14[15] = _1516_ ^ _1515_ /*3469*/;
  assign _1517_ = _1516_ & _1515_ /*3468*/;
  assign _1518_ = inv_14[15] & r_13[17] /*3467*/;
  assign _1519_ = _1517_ | _1518_ /*3466*/;
  assign q[2] = ~sum_14[15] /*3477*/;
  assign m_14[0] = r_13[2] /*3476*/;
  assign m_14[1] = r_13[3] /*3475*/;
  assign m_14[2] = r_13[4] /*3474*/;
  assign m_14[3] = r_13[5] /*3473*/;
  assign m_14[4] = r_13[6] /*3472*/;
  assign m_14[5] = r_13[7] /*3471*/;
  assign m_14[6] = r_13[8] /*3470*/;
  assign m_14[7] = r_13[9] /*3469*/;
  assign m_14[8] = r_13[10] /*3468*/;
  assign m_14[9] = r_13[11] /*3467*/;
  assign m_14[10] = r_13[12] /*3466*/;
  assign m_14[11] = r_13[13] /*3465*/;
  assign m_14[12] = r_13[14] /*3464*/;
  assign m_14[13] = r_13[15] /*3463*/;
  assign m_14[14] = r_13[16] /*3462*/;
  assign m_14[15] = r_13[17] /*3461*/;
  assign _1520_ = ~q[2] /*3459*/;
  assign _1521_ = sum_14[0] & q[2] /*3458*/;
  assign _1522_ = m_14[0] & _1520_ /*3457*/;
  assign r_14[2] = _1522_ | _1521_ /*3456*/;
  assign _1523_ = ~q[2] /*3455*/;
  assign _1524_ = sum_14[1] & q[2] /*3454*/;
  assign _1525_ = m_14[1] & _1523_ /*3453*/;
  assign r_14[3] = _1525_ | _1524_ /*3452*/;
  assign _1526_ = ~q[2] /*3451*/;
  assign _1527_ = sum_14[2] & q[2] /*3450*/;
  assign _1528_ = m_14[2] & _1526_ /*3449*/;
  assign r_14[4] = _1528_ | _1527_ /*3448*/;
  assign _1529_ = ~q[2] /*3447*/;
  assign _1530_ = sum_14[3] & q[2] /*3446*/;
  assign _1531_ = m_14[3] & _1529_ /*3445*/;
  assign r_14[5] = _1531_ | _1530_ /*3444*/;
  assign _1532_ = ~q[2] /*3443*/;
  assign _1533_ = sum_14[4] & q[2] /*3442*/;
  assign _1534_ = m_14[4] & _1532_ /*3441*/;
  assign r_14[6] = _1534_ | _1533_ /*3440*/;
  assign _1535_ = ~q[2] /*3439*/;
  assign _1536_ = sum_14[5] & q[2] /*3438*/;
  assign _1537_ = m_14[5] & _1535_ /*3437*/;
  assign r_14[7] = _1537_ | _1536_ /*3436*/;
  assign _1538_ = ~q[2] /*3435*/;
  assign _1539_ = sum_14[6] & q[2] /*3434*/;
  assign _1540_ = m_14[6] & _1538_ /*3433*/;
  assign r_14[8] = _1540_ | _1539_ /*3432*/;
  assign _1541_ = ~q[2] /*3431*/;
  assign _1542_ = sum_14[7] & q[2] /*3430*/;
  assign _1543_ = m_14[7] & _1541_ /*3429*/;
  assign r_14[9] = _1543_ | _1542_ /*3428*/;
  assign _1544_ = ~q[2] /*3427*/;
  assign _1545_ = sum_14[8] & q[2] /*3426*/;
  assign _1546_ = m_14[8] & _1544_ /*3425*/;
  assign r_14[10] = _1546_ | _1545_ /*3424*/;
  assign _1547_ = ~q[2] /*3423*/;
  assign _1548_ = sum_14[9] & q[2] /*3422*/;
  assign _1549_ = m_14[9] & _1547_ /*3421*/;
  assign r_14[11] = _1549_ | _1548_ /*3420*/;
  assign _1550_ = ~q[2] /*3419*/;
  assign _1551_ = sum_14[10] & q[2] /*3418*/;
  assign _1552_ = m_14[10] & _1550_ /*3417*/;
  assign r_14[12] = _1552_ | _1551_ /*3416*/;
  assign _1553_ = ~q[2] /*3415*/;
  assign _1554_ = sum_14[11] & q[2] /*3414*/;
  assign _1555_ = m_14[11] & _1553_ /*3413*/;
  assign r_14[13] = _1555_ | _1554_ /*3412*/;
  assign _1556_ = ~q[2] /*3411*/;
  assign _1557_ = sum_14[12] & q[2] /*3410*/;
  assign _1558_ = m_14[12] & _1556_ /*3409*/;
  assign r_14[14] = _1558_ | _1557_ /*3408*/;
  assign _1559_ = ~q[2] /*3407*/;
  assign _1560_ = sum_14[13] & q[2] /*3406*/;
  assign _1561_ = m_14[13] & _1559_ /*3405*/;
  assign r_14[15] = _1561_ | _1560_ /*3404*/;
  assign _1562_ = ~q[2] /*3403*/;
  assign _1563_ = sum_14[14] & q[2] /*3402*/;
  assign _1564_ = m_14[14] & _1562_ /*3401*/;
  assign r_14[16] = _1564_ | _1563_ /*3400*/;
  assign _1565_ = ~q[2] /*3399*/;
  assign _1566_ = sum_14[15] & q[2] /*3398*/;
  assign _1567_ = m_14[15] & _1565_ /*3397*/;
  assign r_14[17] = _1567_ | _1566_ /*3396*/;
assign r_14[0]= r_13[0] /*3395*/;
assign r_14[1]= r_13[1] /*3394*/;
  assign inv_15[0] = ~div[0] /*3352*/;
  assign inv_15[1] = ~div[1] /*3351*/;
  assign inv_15[2] = ~div[2] /*3350*/;
  assign inv_15[3] = ~div[3] /*3349*/;
  assign inv_15[4] = ~div[4] /*3348*/;
  assign inv_15[5] = ~div[5] /*3347*/;
  assign inv_15[6] = ~div[6] /*3346*/;
  assign inv_15[7] = ~div[7] /*3345*/;
  assign inv_15[8] = ~div[8] /*3344*/;
  assign inv_15[9] = ~div[9] /*3343*/;
  assign inv_15[10] = ~div[10] /*3342*/;
  assign inv_15[11] = ~div[11] /*3341*/;
  assign inv_15[12] = ~div[12] /*3340*/;
  assign inv_15[13] = ~div[13] /*3339*/;
  assign inv_15[14] = ~div[14] /*3338*/;
assign inv_15[15] = oneWire /*3337*/;
  assign _1568_ = inv_15[0] ^ r_14[1] /*3335*/;
  assign sum_15[0] = _1568_ ^ oneWire /*3334*/;
  assign _1569_ = _1568_ & oneWire /*3333*/;
  assign _1570_ = inv_15[0] & r_14[1] /*3332*/;
  assign _1571_ = _1569_ | _1570_ /*3331*/;
  assign _1572_ = inv_15[1] ^ r_14[2] /*3330*/;
  assign sum_15[1] = _1572_ ^ _1571_ /*3329*/;
  assign _1573_ = _1572_ & _1571_ /*3328*/;
  assign _1574_ = inv_15[1] & r_14[2] /*3327*/;
  assign _1575_ = _1573_ | _1574_ /*3326*/;
  assign _1576_ = inv_15[2] ^ r_14[3] /*3324*/;
  assign sum_15[2] = _1576_ ^ _1575_ /*3323*/;
  assign _1577_ = _1576_ & _1575_ /*3322*/;
  assign _1578_ = inv_15[2] & r_14[3] /*3321*/;
  assign _1579_ = _1577_ | _1578_ /*3320*/;
  assign _1580_ = inv_15[3] ^ r_14[4] /*3318*/;
  assign sum_15[3] = _1580_ ^ _1579_ /*3317*/;
  assign _1581_ = _1580_ & _1579_ /*3316*/;
  assign _1582_ = inv_15[3] & r_14[4] /*3315*/;
  assign _1583_ = _1581_ | _1582_ /*3314*/;
  assign _1584_ = inv_15[4] ^ r_14[5] /*3312*/;
  assign sum_15[4] = _1584_ ^ _1583_ /*3311*/;
  assign _1585_ = _1584_ & _1583_ /*3310*/;
  assign _1586_ = inv_15[4] & r_14[5] /*3309*/;
  assign _1587_ = _1585_ | _1586_ /*3308*/;
  assign _1588_ = inv_15[5] ^ r_14[6] /*3306*/;
  assign sum_15[5] = _1588_ ^ _1587_ /*3305*/;
  assign _1589_ = _1588_ & _1587_ /*3304*/;
  assign _1590_ = inv_15[5] & r_14[6] /*3303*/;
  assign _1591_ = _1589_ | _1590_ /*3302*/;
  assign _1592_ = inv_15[6] ^ r_14[7] /*3300*/;
  assign sum_15[6] = _1592_ ^ _1591_ /*3299*/;
  assign _1593_ = _1592_ & _1591_ /*3298*/;
  assign _1594_ = inv_15[6] & r_14[7] /*3297*/;
  assign _1595_ = _1593_ | _1594_ /*3296*/;
  assign _1596_ = inv_15[7] ^ r_14[8] /*3294*/;
  assign sum_15[7] = _1596_ ^ _1595_ /*3293*/;
  assign _1597_ = _1596_ & _1595_ /*3292*/;
  assign _1598_ = inv_15[7] & r_14[8] /*3291*/;
  assign _1599_ = _1597_ | _1598_ /*3290*/;
  assign _1600_ = inv_15[8] ^ r_14[9] /*3288*/;
  assign sum_15[8] = _1600_ ^ _1599_ /*3287*/;
  assign _1601_ = _1600_ & _1599_ /*3286*/;
  assign _1602_ = inv_15[8] & r_14[9] /*3285*/;
  assign _1603_ = _1601_ | _1602_ /*3284*/;
  assign _1604_ = inv_15[9] ^ r_14[10] /*3282*/;
  assign sum_15[9] = _1604_ ^ _1603_ /*3281*/;
  assign _1605_ = _1604_ & _1603_ /*3280*/;
  assign _1606_ = inv_15[9] & r_14[10] /*3279*/;
  assign _1607_ = _1605_ | _1606_ /*3278*/;
  assign _1608_ = inv_15[10] ^ r_14[11] /*3276*/;
  assign sum_15[10] = _1608_ ^ _1607_ /*3275*/;
  assign _1609_ = _1608_ & _1607_ /*3274*/;
  assign _1610_ = inv_15[10] & r_14[11] /*3273*/;
  assign _1611_ = _1609_ | _1610_ /*3272*/;
  assign _1612_ = inv_15[11] ^ r_14[12] /*3270*/;
  assign sum_15[11] = _1612_ ^ _1611_ /*3269*/;
  assign _1613_ = _1612_ & _1611_ /*3268*/;
  assign _1614_ = inv_15[11] & r_14[12] /*3267*/;
  assign _1615_ = _1613_ | _1614_ /*3266*/;
  assign _1616_ = inv_15[12] ^ r_14[13] /*3264*/;
  assign sum_15[12] = _1616_ ^ _1615_ /*3263*/;
  assign _1617_ = _1616_ & _1615_ /*3262*/;
  assign _1618_ = inv_15[12] & r_14[13] /*3261*/;
  assign _1619_ = _1617_ | _1618_ /*3260*/;
  assign _1620_ = inv_15[13] ^ r_14[14] /*3258*/;
  assign sum_15[13] = _1620_ ^ _1619_ /*3257*/;
  assign _1621_ = _1620_ & _1619_ /*3256*/;
  assign _1622_ = inv_15[13] & r_14[14] /*3255*/;
  assign _1623_ = _1621_ | _1622_ /*3254*/;
  assign _1624_ = inv_15[14] ^ r_14[15] /*3252*/;
  assign sum_15[14] = _1624_ ^ _1623_ /*3251*/;
  assign _1625_ = _1624_ & _1623_ /*3250*/;
  assign _1626_ = inv_15[14] & r_14[15] /*3249*/;
  assign _1627_ = _1625_ | _1626_ /*3248*/;
  assign _1628_ = inv_15[15] ^ r_14[16] /*3246*/;
  assign sum_15[15] = _1628_ ^ _1627_ /*3245*/;
  assign _1629_ = _1628_ & _1627_ /*3244*/;
  assign _1630_ = inv_15[15] & r_14[16] /*3243*/;
  assign _1631_ = _1629_ | _1630_ /*3242*/;
  assign q[1] = ~sum_15[15] /*3253*/;
  assign m_15[0] = r_14[1] /*3252*/;
  assign m_15[1] = r_14[2] /*3251*/;
  assign m_15[2] = r_14[3] /*3250*/;
  assign m_15[3] = r_14[4] /*3249*/;
  assign m_15[4] = r_14[5] /*3248*/;
  assign m_15[5] = r_14[6] /*3247*/;
  assign m_15[6] = r_14[7] /*3246*/;
  assign m_15[7] = r_14[8] /*3245*/;
  assign m_15[8] = r_14[9] /*3244*/;
  assign m_15[9] = r_14[10] /*3243*/;
  assign m_15[10] = r_14[11] /*3242*/;
  assign m_15[11] = r_14[12] /*3241*/;
  assign m_15[12] = r_14[13] /*3240*/;
  assign m_15[13] = r_14[14] /*3239*/;
  assign m_15[14] = r_14[15] /*3238*/;
  assign m_15[15] = r_14[16] /*3237*/;
  assign _1632_ = ~q[1] /*3235*/;
  assign _1633_ = sum_15[0] & q[1] /*3234*/;
  assign _1634_ = m_15[0] & _1632_ /*3233*/;
  assign r_15[1] = _1634_ | _1633_ /*3232*/;
  assign _1635_ = ~q[1] /*3231*/;
  assign _1636_ = sum_15[1] & q[1] /*3230*/;
  assign _1637_ = m_15[1] & _1635_ /*3229*/;
  assign r_15[2] = _1637_ | _1636_ /*3228*/;
  assign _1638_ = ~q[1] /*3227*/;
  assign _1639_ = sum_15[2] & q[1] /*3226*/;
  assign _1640_ = m_15[2] & _1638_ /*3225*/;
  assign r_15[3] = _1640_ | _1639_ /*3224*/;
  assign _1641_ = ~q[1] /*3223*/;
  assign _1642_ = sum_15[3] & q[1] /*3222*/;
  assign _1643_ = m_15[3] & _1641_ /*3221*/;
  assign r_15[4] = _1643_ | _1642_ /*3220*/;
  assign _1644_ = ~q[1] /*3219*/;
  assign _1645_ = sum_15[4] & q[1] /*3218*/;
  assign _1646_ = m_15[4] & _1644_ /*3217*/;
  assign r_15[5] = _1646_ | _1645_ /*3216*/;
  assign _1647_ = ~q[1] /*3215*/;
  assign _1648_ = sum_15[5] & q[1] /*3214*/;
  assign _1649_ = m_15[5] & _1647_ /*3213*/;
  assign r_15[6] = _1649_ | _1648_ /*3212*/;
  assign _1650_ = ~q[1] /*3211*/;
  assign _1651_ = sum_15[6] & q[1] /*3210*/;
  assign _1652_ = m_15[6] & _1650_ /*3209*/;
  assign r_15[7] = _1652_ | _1651_ /*3208*/;
  assign _1653_ = ~q[1] /*3207*/;
  assign _1654_ = sum_15[7] & q[1] /*3206*/;
  assign _1655_ = m_15[7] & _1653_ /*3205*/;
  assign r_15[8] = _1655_ | _1654_ /*3204*/;
  assign _1656_ = ~q[1] /*3203*/;
  assign _1657_ = sum_15[8] & q[1] /*3202*/;
  assign _1658_ = m_15[8] & _1656_ /*3201*/;
  assign r_15[9] = _1658_ | _1657_ /*3200*/;
  assign _1659_ = ~q[1] /*3199*/;
  assign _1660_ = sum_15[9] & q[1] /*3198*/;
  assign _1661_ = m_15[9] & _1659_ /*3197*/;
  assign r_15[10] = _1661_ | _1660_ /*3196*/;
  assign _1662_ = ~q[1] /*3195*/;
  assign _1663_ = sum_15[10] & q[1] /*3194*/;
  assign _1664_ = m_15[10] & _1662_ /*3193*/;
  assign r_15[11] = _1664_ | _1663_ /*3192*/;
  assign _1665_ = ~q[1] /*3191*/;
  assign _1666_ = sum_15[11] & q[1] /*3190*/;
  assign _1667_ = m_15[11] & _1665_ /*3189*/;
  assign r_15[12] = _1667_ | _1666_ /*3188*/;
  assign _1668_ = ~q[1] /*3187*/;
  assign _1669_ = sum_15[12] & q[1] /*3186*/;
  assign _1670_ = m_15[12] & _1668_ /*3185*/;
  assign r_15[13] = _1670_ | _1669_ /*3184*/;
  assign _1671_ = ~q[1] /*3183*/;
  assign _1672_ = sum_15[13] & q[1] /*3182*/;
  assign _1673_ = m_15[13] & _1671_ /*3181*/;
  assign r_15[14] = _1673_ | _1672_ /*3180*/;
  assign _1674_ = ~q[1] /*3179*/;
  assign _1675_ = sum_15[14] & q[1] /*3178*/;
  assign _1676_ = m_15[14] & _1674_ /*3177*/;
  assign r_15[15] = _1676_ | _1675_ /*3176*/;
  assign _1677_ = ~q[1] /*3175*/;
  assign _1678_ = sum_15[15] & q[1] /*3174*/;
  assign _1679_ = m_15[15] & _1677_ /*3173*/;
  assign r_15[16] = _1679_ | _1678_ /*3172*/;
assign r_15[0]= r_14[0] /*3171*/;
  assign inv_16[0] = ~div[0] /*3128*/;
  assign inv_16[1] = ~div[1] /*3127*/;
  assign inv_16[2] = ~div[2] /*3126*/;
  assign inv_16[3] = ~div[3] /*3125*/;
  assign inv_16[4] = ~div[4] /*3124*/;
  assign inv_16[5] = ~div[5] /*3123*/;
  assign inv_16[6] = ~div[6] /*3122*/;
  assign inv_16[7] = ~div[7] /*3121*/;
  assign inv_16[8] = ~div[8] /*3120*/;
  assign inv_16[9] = ~div[9] /*3119*/;
  assign inv_16[10] = ~div[10] /*3118*/;
  assign inv_16[11] = ~div[11] /*3117*/;
  assign inv_16[12] = ~div[12] /*3116*/;
  assign inv_16[13] = ~div[13] /*3115*/;
  assign inv_16[14] = ~div[14] /*3114*/;
assign inv_16[15] = oneWire /*3113*/;
  assign _1680_ = inv_16[0] ^ r_15[0] /*3111*/;
  assign sum_16[0] = _1680_ ^ oneWire /*3110*/;
  assign _1681_ = _1680_ & oneWire /*3109*/;
  assign _1682_ = inv_16[0] & r_15[0] /*3108*/;
  assign _1683_ = _1681_ | _1682_ /*3107*/;
  assign _1684_ = inv_16[1] ^ r_15[1] /*3106*/;
  assign sum_16[1] = _1684_ ^ _1683_ /*3105*/;
  assign _1685_ = _1684_ & _1683_ /*3104*/;
  assign _1686_ = inv_16[1] & r_15[1] /*3103*/;
  assign _1687_ = _1685_ | _1686_ /*3102*/;
  assign _1688_ = inv_16[2] ^ r_15[2] /*3100*/;
  assign sum_16[2] = _1688_ ^ _1687_ /*3099*/;
  assign _1689_ = _1688_ & _1687_ /*3098*/;
  assign _1690_ = inv_16[2] & r_15[2] /*3097*/;
  assign _1691_ = _1689_ | _1690_ /*3096*/;
  assign _1692_ = inv_16[3] ^ r_15[3] /*3094*/;
  assign sum_16[3] = _1692_ ^ _1691_ /*3093*/;
  assign _1693_ = _1692_ & _1691_ /*3092*/;
  assign _1694_ = inv_16[3] & r_15[3] /*3091*/;
  assign _1695_ = _1693_ | _1694_ /*3090*/;
  assign _1696_ = inv_16[4] ^ r_15[4] /*3088*/;
  assign sum_16[4] = _1696_ ^ _1695_ /*3087*/;
  assign _1697_ = _1696_ & _1695_ /*3086*/;
  assign _1698_ = inv_16[4] & r_15[4] /*3085*/;
  assign _1699_ = _1697_ | _1698_ /*3084*/;
  assign _1700_ = inv_16[5] ^ r_15[5] /*3082*/;
  assign sum_16[5] = _1700_ ^ _1699_ /*3081*/;
  assign _1701_ = _1700_ & _1699_ /*3080*/;
  assign _1702_ = inv_16[5] & r_15[5] /*3079*/;
  assign _1703_ = _1701_ | _1702_ /*3078*/;
  assign _1704_ = inv_16[6] ^ r_15[6] /*3076*/;
  assign sum_16[6] = _1704_ ^ _1703_ /*3075*/;
  assign _1705_ = _1704_ & _1703_ /*3074*/;
  assign _1706_ = inv_16[6] & r_15[6] /*3073*/;
  assign _1707_ = _1705_ | _1706_ /*3072*/;
  assign _1708_ = inv_16[7] ^ r_15[7] /*3070*/;
  assign sum_16[7] = _1708_ ^ _1707_ /*3069*/;
  assign _1709_ = _1708_ & _1707_ /*3068*/;
  assign _1710_ = inv_16[7] & r_15[7] /*3067*/;
  assign _1711_ = _1709_ | _1710_ /*3066*/;
  assign _1712_ = inv_16[8] ^ r_15[8] /*3064*/;
  assign sum_16[8] = _1712_ ^ _1711_ /*3063*/;
  assign _1713_ = _1712_ & _1711_ /*3062*/;
  assign _1714_ = inv_16[8] & r_15[8] /*3061*/;
  assign _1715_ = _1713_ | _1714_ /*3060*/;
  assign _1716_ = inv_16[9] ^ r_15[9] /*3058*/;
  assign sum_16[9] = _1716_ ^ _1715_ /*3057*/;
  assign _1717_ = _1716_ & _1715_ /*3056*/;
  assign _1718_ = inv_16[9] & r_15[9] /*3055*/;
  assign _1719_ = _1717_ | _1718_ /*3054*/;
  assign _1720_ = inv_16[10] ^ r_15[10] /*3052*/;
  assign sum_16[10] = _1720_ ^ _1719_ /*3051*/;
  assign _1721_ = _1720_ & _1719_ /*3050*/;
  assign _1722_ = inv_16[10] & r_15[10] /*3049*/;
  assign _1723_ = _1721_ | _1722_ /*3048*/;
  assign _1724_ = inv_16[11] ^ r_15[11] /*3046*/;
  assign sum_16[11] = _1724_ ^ _1723_ /*3045*/;
  assign _1725_ = _1724_ & _1723_ /*3044*/;
  assign _1726_ = inv_16[11] & r_15[11] /*3043*/;
  assign _1727_ = _1725_ | _1726_ /*3042*/;
  assign _1728_ = inv_16[12] ^ r_15[12] /*3040*/;
  assign sum_16[12] = _1728_ ^ _1727_ /*3039*/;
  assign _1729_ = _1728_ & _1727_ /*3038*/;
  assign _1730_ = inv_16[12] & r_15[12] /*3037*/;
  assign _1731_ = _1729_ | _1730_ /*3036*/;
  assign _1732_ = inv_16[13] ^ r_15[13] /*3034*/;
  assign sum_16[13] = _1732_ ^ _1731_ /*3033*/;
  assign _1733_ = _1732_ & _1731_ /*3032*/;
  assign _1734_ = inv_16[13] & r_15[13] /*3031*/;
  assign _1735_ = _1733_ | _1734_ /*3030*/;
  assign _1736_ = inv_16[14] ^ r_15[14] /*3028*/;
  assign sum_16[14] = _1736_ ^ _1735_ /*3027*/;
  assign _1737_ = _1736_ & _1735_ /*3026*/;
  assign _1738_ = inv_16[14] & r_15[14] /*3025*/;
  assign _1739_ = _1737_ | _1738_ /*3024*/;
  assign _1740_ = inv_16[15] ^ r_15[15] /*3022*/;
  assign sum_16[15] = _1740_ ^ _1739_ /*3021*/;
  assign _1741_ = _1740_ & _1739_ /*3020*/;
  assign _1742_ = inv_16[15] & r_15[15] /*3019*/;
  assign _1743_ = _1741_ | _1742_ /*3018*/;
  assign q[0] = ~sum_16[15] /*3029*/;
  assign m_16[0] = r_15[0] /*3028*/;
  assign m_16[1] = r_15[1] /*3027*/;
  assign m_16[2] = r_15[2] /*3026*/;
  assign m_16[3] = r_15[3] /*3025*/;
  assign m_16[4] = r_15[4] /*3024*/;
  assign m_16[5] = r_15[5] /*3023*/;
  assign m_16[6] = r_15[6] /*3022*/;
  assign m_16[7] = r_15[7] /*3021*/;
  assign m_16[8] = r_15[8] /*3020*/;
  assign m_16[9] = r_15[9] /*3019*/;
  assign m_16[10] = r_15[10] /*3018*/;
  assign m_16[11] = r_15[11] /*3017*/;
  assign m_16[12] = r_15[12] /*3016*/;
  assign m_16[13] = r_15[13] /*3015*/;
  assign m_16[14] = r_15[14] /*3014*/;
  assign m_16[15] = r_15[15] /*3013*/;
  assign _1744_ = ~q[0] /*3011*/;
  assign _1745_ = sum_16[0] & q[0] /*3010*/;
  assign _1746_ = m_16[0] & _1744_ /*3009*/;
  assign r_16[0] = _1746_ | _1745_ /*3008*/;
  assign _1747_ = ~q[0] /*3007*/;
  assign _1748_ = sum_16[1] & q[0] /*3006*/;
  assign _1749_ = m_16[1] & _1747_ /*3005*/;
  assign r_16[1] = _1749_ | _1748_ /*3004*/;
  assign _1750_ = ~q[0] /*3003*/;
  assign _1751_ = sum_16[2] & q[0] /*3002*/;
  assign _1752_ = m_16[2] & _1750_ /*3001*/;
  assign r_16[2] = _1752_ | _1751_ /*3000*/;
  assign _1753_ = ~q[0] /*2999*/;
  assign _1754_ = sum_16[3] & q[0] /*2998*/;
  assign _1755_ = m_16[3] & _1753_ /*2997*/;
  assign r_16[3] = _1755_ | _1754_ /*2996*/;
  assign _1756_ = ~q[0] /*2995*/;
  assign _1757_ = sum_16[4] & q[0] /*2994*/;
  assign _1758_ = m_16[4] & _1756_ /*2993*/;
  assign r_16[4] = _1758_ | _1757_ /*2992*/;
  assign _1759_ = ~q[0] /*2991*/;
  assign _1760_ = sum_16[5] & q[0] /*2990*/;
  assign _1761_ = m_16[5] & _1759_ /*2989*/;
  assign r_16[5] = _1761_ | _1760_ /*2988*/;
  assign _1762_ = ~q[0] /*2987*/;
  assign _1763_ = sum_16[6] & q[0] /*2986*/;
  assign _1764_ = m_16[6] & _1762_ /*2985*/;
  assign r_16[6] = _1764_ | _1763_ /*2984*/;
  assign _1765_ = ~q[0] /*2983*/;
  assign _1766_ = sum_16[7] & q[0] /*2982*/;
  assign _1767_ = m_16[7] & _1765_ /*2981*/;
  assign r_16[7] = _1767_ | _1766_ /*2980*/;
  assign _1768_ = ~q[0] /*2979*/;
  assign _1769_ = sum_16[8] & q[0] /*2978*/;
  assign _1770_ = m_16[8] & _1768_ /*2977*/;
  assign r_16[8] = _1770_ | _1769_ /*2976*/;
  assign _1771_ = ~q[0] /*2975*/;
  assign _1772_ = sum_16[9] & q[0] /*2974*/;
  assign _1773_ = m_16[9] & _1771_ /*2973*/;
  assign r_16[9] = _1773_ | _1772_ /*2972*/;
  assign _1774_ = ~q[0] /*2971*/;
  assign _1775_ = sum_16[10] & q[0] /*2970*/;
  assign _1776_ = m_16[10] & _1774_ /*2969*/;
  assign r_16[10] = _1776_ | _1775_ /*2968*/;
  assign _1777_ = ~q[0] /*2967*/;
  assign _1778_ = sum_16[11] & q[0] /*2966*/;
  assign _1779_ = m_16[11] & _1777_ /*2965*/;
  assign r_16[11] = _1779_ | _1778_ /*2964*/;
  assign _1780_ = ~q[0] /*2963*/;
  assign _1781_ = sum_16[12] & q[0] /*2962*/;
  assign _1782_ = m_16[12] & _1780_ /*2961*/;
  assign r_16[12] = _1782_ | _1781_ /*2960*/;
  assign _1783_ = ~q[0] /*2959*/;
  assign _1784_ = sum_16[13] & q[0] /*2958*/;
  assign _1785_ = m_16[13] & _1783_ /*2957*/;
  assign r_16[13] = _1785_ | _1784_ /*2956*/;
  assign _1786_ = ~q[0] /*2955*/;
  assign _1787_ = sum_16[14] & q[0] /*2954*/;
  assign _1788_ = m_16[14] & _1786_ /*2953*/;
  assign r_16[14] = _1788_ | _1787_ /*2952*/;
  assign _1789_ = ~q[0] /*2951*/;
  assign _1790_ = sum_16[15] & q[0] /*2950*/;
  assign _1791_ = m_16[15] & _1789_ /*2949*/;
  assign r_16[15] = _1791_ | _1790_ /*2948*/;
  assign rout[0] = r_16[0] /*0*/;
  assign rout[1] = r_16[1] /*1*/;
  assign rout[2] = r_16[2] /*2*/;
  assign rout[3] = r_16[3] /*3*/;
  assign rout[4] = r_16[4] /*4*/;
  assign rout[5] = r_16[5] /*5*/;
  assign rout[6] = r_16[6] /*6*/;
  assign rout[7] = r_16[7] /*7*/;
  assign rout[8] = r_16[8] /*8*/;
  assign rout[9] = r_16[9] /*9*/;
  assign rout[10] = r_16[10] /*10*/;
  assign rout[11] = r_16[11] /*11*/;
  assign rout[12] = r_16[12] /*12*/;
  assign rout[13] = r_16[13] /*13*/;
  assign rout[14] = r_16[14] /*14*/;
  assign rout[15] = r_16[15] /*15*/;
endmodule